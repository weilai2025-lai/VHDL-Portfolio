`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/iCW2I5Pc3ynM/T7b7hOaXBqwf+6oVyUjUU6ADI1wBWu8pe8sMnAGoYEXYqUc9i
VkpS/m8gOCBO8JZ93wxflthriBUoKF+N5zWKYzm9b32Ff+oU1eAK6oB2cCPr3lnU
9y9SmJmTKIVdfaHYYu3M387TYYvZf+664P8QZ8guZZfLrMechO+Fnptb6EklT22c
LB7Rieg/Ujhor8w0U5ASQjSMalnb7Z+oAo9rFeCPItTJ5oxennszqPb4PG3N9ZF8
lpDLNihgm3NMG4ugx5GGP+x5186OkupQe5ISoB2VZ9nF61q/y/RdARrPxOFotLmC
GDAe51IUWSBZ77wQGjTpwu71MZrI1QDcwrgkVvNkAHN7uyHLWhL/VI5p4Pg4FZzK
M48tBqN1aYDppj0u5DXBgABSKepMpGioq6NOEdfcMw9vaPSgxB6fS9kuOLUcuLnX
694m8jEINhaCQkzneKeKFQZeUhyiUkdKY21/ajNNPAKbGckIbQtMtKzotQElKLod
u/TI4YTzpwwGtsVtpqSgUXD+nrdtAx2qg6aS8dZemcZPy8l3IyifSnmFWb4QoFsu
MRhGD3855KIgv/StNuSMs+5SNHbMdagPGAlrQtPECaeX40IRIBz2BTj3UCqb+WaV
J37FWFEP8RveVFyc7in8Y3jUuQN6yz8p8Tcty/8wYYQhG2rKykauZCVw7QCnRUcD
NKPY6zJSJLauO9GCb3122HVzozMg+HP13ooPHiMvXvNdCAPUqGp1YRWdTUWSzbUI
Haic7XYRQRJR7eE/IYV4WckQ7SJ++IKVC+0TWV4gWQhaXkF7G9Cci/ArVTeuA+Lt
RXXe0LpCejzxcSqhOkAgA/k00j9z+mj/uSBjyi09we88IshS4pCSH/K37+xF9EEp
FJoyr5wrL9D6UmpaRRO5gJfpBBFn44TO3elOXGBxZV6itTxqOrOQ2QWFAMU5bv6X
+4nSG+ZmuIiDGlkEiVc9YpIDwiejLqKxV+/i/l8dQV+LLTgFFXvBp56Im0I/D25L
g5xezdoRDsLOVs0ouWaeYo3KfR80L/gQ9dIBktZ4gL+x+jslYc438s9J5VGugB21
xKGyf4XaJHvOR1T2cIiFpaca79FPr97bA24C/ivVqJUOv70Z0jS+R3GqUsxjIudC
tPqc9oCteX0eEnZ9olMmJ/vj75s6LSbQXX06dWdCDzw5nGCl/rbxAPXws2owJ07G
JJQIVjo+jd1GwyawqVDsFw6zyifpMLvR++HUXfx4vIb8centMnCa6qUWx2QBkNn8
WWPKbgJslcSud/NDv1WwUWu7vVwSsgwQ5ZsX/fHpRgKZEjLsZdgV13iELsT5mh/W
ONSBa8OSYVav6ta713IaZZ+j/cyrV0iB8dah+xSIg/MmrZIa0OtqDnuyK58sHZA8
AjCYlltquXGfzCg7MnzmxcQp+xB1+LF8SJiKlDrlP0rFOgPTqjh9gVGM4xDRWnVG
mLbj9W4VvsjvBY0QNrGLiZ/l43QJnnaz+MWF5cei7x9ZmqeH8df+0S4cT1hrJ8We
73CFSFDAJRWjB9aoR4Vgi/05rS5t4zeA7PFC/9qEKewuVuNejGJrZWdR5wGok1gg
XkVHdh3ipmGzfOyUoxicYjHDEmmFwZf20RAyWrlAfbjJj7N62cPitn1jHEOlcnw8
GxtAE0e6UPAMwXogRG4qGGeP+uTwo3oXzkmg5+a+IL0dEiFWkSBchsuv4PYHmHcq
0b6cWQpoetxQXIckqhP0AFXbfV1r2OkFbglz9ps6co+C665mhyklotpLXYzQhNGu
33MzW4HPWFHl/vxkojdGfHrIsoQkGDLf9nS5LAGpqBHItX3ScXAiMemK4A9tR12m
tEVuiSUgDF5AMMcihkJqT3adY1Caz4BG/N72tk98MeGWTYPPvNpMwRBu7yPEgtAH
34Cpq8JX0b7Xxk9wx6K3QFTYoCMKdIvRSKl5odIWT2SWRIqr4VyounXn98+O8WhL
Scxa2zZGUttzfwe8egjqHWZtti0wKAKqewSbGPexfR7p0DG91XVBq6Friy5Mx+Kr
H4WxqcWmKzV2EsLY2AXWSUg5tTLQzFCXvK0ktho+DZENaJINK94aW8rlPUNGrLB6
6tA3xzlEmiZ76IYeQ8DWZFzvIfrxwRvfgPbgXmg48i3FnCej1WEVvO2hOIryKkAe
Y3bHQ+6rXWnE/0+4jOhPuQp2L3J+FC21onqQw5usIQnSTuNeq52H5coHRw+wwDjP
TCwSwD1FC3q2m94RtMV1hBOTpFCd5thrxmsPO3ROOsHsi4aBDaLJsX6w0ewhrSqq
2yKAdq5Dv4v6x52qrFHrlfyhhcrf3I+Yx7S9xSDcU/mPlOPmQ2iTEGiuW7IKNYdJ
rVJ0aL+/sQkQytf9COLhfOhufqPQ/ASO272gjJl+PlNH3ViQ0oUlpEKG0aLyJXbb
N7RM6kNENtt+1vVcmBG22/Bbtv8TkruM71YIJ+de/iP99xBpXL1wXQPG36YBa+td
CpLVe3o3dXDO/Xo8qMOPzpA77Re6frqzIi+Qy8a6snX8BTaMeQWSVqcevwExZSLm
DM48xbG0Bx0VJ6hw9FhT9LXDbHCnuBkeAwMWzTVn8Wo9IPx3hf0DuTxdOLkDfhGO
GVLPHCwnSSY+/sMbfSq77KROUiGZbjz14x6MnSh55CgsVWzRsH7CKSt+G33/Rvi8
+ynEnqOHhDIQdn5Vr9l8CdHCprhYnkr+KHXxtrYSqAaUqKs/BLTGpvrnD2BdPK8w
RjUTeYy3j1F8QcaUE1z1bYat0lWsOIHzgfQrScbDooj9myDDrRRVWnlsICALB95v
JJyqX2UlbSKnd+9QAVUD58Hj3wPPfls7bduWWh7gl2JXB8R78mvM3bLj85d0JYSk
lLoDP4MkI+LNDAENo+RHHZ5/G1by7w/i8nYxyWq27nIhob9oPLq5bPG3K0HKgso4
hdnfCmbN8SomVC0IcgX6UOZzQEJmLeuFyrpdJJWX1McZ66K1eUuWu3X4jFiwwV2u
C4d18RM+8+072Y9/xbkvCrsj4VY81NPweIcdoYeh10EA8Vc/UkiK41lVlBwAuQ8i
QqVb2Iq32TXB2HIiGkXetvzCKznUTpaqUe8sXLiDF7Ctyzv91l+DEOstnjdnBaIN
ukDDa3tATu2g5bn8jDflD5+bha1WES7OJW/9Yr07UA7Mrd8NC3T17QKitYrGeqv7
nVa961yagkZ3JUE0xW02jUebvbCNJcJDsg9Nk/K9Dv+ayT3ecvvjhEdkc8Zx3A2w
kuQDVpqMgnfJdRuB/53Yf4uVcH/gDM6Tnhgw6yVuP5YSbV/JZ5MAiyKZczZIqGrX
jdAxShw107UMhN05+aUprMfHJO9UnT58QGYhW5R97MH39+eVEkj4U9HVbnE33psK
c93rUphjMDGeDww5PQhyHPATudXoRiOvEpTzqBBMGO+iVtgi1J5ilY/HJlhYo/yT
s/IIIPSaYH70f4Uhq7MnAKwTpuZcIprOzILftT87WYiKMzgfyyuPgboV4hi2MNDI
0+OFyJGKlXg/zSzcemJtQhozkFAPfAoO2iEH3lbcLwHqhL+KQxpJVEiqWcduRWqH
KBmcsj7ElEtCLhtaWGfikML9z804aRX5tMA10r3FAi6HJki71tMzHWWC+GdLaFVq
joAfwMNMZu41k2jMjICMPPt9uFouDBZjiTw+kcKAtQzUuB7WPf6n7Q2bZSLWU526
8mQbtdLEZZrbY1BgWmosrROdR59hsS/4RlGLMkAoSa/gbBRfvz7eBvAQUodTYr+8
nytSvsixsrk+Jm7eQmbX5kZ0aLG2ylgiVsKIffLqwT2/VBD6aweriHO7sIwUzzEJ
F1NffWEPeMEMDwcA5GgrKQo5pkqApgD2UBK8iSIKlcMv7K4oyqFQVSYW8t3BL6SI
cDMQ6+1LitROdczDpj0lTGDafc39Wdakd7doJqoX7m2KVgubo9hVPMm8NEcxvWYf
CsxeoINGKWbDt+ZNalKxKVQdM2dDEZx2LjLs2ryzGS68NYzqPFxNk/glNoqEbm36
0UwcTG0RECSs/60x/kLoG/XgsJSF7k4x2zWTkoVeM5AJ3iXWzlsapV0OhaHUATEe
qSK9mixYuTdZDy11/nytJv1zH0f+JGES33S7mXuTTIWHSxA7o7Uv+7OU6jfhveNr
U7TE8rCfKN2bSku+/mLq/UuM11lvdNDdF57Euq3+Mo/DQ7QgeIrc+Wy9MW4wneBy
tLhZav5VeNJrCZzG7prQMTPtsQd3uNre0dR37Lj8VrO9rnzZDVnupzUxwOcJyX67
8Sh4rQY3Hfj35os5TUHAxmXSBz4qeSPGEfKzPgREDqKkt7Y4EZd5834aDqJ3B00Z
sneuYa16QPRWZKC1oV1KZUq15nLLb7cJ6woSpLemgNkFwDTiw9a2vnL7oqxzH4sQ
IqgeG4v9RlpHUb/aUpb0JF9hMsu7QZL9nJAXBRmFMp2T+7IRRySR9h/QIUehA6ya
8OnGxCR8vMpNel/5BSwDcs+vPNx4nJF2G5fx1NlkmBop0WwME6ar/wFncvqMPN7Q
uyvH3vktehEKFAIHVm8BOFFJ98O7qXGRekjivXPoptSLr00j3cVOl4RSFzsUCbHp
89H2QBIsYVlwr3g33rbWZUst+l0L7am4Uw7mUfALCRV25WkNIJbfwitWDO6Tn+pO
ETJiXD6Qag+r8mHZ8TTvoL33X27sxMHQZPAak35K2X6FbXj5DGIrmQ+IjhvfIp6e
o8nbf/+BGZFsO8lUCepNqRGOYLr3bL+wmDyn3RGd5CeodmbZTBmAr5i11U9dZUWs
3AolZgnz5yl0VU3k/DkEAZt0QljgAedS2mYDDjv8CCmWwBePNnloMasHwW0VmlCr
2APWlBfX/AikwuQcbUwy3zyWQcn5lSMAgJ5zVXnBEb2/8iKVZAGLegcPHOzqvk3E
+LK54hgHsRxWC+bPYHEPdA//7sMlRiIbdL9aGLipCGC+C41ZuN2fYV/wmcnkBwhH
L7P7sQgghZB+swKEAXRaZZeRQyyXqoUTtFbn54E3uKxmoKyi5Kq3Wg9b2Z5nqjyW
l5MH4qRHihRqbYZGAiu1NHw3xTpNxfxNXtjB5FYAQoiXFkIwv71vwl/+KkpeMvrk
4zRKjg+0VYRYasMCC0Wgnfth6f/iRCtdJu9+uGw3qzqVpbQ2tuQvlGj8HtkOkqiY
JERBeU3lDYHUw8zHiAi9GOS8yEqdnknpZvAcCJhLo37crssIgNlIhjk5EJAbqXIH
Q8cJsg6zs8Q9XvYUEoSzz4Iw4atqvo9G8vTVrGQ8O1Jrmj0YjbfZUBcLWBi1ZZOa
CoU5/jPqJb8dU+Bng6kMqD5PR2sc3gGSWEXZXVxIg5meQe7coW61bQX+qAKEwXCx
7YqvzV3BxiWcfFx7OvQmrMCaA7pzCYdmK2zxV9iMI+T7pF7dd/N0ObZh9k6PSBD0
kItJxuFzWtlY6dTjkELK5JQzk8twC+BWNGZmurRKoF1WrXO6QsPlo53VLZvT7ZnV
yQyjYY0e7V47boU+dKo0DRd3vd64x+WemrI5cUU56gNA7ZS8GMMKp758lLCIwiur
NLxiX1h2RYP5t7JlQR13nMVTr6egAPFEq2mjkkyekXVqFQcxz1XZB8mjC+/1y/40
5pGjewcZNH0u0gYo+SzeLQRXgo3NxJP8bgCHhczY8qPDzRh59f9QY7ZckJQ2XSfv
y8G692LkL1beV0PcaMWzpNgptpcEPbH6KQDzioKOrSTuzvornfbzTfNV2Al5Y65J
AdLDI/Sja9A0nby4zQYMTGIgHKH4NSShg6VKiSZ0vHF68O1C0wOLQ4M4Idj8BIrU
htYFVQR9HAJg6tBk+RksANw2J26KijIUXxG5KJFj//WD4ajuhMFHmDH17BJEQv80
tD6Et8a10pyfYuQNeMLkJSy1P27nHCSS/SDJJPcCyi81Bcc8+MgZBfWXpEglV1MD
jZ3YXa7cuL6WryBRjh7m4h4OdnWAd8DEt0wDWHCY34x4Ss3QuDXdg3zOj/lK17jX
6E5HFklvSaPX9TDRHhIFmaEmLhy7oYWi0a5npybMsfZHU4Kqh5q5on88snGiTIJg
r6vzwEJBUAaBr0IdZRV+qnMlySDyILvnvGoHTAyNjfKXcRb4XOft4VcO3iHLkR9T
DtOZBQEeo74xqrbWMjn9YAGYpeC0//ruhdYYJ6pCHukNIBVxEbIROAuasMiTWdkj
ytw1mqDUaY0GL0R+1Weu3G363WrI1wqrxy6oh9bEUkb2QCr2qOVc6Bb6YuY/v92i
8JFceTKWKLzVj5cBeCsgqKNUvZV4O9kqbF9cWZOzacinh5jCJ9nxzGByVkiqJ9g7
Sq88DIzN5/8t19QpcVEk6iZo+v5u0q8VObaeZrBeZQ6459atbD2lJCO4peYVCgCJ
jhjFV/NzKztE5fJVlFzACbTWs3N3Dd6JBk8fFr0/K0MOLLB9M7jt+hrO5dRWe6fn
Mm0Gl3Qf/60vwqSE7rJTs41zRgmbahGJhhgUnxxcliZDJr2osmnI17owvmKUz4DL
Ds2TYnKtp+3w1+9npdgq62NVtgRphNLpqviEidtcUnr81TKuLeC+yO0Yj7yoxiKA
aj8jCgUQK/3WcDSVDB08STBftrAP9iSht8jn3jPjGrT7kqD1HUBCn+2tSs9gB2DU
xEGrGcLZOCijwmdYUVnaQNZJhXfJ2dBFncxIMtRexlat/At/94I+DYq4SOOqBql2
cyJj34PZDU25yPA+3711GwVfdbMU2cE+vzMwhKW+AhwXTZesWBDg95OYTgu5TMgl
BlCDbNN+yCrAppzLjiF9LXBudFp39ZzlJUomM9gMLfReeshZlOim0A1RTGCzZ3OX
LBPeRfSas4daB3fK3cPMNJT/c87l/SWiPaRH1DzEGcIcA5/MNAV5j+knOZGAu7Sm
xAzS7xrNxkkVowoNlbJT1gY0K2eIFNA2JDgTwBEeOm/uOQ7lNpm4tsiA3eXIfAjH
F5QRCzq14LGTNgAt+4p6vf/diTkbCNQUkAdnjTH6JYEexjZRRAOGhm7pLojY1SCL
IB5y88tzWgo+UCcPpqExtkSrGcQVvMEZzFnGvSD6a32lclkjQ0jZdXdudz6czi6+
yeP1s12549MSJwz3pXJIM1zKX3KcLNOW3P3lQwp/67WcdkbQLI6JlM7ZEimDAVB6
Em7Tv/cgKbdixPmUSX8BiHpDxh58l8Ajjq3Zk8ptaLilZNkD7mTdkA1slLATJiNM
SemMY32Zh+P3MN+FO5YLOBixgbXKEHA3NxUuo53Z5XaIdoie1xeig45TjoENwUhY
EntB5pTFSLLivXE3Euhk7vijW9ZIlwsc855WkByI06/M2f9kbgn6noPQi2XOD4Ee
zjy4hN4c383Rsajmo9sbsXW+G6ptIP1BL3eH//EgGm9PFR0PqXp2IPlVk3c3LfhR
wVRaUdkRe9hUgTSw0RdsXMemOng/Nq8q3xzew2ImqW+J/4Bye7KOlcS4WnymChRu
rEIRIS6aHb9t91GuIwApNpR1lQLYcDtwNOX/DKD5dK/6jl92zHEMmQjdQtHGwrXg
XcRzoCLu9GCZrvzc5FLMEWxWoywffM4S5z2TuuusYywRcicRRrUW0oQ05F+jdYSs
mYz5kSSxJU0X64Q7QzcSnFw4RsaMOC8rfh085sZ822XjwolB6vMmgqwIwOu3dOVN
7hJtVwtavquUswPgpcJNdtsPqSI5m6XrnLVeyTFf1TCss5C9hu63bGy4uOXmyxrq
tmSE9npNYDIOxhzyp2yC0wX67EozXXrF6/ibYoiAgtDXlk6Sp6c/keNZI3rTiLOP
jy1IVY8wdKDEHXMGVFTQF7hlBFsXS00zwk1nlIxQR9/gyfR/23LCr55Rw720Hset
GLzJcZzoSd3xzXJQGYrMv+NrRx9y8kpqi54VgZLGYwzMDmvebq9gfHds4a98suks
GlH9OZGPc1OrXJZzM3qlGk6bMaieNbxdbP2b9xBB0it6HbtiwKk97sx+inFod7jt
KZ6PC9PT3SGXE/Q8iGU7rqVFSxotwafwhyfIRCNZO7DJMEDe+KGJfYYA2Td8PMM/
p8sdQmRJLUj73GJFLDYgnLxBnZR+U4VkI75sbLsB9dn/QJbr9zCG+RsUET+WW4VQ
kRftdF6JRxJvzQ3boSlXb5hgjv9kRCGdvZuzaFFBaFjxwsVK9bj2sBLgOF8YfrGP
6fF6gzAdj5pVP/BXwGTwAuZmgTjUEmSUVBE+CNYVAHw2O48w5zDPsreAYLYbAimv
2iFADD9h2Q1uk2EieoS4+VsvdhqzWNcJW5FaMKHF7j+z2NK7zjRAg/gfuBF3rCou
JYDRz3niidwERnlMwcXTEHwtxjoHBA6vrr5a+Qjb31FdP4SQnZYbv3zhjSFtktpP
D4Maaxp+UsNULnmJ5wZ+a2KcjFstFg51mAJoyFtGZ+4b5IlsMzsncxc+Ca0IJFWM
srtY5rSMmdMmupMk4VVPmKtjiCxMskH1Ck/zLu9iejknE9P7jEz3akPYXmOlNJOW
q9UQhs7XEM22trVc6OoK694KGarYrk3McolivfWpbI+5DE4VF5B6+QRpAk5UZEMN
dwARpumdBJVcsmvFXnxLuHLfpkCKlVbzi0ACaww7meGdp9yQuP6v2TJR1O8d3yrV
NqmcnpZLU43VCfsb4uXIVrRW1P4G5RSMOOJqh8tYx4Dw+72gXSC5qYFpqPdz9pZy
CBwlc/0894NsGfa70S1m3kgRjtmTER0DYvOX+21g2qpP33ucO+TMgwxaCngkyVg5
lv6Syz2ujJrX+8ZnmlATSGZVhdjvAKqRQqZ5FwdYqAOyCbly+Juuckdo9nHcF7uU
sudEIM6OxCZs+1mX6UOv25uForUGlaW7JBEheZ1wbHqDrKX6h0q1Z7LJAVWC9LuU
8dgffbCF9VSy/J9xtRTs82O/Esmk+BzY+Vr1lpBCsHHBlD6RBQZlkVZiJ0K/yWvq
g2zI7PeZMPQdurKXNNg1b05+XKEdBnCvoH0qOv95PyVQM3DfLWXakx7ixY38Tdqz
+12irK5bpVZbg4P/iY5UPXZ/zRJxXECpYw2Y+71ERb6EYhcBRhYSlYhwC6VFxgM8
hXW4yTPF0QeWmxduV8vDXOhrcgA+9l4YrQaRDv/77D8LZ2HV46cdhAcOQAMzq56M
V4o14LxQoWOVRZ34m9auJyOf/V9ZEomUtu9D/Pz+o1v+IkcBh3JDLu02ma8m1tkL
Q5RhI2UwgaQuFCu/FE1zkJI9bSTZbY3gugQO0tBsz6lf5xgBPdUZX9H5p+at0QWL
8PNoGwbjkBBjfOPTCo0JDRMweT6AKOQH+4tmy2/yhWq5YeK6I1uehsoONeNp/DXJ
Z+qRyoM2pSNP0Zm6MxbElDyvhSzQIEqMs34slzWFqeNOGEifpI0T5fJUBqlnTpKs
YyusA7mwPBhS4QycE0VIUF71u4yaAyUuRx6lCzu9YAlJejG24FC0enDSnSqNgWvT
6mSttmz7l8zdlAlpEYeHdQcpfrHLAgodXFUwsolEpkHM3ByBI8+MwzgXlvExTDSc
d4+rrUdtRKhe2yFJ0CHfipgD09vawsaum+mDtlJh+WHc5E7ocePMD+zeQDWED51F
m7eUq/SnSKRiD051p1w15EEA/BgtAUu+y3sjC1fY2aUBrS3pETiAMEfcm3+gtlKN
gWp+sr31Zh4LlMHLk4dQmEksrMFFrS+SiHMpju7ZORvdOvsFSUTz93HSQ+u++zPt
JllWx8nlU9/UAYh9NDh2s8FOiXHzG+/25EvnNVKcaPHSb8lGNQNCRdaCA74LXn4N
9f2j23JkNt2wZ0pFnq2pt8V3jePXgvV3Q5nEKMSMUFe7c2FxBEdK1fowAlaHFv3x
ejANoAuNUffwcXY+7tVB9ZNkWJ+iNfxd53/ux+hyQ/1rM6dfG3xvQZ+18Fh+2U05
76jynl3GlxcC8CrMxJBWeinxN3Djkn49fn0ZyXhfsb9GH0FsPB4QFhllIxhVqYZK
h4p1nhRQnbp6qHhjSANmy1bqVUKrjwiXNDP6l1FDSb+In9bJ8y0eUxl76sLX+YEY
SGJV5rsMF2KMrF8iuHXJFPLSEul4+Wemj76UBYA6DP8EzZ6Ags0/wrK/u0FAyUHK
zOxBQgoZS7ceDMjRwMyrjmNqllBt7JcDL6ADVqdhQYgTKBFptKO+0MNCvcyesLNL
SUnGpI7cIlFLivpEdOZFnj332U6zBR1SetZ2RJ25diDDBzIhOZ26WlokY3C59iKh
m97esYmtMuL4cf8vrZy/xTafGjxVVOB7rtWLbZ7qZESERzyYGDYDy6NYI+E3iqOo
R1Ok9b6Rm5JsWOaZsgRWS2/aa1+ZXhAZ6YDTf30ewbFKm3nNV5KT0OO9dNgD9xUu
mTbOdkHRMWJDvTcV2Yof7zTL9BH84eN6XzM36fk/zf+Wn+NRoua05JbEPUMhbyc6
sDezHcBKzq/OJ5OJZGP/NZ/ReLby0xqFzguIoMriFPAmFV4gInePGsBp0GOtJKXE
aVobg4T9CKudUl5Uud00LQSrUDX4DBkJsTfdd8/Q/9lK2HGgr2Zv0LvUe+2+AxpD
e1AbV//1a/xPPdbVgx7MtEjNmjLQQwU7xWZycnQVii9VwDpK+jf/tf7B2RCxH98b
dJPyfC0fIKdL1DLbAbSbqTRNYoGdLtAhh05xCW3eD4haMWValGeDFEhH8/qvDYbD
ZQU6kMsNF/PRfjJKTTIc4/leifp3qNnv4NWxnh+ZKKF11fwhf6abITqPavmiHZ0X
0E66Ce1y7+XyqJCjoEHATIrREz1a881i500zlLJClf6iSl3nWJJSg3Ege/Okk1vd
8MvuyavPGt4g7GvwYqsB+kMwIbA0XhrEPF+PZK/q33X5bnbcD0FjdVtebbk/St3S
Qt0It/zo49KMVSZt6ckqY/Mw+WR60Ra7Zp6Ldhhlcu6ovR+5DAIuSnafYKT4DccW
6ZMwCjjICBzInjXYNkDwMhjxnNpuEbzhtpXGDiGw6n7Or5YflktmlCutD7SeJt6W
eVpUA8qbJ+WbDDtK8Da0w63SLumSu1FHA4r2xpmjsKVSTJrVRs246c6dBlSEobCs
0ve8Pn118XfFXjhnncvsmggoOgyB2Q+2CuDMD9Q2IlzRYZ6DjBsd+sWN+sH2MCR/
nGkwWg0AwiBiKaIOy8A3vjnQWy86D1DxbQnhqsNbU1CZ4earR8lhxABPv8t9yoHg
G519oMe8Adu6s9xSW4vjFI40n+BHrMmlXOMb93KUHR4tpG7XPl/hMoGyQ52fHVU9
444420U5lb+ryHB2+crHKF2ptga0LzQc4kOZ8qarNFSlaAYw9RNXvdyPxM8Yj2li
EYmkJ1eoMoPlu01uDD9tHAuKsuFBfWJwTi4LcN17EhsGMwIurx+6CzS3ZFlLgBSF
WS2k1hN2pG7l2sTCnDuwawmaorT5ohmmrfKE8crSPuPF2QFWuA2Dt9uP0dbte6Sp
ARVeU95v20Hw/CdEHcea3+DwW7A+igOxLLInc/3ozEdyT4HYNs74j3TAAGHgoqnd
60CiPvaVytgV3WkpUmX0Xe3murSHrZ52cBaUNPKLyfhf2a3QJzNCIgb9j/tVJF5/
lYK61ALzOSAqsQiy8eXuzGMiPHtxdNaHTAeGOgghIGUckv/c4WXitd0xuc8FUZGD
Uvc8qj4oBRYibxSEmLHgUZHNyt/YawPfuUZP3SorhIkSya3qHEoMtG9PQVG5laMw
y8cN9+M7kVwskT76Mcsp6XCi5G9ZLelgQv1RtliM+ubJDKv178H7J6nWvAi0X88w
3Xyzfr2Z/WB6m9oHH/Qma9eHmQD2UAb1Ze47QP6gBd1egSntH0DqM6OqZ3SiNDVi
nl7ziu11FCxr7yT1sqRpGC4VdBq0d+QJO0GuoGJ6jIiqwQdWUquJQl2AvdAE421b
Y4CzJiNf/FzGK+m80mb8l5kLeIJBI81zKht5Tcweezw8/xnXfOKcrSU2euij22PT
kqwr1X66CtD+zdwNMugsOLXwbqO66JkNyfQnVR3iH1Hj6X0gtpzjcYUU0tFTeyUX
sZflhyz5IMNXDjn9qjzrXp10Jz7ik90lGvEf8l1DQltlEXtX/QzBu8WuumNjQ1SE
+GpFbW6yFWewaqbRHJfgx12R89FnfwuAkTKssEi5JfiyL/uf3qYvIvSiNuF1FWVg
IRiIXVc8Mtfogs/jYgd52fz9w9tHCaUk12TASKcykr51T/WMTDvmpUMInWP01aRh
cu5pcX8dwsB5bJVFShQE3edr9gqWrOCAsKUQaqO+fJF/aV9RLOGN14bKtNYX4osw
k68wJGB1I5JCyln1JJz4ZlKUzJIjoQezntc3mtZWPiDktvV4ZvTQURhTx6Oz4KJK
1V4J5tu0jMoW29J9hZDWEJjPY8G8LH+MTrELzb0Xk1q9gayi3yh1B+Qg7jx52dYG
hXwNOqSpI3DssuOSh1Of1+tporad0LMv8hG2nDUxYwitrT1oMYnYEyAlYT/1H31L
IDncLWf8KledpslnT7NZ1ebNZdhouDOJO0WiIz7iGVNm9ELDUeq7fHDeuei1BAjz
pqG107AQthW8pg281NJ/5vpxCLEeixs2/LkT6TgFFpmvKMCWbuPGAN1MUqlm+wMu
ajvM/+NK4eRW4F0Tb4ist7/+ghjadz4DCN9cHFO7En7sriwxOWv5J1+gom57Kit0
YGtE5Lfw/I4rgZS6EaiprG8uknVED8ABtce3V4oCUYHFO9j1HIkCl3LXnbhp/fzw
7QAU8OodNuW0s9Gxbi5MBAoGDDXdFFxYixeiuz7SESHhPLVMIaSNknDReszc28OH
zAbA65U+Z7bq2b8IBMjLK/4xFOUA+WNZPB0DkUJRQXl3ws63oMgll8+Jjg+iHrlR
8078pReeagpnCHAV66/Rb4EgoAXFrZtHHDCpex+1kyBbkAn+/ynzSvsqhjRIYwKv
V8xfWRypK7BgYN2gxmV1cSS/RQXArOjZBUN36qqptwOh5Veu7keltSrYFTLMSkan
YMv4GKONn4Uvy1gfn06+KnqhKBYxeNRnCMv1l5wTHSmv9950rbhSg1x0NvCQKp3o
NDYq4TsRkHryKLPnk9hCIATMa/nG9+ho94qM7g73yqBelziCl1qvkGmkLEfeLtCS
prXnYt1Q9pZGc26yLwWmCT9HdYzflASJ0caRuPTNtzQYhzjKxHKxwaKByUrnendv
G+MdK4eoCokE7bTSBUL9iExRFCT9PIuHLMrMg6ydLKnTxG4Li/CnAoaAvIexUcIt
+7qQbxAZuRRmwWpRUgDN1WnXRSOcs7vViYKLkId7ZLYKHcGeTVFg/kIXgIOrGNB2
XWyUflETRYQX7iXsw38mUnqJsmQFXrrWFpuwADrd/DiRgISs4FKZT17NGdwcnUl7
VRzD/OWlXTYI09rogos+F0BQFx3qFJOA46JlCcY4+JAzSQoVZSfs6jU3pX3TTpB7
LMgF9rWNsxlxS6pYw5DH5fWEWBq4PFCDR9r4jhX+RLZSVq53yokjvUcQBn8I0PHv
IK/GNmmJXcuQsrCo3NIMEwriz9xO7WJfkIf4ZLW6S/7HLgDO2bp0l9qvYGhQhp55
2UigDbg5sk9Fn3aSBeXTf36LRX5w2BtSJnBBnJxSBG+EL2z6O5qmIsh6yx9of5JR
1e+xI4QiPpoMxFCLfStNVWDuMXK5CwkUOa8HCfzokaVbgDElHBh3N4y2GEpcRmV0
shFvmNA0bTOU5tSWwIFbZsGSUJJYF0A8WrRQ588bjfcsIewSph0KjDdrAd9KipEr
48Dz++ovymifBXcRjqIgpQxY9ZSpzonJCEZOtpQjxj4Mei9pLRbQhHpmcB8gJ//+
UfnsFkQiGPh3ulhCsIM+vJ+YIKA0MwlbtPDrzYxOoYXUk2FUdyYkxOLwfzB8L968
IKdNQVvCsljh8Z/2mcIt3chGLu/orI4SglAimeLMV2HF0VdmlmB6ScgYkpVYZL1x
mTARybNUcrc7G50eI0QgNgu6TCso/3mzBj9ktn7dAWKNa6AtBfP3ZnjLORcbtYQp
vtTDNKw/Y6r7TpIsdITzVVUGsAJB62JX8JtNyWnVE+H+cF6YbS+F/w42w65SkZeI
c/jyhGKdsuYa1/R8xuNl3ZiTfdfOX5B5BEBW9ODTKNJTAgVJL0ArEgxBTlDrcOIg
wRryNd4RWpstDqru8M0OxQC8G+usCNcM4g/2enliLElNoMC5Iu5E++MwdgqAKspL
kjFoPuukX9GFJkPBMQr1BG3g9rFPD78wMTTD1cJzIIEFBX7YmKA7U8C9r9rRvsWA
3VaT7oHgZfXSgpRXPda/auX4+YGN4WkDstfNSPJtSXNd0Ft18LaNudj4giotveec
H2yDstgtEVmF7a/jFwdvMQhGYZvZFG7Yjp9a3NujeiFf2cLpB44bBURwJfJKs4pP
3fUU0IX6Bg5eEr8xPnn3AEli/zH1iP5QJmfDvrfmnNR1ny2GG/vMDggdprV1UkTs
ZwP2PlsrlvRqhoiDtSpy588TuquWyGlNDjg4cAZE0WP8+QJDZPcuOn3KBFQT8bK2
aiob8ufD8pQA/R2FUpMe/tQ6rhJhXNddq7ZS6xQEDtK0uRxJ9/lewsSV55X2QDbw
U9TIduydXH0zEMF0OnP15oQ9kurtv6gfyxszTZQnNKhP5GS3S2wiV3FU8rwqKBOv
rwCQgC4rgOk+8pWgArecKvNsc7EthhU+1aY1VbpNsgDbao6JcR1wJw+6jFNBNFLn
HlFZ9r09TCzeaB8IDGv7im/83Y+nKpW+avss1sJS7if9mSNWv/c5BSi42uvXmZlr
mGD2ng9NRfo3qzkSipenzLTtTQlv/W7TmP5Rl3IRiw1yi3j6dT7hRVzPlKM3+cy7
4rSmWcdHnNxxJWiCLKJ7IrNyu21XKxmVHPG6AGkE4STau82dFqiT0CBOJrHFwF86
FXoyhcYiyn9Jw5GBymLsEWFQmEf2aSxVb6fwrKno67zmSUkPsh7Npe4Ur9lb1AT5
1JsMHChjwm/37boz2g/Q+XAma/fF176uPXYC1dxRcXygvDj2mybWIGrcDfNkc59M
tZA4yBCAyPRdclsMnZ1PwVjIQD/8zgDRQ3zwRDFEWmkV7xiVt5ISw0KNGbSTbUTR
YYP68suhHCPK+AlTHXdHvHxqYD3bCxA00X06avFC798FRUUpQ9Bos7uIWUgl/UMZ
H3FhQ1qIApX1sYKfVZW/1W/047msO6mknD2jawlft9l+P4rAC8NQAG6ODN+bjQgF
90zyyp3zxhWqToA6OR4et849vjMU/ByVg+yqQ2Di6kJst9FiA2YCuUfNM3pU/Z5Z
acDsmDAfreXbl19jPzQKgpiEoAUP+W9N5ItKXTiqc59qc5mpdEEij9TesKnztqaZ
tq/66h1rPKvHEQ0n/ozwMUgprIS5uB8uIRDmzY4pbAKLZ3y8Bfp9OXuMwmrkS9IR
cOK9OR6u6XHscc3yaWKxFqDRwC3h9ZSDf3IhcHXOVawCIbjD9TcTKwT2+AEnzL8t
4dYY/40kK+3d8eThuoTVt9XVVg7ny1C3y6RcNcCXSQPl6KzqWDvezYcfRWwobRWx
qSSXiRYPSjT71P31EMxDj9eeXothZQpLFjVEntlmvNNnwx/mAPRLRd4fFrA603em
iWaHnE1phEjMML6MkuFhoTmecCmGuDcgesvFkLbKrC6PEV15APWUikfH4z4dRR1+
iSjXulQ5uD8AeNCrod1NYAUsRGYYpaFXK/q+VpMIS4RUCresKqsEt+338TzsySZc
WI85cZRb/lwaT9lS18pDE86w1ZeoPIahBa8zni84d8FTV7Fb6PXLMrSp/YYWn/SU
ne0XeMUrWvcf5G/OS8GzyRC5xd4Cp/fqrbm2U/SAvC+vD0FsirsCokLh8IkYfaA0
IH/641lSm/BS7FNyhzJw8zOyhlxJdhqgY//FpNXiGSOkwzNPivt02JgCfNJmtTLU
bxGCMzOBz4F42R+pZ1emIqDg6MLw9IgDS6fqIyiPlX6xZxS4H0MRR//gOb0jUcVW
7/jizJhXlfyATtpiVRTfp4Q8buTIvyrcysqv5yleFAyJsEKt/A4DkChRED8mAwpi
Hq6f/ncUGkPQD+fazpUafmYi0nT//5YzewTwxefOkpiTpqH6CFHV7HulwEmwRFts
9cMv+LHkf76UZXuJqSYtk4vv38fvRC4xNRUjP3j4svpJPrrxy1fk+5EgowkzfiPr
OqTxpXGqm2xX2aF+jYSKkd2Ut/q8WC7S/h3O7DrtpEqR+KHd33M+l65Whg/QP+Ur
e83nk2mLcbEZvWwngBC/xZOHM4oBzlkAKw7q8sJy4ss/esswZj/A5XfQ4gQEx31C
aFTp2Np0ylmYjTGzt0voE0lYHEYT5ioLo8xPrbi+08WQiuH03VDOvOPlTdPuw0YN
W42wmIibxSse9GqbxFxARsmvUJH4XbkA7gjDHiud0Y/KuZa8SVfjVXk37lr6JisU
JG0ZwMVsJqqnwJcHJR2DH06KRRfRt+XIfAuokhst2PJpJV0t5TANdL/l8DpA55cW
R7caAAUAktBLc0C1U2bTZBMbQfHa2cliG+iVC0k1Zo4lOdigjrrX3fbJe9kszzV+
C2dlUGXLi4ElrCAmQyMbYUlv9v9sFHiGnXY0Nocnb1ZqnE4XI1FbICKrQsrwBBaY
UhvmIbI2XkfBVtMhhp21QVoD5+l12GE7ZLw5hYAKFU/koq3abfBZ2GYRJBWkbfh6
VIzRoN6hllUJg7iQBklFY6p42JOk24Nb44oCq4m/No0orKhf7NwZBAKM1/ELUrA7
56wK3GkgbM/IdvmyZTgZf0VhrTD+kMKS3qFP+lESzKil+v4TvnsBw3QhK1geavWc
myeI9bAwzwEPHoPajA4J4N1lGIgCgMeHPXr1IbMVr/DhwBXFYiOiyLdN8eEMuRhZ
my8zjr3BhfISfstK6ogzgdV7CwMAQJ0llX5wgh83Vm3dbAuETIEpyKaxqRB6petv
kyfGan4DVeG6zoTVmA71mNQ/GU2s2gKxc3dvwUwZ+UTAi8N2fekzSQaPrfmnRLtM
mSIvx4NsILtUmB2mgje83WP01P1R8iBo7ftMt+Ile/XgxlDLvxnEwWGlwFzIGJ6u
qMf9OmQop6Ffr0NcnyIWSt2lFcrcPOmTZ6sh6AdUwuzDtBdokPfsg5o4Y19eg3R7
H+c6rG3+N1PXjrQN8S68dfczFP4wZa+laei13qEtwjZzScaDumbDeUcuqcRouAh8
2JpuqnyBKFZKyVqL5ugqFrjJYTUn4gp1qR3i6/pWoNENS9xo9ohDGcsshQf/+GBj
1fvcShAX95wwyUQC+93qsaYdhWZyAPLNajP/E+W8EQRA0sE0h7zn19Zb/UBvrGa3
n18h9VqPfLpzQ1e4MKDBnyyvKX2fE2rzwjuS0gCz+jthqM9UJHEg7vyM+DEDBHrv
PgqVjqI1lDOQ9RWWkiPyVW9RVtG0rZAH/Xq7ze+dEftOrS6Jm8vxtP2qMDxp3kPO
r5wERQXj7DW51kq6LkzIfyS+jVaIS4SFJusGv+LtDPsLwCHJ+Pgzjyw6YMVaS/Hr
0KhURYlOgx+uG6l5y946zNsUqEto5zRlE/NRCHcPRI9ZBednrY84eUL7mPfheKm9
EyU4jnPXiTz9YnxtewbKwMpIG7TUEBLmuolm7EtotLTjVWlmMAKlsSAo6AiTuvhd
WoNJA7O7bNI1WpMpzfxT7/AteDFOgrHDZvOpMD32FnYkBoZcaulG1N+GLZi2pfn7
HQU/RGGL5AHp7h4kyC5VJKAPXc5fw9zc+mLkBxoexCfiJ6QW6u8ACTxyEU8bWt/+
qye8Dk0hV+EviinJt9fpwBhGxCgVEPFwnwgC0+VqhgABScMatqSfeRNshYOeGHiX
mroe3gdr8zjOOB5BV8GMShNAJy91aa2BIgq7mK8fbp1iM+PTphzIH1pCfuXvnBSY
jQisBCf5ykoMMu/voBEc+FWL7M+H7i6ssokWkc6n9Z1AZXozCPfgVh87KFWaSPX0
YmakeMQB2q4sIABXKvyL/TnWIvoLoonswPMjDYPrO0/683P/SF/EMJYMzGzJm+KF
qke7Wr0XF0A0+o957ceEHCx77OqB/7cn54aIJDlOPYlZgCFolw+dgtln6IVjldp4
Bjul4A/GWLUda3960ny2Szn4dbxKZf8GEB3k7ZqHgbYbsEtHSSJCpOX0AVhoZ263
JV60qCzO9faMJB10X6Ikko5Bb9nolqvvtKZukui96GMdHHrKO5DKEfWpoGTR0r0S
byRDN/tM0UK4vzy04/HDpEkbuUtFJWPpVtBvfydsvrk9y3Mh8oFd8p1rwuCtf0bX
NzBWKugeH1rxMlrEqVic0i0sxJZoUXm3yu7gK7fQ1sCSBwMHOvDdWwXby6EzO9Nj
s8LnfuVEEr9mG5DIXLvfp9J75MGPooM5BcD/xVHqGzuyr8pLabJBHwKxU2GbM+2+
ZYntUrH+FxsNJp8V4Ti64buyMLlH2DM2GH3jRHZV+LVKvKJJ2gg4TZ5jQfQgqDA1
qLOLj5m1Sz9iQfY0z5VSGxq8lu47Vc0ka/+QSNylqcuoMFyBSQxVksK1g6QKUAQF
8Y6wWU7vrJd9xvRUuHia1KBgIlk7D/zXXhI9AtLdpi9P2b57hv3immhMCY0PfutC
J42MEfPU2h7iyZdcH5cL6ANWlJcSfKsUW73MLhV2IY9hEJ9Soj4BSgElmAA1RQiO
7QWfo6oYHKsHZ4KDzZeG67A7kRDzNalJY0+2445n+YqvdU1hyT9bqLdXN84xm9pQ
PJScOg2MFTjw2VXmbILbq9t82aLULrWkQVa4378oc8WADA7IFr5eMyi3RRN3iJNd
H4VGJvGIjMY0jQABJ6MD/h6UlHGFhO8Ol9hdHPfBNpcUojko8cFcuNFmXcT8Q9BZ
nc/EJTyj/Za9Oy94Sq9NHctY5yeOJn2ATusmdDQxi/nrotqUsdkkeZ268VBFso78
1jPZwrsPQ3dWoofdmapnIUYCYTQFXNO4GVRRm2xoEluVpxBc46UA+ZO+cS+0bWh2
bzd8sTWDjudGwPHW+UboksBAT2FwSeWEWBq/yx2AHtF8F2bFPxWiVbZ433pxU9j1
ilhzj1O5q+j+dT9JEZWoOaAJZu6GJ9zr7EtrVIkuon5JUcRZSRZYIAVsLtfaxUnq
p2bEhOKP+MLHd+Cdxh/PZJpR+91KRFymJsfQ8x/QKkpJUemuljqjWXr2hsOEk2mD
+fWmKXtdqmjiehojbdzrvyRYj6D6XTuBJ3XBtGVNyzjIOpbwW6xNSpdAEL6RBReW
za7aXjmQ67lrSoANYTZ7vCuX5NsbMiQNZuYm7AmS3Ipw/ocr2OAt7FUKb/BQKIO8
vsN1pMT9aCc3sFEbavCBQR/6z622/KO+DI48BkWPSHJ3LTbibtmZtRT16Q8Nz+cE
f4SEpgdEQrk3fJEQpWNZmkmHGb+P6zK9zUfOaIUez5pKa8Z633eLmSpKHTJrel0l
5NM6RDQSGdqIpUB+3ZykJZtUoyrYk7oOKepB8GCLdLkuEboejT0E11d7m+X87GCX
O+AgwIWU0251DzmkUzqNWSDyaUE07Ld+m54Uz0hMKQMDnIoQZxO+4No6vAOlc2ix
3p/vubyNt+mZ37XWx0lawYDvKy3LdqW5oHatzo3voXZI1yl9TH33zn2gC/5gn6GO
DaubXajqv0sXYwckdvjbTaC2VTPxaXs8BFFf7/9qJtpy1Fy/fEdpLw/Zbhj9HJjj
4EfvtRVpu/79Y4b6juNhQUj+1cEZb4z7xVO70R+OHnBZgUrGvH+VX9taqZ/baf6z
a7UHpXG22lTbT491DWv9g3ZlhhhVzW8Ow8WjI9ZwtSnFRqXT8MFXs92PEfRuo+xN
ytWkuVnfux7yVnNXLybqlFwSF5LkDrfjzI74MtloDKyfojrwCl6Jic67zshbnwgh
gv0trhJRkY5K4dEquGrYgP4fx8+7/UIU2WZTkBlXLrNSQ8R0Qcwqz8GcQX1RwCp0
T5sGiDrrvftRicsupiQD1UiFeX3KiW48Dhp4EB6+AtAN+Tm6FUiuBln5KFJ251H+
xVG0yBqU7TnH9MrPq/2nS4QL+a7UpQzjghCMVCl4vA23TYsplvgxmORcZr2cySrY
tDjL+rCAkhmgnPxle2tGSjR4Kfeuo3H3ME/nhIwQKmXBmez13rbpoATafBdE7URF
/f+xd7+0pN2wFGaidV277tmY8nbNKw8eUqZKytLF3ts4XO9a5pnf9p9JJ07paGP9
wXO77XPeazyOMzQEOe8mUMKDKCsgsJCo8p3jcRndpu1QIBsuL1u888Oys5oyw5lg
oGsYQ06DjHFF10YOwGlyQ0KCYVfTZzlgPoSgCJoIBABGWVpc66J4karXWYhuBXjX
nmq8i/sbu0ZYlZU/Y/n9t8s6SZMlMH9ubX5PnRKT5aiU/EG0Ur8f0yUY7/ggzsf7
k6sVa0xLF80xQ3gYMaBDtE/zgN5jVY2zl7IhwOfaDCynNpuwJuBSSSV9WSQg6PPF
hj7qZqdBVWjM7HWh3kociPOzjVwaUvYthW5zFt85crRgyBJws2wOi50snQ0EN1Zo
5h6LRmM9WZqRE7EC9/WsYS0pgAe0xWSULPon0HN9Eccja9T8+p1Ow1u2KvQGbuFF
jISUFoIE+/0NMOQgkYuOteNSjyJWd6oJInmon7zIB28hlWcpN0q6ayC6M/WDfvBP
BZ4qLaNWa4Nn1+spUuqILm4gZDcUAj0hh6uVPJkJuMhh4N63qgm+0CHUJSkfAuzK
a3u7Aw75wAK3Rc6k82rxkY88lIGBci8ZswSErknVwIpX/zko6qkIicQEqFKb3Dwh
MOA3TNzsrH+BJ0CIhVyJg1E6CVkGxj26wTGjP7q8BW+CVWFgvL6xytGL83U5IM/u
ZOT92d8ec4K9SFL37MwQITS7FuvUv7uly1CwSm2Xb63pGKHa/vQNcvU3CsTCB4rV
dxQ2PbShKROkgeq0WJzTEH3pKbg7dXNNF1BrrhHga4Dd2SZrdt3GKAgqtJiEOryl
PUG3dB0oAT+aTAqj3uEPoEobgxdG2EJTWhSudRML+OpaxYEGWOVp4YvarHKqLys+
1k0dfg80qMWpiLPXB5MvYOFwSLSO8FZHuFlrmWI20N7ySw/7PrQ+taSwEc27TDX4
C8NbUbYBpY3EX915esyIGkZ64Yk8IjIlu/mC4BkRqjuj6U/095cC4whzWAE8rZTg
dZ/fJzyfTvbRCo7nlGPJ7SfJjkxVqpJRBUkvjhK85UccMUtibCBX0ZuUYNi1KSZ2
Uqy05GR755vIyv1q/NdL4OfXphzyt0NopvnTwIhk8GiqjP1fpL2KRXW6Mi3MTqhx
Y3SmkcK8n0rBY8RoICUxTBQKXumCwdhMWRrbf8Mf4jPK/sPjH+RXj9k+x98V5lgJ
xvO8jdT4h+szqKZNarQZJccI2TwHtEWjTtaLtpdJXUobTMtrN+pRDxF0u6BL0OBj
GyETEAJBDVZMmwO2Pdn6JYdlaJWVnCp+dQlby+G5RnNGuCqaAOKcVlys4W/xqYaP
7CV1pLye+p2kIMQDHNCWl3obxaJPVCu5QG5o32emQ9B68EwEYxyH+zVnr6XWkSk2
WDklWBdtTs40X4Mfs4mBYN4+INMKCL5IKjZZeyr6cDrnF6aL3JQ/l+B+seKFxDQB
v0GzsCXYfN1vVKyiPjW2nJvTOCMF2GlsLvzgycPGCkNFpK4Hwhw4xhTqxqqgez+W
h2vZdnsvj+9oiCDDETR6KnwYhVI+GY3wwkR8rkK2CppbcDMDMbkDENr8G7IkNCQW
I2e9us8DnO17QJrzdMCj5ceL9zTbe6844EJ8uATMIE+0e7ReFVpvUgo9+G83g4h8
ZD3K67D6haOYUt5jFXYyqDfdnVmpRXJoUYHv7GDw2+4Bn+tnHIDUiTSMkCD+WWH3
XcNpNoZuGrOAKndOM5IW5Bxxz8YB9m5G4Plgv2uiuF9A58pNJ+GwbUMYBeAnUh85
MdlB7qMUZOmsFvSjSUOrIiY1r0hb43c/E3kQX0TuqPZ2o89dLAcZyl8L1MFQn+tY
KUM0CT1yx9KWvaUws7PuqKMpXgS4rH1LvSVLYXRGa0XN1REunkn1TxmFTKL+yYFF
PFvv73Ja2C9f6wvQBe0XsimjPdlg3DfhLwFCsuKQHdkMw/oI8rsqBzca3p+5dLUQ
1s3x18B6OHzUudaFjIuWIROj5R9rv23bi5gdOvnfxuo9Vie1ezzpMKyMXoggylWO
2z4UfIXOM+JYhZASI58wmy+se5Bg70NvT5z+kTCSR/30IagsCrEXbiWPjPRwvLNe
Kp06ibiaHKmoO3xU/tY6vXATYNDRWhU3hq0bQCYDG5WPmGl2D1BFbuFjgbPtiCMt
QGJqlLQNlPt9JnmoOGsHII2iAAhCDCwF692WCvrs0PRAA+z9SlUnlIAkbkguzrBd
QnA2+kMod+4+1NG/BfBUC/o8g6RcZYFwfBaxDyzpIlqG+TyqhoYXf8XBs/5lenwf
+m5CqRy917P9ZekUXOMobcbZOmZgQlNBC0Mi92qWq+TC6jVR/nXqcC9arwqllgRL
U842JnREFjMLM3J+oKNVFvtpqBF+S3x2zcDpCOjCwMFhwEdrfaTnmVFvstIFchc4
BmrPFsL17eLsyXOriUeGCd+jxHVwbKmboIjWHivrbFg53joAxDVlk3IFuhs2wLqs
bgfgvGdQBjxnvxEs0tJkvBsFUUn8LUO8sO2B4M8nzY5xhUiuO7yOtf0zWdXnrRgU
HFl7YCpDqMe9dwZqR3irDpeQfpoBvlJDy4GefObEh5KM9+SKc9kjvU8u/1kLQstB
IzWjEMxEJkmSGjhfLMh+/8NZYBrjx/Gk1z5r+noloilpsllaKnI66uIOb0a3+qeR
/RXtn5ritTQSIOt3BXmb9E/z6uYn0IE/DhSglzGB9DRfI9gmBXV1jel0ato2Ne2y
KZCGOPzo+XWIBvV3RBfYKHar+/MOfzcxR84gYSnhZ0sCkZttyD+pbxo9qsGbfgMX
ZvYKUoQWLyTH7UsX9o7y4UX8R29/N4W54lIS737DEre2eB0VbPZYPac1cBOPzee5
Xp1DPwQ01cQoUPWV9F7P2a99iY3lhk0yICEqsdz8zIjXH1/eO2e1SgdBLH3ZES8k
PkDmx5OK07l5+/V+DRMQdGjZQcubP3+UZhC5wzE3v91B2iOhknE/Bfvmclh2k+zP
BDe6o9TdCFFvNqTukZItHncOoOQrDw3PVRvGgMK4leCFXSmtbCmVb2cqx7x39k8b
WBiPhpXKXF8v5vRdvnbm6HvkXLIkmaI4211WZMBSY4Ljo7G5K9ScwqfXzm9CbN4G
OyI0c1dU3Y+LGSHa6pDJ7cMG+9mmx/yG/5a0cSK9HFidohQxNLxXZOPcGlACHwTJ
S/jueGMTG7ffw+rQkeTOOcy6PxJLKbYGghKJSkomRh7SZZSUuI9q1n3ETOQzHg43
njMVVrVBqQCqj+yD2ixhsvp9raoGebcUEDXgSwTOmQ7jigsMKlCcfx3jCyu56QU0
Ka9LFEAqZww2WqglLgIK7VD/mKabMsait19BUNwty4bvglZ66776FRowFCEA0TeE
ji5HlGI9aItHHA2xaxpZ9gxZDsbE3ZshWbbmcBotEdQxgmZOL+5HUWBGGUCnTIXs
9/0YMfQKqDA/L6cS0MCHfJ+2A3b/t2NDneJ01ZWJxl7HxgmU476UeIzOv0Kszj/h
3BR02CroodFk71G7aHu0MnUiqDt0hgHQvhA653VxD2bRxDvxeHcK5WBxi+Mdav/e
lWfokVsQ2n1wq5ZfD/cpsO9VeNsDJB+7RlXEqTgk2MdC4sjdRCdGXs+gh9YoC5ue
ALBzcftvFkh4bm2ACxePXXk2wswZgY60fzomefV8DTYGTMUfkNGOPR1pw51Xw61c
KDohVTr8juvhvxSWo4vbxJVXA/cBKa3qLnrKDEVqnu5D2At5rq4gAFDdGYfBz27K
bh/nLehwd3T6hDksNTtZWFK4jsMbXazfvson42E49/kwDQHCVm5mxBpmbfAAVuTD
o0kNmbXFIM31+MteIn0x1aEkePCEassCxaBlFbpog1/NRgCkkRQVHBX8XkP/enUC
qIrDh77Hz5hFZAlnnMFZRByGkPCyEFIegYjxuHDL2y1tyHenD3Oduke9vFoPRCGm
fQY8FaKRgFrWBM9k5lyXukSms3Lll7UooeAjtd4P4CsdYr8FhwEc8wZaAf99UDnR
IWkMY5grnfTqCGv2GNncKk2va0ccOznxHi3FDQ8m1769M5hlgTa4cw1hR3g3sF+x
zu8UitpYG6P9DAw3Npdz9WyjuW5DIsG37YJ49WA1l0i65+sZuIqKM1izO8GO0QtI
hCcvFlonxZY9ZCDII1N3PPnasCmmq6eGUzMMnnocayZbLozFvH269UqIypKnwMWV
dO6+bKjpE05OpKRSQxZmetiPqY0+CQJqbSr7MZWp6lAXYF1O59DwDubN/Dx62MlR
hRQGsxEahqW/guvyMi8wfQxMjz/bKg7IfdqOIM4ZJlp1xC3rXwXwN9IU+PUThz8W
HJcumK7FHKvaYZDKoNKDkKWSKfegoJgOBRFPqZUh/AkmvhhqHsXn4mMOD7A6K3ot
ixfhnZK/mti7lFjf1T/IVt1YGw2iNNKomHdRbxfrU7y8pytVqlZnidvmTncIZ73p
WAjSB9pzIQKN+BOH3+sPNZp77FWEpGBEVADLJ6o2+bK8x3AwtKxf5n6H516yA1Ad
ogHQ5ukygnTATEF4swk7xY/HEnkRJigixzJCIIMC8a8NZWx6e/qDit6bXaQZa6GV
isvddcagzhOhYmlRCgWj8JUmtHToNxDTt1YmF4TijY0QTQdOb2+n0hLH8J/ue98z
LufKfVTmDqyO0jvzZKVH5BdMYPyuKI8g35D3IPVLcTwZQRbKkqQxDvVejI++SHcX
T3UdnHxmGpn8rNCNH3NfPpgJAr8NhZHyD1yHdDohmLkIkNtVy+nUnXMK0yKHKlkb
9KNQHbfJS0hHPs8e2bkXsxKLNJSL8bL/vHwhc1r54oxkF18fQWQAhYhJXdzdSa9W
5vskYm+nS4y9lfmlns+HCxC+v7CbuqhsEG/4O0vZHYShldEhgdfiePnjhSBa3yNO
jmlhE5bW8t5S9C/H9khuxJ4KVkNyyHYmrLvoRn3ioAT8BhgBEMI86PUdK6YyTSyX
J4FtcmomaJ8fzsODMDjdiwk4UtyjvbPLgouMMlUoV3rlarwRIlSH+ilclSevx7oR
4vzYLJN2X0HKHl8vC53QhfqfjZryqEuarBCDbveiEeKDIfluxv56kuLTQJ7Zgwkc
m+2z1Ag7ch4/aziy+VQbD3ycmAR+WbkhnITuuTpeolaaBksd7/OmcND07QeCjxBf
EtFrAeIDfajRby4dix9oKocmgQyBztKdFf289rYVp+00sk8qQ9aY6kZvwfvgPCym
Jzd8zhc4BuoFQFvP5eKfgvXmfJGdJjCZO6IpZEggxK0wyXOtdHA2aHGms06UD/EY
almOsB7mnxuMKMaXblEGDNWf0ZypnNQggOsN668IldYTGnJl/lX+op9+Uy3CnfEL
HpLXR00AEljrK1V1khDQO5wzE9obhhpSTONZ4VrDzawvBqgwhnfoNOH46t6rPPZZ
JoX1ey3xi+8zZ8x3/1A/Hj30JYRpZSwGxY3IqiwAsG5cWJi3Onm6CF7NrPXv5DSl
WCMz/N97HUKrIBAkTiZCZ1qPpbJfXAOx4awsNRGgQgdRPzvRJNFpbal9f5R2ZX6M
O5c6VRasZnVq1KEqHJ3y31ezxiDHuZXLlqlWVnJ/EVRu3gwQbXkPwq00NZhkLpmS
SKTFAtGEladScGoib6uxsvDTIdzZbPQ/we2ULpyVn3N+TFycYC/SoH9glocNBdzR
9V3MC9ngkIXDSyD9bPHlmVnhs9O3K9VaVlNOdpY8Ea/FgTnYF0twrGbykkiQmiRS
SvfQILtZypJfDXzxR87Wvp804bTXdwtOEnHYXXwvMjLCxiVuhbcPQwMR7OUVXYr2
JI67OdgVGhx3famfIWWQoUWWODumYdLwo4Td/0siQk+cqEKNra2NCqWTWGM0RAmJ
xIefxDhuFbWlbS1rwZKCn7L69685vFcIX35f4HzCxSRwSkHZ7xejBFpkRMcFJtqE
4IxXG4szP/5Lh1nzdFl1UzKoxHs9rHnKD6MQMaEnErHreBmr4I2WZ5Fmy3DMr7AH
R8kJ+3aIyBHi8yFeHr1ciGIM7G+bwDKGfpDWv2LnsTnAvz8Ie2iG3bvdNVBvcuEO
NGJY1MAjIFIfWApkyBSeFlm7ZOWuY6YUAkCmlnFQiqz6xVwR9weF5GPn/DkBKnM5
qpBlE8K4NFxrWew16Tkg2MckOwdBYX0gSxoEpadZlbntdeiQ6Wvcr3uPOPQN0x+q
44orcwDaPmbey90UXdbRygYZ6zuREAlS75LCcsKitPm+OuoU2fH1fE0y7N5BtEl1
i8YdJqI5cLWc+C5icdFeWXEI4LVRN7lh6JqxE84Wq+JsUo0slcJaFVWBUfefmT7/
sSrn9dHrxKfq9qO8JUoh/apxECeqliGJ95qu70ypgtLZL/cfkgV2n6ApquLO1doC
MXQgjIyyfsV2wp00k0Ubed9uuWlRfpKZRLOJoeT1egS+mhDUHNmOl99alvOWVrLw
DIKHlUyNAeSgdIl/loH1JDW5isxYxlDzHTS0hQTEyOuq4O+SdYJq5PV6+HMce/fh
KfPE2j2XTQTPN67goGjWnFX1Qz9tquxJKSOzUpiP8sPbp0TR2V/tmqNn3jVWSqY5
/SAo5AvJBvFmp2Q3H8r2e8i+z1oL+ZhXMpmZWRIPAzs3myjIwEgygX9E3MUu0mS0
2Bbwpu1Ck5sJCo9K54XB37CL/5wU2Vh6QIeEX7ibrKBHKIVUfWYujfPKKqjIkBk3
9uSkV3g/BJ0oHkpbWmWkRXElZ/xzS3mFgmIMDpzDK92DUIxBJbGBOlKkaTj7tf7h
oQ2AKuAMK1AtJj1UUqHtBjWE2ytbV20I28W0rF4OW97cG9YEEIGjVUUawevzHFrC
J0090gBh9yHubdfDV/E7QmL0ugXFdJtA1OWKTek0nfoGqzWPokLxdVsxstEFvxG/
HDCVTxOXqR7jLu4DYzJq4c2alrFD3wyfwK4U9aDiWQw1LJNiwgJGvInSydYl6CDX
Ln2whC2FtDDvGrSrjezlg9fAc2CsaXzN8XBxJjaGtDOxODVA6OKfbBMCXNeyOOLE
a680/ExRU5ykyB02KprsiQvfYiaQHS9sJJXVR92CxtPGWqR7aeeS9DnfrCcGNH+p
qTRPHvek71JOKNwYT/3nhEeV0JZ9kDXkbtqqDaI2MR+VUAc13tJLPJJsfD2s/gRW
vMCUOQ6YLNaK0joBUewHSdnUek6Mf25x+MPY5jsLRFMrpU+H7SV3MUAcd+0XNRmM
ZPcUfnCUO2y/omdLuFWER6UuaEbRDH9YB1hQPooYwIrtYtnZMIjBgR7kp5Q8F7/K
BZMpnul2tGPpuQ6ceOaFUo569atjGYoH395Ns00I3D1qHIQyxynVOQP/deEdIzXw
cxhG/7lyHX5P0HImWpttQksguVS6Wpc4ebeQW7E8w3TN3rg6kwWWCTnvP9X4duxJ
SYiam3g42hDRTcWIXUM8zs0rvG/IANozF9VeTDmlkyQ65/8fi++TpdKRcZIPx4NB
Ng1V2799QsaLNvasOk/qHeLsWRb3KcUbdTTVaPD35DeJdCPB75o1cjGkanWkkZ7A
i/OxrTumhp9vZgWxlVamj2NEhR9yBCZosu4glTVlJhXpw/ZeKz4G/ToFcQNHoT4g
8KmTvzQ+4O0ql5N11AuXlMrEeJETOyUxc5EH0HgbN6oOd/HjBJHJGvk9Ya3yZm7m
4DZfKg0Ybe2pNRvp6cFUvMGHtW80ddAQzci0YenH/TuG4hU8f8Wf6iQcb80xoBJQ
iYiOmUiUeOkrYXW98A/vtF/p1g3d4b6YyfpNbJ9f46YAmmckrz5BGApiXv/DG0F0
EifVeVViHHiV3LndkUB2ZFVV2d6cTLjHj52OUp/Ln1PXRWmIC4gLsfSxJiSUQFKV
FcmqL/yR1NChD/DfdcbL83SoNPYYRYZ4mXSTcuK7Bhuk+Id7gO0noEzlHkf5sNzV
+2TV47Xr1ZO2qhBj5LsoWtRXYXVX+G5xRVxqxLlwc69wYjjbTgptR2PI5r39BF0s
JdJMkBOFpgqtA0Mt/EahtoAUPESQjZQIbZMtQu7NACl6++EetR2T9Cae1FuBSGur
UpIeEVcIb01yQ6zHmQS7wDz1iJ/EG4oXiRGWMl538KR1z4A+wPfbMByYnWXx4/Gc
sht339XkEQfIVA5NsMKcMqAWxFImEILJbVSjbhE9pjgqPdnjvxM4kkpCIYhV1iIn
/Pfr9XNaDc73MG1nQJFs7n8orkbV36tjK2pb41jPVvacZqBkBwe5TmtHAP6dsPus
gRges7U8b/LUBw5UQdka/6oBiRkul8UIdBjgwWQVNl2INaBZNbY43a5VOdtZoAoP
AMdKS8S6IwFDX49l1VI3S4xzjjuZbljEOfMa+titbBbeVEbKVh01UIkO1DZLtNMQ
mPWHZtdy+X+pQy2ZgKmg6yZMMp052Mr1gf+GcEtGmIdKRkHxsNNaOeUZe9qAOLi5
zw3Wh7BHc3hw8w1c8AuFmVHYkwyrEN4vM7Yxi5A0SSPbSwz+EC5W2l/qKP/H7Xxs
vP2QQYlsi5oj+lAZCPiFkhScE+CLaymeJaJb2351k8sPFwhvFipZA2w1njBTciwM
Df5x+jhbww3Qnbtcd6O+64IIMYI6CS3Bu7dW8Buq+I1pVZD9BR4Rwen/vJfSGP2r
yFXeMkchpIsYUNQ7Ubgg2wryrd/Bw/oIBeCMXK114g6wTHc8rj1T1wdLujMAPjWI
wBKGYG6dye+dsWabAP9xE2KMHyVsQ/xrumCF9G8D6qYerJQcXklMbqJ/I6DJ+SJ0
iSIw31IKxvT7gx92ZrEby48m7/mkvlpS9lW90Zd4/Lxe3UbQHb+g+Ok1JEEtXOBE
kB3ALjeDHVlY4v9mr/1o6yMc6ZLPz35vjc1L70KOmg5w6X+0OkivTTs21ZaeTbkG
RDH3wS4cH8+Wg0GdFiV6vdAsBUZ5SzBBe8knNWybr6ARHumghbtvKWinG04WZ5SW
ADMkaOfQQrfoZw1VI+/m7WkZ8PhID4MZgkakYnW0gVZ8+vayjUlbt4A9z2XXczlX
fCDQodZc5VWrE0s8AZfSTIqvfv9WPuiHe/vrxw5VisS2wrjcQilmRWWlyWN6PElj
7qCwQHnpNb6LHOQhEpOn0tM1vr8QZySxj/dYE+mgxrz3ym1SJ5G2df6GOmpGk4Sk
VRVigr7cpiwIg2gE0yLa37ggJwS5AKjH4UU0r375G0iAxyJvFHQDYBesEZ/697oX
AKAyBcmusGojGAUFZ9e5VVZaosd/KoZlamhMYHDBe4+pvbEDTTDK8yLbpsU6BjLn
8B2qexxgpAmvSba1E9rA2Dv5IsVXa3SVVnrSYgUnDqQFfYMh/D/nyj1IRxjMRnUa
q7/QCZz104XkZb4UXRNDdOQKFMLWEuetc79l9xSRv0qWgLqzxGds8WImqubZnyaQ
/2WRe29PbiS/d6WP96dVaJeVAafMNsvjwtc/336ucc6Nh4hXrD0X7ao5iYgMaWNG
6B+Sz/UVA3rbgKhG4ErXNljJtBRCQ2SW8KHAspVETDOBadQcgD+jpFZkA15yjpew
jbWZ8YJCEzMnR5tbQZLECkUxtn4bYQpQttTi7SfEBcBSp047JDKrwvOzoWVVytmC
1fpaKEd5i9aaVoyjdq4XJP20wPO3NnwutM9YDV1eK6h/3BNTrBkP7dd72sghqgSh
aPJrWZvCOFdsscFKCHgs///tXUkujoPWpE7ERk6wd/Hpll4R4td/6rcmD4CDm0BE
wyZHLPH0EPimkhHowX9B0Hnk2vyKkCTBWyOH0IYEg2nEYOPu6vWNpIYxp++HuC24
DhZ02dm3nXQYvsKhSxojajJwVoYTSRY8Gq3nD+X8EqzOvm2h3yPoeFskYiWM+WHP
oXAgOSxa8QEvS5JvXVQyMGKus/dWKF8hZuAOcpG6Zsa6oEVTx/QDraJfZlPvEzbu
d0WBlBuP2/4YLe/o4K3kjVOSyGKRzGWTgj7wn3/Tsv300QUu6MxvPDDwtnWOS3ve
IyGhB+3AHVR90Qe5Xr/siIQyXz9MdS9L2yfluy/TIHIuBlJduF6YDQFb3NaHJZik
dNETmttqnEQd1kx/gd3ki75vteckfl25pmhNiOSLWOBqQwrSfYSaU25YJlJvC/j/
zZEZJLjKNikyOHKFeagDEBsEs87zlBZthraTsmeNfmYD17vZ/sNh12G+/SqP8o69
+NPDnciO4aWAI1HIXt4rwgxpb8u64v8e+ip1kG4QReS657kSMWjZExpvn7Ur225p
2zsXvjbhD03S1U8OOXR6jtZzT7dt+9OCTkGyoBtbu50zcMiwPOqsptsuib2bYkRw
CdHXmENGYt61uM3k/usnxsKGCNhggX0UEtAfSP/2MQq4I5A/ebK1imsbNqxmJPV6
2Ab+RNIafHKKtWAWMicd/FYdiYCiSIscGZ5cR3iMErOafbbSNv4myIHNIixrXfPj
TV0aOhLLLO1AnpD1PrEEDKSs9k7YPWZ+Vcenq7CBoUFMRy931RGUXyxRqCLjdlfU
Pn0Qo4yIaku4MoSC5SeVswa7w7lc4E7pEzIS0tfViKKNuAvtibu1bFlZR2BD0s8m
4Tn9HSrI2j0EzGzOD68SL0JkYQgTxLPbVkogvhC4S9pRMKzf+TcK6ixdLEuWxTPg
8unUNtI2Ezqj+S4Ae3LS3gr/OpifX0RVgDjVQUDfPBt+Y7vP1y3Ume8PipAPLJcU
wjTwaZpLg4no8d5++ZpuqccQH4tDwebvYM6lXR5ikK23/+v6V/0vzUoLbE7QkYdJ
LLYLwsasq00pqIDaXxNeGa9otgi67+2lnD/Tc7g2IEE/x31oUpu2EkDHQG6RoUYA
up8hYJkyydKhd8Ehrey/3RafM2YP7GQt6LrJ6NsCFOuHCffL9NnAieeoIXZeYErK
+qFgb8ZtzLK0o4ART0hJSF497vuH/kJekA6v82KIC4EqIATKyjOyriiGjcdhF4YB
JXKQc6A7HqA2c8psXJD5UQOT+GWgQ+htkaRMi1mYzivvaoH402qgjfspEiPpDKxe
+aruLPPricJKN58jkH26Ga4GnJyE2A1p44By42RjXpsF0lBbJ8di5V+eGhKSSCXh
cNOD0OmMnJbk8PTOUlnGyJmLgFlDtq+GG7yPD9aDmPx3xAvsh39u7h8is447yyjf
HQoCpTi2XdzLVcDqcV4JqyLlZ4UjC0w2YL05Ea50FUM/CrG9CRM8341SOfrK3N3i
tP2VwgE5amC2fOO+KoqDbVPHGAI5hteiz6OPZnBbimlgt1fZk8tbtz+X8HrMapct
+LDrmqCW3HIxVTDx6mgOxa/cwWKJ40+qMqbFSFPyfM74uPF9fn6VA/TnzDosZ7JG
X2vnAHz7GzldZ3YOYCh89FM1MW1zHEL87u3JkCewBmnZSUSeMVgEm6MbOXC8mtcR
txY+QsQgppzKAr2JDNC+kDZ+JGV86eUMJh8MxPK0i+j95OkHJZE4+7VcQxNIf9Ps
GKEooybjPXuul7SkD6mWJqeauwGbYw1zbCrQSuXNLV+4turL4QFRxi0494Z8Q9WD
JCSHVJcO/iY8mUT0V7gA9HUN6W1JCRV5OcnTsOX792OBWszm3Iwd/R/4sYybGC3K
NHHl5p+MRlBXu2nqwlZnQZUH9xvMSX17VnDdBZ+wLW2e5TcSbvrWkR44vyKgbu5d
e8rp/YSca/XD3Ff2lf2TTY5ABZYwnOP43KH93JzJ9MDxi7aeORgo2+WmTE2uma5I
AabHzUnYqHaqS4F4y8UtQ/fQA6zqqluGXqawTYn06oa/mKZmbMEeIofnPGXb26EE
O7b24hY4VZNJMUXwVCG+zBM/nUsTPXIRAXo5ZcjNzsOURPA1q5pEHsTu+bZza6vF
aeuDdgDqnDGqCU6n5P0u9n3UpKjBy1Lv+VPvYwSdfRgw2JwtmVsB92H5DkG/SDUi
cEKCUyBS8DBCzbh5ZaLkWKKtNX2XIsk9RLCH31dQoDZATEhNv6wBKo7nvwiu7y2+
KDylgCZDRhFvnU+2SH2SsMSQ5mfn2o/M1+ZJix4sXuaojvzUCNG9w5GABum6Rnz8
mGuNYTZ7SoQDAEvitxkTQNuyU/RGSj5K4amz0UQbWCWmpSpjpQLDHgSH9h9RvR/1
TpIY+is/S/3r542YYxblCRJEloOfV9jXMn27nq+stHDv+dXYshk1jxhyuWBnIkkO
2JWzATSsW1TAItZKcpyXrN2tdsmLoSscTc6M12SZ1P9rwLZ+5K/Qedm2lpO00xfa
HSPrF1LSLVv1z8whWnrMBFtTmKVDNlgFLbUnoua250u9zeZ/iW+cT+43mypTQddc
7keHhwwzcw9cSFQ8vSBy6CSv/JojEe3x6qt6eNtRKpk7QRR3dSu3kVLALGO63z8y
ZNRGgFow9SipqzHCsobwmXpmNosZnhxZCgFzZ1R/STEZTuMh901OKONZAUsG3GOW
GRB9ctO0XcCnSWiyLKK3e8XFDYysqNL8zZCO98z2MxCOo2h9qhRHsMO15SYjhuq+
xzRAdbGKN9jBs4N5p7pIhm4q5kf2D99FCfpGx/rr0ukFEpnfloiZdybPuZDDnjYX
zmr3DyTJZ7YRWcQnM1xX2E60qdIMbK9UWpspXJQu23SlKUsB62rA6RJHyq/FcqzT
79WWiHlOWpDnzdqgT/b6WbEIv9GlNsp8jnYQ71Ih04D6ygEKlJjhTU3uRvcBVd+t
5x5WQ2peDqVwyMc7lPaNm0Vbbw4RNyNLPQurVkH7lcdSxHGEc9k2rW69woBvD21Q
mGg3S8I3E/wcmG5bnKe3kiaFbmKFzhjYOw9WytHIfk64K+ZyyCNHCYE9VP0UWrk1
G/LY0zjUUIRFMBO0KRZ2nMWjSnPtSUmwQetqyuHQiQ2rqipJtxFp7KgbZ9d+pXIi
vQFcVxqEQyzKZrnwdeFCMzVXxlV7PRSUZzCS/8hoaI7ocpNac8VpFk0qvAw5c/fC
Qwdfaz30fz3591+IkBEuaTWgtgk0aRdulPk5ng5Tv/xOQ4evVLRgrXMDLWDyBdie
TPIYxGjC/lDqF+ZoAPlzedd+A2H0KbaKGbVHRzLANFR1CQblwaKiXuQd7V2m3S9h
aWlWF2z0m8TpSPg/oLfuq9QZ74uYhQFV3jSpyQ4TpJ1lYD3VXfCwyKXrt/VKpyut
1vWCYTt7bLvyDqyr+tR6/Msnq7YIaePKePnQMcveFFdE6TFVGqsK8+IsNwJWUngd
x0dxmdH5b6k0lBBPr7MBCB4J1V8nc1kiyCGWyp0i6rLmJr+fQcEAJgjK1Nd5Pbn9
JsCF5cU4wm3Cbjb0SyorE3kRnklfhEsKWKp4tXyyZKCBMH3bed5OxHdc+u4qiL26
crwPUwnnGSgyzb4oJY+GnS4gDNEhK2l54Y+xZqei6gQ3TCuzkSCiCXSEY0KVcWtu
4gIcf5cTbh0lJ/rkIllrtQcZr1InU/zufgAK3O+JVvkAnqFZI7h+DqeL5GdFseFc
UP8auhHrSFymL/SBewQk8ZHvKJVGy+Vmn3YXNiehwhH1VChTdrRIrYJQGAugn3Bs
FIJM6kuH66OdvHWKvgE9JVvXhJ7mZHZnQfmDMrnz1/Lkj+3kr9KrQsFlAsOk/36F
10l13v2CNbm3F5Jtr2VsOxUkuYZuZuM+UBTseODtaU9sHkHrM8sVa/xueNi5W7yw
P1rjPTikQ+iT86ViU3ufsMC4zSC//4be43iLsxSDkdEE0cOGEvAUDw2nGLp08EKE
qYmDtDr29L8hBWLRWGRAEE32fke5q5e3Ic1hGvoTrliBMQcm7pz0Zie7rCEqxsme
kTj71Dx0B9IMJh4H+EcktIFAEtdSakWV5ewMSccZMEuc1Qx8yFMnNXpCTIJgyB2i
TNwvi58ly4zsKeWWukTfsbuBAFVW0XqrBuWqIc77nVLIBFgD2+Z4pLGlZU5zLJJ0
jsjV+zOzNLA/Vyp5MTyuRgcfuMDf6EXDy63ZWIngTKG2pNnzYP3ZxYhQRgGOrGzd
Ao1LTW80tyn30fyxPXgjGh4Kz8AIqgxcZ6XO8pIAY+KxswZjOgXG3DcQD1RNKkwL
DRtw+vfuPHONdLTC1KP6Ur0vJhrebYH2fR7p4oc8+ZHBQbK7SaaXHRVPhs2GG6tP
1CcreWLbsqjgyNsg288iUZg0ktcLknGgK5q0MC8YkLPHSRg5vBIi1m/BcXvbLsV7
Ht80ike7EB5Y4l9tyFKxdZ13h7NRk9SiJn6RfsUWljs+t+D9QpeFl2kErz1Hzl2S
pJxWdtpoxb32Sh7PxUhFj2Jgo1zQeh9VOPhNmKGo9ygOuiHWnyMAXtT3QKvcqwSR
OOIoLZB9soRLEvsFekEKRbWRwA53fewm//bH4d/TyhwKqL8/JfUeapJGsiha88v8
ginORPNRoO252XXHw4lgGkfq+PiMMkk2kftv/K8pu7vUdkTNw/w58EuY1HWf8LHq
4OqQKdMIVmBKF3G1vEtCUk6ov9ssPj/1sYAuXeKfcGXYgV22uSj+RyS9orjszxMB
qIHmbP1Fbt86cUoARkCjHVARRZzExopd/80VPS9iNXcmqzIu+Rhpfox3Ko6vrxLy
DoRNM4YSU153eBgru7mHezet2e+pKrHdkkbuhS3PcPn+YP8efWEROcOOBpeSY8n/
6PjSWJ3/fmbSMZn3njfyJGs+Bvt4Y9le2l4jbYP6Dt+tMtZt0b4J4JqnWLdZ0RPp
w3tRidERbbZ14hlksZ9xI5xSDIWIuOLps8VgPyWL0RPIof1ITQ+A2NKAnbtAxfF/
9QJ2BjIOy54iKCKMbbZOUhJ7m6gZBah0B66PVUcM/uME6zBeBGkXq//p87J8pQPm
BgCAuMs+Mttg1vIX2eAX87w0BYeEUWAS3PJWLFUECvgxFNmpDxznjaUfAJoXPjgj
n+bgWXX0sYKJ8TZ+RKogfw5U8ZSSD06nKAWENmt/K2e0ZgJvadcfYPmVxt76NWGQ
msPYb56Es+inadfQqYJLGktBEg7C/aNIbWvgQmbnOAF9QfOjmmpElY2lwYCeGASg
iycFeWvDIsCCjSGryaIKCruR1AFcuNEEHh1pRV0cSqW0grGYNYc98l/1egYswvrD
AW6wNSr83MW6QQrf9Qkx2hWGRA6WeQ+IDpFQiypI7rD0/xR5Xm0NT7ppamcHgO0h
Gf/qSSePtiuL3nb5NtnSyfTDCGtkH71y0FjUb/l2RWxjjZBm0OiVGNCsgefCexWM
oUj6GApnAcu/IW6mWhdcNDh4hGvBHT7YZBGcDQTEuW+TP8CL58rKE6+suhDI13ds
KjwLFCL4GFi/lpaxLD7wUW8wY8U5JDZCKg8mLgxcJRYH2dSkaTWm10VEvaBl6TjF
xW1gm60LRg4js5V8mDbnVm9cxIAwgM60BX/LNci4JAcNkH4w0bFVmrHvm6Dk8nCv
5fWgWI/q2Yf9LzoF/AuSgBYZXMLRp/oSr9FqOg6GF3vspOz6czuhmfXCiu4+VyuB
U255NHmATt9G6QF+WLzOHphenOFSeXuGLDRyqkwoG6DWNSg425mfrbtobIIq02Pp
tsti2SH2uVpr/Qjer5uGjbERQM9pt6Qj7dAamDTg+NEKeSVBsTncjo8tDPUeYL8v
N0+CeAbsqjDfYFPhAKU+n5Sx714kGrYdc5Btc1iMLjBle/qvjAzyP2Zmqx31UE7I
WNyc3d0CTU5w43s/kWGMPajMDtinwf0GnQb2/orSJh8TMSKnGLk8LJXbRPEV6X33
v1/x7Wf8Qkqh2R/wfG+pLkBSNNomPIpSpgnJwyvMOxWnNusU75Ul0bAw/XBBQREI
b/0cgd7/zcPUphKNE6+QdoAy2mG3mdnQjysipIG294FQtQziRTNKXc6+qJ+AV8KL
VZv7dNnQWwETxWh9jjtzN6QbKp1GBgBLsv7QPCOXzz/cbne8+JHxNjlroJBhm2dP
BAqtZbRXPvG0+YG0tC3M+bQbCALF5S79PjFuHWm0rAosIy61xbVMyTulrtYgYGFs
k5LEYZDuNiDNqUsr8GI+0grEdinAJTSP+XG/T+voAfuvcO3bF2jrb5eYQ9jhn+Ii
4A1Qsjs9K/Rruiv0LMuT3CoaXXFIAfCWyn/QOBfhMEaWhvkTP4fLQMjtJjOJJgBO
xO5p87qGDll61I7LOCwqrhfbdd4lMsn5Uhg2+3srB2QF7TJc9OhAiNkIjC458pts
NkWS5rc2O2s6PPxdMmkIgmmBgUGLit2MApilgKO+eMUUvIGOw2c+340WJ1uOjqRK
LbDhhZxS/OXzON/NpZtv4p+g9gsgFKpx/y4yz0pRUhIxXO/lgUf5WhyDjFxnNd1b
lr9KmayuYBv8uyC6La9JrHzeFo02KrbEKoklFz/X9o05j3OxoL9RDG9oBwEhG35V
f2uysjYcIVX+sWc9x9lOFFDjFAHmtZmg8KfX31o+B+DLlODdoQ8yR0jbVfjdLR7g
E/ZOfH2ZLZyqaQ2d6ynaWeb6YmdQhUzPO9AO6xFX4omvpASxph+JXHRRvuHeNg7F
cbiGod9pCqZ84AAALxIL7FMblLNAndo5fcwSmNr0EpjyNpSzprHfc8P9VdH4FGY3
cxAcpBHNwYFU/mzX+xwy1ARrijKwT8qjTmkhnOigv8hpRoZnMcEw5SWb0gfRb0vP
NwMJNvFdksM/HWpF1nn4Ln1dfv9LLs/8rbn/maKl/qPzRcLqfI4lw9dtAYZjgtXP
ZlA8VPFdJJAJE+dw4mfL74YVLDdlWy4BCuuOMe/V5QyqRQj+elsKBMggDpd3OXR3
RI/+NbluWf34HT/bki9jLOqp0ZnAhum0Nm5obPgp0dqVj8z0DhetPYxfyeeXLF/b
0wq0qwDh6EikopWWGDJM07kTA7EydVXzFFt9m8QBhLAmJvzoad/oiCgAs6DVo1F5
7vp4GUrpqbV41Y/mId6G8MYRajSDJCpLTdzJIEoHBzlCgASm8wb81kBZB/FVPugI
urceinjoWvOtDAvLELyjCNZTTnSlRbaQ1fSFGF0cCQDbRq34lNdBml3F2uHB4HvB
e4NaCbvEM8DPLZHyqqGwFu+XY4yX4D4AbDZSyO6NAQ+dBwXE+YqkoGUPPW3gZg6D
fOBAFxyyLtH+2xz+QvY8gG7uFKHdY0fnS9Kzhs9YpXwOfKymyZNEyXlklQL9Gisg
hkj9tCHm/pzz9tBUFsev5DUQVx0Dt1DHp7KFAj+VGYce3YHR2PEkgSJrImvWIFAq
vMdl4Ciqw2m4BoCzcPFF4ev+zOUQutU7NXLbLBeJGGd2aMHXPxsNO+MnLuv3ph7n
QdRTlfniBPxtet7XvAgqxke0S84Ui/D+Svw0o2k/Cq3LwmoMj+4Qo6Mhi9P1m5by
hVhrR468wZVnIhjbmeO7sLeMTwAhlB7Ny9yyH0tJEmpJqFP3ondYPT+N75xGn0E6
zm8ODD05JKy2tLIZqoZc60PqHQEnixm32Yu8r4T7Mm+3kkP+BQH9K1MsfL14Q6jt
O/L8sGharaUWt16Wyu/awFG5f1y7ystm94ykkx/QAgeC/xLOXyoOvoSBxG17LCzi
BfDiPun7Ul27UG9ATRLp/+TF5CwPAAQCa9bEyMYNwIh3vL7Qd9iI752rrUqv2O6S
4/PLOEgnhPzYQ7QZ0OexuMfzbsUp8TCdwEAOQIWcbL2VDBnpIltZE8hWtP9i2vs9
5utBosvrWB99xreBk/k5FvjPOjSb4IxQ7pkC5pHQTk1Q8E8/nP0ou0H9lzdHPwiw
KnAEDkYkLdbAIRBZinWm7wWiMJR+sfPfWRmEs5jNgGNutPaIN/G+lDzzQvfPGcmC
3Zm96fGV00z4aFTW+PoF5Q8DQ4g4xk7dFGzBQxqGkZW7+WHJlU0c8d3QfGN+o0+0
J7mgdZ7u7WgYA625/vNKlYQRK9AspD71WcSNcokVJZrkdRaBOoBKnxIRCJFu1RNO
LaruYPuXVkTTzyVy5tCk0YvLXqCXPMLG2mHhRhqBz/DVbXaJDgXMMQoC2L0tkRca
WGXoVe/F77cGZpvzWLPM/D4Y0uMdpE0BA3mhfypBxnf8Y5KSGtzi4XWKlXIP5iGr
qO3uQj8O8wfjeDZSV5H5s9MdlL4LtPKC1p+mTw7iIuQTAb6DFnU07k/dlIlkij1O
nqls85oaI9y/sEbKwWoEiQauFO1gl7Y6UOS5in43wzRr8LCbEW8KVqKeKk1/1YLV
DzjReShmeCFC2GWBoAW5UbmEzAX0bE930IyMVav2mwDZr94j2LI/CixZY8w/wIUz
FTp2cCbNxkH5b5MxtWjDAu39XanHb4LD2TBFfPbHsx8y/DP640MB5vLBcoLZrj+W
H7O15EdnFmxYqNgfV4+y/nU/Ap/Kp3IMLViqGdKcvFHsGB6hv09R4VQbpPby6NSc
7T8vay0YFW73AMUqDOqQ/8j6+8HJNJhnNlY9/fkTQeLHG4cM5/n4Ima+6CjIutkv
SA912lmlo79c2Wxn96lqtEhC0i/h/T3JIo6r019upXwSbO77vxlVEufZEXHjmZgL
rivUs5chRfKySwEbujj9X377huIGb3dYSB8CBxDOu2yu7Bn/JKB1jdGJJ0V/v3sE
2FTfUUTbY+mKbMWDW+nPCInYRKZTolEw9WQwkrJdjQ7XXJkBffWtQxNTiutytdx5
YbCFLyFR6UpGYqHL1BNLxhkCF2goMPbSsfQuMUZI9T5eLASdSTvW1CCAbrWTtl19
TfC0r4lckJiUA7sIEO6USFFf3X+pQORRGk2D4THmQmZWxmUQktcIZckRwGPRqi06
7IrX/QU1Ky5dSCmQJRNV0pJMhp/JaKi1yQ5EFNw1frkyLWoFxVNe00S3nlBLXwkI
++k1PYGWQHbS3SVQQLdaiEJ0524dhkt2D2m32NDINLHlCeVywaFgBenIN9t1tR47
GyCnwzzaMDYkMvrFQ4U+B8ZywSMJVUo8jSIhXglmNX2NO3/3DJH+W9UD/aXwne2t
CM65q9K/EkSZBp8W9NDIV42Jwb5BHZZFAX7xER6oMIMmNazICmHtZrFeBImxfeC9
g3H3jDaGq81qqHUsjsZsn8edS5MkRaV8N0xyxcGGeJNcVNuB9lvVDFn4LgMJIszV
xmS2PwQZJkPRXmIMjJ5cyVdvEuu4Q6/tDXTlmg8dh5v1vfEqijjW4URUtEyFTo1h
EvYU3vgPL8CedFoUqng5gT3O4rALuzxdaWKeO7inLnGzfm91aGD8c88ne0ubsH0i
NenA7eVYHiisTMtqR2MW9coVj1yGWQgSuUbVI8fbT5iH/2Or8nTR/GlC5aiH7uaW
Rv1TfAM+nhxPbrZj+AIYLarGjIffpkmTeX3+YRWodxHyPYQh8h+FBhKe/QgD0ti/
gs8E4XbVUg/5bFEVQTiD1WR0YGBQFax7hGumLvszRuufYKxnOq8KGlXfA3y1UyY2
lxiOQnir05nKUf0waGVmFAFDUoCpqsfjAObA1sZ8mSda9bZwzO18JuH7PeJHAybQ
nGo3uuZi6O3YaKkr3P4pxefdAVm3R4rcJ4YNHegIxYpoGHZ3DrzyLqBtVBVX6bvi
9Z0sllXsgWTI90mNcyy4/iItxvf8UwOoYXeD7FdTUCZZTWtu/iJHitMrqkfu82yV
U3a30KUewVMQSsTDUpOhyXNqItOSuMDKM4kE/mnwiLsOwJPHo1VMCBuk0sCyILVP
9CkIVbM85/srWu3xqXL3xDUhzjfhdWPai6sotRkpHTXg6H01QVVvfnrjOTJW8wQw
s+sa1UiKVym7mWA+Q3urTF5S0oKVEil87iotg4DunNoBf9G91tUgympn/cYK1jaI
I1/q/YQLFssz/BspnUhtXMUgwU42Ou8spBREz8zPkHnSbyffSir8pS10pSGKyQLl
KF1fekiJGMyHEzdOVCmmmAh4zjyOvJGu6mrxtUwTWTc5GhdbmBGIpXIVZvmc8R6K
aAgBRtXF6OJZxYmpY8uJsCLjhT8nAssGrkzIuc7NUnq0+VSdMTkuhHzsblJJpfQH
XQVlKu7E/2e7qCswszXvX5Z1SgfqbIBgbFmEjAMP3WY1v3Fuf6aRNRkVt8yz6xk7
hfWf1U7MaMplL9I2HpAEDzalvj2Oa/SHYPCU+7NiBlLLh0SZpPQdvMJRco6TCn3t
2KjG70EplV11wwiWmTrMPk7ZVBnlw7Mh32yWp4YZVV4kuI73JWlT28A/rPap8UwR
HLYp2j3BjBY1Pphdz8+57lAWrVs21cFGjAuI30wdTftrtMOxVgWGu6octYKmLxY5
E7Ujfb+KbGpra7Iy2YEJnKsx1fqLStMiiZg1976WgCvW1Fk5Q/9eEu7OsyFISB0y
01z1y4QcvYNNV2hviCKIWwnALMM1oCZs/B5WprNSDehN+FBy2lml4HfxpelQxLaZ
x5Xk3o/1R9P9wesBYVKuqiHowuYlc7eL+mOADVxA37L32jMy4txiC6GXq+Z0jaxG
zN4QfpZVCOemkxnlUUwkgZKeL+St72+/PqMRXuh78tl4urgzCiDC96MPAPxXKFmb
faucSWYHNknwDoijh1GpcEFRkjXmpRMPfhpfa/xN2KcMvfEmiIR333S6xCM0DUdF
gapvDW4WOirQA/1FDNKZ8Si0Zzh9QUK9EPD5fVgA92TcKH8/e5kZY8mkgClkjF1a
jBMq4kB2fu1Mn3o6iEpPW9KsC2/Pmz9oXv6BVXve4XzqFNawPPxjf/B/h7jaLczD
YfEbi/ak4PTSEGiJPQxaa8vj9HbH6+lL4X5iAwySI5r0WS32zYrn4CnRfv9eOrEi
lbl5LSRoE/jGq4L9n5ZZ5ygrKYdH5FlVUAWXvphTnZkEb/0dk+YTb/Nt//iYDW9U
6Kl6a2c4oOb2ABp4/16f2saUDej0KHs0auk0ObeTaJioQiA5zr1OV8lnGKePcQ/x
GVnOdm88dE3Z7GLGX0AG3C43FRsY0b5Rg8ftLUj590hJ3ALapa8DJ0aPsBcW3MpZ
EfpmuS/C1Eh+OtfcHMPpdQEKbLZDPlGrRcvX3JoERSvRsFj7ao7MqwhkQ3+KfnZk
N7IWLOeiJp6NQ4MnGRgMcalqXy67WMTE3fGVFN2LZhKgaCZzq/78hOP/iUS4i27x
LggqrQX83gPoRw6Vt6M0uchq2FDMJvci5UcOXJlTGs2PRg1tQhwwjK7WXLIf7V++
Vp10rKORXMOJsE8Pt/j5M1MJE7Pmm/q6/pegIuaSJKnbXcW1Zp9IDzlISI4UTvmx
VZylvWEXp3Fzhfpf8TObAjdTR9s8IiSPqSDlDJYDMAkjsCu3eKwDmwBtI91mOIyY
GEO8VyewhKoeH/h8QD60vCGJtjxfwmRUVskfSywM9BcwggJ93eJLKOe5HRalalkW
YE7BBPTbQTGjjXfj4BzgAsmLfupPkd6hP+3gJNvflBjatR4ivxkeSximXkevidtR
6kUOXTr53jQhxS8L4kEqHnnfmheVXWhI5RFsG/FiW1JSQ+0ounzKpuzLj/06ViTo
+9MFWtFxsmJK5NKjgCO6mYUQcUbfwGQzqcksrwwRIjitLZGwbz40dIppbyXILck7
zBYwcYNPMprd8wCyYEUlZZNdacv+pno+41XwNOvSUXIj1D8D04qNzXRX0dfbs024
rYoZaeoVT5zxw4HyBcToCm2Jo+GJCLPTWOeHs4BiIIP+BQCGS2fVoh6ga3eCh/b1
OWmRIZ2YoUAHBMnPD/vljxJh7w3iEMKRDEcN5t+DNFpamaBQJYTAhsn6WdYOEZig
c8JvCEvhbWYYkKGIoSeT5HtxYEx77WIkScqv+T9C9htVqlvtp/8QLh5Hcwvs3HUH
9sdSoQh0p07Oy2E7aMe6EnbxIjVTkjOQFi4CLJ3oULGM8A5X3pi0B/hXstw8tU0o
zenFSBKI/qhj3bIvm344Awetf6zvK/2g1Sy8Ek+3laHv9aV8xzDbKy9bpmGuO001
lx2wF0quR28TRRf6tIo4K0kFi+n4UPGHwC8sIGQDFaBbt9AVJ4wHULmGGVgeCWz4
YQsehFIgU2bOMBb3t4EaKXBm7fsNP1pfI5ntv/+1/GuaKIeeGqpLKNQ5Yqz214IR
pyyCqOCx+iOS3NlgCrEA07r9Oqhkt342nYSQ4nwz+6Wkf7g2Xh5HnMTTSjJ7Fvpc
NnDH/+Bl+0up6s6KFIfD86GSSulRqo0fhktc2WgtitSmk9BdY7bvxj1xtHs+7EOm
exY7ikFrMLYU8cAv+EmIqnTCGLDUyjzD4+TC6wd/EkME9B40Hsn5Gp12XHEhrhx1
e5+bNQ+qVDqqmSumwjE7thSKiAiEnSuh19WFhIlVNGeWYiMdjipFY93fyLpRIQNE
zvgYR9D3Ju8pkaS1nDiR2hc1JaR6jIL3Ryiuu+F39pP9FwWLvs0R8bcXiHZzGkkM
16UmFD2srTKDBFIH+V3DUe2Er4ulR+rMhRbfHn9Z8niwVMVv1yiMqdU2FUie1b6Y
9Jmg6x0IQBzSJuBb1/UCSmoueSmzGPWY8koTj8hZ5i2dQiUV+uuPJvrHLdYs4CYD
VM8xXKQ4IjqmCwCOjZzRGKg6axoVZeBJ3Ngmk3do42TJn5+2sChqT5Tg3f6uZ0i6
/46AvV3/eK76RWmOElhpg5IjyrTtbTc+FMfAjLXv7dd4xFrnIvDo2L+VFISUi5dv
CB7i/BEDsHZTqHvm4KYzFFDmyzYd5SiMKtvdCr85HNuJMCu87BcSSkUgWstcDyyb
GVdwrLju9pnSlSLybp/VqqhZNKaFb4zLd6Mpst0fXjzqrROSNFIpD9Zh6wDxY6eJ
QBwu/Gt1xlr6htkJRAkjiCYd6iBpDMkd7h/IUm+t3VMh3lUN+wd0Bu8hcyBoj3nz
lGXLpah3Lz/RaEWX62y95eqIPXdkCGt1TXlgUXW9UXoqg5Vtd7H/YFtIEsibPJaO
mOEJxLkTrqL2i3ZaC2yv5NJo9EpcA9cr2BZMjS5I4vFd0v0Vbm2hGuQxXBU8Bgoi
wLMzscR9TvoG31lFnKhRS2F06/X3I+4kMoREcHvczkOTRAWzwSDCrQU46GBztTE/
EtdFFnb9cMZ2lj1VSFGdCFafNybQr/Y1Mw9OX5nyLUXXbjMuCZxf0phRF277HlhB
tf4a8OW0XQpybAfFRqgtgcvv/rVPrs652sNvIGug32jdTIWjLRnp3QSzq3x4kYAo
FMZU2xbLLP7t+fiVwJjRewVXxZiZAvkUG1uLW/i/AXlOSayaU8EG94zRJ72qtt0p
gfATJpyVmOaBc6n2elRdHC/pAv1Y9U+mvy83QuNxdR1dZRDtzCtQQI/cYiqLoDxW
asmPSYX8m81ecuuXLc7ZRtvO/8z1HBy6B5oCXLDDaq95qLEGb4Z3Z56wZPRpC25q
Gg0d7i2SrU1snRn0/CRx3/03QoAvAyxDW0bMghcFeiiRUZVw992SanbOhXhgv0Rq
yj/d3sOnoEvtqGTB3GhzrU7x5t+ZrzAAo5SOSlM26kFuhqLkTiBy8yWoHi121Oxc
5VjuogoAjKZCVZrd3+gyVm5DP+SgPGVlVN+GVE0Cba0qrIalRtPD0osTS3v6sikS
YAeY8K1l0Ir6HhGvKfrYnbVLiWVPM+Vf5ktUbEv/LX4QEwXsrW6Kb8UBZkn8rpLH
LMrXUgUNpueZ63rF5nVCTDffnOTDKPStbYQoZpe8tTJUfMGLTgDb2WbPdT0uWy16
QD0vp2sQSY2nQRuJmTuJiJ8kFmiE6c0p9+XvE3kuiSxc2TVJMx2s068Q2LWfQfme
1WEZ23KULaGPeSbOvzxwWPA+KOV9imuAExYsZpK8h+c10YnlGu6gAbZWdYwWZ5Pq
FW5cibYKlwdGeo2XeTYuUsCtlDpqJrMW2zZM4SdhksSeaIj996hZQ3+TWYembIkL
h/creeugqi5TbiF4HAdHavi+TEe76ZzTH8DJ1H1/LiA5G1/YLwLCJLOG6+/+ZsxE
RlT+T9Q3P4+bbAZBbwIPpa5bIqrZ9hBIALsXdSxH+5uoU8L+96t3gqaq5ZP3zlGI
ddRGwjPfTHateE0P0Obf20jhy5Fej4/sN0xL/zItaKVEXOT35COprLpz9vRArCYa
lxF96/Td6JrMMYklq5dQ+sKgf8DuQhZLqUkgVFuZQf2lMVuhBpn3JrZ1gnvlbtRA
eZTTijyP93M1OQGzkD2+nBpeimu4kJRr93zZm/7dPvxH9+tGS4voyT1UOsJ2weOi
vFveRCVK/GnAH7QAPvwxZmFnkob8717dd0N693RRIzg6Qwf/NX5nVLstTzvUL/Ze
jnbgZ56t6kdZKDmQoxNfZWb1NL1mi0Jy4SQa2BN28MOeFQPP8KVBqD7pNcDkWmK2
9x0IzKybEsihKSTpzWXapJbJWHmdp0IN/AoWeviNomWBZwrS23FXxDI+i2R2EL7z
ndGbknS4HP1pJ1lC7B5zqemY9p+IjPuQu9aiVy7D3YaTU4rCCD1WGXH4fIPZDbdZ
TLkEZnwJcS3XTTwXZYOHCSBNjibpbYz/6llMYyhwDqAY60kMzNMpTvIX3MVmSDgs
vu4kDsJcCikg8YRlwB0NqfvPXDBhsauZIQrHcyj8srqwAew6uAGBhYtFz9Ua0Yj6
TTBiF5Ay9tBpwde5Qo9QR8jClUWfCU17cq+wvcANRZ5IthlFuvQPdb1yKVqaMP47
x/F30T1wUxqMmShKHg15+bi99iVR/WmDCb8yMzKcUkWHO1E0u0y9jLYyVLp2RATd
EXGSy+XXDNxoopHspnxmFdihjccsLyHiJnph5bZ6p1UudinNdRSDV9783kK1KBGA
y3tMOhUBpkBsO1qcbdYew9DkzNveFn04oBtQ3mUc0UAFT5kfFHlIz0kwfK1gvM5d
XoKRv0MMt+xMzlCo5fZfmELt+165IbXTLNuXl/RWzy8wXnYpzYoCaIIEZ8FGdgqF
15Z+4nDMCZTBAH7KBLC73KNqS3In1XXsC/lLb/XuMJvH6CzSQ8cALSBeW5c89sqL
tV2bQDY3eD2BicuCm13H49UHpCLhe2sGqPD4WBYZaWpbNjuP3jq0D/Tjgg/sElOC
O/V9TWMExS2+oZgtSLSZjOt5dEX2WPpFd6UuOp7HAi4vjAihLPxeH3GzVk2CzTRc
X2eIyXQG5YN+VRejnzcBys9EdCQVKnnKdmtWvdSZc+guace0hCQJRdGFDtTZJc+c
PAlNvsirVyiSjUhE7fB8pQ/e34VptJUbY6zrETWzk4bezffLVXmdqN3wXsvMblv+
K1UoXbcnJroPJ7GUE6CBggu8d/LqaBiGUjWFu/LTgw2vZcxKfLEZrY28knWWIu7m
12nl2gbR7tQKr3GxE22LeHdSrRmt0ciDFi+s25B9OS/R52kBqsvAIe89JkmrdicS
PWELwppkT/ubJBJZ0iCkRty/AetbqusiCH7/NW7QXA3Q7QNqx8EgUd8rvPzoj1VD
YLRKiRz/eyzc/gN+nLFNP27HXPKOTx0zrHvcNRcbvnCaQWy/oV136sbkUG9UuVU7
i1htJQh3WSa/9NOtogPsSNpJSaZquZPXtvVbNXIxjqY94g4ksqUffYvU82+wOXZ/
agdXJn/K8v3/n7dZgegBgFHMqLUCtIFxdaGCf5GITKSG1AEoSM18EHx4XEjJYIwu
FH5JwH7ovYU6olPmhGpNRYr49AN5v6AM7CoLqIgfkGNNColGvL6aoY9tIJllS1X/
J+8pX+bLT9LQkAtiAQZWcoeQnYx9l276f2SMc930oBuexnEYysnHgCQAw4EK2An6
iA3ZSG7wTBtE0thCDi50tl4sTV7SSBfawmOaiHfdWP8xY0hmjjqn0UtGqpysl1a+
wlkuUIs8uEJALYsgLFAUHv5tfE0khh4aKeuMCztMyNxD255q/e4ViZt5SKbcG4kl
GIpa6atilzHvM5+s7E1M6njIV7s7s2kFIQBOW/sKmKUyg0CKfkvxKAQ+GPBPYDyt
MF6kvGjgBxPBIEKpagGTRm7JIEThlQJPW/ELbJJmkQza9Hp1SmVp32NVDtgH6Oxi
wHszjvkHmywdyo0y/apVHakH3gOYJvXxuWXdQfqD0egOSita9HvlQIDh6OaasHDm
hA7IlYpAIyVGPKywBIbaPsD0ffP5Ow7SCA5EdlO19j9BKz+s6IiCmabw/PoGKn5s
oVRTnu4EU6WcPoiFzPWrsrxhw5HQkVolcvFdrkcSoYDx6sa+Eui2psnjFusYljFz
DCXU6xyUY2vzuSH/pnM6ApPh20L8ryno9fy+Y04+v6B0P4kgGBx99j5U6Od6KYIk
bW1rzOXyRHYgKfmnUVJhM7qauYX/XmfeneKfsDbTRvZOxdK/TGohoFPUxbQFdQmW
DOss+TqUk28YbSrBGSqyLl57OzUKAhhEamAjlOXcSTUI5PLcdOm2e9I2mDcpDYtL
mcE7xSc9SniT5yH3Kja2pVRo2/kEjULV5aZbkhoVN111BtjFE0rhuCjHqYXe/qs0
T4wLbIfY5vRlh62ml85RY1ZuMuicA5pKxMo6nr0G6XCuIIL+Z1m5MZbn56HuZw+9
1TysufORWYB0k6Dngra2pH1l2c5IG3/W1uXKSS5HXQyPH593KFt/PBAdx0AQP3m/
mkRMli5K8UbROqRHASJUlmtZVGtCgwgDfzWCQwbrX5KLDsgT3AVFI1yjgwJN3iQb
L7A81FR4/77t3/Pk09D6Kwv28pgwGhZbgglXnjcg0LOD7ZnK7OrZTnpO7CIJ/SAM
HsLoueU7vd0Uv02ewyDKWpjMm0g8L1DZq57WdRIrA9PMpsN2CyE109+o38cN8fqD
Z7vqClrVc+wXw7fWV4Rnzw063U/Ta7ak+DNRguS/J/AtAT1eqiDvTW6nFT578HQ/
qaOkw1ab907i+XDG9fYkgNnpCxM7SClLxMH5EoiX52GT3atNH9Y4F+etuqzCL2/S
J8LXxi2PYuTXq+AYvegSHuxlRASAybkpdRVX4ETtFqbdtQ+UjuOteAQBDyRs+KSJ
MluN2lUvxgFKAFpA5Vh65Cgt3CJvIV9EXxrivArLA1jCYV0X3O2NKwqFSLpEtqsC
iLDrHjPkag8M3nZFH0B/n23QsfULZS++KUhzXakncQ8Y+nXyTPMLmzEikcaC8x/n
fW+ckHMqQ7/iQjC2Gt+ESmDt9gir8ke+oCBFGT4rpH+QygDBz5rImqTGwAaKGAi1
MSPyQ7cS0x7GfTLDYFsCwF5WMTHA0fueTI9cJdJynyVcyg3SVvVpUGLbWHV5yb1X
OZ2YEgfXF+d5ISgMXx5ZulgXXQAbs4DUPPoRg9GCFiOdAOS/TkAUwnioZHWE/8hv
HLuxONVxyjbLU7RESaCi5xJIPuJ5T0dZtPD7ROCqpS7xWGo+DMBbBCPQU+g56yjb
o+I6ZQbqMW8UHJMQLOM5CiD2rdEbrEsc//Szogt3xfKNbvIpScn5Y+XDV96a4iaq
l213Tzu5t9E5jcgroohqJx0nE7PYKZIx7h81JQNxZOkkwAfiiV71xgdF4JkgeoFR
UF4Yt/VV7SncnDvESH+02uy2F1ICCr+cff1iwz1nds5m6jzVhBIfUMzveVMIXMpn
CZPEen+ozJ7z/TaQ/mIwsHFgYSX8yMlBPPo8tMUDeZeRCMH/3IEuJVALj2cUJCpv
fyfcaDe2XdQVbr8cSjlN1MIbMmQIlAjyGI6aeDLaEfzspTaeXcWX4mE2EMFoeEkt
lXKpsHhAWC6DnHKETsCe9EZS6iq78goaLmE9t3AHK1lfVPMIMbvBYAphbWMYxsQq
34PQBGgWOgWij+owAy2Ee/xMoua6ATHfbyq1o7SlqoJSl03d2TqqGhY6e6iQ2hwD
sx0yDWNYFClDlG7XZym6U/gDaJjJb0nxzXmKG95bR4JI45Fk47Q+cbpq7nTd54BN
w/kY/GTqiIy++f1JBfCQie7JvF0CBDlvp/VcdPfuX3QrTMCiUJ0K6GbxI5J0XtsQ
/ROCWfPwMtXdw9suVBoUkhsb6k67qXEeJpuKMmimTsn9b4zsyMAZnBmrCK1hRfF6
I0X1MZbr1tbWkV+qM/gxSt5j2IseDxfap5J3D9iS4Tf59NiUcFg3kRdBeiyEJaIz
TlOMr5bEb4tKsFbQnxQY9GQW3OetiWwOAwh5kB9uUGKtzcUjeV0KlFVM+yperLKk
ZWF6VtQPMpihbf57ESHk60uBFH8BuJhmTLg+gePlMeh0PecdJ+cxaRgxjkNE4VGQ
Tct5VzxouZ8IxuB1BDSHBupGgqL01lDVhOD9vb3J/sOsi7wfLmGpgvGxb9f8jBis
9osYW4j6kE7y5Z5Shs4E3kCNqti5rl16FI9kpWXjKTpFzL+haXae3hv2yMUD+C8u
J5EOP/dHRodfRfHRwqwTEHW5CRBmtdV5iaG1NG9g26nHfBcfvYbyjqUqimvcaoq+
a0qdZcR+Yxq4Nf98KHmLE0uE9xUGiwYf/h/VDAZ6qG++SrZ9wvWztHRWP0VQTdXj
yMJswChjYOVyz/IwZty3/tZaZiS5NawZwPdywg5pGHKAREWrZJBzeQHEqNEoDNHz
gcA8B45yh440yB1i2W5rulJkM387LYx7DM7t7j1rHaboKUHcnYVwFGx3tSdQkMwI
Jq+G0pcfbRQiRzYtZH+yXNSRkwEvfkEBGazeoL1cuVB7KnMHL2d6OZd/4cjcOJ0P
wscqDWQQFtJBDFORyX5ucMT0ngI3mWewdX22kr8K6gbOcwLlkDK7BzFNR0ThWi/P
ZP8F8Vp6G4WZ0jL3hM8nY7omHGpKm0hGV+yRA5jGP/8uEygLK2g2/oFxhVPl6aQ4
8TVQEq4CaelPjeKkHjHsei/KHP5HlJqBFKjdfRDqsC2aaT/OODewjy+giCnRcMap
n3QgQWNsSum2gn+yJ56aztLR9ZiREHhjc8K5Guh0N02kqr1e8ze2y7LwAc0cv9BE
dBFB4AGqN13An0uqyTodu+Lq5BMaF4rvlPTp2iqPNBaJ1Lt0Av4K8whEik7W+gUX
QYhe3HMPXXxEutz/ZeiEVW6Rf930LNBf4B7UPHBffQQ2rH64v1t0LR6JZHyKmIl8
oz6F/qlV0IlSaiLZ2QclhKAcFHvnsrsXqsyL9RoVBEzyg+Tujx5bzwdG0lrlTLPU
r95fmVvqWLtLUAo/vcFH9YMZDmqVTa/iRri4HChUjEkhg6Zfc1jQ9hsWQgnYKvFR
fM0ojHS/neK+1qNg0rovsnzUNHUfButLOWyQBzjlpaGfuDwbepM9mumc9Hpd/JqV
8acX5cOEWiKmD6lxdxb75k9NuN9VDSu1135uA4x32gEbQi4War3ULZEPCgpIUDkM
ASpJ4nHPMLpHZGYHmrhpI4zJQayWKQtZ3byunbKoQuSK7UdZjyv4JVcLEUDtyfGM
jB4F7wieXljPnHntQbwZL5lZjXGJ5RLrMF1s2xgLSs9WofoL2cR0XLySgdpjoIns
Rzsj9IxVeCMtzwHnQlBtRUK3Vj21pG1b893H29jme5G2/+ABFUIta1BXYieDZ/Jv
1l92UuNbjPku/wl1guFIhnBxAZYnd1eMH581WrAVJhNJpi+ZjKq56pevV8O7iOlr
RjClu8yGa4BcbqtNCHNLcXBYDKX4iLLwiUFd0u0jfBcVnktkBNHnzWIvYEjixZrh
4hnrxffwHBZN0tZI+ehjXPoJjU35//meCyjlwvlXwjNvPr4ZjcZ95apmI6F9bYsC
1FsSG+1M3KiLVJXzPqLhk80umYjU6NwT3OPIh4aNhoR4SF0RejuYKQQnpDK9Qy/P
NVklKcwjYWlAXr0AYKbKJUxplTXV38ZrvQ2eYXll5MoCVLxe5VEkMHzRi8kNQe3i
M+A+Z2ZXAgKK/Z25+G7iPnnk38xqy0ARDkadXDUv7qre0y79DgWC8XFhv1zwIZaO
Hz30u6+zxN2tHmAIdE/C1QUPuZS+DhWJOhoOuNPIqi5n4zO1h5y8p2lZ6/qb2MZE
28r6wJFjzLajrmtwaQh/zMqKOpj3Cuqls3PQvDZHCcr1/fdtlbw30V11YNvNRSLs
TLU+ddhJwi0C6ZJFyWsNcXSf8Hsl8aoPckvCDy/7oOytAUCIDrI8/rTgfKDjW741
ayJSlSjf48ImypjuXEzHpdmph++LsimWksP3yy8mm1PRJtNw9QL8pPysNaJwWBEt
UsUBhD5PY828lPL8Ilg617pLJWGKIu8ZRRvIJKB5Str4bTTLPZmBnREWFkRpko3t
18y/iH+7yBybiS3LndxsVMKheQOY0HxhguVEI+Zbvtml2AM2efihYv+wJ8uwPe2o
Sf3ObO9CmAq4zPVca72JKF9WpRGRDG9JDFHMsSgs7Fx3JgNrwZoFkhsFA+h3FcZq
Pt1z+FlWvt4LzRkmPuUhCSaFO1jsFlQzyxZOpzpv6Y5fUO6Zy5SxIvWAHFudScy9
/IX9tWl/ZfjMCNCaWUdoeFS3e0N7Mzu3e5DrjiYIJIPJfnZLzrKux1arGf08IDe6
s2eEZZdgVm/bdNrP9jOdRjMwe+qREMp44YfpzpDHf0sO0JcVXrCz8Ku7sE/qDiWo
t7fyQk+6wWR1eB3yAqyzUOq6pCFHvpmDX02n680LUy7+xyMmv9S6/+CGOHATL0J8
SeQOdnRGQrwX2pfn4Kowb9BJpNMKZ5Qc9m2FTZDB/KTxIWRW4ApZFno1tLkN33wd
ovwWn24PFTQ7kuA7Gd1/sRYqJnc0eUPgsaSSNAGWLfeu7eDQg+FzNXP8xmJETS0g
6LvZRYINCZKB/qi7nUUoL7xEvvfq5gvZdKhMPsbka9lmY+Co5oPMLfvx2xs+7x2C
CsUjLIVX1GCaF9qDN4E6JGnu3w14CUYpgOUpNYev26TX54N0l+ToHA/a2ETXDa9J
uhTlOPd0WN70UhwVvX4PBvcv/oJdp3hYAb8H1/L8VeNXofHzh8+i00bMk7szIQSp
7blemL704kRFkNdV+cM5zUdz7DEag06XXQGahdMyA3Z456nwwi0ASNLVyDbePJK4
7p9HvUziaHVE7gAxzXOA43kVPArAgKAydr5q+Gi/RI+TRxlcaLhuoVAPS3ff2WNx
mzrzhnSK5NDjI5LTWSnxIu25ohXGWnmU0A+GWMBmOmYuH2544PSeimj7fKpLD2sb
XUHhdzXjrbUS359+3yZSlHT/894CgMEDJFLmtC5d7fRzxq/51nkckGsjaLdS3Jeo
G8eGcA0VNHgk+6DYylhL6CMMqSY9RYamnrgj5QnAuWNPKTbJN8mqxbmKeOX5+ZNu
v8719RqRl1dU4EhFDyp2qWL9xkDvfbaUsgFLkB47o943gHgXYNTG88xX5x5wtIQq
VdQjM8uiCOSd++thZc53lLpTiP8GmfgEatJrUG6nrq8hk/3g8KD3o4cfNglQSz8X
UNnhX4huV8GgMUYOJJOvKcx+l9E09MYcRrdIte52uDfIivD9JLDsDpjA40++7YFi
bFrtp72Lr0twdfq9F52Ua/NDJEQXAnvg7SGFURrbKxPKODYmnM1d9Pu94PUj3Mx4
8r1rz9rVZoIDZLBQxHbu7LSNePvcC/RHj0UQ76r5EE6lfiiFyvtPa/OoSSpyPIiy
lApGegimTLDWi0+FfwIAf/xVGtShR2toU6F/0ZYsjz3fnm6GMbvWS4nT5DvD8Aar
Mu9Kx0DLWVj365+k59jZPIvbdbh+xoEA9HroM7O4GTIvWv5ob9MZly9QXSQ/Gjhu
DpMdn7AJ3aQjdR0VjUDUWg4/vqM0fGsmwrDcqanCz3v6aWUnxTHOVVsWXWEzPX7e
wzWPgrsr4Q5l1ulR7jCshlhT1YoH8ng3Aa/MBxzYiVAGH2V2l0uVkwpxiePokvtv
pBtrdYkZkdkWVRWfSAd1V3/PgCtVegPdUFiuaV6MqNaULyurN+r/lX57ALyCh5/l
IO267MHp65ii7nPf398s6sEErlDvhaddO+Av3AtuIw++cg6ez3OLUDOC1xqPXi+i
XDgNY3uWOQ6ZhxroZlF7dr5oOS+TWc53zxfcbvukcOr2iSTgFck1uddOat1yo4il
RaN7xMrSxpwYDnYNo/jYeiObFuyxF0JlKsoVd5pRjX3XA7jFbnLZ1CKp0ag+bWMo
ZHpJaC0ABJIuL3xf8QNc/Z+JSX3wN2BtbRr10FArOTRHtDxmeqTSkImv++UlUchU
JmBNSNZ06g2U3VwdTf2U5FOVONbrSQNX2TmaqWu3bHlzMSFf7ARtMYMtGvA+tnnc
uLRHmuD1TGz1g8zO9ybXzscBotmsYYMtNEBcd9Bch8ZhEdXhaU/WBhnJzdWkg4VH
/Wnn/58aTDs+6O1W2WT9iOuTbvOFHmSe4sqoLs9Lj8Da2mejYDGkuNO/knh+NaMQ
xA6KNEGAJEWH6r67RTIULKHxPQZ6DRsqIPCQS6uBaygp6v0zg+rPa/h5L2TO6OMT
ueOIQ7dWuMziVQcEAj1k1HZEgWYb1R81W1GhQq+CIeVech2M1ROC5kpt6MfLVCYK
mQV10z60Inbvgu6fGFDUyh2nxGT4BS+FCPckHcu91wr3j2YiDfzkPI57Ox+EbiY5
fXDHnCuBdlZthXDXgtAy6u/5YI+EYCmc0PgEa797h51IR2YgdgJDXtczrgCn5g9d
34BW0TaffHqetJsDmNsk2MYP9nhFpySh+QLSgEmVCbpJASNsjZXwsWfNUXpLI5IJ
2MvhSHR4phrsNN8fMXD5/AFcugAh3MMsyTyIImeo5AhvNLj3UL8VnONQ25EZeTM4
zd0WL78rwQYvIoAUpbioqGpHbEmi8O9Gu9n1OzAG+a1C6LbLMYQxsCioHycKuGDD
248ytmXW9KGCd3e+Nxs2tRBMhh3RguC5tY58oGqNWzz2/jfxt26CVUdXwXgJa0nM
KfKC+Rn+CMXIBVUUtvQuQKnAsNMhb/zsLD3Xt3jBQnTcQk6KgoeKfYo1JVesN366
SFzq532OO60nRRZghlyJuOXcz0ME+Ro7OgZoWLOA4ajoMdn/MRN0CWofQphD1fjx
QGMnrIotyGpTOByhBPzrsZs8LmKfZWrpTZ1Xa0eSkwqyBDPOzNAzhqOUze1nVcyx
Po5Tt6BKv4cyHGaEzUqJzzFjxf6aVdPg/AXR7C0ijGG4t+MNeX7g8j1/Z7IeyLoL
cl0lWhpqObKqQoUzHH5kZCojLAN5jM0JKpl8qNe5DAEKoV64Idq88Rsshhzir16B
Ipm1jn3I2XP5gsqbftUjl1BEzow0814bvzg73YDIrPhagOkM0pckilS/c9MIuzTQ
ENoFfKEFDdbrrAusXwdn5NqWAnqIMIIeNnzuxXqNDnya8kRxfZlMMS5324gjVz1v
K0Ldi/Qv9Fpxn7UzXeaAg/mMNLTqgzfbrURSN2x/YeuY1XV0X3htlE0YXk9M4JT5
LW5KAVU00u0rO6svXsS7N8jGq8gzjPNzrB2FMWoHfTRUrLqVf0H3YoysPBhs92OK
5gqe5YVQtp/AeLzUgmypJ/1i9oXerumq9hz0iFBelvCSvJpAQpnjoVQxHvBuVUED
DfJd1MhVxD6Q7dXvwqThRdD3rfdIC0IPwF7yfGi34yQv0cKqEZD/biaa9NldcUy+
AMyWrDQpXmyJqIzkrBddc9N0Z6hPXoabPSdFnIK9AzQ0VPNx9EoLN+fF3u3YntSH
jMjgjl/2ahRF3Xbm/WNFnwn3MKstPbQGpToMm6ynQFAUMoTyEWZGjtY186Ojkwwt
xB7CSJz0q2wgiZTCG26xyh8k8vjgqx/26zlZ+vH4nd1Xo4+wNL17s6uclHVZWIiU
Nd/NdNsEG+y8CnP0x5lMT4ausDexTs6KdPCOxYg48PmEY6TmTYEbC2cW7ZzU1j1s
GL750qP5GtXyQcLoCNPs5vSm7Ngvt6RTT57QrQSIBjjwX9FvadepfoMCo1Qy+2TY
gppuWaagmZ1Qblbp1MdoZEkTp2klh18WdKMYQIjf29JNG9QLoTqc3dvw+7If+Po6
nI8V6udutsATPjUjBYncExUJ2pqgt1vv9z5XpVQ5XZdPi+Tv52/Ya9zJPPL7/O1b
e6cQ++E4qkCvbIpLGVLraBJEwhMm/PA9Y0eXf/ALuf4FTQNlA5BWIJAhUri4I++L
GuHofwNnJgZVVRsVhFf4b5XHoJddO0pUiVn5rqbkgePwzTqOX6c++ySB0R0k3+TU
sUgfn9KrKeqU56e1m0+AXndkemaFtm9Yl0S2EmwNuiTctaGyar47bbi50Vpq/6vq
dj3AisrNU48exTBCFFHYnvkfw3w0dQRKGTCe+jZleeMackvGUCAy8z6bv4RhlBjD
ZBvJP89TFtVZizCHa2YvYAQuRN0+zj9G1Vn1RsxhMQF43fYF8mm94Tox5l5oBxcv
+rcLsNRGyf8dAUjQ6VRpvo3JOMRzG0SeyOV27uuWlqfslDBvFRybQv/el3rwrhwe
JH3EZf26Cyw3W9CKW5MXGb9eYPtCjKcC6McfqQKAsYH5I7nOOJxCcLxYlIHTL+C5
0juxTMu1ZbmfF0Z74Gkzgsg6eQJx5YL0Jcc2nKFZGTX+rW9BqhEkt7smPj1P5jO2
KB/ISdJSwQRjZcBbAQvNV8YMY58TULyTc7KMQi30tU6oQmUCaKrTjq4IISolMU78
5lsxD0Zxwpl50KtTTCnA25dMt9Lb2tsCjSNTsn0mIY8qT1/2lCIh7ZSL88NvlMy6
bR4e88uTWSA3HikPUd5Rg/j10MHG1GvL0ndUNT27p30uvWfJd6lqyY1TIN2NLJdL
WcZNw8WxwXfLB/Chvaujs1hM2/Q3LRqpsLQsGL3BNx2yN0M1OjuUrEOp4zR+DWdV
OSkT0KyYTbRtdqUnKRemZ1ZPiSeqsZaGoodrQhFtk4B4VpevW4GMi+b0D2P11/81
UqLtHNGuiG3UJLfkE4uSvz5xH1AxfQPKQ7jEUhDPMRpXkEDzuIBCCWeVDby/F+Bs
D6P5keseAnzM6yw4tlPUJLIjfndmK7aPijOcNSA6FFrAC8kA4YUzG2nFAnCmOaYl
CkzKgLSTYXQ0zGdZvFSO5Q6jWhmL7+lLfDUNIHKXj1uUpqPMgngjM7JHas83l5gd
N4ym319Rlgm2sTWcLU9vNxNYIAr+k15oGUu+SRviZyj4jW4PvZwaDNGpYs4+QQ7F
RGrDUbYP/qwZ7w7G77iXrxx6Ss/J3Sb+dqioFN4EQ+zLT56N1qM/l9+lLD6tDJlF
iTpUyLu1RXKoN+UFj6Do5qN53120IX2fEyEtitKvFoVCzkQEeTJd9S/v3laRgm+U
FYi8gRTrt9HaEHQK+cueth1gebdVmRGTdjLcZnWwZ75JvXXPWD34Pr/Ynva+8Y9U
GFK7T1zcro3pHgSh7QYjzg6G9tjWy24/n7bn+lpFMJwl0GlkJwTcVpa8H2ueEgbg
2Wrdgbd/N2PEYzAm8I7cH03Qq51Xfz/LR+48/VELhQ46rN6vgZ4Al5HOG9AwnZLr
bNi2qj5qRK85Ou6WUJiLeidH0afMYUY/Nj8QNDAAoniYh2xkSME5qgm+UB3ftE43
FBv9U1kBy8p9PY8LucoocMh0gIqvJmHGxQI5dP2R6zf9A4Zw+Hpb1r8P58owKxJi
iXAgqnMDL96WPTH0B21nH2fZ3lYavpAxG4LLbaYT3STCgi0BhKoD+D8l8T/Mf02k
LjeaipFkFNR/U9lQYzQZM3wfx1+JkbF1V5vm/JW5x62LN9/ObcI2jQJYv3SZzaJd
aYzgwA/A3/ksSDW+GiAQbLZGSNh3u1qQemXptqLSIq2ByMzuRGmtGgeQchf/8Q5s
GNDVm4bsx4+75SXuM7Y3/IaGDy/BObJGOOd/FDcOorpzPqzFQwDmaZMBJrGGtRxk
zLnGmJfdjaD5UxQH1s0eAErX8Vvu4BVlnkG0QrJ3zFFmkUAzqlmu/P4LBwUaHC32
YkdI+YPrO5xHYWDYcm5f/eFF6EP6ITKPeKd92YMXakYi8YR2DanDD2E5gxS8Fq/0
nuG8TMlsMeieTxUWV8YMTSEVaxgLH2VXv4QUBt1hbbu3NnySF1M/0us12uNqsbVp
AmE/igAYkHaFqkgEGP0mYF9GVaY1IQPwLNJxalA8Iv4TWtDpKC6Zv1YTfUFBOMMg
fTjwSwknNVJ1YY6+4RkWHCgDWguvgkZDSAOcNxuB/7pgA7ZHOwCzx33tE6orUIn/
CGiWa3tqhuVUWjL6rmDENYH5Jh+NpaiznEvI6BHv7cjhcru4gN6tJxrjUqUOwuLA
HyDS2OBwEenTuJVFTt9t2mzxqo7dkqXbYiNXBaathe3EmKEUFXoGTMBmoRG5/U96
ycO6N8iptLe1oShymYeh3SjwZCTXKKUOGRTdKWO+MLlFOFHBOFfijDjvj5l7m/8n
f8PWW6YJlwZ+PGdo4Rx8Dv+QzXibFHpBzv5SA4yai1OHOAVGzta4GyJWsyzuP0IE
XxYfh9A02omcYQHQ34wh11oIddYcejarwxBAoiCVTxozg6b+XObZnhINWQMFHWKq
mLQjDmVD1WG9GauGICcvAzihHeFXa/GOCAOQmMHTAFQ702RZMGBMxqPaFiRswpgc
19iUGDAHsJLpJP24RB/DRpXZDwttwp2Gz9+M9ODlkMXg922dpn4wbTtBVpqIV/ci
lZc0K/jq0/oOuHjr0QffS66lu0M/VWOmZf0yRJEzkPOUyxUotTidcMPG96QDrOAt
h/N7Nar+cj+Ak9ZzuSZ84UW0EVcmZXAXo2yCeUmGeVvuaSAfFiFeHU5NbSi5sIEs
M1e7LCCHlfkGMT4oHnvYid9e4+CaN/JvwT7wv29+RoNnnHsVNAyz9bpQwanBfnX7
3QbjLGyJnb4pAUMfl5vrFZq+91MJxjjA9KzR0njcNQT1OT4O4kh24x6BUGjmZSqo
E7AGu8xjNZ9Z1r/2hWhK5cw/C6rOz2OQi7sA4p+HQgvzZPOlmbhXFseLwcNw3Z0b
d678n3C1KDoHeWPavCagQ4dmOvK1d8cvfeQm1DANggz2UOjZblWifU66bnTh+MuC
XmsiaNILZGgUL48kf8r1V7pFn+JeYbVf6s0hUlncONClKb7WhOQYcPF3fentMVp/
oKQXcIqvDjUzP2GYKbULKB1rKlQ8lo6S33559DQ3/5l4V1Xvx+dV7b6X/wQ3xEsN
frhp8IzTF6nHMfENGwQmQybf2bKLGEUADQ9LMrmbH/+R/tIAJAngH26KgwqXCNhc
SFkfqzNGax5onCvkXmpVcugidnif7db/K5FO84Jc16Sx5hDwvADpaRUjntX/TPyK
BILVMiJC6cL1lMUefDqpyCc59ljcdg3Iwhnbk180OHMpiSryI7DyWy1wIhPkBxst
i6JRT34LT7DsPq7wgwrrTx+FZP+oe+EZM9vwrlhdEnXIB9jrNVvq90uxaZzEg/aw
mh8mI+hiRVVb4e8vmT8hqp7RkfNm8Jp/kCZeksyfS8+ojTuA4A3L5zgU4T9o1dko
0jR03jb8Ipq15dCndr+ReHHK7An18vXyikn+MzlQMYviKgBsxSxWlmpPamnQgBRE
rFUMsCKxMfXLqkucfwdemsXEbd3N6mg4ioyUOHncskeZ1gc6AWm7T7Rk4uK+Ta2b
LsJ1SzuvTjb5hjN4YUhD/WP0wF+yFIR8lRqL4I+tOEUOSXOV0ED95C7aVL35az9M
J8YH9WLPaTCB6IWJTtWCjQYajYMN5qw3ozcWZgPB/6yYKn0F8Ufup1QI8CvcEapR
mz+SrbkpNX6iE2cd2qYJsfODM/RPkjnYhUFAnilP3sjfx4snUY5lF1/SRtaLo0s+
VoDoyHO+eaJe2AXArs5az80xOZ48qAA2Vxu6/ynh8x7WmWuD0i8SDY4qXXL7rfDq
yUbp7pQqWzggSIbOwM7T14ZJE9QfLIA+mZ5k0XPnfAngegTYbWtaNloNm5TmlbSI
a9xgo2tHtpSWoQ5kjh4r1dJottZP3kBlXrtrpjBj6ctmB5/XjHskWBvd3Ruz0yQU
3a7XXDnVVcyzKN73H+n483aeEKBwkHvoxW62BiN47iyfpZrIy3EeRAkp820epAOb
gPwX7x8T+SWmSYC87axmf5mUcdIqPi4tnvrJmjcMawf1RckpUP8HoeeWfzyUZnfK
rcp/Ex3JamUjcgkAA/lNBsRwnRoNsKVVvGcPiVmDxj3AxNZtyl2Rf85IhaghPfqf
UljlRiziTNUFMtjbNF00ipU/Ejrlbujyglp9XUak22gimJN+v8EIpZGS3FIA7nB7
qW7wddZBFipI14MQc6V16fkX+TnVlH6rmu6fPIYDltjN688e+WkOOYp93Xmr26oB
ZL4h+K3lH+WhP5NNkHfkggp2zsmlDHK5EkbTzVmLW7O1h0ScWK17N37G1c26ZnF6
asb7XJmf60oFBBkjnnSCb1TIHUWP/CF56b9b6HQAaHh9agkNDdK6VXlpCKXn7orU
Vv+w5GMuSSkazAlXdG+iQvSoCVDoA5ePH3ZKchrmJBLh7UisbCo8qce8EzuUTKwx
FhKzyg2atpL9zq+PyfTY1hWLvOy12GgbeV+mZyNydeNM5QQ6Be+6eJhyibhAoqRO
0VR2ikceTDjmrzLdZh/6kpad4nkv3S7+MV/PVUeNiJR4MP3V0xDQO5uuQ5s7EC0W
QR9VV6zgPEQAzQTBpTSypbyRNbq1ukyMO1c66UTFKRkSpz/usBfwBcJrEVdPlOA4
cBAfGqC3dh/4uRzB9nr5qGBUteiYmz9qpiNY/UifF/WYn77pdPgEx1HKK+dSGQBY
vZGxMtLa9lvuOlIW1DNO/nd17wEcEfwmHVFJNERHNGJJXJlmXS3Sd4QqZAvl8Awk
x2HbIu1MFm5foLauw1TVa1iRvn8vS/xvoAwS3OHHjRryZ6kUsuEiRNZCmTOd/Dfh
F172GOg48lq4J9NIWCzRfYbzvtINHPW2nmwlkAqvlsPnGHqzs1uT/EpWkryUC7oU
2rEHSDAYOrhiO3fqaCQ7/UxZCdaoG9J6EdmpJEyWvcImUZmbE03OLdDs3Hxj7Dwm
OPs7XL4QfOej8bRTafxktnhr43onzolodWgJthbWgPgASaowg2bRwxOPrtbz6GG+
ik/7P2dtMgManRO222NtF+JU+E2WupGILKr4uGJpCOLg4pvnsVR4EDabGhHtcdKV
WOw99737iDMNbxfedany76DCz20msrVZWX6grycw/OgpAtMmcqqWhnGDLh0ebatJ
7POLxKN8O3ipfT6wTcytTkdxK36Q6/a/x96vjxxDLa35FnI6N/EFFIcZc847dqXW
WhGlyckMfC6Ywgy9wEN7XWfk95ZZ2VGeCFgdSvIire90bNJJLNcRyovvhj2AW5TH
tE0mDcUgLzAN3idV+BRHaztmeYcW7s/S3xwEXIs5lS0m64yrOFzDpKzvBUYrPIkr
Y8IZ9mCv4JP7i8OTSRMxbI7FvRblt1VjUH5fxiEf1G0AjN7tyqzF5OrORRjuneIR
OLSscvnpe/0Q4i2yR1QBH1YmP4FCEtJGqQ1QwTLnhQ5a8ZrvP1aYN/KNaO7Z+McX
BZD4dr4Nzo4yXgj2V+oa+AiWEiioewDAKnXCK0QCH467Bedj0nlP7fRms/N3MQAg
TXW/NkSRNEw5ZdK3Xii/hBz0juCOOZFLDrhzSriav5zmGN2F/ck58zAWBcmAqJX4
LpGMVxc4E3MpELCwTxj2qEzjrQQzSDDbtmSgSKdWJSBcaj5RAFdP+dS2Vnj3cBaR
F5zkTN/z+qObXTLAXtrQHqFFqdtw3DOah40hGHhusfi6cBcE2s/EPkE6KL+3OYf/
A9S8HKcF85jTBbgckKk0uhpUU2kblTiB/40+sjwLOmfb4nn9qauEW8ZvUUQOZ6XP
asypCZc4YpBK+Wtt6/1P7aY7dw6ClEH/1qEV1EeBR8SIWk+y3ZgI2FroVlLScuu1
qMVyM6xltubiAC1mrN2cCXISDCkgwJpsS/gESUD/CXSk39CBarzvw/eHBIqRD2ju
sWBslV9+ZCOMQR8ua1rMQYzJKA6F5ZdNHWS1fXnV0F9QHfsKsr0w1LQgfM9vf9l9
GdeEq+wEeQ0YypP2nVGZSKQGdzjo545Ep/sVszFj+qv8t3dl4UcQrkN5+/cEqmjj
LAwxYY5UEKoDzn3QkLeoVQGTfVy9f2lCVnyCyRofZiaVvKrxTG403qnc8cBfCfw6
/ro/hJe9kQBg32t4Uu04BdmwMLvEMR1hhvupUkiG1bdNwn9m+XRZVp/bFqr5OvtM
Cx3LW89bIDl3dOHya2u+Nx6/GcG1ZZBffK2/YFr1CoRjQtwCKD/p7OAGDJU6oZUV
n3j9S8VnsuTxFFMDeuaCU41eS/S6rsKsULbnVLuS14SnZaiZLBoCjRX47NYucSo1
6tsFJLY95aM3gSctaytwAD6W4roCjH2HzDERyavLjpdjRA9uvIHLUmlLVL2HGnGO
9lNHI7rMA68O2jAP5BiC1TetlTL1WGAdcZlxr5VaN9GWXpZJTto12hUDCx15iC4K
/J3HJCaNg6rxrsabfHxvssEsKksP4+i/OoSIcoivP8rwniNwcdFp0el1Q42ymWAz
yuLStpk6ps8khxlbEoBvEj3XfdvFmw/R4xu+TE0+3IdqDwuoirslKZhh6GO+NrNi
4NNtUjfijgNsWu7fOeAdWJ6ejIOiCVXmHPb+A/GoL7VhfGim9flmI8pe7iISn1xJ
weWim0uki+knyx7/BItqYq17tsbNnUKcH6xQ7/B6opqkMOWV50aEoBleyPWMy5aj
TbfHuXrphMa1PEiN49WbW27+/UppH2hkaZMxy9XGJ9ydBDpzd6CxRqM6rS86bEhj
E20MNLUSuSr+IMGNCJRGYCxBR3fHN+vPetg2/wvGlQVzWdmwZ22d24sLtvV0DJoP
48+Q7jc0aalUUUZM+9PPbmaMJG9/+o4TsePhSMCKHgejISZDXwLr0XkJ0G4sXDZT
42gSjeNOXL3gEK1EzXRpraG+jDs9grmP17XTO4zUDj/h4IeZYJUe12+X8zRDd9t5
g9fDALpCoEzfvbS+B9Va5JyvKzRfIjX2siYrX/rQ5pT9966Spn2RNg0tCuttD70T
fAvLWwoXRN/7+7HWS7sIdsVX5lQb4NKrNHs+hhPw599Lczs0syCb2+M1cZV+2o+R
V+xWIPoMnsadzLL9UblMMh9JPXuKatAR9XNz+/kYgKQH/pYOv/G0uA6BhfRc2eIF
K1AkXrzgxkbmgU+TrDr1lQoX1vsLqOvQU6xsZPHLxU2HL4P3U6DWGEE/6HF7gcMR
GXv+0gvHiE6CqvVRN5uRgxNOvIOBPbnHzdqE8Sh5AvtQeEbCQw5ztKXm54EawOy0
jvVM+w4y5Lxsv/cMjwHO+EAjLur3BV4Ugm4NLNxQpP/LOD7XO5IAF22p1MSagZiK
T3o9pzh8HxZtqzK+P/Pw16IdtSzsnmUEOv1+H/XIW0NbZOVeolxltiDKkn9cI28U
4hR8y3Gcdepu164zZ0dcj7GAX1G1O6x7xi7ydChdHHwjJFbg64mMsvXulI+RAdc2
UwRdBvjtbt8dDD1L26X6RZSMRmGHnBypoulCfqIEV47Y/jfBVEaN+jQSMZrHGPyK
TtIbS8ohvvHqDwrlbnwNM33RIc5gUblodAy+yzKZhrnNg/oiW4cvJA1jZc6+uiAN
tJni697SOguF7Io5i1hKOjw2eYa/6REpDOKCJu3CcVb9ogH2F1oq2LL+PQGSqrJB
U4jc6qOvg/LSRVooJtd9OShYqo7f8btMVPMR1TFxA8U0b9xGhLgeFUYrdr+uIUvw
5k4poL+aCsLlyAB47auGbLeKvOyjmk8rKHBb1etyv5doLGsVVgPrh0ubJLPGL89m
gSqAFDbQBZskRshckMaK6X2jKAz7nJLuQFTgUYJco6V/2FYWLW6S1SBp+rKvglYC
deddMVG3M20yUvir0zFs6XGzXbPW2jfp1QjG5R+ALA7Vrn5BpusfLzmUgc+kufSS
M/LdNPW3dIFpE0DytSPoLNUOQKTgoCi4hrqlg4jtwrW7IhJL7SmlTlX+jmbqi/+w
CIbWtcUM24WfQ7H4ExBcdjHMDEje4ZMGVA0kBLJluEb01WTWT9RhNwSyXbeRMIgd
WNwhJbjjHnWhcac9S+tcnNPdWQkjVgdPLWFu/udn9cNSMG9o8KOhQ4Rd6kBd9PRn
5uBYlyYSg1n80TC3q6N00/Db4DHYm+c53/v9M+3UVgSvQF47hjjp3gN4OY5B+ZWH
JYkL4Nr01SCz7hKEqmUqzQ7/YduZOViq17QtHUtJEKjYpzatBeBL3CTRKannb4cW
I3NesgEpBmFa4dO9bWBDQDkLMiMdRhJbCEnOwtc6HY28tYTd4XBUHGL4MMzIiueT
rn1ni/hlCJ2WetF41jSE8DV8nRVrX6JUzcWfV4HEspG0zkXYd5J9gJSdb4wIwN4r
BpgpIfCiHhR621wJCkVqcjUZ+HgO5nWdK71CGE4j0dnoAlUoBtxMT42oV6/CYc1w
hARk8Lw1IeaBhhv4nZ2h3FAPVPwwJiWtcJxxeb4EbgjH+P+OUjhDuFRYEJ+p75b4
UnU+rE5fy8CWrVZKtIOPi7nROO51Og0oJIc0Tc0NVcEPgVuy4p3yUS36y5cesOGu
WCl0fX+oGnH/O3MlFxPICsJ4gtsa7LRiF7NXcU8c4pjZ0h6boEtJVgyfYGT96Upw
sQeHiCxtEEZ0a5f7Z1bR+8cfI9QhiT+PLQb/cgnSJ21KEdy8cVPKtf+GrncK1MVN
/ZXYyHc5m50hZNvT6UVdXI8RfUcfTmbYFr2UZvbYD3iRDlcz90KxnLfSV1Ve2Jgd
P2ZWeVFa0fFL3cUM6pMNinOkH0aQt9h719pBTVj1R+dkDngsV8d1OBEdxIkF6bPO
XYw9jRkINpNKTdDcrfZKqrjxLkOBX6qz+8QVgHE40NoY0NrKb/7iVUsV3WLDzvsV
WAwZEXWFkwbCuHOsdPrVbA04GO9ogLufQgz+kYiy8NSCGwuS8oGsfTHPg2p+tyi9
xJxpIHZeMvcUN+JrDrdCs/afwr7+AYXLEXPORJWU6qB2o3OGNrLwkPbAeKHujSKS
Uras8F87hTqU9nSLDOkjuu23k1hyqlyMVddPQC1VHUMPIYpWfUXg1HdpfxVchUEy
mWyTcbx8ie1VMytmAOGU/xmMGnQN9PBi02Yl5fjFyjrXnMfImdd1fLsnLyJlMICt
YPvBNkZ3q1PWQVVJ9NxluKs76Sef+Dam19OrcbS3cK2wVzxUV6qd8DKvUQopm9Aa
Lve90aU/Hx2v+zsTL+byjcYWJjcMyFEuGNFlqoQXVX2eb9ooc0CfdAxGrVSSTisY
f8EWBOfaSceMUIuIQv2oncZKaIJiyzhJ8Um1BamWvOM+EZTpsOOIS7eTv6+Y6yOS
XkY3CxcnwAsuv2gs8kI8xC+LDxTrJiALaYoV/7HWzX9iwIPkmjiuZ9VpwmwyEuV1
QCQRJ8th31bo+H9JYdQC3ZEp93HmY/BTeae5LxvkzXk3kvnBxdjffteGd+8+Hrnc
ZEbtAHoc0W9AUnBfGSAnEizBZPhQ0YNv1YuONC0skYHiiwaYx50wOvwHur7NvpvW
8Jd2rM8fsb2Vnz0uJNBwpz2rv2CCm+uew+Xjj6EEFXIq2c4eKxg/KubZUTdNuPxJ
+5YSKmkNDrS/UymmQzaLWgOX+laE1zAaYhWNldagYUdk6wkrLTpHJuNDCdGOzi8O
qxWabZND4tGzUQltuBs8Feq1AUQrGO7lf6ATt+OqyE/ehwYCPXRTP6u45gFewhi2
LxZWU1yatFkRgsj4AwAKDqbFb202VSzs7ZYj2uYz69MfTBKj8PSUDVaC3pnIwRcB
JIG8RNn/Vp7kXGTZcIAfVBzhJLkk662ryHMqZEwu5CloQzeh/Rim55G0md4vSaLj
RxoF29Sudm7zaPDLFWyca3vWFCpMacut9/Dm0rg3smKVSDsmst9BLh8SnMnobG1x
UCfTtoJPvvB/VBcR/Bqi+fyhKFZH1umhwEuwqt9MOfXWxqxuKl9As0JITxfAczFV
/bgvHI/Mqgj7/80zeS6Uhc7IAb1LlYQhvQO4J/+GUG9vhhmLWe+di3a+cVPN9mlW
+RTNzIxa8+Qg+gBlQy8V2vG+cMJIq1ihg8K+3XuBNT9nqviw8k5bO4Cay+skoXlg
Tsez9BfyyVmLquGDg+Bl9gRHwVsV7ZHgbs/1zFfynP7PPAeApuyfau5gaOSXUYxR
Oflzc5WDKXrKx2fDeNhUnduP57bM83cSoa7v9pwkbwicbGmN53ExsgRPoeNLV0Fv
5Dvzh/YHvsjjlDkrDOgneFOUj498oLD2J6DgbBhDwmL48XuOEB4RmA4wsB/jRgHW
7Up5XdfFvFl5w2Ksjc3Y2YNylawbwWIGW6ZAicoYJtx0UfuiGfvfhmWKMkNeSilw
T8d/DcUGJ7Sho2PWEXxiwpykpfqRDZKaIKx1ki2WFiRvDPh3U93EkDEfD0f2iX+x
pQ/AVrX8qdHtniyISxbe2QZ+j4nZu6ondnSHVC26qdn1nciGXZzheahFvvZll9bK
5uznPLpyOXJyAiwrXlQBdbuFi9PhLzdUCqG6iM/NS6zrDVXxKKjDbNZFRg0jOfYb
bLa8X/7ALpQ/vp4yiY9ECPpXT6wWPGwSBOQCXCjfgqXN/iH8MrZ5hgRdSMBVxIea
wn3bZmFhDPYMw954mXfCa+Vi51vuILEC38+ylLeQvnEJCYiWDjzPAOqycpQEsQ5w
5WHaDgYqbuKYK0MXxTH0D79dQRgk7EAhSvA9U8osOkxj/7gNmv9yGRGMLCjSGgTt
8ZeOILasMxx6ZO0nnxpDrbDv20so3zujFB2LlzZRJASDgifeUjmepJHgGSrltPRa
Fcken3I1SfF5gQ8TO+8brq+vQMjpwqTpxq+Wxe11I5+zzQvSKu3MgcfoL+Tl7eHO
gOeYEZ200E4rch/K8ZxmSwxlFnBSdG6Ol/YzSKJyeYsG2VqzenOi3pHpqZ8sPbbV
hpukNSYdLsKq+BfPyQm9c8RKT1fuvxuBDjjqqMSmrz66iRXavJkGtxMgB74MvptN
1agon/ic47K97ZMpBSpFBYXtoJZyAFUuGDJ1Bz2bGnOPSzYnSGThspGWNjLI6tVa
ALwdSlCw3MBt/BOaR6nIZLa3x6zmRfyA5uQ1K0K9vrV4VqSQREcrCCQq8sp/p2d4
ib8Lg1X7f/I47wIWIhLhgU+XT64Y5elPjM+EKwVqZ23uNVh0jqewsDOQppfXOm66
P6xDxl6p3bpkP45ytr+9sGVuiMM/JYwZSogLyck3MFRrEbnS3h++mLRh5QBVXAcD
wvkf8q+ql6/MwDoRh//gqifnNPqvCRl9FJmj7rXn1MlDzqbNk9wZ4CD65aLd0hA9
WebnufJ9iANWuDiLobLdWdJQ4KGEa5P96RiMWDbQu1TkOcOF8blWnyLo872efqL4
jo3GJaWDHV8xBDzWm14lf+1zlC9ykUAih/nka2+UCQx4Pb9U3utgWYgucc6yJgsq
NndVI5rIfU0XDnp1F5LHNgB6vkrgCwkb78NgqxAsXKV3hpd+q3nJYm/mwNb27Mtm
I6HUC0B8xiq80m3iBxd9cPJ6cG9UY+eKUFLRO6o14GsTgFYy0pXmySIThp9IgGKp
y/jxa55VbYE+wODhOGksmsL0lVXkaEYS3wpn+CmdmEzn4UY4J7hUxAcfxPR7jame
NYj8QbNydU0OykGC6C2qLBHMg9RbyFVGSH2gpqCu4voMrpt3IGNQT47hXTttcIgV
fG5xVM/TL9/rMgGSu3Ay52Nyyr/BONmYNgEVgQCR5+9ljvt3FWBTsJJ68XbyGqy8
D1+YeQJmKQrCMd3A2Mfny+FIvmUhutfjRdGofpKqIqSEBLK9k2lWB1vRdP7P6Acu
cABJpY6UvpR44MJOYZDEJZBbR6pDB8heCwqaUgtrzTwwRGLUDMCJXDNWzfsQKxnp
UaMR0xcEkn/gPZfWkNrzKvpbe1/duOx78PpfPi/cb5evDvrZLQF/XJg3SYBqjbYA
ER6xlIeiHNzrQcjZ+R6UdAIE53thayE8PGiCqrfI+9vaqqh63BPekM7UJ5lJ917L
60m/XrSsLNAkamH56YJcnEIw6AdT/LN82MPD8pjsmpifWHNjvQlYrrj6HTVjIg40
0oUBMx3ma8daZz/DZJKr+x9iFgXCFjcTf5LMViuGjBFHkSRuXk5SdYq7cK+JqFCZ
ezELILSrYdmJ2XDppiT3D6LBrY/BMFKyodxd8BcnZB3+XK8OO6b4Ng7FmsdXJcn1
ZcH/dvZzTrHqKFi42cLUA9VTZXBtECvG9UpU8n3B20ll+CX2CFsWk0m9W7cMzbfD
7xhfhSc7PZbkhAO4LKDWM9OAIL4q+oRrwZfwId4uNTbj0Xsv3ClUhCtIP/3yatdg
KFLFU+Av/XRtCGA3c1VID3V8T4qAI5sNlEB53nqqKCQPvXumcj2aWID5iEtNxjec
YeRtClnyveKw5PhbseczmfJ2PjQLciTz5aUwDZhTlMTWkjoe0WtUyxWLv+gPYY6B
ESTzHchE8fM2aMLPIjrIzfv+Tval86OH0iFgC6qC9zKinTEISQUTkX2I9KkEHA6a
GKFAR+fV6IIEXUtDiETbqDtH6v/34dTRqPxKeioSb/m7oxLc1v1U2/RnQGpw1DpV
y3cataFHD62vTdxi+XXgKNI5mqiqglV6q26MXUGwBxcK3/PISo1yjuPiRicp7ZbC
qs2EvbuSzt7FFT+CjoWzN7OIhE/cc/u4NuK0xPeQFwM+GwXcWnntWe0C69BxZLFY
Xpwu01fnxgKJco4w1auU+0xwlXSu6VlWRo+YcbL8lMEA8YLq4XmrmW9erCjr4eiW
E7zSMsriAXlFw9t7UYiInBVwOeK5gpNqt8ZL/TRFcHbAAI40J0w9dXuBHKKSk91l
UJqqjtHTVWSKiw/gwEpw1ve6indT+Zbb3lxgtuUCGcn96UF+XUfLSSGoulZYgMJ2
mL/khQZILJdQ6nznzQDcf6Li3xlFt/1fLRICD/A0slp9Gy+ejI0cIiY2fIpkopBT
WWapYW/JZZdbQZFW9xopUfE3lzCcbMNY2RWv6otjc4qU/UdDYDXjTqceqBfm4rQn
Opue1J0O6A1CPZH6zct3sXaUZQiEyR7UusZhJz/JgDCRDVTK1KCXu9I6dL3M98GP
+1OK6vNHcPeyPJj5JjMw72lvbw3W8Y6evSW3ieXws0gmS7Jis43GG1xn9UaMOHd/
dmi0K6ulHVHsb4zdI0t0pFH6O8WExKyJqBA2NIIygDMRV2/SxrQKG8Ku7BffEHd+
ITckffkv4Gx6817ga4LrLPooWhV8fJGmGqh/HzFECapF7S11bOQhBkMxvctkIP/b
4CT+3mih9v1038/QLHNRwPn+aSTJ7G624iLS92yjtMghByn7Kh6lT+gBqysUwIKU
rqNnMcGxmIxmhWA9iGhsF2zbPMPFpbwdm47WXRy7PoOTYl+KuN0crbSCyg9T2YtT
oFhil8nXIlnlnPtH67O2xAxJ8OjVJMDSrAS8DXd1Bocn1lQS3sooRSQYKDB72rzV
wbFdezLVhJrylzqJhN51lmCrahaVIhO/k7uP5IBw0UFHbyOqFzCqzbtpa9iG/j5F
S+gMYOGymdsrTawapsLbkT3OT+ts2Mzh3lqLSNi9c5uf2gRW5oMowvoIyryz8aKV
JKLl8gQ9J79c1eftc/ngtWiiHJaJ0JnA8ZnGeXns3SOvi6rrs25MVxiHEW88UbAb
2L2Ceg8VHZUv9En4xeT2JMKuVklQ2IuwP8/r8kc7dH7w4hejXylvvGmc73b05ZIH
GpIWd4JrN7vYq7feIsaoOrDZYfUESTGKvqBq2MptHoh7lDb8Td2oLYCryY0QImdg
DVoPJ8dJrfuaoPN5w8zBZelnBCPifeqY0C4TrFj7pBhbRiRis/WU/3x/AmpIj8ec
a2A3GJO4LnYhfJzNTwc4hiy+MSqpGHPvtZBjYDtitN1q78mXWoj+37RqxVp3uGoi
9RlTv0XoKiVbfFrbZJ25woc300onVNmwLFa0mh76Z9pxlqsydc3TJZBZ9fBpb9qN
+HPBIkXJ3dZNlvSJhu1K/6/IBYWbXp0UDFL+cwIeKO//jUVaiIs+c/CKLAXE50qD
j0Mf5FI8X1iEJOoMtpzTfyUmalsZg6JVYoOpWM1lYuJdAwfYHRlNlxJSR1lkYdec
VxaScm2HeBaXfeXRzej1xMVcnYPnxB8BF2lY+Yww8gkD+YGGmNHWIOxZ/WiDB1DX
08XJWCuhXgj0WK+ywRRo0L71i5s4l/TrjjLWTK5qwcxNXb838/7cShn+RQPmgYO+
77/jjZZ6fnilE7pT2QSs9Jtuo1g/ahwxdPKKRy5kDawTB2Od1MRE16Ysg0zTgzwi
T1eGw16wFjlYtOoOWtVfB+izbNDhs306AYMDxxfolQfArUrNd7QRzLYqOW8RLEfK
h0eSN12kfSbqfwggB+4bhQzwKEKGUoypzw0UraPmSp+g7hJQj9fI3SYiexnHBiEq
S1IQMPVmI1mzs05mse7zZTboTmVnDNfar1DBluNH2EO9/mY6IAcbVpSufv8fabvy
I9NQafpLHJDn7HiuYEpLTaQJgfHUOOokPJlCUS6ybnNek83SCzG3gXzXWAAhlqSo
jSd6yeyOumYwzCZpnZml6kssp2VcvFr69kbtH4N6mzJXTj3mR0O5PRgpqoQb2Nsp
q7r3Gd4/gg/VUVA5O4k99sAZxbbJmBaCAWNetJd3PiazyTUfYJU38WMZBgw6wDGM
kvVCCJ16LLh1oFloVRE56NaU8IFab3hwACSgRwrYod5/SDepIp8+IFh3y1zP1WJm
i5ZWhPXoGXAWzkqxp+QWb6Xz1QjTUsJBYnrixnw55K7GzYQ/hJ9agA9MskbkZo24
2sFHZTbud3WtsMB74bWWd+2tAgkW4STUV5UD4NNcNSN4fbyysfi7mo1xXga+7/7J
LkpU27wNEchq6OdR6Wwt+7v302TGxsqPQ05nliW97WSOzscMOWkAF5Fs3TDkg6in
jYN0VAFOoxfoI8VKUVMvqVfnAQcHXspsbFOV6Hbed7sjXns6zxfExHtwc2IPLQD0
ahgrLfs6JNxikDxxCkJEThLjISujB215fR76EJWeKd8FHzz19zsLF8x2O+e4roKx
jK6pMu/ru2JtV79eo8xHowvCCWUvSj9S62rk/qLiDrjFbVUsgiui+1t9EMJt4H3r
GCm4KwSUaNmFgR2pxr/V4gBVViogagiU03ep2VCalF2ptyZ3csY0qr4Ii2Qzg9bO
fRxpQ9+xJkLXfKI/Lx9PXY5yDYU3RuG/zYgej0Ep80qtEjQCELq8tH21rnk/F6Uf
Idn7ftP+ZM/IdcPi3Nnmq6VSyZAAelvu3KyyYRrVRC+HkzFS1bCh6BaEbScaJaJO
k+SRp/r8IUhmURGUmlKznFCQXN7F7Z6RVKJeqBARHnXllY2KMy5SrSQ+Lz+B1f4W
KVevryNkCjK/sOfh9m6PtmUWEUhpbX9uMpiL0MnAZIVqoww4Fu1KjyDuFYmOFz5J
HHX66zyjoAJFpiKwjH5zZTfQG7UFPRAdb6PJ7H5wX1azRfWWio4aWhrx48RnwhCe
r7X62L2C+Ehqtq647YGDrYdm+DqZozf7zTl2OP8cQCCcM/jW9XkuL9j/Uo+Npl3S
bFZipbVycitbS1zidzDNSdiEr0kI7dtSLM7LZMIPrIzmNaXfC+Iset64UkVxeQ+E
o8AIPZVHgIW2e+L9TBDj5ZQbZZTEpRgtq4l/nsUP1A3Guu6UjPe1I7QBljPwGWM+
fg3jTVIy+La422qwayZGC/rRq79S+d8IaZq55AiWdleFO1Tyk5NSsoktG8ixaORb
al5tQ5NmCDaE7ZuLTv9QcghlDZ2VF37bvLbuDjq/LdOIfU8uB0TUNcaDLRwrkT5t
mOxFOKMAbips1QWHR6t+nlHJWHDa78pFSRd3StJV85TwqUSDM+Dc66P/bxjvv1tP
0642R+M52UUbBi1fIQxeOnpK/IAlaoY9IM86tehX3QRZIKKpS1jzBdmUu3ch2uQN
RRnbtHukcn4OPqNTcsMp0TttHfkwLnIpjU9MNoP6KTRgQFSiFz/oNDcXNkGlrYNh
raUyBmEzHUIZiRA7by46uMDN++tB/PLCsSPTzeyswfJ/ku+mQRtJ2fp0ZxrbQEhD
4iwwHRB4wxheyWfS3nH1gn7ZkG9R4wZo8+DKLwKyur8KX6UdfGqYySH6d91FDJhF
riaQUBYURDztVcPZ6AKdlRsbL51jPHw2o2c33nIewa8p1zbBnNEoHWMpvFWVyDj9
K7Apy1OcSvhI1Aoch51W7pcm6aBPCdqhVT8mLvO7cT8te9rmjxAX5HZgrUhCwwkC
/m3+zDJ30LcI8xgcBe9XY87TmfTxfwZ7xM7P7WF3HO0B1rCjTLktGVrM0KRLNPL9
yKzRsnhOuhiD4UKviw/aIfTZRYKYWjyOrRO7Dzyl1vTGdPtMVPLr02AxUtB9RCWD
Ymx9uJe0N+2qgASWY4SM4jJZrrOJOGOBLarpWndkK51qS/VPnF0ZHR0GwYwaHF2b
m9sLIxhyCweErCtQ/E+kS5wFbUCDtD+aQF0i0pF7HakPUOe1GRJ5CMvpDpyfsPR7
akAtWDC6ClKbUbPsafNKb+kVe3WfiqABGuUZ7t21lr4Dwh5D1GSQmW2ZqenOlQd+
7t98og85BFtNCaNYdPJ2XYiszqA+QLvb4ctJDBZ3g3mZMOT6t6iyILoefDr6s/fF
Z4ChT3m0G1AkRT9ZgabKrzVpAURq60qWqo5G5Nan0/8nPQSpMlq2219srCEJuvTr
9oyjCAMYEoKFfo6M4pfreRvK2Ou8Rw5EtO9sIt0HxV6YTKt5iqpVrkT6MfrZcCpe
nfqWeRdkUYbwdWNjKdU7x7WUujNc7rlukFyAA9+JbeR/IUSjvLA2UpeU35BboWMH
U3ogOYhj8CekpTkc++M5Iu56HvkQf4KP6cBk2LAXe/ylNNrL1tahnvKXyTcl1tHg
BHvQUtKZmDtOfLCpfRTkQSzRiI7zZxr5g61vKKfZ03zOoqlpR3PQoglGVlOXwKe3
2FnsI3SwNGrJxkzXbw3sZprH4UxSjVMwPbl45kjDf4SHZBPX96Bl+wBGHd48lDUM
hArCVUBdcVmbaONija3pudQHDvbD2vixnB/wFa6AT95WtmrrkPc67HXGH59QVmGX
5wpgP+inJQaEV/8WowOKLQPrSWdiRqbPts3aQKNHp0kFevI1n3EgcUNI7iFeUmn9
Jez1mbotfW/yoCgU3LXZQQB7W+JQZCWkjNdMIQp7qfuxSyBCUULDWAJaA3TQXlff
e45G6k5gZtJ/PZbQIwFZBtkJbjo4dS+UkfAqwfMTt4OItFxufo1xdQXFXtBq6jjo
BQTnlXmdPvPmKdAI336WnbehZBtkHGoceI40xxKxVCxSYjX8afHv7Qy2R41rASK4
fYdH98qBn3RbN2Ar8gW/2E7xHMuZtz2aOf7snOlpHNkV5iwo++nhXo54uSjgd5g/
GD9HiI0KNIbSLrYmMrWVlwtwKqOljKdiwKuODzxhRt7SjxUsP4HF+u798NlkwI8n
Mtzc6GyQDWaDdzAojrhm26anuB/g3sEAoD2tJonIK1O+e+WqIc+lCUlWRCawIgXr
vOVEYT4ql2E7M9gJKhPuMQnbCSdT0EZwLBsibmu3UrnA5U3/EGFfGGqQ9fN+lT6c
k7CGtZqr+UMw7cxwzydfp65YLHBGdslglrm/yojzd5SvTL5qGUA7p4+C3FUb8RD8
AFZWAgUgUQCAGeA70xA2s21r+8HL3tzUsgDL2r25V4krd3hrAUyk/ROFG50LhIuH
uFOWlMHTolVJq+QWKzopdeT4o64zfdXPBou3B6+wGJtblJshFCOr3uj2sJOmygdD
3ovAqpCUK67JUbu6iPOrGGaIUWIlRLsUdNHq6QIwAIvxRAGtdFJjFs1MggNNsHnq
hfcXX03sZc14bb5blH5M9NTg+bBG6Z+Fwy1guAjdW5zx4RTdSo+QJE2y85bXC0lV
BkbQ/IbUk/swORxQSoj7vvRYBpDZgKc3JJUqxTk8rK2nVmB7MvvMKKebXHzUUr+m
vVuWGhO3QEPudOFQXiVL9CBJK9xuQHmrSFOzhTXiKfZSlfXf/PgY8+nDAebvveXD
WhaZ9F1LnRMEDGiTRRUQitTC7x25+p5JuEYlW9m4WmydLP2F5mG9KzqzUj/rIC0N
AU3kKBz+yzItHjkdL0/55ZHjmvDD/+Xx8L9h7sybMnxNll1F+Ng0oztaDXKmVL+q
V1aeDqKHfakLGs4g8uAvb4HRWO0WyTUgLuP4CNBMGkTWVD6JgkSofp3vMQlLmkLN
AhJm0tVEwkEVMNlWfqDcnbwF9sVi/n9ezEPZ+ZEFfzkaJ4QqNWDcYA627LpoznFp
sg9yS6LzwnYNfgk/XLm/ahdq7p9pR9taPjdoABoh6sFVZWP3dY2JXvZZmBV97hR2
L98dfKC2JjNyRkd1jLXLWCwdvzT6fv4n3xsBB9XsA4cqKfcaCiAVa3BTQz50kFtx
tzCSPGZto1hXZcMdabBlxpsPbHy9xcd5NBZgdQ/4ZlQyG8g/7Rk4he/B3+avIuxI
lbj4fKU5Tt6mkeB5KA836+lqNWpfyt7Q5qrTX5H7i2j0Wjk+bAEI1hrofSD7g/4Q
2LMaVgeQDuUcuMvaByDBF4mCFmKKUoPSCfzaNP9O2T5L5FjkfxzpWx5yIC7NMQU8
bX04Km0xMbKc5/TSxmXzol0T1IvwOdQM+0rj0+2bkfHXqlD3srtOzbQw5quagmKL
XVxpA04uecOpfCSNoVaMyrNJEsYbOkN2BY8k0Lh/kYOb3uxrn4zidWllA44SesDP
MwK37Yw9zFQHO9WwPfTbdTl6bE20sQNJ+H+GAHAaFQ57Ynb46KwQaz+Bsdm8evn6
isODYQpV1DjRU1oL1ocDScfqToyU5N8klAfTQL+8IG43MOxl+gytl53sPi5HfuAq
NiRFYSvHmXnCbGTS/6z+W05ZRDBzZX8XY/CaUWOP6aCYbfy/7y3MRjjXPX3HMSB3
AbCAElCYvXLWok9BLca7bMY5NBWY1QXfe+eNKnT2Io4wmUP0WxOz6djdsi3XqJyn
vmBk/2uWbuhOjGBQPVwtd8nxC8Zj+l+Fe62VFwqQqPXnjzQzN4hCKL72rfDj86ea
fpgGvi9FIHzygVSW7qP/+R9/3GCuJw8MQKAwgEI3hE1uwY7afxovdNewiDBDXyVy
cEc1SADZ66D6Q5gmGVJ3nj4VI8ULiV+kVpoRFeVfYLrqmN17tq9Ec3w0NxCbA9j1
yYhJQ384WouWFS4UqhH+bVF7aNx43U2kqni9Kx2/qFO45svkDDVMS0KVsasJsFdZ
2GTHJOdhSpLeYZc4Yh/ystN3dc46PpGyL1GrUICQNuVL1VTPHiKCPHSgCMvPCjXg
vrYJEZQCK63whYG4i41y5LCT0uZQYBnOi6TiWg1N+HJyZBSV60HZCL1CyJPPsReB
/Xkid7KlD14MVk/FC+GjQ5qlG5O9ixJQpQR9iFVtvYa4x1nJARnYhzgEEEBYB3h8
zpDrIpvR8j9ZhBDWaaMicmEPV0puDzFKzEPdDt6j3vPEBrt9OmfgQZHX5MpHwNcd
1N/OYqlO/VQWyNk7Dfioo+YKHxwpVLNQGw/t9loNbng=
`protect END_PROTECTED
