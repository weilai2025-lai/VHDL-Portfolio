`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oh0gJ4K8lrvxX7aKIvTvjXPyFhTtVL/4h/5EMoHQhYCnyvyH6Q4c9oUru+Ek/0kv
E4br0FoCy1ygQ8nQeSbBkpibdGeD2wlQN3TfmCrAtksXg4Y4f/5HpsRtzH5yHFSV
m5DWf9Hu56NLRoNQvotkBR2McMOLOH92TTqFA75LHAIGMuWp/RN6KsEgCmg9dQ+T
YV7lFJIG0IXXEBCq4Eg0+A==
`protect END_PROTECTED
