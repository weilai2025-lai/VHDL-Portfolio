`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AecrA0dCthe2JYackMsUU52AquMJn05nb4H2yJQPpT1cfMUdJ5p0HfOhgtYDlmuA
QstXAzZl80PpcNQao6Eu6LnZx/+/OBiYw2Y/w5HnLzVSWMWl57sKdF3hFeYoYFxT
1u0UqyRuXxPLRegC/7S+KCjK8cc3+JP+dq+5EIq3flkt8uo8V98GYvDGMw6zfSWk
b0ttWtj7waKekHsJ0mVxAyIUeyZp4vHEiM7T4CAaZv/CWdagisnUKN2AC5GFKpBY
X/CXVbsM+jt8KwH6MfnmOIIwbXwTF7HG1ouVr8mythAXdnJc7lOcenFoYM99zkzR
c7DeZxz/JghxZf1cxizSCiz9OfMairn0Mw/xWjCHsI1dDVgNn9eetpgKU5yvkgzF
IpKWRf51MXbjy1mxyQKl2cMja0RUMy0ZyLYbPxzfVCYhTXomjS6t3WnI0uz4KP3I
G7djkV+ldK+w/Acrz5BDNgu6E59N9gYtHj8bji7kkvyvCWc+bvknw34s2TiC5jKU
PGra9sTJAzdZEyS3qC5aiqaGoarFYw5Gq2KyhCcPqFGblh0KbdtoQv9zt+lz11sH
hkK9BMSNMBs44MfZKTLvn56jxUfq78Fqf0ofkcdincLyZNJWL5BMtEK0735T5AKf
pIiJOYovGKXwwFgYRfelteV8rX0PMG2KcdSumB5m4aU2Niph0gmBt0a+JkJY1vf6
+DENyLkNrD/MCJ+snppd0aIOwmv1NGizJbgEM/FUsmF9ZFq0yw4q5qmv1Q5PxT2U
wCWzodPIQN1wOdUIVtwi5FMapOpWWEBwKYpanEcrn+CyiwU5AFiX0ZXjLqqHjJjq
IEci5Rn7to3utKy0vHPxy2ZNTXNQT6sBWX1IhjE7IvQIdNBCP20S8o3KGzN7OwWF
44kMGyGcYmlTcZ7PptlaPFdME65L+fPBfBDLqKGXOJaj9RVcl56DcsSClQYnmq91
gEGtTbhPuXbzEXZ0tvm89B/5iUoSrtrgb7VAJ4nPH+s2yWi6KZhIx+oDAC7Rwnbo
zgzhfk+pbEUIwdj4M5OZGOWoIo1PPLedCx74xmHk9sfROBacF5QijtN+uGby8OEV
p+BfnzkIJvZguK4MyZd/NAsEteY4tq3McnmR2aHDWJE76Oa4IMYefRebLBJRW1vR
xYRhl5yv9t4EXsYU8X+Vxoipv465CZPBF0r2uQPkyJbmhQp44Jnm89H/opnbBTk8
CuT4zX5bqd6ovr5GXdJbK6kgySzCJZRYocTvub9yoMWY2P4prYhn846lYQxj2odY
rB1Smqrg8lwhUHHE4wWJinAgcPynByklPNn4WJr+w9iKfsKG0HauU0zsVVyzrBoK
00T3fhVwQnkUgMDo+VQg9R9LPsgAb9rRyuublN4gd1E8JI/k7oZLPNzsSEZOI3Tx
Knsvg5ik2/qkxPPwkfr5dhUvUarKErUXP9x4PRsiUfgBsCVY9lomeakcf582xNdA
FdGrjDR4vfP+1WFZX8a1XMFtRTIa44gwpuJUMuvtSHaYMUbyP+PlnZEqFeFAwDCL
3TpfsyMTjDjq44VoO4trJlmDeyYB7cu4tr3zpkv7ZsxhCg8QiJxWOAP5F3VWSrOQ
RsKmPe5e1WoQGiwPezSvBF3YkAixQdRJv3zuDZIrXrsnfFYQrVNzyE+sY26WHy2i
6sjqG1u2tPN8j3LWWgkU9WB0zdNJRpV/YaDbhXbtlshed9Ph0KR0jDp1ax2qn5lm
NRvVgC7vh6+pQvpAj9CbiX6lag5DGDqyGvgdgWBUL5D59yMMCAKF8aoCHCX4XwKx
WTSwhLgQp9qP+/7pOrP2uoHlCNRx31PmOEpUo0sshQutM8UeV7TZWGgxwPfX/fnX
KhjnixtMumShhj83bX5782PovzWNuGhJw5RCQEN7nWJeitwOTunsL7t7C/terzsP
dKWCRclGhxv5iZFtIQNtU+jbTAssPrcr4YSFGXW32hGY7BaaVU1Zp/bMf8REtsgR
HjtUwLgO7CImDj9ZLK8NdyaU94sNZMD2kfXfW91AvHMOpPNfUr3gd+fbaSBsGVwN
iGh7xG18cm7AitPiUP6uPuSIob5Odf7xvoUnhSiUWGeko/V6aMPYrcL0SujBy5UU
XFlVxydOu5jYNtGxAD6pIlB60pwxn86ZsyuhEbOojenSQZPM+ac4E5LSHXEMz54o
TTCAeBOFOtX/N3ObzpvFOiZVCTlfqRjeVkEGlwq8po8ERVNAoIfvmRXLBwkT1VKu
QtTljamXS/aDXMGIa+5juTqmCrVrEyFQQFAnsrJW41XfdqNzHGnz5e4dD45vlxEM
1vog6df8K3PAxVBt8jhe3Lv3dyWI7dzttW4tNIiIDAj5TE7V+58F6Mopda0uDfak
WhcOrxwSFkPvySrWHBkrwVFBbnS2Fspp6bWWjc22m39VNOwMg3gM43e65U32qC9y
b3tIrmeqhazTojb6xUFrw14zabnsiwSBY99aVhk/3bMOtslBgiTXZObN2i8ozQP2
13mYY5Fe//sOHRddypqRx8prdY3fMVptCDbdomz2UY6Sl4Zvw8+qY2tr+8+CX+z3
07zM3+PwKj9NgqBUCA8qOq4xttWociolTmbC6tqEgyfgsJa8hCf1LVcdGSHJMHDe
5aqLz0Xw4ojQk+PNSSFzkQMuqn1afTF+f3391r5jKpHR8kNXV9Udl/PU4NlIJqL0
fZgaHmtplnqCB9strFDybqZLSJLElfiiSoN6UdT+ki6Pym0EVlHSLyNMoyelk2M/
J23oHrD8vPh0uAWWeOr7eIaLPum6feSKX84lEOSdsCJ7OOoxOUsS/OoM1Q3v66z1
Tv1lZaugVsfqtpbpaUQ51lNYjKvbCaCfZxxXuJvt/gozChqIaJXhDxUxy5AkC8dI
QRMqT9K1fmIrnNRVae8xUKdEN6jzAxqQ1mjIgLxffGfZgXWAOGHDN+jaDbyJMiJI
F/zPEHm0ZrXx4htl2asNQzm/SOOtVZRDnZWUIyX2hxufsssa6nk6e44pMufjsYRR
v71jxDqSATGbJca9h9OfS3U4qQv4doIjfNmyNH8UifzATyaUshzfK46KIGj7M+Wq
erVBTGTpr0uYIuiH8qSGp3n8pYxMBCeGiMR79py8rFhPwt+tgNBc99QxtZKqblGN
lvWrkQuAGyyFRPI/8WKCrIvACjV6fSfq25/67nP39y2zVZHw9C3kuf8oqNE3mLp6
JNpP7pVrFHpjDgKz58PW0Jq2CJsRUczMrx8iYO6d17MA/6c3UG3pMh6+JhLrgS1J
ndgN8vX4ExbyLn+7d1gAvH9jdHWZrTpxBy9clhxlQmeLvq+sJauPWNFJZYTg3TXD
jnwgB8VQwFjSxg8aPQdgPIOkdsLqEsSv/Y4SzPGr4wcT/BKQm3cKzLyKx2L+IJTp
yhPpYYF/ebHU7nzayiN8WRdO/kLb7awR4d5LS+Zlmu+HchG6lbKrU15+DIUGvjTl
3gKMreH7JPfh7p4+TA2LiqBHfwzJakZbGrYWvS4oBj0KLpAlLiegrYnrgIjU8pBZ
TBaESaSGrcw418agbEdqzi80UUVgsUR+8jkHzPbAhLYVCU+wr+VOYVVu70mUNQc1
g4q0R3OtLhFt2wpVAmvYWkaL1kda3rJVIEYJZ8UoLf1wAuSHFdOMJYa2A/HM6To6
fmHIbJJ7khNhxUbGbxTt08qngXJZZZhjd9AgaNaoE6vgS0OHu1BMUwIW/3tXh+vP
/NJqsvR+xpOeGKKCpdeI3GBff1NJ3kNdh3owJq19Rv8OPmD/JQ0bjVempMUfiJqd
f/IVRtNDDE0Y8iy2zVYUTtFRqzbmhRH5ajV7DfFjmW4sJhibeJBmPdi6F79N69dn
gCN/oOD2Nbwj7NravsIfsHEFlX1z1DhMvPv3lPsxmG0VdRCWjhXV7hEd4MfK3p5V
/1u0zOGS2kYdbvBpPbUxPlCayTwxNNa8KQecqbSDKl7ame2Zj4KO64L2gLCHbv6S
I356ORDeE0T5myBRgKhdigIuRffg5Lxr5qS1AI7uXb0XrcSpu7+u8VMxF8dO4ATj
qqmouXFlSj0G7GY7bnGKVLkYXeuUqYq1FZZ+46qbdhjm57h58NQgSjFWGL3f8O5w
EWxAFdYGKIc43u9VJSnpFuqElhYGDYwIeXyUrR4/BIXsDpxDKDqPGAGyGAvvcwOI
d8SMTPpEKNoQkgD/wDpWvXdwTM0TtY5anibRkmk1G7gILYl5x7E5bbvTo+dEfNnX
RgH1hr2PChhwp2QisEcZp5ji7u4zbVF1W0Uy4vXR9IilbMygJpLJtQRMCP4KAzbM
r8VQJjz4KgRULwTRsqUn6cgwtRMQTgeR98QoRFJuvlelMBRUQ8rO8KGV55NBwxol
tLsjbmkv07BPVoQfmw1G9UYRN/BUtuNSEuWHUjUbrAq/p0kcsgsxBoHNOQIVSLx1
ZsuFMD9wAwm6RzOElZoCjMc72xHbkTPETZ2YCirvC4PXIz8yxG03318XtvCpbnAM
LmzxYhr9EaGhtTPnF7ec2vT5vtFD/yJJSveB5DwnfJEQvtYeoovNL40yuaVW2qML
vn3CCi47FdHXYY1R9dx1hYwBwjNpd/nl8pkxbvX2TVvE31e4AndDWCogd+o3O3za
JQsRsT4adggiZdYEZSJ1CfLfGIYZHK/BFw/eg6JdgVWVWd5wD3L/COgL/JABCp8Z
5t6zEhJ8VpO7k5CB41Usj7MlAxDqGrcWRXLGSRrYYSjMAOx0rti1tOzRzgpSD0rx
ZXj24bNjTtIGtKY2391UfoFjB5EobkXWEcsDSI6qlggEjBNCQ46GIcUxT6aRTwjb
Ky3oKBLmJFGWKUkLq2kQjIdN1WiNAOcD/lPjTCmC1EfLxGCy1c/V1/eYsEruTR9i
CFiTCnHSAkSfemoWWCwS3YtcUisV1i4WJrUkJUVBmQQbOn2SOQfsMCxP4BiMhVld
wZMglYFhUXFp6WFkB+Y31rJVLvQzaubikBbgLlkUiStDdOkhveiKTvMHX+8emQWt
qUzt9ZJm0XvMc9QTpmK0J0+975WoJRewn7UKMZtQ52QRJ2x2rQbUS/C4piZ2u+Qg
i97Dv/DZuD2Mls3KpDX5d7+KxgfEhI/PzHxoXA29sWC/NvRYhibVibZwK3m1kcvs
1ZR/F40y7hW3dueBdYZ8++KS7pSIDi2sy4DtoWKzQi49rPxMQzBXAfNtQZhac9kd
PrWcQWv5+4fLYTeZFh4ZAM9pVaI2IbnalYsz3vVjCJ5ksrGUGqFKYkcYmfVEZEqM
DYEoaZAmC6Aqy3R793vRybIrag8sq6OIusLv+tCeG+Q85AJb06suTyVLlobMLad3
toqtmtvhg4YNsXFDwqJmDVpw0WwZwDQE8ZR0gzEsLYNj1FW186/87VmiZgwFbNZO
J+Ouku6ptptnbvrEphon49Qzt/8X/pAxig76UvBRx0KC/itQsYv1ovk7bQhkakcR
EEgIqx3A4vfXeJFyCu8l7NDHtDJ1K8OoVAYVhRPURnvJ2UQ0GC89orysGEQ44vcL
RwyH2vuDViR+gZP4rIFyn5dTgLBnLzNsR1yYriUKy6nxYPeVTgGoIWB0b6YHDymH
HMNj+8VdPV7M5w9TWt7tdFKEQhgohTdCXn1ykFV0m5hfT7jezQLHL6vFofY+/d1A
de4qH08A5tMMs0WVIb2jRAhUuHywiBfZvVb98lbDD0Hw3c4S/08HXMCA6Z7Qfa1m
5v0aTJwSWZDxFrG65H/4sIFp6KXRyyANPI1r+Y8w3WnD2/OCaLj1KiLApnI32fZ3
31iaCpdyihkB8E8t3REHiZcBtgywcjtfL1ykC3k/lOwhpkQlz2pPTWFVYlWSzIc+
hvDAyGingVrDOdiQTKAUtFdE+0HM7+pi5n4QZNvlAnlyB9vfbYHZpZORl5UZ14t4
JftRy44cQGMPYoLSPfVw4c2PjRnJ2UE7xGWDt/JoO30cmyR73WO4ei+daU6EO8Jk
P5Cr00TrMWplbto+H0hFVt/xEpt5eTU3RlDBJSFZRXKTUJSNPKhRytGoHmt0Sjcc
rL0DHoVmtBrSTEl4vepnmkztLS9blagdTtf10zWnNjXUXYycrhT85HOgKR2HOowa
FLUjqSIzp2QImfexI3gatq04BU4tuHFQolTTQhvcOnJqO+WqCtmZFQBtFh8UFtiB
vcNp304/Vkx5W50SXjzcCAERP2mkeahDMbdAWYJGQ6wZ+BdYH6FPHyeqNDTBCF56
GZWQy/+5Iz293LXiJnLwP9agIuMFfioZE4KGYKelovNFu/cpF05bA8H9kuAenqCW
sJHy05DuwvYrGxz6KBq2muvjbYnTDEqwJhIR7Drn6TJw0Fhf+TbMTU17Fom2zL7y
ny4HWvOlUCNtgJxCirw6UVslFGvEZYWdOkuNSkSUEA1lsv87NV9soWOxJPTUYEC2
1grDCN7aLuRb5zSqPiaG8EEhu9k9lVG5hSlu/47vExhgZCEkYIq/d83Psj780NUJ
APqv9G0ude87FQntw2kN07GQ8vhFNhv5IYG9TRWKszmOVCS82+wKCq2Xf+SauX+/
3Q2558LMQ6F1Hn/oRgzFNkmUQ2vjb1oOWDTHK+slMIBf/vql7389x/H0cPO+3PeJ
ljKlM8MQu0WD2vX0TuQ/Pab8sQoh7XQ+er11Np+vfGHSoTTHD6Rf4ElCrRP+XLMc
8YLxw6tF/+gEMRHt1DYQaDsJhKlxmP6jFECWdFuYFJF/uK0S59EEt7UmVgPyMqmo
239Asj2S9gAWGM628VWGx2LzVA2cJfomC8xBuz4XcalucSTIebFGeoiTCEdVWav8
GyO7el7qTAhQeZ02kcnzUTwwwVvk8fmS4YG3A9L1ODQUYKerddOaillI38uC4jFJ
sqxhSNCNeZFjnQrwFemhNDT8hbOtnE/0HJqfAIaPRGMrQlE+SY2Jjsnk27zcNP/Y
nC+SQVh3RX5vUcL/kSiDq28gY4R8wYeeDDFCff1m7VKBYbmnFuIiglyK+CeB8QCT
KcwdQHIcsyjP3aX/Y4ij9s7nYGqsyEfF0xk2fFPJiVghSJAjLyhZjkabDksvNBxu
ldOq9+a7YzaYri327Y+EWV6vWAjbULYEFsxkHJrft2rWtZHrAhPeCocdkfSCNPPl
nvf/gD6HPFT2W/QbubZpC/MviYHahzUvKC7gWqdvXOTZL51YA8cGWY/qdAfln+xe
OFPfd8btBKJ/sImlgdX7A1wAOOOf6nzvAQyk1VipNRGzADFcTqOc5ZYiu221LUtb
eZn+HGMg/I3CZnQKY7SxMfBZHEdRUi3JFUgVBWlxIWBWf9A0YcK2y+xACBvzuEYS
Ss2fF8qEUXKSvWvaLhRWfFexZDVUxwjF/m4YCyRuWlXrv7qrpjRFRfGA8PgacNl/
XNja9Ii0uMhj7CM1RQjfz9vr8TGeE47Q78FjZ1gplw54z+ZZ5ytK8Rb0ORfofhj9
5pvzqmLjJngVG4Y7oIAeVqmlDYYl7C1ROgi65biDx4vmz8ejpuAir6CT11ZncVAB
UTIM4lUuj+EiyYUtEkew6fgJ58sR4yopQCcH2eQRriEXZ9esgGpu1+BpO5sNNXqi
bz5qlIFGnXeYyXHmi7IgN85LQ4I9vXbjIhyXfxZhaKELRplt7EE9A5VCCUTF1oiM
RXQYAhDn6JfIi5gE1K0Ha/RML8FtpU5exGhDhPu89R+YMakZDW2OkhAEP4bHKKCP
SNLtpYpTm4g/hw/sgj4ijz/wubVXwS9PtzYSVj54Pf2VQEFRdp40xkGkBXgFlw7g
JBT1J8BQHJDj5RnKnIifL2jPePu+H8o1z6hmkoF2g6NZEAPc+HPVAu/EblAe6HCA
AcU2ss05shbQKLuAqXFBeZ+SdyWXjOqOgK+F3ujFwkKcyhtFcrUqV/cJz85Gya4z
bmSXYu4giw7WwtszbbgipsyRAW+GVh8z71Yyk/sG3CUESMLdBD6akSaxv1GPHWC/
X4KywKo+n/I+DTvWuCS1RMrRoIMO7Yp1wRdtoGxaBqlO8O5ZdS7ulZPeFTr2w/cb
6gF3N6K0dXFNvfSB487cCkHpZFTWtaw9wix6ablBaAjk5Kni3GIdIx88YoUN/pN4
D92c2BLYRIgguBQ08Hc1f4yG/Q8/6Ym2oB97lLllQ484hkY1oMJjkk9nYT1NSEnO
tFXPiwqv7tBDV1C795zdYsHaFUiOsydWZJJHVJ/sfDfCMq+qVqydFFIT5xih4eub
X0RAcheZy1Hi4B5nX4qw4FJzkJshHbizZn6Jtc/Sru38jMlguVpJEhQaqqCXx1tW
RH6CZjjJ68/lMfk7K0WJH2e0iMBfNibdf87dbVbWcz9RWqClxemN0/0pl37HM4MO
Eb19iToLNUKDwK8iWBhVe1UIYESfg4xD5CIR1siy9Z2OWsxg59ZONKPHK1NlNl1V
s85gPDfIJTfqFMRtocPiei9qrhQles90Xcvgg9dsDW3T4teH/Pb0cWCylEz2JIpP
h5O0+ZDWoo1mJn/8jhuy+Iyr6kWmOEcEmhwofZ7cz7YxxlO0jA7k/VidsglP4BXD
Bomv+qChGJMRT61kGJstQwWci8PNq7ut5cakmL+5fGS1ssU91fyR3QKzcUJhElU4
DhZYoSUbYhHkJj31YfOFTlM4QOwv0XroHXtYYz4asH11iXAg4c0/axexEBitxrEI
Jvk25WAwBw9PZlW4JxQxdrwkEF/pZxaVYs46GobGfadOMdzZZC7ifZ+ScMtVwYO3
9NmexQvkNtZZJ4VsObJ1zDUGYxPKzLTTmYwNCtpxpPEY86IKrgqhJ4RyJzSfMHtu
Kv/CQOpfSpY1a0XCHTGOyHLh6svRNGml0cKYCAjc87nnb2NWZ1ELNYhyGfnqTzPM
qLmL16EeN47q40LwKlws4irX5DapxUj/Gq2y1uv3mquyzCMxtB97BvUxJrrf2OAz
VGcC3C+B4UKJ0jHLpSqXU+xTXF87Gs08+yhYheQhq17SPnOaOxH3bqPr389DaYcp
fD+P1iwVAkR+4ul1HGE7bnZQIXrvFn01cRpxxPZ3c7LcgQKgg7FRx816Sh9fKjJs
5gcYAsLElZEjajz9ytBmokBbHQA1djfW9JbCSlAK/NFjbhkZF/QcCaKqyKoLtvP1
n5m+hErOQowXkRkD6v/yT/PYUVsWCEY4X43N8OkYZVL0mX48/xNTviAxvxIth4DG
Izfz+eMPN30PuhWbk2XnStwjghFb40UpxKlNfJMi3DX6lhH8OeDao9vWbV8HuRP5
szq16CxhzU+y98MfzohRDiVj9KPeKD0fOKFOG9uQnGPHpnaYBcXcgtdcSyfGXq4b
eNs01eY6pd63ygd30iOQXJxVCySifdN3nFuPwup22+VkYc1/9sDTVOpkmkDQ53+P
gpQxvunB/U6L24+WxqgL0HyKKAjtQjjBQClG1PNf3PuM3bXkv09uqU772b/x883s
jdvWr1G8uaqUBND+SNGWrq/XJSU76D0alWCI4Zh/UQHo1CushzUrAQa7vm4vOBDF
Hg7VthTW8dOb4OqfDReQUr4odnfnWXRj4zqjv+/mK5RXTTM1CuOG5lINyEFEVjjJ
8p15srBMAGiAab0Vm3I1TWkuc1Ba/TUTxGf4PxhAETr1cEF9GVbBsGBPqkWiuSZq
o7X/HIkBNuG0/CGIPxCgnp7stRhQm0c9qq14L3oYainqMqN6SAYkY5zP9s+Ashlp
x+Uh2Fa8OMy4G9aMbpKrFKYitvQm0UvhOJ1WUUymnLlHHKTR2SihzReK661NMn3n
CxfGLnAbR5XerGRGu/YfOH67dJqMACiVikO7iYV8mpaI5wdnPyI1Axsp+nfCqlT0
XTuqt0ef+p7Dzz7SWJWdIKr3qoVzX3NSGwbMzqQ0T9qkaLW20pPiPtO+N/lxYV/L
qbJViDqaQwidfFcE6ZzquLaw+tr56jLP/kwFUpO6lTSQGDuvSDhnOqhP8cceuK1M
DPBWuAp2xh5t43Y9G2nmdTOQtlnl/7RuTfC+qjPGPm2CgMq7Ox9WfjuRbCAdqvYO
sKaguPhBvO+nsz6gNL6ZtfUFmDiO4nMNVDWSSZtFEu6QPlkdH1Y9HaVRqByhvXN5
6t41nCJG67HkDXop9yihygsPuHEWUP1TZRRba25G05eMU/gQI6eJugfScy0rp/4o
uZMdTurJfxwSdjL6QHpLCPgdFQxmCpxS8cc4+TLDIJQUmQyKzuQw891j713Me9v6
ogaxUyxZz4YsaRPhLFWMdTOKi3gv52SYZ2FeoQX7pafVO5fG8tu20rix0e+ItWc9
oRVh33ds/+oxTmIjX+Znl94UxppI8EStAEe6WAzvIiVByEsKQPOvb1iDR52WVfnW
4P7mMQP/C/I+8NzJ30FJkstr4MMAjoEakpSJDN4AoioaZiFb64WTuIfTuGb6rJQh
RttJQbULqj6lQT7Iy3CrHMUKH5jilZ1h2tEg+zm4XDP7ik34q5WbatjZQOTr/Yjr
Ta6N4JVVBePs5hyo92YYzu3iiOqt2IW1Iiroj9Y5iGNWRZvNnzx0mvCTDk9VcxGB
o+515PU/8rkB5mnt3ZCeLEoMCGUZIUHQzYXBBXIO4DLRlqhmumT7alkl+f7zgAN3
UHfKzABySFq4PAbMThJSZXi/AoVSUzj5L8PezBOpGRXLoFxlFwzcbYUgbon53FO8
bP8xjxc7EGz2UaPgbLdxIqGLVY7zIHSjzj2FHT/uiUGMH7ChO24uvGykAGfufzFA
VyBUOfJOfIU9hpTl2Drx00ODfJt/Mr3p07dNLU2hGN4d/KmSM0mdvOBAbjCHjDyx
R0u8ECg8eebBogQVVefp46cgT97GIIa/Z6MKGFe33PWPo+90UlREBnQanrLFx6FZ
mnO3RzmgZ0QJrJlkqvItyMt4a+jWPrQXARKaUmyUuCcpvY27hUW9kgFCiUKMO4k/
ZHkdXCM74TCFx5PQW/39NhnNxviqj0rNMCE0bfZFLIFwf3Viaxck2zbTksOi+r0Y
pyep0YL3h/uoQPnlyKq+4pC2Wwf7d6nM/5IdATYfCLmKDUF5ZTc5PQ/jhdJxAum3
YudcXR28NtJM0XnufhbJYz6RLtoLRP5qN9kxOw9BE7QZfZ7uz/iy7hgKCZ5l1enm
tBgbvD6s+v6SP2MDsCYsVJT4VOIVaoyAD03Jtimi7xzI8tAA1zjGVj8WX/NmCHh1
IfNGLfWsCHc10D02jneyUkpKR5frwAtKW1ji2pegMwvqaaCsNXcnqXREm56ohLjR
nRsBz80T0veWV3P0sNTrR9STJXJjI21XSdR+EMBc8PaIIhWqAGfuFieCcjf0U4cX
z3EM7ELX3UEIenodeiVxBVzKbLPyxwZG2Up2hZ6P5kpfi6XYdg9WjEhClQ62cb0G
V4wan1axqUr/9nj2gNB2096jJnEM5ENnpvU6iPQHEOuCqcBxqTCUGCq4nRogBvKd
eir/oO0o6aWn9Xh0zxJAli/tg/STnUJ5xNgJ+tJLxLh5B6yNB1h8PqONmY9DKV+v
m7HVSvl8gRu+Fa4PCTufVLxKlUlbtKACYFW7Qw+6A43txXrIEFPTFEAgTKVAAwoc
9tEPeR+t2ZDYwYU5sNaxk/fq+d9UqVw9U75YwImeULFl3Ric2XRrVeaNZ+8Q9sAc
D9uZsPJg+P411YmudekVKhtwWNp0UcF+UcTuA1g9CAP4nsRv9vMhQdGwQpFysko5
4styOw4P+n28AdOyk45N5KjyEwGkNnNNz4vnhfjaVfdF5BU3SuXqmvJW2KoC3Fz6
+otkIrCbYQHshQ3rSyNn6C9UeLcN8vDD/eYs7j2i8J/Nm4x1JqRExeKAB4Ce1Wk2
hpM7qiELB1LZ4e3Esgc7kvJR4aoySEpBLOclScBJ3USGdbYoxq7cS0MS1M50vvql
x2qHesVVB98yqhU4/3uJlxWUh3EaF+oougbpwhVXx1LwihbRadUU4KFIk1Ny5P+/
ncRYLywfhXRsS9NVYxRM+s6q7ND844zDT4ayDs1fm1lkIptSDAS/l81wZ3iOw09L
9ClHMQU+1813kWyQObFM3/QDiMDCsizLYpZPfy2QHIn7FjcSGpv4BtwYDHG5N/bv
N9YMhEE1jhXuGjRciuHZnQ5FwvYYdDqIU+mT/C8GGSq2EhY0bAElY35qe4ILnJKX
SpXC6owG2C8S453GwwkPQAQyP9m1eLVAUMloc7U8wRvAV0EvVMBHeF5SJJ4vSYcE
UEcKxOfGSAQJxUtdhjC/gkDu8p3OXx7Ru4G3Xl7I+iYyHlmZRcoQ4ixuNc9NXBxQ
PypaKCtB06Jdn8s4w/xOD3SOPajY+R96sxAm57EMBjwBQZ9tBZYyQE5L+ICnJzFB
kmjxXBMtY2Zz+iBNqKIT0OboGGR57xLbU1PJqdO65FLoe2sFK/TO9OKGcsb/PsbK
TdIteVyNLJ3dqxKjhKXSRH7Gk20S4Jx2fwtSHJk7lCNSYI7OtiL/c27aWyjbXZTa
XpyxNvOfqVNod6FP4ZKEMMI+nrUrtBgzHXwzROPH3cCBc9nKIwj4vJpNF1k3TmxO
NMfIpdmGN68n0fFPItdErAkgEFqjaQSoOC5lt7JvoO/ue7wXH5NxlzrvwMsqDkev
ca1YtTvzAkZ7JTPZ9jCuR6g9F1YDB9pyJCAFhdUWsthzrb2yL+lnOXRBsf9BCaCL
nEMEKl7ueLg83aUlgIRlojhUFv/AFMVL4vwX0mMGLm8hLKaNeq7eG/mp4bLNTo+t
qpK768PjFGRjBWBgsTQTXRjuwMVXhW/ZXdTQAmRQlu6XyxdBKmoYLtOm9eA5A1NZ
5kLGo8W3PZNVEOuSPlewwd42H+4snUX60YVLdEFDQ9ibS0CG+O97oI3Wy5CMv+xA
CFzEkv3HHY7GYnQ/JfPQw//JvldSW3Ld7vGK+Iqy2dcui8/B2WpMSr9qLrrFgymj
tYffkYXl22bmyOj0yNTyzYcOE3lQj15dI3Ga4q/WWkyGARZZNVpQixYHKn/zsp7D
BAQCCA3kDFICKxLwTLelgoCLk/kqdVtlRQao1V9/pw5YVCaMsH8NcqExll1Fdyjn
f48Zc+u/LoNriYaSiQejnAyvVh0FBmn+x67z+iXdEnAL13zdfg5XYeVrlmIdiOEX
Z+279wce8xvQwZ4jRqavjOxgTo8p1D1few2S205rhasit3jBTnd/gg6Jp6d9DSCZ
7/Kw/kwzvWiPLq6n3g8urbZjiLrdjxcrclkw8nMv4q0Oyx++/aNqOl9wNAzpneIB
0X1LBnCulCeOIH/9VCrswp/fh7C5l9Dsa/IlfS0TJK4l1u5m65XEavQkXeVvZlK/
A7lGFi9py9f6QV0x0dgcc02uYBBoIclWRVHJuJsKPn5c739xhDuXkm/XsiuUQsJu
nvtkSfSEYjvDWDLKp7pQAxTMKTvsJyUPi/gmz7VJZlbsLvH/pR27GSYacutDekIU
hom1rkBFPYiptbhaLJQ4n8hbk9OyZLkEsrhPnVlDQK89s5deMTHxt0o5tB86mlxM
0I+B5HzMbqBESLiiHScy77bF1ADtmvNRP76TB+NIIIenh++VxQHL0OIOjBJmyN3m
LIPOLC7BRgGqFlfhRGAoIoLNL1hhZChwDAVbK2iB9Ku0FbmqKMK2E5NMxIKTiWqa
cToOvgTjsjMcMIEVcjxQDnc2Xia0Nk6DrmpZg9+oSpUsfn/LJ2/P49dW46cetfz+
XQVculpN3b0Xi82pcyUczesisrqmtuTsC9yaQCL43gaTeRUnA0b9hOeefZ3d1zu9
9Uo2wC7/FuwuqxX9dI5SXmepE6CKLbfKC/A5TpdxAdHWvyI61RgNoVBV4UOEzrNm
7jBgB/aXTG/1kEo0XGhbVfoawgvEy8rSDBSy0SwJ6evZqihichxJnPOyPmTl12qX
xp1Hfq79RK4vIpNS8KX1zOdWB/7DEhfqD49DFn4zO3rrriVZDw1FrctwN3gDgMiX
8mccyX8Wysi90hqJJe8bVmygHyIt4eNagkACV4LPMizWFtLblrNMoeuLSwQey6aK
NtP/ZLNGCMOqjMZ/lwLBb6aMoma6STm455TltPUzUeovd3Xhmq4nU/mDYfiQecHp
e9FLPgtKb73HoSaTW3wPRvbIspn1z4gwm/oP4r4EZ0tvXPHOp+lCP+gYWut3BDsa
CP+784kYFWaVBqoPYy/u2pRCp/tT5RM/ckt0m82MkBtRNH49bX1qHxzLZXZekqQm
eO1K4tKEuAUvu6JQnWt5nSvPsEnxvM9Ykc0/WYF3lKoeS3euMONeTsq9fideSDYN
POnRFIFeFzhXm/KG5/sGflQHZV0rfQG0NaiRBr2BCnv4QTkTABCEDn+Bgx0XghjQ
n43a5tt+zRxbDyVQ0i2wMmZ6okdlvvvxVap5i9G0mLrVMA9Z1ZBhzSNpUc2sRzHX
0Mbw2/UiPwkKL7Wt/LM1HZMOlOoV4zt7tdTts82sjr6bkXnE5G1W6irgz0QLtbGv
tKNHOUeYn6hpoe9fuBfO7+TIozfWsL5Bjtmu4q8rZa9j97E5vtKD4sUkfCHUorar
BPcgFgrCXu+se4K/R4YdNS8GLWxzMZUNipa/RnIg0VHDV/w1KWton8H4pfz7sAfu
l+oaa/9vr0dgyGeE4s03+jJdywANHfGeE+Z1tNKH4sbByYlK8qRIkKqp7deeiNrQ
9gsmKvXsrOf5oCXcNO9jwXHcqronwUYOCgjcdG+KHlGUPda6oRBgNiPZwGKmhDUq
bIEY/PrghMUsQs+UkaPLkinbt0SYLgAyfe6pfs1eHoxtvvEG81Xafa2IMFs29Xoh
GMSGG4A1z16Gkx0eSkFwVOgAFsonDsLEdzuOrEnRnP0NPjU/N8/DNjC4kUoJEGE+
GbYHazBv3Yw20DX5ngKa02i7TabpdAmlXEHnBByAz25jxjnVVyFAJc2IRyXRP7qw
v3Mc2GqQAUt/6587c7x+fyyqMNNRtDhSvYhxxhycswvB0EZ4xJLgysh9rECVlAGX
7lghqFXTjkc78k36Eq9beokX/SvF7fYQW2beWIDiqwFf/TjJ4vOZSXfHFc6tpM35
dP9RIeP1bxmaW5YZsv/RAvUOnARG3H8DA1wsAhaS3D/A/jeRa1VCkf3UhMCH2B7E
vkPFdenBVEIgBYGCaeVauDyz2aEpbNn34JeyyYUDw2hpiGvIZz9Y+t4gSyVeHfEl
UOUxxqHvMGkHaOZ8+Q5t9dfzbrBnF3AkD+knfNh/xIs9GmxibJhbBx9XjASWYV77
lVNBSrxWeRV028w6hrJE5fDhhVqVVgMRRGudV84lYW16suJdGJTmPdpeejhLAtmv
2Jz8IhLslFz8JbHuj48XQpeFd87i11Zx8GUPsIwISwk9udd8HHUV7WSFWeQaCk2T
ESy5EGsI9KLivdbtpWO4h/FBCGD1nqTuwqMRdtEb9RdEVSlYfE9P6W+/d1bgIkNU
blQn9RjovMN5Xyl0IZob8P31dDFdqIC27rRYqWFk5wIUhFOZL4h80Xvb/y3mppMp
YzjVR6jhNHloQXg5UgE8vqd2HPQYNyLeBQUUKEm2BGXNSOigUTt4JRJbbCfqSz6a
KNnP1faNtlBFEr+9f4ZT3IsM5LsHvpwmRzkmkASidxb/FeylN0LWIifzCHJ27SQG
1vc5tbJVmNTBxAaMoHWNWw5PVKm9y2uZjgfXNBIZZONrczftVKfE6Kq96QpeFcVK
aYy+eRzhrPdOn8h2qS/BIBtEKVcFYDYsbof3oDlvrhY0AkA1XOs8rOPe0riv43s0
yyNHoQINkxtUBSbgflc92EVmUtCr0fTkBpyUz4pj2Lr20AuxG71/Nvp6Oqe+V/lv
ozouFWEqheg3u7vKk6RPc+QJdtdma4rToftD73YhVhGKP67e1o6JaFbdRkApFDqg
brhX+e5HBBUqselTZWtCjnrzZ9edQ0N0ZLKe6I+gww3yS5jh4PnmA0bs6buOrtZm
e+36dR6o+cDIr9ivxZTDDvivGC1551ousToIPKAiq8PiyH4gqgdcUIsSheV/L8MG
Q8+R5qsuAjiy0e8rsKDmc+ZOf7HZUkoVsY/mPT2csNjLk20/oK+/cH64gQVUy0WM
buRIpxMBCKp0eEUaiwr35Ym8ZcT75k7Fqqp/JK5z0whElpnu57FqYMTb8QtIIWeu
AaB9rWFEHDK0pvkThK2Zh0y6LqLmoPk57OstSDO9dw/dJZtn23h4iuQArMgLi/ut
2et9eX0DVzTW7omtSlvZMegc1eVbbLuKLs2D3bi/gJ2R+WwKgNFGv63prkQnQSQp
dV0CZ9QHEa9vTaAGwGcSw4xS4sKxmwqGcBCGi90FV7AW57ECNeR1IyVuhjTKaznt
zi5TnzRO2MRIBvKeJ6+fAXCfJAxnv32kiTOzekGNHOlGshh0krKHV1Oy3gA+g+Jb
Mxz1zhtAWQU5CAYZ+r6xwtRswuRVf0DUCld41bwAsgD5rhNGR+LxN0Vg4Cq1X8f4
5N2XLlPOQBrW8vUEkt04HQERM8dSqTjHgdYfrLP817hCQgnUzzvMFtyGbizjgdN5
ljJFUGNQfJSO1Wv4+kBm/agUBVhc35RWGGRZgn5npYKLlrJRR2h5WIVNTyheAVDc
x+e5ZmJumjko9g4rHrQ1LshvZLuqHCyk97oLBblu323S2XlyB/tZ9kbHaRLMe1et
TXd2jUvy0+n9qrHux2k2WJ7zCyCYxE3JIPwS//kob+PIaXNtqtjT19wlyy1sDFRc
9L5WY7nwCY8Oj9xpu08d0TPaww1DACpBZ+NGnsmF+TCYmW6jwXqXsQEtZeCWuwfQ
jwxQziXAN7lz0tVfrwuvoQAzQByx9QfMUvDkvxnTPLCECWWQtT2SB9QH9pXqeE9S
/WfxOSFXxp1fGTeAQ66+SSxBdL5JLMynp7UuR1lHzJ0/4Ru102AiICv6qH+fOvU2
1BA8Cq+4yDPhfFy1gSdrG170N1jMVp4QzWcUKKtT48j5h38OP9LLPXQ7oKAsYPEy
iwpX6ZBxutqxLBB/Xh1uWbc+DF54tkz+w53LiXjADw/FEegrD2uQvRrMdW+2cuJ9
puEyn/WmkqKwVJ9Kw4NNiNSKEf+xNs5RU7+UMMzY11YgkehywsWR4hgkFTyXKprf
tP1PDora7ka+q3j+DQiG7zZi8H+0ULtkCIpRKdqS+IyCvNYYhHmWs7s1PoCf7Y98
ubMFd7zuGFxwy4Khfz7ReVYzdDFUyW5hbwtmllyHuq0gNK5xYdTiRXGOS1wyIqbe
jNlYBtLENVihuXJkYMWYGXZZ9NfbxPFSlov4RWyqdLz3TGjU2z5FabRAwHJqzo46
eJ+wcrRsk5M5Zh2SZT6mMzBDax92lWYpuGhMPr2qxWeBawy7GhSGLHZ+3Z1vWSSy
+Pcprz/u2QfgYCrquGx1QOXlOmO0zzRReKIpAh2F5iiEk3rt/0D3iaWyuLGR2Mf3
dTFdJXfBIGv5qoLIwvNpk6IBQKIND61Xp5o+JszVmEVxhx0KNOUKcXihrGPCLl8M
agdJwlibXjeiksh97An3gVFzPnq/HTEBkKNYm0C0NaCIELIZXs8MPkzFfrTBR9UL
/YrorbfCHCYzBy/QCB3Wm4WT6VIHdXmkiOVEc2cz9Jt+iESsC9rwcOs89Duk/8Z0
KN5TnZoUkvQQ5UM1uwrkSjj87e5uCjIXcfLaOdUzOMzmRfuX7xIdin8iNXm+1Pl6
z5i+UfMhg3OhT5VuV0Tn+2G6Qt6qnqgD/r+yVFo3aBOLdl9MtEehvbc5N/m9tu0c
mqhnA6A21k3eANEA0tGiEec5pHi9QAjDCUj+3282cFjBvEICkYqlZkDbQRkpfQGI
SlYlSsKTL1VfM3opZMRj+IaHiNPCGUNu53u7J18J652WC21lrBgLBkJ9kvjsQgXP
zl8hemMkymJmoAUdCNSDvhULfShH3Rf2Brrml3qbpOY6vMrpjI5vlxEBi218Q7WM
JufMfMRFBDoXaoeVFluFFgnTokqxxdZDQxeIOgrew1WT0vtxEBKFDX45h8BrVc+Y
JBcG6SLUvhIc4KnqmEZn7X/lwVlQXNIbtOSerkJ1mKjQKXRYm9vEa85GKxEH4TWg
pm0kSt9x3ob3dMwt+fLbsDI6A9UUICy2Q0ubUJ/eXY4wBtiD2zb8NTWCl2TvkzqI
5KXGtftPeXDi+s1VhckUETrfME4Q4aCnMWJMg5yEA5fwmCMDc+0v1JY4gGYAtrQA
JHnDeKE3rWi2+IW7yfbdHC/GGEYp4lAm+q2hr2SlIYeKBBpvGvi696fmYb7TWkku
KY+XOTrh8ho+oCqPW/yZTtwZu9yvSyirkzmgwRWc0ntP+IkHg1iF8zrf3IpbrWN5
zqRmYHf5pqZnRvZP8CHKkhiuxfV/c+u4lul+BfQjnVR7zTH8tPobnjFLV9L7NSMZ
r8ziZwv0C/k5qfxUo5TogmX4EpkPNYEoDLup/qbCJf/I2BIs7QiC6dokDAAPBqkZ
sQnFD45vkvKgVGnIN3ql/uhpvTD4Jrbu/JOorhm+zusNA6jQhs/J1D3kSRTNChbn
lW3iHnPYc0ecB/WV/92dSNlZ3+zLH3l7palhUQ413IKjRQF47ruHfY7fZgq/ShVy
PTmbxD1fQ69s1iUxhRjVOSILcBnHeHfzznThoK9LeCXBp2JYJ8J1izccvmPB7bKk
fLVnm9siYaF6HoO/NJxFOGMlHdmlmcyftc5xA/Z5iwrL0pmXXqwdeTsXdvRMJU0G
Ufui5wLmDvroqVpfDZBDq1KvHINmOgn1AC/eqKCWmyPoloMie4wVnKPeOOTVZXe1
PYunpJOfHU13q0bsuWvEsUq9YB/Xya7MRh6yWMkXdd0RtjZoE4bsr8MiHhkfIx0/
5whOj3odlA7dZd1FyPhVwudJDFP92B24oRktRH8i9KqMtb2ehgfcB4wZEwElkceq
BP2PrX21Kz/AsbfZdRGf7AiuKdnjj7OzUBiRjzqdS8tkCgXlBD5rHTifHQnxt/sj
L0Gjm9RiltR0Y1wjsBAruMZFNujxlC+KRkmRYE2j0vaxAJnCyXg94FaEk1ulVPyT
XroZ9dETZldB3wi6+u/U/t9bEIYrjH0o5H582+7lV9h+3FeINXD5oiP9udgMJ2SR
/l1Ujm0LGGjMkauqg5A/rWNNWidmHI9yPjzkk1DOc+zeXPxrWgQF4XU0pIsIbVbJ
ftiWhlesDe8DyRInSXu3nC0b9KXP/yxANtVUUSi27ixBpxxozgFO4c9pKIjT+8xc
76BGThTcUKwL9zZxu2rLa+dihj17dkTDx5QCBceGFhM2zVZYuj9pK4SlwDZnKRDf
i5kFF3WBCL/LKB+XV6EHJpn0VKj3HD7HgOYDBkWcWlF6lnX3Sp/R3d4Vcq3ZiAMg
8CUUbzwic9S4dNz7zWHZowYNxhMRyeQ1Lc13bXj9AT8Jg5FQ9lpamTXTbNuzAL6P
Y7tCywSlpDFS9X/gYtaPswgZcdo15rBj5tp+SPdyHLU4y5t/txo1MUim5XVNtb8I
q3buZqOC2hj7MLcqneeK95w2H7JTclyQziBYK1vJ2RYGDvBHs8Z8Zgbqf0RphwH8
y4bpQh0qfZiy+PKS6yVatXhXH3+10ykgsQy6pZ5SL70jOOWV02Pxxi549wFcTV+G
nQVjiinzS4Rive6U0OxnoQp5zuUtvf92cCnyP0St+y/tblyySQejLw9HQPR5hal8
+3Re5Igyih89S5UeGdkhbRrVmCpBF7yZgf9eD7fpY6AoTzHD/RfVhZyh47AcIalA
QYf1D1onMYu46h6bTk8kmfrOSUBBkFUs0cDBLapK3yfOvClaWh4PvPzZcdZfone/
6LnRi5vwiJx62+0ZX1Ydy5KRqOiTuKBjVjus3O4LGK2wzIkBcT8vZtIz4T3frXM1
hvjHw0WDY4VMVPlibOqaS/hAy8xsC28JjaA+9SDhBxUq65G6+5HFdsQhWtBUa2fO
BvC9cw7C2X3QSoB5NOzAeoVOuL13hPQgCaMg23X7BZUUffre+BUwG0t0+TX68tvc
uhtg5Ek61ywr8b/xJ+BHgD5OFkxuZIPRMDnBX7zcOn7HKsdN6eGl+z3inQWDM5E+
USccxcCfK1SmL1dclq81qu57qSvEDcZ1fAZwSIHFoLASjUz3oYZFjrqwvyuchcCb
063wLixX7PRd0nZbYR2dZHeHb7+rySt+TfgNZ4BnHLzZb7NeMXiBLhQfy8LYx+K/
fs9PxJhY8FjCjdqxi82GtNz8t2tcoruiOvB+qaH19RBnFhYtxN7191feFzr1a26c
PDWPSX4oNdgqCDD2zuaQujZR6tb54sQiAlvTulpY/ddvqGTP5uH8zujz383pnnPP
8WnJrJHVPVcJyxBfleimS6bR8P3JiclPXUP+7Z0Xy2fMYRQdwGhK2cGbHWTc3X9k
Lk8HV01+5WLgPyWtYK08QO+XljBfsz4sBofY7rrsiNej0eVZ6v+0vaZ5BRaMl00/
8g5HWS0GppUA9n7FKwXNf3N0bmHMWyd37ydBPL92VAuPJgJSZCouyaXB3m5AZBCm
6kYXI0o8a2kptkkZTKvlwI+7cYnwgCUdb+CgqOATa0aWQhDRxme7mguH2rjcNjt9
joRtMnhYdCglLlb4z9RzDt8fVwz3IYrSPyxG7Wh6wCKa+c2iu8KI5T3tcC1IkRMW
bfyllGP6qj5NJsm+rSWjG+RAtxAcsXAaeC8pk/MSr2E8bh5uwDkEDHoygW4L5j28
4VrMiio/e938qcHBsemdW3KEpe/X1DhqcwL3v221LRWZJ704JKZ+N5ZFK8nMdLEc
MyoE0edgM8JgLg5sjWyZQwj94LcdfqTL2EzogrRgpS7qDin/Cr2zUNUJFjrfbyzL
nXVmtX4rqCdtWI7nbyw9MncO28znDXmsmikSvVz0NK9pQf4Yhz5fn93JIQJisoOq
+ln3SkR1jptgKIV30LSoPDHgrHK6wHcrZ3tAWk+P3vXMVE4I81R/tFQlstv+nvno
g/f61ugwVR15Y+o028P+gEzk7LkC4tA2e27Vg9REl0MOa6MKVr3iQGundCpCPCBd
/9CdBCb/sWYYpiUimLe2g6VuEwF9oQtGcNMWFDZ4etk3NlHeTHPQAbCAodHgFw5N
bvDKxumJYQBN8c7nTs8Z7pw/CnAC+GbqFuTupopFTx0BFEoeZ5WELpr2yZ278YRx
QvYzP4Vxv26USAx9v5MDPLFsEGo6jry1iMZ+k7QKAL0dmrkdtZLMbJLSu5/j82RT
i/kPKsMOG099m8badvQKGIECzeCs0sVZWr9mQTRYLn7mp/4PspCJCuGRhJIjXVz3
St3mTmHDPGInvaWHFHUTXcR+ibq91Y6NIdVqdY4qO7ljqPUDlVQNNNPF6TxvjRbt
gROzowFmP73HH+ocAh07R7fBwnqvZDiXZys5xw3d6qGNtMTFVQPDZ07w0iL6g/4Z
AGWTWzRJTFlb0P7qTVzALn/WWiaXpF5NWDGhO/jjDplB27I2Wzxc0yfmV0BTumXA
y51SfWv/ov5jK7Fxdqi9bx5q3baETONtsL2eztOcGTuUwa5r5cSyji25kiN0m1MD
FtimL8EHICZ7dd2pxA+cHm7Qbwhgs8/9U5IgnG9UhgSa0d1Wiv33q5GywwRpvNf4
/Xb0RkGgC3YiX8Zt3p4gH3EMHHkR1MAIlR0YneKzGaMR+4Hk6b2dtPxIl6FxILxU
jzsA7nx3U+SCE8wmR01mbhMHYNBG8qY1lRqsiwftdJnfVsoiMqM7Yk6Jwr6kTQEA
ipFcoRliy6lmfXrYRu5+BQNPjLFv3Dnae92uRialNWnNfX9PtBHPtB46vGWZ4auZ
OQPcPZ0+Guh6mb4A2Sp/ZYi1+YeTfHovy0rLPwDGj8Ht7ZlW4brS6dhUsMyhkVM6
HW0QnK+NBymgz+rcy3yarvj6CW9Dv/LrorH4EBAh8aJ0QL4HULLF7OFNm7KwhfZE
ixFREpG8MiCSvz0h70VXeL4NdQq6OYIx4jIV5n874PfJ45zxjeGpo6n0GR/YGUfU
7g4A4Dx91nilGDWDFVH8sdQdoGjIpEuqZXkkLCdzr30jMFXEWzWzNFSP0zFhNCBp
tWM31M2vZE/h9vfozTNlQg8I4JJHyizRQI/w+RqKYXaPDdFaIso6NXdiFT7tA9lt
O89JQoZxBRVGYbvKDy5BnH/b/pHLLya2gmPEMWaEOUm4OltHNX0mkFZvfN2p51qA
Eu6gW36LD8tjdM01i5fXbOiIUrRlBzlJo3R1y42yZv6iW3ZwkBAYag4857/M8tO3
MZbN+P3uExIJ6cdh/5aegKxVeE9IswKfUi5T9HIxd+2fAtTSMxrRh4ukwF/6ZCjF
FyySBW7kq1EHBfUhIe46FLBwjQ2IxszSis9PzEJU+GWN258wwLY7FUnq0V123QPA
N3/dG8zZYM1J5jgEMtjFnWUuTBMDTxBU3CfNDps6/+JUVSLGh8qIQcFLmiTJ/yaM
5EZ2SSbN2UM9QBiv0TV7Jyc3HlmUqC3M4f+OTg9gpFqg2J6yWv6fZSK7pCJ+Rzp9
wJaplRoMs+Mn1OMymxnL+CciQ30ar6QCrkcUf8Lj/27+2FPWyMjzKwVyk9qQxW4V
p6moauqb8Vnd9RLUlq1bojEiHa99m8QEAkB8T35jyIdB4FREQPIMGKDONGv/ca7c
djlW6Ra0xZQy1HMcSLTOYZ7QFEcDfOvjieDZerdk56wDMuFyCl3qLdqm4jatLt6N
r1nkgi3ize0B06yyiBokqHSWxgTF1JCbLLGIMADlFT6oY31ZGMqva9II1CrwxTuU
hROS+b+WMrsnZUOoRONzYRJwkZ7FNmh/cvQVQ4DP5ri1rR6+nTEctFYDh42rIdLs
ll33YGxvPZg5lSvRg0HbSAOnwPV7+oex5BKLAqqme1adZHkebQ1I0/eiZ60gu8i5
Qag0mocWfD0mY7V8M1C90YLzNDWzKhDDi9PuNY2mQ/n1uTe9qbM2zzDpuim42Ubm
und1KWyYyFcPBzcWnSTRIBDHN7s8E0QhayPqov90vBMjPrT9LFdnFyPSzlbCjoQW
J/mvHzrjacEVlJk0tJC+al9kCofkkyLSDWNvsk3uEtcNUxQOSh6xIqIWzjiLTIGY
pLqqhjKCUBEM60uNJvhGWokrGJkyTM/+AvDgyM8DfFljQpAnyGy2GZCNE0ZqKUDu
3Qko0LLAfOjgYG6jQ0ZBDVwmXzfw8lyxHycjE0wIpzuXQT0sGHjRHveDl5Qm3CZY
hmd2H/J+tzoeT7dfBZ4J7U2dc/hRseDTj3AhU3kaJBYEQsfFyPxrARJbHmtN+MTy
6NWDPahogX2Y1KRmXLK9WeCI5Kf0+T+rFObmSKmDo5JnTxW8zBs+v8onA1sXK2aK
oMXd82kElADunUZSUH4NaVXhaqOUNRSqkInu6Kfcg8jPlGJ3062Q00QOyKgHGXUw
bQ+U0TBonDhVCE06WQmXIXw+QPdAyMV438NjX/XD/iEPN1pT3ApJW3vh7J+cUCrS
MEhUC0vqNExixfHIT9cqVsnPkiY27DlXjURogLUR9MC4Easf3NGs7mbJo1YrdKGp
mQYzPMjyDO0DfB9BR9N1GO/JS08hsRqugF+81ngyqvYU0BqyYx0O9QsaOCTU2XFf
Xg1Dm3OkazZmfMRQq9GXdZ8uQ950of5Ek71Eo8/nZAwO6HSgs6cWIr+Lg4kQZn93
8iRQg6Q8Zlj/EgIzlwYu0xE+qN4+pyvNWlaNZULuxbFgVRwPdoSCjd/XWM9bmBKP
HKyuibgAF5XHTxWjRDtCCEJ1kKJb6U/QaX1dgzMKMfDp7bVLO3+GhaawGU1ut1H+
f48Y+w5A2TIKJoUONb+HHWj0jZrF/qrEFjSpNf6fJ7WyIxrZWO1f6wnon8TtODRl
dBCodARrO03qA+1+GX8QJw/SKoArXU4yxXvTcGRO5DDsGJpikCj9OtWJ956axygk
/0rBBH1IYyJQG5rJHfuXmjJVaaKj5lQU528E82izVs4pijz8/fepKdWRlk5K1E39
LT++MXqUpEzN6YKC4Jr6JlG9Zoz3MLfkb36sLPV0O2Z0ULFvT4x7z61OjDmKu36z
D25XlOYaDB3APkCnEY01qIi4CXcQ+txoXazJvtvnB69Q/999o58PGamLnMxZu/uc
005xUufAAygOGfxUGUs6pYFEnL9akEH8OTs2270XuCPumUfIYh0HT3xdSCWAS6k0
8axhL+C7stMMt5HZ4B3YB/Y2oHI3GBYLKKIvVvQijI9fan4qXD0UBvBcP6hXSYR7
7/5FI0Hy6vlwMjiLwwUdUd4DRNObtKBlRLNeFJK0caNeGYlWYzSrmsmRjPzOb/2a
pkcFo+A/9SUjSyUz2KBP5C7BPB5L7pVLBXbuqfS4iDNLewv+hvfWQgrmjjT5qXLm
cs04Rm8G/K6rbgV7yX/mPvvIgJ6J8a+pcWFL1rHGz/F/Dhmo6n4T5ktmpxrTjSoX
fbJEMdGrxxvTamz6FKegAv1WSsBJ4UVswxYaw3EXntGb/rlF8Hi64cWkPz5Hf2gN
g/ZTRvvj0q+TSCJvJLlACR5rF54J0MR09juv8gHAgy7BCp58E78AQ2ET4hsj4nW1
eI6YRqq4fS/Gll4sf3tl6tuE5L1gxBaUMRwNyHcjb3Gp5Znj82k+j5DzLbRPOSGL
oKNyMuLJciKPeNJOq8/5730cY1CWDGOI0qR9C7MmfV4+/Q+P4DvntMwC1T1Gtg0v
Ew3xHCDCs7IgkbSZY5VitmfnR6vazdZY9nuk90wkryhkVHXKVJUmLJ8jqMq0+yUN
h/RD/mVX5yRKV5nqftw3XmutCeqDNbItHpi7WZQ/YPIt6YMbpv8sygFs6IMCJpT5
Yhgukmd9cmV4rL16qEtNgTCWvQxmzmxKnO0QrqlOjIDqEe0EgOVsm6LGqPxU0YVE
zWhFfsIp6FVkmIHLc/a3//lXrFIm75NJOKM9P/a3XVbU85EX0P1kJoFemDcEd0vX
KbFF9qCuDssC9EP8vx6A/6c4nKeITEUzPUZyXkQqjDKdbTWDq5yVkj0HNGvI/cSd
X/6pnJ0cVSq0kptS/lbudKOS1VhZSNxturJLf7uXp7nVvVmEEDtPMeRsN2iz9o0l
h03SuzZ2Y2QPXeLprSKjWt3vDuQf7fRWTql1D3jEBAImC7PfEzZE+IHF9sBlhN2n
ssJ2Wm9qeYt95DhxTcQWkD2V84XOjQXXJcd53PkayKHf7Uw5lo3aTc9X/sHMAuRB
vwM7C2/f/xtzdlpTwVLTmSqqVKCvQpW7XJgxmvroOQqmqwlQ/6wgUSPsFwbZ0rDp
WiwbSyehO1wR2z2nK/wqNgqoJo56niWxPJJESEfeTAy2mHGodyxCHFuklqgGU5dO
NvlVAuA2rXAn1L0xobvH2skd8ncVI4UJ6KuEkBJCRsEvBNp/JxlvSSsyitWljcsm
sP/Bc9SKqhrON8gWYZRUBfxDngEwDTia43lJnEo7uQkNKUbC0SkMqPRe7Ujw4F5K
kGDEBfOnGcUgr0mYTbELiwZsnRsA4DjgtpTit+o/XJAFGqDQukMOZ0dXUmvI7r1l
HcJN0JQAuIIaph0RumtaBHpz1sA2gP2BRsZDzB1NgIRjAbrIHA3ZuTpR/TjsNZCr
DHnBxStRKSXIRkt4wcOCTsTed1LDWrIN5Zf0eXGsw0ziF1CSCHLcMob6mrfcN6jt
7deD3dJGw1ZvdAn1fdZ1GRiji6NfeBkPAUS627dmJheVl3O7upyS4E88AaXI3jvZ
jAfzgapo9BGECnFuGx4cXG3apQomFnmj82jwrhJo+KQnxoXNE8KlpSB5uL4wKW3d
hKOLSnYDzPH3apRNXtwLqbGGqOUu1PaxgtY0ZIyOsaCxTGuZ6c0pNGgdU10jP7kc
ESafm+T4wbYwZeN3FDjUJEe6qFz1DHi5q3vyc8ueX1MI4OdMUamYp2fJ/AxZCx6c
q2qW7PoujX51XquSxPnjLwMIdXPrNaLQmsLfNa2da4KGB23uwRurnfUkgaJTWkoZ
2At6CuuoLxJs1ZxPLM5NXtVv8b8LXjyIlvh6yRqszykby1unc1ll4q+hqvtjmJhH
xydG50TaFZdtW9KbH+xq6lOkJ/+dy9JWaOx6ViWec0h0a2Un2QwBI0PNRYrcZIZg
A7ZUmbM8k851MGxFKZNjrCxX9eEx809GWeLCVzxDI9ovj2LQrGzjyU2l+jADSa16
rkFQx5uAI7gqVQaJlTF7x4/nDqR78AYwK8ZTDRzb+CvwumbBsOUs2eAegRICrbpM
9yzjOqYOh8YK19FmXYFnzWQOe+nT6WfRcPT9tX05CAIPwMMKjqKC2hC3ejfOf7IZ
K7PEEEANm25aw1LImgFT6HP7pYtCcGGVsqKnkjS/VNx7sYw0jZrVvctJsqx3G63n
IVt/VTFJV5qmEi14gov9oN22R6iTxDz8KdiBEXtR9Yc0+757oR2xw7vdqHQEqhcO
3XMjPPjXzUxHwtq9oc1tZfRdwyYIWXNzxyGJJ1jfa/Is2W5piF9qV22OxkZXEh7W
vOxZfrM6tAnTpI3nq2V4+MY5oyKcKihkC+7TD4vT8rfN62KfZ9s23vxhET3TA7Pa
WbCir6SYiCz2SmKJj9watYuQfv8O5ZPC7TvGdBHxqWyJqoGt/TzmFvFUql5RkKhm
Qo91vg9uNPODOZTzr2u7DAlnFV5+tyWFz6osfP9eLztd8lWSVmaCOQvfLPGurxRk
s80sfaAFCG2XO2fsIZjoMSbCtQ+YvxOE6QU4MKjqilGqVnagUCrsr1ReQkOU2kvf
b02DscTYLfKkjCSxBovRWGErccu88Y98Wx1wBahC5KOoSqlHRtPrbGnW2akRoNeQ
PcMPFlgXN+I91CHqW4c41m8mMb92Wor4YXa/u3xM28fDRE7rKSOWj7MAfjRRmVWz
BcUaP5Onfu1Q95J9DMMHi1I+GdY7+3YuPN1CwVqZTHbuTpQ9XVl2KOlPkSiYn2nw
6zWD2p98MTKf+Ea7BSVujI88UJtqf97cq0MFaw9LJarcTNDMHRzqp/Ppv6/lbNhb
KXjvTc4LklSBxUpSYQ5fVlGBGWREuoyMTlDrWqzJWjSISJJ05cDqGW+1OcrIXeOi
pXvlZ3fs2FFLnnu1C+GHYDjgITmUxPZILUD302Mvzs+cJO9iPqOQBSjxVo41mlXK
B85Y30TfhurOPAThT8SQzdXIwkozZucpFlTxb24r+zei4hJr7rTKUBE+GXJ9M6vc
JF0yjyW4mpCHw1xNtTMGauam980qbXP+gi4WHgHDHwEcE9EXHzyBjQp7XSyuKJIg
6jb230dyIpZeKrKMxCr6K72ZT9NBPFVC4ATywhVtlUAkf5velO9lcNi8T2bVAKB/
d/lREOyAlwrdBf9/lj5kQ6JvEA+Un2m14f8to6FuvE5jhDJBTA96eL5ybo2nVySF
50SkHzSPB1PuT25pir5ygPfxaZYeLXUwV5h0vh6o6n7uKhEM4HY9ThDodsKxuFdy
BMhwvJtEw8fPGtv6HoS8rSLxj/WyPbGQESX1O7/QdTNMVcZqAlRp+emcwfE1cVNm
EiG36R6NXn5ZB2xCcguTs2VafoRgGkjr9Bw5oGE4FgHVGkY5G0tw1Fk8AhtlSRPC
RkgjOUHaAJZqhPyDyg07mIOLqSm+pxHI5CGwVLKMOpc7H/i3GE+FznCM4HHVpeew
Vdnr11pqSWMuCzKHTSa6nbkDhds4N8ByI7JLp3B7PltQ80zObRn7LR4F2XyL+rVC
vLn/NCJ7ywVbmJcVctVkPhXh4eAFhXKM4tug33W2cKgXDi9oiwQt6XHmT7bsfiD0
YhdZsPvGZkNV7IsKSeKHB7tiXsvskIp4HM/ur+7UHj5gJzX1kIddVUhf9tBO6ItH
qMTWmGoaPLIPZde7r8u9aPj5KNpdlNvsfZQpXTpB8LvJ6+NtOEyd7g1LVdJC5Z7Z
PYPocwFkBNJ6s8Pec+rnPCJxoB7HAm+9JcBcV/iRXU+GabQT/CdYMspFCP2QCitX
di90DS4puRedLz2jQhNrzaurOUTw4dAsRGi9w1sALkXfsi7oFlFJaRns18Cj5aS9
MeQ/oK0Cce+ohBqL9cBCgARAKzJQHBcXeZUpVn/GbtvzJ3JDLGuLidzdMnLKbejV
p2s2HFo0dCTPMP/e26WGSMIcb+8pXay2pCTO9c1XdA8U4EY41Jujj+41VQ46EK0Z
KTfVgrZ7cPzQM4v7Hj3ju9Do93eF3k2aEYHtzSBbHI5K+kQTjfjw+zway79tyVT3
raP9GdCDVLtpK7Pmo8VhDMrShQKuXduijpXJJ1rr+YwdShAZHZsiAAVGDlhszDGn
pmu6a1EQMFMKzvBSCHSAPoqkUfzumvQui2h6FTmzXT+6CCCC2xusB6/u9McdOKDl
Q5rr6+9mvrCjXRme3D2Sm0+wDXRUJTLGz1umvgIoT2rfKvfYo7qJzOxwaxlai6jx
Vx2B1aM2SmUM5LNNkYS+P2nf2FtemcLdTfJkHEmTIn/keB4Tb+oGSRE6KW3Yf7IP
xH1ff3F4lovXhA+ySszDixEBvYXm7s/KzFpjmeB+Kg4mkdmag2QUU2/M0JO6prpt
0gRu+K6Jf1WeZ6layFVkEOwMu3byQpBi7M6u1fLm4IdAz7Ynwdf/Z+LtwGyKBw/+
zJQL89NyEGttQ3BDBSQgE5FZNyUvl4ECvjFGaykjqDRj6W3aoP/GRY1lRnzA7Dp8
4yCqBsYK5ULWROEYC9udu4JFS2nMlAvdtZL5IuhvaLfIG88lU5eWVARbHgjR/o5r
LKh0nwnM6GotKdbUWmM9qWlpUHu+ff+eRtoCioeOQ/POX4OoyDi1xceG3HnitgaU
Xc5oIqO3SeiqKLhTMpzWMhOeFlHkCD6NSIt2ERqz9ciEbjQyX41kmRPt3+uYssQ6
0qgljwuMM1+NpnlYo33r2uDow4hN4lEoytqDcK56LYy/S6ZPkExXAUS8AcE1voHL
jKFM2av3M0nro18+sbwG38LYNbDpChOjT9m0YdzGaCjnSGDLf6P6gFhgEY6pgSnS
XHAe9Q3aIU8Ap5NrLEz6FeuX3BNww+2qHUW051ILTR4tXqE5PJyOAVTnTInVAwl3
20/Xd5bbSK1PAlmVW6GU2s1pvOqCOMzWwXpbKmAtDSahdrQw7hDgqPyC+0EF1ADa
5hQWTnun9G8U80Qd1oSxpBuFj7f6e0xdbdVPLZHSXoSluLUU5C66Uzog+D6JydWw
ZrF5B7MMwQzw0Kh36Hz/RLUPINp/gZM/KVW5YUJBp5/WwStNjGSrgJxYOY50ffIK
td5MHsr00uatPUsbTqdC66ssjlT+kmdEEQB6Sw1J077Kc1C9GAO9cN5GA/Mdns1U
yxTwV4qL/Bo2QbOCbNCxJ6tupxRLDvFak2ULR8B7wEC3QlKa17jq6ZNgNVTv3Mqj
VH8ihVEZM5U6Ty9EAC/zjHoFzeIpm2Xsz30t/i84JY5BlyX7HA6N0M4RjKp14ygs
VF4hA1eCedbSMrhaJiNdtrarnu9B2pZv6GlXz5TmqI9R6mAyk5GEQgrar3uunXVt
MTc6Bcwn2ETyVi5B/YhtAX++nD720d9d/LdO7AS0BIeSP3jm6IDU9AI0596JPl7X
25VYyii3h8qcxWuZfwY0Kt9C6bTeHW6soeDYcm3757fdG2UcMAJPycRXm/B+UcUZ
0hb9ovEHgKLyqINiVrtMHho/7RMoaH8pWhkoWd/pkv1fZ+a5glC7CzvPEHXRcNsX
AHgFaiQ45ZxUEsj3rxR6kGrwXXZYRvyMaytHsnyz57gK7+kQ1mAXInZPMWUEf1uk
jWujJgTuA3b9j9bBbuA7B8glR0AsImGB3JuogSOVgkwfj8CSn65iWNrZL8kGVzvn
XCKZQBgMbp7AZ5smmn4xPvnobcf+HM8HXKpS46DY42ApU1ea6DUFCg0sP74qeWWa
9FpmnY9gbSSFoJDRMv/9CxlagaOLM4/LFGv6W5GQ2VFpzH0MoRAyzLs2h5LpyI3D
UPJfDGT1+lVjz3W3YgjgtjqqyI684aHB4qhCv9+ArpetBpsxhyKt03Df+Ri9ywZz
na+QiTn6Fa51C+a8kc0EWqeFigxIcVEMCkw9TJH2LRQPslEf1lVkcmnmcLltAIhc
RvxMuivw30LehIevb3OiFiREftCxTlq0C4ezXPXZ1284cENgbX36SeWwSjAPX4zJ
/152fha2RcPLHnUf2FEF8lI7Ckd3l14n8iNPAq1Dayjh5mK00w+K4BeWn+0Usj7t
HEOVebx1gp9EqXRDCuHAvKxEihMZ0eg8YbmNxAfXvO0CQqpKoY+vkU2Q0nPeVZLb
RYg9bIKA6BGyPwpNEavQBD8gO6n3A8T/zd7/TFfd3Zte62VoaqbcWN8otM0Mh/Fo
0guRJlzAWy+ht5Dkl7Smn1GwCP6z+QyZgO/S7JtAmv5q6QL1iXUekkklWnGPT7D7
l8GE4D/xBSLKbzPdmafsf1IOAIh2x/t2ErmT427GgoRSfjK0QJObdtBucKswN7pO
XhDYqRsGyjWFphcEre/xYPRHV0WIxo/q1MFuxkYaPrrJio6hAdTONcEYuBB9qn+0
LcefXZWvyXgjcuNtK/Y9sUKlxbY3o5Q1aCIVs30Od7VtSJ5qBQrjfpawLXHiaolB
/ZFAVpuHkbMdanuAXJwi3AucTNSYAIwvf5P5ioGjjYUFVwiwFxEv8MmBVFULD7mL
0gHsYwpFvTqda25ntsSriicUh23tkOU2eCNd4XknGOvThzuOasJBnoKK2bPvvucd
5nUYXqMus52OcNOFNRweFVZXtXcrQhmpb0EfmCktuKIQ3TJ3qIG6ZpuHOtVwO40k
DYkaCQNt/9ubvU9fPuOUmSglQ6dgRyaFVlZkSobRWuJo9rZuPp9EvtFosB0dbKt9
+RcraA5qjM369f2GuSsFkTIJI3zwMECIEJnu1k4U39eciO54z/2JTsy2iG3WSF3m
DUwCwwJNn51WS7sPDe5XLtRdMsLc1qeMaeCcMY6nPjqKDwe6g6kRECuZiUMIJ6zd
e4XCV/c3S7NPA8tuQXIbnMXbS7TTcQfv5eOMoTWw5UkSawjBF3MR2dMr+VvagJ3P
D0M0csG0k9Vy1bOVnUg9v1BCOpX83uYGBur41saR3vUjz8dz5HkzZhLSBdeWWTkg
mmVgSUh/XgJVupnpZtwgKVOObxu91SqHGDcCAamffaLZU+4fsEtCV2tDhtDqbhTO
0XkGDoN2+CCETLVDlOAd7SnTIIrHgToK2YXwGePGkdfQQ/jKMLXTT7+5sl5bdNVO
qzppXsaDk/HUwS6OO83uhUei+xaDusr6VPQuZ1H9YW9W7uKji/yy+9QYxOw74j7k
D2a4RDXYIqlcl/VhqREMqDuz6ruwrM03JbuR0tq0AZjrZnckFWoXKQH52A2JEdCF
y+I8OAYSz94wDuTfmaz0uOEYNabRQkHYCS9RkU4IIj+i3aWijgRSz3pxuy8g9APj
OOfpazWBuWzjTfGkOmxo4Yy0qAhiEpqT0nZAZKENimbaseiHoH8WHTiJz2Ez+DG+
uesPmevwa4OPPRPvWOyf159uxQ9NUWU4nDuTG1NEP+80GNG5kugd9HpAzJyCkjDh
KKpQsslSnId7VRwNMPOV7PP7o/wcelwgp+tR1Xn/e+hNtlEjuSSUkE8cX4cNdILZ
8/DUqpe0NIb/Vj3MT51zr/0j2e9iYPpHmYVTyTcVpSKhkWmirEf7I3n0g7ljLrOT
nOUMHLXtQHPbmfZ6zuDp85qfSJmKVhDBjc91qwy5u7OFv8njaMYmzWrvg7T+asls
q4MaZC17xIx8VI8SJAwbIXqWmnpdeAs3podviWUJAtmuUGPKipGzDRHTB288qwC6
Enzyy8mPYmhtXeKM5jQ8ZgKQzhXR819YrIPF4qdetwr/5+hpDC142UwX07OmOpkw
nEb8sGvc7tHJqV82UH5QiQ12ur2MLQyeajS9lmL2H3nhzXzF7Nrbras0UyBCD/MB
46L+crtv4mPyO+tWCBZOoXZiW7gkSYjU+lik1DGTDVyyPWIu3/RQC/jYK3F6EoNf
HSnXjgS2Ohanyus49jJVcFq2xp+8d4ItK+/T7rFsui/eQUE+LWY9fC9MGfwdc5uw
IdR7MoFHB0PJFZj4UVsbP/fcvJWw6zuSTfDoxqfLrAj+aNS9ASFiyP1aRzID1L4m
xaCu6osX5q8LBuvmuiu1WEqAb8Gpn97NXvw96oubQzIVCzC1GqJrvL36gdKVc2vA
bJBhovndbfUJWJgqRMCS7zVCyjv2HTsJfcjf8VfexfcT0MyXFx0FxN3d2x2pdDoM
AygzFTr7/YwQjeubbSfceT0DvuKu9veAIESvM5k10AY9G9W0d93YelpwhPNempAd
DjL0uRHaOGrK+zzWCv2G0w0v24a+8ARDCYnF4R+WJrNZeWgT7auPGdYJRRc+z2TO
Pv2d1FWabQ435s5XFmG4Un6dS1bGxP0dHndWGCqVXyWiP7dVNUTh2LdwrX7tbpXb
1YedRSbkM9AZLs/94MbD0gzn/kWnmg6JhWGvFKecnszDV+vDv5km3kKgPoc84l/j
yhT631NOXaGAFUc9FDOyOJ+8Ilksurq2y4slcE7mWPPW+P/dx0pI9qxXDdTZJ3Mg
Kcn9kRsUnPsvz/NFcdEgG862RJWIjJx9L96XF5YqUw7/bX8QYGKDVHmfFF35M+yp
6FZa7QTWLyEk3fwBvl+ham7eLI/OUF4g5DOmXniwCJQ+el99w3iz8pWgDELtE6/b
4/kEZcUtE/Z+XOVTimWntiEFDjFyjlyzzjwmvYex0HjyXS3S+whK9RSUWtqlPG9c
w4D8nhNXs71dIEKkwIKLhelM1bR9LHxmC38LbRTnXa/NRue1ACEjdguJ2ZiqZgyI
04jV1B43TAXBb8moxPCaa15mldGLKxQpmFFcDNAtxL+CEsq5L1GaZKTvxj3nwcY9
Fxr4vQgozIKCtBtWHy/PebJ9gPs3mMFM8Q0q1rJWazjowjvsXWvUrn0/CTXgYYUQ
c8nYrSSOWsjfA0ZjKtCEanzr8iJ6+NGOxcwBPKULr621D93KBn5O3uhH/w6QYWO7
jMA1a43oTLwvenYd8ScJPBa4C5l7UnA0QbbFISncuJf5x6XCA74ZRBT9B8HxQG1w
ufq9sR7AfvTY0o6uJcBPXZnguGIuAj1WfbsKO1FeUJDfmCvV2Xb/IAizMCEt5iUE
7HGmGAc6dEnbAJso4qYosei9aRoLlIpdlfuyPG4WP2OxEc1DIPx+MoinE3weESRH
X6ocbibGOtzkOyOS8U+2PIhMhED4MWLVp9EIyQHQjg+fC6SDo/P/C7THm865nHZ/
ryfwialzbD7B/C9A2BAbottHbGgo4XchKS/cSE6G0UG4WJssVytNzhHYutDwY8hQ
ASkdZA1/Xx0Tr1jld8/7cY8WqPFbbBCVZVjE3oMYd2oAsHsSstvPE9OAK+/73e3J
qIzZRNxQs2tUNGy4X71Hjq8DRwFC81fL9HiOFCaQpmXQvi9cPKPWASDp5sO4PDTx
uV4uIm7iTZ2M58GPQdO5THdv1ZHwMGrpjKiFpgJMC6oZV8FDVHSdMCTU4OKyDmf9
6Oye2+askqCpYDVC4UTADk/MmZBiZW5YhPvz6KU6vncut54+kgLJ5UfvsSLzDUzm
9uMRa2l2d514qJPPDoHM/YOa00icDEqoqxJh1K+wNEqlONtgzvqXt8Ibr47vgyY8
EMSxB3WeDoy7j3lNannJhNlSSF5MzKReRRpuDCsSfRf90qIh6TRQ6rFhOFu9uOBq
rlp4PEkG+q9iJPZdp3b/0V8A4xGNB579SzzihT6KrVlUkZRQhg0Ol4IecKwyhWME
AcVXrMotHapHI2BU5gSfkS/UWOl1YSVR4oUr+r0QCXBb8GLj9KIqyM2EFb910GCP
oYjO/uQMAdZiyI48WmniRAilR8bj1EsIt7hWeY4mHj/mVcvfyTHvUbj5hvHidIm3
QngBwqKvD7Be0npUD1fehKKE1M32vHP7hHmp1UlMQdNL8K8ob2yx7PvWkLzTqgUt
77HxjZktqr5/di3GI5ftDa/D6WpLUCjuS1g/uOfwhBEcAWT5h3+Th5itSKFCTcrI
xBhXO39JRUdbpWetfIsd36OAK7dqFHlLaI166UkcD0ysohRPmbxNiiibSOFkrJEJ
Z/WxQdwAeylg4WS/hVmnu0xqDSt4YbC384qPzE/oI91aZa7+uWNZQNw/TeNlnvqV
kHnPFJQoaU+VELfuLgNFFfR4DfmyKXX+CFl1HTLEEv95WeS3Ck/kyZ98JOp0HIEL
I1Fn8vYrYbO1J5pZOva+AJa0FtjM3Ne/x1JnY47vcCLaqq/cJvDLjeF9UGmDYU1b
1o/Q8hHS0g1oUn+UtVhTHxCoR6pgina+eDp2mvnPqpAm3cjevsAdrMMbxeHcFmyb
Mg+q/ic/NSwjRQmZ8UJ35rgxxtBdGdvHSKldphi9KwRG75IWpC27zBLLy6HaeCZD
toV4Gzy2W1ZYv7C2KB03GQEZVn7ec/EkP7YH6ljPIiO6MPFx8u7ZEO5i7W/yVriD
vL9z4P/r3/Z3Q1myu2jkM6c0BRKFAKRpPdfFPNqcQtDtzHpDNtW004OJ7kVd1rCL
FeSxeM4/LU2ElD326azR74h0IwzDXl86uSHliKrozHDYnuav/gX7hdLECVqxEY0H
tosexES2w88sCEnsJYYFkSnuRXHLovfIYscfaCYL/H7I/XRT2j6bBLKqm/3jwQk8
qa8mfuJU+HF8IFj9wlb9l84I+LMDoY0SLfLSdvwN0uLTLOuNsGDxGXpMI3pd+dRb
sVAa2+YJHHSiKEz/mhT3TyYZwMB41vmU0blOFM8EjgFiIFmfszehys/Z9xWyNtle
EQbtsH7mA3bU4xebX4Hs5AYdlM2fCtC1XRRoNFul+esQVRr/c49RkfWuzHgnjGPd
pTQgXXrnoc8dUHnQj8nPWbylZ9ytkm3oGpXzy0NyT1kOAWZW9y8Ud6FVxsHWylwa
LEOTI6VVossBLibpVAD5qS2H8NTeYJwtapgFGHiJ1qaBwlYLuj4fFr8nqRdR8DOM
klC4GQ6WKjAEHvZoXQBzdaZDPUlot+K7mScLz8Ws6/GhnagyxDXiDZP3oEjL6x1R
G8nR/RPaJTKhOHCHDEXBq99YobSeo9m9doFiN1Ato1yDe6JxUr1n6eBHr4D+BMET
rk/OkkD9KKUfOJc2rFiot7zwRbVJd/DbmltfYD/i8Ogt4538PjrpkL+ihZfAqu9C
iFkWoEu8/fPbvnlr0ZAGNMVa7v/QbSmpA5GM8waZiJnUE40WbuUA+FyqI4TU1p+6
1vUjBrh2BW6M/YKQepY18fZkxtDSDIAbKDlE0jceHihdJ9I87VsajzbczWxOQBhS
XV+uB1Xw5Klej6JHO6bZJy3yH9L2NhGU/8smbq8TwbHaUgRiW+QWI+in9UELFh0A
xHJCm/rA1pY+ygwCRR+tz49hE5MONZiD3WKtVrTpoeYq4sfQgND2wF5LcKjf5Edl
6w1zdQ+1fUs7P8QrNMSah46DnUpig/UQ2keQKX0Yn0zoXi0d4b2i/rvwYhxnh6Rq
8Ok9VrPNI71IYn9wZhnHRUgE6BRgTul4dwPJXChuOeQ5V0KxrF7lY9dvDyriLztn
dFFTM2as+eKG5g8QO2nj6/ek5VjBZQ22bh2aFocsS5mc2vp+0ORCnDmSXtHYOaTF
3ks0pg3FN9J1RpPml57vrWDGDrBFjaoHIWUPq01nam5RGchyEZM8bwFq3RTps7/k
FCc3ZTGdN+xOWte1MpUPy7vo5MVcc2qPwq6qmveI9xck76fwymaWh9HaaY826tXl
4oEJU0AmRIAvGtIhUaaW7Z+Lbi0IgO+WFsRJoCXRbG3HsfOE3iKxlQSMDTSEqXWq
n0gnj1OKpAZJlff9D0bzkekiUdHi8v1hk/JGeppzYT9aZaGnfc7PFG2WCGDsAsbU
8nthOG9/vGSQg9aGF2ptwrCHnUvWi5p0S7OZzITdTXbjd+e6nJ6v2yoRbyPHSMaN
0+GEoNG+r+ogDnKVcgOFYkJlYZGHeizPHr+kl+OLECxyQXN8IQSkywrbhKaOhTsc
yUedv3kokNytCoQkz8B9H5r+jSar1ams4fTnJRYTVHeNF5IBKXCjMUF6Beblkten
1JdhrsxcilP0AH3cUtGN7UNsW0b82b0ZEq9fKRNzyMfc1Bj6hSl25SpOjSWAC7K1
JoCNx/2aKP1YlvllBSh3uP3KhWXORrXBURZBcsIxRGDivh28hjvRLa7wWUvdgr/C
RHNVEjaBxnaY5quyekwLlXD6VV6VFBZJTrxevO+IWd9S/05awjef3wHHN/T9RGze
7LUhqQ9spn9oapt20RRgLeFNHIHiV3NQiwZM8YykXP6IQfURqMsQ7abUGo7EtFIa
R/GD5gR+f3jAXsXS4xAMgP8sRVOdnwrlfYXeFaIFsBb82hSm5Mg6wgTag0bG54Xk
5dFALwvaZQJ1qKntSbkGTKbTngiMU3aaG6FvBuCg5DsQ5BFU6mpRBOBFXPyPVRDS
I/9vB50UzVifkAY7doYocLgH4PRgaEvaGDQwhLfUmgRL+iwJoMrDTZhCWR7cP+i0
UDD/2Kj0xZ20WeC0nTv+LMhtY98F+A0Csx6VPTRXyeP7r6cWWjWGZI8GQ1I2UuXs
+kmEUtG0uv4IYE2+fHgVs5DWlbpBhjEcQO/IdYJsGfY4TK94OH1pZ2yqpxG82JOZ
R98J5dxgwHFfnf5itrabL4feLhANNLUyMoBGw+o4UUgDNDXDTefkJ9bQ6bqrzrQF
rLcvyZy3DwkRijZ2QE3yywYgNdVewxKryNTSMoCUq5V3V/igiBl1KCHIjRoS/gFw
5FKnpn9HWQbghvYy3MF+bhgG6g7gjiWmv8+RnZhzzlZcvWkk+wcJXWnHqfD8XKia
1LdOgM1ChcY/JV8kmX0kI0L6JRNlUR6W+VdkkYDQY+DatWSdlSynw0b0NmigEhNv
4e3tLJteu+TB8RgF7CRnmzPePuDAB+XW6Wui0VjlJpHds8/+vluc4/OvNug435Vz
gV4nlAs9OTFRfRrl+7LMwxSszzTci0BRD8apxm/PC7osLL0w4zDsuzbT/jbUzQNT
IwU12j/8ek01hu9x6j4oRdTMQfNSziocppwIvGVvA21T5/KBSZRbnRAd4Fbw1d3b
gR0sZjxJVAT9uvdXecrQUjA92HL/jJIClAvyjw9xfBOkhgU6VuZGjtV5y6OAXaFW
0hAGLrYNp14E3dugDamZVcYbow6W9d/ngZsX6faQauPLBM+ZL56DXmfiZFoAJu1F
k/Hqs046qFO1xHEWFwN+JNpPMtyb+SEjbihSzLjsHMwWImO13ryudGUc/wAAMEcm
RTWI8w6c9GherWjZJYN+9r18U27EWyf37vCaTWWnLU3kby+kFZlko1F4aFb6QgtI
KjW3U4G9fEcU4EaKOZTf53/iyTBZDDj6aFgURv/JdAxMJxRq+GwigUMiLTrkVXTs
+E4AS62gmXXrm3Qrnle4m+Wi1bSCdgSNCEde2xzZReiuWgEivKvAcJkKz5PacMOA
BZqZq+F/IsJyK1OSSAoJvqtkdSwEbIOKZ5iuoWpMOpXY1L7otfTEtIXG6UBEq5u1
E9JLXenlIO8u77KUY0TKS8EWCgtEdCHnck32LPObUovYo860uHJ6oLpFLbOGalJm
mE7HGV7k83MS2yVFk7ncOepcNeB5R26VJW7JQCWtxlq6p2L8jKWQDBEWmmwSIO8i
96T1jwYq1MpJfhmCkE/Yr4aRAPYLSoNWS8NDpRJmN/CROo/2W1aJEOl+xwg/VS9B
Kp0AAB58BxlT/jbT85swNdbYW/fw0Vxtdd5BJuBQbluUAGadx6pZHEBOQGm832id
JHrpDOuUH9YL1L3vlIltq+uChWzG+xf6B/eEvBtKPoKf3cwglY7u0dT9BZvnT3jQ
S1K40scEnRMqpglbiTkk02oZ3A5+MXuaHrP4qZzS36jt/9tSvJ+SY5PNAnMAiL2d
NaApuTwQoPun1dCunIMjlXmp9onVEQT6v/bRk/vpRplgcm2bHimtAEh+ty+wDs2R
HvvsBgjSc8cmH/Ab6yAmGoBZJZRBgcx7eXey05W4OFtKuRH7YF7pXXNzPcCdoNq9
D9QBVSAD6/7CqXVPP62Ft4ncDlvb8o2XP5C5hu1eD0sIypShshKECHccEK4CyyWa
SpKlGX1iQCQVKBfzQd91kbrI95CcqlOA+YPl8YEIlyyHQJyrYxXvuTDty0JBcWpa
fnXu689lHtNA9CysQwXQV1mfQ0bMyuIQogia2ERqDuiRULGZ1Hij0OZ9kj2eXSWw
Ieg6v5N0plMOiIY0jqIc4w+yMkLBjVOB73hetmtGn8+tp/NpwOwQh/U4b/q+82X5
gKzbEpgq7a0m1gOYV9fnt21rVY9OwFoGnznerFOf7Fvdg3jEqTY0RL6Aj2ewylCQ
MmHQrhFIy4KYEjdS3Zoo1UKdloSQQmFtZJjamOnQqlfpmH3bnCjOVxSGpKnQNwbJ
tfU80RRJ0xkC7w1szOAfUx4wUph7oRSEcmZXBsk3s04Q/J3Pak8SzAD0L6q9K+gk
CJZv78MtXNYKPUJYeojXI47HaFR9M4Zp5dfeLUXWnxr9MDURGOKfVlN84/Nn0yke
0cvKuLb1KxmMXx4U/jir+YJOJXEZLd8ZB3w/Hkkitzj939z0zmSf2/GvOxKeF4/Y
FrpOkGWYPlqaWvfQrx63JltudjpFqD8i/zBraWQ1376/oO2vsrLYt5Xhcy7MPATU
e+L7eOjnF8Eqc5e1NwGVdTRAKGvj1FarY9MmtLcYFNHqB4N4tmc+iXBLGalp5XcW
tvsUgg/UtzFYJXZV+Ifmwgy+b1WXaRbZ0YrTZFxTZXyvrKBJoVmcwpDZlde3AwDF
fGz7geSEhV1PjgcD9NQ0e0d8HN2tPbsbE/hTtAbwlhhom36AM9rgnpPx1Kh10yiR
baT23g/CeQUgElySv4HwPEQBbL5p7y5Z/bxjvYWvl/gJtmkZJeyGp0I80ReCt2YO
BaxwzMSmz0u9BXAHLTlg6UeVFFAkqb83WKOaDSEodCQKAQEINTLFZYkCmQ7Trnlb
Q0RJJiCVTeFRM9WMlfuY72+yWD/a2O00yYxuKQZDz+2xf39CWNyDJw/3chniLZT3
wGpCfwa3uUIoJbApU3iekR3+mD9s+Ef9ndWc3KjveBGJkEXisZXmB0jMU2QyETwt
QrViynDLoPQYfI8J8glIzimUQau9RfdHeDwDuzQuizoy4o16JQGgp06KHoYbJcLg
nPkTd59h79h+UJSPRsN7w9zIpACmAN+PKyBtRY/V6bG1Kgf8zACDsAZXs7X6mId+
iOFssn2Uq/V9G+30XYtjiuQmb5SpVaWIQsWCZoN7ho5c+ujp4uMOfEoD1i8GYZ3+
kK2mhubXpLoSUSkYL829mcfJM6uWS5jWR/rnbXFmvlMFaAJCil17n7z28HtQ3DFP
XRY+pCf9EzK8xcgEEELOSfmVUgUhrDBUmhZ0xak3/R8b+heNY0Nqg2xwu8vvgubI
+zAb5vjnJRbjLNkZ7O5J6VejCW4CH5S8cSQlYCXQLxa5M3O0eDYeB7ZbwjK0EkG6
CWCmmq/AXrraNuF17TIMHSlLlMNzlX/vHItkoYwcf9TJD3qwKg65jAkCi0LD3hj7
y2aYXlLzxrneVgRb2Mbn6Onw8zzuhLYT61YM9Xdb+uu6Fb628LA32bx2GH6ghvgu
aszOaYkPeqYj+cSR7ByUmwRrQhDYPKXyItynxMeDSndnhmP1icDGqKQnLFjuctrf
e4iyfAyAkJEerPlyUbfP+oVv4CK3eyAimYhoakYZxT+EGH0OOByI6ue//dAVsji3
Myh22m1ef4zOuMvXKj0Ii4cdjJUmQEW7uwYJbMwWuNoBR6EsJxsRdUfI0V354ldm
6aJat/0sklp/V+7Q041vc34ZmXkhajAixZ6YjJ1GiJML0/MCqolRuTJunO9IvIiE
GQFvyvZ5QslXV78N/JFAxzXWbh1m+3Yp1Hc5mV2qQWUlSOyrxWWI+uiw2NoGX8Mb
AgqbakoPxlAyJlpUNAgBpkVGFVk+ugDKd0My9GDYwTsYrvqSYiZkh9wquCmhz2LB
Itvsyw+nnHVC7j1LGdsbHgG+IF9D5yAYbdOyN427CjSGIE5XGxQUY96GGXlcz/On
Qqzsy+eliTZ9flgusnRcERICj0agGO0U9kCZHXdUgAn5EbgTvZhWTAyoIrNGtX2L
f52esndcVSqO1bc3mtl75oXPeomEsKA9sR1q5mXZlR2OdGc+SrrSXkpHzw2Jxfyy
Qnv98nMRCCO//9f4rQxSZSgCaggzu9R2H9K0ItP2tWtdcX+aEGjEOzjofBbXT63f
BMY3Jcpj/KxlXgX7bFkv+KwYD6S/G3jK0GYqb9ioKKi5pyHDaQgIF0GQM23LApTw
R3Y95aV96c6MVQD+ItwMULjPufl3eyJqUjQSpGMk0sZs2cBVfolZTJPuS3yFbr34
BL+r0AFkm4u+wacFnJK29Ed39yv+s+DZZvNHuqs8jAuQl2Zy8mxLHdVzJm2eM9tv
CUbWpCigsNVVmH4/rAvvadkbI0UIkhTo7/K8bJ9bf1ZmGOZM10KtRWfQIuUIefVx
wNNr+FLALmzvbUIUWPESrSJWNm0NQ3Sfve2YULk52fFC8HX8FsKJCDEzFvIkU8Wy
OvG864nYi79RBkJlhUoiSHkO55qTLO1YNUZrf8UdINXqbf594eIpt4P5jFGS+lQm
vBaz7C7Wra84BIlu3X/gdz3cSs6fvUUMy0ILT6jE1Dici9VW3JPdrE6GLvckBXEw
lf843jZwwtT0RuLRCzqvF8U7KHK+qDpBeO6p+PGibxXl+rngKsBtb+Ink4fvnE4B
9fh0Lhy37P5EpAFPfqR9oAUcxKLbuNW3AjBFfDXiGWwzf4NDaYLTYx5ojod57f6y
DwxAL7milt9ydXV0BwxjGwuBLp3rM4ArwUEajHUnVCypS/6Qi4YoTZZF2X76RjtY
A0U62nUhqu91+qfer2Ws7d3IZEpdnCLQT5/KEVFWqsFNqCVy9fEFm8v174jAJ6hW
sldlNMM934GdnACXQZO+ajyBVLZu7Eaks6tlM6Zcqz5oIRL+FPT5IDqDc2DUecxr
ExD2P+FCsRAe/DUNo87jjwjKSzGFm09A6VbZ3AKuryxe7gimxv6LxcAgkikZt8HL
v1H/Bgsige+HlZ9lmdnYpwWqz7gH+4X6Gp4z7joqULkMlRW1Ikf2DZjq4r9I75Hh
/H2F0+n1FJ+EiYE1LjaSU3uqnNiDRbWUjzdTp8F6K5gAL9uDxebmpPqYs2oDVTGW
6C3oa2i7sPOwXMKI04t8ve/6/Sc6s5rqQpJCa5lUYqO0o6kDrUIZz0HabY0MwW54
hSVktgXb8lAfL5qG0GgtNVfK6EeUHcb1UA31lE71OfUBZSBpCtWLsY28/GdkuQiJ
CD9wmWgbHk9xn3LoeBpViS/rhxEif5HmgPA3ycErwCQuMcPmYC6x4O+bGbKlbHAU
WeV5M2oZ6Ilk6tGUrRbBJIcF1zARXv8tHYmVpDAhpOHh+z/bjRgWRaTIK0Pzfwuu
OhGMgAbP4EcfLutvUjCTIof0G2sbD0mCXKJdEDl6ebzZ//hnrIXJ2o9PClZch8lA
P7Zsqv+I/OJ7JTh30kmQYxtV179W9CJZZpBgnrzBXejQV4/ELY0/94wvTD2bJ4NN
Y21a3/TX8wZWwCrv5bkd97iBOoc3VR3E2r+aIIZ+YjnvtezufKNgT25EwcPC2v2l
S3ikQh8s1jLyj4etJmVMwyl26GBwTW6LRRipiBwSFujz9xwzx/gO7C3CRfAP5Dg/
vQ47uA2hx/soeb7Fh2Qvr4pNKkdjGWhx3en1+a5L/3GNdtYrz4UhcnqVjPX6464D
x+rZ/O9T+nxul2kFYr4N+GF0wzETHuSbNXfGJxRdAQRNlY0m9sFuPBWvCEB6ZtbK
0cuTNPvJEkHgyRmVoz1BtKG7kuDaP6LJZ1plnOvsoKSQS5Ku1CYbVTjwu36pqHxu
P8wNWQOyK8PUdZpapLs8UNyBqEAv92iaI3esciMnE4040typsNOLgdHD7VM7LPXB
ANIU5acsaw1icPoPvfTFJwoklBmqYD2dvKzGykPSVh5hyJkl3sBgvbX4R/ifexc5
J6Fb7XxE8pQo8z+jzz4MKIgv4MqAjslrXCaxAnEfTy3biYsHJHGs4OV9u4iwVaTZ
44MlSr4y8DHxDQsU5SEd/iClBwglawxwNd1YR6qwojbR0jUPMbY8m3b+y7/dS2aw
WS0E6uA9KlI/BW5eUWgjF10Pex4w7eakRMHfEimRSTcUrm3P2Jtv+AwcOU+qNTGr
4ly/6a/w7GpBZbIP8E4EfYc34O1fLG/+nbQYpEOho1GlXd6Z8nZWKBVk7r6Yzk9m
obWIGp9ahCCc1C78iz1WJUGFJqAwMSC+D5HZsv/RtRInCOc0KmZ8NKt7rBjexLUg
F/BffFymY2wjxqn1F9d47m8aQpqicBHmg+hG7H9ut8I4tPBU/y9WwiWLKGPLG75W
no6RmMv33lTlAgCGnVTW7NPPFqDGTpi8HRWGx4OVkSr5sMOcMirMeLUFOqcFnKhv
f9YfVfWa19ST9cW4KyP2xVQ9dDJu0+XCwvl/y1Tb0rPYV7nsazviYRVEzWam9xVO
xhAS1Yp86WpfOLeK601pepZYKk1MSxOOOfs9DxFMogItCBCC18DBe28sqVj3yAA5
2Iia+G2oPgWzXu2O+s/YeBn12xjh5wT4e4Tc6MN+6186aV3gJJBjNpavnStSTtM3
gp40F1AWhrTe7X2aMpVjapVgMqB8M0YXnn2dEHhQvE69TfpVgBU3vfeTxapGJY+2
bIw4YJ3EugrKDKglkfdxaGFql9gtsPO/rO68pxJqjbOZpyJzO0Kr+YCvU6SSLsCN
BldJCRvtToxc8uBz8ow3yKP4vsbzk3YhrqLO0t/YCrrA2VdE7X83oG+6pBMA5Fb2
jYoTX7C52AVYq+7sEWQEc05WSZAYwBJxLKjWchIjWjmCTz0tHnGbZgyYDCIgla4D
KBRMGjCmlD7/SsnitAvpiV7Su2TY8HW4pthuyhTd2BG1DWsC3Qv35Xo0nZwnAh+O
pVoeIiv70s7OBInMi2FCdngdF27xOejXSfFGRpXWYRuylwhhinIKc5+B2Z9oF2/u
d/JemtaT9M42DWq5oG0IjMODtJjsySmIoD7rHmQl0t5xRSg5BN+6M2tj5Qa6fjI1
dn2UgkkWCD2tM/AFHfUGRQwXXI40I5Hdcqe4D1SJKyM8KZDOmzXkvlSZt+51udIr
3xM/VAERqTy3T0e9YTc/Duvuh0hicH9Ub+vJWTerZbEGuQBwFYLhhlMWrqwBqEch
v0E3vow1aZK58bVjG9RCZCssD2ugXMdGcqvtvrC0ijzqPNyEl0tyD/HXBeWXxRwP
y3w4ljUOlcqmmFDJCqFBZp5RFMCS4wHsc3kkoUpI5hhROHKJsU5R/tFOuRzgSN1A
o+2+XcEveCsBcB7hivqk/3GEiPS/mybLG/71f7iFrXKo0oxlWFuOVnLY6+jcw6JC
AJBuGzXkgNdEQqOhMVTD4yeeJKqUHrpsZMaztTzMRmWQQWWqpuIMxPJiHFCFQiYy
53e3ZncC/0PCQsF9Atgk8X5T2UPV8GjE814fDpD4BydL3zUe7E28FKBR0FrH6ct1
Xc+DogMGR3JsaxTHOvHxhka/NsUw3LZ785RzvPKodpyLgfZkq7odMDt4wijg/rOG
xlZNTHn/sIE5kb3r++POyUFm8eUOM9p49NO9gXAdw9rPmf9GnqCRC1NBkGj18BMt
gcUUCqCBbx2wDZqBPjZKGlW2XxUrmVb+yrI+8SVjVC/n/VpVyxVia2hglFeAHaK9
vu4SyciBgvseSM/0kmvTWXEahncq8nW4kkF8DhEcGKjhv8OzCCzGnAdSRWlJPgru
lvQHE2OUXM+aM/HBbQ+t0N7nguS6n9ZybZr/P2001cwsySfOoVyRkT591wHVkTfT
XCf6e9tVfdDSyC0tb1DGWa3TtZtAb7vjaRCTvq1CCB2ROlpvFbs3Y7v+QLSaLtoA
zmZmidOJjDhqW8Uo/prLOCY++PvuXxlu6p+1Egbm19EQs3dw3VmEg8D380aq3iHN
jdOjJ0TzfxEZnk/m9mTsXs/Zc9RiV8W5w4DzJfxmjYBti9z0P5vBFSBNJg0IKqJp
x+vVKDwqj1d/cX6DWxVlE7ETT0alk3+4nneNLHbL0ez60Ubos1NAD5+kIRpsc0zi
A67bxFfThm/cBbezxm4x3kG202inoJDDfhxKy3CFSminbBOUMsNBxydrTzDsc+jw
FHQF3uen5hUZrriECWa+lNVjTBmnCIXbjnMndbWorySLnRLNBxpT2p+g6IMVYvfD
JdxG4ybTq5dUJaNUv0KO21wbHimEATEcd5tGLj4iBC80I+SnhM6zbFo1SrP+lDsE
KqD3QZlZuQ+EU1c/IwZUyui64dlS1OM4OuC5dV1Lz1qGV6g9N7zj9R21/adxP0fJ
f7DaSnlK8SGS6iNYpO/97BxLvYQ4eRqzHpAwAZoqwmEkAxmWjmt8PJVWNlyGCkvu
hlK/qNBe2N1+Jr1Sz0bvD9Jmo8oXEJg7IJCAAgslWxctJiEEALQi9r5q6UAmqYMa
G9YtGCCKcQKFi1c5VT85TRCHb7r7hoTKpAKZFkOQXjLNrGQ2o/Hrkb5gnhl1epab
vyGp52VircfqSTkJlKaoj2yBJO7cBEg5to1KPnQr0Vt5H1UPIxSxPUpo2FpfQdK6
7wMSu4Mhuy+oWEk3gBSaoR1QgkUrXybgABIcubCvobzUnl+dFHCCEMIv0eH3Qt3Y
TnAiq22rZPfKslVHBZaaAugYadwT7Ugz+2biPGt7Z0F6ZSKI1FnFBo+ygjzFtIXQ
w4/Wu0pmjrBQ/xt6YK9+zzb+YaMmrGe93503RuSbf5wCAfIx/Fwe7lJ7gGLTCuov
B0Ifbg8z1+cnFY55xEW4+wVG8HXMVfI85ybDYd7g3pG3yzaDbbpIksusUxrZB/Da
8YYkqnQrV6ME/ko2ttF3P01Fgcy02akBxWWjRXL/1y4MlGcft7dTX4l20ztV/EdI
KTTdktHRCOopnBnxhx0ykSXzqCCSpBQ9gQJ+lNJiujxRXqmBC1boStqv+2FwYxX8
xO9jqtu37CHWWA1PZgeIVYAK0RrKqxbMT9zdGzKY8w8eO+ZCgRXx4HX1vR6e6t8r
xvbC4Lzi5fFuPueG3Di+IiBd35+O11R8Fj/QawB8SyDyl9IpuG/PhKAM8daNzotV
n2EoQYAyD2w1OlEhUD6I/DUcP1MOSVApc2TzEB4s93nQkdj9n16s3BnbPrUylNWr
ANmn+WiCk+5kiQQofkeZz0PHPe6F9DmXfYwFN5/8wPn90C5N6fKtq+vfngV/mUvN
gpTyuyjVhJfU6bLj+2d/X9N22w6rvssRkP/fh4aGRxpFv1dvHryEhleQPCi9vjP3
IgXJOBLQcUaijh1RSutStH953K9nt8rbVMl8NeQkLw2FXjUflT6UJ4FrNXWmtZJ8
KjkQZumrt/W0zk/6xVCFARAxp4xiHRArUcdyj6kRkpRAP3/2dQpSjzX0vg5HKCcQ
2EDqTiRIffLmuiDBW3Dynw9JhAn3x9QS96du5X/4en8E2iGUARGyGLxFhA6EZOjn
nXAgoR7TIfvYxJsZVjAeAQo6zODlm+Edkhak+bK/LRSDnDiATzEHbWQ3ANrX+1lc
y1CCNXSuLy+DTWCnJ/CjDqk1Fbz6HMqllPaSL7diryG36HS340069q0L2bSNsqrs
8Y4ZrPatUiqsAHKVZ0esCmqqHyltNO3+E5dPPWe8/KRzQjGGwuKFscOBKIRvmNX9
DcwMV0hi1jDFuqVZ1nqmT9u2n4kmagi1RfOl5320l6fbzCCAMvyviYHooPkgwRUF
aHQ20U2kqvVtt9zvtWmFObom/0RTl4aDg9boHa4FRYsAh2Po8k1QktD2K9Giaji+
fIjjfuRo+OMdgDIpSO9F0Fxlbvnt5n/QQ6kGOkADnHP6XxE1HZ1eXnMw/d0Sjoo0
Fw71KduZeGr0fnUljyTcf2RWoZwKxktmqU101Trx451LuL5Bf5SZ8IDmmbKTfPMK
Fdt59DNx6BILLhmEx/9cQxTn00RcTq5uBSYIGntLLXFKGJrsivw4jVJKYyNa2cAy
qUjKhvKOP/E/lQhhgw+JPnOZekDEMCBcVAOCaXE8XKK7aN0QZGs4L89cuUAzOsKx
7JwNFwo6Yu67ClEmCN5aPP4vUhpeAOtNhSOmyznYaKXtRy1SiUUKhuYa5z8kz1GZ
u6Xjxp7CUbw7tKMUYo3h6YdirpZ3Wn/6WXyQREoQGOyCSl1lf+cydDwNftX/nTbe
bZEABnlxX5DFh80zZB6dQrJUEHAmVSy9o/Ev8JhT4eYG5/quS6twGsB9MWkf6Hk7
rKz+03RMLwIQNApPfudWGVuRML10x8sT7/ta323RNJryel2KPdMjAE8VsaAfnwWd
FYEUtKO8d4vcFnIHjrfu2bSTQ5vj5VZo8lDpCDfiaOVKLULDG5i9KCGTI4wrkqE4
GwYdPhHf7bDZx7gRzRSO6jpziQUGMqgWBsDKszDNmhu0zscKtcVK+HejH4rd5VCG
qnG2/RhExjdBg/n/BE07Z1YnlDvt0+ESAtwlU5JiuvlkN9S/TLbrtsg6zycfl4fv
djAY5Iws0+wh+sEBfq6bG5xAvuOKZApqhWGjBdGZvHH7oncap+YdAGryU/I2544U
o2qLnhtF/oPCX+S9uK9t1PNBuVD2kp4AQto2db+k7zFIgSx4e/SsQGrpHJLpA5sZ
HIEAuEfulegr8epvLCWn1AjaHxjvouMXrCHQ3ArvPhjGxl0heyg+I0A4TEkpEfJp
OxgAUYHtHe/ekQ2BwjN/6RuaTbU6jER6jXxHFdrfAymEa49Vi63/VlYbBgmXLiSS
o1Cfp2YyYKsUMuvSKQPaTIT5w+TVlqbZJTxyBmVVkZt1T0c4FCylGToW22Z7UUHk
7h9Fe80/LU9JqTBLAtYIlR+lJF9NpP8gZxin64bqPdYvVvmFEMd6RlOQVAnHr2yb
6WjDJYy9g/ERjPe8aXgAZBf/kqcUvdajQsXTlLRtBGRHFPSbq3cD8GKWG6WjtJre
6VRGiTPwDa5Jf9dV10JxoZZuzTlJImo8OlPK1/p+EXylNokQ8fOLP+rXrh7gujCR
ty/I9W1MM1taT1MfOJ6JXP1Lx9RnHGLSl6MfzMzJQmy07ZjbpPNDwgpCKe8OK70i
bNinvL+bDNNKj3ZRMAGKYP8cQLUt25Wn4X2+8rIludI5mms+5mK73jYY+b1qZLRh
9M9UotY2fOPBWiv9Bs+9Pz0pLxNrEah7pkSKIz65jKIpiONu3wsqjwr7mRaxPwDq
3A9DKWd5fLAw8sz4elR6rL6dAHg9twp6zG+22IRSw+vocB3NynR3g3/+s6WY3+UF
o1J8BtROej8U2cMrb7g+JkQ4XyTAEVIZfCxX5zGTZTrjrmmk3VuS9mzwc9EL0EyQ
Oz4+LvzGhzvETLtbUkOSK6kP9VTQFUDdyWN+4M3hBwaqnFyHqHteK/tL3CUAOTW6
nE1N92Pwcdyu/DMYEMRXohE5AAzoUPSiv/wU7UE2/hxkRSYc4RMozn592JwRRUMf
elxkW8XcmQxKlSvoqtTGAmrFpzAeqQ8JNs7snISHbh8c8RMyzsHLVFmQFU1+d9qg
bHQRZgoObg/w5AEVvtLLcm3E10oEhMFJTyJpURKvWx57q9mzbd5gG+wYTGwsw7DX
aPplK1o4y2CDEgkxEiL7IMN7CgcPI+B43sP5+fQpCi3CVciCKe6J7IWJudxPjUT2
3KoW9g6laWitXw4PxdXqh4gQUAhGkcGdJP6FuLG/BywiWjjnkO4C7bBXdNskX/Qa
hQoTIvMRRsgvrol8G+SsQcyN9+ITsjslzv6lNZA01cmG5moSyOurEi9Teo1Sh+AN
B0LcYO6ymnhg1GnY9dCYmpbjzItPKqr9uBFOdiCzgTt5K8w6Ie2jLiHKboIcOd3f
HoAL5Ojnr6EvsDBaW6BjzYClR/Gm18Tm8mr9mJkkLbd2kts8JXWEPHk/nNAg0Nlo
SrKQyV4MnP3pol/Wwbt6Jx0BOSvkyq2Cl5609eIp1WCc/9wuUveTdtRkVDmDCHMz
je50Z0NRClMD7XYr04mxU72yVdJ/D7sMyZEMwCR45FvkD26dE+S5KhATmtvaZcdF
jt/rxJ5rN5xRoMYLxs633iKQLZWGvY4Y+OCsz96qF2+dlirJCZedc2FJFu/vVAsV
8KNfLz9Kv71JZm8wlSwMbHYJlur+vrhV4+nfIlpcfXrveCa+LaXQqyI/iQfw1ORq
nOkR0o1hJmgONk3d8l0r0R7bw98P3lVsJk+BblAxhABF1VJxCOYDZMporEerZgcL
qPOgwsLe1ZJ2IYusDbalVs6CHaIQaPbvi3bfoVYanNdWstQcwNQoLeoK4khnChEV
/KVQf6S14ITrV61Jz6E+tURrV2S8TYpB5emGm8H757Mkw/GHbA6QD0VUhiaRbuKa
9elYDBaTYjppVkMnGpJerMwLkEakex34vFByTioF613MjK58iJJW/mftzk50AdlD
TNzBQzltAsJDCfiorS0YfKNwOfjjvfcIuEmn1FJDfolSNSSkUdQsf9h7GkYObNjy
XonPJCP+YnZB3ngNRSuwV8vM9nCKxygHUNxO+Tn+t5Hg1JLpcr+HPLstEI6AHbV7
44VQe1a249Cyce81lTde10IqQi59uRtLXvMgxS1nlVBttv6cknVqrI4bj2Skn9Ek
c24c+onpUnCdR1jXLC4F0ZXbLxQWFFdrfP8JTqc7MF5/hpHUXjv+p29Ea4zhpkD0
HVYmeGo3hQgVCEFb7F9Rl/yWHa2+kfHamh6ka7drC5gTTko20PFqUHx/vKCmywUz
lzfTClLc+V1WoGn4eQ2KzRoSoj8pyr8R46H0OwNhwWvBHLP43xwbgRAterDkpqja
EVCZGFywUQQaNJKwZN650YqHYdJEEYK6I8fjt0VdFBtP5WsQaYYMdfDUxkcGj3i8
zBW9VBfc/qGBnk+Frb1oAQ0LWcry3L8eg/ArOr1IuObA4YQW9PyQcRYkamTUr29+
tD4QVuODm3Jxx6wYYoCkdRmVWiW7AGZQ8MMVgbE6KtR8ASutJVDMgASrgDp3RmR1
e4Jf/3iAFsqI67CfkKm48NnDf6Qj0D9EDc8TApxqKEN1war4qnACqx6yotQ9Y09g
L3XWi0kT4jeKJyKSfjCAWGzmLHmzNc//XJYnptO2xkTeRGLFfgspXU6R9b8HaKRf
1e7d/1tfKC9jqx+zIUMaX6N4SK0aDLFtr2of9hVhV3tmk2uvHnvGKsJoRrkg/CUL
+uXTFh7FCUp1CSigA7w9Z+tIZzlsgrT8eJwOIAh0bj0pQEufxWMT0VwmgyCpGMrb
BZbkV22mNiTUGmueocPMnb+UFF87XYZo5+qjtv0BtMYo3gayYXQ7dltNkzYgd1PW
ivBsqnp6l7kq+3MZDTzyWLznRGfiynaSk74uVaVYYI9eJqN7fADNyYx586ixeDqF
kq1Kz2nKJg9bNgPPtGanWzkvHDbeGqVHHl8k2qWAvytOk1ShyI/WIcPGwOi/xPPT
RZQV/PvugB0DZXk6syMBx8udpuaH8lA8FNnsc/BsDWyRXqIqkMov+7cUlUs+2WD8
/6X2oev7rB4tTCxupZ8s9RdueNgdv9i9CbxqJmbN1QZ89CyNGHOroMQNdv52gwCW
RnWvfCfL94sDOPucSvOdJe+OIMHK1riAN58VrKf7jnj1f7iXhtnu4GsSrL5jAocu
PzX6i+mzUMo3X0zLpZnBNznzPHFbOFpFNHCec28cK1/lqB22bqg8CHD5ci2azcYe
tC3HDsOBCvVuxbHt6lYdxsNtaLpqKL8fEqbDqKpKQRg6IMQEo+ofWSc4H3l5Jgd+
YBcZMcrCKKGUHxGZ9ip+QT+qznlYpTcbGlnKk3hfbvTzH4o88Vy639B08Irn/HFa
HCMn8qXE/24LrZMlHeJ6kAoxBbulsSpQrE3Jr87cZdGF3bqJOf1xiisV7MFE3BiI
mbtmKD2EzyqQr/px2g0/8uX6E/Gbsws+a8x+tyb00nWOGxLENctjjMsW4MXsSLeA
+pBFF4yHRilW7gf1UFTFcRSUhtlhPz33rWhxwQI903r2Wfw0GNBcG3Kz6J0Yrmtl
dFim7u4cJBTTKI38XzLWCxO9zwm/YVSFxVT5Xfly/s0Ai3ZO1JOQj225GiOdS6Y7
y/EX06tP4GukzGOaiBtFaDgOvLt5781Iz4qSTPQkQH0zfIOMW/3u+xKOyS8cvDVB
3fTTW/n/51NO34ygoBsxA0EIr9xYLWJ4X6LxlesPPiTTeH1fHOKrH+GGuAi3eK7Q
vdQjlKgdj0d8ykSB/Sjebrrs+j4fhfSQrg1AQumLZhZxLzmePgC2oYpW+2GMjofB
eVs4ES0qqjlQDMjoydMMWhXNsts0e+NxMy58nB9F8lbcztTwVju3yefaKoqbYBI+
hp2bTvvuJSbNMR6zTXzQRle+vKt9p46hdjQLiM29K5M02hW4TbldrFH0mOxj4A5M
suK1Ufu3DxeZ9HenyTETITO/ylPvKgEtaoPnjk6qjh7MbB5Zf4+ZsN3+klZ6Glfs
Q4lYiszcwnzO+dhha8aYHXYd69bhzQeV1b+N3/K0b5Ldu86FWQrOuftRL/jLCc+c
L2aicba49xVr83zLosmJAfyQ3/mN/wu3yJoAhL/9J8gOBzYV/QXd+XHxsNcGMKGg
phLmhPlBVn1jT21O9Mn0YewC6843it7X2cvhozg4nwc2PJ/4byuIl1wE/TNn3jPW
FbI5/D9xybcdNthojOBCJbxe8ZISCoVDA/RgYHRyjeRq2TE7wMSLSp/VLjvTfsgk
95qkcInSefLKAwgv1yAPRLewFf7wLB2rztD59OxFYEKqoa4oUQh0ZKiCqhPqCiy/
+6h2VPdGG2w95aV5x+WAwYkSumAKWyS64nznD/NRZTCpnMd9mfWxqk8SZiAYmanA
BhCb0xsg9EbNNMlPxAdhzlBzAXVcj6yIkXd64cQBoLY4bYei4bGi8448assT/6/J
2iYn+so0x0bN5O/WwT9LC0/JmlrLt72cbqEX6ogS8V9hhVU+ABhK7PiUw6EJqT6d
1XS0vFOuFVYBEAWgFrF6zM9BWIijVf/TpvcMBXfjfyAG7t15gCI2KqCsNYwi38vS
Yy6n37G6bMQAMb1XoJyj0TJWQq8f6cdLDELvDSwyOQ7OUeU3f6QxbR3K8FJKjg40
zJKl//tA6lv0DAsQcvYN4xDcMTj3EL1bl2guxBOcjsD+ycUFHYrOTvloaBMzsXRy
koN+OOoU2o8FTnXxEPVLjzsKwB/RZAcVel0c3v+xjPXNeC1qM0GpthWfap+q1hse
508BiFKPE5fIf9L2dpwu3c2fPCwkI+VQezk9HVU6wTD6XPziaJeOeJ2vSaD8Rr9C
LKYTIhMmT0mcbSTsNvHv086h/aFfYUjfQxnfQ+s7KV+JdOFZzAd2vGnX3eUapG+9
XXYScI+diqCNIVUilMEL8AaoNO1fLUnDSh/8CPI3YnG4RjfyeEgHdujHhLvS1EgT
UxVF+bDmEOog764bbJzYdkwMwX002E5td84jMU50dsF7VfAlnRrs+VzEr/I2bzt4
1/wTE2VysnkA9wsJeBJwKEb/uEvyy5wJbYUf3dIdtPSf1qRueDmZy3FclNdt3QeT
mb/6EQ7F6xBlPTuECFeJCCJCbXwzOSCWRkrNmbn58a5bexuXr95gMgw53XrKphw5
5rgKKFpzqslUkrJNGftOfbv1MfvSyfaShxI0ipvG9+wNHYbf8IsC02iNwrwR+rtU
18KyQ82CZ5/RWOGQ32UOKLOOYe/AsVCE0OONUS6FmahQ2VRw4S30TNtfxwDLNKDZ
l4h4Sc+gu5B2bHj4k0oBOltM7d5/Nuf20Nl353OdrzKNjwdUMcOaVI+7AwTztOPh
6g04mPgTh+BZzuqFCIarIX02jdhkixijezXqEnLrB9BVwE3jIe3j0aaoBaFDW5E1
CRBiYTj1m2rpoXQfPEsgDyF8pAHm37tIUaizB43ZanBDWnhKDjKWgXTaPzakXZvp
q8yndSHyw+eGGTAuDBbieTFQ9HGBek+VGe85KkqBhjCij0hjSVKbjlQ8ygSUXZ2q
vv9qUW1TH7HEyPQWrirekIrRLvKZ4tgzNgISlFzU5w3NqgVY56qszFotLXWmL1nK
Hdo2GD+A4Ed14ZTKLF01lZQhFZaUiJ/zqorfqkkCaqSjJ3BIVxvkxvPp3T6p1yJF
aYIkATkwm2fCpPYdSBfXKwuCO9bIXBh+HbxPCxVoqf1xodOzOIDfjRpjWzLKHYge
P5IJsrVYSvT44H1v/7dxXQBwmW+tqFunXvU4ZVOuyKctJEfzUOpFq/8kg+QBFlYm
C2SR8KYxl18N8CK4MeOiIjOQ+qvf7VGuWXisb305K8s1XpblRFH8aK0mqNH3/5rD
zOWctJ4DfVKpKcNERp5pxbydX0QLaGUTPQqjhr8hEOmWTmwBFKgUSfkFYlfPNZYl
tdElN1X+hSf39dvxH8tryR0UXn5lfBeRBgiTYMzgk3+xQLklBB04B9FUbNeMBH5Y
Xf66Lqea6MIph3mfqF2jwpg2YWEdVl4WUCFiNLUksQ0HpJ/q5f5L8a2WOhY6gK4v
SWWqdozcMRQ1zU5WdJ66Xzsvsf8K01ABRQ7SOQ4Rs+z+3Hdn6WTU+toAelo3DdNX
NraA04/hXhTfVrMm0o11D8TfTqpzSI6D3mgp5pBwyC6ZZpT74NBfZVsH4nrge0jU
zXmdhzO6WPNw/kISEY49dgUVTgJEiWNh6IPmD+NYA6tlAgjIyF/+MGkyyriU8tuI
vkWPhNFnfUvaQLjylBU/GDrqaS/VHszm0/CQ+A2YZFpLvL4SiF4HWietyHQFslrh
fopyLmukoqpilESTsMZZvkjkovKLSv7LmeXqcajHdldfLaCx6k1AglFGYy98nnFD
x+DblHGaB3HmqkYkl6KenV/vMg1XwwdFe5XWsmRZ34HCyGclDmzGx36auuCC6zfr
TAsOc0Sdb65ryolTkoqI5qJ/x6dGvn5egLL0XVwVBXtTIgITm3Pta2pdyw1U7zpD
qmVyrBaSdZnzytshCViUI3b2XnGbZ+AmNiduA15ugTFwsqFAB0QxAbP8ddPFlMz3
gDg0qhaMlkRfaxx0w/GSniZQwF4rDNwPZozurlH0G0WwbqM1NvyIFUAvkmYRRyry
LU5LnKqWnaLV8f04Ftk6Uhi2fvyGvFrc2gaju0YVcIf3jje7bo56LW+WCTRi8PiJ
istJxDwJ/D87HaZiR9VEG1H5vhYKOkNN2oynUDZdsqTq3d4bcr2eeexCdhq8H0HC
ULPYoei1Ic6GmNJ1eP7A0Mm7TGj+yDOc+uoGg68qhj3s+dthLOjkZjEDVOqUWqrS
gdGXNpWc60lYHYL2P+4GFYkKdL1zQW5ugBaNRXDjPzody43TQpWwCvLV0ThvoEQb
auCo2V+zmqhvZoHyF3Zv9P6IBrIsZ/bxL58M1vpY0EJ0PmjhpqnWxLgeIYHY44bc
JIaVYeVW3e1yamEaTVN+J+vtKiHeng5BQGjhbz2wOUkk6y/ZxesqS0lBrlZ7Trll
dJ2bXyG3++ycMUtJJi/YZOxlyCsRd/0EKfMzu/UidD4zKbGdvfpCl7ovofgNp2LQ
6LIeapN7UExAA3mSsSLtbqvqC1WkuALDOljIt1YszSe43xwxamwmPQSRsREbcRTA
jP64c/NgTkW6PP2/jBAmF5sos9reeN9oN47FHNx8Rd8e1aTW1XbYE/iHg8/v/fYP
cyuai1DsGN2EwwgwtoazoXVGbwUcXLWolgkq+HagBuGXkn7w1UOxySI9FJiI7mJm
BJmEWWprV95nI7CLVWOwyHgE6Xk0c3sYFYsnp2xC7PO9Y4I2pP54OU6RX6iCp8+e
7WVaCDVkg59A0qwUH9/eTwvCGn59GCAi86zdB8kZ5Qszo47OPEERFwt9yXUR6szp
KMjaJffXl0fAqNW+K/JQ44YGoS8Jn36iw7v4c9EfWj1E1YlT036bbH36H5/iUdBA
I0gAedKzbJN+1eCzwBZoY+6i4IvifzhdHmEgWCpqZWLRafqxjoBfKpjGEuvjUryw
5gnRtqjYj6bEiFlGiuSaZRe1GKY23LSp/ZOa2gKPo9w4txuZPkTBCOZUHiDO7D07
Dz1l96hy5ILwERISaK7AExg7xuJVAC1zxTH+gTWqjwH6pbQhhSMbrCV6qq9cmdM0
nxIpchdUUyf8Ai4xAX8u717N2bQYB9BLbRNPBfgUOrRiSExvF2kilyYq7ThEW+F1
CW4+W2efA7OcgJfSdsT/SMXArxMVk4cNmqNZeqmybYOEkz0Ula+b24LNm8OSsemU
hZ5mgGLzhPOc2+ZHUs0nP20j7QzXMUKjkiF/8LtkzeRXpybbPpBYDV7WXrj1LRX8
j9SI5Xo741IAtG6uoZczeAsCB3CcLy18Zl77XFys0pBJoEWSOCFSsjbJyYFmMaoo
MMBWW9Nc9TfXS0XqmhAaA0YsHCxo8vjWDliFv9r7XNw+SsaLIAgBolhWT1t9qh6t
5sJ8ip6jhPlDzuOPDiXolwIr2r3zMtL98D97q/DbMvPVm5mnTxQ/bmdtCL4hWIDK
voklxFz9qMAnSL56YUIXjMHCZhdXvBpTsZ53miEUk0EZpbbVNAj2htepVo7egRDW
sFs+/Sb62Qudi8+SUlELk4ztoatcCarYFQdfYKHTzz5qA02joQarsUTaJr4Jglke
KD1gWyUOAysyBOUsrWAQdam1gFZC6mvb9966t43y3wiseSnlmUZrSGQ9jK7shaQi
zK0XQ3qWYSQC8cmfarULrIhjheYH2CixvDCvhIea7W7OBFhFvPOuL/grGShux/sR
0iyYlJ5UD7tacFo+87IqF2zv146nGlHzaBrgyLxowkCEyqUaJfs0sGLGFq0eX0yG
D29BrVSw7g5pWdKm1Abrcpg+SccsDsw4oQbTJah3I5bc+KEtTja45sKhafVI50TX
dRYo41144vMgjYPSO4IcMZ19UKqufGv4NmlyaQW1tJyxhWVq2J8tN+g6aF1Csce5
ikim9a/3k3gNcZO0unIaNSVWBXKekm4DgtwE0gA48aJ/LsrfVj3ot4vU3F8fU0IL
ZVw9Tl71zyapKFMKh2n+8OjhoC7md1+2sIQAHPS1ftmYVnOIa7jNiTWmLBwEep0T
1ccIgtxeNwKHJrrKJLHvsfYqb6OflnU/n09bvzOcwjo56DUHEClxzRT0rfH3R3Xl
sNwZHCEkpQsbmlK2r+pMsNQb9BnnsG18La/hn5sCVv23l3xj6TotYxpUS+0BVZxx
uaeq+X48hQGJWtiLAB/2Ln7nLuhfPl+49P+CLLIssDPCOzD0PA3VqgoRAwWQ9gbk
2AambY0E1YPJj5SJRT+dQCLeOAfNrw5IK0+uQtqZro70VSnRKZ7b1kNnE7B6jzJT
AhS5IYRu596N+pws6dnAZKqLv9BIjwgjyjsoCd4ILfPGlq5nyvUsRA2sjW2D10ow
vmWUtVeUPZyfsf0eNudxeOlGbD8TO3V4wphfAvkg4OW97Om3uQ8J5SyIeE/gingF
KhqsWNVd+EbUbEmwcv3FhOzOd1e9ycdQ1sfza+dvj5WqOyXawf79NKLcKNtUocix
3aGy6uPsaZf0KHaEPInbmUiF3Qi37/5QyleDQpxdLvOJb/JqmdW6A5dTNFb0dGKr
qEIs5zD/WbsZxmYXQdqLdfyQBRchoDdgxxMW/+QslqJiNy71s9f4W4+Ps+ZWTGfE
wQs07Q0cEMLxOBsyj5VRcs2GX5rmGf+SehYSCmro+z/cI9LC5rdkIZlLuh2jiGUM
a6htIqVsztJJWUg70Dw3yyYxg6gDqZSCiDnUPTlYRUEffJJ4GI1v0a+fLbxOFKn3
HuseSJKmpbb4FYw3h+G+Ejvvh7jyK8nXZLyh7Tv8KS4P+KA291qz8nFb3dUekGav
/0XCqntA0GIDZ0bvbyaiSeUvS71/VmtWJL8fp9+7nbZe3U1V9dBid6b6ynxRBeb8
j3cVZpfql4OzLZFunCJvG3cbyF0hzU8fop4B77Yl4KfyLucT6n+fu1UxLPOtEnH5
EMuvTkWBMdAz3tjyYh9RoYnIXotAjM07sEMz+guhnqeamojSBG4XXN3P/Jqg+u8P
ATrGIQFq55vg3ZDtNEwmmmCBydZM1EPHALGwHpjaZOZLNVJtmSHOlUk0ODmRvgEO
XBbBqYRONLRQFlKUdW/Q2iyrkRfNZZFOxirBX8Ajd2KoxA+kGPlezjE8dA0cogyZ
pjLClKwHGD+GO+d9jbjXTRQFkewwVrKkUdxv+c4k/F0Qi48IH5eQoC7tvbvEjNJD
J1UDFZFNIdAOOJSfmLqLBKJqLwBhjdKkYHSNeP307ESKFQGEWXDPcd9vVArKBaIu
6wQxlf42gBnVKtyDmO0Ao99PTuKBAzbGLETcGMStaYofQlIOaI/BWejZydhq5qsV
U2xU2BnO30NkBjuhonmO9tWVw0RnBpVqLOXziget7Cu0Gbf3/Wx22S36tsarmXAe
bPcQF3UxpCWdHCT9kmArJGsMjtlRZNnx3Ona89GKpQVw5FpW/vPp33SnfyFiuuSF
cNYUwjoASIM2XOS1gQB3ylch7rLdG+n15sGFMsN+f5WTxY1BSfulU+T2m0eyGCB2
rpHZUsuDp7wCv8k2B3LJ89l7PL1o+vCb6CcyuPbjERhP+vJgdQddUSDjKr6YYQkO
w0pq/wtYsH0d19ZnC27oBuphvAM7P45WZTPzcTw+XxZDc8A8Vsm4nU9VC8+0iHIP
MWPr7Nr5U49mI0pg8cgeHK+ws4i6iGQib5Pw9AcXTnKjjQC0IJ1s1BM6V9cOcIm8
4Tyy2PMyKONnI9M4AgWoSdR0lR6+gIOg5X+0z1zdfj4PCcQSp0I78lN7g9Al4mca
jnQY59BcE5An0gT2DudUYXsb1APvcXZuAKY3WjbaGanqPSPAEgZRskdW53RnE0sc
KISnZA2P54M9zaEIUbnJ/ADTnXgVxWqSX6d21nz2BJyqGc4vKSb00KATBq/UmZxa
Cj/9dPHkNpzkNTkGHEkN7UcE/CcPKHEGh1ul12JCF7cPhi9/khG8YOGQnJZwTIqx
6/oAX1K8O3SfRo/OLZuSlpx7aTRtZxCAPEZlD+GrDCXmtxpQuTzFv+CHAsyILGa7
LAsOe3k09pLTYLApGZbfcVnJUIYB2/oXSUvw58hjixOHaRz4zxNzwxoOx1/Z2jEG
KcpBX12zdOxmvTGEcm1uHbMiPNCKI7H67fQ5yZYaVTZMEd3MuNVwndvRkVkL7JjW
pD7LPdLR+WRh8QJ6sW76F9W0Yyij2DBQlpx8ZijI63u2otuU6jRBi+fRBaLBWq0T
R6t1iM17HMTH87040TqiE+etk8SC05lhYyNh7bNd9ygmz3mORwaIOzWN8PIgMKQK
4pfAYO36gcUtGs9jgdDjnlDE4u2IeB5KF0O6qlS+d27VwwjWWXuzQkxH8qzq4Wbr
lA3ij1Yw4trw/LxqcfhgJopbaOzfq7DoramjGcOG3SOWcHY/chbIMWmKaTmTuCaf
hnF1tBDzTtvhi+TI6pys7qypvwFGWVQfNNcOTF3HOMlc5HTpzO4fXuRRvGjeoE9C
8Li0hIVCw9Dlfs0XAdAoEhwbo3POmF7fvbq/ULhKYVV7yQDs/U+SVpGdTcx2UJyL
mqAbPye/0GTKjrPPA+y6tFtWM0LJOtYI6c52VKXmzHSp56/TlHAFMcPhF+vBahiq
D4aJXg44KmOY6NvrV+09gSWj95gOt/yTJ6AvQzPhF18M82FtjHVXDup7pPr3P7Bt
h0EiFNFkDvXFjDVJ65ypLvFhL+dYi3wQUQiodrTnNmIHaNXDI0fkkoJpgI2VGsmp
f091SBs5CfgrrYGTQwDT3mChSwTxFGnBaQulb7L2axEU8iHmW1PsvNRaNfq55DHQ
g7Yk8ZpZTnnAmhQW6AVAKxTXvHG/40gD5zlARhk94tDGLdJbDMO4WJPaufSMzOpU
iJuSZQ/RqVk/KVXP2F+uMub2XSk67IfeCrgAX59KLGe+GQpeTc2XBCJOTIffL2ae
EyY+r2slHv9U1OcELIzTi0evHuWGwcfHaE5hGiVJ0sM32NHbCOuAh1Se9wBgMCQD
bB9p28pBTFKM1nsADDkk8r5N5z64w+PDxZz5oViESv/jTtop9gBONDjxJC69wXQC
C/ahP+YUfoyi3upJnQ05oKEZp/s5o+ddBeDwU40dbabcCgh2BPpG+x0736MDUdUe
GDX+u1PWZDr5PHwXxh22qR/WtCVlSHfMt+U0T29wcVo5K8m7sSj6IJMOnnmwh38P
AvVXpm7zTn/i87YLtiN2L78GM4PvR++TKoa1MAWhYKHKVYzhtFlEEaugQw2UzvTj
sbMf8DG2KdwHsFNfdpfzMpARhdxaJphT7+aZ7OEQKDGHhjedZ7+1/7DKTgg7i+Hx
dXQ7xd8mmMFlvQn0MUFYCtwsMfJTu6LTyz23zpQwBb23we+A4z+pN7dlXMZsyzHk
sVqMqJnACibXmNCGdPuxSquXtN3uiOayrMNw6bknfbQIikqCprs+GqNmNciVUnHq
VA/Yq1zv/cF+6f8R7tmZ4EoPJKDr/OC4WmFOVFtCQDpB+li+gAak+zr45qdjtDh0
ZHgk8jcAC5CrUR8F/c5LoqsBH7Ul+6bDL4GpdexisL6eWigm5LCuHt6gPzHOD3gg
mqajXIQux7MrxPwC7LnK7DyQK2+xPM9JFagHPQnlM+lye/ClRHndBCoKJsqi1JfT
1v5TF01kx7TITTDHfE/TpedmmK5gQahLvr0o6BfLB21pQTIcFcyUuQ6iF2DXpAkI
S2nWFyhgZ2+nM5PPvJOZ+GwZ6kL0hSIyXy21j18HK7pjzUIxD+s5lcc4rZAecdEb
WdN+lmo7B4A9Vu26V+Lm9doMmsXyaohOZNtyCuxfwwsxMRyr4KfHLjNGvcpVUqly
Lp4hiK1UDT9TCaP9T8fzsgO5qYVVEE2RG+BVNBPdWubdk+GBSNu0E/TEoCvP9oMv
A5mG0hxGxtJBRXMaODLXkrQo/2QYtvBudr42rviDWm0vdRr+C1EElSmzSqkOw6+v
b2T2pByspz1Up5EcJjdTuBjKhhbqztzYkXqtoASBcoByuZV95NSeTjop4DEEbVCp
sCbei0kPgx6R46gm24w4RgQG+ekt8t0S+PbhbBRT6z9f184umWYIM14UU7UkhjI7
Ba7bwGBkQKsfwd9zLogJ7dppkGKkOvzL89aVk7PnSrNtUWPWXa8Ufh3HHApFbcZp
2Ja1wVLdzU5uHSuyXe73XfYm0Q4VzkwXoD8Swvbc0jL1AAwVxWuJ89TLMNFC+31q
4H5M+MTc1OdJrYalJY5NIfkzih8NG16eONcpTsLvHqEj+acBQKptGond4TIrxVtC
F6NAFYWmWPMAPX0p2Zsi3FT9Mebj8F1tuXQBPBA47VAQ0TxqlCcmbcJs5hayef0P
WTEAEACn1kNLfxqd4e5yhn9g59ZXziuTOq4l4+cvflHL+txinM7koN9ZUkk+otBK
sr/noLrZkpGb7mEdH+IcWcnAVBSRigNas+QbKV+mhM2NRy+B0Sc7CxT0wDZZj2Ub
A0c1PTZN9ahnrejYDbDBWGLr5qbeXnTqPxcvVFgF29W2Tw5YJp9njxhCQuM/9/Oe
8MBXi7rn0Br65TqvAXjsQomZW0T+xW7wyCXpBGeALhWsDvFvA7TVwFysLXJ/+HXJ
k/2tpEKzzb0op+LMERISw0uIimUhJ/8nffKBjBnP2GkWk23vIDTatAZp2ksnG91R
T8S7NJ+W7CYUeX64qu7Uj/hM86f/BU4hJEG9JbWHVvtMCnWiJT7EvcoBGcWmjGAb
opDrGAxxnFsVa1uyOklK9D+oaukNwT+gl94511MH+SthRXwlTvqhPKuwFSPw2B2l
7ibwT35cruYrogMj3D7HjUS6DoPJh7uZ2vB7p/vXt0MymHhEEIwh5F+3SpnPcPaQ
tB/Zu9ZBu4hW1F2QnzDzjJg3PjgX9LOCz2sbxIILH7Otbdm2EezRPWiMBAVK1ZtH
Bpi6t3/F3W+LuPgHJkzL9uPxDSURTVnKM3XhDOzrrvBQ4WK09tCmhbBvSeKGYtoz
QlhzR4UjnpVpKeOUsEnunmQiOHWTPs72r/6sghglXOtLSjqHtXy0/7kWNGRn2Hg6
4+fsG6JBMWu+1jFgW8YJhUIulto91YfOhxC0HrV/177ljEbnzfhZu77hIhvuLygY
bY2Yhq43Yn0N21TTQcWpgzTuhfkEalDya26rwpD9o91zzLrCASQDK143avQcTCRl
C0U6uRc6MexWtJBhGWrU3MPN3rIx/eKd3YnQ4cd1AOa2/mYtiT93Vw3uN8rN0LgM
Gmsgldn54b0TnS53xqu5MnKl3g/ZwOEppp/5nKWoG8sWRn1p+GIgaTbWGRmw8zYX
pi7CrnqiAxg7AHsR6y86IJYlHZFLZetd3BHKZ89UJQbWN54OIHmGZ9hNprgagnha
uS4AUv7yPZDNKA8rOd4zghyp+o/wPsatwCYPVbbwE91NHtVdHMAqEhWwXjuxgqAk
pEKuspU27Sg2jvvM4SHSMtm98JTemNXAoppvCcHwzvAR+nk79w2cfL5e4PmqOEwL
sVc6qtLQU7heea16SCPAuWY33jWSbZez7JTWUyWnxvqS/t6lxZr5i6BvQYdKcw3I
xuVZmDOaMFQF8mqpd2MnJUfJh6p3FuhmDeoWzhyR0JTzuQled9+muTmWnrkGnWYi
ZKScg8N/ibNHmZmpNnUGPh+50LiqLq3WPuTmFbiDhVm3fncRIvrN3Yh80J1VMALC
G6JRHkv6aqhWQi0LyUswKtJwkrMzp4dTfBcC5a1hubixAlqBv8Cb2fPaQj17GJr+
aQCv3aD3RpF7kyXAzpjiMqy3HLWnm+eJtkfRYkB1L01mEi/9+ngmUgRjM5LG5jU4
vvOmTTdK1g5OhzY732VaNlKl5n+1nqTPqn6yfdGwt1IN7fLj5piQ8IKCTXfEjqXq
E0xYDezUBh/4gLp2Ip68iK9Dv9rFecSNeSYbS5JYAxvIxtqOPms/mjZPoz87FY6K
XTxkRAnd2PBqAie08pQ05seiyyirc8bJofIApuFjmr106P+Y6EOQIj6RSd1BHZAJ
ydrOXQj8e+/PJiTpSfg5MjpjOHlQxGJFhSFMdKeJCMd1J+xS5k2NgQFaalrq2tKx
xdDustflBtKlaAbsG0jGwhneKGkayK5UfKEo82Bs/lBdussdvtTm7gJgVdpMIplf
/O1rY+jmXJg87ryJY0ZxLSl9m7Lz9o9BGSVFPXrDPgibI1gUYgvATHoOUIX+/5nn
VGVqm7vo6IWEgZ06NMetIQew9eG4klZfO0ysBuvSXqQo7vxmZ7PPJk7snqphmybs
CiiJ82GxC3l9Rlge/DepeqToUoQRv2IG5WBnhmeflv7Gw0oHp1zIpFwtclgaESrG
MOUH7cVmlrahHu0QJyDcgiIIIsp9ylNF3xxai29in6Q61vpiGqL8ppqiBHf6NGfK
CMIH89BEcw8GK4JvgTnHyeL03VyqEaMm9UB9iEZ6qpymBzCz7YX4o008+HESaTYk
aFH6PiwfhG5QaVC5ox2UWNPLqSzYlGYinJaDuab6lCdWPJPsHHF7CZEMDZs7wrDy
GJbIBVGudc6PJkITwOMA7Y2PtUP9OJGpbLaf8oCzsDVEWaJnIA8nEV/aaozy54Zu
TCMA5Z5B263NEhqqEBYA1qgA24PZtjJkBGYYQG0ar3vqPvgeyiJSR3MMonwRx+nV
fXIF7qWnkFNhp5hzVBk6NHfB+kNNH4aREN8ZoFvGBCFhocMBzpyiGIw4fJggUMhl
OPdPUHKh39BHQ2qtAswAA82PeNbrhFM5Zl978c66GVBCT2PXDspnnCfQ8QW7JXEs
BI5tmnVdcG0vy+0tOXXkfDRorutExEKtLMHa2bdpQrIPH9yQ1gQkEUua78grIK4x
lY59faqQqS18q78kC6f7F37qjFFEDYtmkANV66XlWWFoAaaikO61fj5M454TGNBU
eiiwKaF3oefoZEOpRjMOuMWtBvV4aVzVGgKXwrSxI6wRRpenNMSTI4oo7ThsR0Ij
4St1AiigMzT+E8vRIV6K1t+xlOLjF+UR6khEg6/v65Etd28kjXAg1kadM2amefrn
Jqsv9XXGJiWruCer6t/whY1bzgGsP488URRKEFNvo3jMPn9F4hqzskeBrzGZseDi
gHeZD3llocF/Oz8zDadgP+rL45bNduO/YAMKvvZ1JtNcnNfoWMUxQIeIq64Ky19O
vcf4o1NnnOwBrYMIaD6pkFHeTBRj6TMys5x49S8trzkP9TF3tUaiMyVcIqAbKY7m
gb95FRgl5bbIOZB8+ELfM7j+VLaFDrf3T0MIrfhD2pvJWE4p8Qlnniro7oOjIFjv
hI7MBcfU/wKMjtI9JKf5+m9tESDWJ05nKYv5pwFeHI0+b+IRnPFNfqJXbGkSqzLP
qPKEjfQCQu9NY/s99TSgWYcTbRqKNpL1x608CJjNn7FgmOYAzhaIYq55kgk1Rt+C
La6OaYp31VxdkjT0AItkQpxYDZITtiZL0nr8swy8J7QjATlsfI+oLpKBEuqar6WD
tAlSIvnTrtmRG8y/Zem2tCy/fiSdA5P3Vknhvb2zdQxOuHY0apN665SKqNFDDgoa
nyBm0cA+Q4vHkpeo6inBXR/z9Obwdocjd5qZzKMzYYKuqzMXX1Dj3X7zly6HpdqQ
/a22iUC7XIG2zQ6TSfFlTMr9Jr2pnsWGXJJWeahStnRptHMcTVWWr5zl2kA1kcF5
wd5LGRlAWnTLJ0UNYA9MX7f4hgTegWk4UhZ6B25U2p2AsvMfchpoirL8/9mbzLJB
EXWy02FqtCnYzQo8wpsyZ5VlxAF2gHsm4FA2c0b/yupumcRAfn/lfnohLA1HRPNj
F1o+si2ZUbGgbc7/+b8uNcAKofETPQHcXDa9dspJE0SvRBQOaQphjG1V7Rt3IkHk
1KPe+sJ3QQr8MVbM+9cUVQYyhG5rsKYPa+etfxcCAjyeFDEvyz/qA8oh1cwX13Jx
XMvju60h+NBWvQV1e2yuZwWvHtJ9fTvGpIPgsyKf482buFOfGuh/tE6nMBjRwC5c
rSUCByf6i5Yv/ZBXj2be5BnYtHTG2QZcsIY1awKtdiwElB/9suGTGZ6Mgk4jW29W
NfWOxpJq9KkTiuBDJveLemILfhSheIqtVAssUuhSpCEIq4xWNjW+sXqY7Q2gpfEn
Vba4kmAoeLsV9GJTEy5m/gugC/h75JKQrb6DDFDt1IDdlOsP2XzutmWwae7Ieopq
DeYQDMxtYMyWDBx3Szrzb4cDdSnsCF4maulKPImICVudVPIT/+ly9F3oxGzvysv2
GqBb8AI22KOvzD56EJleuBx3JshlPkK8VojQzyVwGdtkJWDlvKwZZHUOPxQnpfu/
tLEuENwEbi1vLMbZ1jfC8b6PXig8ZvqR9soH55Wpzss/47UyXLwuA0dJoJZJrwiL
FVaGEB5lu5kgFvC0sMA/TTCk880g58v83uy6hZr58EdCNKPpuv7mG8hEwjF3+g4A
bqCmqyKZV9w+RawHmipcYo8Ve3PMT9JVVRXohQXLImqjtX0IODzeqx+55LfJs2Xz
hCughAwm8YNhlwCySq0XEJKSuG7m4saVcCSm+DtF0SrrZPzg00084RjgmuOoZD+P
kPEZhALLVsvPKaAyF+qFtBy9WKNMCHX2Xv9ZxsfnH5prdWVDVewDJg2nS+dDf754
UJtInuTA3X2HM0iegCIa6XANFS5atNbCmP+pDBgZFm5fZJnvJlohvc3uDKC/Z+Db
GyQEXHJEqupyPWMJ2QZrl2GI/62zCHm6sN3i6Du7dFhWrOSRGt3k9wBKu6yg7Fsy
LlkZ1y4wZPTz2uU4RVLxyTSwo1BIZHldCY7dV5E9ktIFcxHuulKHAi0FT/9TFVzE
fwy13F97Ex39vLuKw1Wxbswd8gQUJAd0gghrLm0F6dPjIxTge811kXoC8dCn45oY
WO16CYbcseJOwk2LnOlZxjRLzrza27EmhFNN2kSKtlUaPZGJYHsOVDhcwYnXg8El
2b4Yamzk81Bugqk/EzXuYqoNnPCoF3L+9WY9vRhCyghZ0dNeeoi1YNrXVPE7q79Y
oLBH8yX12NxtRe4SLaNOO01kZZ21j8XAAgK5ZIhpIxMtdA0MB8XDzvmeF8Z5/jRo
twMLlBTEkfAGohPfk3ecp9bqdRpWgTQveWl7xV1EmiCwWGTwK41/brpnEdwpjb16
Et0zGqQTaKlag18LD1eR9AHTwDNIloVltQjnvC+1gvQPH/znO0bCHnH/sSsllkIZ
4aWHtT03hXmHxB63GziF+i/2N6Rh5GUgzYXP+VRcLruVBRZm+3Ea6/o1YfZz6ZKk
RyAz1dmJLwwnHKkwfGtDJzkHm+bowtcNtjbUsk4maw6dLjIS0d8OWqUuPOSgmZ80
7Or1hUj+Pwo5d2qiP/9r52hwdvVkHZQVoqMZ0LWtM2lzOT8sqKDlgAlCv272mFP7
8a0/+L+Qp2msCwm8RIr+78rzWaS7i29BLpJcM6qCs9bUbklckxWG8FMNptB5B1IE
KHEKrx7UzQcQpmX21Zup2u4b8tUF2Wgk2iG22zmqnJdKDT8pzkS2rRaGz/ry3RcA
+x15DVnzfaLBDfRwqlmq2wI2bo7HBTlIKdyTK3EqnsSufQJCW5HQyWOBkonmAh1a
geCmRhL2BvDZUE25QVArZwsAL1CbzKNM9nrTJ1e3gYR3ovpoE5cpHt/NY/kt7Tn2
oj99mR6aIxFbziLuRGGW18ufaOA6DTCgcmaFM8X0o8BjArESPm9pr+LFlCZvMqan
jJzxRqdt9n8nr2XbwmuPcJB2SIZBTG4N1Bpz/1iWbRTVzY94lGdmiBay/AnNKPMe
NCdFsI9tRQDZ88wC/du53Y5rtlfIdDVqfF/5xugif81P5HSiUrcoEKeYFJSOgUIs
wmjZWfpWsPjVHvOplyTKLTKJRxTKOhqzcgZmiY3y8XgkVDv3muVlJKxQp/SaR7DA
CrjS7LX9MDt4ptPJnyKSnaX7iYoVmYodpyTogJOQ1hP6PHKzLOSvUlh2g3XSffHL
YclRJ4t+F7oytDqq+cXZ2RTIdEuKYEZ0x4ynuDgqrCZfz1tC57e3VE6uHHDpR28R
uWVV5XLdyK7sj9JIleS052iSQCKSP5qIwzAHPOXpPytzEGGHZuj4mmQ21KOBUV3b
gPVwpi/9MShyeKtZpUyrFfv/6z/PF4U2d63T6tpxWpRDLVpXlIH9uSCRD3u5O7gx
yiBJHYGO6xghvroqfvepgOMH1uaZj0HxB0Vd5fPxeB+t/8cqa2llKVr8lJrXjK6v
wNV3YcfEEYr8tMzQCzMGwCgdT0WdNEsYkLDlC0A4JvVPa1NNznegRSdzHj7YlKS8
EtAx/Zh723Ae7owoniGf29GT1Erxp7z250j1ckM3NoxkQ3YYROtQVbTHXsrGVH/v
GaJ8Efyq+xoaqfMIehSBYES2a3cuo5Mco03gcToHal7VJxusogPNNby9txyYuiAS
arwamG3bVgwngzoCNVzMYIAby93hSdU8Ow7QFpzMEu3QXQ9EQDW9hgHwPX1sXQXf
c71jeuSluLyEY1aFV/0H4nGU9yt7ROd5xxNGy3ylhGn2IySRL80UXS+A98yzh82o
IM9hDIRrEb/emA773Nsywm2eeTMMdxhsZSNgv1i3seAILOkX8BqN9Xk8nwK+9TPZ
7ypWwurGjbfDm8uVoaW8eMpmPTsTRDFNEFAi2uNiu8bBrCgfVC5HM54zT+x+q0NE
XQqQ743DlzHywVlm9Omz64pcdOi7jkZxpcbn2epSZ98UJQQQjmSUisS57EEB7sq6
kBhRcjKwfimxluN7qKy+9Tn5RB+CvqnsRD0MmKUeqbBpiJDNm+KZtaZk6K1joPTj
fGwIl1an3M3Zd6etpkdncwivQRhcfmgbgRWy7TK1E195QEw1j/rRyNJoi0sIpPpk
D2ssetoyoJnKPZxW7Wdodw7ZhHa2A0x85vWq+ElJ8zcilWF3wd5W+JP0wdpk6Q8L
GCcr0oHq1dJEHq8hUIcDDZcVosny3iKtMABqreONVVM2e2wvL8lIGy1UAout8UDq
s2dycfCAP/eE82yVvHpKIhon64rQcr+6CCxSOPxdY6alogQVd7cK7quWNctaQkx9
YG0FyP3k3IrU3iXZi8jOXwI2kx3vRo95cieFy1Z5Dm5xqR4F+JpeDeu/p2FCwn0q
STMSpYh5OH6a9WwadV9B/6zZJTvpC5x71cEZ6ThATwMOXXlnOkqfSZsfG1Lz84kY
iPKemGEw4iP6sZUkSdYQOljV5ssWjppI4TUXEc+JC3SiBmypgiisoa3Sd5grTX+B
jFzfPhH8Uyii/2eR5K1EAsWNyKbnujMNzhOPkF1KV/gMLSlVSCL/jdhc2FxHIOOz
H37urdG4nuo9Zp7rbaDA6MZPnk7sa5djECUkDh6yXeUoYN0JJRB3PA7/qp9Gies2
V1XXHMF0ZJpVOOylm2l8AxkEBhlVLhma1h/oarZnaL8LG+zgOYeoDzItpO8cmK2r
X6pheDE1SencryjhO2oyqbZ/7fI+Lv6YHbFx3Jdot98WQZAZAwEhnbwml7O1dhCt
F8cm0xOICNNCEofqUV1oTY7wPOtFRd9HJC4eFMkh9l3URLwEyyXYlT5w3TG4qA3g
umGrfRBjI7CyUkoaRi94FsGcOjDtysKoou7YbeGY6zJOtBgqr6k7f/5E5FqVqtnk
qkv+6/oT7fPJ3JO7vmhWxtk5pPO+U3g0BM2JE0rt/b+GjlVQkE7D9B52/QBCPc8C
b5E4/10kyu4B89xqzLBDNaYl61hcO7KA4jDsJ6L89Zkvtacu6osSGYmRQ3YSM2x9
l5Oz5BHzblYVw1QLxBNRCmBb7usH3zhuPwpFxK7feDcUe/R3h4fruo197V/U0kOQ
bqFLByFLc1Ks9FVuiVNYPwCMbK4Gk2dOEZPReXtUFoBEc6KhxxsNAW6Y3Vz+xZWa
w94pkfu5HioRGA1QpHEfWSdqN8gff9001ST8Uo29mQTNbasUOM6iOYpWiuepkjeJ
MEgnWNa5vGW7G881HPMU1QxhHC8RQYJ7QAPcvuXr/3mAfabi0pbA52pQ34djGFD/
WpaEj/2mAanz8yRl4Hif+kkkOSG96DvSWWBOk0UVNCobd89bZo2FybUXvstiDEsg
Vtpl93Y6biFSbt1Qg6ViCFnQRaB5vwJ6WJE4dbZLylqml73vjnXHBSMV4GW56Tke
DvJWLiWUNzSR6Jad8UEXogjUMesVtx5STgO3q3W+BiOu2ASGRsIasIqoDdZI7zeb
d7eUEIqs19/F0sCjTKs2BnKQJ78yBM4f2y8OSHfwJzl5gIo7wRWCqKXjRLwX18YD
vt+GTGqVXpIu8tpwjdHsss+8xyzYd5hwQC+oha7o5o8ZV/Iwbi+vLXF3a8xx8UMS
VyonLS17o4xaGA/LvkWJIMipEu8QzYI7l7GkndL6Yy3ajnKvei5aAEVUole0mOuZ
hgcqoimBQ7OFJburo+2X4MWhFQifyz/lViaJD/nGB3WdrDqBNsuHAlbDj897d17J
AXLDnBYDJ9vjFO/7xt4fW8spnW6oq+2hf1KduBZLs4I7GcYEV+WdSH+OQCT848OZ
aUjF/Z8EXs84aX6NCeZkTtchzgjQJ2At56sUmiML/8fZMohP9nPVsqZG7oUheEWH
JGvFWzCTzzfH0+vTic6hte2XM3ITZF98kxw/UN+Uf/xLQjm9uOLkjxqk+357Rn9v
F/XyoP+iTpzyqFJM9VPKoMfrZFzYT2rsmbEcoDvZtY8zByj7ll3UNSKooAsvhpYr
9OcjV8jWdL9NmXRp778CJeiQo62w8K4GD4mQ0aESng9ctW5vRQHbFZA91vedF6r3
AJXKr+Mauf7WOfzodBBt2d9y8ozXO1Hv/AvmXDMjZsrpHDk7lTLAZNOopbiZYNaE
t9ifJ0OjEWia5KZTWbAvczR5u7+UuucuqYawkkZpPPXWyL6ig3EkDvMmRp66PccT
vlSd3gzpO0JFYXpyRsxLyqR99OC7s/Ee+ilCUuLkMBJwjfD9+4z6PwA8ACzI7sJ/
+ieeR7yzCAQUt5nNkZUpvIDNWQmbvL3pIXWKM11Cm6sh250H5Nlikox+EE7uy9w8
d6cM3xzR9z4IAzyzQKhqjaeniqQtep3TvpF+c9Hqcti7iO36JpoCVgDKMl5PI56p
l/KzRLWXPkD9IY8DiJEKE0F9/KZEguxopb7j3tcDq5nYquWWykSOhnCHdfiGHSf8
/faeoJBg6sEP1cVDYZvxryDRmQKTBwUw13A1r/RVa/lHEHGftOmALswCapK+k3va
xYDOK++Fbz96+hVrk94lr6Gxxz0N+1f0ucG+WBgZ3tlseL2yS/p1LzkAQbaT47uF
qw35IMRF3p1kBhkuxcLHul/tg/R0VuAOfXx3c2nIPy8PTx8ehNNR6LdYCgUGd6kr
OX5qYxsTnAcjqFkO1ul/xhONXM+HA4J/Yt/K66DWk+cwAGFgp3V7VwAwgntf73Nc
okEcmdorcraWadJ8wBNegylzRmqyhxaKqM1ub0wrkkrlBobkhdQREsf6LmHzz0dP
tmjCv79xeHxusNHT0pQvW/Y6vwXHqY5nII4RpZSzM/3Ksm7S+B2kIzC07EsrtJWj
bhsEQv3h2jk2//iE7xLGdZHn2IBEX6UENNpcpC0ooro3uoRi4wZLnmGEso4/EkPf
4u30iRRIkpzXpw7uDssFD0pzzll8Opkr0mtp7evgMN/ogIlJsrYNcDMkhH6thfIi
Mlk2OosstXqU6SMjQxnkjD4xNOCYXSe7/HEz8GRFy/exR9vEgBuIHIu7btln7jrO
VF6O1wUimBApqSQQn0rhsNPFmc7IqZfpFWt59c7YE0w3mF7ie0yurAvYF9rFNQt8
KBJO84sHty+nr3e7bsARsLBxzm0NosY5g0NP6zIwdqdTcGByWW5mFRsM3M5HSKrE
dSGGA6yvQX068ENJoSDYcVy8yATvSS8mVotf9KfMOVwTrKUpTB2CUsXI/bIrzGlH
RCmpazOFbptRGPPEv5akvzmZqQ3qXy4kEroqdGKvYCO9H3dO3VVDCWNONvKfGAo0
PWDfGYg6d3+Xu/acoRM0yaL15F7XVzm8LsmdMM/XHrLkp44dtHMsgfl2Jf/naBgQ
C17mI89KrUWIkc/fmLu2slewzVy7KrQnJStuT2ldY7F3NNmZ3Cheaq4EjxMbt0JW
puF6Ggq7YB2Ly5HvHj+Tom8owoq8kOYRkNA5qfe6551qnDPL6MmZuzE94RYWC0qV
/Fp80W+AWktNUIvxn9rNNF+caacty8/NyLd4tL8lJ+YPRaKvZv36Am6nPT/89KrV
tFANuTxEhgsrgaXgLsYnb7g1igbMaxPC+I5yurXlKBUMBCFn7o8BhcdtfL8ENUEd
kLi4TZ/oCPBxl7WqhShIjsAd/Kl+orm4UjjcReiVE/ijJZID8F8psZs/QPgs6jn7
gfD0wIDj+cd4ZKRpKcwlgFVGENp9Vcf7V0+et2I1fytlxi4fdSklcj5q29HrCjmo
QJaUyBKMo8YM7HyCUVZzaOzLDxEiuUgL958HaNj7o9qxrekA6agMxiKej39U6ZFj
6k9/DTvTIZ1DoR+dvRwCIf31QE7e4lRIlre6ZEvxRlBDpAWC/5mvjG4ssz7OhXMr
LotubtrChdO8Sd6WvWeTTCNhSWGzoZOLtZNO5KwPh1REnKcA0PZ0CQpoStzxuSQ7
Eq65DOSrCaz3Ii5FQUZyF4oe/O8rEPfgulIM7SwN14f9L8yN97nnH+NLAm12HBhl
SCxrJln7fhPGUVrZF6mblPw3m1fGPnsNH4eQ12oC8fpblW+U9d30s0Qwn6AFJeg7
qxqku+jwUxKiQlyX6U1CfDNGEXD/8e7NLmTmnl+FWhLIvVxYxS1EQCwQPQc0PPlZ
pu0D0/b6CAs/oaEVYjEHrwxi+9j7A3KLg92lWcV6UjumL+q170skoG5isUpuGoSL
fouTmukqMibVBkvVoZlXHeiVR2QOFOSkT2ixxo8yyuzIajZ2afsbhmkHxxG5UoV9
8V8zOsnfg2CAKfclEAi6eoa2xWjBEOAJaduQzzPuXPqest32GuOBrIaVRj4LGVp2
qwgvAXNaDTOBgZQfo7nEdyBwZYwhYY0PVaCirnOyYQ/ihcUQSBWmO6Kjoa+in6He
zgpB06H/02ErC/CZl9ENUHkcuq4xDBWdB9z+kUHO4Hes4v8QUYDh/aEJVx2U/uSG
Wpj2rE7LmqyzCiP32vdpAdDTCpe0V/1D/9Yl+q1l8uas4NAwftv24QI2T3wvys16
HlVbLkg1luZUpCocp2QK2doKUa/dklhLAjK1XNSs60c+JJkU7lwo2vFiSjX+QftI
txUqSZNxKn0hJzWbYvNUrq4upDnUFsn2pKwwDCEW0Nmn6FsQyzgtW0TPydC1PaB1
FTCp6EBdeU/OJUWvg/haBjZYTphq4hVgGJALjCgKe4keaqf6Z1pu8/3xFjbP6+a9
XI/dKItepztQZGlPNtApE9NnNPjpxR3lRJGaR+YTVGURbG/cQeSczz76vI2Au2Su
CxXLc5A/tkvBiHz5Ydx4oQwpQdaNvz+MjC4Py8muZVI4nV9y6LgrWHrV8zEw3zmi
MbLFp/ts3lZXWi8yG9b9psLNFsEdQ6MJBMU9D1YKZ/CJ8+m/xf0sVfHNeFTbNU2M
s15hVGCJlQqEnzGBYyLONE4g6rg+0ejMVKKS74BHIou0vIZkv+NG22kLl71UtV/H
LANcs6+CR8Twc678eK1eJE2v+Rq+Ds06sVO0cc5EELZE1K40SqJUwPpgx94RrHSu
+MSLU21LHuTCjF/jS2Q7IPUSf9A4lNU1gKL2bYJF2TW4s3KuNCdDXGzOlBCYEJ0P
mfjy6p13DPYTzrMSK/0/ehHtOtbePdi/tHvRQF8E5/KEQa8BkwaBqxpju2z8lIoE
6hT8s2vh3HJBwfkd+SpNCiBlSQFXzEYAZQq+aNBSRLcAxB0uFqr6nff2DvNuXWWC
ysJvXrK4KQs3IqzFtF4keNII/7V6cOzCoz3GSOFrbDgzMD4KLDMsboq/B16RAoQj
+c0Sr/Cia7Y8xhEyNLlfLXorWpuSobSJ0i/9tMERdJ7y6/aKBmh+D/9J6NWG6qVW
/gMU3fO6tUQCRukduihlRYecrITBHTwwHKVTid9CnkNabooHxrI9yyHpERFJ91Ly
m/gYxcJohDR6xEks8HvlpccKUIVBCQEbKslBU8drcy5H8xCF9z2WDUP7UmKyk7qJ
uFFfNwBjnxNNrQUaEWkRkZCCTL+i6WK63L8Vsc1zlY+mjpX5JRyaXp2Ra7pUBI3j
t4sLUn8hLBxxHxoA19GKMK/5KU/GxDJrXmHOhJTkz86+sBDNcxtZQd5MfsGyAv/U
DyMDdvosONMRF2wc2DeWGYdkc6M2NiKr4mJXURvoCR+FNNMz0skHX0Xl2YnWAiJf
gUyjruMHslUP0KXngInlWbhpVuwMT3/U4hZsVxj6d3Y3FgYebXt3ybmcj2M6Im+7
Mq/nPy7+eZjkkZdjx+P0hY8WYDIXiSWozm0EosBufO520xjZPgQg1NDv/yg6fNfg
sWWJddW28YvBPPQla150JyAksMmeIWlGoYBYwpb8cfrQzWbL8pDp7+Ax5wB94O9F
PeXBo9D3k8ldH6WfW9LcVnMhl1ee4YWF74bLqiYyDTfvCQR1vk07O5oV5ixi3r9M
k8HfyS+DMOY2otKp6PKzkzziffgka02Ov/Xcotj58zP70unGN4pH73YkDXSdpXNN
XbD+2PI/OSkpFNcqsyB3sMHbwluc+F4IeRlXVD5CkNlGYyr/SKRl6v0ZgJbNd7J6
8Hz2iAfuhjoomPHuIUtb/lYgV1hPToT9kxSN21/67rz+A668H2ZeH05VgQ6COI2K
uRvIWZdUVYzFC49EjjxeWgHgm7B7isfFb/XEfdtaepe/40Q6Mo2J11U2YFEQP1HZ
kDMMpsKisp6O4AosUdbpnuf6dg7KCbGXblbGmPzIr5T3z6um9YO4aB9Fi46gsWpb
XIj4EBPXRaJGceNf9EsSuTU+7yieAeh2Gw55a1wlQOJovqdGCmGSmAM95V7X7BIH
aTqDSkjaAd58PDtYvvXacT5aNr4o16XjBW4KGrqjLAZNTnzreGUTkAW58uSEOlNw
fUq3SVI1CbPKXB6ZIbvHiWsqxVJs0r/Q10KYHMsVY8meePai3hk/Ok/qh03Qi+pG
r82/fwwataxNfT571rQn4fLwzMUT2IOnMpoLUMgmUhUBxmmRh5frnxZQiXr+2lj2
PWWqH58mTicDGJ3Tsd8YVhHJYQ4F/iJXc7vy2/w3/d9RovygdPS+Hb7zZn4zf/Sr
rY+GPLfWKbEVRKd00EebdMCQoQ4SEyg6VNMoL1ag+ruQojh5ash9gKXnQmBUKdZQ
AJE+DS2VCIneEXX/7/HhAHrj5Ibbcy4l6J6mlIHH7AqREBYvJcbFi00d1oUoze/X
wwtQeVSbkRP7szAJNX3bGuvfg1xt80+Ayr684WoVLrummvY4W4Vinl4rXIGucgpr
emHQMEy06v6jx1uZwq+VOHRbtnISMNwyPz2A1NUhxZBICnqF2xQCMxLafwEYcPy4
ApZV2chvUKaDA3X0FcPVuP7c91vL7ME5I1GVWs2JPIGQfyWVwa4CsqsCMut3Swmb
tP0340LJ8uUuRjA0GT9FQ26t4vo2DlFQwmk6HgV/cFv+eUSM+kMf0rCi3GJKLU81
91x7HHtoEdTaOXNAiYR1Akla4+wv+FL+XCtI52vDWTnazVapmjRkCEvfU9FqSXWh
FAa9w3qkONGGiGO76+WAC0NFsEogFumXSl0uSkOPmqmUfVAX9iIm7kJb498vgvwi
wjAWLvH9bjWh/FHHruChvvEKUY3O26JbLV/jkLr0UeUmtbJCiFVjzOmDvLXk4LPu
ta4g2C0h9zKOqKd5a625NW/rcdYgSvxowRmAI4Ye+haSF7N4q8qj47YhHimA68SS
+DvoZqEu2H+zbuNm/fmpHyakT1jjJUHJZ8YCBL6GQxctDk5rsjVo8+tqmW1NVLFj
JPeFUFfjbESK2dR+v66Q6J7elSS2wnMd80Yee/h4YmsUntK7AbKHB8qVblqOpxQa
fLxN1Lm8ALF4njgeFluqvNwLA1CAjIHnd+UGIySfcUhvt4gNEWjf7vEbg2ln/kNx
JDfqDX8lmvxVqm1y+oyDizSvpQqIHuGLHmHVIuML8p08Us3j3PA5fbfmzD8p2iHX
WUcVyK7AngjWCWN7k05mNSJFjlTDaKDUjWB+3ERNxJsvXKpq87X+jx0PfYGLArfv
Kto9fKn10BT14XGf1HI+PM+q/M4wH+J6j4Fyfl4gH8qAZweQmcfydWNASHVpxev4
2x9edmOxYbHwuMl1ZtB53sncrXvNVB0Kn2nTD5ebtrZbWfXjsmPOUl1LuXR9pBJ7
P5KC0a/iKsybxfvlvz8I5+Hwh6C/SNSxKVrXss7+HZ4pGx+z7hefyjhwfO9jDTNb
DekUBMykR6WXDm7F2VWOZ3PcNkdrs7p/mCPROMUC9b46zsbb9maZXJKIRpfIe7sv
KbxiVaT69Ma+Bvio1vzIIu/Vx7Gjqm7l6ZG5Q00nGAXFTYfINReP2IJT/hVY5iHO
H3+q/V+WLTZi7BhgfnFu4zUti6+SQ+6H5nt7VDD7K/q3ihRQWBHNa7/cLOrKNc4u
mgNH+hTnzOlCAelaoiIQcY5hzVyQVdAkBNbsoPfMV4XUdf2pcKnD/LPVEDF9lNfO
xtZoEBkM4U3HG2KKThuWvOUR6yTXuDuuU0P3Tlynykw/nYOPM663eVy6ft7gE08K
O3DhykgMaF5Q7MF0cEWJnSatCtsldBTGF5M5nSAgffsCKR7s2Ws3wJgq8BpsFYrN
hcn+Y97W+l/OPB+RCx9TdCnZuU8gZz0/YY1SNADRFxElArj8a5hw+aZU6rxpdjWF
TbSfgAm8fLI9hbG68j3i8eULCBDFW0meQiqTFv615ep6RfV1SjHBtTKcxxBRHjHE
rmrZboC/97IicdgrbANRc4fJW/5TQfOoif+GNXmV/jgK/GLGjoqsDbM/YZp+lvBc
xQqWNiU+BMGzttO8ow4WBr8s+hI6PDcxJsN/jSIpcZF35tk7/0GVuyGjgJUr4eOl
8gAKq0NX1b1r25UCkG9G5DqCo/XoLENCaIfWcUWxS8Cv0mzOmGbgEHtEjiM1iH4e
i0uZ18Ya5BjT/pvZETwi8CQ25RCOnJ2AjplwMmnyTE23Rh7gNR8ICu/ajWf9P5iv
txmfxMQ4+rZdBMeQ0VcDURXX9UdF0pLfehUZGGyaIgJUBRHcIXmEc5oqDYZTyLqZ
P9AmMLo0bjJDon/g4JQ6OqJl34H/j3bz7PIvGrEjX2fU6B5YN8YBuTm7VgIQkd/O
54bQj0Ky6kQ4G7W/p1Qnuxr/MJDMkvq60kYjm23QzmstATuPzVUmadTyM9eqhFf7
wLUYQ3pD7kLCKN3qAOkNyp2c30fM9oW4np7BSX7J9pD7S6g9PIZDUI8kdZ88ytN3
WkY+y4giiIHqZm2TEZMs723RFhLLduVf7kTfwIwkc7rlG3iIJ5mp4pbQoVY7kRbp
Ka0rzMOZrq411q+0irgzjn9u4gE3Mx4obe1Ic2rHJOhQLW0jNaocPF5fC3grBSbf
fGYxBGrkAEyWFnhxvzQW3okLhUSplRClaODLueRfMMUhXVXlda3Hb++S6XZRezo8
Y0CaDwYOT4oBpOgpqXg+TFVtnZM7cYPiK7juwTPiFo071NKRci6aEjQyqgdJs4gW
RUpL3HawRQYruWG8JecttAUGwExL0IRlb3Hbk8+8KuJUAwwTa1H4bpBy7Kmk55z9
/QAArVDn0303x8tGrqI+vrpQeoalfPt78qvjRO9JjSj50wlO4lshZkKDoeaFaOqG
uY+3jiUmZeSIoHWmuL1QOPVzb9taMNECQmRkiLuo9BbgxKdzPqy0W8rnldBY4nvM
8llEp5vdPGIHViyiIcv8mIrlBhpTahM0fJ36ER6RTwppu0Pw/UcOg5OhDOuEc7dp
AnTddBnVyvmUpocP/wLTk7urm60Bh1Pl4RtR4kHppGxcY2PPXVvtE1LI7f0C6fZ6
ksSmQbFWFqkGVIiPIZvUpPV8VtxdxTwxNVauTD7SVfN2aw6atYYWEsYX3lw6W2Rt
XjzHDkLsV2B63OJFUlMXrUtbJfjz4zPdahLpIhlUZHbKRtq49YhdqvH4xRid/8+d
kF+Q5JNzqTF3l5SuWBt/MATLK4KqRECFI34y+NptRB6kAxwlgpSsNZ1Dog8PjtWS
j05AuJkfpC7ny6UE9giDSsDpSz2DVOE8qHc4/OdvO6dv3ON/yFnyrw8hXDCO3vLa
696VmUZMSMBcgKYiQgP5GbFsPd8Ea79u3bdUwoQekZ4fJrf8Hxq7pnePTp0OIBgD
Ee6VgIwa06rD1mlfJsbd958KZh9sAYGf+j/8VW9FbIbBm8kHHTeihTC0vKE4mwMJ
WffR7FdNJtfjrOJUO17BWqjtLfI/5DOKepK6ic3bvjuHWd99feVEyDyPK5vcTm/s
7Pwbq9QKRtty0UYk6NrZf0MBtCb/G150Jo7Ev7CoDYPkl7whyG6sPqdPXSnPFZu0
dV3vYbU2orYR7q23gE510wjympeJLu/KZr+SF35ut3+O4nPMJkFDMad8WlGVR9We
hKR27RTVMx9OSczK7NqoctExcXx6rbbJBgMcUOxQPGYxx+elsh1vgbTcw7x0OnqW
drXXdMPi/FFuCexjSzNnmMoZWzLRPau/SyP+JuV80iHqQjJ6AwwiPDLGjwDwOlEI
tlMca7eUCW6v3wT4smop89X4HkLMw5e7RtL4ETGIrI4YTzT3LNw6aGxmkGc/mPef
c6mJ9EOPKvF7HMEWgkG0GB+MksChu6wnQbe44XK2JEf2qe6KasKFcVctkP1wWdYv
uSnLDdC551DQyb/ZsgfLny+tXRyP4vSNI+S6Kh90EBSl70tBgmvnjIKkYifo/Ghy
le+6rcl071szeZBGSxcDOADRfLaM4PCmrTmLHon1UeEqZUUUX1M//mLuG1GjZgN1
j+qSbk3+I3Wr0lLt5/7k8jj7XTTz0zpeYXOrpObPz2C8gJQ3WBfH/uZDeFSE+fTb
q5jSngkNROxWxQW8f8PcyZvBZdz2JywWSvQPxlOwIBL/aS8vxmdBDU8CYifRYNyB
PomQxjY9s0fR0ii1BZvsLkcNWuRP0lH9QkJFaaEfsOk7ywq7VLVlC9N4C0JZ6xBV
61xZUsJCbPEjUh/z4kQh7sa23XiaAAi9c0UfAtzpqAZ4k7DTud4qIhbMFC8lux94
THEK4CYIrOvU8aMHpvD2vgozF9/UK5c7NEJrYnAFGd14T93ypQXusfjJgtFnQj3M
BCUgZSY35W26gEYLkpUKgkxlI5dNI/SWMSQKW0TjlHBpsQzmaIBiZ/VHQs/hO9/g
WrlI85kX0/F7LOv7+uHtqRVihagHxujanDMi3su6VwqNMoU9MMDAG9+T0DZ7Ze0m
MI1gfksnGbOOd1h2bGZsJqdY30QOt5RNwIMrzpL4BOLBde/51ZXaQXoipIhrocvP
wy3fAmG1QzmDx0We3r4VlKomLysSNnWpLMioWMWaOikum7A3MZMRZqN3ktck3H02
3w7ax4FsPJ97YDOf1PAm4KFj1BsQL4GmgkUtWGjrSK578lZxNRQELtyXe9SjW+ty
Ax64KXemriaqbT4m0bs5gTQSa+k/J/Iux0D8Fr093nt6Xgi6VEwxDop9r09gDZyN
bYcqF+Go8PICPIBcta+RXIKYs7tQNut+dj15GQgvUaZNfLR+mQjMvAMQsgeA6gzq
1BqljhrXx50vZ3kwKjMmXO+igwxgNyPHgm8oQng9ia4RSpvhp866qDyEpSx6CE7P
7pwb7O050BAbe9eGbl12IVDqc7rKHNYKDOLcVQPMmfUf9xBC1ybZ7PW336w+IREI
kDx3UdK0E/jQRCeepHeF/Ztzkndg3EtU79GOsobkGL4ZqfkU6it68dqrhnfAbxuQ
wQOxFLqk8PbSTn1HeJIVmCC6WcTWzQqqn9t/vvipfqrxgIzWKJndbXq/qDv7tgSP
LOwCDp4PZFGwH/63Yr8wJk3eVOuy6rECNYskuALTGB9ONePOqyHLOP2UGVtneuzQ
2ebAKh09LAnoRD+7rRdq1TjvhrBfX26iMfpBB+1db++/iDc7A8Adp+TDWQoon4LX
CCqAb0e47wm635jZYbd1KbvJoLXXBubtBgsURs0bchcVQu/04XoPHhgSuBLOZSMl
rB4Xm8WROBhAWhQZKUJdEwTpnp546F6qVY6xtkGRoxf+EQopx/Uh6SxrABhRaGf4
HmbQ6KFK8FfPYDjVhUrlqpComnnsBrxZ6Q7RW+TIFQVvxFA9qFbV5JYOPC2GRuxx
8COtLt7oIOnm8Sldzy8rBpB8azYNE+hTRHiiKkPJWU6KOfP13y/G38gR01DEr8t0
I55cok+n96oV5kQVoSMcrBVKYUMvqNq/t72iqjJRS8dFGN3wF8Sgji1a+AizTJyK
l9rq4MdF7pAYxVBkQix4QGK7eYPTU2mbYrSeB7Xn0Od5CL9bSMJwEc6WDRRLYlMi
P0yIJEJJmMfxFe1W79ZvEUlMBpRvxYaIFY3QGd5a45kYITRP8OV7JS2z95dHI5L0
pjVGmj9J10rq5PXDxtehi3WymeASMHgkUwNuFZsrmiovkcqMMcUgcCPBLWroR0DR
PvnW7dkdi5lfxuQaBkypviH8QbKVu1tj19dRxHdGj2sViwm0v4fjkhj3h7bOu9/D
OivxX+umumxmHkGkFIIXqFMANds92cc/+qge3pLcnNVzD2YidtftZrWFrKnIFF8+
labreZNIRZEq9OXSbwsw+JgBwtb+cAtngPruXlksW3VWre4mbd7MgWeC1WMiPiPO
LFZHHgMLxAg9m3q8nVKWfGfjygVYrpq2C03m2B/P3GI2cA5vD4c0dFZCSantgc+S
rngzpwcjfEODGElzpIsv20VAWvUWw/xz0c6vU0Vs+rNfkK1rtK4gMtjeKMRUPyoA
zQc4jBxQpxHaxB0FuQdPC7mYNZkhKig8FdBvbyn+5J5rzDtAz+GccDQliRUdBdXR
jy8/UfYg2ju2FNEIwYSzAAw60KBMoDH4K+RkuHLD+Fj1aOy5oBy407zONClDgv5W
oBKNwTditeIjvQWrfZap3FOQ7A1XjINsmG+FmZgF04+gYZEYTAxFq6kmLHT+TuiC
pvwsVudn2TZBtocj7U1GuxZbURq6tn0Z3zGAHnIMpS8mTHcld6m/6L7UN6JL/jvy
1Yd1CGasIgpd013hNuOSpDyy1u74ZjwkLW8u/g/KM6WqX/kqHC5qRZKmhQg5oa3o
ncstvt7Kr37mv4nfX1lzEAq2Bfsa+kZmhvW34+xO0JnJYmvEtB13CI7EtusSGGV5
cQUdYRqtUMBt34FXe3sxFizKEjuAq8kVNjbvPxHXWLG16vvUMHdDIgajIiaapk+U
KuHaRJRtEB12INTHtRO5SiiGJGCxdK5dmATKkyt06Noy6txGIsdusPNqX4x6mnce
YEwT2xML9gllIViqyPRHKF//O23AGp5e+PywnaGvpX8CgVk4IktECmqCoBsrOddN
m1P8PwEclvjlJsIw7yYz40CJCJBhqsWvraIC4oq+tivjETel3ukLz6Xc+h4TdFoV
4lwvudAAP0B9J4mi0iJzGKT4DYEoXB4QNePDxL1cOS62Qm/F4vNRVFK1JNuR0WSg
g9UEL5qIfaKlJio1oH/YOsaG4C0GFQ/V5lMj/hQ5l/VIMXwZCxglMNLTtVGVFAIS
BT/at0uU75y0S2x8dQHECaHVcatkQAv5zb/lpllyW/ilzwFJ8+ogWlDzBST53vXm
g2vALJMqcOh/4cq7dxquXdNAmksK1fpkEXLcVDZ074HLrirc6cp6B1cf7b7ZVzu/
fxU5jasg+eN9CUamy7WS7pn5XuZ4bWAbPIDUrXcSb7kZ4kLiRZBckUYmasUpeYab
U3Penbz7kbBwh/QwnzrSS2Iy1foHFmhfYq+f/iFFDDgg2nBtmQzS3PyGSjK4YYSK
Z+1dLmAAuWCxb1/St4TauFMbJ2M+SxI6hDUKyht+UTXrFOR2O22Kik/Rva+ObenE
NntTMv8SOfrmnBg1XZVyQQjIz2vBUGD3pzREswxi0Z3s8uJkfpXs4Vg0sKITlRuC
EIauSeecIHYz3wGpflYubXCz69MLloZw1Ysz5kvCc1HszG3NbXWskOvLhweD9IJI
hQvXZEgPwt0WjhgUYqPmDUSsrhwID8cziHFg9lA/lsjVmiqAMpApYdiDEaSej05x
QGaN+3hoFfsez2sTiS+pm66vwtMplkK72kuAcsuUMre38HJxvXCHeQMjlkxDRRqh
GKa5cMahX4VH3S3UP4cLn2weX9bTFaNZUU+Flhs9AGuBGUG3qAi6i++1M8+nlIfx
KfRCabGd6foRmmxzU8joJjQwwlyjMBZ33HQfi9KrdAJVuAqVkcQ5T/hFHfdv37EI
+ScAVtoBv8WTXn5HkRNrcskhIjuSaeTItdWNK6VsG/9+crq2x5kc3Cnis0IYzK81
jUVabD3ezrz6thmJ6ZccbC8ZDs+r398X/3O2bFOZ9plhfx3OdH7rWaAhlCiaj301
opcjgdAoCY4PAyLDTBtB362Vl1KWA6OWTOIYVizYHzxleEMGBZUdsl9jzCzRuual
oy5Krlyb9p+XZECAigBs/0UcPOByPnd68JP7ue5tUSU61brLIDOLe8R1HejJdVQ8
zYL8JKNqVwmJmvlT3p6AmHkyqcoz2JEYxgrCRxFbTNZ0vVEJHEP0pRUCv7RkPTUL
9ndIyfqS7/l5eTOPdCdk+6dUhqg3ECjW3+r9cSEfn6AJxMs0Dk2gxZSufq+nt2Qe
T5P+JL/HDLNQ4tvysWwpH37Hy+fNsQCP6VXZVwakFHJjotlXeSGXchpaj9GrwQOd
YskWDmujKWaLqXPekxDeabUjvctpBsFZFMm6lc+re9ZNx1BrFQQ4xi8wpREIDln2
4fY/9zo0usHux9mOpGF/3lSLPKTBJgecmTkFOfZTksZL1NhxrlBfrDnpm2EQeyNJ
QMKaR3U2N0lQjUQmX1feqfiNm27QP68fdIXzQ3yhAJJIgQDBvO1BmabdImbaqSqT
q6NT9uuPv0wM7DVWoE5Nb2bIyoqcP178tHchrZCMO8dLgzEQZA/pwBO7dXPyJiUk
ZeYIDcnmlRt5DOYOhnVtbQ6vHqC659Kzb8kmIssKSld6a9EyfkyKZtuHT6aqaYJ8
luc44bFAhQBXJLuAXt3j4Q7aHuRujV5JIsW+2+P0e7Ipck3h8dAo7ZVJLWGbhk46
x/HOpSkywOWP2DrD3zorvOUOG1OAXf8VuJQGYDmZfZgTu9rGuGtUcPxa8LRRB1rE
44bED3G8smUK9YmgEnTJC1qN9qaBHZ1wOtlug/jJO2Xm0KlNc7+Uk0fkIJFp6cG7
MUU8/M6UqopEmadgV7x1LDhGZ4mp/P7ChbLV4tST6IwlVkm1kewl2cgdE7DfGVvV
g8BNXDHQyMLELbm8CJu/4V1F5iXOq6P8T9TUt/LIGs2LNBj//h7POXbaQOsCaVOt
0WTrmgmRUIjbcMRJuOKTU5VYqhnSwnNg3IsBIAtuKXg1YBVKoLWC4D2kSc35gLX8
AYPdbbJAZdnLKzQWBsSj+MmznRw+fa1Z81R9ACMrimwbCkTiiFIS1XB3GwMXGHAd
19I/Yqi83dcp64AuUxMFJOpxFcao9nRhdJIIUwtgaki0XfRdX9htamNR7oEQMfg5
gQDbbfJzusMIRlPCRKIN5H+SkH3Wsm8klaAMmahd20Hc2ZCfwHqX/VjsRuQvs1lR
l79ntprz9E1UFYEE6UlpuTo/e4oUSRZslLHMf+aszJOMn0M1OED3EsvWWo7Gnf6v
HfsvG28PkQ3c75VkGN/L93c1kpugW6JSi2qIdVwgXMjBehAYe0RS5mip+WXy0rRt
I+e3cCWlTlILf3DAubspwmXaR6zDcGoVENpdIq4LW0kiYQiYAPnAY3g/t5rANu0m
8aWrS8HwhX85B3nN7vx443+bzQCaXFoXoeOQWXnos8/9vplYvZ6uUgOVjr0iRtJS
O+B+jN9giBfJprfl+pcebFd++tqUmNKC63iUrHjWURvvbeO21kc/I0qcydgyCNSt
N4rtwfobHRs6j6kbbIL7h5Mf9zHNK/VsOhHRhJMam7N3kta/3KgWf0/CNPFL+8hR
ku/5i/rhqD2NYrMAwXpd4Fo77EP5xs1oQzwOnILmDJr8RAgo41gVRH66TtYw4rMc
BSKLdgX1/RPYcMqzBuDq3C3wfAHdgax12p5BImGulMH3ibXtheKs+Mm//iBW8/9t
hUtpoiK7zcLlzwz9kgXq01WJ4Upycyg4psEna7iisszEDX6F7kRvsVNnJugO0o7K
oPuRO4SJcc7WbFiTkYUNg8P0as9EeZNKrk48sK9bvzyAPiKciQQIdlC8+4Fi5fEL
D84i3zlZmQ8tPQNzACr4eDjWPk6p5uLLBXJceYd+do+c9x09GvJ2tR8NzrcCU41Z
spFyuJyN2AOUcNJ8lIiivdlt6qEHwo1ypXRc69hNveSPd6R6afb7VNkZBMAn7827
1SZWo4QCarcOh51LvLyT2hjk5Es3wIgDo7v+8dodnE49bh0Vqlf/CGi+nHVgtHTd
xs0u/iSr0dAzbNXvCqnYM/auMZTAVKLJTJ7xKnOCpYKNVTdmlTbRQNfFGkEFpnhy
D0rjd8yGvda/TVl/vNwhGVSPmhX5hN+PCdUMpJVPvCa8fKUSrxlvC3i1WB05TMVr
KrxXM1hQo+C3FPmJCa6gnXhNJZKjbbG+PpRvL9/MRaTG195stI6gOQCfWSqCkOfq
oH5JyhSu0GPSwcGm3zznbL0W1H1vCKs3T+mvKB7PbuRZ3dzl70dql5BESW6B7tIg
TfmWKHZDIx0JyeV2EZHRNjKRx3eXdW9Ga7C/kmJ4J58hgE5lEMflpLS5YPTenqiW
Qa7grAnlrmKKnpFkkglOhljXQF4pstQspWt4t3lqE2fEni2f9P16uitmiqVE3Kj9
yCErSRiZ1NrRgv+iYx/fO8XD/S2sVHZbIeCL7xMl6lCTHdGOvg/DIZFXLMRO1pVV
baga60I5K7iffZbfBqoY7Gg0nOqp7LKzWirRb+i12kktmmqjpsQALBuopOTjxXjD
IPjm+l1037xTHim/tNEf8kbHP0XD0+2Xge5mxXmp73q3nlr4rXYLL/cboWcEmMW8
tX11A+qL3BXxbZSPBEnYspc6+GCabjYZbVutv+c6+yODsohJiEhp9MbDUo5Uxs+7
JZsuLiW5QFn1O+I1rTwklOFsDEL+aTNwZ/8WMjYk7gC/spJsLqiaVl7W1mNZB9tw
fhr94PMrVHkVVlAt0pundeOuHCad381l2Bh9Xues49aS+H/Fycaj7bql45kqYtca
0NAmev1fuhHybyjw06rvCnow3HIhPDx9yhrA4Xr8PYKOAf+0vOgSxDYDsPkDs4ou
ez6h/uEVoX5j3oreQLVx1+CKjGzXeovtGMqlF/14snES7h1DVjfjiB8oeJ5/C4aU
wjygNP0a37GcjyK7VxXHKZGtmXeAea2+wPK0QB4M2XZup6Y9o42D1FJU0rnpYW7n
FeHkddlahjXsAb4u87EFxDegUWaFnEiy8rJW8Ig8K/hA4cVcVz/GPhcxVa35Y71y
7uzeGvDS097a85t2YFTF8aVgQac1Fuq2H0L/wQV1HkSvwoLEzUGDvL1srEPYH/K6
7XoJwazqEZBXxhiJ47zfKnsBu4wY5+XjyNHbbBCBi8IKXLsB71cLokFQhv8xY/mJ
EfVHXkMsAWGIPazjU2gMKVkDXhY3AjEZULriXD2OHH6iqBARZyY1mVSUys7eQTRI
oH7Mxr1ZTQqB7Fp291twXjw4XU1pnzAyncba0Ou+YhDORsuez37+BCtH+FKae8GG
bc2LQvpyDhv6rCWewdppHPJ0s5XcZm0TlTs8fXkHcnwaVZv8A5YJeyi3GGxb/R2R
I3x39gs8d6rAXLuuG7S+/XQclQn4zZUpGFiBnmvfx4bk19PM7DCNqrfcvXx2h98+
wVDh8+BMruHv/FiOMNBfD9Ho7uVws1QuxeeK9SaeKKmUL2Yp1XOLJzPA/VLKOolV
AQPO5ORG4Nv/ezH9Kf2DF0LZEaFW3bOvfiEbUWQppT+vDTTDkO7gtf9MGttQkyY/
KjvNbqngTSHJRAgJAuDiQmNHjvYIT4XABg1PeSzOZD4oCg2Em2loaPjYcENkLab2
mGzPXKKyjO08XNnL9KUNPdcGj5oUUni6XscFcj7DEuyyxDiSBDDeEiv/6sZhmNqT
artjLuhoWzxUPHDCkrKfZpIHqv4jVisxiI2vb4j+8LeykEzivmnDA6vamrUjABHw
ur+CKjbli/mWhB3sV80OvWEiuTupSHcLC0Arrjg957y+PwZMvn6zGZ4szX9l4s6B
YAKAs/P0JlSBP8bakNZLfh4XMZzDV+D5KIFj5iELFLlMSN3zEbC4VC/0XY9ZAtuB
oQkQGcrzopps28uD9xXDq0a/403IJpjXgFnSMMkgkxkwKfytD9eEqNjU1ME4M6Gb
WzvrNiopVIzMpKhgftW7jLWDlLUPFocKp06+fO0zF5fbzU4FEoXZmWhOKBS3OzwP
kiSpU6I/64eWgMJqX26Vi0dqxj3NnTyAJH1MplNaGuxhxKlE3gCPF0XF8hFjcyH5
K9K2vT9fWRTzm8PrR0/jXy/UIDZVaas2DfdE+hlCZmcEiLCoya40nqbvqKm/4ZwC
d1vLZ/uoBSwu91GMWNTvo5cpXfv7BF//cpYQ8cQrTebMiYK1wwnGQ4vTIretvQkR
fauizITvf9SXBdwFKAw6TlBhwnL70iS5HlXP8F5Vy1FjKxJYu1QqM2SEqTME/7fE
2ChWYdyy7ZlRlKLRC975eStYezUirOxkFLNGy3+x5Hfz2oVxHL0wm3bMIqC4r+E0
W4Zc0ZD4/DmELdlgzV6J7iR5hZo8q4brsv+n5ScmUeDev1OJiz8NObaWoeQd7oAM
ZIApv1EzF45GXo4NEnZLHIU6GE5VLVWaqP+qJCMRJXLlemrVMj6HWKNxSHiJABgl
vljG3TOhF8Y7M/VIcD/wKfNc6PQVUj28iTcKcvoTyGkKq7ZizM6jqquVrD3VzS+x
pKs1KksHxShe7L9JGNDL+d+yZWShYf8i2+FmgmjwyBqR3yJt/0VAjLX+ViKEgswA
lnkUiAt2MBYXx/kLiVDIsYNMN7YqH+IBB6SkHus6lcTOwLi5IJ9VjxHq/Kbt+HDY
I3zilNYgymMeyla6jSL51bZVx8c4SB5X/R6DPnDI/afcgP+lbEmVDcer8TFZ9nza
ylohZVL6vrjmS91SIRupoPGILlfUuNbv6LRrdTtu9f1xb9lBd0BRs+sEfyEmrHMO
9Pw1HXKsXw9Z069tlpdlLjP6M4RmMqEwdCvf6wQIDON4r49W2MojMB4PC4Sy/nQj
Pg6udLClyyOpkMetjhbOB/KegkqSjA30fKJXIKU1aHfQaQxAja/Wy9qxBwjHxt6z
hRdV0OCXORqIkmPDAb1On8lybXv897FuwHW+V2Bp/u+2Be6eLU1F0bouEoo8MfTs
a1CzoMUuidzGg3Xgz3GApJrHGtqXfFW2TshJ8stfSnExtn7dfvosHzyJ4Vu1rwmo
8TINzj2+we9tjqA4At+1c1yKjbkwmOQDQr7ZViXN0xO2BqHZiyBHGgcndzUEHV3b
22+d5BckNjKxUTfyODTv6v4ybxvsn757hteCPRYgW26mO98NjslGO6qSvalhBfcE
EeX9Tg/gVyYDwUk2ld3NcSmT2hC38GVKtdcsbEh5nyM9IgITTgdv5SSJcVm8CPrd
JaorQAY+Y9lLdWtjImE+mC6G/m/jWnLAHnk6sfOpwXjHogBhmJsDmJ2r1KH/pHtf
mNLiM9swo/9DM0OlqDi8d5uXaG6ZAQIjkyY/ouApZYIcWEeDBwC7eHDytlpwSH80
NLU32gvrkCb8QTRCW/PATa5vKOvSqlgJDlhNEQY6SFN4qhZPTAyPLEG9nIfxq8nX
8c9ImdP7zY2+238dduwmCev3piyn4g53gILXR9Nt6UW3JA+xhY9XwXmfY1ZFkK71
OR1wTSONjgtCEg4+T0cPzEgTpJRUolDW31amwPVCVKaJx/+liO7mkjJA3EUvr3vI
+cMnX4vikDmicCSax1Za0FbREGl+WpcB5UDwCH+3H8miFbnmy/rcpklOtA800NGK
fu0X37Kfkcl4evCKk3rXfEKQOMepC0qzBfXNEeQM1wxAwybO9k+1a1azRzzq+EpJ
+KmDiO4RNwghQPLw8WJKP8Yu4qcIcMH1tsJrrAsRYOGZHXDMSuht68wJS9hLMRhp
jtPwu0UaSzVNVBISZtfIVOVOQln3L65QvdzrCO3ImLG2bmdVtY7WuXQi7z5ns5M0
4GvKWeRkq09PhinyFmdwMiU/XBrOIbz9jP0N94o7XGORunNQ8w2Wk6xZZfNyL9Sc
MBvmOb/ivrIgUdpY5ISFFKG9cT8mcThd2N0efj90EOovQqKSO33rW1S5M4PIhfIH
PiHcMMKflmdo6TDIpSsyi5IOqa5+kGIfY6f44MMBJECHFBZYfe88w4fYbCs1fiGn
7JZJyEF4Yc0bAfMLMAxGws8rX9ZuyuOrBj5x6gtquQb6t+MiIVYmNeMbqNRc95+2
/sFF0uqYMyrjg2emKS1nN+KWR7LQ0bNlmguZkkMZg1rXbRo4A0HGnNbrdibADDH0
RYbRuw1EsjzwuWRKa+UhC0gMhqOdLEEVRA3SyVxYuZrGOT6wiemDHdIe8PoEwe+R
2GywbQJ1QGwt5qROZvF1y1gdK8W6375mcqlbqzlU+9wIMKR+JkhqrLpBkKfKAHZb
KpsoyGt2hQtY9G2m2ySwAi9gH4ug2AEbsxE8LQb7k00ybhnOX6soiy4TEVep0zJz
vIt9L+AAeEhnSFCoEhShu489alTGBmaWGP+R6chPuK6MwCzzD1DpWXTB6aX+6nOm
4JyJIU5AdAieo1xDvS7ZCJk6UI1nlJ/T+IxOEYkAbJurV2zAQb9EjeeJeQs9tFD2
XuuTMmQcRcwW68Wny7DBEqL71Ri4xA8T6sD5w5PqSby0uqVw4cFC6IpvfHg0+XZY
z6xB99FPohPbn+H1nbdbVZkSmo+HA8wn1b2T95yuwRw4uiZ0Q13whGmerZ4AgSil
oL7VS3X1HE4AvVdfbIZEgTVolLwxF2ecNg1NwjTIwRDIL/yXOZ+DNOV95jT0wjDg
7R/RPItTkek7OAQFpAfEy91RQXbY2YJ8YhrRNH5vPx707eygkZU5hGNmi7wPXSwk
XhPnN/cTl2hEdUxEV3Yi0dOr3kNKqQSE9To1PaWPbPBXPL5Y+bhYWWEF6Nh2Tpli
WUqi+kUOetia+3ngCCU5jdFQI1ZUoMASU53fLCM7REnnUABoE+7FBYaQZ6jDlvoO
cjwkCKTQBnI4zbp+uLNys8wWXBmCZhptSdhZJzlpCxEJRkEQJzyd7RP1TZJBU4n4
dOk5awknEYSfAQox4u84q7c0eCc8yaG2pscx5irZown/IPuqSL4Mgl6MEkq1vdwo
uDyIHaG1VGrHMzKzZv5m6mE07uxzDLb5TxYWyhuTelaIQpG6nd+ttjnxHe8Cwx0N
qX87FC/iXzen6FKMWWY53mMAFtzYw1GiyeRaMy6/F2cmq5adA+dcBKPCWSaLgIIw
R8KyM4nXjeSgwiNF2UT3/YzBft+JZUys/x4IhgLF0+sQiLCi4PrOwJ6DOHXV5ejZ
/OKoXb7gx+ZYpw+3xmWjs5lWVYa1RBqMRqYROujwhDyapfK8Us8gLwqVSA1Tq3tb
BBsPRWDw/kBTKuG1DHgyXBG5ggHfQ4tFYoHnNitla74nuBhJA7+Xia7baInz+r8B
TjFL5LylOW02EQ6tcNuQdU2bhHSdHCXZcJr1caFrN9Wa5EBSC8hmn8OBqa7AHzV1
ICpgBMEjZW2xfvlTUU5/8Dc9/5JiJ1ikTpkbG2tV+U6F5DCPERNgAy5neBy8B39x
JxH1D9y6Yh+sWWA02qVmZUHfdy3t2q82p9Q1PVIjbIWMDgTT2c3YYZVvxcMHvipd
ezJdio0qDhRlJJZLS/A4emRvsdjf50IXvGMgUE/rNLQaoTILGE/Jwz1q53BeJqY9
XF3fKyC51ozmuZZArnuo/WGi9NjTrBbqwUi0RVzMI8XPrPHI6iNE7qdwTt2iI84+
ozpBhCpEDXVHtecKD4NFvmh+0Crifo+EfPQQmdyKiQEOZzBZZodclknz/vs4qzyH
Kp0pVxm5aXDC61xGy14XpQVPSGolo9vhOcOaTCv9RRVb5PQIlBi4mXJnRwB8gbDv
AJeJqCvTftez1s53FDeqUl9rtrsu0nR13DRuaLDdxATXFAhiVOuuf8qI3zoW200Q
euvxcoV/+53rpwLUrpKav3GD8gEpWDB7Ag8Fvw6Zh6r34kvrUfOZIEg+5JC9mIa6
UyaKqIz1pRreYChjaAkWbQ25XN7+rs42+h6plFxcqVNn78nNSlVJQojd5HDmS4qd
ghHobRTFrCHXqRNcnZYalkaQjqXLcxElNgMTaZU7eiB45HV1ANg0O+CG/1jaSvGs
FVmTsRz+p+imc5z1SJhmebph1g3XKyhMs5yXY8fKIkw+WHIvqL2HQHNna2TN31X7
O5BeIrTQv4kyKmUzZ9zowlSkqDAAkjlzyFagxjei/UTPfMT3U4Sk4uFKcDUbZwT6
xsV+QEAGtJDu9z5cOgsWz2mRXBgYuMp4hWqM8aYXMQ43GEIIyGPXH1KjJK1aBm/h
F/xZm3OYSBCW8jFD8+OgrCgqCBSGXKVQZaRGIAnCl+xv441PP42lbeahYNt7VH5h
rayh5TJWMpLb82q9zY3l0v8+jJt4vxaof1EtWiTSEajnAs9iL7xmjHMv+dnsTKH3
ZWIL8C5yVklcQS63+1PddPb8vdqEBgrEGQ/ov1UEC54SENGyVGyBYkYfjnhNqVHj
JUYQVpStFUnSvYCtCv7JY2Snsq7vRmT7fsvha++L5ipIBjGmi5vmYIMLNLTqpEJo
DQoKvIzt/uOpoAZojgUfM51ts9H+/QrA0vdQi+PEfxkDGTAGxiJvhhhyjqhaYEdq
Xc+BeKaWtJk7eA00dKEE0MQR23cbR5sNNcTVAv9z/SFWsIzlTvvrChVU6B5O8fA9
0JSbSDx/UXltkzdL1+As1FaAM5W/2KhG5YvDpi8NYL15uhZ8SWiaLrN09TssXZN2
Y7BIYCuLIVAroTgqGhUP4FeV8QD9nJR17PsKYooTBcWHymHJUpe0CMA/+ltBFjGc
rgQ4NklBO/yFzjOyrgebSqt9WrEVDQ7DbaAHTc5rU3/4Ft9qfn6vwWl2JWdLzg8n
f1El1O+oe4QefrzzNWpX3OoQW7XC8FZn/zz6KxWfjgVmo5y+Ka32qrH++EqTrslF
308BWklkI30vnPW0t3qliB+wfrJLzXSlaxpWULeH7PYwRyYVGQfI8epcxKYylZ1X
D2fIjhDvtT+9BYP5XjxXNo6+idu1m/twbffFVD7CdcNdjkDZWHMNm3swjd9CiGzT
AzXBjanh06IddL9qX6rwf3h48h+aLlFIImGuZMxYIg+nFmaxHUPzczcSMMPzXr8d
LsXHSuCZV5WP+QICgBYvYak7jc8hn12i9blVYj+A1Sd76IeSNMcJnvqmjsJeVG4G
y3V83NFOtHR2RZsW9sRFtf91HtldPEuIgK+w2YnwnG7uMl++EW0EsWLxEjbYzozs
5+8EBA6sEZo7LguUgEXXPemIq2AT3nbfvOWce+dXNqnfPEvTXl++qBBKMqWPL3P8
gnAQPgZ66BopY2PaaFw5wtJ9OSA2o1J2+qIxuJufJpM3H7a8B7bLgfLwibgQM9Y+
z+lHBuJM0PKGMekc2oODq+66BZeE7VYOHVlc3zCLAOw1JqP3Vd34QpEUuOI/T79p
PefdnL+Zgpz5QfT0cyur3LRdc4ewgWio8TfsYwbC6Ff9mc7zPwMiWZe5qn1VJk+N
TAAY7v9xyyc9XRe2BwmUrd2rU6d7gXnstUtrinmpoQQrUGlY8cRpPJHKoR+7wZU+
Nxv31NAi9xFLC0Jtw7M21SUDL6e1ENyeCEM8qA1o9qfh4rM3wRlgxJjPOQTh9Q6g
Rn9W6k5ZIhZzIRxvMi77Ss7U0hzrIM/g+G4AGuGqjRjSZGT0gTMnhDexOUJSjXjw
IlqBioTfMYLnj0UR+36bWnPhtsEFwhjicZbKcDYO/RK4Pn121bxu0eXwRMvB55UT
Wcvs28102JfKz15LbS656GvAS52hImxOqfIOYosRMChlyd8urM3Y6Hcfvhr/8Hsk
V2iV4ekjwpIpyICd6YWwosRabbW+E5E04ivMJBxKZbvE3mGOaD7IoFXLyu/KPGz0
PCbRT4oQno9WnVxXFHJ/qyuJBKtbqgwyxVPjrmEmcbMz512OVQnTIVn5TVNvwRco
1jx0f7D33+MkzUu8mxchAlWM0sgVkbtfosUFM+qIdBKwa3oOaJ7gQb8FL/CN9zfc
o0t3YD6Oxie7GytHkCrQm1bW//sjDWpGxpVpmeYZzkGTe7I0Us63rk1DqheYSEbo
ZyNTr/WJFUN6U6bKcd5UgHrtp9C832sEn3iXKaviYyRsgpttFxK8VZ1NX1I2McCK
f7/qxfv/clg3hADPkRIOZgwRMPVidFjquHVpd14OopVinqzagsuXe4uJhXNB8RSY
xyfhdToANDhxdQJJ6sGcCcfOr2DqQdEzqqjCBz4T0l7Xhn9GqzWIDi+d4WcaKsuh
ZtY7s/iGNCI/0n9SiFRfC+bhICd8fct5ImJk3Zvzx33dWBT0A73qC6L2oyx0CiFf
BxU+sqSPOk4H7Tu0p9cKqsJLyzaYNn1J/635sMfLH5U5PW0t6znIn4iBs2UI8XX2
4G0/0nvuHNi+ioifabhjj9oPNGFPQVtv4QVrmusN4C6hpEzha+AmvVddbjumcU8F
zp8THQorIxSw5lLdUkL+5Gjb+kIxObcRbNS5C9t+A2OJW1hRs1L2/uXdDKZIffyH
w8VdLQu8mVfRX7qR2El/YF1mVU7CwFE8SBR9Bd51fh/C97hGpWPS92u+lVNar3Aq
vWguRmr4Q/hJWYFVHNsMm+dyN6Cndzvtke0bHpjemzY+AZGMezHH5Xx5LDlTku05
XEJu5vB1h1agC/Zq51b2VqsOluHFVNuCR2v8XvvJFozJFDgfoHZJt5N6AM1TF1F+
WsHKMON35jDooHOAXatUinlsPzTVA+bkg+421MU4zmj6xkEgG+fXKcG9f/X+RhdO
PaklGFuXpZlDt4couEgq1duuvyLCwHFvfaPeCrgeIfxu/IAxEznMShINXGu7oi1F
ejYEW6EbgdmkEnBy3FtEGPqiY0mFNHDQp0DqXlN/we2/jRuwJo+QcUVuelCZ9Rt/
BK+NxO9OU47jAh5dF0Hw4H5ErAU5X5PRWBPxpP8wefE5EdjPdOrjjGXcLwMHwIws
o805uWdqIyRVymMhXOtSwx6KfqHqwW76xYaQoMkcLboeA5W2sQ7NNug0a0b7DYnr
Js13N7vcxC5tN25toucl5ZE6tMY5LT3x9WfCzQSSES73XQFy/+9J/MBj+WsZw9/7
IdJjWcshIbT+mQYKtSVv88E3XPWVCKBhZu2FuXYx1aXWlHTK8osnbEkyTR/fdgiG
BC9dFdJp1GkrsuYC1O9ojhi/3knoFWA3l67M4U2mEqX6VhD8anoOftaqXPhQ2V/2
Ivaj94IjrJcd2+Jfi5p8xg5CRls7w6X1kfzXD/yGAfgfP4ZpYrEN9f/x/ZTmqEVi
ganTOzdMm8aYZrKk8L9/s9Qo7D00tySD9nYnH1LP06rB2TbihV8XDOzFivvDIQYH
RTLDSA/0g3zA4jMrQ+7gQhA0QCaAzaoh+xqIZwJPEHXoHdjlUV+Jup3A5gmjU00m
lzioG3f7p83TXVZ/WPO3iCFy7RGAF/pj2B+VeyY7sU+MOywU7DqO6e0aVglO+eE1
k3s6lOaoXaK/7Bds6C84EYDaIhPwPfgZoNxsK4wc7wLINOHSFkIKK3vVTCF7EH2B
L+UWCyHq8dIi2PytVpGF+4QQrLdAwI72ZmLlRsj7qPaCtXgjNvfhJa6TAg+iEEPa
RAWTQuLzYCcxGBLNM6BqNXAV597saLJFMjxMpdriF3e7fIbSIjEVyzUCmqhVr+uu
vwJRD91sPyNSLGsqJx74lYJXZmQs9WNjfYwZibvmf4FisOMp5OSe+k/sxruNc7L4
hbPEPFSn01j3LYGydG0Z+A1Wwie/kvZaIbzr7SfIgp6kYrNdVBAhDQ5OGud3tzJY
zO6t1Tqg3hiJ+dEhCXNh9FZcF16E+fcWOjlP9D3+phe42DD7F17hpAK4RDTqmZ63
hg539sliOkQpR72RMT2kliqudalh3QcGq0Y9d02EVM678epbJblKtYTQlKg2tew7
whyLXj44Ie6xOL1WGEpCLH66Y2BT/a8Zqsfn9TOUsScQizCruyGokKouP6rFa+JT
ok+CMVYbFcwtQQCqNaySwcRDxyVTEqDucyp9WnaurCQwIFq8TUsMl/tXSiVAPgAX
nutdH5aSMAM8u/2l1GhZRpQtQ6+y/JO3aOr4fWGcTdoQ9uA2XMg9OiuKjRrLT6a1
+7lQm1XUCsM1LyT/D389+j2aEKQ23JCRlyeyLA2/JgAgbEsrYRMVbkRBWFKdAfl/
OfVyMF9Mdmpad+bx6sBEd0M8nDy71ZnLtP29UDEM7X0WQzzy0wbNRRYfJyqq6PFm
hJ6u/wHWkUZmohr3URRwLDxyvg4hbCeTyh5VyqvQvJTQCJbnmm6kLW8onGBHhqjg
ZwEU/MNVMOWXQvq93jqnkariQDUZRvx/dfjjiLDKsVKRvKrkw6Tv2QsLpyBDbgM1
vVN+q61zbOHJ+c3azBehUtfW/0E1BctdlySVnxM9sc6QWx3Lef9rr17n1AesY5RY
KSSKXEkqY73cJa0wd0MHnZtfVXwUiv0Aj2uF31C6lCs8PY6jfC6v0lAE+KwhmKHQ
EECFyHUnsrhXD8eVAWDJX3tqKThcjTW8WtfG4FtF7feqXZlg9PPxrGk9RQa+g6ex
M4VGqmnBZ+afVuUZKD6z2k0FNbNvFcrjRybxOBhGELvYrTaXYiRzT+dfpeHeUl8A
44OJN5sJQ93Y8YyLZtYfrarcN05OARsBj43cZYTdygtzDA7jZ02kvVUk915WW0+u
WG1JbhiXlzj55gHG5uH/mvdKCIpzmTWYIG84wAWDEfdnu5c68tm5NdZlaGVg4MEP
TYeEm4P14SgBtzmVDr/261CBX6BCBRm1S0ebYLF3oPLgnX9anymAwdp8cxOF2YSq
CFWuoo5HW4nXEU02q5uvR908qGlVwKqF81zBk9OEM+CRQAUZkFFXK/BXJUFm4jif
bmyLyLp78cpQjfY2jtVr32TKN/6a6QS8QsegxxXJwHU6GD407O3pkWScOQm4jhuz
5EJJJiUeVn/tfm28W2s8QetlISWwh4bPleBGY6KcWB6NgXS+Y4INeSb4RcpND/C4
XCwUmIXeOvqtASqohtBLXiN3zFF+USnzw9+yfpTAZbzYLEIJ14O6/PeZ6hb01czV
uz+OjQ+mbo1sgyY9NT66LMVGTRLsCVzIcqwVpGziNhFFYMajSMHwo8G1PimqCy4P
0BoqEqNgTO3nCo8QJxrR/ILX7ZSdHPjHKO+KfobxCJLbrCVxvd76aiKvHSBVtcAD
VayriuGsrqIlDPgS4H7SAuUv4E8s2y07DPLn5WY/JS0sOcSE1sHwiFA3ecCt2x0N
XVmpupAol3E0Mq0hp4XtQZUtvtVN0KUbE7WvNS/Q261OKeElc41rzNdASuC0dOLk
pAVxzPT8krNWXu2teOYGH0ZGxh8YWydL949hAFCQTSjIDEn2nfEAfYI1Sxax6PI5
0sPNwJ3vp7gWH67VdWiU3Cr7Um90Vb/hYRmt7TaBu/V/AcrrMTQPAGGFDslxhv+L
QxwO+85MMLh6M1GMOm2fFQtbTfjuYNgOGJQGOVNJ+j0Fkgypnmz8fp8Jqnw1Mc48
TLoQJ3wQCILBoZo77Fsb5fo4oQhOilYjQ6kk1f6DfgioMsA0Fn/l+8ZRikBVYY87
HRbE2NSrKYyppl6xP2FGn0ibR+1WJoFdrIjxwALY2uqxfx9xEKzYrLDZAmBQBTDE
XD7EO0miEnKI3xlRY+M9VXKA6CSHS+0Bf4eNZk+8aRPD9i3XdSXTHMlKlkJhVlrL
66I17c/6U9qHtd+Jui4Vk1wXwuKm8u9P4NaeFPy0xx2vcDONL1GUaocDtOuGw6Nx
8pc+UNdyVRhqyrM60Zq5Xyqzsr5nOpRkCvyxElSQYPHy6cEnetgQZTPcATJFHPB3
nHYxhrxZiYjRzrD7thXmTk7+NZ8PRykWR/ipKJabBupqc/MSLGPpasxoaEC4pEV6
/yOfw0Zzp5nHKxbSa4LtFgzk144TgbNg5YUO50YG9zX6RbqdXetEXQ2w8kGU+YOu
JwnMFyp7zzjv5sXtBvJojWyhO+6xaAyB+xKjrquNgq7EqMsgzSkldOcizS4fLv0a
8Mj966ifiWiJ30wDWXrLbMdu5AT1gP5puOC1mReMxcq52/Ox01YcpHB9rPCHAhUE
aO/Kp+cJQVxqdQBOyHq+7bsNH4CvvUd5stghr4gNiyAGaaw/mg6DfiDdTeafgRiL
htQO8N79JOir5bOgvwBf+xwC++YSlz8VdJTH21OIpdymF5y9jhrtBcpzWnZvu8fY
`protect END_PROTECTED
