`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxjv3HoD5sddz407G03zsT9HSNWEjwhraGn0F8ZEYfg3shPqmZfs2sZkndjSf4rm
efJ2Mc2TRrU7eSGpUfHcw5Ffd9t8MlyiMyDTyvfuSxxcyn77yjPplxIr4pBTEqne
RhBmFkhhE9m6BaPCCO3/ZBJ6IKsGo1POdQLHmsuaCPofEq9b+ATUR+hgBYRVVp1X
Md1t655xgEUpyeW07Z3czdsopDQJ7PAE925Vt2U0MmFOdNNF85eM1gagV6mtp6kX
rQ3WDodDmfpd0VFAK9oVYJb42oQkJNx6I50Bzz0zPkFdUP2CrUwlm8NvLtyJ5scK
uctYrznaXJ8ATS8VM6sLLjgkiYg2OMbsTQG2aAYPnB7TDFNkBk6kdA4ESQ9EgOh3
nTM3U4AMFrPxJraZckaenfMPizBrsWq58NSo0Roz0sYeExVfz+CW8y9cr5wn0UNX
+ED8AyTwRz0OaJbMgMqRuzpIoTVgTKmmYr4yDF/7LWCMn4FAUZD6YPzEvhFl9h3g
ginrlUngxo5DXlAm7vIjfzhXpX+jby18WCrd/Il8pD+hMpNynO8SpY19GX1GTAa6
ib1EMxCCyZInPfRdSAxJaDHo+UQpDLmJSmduH5OTtTSuwsN5T8+0sSiDpmnax5cY
LZyfy7i+CTgu+ShcLNUZ8AbR4k5wVMcYVlw7WFlcNCzvzjhDnwTrKTFkJSAMFzQE
cAithGL3JO3XaNH1i8VgOr/K0WH8XynS3dhCKyiuvDoVzOm+FHtgK6nOXJnNq3o1
BC1WYt7br4RGcVUeDyeD/YfACDZko1UuiC24MDDXtmag7kjSo38owonfLeQsOteZ
8ZXcKK7isNXAVv/KDkC/u1ZV7ibPGNPYMrLZCyDHeyyAfyRWpUHXl+tIAU/4zBvw
A9xRavXUKFeUWPYRhAYd1obhR7u55fo3ohD5Wn3iiz/BZLZTLIBUcmqxbc0yFy1W
dv5bYh+PBOXQK4nB8Fsu8lJ/RsQRhKMde46QoCNDDt5NAG40EG/VYiAWLRioPRol
cbkccXVy6o1oiAgmvtaKLt/eR4k3vRJ/yYsP/pJt8SahV00QvqVNY6WNEjuadwVd
jrkDjjIRWRL5Re2QUrFcqdtFGE5ZChDQMG9ImVHx0ssVf6l13QridcHlJqNPJsN7
l4uF+yVCj8GKCnHPxQu2vTfdSrORFfu7hRKGw4RxiKbFsuFFAOaEuk3cCHPZaRNF
V8dk4pfRYqz3hC5hNw0+z9cSQ458XZpsahZkDyoPImDApYw6arBKtwrictCiTHLo
pc4nlsoW3FVRrxF1JxGS0W1FcstDZBG+Ubhg7iwXki6y0hX3kRS/vJVUOM8ap53y
UfXgzHrGwIo6LGXTmsvCtVRcRzH36KTAOE/8quI3RMkpm0xm6Tl/d7sZ6jzH5WG5
QScnraRf12WUobLo7Mnm9ByZ5NqxeEbDwkfcdiMFsnKExSYBCL29N1L2SSJ3dZa5
rc/RbesK8aTh1LxzFBHKWjOdJ8Zb536NezTOOEXAlQsHOUxpd0XbsyNfFrxOtEiV
E7QUHEmid98D1t99AphUphupm46yWEqx2/lgqIygk/7PrkbQcg26WkQNBBaBbrnN
6RzM56YfK4OZBcl/s/vciakc8BwGVpVmM84Jt5yUhjUmlSXLbK0TamwMKIbOLsoB
ILBoK45TGKYYW6jhT24R3JktG+w37O6URC/COXXBPXvRY2UVplhE7NKHDpcPvpri
vp2yFxfL+VjkHrOzbES7sBcqs/GMUVaMqj6rrF4hgEFIODKVXoe6ha0aMHyWUAwL
/ObEB/pKiOZbM8AqouJ7qASdhM5NNWTWM3GqHFUHALXDhq+vb2sTNk0bl068rT8W
0wr6RR7G6FWdmqUjp9P3C5nba9vbBfMyBwj4soQwjxvc2SddwigkOXcseom8A2fn
9ftPKSbxIiA6EET9YqqKPikM+CXjzaxhtIWMmz67nXZeWDFe8Gi4gk+XdbTPjylj
ZDSRdtJcXYLQIzy+SlsGTqUP1H5NgFDD24gv9geJrcMuovIbUOwVc7pHTyuocRqQ
0Ft6WtNW1T+FzgnhwKOXoc4Pyo/NF9H9I/ytSsR8oc7ZLr0FsHd8PQEXN/iikif2
cI+VMj7SmTM9lQ/zFovysX66VoqdhnLmsI62wfUt5KKvAYxbAgvOrPMM7AlMsX7m
ZFsGq7SCrHri4kmC9vYtgstsL84B2bvTZ7grLpHJvc/z23qHPAHWTM5WIckVlWek
ROO1oeQSEM03QKAZIEgFHBXdNzJ4YzxDs/tXOVnJK3omiSrg04JpOSCWu37AlEgt
18QjAFhOTpJG27T5NiM8IRRny6yLAc8UyJTLWtWeROotYf81ExoBTvuk+0ffDhgZ
RhI+o5kQtA1z/zYA/wN9jrNdPCybG7+YwxojTpzv10UGy2RW4x0j9SXOqjBooezy
2bB9osb5BYPEsXjoadJfb7UtZiiDaYr9N8AC72nnZ5QbPfLWXPfNthKRXB1t80IF
8MdkT5Y74YU8eeFEN6bYNqy71VaWJcIfzle/B95Y5yR2YRed0JJM1ZhZBoSpPj37
Yx+FOdHGijMQ6AuMW/fzKlmvqVXwmBrd9JwOC1V4ZBYyh1XW4+wKFTdWhoIyEeDx
OhRhaAIJ5YVOacJw20lZ3bK0otdpKZtlEp9Oi/7eUhqKff/BjvPxlUCmx3i3Ii3f
0QBdLkKZet3p4VtGwpA2V0ZDuRLynJCM6+bfIHYFp9sZ5WfXwX2wTy6oVAAoPjmG
768D/0j8RhfMDw7y0N7LVcg7VHbRQqrxCInYthl0ou9KDrLnu5P6cSMbuO9hz36Y
Yo3RKo1emGW+DQ8jf+5Tdcy3v/0sS7adBvyyk38cDKm0A7E/W9ccuYBb8ryru+nw
1aTxQnmFC+zYwxFe32ludLfOGyeb/k1W/JWSymjrjv4vCv7Hl8nF7WLHvevb6IE0
2Q5Y0MyWssd1AfvQqSb/UxV6g306Ve4VpIzhl8b4LBxePgFUoOtP3vV4BioWlFJg
TfVhQKL06c/3LVgHpBVcNzlfSnDYIVC0hXgb5RKaEy7jYTxkWcEhzfstylojFlaq
CnzwoP0rmgN/+4OeEKSq2lffS6NmgLWZwxbsVz+uHqs/ieyfeY6k6CIEWA/Re06m
l2VDBYIU4RkKoVHmlGeMHRy2b6JYNzE4/rsw6/aCff1x1HM8lvYFFKzQtPXDYxW/
8KIiM550l23+rxm+oTe2vu+CkilqaoqLxEHkz4NE75c5TOaDeLcQpcwgQYSMAX89
lOjDECA6qUCTvxezDMsqm4qf/a1G9f4DDcGXgM8NrhKPCq/g+4DIzFn8eWz1CiFr
yZboQRSV5tmOWNHXvvdx3diaYWv1DJ3HTrpI3HFZDTPW00YWvydUfiAac0UB1Z07
SUnBcAzOwi92Uara2iBOFmrfUJRXjtZsJDBsYm8S/FA4NWRne2rKOrks/Lt8Yx06
xx9RC3/RDuFxdUAV4BRaDXAgk3dwA/GRDcvjfF28/9OswXy9LPR6sOv+WVDLeCzu
KmxOO1A0QJ9EpwPGlQzv3ZxYAK+0CKG7bwKf5NZgAslmdLGgNc6B742zkJkh4FHE
dhjr55l2f9zY6ErGlwBNCibRKuYXy+JsIg6kbCfvio50GhI13n6S0HtixgX0iJg2
IyxAEY7uWqWmizOIn+0FXjABLMJTygEfSAvEChigAnGEqp7FRce/hAOscJouZS+7
mSoIgOo/gB+zPHWvX5rgoruj5fjHN7/EXvPu91JIL28m1dfbhUPuC4z7Rvx/e1Xk
D3JppcwkpMRb07r4bw1JnPSmf/1HJD36Ds78PvA7HxYCR3Ofag4nSIFW3wCrbxMB
TAz9H6mXP1ZGqz9o6tHnR36nGhWMGZD8wxAoakJxEFUO2OAVyKZpzj1tbIDde44b
f+vU5bVQWI+wOpBD8+4nR2vsmGVfGhmXycZRo7xW4NMBl/hDI1sWgxoQcqvovwuC
EusujAztPBXpriL3Y4E6mVu9lTL6Vnzcm28HqVL6mcvfP+9MmkokXMjNa8THkmNM
V1q0JdROp3+N2QtK53TqqbUUAiI6nHZokS7wCBJG3RapKh9rQiM7yvvvJAw8OnN/
XLUtOKldPrIppiuHtLsfjdmysch8j55U6zd2/4e/qnBLUB5/RtYO9RmtIS1LM3rA
VpWuzqxqpm2bFqa9twkgoO/bWKj9nfwBW8E7+HbcMBK/ALyV999MaOZ12cAHjOZl
PFSAQJYTW4ieyiKjguNWYAWzWa8a3RV6ZesZtWzzoRxxIW+ZLgBwHP2IsjolxcaN
Zx2YeSiVLbhJoAEO3x7cGLkNJnPvKfvIkss2im8zgrHpTkZajuW97DTbg6GyStFd
SNdfZKHprHEJXLWNIds7nH2oyTDJljVBFrfd3DXvMsAyVs3OW5bDEZFVKMqyeL9m
ir3e25mh38GRpYE+UwtqixF3jNWjYevZ0LCtBFkjhfamIIkun5h0jxwDbWd/En3e
hWU0kcex2AVVvpPqFNKHMtD3+KetAP+ewSuTkjKMzs2d1YX4vLUisg8MtpddO/B4
N8Os1sPE6gBtNSUhiOxXBQOTFoziJEt2G/oBlYbKgMSnq+b1mUeIFe0SxOxkL6tW
TLC7xlmqkMfrmMIvuu+Gg5IOPHEIQWsYgvKxQWiS3Dc+0Hu4WB0dgPE1LCQdAD11
Cnf+zE50/56QgU48qkcQWOTkJcpZQRL/zCD/2tB+gONj2AErBb+jfYWCdldGjB5R
6CkVMh6+AmvWDb08FPDfAWrRnAGTpRjyjc5oW7tm2imTXsFGDzt7huIHNmbhO487
tU3LIihb8iWu18DSYYbIAwhiXy0DNQ0CCwlAsSVLsftkAf08FM6kSotdl1witYPw
sLRK4ORp8lX3f5Pf6ehMS3GLbNu0rFtMAaa6kiRtol87GOsTf5w/bzMELIE1rjGx
6XbLRefE0GM62u8krrOYkpc9uX30zSyl33oD6fQCbnlvvWQ438rocrqpYeY7rvEm
ghLXm4mUtPUxfBluk8vxlPkRGxtWZBGr1ElfaYJHlcDf1wV8c9o+TCRezZpfQK4c
31bEodotN4X5PEjzc2Tg4+sb4QefMP2l94zHXwW0Igi7vgasuYcuHhQjmBf2siX+
HAMgeEKWy7Pt32nQS7/VDBKpzCFsyfrEyLX4WuYoMiuBoQi8nnYZvFR6As8lJdhz
uG89//KXAg5VrzFBZcFCoM+9Athoh2qQaVH0W98z2rNeKWjbjhS19qHqL/pxD42w
eDEvND3iChTZ3YwNwxCiT8TshxokD7xqlCmSbORFHB6d09FvNw9jZ8RatSMedrOQ
q8QCx+mKkbujFGcPgS8Pffm+PBCL0fX0fira353okw7swCaUUb0Lwb/6whR+XPzR
k9j/UHF5bnvwPpTXXgDw1s5fbbJScFVxuZL348pwrANFQ3Jeu1yNwMKqJrxDZttk
yCwSaSo35fzOtKYa+P2GyuKGW2F+M0fllcqT+JacqQ3q1QZmrK3APW4Tv2dpQzz3
NfLUz1OQz/qHqI5lSqFImwOJSEW0JHg/v4V9xtVWLtnqRLHH1O8cpvrzCLUyU528
MEMKffC5b3Vm/E4n9H3uirb5Wb53/y4zWI5gUrLTRY3Ukyn3Ak27q00P9mDH49kq
+s6UGN3XUBXgbYURMWziCEHXueJIRoEO9vcGHv7ttxgu0gIE4tdsFU/JsIxhYj4v
1/PFoSMG4i5FYtoz8EH4cwQ+9kYSVkAnthOhmZFhZcGPUOGr0w1398dvCk1Fv4dR
vwpWcKkz9LjVpXqw3ZAn28X/ysbPoZL7GYkO2Qj4wleHDVgxz87v87Lsq/hnA/DE
NHgQVOZH4r1Ulqx2Qh2+r+wMac8hscNWfpJZMiboZU42bfdJfdMONxJOqFyBCcQi
ziZSMyPIRoK+wtl0RIz2URYWjNSHUhdUx4PmihsPUJFPKEBmCRLdazSjYxyAjFly
BdvJeqPGQZx1sqzTxCp7khuYHZmtb94VftvwozVdgYb4vm/vwWCxxiib+BCBphCA
CQ3TCjws/Bshu3X/aIW6cGq6PmIn9getMZ+LPdNCwwK3caFSzZ56FJYGOkb/s3sN
njXsY14JgMkVuWX26SYFw4XPV4hHy5l8RV632zTMkCJz82DqiwD3gTb3yaqh93Rh
JcUXLqxbi+/hlB/8WFVGK6ccFC/4ir2188yCDMSXiIGNJEzU/VjNkRq6aMGfEwBe
fHqA4B3nxSziSneoNOshum5nO6RO1yXqRM2sp84mg4D+lyOTBNo8wqn7v3eKh1H9
ePMmgNLR43e+5M6amSOJPcrQ2J8e0p/xLSgviYPZHo7a4yH+X6AMUVGfw5iD3GfL
X14TsQWbTQ6arxJZ7WpopgML0aEutRasENml4Q4H+NM4w2fV1gOwioEUvYrm5478
WEfIPyMT1RCRASZ3UVmn3QIAaIELsg2JgAb3JCRl2MCU/rY46/zbwJfZ5ga9pDWs
/E9gRKkskAJiLXxcAbwQ9MPXfD0ugI8xvUixOD2EwulD+OOngg7OgNB12G3g2a8g
kApF3XKLxtzCxvzCQc4uIb0l2AIZHyGsaCsdf2KM4nuNPXLZGTaI94CL9u0/wReK
pQ9Bx63mHdWgQyEekzn9/fbS4ZdjEoIUsgdfnXIGf/Z9XxUpCzttq3OXa3A3QM0U
ojHVNUx6Y5Rn34VjzJgEw5tlh1RpWGryJ7iV1aEy1PaHb0OCV+uZIRQ2pdw7Is+S
QZTBiCsAIhQI4MfALsL+ZoqPooOtO2x5EWEivWtlwAnm9XhLF/hJCRF1ky86/UXm
uezzpq2LXSBkU2KsHaLcLvrpEu2isArzNcpOq2juUm9UbaiRC2/dWMCI/7juyB9v
jCnHbgXvciYb7bC6ehXvAmNHEkmFm8ezD7gkxwbJlg9YWtxZK/9JcLkf3R0mniEo
fxzvVJUPZYwenHWAUIQT943mMRFyXloeEyoeagFa5HfA31z2Zh/ydcIq/Ye6vIVj
gMqLNTAc7jksXYneqA4pgsrF7weymFoCP+l/C2SzR/qkJoobcvKZq+/AT3UXcltn
hELilrRn1exILzGEBwBz0N0b5/4hehIv/MnFVhPVEQIIwCuU7etToIw2u7JaL2mr
0q+bEMlTy9ErCIwn/wzFnBW4tL4DytyHqm/8WH37vzTG4hP0cdfh2fPsAkkQ4Rag
jJ9ewjgg5d706ljD9cEb8HirpdKO8GgjHeeI6XVAUqBioKJWgksf4QtFoWQ8pGxv
SU6VFl3SSwaWpuScC8qjxZfno8RdBNCanliPhgAPDNwK3yywOlEb3V3j1Ys2gr+6
Th4WaSf2gbfnJqar9j8Z8vQdOrRMBz0zY46mcDp8oAw4KA6/q7uFUtNce7VxQUUa
ym6o6j0sWnaoCI5Qw1As8Vjv03FGVna7WHfpqjV90DFUdxwDeUJ9UKclUC2hKAiD
f+Lry7Vu5h00MAcF4Q4yU/on2Hti3DCztXTmSwx8/N5F/s+CbQQoece0JjedM9Ty
BBfs0KqUMq+fWYkR1eKzrnAtBgajl5gyHzY8gYTOv7qJgaVRifTJoqE/u6AVnm4H
Vcu+0Kl2Fqz3LqM295IseQOjuo0t3BGORQfA+ii51CmMDs8CvY4DiM/UnpDIliFS
M/+ybrnsptuYYSStJz/J/TTG5Wc7bylLbwHhmzSNwYB6fM7aJzFCXR2eOL6AgvBv
FhJqIFBu/PFM3gnFdrdNQjf5sHPJvNT8PxTuI2FkheNaWJcElhx9DSpOo7i9qB03
urH+ZG5A/pl3tVW3nCW5jbXkIbyRt5rIZllIBdMwISbil0mok6aXMyUJXUS260JL
wZ/aj9tfg8+zlgtgLjANQBURndyY0kfBuVic4wrRbR+G8lqrLKJ2rXPFrKHYzvao
6jkF0azrbqhvJzU7fZGpg2rm1OGecm9Nhorlh4pA1N5l+ZrECMWINgOWeZV8Mcep
FEBB3OrU5n1gMMh5vlJVRWThlb+3nX3Iych4FksSflKGejo1Gt6Bf///7bVAt3UP
apLwrWAWq5KmscxLzD9b5RfdSzT2mELqxRU/4JuYIouvwD20rAq3de9xuA7sLVWI
viSPkvMHxuael/NDCinAPxy1fcvnFgqHhu/nqE7X3K4I8/JBRG6NEdFVpZfJBSIv
5Gv42d/mzbrUYU6c9mktiOe/cQ/OUAVBN6Cl0htlhWZSiKZu3KS0msJOFhO9Vk6U
9Q8Z7K/9GcAViH1LJr+u8cdk0lUelkk5OPu8Hic04aVWWGglmUgxdhAFbUhFjO7S
OCz4ZnSwmvhYu33DGq8dPhUxXzpR4evI9R+wXNWP67q7pdY4m2EDa33l5RJq+zRM
vijEbZu7ss/7ho/MeNRGjnhMQv0rLv8yPptv/ggcu3q/biQSecAxM8Z9r9oT0gey
BEcSiI7ACBaD/7ojjAwDO39jXdUdenGkfHtgdCZxWlkkgw8nKYFIeBJTtcUnS8RK
Tf4cb4DjGNRS3hZBvjE5uzKl8piowyvXqTvj7OhkKhUtKLtJ7NpAtq2UWYljJOFZ
9wlBtXht2tSB8thuTNoWkPrzBH7QqF56tD//5ydSbLlv1WBeQEH9p5t+DqUtKHO8
gXDLT11W3B6k/w5WxnkVlzIwnKiYdPTn2I5Yuno8IIsKkOyUnnzunQTerkuYoBWo
Zg6zBHW+hdlfpLgsyTATb6AnuxtXFo3iFHdlygMz6X0mCEIFxuswMsEE0KLl0GtR
lTUS2xdgQ+wJ0EFZ8hnbk0kJMhYQL4RvzC8STPz9NYExgMHZcgH7K3hjF+aMSovn
7M6gaa6/TfUoNfu2BMM4wH+bs8EIBiEgMPiPOmPwDjk6esHouONvvQQwayuI75UP
l/f+5QjlQvx82re5a/2McXNLC8ppqdQGIsQVvxVk+X24rgMw+OXyf+aQIDqGEZZm
yly+ZdmbpmIh1CrMFNcVwkLRa0KHd0kxj2kwKJTfLcW9QzvLoPxXj8ZsHyeTbyUN
wa31fTVTmxUxdce4Al+0mUtbFiD6VRTY8tTE6a1jU2v0QKptdIciA0AX5OLTum3E
h4N5+vl31m27dPmHnckUfJiX0sowlxMRpzSgjp3ghJ8njzcICPWMS/jfnYG1iBHv
1tvMczbJhsl17klTsjV+ltVLqsaVNrK57L/7Mh4CB3aG386HnEq61NuW+HEHJORn
L3B/LnzTKMHA6qJbQxltUGx/7QYdT3LXHCbVuP3nmuhaSw1xGgI6HoMYh6TZB1w+
dbfmFldr56v7f865kFs0jbbQSkEcUOnLvRbyUjKZ+BZktpYHMLMrXDAzuavSM5Zw
mt4T2irAUClrK9mLvqkZPoK3A92usc0mgAfQc2vrmG7dMaAq/p7AOgQJ/PTqRrba
ZWI3GWM7a9KTdH7eGJgqssXbAkekuHfbXfBaULyKHaG11WLTWA67TjuuhgHoWFI6
l1HExdSNjrKQpNQQBbguxbLWwjPyFaXVPiQf18FnBseSMW9rbDQ6RadGc/Wm7R0y
LSrXGzh7iZiR443/rdWfhIatSV+jWeW97Ry9J6gag2trH3bwrgN0LeHQhmDUYdA7
6YZHrcoaU++mGlIpJFqgSk52HeJfWw8M7UUTTtM/xFH2yt98x0qT/nZdk3aAg3FY
6fDl0/3GI4Z9RvGHgXluDfycmrZiJ9Lp09Fl59OMA8uhlTPcqvmrsvqhnxaMLOMJ
ZKzuRHb6DkH3X0yhJ0KrfFQDR2m0xhIwF9I13I934bhWR9PopLVkvxPSRvEN2k4h
HgHCuzCGIiccmg95oeH6VswlTtbrcoMSEmkbQ1h7yq3HhlhBVhCclowF1sx1cchu
rA/ISAvrHce10x7SFCc6ZvW9cKQeAB3OszKmHJfAsm+p7k/jH3Q2nO++HgXT5NQb
uda6VQbjgyzVMlmua2SYLfU8aAYAbPgKVDmvlJcv0om8BqoX5XohuCM8jq5V/RQA
oXFC7SwXMEdeli1hIjGbJ9h69n7idN9H4BBB7CRDmt+40RPS+x3s1N+/07oMxEwg
pfBIGI/87IM9BRiAkLGvKKJ8NOcQRY+u74qZrzK+l1cd7PdHDggOyM66ocuLyRvm
MZu+gZgw09RoXv5o4U1R6deTBfyuCDgKIyIJ0gHtgzFsfcN3qFPBnnhDkFWOCZrN
AOGep2GVDjcQKdgcePOLbDbtbG9pGnmcb5JVL1HsV0hdk/oCC9gnHBQ/OHTSqOaj
z9ezhgcA0wDnTqmCBQ4hBs4C1q21daaG9z6oqonv45/yWchHx5UbznW5rkb6HxSu
QiErwSGP/cR+uL2V98DpzZO7bLQcLNS9SZxIlW01JZb+QQ/AUquuUM/4GQzZ+CAV
80M9+YmxxyPreV9K4LzIkiF/zX/NiKgkB3C7H7v1tV5GguW7MsNz6u6qljp2Nmpw
BN+Hg2ZcZY9aD87Y5V0f0SKctNngPBLIlENJjq0IoDFULUIHkhPnbty3rcBPNLQf
I8kFlQXwES9vsYk73L0v2Vz4uegPPFoYfRa6BjK/jKR7h6PZ7opBc33eC4ljVKO2
niS3cJg9EhpXcpZ89wvymMFE9a5jX3grt0cIgokfa0MFmEfPMkDbJUAmtm/WH4Xz
dsL/1R/ulz/dJx+aYaOQ0hGQWPPT9nQjw15myjuRbgWqNv8IxO4q48tohayAHBa8
sOVNK/XK2/sjyYT/Hj9Rqw88mco/HUYHPOs6Ue23OwGqDjAZkguvnhr4Jq0aHDdh
MHAw5nzbzdvexbhTz8G2/sm4mEqw1Y7nRUBigFwgV+o5tukmLZK3Q7fBGzmM+s2Z
gLEPlBNOdBoBAqEDnDzWhsBeXqCzNMZtIXx174dSvF2yhzQtxFpqMf2HoKNnA/nU
BVfSh3RZr7x1BsE/MdPYF3Py+iEDroe5xOnTGk17jQEVX7DMeRGHY9yvh1X7b2Qx
arNWplD6GQidNM1EvczqN0oOfbLdWSLQChjWjFa11L1qFxqvPrUuVOAWaRH51FGt
hvv2FzNSNp1+OfOIC8fK2k1XApL/dIpc6O2Lh0SKWO0qftehY6F2X6XsXa7GjJAj
IC9moE8Ryhs09Pf8L9t5ih3gxZCUxFx47HWhURJgb5oi54m/7ooN6LnBZ9fTpY5E
zI1c7TMBHezeHxq9bqd9vXONPR8MVms6ZkEcDg/abhgW13qMAgqdih/ozytRobvn
YfcrZW9ZnfwtCzGOgqPH1yPq1yu753A67l5Vb4X40+VV2q3jYm4rfbjSZ+xaLdKB
WfWgqsr9R24L8IQuO4qsf7mD3hwtbMgx5eM9jfe6VU1yvC8f9KgWHykfjY08qbZI
VwJmUixEp1m9i6xe5G53G7HLAHdZQ+2Klnw9T2eCnaQzJNUOuq1R8kbAO9it8yAG
9t0BbL5WRNWBDw6ndqpJkYW0qNNzE4AA/tVayzh4ZWKihF+bIBxriKLxrl34aJt9
HeMqeofE/3kQrPZECAs1YCjUeRnC0FOiDR6KpMn37UknsvBUI6WdoRyJnNwEqWri
DjOtVkXIJviXlmfahsJszebcN+R0OaDEhJ/vkIbHvPROUIcrLQev+L7tMGGVKk1H
zzVQvViliJashe+nQq5wB0c1mvEZFvrLa8m0EIfbBqX4+grhkVYENMsuPF83s4M8
NMT4d780SyxH8aPYF7nz3GjOtjWEmbBlFiXVBccxeT4Em/9VvMibPU5bRhMdEuDt
3+sAk1R4Kzpp7xEu1fw8usl1Q/x7wxrbasWRN3xoatskLSPQmY2KDb5mgoluYMvm
3nDuY3L9/d5o+vR+cq3boQseYwHOaWq/CFMK2p2JilbiO2sbcuNZ2pwQit8e4fRg
n/R/DEEBVDvq8xqfhpz3uu6aoow7y9/l8HEe7tq4n0Lt/vickI00hfznSYp8qktC
EmMKgZztCifP4BZlneqMvulyHKZ/Gbf14vlo7cK5DiLAOP/prgqBu3aIfalnWB3U
uer4aj/99Gr6H/dlVNc/4ECt6UGP0ShpIy5O2/9Y2x6jq8kwZ6LTVyauEODzoqlF
0V5jCfvSiJCBUyY2UyxUGFzyRbet8x3Ig8nVqaQjumn8qZ1msnbWLuAnaqe0pkCK
Bt/oP8nEjpGYgBcVtOHm0SBAhH1W6OBi8v97LoSq0TpDxAiM2ZgNnNmPsrwkxFyt
6M903wd1RvxENVCu/zdvuLj6mkVj1g4CPrNMqonLVcBPLkDvKI7HJG4nQADiFbY4
MXMAyzDoNef+jp1kBU8Dq2tEzv7yND5llgtfBkCy/lF2w5ZVAUKqmpRZWssx9OA5
9BsI/WS0C/9dOAtF5R9xhgtY5KtJs/ej4VNAOGGu45Mra8wQVGurOwC59qtJcEjx
1HSh8Hz7JenfFZ67d2zMuWKZHaYkx3bd84uQLI8HUV0587IxI2WL4PBi4n3t1f9m
9tsMF5JsXkzZEFbfvUFCvzaKE6xrO6ohyQ5Blt8L5zOWG31+wrxaTEeGB1sUu3+e
Q01ZUIil9mMwkoQhCCnlpLekV70qK04rqhJwo44G5zrqeJLImTpDdnK5UM7n59XA
A8Zm32j3L7+9MG9hN0s70K2MvCyxoY5urcbe2PP9sCdXckVeBCuRRPeljz7l4ih1
DTcOOrC+jeVwnKI310kQeGahsRDRzYBuLmSzTO4Ul1hRQmhZjLmO0gT9RxHskSVo
8kcoUqLLQ9R3x+kPpDxbgogfm1iqE9bDwxkVhbYD0c33xNWYBRDougvFl1VwMHSC
LTxNX1eRsphQqbvy4qkpEA5YYVS02eitNbgaK5i6W5QDx4QhoZYRuMeNoiUwHt9P
e3m+L9Tjwsd58m54aI0YkbO//KXsSBWFzF+uYtKsjAhK20XqI3uDCrv+4zQ46iZA
uSwHUR4ezlwL4GbBbqsdchiQNd5WC4Uzf2WDRxgK14U/l1KavBzxTdUn4iwfjki0
YlZuoSaZPQOJaRHdyYs8eXB5medVsa6n2C+dfOtYnaBct4nbcQrPWuzRqANpXekS
Br+qYPylI3civJxMcl7RcXfPIL4pk9lB4BHFXnHaRqBFGfcRhQQbkZD71aq3iTKa
vLtKiK6Fm2IDSSmrftISt05TswItEyrcxuNTLD3hAC8nLxgh1OuSrWdKNI6f8tHe
ytUWX8vqiEDcQGFaB2iOPL/e8ZRvhgLaNiEHEhMM1HYop6l71zB4fG9xJ79nLZGc
YCxlds2w8lc+GBtHPCBp5UJ4qeGw2NNJ0FYeCzJKe/3QkZQYClCmOR4eqRVCPXaJ
KlKiYUMGDB4D55ieCqQSoxZGwjI0ko6Z128qBK90jnUomlI8QrUotbEOSXDXwbzE
/YIul2cMSmtAvNms6L+Gr5wObBEc6oZzDeZlpvomZNOnO7oRM20qRC5Vf76tmDn1
Jv++5N5rY1Lwu9b5Va2JywLqE+qrWVBvfyz4jJiR2VRL6rkpwCP4z1vUBZOQsAp5
TkBAVmkgl7legke5MjrpNhqFp2s+SWM9PbhKThDoK7PvsBCur0PNvEL7D+fi9c2X
Q7gsmvGkPGcUC+nbr/ckFUHldn6YSofcM7xXNx6H+a3E/Z+mYvy4hI3nhgcHq3eG
Ff5lfu1L7G1Xqok9uOnNJXHr7ovvgnupPb65TPUV0nu39p28MpVLBO3L92yftA/O
5+1YCvDa6PhsvCfq2eH6U7Lu/xnnEKn2/KhTF/ILW9GM8RrnO7kmHGAgKLQ65U37
q9fBhq3yEKnr1+wYPDDHkS3bVRwNXLDVzSyLsTxwnjaMJj4SL094pti5lNqVuVuD
KWmk4bFfB2eR02Q+MaFc9hehS+sficCT0pQMZQXBabd3SZO3fAHUvRWWL0kzedsc
QrIbtGZZu7hzlDvk7xpw/Ei+kRkxxhkB1xkAOaG6o9q+2yVjz2qJBXhRjUZgHxmK
xvOk0suhe09Zg3qxQQLVD+T9DY/fwSbHxIlYdsmSQERxg2eqR1FuV2YFH+s1UDFJ
xnhZ788NyHg70kmXaugF0RIz+xNG8ewsRZ/mBE2tqkItyEL31LmRA5XNSp9OE56d
3yASdu+35hQHjvwTpL/X6AioTlR3GK3nAL5/dYjaJSvS1RtCAnxhtq/AFdn/rNCS
rHCVG6f5GYtDxt163oQLGRtOQXk6AoHxW3cHuSYEbGNookBKF875k7jYIOBQ+Cch
R8jtd2/pzpEkQHxt/DQMwlCwth+/EK/GEyjMfpYVzUiFVF/1mH3BBqwk5Phd1xeW
SAgTvDoOYN7R3SOqD7fBv5Gb3nPx23J1Xm3FSXOet1K4QZ0+k75LJW6bOSdDT99Z
mnXMffPg7SvY4/dTbjEJbtJJy54f1LAgEG9zUsKi/2pJuIFZ3dFQPkIFshFC6fSc
cG4pvcydI2Ymz3TgwkkGmpBgkwpZm8U02Ri22IcPs17apPZik00N0k1O8yFcjhaR
YYsCeloRUZvk6IYdJWLbu6GDl4gOtTGu77DAJi/y267w+wo4ehWlfusmk1UM6RtF
Fb03jjY/R4Py4jkk7lLTtf9/3wj7swsy22Ym6Gd7FkLNFybZBhpuSgyyZugKPpyj
HvlNEQbgb2r/uP+rvWhe9oVetJtNlYpYV6saqUD/6Lgl7Y8LEFi95GZVVa6cXpee
FITk+miuofti9c73evLoerwr4Ok4YPLGXZ7Nr8csoJfGgz41tH87im3SsJ97Hc4t
pdCExNRHeDY884wBT5XQeopNqmDX36HAkxarXXZYHM4vaGSXYgaXYmTlNmsNYLUy
qsknI3J5E66Bq/XgA7lfz9ugPO/OFzd2L6DT+uSdUjXDB0+aOncC488/y1C+wxvR
x2mTtta2nPk/+vhLAUP9D+1YiD6X6Lj0MhIT/UxAG5hEbSNPuGwf8Gw/VDWWdVpt
b2cD1SM7Nr/CnFOru5G4xUFmw1ush/epc1rOHJ7Nk2mt9P+1Rd2iTqiXaD/C77tp
TctVyRJmYAALfQ42GU7ndBAmmjmd+tow8kA6j8CcQ91zNw2C5mTRVY790LJnY8Up
YwjKoNOYytLAty7ZF7saL5Ph6O8nZN5+Xmje4Px3rIrYQPRV+snwh84+PxCKKDha
F0XlpF1PNIhRoIXZ6VKWkirlyqNz25T8rsYgSUztu87inb8iUmyGeRoNuC2LcPCZ
YhIElnBM1Y2B5WAFnWRkVK/4rIWa03dp8RRqOs+GDgb3ylKPnr+yuvHARuBQPvj2
UAxxEX7tQLerMUf7OfYsDITA98zvirQyJm2iNu+O4t3uae+DE0BiWuTgRjEZPmq0
RzYxZCnRmZEcOG6U9jgUyMBEirMQ+TIC6ACuaUkgiq/l83fs7UM3O+UqqkLy7+ub
fovtfY4etTp9DZiugL7t9F6J/rv9DBBj7GocUzVMZJ0CgOlXxACt+qhZlrCkyscH
aB9kG03IS6TNx7aonBNA8r2S+wwX0W6BrFygtcWeYhGCqWajmYt0VEFWzMlaaOP3
LvvA9f5scW9G+g+nhwANGmY9ftkHEG/1VZ293hnCctTRg8p9LDlwvf8ZiZqi9bFX
ysLe90Sio/hRc2b1Q4JuFxf5TUJBPlQi5Tz68sqMZ9h2DahK3Gbvo11kqVA/+byO
UXdICzCp8njqtdr6H5bUppBmgC8glQqfEDClNvI1uLJRVxVGkRjCuOZZUVRHvMEO
8l09QKUgc0c1Q76PjvM3r2mhWwMYyv89eyuJpud8attyNGdD6AJeoXN+CMZbG25V
Ph2kqyaR98ql07K7BIr1/KcHV/rwsC7/eBqtQCi6CNgayIOHHag/L8JX+DrLjIVQ
IOGA9EN3Ah+GppCIUdtKUHSRBKrc5r0Yhf+8864ULyk7t+KJvmaHeAcK/V9d+1Vy
zascnEMpyvZuQB9EFs/929ysytEES444LkxYgVbO0EhAwYG4Z9yzeDB2nEJ3U9Kn
Jf2zm2qDS02a1+QNNN0vc28u6KnzVm0FARWTvxKD+BA3oMT8gkT7XYIsTEEivd7v
LIosrrn8avIER3kYd6PreH/h/4wr9zLJT+ho/KCti+2eRoOKlAjaVhXxzTAVPjPk
scLt7tWb9i0eYVoxmHjQljT6eZ+tjOZKvlWVRPI7fKIb9QrgbNZMK5eTiPV/ixSQ
n2GTyDfREJq0OykMnbaexI4OX6eTuj0o6LuFHMev5UL3sLXrcz4XGADoPAblLf5J
N1JOLAT3brTWPNehkBBeE2S6/K9jN0t506xHz2i1Y+59P83pNP71wff4OvzSZp3e
FQ13XVFrA9e97e9Ho6eZzcVUjiqzRFJDdXwSUvjUcebdr9TphPCfurv1aNDbqvGy
CDrM01DitEW1KCuNs5+HY6xCnqYL2CAyjoikKTcKdM3HHYP3/U3KBQLCDTBNbz4R
SBG0X1RFnyU+gCM+xhMoyVTye/YURPw68T0vKO0KxjDoZ+LGwz+kRpqJp7UrRmeE
NUs8aw/CoRkZbXUJl6ryhXN787tqjMXeNy2RS2i7bP1BlJHJBphoKv53AvYnHBBf
+rkhQzfKXYbCnPEXVcGE42JmlQQ6jeSVaRl8OPiCAnxodvG6XsBmIIL+vfSKPhE9
pqji2Z/paKKGaSnBV71SbJ2B/imFNz7dSVt8OQD1CId/ulIAtLrtn7YZQlFuCQym
RbD/NVtzxDI7JijzNqIEqBK9MlZQZfi70t7pgsyRgioUKxgNHmCUJb9UnPmKycNe
LNE2VSFRdAQ3MX3FzA+gxlLzwmO8fwdHd29LHsvLM/vfXH3iQZ5aRcmX+zfcugnl
Gh34d6AEX90+RCqviuiPY4E5S1PitzzzFcYuH6cr4WcgEuncrLo1mnrtmZrhOLbD
SHcxVIneXQJRxRNvmD7n8GGtZ277zVKJcWqxSbsiguCUKWgfQ5ZzyX4G5BBJ5uxC
T9gaFGlkGUx4TLaJgcSiS2YKr3kxkqJV6dCR0gDDevav0VXvJOz+V7DZDgNqQ/rd
rMdu+Fj0UMxqqHmnlEWJEluxauj+3kIkeDIOCafQ+lm4pVb4Y6CNiOUWFGFn1D1W
KCzuPraonN3WEi7QkRKBMLC0HxDnP5/SoSS66ivw81RvgjURbeSfmKkYSOuoIltD
+We45Hj+wgcmf9jfOrY7VCdaynY7GJOlT67+s1MvDTGJC9f4BycetVhkMxYsysiL
iu9wmgwT5tGUzSongptsv63JdUvYzWggWzd6ZUdQRB/REJR73ZjQ44AqalkNH8tP
hwJb9LiWcVjRc8KEntqHNntY/3FpUE1pLzVglO0Rln/C6WmUSZxgkRFyWbxQTLTb
go2JwZss064hRrHsGJMHQVS8Ugj1ElBIqVq1+u8Ya2seE9bSoZvfxDWZtONWb2WL
QJQng2kTWYd/j6G920xvBaEV2uV0zAzhLv6Hg4qGKmT57OpIyd6cwDXgWfqu8apT
cP/gCk9gwEExHF1mINz46qEt+IOLNwaW8nX8Mvma/FvkfOz5AHaovqVValeuKkzc
BQKuCsBoT3C7smHNJ/szwXXxeUsYKfj4SRxT0ZLauBBQ53x0nVkd3tP/5SLwnENr
KncfPcVFT2zR1CHy326ODJ87rk2l9SWScKXyQvkdXCkEgXvyaz15mcL3eAKumV9T
6hJ5vGGdkU+ObXXu0nSfs8FmItx/YPivbeX4uvOd/Pe3tCOCxanZIzR6mB6ocSkR
Wmx/MyCzA5c3b4iOvoS151UKppYO6IUSMDVW2S9O5R+QvnrLI93qv0E7oJwMWa/M
SZarq6djJuVnIcfbCQNng6dDXZ/fAJytAz2b3ByWTcWyCUII1MKKzKJv62o8QPBn
83rQhkTacPnIDrKq+SZBkCPI0lTRallbS8Io6C0OC2gFSovG4ni+LZSmX9tSi4OM
EAu5CBW7L96aDdGG94OJ3ZlhNourjUohK0k1mvpqu2rcQWd0uqOUGTtwZPDGk5nA
tvUxC6wgxBxa6YItapYQaOfZWbbZBc4iiidg8LirxImbDXaxN066xeYFrNOMlodv
TW1o94u8TPoZomumhiwAiGGXy1t4/s0ozPq5/NwUk4QLPkEd2Cgil9IZPaK+IM+Q
g+kLKYFGAF+1OSNm2pV8kQbLgvO+hJLT/ZkaoHkyJsx7rh+Zvema4kkP+OjkOWK3
W5EwQNOYTfuWBx9+QCpSCbwTlW59NbDSgFvvHgbMAhfa1AN7QI8x0KhsepZYPTQS
GRTbu7/7vYRpHhKGtk7Ux3IqGi/jiO7ShnmqfPKrFZ85vA8V5HKexvSaOS5nlKMk
8P7yVZDtOeEQtf1pA5wT4ddvULK4Cnu4ZA/ceHAdUyTylu6yaF38DdDkvlGWokvH
ag6vENsO4tJhhn5BZZXRGPSBGbXn4mvd6h0UYmvvrvTBfVnN3vqljQEb50OvUzsE
0sdUaQLngG6A3nr9MaklaYltmjvbQ9uALGJ6dpuzT4LSwT4djf5BFD8XyG9mV2RN
mMRjuTwzIW18hdDCoujgtSLZPCQJlNX0vOwvKTnitp30qjCVGtmCwz0msIxF12YF
89uTFzDQBg+fU2IjuNiK4IOevROJqMdofEv5slEVh4hRkcRpBVlMwr8t0FkjhNe4
ASRMt2LH/Q/P8brWo/+TvETcUODm9wAqmnVw0YuoHH0RbSRNKsnMuRw49caiQJAV
g8qI3ZS9aVmY6Ib74FZga+saN11E6L83LcokYbUp6rYjfAz1bvDCcTK+5elzYDfe
a6lZUx2+oOfdqF9IiQ8QoBF2V62KC09bKiyQVcsbKnXSRSJ1wTRrrElwmk/lkEv+
CUsxerNXX7Nkh/s1IzwGF07ykKbs5OwIxAyNLT8iOGB4bio3q8Mq8WWbEs1Zcp06
eQQQU2hPRQpHmXX3kaH1RXmby7MWlEdAgw6myfe+XaL7HWiXO4JDNafdpvfO71Xp
+JbYLnkqrqydItXn/Ff9t1HkMx/1/AbJQKcv2+RuucHIsOBNdbfICB4jP/bPDg1X
KGet6XJMZHaaeXqk8t9WXa8Kh8J+97HqnD3EnmgbcX2/EM4QhA64ZcGjfnUQLQQP
IyWiuSGprLJPiuA8P66OKIEfw3mIInqvzCTb6KJLkupoDHzPnuhTm8EuXOMTIz3y
CWPRWLX5G4YI3sNL1/fbLItm95lGazNwNld4nqR3aM9Su2zD6GBZUlO8L77vBEKE
rt4cAKAYIutJ9Z7Vn9xchWMztINwAigBqRn3WNW4IZr/P3Q1bY8rPdVqVPuWUTnC
GJ8RFFdRQ6mR3PqI/RtZZcMu9JVSE9PfpqQNntZo4ECdlktUQ4HZCA0VmBOXja2u
EqRUvODpvA5IV5oXq7SkEzJ0kDTWJf4pfno1j7wMhrHhU3Ehr4ng1pH1DoiqbaTL
INPAoWssyrT1DfRUulmGhkXl6l6f4Sg70JMm+a01VGRFDb4rtTqxmpM4j7fwvp/L
pqX4DPyMjIRM2yknSwlnYJmYdrwj8wfpvUa3FabnhByX2RnX82dYnciYR7lFNPOJ
WHg6VOR+Kdfj7EFiQHpSK/pradlRokKQSM5ykYotKpLT5OQa3JY/QjqQalGA8q/Q
qJUAE4r6EiJ8F92jsmXtnudrwpnseaCRLKYWh5lh8SUjHXqzv2TPWEo62hdYvnW1
gER6ybQOwQNbT8M0T4Jj4rRMErvUD4xrpbDvka4leYzmqtjeS4IamPv0GA0KSKqW
z9JlAIhNGRpKwvFhT7BGkZvLGrSunsGcTuejXOaFxrY0VRH0+mrTM7gJYuigc4mr
D0s1VJERkeJ8ByF1srxLhY/MHi+sula/7SstyGVvRBdCcfqt3suA7H0LHp7lVc3m
lj3vbmtlIQQiLazcBPeWQjSNhm/11bTTIfQd0tCwuFf/7hERBAVnw7JESWRwl4Tl
Lfuq62oqhsFRy2v53A/Ba38cSkLNTEPdf6/AIGHGc8l2CrtSnSWcJHV1VTelv0xf
aIuwoGMOsyIBL8a4KGfXdlyVAvDCZGGn4tx3w+JVINHqKSM/Ipb/poJgSyqs76V9
3vs9C4LVgHL4bx5h4lf4+kXlpTS/6wwe2BKgLqhFJWp2hzA8fSVh6SD4fpSqviOw
AUxFntv1DpKrVlqagrGtvNrb6W1ExnqLk8WlZOeO1yw092fjPKvRcQNcjojcJtp0
cHMhGWeKCjXEnbA+1DC6kb2hk9m7+a5pifxp7XbtTzGiw68nO18PNu052n5fwaYU
q9M+4cyeZ9HvRCu5mY76t7K8+avBKr6yjaApwQ/Dtik7myCF5snqyZUky/hyvztQ
aQ1XnBMipgrumu2GuC1VGzroWbaDcWkYJl66g0px2IpHSioACzlXqhy+sk8cYomU
4WZZtb9xpUN037SeeFGPAYXiz/9nm/SBd0U3QdWem5X2ty/NKruszMQFZLLdDhsV
IQh9nvr7OHrMwlwSRPtKLoFoaTYjRnI+8sVeeal3W1Lg3hwaQ5oW8eIiUo6YKQjK
e7leco+4jFWevuAThObhg229SBkbLmolJhVUzgH5dxcDvVQ3lx7jtPbXLT6VK1ME
H0J+hCJ8dpuyeWlN6sWok2BtGFvmhZUXfnrjh76VYFgdBupJrg8Xkl/VzajjtNJL
QehTOpcMzy3GBIfCSLpvuDDSy43PMAQFkDVV+f5WkKcGSqM1H6PnLZ7RIBRSQdHJ
TJR2gYJH0PUaA6/uCjtcWGASQiG8l0wpCjawk3ITy4rpXcV2+vshfDbkzI8U1E5i
Bp0fIkw4h9aio4eSnA3RsrT3TH6q3hhIv5kgDR5Ls3Jtl+M0nGRLoo026IV5/wes
cZfAr1xXL7tyi2gcFuUcG6lEx18eWS7mYtfbdYEI9p0O8OLmOH86G9Gd10/LDJSJ
l2xt/5oPjOEaVvZ0M1A3b7vMoyw/bdLkMDaFleGgq3bF2ObhFastbAsMTG/ah+vs
oVP6S8b1EFeLKqsBhAUchIctljmR+CCZlpfpNl94eyz6mtvHdxSWJXJjN0noboXk
Fxs8N4g07acKEsBG1+3h17Fp0LIRk5i19rCSlBrJ0reglt9S3+U/T3lhWB8qzayy
WDtXHxkStPJSDip5stwE90johnOKrAYaKlpTA6UkiQEcjog16rfMUHEhzkw4NI6J
WbeEDLAENbauF0LvLtJbJ844157n1WuCf5sPLLVvrUHCrKMaPQlZX9FrelHLqfhh
AEB3H+pL6vufgNLQhxj51Pap3l1494g33fnZaD3sn12i+Ylj8cgsl/Tr8RO5k8YN
kFAknU9IiSgfby3bbWxsab0q6gN8SRkGey2Hzr0s66Nld3KgQ+/EQVc65D9KIdxm
5JxiuRtXi4clnuWqeyCyaHADvK7V8rrVnmt10q4nVjMe8sbfDSWOuBs+AH3dS9WK
ux5VwACNFMztEZlnPVusjbXQNH5x9+1QVKleaW1p8KLysoTutv3UomzxbeTkd2W9
63o7EIq6SGIYHzCwIdhgkwY8PbjhGZdoaCyVF/FgxFhBHXtkNd+kAG3fGJ7eDcMZ
CNpsbbq8AYwGIiTgUeZMBONtPRR6ACJMgbOdDlUO7t8O/2YNTx7cBPhrdV1VNa9c
xrjeraCW2KpLosgwL3RBXDDKml8cLbDPANbtfZWtY9WbBGgWwydL9r7NDeMk8zSx
NAvjNDsWUVKGwJ1yoM8SGF60HV7mVVQ7ZGc06kxUq8wjhbwjJHazD6uz7uY6vYV3
F4MeatAIZaGxVot+lKYHab4aiTNfjVOsOxefwt+N8RsdVqv+pDbw+YWWR7KNnKSc
hz2xNFA5HDWy5mJ0993COcTRfTRKPB5nkPqA0AeLp6azn4exepllbsGZXZ6TTXng
1VaJmlaZltjt42/VXEt8mcZKTjB8rUrTJXtDXnJ1KtLNRJTuTLDd25HTAO+YsUCb
U75pP3iJa/6BDy/tKIHtc2Io88oI3YEI2bq4FOOo2lKrR3kjoG0bV2kctem7rnsM
ziIR9Dqr1usMXy8nJ0Ls7r6eF9wX15U32ZDbBvsGl0HY5fbGE74Vdpt4jlbCLPPM
idGIJ8VpmGDp7sLaVCeIVwQAEesvwoQyPlSRrzdyF2FfVnkq4OtevHnqf+Q0SHz1
XA7zFTWtHJxeK1UZruXv2BKlnaMsr+aZZCZkT0OcbAv3z4NLxVDxoYkNjmWC+Z5z
EqJM8H+MSrbQWQ0ht2tFLlu05hfB491LOjQVAyFbFuIO/UgLtYLQ4PD2cZ0zO84k
Q4/GXux/C5hCqjuRvLXluiI1ZN/3j0cmNimed8bIVHezJj8ARSqEOSqPRVp0vyCb
iWfPulhaTJG7sIeXp5zWsLuE3m60r2D7/nvBpPx/wXTI/Db3GxdO+s0HVHBLSzRb
WV5vv75SFjcrzcTebjjNNFqSHzUCAg4+uhGTPOFiUMcigQL3uUaSXTYK4qPr4xb2
bRUrCHq7eLrOm6o/u0DpvDYBZa8puF7SsUSeq4y9NKGMM2seRJUJjjX+DMdRVQ4j
H4dgZR0jJbQEWTVPi0Ou2N6oMJhjWSzQOHBq6PVeblBgpfoLmcKL+85HdV+xRIay
kJ1oKbz6ejk/tab1se9Ax8cksPOAx7FLwtmTr6cTkcRZs50huzL4TD8xFfnXFiOg
Njy12mvB9P4evdIyevHFEq/u/KRlSQebZllvebKkRmzcNfxJrr/EoPIqbqSo6Gtm
XPSjDrkZCZx9l68uPGmuWSiNVZzjMhP4b+XL2HwEkrg4HW8qt2HR+3y7eIxVGVd8
1IaPVZzNYy0j5eNGNuhXnHRqDMW95pUqITzPORhqAzOITxAFj94jIFTAkyP64t8n
q+maRM0QFsxOsAs60jY2SOWyvaB/jxJMg9oRNDtYk+i59nPbK/ftmVGgNdc5S6wB
Mpytu44uwIRBttq9U2+BW7fuJlQY3z2epkwNjBKkdRkIM5xDb3+dRW3GmEd94/du
offo5HdCpUS3H9RzcVH00uHMk0uAracdqYvgefLJVutOwQEzLaQA+i2a0ZYrkbAs
QRO+cOgTWdE13kcbNFOrQqy7hC1ZBTF3jWtafMDasC3rsssAAib7RKfl9mCCE9Ws
ggqC/NVL67//h8CSK+WkW+62aNLoSeir780zB9pPMidx7fsDgJXNfamvN8efGZn9
kceQW+iaLKOYA5vqypae2Ve9VgLOGxPUTgoMAE/9laCR6xEERnQwpULZLkfjE83a
HdCg2RCNfjyczm8EL4QxQjdL6Xm57vEBIKi0bisWm97rAne3iqcUgzzHzHH2cm/W
BI/2ZBEC916HA5UKq4Vzw15s1PuLsfx70yyzlKVqiyvvTLMvTqBTtLD+sFPg+GTa
NXigcgrir6+XQDk/DvUZVXy8XRghDFxE/ToZ56DkeVwhA7TqUR7p6OKnoGo6gcqg
ktzR6DCO0pSoS5wMihR8QtykcEv0WbpwEP6AUAMfsCbSLrlNrCy/twqWZMNnVFPU
MZ6So/776gs/aqVxUIo4Ka8vZt379TVf20tKWZC2beXQLqneAKAmhGdtDbX9dd1e
4Dc5AvPsLhqDIuenEOSZV3IT5XzzJvMZZIy/3enEZyN/vpHMlPjDjKmonOWjDOpt
K6pxyJamG3mkHvrljfW6zA48xm7D5RR+I5d0EQG1TecEWz2ZkKCcDjPYonSRAp6/
WKY7zoPNesZXNN97dpNypNnNyOCHJWlInexB/70GKbLvOeFyISjXjBMWR/3rtgR0
Tnj50Zz6f1Wkd6V7watbYKz41B7VPViqRBhzq5Uf7oxoL5irFi01cJO9Dr8K6yw3
lPHG++m1SKS8T1QepvjegZMKcmZtS42Um+p5UfoS4WCFg5FrIk0bOVckkm8lEtTS
aLnSXAI+XOf8DKry/aOtEOG7PzOREQ/mRuap/LSTvJ8sFGADbnH6ImwvrPWnvsZK
c7d/I27b67F/H2PKQmkxzg/g1kqM2hzcCif8FhHWcf3xoL5z6BsnCjog2CB5J8uf
2hhBcEq5hCiZHvePkJv1tKp2LFKWG+9AHDe1AOXCIVsMN20U5N9yXNzXhduyXW5d
bGEXooHE0KbmIaDCpIATnUbbxFf4zEocakCh/jtpUildG0fP0I6P9miTFT8eodg/
KvnmZDW4NuL1FgzcoKX1lzwUsMPS3wvkWLEy1hvRABQpkTJS20mIex7tPyKbJbx4
9SIw8N9Mgz/Q7jbIwOYbjSSdk7PcXbfXLGinxErODr0q4SVkU4do80glKrZ9k4v9
cB85+ja1pp/Ybl8affbqp72hxl/5rgILOC0bWIKe6JCAzEzSnIgvkfL+9iRPVPSl
xVkn/WM1XC1cv7QtvpRNJDVjXWc8NQwJtUACTmUNgDzmixLIAY03dmhqPKYlJ4vb
10QNQmUCSlwW3p4ziAt/1fxOS2/wdeFgvMz4xCYkXA0qble865g1tYRqVvLCEoKS
elO5psjhsaRX+vysavMWgj2cAhFC1ZlCSm+A55cRU93IM2e82K4b4Zlswy9SRPFY
8U8pbjD1MHlSmVP8f/qlrcBPT3wkQtRyXSSAVJoi6UvJvSh+IN4mir/+qHB3ywRE
MS1Pzf0bI1X/L2iOJRdtQGimUCVCqLpHxtK9Gil1emHEBYnPkpaVv5p1xBdKsNgc
ziVxIQdKaxreJ2n337ZLx3StQmgvyoIrgxuJwMO+20qd4o6koQAMYnrNwqx4anpa
/a5GT6wZs9228rgABV7wFNBca9ApZxHXbSPB4zhkQvhO4hW8z1H0RWkN/IvsyQmr
DVTDR5zr6OYRAa5OAZDEBVZMlKf5MYtMSYfceoNuPMlODaLzcFDGPXKsbN38T7O3
MrDwChk3+i/GZIBFNVkqFPWtqH+bXTzkBD73//z+mz4m8ELmrt1ZDu4rxGfskEfI
6GWY+FKBxEocekWAxpZ9TQRhI7W9girwQcawG/xrPeyvPPp7a3Ir50iyquKPqhzk
CDTV7Kt1mtBvphKm7yffnLs2kyGD5bWOYpq6zi5ytFKTQFvkkrZdP0tgv+wIZ2Qh
VZU97T3BhZPCzWvl70mZVR4mj8khnRsun8Y3niJwjbzXhtiAVlhPJg0DZ89yhyMz
0Vp+r1wgPuDpnfHBVZoDzQhQtRV1IQOm2lz5edX/AVnMzHYnqy0z16SOAhhyw7GU
9Yenuxb1bw3Tk5VlNHvlFm6RKLkFswPLWRN9H9R18MzrQOmGcdYR0TlNRz6o9dYA
CLq6HKYskoHXVL1zQwq2oLMjRPztYHmv7DkgD2equpfgYjeiaD8mPrZtMQFB8q5i
wUlAUpQSObASpIEvKLHI9j0xIR1vgkQzih7ltBK6IAKbjXcQM9CSykBRG9caMbTL
f3Wh5L6V2k8xIGvJSD9nL8CAYOB5Ly3GPQqbOQXOmhIWYbw+lIMmX0oSTqOpGNUj
4lAD4d6gOob3I0Uxtzh29jYxXQSd1WwF4wATZb8Tq9PHOqxQ7+0aa+R6nvRQd3MP
V15vXVsiNGH6NWN04Sh3KdSCMtUn8oT0KH1i63m8bh8UcxAOmoWefp4FICwe8b6l
2EwGYPUZizFSE/WkfmV2Rj1l8WNZO0gqI5GZZS6y+jb5fvzhUPss2xRonkNkDQeG
bAADHfPdw22TLyoJW0j7U9DDs4GVvyGsbzNaKKTZMmU3NVUW6Vpm4TaAvfXROVxJ
ks2MuoCNsacmiV5/wVr3+larp97WQURafo84wUXSTX+x/fnLkj2GjLNXu47ogxMG
VPXHXMIREFvwHTMDu3sdQ8sr15QwgX8eqkd3AsaT7S9a5aFaTsTudDw24Vto4b9w
bMzNZOtdsGqQAgzks30LP41k32c+0re0Fa1DrYm06TwNhP3AYHZCIrrOkUoR0Pbv
/J8z39zhIpxG9rx8HcngVaY+SodPWM5WYrtk2YCTZGNt9RJS7+ReRbSsxFHlE3jD
pcjE6Nh/SXOf2vp+YZlFpskS4mFu6FbfD5fEL3kkDpINkfbGwV+Oc5ze/SK6qcDs
8eB+n9s7ZSHnFpLB3xB2v8C+pYHpXBKjVkEY1/K/gGWHa1ht43c27/vCx5qBiTIr
Snx95K/3SPquZfVBEQwCqJLZQN40F44pKA7hE+4qt5uc3w4CguscdCNwtvbMAKkx
Th3FY0HK8r0OTzY0CwUcz0bUPoEbvbuG5R9qPTJrIXwkUu11K2tnznzyxl1rbb2s
Cqt/rem5XsinEUv6VzusoL72y8ybFXJFTIV0G3rQ8cLJY+kjng9YSa4+6Dy2H748
nzW9pjtsbMxMfYdG+P4EHtKp41lZ7eoY9qU+xWmKn0nmwb10BXxvgK7aM+JKcXRl
ljJYgn519zarP5s9Yq6BNZzaHTztuBYjnb6ao/ENDZn7udpKkrrRCtp1JtJMMHX5
JKJ8Cow/j8ubGiwxmaR/N2WFPxMR9DufyilKPBxgtVUh8bX6VmOspTtKNkug+cxW
DvasVm127pkfCfdwU2mT9B2hYxN4eV4oS4GfPGYsmZEyowzTGt5OwcDJvDyx6wVC
8IhGYEQ42s6UMxhTkpDYDof9Slk9Oc4ICiNaNwo4oUdezwaTZJHfht+WfPSdCdmK
ADjDtrYGGBFImWyz/KBeC5C8sQer8JBculTShOMMWCwvKRq/HgFzAGhogxzReSLV
9gCAx4f+WTGaOGYJjo8NUIHG4S1T/RZRryGz9wImKTUYxshFZT/kGYtfF9GeRrY9
gAfPjyEwEqzYOHlWXRv772gpzuxiqVWYVjwDV0Ip51Ymlm4SYWO6Wt3V+vUMs0jd
PvTRHpgFMQP54nhDXtn41maGrp9nyLsfWGwctfI/bo0Z3UAZtntzo50XvseNTDYg
1xDDjshFOSEr/LIN4qbh5BZ9BHyhOb1EA810k/tMVOwmL5GYSN/MZBUub5V/OGEi
YsqeEmBLeDBFaF/2TyPu3Jem+ydP9X98dcC9GI6Yr0AJu/j0SsMUXP8r+oFlDXJI
qc6ZuzBv9fNnM6rzszzlMyKM4vrnaAvZun8kc/13WbYPv6XzkOUZHAgblA8nBGsP
66T436iSe5FhY9Ntkj+ZFQjvy8W4wzAziV/8n/3Za3TXOl18emegNSghm0XwwQWy
TxPoydE5TH+UZBfwRU96QWKCTLnMC0ciQYFAa8PoU0UKfdUpFl6q1wwVqpDS5J0H
IzqHkDJQuBbe/wHLRuCgFMUESJt7ClinTLQfzYUSzKRglm8YXQIlHXzumtP8Ntoy
FybY6nQHzWt+UWzdlPzZ/Q/CVHferQhnOSg+LLZ1TTprjRHU++POuNOqjK81dcz0
hN13dPsgUZ95XAHt7u2+ZliUwMPdY77iw3czOJN7g3Jbkh2183k4g87BALb1UU3p
GvtRLNvsgMqS1g1nVvmNjXtDiKMrw58Tw+/Vaw54YrCxhfDzkT5GKSqTM356ZqwS
k1sImz0Le3BXL3kajUzAuZfsAJO80MPg2ULm007vY4BKckCdQCs+SMokQOADy2VK
uCtrV7THdpFCyDaUUdAc/uLw/ZJz9t42tBrKyvvp0Iyp11InbMWXQ9Xe8L0P4hHx
es4PRL6cjh00HJqOixFGwblGd1c53M4HECudCjpUVnd644Xb7UfwrkXnZeaGrdPq
Nn53BxGI4DJkdw7f7AxMyRJA4qh+yZR8+Tj+r/aNNg+YpkOy/S/YlfLO4YLqvfId
0Gmj0G3P9j9a31K3Zu8Z+rpQ1ZUZsAbrF2kIEzo1gA2//NrPcrz4wUD1EAjWeiO+
+3liCmOlWLmuiGv8poY36cHMvVT7dAXCOgCdOmd9+p+0w5tHTV1eyRTeDloEfUJB
BTgizHmHoA4h7eYVMZChtWVNdn1GV6E7vKgHsSyXONVXOhShGZ8tIMrnS8peTdPe
7oYuZ33uCnmn80eWx7EOx5DW2xBiTT66SDhhPZYjBWiJdkLqPufFuq+68u3q50rZ
VxocSCubq2tAHr6Fw0yAx66GJJRNJ10Vc8sFLryFt36iZGtgsySP2vph33QAO596
hEjqV4DnnejxU3GuAmBSpromCc/eb7uKGyVOeejdAT8saJhStKGQyk2fPfgBOe4P
SmTSvzZmY19k/3EDGeqhkDrmfsWfKmc6YA9h0McxLLzjuIrvXsXgauVJVKQkSw7C
DO9/yePX6qnumLSu4jutwUdOE0md2VHXMYsbblLmF0utpD8TneUU7MDyQcQBKBtt
jKpJ0IRvb0GUu8FLk6tck68tjp1L+0TaceNlbEgAnUxgaSlbD20kAlsy+gIo34Yu
rOZn2fIsmWuhGNINmvwHmpR71bKKwWfj4Fub3TGKYuGmzcdLCf1DI3QRO8Ej2x5N
YrrtrYUB7DbyzunzgklYAgqUegKKWkyefCTl/GkSuA9XB2y/lz3t/jE7O3ZZfW9w
ys6Kj0QkTQfCt4APbgjf5oZEu4u3CEHkRWOBtUakY91xMLDdh0AbkXI0YFx30db9
QmhEzt9GrTtw6mluyWIPb/0DrQEK8XZTwTLf6ytTsqus0l5NaIX3CMfgHSoRkqfo
hOrKTbajXv1ad1RTiEx9rtU/dIpu2r5l0Jzt9t+JirDGNggyhUinREHrdcb83GjH
wtc7+MxloVyV1iLkGYL09HfMlrY10wZy6/Y0l6a/xubIQJc4QyQpLg1H9dc9JWnd
KkwVtyisKnYZH1i77TuyUcjmnzJ14rJJHl78s3veaBNG8FY/s8wehjG+yNMutN+a
OvSuXzuKC3GIlxtSuRw+tV6y9bwUQ+5FgfC4WxiW/RJY0v39M4wjNzO+tIv5Ag69
2QKbNoXOsrnE96Ssxtn13FOrOEWEsANrItdE3P/D0tzibmsqIJzoj7pBct+oy/z1
s1Vo71/8D2+JfRti9tjyEo1oCfA0db0Y/gx76vN9YA64Py3+frtS4yuHeH11BToO
MmUrUKrUrFy4n3s43sAsz3jKJNkyUMs7EGEqyYE6DzFMB5VLwhKNvpe4Kot0J7mE
SU2lljX0j1yuXCA6HGbU/rid5nfpwd+/cZ/ZyHohSA+RlNyJ7wOvr68DmmPTrWx9
bL6vTZ3Ah6ocE3ZuOkVYq4UYZufK2GlkPcF4ovct+1CobPLZEvoft/5hg3PHw0He
+zzUNHU7hk/jScw3lEYg0rymuuakGa8t8LCfTR8Hi+zW04EVghrAKvlv2JCkRk0C
lBG+TgSRyRV5MrtHyOCoaTlitxEDY627RcLiFPSldHKWOv6F/1F739ib9KnFOLRb
A4Fz9F3QSB/T0BQpQH7hXUrwQKcB3+zMwT+vxuVyhR3Qf6lHYwCpQGdPSN/PGL7n
PdNtSejKF2zS3sAT+o2EZWZXk/XWtXa8UkVwSQVRue1QRbCxAZ7nIxLdd0E6q9Q+
AmvgSQOW2FSfUImbo4q8V1RdJ5CE+EHgTEy06q5Ma0eVYlmb6U5Js99dnSgdrORO
uN64lAjizN+wvlwg00hYbteuSSJBtOgDR+0aW8A2KmimthGqmmcpZFq9I0b6iLPo
K4lgXYdy/7A8cjcL3Eus5RzZO/kLXcB2GZgcVWS6ZVQhGv1RvSYouSGF5I3DhUam
r9gqbJ7jDxyHCyMnC2RaYk07SSuD4RXltfnBsKcBprS/Qd8+LfJ0rWtNewIHhTqg
qRmrdPJClIigVPIjrsfVwSs++ub8RGxd2FrRvqIM6RWqxDEBbHhGx+YiUuenXouK
0VG9CL559jnRkl21aLUH/TgvQgADn4/dQ83gv7K39w++TpnQhourNpARjYKkXIyA
3NhhYxlk6SkNugdgQvXoMGOdZznuYqsIZ7sw6oFh2v06toI7mdOrS+VwAxHqsFEA
t08eKYUEAtVpSG5h1SjSoSK4ef3wVYoBW4/AgPtzVzrerUEuS7ve23auVIuy+Nh4
yJiuVnra/icur8ALyfmeug3tSnu7TDmKLSqbQDrZYh64PjGcyBOEFnJn0N7Eb+Po
JjnJ30/qnJ3SKMPrG9AKyTU0BReFvEy8PpbynZU1U0Ix6m/wYfQgFgCNd+FJ6H3Y
9k/P4R5+v6zp/+9v3N6bnELld/D+oB/hrAipQwI3KAZ0zK3GHL+Z7oKFPF20Nyej
6ur7k773EwLhuPr19YTbG7XlkAXQYm0pdODEbHyKO66nBSfkWelKljiIh3Cntf2u
MaQ0U8pI+TGU5WmOh/Se9vOkf3ARtypABW1yeFxkxh6byIL1xzAlySuce5ELQo7z
tUOD5j49x8B6A7pRAcxSYimIVmQ3qYVjPJG98mXvFY/ChdoYWhgobrRZ6EOzJ5KG
bmHWqspLmC6+Ip9I2yXpjJ38X2z5PR6zibwFEmLJC/ZQOVWOz2iaEbPxXK5K7rPW
cfDcxaxgy7BNZ2uq2tufpEqR416/fpq/JuFT7F5+5v8cuCGCRuXcKLe3JcJnoWSg
OHpD8dhoTNs0DNkw6hhbt9HEpS6cnEFiQXJDlRGNZsgUeUYMcPT56lA43MYLtR0Q
Wr5CCkzWu7IJTEDDhi0iz0K+ZkbWKqXWGnjEsuuR0YnPjoLjgNTTQsOYPSQaCyiM
/9sgIyl6FsCRY+5xRv1NORcZcdRyQUjjejEL+rPQE/GJmoOLyYEq6yDMWr7jtuTw
UEBVArFaclb3Ntg9Ip/UqpObFVMktefzLI/GLIq0Ntv8xJGCCo8mVz0DGEJx+7qh
s1Sh0lx1RJ71I9Qz2cyyrVQQVt+DdbWNsZpMZovkyZvhUIfDXTsHQR05a4Vy0Koi
LUMnjkPMQ0DnmZjKsJftXraMViLzAtW448ZyuoAiAEGeMDRxmz+6BLLvD1Qg/4G+
D4hLQJGBXigoSgfbM7bWl0pOnh0Dl4+WFmkEXHxwY4szD2IUxlkWGU7XbDf/0VWU
qMtzUPHlD1JryAUkwR2ek7wpBTaAj4iiZZ6e7BwN7AEQnOM8HmLVZDCfCkK4Znra
GeAP5BZLIEFFIkv8r9GGBC6RkfWzLoBucq9uYq1T3+VCBmhWyA2ph7NP9IeplALo
NIMCAwnTs/TieYQw2j32iLKcvRlPLm+rePzT3JPfyTYECr5CwghrcFE+4hpIW0mQ
+itzHlvVPBmjC+hsVhmvzaaVa4es6GyP4U3WpfNHixob8aQexAwV26356ll4dOyG
RJmLSKrShbbLMo37TkbvK3WdEJWSzlwEeENpWt66dAPO8ApAyQXQnW9dzj7ER5Pf
OxJvpeV5ZllczzDvLjYXQ19qXEqd/fGP402fNcNl4NrSnrLgHlihW/uBZEUlbHcF
fAdG+bOE8XItEpY0KCVsbLyWe01Jz99XZtWJe3DsP9Kjlv6aKxeTCyJB+KiOjVa/
ce/w0olGBp3PoH+r7QH+PiMIDD5NXA7pzxAQ14w3aJY4WuXq4aZqoD9qhQBi5r7l
kwSuOa0YCmjEVk42kHVdXgXEkBn6NMazL1ONbZbeVkTg6n9p6fb+hOJlKQRFfaef
pw9fHLNqFDAIwZaXeksLTSzZpI1EKxtVbrbFG5aRg+VmPTLMZY2/cNheFKX70nTU
OrIaAhjvy/j9Whrw0yl1gYgK99af0YmP7X7javpcvgFFCg5KbFkdj5ZVWzxnaRmp
w8TJ1u7BiZL67qp7DTE4WG5k19AhzJ3q6x0OdUA1Lx1liIq9ODpCsPpD67rgXXRl
1KJtbEwI50fUOA7sJ5FhPHcKs6o1J62QubLDO5WVMqCiT/NJsql81FWtKsvJLOFY
kNqxT1B0f3ZJ/XAQcOMgYHL/TtED+7BhdJCwpdTodF19xFsVdVchj7D8ceqprizd
ne9CTRC3gWEihMpeNshFSUZT0VClBqG66iYer2VVTyic/d5WXPPz2rp5hDi6ZKkn
JGGz5LqVnMKJ8D64uUN1Ux4UN8x6kJHAoy6fDlrMQR3wv377rVXJY9/+Y3esKX93
f6lOgcocpr9t0U6wd0ItVzRqKImMAuIhgvUVETeaf7EKI/7pgCZFIw9PJgX4wYjp
b6jdRJRCLa8UU+cFJfAJEcSosaxNT3Zsf8OvxfqHf+ejOD1LHTbryQ4de5FoF/TL
O6ARf8STiEjWvNvR+VgaLhPO2f6305tALMQxRg7u8fe7L8pgL09Xv/yx9Nf8nA3U
/xcXfBZ6yHFJe7llnEeOgGGey1rgs90yRAymspXwcsdo5v9yB3YF7dZGPkx+wJoW
dxvwOUfCe40TBDSpnyrgf/MEXlWi/c+GvHFXkSZU/WZJXcFQYwpa1iyP2FqKgERF
ZfcyYoBQ/MZKaMmP4NnNcbQDrvXDJa58LNqvgj7JXhQ=
`protect END_PROTECTED
