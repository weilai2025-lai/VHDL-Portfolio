`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oToS6EMZjU5HnvSYnQ12DscB7GPFX143EO1ykfK0tMl4FbZmolKTeOFmwsL9gpAR
gvzYd4Fuets1/ttm+BHS/XNlSNjGlP6fmJJSuqHIsLK9QTRu7gb3g2fTkJrZBpGT
BO+GzU5AhJ7O3r7EfkpwIqtlQcMg0E/6e1HlOlMlHdbOitNnMbWqJc5TyehgsRH6
nuWs1mz+Q05EQL5iRbKxaKBKP8B9L93fzf+UxhX2hDu+mAIY1cE1jXI3CakDPWdd
hQd2+BKRWG+GybhPAECmBth4uA7uw6JrEx3Wci1Lt4IaOGdW8qlMQ9pEBdaFbakN
kElo0uc8qlnW5U0gYzZzL0H6P4PcmKbaGEWEe6x/XBtoI0uiTQuNCgAs6QQuMhpm
dwHXIIwuMYalfzKmJJ8xHk1UhFbBRlCCjYz5xKBjYuh0cXShvfQ71WPnv23YAWDJ
t2V206pBhRGI92tk6Ml2tVsfBEJ3E/8cvRmKmYkc90XllZ1j9xG0mdWJebdfeMvo
fL051FLUZtHxfxhkdZpWuM4q2eaanMUmcnrmN3qe+pla2fWoYkwJhNLFpWi9Y+sY
MNhcTkI7mWefivGvnr+VAgzR9Ay1t+rqOPFJOzVuG4XbBlMhN5eBRBwq+siFFRUQ
p3j5zqCx7munJXHLhn64XLjjZ9b5+QfJs0c7d666Yj7n2tPRJ1A3FOcxNOTNVlHU
UA/a1qBLRky4szY5L/n5dR6EcnXebb6WZIufkXunhqZN1zowWfJ5IdaE8qkqdGEm
f/mWqNsyjgP+/RRlG8FyjZ/1/ajgGOmfqcQWT1qJ04ro9UYdaY/ogOICNgMFgQmz
aW2zHdY0L8xfnghvafD8/kZ8voLGw5R6+4GOmkooV1FbN5bfrOEFL4ocPQHDnvtc
sDvUEHkHgF1+WZv4Rgbbw/0jzM39EW3+PaHVnCNojsyFHFltFV4/ej7KC/4EQ7HQ
EDwHBd/p+y4Hx/7WN+mSI9FTsB+cQp4+oXxshNPcUc3fXms0CTR1iukwsi68wKh4
QeXGyxCzzgo1425JD4a/B4WQKhqLI4DGYMoqLG/vlAJoAqKqFiUCN+saTsFSWUIy
CRA59afPdPWLPtEBtfp0XPlDIMsgtampNpq3TsFEfZZ2bMHQHjRwzeMze3dcdIXq
e2BUt7HtuF5xx2qgyKKF+rnPTUbAwflXkg00og2B2IUJCPa/aiiFJVDzmAnL8qvc
YD7U45e+VIWDrCRz5asRmvhvV7NjtS3f9ikrlvyuWjAihMyyEEtxOVozr3GTHlYf
O2F3mJoLxVqumua6Orjcf3EsMvH3WgF/7MX0bMnpqVwurNuVI2oDVvlbrJc2k8cA
GDHTSWV1siQSwG4oHHhbBXvUXxECvXfB4xruEXDi3kLs8Np3Z82SHO71FYC3tLX1
RPjznOKCz1k5/70EEnPLl3gjDQmsM25CBoZQ9N/GW6kWRGXUt+8+XA0F5Sz1mZNN
4CcRGaYGLFEvlyf1+rUDQSQ561aROOpcHS0ZllHlvK987hj5pKYWsdv08Mq1HiIW
1ZApIRC/6i99A72dczyCgUIdHL0EX3jElDdcLS5yiuV4rcwTErmZ72UylEeaZ6J9
Yc3vbORif0by0JttMmrDc8Uynm2miyIh5ep9+trMN3JWBCDmr6lkmXIXl7jTAijY
0ozu98fCcf3lASGPEoN27SGCw0PBU6k19iX8CGIyQePz1ZRbl+Mvuk11xHQAjUux
bdHAApYySqCvjaEG82GaVGp2ZZFOBpsZrRSDzX4WSF547QaGKUTE2BmYV4wSeg40
euvHUy3r8gsweu7Blcll00BjMTf7Am7VhV5W6rm9qS/iAj0hAKbKGAna8yqGrMJC
o+l7cRhzlSwYGPaui/OeoqxE60oVcwaiR2W6Jm5Fex3DXIJzOFTx351VM7qt66PS
CjWgynjOsOfeOZ94OV0D1+WbfSqSmDY8u7kAGUrwSBUV/Uhwg3TezlM5tq8J5yuE
2yfPqsHtmyWG2S6VS+pzUc1AkEquHoIZEaCOHom8Y1ZnlD5n4xelCFIikMPYm3mG
zmM0yN4GHMJA19W6pPrLxZ65Lq7Z3gDiPYUf4oKeCCvG1/qqfUp4DQCylMXl0hp/
p/VnRZNt/NuGNeeD2vnE3gwEYdsFdfVjMoJbAzXbREKfd3STzN5L5hMGwW3SdqAB
sTjEP9i61ppp+6gKjvY4MuV7QArvTw9u4BQvjy8c68BK1LUFOjQ70L15jHEMdC3e
YvOtiJr8rK60tXre3MiWbgOBRnIBhqN1TOevCUQ3YqvphwMoFZ4CjULiKdA+kDTZ
kCRcm5BpeRnsz2TL/+Fp3jacwCr/DY0tta1qpoAQq2neys/SpZmqx4LcPld4rquY
gBypcuUHaQiwBsMPmS/1N//ABDzMRkjSQk0WoewpCbnra/JBiw0bL2JwFRRlJJpL
bM3pFetMzUkerc1Rx77FMtPLCXKFYVosx1dr5rHTXaPrnOYFF0zRxJZMZOx27e1D
puQGWFA3uXBi1k/aUH+JNDA+C3Y/RfSGqYziq7C/fJIdhSCDAFKZJYYTF8lMcHOL
PyQVuWy8HnZNW9ySjyNwr1fE6cfcr3bAgbCeqgL1IecDoAC7UQLaIxVmv/sbrQ/D
AeIEE1MQXamwNkE4RQeScW7EFFAbkgUIOMifVB60cXnGWSqLo56fu1T2CEERzIrm
96LNqHUGfxHKBJaecNRJe4eYJWY29qBx0c6UstYFyfyrgsUMKHHht6jYZI7TC2Vh
6xmAhZ1tG3ISfLNo1cnGc3K8ZTSUojV4vhr0/JEjP4oAT1dRbJKk4jdz5Rqleu/N
cbgtoTfFpLBGxo8/DUXpMqJuRjHTizcm+60H6Y1nlGLO68X8OI+les5gE5VmL1Xr
wuTLQvtFufdqgMO0n/MfciZVHbAyyIuEhLiTSvoqeU/z02Z0eSPZhbyfbqEWk2NC
uPYWZv/8EIWxiNaajd89xbLKQZSqyF6MABmoY8a0NYcpXTskXlFigzQA8qZwophx
lg6vsqNzHNUc8X/W7PEfnSZufCmGp6FE3ERsuAD4k9/DNL6unillWT7fxWI72Hu7
PTfdf5fpHtbPfMf6Rwh8FJNJ8DXMeagdq0SWvwV7P8eKI16640AapOoCXeA6pUvt
BSyXazUfOCikk1NTWrZWDTqA1rDSTP5Afvwp+dQNlMCeFa0awqX0V+3pdZ/M2SJk
qvuKwCpPSSQ9D5Nq+HPGZvVmqXwWkkZuGohWuweBqH5HfSutAiRiz8gN1Tl+QEqO
xz846VY+3kip0DMnYFlctACuRmaO8Tu8s73sbOoEXEA=
`protect END_PROTECTED
