`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DePjE6z3AXXZ19ehPfYfE8NS/ypD+gXS6i9u0LD5kf/s8v0LlMIXgtCkVV6FjUt
SVjg7se+sS4VFPPzq1d2UySoRRYwhJIF0OcM4CGUlCIN3p3yGPZ0NIauIRBAm0Qv
lp6bPspSEyocHow6IqRgda8M/hCQ+N0PquV7od1hnW5BDypZipOI+ul4T9FIz9Ob
G4Ie/pW+McYDOfwZCFcRdxahm/WhU+XlQ93MhEL2gUUaeabVsNnKsEUmjorSmZ9p
C9Ig9NHAIH+8p3g37QYJ8IfaiuGtA6tOmBEthaN/kOH87mgS9bLfxi9TkqkhwKLD
cWO9fHZjmW6Y0fY506VcrhgbRthmvmw/wR5w2rSLzHmHGl0ySmnbhgNjd5IRtl7x
Tq6aoyxoZFYNiKee6f4qU091a/E0Gwbq77eMyCSiq3qIWRgUMSPycWFc+KBwxpsx
6dbg9i2/o2tAcjKrUBjKCXj1npXTZq+7NBqeCX7RHs/KfcB+bMfRMudDA7Gnnitc
l3zM36BfLiBFmGv2wyt/SHVeYDbYe7GAeBjV4dYsT19UH0dHKPNGC31VWJDTEdfy
gZ5ND5HQ+Wvu5euFRylIRCwlIuk55Ye+WanRWUVJOE1AH+Qr94jsY/OA9EiWJ0rB
CQ/VfRHyr5SsoIFhOXj4quY7wbmDVdH11PdQ9hqKJJqkCb+GgXnkz+QBBHD8GN3G
Ik+x19H1gf3q1zIQX5AUD6O/6l0sMLg88MNHmTYBrQB6rfPLhcWnkfJjz5UYiwPt
06ElS9vJ7kE6fphcq9gYzTSyAARN/NAZhM3YyEiJHkriS397F6A937v4Whbgqq+5
JQOZMlL3mnO63Gvi7qvrV78q7ajZ09KpKMQT8jRLcwQt4vqbKcS7dtiX7yNqdrvd
HWnNbKtvdRWBa6IhNpv41Kup6CPJBT0KUy9dKMXFuzcIXfn0LK+xeZ5Pt3V0+L5h
mqvf88VH8K+e1c9fsrO2QD5WzaDaB1vo/PuGjH1oBOlrxoy2bjnRtHMzVVzA0Efl
I1XAq9yJINmjZQ5DkCI+6Ge7M+H9tNzXeKiXYoDkMBTmCkWMtART1IAwjJ83wZHm
7pQg+1oVKcZnyRCzeUoA0uCZ7wyf4menHNn1P4dgnUQs6/0+uANp9A++IQUvkDOH
+DLLh+c41v6BNYShyYjqzN3FJYcJaedThqcyYeqnylIGN4Od5Dcy9jp3Q2NNcA/V
xbWbS1AiblxXvDD7q8PJ1Cy2uNk8AvXLVbhv8wOR+YTypNo7YtdH8lCS+RVWX/7g
T+IoHRW0x61G5Fmw7Kks1Q1AZ/+Y8FWRGhT/tvy+GShkwIr1VnlZlH7spkTcFkJJ
xfiUxAUKUX3nBqOIXVXV6ws+m9z5NttNPg9maKPHqEwayN1HR5etyiqW4in2ImMy
yfbFidMu0jV2gZ0GyqZXW7L/FAtM1mj3C8zPM8uwvcxRRUXsqb2CivFdJzo6BHMv
`protect END_PROTECTED
