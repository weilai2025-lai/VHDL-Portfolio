`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VWwGH/6OEtV2j/biYmHHuBxpFAXmoPpuJ9kKwETmyKUEJJScWUKHnWBhjHz7DuMK
ajYoowACDyuhszP+fKyv8YfUQi133um9Ju0NFnbaC4UV2h3p+ZqxO+NARFcNynW6
7va8FL3565iVmPE6aKb1b59rKnlTxjJeJ9zjalZXjh+k3F4vgQBYiC0j3/bdw6lS
bPC0pg4egQs41KMGop16QPp/YrBkPxbkXK816BdkdgBtMkNm4/jTO4HdWfVR8Oqv
LZgox+hU6YRS2USoMY6V+KHhv5MYatbI6H46vQLJdeHXkazcHMBQn2Wv5HhdkUpy
NSQONS6sNhTZe4qb/Y7UeJ/9Gt+0RV9o+7YmLLRWeTW4JlpqbfVLGQsYeTQ9+Q/P
PuFgkJ1+p/6cDlBRruqZPRUjnExaqj+AWh1IhFJ+OJNJMCW7K4rZ1RQPMqXTqngO
7nQ8kpnUKdDQQQig6lN5v3DSHf2NbxEi3sbCzapmWbgrf34k90pvb4jyfFKVhj3f
jUEoCan1p9M5ZikSHeL0esb4Jp2C1W4XlCT/ikOdooDZCFkfXZLpb7kirRzY6xzJ
0+JnPu1zWDdXFk2UkBXW7rnHg4pgaeWo+jHjtVoAT4DeVwvVm1jcMLpgFn/6vQyC
4oWJEi0NuXiIW5jM4nXOvQKzzFzTGxTHStxsQRNAanGoYnSRKxVAJSBvIjHhkSH6
+e6WlK9Cy1NMCPHFHRtjSDl1yxJolj5j9+jb7lQ1Bc18vaufQcmXiJDhOfRnNrE4
gXNKCQBIupPSaJwaAEl3l4SWZOXcW7rqaIZZYspQNWkE4pOPxZaA5JK6CT+B/xoN
R7wV0XxalYBpmeW+NyMby2Zg9yr79rtgmuQ9vfCBvHBri2/8VPjY9KtsCAudNjZr
7JiUnB6gsLG54yBGXm9Ve4G0BHmArdgfCBErhcYxVSxnjkd786QnCpRmtTMCBgYV
OSlzh8PDQwjgDA1s1terKrV31VF720f3Kq2xMW25K6pLgNjZF8dj9Z207+KzrlyO
Xw62tYt6D8rh//i3JO6Nt/VpyFOqNYC9Ki6eAiqUpIfl0N2HLpAdnUzj2Y15zAsW
zUCpbg1GWHal/OM2BsGQZq00QDxFuWxWU88J6ib6XqPQo1gHd52XVtNbtr7VKc7A
W5RV4FnGvqp97AmjU7lFGaJD0/92ceKD4kVcaJ9PFCtywOi1CpYEyZJqFW/DrmqL
g5rLmLXDSO1ZMzbZA/lzfZYNglBoirFhjzq2xpTnYS0OMaUFNUMcINlz2E3a7HzX
`protect END_PROTECTED
