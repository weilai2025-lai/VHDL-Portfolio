`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh3zm3mhqYIVxbkTeymByH4PUU78B0qq/+ETKsS3LJK8LJLqPHHxtlrlQ1STenfJ
F/8qpSAJJpT0+YH7ZZxlfXfY2n3jywF5Xb5nO2Efv9TqtDczakJoItkMljetLdff
ChQa95otztNrjtz1oufik4vX1W0w6R0GiOrDOzkktUuEy/VDKl+23Mpny9X8usEd
kNquNoDQ+earlhAQGxNsxYt7t0UvhvhNON33I6+zDU6qhI5U4VLaBD8tLxpKD+OM
Ulftwc+eUmpRMGlCKJ+U2AerN5dUuQjw/oUeMS47YjJJaTyMzfNl67hcLLp7Q26m
5w6pAJhLh+haMJgqvtni5yOyGl/hTihfV9O1L1bd0RkTal4lU2ZbzeUxvYk0cTSc
`protect END_PROTECTED
