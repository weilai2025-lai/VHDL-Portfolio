`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WiwPifuhIKC8bZRcoG6y2w/6tSTyqyVlSJaOZ6G9fB8lNXSlxddeOiYb/hOkr+sz
pwvFteh2Ami0k7Cg8nVHA5YWy2sUQATtrq572Dg6CWnB4M7LUE2GKwGm1YsE6eC8
Ohqyl9YuHBKGPDHz7EEN0kALVLSsjvapwkE4eiie6nxBObfECXcMbU+hrbGI1VDZ
CRMAj8NvvyUv9VtuCTGTziwaCVdnnMKS1Un6xFgT/SbH/uNbAAmOyre5Rz5V7iuK
lkriPLYbKLyWbHJzRsQk+Wb5T4fWykg+/fItLAz/xRlqpUPz6qF1srLWEDZig4Sy
jJ29Ee0zHXczT3wLn0kZfo/gIRdIFipi36HYQhwzmWTVAA1ehkRJtjgTl0sXMO/D
nhC07GJZi01oUE/6dSd9NsW2AIwS+31U07OH/572vBXbsCjGNYOTkX2QFS4necaE
W+LgePKAJSjKRMwTu1gMUkoG9EsgSH5QqCDsTWviwphCTvCa2ypsOOvZWN0tea1U
8gfYavarjyFpsvtlwF8bSlBIXizVncxtORgQZwNYOKoAVyf7FuU4bBXuCFAIITuB
l8tszOqCP3Spy1t707Sc63JZXxlhNHcWeg3+XAiiwgZ1PSV9bVOxeFFibah5OQkd
ECEbV9N+g+q1hkgbZ6Mu+QQVISsOGMurzLhBWp/xhKsj4Rf40fpVvtwcEo74zI5A
r4Y7cUkrF0OZ47t9q5gkpi6x4Ly23+XIoyyu95l5jYZ8L4G4efOA4Q1KsiuKn3xl
DZKzCIuXMTKAliIgHQ1Q+pssjJ8IvJyyROGx4rJFb0g3N/Ann/7ryF47q2dGmXu2
4lkRLAGC9hq8eZ/UvuB8dovQEGcQNm1fypR1I2pA4G9teKLlaKdorEkxWog0h+Td
nnUuweWXtf+NB4OuAMBQdNWv2+/gj2M6tbJ/fZgZIN0X4xUXBxBPt0fNEJ6QjqTr
n5S2JWt5TFN6qGb+vytxqIaWqnT0VFG4J9KjDROP/L3Zo3pvPN9dTxiKiYxWplvg
i5JlWFWtpRWGyDwQqlRlJhWkrTcBqTV5N/6J7qMegzdWhw9WoWxsoq65Ctb25peY
SQewO6yk3y9DWOivxAFMnVchwfh2ZeQuPJ6TXG8S8D1fVYCyqX7xdtX+l7RtnUAq
m6163py0DfAykMrdaH8s2L23VCRUdTfdGRV+22X8pRR3JfqGRrwz2Z2aHyNTvR5L
BHuG/CMEtL8bktXflDKB2bwSu9Hr2F41nIRM9maZRcn8ypqX7EQbQcRFDmbMe4M2
ofL7vG4fqJasFLw29iZcpM7k+9HW4CpsQGh/RRl8mKS1R9vXbmB6H2bhvRH9IicU
MD/gxta2M70LdiJMMho5LJIkK3nB9UMjlZzKkQAg8lNcjSyEdoXxnDHeaZeiPUK8
HwOT1xv6jaxLrgSL5A4twrZFcYl07qFkChN8elE5oeUKaH/uLbhK/R7qjrnHLqOs
/BUXgHkXwT83uaF7uvd5rHgaBdB7Mzr2x+rnXk/wfHp+U5tLudFoKsbAKXWtcPXP
oRwRf0AYXPIEDJFOeAtTu/ucFqElOT+Nmoj8bC3oE4/z3p3WFpJVkuY3nc9H0O3t
Y/DN9aFXdGRKbKhtKz23ZkoOulEPa42X/Pwlell6AOE2lrwiQbZscgzqbES+0cxe
YcVyQWloUQ/4WmAeQqAwPhNf0qV6wwAS14ExwJgaWlr0XoNP2THk+FZ9N1T9+fN6
OqVzcrfMPMW19QaKrBGOw0LS/wQxUTTXY4JH1uI8W9Eo+FhBavkQ8+yvMBGzdXar
/7fc7Zy4kDe3e8sDI3OZNiZpkZXvlfhkqzpsRe7ufqdVSwdsxqWKq7MciQVVrjnp
8cbmtnbh4qI37YvyFNiwCnuzq8dzs80m9zStiCtaPWWt24g5LYPVeoHi685kz5re
Drwn939WoiIk6oHkPNdGtL6d4xa2PQprKBXothYRETw2oP9BXsPj05jhgd4ID0qh
OXOO4g8aM6DP/K7TmqMbcYYI5loZQ19+jBZioWdy1wk4y2H3Iq8XUDbh6S+ALBua
k7rlMZKVxUPnguv5V5o2+R//jXFtQzOArM2PmsMshlROK5sbLXGLDX3IhCChUIUO
OFeZa/1kXie+qnlm7KCgVVI2Z5qCFYcocDsSth/LzuP01uGEbVyUzfeaiwL2n1Me
2gpr+n1WsLKxmhYK+ZjC0hK4pRWdTsbwmP7PG3aPfCQDpDco+h0YGKNfPtwsCju6
jHJ58gRNORXMNJKiDaStW8kTH031kmGZhT55vnliffKtZTeGaKz74GF+D83m/TWs
3c7PK2StYzFUEqtAm4WS8Oeav8dxPjhDKPQqyEsbHYbYE1vY6+NKorPx5BwZ9iEu
dQouE3mqV5VT/Fzw94NLpHaBkJtr0NmF6b0Sadcdlu+6QjFuHh/jRrlpk7mswlTL
GSMc755PYsSNpdT3tjvgaQ==
`protect END_PROTECTED
