`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjhV4Ihbc/ALFj3Tm5FQKMlBtLANOPnhF6nS4XXMAlFXsgk7pBXs4M7ZGpnXD27n
5WxsU66pMwUd4zOuMgys4fLlYEAWf5BUV1UooxUWznXkEH2wHnWJUZPl2GPcUCf+
/CKq/JrA3qT4BUEEjT6Ye5SZKyPG3K7wKZKDNGElBsykk5DC5Xmnmc3+Z5XVjNEQ
GWez+yjFeHOsbCgaK5c8rjZKiMjaT1303IXUuhuDbDX+lDm9csnUFP/hjh7GUjl0
cy241hgyOcLVrx3uI4LBGBw1MNddkIEJJOs9yXGt7N71p8pIvKiA5tEE8515PYJ3
y6nEeFDHXEYyBYMMjznDDoN3qwZxtxxCnoTUCpkk4FhLIw9hASvNG7iwa2YRi3xf
VhRGlamWU8yBvFz3j362TMef+NpsNW6KJq6qTvELxKWrRyeeC9OY2Yi626DuJ4hD
vLgow1ZOPp6eivfR/lAKW5Ri08m0ZGz5deBgiMnY4hZP2s5rPg5FSrnW1oUEHr+S
Pq5slexkYMkQjtTnNHmKw6I1HISDQqtMYkCRg4VkF+jws8vMlEUeCJbWOO3HYKZz
`protect END_PROTECTED
