library IEEE;
library STD;
use STD.textio.all;
use IEEE.std_logic_textio.all;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.nn_config.all;

entity Sig_ROM is
  generic(
    inWidth       : integer := SIGMOID_SIZE;     -- 例: 10 → 深度 1024
    dataWidth     : integer := DATA_WIDTH;       -- 例: 16
    sigmoid_file  : string  := "sigContent.mif"; -- 模擬時讀的檔名
    SIM_READ_FILE : boolean := SIM_READ_FILE     -- true=模擬讀文字檔, false=合成用內建常數
  );
  port(
    clk    : in  std_logic;
    x      : in  std_logic_vector(inWidth-1 downto 0);
    output : out std_logic_vector(dataWidth-1 downto 0)
  );
end entity;

architecture behavior of Sig_ROM is
  type mem_t is array (0 to (2**inWidth)-1) of std_logic_vector(dataWidth-1 downto 0);

  -- 將二補數的 x 映射到 0..2^inWidth-1 的索引；與你原程式一致
  signal y : std_logic_vector(inWidth-1 downto 0) := (others => '0');

  -- ========== 模擬用：讀文字檔（每行一筆 0/1） ==========
  -- synthesis translate_off
  impure function readmemb(fname : string) return mem_t is
    file f      : text open read_mode is fname;
    variable l  : line;
    variable m  : mem_t := (others => (others => '0'));
    variable i  : integer := 0;
    variable w  : std_logic_vector(dataWidth-1 downto 0);
  begin
    while (not endfile(f)) and (i < m'length) loop
      readline(f, l);
      read(l, w);
      m(i) := w;
      i    := i + 1;
    end loop;
    return m;
  end function;
  -- synthesis translate_on

begin
  ----------------------------------------------------------------
  -- 計算 y（同步 1 拍）
  ----------------------------------------------------------------
  process(clk)
  begin
    if rising_edge(clk) then
      if signed(x) >= 0 then
        y <= std_logic_vector(signed(x) + to_signed(2**(inWidth-1), inWidth));
      else
        y <= std_logic_vector(signed(x) - to_signed(2**(inWidth-1), inWidth));
      end if;
    end if;
  end process;

  ----------------------------------------------------------------
  -- 模擬：文字檔；合成：常數初始化（不再用 ram_init_file）
  ----------------------------------------------------------------
  -- synthesis translate_off
  SIM_GEN : if SIM_READ_FILE generate
    signal mem_sim : mem_t := readmemb(sigmoid_file);
  begin
    output <= mem_sim(to_integer(unsigned(y)));
  end generate;
  -- synthesis translate_on

  SYN_GEN : if not SIM_READ_FILE generate
    -- 以函式回傳 ROM 常數（綜合用）
    function pick_sig return mem_t is
      variable m : mem_t := (others => (others => '0'));
    begin
-- Auto-generated Sig ROM HEX assignments
-- Source: sigContent.mif
-- DATA_WIDTH=16, DEPTH=1024
        m(0) := x"0000";
        m(1) := x"0000";
        m(2) := x"0000";
        m(3) := x"0000";
        m(4) := x"0000";
        m(5) := x"0000";
        m(6) := x"0000";
        m(7) := x"0000";
        m(8) := x"0000";
        m(9) := x"0000";
        m(10) := x"0000";
        m(11) := x"0000";
        m(12) := x"0000";
        m(13) := x"0000";
        m(14) := x"0000";
        m(15) := x"0000";
        m(16) := x"0000";
        m(17) := x"0000";
        m(18) := x"0000";
        m(19) := x"0000";
        m(20) := x"0000";
        m(21) := x"0000";
        m(22) := x"0000";
        m(23) := x"0000";
        m(24) := x"0000";
        m(25) := x"0000";
        m(26) := x"0000";
        m(27) := x"0000";
        m(28) := x"0000";
        m(29) := x"0000";
        m(30) := x"0000";
        m(31) := x"0000";
        m(32) := x"0000";
        m(33) := x"0000";
        m(34) := x"0000";
        m(35) := x"0000";
        m(36) := x"0000";
        m(37) := x"0000";
        m(38) := x"0000";
        m(39) := x"0000";
        m(40) := x"0000";
        m(41) := x"0000";
        m(42) := x"0000";
        m(43) := x"0000";
        m(44) := x"0000";
        m(45) := x"0000";
        m(46) := x"0000";
        m(47) := x"0000";
        m(48) := x"0000";
        m(49) := x"0000";
        m(50) := x"0000";
        m(51) := x"0000";
        m(52) := x"0000";
        m(53) := x"0000";
        m(54) := x"0000";
        m(55) := x"0000";
        m(56) := x"0000";
        m(57) := x"0000";
        m(58) := x"0000";
        m(59) := x"0000";
        m(60) := x"0000";
        m(61) := x"0000";
        m(62) := x"0000";
        m(63) := x"0000";
        m(64) := x"0000";
        m(65) := x"0000";
        m(66) := x"0000";
        m(67) := x"0000";
        m(68) := x"0000";
        m(69) := x"0000";
        m(70) := x"0000";
        m(71) := x"0000";
        m(72) := x"0000";
        m(73) := x"0000";
        m(74) := x"0000";
        m(75) := x"0000";
        m(76) := x"0000";
        m(77) := x"0000";
        m(78) := x"0000";
        m(79) := x"0000";
        m(80) := x"0000";
        m(81) := x"0000";
        m(82) := x"0000";
        m(83) := x"0000";
        m(84) := x"0000";
        m(85) := x"0000";
        m(86) := x"0000";
        m(87) := x"0000";
        m(88) := x"0000";
        m(89) := x"0000";
        m(90) := x"0000";
        m(91) := x"0000";
        m(92) := x"0000";
        m(93) := x"0000";
        m(94) := x"0000";
        m(95) := x"0000";
        m(96) := x"0000";
        m(97) := x"0000";
        m(98) := x"0000";
        m(99) := x"0000";
        m(100) := x"0000";
        m(101) := x"0000";
        m(102) := x"0000";
        m(103) := x"0000";
        m(104) := x"0000";
        m(105) := x"0000";
        m(106) := x"0000";
        m(107) := x"0000";
        m(108) := x"0000";
        m(109) := x"0000";
        m(110) := x"0000";
        m(111) := x"0000";
        m(112) := x"0000";
        m(113) := x"0000";
        m(114) := x"0000";
        m(115) := x"0000";
        m(116) := x"0000";
        m(117) := x"0000";
        m(118) := x"0000";
        m(119) := x"0000";
        m(120) := x"0000";
        m(121) := x"0000";
        m(122) := x"0000";
        m(123) := x"0000";
        m(124) := x"0000";
        m(125) := x"0000";
        m(126) := x"0000";
        m(127) := x"0000";
        m(128) := x"0000";
        m(129) := x"0000";
        m(130) := x"0000";
        m(131) := x"0000";
        m(132) := x"0000";
        m(133) := x"0000";
        m(134) := x"0000";
        m(135) := x"0000";
        m(136) := x"0000";
        m(137) := x"0000";
        m(138) := x"0000";
        m(139) := x"0000";
        m(140) := x"0000";
        m(141) := x"0000";
        m(142) := x"0000";
        m(143) := x"0000";
        m(144) := x"0000";
        m(145) := x"0000";
        m(146) := x"0000";
        m(147) := x"0000";
        m(148) := x"0000";
        m(149) := x"0000";
        m(150) := x"0000";
        m(151) := x"0000";
        m(152) := x"0000";
        m(153) := x"0000";
        m(154) := x"0000";
        m(155) := x"0000";
        m(156) := x"0000";
        m(157) := x"0000";
        m(158) := x"0000";
        m(159) := x"0000";
        m(160) := x"0000";
        m(161) := x"0000";
        m(162) := x"0000";
        m(163) := x"0000";
        m(164) := x"0000";
        m(165) := x"0000";
        m(166) := x"0000";
        m(167) := x"0000";
        m(168) := x"0000";
        m(169) := x"0000";
        m(170) := x"0000";
        m(171) := x"0000";
        m(172) := x"0000";
        m(173) := x"0000";
        m(174) := x"0000";
        m(175) := x"0000";
        m(176) := x"0000";
        m(177) := x"0000";
        m(178) := x"0000";
        m(179) := x"0000";
        m(180) := x"0001";
        m(181) := x"0001";
        m(182) := x"0001";
        m(183) := x"0001";
        m(184) := x"0001";
        m(185) := x"0001";
        m(186) := x"0001";
        m(187) := x"0001";
        m(188) := x"0001";
        m(189) := x"0001";
        m(190) := x"0001";
        m(191) := x"0001";
        m(192) := x"0001";
        m(193) := x"0001";
        m(194) := x"0001";
        m(195) := x"0001";
        m(196) := x"0001";
        m(197) := x"0001";
        m(198) := x"0001";
        m(199) := x"0001";
        m(200) := x"0001";
        m(201) := x"0001";
        m(202) := x"0002";
        m(203) := x"0002";
        m(204) := x"0002";
        m(205) := x"0002";
        m(206) := x"0002";
        m(207) := x"0002";
        m(208) := x"0002";
        m(209) := x"0002";
        m(210) := x"0002";
        m(211) := x"0002";
        m(212) := x"0002";
        m(213) := x"0002";
        m(214) := x"0002";
        m(215) := x"0003";
        m(216) := x"0003";
        m(217) := x"0003";
        m(218) := x"0003";
        m(219) := x"0003";
        m(220) := x"0003";
        m(221) := x"0003";
        m(222) := x"0003";
        m(223) := x"0003";
        m(224) := x"0004";
        m(225) := x"0004";
        m(226) := x"0004";
        m(227) := x"0004";
        m(228) := x"0004";
        m(229) := x"0004";
        m(230) := x"0004";
        m(231) := x"0005";
        m(232) := x"0005";
        m(233) := x"0005";
        m(234) := x"0005";
        m(235) := x"0005";
        m(236) := x"0005";
        m(237) := x"0006";
        m(238) := x"0006";
        m(239) := x"0006";
        m(240) := x"0006";
        m(241) := x"0006";
        m(242) := x"0007";
        m(243) := x"0007";
        m(244) := x"0007";
        m(245) := x"0007";
        m(246) := x"0008";
        m(247) := x"0008";
        m(248) := x"0008";
        m(249) := x"0008";
        m(250) := x"0009";
        m(251) := x"0009";
        m(252) := x"0009";
        m(253) := x"000A";
        m(254) := x"000A";
        m(255) := x"000A";
        m(256) := x"000A";
        m(257) := x"000B";
        m(258) := x"000B";
        m(259) := x"000C";
        m(260) := x"000C";
        m(261) := x"000C";
        m(262) := x"000D";
        m(263) := x"000D";
        m(264) := x"000E";
        m(265) := x"000E";
        m(266) := x"000F";
        m(267) := x"000F";
        m(268) := x"000F";
        m(269) := x"0010";
        m(270) := x"0011";
        m(271) := x"0011";
        m(272) := x"0012";
        m(273) := x"0012";
        m(274) := x"0013";
        m(275) := x"0013";
        m(276) := x"0014";
        m(277) := x"0015";
        m(278) := x"0015";
        m(279) := x"0016";
        m(280) := x"0017";
        m(281) := x"0017";
        m(282) := x"0018";
        m(283) := x"0019";
        m(284) := x"001A";
        m(285) := x"001B";
        m(286) := x"001C";
        m(287) := x"001C";
        m(288) := x"001D";
        m(289) := x"001E";
        m(290) := x"001F";
        m(291) := x"0020";
        m(292) := x"0021";
        m(293) := x"0022";
        m(294) := x"0024";
        m(295) := x"0025";
        m(296) := x"0026";
        m(297) := x"0027";
        m(298) := x"0028";
        m(299) := x"002A";
        m(300) := x"002B";
        m(301) := x"002C";
        m(302) := x"002E";
        m(303) := x"002F";
        m(304) := x"0031";
        m(305) := x"0032";
        m(306) := x"0034";
        m(307) := x"0036";
        m(308) := x"0037";
        m(309) := x"0039";
        m(310) := x"003B";
        m(311) := x"003D";
        m(312) := x"003F";
        m(313) := x"0041";
        m(314) := x"0043";
        m(315) := x"0045";
        m(316) := x"0047";
        m(317) := x"0049";
        m(318) := x"004C";
        m(319) := x"004E";
        m(320) := x"0051";
        m(321) := x"0053";
        m(322) := x"0056";
        m(323) := x"0058";
        m(324) := x"005B";
        m(325) := x"005E";
        m(326) := x"0061";
        m(327) := x"0064";
        m(328) := x"0067";
        m(329) := x"006B";
        m(330) := x"006E";
        m(331) := x"0072";
        m(332) := x"0075";
        m(333) := x"0079";
        m(334) := x"007D";
        m(335) := x"0081";
        m(336) := x"0085";
        m(337) := x"0089";
        m(338) := x"008D";
        m(339) := x"0092";
        m(340) := x"0097";
        m(341) := x"009B";
        m(342) := x"00A0";
        m(343) := x"00A5";
        m(344) := x"00AB";
        m(345) := x"00B0";
        m(346) := x"00B6";
        m(347) := x"00BB";
        m(348) := x"00C1";
        m(349) := x"00C7";
        m(350) := x"00CE";
        m(351) := x"00D4";
        m(352) := x"00DB";
        m(353) := x"00E2";
        m(354) := x"00E9";
        m(355) := x"00F0";
        m(356) := x"00F8";
        m(357) := x"0100";
        m(358) := x"0108";
        m(359) := x"0110";
        m(360) := x"0119";
        m(361) := x"0121";
        m(362) := x"012B";
        m(363) := x"0134";
        m(364) := x"013E";
        m(365) := x"0148";
        m(366) := x"0152";
        m(367) := x"015D";
        m(368) := x"0168";
        m(369) := x"0173";
        m(370) := x"017E";
        m(371) := x"018A";
        m(372) := x"0197";
        m(373) := x"01A4";
        m(374) := x"01B1";
        m(375) := x"01BE";
        m(376) := x"01CC";
        m(377) := x"01DB";
        m(378) := x"01EA";
        m(379) := x"01F9";
        m(380) := x"0209";
        m(381) := x"0219";
        m(382) := x"022A";
        m(383) := x"023B";
        m(384) := x"024D";
        m(385) := x"025F";
        m(386) := x"0272";
        m(387) := x"0286";
        m(388) := x"029A";
        m(389) := x"02AE";
        m(390) := x"02C4";
        m(391) := x"02DA";
        m(392) := x"02F0";
        m(393) := x"0308";
        m(394) := x"0320";
        m(395) := x"0339";
        m(396) := x"0352";
        m(397) := x"036C";
        m(398) := x"0387";
        m(399) := x"03A3";
        m(400) := x"03C0";
        m(401) := x"03DE";
        m(402) := x"03FC";
        m(403) := x"041B";
        m(404) := x"043C";
        m(405) := x"045D";
        m(406) := x"047F";
        m(407) := x"04A2";
        m(408) := x"04C7";
        m(409) := x"04EC";
        m(410) := x"0512";
        m(411) := x"053A";
        m(412) := x"0563";
        m(413) := x"058D";
        m(414) := x"05B8";
        m(415) := x"05E4";
        m(416) := x"0612";
        m(417) := x"0640";
        m(418) := x"0671";
        m(419) := x"06A2";
        m(420) := x"06D5";
        m(421) := x"070A";
        m(422) := x"0740";
        m(423) := x"0777";
        m(424) := x"07B0";
        m(425) := x"07EB";
        m(426) := x"0827";
        m(427) := x"0865";
        m(428) := x"08A5";
        m(429) := x"08E6";
        m(430) := x"0929";
        m(431) := x"096E";
        m(432) := x"09B5";
        m(433) := x"09FE";
        m(434) := x"0A49";
        m(435) := x"0A95";
        m(436) := x"0AE4";
        m(437) := x"0B35";
        m(438) := x"0B88";
        m(439) := x"0BDD";
        m(440) := x"0C34";
        m(441) := x"0C8D";
        m(442) := x"0CE9";
        m(443) := x"0D47";
        m(444) := x"0DA8";
        m(445) := x"0E0A";
        m(446) := x"0E70";
        m(447) := x"0ED7";
        m(448) := x"0F42";
        m(449) := x"0FAE";
        m(450) := x"101E";
        m(451) := x"1090";
        m(452) := x"1104";
        m(453) := x"117C";
        m(454) := x"11F6";
        m(455) := x"1273";
        m(456) := x"12F3";
        m(457) := x"1375";
        m(458) := x"13FB";
        m(459) := x"1483";
        m(460) := x"150E";
        m(461) := x"159D";
        m(462) := x"162E";
        m(463) := x"16C2";
        m(464) := x"1759";
        m(465) := x"17F3";
        m(466) := x"1891";
        m(467) := x"1931";
        m(468) := x"19D5";
        m(469) := x"1A7B";
        m(470) := x"1B25";
        m(471) := x"1BD1";
        m(472) := x"1C81";
        m(473) := x"1D34";
        m(474) := x"1DEA";
        m(475) := x"1EA2";
        m(476) := x"1F5E";
        m(477) := x"201D";
        m(478) := x"20DF";
        m(479) := x"21A4";
        m(480) := x"226C";
        m(481) := x"2337";
        m(482) := x"2405";
        m(483) := x"24D5";
        m(484) := x"25A8";
        m(485) := x"267E";
        m(486) := x"2757";
        m(487) := x"2832";
        m(488) := x"2910";
        m(489) := x"29F1";
        m(490) := x"2AD3";
        m(491) := x"2BB8";
        m(492) := x"2CA0";
        m(493) := x"2D8A";
        m(494) := x"2E75";
        m(495) := x"2F63";
        m(496) := x"3053";
        m(497) := x"3144";
        m(498) := x"3238";
        m(499) := x"332D";
        m(500) := x"3423";
        m(501) := x"351B";
        m(502) := x"3614";
        m(503) := x"370F";
        m(504) := x"380A";
        m(505) := x"3907";
        m(506) := x"3A04";
        m(507) := x"3B02";
        m(508) := x"3C01";
        m(509) := x"3D00";
        m(510) := x"3E00";
        m(511) := x"3F00";
        m(512) := x"4000";
        m(513) := x"40FF";
        m(514) := x"41FF";
        m(515) := x"42FF";
        m(516) := x"43FE";
        m(517) := x"44FD";
        m(518) := x"45FB";
        m(519) := x"46F8";
        m(520) := x"47F5";
        m(521) := x"48F0";
        m(522) := x"49EB";
        m(523) := x"4AE4";
        m(524) := x"4BDC";
        m(525) := x"4CD2";
        m(526) := x"4DC7";
        m(527) := x"4EBB";
        m(528) := x"4FAC";
        m(529) := x"509C";
        m(530) := x"518A";
        m(531) := x"5275";
        m(532) := x"535F";
        m(533) := x"5447";
        m(534) := x"552C";
        m(535) := x"560E";
        m(536) := x"56EF";
        m(537) := x"57CD";
        m(538) := x"58A8";
        m(539) := x"5981";
        m(540) := x"5A57";
        m(541) := x"5B2A";
        m(542) := x"5BFA";
        m(543) := x"5CC8";
        m(544) := x"5D93";
        m(545) := x"5E5B";
        m(546) := x"5F20";
        m(547) := x"5FE2";
        m(548) := x"60A1";
        m(549) := x"615D";
        m(550) := x"6215";
        m(551) := x"62CB";
        m(552) := x"637E";
        m(553) := x"642E";
        m(554) := x"64DA";
        m(555) := x"6584";
        m(556) := x"662A";
        m(557) := x"66CE";
        m(558) := x"676E";
        m(559) := x"680C";
        m(560) := x"68A6";
        m(561) := x"693D";
        m(562) := x"69D1";
        m(563) := x"6A62";
        m(564) := x"6AF1";
        m(565) := x"6B7C";
        m(566) := x"6C04";
        m(567) := x"6C8A";
        m(568) := x"6D0C";
        m(569) := x"6D8C";
        m(570) := x"6E09";
        m(571) := x"6E83";
        m(572) := x"6EFB";
        m(573) := x"6F6F";
        m(574) := x"6FE1";
        m(575) := x"7051";
        m(576) := x"70BD";
        m(577) := x"7128";
        m(578) := x"718F";
        m(579) := x"71F5";
        m(580) := x"7257";
        m(581) := x"72B8";
        m(582) := x"7316";
        m(583) := x"7372";
        m(584) := x"73CB";
        m(585) := x"7422";
        m(586) := x"7477";
        m(587) := x"74CA";
        m(588) := x"751B";
        m(589) := x"756A";
        m(590) := x"75B6";
        m(591) := x"7601";
        m(592) := x"764A";
        m(593) := x"7691";
        m(594) := x"76D6";
        m(595) := x"7719";
        m(596) := x"775A";
        m(597) := x"779A";
        m(598) := x"77D8";
        m(599) := x"7814";
        m(600) := x"784F";
        m(601) := x"7888";
        m(602) := x"78BF";
        m(603) := x"78F5";
        m(604) := x"792A";
        m(605) := x"795D";
        m(606) := x"798E";
        m(607) := x"79BF";
        m(608) := x"79ED";
        m(609) := x"7A1B";
        m(610) := x"7A47";
        m(611) := x"7A72";
        m(612) := x"7A9C";
        m(613) := x"7AC5";
        m(614) := x"7AED";
        m(615) := x"7B13";
        m(616) := x"7B38";
        m(617) := x"7B5D";
        m(618) := x"7B80";
        m(619) := x"7BA2";
        m(620) := x"7BC3";
        m(621) := x"7BE4";
        m(622) := x"7C03";
        m(623) := x"7C21";
        m(624) := x"7C3F";
        m(625) := x"7C5C";
        m(626) := x"7C78";
        m(627) := x"7C93";
        m(628) := x"7CAD";
        m(629) := x"7CC6";
        m(630) := x"7CDF";
        m(631) := x"7CF7";
        m(632) := x"7D0F";
        m(633) := x"7D25";
        m(634) := x"7D3B";
        m(635) := x"7D51";
        m(636) := x"7D65";
        m(637) := x"7D79";
        m(638) := x"7D8D";
        m(639) := x"7DA0";
        m(640) := x"7DB2";
        m(641) := x"7DC4";
        m(642) := x"7DD5";
        m(643) := x"7DE6";
        m(644) := x"7DF6";
        m(645) := x"7E06";
        m(646) := x"7E15";
        m(647) := x"7E24";
        m(648) := x"7E33";
        m(649) := x"7E41";
        m(650) := x"7E4E";
        m(651) := x"7E5B";
        m(652) := x"7E68";
        m(653) := x"7E75";
        m(654) := x"7E81";
        m(655) := x"7E8C";
        m(656) := x"7E97";
        m(657) := x"7EA2";
        m(658) := x"7EAD";
        m(659) := x"7EB7";
        m(660) := x"7EC1";
        m(661) := x"7ECB";
        m(662) := x"7ED4";
        m(663) := x"7EDE";
        m(664) := x"7EE6";
        m(665) := x"7EEF";
        m(666) := x"7EF7";
        m(667) := x"7EFF";
        m(668) := x"7F07";
        m(669) := x"7F0F";
        m(670) := x"7F16";
        m(671) := x"7F1D";
        m(672) := x"7F24";
        m(673) := x"7F2B";
        m(674) := x"7F31";
        m(675) := x"7F38";
        m(676) := x"7F3E";
        m(677) := x"7F44";
        m(678) := x"7F49";
        m(679) := x"7F4F";
        m(680) := x"7F54";
        m(681) := x"7F5A";
        m(682) := x"7F5F";
        m(683) := x"7F64";
        m(684) := x"7F68";
        m(685) := x"7F6D";
        m(686) := x"7F72";
        m(687) := x"7F76";
        m(688) := x"7F7A";
        m(689) := x"7F7E";
        m(690) := x"7F82";
        m(691) := x"7F86";
        m(692) := x"7F8A";
        m(693) := x"7F8D";
        m(694) := x"7F91";
        m(695) := x"7F94";
        m(696) := x"7F98";
        m(697) := x"7F9B";
        m(698) := x"7F9E";
        m(699) := x"7FA1";
        m(700) := x"7FA4";
        m(701) := x"7FA7";
        m(702) := x"7FA9";
        m(703) := x"7FAC";
        m(704) := x"7FAE";
        m(705) := x"7FB1";
        m(706) := x"7FB3";
        m(707) := x"7FB6";
        m(708) := x"7FB8";
        m(709) := x"7FBA";
        m(710) := x"7FBC";
        m(711) := x"7FBE";
        m(712) := x"7FC0";
        m(713) := x"7FC2";
        m(714) := x"7FC4";
        m(715) := x"7FC6";
        m(716) := x"7FC8";
        m(717) := x"7FC9";
        m(718) := x"7FCB";
        m(719) := x"7FCD";
        m(720) := x"7FCE";
        m(721) := x"7FD0";
        m(722) := x"7FD1";
        m(723) := x"7FD3";
        m(724) := x"7FD4";
        m(725) := x"7FD5";
        m(726) := x"7FD7";
        m(727) := x"7FD8";
        m(728) := x"7FD9";
        m(729) := x"7FDA";
        m(730) := x"7FDB";
        m(731) := x"7FDD";
        m(732) := x"7FDE";
        m(733) := x"7FDF";
        m(734) := x"7FE0";
        m(735) := x"7FE1";
        m(736) := x"7FE2";
        m(737) := x"7FE3";
        m(738) := x"7FE3";
        m(739) := x"7FE4";
        m(740) := x"7FE5";
        m(741) := x"7FE6";
        m(742) := x"7FE7";
        m(743) := x"7FE8";
        m(744) := x"7FE8";
        m(745) := x"7FE9";
        m(746) := x"7FEA";
        m(747) := x"7FEA";
        m(748) := x"7FEB";
        m(749) := x"7FEC";
        m(750) := x"7FEC";
        m(751) := x"7FED";
        m(752) := x"7FED";
        m(753) := x"7FEE";
        m(754) := x"7FEE";
        m(755) := x"7FEF";
        m(756) := x"7FF0";
        m(757) := x"7FF0";
        m(758) := x"7FF0";
        m(759) := x"7FF1";
        m(760) := x"7FF1";
        m(761) := x"7FF2";
        m(762) := x"7FF2";
        m(763) := x"7FF3";
        m(764) := x"7FF3";
        m(765) := x"7FF3";
        m(766) := x"7FF4";
        m(767) := x"7FF4";
        m(768) := x"7FF5";
        m(769) := x"7FF5";
        m(770) := x"7FF5";
        m(771) := x"7FF5";
        m(772) := x"7FF6";
        m(773) := x"7FF6";
        m(774) := x"7FF6";
        m(775) := x"7FF7";
        m(776) := x"7FF7";
        m(777) := x"7FF7";
        m(778) := x"7FF7";
        m(779) := x"7FF8";
        m(780) := x"7FF8";
        m(781) := x"7FF8";
        m(782) := x"7FF8";
        m(783) := x"7FF9";
        m(784) := x"7FF9";
        m(785) := x"7FF9";
        m(786) := x"7FF9";
        m(787) := x"7FF9";
        m(788) := x"7FFA";
        m(789) := x"7FFA";
        m(790) := x"7FFA";
        m(791) := x"7FFA";
        m(792) := x"7FFA";
        m(793) := x"7FFA";
        m(794) := x"7FFB";
        m(795) := x"7FFB";
        m(796) := x"7FFB";
        m(797) := x"7FFB";
        m(798) := x"7FFB";
        m(799) := x"7FFB";
        m(800) := x"7FFB";
        m(801) := x"7FFC";
        m(802) := x"7FFC";
        m(803) := x"7FFC";
        m(804) := x"7FFC";
        m(805) := x"7FFC";
        m(806) := x"7FFC";
        m(807) := x"7FFC";
        m(808) := x"7FFC";
        m(809) := x"7FFC";
        m(810) := x"7FFD";
        m(811) := x"7FFD";
        m(812) := x"7FFD";
        m(813) := x"7FFD";
        m(814) := x"7FFD";
        m(815) := x"7FFD";
        m(816) := x"7FFD";
        m(817) := x"7FFD";
        m(818) := x"7FFD";
        m(819) := x"7FFD";
        m(820) := x"7FFD";
        m(821) := x"7FFD";
        m(822) := x"7FFD";
        m(823) := x"7FFE";
        m(824) := x"7FFE";
        m(825) := x"7FFE";
        m(826) := x"7FFE";
        m(827) := x"7FFE";
        m(828) := x"7FFE";
        m(829) := x"7FFE";
        m(830) := x"7FFE";
        m(831) := x"7FFE";
        m(832) := x"7FFE";
        m(833) := x"7FFE";
        m(834) := x"7FFE";
        m(835) := x"7FFE";
        m(836) := x"7FFE";
        m(837) := x"7FFE";
        m(838) := x"7FFE";
        m(839) := x"7FFE";
        m(840) := x"7FFE";
        m(841) := x"7FFE";
        m(842) := x"7FFE";
        m(843) := x"7FFE";
        m(844) := x"7FFE";
        m(845) := x"7FFF";
        m(846) := x"7FFF";
        m(847) := x"7FFF";
        m(848) := x"7FFF";
        m(849) := x"7FFF";
        m(850) := x"7FFF";
        m(851) := x"7FFF";
        m(852) := x"7FFF";
        m(853) := x"7FFF";
        m(854) := x"7FFF";
        m(855) := x"7FFF";
        m(856) := x"7FFF";
        m(857) := x"7FFF";
        m(858) := x"7FFF";
        m(859) := x"7FFF";
        m(860) := x"7FFF";
        m(861) := x"7FFF";
        m(862) := x"7FFF";
        m(863) := x"7FFF";
        m(864) := x"7FFF";
        m(865) := x"7FFF";
        m(866) := x"7FFF";
        m(867) := x"7FFF";
        m(868) := x"7FFF";
        m(869) := x"7FFF";
        m(870) := x"7FFF";
        m(871) := x"7FFF";
        m(872) := x"7FFF";
        m(873) := x"7FFF";
        m(874) := x"7FFF";
        m(875) := x"7FFF";
        m(876) := x"7FFF";
        m(877) := x"7FFF";
        m(878) := x"7FFF";
        m(879) := x"7FFF";
        m(880) := x"7FFF";
        m(881) := x"7FFF";
        m(882) := x"7FFF";
        m(883) := x"7FFF";
        m(884) := x"7FFF";
        m(885) := x"7FFF";
        m(886) := x"7FFF";
        m(887) := x"7FFF";
        m(888) := x"7FFF";
        m(889) := x"7FFF";
        m(890) := x"7FFF";
        m(891) := x"7FFF";
        m(892) := x"7FFF";
        m(893) := x"7FFF";
        m(894) := x"7FFF";
        m(895) := x"7FFF";
        m(896) := x"7FFF";
        m(897) := x"7FFF";
        m(898) := x"7FFF";
        m(899) := x"7FFF";
        m(900) := x"7FFF";
        m(901) := x"7FFF";
        m(902) := x"7FFF";
        m(903) := x"7FFF";
        m(904) := x"7FFF";
        m(905) := x"7FFF";
        m(906) := x"7FFF";
        m(907) := x"7FFF";
        m(908) := x"7FFF";
        m(909) := x"7FFF";
        m(910) := x"7FFF";
        m(911) := x"7FFF";
        m(912) := x"7FFF";
        m(913) := x"7FFF";
        m(914) := x"7FFF";
        m(915) := x"7FFF";
        m(916) := x"7FFF";
        m(917) := x"7FFF";
        m(918) := x"7FFF";
        m(919) := x"7FFF";
        m(920) := x"7FFF";
        m(921) := x"7FFF";
        m(922) := x"7FFF";
        m(923) := x"7FFF";
        m(924) := x"7FFF";
        m(925) := x"7FFF";
        m(926) := x"7FFF";
        m(927) := x"7FFF";
        m(928) := x"7FFF";
        m(929) := x"7FFF";
        m(930) := x"7FFF";
        m(931) := x"7FFF";
        m(932) := x"7FFF";
        m(933) := x"7FFF";
        m(934) := x"7FFF";
        m(935) := x"7FFF";
        m(936) := x"7FFF";
        m(937) := x"7FFF";
        m(938) := x"7FFF";
        m(939) := x"7FFF";
        m(940) := x"7FFF";
        m(941) := x"7FFF";
        m(942) := x"7FFF";
        m(943) := x"7FFF";
        m(944) := x"7FFF";
        m(945) := x"7FFF";
        m(946) := x"7FFF";
        m(947) := x"7FFF";
        m(948) := x"7FFF";
        m(949) := x"7FFF";
        m(950) := x"7FFF";
        m(951) := x"7FFF";
        m(952) := x"7FFF";
        m(953) := x"7FFF";
        m(954) := x"7FFF";
        m(955) := x"7FFF";
        m(956) := x"7FFF";
        m(957) := x"7FFF";
        m(958) := x"7FFF";
        m(959) := x"7FFF";
        m(960) := x"7FFF";
        m(961) := x"7FFF";
        m(962) := x"7FFF";
        m(963) := x"7FFF";
        m(964) := x"7FFF";
        m(965) := x"7FFF";
        m(966) := x"7FFF";
        m(967) := x"7FFF";
        m(968) := x"7FFF";
        m(969) := x"7FFF";
        m(970) := x"7FFF";
        m(971) := x"7FFF";
        m(972) := x"7FFF";
        m(973) := x"7FFF";
        m(974) := x"7FFF";
        m(975) := x"7FFF";
        m(976) := x"7FFF";
        m(977) := x"7FFF";
        m(978) := x"7FFF";
        m(979) := x"7FFF";
        m(980) := x"7FFF";
        m(981) := x"7FFF";
        m(982) := x"7FFF";
        m(983) := x"7FFF";
        m(984) := x"7FFF";
        m(985) := x"7FFF";
        m(986) := x"7FFF";
        m(987) := x"7FFF";
        m(988) := x"7FFF";
        m(989) := x"7FFF";
        m(990) := x"7FFF";
        m(991) := x"7FFF";
        m(992) := x"7FFF";
        m(993) := x"7FFF";
        m(994) := x"7FFF";
        m(995) := x"7FFF";
        m(996) := x"7FFF";
        m(997) := x"7FFF";
        m(998) := x"7FFF";
        m(999) := x"7FFF";
        m(1000) := x"7FFF";
        m(1001) := x"7FFF";
        m(1002) := x"7FFF";
        m(1003) := x"7FFF";
        m(1004) := x"7FFF";
        m(1005) := x"7FFF";
        m(1006) := x"7FFF";
        m(1007) := x"7FFF";
        m(1008) := x"7FFF";
        m(1009) := x"7FFF";
        m(1010) := x"7FFF";
        m(1011) := x"7FFF";
        m(1012) := x"7FFF";
        m(1013) := x"7FFF";
        m(1014) := x"7FFF";
        m(1015) := x"7FFF";
        m(1016) := x"7FFF";
        m(1017) := x"7FFF";
        m(1018) := x"7FFF";
        m(1019) := x"7FFF";
        m(1020) := x"7FFF";
        m(1021) := x"7FFF";
        m(1022) := x"7FFF";
        m(1023) := x"7FFF";

      ----------------------------------------------------------------
      -- <<PASTE FROM sigContent_hex.txt HERE>>
      -- 直接把 Python 產生的每行：
      --     m(<index>) := x"FFFF";
      -- 整段貼在這裡，就完成 ROM 初始化
      ----------------------------------------------------------------

      return m;
    end function;

    constant MEM_CONST : mem_t := pick_sig;
  begin
    output <= MEM_CONST(to_integer(unsigned(y)));
  end generate;

end architecture;