`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35NMxXJlaGDepjO0V02kjPyx1l7s2MfC8kiAC/gMzSD9GdfGvoT4MA63eIW7bzc5
4ePzhyCxjSh2ZIzQr70Re0BLniYPzn25W6XLQaXDogHhmE2W0miG02aPWXbY9IPT
0cBunEtdYrL4VuTGi0//7ZHaX5Wf2ONnoWdbm6bStc3ZH8TsvguHPGgc6jzN18WT
3hlwiviqlpVklm8ikUBAo/zAXQqI6RkdMrw3KynGqo0tCE0a2bki7kDNWEzPG2Kr
8vpnfuvwuppDh++oAoKHm9d646/bWeVbNLhrtskqC3527LW5YbCNfAv3cDlzkXOd
SdPoW5zlrEhEK1+pRXvUj1VTiaGkSbyOuS/G1jxHE2A6JYTsXYJXRUi85SYUpOoh
cdoF4QDCad+SOrEhI6YZKjZUXm+9y1/X7nF4q/L0mGFMljRGwQ8oQ3ue3SP31QtU
638GMrUCx0l+EFtHPm+S0gtC1N7rGlXGUtz7LFJ+ouHhiUjaPLb9HdfPR5i1+3Eb
hQthFZJ5FhcYqHOCKBKO5cSAQ1zkK6MKNFSSKEOwuhLvMt3LJwX233H835M3349w
sCA27UDdZbQn6NDyWWcDKhIY7l4bjjAb6nBjUQP146/RTW/mQDtmsIPPXn355sl5
itAKVZ59CfGZ46MTaC4/D7oduwfYwElpRBgxCJgc/LuM3ffGuuWdLSggFgyU7PbA
N4OQKMCJ6zy5ynKhNY1IkyQskcffTWqA8PMgssmgkEr+oZgoQnoI73Uwpcr1leHU
KI4HtCa6551EOk+sJlpgTknwVvfSyKAdfBPVl9wC2ADxGafv8sICnbYkg6l47JC+
/NTcKakqY1XIVhMIYuCVyleqmqIlElXzIOdcEosydxweS3f/JppeUNdZbItjXF0E
/kOY3uqnJou9StjWQSgdv5wwvc/2liPUtXnfbq+T3LJ4i8as+UVFEn1rLIw0ZPWf
`protect END_PROTECTED
