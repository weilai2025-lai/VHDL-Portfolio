`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrOJ4nNZ947UMAM5jl4apwDc4udh5XAefE9yL+thPk6urRAxKhoFBX5EtJyE3OEl
bTucyDKlQefabosrv0QUGl+am8eqF/MLEGBZQHPX5iYbV8cg5EXShib3pBqvCVr+
tmdRqkwoL+sK7ySO7nCKql98vQXA2iQmCykBLuJSYdPFb2tTGN+nLuuMzmYS4UP2
PzuMyMmYRnkByv8giekfEg3zbR0Cx5ckjmRLohQ5BfPGzUkY0x8TrjLVhUlMyrEK
dVJLl7k5SusaWTnjau3DKWBDW3LzMyepv6N2QwaDXM4Y5Z+eKygJxwltbRULdYfG
Ak7xsa+xHDkxlVzLkhQ3CvUEtfVq7LsuO3R0dAtYmsTUMZobobzYloDb6Pns+gvR
uW004wePrD7ddnMMFDc6MGzxI+b0JWcSW8QFxAEtrxRJJAmA6OP9VjAEHJymg23k
zCVE7+Y5mb5cWPg1nynv5JGO0SaNOhuf4Bvvxnt0iPnwy7PWpbVhJ1NRFfBvbY/y
B6hSlBBotiGgK6OCrfZgh/m8FdA4XBKueHsAXXmm43opArkxhrsHGjDdKPxnWmzl
VCtFv9jFzTLTkuADqZKZqub2gNOoYKb1SUcnWQdUXqxapTOmaNLEzuFKDlXkvbuX
a1cw8ebvOxvEEXvQf3i3gRHUygA9iWKGyJD7x1kEmkp7Tw3W0CNy6bTWf6zUsCz1
MwYU+tN1gQg6gcCrRV8wwLRI4pQrep4NlcaQHuYd0Y0rwupyC370zxYu/RQr918U
cmTN0xpwol9FV5vYu41pC1bjhWyFnIekaNSZgkUucYrtoArSuz/5FtIiT2R+Zc8Q
6P7kl3Iyself6j6iRQbzlBROZHOmFciYxHnry4ar91BV9KMJl1vJECay5EiIvktf
UlaAdcMF6g2j58hHpFdh4o8A+gd22Ee7kBC6XaH7edXWo4zCoeu7KTe70F+TMmaO
1pgWYqylpmq5Riy9FXhn0KPLZCn42C/C+/eLL8wVuxnF+ikZGCwLQ8vzBH2mQkIm
Ake3ak1Tc6OaKpVfxulEKD90YB/sumjyYzSJrrXvFRta9JACYHKiD7pgaoaWC3E0
2+OxvwOMQRERIMYwxlVI+goR15I10KfcDun7qqHeaBSonuuQP28KLUGKsSAr8kXk
X7o16kEIQtWMvTkDP3BkWm/tJpyy5ER+SM0/u/Qi2nYfeMnUEQVmveNguQN8GpjV
8DhTele0qMwgVogByeipuXJ8TCGqb070NrEYOVi6zbJsf6LT/xk6QW8E1yinrWJU
c3syrwR95qTjueh2+egm47w5kGpT5EdeHKjbZNy83m0QhA9vmTyi5eXjvdOLgzai
dJ0TSaPQrGcngdlHi3rpGeMoTIBFSmTqhINbDAMRpjwO3nP+hCsIV0CLLkYYg+nz
A+4wRnd23S9cRxm/GYjvfnWpE2RtfRz9z6TzZRgnEj0I94ecxEiy+TW7t0Xr6IZn
U94UvM/u+gHbDHZ12ZOKGJd1TzFSyWMPr2G225ato/4/eGmzqRO4gbtJoJlHVVdn
ejh0IoA13P5hOkQ9Oa0tIgtaLBWaEA8keaG8FCV6bwuArfSAKXgnbQlqnzsfSZcd
fmZiYo3C1hQUQzbZHLzTwbg6hVZcpH8oi3JNo/A3c631S1gynJUNLEDij7xrO7Yq
FBOllNfLHrwkFMA/rOsODKq3455mAldrcgtIWTNpXpbDIAWp7b9YD+PTCkB4P76r
VxKH2YrjFbQza7oIwUm+X16siVpdZp28UKpfpGcKH9JZxAvdzHml7fLJaXrserHK
nC3i7ekFKeiloMXJxQUNm5Ro83DcUlzfEkvgEMuObrWwsxXTnDric2yeNw2bzc7U
WI2yCqMIoulqcD8tIolrmaJx+i61gAY8nn5bQNyoYY9i/GZPvIyst1X+jvb8qobJ
8CTrHh/8J+ojw0FCZO8Xmcf3qgrTQHExxjcCz244rFECOegOkW8DyYoiYpeh9ZJm
oBSP3D8BmhSU2ZjIRt8CiwuUgdoCvcZYjGMEI7b2Rzgj7xnrWb+C/ET4MPj2F/EP
QFfrCKc6yDBtLR8f1FyjnoQP4lVLKrMhaB+L5bgt0ytBElofvkNS9HglLsY6TzkA
ByafR2YN3K7YbFdezYm38jT8ql3HYOnveUtMY82W7kZHNF/ii1COwr3i6y6kirED
nLHldOe8flc/hpEOgvum4NVEvITmYI2HvjMBNPqLDfjNEo5yb6+zyalelr6p5jZ4
A6yW5KEh6KpjKIs8FYdNgcO7qe1VZu4yc0/5/AZ/tOZeGbH8XoU9ILMyYT9oic4d
ph8m/b5Lqw1uz96S2B69ui7dvGX1mEcTVDmMtdmLKHRAbYZzANYARYGSOrAaxp1d
HtFYm17V0gAhm+rObyQ8t9c6Vl6M4AMLxdt9fSmsOHhXyf3+9Q5GJDCAfd9o+EQ/
awuFMxBmNWKkPT5R63Qh+3tNOYB0Oz2e4tJFYcQLK7xjm+dOgbU71kUiNPrDeYZg
BiHQfxhao7GgX5XnTqWDE+/gbx2uWs9iI0lGeMxlvanWmVyrAGdE8QcEOm4PgrhS
dAiOzNA3ZYmiS+eD/JEgtnntzEnK6gi2naILACnqCeWsyW3Bsiwah2RK2xz0pp0S
Tql9BvV/lDTx3LVyeW8AL4lRo7kRNb1B2vFjhjqnXzECgv/S962szKcEjcR9tciy
/M45g4T6YmSQUt1Yomlo+UkZyHEtcAqOuTpveh5CtdkhIE/TaxdyusrFoJ1UdnZX
r7+/P2R36s+7D1eaWROQNWUXjSo9FkkvKN51xv+KKVFBqTZ869+Hg85XRF19ri5N
K7/5z7b9yL6ZYT9vzQs/WoOz/+uUWcjXlFQhAEpRj60wVMN1OWUDChnBSxcwJEaA
4oQBjFfIHZyisblhl0O/rMyZkBakXisMQu5wfdnsFNwFxEyJ13enEQE/OKwQ4TDy
d5DLdNFSqivkcvepxYKRrDNllqItxKlfR0+1CyoatrDzWqwPZg1HRRYq/3fVSk9t
4T71495vHc2jg11x2D1/nC3BJhO1BsE7mO2gSzli/ddHVDyWfuTqDobeHjDTaEgr
7u8ZFchiDnJs2TOVGHISzC/r2uYuC0XNxiwJqUXVcLRqtxr7fNeyWxoSs5XfIXMT
o4Z/Z6xH1lKCozOmnYd4aVSPOSagCrmwo/NFofw95PBdyTlHbEpHgOMkvpRDdwmO
kKymi7gS3wZWilLoiO6LvwLAjy7at/QnYM8CbAsGwGfKlT67sNtE3HpdetadE/Pu
mDOGlMSSnPSlgWv6srmujfOWgtkxqgmVIVOPKxL6ze47gWtg7xgR+qQuPXG0VB+t
qi/qXPZQOQ7H6h/KV/vWUSs3ylt+6Z4msbTklF4VsP6zUPnst0h8K+DB0AxPjDHN
SKan+HPsT2XCXc0z9fdovuAuazpJw3UmjX/QEWp2jyZ4s0vrz8/Wpb3mBfi7gRCY
cjKtNvm3jECZ6nd3CUOFWzRewbiYrkoT9Be8mJ1Z02610riLGUH8lW+jBegAs7oy
IpmEMLDp4D3cB7d/OQuwUjqstJW0917ME4gbfLD6vxBg1iYducVMSPpAY8DW156J
7pZl53dbw9CTbgpIrpe44phD7X8fG91TaUqkxS8KdwmCyr6ZNMjgmVSm7qds/Khh
90PvFkpQcLJZyFUbYoaLSsygehj3RxsheYd3QCIyEEKZ7Qq6CgaJUBI+xLp+qs7M
JwDiRpLATMC9lkk+d1uWuwsm1nnEXHT2CTZLqltPurw4+42SEW0XPERkUTZGpEHS
NjCbsffge6yFisQOrsEz9ebytYqDwqNjKN8t5xTyUT4e2R3WoyDGtyr7aUw/Y1fQ
IWTzMUZN4MG2bMesSSNErQAyCh5EOj1nb4QvDkQCQg87BLcE5LSlhtgBe+a2YEOE
8I9Cb0RC668KOWQd7cW8ruR/E+fZcGFmrLf8xA4HFmRDn4DnZR0CgFMGxrHbGNYp
vPGmzshlFxrinpMdxYSBJxHLRGg3OjgYwezGIRxEW+lj1Etac+StT8cB6GbxHt28
X0XyS9iNzG9TLYuySN/X3RmqyNdIENcCM+bi4R+xIrBzF5ehmNFLumQX5G6Uohcg
QajIIEe9lBXP8VTf62B357VlPZHLcSe0QwgUWhhO6/wzciHhZPdTc7tQgSw7moM/
JBEo/Z7Twc5hA+2dWtW7ewk3JbU0K8m9X0EjNoLwg+/NP1/4DD72ybx8FiJcj6+F
AzEA6ZbZMEr8Ji4TzKDePI2ObLEqquvezJqT6l9cKsX4HJ9x9+MyvBMs+oeu9GN1
MQEjfKWaiSk9G6wbSoThURTjpjlqU8K84q6VbZXY2B3DIUK36Tt9CukXPp1j7gJ6
gnBIgX1X7xxH/YUusSoMZjfsepYx4/yHpzL5a+mYrKELTEso2noXPPy37hkjt8ly
8XXrbSPQhiEgAb750kC+Bdyjtuh/ZkyKdOrU5q7FBwwG79nczTN5SQNgZR6Svtyi
IrbxOVNUQmejEPSUnuMQmCvxlrEzsGBrvU9JdW1AJAzrwtV09eexXIgloq6zEvB0
354h6TEbTgtMLtqFw9nV5ITdBKB4RLztsHAdYlvkZghNhsG+lY8YN2viJyk57qYm
71Si/SDMJhvzWFvwiD1k4+PvLtmkTGZS55jkBrHB99iY0Ao7EETrZRSDMvk3wA5u
CsXPD49+IUHM23l9uDHh+nCSBO+a++cNR1HKGHGf3lS2sXoXvsgqxSYnjYn/uMTc
sjhfjxWkNmzNJGE+9mbd3kV4b/5ijXUBGi4wu+OEOVvsgBLqHadeIIzhytGqGLPH
R9v3qvxCKrUdQ058IQ3ENQq7B3yB4pU695fb7Bd2mUND8MdyJJFxjzbtd0VBiKYi
g0tfG0gT+D3ryIwOVC8E2TASDht7HT/A4WpZ2z+Kmc5q8UBboHNoSnPhXVp7H5LY
WE9N/JQa0XM6lKpsZbLUTouelupnRxQj9iUuO1Am1RjcEwowNxceRGBIgaZtz0yx
+HhquxFMmOMgNzFdabb4PC/2mSCCegw6V2wuoptYt3R7felbsvVz3ScjwtLkj85Q
2ojWn9QsfbzLWmwxGhd5j3y+jesA2w52fl8NvO23R3SAhfRC8IG6DksBpA+NtuTc
L7g+soh8NweRe4pfdYXYEtyt/KEozGCYWAGPVvLjEXYVVnmGTRF9hBr1F99A3di4
EA6X6/lkhAth1818Y/9igmvKd3qiTApWq+e1StVoYr1OD0njjNo4XxaJUJhC7nSJ
8i01TXGOe8k/26FWrYXxfPA2wtR4hgkqeOaq9UHt+9tpYd+bqVFGb2ruhFIHBbQA
75nc0FWgALY4B6ZyCGxeTnMhunpV0Ja6BPskeBRHsjXQtctSz42vgOUZcYeGINNI
ZiIi7aWuNS1R3UoT80j6ktlddqpieTsOOs964fNNCioBUElPE1bHU1BvR8fcvC+H
VTnxf0NfE8exPhmM0tp2LSWdB9TUgHBVgfuT3TH/4GzMoj7ANvSC7u1AK7K95Ian
BIFl9YBaNsLOPP7QmboVPYYOLeOvWM4iG3PLyyWtJY9lW4XJLEDSMTWFQtKT1f5U
ditnrSw1BTjwKnfKTwJ+uRNch9MZemRr1EfuMXVJw4Fg1ISKMKVAoILBz+k5wBRT
GqE1esZSTvzkl2ydeFUx//B5xc/j5+YfhQvWq4ksnvq9PzKHC+JCDiioI6G8s2wX
9huG+UU6cB2rd6E2wk1MpKdUNsN2zQQ1oZaZzXCxWSd3UKeaimsRgw3Ce+fTjPkz
nIYkUd+LAO4G4nBo/i3Tn4ISuhVzlB/ZGQorJkX6TbgMPLnW7GriqOMOF5r+1tIx
OmfB4QT5Ni99BIJLhoNkOtMxHLv2uw/G+0d/J77zuka8aJ7wIDl5da4wz3Dh5jRC
jLxLT0LI7QBi8usvRYXJQBcI0sn5D8hxfhXp2vtZimsSeJIiuPUTFPPejPH2yyuE
5m8WbjNW//EsSSJUW4bUt9/v2U5MiGyLP7BDf5a6b7azPp5boB9ums/PX5S1cbXA
JNNd7k8k1ZXMin30Hbvaa+zsGeoSxNFoje/3kcHagii/boeduKOByw+abUARVKQ7
H7qfmLFxeYClLakiJOw9RqokJDPHSM+0iMcLDbIb9v2cFNRo3Fmpe21LB9W7UHzA
54Zouy3geNZTQb1hya77GewekZN4JCsmawwTfPtaH9mmEuFucKYjpvo+kB4M97mF
bO++bbQFthry64CKVExeuy6IwmPdJs2C4f4ZyOqNWPmFsrZZfJ6P2luXToaNTima
0FJXIdeft8w+8bpbO27CD+xxRTG3cbj6Xg7Kd+7Oui25l+26HJI2oq23bEGkEM8Q
jQawlG+EY+g+YtHP6GKMhMlBhybD0Jb0vf/Q+mwiwQj7n9gcFnrw/Zy6+eeqUKWY
glJVsptz7go5zhNFz/5qh9Vy0YZbAA7Nezoef1fQnALWwWI7FNomeZw/uVAIRJDM
rdqIRq8ZbmUcjq14aWxu2YPMb9BWjEXIWC8QXenclKbExnxO296BdvYtJ7DsmFat
Z9kwOP9yShOZPWvH+CHCGBix6lUBz3oQgXbr6gR555AcaCb3A/lYYv6vltMujaxN
FQazB46D54k5+mo0Zrq4op2ZKmGR2nxBPsChrtiWs3GQZFeTHTbjeqRsWN702XUm
CDAn42SmaAto1UpNSHu2fXH6jXsIGpGe4HmLb0OVMCrf4cwDvjPrHStEYyc6hv3u
NhG3GTBs65lkTFGXmlyss6kXjbedRfTicAlW8wJoKWljNAkT3HKDyYv33y3br9ia
2bodht4QL87zBZzN5LJeVkH8+4qwX/gNDKj6ctnZ0D5+Nr+limX20ibkX8YaVkUm
QtlLMEybdd7SeRBAKbTwvyHuripiZGsuFG6GruHLw7p1fYGUWrUoLH0syGCM6c3T
NGFm3rePwlCjDeW/GYzyEBxp8kM20RWkClefTbOutDzXozq5Hxnj7nV8jQm4PSA5
yw5ME4iIqha1tCqmaHEHs3m55iTQqpIRZDrpvLariqChQ9eI7YppYrvXyHRIXtm0
5Y/TecO6UibKwRs2xvu8pnhaIisl4rnQj6P6aTgURhoVkEa6UNhLIsaaOXoh/A4J
CIA9kxNGCtxo9sm1ygw/8yffdLUtPEZioS/v1KhbzuUiJ9j6B19FxWjYGM7kZsA2
OPuZx+OqSvol/jFM6h/lNGB5WZnDTSQAiuCclGHpmPFjJc4YKQROMorFJlWhhUvC
ZnFXqze1XFQfrhzQlQOjqvZTsTUueo+phXVXsQVRCWS7DqTVgQIUPuajW/EQYcIT
nT9LEgO5YJI1YGDJ+K2T7RtwP4kph+f4a0hEozEyB4TnbA3jMh4GrAKt0UwxZLdz
3rt5eItjhZ/5asL6phXQcMEKfYp84u4GiC+KPFfSeAUrm0hq3v48EVNSWVGjmb5x
L5OII6nedc5UV2+mWxui1D71koScjBBIudABqHG7PfgRF2dLH+1S3wv+PcqzY1rP
O6Mldzj/BqbjHVh3iaEIOejPbMc64+XYEGgfdTa/CBxbdLqpMhJyUP61M+/W0h+b
l5JfpAHjqCjfKoeOZMC07mkSVh+PvIwx1GBplzYa/cTvRtZrFBbDtJ8vn6vNTsqn
V+Onah0/CnAJJd3rIBsAQG6m73JMdnxcRf/uQshWT9hLoBqCGAwdmEzx1DBbao4P
UDt5iORKPIbUfavaWPTxjwnKStFVZpFXgoP/nbMlTtRzjfLd6QUvpno+l4DmDbqA
l0bksMtkcFgkk/J57LZjhy/76DylPo+rPlFLY7dzj1bmp6wxf4ruh+erP0o6wtU2
rphNHPxZcDpmfadNrgLsAwahkEByGTaNWrR8QSptqUcdTvTKMj9Y2Dd+pODjYE+S
GUBVYe9O6fWYkth97q3O/lxfSltIJOLvLJflbLOvdWGv68GMyrJoYPQa4MTNKqQM
zaibPf6gH4/Ijuq7FKAvOSuQOfvNig2tUPlRZv3sB2b1YRKJQeaQw7D3BNy8HJ7q
dq+yeR6L1/1wxJs3N7R/sf2LDhtIfS6JLpm0N5rMXQayap+V/DXsFka0BS4UGkkE
HtQvfxMw+1nefeVTaPPO9ql48GEVmPZJhg/g2CC2Tc3EKoU7/NwXdxMmPjEWlu5R
NEAN1Jsm8FtiAzK+/09Ae7CDjRTjFx7bBmL05AoeViBVZ4VGFFb4vcVjku85YFmW
p04gHthNmDksVycGDO5LwW06SJqKFybr0pwRJjIxOodKBcj0p6ZtiezpRAOFFz7l
Z67liNooP28tOoToMeeiyEUifY3RrRKdOjblQy6rdy5dZOCrRi6F5yW5tAeCtgys
BPotRd2afAjgrPOUlR4Je6LREHzMN2uBUE1rYpi4DboiPTdnMe3mNWcNRCyn97Lb
Q4b+kV8uN+zk15sEYngHAmfsphH3+3Y6Ll7PIUSia4D3OZRpWgMBbC76Qz+X5naF
Knpq5S09EZ5AtKidG39/jYt6jkFOBBiCmSK/EzUTgBkqW+ZjxStPXbYgKGeMCode
rlykFp8LvfN7B3X/F8s7XXWC8aH2azTSABNksugHYkS1qxJEdsZrr/s5y37Ko9yF
1rkgqwrEuuHYApCt6O+teaW5jqeITJOBsZNpIiD33iHuOYnBmrQwinpF2gVw4XbA
WJQlG4H50ZR05xRy/zstnOCU/DYaQHMhxd5zJc5hS6WUimnu/0B5HTDa5/FhLlqD
4tU1xkc6msSU+sxah+GkTQ680s1E/BRHcs+vaw2gpQ3y7axUG0cyib+ixixIAuyG
SofePXMmOe7Bdk4jI5lhnEBTOt7yF1sReHPt2V1ylVjlumhdBG4XzDPkQtP5tolJ
uQBh3X2eCYVBHrZ9HIdyEavaUS0QeVmWKFWPQG6riz0IbIXJiDUkE86kX0DHaIeL
Va0zAPfXUaQk2YUFdTEyeJSrXx7bwUPUve8N5uXfFOHW27tToD0jXhXD3S3fC0y8
wt2EmZQf33xB3r0Dm3QG+D8nRiMmGWlOnR16MGX5XZJYIfB6SBjkQt+rVIsbJtHF
sgD+1tbtuLvnkUOXgKmtFwgicRti514gs6A8HdvSdOquRxFRRbEVn6aP8L7Gzk3S
M2enldzjzkTa3sYwzltLbwKXx1ERjuJrZIozkZNFbyTB0d9frDPmszcgKmMq8FVH
zB2uC0QSr9T5cUx/k1DUML97FqBCtucDTaGdJSYWeobsT+hHXk5rCPhjC20tzVGa
jjRb7R5eOiDx0u+qEWB4o4dwXPwSR7v8phuomt/b9p82RLU4GIlM/2u2igOzHajq
6IxIL5rZL4fECuQwnYfMd6FrZWSM4RAU/QROQVKf8k0eJ0/MxRZjnU9t8afe67/U
lf78oneUf6jlthTT/Uv6V/5Tg+JFPJWDsgQP97TvEJ16C9epU7gNhJKYG9c/cgdO
qkbMdCnTNSQ4UXiKBbxh4Mee93mf3x2rDaGeAPJbumDsLzGVIW7q2EmeFPz954N0
efr99id/1ptCf1ocwV6LQ47QEc1o9z6dz03lHAFOHE84dRyVxz8CUpMOzt1+Lw9y
fUm1xonmVksG4VQcitqU6lVTnjPSxdiMWn58ZPshYZvkzh1TCQCUPlzjVTGdtPuN
33IuqrzXDsnOkaGJYhVVyenFUCUuY5WhsoikBPNsykldxJNkjc/7gxdrHt+nmiJS
xEUdQdb0wnmQgqKzlxk9K79fLPmDw9Gw05KKMY3xALJvveLsuMQlXusLdQVPOHG0
3VJamRW/w0OWdfildWUduUxhH21+juK2ijK0dWO5adAHK4lZzHGBf0lMOF0GTDKw
Avs2BuObwx86K9Cfu/sKQsr5F3UjqpmyXlTdCD9WUuqA4d0APSNcw7t/9YnUEN5p
TFKYOuXsQ8xDZ8MvW5ct/MBB1Jd5GlG8DUYsVUtXaQnrehCac4mg2xNg68iMh/9f
lUz14jXCXRFhXGH5RtfgNb+aYVKjkW2YI1XIKWQxRCUUmbp+kfaguc8lCYiTtcfr
sXQlhtVw7OK5BaHpNC5ufQcnsRmZjH5mlXOZWo0dj1IFajOZTrfVbS8hwBba2W3g
1+pFVeHkvs3Y4mTPqXeMQX/dTXLTSGY/8cckP8NIR00v2D31wE1RY8QP2pQksOOB
wbljUvTj0Y1T85rgG0WdsWh7hXskcqmzvb+YdCR1NquTNOvtcvacUCZ+MqC+NYN4
+LccpzubxZOtZ8IgxCIE+yk3kKVpzlNz7xP5vtAFZtwDuqqWpUipCslggmYG0tHH
DRz4wh9rTeu/4eMvxSRaVHWOT7bESGb19/exKRS8tdTUI5JUl9hBbKwuKfIRYthg
ubKE/e9mCOKvgbPFHyxFZlNR/q/yWYK3DqZ1LC/wh7pJYuV7p8+R9te0NTA2MbDM
aJYMPK47Y5X0kREH9M21EHV3A9RQPXXCXS5kGOF0cCbLJGHDHKHH/UHiE/LGnF+K
cOpyMdbczwQ9+cJVbsTAcrGjXP/2eDOywk6yx8HsiLP58Ip12DJEP26Wq0+xDnoL
nW5FabWUrgcJIw1izDoNwuYOiiGwXle02n7nEfJ0gcXFT9TUkKejGK/5tPd1qVHs
1sgGxiZjY7NDotRe+r1RKHBixMjVEk0g0cf/+bBaEDWMJYe1YtjGjVv8qTGngKc4
Hyi8wfPgVUZd3lOSEE1hpBlUqHFs52LpxeByVG6skIXtEKOOF9nLI0H+G1Vp5+9Y
OF7/gKFUCMUZaUsb1yqey8IkAJShPjV8CtFmogAbRMr1ELfU9agVeAIqGjb/Zk+1
i/jH3t+RMFoOLCqUGK8lIOi/zYEy+drxkM5Ii3Ur735r4xue6Eyem6bcqU1s697G
6+0bITz0Qc6H7inGkNGi2YwmD2vD5hxG6io/DWS2F9w=
`protect END_PROTECTED
