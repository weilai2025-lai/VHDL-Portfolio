`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8l0uYw0BaqiWSgPmq74QgE2GjPYq88fzO4YS3KQBw2G9m6aPvSLx+gfHju6qwAh
WTGZJVzdr9+Q5KCSglYpq9k63ZaI1q7ujaelsICAttTWKHmSbpTl42pnjG0nWDpK
lAwF1arQCFjsekiX12Df3vQEGbA/BkYc6Itf2Tqru+0xqPCL6HdDOnkisNJs6qcT
WK3NIzc+ka4S04lKOj0gc55ldHlEpHkYM/yPAVATmy3F43X+2nMlQGxaJaIM8QIc
Oqz7hZHPlPKBrzmGPhOlReyBlhXB66zvQUcj0xNI8TehonIAE/eTCffwyR/QEaWa
FCQHZvfNxMZ+RFDohOFGdjYzF1dgx6jCpjx7eTk3MiAcZc3SoyFNtpdhHY50dYcz
nwF3CFckxR4vQ9Ta4iaB5rpnXykyi3TMWmDGNPNta/sSA8qvu5I6yXVfGHyc2L9H
DX4baP09qpIT7RBvhN+nhJjm8JyBvfxncRJWSmntT0g4O+Q8uRTmBevgT1Ynaaon
Q3pjDDEfFCTz3aG4TUmoHXKg4HB3PqUuYl9bORKukpAFPTPhaNUNRUYxZRMHJI7k
bUOEu9sKqHPHIs95YeGyuIx2wijG1jqOCD6zc2Y2NRoM1JlwH/J9ooxaeh/tmHMw
xKD4teE35jTv6MU8Al71GdMX0HSr2ncsPxoC24QkBmInyVn1wgHBvfV5td5CGckr
9UeMsY4G5rUndO7P0hbE++LvB3doP+OGNXIgZr3dZxBz+pvnSzRetGUI6XiaoGu+
lXunp2RQqLjxRCu/YntXJRClGAT9yVywpZ7gTiKdnr+KYVQp9LOO56qmiJ3Goygc
I5n18NiYY1E4UBsoS09FcMnVtyznhanZW1EpuLiXanyHnqeCDOOGHhjeOK1fR8QQ
9GMRFICXNfDaD+UrsssI1k7YBLqmEwLVPfv0ZczyL+1a+B6mSrd4hpe6ZWF315V+
Y36sMiOtDKc2RHry2m/ovXgQErEXepPHouv/nqm6a0lE3gyJM4nKRT8OTeyDBZ4k
2wvxJx2sN4pk2ugGGlx8zxD24NDjWDQ9CddfDivJ7RKr6rI5JF7s9jQyUb/JStYn
5h3YEu3tgIrGGYZkcyRJD19f+Syyp8PPpYwf7OhmG3K0T+hh+ypXVwKbuHcGYVP/
OFTEUF7qK5otmwj1br5yfjsfnMjkfv1i42gBA9E2wiaRBtclmQqxtxa5M+cbTghF
YT1DNzDPvnQugdj/CuFwL16XlzwHamSe7/xeSb0EqUA=
`protect END_PROTECTED
