`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWUC8LjxgXr1qHQBWoK9ydvzyedh0b/6+PQ+sB/w+XQZRw+eK9gWZbzRWfGPgKgX
8YcqQA2TE2UrA0eOixTxVADGEnyPRCTmeAzSj+ALhlXtRPSE3NTwJBWE7zLlIpAH
ozL+sKm6q8mE4z907Lqoc2ya0EnHLSFycheOJNjQlwQi55KvLyn6LJYJ67EuK1Az
9+Lm3qJJ0KhWsO+GtuiIdyewwAJ4UmqQi4MPGo12PJNn4aPFKHFW2uAbQmLKRMDD
ysLEPIarTjFNyFybUS9HdobCGSqJ+rUrHtHhJcpm4KsdO3rcEQyFApMKrl+lDF/s
zu7fwYBP46oggir3N+1Ci9fnNY6+VIS9SPH7WBhVAKjRPuqVkMbITpVIZs2OpMOt
GdqhZ97o9bUh3yeBrVfXosCb+Pz4yWu3LO/n6BW+KrrZkDYIt0gOCPempcKhELDX
sE2bR1E5dX5BtrL5/5UXsDK5ClTgdFCrO/uclZ0QMPmVuxPFM4HSkaKNeg9yLYVT
GuDQOwincFWnVOd2zUIAOWTBMK0gpfLmMQhFlS06qlh/i3sm5onq4Cfnz+NAtcnF
vc3uftVz3cEJRiTF4RrpdXWp/Y0Wn6s50zrEmHtccIjcqR0ttujch6fe+lENGPJe
PZBG3EAGRnVaJEisnjvfGPI0K16wzx9R4liy5mJmFgc1/sRM7AKh0si5rODfFIVZ
99+D6i4ecY1zh36ssaLEVLJ5DcJ2ZtZkr0a1rQH65QBDlNDnkZ68UU6gcFzTvIsu
1rqmn+wtBNMccj0fK3S/tkqXHCz5FBknwcsWSqvFa/pw0AZz2Ect/I0PyAC+TNPy
DWGOe+OVW7bYF+83S1g1aoqL9DEMCxFymCvSrum1RUY=
`protect END_PROTECTED
