`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3xHE3L9ZlaaXgLqF1Y8vBngVNng6VfQCH03JeRS77+/4zINoZStJQWhyRkW7M6N7
P+2fTDMjiV7i94EUai/7ILDYY9VVHPBwWAOOD0ECCZqYf2FQDFc4c5mAM0E7ih0Q
MmTDeToMZ9yfYEreWMKlVmY1YGLk0qUt/RblL/Z6cEmccqvxVLerw9jRKYicB2Tg
/Lksg2EMRxPdFIO3k0hP6zUs2fUzmbr/wZlK0KizjOMWBzKCb8qDG/8afLDwS0EC
bbfeuBKdy+YNcWCVsJKO12m3qX9anbA/oYfe9YJxZJUuEvMerv3jgUmQMB9Q6VZX
jEJGm92gERRoHj/7sMTjckfM45NIpROyTaN0jUcGfoT6+mPAybYSFU1GA153rxjM
yG6LH+mFI0W1FCjgsOiK8zb/9mOzov+zrABcTjt/JkZ8vo/wA66c3XQ80PW7SAsg
Glj0DYvLyLRKeNjTRIsxQ0nCC+TVDVXwNKnBpDf8JXUrATsaJSf3dm3JwAk3qPIz
6f+D9C3uUiLt+/r/PvSp2FdTZKtQIwOZEMfuS5ZBmj1l6vJZKd4Heg16IiiGJOYI
tyFlOFq7eoxR8Oyh880WxZq01+HreYFNDNus7vF2QcyBQDRJ/PVgb25GMbmjq0HM
ojyhPSTapqKcf2UnA5HYPID+ECz9Il4tRHg+V8wS9ZuEu9GrqUogqDQz38gZP7W1
q8Y3PPSavFLdm2gLLLO+SmntW394XSZdFrHGdRADUuFJ/lxWPLIEWktRi92xr3xy
qGnl6t4U1CK478/LjN4E6jxhZxjozU8Isq/+rmn7NREnJBsI48N5yqVOJKXTc98A
gzdr9ErcAD0g3OhL9YCdt5Bdd4G6xxmrmQH5TP1q4veY5ZkLM5URAcY0SCJCdaUt
N2W+Qh1JLAjeR24sNA0BN3Vc2wQ376DJXiOj8V0gM9vepwCNcyCbVV5/H70faI4S
KoVJ7gB2szoVr5NPQRdiaYSvnrEsrVgpRfDB2YsI44MOB87FveInoM1ujfzpdeg1
RfzKfhu/eSXhc37RjjctCfcQN00OLeMkBcjNAFyCXSnvbnaut39EZIySKjORXxzK
xYR+NSEDZmw3ee3iqj2hYNba0wt6RQNkxQrX/uTdam2gWenqIeiKNeIyXFrZUIcw
Ki77EGLVEZ2hsT5coqXtjUMrk0jKoX3aU/I1Me4D/8uPiLrD2sdxL1hZcVFFqZAO
9tUP48AbNULVNh6r3QIvOPpYJkTu2R+Y9dWjbP2cDCs=
`protect END_PROTECTED
