`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHJgZtimnYn3J0aCKklN2xx6lmDbU4ySdOS/jr1LL8s/EXNPq9Ve3LgCY1csCdFR
aaIaS/52BIqgWZt23crXup+1vq+ZCb+n8LFf2wnDIKZtKsH/bfOPA4pFz0G0LBXL
uRGhpZuFRmIk2DRUZpdOXWAi6yGKrXZIA9x80zWqcyrpCTqhuxxD+pWupuueGdkz
QhAy6seQpM2ksrD9aFRL4nhvVWjTIS8MlW3B0ICAe52xaCixZmm85TvjoiQf7UoF
EQW3iAC+1+KbHKyuV3VQfg7rIBXGVcUB+yasso6FaF5pin4NlFZC9yzoVsv/FJ2r
VBp4wdZZoHpcU5PHmuw1FflQto0Hu4My719F/LyuItAoXH/3CZjp214Q8hncDN7c
WJCsXZQuUxKCoxMIBHbRvUWuN+Ag2Lxti76YgHul16ZAMpd4WaJArGdh/GVLiMPH
6bDFPgsmAYYvaZ0+sipU36rb93xGu9LOFv08U1L9V0CR9gXVo+MKbu/2lllXhpq5
uw3VTc3jcJoh36FJx+17r29B2n3D7ImQmgem3bJ4GKdVefVz4UQ3tPUedrqeLTH9
QfAPxyMvXOTc6x6W1P9HXtTGC9lOJ66vLIHBbmAQi4VV3Vfxw84weSMY5oud+B8s
w1ET8Qac4GtxPakygDWaIjCdqH7o/mYWjUM8EXXrnLiTA0Yn6AtAhfgmG5IGDPq4
QSyUPYcTyWaF8barPs8zVbJMN0Dw3X/VTljp6fhMGSWUL0ZftkUcOkJVh7y7heCm
ivZvTld/jdNFaxaev0/4ZSKlmivJt8gbVinZvsGIJ6IAea2GYTQKV418ZiNzWIVs
6kwaHVYoqM1jEHwe2aJ41TnLGrBsns0ydGCZ+IIgom1Rz7WMfJcFrrRtmmA2b2Dh
r/gBRUY0OGIcrpOl1GyRqDYswRrifNgc7rJeZYqeAZd8RgqTF1iSFGF/NVUTjhDD
cVA0WC5cGuB3MpODNR46cCud+SO5OlkXqaAfXgzrxaLbiTQJR5fgaUZunYusIzaL
zhnmIYyrsYH63q9m0Aifl0UieK2ivcIZ+L2V7VKx1G2fMezdnCy+5quW+MVka7dg
61AKvEGDWNZZHfV1MB6w6Lp6q/eNC/ssqsLp1PvElXu5EDkaOEA6qQ8bZY+JKqwm
UhW8M2yQWdllNKQv+6UKyZ1Db+RX8yIKoc+k9d4AWs7SaCZRaJYx1KiIy5al/6yI
Mta6sYcBmUJYSl6Z/EJrrg1LOpmUwLaeT/aHGXo4T+KEQVFGAWYMdeNvA3elS5xr
DTxZdWQozlwJTx6PawMLG0/6FK6hG6lApBydeJGMsOzAfBPYEMIKGe4wYEf7PqN6
zUOLiNeh5lSEY1YG5jGge2lw2AsuVHFP/yWxS+6lTuOm8/WDFPEzDi0tWucoymbw
8Kv3nONdxI52DR2TlTEOMW2LIQGTFTTMk6QTJqAIE5GtIG0iMvNF623yQe4ZEw7C
GaMazc+Aip3kCMHJ3TojDruLfFv9B9AUWY+h4v2xhIPnrMr8JAVCrqLWzq/RnlgN
nwphpeYKVaA/pF6RkA6btGgoBULtQvp14QpJMuPw0Sks8jET7KTV+B9k+EoHkjSX
7r9Vv/sl1PSZq/KD2UjArK++bTTXwu0oRmMW7F+R18W2kbXDU/Y+RRAxeO6WFEp5
PAi/bgmfOJkVYE7o58T9s6I5JlU56JngCoc4OLGaKIs+A05A45g+vA0KowcgGZi9
Pl0UZtE6ilW+yPvo+afXlhiD/LOm5DJLbfMnQxM++XOnokTjYx5aDnOxmWh8R17t
8Nwm2quF+rjnabcjGNo/l8uKf9BePScHDgVIr2kJ6ye0WhrnHhpXHssAVmDUQjYq
x83joUnZDqIxckRYklZJz8rZuKlk8tfPFZTywmIK+R2iGwUGIyjDhKRjFZFUiakM
EWnQ9SIpO42/CJVVnxfIjaT5o+5owSmbgF46uQHr822K8Zg2S62kM2DUMsEPBPuH
gtDMPpEN+UCDukicqbYwEMVaCmRfnO/mwYDHAgSLUCN6FgddA09/C5yndv+HVd42
L4AbgX0oY2Pd9q/NbvAIldC+DiCroxYtC97V78FViSYW6CcvtBo4R28ycSo0uppj
TEt3p0orTHhJRtSTtQjaU+YaBw1nkdqRN4I9mp+qw/KT9aoeE94/1vhA2xXz8Dvd
ya6FPyT6iEtGieJww+bCMOTRNiAmynC5aoqcaErXmu+woQSs3Ksxd6q8Sr7TODKD
jXe3ROoieLo+sgIdnxZ7exhaEaxUxhe0zkaVUM/o9kwzumxoaB/5mCZ5qPeAmksg
9IegMprBrAurJvwhFQMqiqOulrMG9944OuaPagRXPRtclkoOR7Sa8oUwwBC7yuwM
kIMU380qvbt4F7kz6+tGryRIJ9n/Br4y6XiKZT1Tlu32zUngPWLL41v8VFxjd5Xn
er7/2b2o3chGU3H6WEIo3jjLL+4qemcD8w96JaIai0Iqlr5Ms7/oaEjmDP/8xj6C
Z/6aBF7d/g/5Y+mUwHAXcT6+QuVBBzQlYujl88XEe1OePcSsKsO5G/7SAuIIyxrS
w6q2h09M95cGHF0V1lArktnLs84WoYXvJQgnW/WMnbPx4SNQkwxs4NOVvsoXSt59
IW/GRkp4tEo3szs6TNLgertWZN+5SWjnAXsAq1gZzkRLtOsKxoQ+F13Ai79bRNRp
5mCYPgSR10+CMJnyLLLkLfCoo7RnyBiz0aH90FKZznQE3qZtc/VisHYoS1qwt4EC
8DBSuJw4jH612zRMPvIb1BYIocpE5fWExmve+kNSTiYJz6q1FRXtTs7nwnBPHPc7
CUHibXFDa1FEg17LP/2CyLsmQ6+F4xNVBx472aggbNANB+v6dbm9MKdA9zo3ifRi
5XnqPqiyEbc/3xThwFPoP6p+7nhK5E/dTLPhI4tqtYUeK3z0nV7X/SuQbiDQuDXb
66Gc6bxB3NcDCwbXCXOItjF5xHU2j9txS6P8NogCIdsQzUwHcnvDmho/OluZPHGF
/Km7lJcGpsoBN6kHpKYQAIriew9kJ0IEHqoOcDsBtFXl1/PDgzu0wyapkiFGSu9C
fcl+9JsGo9N28uWs5vwmB+XSSa2ps2LYmXZGDGIrvq3vJ+ISNzgfn66RxjcIoLgJ
kA9qdPhF9s7aF+e9VoHBzS27AOMoEiD0ccku8qiIFNVCZG8l7R+c7Sp8J3byMIx/
CMSpcOS7OFFVkYMcevy+6+XxmJOW0FBwAs6GmC9PwAKfltHAyRZzIqQ/3HuVYQ7B
Y/6W2/Rfkd5+xojU6XzoQjHgP8bCyqlumPDih3eLaVG7GRFjVwbfQNVKxPA6yftb
RynxE2Y13iJ75GSq3A90syXfKg9d7Ko230X9RjIaByhJVT8/O18bgWVlv6regHg/
16WdE57zP1bMs5KWjCOENGrhma+wkK3DiTBJznyNxIJKWwNeml9ZvO32pbiDXKJQ
9NpuvWMEJDrXTznTBfW0ys9jw/bXOLC03LeJ1DYy5CwSoc14mSCSXvQFeGuSAVMd
R/9YBqwli3wV9/wf2U5QkDZCAEBgPVSFAwiewfQBjCfaylCj6nc3RKFPEYhzqyVv
5OJTufejc4l03ujewqyvlpi3fLBXTPSSfbSNTZkgbELTaKehWVrHDtwZiYeCwZQr
Tjcdf+NixBsy0U/twrA/gjoWPOLGweE5PL9JFweashTe90Abtnz5QlcFz3LdN/8e
UQcTipHWDhtylvxdjtMEteUGnL1kRtge3rwo+1jRxAyup7himCktsi2Vhy5ldIls
zm2l4mnsuy/7qqYB0utoLRdAIV83XFnaZafDyLjKAGSlzzKpUeqDRTzKY6f6smoO
jTqCnt+PrMhGTQ4fte4BPIw9sSpfmErvk6hVZWAs0VPf/y+r/5wLhalCxgUWBJcP
8JHUpV+e68cYQ79H6wEGmlBJA3HdJFdB+jhkibxrsuxXUzWLABXRt/JRgr7Nxz/l
wcXz1oFSGfNatKvTNMIKR990AJ4JC/QPlubsmehQ4TsdL4MRiHnAMakKJkhXF+JE
LqNIZUIf5e2ulIog4AXFF/6TwvZ+davFBYR5G/DoLrNrywaGICwbwrbyr4T5gAP/
zDNqAroFfbiPBdHW3HwGrdNygweoOpUWe3Zk7yWKpDu9plBytKIUfEW1EIkgdT4M
GxLRUIi7PwAXdZo1IHhRayaAiSCavRU/aXwTaO32MdAl9/mix+ghnRx0A0YZH2o0
gb36RX5iw502W1mV9i4AJJ2NpSduS6QzlacCHDFSltJ1+QsQu9F9EpyIfFmD0j/z
vqpACe4immwkzPVqLQOxWQl4Dn4SB9IVQEwfiqNaug3/Go/0hIt0MRxCfMOoPiaE
482dIgEXrhNLTxdjCKKyDQxC/Qf0ZHzSs3jhhA0KMUbNldF+w2c1YCkJmTV3T4x1
H+cBixAgBLpPu95YqHyZ6/BkmGnvaDEVb1qE56rRp21DwdOjjTT5ixqmcUVLUjSl
fy4EilQgNBZ5/mpQrDWmMofj5XpuVTJ4V0HiqKDG0EL5Tlpj4lkR2WZCLQHNh9a2
vDUG3LKVkp0msLWbQq088Lnh2kQjig/e09Mf+jWly5NQDpCXJPJ7Iz4/W6kJcolx
1+BpARZOUYnph85MHQ4Amkfx2rXcqcdEI+HN3cU91eeHbarInVpupaZ/7dJbhvrT
WUljGFEajxnAU/cVY7zCMAAIXiB6IIwPChgqbKCNw9zPhz35MHwXJUivoAOztbuj
uCxuwJkbNiWmP8Qv0CMxTa59VuN3j2j7irNE660XkbZZwvN13pnKy9zFXTRLA5St
QadW8BWZyd73ZNHF9xdEhjN9qql3RT/7zvNGNUarQI4pz6mpGEwV5enOsbr+GG3A
QPcihcjIvcr3MxBsAAI7DuvhWb8Klt/bFZXocokpEIUKKlCKSULLJhmHi1n4r6cf
fkraHbtLQR9S9QQr1MNypH+N3nzMZo4UaPnNYwU78n7nfXE123yQ5eRJXSmARmvy
BSqg8F9SXmRXiowl4ESBf+lUHEqi9Ag8NFZsmyehSVSN4MSIx2V+84Q2ITWoIiyZ
SRJUjdy+imt8MpHQOPmlF+8X8Awe0el/WpweOi7zZlMwZ/2LYCafPQx350pmdyN1
/l74PVM5SH17yz3+Q+HYyN7ezMISycwWLVB4MM3dxHvH5+MJXLK106pRpRwqYh55
tXdCqYI0mfDSdYfuB+bHT04mjebQBZSKjb+LSA3v57U+ibbvb1LD6Gj9gHtHl8GY
+DPm/9d88I4D0cCfBxIueyX+aKJ7/57tKIn9A/WE3O0gY0B3hWE7GoJ/HzGnzabk
1fya3mOKpiyhxHfCXA/bFR2kCiK6oKKlt/ALPDFGXJAXqFGK9hbA+3+tr8yNa5RR
RGY4vM0p1ItlyPxx5XK505UgNDAnVXkg683o/v6UlRtakmT8kpexIxrFDDXJwMse
+CHnCw9lbEX6m869o1HaYdAdr19utI3PlPoNj+O7BYVn5bq2WM7/qrO/s+P8WwIU
28Gk/mB9EN+67Dky8YsSRw0/L+HtxVuZiMx8QWzl1FV88QYIZcfutSMyYD0NKNRa
yRvw8yHftCnQJOaCeyKhD5hiqfTyIA+h0n/IHaaRV/LGcsF0imNnamKiloJtdMeM
oto05B7US14Utw/1bZ8FL3EmCc5mgQUQ4H9QOVNaEY3HFvCvcXAn+cMlATRfTYef
cCQz4cVH+voe2lD026VnDfuaOm7g/HYZ7/ahK9UqWcu2Sjf+UiUQFrAADEOm8aJC
slly+w0JiOYnsX0BPbDyeV/MEq2DHVHJCSnC0tdJKom+0C+qs4ngQFJ+qMM3u5r+
YXfimxl0Jcr60CEzldMBeEjJMeVPK93nScJOsO1QTKMp2Yfm+7ilpeCDKv76iY8A
l2t+8iBweNKo2DF44mndaNMKCdrYUfGF+796i/UJkIfiCQkithg6QxHr+R8lg4Ry
NMlH8TgVWvAxOxSoEESHZT2e0UjJ65q41kB1JWE0Q8iZTTwQWwbqCnyALcxhdfB7
rhoijOG7klMWl6mHJ1mak/07dvT0ZZ87pS5djqpuqYYt4aO4thuXeFOwyd5b47jy
HhJ8NhSEXLW1w1AYhDRN4njXJ5Qrsl93qWIXHbjIwxyJIv2vNPmpJ+m8ODDxpspK
EjeCgLxsS6kCDhI0vto5t2IMm+s9wsAjAlkYXBs4rgbhZmHJ6ToiPD0g7fMlsYoe
ORlsozjxEBD+asfczAecvW++pjRZW+N427cHJ9HL6rqexMAlt5FXo1fa/c72DVl8
ZWzqp1Zt5HS8OJ8g/W5FVgOl+GMUPawSBCSmAoJmpeQ89N1VFXKwRDmqRQ604G5F
u1bX77+PGDoN1JANVjMi9eP6PYwvCiAn4NIWm7RYAsCEQMsXCnLQqaPGdnsS46T7
39wBcegQT6JcruSMOt8HxHdyqtN+zM/pKKUt2T3Uv4itpSW3QnJslKvOvr24nHLQ
WkfjT8tFnLxa1fts9NoyTpGV2Lwbb97+AuX8CC8of5MqRg0k0+7FpjheVov3Q4Qm
qKXEwdbdJhtbtL5qzcs9hcC6dzAscpqAGxngas5xeEbglrVv22lvH9vMdCiRtGoq
uYiZREwasdr+703jXvkmtK23+NDYHHOq+ISoZ51kgnNK9ZVibEhtMwIJPO4m3eSM
XkLKImoH7S+6pFi0GT7uZQIZLC9qTYC0oaXZQeytr8nePJXsjniLfnRQ/GJhbiot
1uUPtpe/diUEnw2n0RujdnRK0qkLzx2SxwbsN5w/uLCm27lTeMqyuHWBs0QjTqHN
hWgasT+0M5R2DJIdVRvjm9kolk8gFI7qtZWi+yCROlWVG/i7tXm7THsTj+EK3dz0
nQ8i0HH3zcdS21eLGirJKHyrmLKzvSVPbNuq9LrTt202qPbGuMALkH0aogFx+L1l
ZWDTMb7L4sIveYYKaQ2RJ8cx74hyfuoGSyESsNTWcazD8BUqSTxs+rnZgnQbwiEX
9SK7AL9TMLFKFJpTMFXRJ48nXCmFisWM8UcQj9zaBlcBPPfzOTUeFxfH5cARgnDo
Mh3J1JM2SwH+Q2FNcQDgg3VlzCpyj9Kx+XdwsUcDeTXn0uJ54kOZFX7yl0emNz4y
UQCobuwo64PfGByKVS/7766lIB1Xdqir9SjmLJ9xSYLgHPPsW0yAGEqaIi21CF15
tmI+vcZbZGvPY5sLUFHPCiX15uc90JjuqQ6W9JDOMNVCtDJn9Oobvys6AeJwT9Yq
hQYOHnnIyVD1z40Bp8NoTK9RM/YHFgQKElXOj8hehaffXltRijh3ZPsmByvP+pFi
vCdzAk3Wlg2y9AiPnjraDuY3Zntwpkw21UMU7wn8torstDyJthX63sQ4Up32R+7z
YD7+enez0XDbJkmzWW+USzmCGYUg8/Uc10LfvIRDIS1LiJ4/fCXWowxVwLz4gmIC
VIJDduNPbUvMi+Wdtp6bTXwfu8zpBUPoAG35TufPRsr5T3oFa4nlsnoZqvOcgll4
9qIjbUFSvUtwI6Y5vtFpObxBM66sBA0e1jmy2CELw5lSXQbjk68WW93hmyFLxiX+
8w5u1VYs8Ei9dwmU7ZgoBt9aSX9cYV3AD0g7HF6Qb9wI2dk7bhcJj5jUwc16rC8R
Wwhs7JH0hDdzeC8nuzQDlykQXoLPHu+wEX3i3rDGHm+s1t2Wi6wRTa7y/uUd5hvF
+4GY2Tv83ze5+uZ9lMQF0OaLukZvEGnWQ22nk4jfBzLNAlck64Q4y7UPCxgHFkXE
RybcmP6k/7FyOCAS2QigaZpPwWVdpCpJBfjQcD0S7ls59VfdFUUJtEsr/4twkzoO
5aYPeH1JSYYE1uhoaiMpjfxMNcZTxmB+iG/k1kUPv9hKtkX3dY5IobWNtBenYcIo
btjvDC3EFFIv5l+sCWHX1tiWGbAIs1Su7IcIgAQkwcTijjAjUPQGfKv6dpZPy0nz
morhXZUfS/wJ79a3E7viiCHiAfntvEG+4hWX1casN6F34DfNQU0LGU1pFdF5+kWD
xuQBuXOrXSaH06MV7ahjRVhbyUylrgrFf2zN6PUECakje/HqjOu3ON5sSU3O7S53
E3GSFWo7bQaBVRwUAfYnqa7Jy8yFxAMBdepkWv44Yho2rH0+KscbUd3MI6YGs/Ir
ONIYwtx1noyd7BidOdu9/QvX2hj3hXyLcCE4SdaRqGVcB+77l0KscbeJz+HHYbs5
qSht0/2dtyi7+YnqYrJGm15Skv7fYrhgIX/tG67hPv0eai2ScwRm4OKcmxqcyrmh
+Xs/nXUS/1/Bhr46vfqiL1yeqsjqDmrIZEpsZkKP0gEkW9F7y6hYidXpiC5kxHIs
hIoVf7+0/zaW+qRg27HG0SmU3suf7rRAsTQg286KYvO5FvSYia91+rADSEGeJwCr
+wHEEOTCgzbanpVL0YWefO1hZgC0QtC0eSdzqi9zn978Q6NJSDWub7uo2kTbV11W
kp59aR+PeaZS7r+iKEeWSsvdLHCvdqkYaToOuCyZO0j1ferFDEQvOzLfZR6SMoOC
eP+z3z4hg3OQmaUu6UbT6RUnJfcSvYEltdvU8N+jTwJ2axm60KFReh/I5FTa1QKs
P4U5IxsNxq92tYiz3mEfNWQGEhPfP1Vu/OAgc5oncz738dMQ0Hgpd7+oxppWL//j
JpWAIOvTlRFO1XYQXtHMFQ/cVaU7+8PtK5bSidE7nUnXapcg6Igq6fZn2gh+BKKK
AG725E3DNAz1kbJfs1z4HU/RTs06NsVdWUCG80isS7HDMgLicauHVxBY0cYFuy2g
hoezCmdOafMRUK/hiD8GHGeztUqIYf5yR8Vm+eLfuCX+O8PFBlBKkuENrsX7gUdj
/VBw+ar7VeTPGoPN0+sbSqC7y/ITZKiHOA5pQjrLbmUB+NNJAB7uHkkonFY3KS/x
0AxKqz0iuHTWRjdq2Db8kDP0NuWhCxhHKpSxbRKMXGPOGVP7nFo6qfb9/RSBM2mS
WqNkEsZCqBvfcX2q9B+8s7FA+RYqL9Tw7mveTpUQtF/UpiAaCHsd4HHm7ju3nXaM
AfCjR3rRRaQSROwPCk8aawrWRYOscnDlSuHW6D+kT/SEH9EIv5m49boeNb8LsEZN
7qyMyAYSTvRPXJL/7WEHfYfwldZ9UhyHDSp/P8E76nMLemdrM7Zgg261ppTz/T77
3Wj5jdDDXk+7w9lEuAEJoZohUfWeNMuVNVrE6gv4l7f3tsKzm1UnFh2gkhbv15Fx
yE85vLon7/fMx3vM5GKG84dHsjnxJsJ3EeIr0Lw5vy1Jf+L5GvGUGyqUy6aqqgKh
+mNAbVwsW7nDsmgZbh50hI3bDtD37+Y+r08MZu2gnYL9uQ7692+yMbxBNbTJdxmv
oQjPQnTtT1A/L3K3NoyjuEk/ITUPHU+tF1MRVvy1BLGfaJc4zVAu5vjXDDl+hyvA
JNy6waAvCLqi4sc76ZpJY/yi4jJaj6ItmqPMtJviFEayeD5jnlsL/sbVULakbIqU
`protect END_PROTECTED
