`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eiV+3/F1p4EMs95suUV/IxStIHh3kKgf6b86ptMfdXjRXEuDzgEaBycwF74WfcW8
stDvxIrniV441YM2Z4S02Yra6oWH+YJWQenQe/j+FDZTNUId06Ba1JeF3Rcanzhq
cFbBwOVUAyn8xonZeFClTrUakCy3yOQ5hiZ91JPrMM6Fbtre/QsXNzZ+aMSMSisr
OGh3kT5qowJMoLf4VwaBSVE1xrJNH1mcGtPY0wYZmann7iwWChRVDUj/KT06/+ZL
BCLlo2gf6XYuqQ2QBqOa8Rat4VlPV5AVBhUNlVHMV2goZGxf3pCaSbvkBE2FJe+x
u55Qvp2xb/UmhXGOtZKYjJgVMkUS+0gBRji6dsub9VSkuVfKLkzMwTM6Z+KzEnAe
2gr5bIKPCxbu1ox0hYZ2Z7whueQbH3jDv6Ekit5lBCkK7h5kIqpaF36+fhHyHTmd
bYBMLXhN0nfFzhzPGLl76Gc4jgWA5BinkKPI5CFYkQQP3Q1LSG7i1K9OX5X1rugR
uixE+9FAwOO4ZaC0x4/EJxad7b4/Nq2PEMNx+lkq3/Vp7vIqVqQMpg2z9gInYflN
btYD25T/wNGlROM70dC/KV0iu/HqcTpgwC0BrDI+WjzvqiOnMXTwukl7DsstdBX9
RXsKoYvAcCWyKrmW458uytjfvejttjR62Qc7GhtXDH6fGDYVPv294cTWCzwQ2Y+R
PeGRForqi7NWmA9bBYz/1oBIyouvr3K13uQn7run8y23b5Sj1UkDjAqyCXHUG/30
I4A0hpmPLamNGV6kFmvLHhg07sb3zeLSsFMog2xGrGyoE7TOKQERIukzCNnXgLUH
YItPfQZeZ+8x892dafrhQ0DyLGhte8obAOFYwzvQO8aW/9G+u6du22PLjoNnd4Sj
4fMsXrC8YVCoaWmGXX23MQMa8R4oCdph96wk0jpEa6GLn6pdTmmC+KNxbob+rIFq
2Q37wFTQnKuoVgznPQiW3h0SlB+oyPII0WV6E06L19svJpVwgWOvZUciw7fqNRdi
6k4rp+GUgIedK0zqk0ZZojbbq9TkR7EE5xaT9bV98bSqYMb5PAre5HYQSC2gks0k
uUVTyDiPmF0qaj4WWJfx84G3OM5hAYj+iTo+y3zKq+jUVmm8mE0GNnWTjEx3M37q
710kgBtp0POxjgyzT0mxiviANfFRsMubNrvrCCiZ6S7td13A2IxYvDYo4Yi5qDHo
3WYbhYMSCeNJ0ZJityOhHJ9d1H8BT3H3SmMkD0lbrLLFH6bkKQZDR5/G3+7D7g6t
3zIx1zeW82Hxhwa2F9QNA3r5Cz/Q96Zc6vpm0Upsih6FSN/C44bYXZaLogiaf0i/
zt5dNFSTZSYDR/APW0wPJelxNhbtvwxWpjhSwB9KRm4fSc7wdcLTruO7hV4NdC8v
MXeL56K9DxXy7+vsm15l2ClVcBY9sU7xZXkbsbrwrCTXsErRPtSSwy/sJWn8DKz2
QPYHM9pKvjAQj8oocHv2HEnnfMZFQO/dPqtrdt0A9nSAqhflBScYQfu9Ipy0ZmOC
nJNpEFgTFxsBDi0V+4LeRrgqNUY2hLT+wAXi+6qG6Nk3hRSPU4qNq6QHqABpPbnc
37XSwN0/M/SY448QpUVjvPeDqQI+yvXIjrt9UjcLGmLu9gwt+WLO/rLC8UBoi1OW
RMTpykz2n3DtikN2u7KGQkQGxsZm+f6mWb2TK88RPMlJz4C2QQlmMbuqOLyOp7QH
p1aKeD4cPZgQMYPEeh0H0/Yveo2ObfnWpyt6PDKlKJ17Z5XLlCYvCvTWf805JfWX
FLLyyDbJ9U1gispXKaNHj3x/72n2hJLaKrgftIudDaQO0RQKKjJomZjonwJjWMuz
27ClbsMCRCrPv15yunvicv1p1g57uwGwQXfA8116LE4FVrfKH60XKuJIDK23KQF8
71pa/tBISwvFMEooZyyqrp0egAGjqM0ydgLbCtvKTPcge44p+4IGHbt9Ub/s20jA
Y1+7PKkTWVXCgNBxY+oFkEas2UR0b/CvystZu5LAtSnZsDN55MYOx+6KcYv9gcOG
vnOfT8wCHO48b7R5VEuDUzS4SFaWaa4RnKI1VaUlv/BjI/vH5JHGhgUHUtjcsppU
mYH3qrIaqrpJaozc5NKH5tHTSkCkO3HT45pI7+jkAzGZxSFmED25l/1eAzX0PHin
ZnaczSfuYz5wVDGMUoKIXuOrAxRmLaGxPzXCy7/r2cPxlHPJeK3dGNpki14fGtFv
bMWOwXLR5dumS5cSRt+Fl8fpyildb8WuXgEa1Eim80KzFqI1O4AMwmirPDD8JGzM
vzCIH9LYgcOvIbQ1/g+fHUbj/Bvxs77PBzXgDiGKC4yAf0BESI5gl1bv9pwX5OVr
`protect END_PROTECTED
