`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLjhaAoDSMzTXrBkLFBvf/Yk0ZJbMgwpn84qjOFyVytITcMnPvrUxiTRp8gh0vTc
naS3FfVmuwXExEvf6Wc+QbkNtL6vfnSnO3cMMY4Dk0WE/gLw9oslwHFJ7Sosbmfb
FbeAxnQ0o1CnusxoaLUokI+wbk4/A/TBQ/PhszPi8Teklpp+eIc7YgGcaJH0JWE8
0eUYjMlc4NuhGBoXLqOj2rOZEJe0B15w7gPRqgqOto3leuPDwVUna4h36DI/AQnk
OKnKfzoc3IS7G3Ti+dJaa/G6Po35Aby/EU6F2po7wzRuHdZv/e9c+StJmOcVN1Xr
RfJ4mkixJXWcYR0h3ecM1xsizDqkbsNalAhfFZIKD1/UlX99TRkgaJgpLvBRXx+t
bMBAX0/wBEsEhT9k6X5NdxCItYNgIpe4ZUV6Yx4mRnErSRr8COJIN1QIEUwyrthU
O2RhFya93oP1r1QhAbJPbvpPa054kapVbbLpb4kHLecUx6E8vODhPEVdZUTNPCu4
Dfo2is8SSRrkLNV9tF9yTBVxV86M8LQNbXtv1H9EywkE7egaZ0LZPHoqhQcA5zM+
c1lAbbGFLuP/iTfOTvmxD/gwTt+oncEUK3J/dJOZuEEVzjEXBHp1zWsM1q8bkEnZ
7BlH+vljcu0F4TzYt/lE78YYg+mJOR64Kzd3u+O4ETZAsaGh+WhMtOiIJ+eXeZHA
LO0n4C8fTKSfuxgH/YVLZIBVl0jk2XVBYisrLn+IppdOQPaG/HBZQea4m6yrWciu
cJDjqFL1uwpWjw62sw5r4m1l84gXCTjv3XBZti5+t6fk1DBNKw5/WvBmjeK1kls7
On7gfDEczy0f5NPLpzj3NnAXWpZ6boljjRH1QcJ+6Iu/LttLeC3FU/xugPmfooMH
ZxVKuiwf8uEt2wcWzvi7B0/kUH3fui1ahPpbP1wDcTzN4dspeRVHzisAPkOiNXyR
Plt+OthVYt1cuhFkBUIslISn97GXLzFNj8PMBuz+OZEtvFZ78eYqyVwZn7TEpOjb
hEA+dM/bDP6sDGj2mXOHwvwxCC6IyZ+E2Xm1Dkp5e0cKn1nbzlBuBFC7Q+FQppvp
qRs24YhxvUt9QesJjE5lM1YlcU9dszxHC5m+kA1hXsSwFIzWGNXtmo8RAPZJzHzi
Fz2tNPeH9cwNNU6+Rg+JSzKk2PHE0V0zBkr4MkScQo8rpytnFz15LFK512TnuULI
uYk/DemQYQPfll4wMXtS5WTzWqjV4cveUj8XeY7NYkPU4fgyXsSijjvH1rgUPHlt
8ZtufT7Qrqb78aiGSJjj1WXvIn9x2AOgp6f3netWUEkPEqXqoQMhCIFTaa7CkaAC
VV64rZ0CjnIRVMI8BpwIvYiuffwsQXff1ZkPME6N+gps5EMH778dDXpORF8D8G/V
JqUrsWLs0kAlmxhfbYHKRvgnhKVi2iPuQUqtdOYBgtzdwqTa2/RdcbZCM9wRU6ib
cd7NqR6O1A6lJjDj800ZcKMfiYDhyCD0xTUKUAKKFhF5NhaW8HsDgG/9rbDFivSH
zgEAzytUg7xT5n11eUAPVl8axj9Hioug7klXf4ESelZ3JtkTAXBjsfspDkvKoHji
AyRKaOU13NiFcxNIETBWy6fbS53LtfOMmOFdxQhk+UkOW7dKRCA67ToANqQXecEp
Jo8wvpS5hyK5PvHly6MCiRrV3kQFbFxmvVsyVHpZxR5oAxoRkJt1ciBfAr2Rra5b
8fmqx05v0FWMFe/rg4x/NANWYNUOT+eTEa2Or317UXgA9xyMlalGnUf9eeS9euFz
sMOg7Cv3KReOFVLIr+xlU0lArW/UJmCP5sx+w0MdoI9EXBZei8QyQHFgHiFPyeBz
dVjJ2M6Nh/5nRJ0DDghl7X3jjcGiDGxLZJS+BxasOLoAskK+QKKsR417lkrjHrXK
M46M36AeiG0pg3lfmVpxF9TpbophsN4mFaN/FDRDlhDUN5vd8WDUTIYgTM7FodkS
Dy4PMcsdp32zFpsSs5hrvGm0IeK2fpcHjuq+irT+onXlyn/T/jkqVc4KD+ZHZexb
x1Q+VdUqj6/AwMuFQQdR8gVav7oaLupDXuo5g4GuyFNF/Lq4yRrX+K7eaVdB4Wl0
VKfs6Y7/SGUQk26TzmB+x6fXKf/J0sCGxMK96Kgi2GinKnn+pqQ4YaiAps2fkaO8
3Mg8mO7nCqCaTe3DJrDTy3g6447AUYsV1ZOs0SmVRLM=
`protect END_PROTECTED
