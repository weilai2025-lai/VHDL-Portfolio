`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5XxZl+XYuaraUVeM/10KjxnnyoZybULUxCksh2Z/MyvKC1IEI41BKpgpH6Qk/jv
PHrPlm5rNDxShD16/69mkvVPopw06fo4rMccePFD4rL6NKvfe3u91gCQ1++imrFI
dgZtyrqk1FT51aaFgacpYJ0MIJ++h4qI4Knbaz0FXqNu5nStUPevsXJN6D/uV8d0
54A9RXw6QiZVIoVcFLWBQFF6KrRSVzCzUKRzfL6UMOYwO92OR576+WOEDeLCvGrZ
iFmYZhoIlAClG7hUncAU1ud5dLn81mBtXJCbTuettdfMcPwle3VR8JZpOzppHorE
5N7kJYeHMciZ8dlW9qsneBY1oHxgFHGfuFQxa0OrviimS7rFUQk9eKqsi8UKGNkF
jtgN1/BZX2XDp5Hp1vIaFchOAmHBQqqXkF49Y+jXEsut3okrgm19n9iZOO5b2msS
VSihy25Q0oENXxT4/ZfOBQnQwtdCv+SXY19cd1p5zY2JLpXOelHr2a378RY1IpN2
AAgrGaTFqNfy4TzupNnShYQitUfbI7beXJ3zBF66oXvIqZ8IhnSqg73uDXYy0OnP
lzdnti51FjBO1nbVyuInpNgZHK1QiaR+e9b7dLwb3BUnQBTiTtjp36lr5OoSVBps
ttEwwOHJhq/cmqU6LGt97lt4lwdXg0HqmiFbiOwdr2xC6oY33pqanAKtRN4mEtly
WPD/UCFMoUui8YKukt6EVvHIPj/6kAceMusVC02pT/XtEmOkNOz0HSbkB4YcdmlH
MzaOjEnHhForCBrXKoSJEL5jMiUtYwPTEzAfXVKYN4EgbdVMpX8NsD3c1HNLhRBF
jwdkgLmVAkqmm6o2NPbbiLPLFHAeYryFVDg/JYk1/3XiTnkb89i7UagStFp5w5DU
Pavk4gUkCI9G6Df7y2neB8DBlhP8mPNz2albjM6a0mZ8eUJuxFJV5KYoWSt04z0d
81mof5d5B242JhhQM3Vq5x8k4qhf67OI8nHTa3f/S0zJU0s2zl1vkwahPdFL66QD
LVPdvp/7gZ00tE1XC8JKh0rIVmf9sgqJUosZLrfcQOzBWCK4f6ImNlwhnfR6YWCe
lPXqUyL56TIWbVud3I2e+dExxk+Meb1I+qLWAVg8GOeaUspcg6XxvPGs+DtcQ8aT
kStCWiwFJ3s+385pax13SkVkvI1OtkYY1Y2nAkjEG/GSLqVboQ3lhAOqJnsi9tkd
VmldPnNu8UQopeLupcG8OYVcJnRAhp425i98wo9Dr2XbiwKwZzFwcSxoeri+dT2u
mJD0Horb1cq8HaQcVEYmi19cK+fnbQNQMfK68NJAGBDrnMxYZJz9q41WmunN23dH
5ymZUL6hVnZWCGM4Oc/aj07GtzOcftJVvb6yEqiBSy4BGdsUwMDvO1UZDMXKRmHQ
W3DipKhoz8bmKzMk0d5U+vWUB9dPZuwdwifaldCv5+rBMRtfjpcfeOz/0Y0/hZ+H
8QqYZIe7m/o7hkPIJxUiprvKtgI5Zz84MnC6c1ePCLthS20jc5Q0QR9ApJ2kxa6p
VwbvGeYuu09VvsuOXPm0i7zVwAy/yz3S/wBvHxQfCdpHT1j8onocfJOG+bwtqL7M
QS/ARKO78wUCTindJ3Xwf3TuTR+WaWb/x7Pd/cxxXMnSCeH1+mn6W7/FQfNmViaD
N5Dle6hDYN3/Uw5jE4CFFaLO5JNnD/OjHkA8MLq7oqq987ueViWiv9fChKMXffHG
6me27/vlbsCHmGrKNYUs3xn02lKuiGSaZ69iGDIKO7SnflyGFb76MuF5xbSUl9G5
73QBCN+mGe8bWlojbXmT3BsV/0OH6H6wF9ssXc5URc3ST6It4bKG43MOGM/hqDzd
OyM9vOhaoByNWecGBJkDXxtrWIQ0fd1s2uuweDF9vG6yroosHaYSqNDwtUDd3PhV
/lEnZOds4C+orlx+HvvOy44xFuyZJs50qIYfII321ngja3FzmAjsFVf1gkLIAVgh
GwZafk9asCPGFs+1h5gsIeGfr2W7DwywdRFCDsqKQPVjvxVxgsX7e4SZ5SIw1BjB
eGce2jdxUt0xIC4HPIir/EMowguKJu0KAUiMQrJwTxHeltxLahCWzp6CWEzDkLY9
Ti3u4dJh8ZdLeHrfI+1px9sIqWW78CuqkVKXpCtMMOAtMe6XTVFh34TW8OWI8BI6
2REtcs9UGvLHMEPq/U6N/2LKZDpzE1B4w6FCjy7U0S/1LxGEyEkDARyu8z2Rnci/
ICaC+spCkGW0JqU4f5wetJeHiGGT7yhIO08ncBuOyTcPebtCDHwLbGeLKVjk2+CH
/c/kjmh/lps1iGUFa0f5HqXRZZ2AxKc+9d1yFXBUYQNxlGJLK3XnFWKRlTh8J6OP
ID89fP7dRixnuaHykml6VcN7JlC0jJZTdmv4T3L37jZ0oH8c+4ypnW/NA9nhShVh
sYzzJtHaOLEO1tm5f2ilrZQVM3Hb/bj2gahZ6PzFji8nNj+Jx7fl02KiM4/SPTdv
03dxrkjyhIkiXQssu+ou9NnPPqrc/YuBpDhQF/hXfJEG+7yYuLL2sCKYzXItSAAr
+jMgvsTOLXtOXKfka6ix8xAIl3s66EcFt9Ptc0zOArc3HZwrfmcSkeWZtsAFTxHy
gtnAmwctCOrGP5ze3TJ/xLIk6n3JKz22HdoYmaa+YLp6h0a2GGCykhH6NDypQGX+
EBvEjEz/bKia62OAgte7Y9dgasjvH8was0IbDYbqpu0SBe0kjH/vy5NgQQ2/OVB1
kzp+re5pBHlHHZujwWZ8fRSc61Rj+D3sPQyPARuSBOQXsyPrVaH57ISlzLFGspcq
sQFqxT3oNGUwZNkyN/Hn1X0updG6fS6PpUVgKv7S8ieI0jmN8GAzx28P6lBhXmfT
8/xEFOR6nR/vr7otxNL73sQgJuCrHYjg15jp5gTVGjuRqugXhPJdSw6HyI3Wy+Gj
B7tQaIgGz2IYy04SRvnSmzUM1QJ1ui46gbpJrowp2MMsynTQOG7hdd0lxXRk5kFJ
`protect END_PROTECTED
