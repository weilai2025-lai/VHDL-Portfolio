`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwYuGOG2lr9JaVjg9zGtml6BcDpmd+ttzF5kJpV/Wp08NxYrjKU2FPKxtRMPQlM7
xyuV0MLtNFLx7EQTjZk4soLFKE/yW6VOUtBv4dRprcN/eo2rEsd2zL8Ry8+TuEjk
UfPc8GbirwvhT+n+z+5xJVqZ61PwZiZ8EfyxeleGpdlbMnTFvavHKO+BD9cnCp1m
zE1ziVJJ9L8VR862+dDxEJnfALLWvn/ZnFnz6+TmfqcXm218MNHXOWrHjnNbWVYl
/Ei3X12raIB03eMG9UErRx7t7jxfVlUVbBQuGVmfxdm6Z0e8NgvgZNXxPdPSrYfT
+ipfvAzAA7qjcYrdlkWSrfuMreftgl2Ekr2OOhQZGqeUVdkdA5b3hsV3zyHZdqNO
MhX+AxjQxfDrg8K2lV5yYk8oNSr6bnpVIlWUDo18ftQXbvpWKPX1knVArWdbWbBB
1g9/pbk9kNTcH3NJS4tIEyttodW8VcoFj4/puRnS8rv2x2q4eEqMAcUvS68TaT+K
r+jZhlWN7f6wY8CvtzCov9j/LbcLWrSFqbKrP6tPtSr1xYGE672erJyRg6VDtZ4V
nHntzY4pYnyan51hK62K3vQURY91FKoe5dziFa+PqJXx7HeFXvx9I6hRll7q7Qds
cSmU/k3giZVCT6hrYITpVRnr8kQTQZ0D6BJaJ1+ksso5gc9riq3LAHD72HkVSyel
yWpqAVQnlxJMchux5rMDI6fIwCzttgOQqsDsBZcMAGGwFqzB7Na5z/LlveJvzgI4
qDkC8jAQywDeyIwGDhFeay8z48CMjra7VY8cCv3Tmo+0orIgTTQKLGNfP6pNImoJ
0Ve84SlWdFrzztvGcMstLVxCD+nsih/+CCgoLFT+uKu08YM/v2TBxEDubaB8Kqwm
xVI9slheubFELj291H91i+XGxT6kG9oJ+z2dfO/EjNb2fIEVzuIBBVlqCl85Oxt3
uhleb/L3pn5+jsiQfdWKfOBHF4B2piWx6As6NQx6EMOAKp6oCBAW5Vl1s/saS9NB
2oA/mBhsbtOhuppjk5Rye07wp7iHROnVrvHQRtNvEAkRUHK/b6ehpTWNj+bEvXbB
HD4HG0azJyKOIC1GEcERpAgZVAhS5x71jii0H3pbUDjTfSoLRYDYE4MdBIDgy5G6
14cjt3QFMGFKRcUWfbC2r/FE6feI4HVsiAg+6B4u9TWMT3ELA/LCE6ab1rE/fBy7
6UdQ4g56IUvoOsZj3wQRN+iPYJEnPPJS1GPPzipKw3YrSWJQXT1Fj1R9abwEI2Mn
8e6/ez83/5wocoBEiO4eQJDFLNBrzkgP9Pe0clrl0yZkTypFZymX5ArsLEhiBi/L
HuyQOjzb0v+J+1Otjli6qWP29X8QUHEBHs+nd8x3PPD3JSSx/qhTwp1Ywz5ni7JI
QTX+8isZj0VR8tMF2+d4nGuaMunRbGTM1sZapVVRN/qk0l26OVtKGVi02G3Z8kLC
9qSFrIxgczV9OvJc20ksNKqJ3rqU/u/2h19z1i6aDYvzYhm/DVCOvOUuBP5gGJaW
IaAsSsCoMC/oF5lsej45g3A1ijZJx22N7g3cKLPcbVe9L3i63HUJqTx+VSz0b4rN
iYdG18Zw9qExQONNSQWZHWEZ6rZhFwLaVgKDU/7zU212ZjJuvq5+yLeAnJHckN/1
bd5h8F5Epni43KjUhZIFr89B8cniZsc5F8cCGTYMqmij4/UamFkYF/rO3tv+Zowh
ZqJ+QzNWYwnL2dFnjeO+fXNZfw7QvEKI60JxmDbN7rUj9DdYRdvC4LTofMv9ARD0
sIsFvvGzYjVVtj8MBxSty5JwgwKVxmz4CaBP+QtuPiM+9beYZN8FBn9Ko5b9qdVY
gl+yZVpYoKaSwtzxOGu83jLxN5Z/7xkNBBWcBPBg//omyLSbmIkqseKNkaC8N7zK
AEK4RzY1dd0hhb3pNa0eA55QuJL8RLA6vNfrNyxPhT/AHFy16D/IMs6o8hHh2coP
HtQTciuUjFXTjUiMLOOvN03jdbDmFIyUsc+HzohzySJd8B8u8zclIlQRxWtI+s3D
CF0kgNV/wTjJ+FePDiCmfPJeVHs4lWN8X77CpwzLSVzrvvLQtn9Sb71Op1wSbAFg
PpLTcBEvbZyOOIf241xlYsNY+5MPraTDv6aFv8gW6fiBQpi4+DvzT6DGFsi1oQ8c
Q6IMEVGN2HaMUF8VlfoG/KheLLPPom7+GrsBj6L9YqottJ9Bv4br1ZhAa66Ug2Hn
2KMgkqS1sD9bIIEHgEUPTIxvpjYjEpF76rGdMoK6EzTQT8wt8K2312eKRQxKXL+n
G0CMPwhvrgq202gugSBQyHiJ3UoHSVTBoIudsIpDUSxN6Ug4AHoU9McyMQxOGHKc
aZrOWfdFL2rEXArWBWj3iA==
`protect END_PROTECTED
