`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EG9RJ1ZsZbNqM/4AN1mU3IQVtPkLc/RhteBNzMyibt2xJPZMAfo/FUfbz8Z5z0Fe
LShNn6Qax5BNETg96CMYpqbrpLvxcGKvCaZ5TxJW68OQrDoQT68xZxYKBpquODNI
mf+NXlDCse/zowuwYIW5qa3i7ptgyCjqi4QsMgYfPzpiSsG3Bqzk7UKIXtNS4sWa
nL/8xdsJz58BwAfXc9FQvRbhGPaVrtlnAc2d+DgVB01PUC+XX2lteEZQlSP/vcZe
PGSGYR++cGBzGh2A1e9TdoQ2kXRveoYzJoKEbFEuGKhMU0gZ48yY6jfsCRyReKao
mBoQuzIPQ6k0vCMQBok5nccY4w0JTGOFTpR0YpWLOf27jn2pXuhzIjwN4ktdbjyp
QPZceRWGSJsRArSqYm+8wK1fo3w1YsMVOriepeVBCbNFRBLCYaaxdS0/RP9AMiC0
`protect END_PROTECTED
