`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+5tOFteyluWgm4kZvzbFMosHus07NyFbEyGW5bVbCo0n9zU6CNf33bGZEp/pol1
ms22OgZiYDJm1AD30L8BG1DO6Yw0o1cpcejub/7PEnLYCOmJQwXnviTCVLXoNPov
rz6WvqKLCmVCD9SHYR5dCkWqGRyaoVV1M8p/Qm3pdS1Vr7uvI1b1+I288mq3g3XA
BYF1lMXetIm0qcYyLNzedaZ9c4+/ogX510jF6SHGa0SBEyJsl5KDAz5gxoSnaZx0
INtbiv+yKpgenKgTEaVad9eQ1PPZPOaHsgLKrg5n+axIHTFLotHNLdjGcW3yICTi
JQ1b1c/sSvVAqwJjNMTw3r1bORUJNU78a+CtdenfZq33KA6fQkIZXTiK6y3XBivJ
x52gwT43+DxxJtaXvIWWWJwO18RZThapBbK8LNhqlF6n6BbAx0132GTlhGkeB0xF
z2HUTET4yFN5X7KAF4daelkk8FA7EOqJgmtYdkwp0VXrgojlLZ/qdwUH1nb9BE2o
beUSdYgvd7L4AYD639dMsmbeD58syNg2U9/PgKSy8mO/VGs7twuxI2etQQ7lZ6uE
CjDdir9e8PzP2xgiWinoAJOTuPDy/aeUNetvv1/GXqoGyZruduUDcChpViSkvwhe
ErcX6GYzs0WLWpRd21+EfuC9wbTiSaZS7WN77ZvM3BWb4EwhuS3ZCEL5HeDlu8hH
HkHZRcs86FLgLmi46kOavgT71o2NVA90vtRCgm1HAAIMDEP242SZtP1w4CYjEmS0
krj6VuT/jKByVLm8jig15gTWrPmqjEjBh8ms3+ia+FJafMn86nCkq4PEyo0m4sKi
8iZgX1KyqeMHpk1WNlcvZ8mL0SS7PRcTe3h+5c/m7+uRRNorANMrjvwSR1Z1Dkh8
kRxIL5xEVdBuUFKRbu5jzah6njhZ59D3RfEVVx6ERchYamq7RDDIkOckWc6Wql9F
Rq0BizRdGDh4aIBBFuxdkjgZPG1rHWT/DLCQlbejYhzL02PwvioY118h58CV9R15
jPEyPUZJc3flFNxGBHjAwZdfgkkcxXbfAM77cc6GPQ4uv+wR9ZDsusszVBwWQ746
o8fn9rZrJ+BrW7b1eJmWMYpdYzOtKVezXbZxzNpNTzbb5lmjC55CqtEmBiVNldGI
IkrB/eo8pPyalfsB0hljjOjvg0HRmM/VT28i3lBsF47g2g/u96Xq1gbKc9HRXYAz
etRpfOVl8/0FJOVvSirqJPgi2tiDGCOlQI4sQ1AFc4fQPmbl6rb6r5X7m0q3nPPP
OI1xRtaOPgt7cij3nU5ldfeZVedRUorCb76od5NitrkzkR5K8Y/+DDkNsvpvzAVc
m0unc1jnddrSqYKCD97VoXFwY40kA2hXr5nKIslgH/KjzEADtbQj9rsaQe2f3z+C
paR2RjeQ5XitqvoWAUHG6DhQmsAHfoaVZJ9OsXR5CR/zTFYV/LoqaTNJMuAhulDl
uaWrGX8fgt+Vtqmn96DXBJ/nwHaR1LgknLQvR1A3jHimpbPP/tJabYmqRE1HAr3m
DNVZz2wRE6T22F84URJgP0eqT6tXDR9KbRX50Jvl3UKQBRH2Zf5QAMcM9qVVI7w7
AzW7BCj6psuw1KNIdqKZVrC1oXr7VhC+PdgHgTFqaIf+SZWX2avHMSb9xUAsi/bd
zl2Vl56xnaAHDXY5cDDmDhfvbelbgtUucx8sBAJfyZQm5mVNx93jN0/gLgx0vL6x
anv9n/Z+3zrc+xSWayrQ7TAeEOg6M+RrB7anckqeyi1jzIcpF0aS8I8Ib5scVzO1
pGS6mIdn2yu6fE1x06tYUowvKV4Dt7se1pnq+tXqZ9Nz5Qysp2tWvrbBPropS/TI
S7jxCgyGHif9ODbRiog+acRosWxfNQFb+zc2++Azrmx1cHID0DjEyzuH8LBn4zuC
u3k1ezPaas8jR/oMn1psuFUIF56YLGIldGa+rgADEQRcUV1OiXdfP2EkKL1lmWti
j6h+1xB1TGUG+Di6VU84L6wOF5+cw2Sb9rBtuuJ5CFdMSZyAKqvhlkXT33/huqNQ
O+gPissNzsquq2Tekih5GcAisZplqt1J918D/2beNGv6ii4jyrp5zV0Vkx7tupof
J0CGzo81LETkEFV0+gQ/Wt7UoagDIuZizTFRJnOc1d16c4Un0bNGgEdavZSTqtxc
u95YGivD/1qTvWiPFdQ/1KE8bf2dPy/7fW+yW0cuUmhQ1MNoK12ttrtIUjS+RSBa
V2k2L4LQyu1phlVO9Jof6dW+FRo/1lsf+OGJfi3gFDYN87X4QclVQ3X5XQlHGrnr
C606waKgrRYEAj1UcWy6HW9AXiqwCcgx06Uzto3XljXBDpqizD74bysLJElY+uwN
lRqZOncUvYXKvk5Vodki6tk8HC6XaLeXMbNqjm/4uyBUa2mmFRj5e7RbglPv/4Ng
P+Wpd/uFmqO2gl9F9DH26+1vWjeVUouHa+yka9o+k17Vqexmg9npM/ofI8NC709U
bTBnTjm8ITe2ntnOsU0Afezd9mTJ73wRNEagFWGXQm0UrVn4tJ5KlXP6owUNbVuV
5XJnozK5uttx+svPkHTMsPTyfFCKqNC8+A9RBdtSMSgouL3VUsbPEklR0bvjSbH1
prf/iHDc4AyR13KqzpoSFOJnlrr2VgaFywyZgAvu9x+E7JkIOQXY+RcO6n8XTfNL
YWouDcE5vOO1VlFxFVnpRqQMvUTAf+KWn5KPKYxV4zetS5TULZvnstS5bm/7VAMR
Ttpyne8k31ZJV/rUEAN1JRY00m/hmP2Jbw+4irBnQPEzdztm2TsRhAuqxZPUwp4f
9aevxqaFU6qydjP5lmwaIgBHlyY6w7EGKx2sWSin5UAHSdPj36Dm7cU27r3N9Gq6
K9vr0kfLSytIq3k/lJLPAWIt2M0Sf9UfcG9w+8uQ/jLSDtEHCcGYAr45Ewt+7KME
aUBkryr9FEFsw39VXdgc1HSXUPa/HckB7UwspMCwq005iSR1lkkejSRwnxV/sguy
O6bmOcJXk27oZyNCHZiz0WJlYRdpj1geI/UWMAzCaj3mjsqvNzTGkFie5YTrcxVy
3YJ0/IrEpZnC9fdXMVRbiBQYXjYIcGNLv5hahDPwsTP+QUIMpxYOx4MzEi16X96S
8VMDunph+s7PfiqDKahfX58FWu74QtvihHLU2+XeEHm75UGRwvwtkbd9Nno6jSBK
3V4EqrNSHUSQpP9V4M/7dNVFV6KslpqYSeSpEa+5vMoTC7zW5SyOFwLlw9bOYoOp
qOBaecotBoWCy2jfeN19KYvTQT7fQd4gPig6ri5hybWFjiz4qmy2aJ+8eOkwjXeM
VttXB+JPXuZbsFLequMxXayCLtZ/7S3fGy8IFHlS1oqTJjSOwkISBkmz1+q8bm7n
uYptS0N7n2xCXga4V5j03nay1fKBcuHf1oxYpN54EbosStTQr+6XZ9w38NKp3a7h
srRl4lZUZWl2V8efMynIGzvWV0CEBOeHDJ/CTbu7+MRO2sZr/I7792gP84BlXW7O
+34q3MoGjkoSJcBKtFidmGsNAU8AYDK3yeDvMpPE4fpGR0cYF/n7RGaTyHRuELmx
WoXI6rRMfaJ7lGL6Ng2QFrIyTKpARK4JXg91B4YJTUWr1R+kHxcj2T3pNxPp/Nni
1RN/WUeY/DD/PGnfas4t2tH/H+uosnBcOcc/I/huSgvLmWJLBek9qkJ8nPGgoSuE
qgv48koZiW2KO2ECn4bBz8LgvXctHEOYaDkpM0igDyChH3J/0j0O8+p1OwhJvTua
sJo/vQlVd4ysKnw/8XkpsiSoAD52qVwGkuw2+u+m6KDfA9H8KuIjvLhs+lq0JqwQ
VrCiGIHOfA8O0baL1GSBb9VT27NDCtA8NWfoxdjVjcqUvGtIi9Y6fvs0/9hhGXq7
+cToL3TsWT/ZSSQYapKR96sptf7xs1RpOTa8ABBC52Vn5a1lLVsZBCSBSWXY/pfT
F0+oVct+MUGMLQVmQ/j7v+xZ1cztwzi7cxv3BLV1mfGIAyFaGK0iQ2rVJh4EqQf+
ilxbYPWDpuh6YjUYUtkWXuP5lF0myYgEAmux6rWMNTdeZJynvfvw/NSI1ijJlFGv
6DsGULmBsGmypGtw6+RQynGaFNe7DPO+neRLtHfuK1yZV1xCDcsmL2udCV31ZO8p
VHnyT6isXMrcpV3USoZGlxy7uIteSZ0ZvplH8eqe2DwAK193xY0ZMBPi0RF9rr8P
Lo3EwnhEEtQFM4UK+KewrW8RLE5PAmowITAyTDylW+7/uFm42ADapjYejXvbfmgl
iZQ42M7hgSSFaYiLM2GH13M6ngovV89oYSb5sB2GpyG9GilIZMZzTiGDZ6jeyxz9
6uT9Mo/uyAm7UC3huQ2vsv+j5JmaGeoZVPkdVqqt6oFsaY8fc9YGVcrMEdjBH462
ptzL/j6lB4LfL5W/8HLzP8vLCm7H+4HMYuyNPCjNsruZRoe3gDBG8DLXVErnOBfV
QZU92rKKIP8IlongGABZcEG3lmnZ3lOAsZIR9AWIIqG6/CNOj3HLq5pI87I/0FRH
sa75ZbA32sVEjpAPxiR9F0Az304vhdfTYTviTkSnFTGeMTtVT6E70+86LPZVl2jN
462blzO5CXue0s7Ap2o3Lv5n4eauxYX/usUpCMuayU/ONg5Pt0pAooZkalwsMjur
BCHNFzyvrDOMKRpOI1tGoQeVxIDnUvW74XTBvY5xJTVz8/yoa69mKomL1Maf/p5f
xicfRxCKYmrFWWUA9PXvxyVmyOQ8iH6U9WFelxb4xdAD5sd5oLnr9DPYyqU1c9ML
j0ZFpjSI9664rOsCjqOjFVxfuSv58dLKFAyE0tSEscgmBBZoqjXNUHfxk0z8l7Jq
FVf8gkIE5TbTyM+jexCQhG2L85S2zaapayLHmZrU5y3XR4JAsv5FB4EaZEnX2n8H
u4NRMG/dHoFuuyKCbhQpGWqfVXSHkey00/D8OJSG+K2uyYh2N4Ev69MIE4Ebc0wv
7MnY5rr908FtDZEQlcCsnZVDTcNsikr26yyJ/eB7IrYSYpdpg4QzDq04qTIdmMJ3
9eo3JZ1ypEazQq4UqZOn1yQqDHBR4uLENKJlXW4NN+GMtUG17wIZiHAIy8Q/T2dL
eTVXUSxVqeoARvL5s1mIj+eGQy6RYNWpABpraRGwVbFkiyRCIIUplOyKqypR24bf
FRTGdhu/GqSHyssPFcaiDEjdoVqwHhZnLqD07oKHxFIWnwIkInqPL01fwuSAMQt7
cpTfqnaxJ8Ou4FwCXpEN9jaLNTwlImpRJIKzCF3KKVYm4wQnMgUmPIdGRPRR7FlP
1cPF4q4zqTIfrUrI7N6vEKVnP8iMAv9Xxkg+ldIAHAY5oTuogbQbv7SG6/KeIBps
4itewgtHoGk9XT7iPcBwRKzw3+Oz4S2dfps3xenWnN690nM1vhxDuFgwwl6dV4Cw
j+HvjyuxHDpR1b7JBNR0DcBxXKEQHFWEMIYkgPQ8FgieSWpf07MjOR2FtwxszRAo
/GXaJMeE2IbJMDnxQu/RTNnCaRaKW5EhRKcB2iVkeAYGeoqtbpzU+8ah4MxhITUV
/EgiQa5UXG8qgvl7rw0oOkjnMdVjPwR1edNUwKgjdLGOmz/zlZLlZNIG9Mfw8QZp
Gc3ctNDp+LXvzXh/u97eDcBaC+zUFy5UJqAoe4PSAGfXUQltX7xkr+PszGblO4XX
w+5FU7QwnGQTirRYS87PmWUeaaGv5yllFkkVXMw+sBvEn7voi2u4MZBC7PcBh58D
ICnh58YXvdA9yUdc6gVTJuz5pCk6SGghV6c3DgFuwArFRr0FF68IVG2b79HmWth/
3iWJUKU5t69+0WTMSACR0sqtOi4+xzD/bfcKbrLjv4VsFr3dbrOYPsUea27xTfv2
OlUsmHmuY8OpkgZJybzmi1jTRlST/S/Ll1j52w0GLmZ38ezI6QWkAyoAfkE30e1Q
oE2HgotmIF3bJyK7q/6jJuxBTHMd0QvBE8uZYwLFBqyv3ykC7WE+7Wvp+odIXGID
hprQXREIJKgLKnI1MP77FxJGf30QYiZiKNobF9XNXm1FHdaFOs72AbXDgADGBQfs
bwycj1YwOXkNqaF4FFmFupP/sXt+sDlKxyOWia9IcLzvdMFdvZ9/WfPZeHQb1BXp
MBfnk/p/6FjJzckZsDu9s9efbqbgOjy6+PZ4iOS+KdxylIOUSVctIDTwnbDaG+mA
BK6zkbJLtorWYtdCcs8KOFdJNOnsZFjexcoVpVggguWhFuf5VYmX1SS8SMaEjRdR
X2uNRtl4ZO+qnH3saYMPj7XN3rGmG/ROIeUedJdumDH/kUDOhTcpXXAxUurjKESr
CUmfgNmuKfFelFiEKYV1tcMFTzx5YvqULtynQ/9nXNza7vR2GS0dQTCVdogAELkn
XNU5LywEADbIrUt6jnvjTZA75ZSrQXLOeYF1JWpnpxiXMEEITPxMLiKwjhjr+ny6
2KwJyI4U9Q2EJ0X9oC4A5FqTziN+BK6M9HoqWt9hk6Xwq9q8a9eDk/JH04rA3zqa
FejwTZrM7pK2CxD0ljSuLtaPbS6kGm4yso7hQl5aylNaJTQjNImgNFrZZyqcFzv3
vx8EtDkVQSKoA1FL8bkzZG4jCRI2RihXlSamkHFQNainuhdWCMQAL4FI5Y2R+cw7
++QJIHAOppKubmHod0rzDINCrt2OLqq+Dm5Eg+jkCA6Vu5wky2ornwhfzLVIYEjz
fcv25kwYwoJkNnmp54o4L+lwwfuQTkNaV5q7S5N+HvRYrGOlyLJ/Lj+nfVy1S2e0
88v2WcRsEyGO6dThNXdai/6cSQ4t6Q0Hjp+3SGgp69xF2CKaUx2OoCRCE17wzwk6
kSazLWrA35t60rUWe70sHg2Y2Rf7bxrETzQTF+FGuV4lb1oGzLnnkyJoqMNiejpm
zRrdlv+Aqy9w8/ekuXmIvok+YE2GsW2AABI5ZN7p9URaDNF0ZOz+G/oET6OO8KSn
oRqbKYPjcN3Wwlr5oYultWfjNKMRSHL0rjg/vEBkHVBSZYFAGTdsDLyMkzN1sr0x
rduUfh1epq6XyhRwXVtdoOrUvg8rm+5C7dfly/ToiZnwC7D95Vy2UUrTi7wPQKqw
YT5bxhgCTJZhwxwVwg/9sKRPIhtpL4yKVRs2+QxMeuuA31v//H0H5iss5lB7FckJ
C2/kjUnmSyYyoYyF1JgSLVuZ7LzecIS5mk9LE02VZzpzvIQ1eEzc48BfgKuXDIP3
z8x0nTstMvFzCccKmR4OQgRh+F/G7hRhiPu9mwr7bm9sirAa/D5Srr8swCAa/kG0
F0DFNxLA265YFHuCtiBqGGd/X++2zrfC0d/M13nSAoVnX9kK1eJjBlC/vFOrwq8N
HzPC3KbIGaZd8fXXGINXucdGoAoxsb77Fj1TKPywohUF4gwn1cKa2P8zJOFMr58E
rGzJib1e/P/dnTJgOYQ32IbRf2K2RvAES7xiqdBIGQi0uF/M6xjFJcXyjjsJk8Vj
PxGdBAjTxFoE+tSM3LqdmtM6MbbLYF4UbFEc+ezV++3QcpXtkvUDdgIYnKLvRPAa
Fymr+sWIPTVkBRTAm9SZsFcAgiOsZ2lmtdvMUVmYdgZ4X2XOYPbZcXiPfXExcqxg
iUxdOWgFi7OHrlyxWZZbIgNIOW1B3hLpBGC4ISLIsxuyRk58EsLeWtNabEBHfIWU
ExKkhpKgfn4zRnks5X6edoCXIgQ41W7KIskRHHuViSZA403bq95fujX00s2e4wE7
O67tkN8LJE7MOIogCLr8u4o82e4Tlb6WtA0oBtM3EM7vgKAVjcar92YYR2i5rK0v
Pnnemd+lukER+FIPBLjMrzI4bIboS/0mZdzLUk6LJfrHAh3VIpfT3aBxw7pN3dOQ
QtPaBRMWzbD0cQWfvpEx9Q8PpQjjYDnEslbHm/YG+z1HtZnVpwWW1NPRFxw+4B1i
rgLznhvhCvLPfznGAYZRZdDvAFeSoXLDRZP6+GjwZxyAlp3+pP5GYl9BsRP/0i/F
NC5FTxkyVzlB5Zbzpj/wa0riMmNyD57Fs709ziUVkVBBqKtRB6qnvWfL9f/Rxgzg
c18WcmyYXDU/qJSevIQFUG5NeG+Ww6Fvlq9mGbfIiuZTlkUGnL9JxGKbCe8+6T8w
gMV3HIBfJ8gCbZATDSsQFGQ1ZrLjE9qsOrnOxzzthesTHH+ae9y8mOQv9B6febMz
vaPKuen9tNXJAOSo5qtSVVo5cleT5rPqKA9mcUduC1gZoaSWStrFnLBGrM7nL6HG
Txf3tJhGKJHpyk4pjxEhF9shUVB5cmPOlPmQqeHhwR5UZfkJNG+oA7/mYmejtwow
qISN5JiBOn5LN/usiU87k5jJgkN8cjepO1Go0athbBTI1g8zaSVqkDRJsLqzun3Z
ZicgW3ApWzKh7JB2NSQf+XIczWwksRrk6GONMagIfCzUYbs4aIfPqHEK5//rZkcB
imAVK+QUt093Lo+m2jcd9UOX8HqAuCYiCM2CUTehlWRsQLsrG7rnSXxQVLcaqDy5
1+85ltfYbGzJL/GcxrjSL5RqPsBGIoXk0muVl2DVXgjQYf2tK6C30hW3RBXhkHtB
BPYN/XrndF/FXfLlzYIkbMHTgYdXh9SmqJ54JfT0RQXfwqbjBlj085HW5Jm4zk7n
+EFNYWXCqMT6KwJZLGmCCzi6O6E5E9kAamg71LZ/apiRy3mLDHUxOBSH26FNxSHp
Ldj45bmPRSUnAGpUf0zDEmzuu6NEt1fzaoyMY0YNJw0L1ie9EYaGrkhteeiv9J70
8DVt5W6hEaaIBae7if0+urvX0Rjd8IE3w1lKvDaHniMc3drbf/nd9k/cryhab7oW
hIXO1sw2nQcJh8kn4HJEPqVB7tZ6YCBTgSLJFp9NspH/TydU5eLFqm7j+DPRSlmc
GxSiWsggBmHMVsSfZ12+56WOGXxbledGe7XhfjNPhYN8TEjTWBCc6ENw8rP4u6qX
E9bUvZz1ioVF2xmotZU1SBm3MdJ71zOza9AYNEfKw2PLjBzfBvMVEH8e4w5wCih/
qsagBi2DX684Zxg4zMCOzVpg6gLR3bS85h2Fe/l8zJgVQeZJCNe+QbU2PqirOGRB
RAKgFoKUd+Sgo+rU4nGmIZzNlZdYzVGixnnEDwvjmJHyqweXNh3hH+hW3uVRI3rp
Vjp4fa+nHP9dk8CiA3V3t5pVH1OXUejn8cTtctsOnt0BfV8iKxE5QOVRpQyTgvfI
aBfM8cllnBV3nyWe25CHzMVZtRyTVBNTMzPqDrK2TUNyt+rL9i4RFDo9DRTnvYdF
DxiAvlOekp0dEg+IWsFYvsgRv+OjN6E3Z6824in8ktuUwevTjjVcSjiUAJi3wuEL
FDZQLDxTf/8tVpqjEesehoGajsIggKHOaql5fVvT8D03LUMchl/Y/x15rb6YXFtk
dpmA2Js/73CjYPK7hzi8D6Tq8tbMfGsGGSQJk1bElnNt74/G6Auto0KhHQJUeA7c
mXLlMdQoB2XUm5KelLoQrC9HWNNS/WT6rCsriVlHScsp7g+HEucregQTZzj4r596
3omueuh35RUbY4nwoFQ4cSOOAED1UJ6TEyxRGUO457NaGfV9xbqEVgqg9tCynpjK
pfoOyyYSe6+rWEjVZxDMlCdl9k8CwSxP+t5VIR9FT+OaCR/dYi/oE7ZvJl6kUYJ1
vOTLHyALaRbfiOK0JRaFCULHWLAIwHU6RsBHSzu2UJ9cuyyv4xCGGrr3Zxp+YtRt
0qN8OeTflGB50fRIlhrI28saX6+iN0px6MgwPCEt4pgzoRS0wibGc0MkJZkWQ+Du
yo8FPDkIaAz+HTtXpvBqGhfKG6wCFVRgEvEzCg829m0uxw0mBj8Qv65lnTnI99KN
HYb3VtOtsgHo/JCCjCXVdmtCHohE9kt8ybt4ML8zQ+xs18TUI50+FS/MsVh5vJip
GgGtXio/Iqzx6NzlmqA8dALqinbFDajcwIrjfDCtSTPGBckkEO+l6BmRLqpc1wJx
Hyp0rFii1txZE+feM1QXqS+SnguquXEdK5fqbG3pbnUOq4Kc4M5FOysB11hsZdg4
K6ZEWl2G4G0C0TnwGQm3UfqLgZmBleG9A9jPN55BUCS8Z7+qV+smnxmDioxhRl44
0UCQBfhp/1fneHUYZoh17IV+84Vt24Mf4KMuQJAMTWDPraWcUeoleW7l1eCKoiUr
rwiPFeNwwkXJ4NkufT0ZEOuD15XCR0utwGShL4mfIGQUPk/pA4n1xzx4qjDefM3V
GRtssb/D88Z4Bbv1BVLdZzwud8EajM7vnFcF4hnrlxLawQ8JH0s/W8VCPd1Jo9+0
crIhpW6s1zYvLOt5DOeqOXFXRnNotZ+MubS2od2UQ4wZ4Kdh+3AKlINLMNEkI9MU
HHeERvT0q5osEqXFNfyfShwnym88Va1Y1VJyEa7sTK+b0cobwW8SVGNsYkUb6Dud
+SaJW0N/fJ6dDMKTBQlsLTgr8CES2cBB8O8qLqnIjV9tbKJxhoKcOigA3ANtygTC
F7/FN0xdhAcAsALzjlS1Xo9Eng1MVm+ZhHw572lnvJnSDAB+lP55dQBEXPBOXwO/
OBuM2osYazX4CE1QPhAZ5vI+0vYTThcNHYA4IYz+Ws3ApmH+O8NxZo/mQ3MD/R9c
MFhmirr6ZykwegsT0tkGep0I1es7R/CQl6vj1TmdpawJa1O0fsGtU+CFN6S3S0Ay
kAf57AyA/kseZFJgirbR5UOx4KBD8VrY0ZbKpDc/Q7sA1R8Rrza1Ogg5+iFCaD+J
SZKg4d4IxbMy3zuSCvCcibnnFAcIGrj32a/GGOASprSU4P2a9s/Ch8F/4dcgu/ri
bb40pQiNyuLw5/tqQS1Zz932xGCoY5RuIEcUZXKXBsVGTNQ1SnCkhFrRo1Sa7pva
IPCoU/6SCOtKsrcAbZuBpNY039wACtEbBVvQKJm7C+c=
`protect END_PROTECTED
