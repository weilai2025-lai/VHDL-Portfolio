`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lpsFSOtuyOQsfgHOBk+NH4U2C3LtES0lt2OsuLW9qrNrM3j6bR75698mSeRKjOow
QOwQ8LC8ZVKVRMNvFBgMjbbYKOgTV8BSp/pmo2nCBrjE7bPn+yPe0qFWRViANpZO
xBA/8RgwhdPSF8ezBLZfzkvaonSrOYWDlueMq4EfbPwFWN9Z2mPJsI2nHocXVLsH
xIjC4MOZ137mWkQbdH5AdA==
`protect END_PROTECTED
