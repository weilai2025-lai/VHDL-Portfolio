`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bz+ER1rcHQplcQeus/dMsl0EE+H3Erd3eHvagh1DzVDJvBG4VVZMynZO9bAp44bL
wSj2vw3W2gxPqMxmcHvRAsh5/qAwOINinrSoOVZF4C1Ux6ufDq9NKq17sRMLkTtf
j2+NgxRHqi+0y6hFkMdJCkE+WY4hQ7d5yPrG7pGZJ5iwdgZxTwVl526tupcAfiwb
Z+TNsDl5nqdxhXg1FCSEm6pkn7F/+LfwvcubBHydSzUH4r/3GS/Lp1E5Z1NOjNzE
vXo8e2dlQU5nbHJiOsBVYbJRQYyrjI+8f4s0i77GBHKqryHYny/dArfYUOK7dOwu
YSyHGpBO1UBPz4VArb32pwz/V+1n3vKBTE0abDxs/GFFuXnvA9CpOO9vG1D8vd/A
YwS93FuAQbGiTaKJp7WEvzVdFxUE5FnYaw4CWNOgyHteGVyHM1bE1C9JBxivCDuo
981f49m+MzLQtLB9qdDeiUn5xhilgCNaf3CPF+6xoFsyEJfqOMT5NVSFlGuocuL/
vvdq+QSrO3F/eo9t1w2fJuIf4FqkoSXeQ2eLnxN60R/gnFMuMwTkgxdFC107cGvK
3FMkrZJvs5IjBiBGA1NOWaCwYf+fzvV4+/Vu2FySrQopKpJBWpxxpPrYacXhhgPY
Oel2ePFew/wIAcWcDsDhVcxEtXR7goE2eFwhqLN5DoLWY4P1ViJ5NFZgvHX+M9U7
AfcmeLevZm7OubLOcivMJxxfdo0NqngHv3KW2jRe3aaAioFbCLbMpAvhFh3WPElg
Od6rKyoqEEikamcYGpjdKLpKLTsHhY4noEZaX6tTYzrVgP1NFNb14mU3yD2gpt/9
f6WU47ycHK+FA+lboJYWip1DQPcHGADiw0n1exBdbc01EWxgpNQUFFIeiaDUhO3+
pw0wqckP7b2OKn1PCTP9ARGHr8ImxNnHNOomsIE467vqKviJu+S/ojMXq/7FxG1j
ZsKMsJZzNqTfWvbBOfDCvzBvxrtRnVnphXbtuJmSCnROoK3HMEy4qv/up92wlMbR
S40mczX537mYmOoHS/79YJduDKdvogbLUD8TlsLIYn8/v7593H1EA3qSdQpQFH8j
Cqzep5ABuDjvO9wq1lBKCqbc/QPagfZq+Q0aMdDDOlwFWYnvSLGJkUXfYpslFUyU
r/kzcSpr+FWFkLXBiWbY1vfszdXOi4DncTLxE/oZPf60HcwvN5ze3hhU0tWhZQLE
VHWXn/cyQzCdjuSwQsNnok49Rd0X5XT5W/epTsXJlgXsfUFq0AFyW96LeqDEBd/t
rVl6ayO12gGPHKkRiTjEwrpYxyTqrDUu2oFW84B5EzB78uvq2FyU0WwH9KaKi011
/F6InLF+6tRrQQdKDSudArsQ0Uo9G8C4lyP3QAitFTKSNxt6Sn4bgXvfSMEcNL/B
lOKmNZCyg6f4aZqUmhRqV1El07WjxoF2oJYqKMVNyIPz/Gtv465ZP+NGAZuU3jRg
UXf1/+jp4h8HVhRTScwqvfx6F4GVpGrl/HqmO1cTa33Ew6Pl6dwkZUMnLZedCc7v
qtlwAJk7r/aaMtiFiWcih4W//OtKhj8wQBTJVbJgBCxqWc31tj+Lqv4UwRQuipmf
mW1tTVzH9rVA88unHWMxdWf9cfJqZARMgXapwm5G37SLEebW5QR0DrNAbTBRy2mi
vCDHx9enAywHIIZK9D39c/CcI7kxs/N8lWDvRUhxUhd7dvaIMkgHXLmFiV4IDHGI
/+ARrq1fZvj9rAb/GeOWxmiY8hhZSNOnB4c4oJhVmdQ2cdViKYMkQJ/DPBNNdsKu
PEYEUxm982Xd4v19XXBRNGTWKmLQWhDHiwb9W/yynLr1CQS0ZVt9egoffJFErkqp
OhHjVgZ7WjToUFqXvZhPW3UHOFSfDaxI+t9iwvkDBQGfPwBxKKC3ks+W1Nsyko1z
IWw5YvjTd4KzSYqOAYbYP5bMEBXpQA+vVuQbRoPE/9rgCkVwpZoGKOQFB3mZ6eCo
ZiTGYp+rY2NOasnuBl8FTmlf53d7Wy8mzUH1kXkCNHIFwj7r4j1WuAn4tWmuoeoy
fqytE17d33k8kCPAgOMixhmK+eJLa3qRsBA66b6kMYfDeXp0buh+QynEG6JioWi1
3yRsctV1I7OSJdyV3G1Ek7zHu0aipMPNIZr703SU4lhXo16bFEtAfuYlGgP9RswW
jHBIZxhEA/3H1s5FE+5PXlSLFaujRFPDX1IzLm8f8NBPqYHTnUQsuw8e94QcFmWt
AY4cCnx20AalSOYE0HXTe8IeARPEuZwz/OrtvxEUK2ROKaXpW4HtZAiMFiVPcEkU
blIRKNXvHovmYrzNvrB23iSAM7ej93l7bg90N1XfzwmNkuTBR8R2vAbNra3Etpls
CysL7/kCr1gjFn37mFGAv3rZk3+esY2x+QPurnYhpQnHcKNp5ktJcNGOw3bZcsxZ
93AA7+RhT8Py9OS0eMuJTYM1hkAA4MKuHxCD4pTEjf7wxCsQiU9Q9RnjCMtYeihV
B5ZeximgVf8ApqNZNShFYAB+Q+aOHVVcdsFW7ZY8PqTQIy6uCW9vV5I6bj3KYrKU
vAAUlLJBAZMY1h0tXeNUqBMbqjWRKqmZE4eSG48ez4XJspfsLfMbaM514NC3JLu6
kwMf30lbyL6Q0+vL5NmE8YKXW9woCCEbY26vTn44feTLz6VkaAcSdBl8EIaDYI25
EZRz2abKz8Sw7jH6Pd5+NvWDPgxOwjiiZx7Ovl+5b7tPkCH6tDMoGrNjTXyGb4Bc
xzzXvRylcH0zl6T3FLTBFrSXwTAV61RwBY9FtWCoLJxHfoDLZnZeLN2n5N3qGelR
oECRKQGOaCGTZxBSTklVe2ZE7rR+0M/AzuEtdyqDnQCo7gTnANCD3kab0okCXUmH
i2J0joFQhIwcE6F55H4VGBOE9Px62pZoqoS0IHQgGmPAtX3PelRrR5SVnko8eKVU
oRbO7hoj7Ctm8wQI7NB5c8nQtcJKuHkH69QO0k4OMcaXeTESvigEOL6dWVd72i1i
a8ATkUdXKYxI1a9A0SFBJOly/SQA+VC1Mu7Fdg3ego4p1KiXryMiJDQgNKUnAN7L
pYeDsEyC4Jc45NQkwpVVNVtjxHNL1Piid8u1mMQMRi13FeG9e0Or/i6T1R38/qYo
3tCfxQg6hyE7CMYZYDyTpYhMqg9kbGmRANBAe2i114RzDLaFvNkesqW+kSLpw23U
LCLAo/3Swe6ayAYDqxkXbmCgKBOuqdyRVlpRlL9W6CiXFPxk48XUwzEDLS+p9zr0
rhBkPviymzL7M0uGNkodAzffOs02QmuYWKVFw5ow+sRrea+MGIEZhaveoomEudu2
sJFp8AYp5jsYN2H1D5i1oS9WltO6afrlEWbEvm4NiaPSJ8jRCFcajVwt6UATqZdm
BuYUu2v+kyrJ0NCdaJI9CrCqgdM399cl/Lr7lbOJIUM4wXWJBH6Zk9KYX4PGLD2w
IbIeWavOM+pudgKQNb9E3rwd53AZKiu4efphI5R57qb8LRUvHe88sVGgHcakMbAa
j1yoNPiFQilJNTix3DyurTSIo1rbaRLIRhxnb9zqD8kQUj90q88FDL5oNBuGaXIU
AnE6yvWRWQYOpYBd07zWEiDcxaOrOltkr9WMTAdaY/eV822AkDy4W1zTAm6lARvs
MbMZ+dkDRu1Q4E+/mOhERaG6OLntdsR4OxMysc73jsUdK9EOs/E/ZxEp2D0c/Aso
9w23CGz8ULvJ/8DeI0SyycWhlzqZSogxG7QN1GScPSFohE/3LVy1mXQiw/DGAwWC
GRZ/jp25RFD2JyK40V6WIfyeqjx92PbbggIEG4OQv9/SgxSrxOw8mY7+i9MNHl5l
6RzZAdnwFxye61IWV+nlAaJxg9V8oPuj1b5fgLkg6veOl+9eG8LA3CrszJYWRhs8
ans4ich9jQgvkIl42gJSceWxAHENzz+6MJ1hTXgcLXc76S3HuyLRPBizm90d/Mfp
zXcdwCTosSG63AwVo5fFmMVqUC9sTKkTjhKZcAHSlu4YQ3YFVg/lmXwehjjN3Rd0
XTHKVXxGcGr5MpRFRu7UUkAiXiGAjTRjnvJJhfvbAU7PbOq94dX0Gb1hEsQBGWLT
koIIE0oqu6kezgoJa61vToAVCQaCQ8lHPz6lbUAe/ZKxpkNGu8k08iA+HlDX7EB3
NhKxGx1OV/fFSuapmErJQMIyCGNJZzuAkUM0Wn3VPdWgxG0g0Z6p5xiBnELeKbx4
xYXX7Q1ipA6WLQoW53QYcDFOmK2/LMrtZ05LN43b/XY2xlr/53N8hg4iAfUxDWBS
a2MaD+fG9rLSfdgZ7Do4hRo29xhaUyw0UFUJMy2yxIfZsXU9t3ej2/mw/riUNTEr
k4vTf+sY8yNdkIt+pdOnbNhPsddvkw6Tyw03GIPLX6Y342OgFT6CdmB01hqzYs8/
BcHcRlglANwZSItmm+9WhAliCiDzVgRGZ9M723SdB87ejBMn2gCGUwtL8GIVUs+q
mfgxc9sGez8oKlmQcxJ/Rk+ticHHStmYMAnV+MUO8ukwtF/SitM+FM4uUTYaxLgW
ap6BGmaFT4IvAcvmshTnqN6Q2yfrmUHcZNNw2RFAO6bK5oD2V1rnbT2cKPLzfz2m
CEuv96sgHMtGDfzwm2/EYdVMamQIrQ0ZXlv5xFo3DzcqJdyyWJ9WgzrRRJSYootM
sGOubdtKuvsNrHi1qQATt2rSeCz15VZlceds7y3HE5yAy8yP4YzHqcF3RUKLmzL+
jJ1fruq9qZ+cACl7xbI2Pisf1KVG8ogvhN99aJk6CuJGmknpp18DTVdPx36rjEI3
+GqrjYFtJq8FI+q9sr3yJLUznMu+bvHRlksJRBOImgnGxwUx6cJjznP9nYloHEJO
bYrcIX3EJqMAralkuC8W2QBEwVkR6UUEsOSkALmA4/Rx968Zc6w71DsX7ETB3O+g
dSLorjHw4I3pOy5wK5qFlBo1tMnk3zhrCsnyN6rfZInM77GiKggKIVsUcyMqSoPj
ZqbH85mhaLKy8WjiOZnDeEkVh3tiBl/WZgCuOSA4aFV5EcDk9U+2tUYi6o0s/taP
n/w0sbmXHeWtj1W/PktT64V67Qa1m6Xndy22zXm6MrzR8bbROVRByK6ayblVZwm2
5IeBfcrX8Xbq3FrLJYH0j/mXpPU1HPAdtAszQ86JgripFqj8TJSdXVP0G0O50PDL
MWoS2mRBMQ/aXza4V8iP463jzIdzf+Npot7gxeYjet3nXboaEEeh+2QFj+t2f8wy
KN5CHap8IuCVV8wGZzI1wAJaa1l2VFuIdaumzpgyjGJUmSLbACxAZrgkwCn68ktr
JQYJLB1Z3GyefXY6TaHbxV0FTMfxoLZZXShj9LiARLi9T6NkK51thZDhJvizt9du
FShrOFIgFBca1Xr90ubXw/cS4izR/e/hqbrqseM6vTDAc0z2yBPO/1puPD38IpPq
bjIVTIo0Swe8HEDckVTWhWCjAwpC+189/5X/CAB5zGQsLjJSEWwwA4W45B157st1
qZKyAO/yIVCwZTEQ9F8S9jA1PObKAzX7p4khfhlGRS5RjJY/d6tRYBxALhbJXxVi
buSMRm3aPXN/8JkkM26KcnozCNKExWlpeR+x/hDo5gfTiJgK5LeiC5hR9/A7mFcJ
vQ7gp/KScPlJBt+jRSd+HD+bNDyv2mODLaTP548NoOGC9B8Td7en3OWrmciFd7VD
FUw/3bIH+mhliVZUa07Mg3YQRh3vsubOytpzf1kcIoNZ4Xxytr3sVby7m1fjNFKx
+bURNyS3ZIE47UMXITPNIAhIu6yStcLU6trbTyB+oAbaZ40d8XXHdeBWNw0b0RHZ
/Y0fm7OdgHE+yrGCnIeKkLJ6UlbMg4zAU58xZ0YcM7y1Gu4LVhiS50i55ZzW1NaC
z0wPOzyWXrkq53/cSTwhXiHs3Q23+NI2e8YlTLVNhdwC0HbygxEEyklBePPYcDam
ap9md05POjBaN8DixPmfwXrEAF+LS48LHPBf36IQBT873mttm5hgCOVQnHiJAxfu
b8mH9LsztAi/9KYoY22dg8WOSwP1xupBg5+ZwDK0N4DLG0gclJGfolxdQaI5QXfe
9j0KbW69H22dUOSgF8TuF2I+MIaqJ2T1zMYKhDmDW9csU2DKgasakkSQV6UKQhFa
OWAtGmaXoyAjVDSS93bFSm07dleTTa82tQn3YW5mRhcnwoO5L2TBIMj8Kbk03WSZ
LtwWt3WGkEcI1LGirApGKvgV0yzv3ubBJuCD5bbzAHDnqMn7JNc0fEv2FoeUHUqL
H0z673fu4q7U5TGwjUx8Dnw/nHgLIYDtM24wifCIoVktin6cHAQ4cB1J9X67eHPG
UHEr9/M3oE4Hf2q2syl/iapHu/ViO4Q0w+Kb34gHl4bGVnKqqz997iuVssztCreC
FgEg/h9TMUT3uY3a1fxHrtjVZ9mtceGIrBBBwZKEg/Q1Lb0vdqkxqN8w9BoQ8EOI
S/XW/5FeyRb8S6ZKnvFja9LEq987b2jId4DaScXFYidCdsi3BHyiirYoYfNmpfD5
5K96/R/iyZgzP4dzDBvCKLOnsPW61LGy1KJYWbpI1jlA3D8NpNKD077dC+DC+keK
dQLalKK8N4HA3R0iiMJ7246TLdQJGwHKARd+AWwQzYt52r/VutmG2WauMb42Oqqh
pRxYT+fnc+4judUL+wJDnaBrRU45+YAC1kWEGyCY47KeP/g8Jo0QfPP3Q2l5csll
Jbm6yzsUNe9+c2T4M7mhIykkJnQ585rNL8O9YZ2C9CZRSZ95KOwNdQs24LvAc3/o
Mui89smRcvJTRJtb/K/f+oC5K58nIQHq10YoEpjc8+XsYK34Ax6JykxZxfyyP7EK
rn1gBE/raqBWyS2rkzv7HEKfc/C9aaXmo/FYAAUPQMW82a8etNVusAwtPMutj531
5OuDM2KrEXEd+vKoJejbs+kI9hyAAkqqmBq2Lk64vxa1myLv8kSHs8sduTUrRcXB
Gwzi0mcgvTj79xBqG1un+hB6RRWLXup474JVRHVe6H4NMje83q2vbTtQYm0G3+61
6QDgWILdZmwHeFuPqJPegA7S7AMyQPIfqUwwCMURQLu/vi/zQB/h50HcE9cBBuvg
D4ESgvPnPi90ayiVTBzxBndYu/MibqXLS9jKD798wQwgT+so5Rgg3qwTNP0IRu0h
galIHJm2Dm/D8kzOrmISn41fQzKHd4pyMjuI5GpOo8spQC3A7jzf9XcEAiCrtRw6
faK9m2XJPbJX2xbam95CV/LOUi1FvV1xpA+lQyJNi4GSqi0S2GWLMAF7w3ZT7ufH
UKyugxms/w7Cbj96UkcRHbhpgqSRyG/Rrr+w2PDvsIY5NzuQfBI8DUZsMnAlzcPu
E25XbtHEEHPUqV2IXFrAYkozjoCcuo8isC6wpeiRVu0dNlgOgcBiRyV5Fv1SgYch
fetycA+6AeihVxNPNh+btdLhbTyfJ6WvhuwslJ6qN0S28mW4sGd/WWxF+Yt09A+0
XGAsraG+x6Qd/yf5PO2uSuSqiPuPZFNTHoiiRzxYVsV3VxX+kF0EAGzb88nOF4X5
MRt4uJxILEFn9saqRVuHpiIWg4pOwSJEnfYYFG65xmq92QS3Q6Zv8qOqadFqk/TN
DTR5Kvp5L3ZcPwEX5c2LeTExPE6LG8oZLlbYOiVadbu0Xh9a9L1YMsPOo7CSHR9z
rs/64cmvmWZNdoaGOHHU4csvu1m88gOX73la4O+s4TfWNTwCQhlshwB71XWD5E8i
B9uGtyCgM+WTc9Egf2t9nNjznDSylJ1Dl3CB+kuOE0+rup2qHDN+GhkqXiOBN4A8
/Cytb7/07GAP0TA10JT5LIJEHld7p/jSW1JgcCowWoiIY3em1F4J1cYyZ9SzKJtc
hhNLywX6YFp9LMxrcD7QhFkD5Sv02P3BuKCzepSSYJbfshpXKwvv7RXj51DB8qYg
47StZzJHqyNDdv1IIHWqLpHbFCKlrl2t/nXGgx4FJi0ias4rnL+8FDKqXIIGV46b
Wq8N3rXYlvXg0pc/YSYk1SZx6KbBKcrPz/nzOtETQ9iJLJza8RAVH3PRuAOP9qoh
DysK57x1aOrXC4uHopQLJfevYp4Z3b5rMCxIiPAmZHFFlEZy8CFVJ4EtxDzjw/zC
VFMcEA4wTXboBEBeX0wF9m+zCxZM6V6yX0pQpIe6jTfmMwo6TimDGr16NfsUGw28
zjcXlx0CjKxgdKLITMBk8hlpA30SMixexTpmVfP1pGMi3zHJrWMieT6zz4NjiCid
QeNfyKUp3Lqs35iw8GdiWG+S8vMib9j33uMl+finRAWBrpsXvxGq08UxyaHKLAvo
NqUk0JYauPFxE26x+uanZbwC+bpOw34T5gkWPEceOuasjrLfGex3fRAA+Cq1fIrV
oBOTdZPHGzqXGyPuoDhDm42P9sUyiErr+pHDULSfleoy0DhArigj9btr/d2q7o+A
TetQ0zFs5mgTuNCvKvednrkHOewEpB63Hyl87uD0QyxxLtprYOH4u7E/5Y0WFvib
v9uQKUHD4AwS5/ocewIMxz2BRaVn2CR9g6wj3fttKTmGpRSq9920yKmvdVNB9W9S
Qjyo3gYcUZz9afVXblYuIEPIo+EZmaZttYHoWvzDtUORzUKik3uCxulxoLSUAJzf
huPrw6AXmSQzWnfNma9bE2oPNhikxp1iuVLPzgvQDdBaECuZTysB1Nb/Qc2fCsUp
d0nQQgjtcswd8FiKmGP5bJw6JLj2Y2qv6URZRvHjJc/yXs+8E6HnT0i+jgTxuAWg
t8aV7VmiwT+RkNphKNO+leGAiNYX9+HC5V3qU8jojvd2373pmyYX2KWZWyjAQNgB
CwEYPAURX8thtRGRsLk3vJ7MT6HaeNT71oOM8XbU7mE9EAuCRapLgk4neTpnRPDQ
S/d7SxjdCLPsrz8fzi1ACc/lv5Zn45Xu7W8a7NWjZQXOvHNRSYy3VfBl5l4iCN1y
KFW1L8egicfzD05ODmTFMY1pMaKoYGlCH1K3xuFIIp8sSTHvaYHcXqyg/8evLFmJ
AZ3KYgSoal5nmD26CqP3t1qpa3SPMF1Z4k3LFySGsYdA+KcNHFA2+gWwqrjTKe3J
cwb78Sh/HHNq6Tfn3vlIm2iaEiv75tsrN752s62iaZLFEsTnn4nsdWwPrjhIyCof
//P3MyUaUxNM0O8O2TJ1T3Rj5UyaaqBw4fcEHtmBUD9fmAMxmvEZ9lXfjk2/QfYx
9kVcQ1axNJuI6jFJeS2Yf0Lt+wQaUOtkkhPFC7Di0rZQ1I/pP/SjuVL/2ZWAHxGH
RCvaNhfQbtpJcOq0uF/NSveIZ9Ksmpv0qBTrpvpey+dduxR4D38T3/FIjjq91T2S
9X4SjVHyLwGTV0wTcXoIO3H0puSmrzE6JTPzCN62WsbCJoMHdlzwl3bGuMUJYM2X
jeYUYzoxaq0pZi2xpHecN7QyhxEHeLCH19DR/aMMcZ3bsoimGBOr1X7563Ik5zrR
InThbrrVyikRUVVhunhFKqZxDEzI2Fa/ttXuS4FBQfLkb3gcf5roCgwkYaBWBgUd
5FYSqdmpcVcaofo1TOGCUCvhkQ3UvQOfBPmXGlENNc3e1oLit46aPysUgzuDvF4y
xyyL8Ft5Kp1qe+bHwuGzSb0/deujSjIeh8HqUAhTLmw+FS6G6L61S5fHGIG4S1h1
Uf6WeNvWji3cybJDm3fZf6yVmSP7nJN77OcWtcdkLc92eb1fEHff/V0sOggMKzhb
bYfWqKxVmyvKHRRa2c2/rNDuV8Z0I0eanPDTvARMi+xr572SO+Szvimij5KH55Lj
B1erSIGBNSGfCz50T5Os7fhBthmebJ+QBdAk7MZB1uWUTue8OERt2wRDy3L21i68
s9qEM5fVwSic6WruORcj2R4mh8bIP6xMZ4ZPMD1dm7X/bBxBsEWzfglyQqZHGbTl
YmkGyW8yLhV7DZ1KWkxrf6tA/AiwqAMJZtuzO0ld7Q/c7lvopERbqHS9utVJl/hv
tymW9V/SjwK/hdPfiemltclSCw0oaUwsVJqqif1xA4DSZfRkvoWRaJsaDAifjgzn
fTRoMYTCP36w4OcalI2UTjEs85Vs6atxxfn5Sp/No9g1xEdbBSicLFLH7xweRxUQ
UFWxB8n581ObtspHk0wYFhiU9S3K9PHarbGEoRZs/IsGg0GCEBS/WAWfo5P/iiFV
HBpW+U41U5QVAVP1n3KUnmB5N9BLHqgylyQJz0DSov8NlvyRuIoHR296XzCbgWqr
pfBiHobe5gDahBapVlpJPVZfga+0IXF+pRnhzuj/1sXJl8DEnjSXP0GxdrKnjnve
4lSw78k6ZLMWLy8br+K96qOeSYvDth8c00cIBKdnMa4/Wv7/8QYiVXk5FrJCPwc2
wxZ/oCTSWFvoND5zFICx8VETeVkZplcsFm0PmmTJTpxJrLONMrB35F8+T8uxghug
Gc/GoiQpte15f1L2uP+J39FSBtus2fu4po/jUdjZhcUNeHfp4AxD0a08h+eo17HJ
DZAfwUjGeEb4P1f2QHUs4aJHFFPzcfIrKWe2ylYOiB8wv7wnD4AfBPKHv86aoeqS
AnO8/0XY0BvNSL7HnJFTB/yhLQ6XUQ1K+0/48sPYSsUMfetIXBTdeRgXMTzRJdZ1
qCPBge4ylYDlLkxejYjWf+meZuYiVOTZohh4sFuk05ZVAeBiJzm3VhNEJyjBUu/q
Hibp4on4dJhI9/zyQezkGzynEVqZOW/xr7j1l3emcwdbhc9B4qQfZeurGTfKN6YC
czjTnzpg2LQrKEr1EaTRQUlFSJBkNOqlQDsG74Pt9qTCR+s5+5FSOqtHryUkAFMH
c6pqb/jiVrBYPtvOzk6YlQTtvzHxdMMiWltr3KLX5+a3aaV40awjmFwTS5EqaKWJ
R54IsJPOo6Qn4JaN5zGqZfv8+WEgQknfYOkvDWImoBU2S8fzYWUkbLzqCYpEjws9
Vlxc9Kra5jKMYx93U0SWmGw61+Vj6OQGXp7dTtir3kI6j6+2sYcVAIPF2xvCZT8A
1yZIkO1A9Kez5nzR6ENKD47Ot4SjF99BmJXf1JT8sZutfVcG0W4rQ7ItoMB3UmKz
lCp25DDPSHsKrPb56AqtB9DM0Rgptkiyh8AXRs8JYcJ6xWdbMyAqV0/E2K1LfFAA
Ox2+MTHW4C/MtjLB1qTBoHjgKLFetmWGTVviMGgmqcAnyOjF29Oi7LEFTSd1XSNM
koLpXXLG3xh7znbgXIbSADs5+kXTX7nAaerq/ytbillJpoY31q+SluydRyP1XdmN
N3HenWTM0aQeMCXCcDsMTZq1M8y5K5sMAcAEEg3lpLwG1ojYnnlUfIukaLnaEj5x
+pW94NwoiL3HAIXF037LHauC3IwAHTFCZ/ahlfzDVXYOn1agoMc1xF5/sD1X1XeC
vI9thLCP534NC7fjzwA0J5OZMIDweZAdRRvLa950Pgvs+g5ySAgdEC1iy2SRh2oB
gMVuR8alZKq7Mxha1eoXcvcU3ViCLb8Snjs0NQg8eRAO4jnKh6T0BiGruRs9TAwz
4swy2o6I0rhnBP+ypGjxo6Yre+I/GAjBWwvCYWJ1tc+x8v0Wt2jrBGiCNiWjAXBp
W542b1ZOY8pgo/1W/7o9Gih/nSimgjD1JqxSXQ5owjM1+h+TBhZjkIQManbPCgWf
DEnDJTfLMcmnhTF+XCh/je+iDD9l3U4LmopuaZsPvQUoT+eTWso0nL2J7H8AkQ8i
c6p7BaI8dn23hu5VoIVlxdL/qKncYI7R0v+uOcxsDND6RiVy5gOyvLRBoRq8Vttd
fPV3OCEo0ucyCBz/bv8X65ZOdZ8bFKmUvrSF4t2SU65mda+l2PTYnZPYF4ttqoMA
MumbXXkzIY+Zn/kx4nFfHRnfbgJ0V1l/piqJsfpvKOK+4psnRGkjERlCm4TdsNxC
kTEZTI913rxYSCUmXBnP8VApj4sSR4sfQpmGHiLuVvEgmHZo6Ol0xzpJ3jkjyDZG
8D/b28cD80FtLe6VAC3Ig4qSoocIzwKk1uDDDzOCgw9SywrG3CDZ2P0mDTVnjYHw
FXFDcPqN+pM1acw4Ih2Oc/rrgZXFsczhkhycs6nDXeAE+C/HY4TP79G9UlVdViW+
bWgkxxOJRnuzRrMh7gHzQ9iIqzZ+r1Uvw7E4299/8tKJus3GS6Xl94faGhQmhQo6
AKN4Inx87oMvBIcGtRvsKhXWcO7hUbiLra2xFpOeR98HjKzNYSDjjY2vlZwICoZW
rMz2oA1QlSJVtQ6b2SGIzI60nfn+uIi8I9UbAgokeB0pc80sXGJ13PN6Jzpv7TM/
KH+EYL++wl5hPf4RG+MgSW4ehrXdPdwUA3JUcUH/TZNZcSvKAKtns+cAn6NTw58y
Eoa21//65FvMJ9JPfyRe9OtDpywO7MqbaZep/oXhiCMVHwRef2eRzaUVOaOXiRfo
BnIS4IH2eHdf7/Nuv7SxKuWnr0phV+4Ck7D/o9i5epZ5dGkqrOYXtgHwF8vpFIN/
RJHw2Js+0aXoySsQlYNZEGQiMy62oXmYNuGOQum4uF5X6rGgwc3IciOlH+mSI5+w
7TdJQ+oLqb9PTMYvMz5tkle3G2G2Cl5BZPZBvlMsgYitRt0A1ndE+T46ACJqK8So
uXXZjhraY+suXbfvCmmWmzwOvFTN9lA3B+99/GHmNHvVKBIdhvMefqQ5ZLUkdLOW
i24nYe+y/khmZzO4lzutzlsyHcflZAk/LFGB96ww9ptTSVMB/gk4YfprfW/BdNKf
nJggMfN/UzQnKxTHawMt/zU10x/HkXNapx6Vk1lggeaBYFYifk4VQZjHjBiHJnbs
0yIuHsNs8sQvr3zVAno1ByBUnWWHYDUPc9e66+ocw24pgt53SL74Vwm/Zm5nrDDs
ech/E8/semBTasF6bIaF25nWaiLBgjBlZzHqeavtcFdduIa8hotPu8MoAFrKt8X8
D8cALiP2vRK/BCHqKcZ6h8l7F8eDz8PEsRuxdYooLIKG7oX4bft7mwqeOYMSGVT8
SBrsGNRyC2QYB5DjDGolpE+OJyistlgxClusK8zop7R4xPLik7qXT2NC+jxLjLa1
rWSWTyCyawJzitRcI9P8/nki6vxwu59radPdhYwW07ucuX8lgFWKWdSA/sIoFMJ1
7iCZGf62mjwP+bWIdHmoJHdXH8SGipdlRNoHamEFlJ8vjLwxkV8Hz7vqYO/2Uf8k
2NS0AnWYQocB9CxHYkIZm7S7jBLdoeYWXUsVr+p4vyujul45zl6iDQJ5a+RgNRf0
UGA63xbnipYRpYYCla2Qz94068ka9bBgUIEzFgc0jMGUqAAVjtJNTrJD9olw0qbW
xcnUPYI4b9YS4aX0/LjWFwCsCTu6w0jxJwVROLz7TU3PspKw6E3isnzONuAEn2R3
XNZ5ztp/iIx8PlMUL2CXd/hxAJsV7IU/cfBapHWmWg1tFDCe3l4lB0JwuYsTIUXO
yZb0uUsBN3t9puf3ScZfocv4u7TDqRhGtxpx/ja/ET8VzSfr1jW1sXMtLsA4Ty+w
Q6uenL8jqGawFeSqAUCmUJiQRjOAoC6cSHW9OQGCdl3RteQ2Bvi9BlR6BcGUQslJ
RaF5BgLxRgMO2YGtcAUsVEe+bJzMAkt/wmo75pXOSb5tXmk/QRbkGuUDW0Ete+q7
NUU3+z2viehwgGtNjsI/uPKbab5OJpGBdTg7ZEZ1reFKaFnkvJMCcTTYOBR1NHAo
wS6hyRvApBOkXVgkJtuostP+F1p4BovYbmNQR/2WMWkI+NAmuN6EPwexpPVnn8T0
VHUfisqZeEOpYE+GZagSw145kEItTXH9QqEZvzyKp+TA2WyP/zTfvwT0p6tOEzZ7
AZ17po7J7E5WN9GlviFnikHFIIzR3Nh0nCfuzWBFcmcdwg6ckLPt/3fuWsLoZZ/z
b7zZ9LLQBrmrPUVz+rLVwujj9Supjf5gsRm/oUaPKd/AGRvc6N2S9EIOozHd/jK/
AOnpowUIfs1HrhRF99p3edfk9ZiFEcu92Obkqcl2XW+guBF91Ui6E9Wh2rI9IwqT
TCdH+vLr1MBDMa/pVyQj5b4rLw90Z+E+ob4+DoGnecsMBqkwAJ4Qff3oU7vZVUIX
VjBfd6UwK4S32VGv/m3hfW/EkPyDRG3Yh65w4CgK4sbWDDEqViZBq/FdJGRylVJV
Ot1HRtAxbGr0hxXbhOMluR1GIFY7sEdAXPs2xKvDtjQqecZ0qs8kC/lmWQAt0pHv
gfn1JIXQ1ZXmKwlvf+gWK9fuyKln6MfoQZZGMh8Lcr2rk4BUQzIsfT1yvUGAvkVw
F1xFAy/R9vZUFDpoV94Xkpbpx3k+mzqHj9tohxbMlfCrFKFFGWEjXXC/kijj3z5j
Me+sNddHHFiaj9JD4IhFAr7X6YJqZatOcoJrQaRILUiHjHVHap+nx0/7b7Lu+suF
WRYrNRJwZDt+13uEv4fibBxTPQF1776hzCXyf40EM1dPrOdLaJSC4Caig/8HnT2s
4SNKk3toZGYNmaCTZ6Q/IfhzM1R8+9H9MZS6N4TWge7sf4GhnDxZ81TmFOiIdXyK
ajRikgWGZtx3syzbSFkVDEdNECs9FpYoEsNGWlZ9OuZq7zfTiBP6nsBpZIy2GLMy
QnHLcfPf1M3FZgKnQsJItPLf9qkhIIe2+ncYva8mxBeiEnJduPIPAupVKnn3TdXC
5r41QbeBkhRePnD7CeimtBdAoGdy03mP903vhqJ+RHufOFo6C4McQVWoDLjAMcBI
iUo/2urPNGGj8aTFJqGdT9+7dP+cZJAlJaDDdr9Fzzam4pVHwyeS9A+cdE7NH11x
lupZ0M9Y6jQI4RVGkTSuGJlZ4OLxI48Hdf0l+EbemErUNp3Opr+WSaMgdWXW4pQK
cmPHCdNQycCjIIt8p6JCCYu7IkjLO6SXqKBj3StEE2Syu18Cl3WDo6AOcdC8EQIF
zVBbGMdlPj1fpMB2HyoXix97t+I7+AScX/4v3EHvl9n4DxDFAcL8i+viPZuTHkwd
BjHMQxnujNmO0r+h9Yiq5KLlTNvpv4JzC+fi3YLRxXl4pX2eGov9nlqhRNPOKIHV
QHUCDE2YkPzyjyr87872C7DpPyLwYTWBRRGJEFNXIXZxb8nO+wYkJ6o75tuDC26f
2uk45VI04QgrXolU+5z10bCKcCj4+e+s9Z6/fHHi7tPex9Rt41GZd1noUOr30VIR
1HN1wGG356bRJPkikwVpA3uIHkKwaoseLoE/mX8iZgQm775WAb3bvKMkOJKMsLeA
h5bi5xH7Z+hITpOBE027ndJHYR65eI3T//Gl0/OIpiGAAhnJUwsMRGSlJrfJ5oZV
ZclfTLqyOjeNwqcDy0wJkO3co/QplXhuAOejrjCppg/T+UF40bjGPY4WR7nwq6/F
4jaIGi2ArHNCwpa94ZNkT3GIZ+DGzvQmwIGKxwDOfEb0F0JTeQHOsBPEgl8DEJb/
+s0vJMVgdICCcJYKrNha2ogQdDWWSrZInu0IaGEJvWVjx10DgziW+s9R+v3m173h
iy/hbQlUkyT2a/PJHOIaDqnHCJgarDvZyhrPkO7eKeh1vCeShnITeP6t3kpB3Ul2
/iQM4QuEDu3eSQfszjkSSdmQaB9PMGpKbqa7jqMpqHOh1x5fYQjXzv+M0rHj77cN
foaCuv2wkDuNw1kDOofUcFNlND5xw4nHZkeEuvzllXVLtq3eEFcgB0Eh203ZTFKw
VwH2N0+HitmyjHbglznaCRnaVWs2YBGX6MiaUxq0izx9TYkwaonxtnjxwfjR90m5
eha9lWBRlH84bkRST8SO8eWoi+282V4zulTry50X+s0R/9OL8qBkeYm3YLGe1Vwq
yV/0l+j9hAQxVYPK3cY4ja7/JTXGkv7OUc9xdXhjtdpalJt4ylbRTIO0WpgKSsAL
0DRE8G+tSdjhXsdm6c4xcWFc6Tg3ZGCWbhVzFrAxGGkSdYdcsUgOiK8OqHm9LKEk
nQZB64mDCe2/XQEWiUe9AX2/WOj55YgxGBHcQA6BLyy4gU3sk8dGStgN8pSeW4Mo
6bdVflYmePdFa/GAcEx7ZA3UH1nFrFlWMTrJQF3y0YMGQxD6Y3GOs1REBpbEz+hY
L8+QKU7aQB038H0svvrkYA1aqsteINKiPqeHu0LsgSGPWeuqWhn+pXr6SXVhnm32
dzjdPOXOe/fMrF6SaFp6kSK0QXx1FV3Ej5wsoLN9eg4Rk6cs7/To9RVkkSF4gfRC
IF5jwuIjGWwRx9Y+akAYS+5PNvFcKUVqtEPNORIoM8QTLtGL9UWS8Lhs1XZlF7Ne
ZyX7+VWMkd42vGTXXwXhs+gYnCkdHh2ugkXODxzDli97tmIO0ux/4PE5pLyN01hd
W15M4AusL+CgMS5r9ea3pIlxVRGRU1IAObFyZUs+Om3Rf8UgFkkHt1We7Ic7ky4D
GpyYl7/h47q9GXWqlHOa2lr69w33fZNSrP0OM6dngCQvtCmvhWI8p3EgH8hG/gtQ
Pgc5+dIcizcylq/qlyj+QfQ4MO84vyrD7gQH9xo/9t5RLxm+/06ravSoTaXj2BGM
5652kokbOCtmgKqwC8ZW/0crEWviHE3SAzpjZBixRoGuHnFnubN1npzp3MzqPvO3
UCBprc2+WTxCVMndHaa9SSP8IDODM1weaK1gV6Bl4mZaQ7aNzGCfE6RR3TXuIssm
itZvaBBy42cUsGAJMaQi+OmtgtRagZ3z6dGVoeonwb5i4DIemk/zS2G00g2aOVYy
CusLMbfti2AZrkhnVd6AaYLO+f7RTsNs3rl5d6it0LS/hKQg/IzyN2asHmnUEEbH
Af7oPtgwGCruZCM/agWGoxW8y+Cao/H9xpUI871qknvDjSkum+ZMpl83EBikeIDw
0eaKaekKNFr8du09A8wES8SvHksGcTCKYgWVi3ngsrA/XBy0qxGCUPsBoZdlV7Di
/U9mp0bAlFw6GfWOMiSQstojnQoNodyT1UXIw9Nku33/I7ZnTyKOFBxTcLSKV6qu
chyZvMGE+v1FzssIduM5g7vDi3ATM4qyS9gNBgVaKrEb/1fnYmFB69MPor3XenFB
de7yb1xebPsdp8V0Ib1qc1iuDBB+VQC7MUjKhj5pFh5/YQNNGrokx6tMnlVF0gDt
2w/EL2KIW8IW2mc4+l3DlLFbl/nEd4sSdagiPEc0VAQlP2N+Warmq+Gcn2T8qaGo
dzKPrqnF1enO7XexR+XYXMg6GhLDcyee5cqiDBdOycAfS91RkKyRXd1ZhYqr7FDg
6hYa3brGEsEsR786gqPfpRSqwWQphd0fUtfJ3pMsgtnKPtM1W4GLE0gZ2wIrUXu9
Wasg7rXQsLdDRMxOaFZsgfVYz+YoXfh/0+x65P1X+6J9IC5Gz6wl8egQvEQX7SNx
QO+nGw0muYjJajbcqawgDB2mQJnY18D5762uEPHfufDMhcSOdxFRiOWqg3Auf9i8
LSO4DLSTScpMAzB0mXPVu4PD2SdDdfqDtnaiZbtzZbqbRlVbWG9om5LzH+D49ZC5
oA55/UTmb4Ci39aIKv3Z0pVnsaim8ufeawoZxhfrXHKkPjMugdbW/fVr05mdyCGP
4pbo3kyH3ntfB08b4/al3L5POxVFCauKYPrGZhdB/kIyMM79NZ/4RaP/4iu7v9rF
/kI2WC14VuiAta6o5wwwYor17B2YhKajOAaQ9KTrS+saCVKaXQ3zeIqc0ztDNnKE
vBNtQ6S3W4fZ0AoEjhuYjvoCJzDp/Qk2MB++Xj4Mzdlt9hyQFQTWcaMz1A/FpGru
XEJzd3RCW9vKHTfH9MjIy/dTPDEZmn+u0CMLrcvxUOi7kcEWuNveZBtDbW6VogHt
eyxjBNz5WtyAOdaJwvMm4sI6aq2Bfrm0OpPb6AOLHqRWGqwM5sv+kFuaHhW9fGWu
vDsfzOtabnGwmJZHOnqX350ttyz8ARRk5gq9n6H+HNDDa2zOpiMzblD/2oMcBYmp
ypqBb9uvNpuB4zb0l5Lb6IInqspqnekv/Vdj5Qf14joRF58hQUShXaBLJyH5YgA+
NoHq/OMwM6ydZwJL7RdKp9vjv8czmqOt9ZplE1YpGl0R/aFdnuyQWh8nH6fBGXkc
LimIIzMpNgPp0H3JAjNuiT6cEg9m8qaAPeohzIuCv0zwwdkB035NdAiR17SXKCf5
IhoXkRaEqMITo6E0V4NgoxPmNWr558s4Uj06pSvlU1BRuSc5izuK4vthWD0e5SMi
L2kQbShMu0MvLSv56pmwO7ry7QbfHrywBvD3DsLKEcza5np89NIU5/z2pz/mNLpE
Gos88julSR7iLZO05h0VRO2Ig8tsnBgG50A97lfaKLSIu6fYQXSHK2GCIPWLtw6I
d5hZZI81cmkFVUZEqzBbb0ysWZiKQ8Ko5ZkySxbbKGDe6jenFHpikvZ6twOQutcI
H1d/msYPsgqi+Vg64UhUM4ksbyGLviiFGmwLc1rrZW1SzXJHKRZCxwZUZTBbUunY
1BOkKqcBGCspgiL/FL1Dcf7asLxeRKCuZevtENrGoPpW4LHznY5LdK0/TZ+DlrNp
3X2ujvPPiVCXc4bF9sHIc4Jqrdld9IGLZimalXy4EX0zn5e/ZK29jqb1hbveKRdQ
AZK/hWqpL4xTe/DmNRTL/7QXypxXEDDXcHqEPZMr2gbJjShEqUUdmvf11kxe7bJw
UTDs/agU9d7S0sfayoVSDU7csa+ylfDkZ4RMnPWSvB+sxFu2ZRbo8ykbj+47M/fT
3fA3XKOnFREBzhL660/1l7RoFuUHnVTSuez6oE4fdPVIxzPNnFI9ZcVC/Gwz+etn
WTDXw944CrRqwqZ7uvEDJH5Y5G3K0Kw65KYts6lmLvdKDFetmOlpVqKh2iDCdDkP
4rYgdMY3uyCoBU7z+rXlUDsxQxcMGNibN+3XWFUPZCg3c7QVTkfSJeWXNi25FwwO
WyNx+FprjiyDJTr6RQQlSCid2HcY6te5coGLVcmMWduORlmJI+BGfFYAHDHA4POp
HLL6L0uLDwLc2jNhBXb3UZIXoZIz+hlvNE/jDP9ZK9LhfDMBfjc6gW5id4VZJ073
BQQzETAmb/8BI0QniNepC7Bdletg9g84j/S6wwrdaoWO6qVvZJiSY9OEN9kKusj0
U6VriDRb4fMyikAEclfNMqlKVo7/pG29c4XpVDkcILaQ9/diak+V/ZzehTo1aQnE
QoIHUsyKZknbaStn1TQbgiYMeSVyzesfExmjMdpC7K2O6slPf0IWHmmUl6ntt0sx
r/0b8oSDUkvn0RN/IQ2GH9VsDm9QaQ00FqYiRFgG8dZmDLIkdmHZNjyOd4XCvIcx
UHi7+i3/firy3g4BcEw6LsgNEGOWtXtXb5AJf5QDbRQrpTs2GRSZXA7VSZXMmACB
h8Fcr8301EluO23TwE0sJ4cML8oXjNou9I4/csiSTTczPqAWnKPKCliWS+Q+8vCj
Z6NkpCBg7uWMWqrXwTy7f2xyRBwD76wcQT5AQTEtRbe53KO77BcRuIQ3x8UP2vWn
XBbrBAaJ+rI5I16/Mn1vULgRH+xfG7jOWNrGt8n1ogi8eWdnfhXne8QZ0rqKRGbP
wsZlattGVjFLRLUhlD6aTWqP3orXFid96D0bejhzthShBnfGwSFRLsa/pdKOh8Kg
ZrjIsam938sWFulFqMpd8soAT4qBs2rOR+KzWUw3kZvS4jqHvxsGuyLIIs2u9wzh
zdBBfh3IFzoBf7tS/mPP0BQhG9mzUDDYWFWvGlyXbs2lpT8iRm7m16zV5x5ZIxjy
RH/u9UnMuw/e1aAFQK5rz+Ugrkyr0cTCQQC49Mz4uhtYqDIXA4sA191AjKlQILy/
K+k6ylmXreWOmpEORpPPQkN880LaTC0b9vegRw1+bLoLNcS/FStsynAyyKldn1aK
cIydECju5HZ5aAY4i/7BxDuJiOsfV6KJh34ELkMp5wqaUl24Fo6Duqx7NpHD0BIz
4FNBvRTPyJhUTZ9zNUn25tTrcAsS4+iej5wfom95S7Wn67ebOCn4OiptjppBL93w
UDMfXUE8Gn8xSRTRcplDPFwMbMnD/llXbq7ymYlgFA547PiP6PN0N1uaIx7r7rR+
snD2t2PG0lTBS6rHx0Q1NRZOveM0xLEf0r9fxEyeHzAmLFqFHgYO0EWxxhHKZrEP
kxCsL40tMohRhziiipCz8c2uB5C2nQEiFZF+W3M4sT2PY4sNhlKZ17rhQF/Z/OUI
RHl8fsnIYFXdSNU150bz8B57IFwW0w24+ofAUtQDmmc9ImB+x+1apBq2myfDLXyl
SyWD1a2NVT1L1i1wSJv8d6HcGgI5MD3OOVhjdZitj5yRkAgF/2wMaEu2EJQty8bP
Kbo1rNXy3pA2POaDkF45i2CINFDQwC4fUq5QVzW1+gW/gYF7BHOT9674mt3iKToL
I+aqSr+exwI59z1IqGJ9TAObY6UQBTzgXIwFtvQwF5v65PFvda6PvmRa06E1zaK+
IRw8ErmA/sHe2tJQPAomCUSJeBa8rTCOCIGnJYTQbmRRk2Il5yCv4yjfNMo4kO60
yUNfve0dGbtYfm1D2FaZhfdDaG7C4BmWkwvy0g3sLPxTq/q9pALhdrW+ZcLrk/DK
ZAs+x82bYalB7c0KQ9Q2mQpxJ3OopZFOZkv9MDbooCNPJvR+bO/XmDntli3gm6aG
LTJ0qYOHEZWCeih2MG1PpBkXl5b2pmhv/p97vF2ZUjvsPWy/k3RKCFQ9ngue7iyS
/eS9gpxAwP5A2NFiov0m80B1yvTlGziS9MHTR9qOwT2v1v8D+QVah09sEAp1QlUN
im6GMoEVxFfpZxfoiEJSXP695B9krJm4t/Jdp+tuW/mvVpn9ZeyHVJSnyC0nKZGv
nFEqbkV/oDzCco+/AquKYQKPFtiBXex8c2Q/rZexo5EnnC6Ou4nMnT5iCk2rmWwO
gRpSdMN+h1YqQgYapKjjQ/gCg3r6nxvkQW1io+7oNbJf1o+hAS1G/LtofvUX+lC7
BjR9CFiqqXNb7rO/lsVOX7sKZaqRJvycIBwnEbTtLp2EB0uWLD8lITonOfmNvovi
GPPIe3eYm9n69EWUlIB6MJKV3O4vOGUcVMhv6ifAQX423DFQscXjcFWAkKOB3B2N
Y4h2WctQVI4jkhNoPDMA6WTEj9rpxd3P3IQA56eRqhNJJzEP1PKm4G+jhLbKX4zH
LmedwlFe2SMLPyqIMv2fYEJkfpJT5DubRp4NNMCmpIjWqj1ApmG1ZZcs8dH7lbXy
V3hUfQDrLe+TXPPEML3Nc/lFS4+GPzZ2nfa+P5FfaGWSPbSdMamsYWQMtnvPuOHX
S2n76MnlSlwu8tl5OsBZWXe707HAjaa68jzDRfnGTZam/NwgqnNfxT/Z/X7Tuy4S
1RllXKRQLcWjBZgAJkntxHNXPSqlhFGekPRGeg/BySRmtaO5dMeIW4oR9IkLyggV
FXwTEqBik/DIe7FmA0C272JlE5Ip+OlJE97BLiKVQ0gp2GZ0jnRGI8x6DnMFZX88
AnzMkISvRhOKiAg9zF3SUQGrF8B8hbC9uHDahC80pZnM561+IghzYIFTc+sMKhQG
aevW6/BRx9iFjKRGk1au9WMELyVYz1m0PNI2Lf+EC3Nj2u82P+pzN+K+9tvJq3Pa
D1ne954i4H0KolJpJIgf7DXMqvDr9m/4T/jTu+uyF2xFvK1W19SzjhtsApM3vB7S
JBb/gzMAtuHEZTCchi7EbkIvvZAKBI6smGo499yrZtiycAHURYoV2tKM7AT/Dgsv
EeGBMEiIhIMjViDSintZKtuqJCBAXp6DCMapIRQ+CtUKf/q73OXt4WB6Q7SdK0Sk
LfEPjXcoYJeIeyi+KGAHhx6/aQWDYcymAg9Ey+TOCeW+Vf1h8BiI+5JQynbbgbvs
UO3kdjPNha/oYtUXRz+4gN+HcJTug2YRrlahCsFH2Gjr0hqUwySjBmjWf7KABe8z
IkRLift6ygyKKZwGJKPofzNqwzWWvaupRiuDMCyTz2TgKSfmNhciLSPHySEHnuEp
cykipn3/W0VuIT4cRQNBg17za4lTzqllp1DrzIV8QPsLB+sAaDfVxLJedsTfokNf
q93coc6B+z8MY6Zuwe0FxRprS3ZQLUjTRkbBLaGMFb4D7ssTBDgfV9zfbNiYqXAK
lb89gxEdSnzg4UPpcoQlfbRmf6fZlae6uXZLAbjKej77cWrsvmmxJXwgj93YPJlx
8tZdjO+8KRHWaf3ARZXD26tt43S93yTKLgkqQN/WJ4O1TT1OPd8Qf9pk7rMsZSSr
0sUwiJmf8VG/CVwntHBVfZQPI3SvDuRA6nqFRFQQq8UIfuhUNzPsWOWA/OYrqXtp
Mw0tNrnpdl2fGqDuz4bUtfmRgaNPTwwemXxAV7rp5webXhWu88UOFDl2kqy9ub/L
lBYdqHj6s3/4CXwMRxBOx94PFWxaA7HrZsRbrkv7qPCTZFDdWwOG9qdj9SoASkno
Duhzu0uua/LzhUmkCsWJsM+r1PmWCsHhnRH3ARfpmDNFK46XY43Ke7vqEsskz+RK
E6Y8oArNdX/kH+XDSwzbvg+N66bhDqtAnmIcjW5FNY8TCpu5+Z9gBaa51XuYedei
WoznDT7TpP6Iu1K7a0sKwbEVlytOq/JxJpN5VdM8afeYFuyiHtNojWKtgP0A6WiJ
9QxtVIXS4o5Tdzoyz+pVvCcsrL0mNnEtNzZw4lkvYEONsra63jsP+AW/l4R85c67
ELXnQnkT3tSu4ySgPuVONCpsroKVMQUIlyxG3ynZDU39XZbDejlFJirMBIEdHMvf
yldJDBywn7OBaq1kOZtR3maTdN0FSjV7uGFd/XrCh4TclUF/6jSv+8qJgjhxv1HT
HfAYe786N2DdNLviHa6pOb8f2CTqJwq51EPzvTxGFQz1MyEaeH5t7jO4yLpGTVyH
TrUi8u5/zSHL7hl/lH5aqpg7m2VEQ0jLdcYV9qNETuB66hSUvSFvuCJ0AbrNS+lu
WKHXgx3AlcQi0v2KNJATm0hoo4XC0exwdJrg/ivRbSq/C+gpHqHG/Il9l3+vhrC7
L85w+xkQuUKRWpx1ostuaoVxmTlxf18tnpLa72LXJJ0JzdA8G70wI0P+dTUTCNET
D8kCvbV/JKMrGhJqFugwHUCH9fzeO6zSfjFEA/yUIzZTmBqq/uvc2s8Abs6fzbj2
qa88+5QM/8uSLluZi0QPBgNOT1epAsIhzL7zfLpJsUe9r4EvPeid5beBXBSFTF3v
MJAcwCQRhXA4yxc1ZCqE0xk/1cSlSLTVXi2RnIw/1peLUnIZMBffjzHbN5eHNfSv
LDcJPoy9ntk3nCFDp57VpL90+9EI24zL/rL76T/egW0ou30b0t4y2sDheI4Halub
/n5GJX/olu2QOcy2bvQFh5PmTlopSlrqs7igfBIc1Ta3Ns99lrFz3GaURfSr2ktc
VK1ZqKisALPVZI7axm4dXAIi0ue9xae/T33gHnrDhiOGEETz9CAaLbSyZGtTdpWP
gwq8SfH57VRc7wN7nbYGKLU1Qj7eydkJ1gyYi/nsaeiRNWAhyak7m5SafXSGwN7I
ZoWF3fygWLPre07f/e2V5H/jILzT04jRTihuHgZO/WoQt1T5GZBMbxREX9zuceJa
eMVtpRFYa+q2TFjmbEhXWDvVwvIG25ndwK0c0uYxTmXba70lT5TPo2iU1WvJOEDP
ihnZpk/CddnwO5q4NPP7Cldl2CS0xBlbmfd8JWWiOXsJGXmfm9kp+LVhgFWa9Z8T
ueYhGQSHYUbnXHhL8pV/BGMS9oQcpv/kZYkyL09r9nNRNAq1HgXRrgKw2e4mmpNi
ttk3VPkZVAQFIPxbUHKG1OqQcHx3EwC6KUcmWgee/Owo6rBMyvZfKciad0DkbWCj
bpD7unF0yLpCRWf6Sl597FcR/wSGkeEbU/ekikQGkPbMNmz/eWN1czonYhp2rRNS
Ri32zJuZJV7r1FoArRMearwhCTizm4X7fQGM2xtIhLYAaIoQS9kd0L0WlpPrh6Ma
FOCkEX2VpWNaeNUX9ZIpPp1bAJzrr0cQHPE6xeIvaClJ3NZBZ7kYQ9YDryyXYUcR
R8oHOZSArOBxzZECQhRn2P82p2UAk16qVKsNABJH8KbZHuwD6JB9U2nmU7q10Plo
y+Bi0+BGH75t+qr1QSyyIUWdR12s4DWOdvy3Bjl4raDJuXTfJh4HMuwJWhrtMN6x
BcKI7bUXH15IrUhqOT3FERq8C98NoWHQD4iagLaGizYXL6l7oMzeT2lXORR5DTk8
XLvPwnCjRsx2hfKmB9BSzTP0ftWS2r5jzTuTsF1m3tPJBupy6gA7gD7k6DOMpQQo
BPvw4jGSgD4ACkjOCeZE6jGGdo3VY7b2zNJf66XsHsmoT0weo+EWuoIOF96YP/Nc
Uhb+dkrNKa25PhvdW3tUyZfEx2rlJHPOaZbdUs1EDeENdSC+PNaqoPiP3xnDCCo2
QzA1PqZI6eNMDTzHwMnGmq266955A/tJEkcLAnQ3omw6BFtSetNJvIWGaNd2nBpb
bcIpULLQWgLkyaxgOFztmlsjXxK08f1iGq2xIljm+NMneSm+8KCmBBkdJFLtzHfh
wC1tkVSN2AwWxJiBuSDair/hiAV07C1oIndu/qGnwrNyM6obAukKOTa5Dlm3NAqA
NCHKxZ4Oqj2TE4gnC4H96z/xf411D+AnHRbw+X1EJwLNWoi81jvcOyJSGfh3QscR
WUSUD5D4OnRLiXJH/rZgV6yV38hSd510nonTwX8z8lndz+q64tajJkXVdi7L3xiN
NMo+rBUBXmAJhuZDbSAGvnG7u6ZJuucInnxp4lms2Mh1UZmqZ+SK5sA9x5ubEWQ2
11yITVuikficJGmuYSDwi3aJ57La2jFavyY0Aj0K4L5uhraT5yVGHAZG0gl4MlJD
jKkmexikXWdlNAzvBIVnp/LBsqZ92dKJiyW7ji1LdxO3NpGGhucaJ+ZWB+6tmqp4
8JCu/tGER+sxrBhUDAZk5F5FVzU8JowP+LVx0PFVHOeNFnRIoZMTPSyOlWqlUUPv
elgpwa1Bd8XtVxPrqaBEwLiJDOny/oL/gUxf64sssfJk+MgTTgfYQzGHPzKvNVMT
TZPWoEhKdbD4YoOVZln+3bvkhaNIcp4vXzTfvhNR8TZwfA2jviV/Yv1aVkLdhSH8
TaAiRsvFF/GsUI1fmG3uKhaVHzXsU3Iu3WwQmZfpowPegfxLy+k1CL1xmfF1e32K
7FMfxzkzbIAArhMP5YLiYHDs54I/m7d/PGLsLKbKwP5qJl9gp+EsIMUWl92ef+1k
5OC+iL7jl2hJVrfiAUE/0Nc+F2f+SrARuyy02QSJfgCeTOcoP6+GlOrE8rYPEAKV
uygu1Ikn3wYpVNJ9e6CXz9qiw1h525vbsqmGuLwG1lMoxsHINkYINwoX9738mjm3
AeICVXCTycQWaiOWbwchVCNnQTRBwlc6Bn6+TVHJqJNfELqx6LLVa9Klt7SP8DiT
ERsm06wBbP0YrxbJS7LJ7Y9ajTnQu3M1TcVP7k6Q4d8T6iPIB5uaevTLRdiFyO3d
yPvhmlnt4H0IHGrqmfgPE97GAha5wVat5JrR+nqH1oP1b4rpIY1UVRdYaWRHQktz
LZ/otU9mk14Qg/t+WsuC56wCOki/3ut3RH5DLV7z25bjPCfV0+TEws+jH9PcuLtb
160CXmAbKxh61viPZgjQzqPROodDw/2CzHlNQzceGuQ7v+M21VD9gmJ/LV3ag7GL
jycMRtrNS6Mdkh0cgAwyP28BDiQc/u46YzECjRZ7NS/s6VGpZ0k3nL+I+53en8y9
Fq4V8NhinDaBUc2connwbcQZjz7FqTczB72ER4aLzVN/cJz1xs79oSGQ6b2nOVty
oFgCc/LCYRNzg2NNVO3u9KK37I3gg8MZiwMbRiSROqAouJ5i+XdYWkD9oeOgqnXy
VQzN2vcZydqCOQ+K+eUSVOuBklYIxb6WJHea4s7Sn0YIFDt6P5PtMcClL6EbPuDs
PzPb8gKrPh1R240ER7xVqJnL/lxZQqn9lzfDfsFugQyVmtCYMEGTAcx84YWkGNqb
xpeSDPH0jUQ1piZ5avy/5pPe2oaW+uBFwXz1clbfJFQeyx5VBaDsfy0gnSMgPTw4
RxkWsbmhkoGO7mm5NpDkyXOIKaATWzE5buSwerFJVQ9VXnb9GZ9AJi1jLk0xEtS3
xQNKBYec/yvQc+lhw77LNnaR7fIOQcjjtJkAe0y93UooCKL1fgLsC5eL2cTTJ9IF
0+Nce1sGlNlYPF09VSVg+sKWLDES9YY+W75TyL7RJlqmCJPFAx4yVmsiKk0Ow30y
3E5l2MGqDMNXJMIjbWPWdUDxk0MTXqJixXo4jsiMjOfdNXLIvUL9ChJ4m4KkKjHg
K+gwhjfo12TUMxd+oTYjM+Oqt4y9nSb3/jkz39ZASYvwQ3FcyBjBtIK5LxxEMnDL
yobfVajAYXitDtuC1qw018qVwpzcxATZXG/Iu3Kw9AR0mrw2RLJjexB29iVubD20
3iFE4P6Gh5NmnrPZ2AQ8tDNb9o8trhD0A1+He09N3RvPJ7ScVHe7otQEdortnV+y
rMNl8VZdWkIGrqZpZ9rCtTZ8AohyZdg/EiyrmpCQTFQEpKVqNoRuH7J6XUaZXspp
fP4zMr3AgrSIPe4LUN43853+FyPtYJlSsygEqmgwa6T0ODa2YAsLLsQnK/IyZw2M
dY7n3saYYjJHYuY3hO3unx27xUBeSUDuKOgmybTrwiGW8EniAHdiK3yDEsM/AhTt
7hpL5DmAFbw0+5hBHvA+vfNvbmFRrj/OZL5HPYDQk//y7kjtyWrfGU2kCiiXZjqf
zfoOgnBBb+Yt2lwLgzmxBqlt8Qy4LX32bx1kWzMUhOu2klewZB65j8LU+YT3Z7Zh
QaZFf0szOCUaDiEUa26cmJxV/2MqAjcwW7H+/+NAtegEKZ2xlXDYwdHva0f6iLLb
YmaVm+r8bRIgRPkPUNPycl7/Q76+5sQEc+qrqwMBY9mLfqmMBU1aPxOZEu/JoJLc
/7fylxkZLIGzxPZVUsG4zlbDi2/22lWm6KIolFtA3LJvFIWw+G5r0X5K73Vy7ev7
VjLz/p0LRFugLVrgXlzirQNsej2Q6QyHWp+f8ClpkzGlgivzeI3OBjWkS4UGuqSv
7//uV0a26fVmcCLiaL4MixdMZ46WOPeu+h6eUMdoOQAoLZTEIGoauv+6DXxfHrEf
vQd8LE2X56fPLd+q0UVeeAIAXR0qDqO34+aCWSh3hUAoguydwjpPAL5MKi3JoyWs
iJ8otDFIXj0/zvUFW/Mvr57PmbeclMq8BEvyk5hLk+OsQbGzQG6MXY3JAZqKzk6d
1JZyo8aUlMKAiYO5hXQprwok/T8wfR0NeNYxcQQ5u0vy/WsFR1LhdApmqY+uc31n
mm5oIv1lpXG8hhlFLiZzTSIixGQy9pv6zsj5JS+ZmSgPmXp+Y1JLAnTW7ZnqGjrY
lC6D6+UIFINZovTlvAeRX+2ydLFYfhgTsdovwnijvybYy3NPDH+1a2d+CAT4G2W+
UKdkFVSqbiynNnCMD/0VFrRfbBeMxwBUp0B1EbJkTJdlX6rsDH/YhK38YfpHxCYl
QJUWqu8wcWA2DTutZpZNFKUgFGJq0IvMmDJTHG+YpHZ4cmn+bxNC4TCF+kqTihV+
6Niq4zniWKAWOHtHqVB4wRczreMqs9WcGlYxpOjDqXh5EONwzMKHC1jR40C3y5Sg
jOFrtHEvI/xmyMJn9uuUxkJSYdun3PNvKNAKt0ioS/pEBLnAXT18UlVFTvmcOEro
A18Lw+qLk2LV7G8C1bS6iqKysrtJ93IOjf9++jo/0n2PRV/F3VU/gU3xMQpZynpf
ghaXOtncC0i2tL9NxY7YNpXHQM1CCne9nSeqhlCF/OL0xgzxvWR2cpSfMxPmT7VA
5l9tk6BDZzM10FlWQbKkhoXhsHDXdwLzP8U20To0ZmLyea/DbLYrzRpY5Dto89Cr
t0MPckovnhRqkodKkGRN6/+kVEcIwQib54wkGHQJeUyZaF8zprFyvTTvj+oTiw0M
IlkfuRiLA34NslRN9bBD1XJitcnX1zT4SWcmLnTIQz2tZtNjwjF4vgPNMS27N/6H
fcxNV/hNXbT0Zyu7AbXvrul+mhQ1vYdaHHuQ+xJm7K+R81cnss/YRJFqMzq51Pqr
ZK1F7p2vltA564whbv6cPl1B+9vpB4qDJ7z03+vOn8DrJykWRtrSsPFozMIx+psu
kUd7Qotsezu3tFZpgXRpKjKw9OpZUAIy7EVvSPHNnjVVVGDIasYcVX6PHWcsowBc
t0YyjsGux1qcfftECX+/B/FgiJNy0KFMoTc8Oz1me2w924xUctTTr/2MdSN+3a/z
18XTfA4S8ymcSHDt3H86S79F5su+NsM+0Klz0BlHEYgSwiGbZ5b8TEukljWAcJuo
1grQksBLpKxQovzhMpA0+LhzJA91pPekQxjlzruxMOBRQMaRz/Z+XRSqCgPBXagY
TTmz9+PWlwyiauUi1ldxNxSEyyC4jaXM83Cw8MueTvZ61RSwnSF5w/jHTLinrQzO
aBAqq39gNS+8oW9ffLfTFHlf/t+3JpNiMle14f2U6es8GRuB6JHEYkPrebAyq742
QE+yRrKn2ktofp3NsHrErqGBx86Fwe1eHDxkGpEio3BzteqItzKfQxCJ8jWihRlm
6uj7Ws0pseavD2/3YGcfeliQP481tXdPWCu8pUUalzLVTYcWgTYQsnU1bDXx+NYw
Wbeoz8uisWDmdT0/z7LmjVtNyn62QIrV+eag8Ed4C9GAtKVMEhZNpJ6dPWrrHgai
2IuG9hE1vT5WdEItqkJi8CJUqeVVjw+wMmb5hAuK67cSBz3OqG8Ks2mOwWejgvmm
XazKh2GrtngWPeaP/lZGlCj0BxJGpSelF7SfS6JFQCeVf8NZ+49Ad5su97GFfhJx
6zw8phWd6Hn2AQedOApbgpDij5NQj9EePlCmjLEhHDcRP5unwFC9xQ0TKj8Tt/2x
uPrBD2guMcUF0JidTCIREiu1x9vkAZYUS/7DzmpD//kXWFgVzEO/tcMqUzaAO2Ni
Rq1nOq8yTgJ3WfEjSVVGtH7HAY2dj/ZTQHqLgZLMmzGXG/ALySkNLlH5MBHHKvQD
wS/rsxkjndiNmtpiWD212SjDx8odeXDwhV4Gdw0owxUHBic9WWFYRhEpBEbioYOh
N7xl99uBuWZ8+o7BGjHEsWO6Pp7Ns3AxssGr9h/3fL7EckKf+dAvjfgU8MaOrZNt
hIpuBtZ5Ayj3bkGexWKpyL/OFuS5mPMPh8846HnxXq39jyvkoD5rYHSUYKCZED9U
i07QjmWrjNQ3ixVF1jSsgA/0+75a/K8JWOrOMkmLFYr7uVpRelP2BoMPoGFSKGS5
sK79plcn6AnEfLKAp1o+/brDNsZar+vjawtjK4lPXUN2b4gs/Fx7IfxSTDILm8qH
vWWS02Msl+VzyNC4bhzsqwEaeqmQ+MQP77lXNopLJjBTMahJk/HlVpN6LamBoJiB
Aa2xIh+xXOmozXOKTRFOw1RTFD8PdI5r0AmJZ1AKl+QiraBL3YSCekhS4Hro0cZX
ZjwFA6GFn6NBnR9Ey2aBHuFF9DFeVbPMilMvy9AlNPloIwUV+P92vqQS0DMrQWv9
pzUQJC2Dc6uPsyxsz7H+IBQi2sd/ZheXlMv/yj/9/jJ+w46SV0a8wTvlv3Vj7R8e
/SPURgSMUY8GLDKep6FwPXrDPa/nsA3s+OPIGT93xAlAgjBNef6xTP6zwgcXltxk
qr+Yj0fMyzNmgPtMvYWOA1wSaewvwxO63LAlYGf85crdeY5R2JVUQHMcSDz9UQa+
ZBghKIboVawjojfqZemu9kaGJj3BWk+Sa/Vb8RzTEiti5UZxka90HMYO4VIYWyNv
mbRKPprn8eGYDGc0JkddrMgZT1kUGhVtG+I/oMhy1SaZQQfdC0mnTvrp1kLeCWVS
5RwT7MXYvXCaoVyp9Tg5RFeVGQBylXQ0jfcl8IqNZenG2pfLIeHC+KkcWl7+roUz
qTWwOPjph0vnB9XlcDP9sYsKv9HycEf3GIig43c3x7gbJ2NU6liKmJX82+Fh7JZi
KU2eWHeeDXaVM3/QDMUmSCn4aYwqYfu5/awO+1wFpYrSePtQuclDLoSDYq0zijtV
pfx2wVsMW0/T8q15k6lgDr/Gbp82KOpRcoTU7wX5IPi6Q0UGUyN6gbdlDvILyElX
lYhF+Ff9WvnqlUgoQFBhG6s/fuHhYKmhe2+tEHLcH2sVwKPVS2/Az8Up5o0RGYNd
oZQ7xQcGtdh59w+jGUxzHUhzCHM5rKo1bcAd+Xdl0ook8s4YZkSoBv0Nsl14hUhT
3OsRP/EGQB+LK2Pjm1pmX9DXfVPew0dVcjBdRNyBjDxvbpy3f/F8KsE/XDrRuzlj
J1Smmz3moB0x1GfFVcV4mj9P7KL4Rp/OxkMTIFlQoVv6LYGz9wKM1riV1yJgvclA
cGXweKYLr7eQ890LNV1OYmdPgJllUz9jrcAoASu+o8wZYIPH8PAS/CCp/gb7a+Kb
oBQwiyAm4HFioJqHUFyRK1F42mOeHvo05egSkRjFeT8tQ74K+DS4I3hK3IJcR1RC
PbnNi3/e3hVos1ZxaBcDOCA+cqZQOVUqBuL21eBY9BT44uFj6koCITjjZ0mwZkZV
/n+0kBVcoBRvcDTQmlEyeFcI0rKGbgwVXQxWuQlmrjb7oX+k1jdFtYMdsnPhhjpR
vt2CVfm/uEPjW1aE7XJdFwGkBCG8gVxqhv/NXLKuHQl/8NNpzxNeuj6WGIKDfp37
ngVhQmi2pYCFg/AJXO7TLhvPQ0zZKgb50kkauvnaYcOX56/wVi3BZflUIyr7jX6y
9c2QnUHj0NijRS9L1DhKuU2ywMtmRy3RpjaprTwhLxEk+e3M+5rR+oB6c3+ubEF5
LgG4XBomtM8A2HlpeBdYlLF+tVy1tZGqJyj/RuCmMGfpCN5PUxu9+6gy9h8uV3v5
ndsqnhFLMMjwtCeKNEtX1A+a3prkS1e+kLaQAv/mN8jrfsN2HUxvWH9g32BZPlep
8KT59e33VBmX/xW1ms1+Hs5V8pGsad49kPzH947YKjdP81KCu2t5GgOpBFnuEND6
A0mq4A171G84hkB5ARMZtbiMqiGMsC4Y0EY5VHEeLc5ebPm4m98nd0fn4UE64s+Q
PSRGJ7/aos2gmDLOcNFtHuRye3fHPe0ySvSltlQtryMI8FxSTCFfCW1xToJQJuEV
Byfy+ngqg7PAmx1+KBa2jRhjmNbcSbI+46bBXTE11T3azqcTo7A+zKuFCIT5lJlg
rxstb9kaYOI2P8jeJyZ5k+kNNUizYMVzcnUnwTkuj1+AaIpp2IDmY+OsGly2tS/i
sylaJM/7O1tHSQA9gC+Y/bZCI3P0NKPii4oFYwHpiSV6uJTbmeOa53buW3OP9Tkb
nYeKZWh7j2q10ifmc7xefhZeqf/hEkNZzPpt9fFTBWCBLaO52R1NqCoqn0NHHtPY
zvdrGVAikIJyP9D404M3BpQFz1IlRWHI1kp5ydfNlBbiGM39U348pVYwO+EQgFhO
8UPEb9lyK65EC7v3Jpy0MOWfbGYo0Sys864JfwZl0e8JfiILmpnzSUblK2HwlhdJ
ZSBSkKphfM++uGEnjwvsmxS653rwa5V5Y+2jFq/CiF4JL9/h/VO/sDjKrbPYfO7t
ZgaOS1+TGfOFK563c5Tu2S3edQQztc238h7Nz7bfp1ozzmCpivgvqtD9UV+/MPmV
qL2BNt4xXF6lgXwVKsVhaaOB1hFi+Ld4pvXv3W5jG80vSCkd85G/inis9DOoOz3n
aFnaIMAlsol6HTYrknGTRSnYMWMJd3jTOZNdkYNcZSJrKmnV7FxC+py+lQS84rH8
uiQS6dPJmSuKwL3F+R9xVvVsletqg4/7pI91PhGcNqsLVKxRrQHVKynmxe2kTbY1
L411bhwy6k5BPgpuRmvdYu8wQ5Grs8upClPCvmP0772foIFkMBAsVYjBVdPtu+5A
ae9LWm1q1GkPjclEz115SCJKCVlCgLHy50WTn05Qnx7nSJEyg3cd2m+6BlXMuSZD
0IwPTzewV9gZxR44x10TneygELn3d0Sdv2y2vEk7UpN39TCDMj31TRuqh/PB2Ali
nCz4j+EwG6F9qxfobTtG4VyYLIDtTYCJ3JKzDs9E5kUh0nfk/A/O05TzmRr4y6Np
NLHxMbYswph++zssZQIexYbabxjuduIV/8T9yD6CtHmSi1usfWLBzzRLRDknYLJ2
lqdDkyFbPH/siWYdE875QFWa3oG0fBAt62OowKEKc7l+szWzgxLXpbjpK/cp0Lb9
CzGFYhAiR3u0wfGDKiVPO4NtLXZsmT8g1hw4IhWkn5rxSZoDZSqLInn5SEtMa/ZJ
mz0fN3YD0ygowGHAhVPmARYXv1/AENH3NeXeJEB7SxzD9qJsx5cAgZmjD4A+DFg+
THW2cOjVppbymICmzRJL4i6iFhWOI/ZMSEvuolEnawCi9Z9MN3iHHv2NOTg9B0eW
K4iDpyptNoaAqVQOGlf3FkUifH0faBrOdyRQyTM+gmiLcHcpG17tAW5y92gM4NYB
371Bca75XWDnk/UqBDEWU3p3gWXDGRAhEB+R+BKP/ZwVpCpCbg0yakMABQCW2EFi
ZN1SL0X9CdbxK5HgL9YzYd1UF0yzfElzasFs1LGFV6MZ2Z557b+62RCGuD5ZSdhZ
3mLX6OrzNkfKFiBHwUEN9ete3HF/E2T0f9jKNWjSX+cfwYolJ59zmLW95eexWQln
3b3E9DxEM1RwGaq7NnSGqzPDMu9kt0TwinKrOxVk8+iWWrZLpYDlk1coY4STpStP
bcVaEosVR0s4MhQYhylQZT3hXxcZhc2dfp09SWT93kicZXiYrHDNl90VX5oT+XWK
DEzhM9RVj3hX+lkuIzOonltYc7c7sMku9eM908e6bTNviTwGrl7LFhhRNy0LcNdi
Qeajcuf+ZMXdEcxmQhaPZDvbSV9jo51U5SSanhqwrkVwCAN0iMiqO4nkGzz7r4L5
GA2pR1NFM0okik1I6k7AFTRF2cWUqaNPjVoRdXAUtuPSA41YW9TOG17EaACYkJ6s
7qqHZSebueYqSGFb1/XLE9JOHcQKhPlxm5TxEE2+SYfum+h7AJK/y3MsThjt2+7F
x3N10u6VcaQ8VxMKwhRG8tAsv1VaYwsL6j+PDYHLdmqv6PufMLt+43VL0RrJTHGU
/WzLHHfYfvC8x9zT51wFB/AgwPIhCJq6EnSZXGi1n5OqEr+i7AmBUi4QbDJEiLXZ
2JNldwaU0mB8SGR9J8HHqg70VOW9MP0Y8A/MmTgRHLhvBbqH74U9Dt6NkXpyrCTF
tkbzEOvE+al6E7ekE46J8v63X6pMT9uBR7XKWK1weDWjuLp+XUXC07Vi6hrrNbkn
bSX0n9AIO20JkoeBAVn7vy1ArmA7sYV1xIJ52IfRmfwDwrt3cw72NOpXk/2hSxQA
FNoDZd10GuUda1OgdK1Lr9BCHYWm5a2esvzom6Vke+vrNYXu7I3lpumX8V7zZOvF
7FyEdW4oOtDxwiVlVpAQD3db7cgDBKhZclMQ1j1eqfjuBoiyB9YWRMBZdcps6qVv
S73lRGwtQOppCoIQ7HdjX4W0+hkPjT1Tw5KOFl970Km6vE+F7hq5LKrOUys+3P/U
yvtnvDdktLZGlfmhyvIJc6iinTmsNNe0PhFFhqQR7jq68oDD8BvZWOo4R/OCNik1
P/6vPNOb3/snCFud7rGrkGIexOO4fzUiwE1NEur8jdgwtkG7JvMr34TjTYNQE1t1
ipk23tCSrkHWJo69JARHZN6j/28uSKdx0r3h4QhdUpNVODZduUBsJUHIRMHk2Pw9
7KJO/5L/wLLA58k9rfocbmEoTcczaJEvfSbY0ioz2HDolmpW+2fpeJyNtbIhxSoa
zQTL+NITYjat7vTH6WqvMFqjYszMPvYjeoY7sF/kcHM/lOgoqVinLjGhxFp/5kUT
6tpohGsc1tW82d2Bpq5nr9R28WU/+DgzeQJkf+x/ohVFgrGFw3BD8kvaBXuAX538
R368fQfp0VsbfaF3xlXevp4N4e7x48NBsMLJcWI1zy1IyqsTy5mDKpq8GxC40Puz
z7/k1h/uw/XsPLSSxaP+WrGEJXGUxx8bQiEtMlvLdkSfzZORBOyVZYIUJvJmF+MT
lpmjMlW/wZujQHe4HRECbTqoO+1dhX2H1C9VPiZUxCEkX88gmBnZsYyL68gkiqGK
B7j8OrInW5IgE28uCAU9h65W/Ss3MWtQc2EbcypgfTsSEkFqthi+Sl6keWHJx0ha
pMt3S4fAV76NadRr23q6En+DfRqbJCxmiYhAZJsHM3yTjFvwiq1pGGyw/a5j6nBJ
wKEmVUdgPbwLGbmyEF6iC7C/MealBHlvWbSeVZHn8XlAJ0ytW4yAJzMxl3GpkfpD
lBw0YKMkRbqedwscQawddgN4N8noIMMYNACN1WbrsPvsfGoVb2mvkK9dROAwTSoD
FdrrBf1AgfdSlVFySc7dvclg6vcTFKa7Xdfqj/gvv7tzhHiKIMrqlfrpT30c8ggM
a8Z5z3G6T+avlfxd6amtcZVGfXdHEhOZBkNcjjM98GAbVPklRYmLE0DHmi9Y49ty
P64f/It0g/SNE+Jefs8W7ZSMjyvpmA0Whzfj2kNlsywkUkMb3ffmotfr9jsCYjqx
J4QsXqn//fgREj8rfAs5NpsDXZIwEMyci3ko+kl1wzE3UyP4mXuJRS/TmTliNk2h
o67v6prTvAn/s/jIa/XG1SDX1ME4QBzpxtepbi+9mpe6qek8Uxcdedf9OaWGyS16
9867SMRg+j9Tpk99iR54+cVU6Gp4/E7qNF04OfmQZs3cwVhhN5Xz5mn2pIcmRJnB
1t/Jo2HL3Ilsim7eFx6ItrHG3o7rA1Pmp/8OBKEP5CgkpCHRitboONh7NK15JOo1
nYCnRamWuagwUL6rbMC5nhFQ4e55VRjQonU3KBda+M5LLCHVjc+/USslQZUCMChf
E4ht5zU3k3hP4T2TTMzHJnypn8fg1AJQuBU9GhWOXWZpf8/EIU/Ud8uTi3ktP/H1
GJTdaA9LWkFoJzQ6W3u6JzehzsNJ34npE0CvIgo3IcjJj0CGubDhdonrMvpJSjyq
ydmLFdxHNZywx6EQWgURNNRQlPVunriaoH4CbnspA6sKXPZj6Q87NDCudSAbP0Sy
4P5EjPv7HSatFyfjYOeMIVYo+lY13+GulHMP0mafFBeyjulz61NnS2Iufsa3phsw
ilnp8rcEW7ZRc4dC13VMIa/sEPrhS6RenQgC55MnO70k3eoy4zaU2ZGMju9GDuIp
CVhkFO3xAWbO0Oq7LzDDZI4CuFseUOGAk/i2vWjh38sy8mjLZTRp6YrvsweAfvPg
8SBUNpIORT9nu9dowSRU1f+loGPjtxJbDnliwvCgJfcFOHAtThN1QewYKXFi/SoN
oqluojb/41jD2UgEv9LXmoAxBj3rHiS+cmiOnnmRNHcjtsL3C7JIDThd2cAHTLjp
yBFx6KQpeMz6Uf9qnakcv9PITwKxUanUiOIxpaoNbq1wCGTuaQxnJQXTnpxfP02G
mzHThz4gZAXI8dp4AAEM8NaFuZO90MtfLA0cr5GGGJa3mXHR80rjwvgwS76TaXAn
pT8OCE08Fek+BS8oJiCnpE2ol6X6HQKPSdsJYwBsjtj7dbhSkaFoIoUYGAQexrd4
IMeWeLafU7+v9Vfhf9kRYiqccGh820z4dY5wQnMn+bddmfCmE3cO1w3J8BgVgyPW
D+ewy9+pknX2RXuV4WF8LPoDOv/GX0ODbZkh2kSUkMEeJrAfh9OY+kKVEZjK08PG
ro4w+i2p2GoWzgQ3CvPreT3B/UN9bHdxCFMkoiFGDP1zPcZxSBz/KDA4fEKpwz9u
NFkOrre/dFu1BK2d5ISaH6revfVZqoRZPSLOwUv9gNf1+XI7jukiSSE64T2hyUwF
jzGFxBZCh+M+oGkqYYbfUg38bbpBNrQ47HFtqCdcvh3Zevp6iEvuQw/gx3Afek7h
DdxgCSDIcg7bwwjRGMAHNH2xEXp/3v9Ifw1WD0gE+x5BBgCVQFYZxYUg4/yEoV+z
YsuHkD0iAhSV7g8Cpr1ZF6UH6ywp3VgATAj0Ix+Vo7K+jsPy0EUUHc1WaKsM7yLA
cMxQSsbJbRuJmyw1t0KtKPrVo/8FDYZgX7eqRIuMBVGW62w8l9PTPFOUrI2BB9Hr
ojUKeEazDbwjuaU32fj7Fs841IS4zcj3LGBhNurDQWFKV56451vxRtyvMfUXDdTV
BgJFJA4aYqUzxQJo50pg7+7SEFfIebZFD97mYHlHg51UXsB7IBW59Rnce3RpDqaZ
TN/0Atd8Z+joQkcenvdfqxmgEHfmAN7ZLW97WtzO6NaSS9UHXezM10DHSzXZX+pY
tFha+CRCg/fSC78cZvbExwifg1W5jst5+WUf6sbyYS2S17XS7n8NoYAuS3cVRmLp
RpV606abqZZKb8k+ABiBdMBHHc1/FBGy+7V1G8T1jeya3VSRGQEClrUn5ESeJOx4
OeZjgI+vtaysAHG1Nqz2TkKXa8R69MNiloNyA+p/Je0rSHwV3ULBS3/LDv23oelJ
Up3XZrbLPZW2eF89hvxFqV0FgNoQLlcFwvIglLFp6Y8L0sGXsK2T5cYTHheiv1S1
Myt6mexVlcIClKVlprOCMuv7WetXMBf4w612f0sCoEuhjpKutXVMcnhpGWI2XF0T
+ycmn5wTku92BFrTRDL9G5wHmwZq7jcrvndfB03G6tlLR33nw2fVxThDsrzBEjpL
tbDviEfc7iXfzrg8usLAcmnLnXJvMKTUv0cVJhxVBlEuCVy/PFFr+whjuVU6WMy4
un1IUVFfoi8P4tjskYYAL+7eb952zJuJBLQg4LAYbjtyDC0+pHAG27c4PEDZ//wg
c+g0wwsHvBBrGFEJ+Uur+vW26htPTgO+aRfBRkDb/ApdpN9E6bF6iy1WzZRfHzpi
23hiLSTbRfjsMlWExbuPpiPckat5pdGQt+Oj2F45WEAK8MNxQlMIM+TMIP5VE53N
FHD1TCSqeF6jQ+5K5d3KQYtuMnuyZUVyOTusbV1l3NJYr3meT9Oix9imZmelA/5c
8bY5Haq+mJp0rRmPgibvIDkcfvGpD+WbJTRBwezrvcbLhaI2rsmA3P4NNIpWj2mS
vqetjkeOYBl8SbkEdKUAfrXump0iT29SMzL8OcVkf9tTUBbjUO6SKoyuitkpktLV
1GRTfGpyR3lJnC78XL7HhDSek7CucYHEve83JIAKnPODDcy3zwx2EdgTPIHWNPkN
E3av1YDbtPy26uCS7ddqsDuLnye+4g8auuOiBvvEYlJAeLwJ1AX6QaAjfJwe5Hdn
hiIXXn9rUxlqyrS40yk4nQL7ZlcLb+lr+VCy6S1cC39tgrpG+9qlgAx7VPc/Ph4r
0lyjUAcfFUMMbUL1ci/MyRftuIUWA47M1PQ+hPcTzMBsIQBjpRVNyBle+SXK/ca/
EJYairj5gf73mpN9teulbm8xRrpsZsfTdVPQ1Y5wVBQg/1q4Wny3aeoZH1q9FiQZ
nWJ8s5teEJ/7HQ7kl6geru8MDr935b7nnfIDwk7eC6LdiGsSrpO1INn+qHweiKkt
+TeldFLHRH7HMdTVoOmQGJOtBZi1xPXcjSVW0GAmSJ/N9j+RiPYZXvP+orEruxqm
LBxphjX8eahXIFA3lbwEIfPLCWOEKv3ugww8/mW+XvU/9u3xKFTGxFg4lwYYHAJY
0HK0QKkmHpc3p10b7Ky0HwyQ89wNuhLqTjRf4lpiDsbw4JnMJhos3AO5KMqAsrXo
ZJRFtBowR7p5ftjcl20TCirrCozGFnkcm4McPfLNaxOrvh9H6z9ibEWnMmK9sFcK
CdBTO2Dvrrafzx1Lcxy2PLSbydQAE5SHyzS4PCxHraXZIFG/pU65mljrzEwrMHPB
dIAVAPnMHPyXLW1dRa44VyD6e/CYv4A/rzCiIHyKApw7q+ZL0qyi+qfMzuBl9Zxe
MzLpzUpGOZbKqpMjLpjz5woUt7phROW0Z1pC21MbqDsDuGsC+Rj7/8cD2HSrEO5X
738aZLt4/YJPPcUygCQI9atXZ/w3AC96MbTjBmgkjVQgHzNk3nHwpCgE//UneXP+
sZ8TZE9d8ZFOIZPBvTC4N0hPv7Z81HkTP1IPc7pQtRz5GkJRV1JFmfP6CcfCjH2J
HVV0lqWBiPAOUlHw64TMX2ue4yJp4RO7EljSZKgUiwcoeBLUZYa2GNPLTWTqLf5e
lQ/Ofv1AQQUJ6jdNVrFNqmosAxxHq/gS2ye/xszKIHJfHeuR8K4cb1gEdlUS92WW
59tBVfKKo/a1aT43uHhJVwMlfiUp4Xt0uMfDw+r8onj3jqK9y3TY83fzYft7OnaK
r4KbhdNvQ22SCtvzXRcuEM9cRBShweAYudm3RBFJX9aNUaVB0Wt+mkkTd89/fYDQ
4oEyQMdXapqUbpQWXuvItZaW1ltKyrD5p4pW6Q6oBA9FYfSjYdzbVogYj1gVKzyS
6FTzzNn9kUZU/PONnmoogG2aqnNA8UMu6TTV74+BZtnX5jeWe9hMq+hh4/iUrMcE
pTQ2SIGPrLaCYsF1HYj0huZkQG+Vgtg3hKGzzsx2RxB9t5IpIn++B1zhpUlnxM9u
fhZVUzLsKxeOSTz36+A982aX7EKzg/VscfGeW+B696HWyQM9at2lI6PrwhXeEWff
VfI2AUhoCMIo01GunLydzbLzQbksXYUac30KLEp30GeewINczsFsVCK10pXL69vB
RJko0d9OsZiE87MIlARgLuRwGQAP/MvVr/r0iBey9+DCcewMKYAk+f/esIgpkLVt
/HN2PutLCP/Psjmi1H/1pL5vfJ9hYd72EKjKQN/aYczHantKQcfZDC5GgZgZdrXp
tFfwECMa2SEo2RR9kAIyGfkUtuzKoOFHcrzapwPP7TrY/ooNGLXqYHIU1nqP/6Aw
iHC+IlY9G2+dwsb7pWXCf7oegz4+AftJSmjz0Y/cKUuN38gZ3rz0aipWk35UMJo7
gF2ceHF4CBlau+O8S5O2GpEfzQdaCe1DV9tUuL6byzDss70d8yH8/1sCwQJ5wymc
oYV2BM/yY1Pra9o/2msw/xWppxOBXYxNxUC8tflKyIpS4kIFMgIW30lK43qom2ew
5HxCrZVvSRDHMmEa6WBn5syM2JPNeJut8DxBmTkXCXIsLJ6x509dp1uqROixqdf6
c6gEBTHVfU9v7uTh51Mq2ZD15NdiA6zAQSay+zjtdY9jNzniftIN+uqn5YnCCDrQ
r8yNyHEC/t9DK9PD+WgQoWdCR7Xr0cckzEQQVfFdn3ZAnN0rfgyfnPCEIL06csEu
s8yuxer0QNlZ2dnSu5+emNpcyzh9yKLU6n7e3ly1NoreuYv0puEvhE66q0EVjSqF
E8gVlT20gsjJoBlqyRWNV7EoGkSia6suWykshQ9T28IOEjBUdzjL4b4gFSLXJjPy
a4Yi3yjm7HnusA+Pu9tbOjWY/7XB4HZr1kPhs4UV6ZvPsxatMc3EculQCgKjqtwW
3hSbdQhJVZ0Hq+R0DHnExGhC53hGra4UiQZ1OQkklyDx96d3qIMqr4kNJ9DyT4ea
6z/aytFogUN/nUx+aA5tNEEKa/rZpXBnJSaRN+mGpclw8XTMpAc71RopSlLPdtK2
MnRhl6rvg7butf9VHqxZkFrhUhXLoGdn1HdL8P6qhpBJFDn6vPnxEYQZ40YpPW40
lpi+X4je7ZjzvWfVx6AjIqnRd++3ubHNGKLi/MAQWzS99eTrLb46afu9IloxCSTW
iRXaO4v1dFe7PFlaVM562hvzB2QWvnSqX6hr17NQNFreVH6fD0xLxT+TFg8l5k9D
dbKdEbEOPEeFXlPAtTm405UbjZz49cHgpa9iNP+Xyx4jikdK+Uai2k8z4irDwMX+
K2QnNDna3KtMNwyp7sDAgiWqzkWnvU1KCO/llv25Bivr0WFbFusv23YP+JTtvN5X
k3lOEVZSEbfg0M8j1T69YL094kKUdUIPoiJ29+WWLoJ19YwFV9JK/dlRfA2DQ+Xy
rloB3uNXehqGB7xQxPsrG2gspuAKKI/Q8DPBT467fuq/H6qOn+cfGkmdeR0Slj5m
hsgRRK7Mnr0VaIoIZlFMtUWqicqPq+7u1xgygH83DJZ2vaBGQzYZKhZOuikG6EUE
Of9blh3Xl+vnJf7IzBtNbCdJNq+u0ejkkrQZEWAVA0LDi7zazjx8nlE9os4NyPZN
tp5VaQyozZdsKu9R/7Pqw9wDlcpdF1yD1egvnZJ1kylkQmyewtNS+jBymEszGM6R
bibFV7gLO6SYlTDvTi6vo1T3psN7dZLjcWP76UHZ6ty69zu15dMu5HzAPaOGApOX
KxIX4IesxWTQBcApgK4f4ck3plClOoUVXsOv0P4nTvddMvKaA6KC/owVMzTg/lhe
mX2A/F7McC2evTps+44uBJZ8huO2QXhJgB6pBwdRFKDts5AmFDJ9emEoZQfd+Ku+
5zHGFTRzqxdVHmFaQ014fl/irULcahR+6W7oaBEeHKGWZkXyPsLuE9tIQ5XRJv8x
Kna3ht0T+lmflSBi5ynAg8bsVaR+Y7k7jshsRktMMvpccT/OzaRS8aNUC5kzkYle
aFlBNDuaEbaljsncaw6BI6Prs1BlgAioP6ZXqLulUfP6jkrEywdv96NBrCECRIQ3
TAjRy0SszDo2VEpFUZ30Dg76B6DjgweZQ7Ma16hArweFaORbZr5ySiMD5Yc3EjqM
lwbhKA5pBXTVK+EcSg3lC4rEYaSJqWy6U0erMfC9z8iqmUSwCXg9PPfNFId70vM7
nO0ySfyq9t65Mv5yzDLIqpYtCBw6fHgsvNZkqvpza6ZbaSB1egR8PVMgSUn/58QL
IwiVn6J00YCroWYA8GXVJoyF4Xncdg5v1SxF62k3nt5nHUnNpJGpixbWBPvBhvPL
K1BJqhe83gMfhcoVTSpKmWRk1+Tpa9tzmqIrqufi6krDsZqj0Lglv3wJkV58ZK8q
85FlvIwSYmrIRwnA7NM2uoW0Jz2dBIFPIQA7w+epJ0Vx3LE8/bpzoDtxC+kGeX+1
XgdZsoVUlz3bqYs7JVIWK0Hi43CnxvqpFew6Y61re1iQzsKqE8ZuxZwBEQik6Rlq
E68oUYFMUpnlNj2VBFJIsvJoY7PO6yRVr26PAhBYs8rGVSKcuLH5erMQGWzfL7vf
d5/TDQCPAwfHre89PpLUnKmkhzu8dbXRLWMnHQSjhoCblPPRW610jqtmLhlUSs9H
y6r3HY55n5tVt/KEAjvKn9llz+iSm7wL5juRotlBpAHs54BS9mi44fhDnhfwarTm
NtFfKDTBi9tM+TLXKJZi8kHlGbta/Dru+LzvWoGs4RIBlETZ7D9Iq+XCCAVbJf5E
Spp2FZRi8cYY+hAdvRAHhNmgo7iPu+Gbyoj3qrnMgOJ6OMkw1H0umGwq19EwOIV6
FVCDSbbToh9YUldhJ0MJhKjNxBaMEf295V2BM6a+O03EdcnoFGC/dvkRuaizcnkT
5HfEAgw21S2w2H8kYsA3mG88jQLaI3DYNpexzvxAY7XD2BVopWFhq9oDrhAxUCJL
GNrHJnBdpMiKUIwovccye3ns+R/nl8PC+iMBQL7MFbEMgPHzhZRtQFbtgq2FL8xi
YDdjt5WTWXJv57jyi9yKy7GgaDJP6rVthOeARSTPl1kceyHgsrQ7mmHGrlLIAydq
ZZf7KsTx9n32bfO8aW65FCpynUG/P7ksmIFGlGtiVecfVe4DVe/mmzIzATrzRrgr
L8FHLrMo92uhDCD21BDHdvxp3+cK3bargoLflIB1xfnktni7+mdK9QCRVz2azPIf
UN+K77mgzOtgZKNKkOupF59O6FFpWmUqF7KQDeH0DcZ8DT5Di4BGKS1w+p0IZtHs
JI2jazipnl5NNcd8zFbRrpZ+iXsM59HWqOT0oGdTqsQV5WCAZXZfKwtvFIP0mi5U
aN240fw5uIrMeZqG+QgWvrTjSJwxxmnGDNGpRg0Bsyww1wiS1EO1xf53xIqBU2m+
UJytN2fsI1VWWgpP9Utw547/5T2gRgzVUpcxgxndmV3PjJGZg46NSoMP7qAyAs37
WQXNwG14H6XqeLL8CWdBwONHlE13J0OST8T/8Lrfwcm116sPjE9zJ0UrKWG5Q2xl
BXHcGii8WzoUQpTrCeC2xOBKxdR0HxlLd3YpZY9uWfeGhyCW+VpgVIxD8gUa5EQp
GWBBwfuzdNUP68nVNV74oLJnyAsqPh+srzKuudFL65DHKB0dEhtE3UNPmkVfMKxg
4mWg5ozbp2THvv3dGG4+ptnfwsPZcC4GxM2PFH2CgdHN0FeAItJ8DTXfDOn7L660
LTtd6QURPGHmQz6fyKABzYJRbNsORx09/G0JSIH0kiWl3rHhfGgJTm4omwpFvquq
TPHd+w9XbUhn415FKXmX97+ZQZVdaqye3pfIdmtsaMLiwtBanafUgkJJDgKIxs94
iy9rXNVH5qfJ6Q7REWpqtmexg+DGa/XO6w0WkknBj6GiRvhN7Dy7HyNAzJAZebKf
LoOH/iSJt6kDkSEBHfWUlV5nzlog2186kP8XiOs0oq1PC9VmRFKYAZ38cUj9pnF/
fKljRRvqPs56ysbxJqgN3d4exVN1iGfhnAOerbr1OpSB7tFWabyDYIQ+hrCdPzYV
/NkrinlP+DLLc5+f2gm8/Tv/4cmR2lE/hgsPasZjCIFUSpVYT9SUdkjMC06rBqM3
JRpA0VJ2P/p2M3JT3NHsd7ZVhuKppCWisK+gI+V3Iw9MkVZDStPbOKmcC59cKlMW
4vat3V0frPhZMdeou28aezzJYNOhMT8cQvKDNSpG7JCz4L0vLdOyut2RzUjjzfuU
CkVFR2awWKEL2m9xl2zRyzf3NbOtKvqdWk41EhHI44eUhv73JNBaOSfqavTY2gN2
0vpZfTrXOMMDzAT8VC8oy1RyWAddg7mrdCpzsKxROyPvH3zglbHcwscCckCtv8pw
JmtpHQrg9Q0kvU6NVMKRkcH6JuSZ04N2Xg8N8hLtBxdU/QfJCW7xvSUk58klpf+H
oiPu72Yw26ksEUhw5dOfC18LIX/wlS1xntqH/+9mYlYWxvF0IDOAnHtq6QodrbtG
5EpmUCXyUk0tFtqzASWwPc1rFLgTXu321bVJ70gqpzYdrqfZRxQ79gx0ogwDYI5G
kGp5dc9wa0kDYLOud3ZvM+xX3Kic6COntY4+x4uZ9OtnjT68M9MzZ6P+DF6hLYPb
lJLQh6eCRQNM1ND5N4UEVGETN+r1C8jLUYWZkjdjRMrYvxs20PvtoKvloBb/9WyU
AScLZFgUl2D3bDXiDDp5SSoPRV0yMROXKjo+KtmKQ9IZHUHRcK3lBaKq8z7Zz0lL
uJhDOXZiGENXsCKaDE81nNC1SCqNa7X2hTPDntJBChbMpMcnn/x7cGkyBNA46Qr1
F/eapLNCMyf/IX92sw4uPtd/RYSjYujSrlTVQHtnZXPKt6atzX3wTNk0wbBZMWof
ggGYgnqDu9nUGBPtVkd/aLENujdNlg5vp/EqcgmgPp+sqVeahSVkBR+eu90vEwvK
76HNMAzrBJIovzTGeEHaqvBgU54nAY32YnPUBWkXgSdaG3j3grmrRw1iAOy8W2GA
rrQrjtCTH7GF6UwVI5WblzgSUF8anr4gdPOEu8/+2UknU7gtduGRvjbZQoorYjVW
Vr0lYiiZvSklztHE0zP9OEs9DxjmPc8uo7mEK80Wh0RHgEfWOP1H5ua7rwMDCpte
IRK1ksnKgf5gShmSS2FPKZmdt3egy7qkwvchKyZ0Se7rEmrKrHBFIqUIwQHSAqfV
+IpNODr96GuyOIi7aw6kGNyL9hbqE7OccoXHvRWT4nIHlPNZFFBuNSFC/p5ejjq8
7odP2CgEf3wJzBtnkHWcgVi1bZT5W2Ny53vk89y5O3V7CglwarEXFOJ9b0s0V/I3
ICv39JL12qABSdxRXN49N2gw7tRN1sE741gDXXcai35XWocxn5reU8SdSZOVlc4H
A+uLLoS6ySpboNGMDSC3xvVj4FhCGczXeKawNrz3vTorJTodtwD4kWx/xSfHkMWd
cR6EzUfpRKaPWjgDEjMenN+RHuEK0KVWnuiBd8/BwGKMOL4puu3ZmaNpitbT1afr
xuJF6fv/u9FRkOD3TdmyGRpBqEtH7EFr/ckS0+QPtKvJprAvOqInVYJox0qluLFG
Du2CbIhXQQrbuZzkJVvu9A==
`protect END_PROTECTED
