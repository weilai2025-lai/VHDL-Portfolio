`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4M9OY2Tgd0ZFK/UgjDKVUE7optiwFhJb7a5qakUzDAl5LtYFDaUWNiGN/SHBTGd
KhQM9jqPbekkH5nqIM60lfdOGBLS6wHtDads5ldvb2VB3JeCvmr+dZm9ufk1kOeT
0z/dALZ+mKvE+uHHJsqIKradqrXgYCu2m0F1sHth1g6LGN/LrLZOHjW+fbu6TQkF
WhAl7Md3/SF5ZBUdVxWmqAudOvs4UvRIp3mQ1C08h4ebikK7qK4cRK/K6bJ8JzML
/XSZIYRlN9+Ybx9c6lXMBO9kZYKTrJJFTh7uSI+x70dioylWj5ffagAWqSzgFe77
kBDjs+xZYn4FTFCPcO4GoCOJyjCAFeC+S9AOQRTZBCRLJGbAl2f2gTb9/hKmpu5U
+c8iJvAyvJfdbFokc0o4zwiawokJmoW9TOIAfA2KvPRqRwhBlYNrsO4yLaE/Le5c
vdhjZh3qKiE2KzgAvIntCFUbg9bwXMiw1wWj1tXAkkgA6hEEKpubVOO81MJnESn2
Nz7Hj8oy0PYk4ZalYHynzqCeUCU7LWn7wUi2ja7f1/fcjkzqxcQIWmJlRlGQ556g
SjfwMg7iG9TFFk16xvMCSc4zjb0C/xiVBBk5OzcSQrFqVvF9HdlM84BqXuvkquDQ
PInnW7V5Ro5NVAPK57ebRZRNdmzZjsBIdJ26N75d1K/EzROU0owLe+VFugP85qQ1
R/+8EtqgVHyGhNr8o1Nwo4nIpspGHkRQ9Fkm3cOzm5iN3tUYnxps99vMM6fqkvFl
JKFIOQJ7of0Amfp/BrxWB8fq9n5K5I3xKIgQIbEwbwv8SZHSG8Bq63xGRMu+DJQv
A7ToAivt3/y2U4afqv2IMY1S4BA8hgLy3ewYXsgC4aCIInKhKigFN9Mn51pY2AIQ
GkR3zKkRkec2fz2GaZYwE6qzBGwCen+sSL71pZB9GYJt0wPAQ3DdKBa3sMJPEQBl
QVtD9cQcqQYwWstHkeDCvbJ2Ha0Br3l70tEfR6xHBkuTjZhMybMU0YizHlqbk+oO
Aah+hJ6n0C7dXk2kd8ltqbprFtnLaND0SLBnyRSl7uhDP0GeXrYWW1Q3kkSi+ZLM
7dq11aF2cCUDSDSK3UggcJIXmfKapk4nvCv5s/NK24Nt2wHsocwx/ZBhMqNHPRgE
Vy0CyTTrblT9Q8BjUd0uRA4wTFfmilWvmCFnUdgzFnK10elCwv/wDh3wgxNGUCm4
a2soQ6H6cmiZl1XEOh8QfHGUiNXbxBN4zDXd8G+2+22FMvdr2P+xF6ctVsu6TjDB
McuNOcC/bb0WUeec7laXYkbtmMp8FvPOi59kwyYk2wqoLvQzbDZlMJoC/PEij5ol
jEqjCoSL8FMrKBF2K540INanvsk/64XMuuCdoY4Lmkvr6LZA3CGA3jmcqNqAkSST
iARC46upQ7qT30l7tm7Q+K655fJ9XHPDp7BvxhBh4eDamS7plRVsXxGO87l5fhex
jEj7K7ysiXpLDLnNxqHdY2qx+nB1Y+fjQ5nOodcZND5kdbSr1F4Uz+pbKAQRH6op
NiBoMmtvwO1I14aaVyuF8ow43oDcePjz6T5mObD9HXUJPkyKLHMM7YZlM0tS0LNh
WLfoPcqYqPgTBgfYCl3p9VmBPo9pLcU/P1pqHNoNUlJsRCIXm5O0XS2HOZQO3y2X
eIPv+GBMvGOMuFAhpjBG9MRy5OWiT5OvW0b/GPubvsDdoMVx65vVceW3bCaMHE3V
OO50Grj3C4ZoPsglko+lC046BSfNtyUSaijj8riNQYolquqTjh01eljRs0xBsetQ
2nWP+A8Xbagbp1d0M3TCHor2KLXPgKRNcY3IHBNrdjqIQNDScTx4oZJX1FrgbZny
1QQU0U9rdIkjjkLBszraJycXeS8tioiAMRHEcQSqxgtkJMm/elGreqcDuEyR5GBi
Nsel/xTCOn/YaY6LjGZ+J2BCTocYDNxrziaeqDZOiGjlk7LCDWYCZyPheiZqX7Cd
dh33dNZN3Z75oWgcIH39KmS+uSWfPC0xrLskj5H0NQ8iF2eQ6KGI7Fl7qMQh33j5
4q93thKdEOB7PdNTYDTkm8n5wu8W9w+9SvW0jXIrD+th+MUKK7YMxILeJG3Ubtzp
ClXGSelWGbX2lx5SlDm5M/DilLVNHjZ3Hx6V2nlqTpMHwt/he8bF2ePWf4yQX+dv
gSzbYUHnSNrgYLmtA7uVkB78/MDWvso2nWoTCTkavWm+8YeHaID0/zimdtYqktvd
aZj0RmFdc55KaseQsu9SxOppVYMPEiTJygIkhALBQb+0jfjuvgiCLN4ZqsYrcVw2
vsr8w/PPutqRpU4zCFukTPgwatnnaJiX6YEXXSeKSNPJ3Zwr35mrNQ4gCCdO55In
T062AzlUTkc0EFhwClKVYuRyQA3OjT8bnBVqFgV9JhXh9mf9va9EEJa8U3qOtU46
29e6MGdLKUJHi/vN6e1MB7h4Z6ERlknLbkC2iGvc8191OdJfV6Fc0K+4H5HNlg9E
4tXCgVOmWv8N4xynixU8nLaGeSup6AZJsh7+F3imhBDeTis9kOIOjva8hqQUPjHh
7PlDkRG8H9K/ID5J4rtHeGwyp6TagNk1VjwocBLBa8+DmhmlIisZJ3qpdk+QaR5n
hL2mP7/DG/IaIi6toBbU5EitPIREHnEUPzrkeaVmdvSRWC/rLeu6QWBcD5fIW2Wr
wkt8FAg1wNd/rmNPhsAAHGNuQ2Dq0UahJ1htg+lCvUSXhJhMq0rP46BQaKEdSS85
kYcTiKvaBLPWXeKEdzkJFJCdj3HpQRPFxPboiyXy+ve/U3iy3uSxTZjwq7fvLlux
k1lCbTR6KO3olSG288tmXuLRUaJX+MRvYPxLhnIIP1KdtjuVvnQS/KOJFiunyU7H
HmhbSjVsT7F6j/ZP7uYs4sKGfd6UEQDpE5F+YY7OfPvSQ/+mPgg2VfCqMUBPYWxb
4H5H1OsxKDZS9tfiPamHRT8cq/2UOYbJGsOP9ynY50ZDl2ig/HEqJZbrt/j1wD0y
XQOD7oUAy7jHa6c4szA5em6dXPfBbpYHFjaxYCyBAtVyCFIvKhHEO1/7PIMefGAz
Q5vl6rO8wm7KfDQMt2O4JpkNBtjVSePyAW+FcCLpsN2duTEhsdWxZeHC7F5f1iio
f4iu3qPKXxZtgXpVirDwKm/23e5mekkVDvsiErVnqABpVO2V5VYsgJ/CPniAiq6F
cThVuLnkmsPNTpQvT7XNCvUl+J7/iooFGUyXrztWW7xYjezt2oHjSFUiQakwB00z
NfkDCqXujkEXxzctJgOWvUkNiz+WvGQ3CYy4aXzXhm820mop61yARBkj2x64pLxa
arO3plqJ+qkBojtmlO6nfrt+hJe3KSyUgjlRqKMECk6EYVAKxiefLTXWeDqf444S
9gS8EIvERw2AsoWQSAiS4u8a67CXI9aleF6DLIfpoj0pZw13eE2VoPlEsOd9xdCt
1JSXj6ToYJVU9gtyjnzgNPndTYcCl/8+MKOeygd3uRscE/LaHllwIL5HkPsGTuOi
QMCJCLqQLDFpFLehbox7g27Hz6TZ8cLWVs9zy4eeYeWfCSnUAUyr8mKovEgGa+d5
cHuuHRulCKmJsdUFFvgNjscxnpZjEXHIPKkhiwP3XHT9IFf29jiX4CR7DlVbfMjr
JiQ6EM/JmFdncX/3giZA2GZmnFEe9RxO6MOzt6PLFSAC+AkV1p0oZElSSJGZSlgN
4LnkQMxA99eMpBki8EaZazHt8INNOqpCZQYPPWgKX3TUT+62iKp9cNgQbf1OPP1+
BoIca72Dj1bCgLVUfgQ0Pmsq0l5djjao7ZNnF6t/zVRk4m93QbDyl+1XjfbcMlv1
JtMyB/l7J/RPC3aeian/fc8wUyymAyZPHz15gtDpwAkKBDOVcuhveZcn5EK/c62b
tEjJkuKc97X2+SDVarTxm+XlQ7Qnpbu/DUBiXkyXmnz0Hyum9kCw8qU3rHorsgiq
6SPyEzqgrWU/TTktI2FflMtIP+w/e+owCFuHlg6+mPZmjnnrsSAFkeuYVoXKnxcg
7cU2mhSLm1u0lnlmbLPA6y+MHjAKv/4iIiGzM/aPSd6+j9TOdjOEO7PYdXu2+svB
AqA9ZUiReSOQ6cnBakazcXY3g7gBLT4T+9P0p9pmTSrbYsZXUOL88e0e1PC5h6g+
yMp2sCO3AVw5Y5xPFSQjc3feMhuiTQez65MaLWdPsNKTveoIHNFae63yA74ODdxF
0VxsK/MpWuhqQAl+UpPfgHrCXsg0DRUc8ff7J3QS6CF9sab5iiM9X/AakQomSlU3
YboBJVauDyRga/jghkmeyFrZOLbwuKoeuuEIQMYtpYGla1GeXo9YVMf9+yzfnQVe
bGWjUhG0MRfunGJic4lCSx3DVu6NcYZuLC1Y2wm5C8daxihE0vpa+tB6njavN6IJ
WEtoNA2mXijmz18RmWDbRTstkpzL+RrYQ6YPZcC+sA+1D0bvJf9nEqEOYHqfi6gu
vT1IDsF8eamu/FfYgENT6Wm57rnE5Ci5V5DDKz19Xm0fK4OcTa/J0vaRJ/PiE120
9VHHyqJGBkv6aGlmNn+8Z2GGmqJK3/hZo2XH6cpcWMBq3AmMzOC7gr/iV97rvaCW
Y0jTZcuW63glwnSHMm+wi+FwfmbejxyXaAYHpInY6okKXGTlU0N5FR2X6D3XMDIB
EHqgdtv9vrZmjPAgiC+BZ/bJaWWHJYBD9qDSOea/zRik86Akpe05SE5QXE6kNjMn
Q1UNgqVcSEtAr7xJuFbNgpAzPYnprYiHSP0cnIW/6PZW8gQ0BiQXeoGExuGan2PN
knB606WIyqEtBBIbJqobgrKO8X1Q3nBYgtYEu7CTOfPoEkuon/E20a6x+pI7/w0U
lRgBS9V/Z41h82WpF33dDbZI2Lec8Hp5xE5JpGkmbEAMJSOrCLP5v1rVoUIpljsz
g1vrmJNr68Yw/3+qSZurViUTVsXeGEhvLV4xEFZZ8SG2n7xNqe3GrkF9ySrEmZqD
t3glcVpXjeUXAaFQGN+kgWWBRq/C3SIjhdtQweErDTKRVmC3qbMIZ01hv1/Nzfvs
5YOBpoY+7LM4h7qVbQVwRUZRJcmj7fYhakht+72Q5SmYtt/BwyFcMjg18WXUniO0
nwofVE9tZ2UiMZFGXysUoZcgtNHOKxWj0f540FkDl6AcFagh403pGzOuGQK/dZaI
ctJW4RtGAZ1RQKbyV3ucsSTdf1+PxrdOvFL1nO0ghntdWvPpEnkdjeN271ib6HVP
WLk87XAgNBfmw67FlQnfvm4BvqXRtseW65WyzCYH0toOuW+X3eH0h4mgHph70ifh
vCUePup1q//pAavU3TDGo5ijaYywdXOlqILtUMQbTrSoR/kCTxAWnKdcx7tYzjUm
e1F8Thhy63cxkPTlN+4ZA25OItn6yhufUU5HjSWyYDIQhOIR/yTynYfOUdAtfw3x
5lb1GoM3kONke/mm7BmlTkntA8CMByt1cHoAzSLwir34Mj9YF6IuSQd2hgQyL6XA
5MH5voVTIz/QPzlOIAaW571/02BqDlzoOXTdJCFULCXEeLX4Ogb8AhxTnzFEWgma
XNr8/u8DaslmBF2yBW8Q73G9HLKSTxD3FP2Bi3jE3mNhK2fTYwxZsGO6nrIFEnhp
/KfT2LQ2ePFMZj6fS3e3bA2WUDHO400V0MgY0Ewww114bzcntV7sNbPJ/NkVgC09
3x6WzQn6V/rnELVTkd0riXzBebeZC/mFoOoaK82qji1raDzCSKpWlhNufwiWesOK
lNlGc7c0QAqe1hyxNO9J8zKPhrl0DgceWMbws2J6ud3kLk5v4KKN6XsC3JdlH8Bt
XWndeg+GnqGcyq4LB59dt7BCFMTnTF3zM8/Y5ZPLWA8zx10ZiGz9kEIeFR18Jahn
Wu1m/jwbPI74pmvGdnz4VInfltrXocKghKWfpkw+AayNo8zBrjsT6aLS+8U9g40Z
cBhxR0z+se2vUoCOBNNSfTa713eRJ+mqLwmtAJ6E5iZe98QGb4s0iApKhz/1PJ85
ZDp6+pvuBGQE4nY4AWUxbKZrA4rEbdfi7KDltbS7S9Jxx+tSJZGdmHFm1D3C7fOO
alf7KoL8i2hcoNWdJ5sLuNoKhdkrGmy4cOCyDoETb2d99aw0ipUeZo8tuHIII4WZ
skQymd+SK5+zo2gI73NMJvQrLpdZtBGX+VM+fttAr8NpjNuBMdHMTyye3rMRrYTd
3O4abnwKezO3xsy/rrMBeFGefyiQb3Le4t5qYJI3fPC4PCkv3sv+MD7Uc1jlFlGp
RhOjviQhmtGbrSW78bQ5EVbRjvFesjRzKrdaYOwL0/dpzvx9XRbL+wZAMSi4hsq9
kmJ1GpP69/ZtIYAoJjJFcyJqQqJa6kKbGAjzsHCQ5eWheL7pz5rbv/cJXJAuWFkE
pLRIkH/lbMRDpKhMbRVRhqWgrVqivluQ2ZNGDVOU0az6c/qCZ5HSnkKXcYDqmfVB
G/FkDCYNVWNru5gQ1x7zc3mbTyvjmVHA8RrqWh8bR4drORWwxU+zYPYvseNKUXrA
gz+hlHcuriOrS4WtVUebHdulog/rCh9fZVajZLwdesE+NhsBsKbpfdBq68xpCQ8E
z6dcqrB5Qatkk5jvLW5XNHpxoTMzFvVflmNGeW8PjwLyqzdny/SEVw8c64Ntu9ez
j1o5V/SFIHCt+WfWaulgqs7pD5mdYONp9Ox72Ms9ABldZOiX3GpxmjutpHga/0u8
11TOF077mNYCOztYK8KXEkudN8IpEcGt2+CzHIIkLV44xvKm3Cnjfi53XC3ITFJ1
tIUhDaUxDUBaN/HwEhgn4YEXOWRobxDSLfy8haaT0pzIJfI303dcWU1rEGAtZ+g1
ON/41KjcLJhHtKgKYPGnlWeTZ/QTluTR7akV9+WedKmpQrAQsJJLekNSbsYOiWTL
FA+gOsVaxAmDwNBtdYjIDg0+AEo9QtWoqzyufDJSNwLc9c/22ZDYPANshjAf7f2d
8G85tNi2qy0P0nKBu/aogTcpphr9JZZcSLVE+g+mxPjvqiRZ0RuJOr2r3ypXDh23
J9hIBgEq61gYxXWOfuLqo6u+tow9lMyayl0XSCndpuwqvQ2hrmrh6+taqCMrOl98
9tsr8jWfvG9rZSxiBDT5XoX0edRCBSoKGaBH9Eul+7WeIWWBuuLYa5Hj2JPhj7Mx
zlkdHLajxFffJ6lfCzdm11jcf8ZB4bydGmgDYxcnRCMc1dalN08z8Smuo3xV6MQ9
kVEcfXkJwJ+Ed2i526r+yPxvwsE0jV89r4oIf3eRmy2wT1Ukh+MdEsglxRvU3k/G
YKFOOs5O4Uetfda4YJJXG5OROg0fpVA4+Lomn0HS+LcRM/E1Tc3T1TwVqi0PoxIe
I7g6IIEOHGNNITr5OlSZPN6Iwq587YdXu/CwEB5DOwyWmpD0AGC81GWsgRwhNXDI
1TvOKHHhvjWEYdDuX0xkRGEhqlICp9ohYStzxBs5JqW3oX/7smosoO2a0oq1jUFb
21Nf7OfQfoaGCxgiveb2ZDQGaDc7xSqRCWzazidwhquYSv8BpkT/PTOA3pv24jcQ
DbCle702Vo4yS7B1xx5Lrl11jIwtkujpHk95nK0KVfG5ptDR0xbNmcm4Dg+TlPyH
UPllHUDvRCPo2DxJIyDs+a5/uK5ojd/rpBeEl4jAQrTtpBlL4GRf5JAPVgHga/93
w6KCEJAfzd0zPMxag2KtMzkPgnyXJXkOP7PWrxCrgc01OjooJzafM59TXMRJdD0N
OvCutCVXRoSnyD5bRSO1yTaMZ8/VFX8rOl6iZVX+2A/gRQg0Pca8e6mbuIK5aLnQ
T8DLCIVgDBkGI4StOrzkx1mR41W/zhy6t5dkmCcEkeIjuobW9vDG9yUxV8hVEMWL
Mr5gMwO4dUigzvj0aZWaoc7GHuzjmBApaznIUhiypSLG/sA7Afx3QkKqd4xuPusE
Rsiud1fnHlLvoyAKV52PokggC0N/Fh5VPRSxFmAQIjlq3tRK15dvgdSQV0+G1xhY
wtcy8DizZjSpGeBjCZuza+aa/UCICvHlntcXr+eBWfVthrpY9zNhxryd5HPJnDku
ivOBFFTb0s5Cs70AGuEiudvVS+v/FsClphSeG60YREgCtrCpmt0QS4Pg0+/wZInX
f30DXn+D4ilUWeBQkJOAjzGuCr0wgQrP1qSojXKNds4yPSy/vYsgVPgzZIIT5Tfk
yFjEQ8MyfMYYvZuLKFESurCSwu7SD4mB2EznQ72f0glauFeNXp3u27b1V/e7KrLN
kY2UdjDSDEl+gANugkcchF0Jt7Ge1RWSfvKDh0UW48PtNd2sRbYIkXW23usSg0Ic
44MMW4BsjGj6AJezGa1Vascv/9/N80PiJxgpq5L8UEDdZEFibqEZoORJIe5D3R3L
eo4yHvhk3KkD/3JDBWmH/qCP8PVjz18aSpi1peh9px9Y/4wqlz5OknRZKlHkmN4u
xGqoVmJazfBj1zjV5X8Xk5frlyKsidIwnjZWZEHZlJg4w+0HbYBkefUzQkHFTajB
5pU6i5mjOePIP4pksqTa6X1RUOHNqiME/N6QdaW0hK6TxsaUbRe+zAbMBRej/jJj
TIDWIBXcLpx4QoRQg0ZQa1AOg8fkE+gcHO4snK77tVrjZN9Twj38CYRPoHUWzGlg
ePrL+BJLHN5vDxlnbZC8o5tVRlNbE29fbgDlMTro416PPZZOgsrhz5dWLplOfz2P
t9AB3twU5OZFuWIO/CiWjDSFQ4jX0+/3mdFyO4bdJi3A0v9o5hVJ0ICFkXyozbGP
UNREkPes7xSKhtwlHDSVMTD+/QPk8XnVi57l6hV1m34P3g3UuPE/q3ZQOpOeAeEZ
qdCLGwXGoGuT3OEkusAkDtbMgtWsIhirl0fwupPZtLqRFltpnXKk72JwLhxEmsBP
zOXlKdiiTfsaITi4jFyETIR1+Uuyeb5EFzX5Pii5FhUWJNvtCnHUHAHcV80kfa37
41SsWZtkA2T0DBOuZ744iqy2bIAUksapJBRRjBFCg5bdnwgBdP/FjPgdBLWIbFeA
H6A6Ur4QpCswlEHBFlI3fQp2Bnjf7t7YMsS1NVaPOTIVEmnjxjQbkMJuEmfD2XoV
mpDHlRF5mJODP8SHQ5YqrOc5rIST8lGU1podcOfedd41ZfCoMCbPmjtwVkVJ2Hbx
pLWT33SB2TtyPye50WEL/S2QJ/7EpQPukzyQxFgMxlG5HGcQIKGQ3RjEymYyS+CC
kAJ6Fye8BxlKYiiWupuAxhr9tHizgO313KBTMIZsc3nonBNGG8H27xsPc8Yb3FVr
LqT8BctKA93n6vJog2iTQQJgmi5W+jMyPt1sFFhVOrQKYhFk0X5EDITx99SwNzPX
CRsgXTtsy4qhQO1BKCtu1Ds33jgc+gfZuvxWlLtZR3MZI1+0yIMPHXtpa0kXB8sj
8vv/CLNGchc8BE4zsKic4ZEKYo1FHlLwu5hjpCcacQek8SgoNxMaQnlHQOXK9/O3
i6d7FL1NPubcCTZjhsf1sqzLm+tt4kCIYqAOwplctAuOzcGSdJUYHTXvEECGmPPS
9z56K4roKks9tga0zKk3v2Bj+j6kfDEzEOZpGkqdd7Oe675yIlirejzyO0lWTCxi
S5CJX5kT2PiZbTRiOLbB+U/QqTm2VywXHOenYa1KTG/DZrKPw0IQej8X1nb0H/Vf
d6+fu1QCChAITUSgiZKCZq5AFeWuSqrfhgYPxCIwxqhrmKjRaJ5ugKAHvAlz2A9/
hppv2dkeRXIL1+p/QzlspxpYYe0XsQULem6NWW4KNpgKNAlyjS/6ucpFTdylexuC
fJfPJ99Kq7j+kBx061dbKgnrMq4r7dRlKW5F4yceI5/Oyzv2Gn4nGfIcNbo+zVy/
li1XqeriUDJhda6TasBHHPG/0KSv5Qdu3jEJciBioBs9+sjrudZooTbelGaEoNsi
qDJs/4FKI2jjKfxa6sElColFXDIC38KxAHif1jLCZtOM7F1kiAefR1CzBLivtrmk
kBJq2S0NoxbrVVhOLuzZiJFZMLTLaIuXxatK9nRv1uM4tIccwOCg23avSP/Uqjgt
yjMdhw/N73ctaGzaeArgHcxF4LOO2Z6V1DvmKlgB3NQSMBQYbie56nSDD9AiTvBW
MhBXbNoInG/+3Wqdp2eAKaVZMKRKdULBmkZQlEvXPGQnoy5T0LPJ6t6cyVs/ItP9
gVZG+5APvsyiseNFPj3+Euwah/mHmg5NcL6PbesPlHPNV5w1qaqfUF0BXOFwmMOW
gfdByMAiC0qMdZttnMoWTVWoxXew5I6WRTInRoEDEtQ/OLcn/o84N2kiypvRm/uI
TuQVGp1ksPG2M1E30+7yhe8ZNj+JUmxKg1LDcsa97bILzZxn6pgmrgtAhb3+zwqH
N9+gI9sAvvNRquevP402xGU3rg/SokjlUd4emUBuDajitskXoUTyGvKoz/YCwl8p
c2bqpIwgjThnsqYUfrBdkqMuNEWUgavQuuhg4zgtp+II0F9tYoF5oH8YiPj2KKJa
lVn3FjYOhqWzJK8Mm3EomYjKh1pVk6xRzVQuhmMQa5RLbxYTSu8CLRmPVlnhX0hB
PfH78r1SUpMmkhImcYTu8daeKKKlKPcisTfvLcUqBDmKlzSWYf0qbBplLmhJ7A2Z
C5D+Kxl1xaHv3HFnLxV4w2PJ4TLfV5k13B0xM4ZxrHTsZsk16XG1yN7z6gpQZyqs
EuCcB0mhlY97O3WdBEB6iWtRyl3wa7wBlkuw1ae8LK1vW4xgBAWbj4iYvFy7SCUo
S53/9/9Bb4oFqSnRODMvtIoFPP7F1QzNC5a1J7p3ajEo4n6aSBa+lr3Z2v2/vaH7
sLQVM6oRtUDsFTMzUnGOLg70zK28/JFGupWjN5B7lXBW2YTGO3LaezewaRl8n2YL
WrkT28WRfG6yN1ReRg3oUxqggfXqjLl1vssWGMsl3AqIaGz/QomczxHXgCeisnZA
5M4ouJ2WBeCBtZ79SwUNceaztomwufWpeN+hJwFloHVSWdBZEsvnlRx5L61xB+c3
Ty1Gsffwt7X5gqyeVVFx0uQUSsnwLqCrqqY1mnn18OkxZ+kbeeUVl+z91fokQNpO
BVt1g5A1WJ3OAdYaSq7WzhFDP7KsfG9ytf9kb8fGi9iHvUI/ithA0SDt9VSB49BA
HLjcD7Lk5oXw648VYVUegNEZK8ZWUwp+NkiPejV94t9mwbgP9OtBEHt0SwA3KQmE
t8277wdb75niylKhrVJw1qkeTo5+W1lP1+gC/ySNfLQBZTGFbA/7QvEj6bmmFPgp
pdY6xiKHPn7kn4TluQKDt0Idii/e58L4AOpGkTa450Ruq81A/JIyC2YhoiRaVh3+
CKGnQeHOKx7eOkUcR7v3HjJKc+tPGWkDFb1URuyATAn1iJe2ZUjldMUfWDkFwD/6
zcPTUYaRA0v1XxokrI7LSKnGdwdfNQ7mkhhZYvWtNgTLzIXmyyUJgyutl3QsOoEN
o0pU0A7mGklSCrGAgsaTvw1B/ZXa7/Q83bEsqhs8ec9g1mY6tbEZFvZovjsKgFQv
+ohkgzIXg55L41IsB+6XP5fd/TOJrLWGeREyN64vRoiEf56hYFR81YsdmXaSgL8O
lZAulpD6jZdzsR/JScGhu4Qq6/9EJOp6eMPlDQkvEabO+5wILIlTQUOPmejvWXN/
a1Swya1MVPDhH4YbvKQRiNUkctPHYHs6RQlZx+PTd45wyJh1dw/eWvuLiH05O+aW
5ZI6OFb9NAP9bk2ciOPgLbTJRel+waEtWYod2NbtGBiMG7qokwZbvWwxhKRnfhQw
wWlbYFixJY6yvLDqNLvgcId6SpoAvmQbNCPpElj5JtPAwwWTLeEzgta0d62h/DYZ
y0YyCJqY/RVFKwFrxSGY9E4kfoZyx0MaF6zFES5zCk/tD2zAd/Fqkcyvwi+yGJYv
M3yLm4X05UAOGbzF/2Eri931WfaqNJCYzWG1VsGxtDHIQA6GSZI6UooZkxAnVOZ5
L3WK+HFSr8iH/AmvC7Tl0tIg66/rYNAeAWzLervQrYqqkE1pbgPh3h/ny9IIl2rs
97PAbA6iULR9H9HTLoPxg3LEFICgCtR6I9tKNWN3F5IDWVT6msjxsmxqU86qGzu7
U5KaLLPD+NQ1o+Ss3MX8RFLcN1uts16TbIUo//m/l5aJS+nOTr7J0ziQWIJ0uJn+
jW357CZRnlWbxa2MOtzMEPxqAvN893L5y6tRLh5gzLRe5ILOTm3l5uL2kEZ0hIDo
LlUvg+FpOjFQuuZ2JwSihekXupFUStG623zXFQ+x+0ag0Sc7A4b2tCfg7bAkMagf
UyI13pBG5HuFR1aK9xkzisU9qWwJlQgualqsJaoykHrLCCq+Dps8ifzpg+6OSLUO
XAGvMNZKsRAgNj1Bk+Q0U8CAvkpx3NKOtImKwMAXB/IRYdVEEHZpTXqeoW1J3wko
g4FkO27PyMIxA4A9t3Bat/pOThOXChGEJZfTcttK+CZePcJfmNM6QvLLzfwa6U6/
ejmaB2P/ZHgypB3f4KkOwDkxtGhLdeOsfrGB5919LUs=
`protect END_PROTECTED
