`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOgkDJweu6KLKjZahR3XxRANn89WtaGY+3dVmSz4SsZ/o9+ug1bC8Lrola+9Xlnn
qH+eif0+L7iK2Vv/fZwJoq1+HVi+IjUI7fbfrajDyQkTGRC8vrhhPrjCxjQ53+6T
CiRf99kO2o5a9fPxEcaxnbUMx7zcHw2FG6OCxJDk7stOmR7KsHDYUI3YGKa48Fc+
msR0K41HAJ27OJ+7UMpAJLuYC6PhCiHQrfMpySZDfUbCzmd1HG6639kvv5N5Qr7Y
644JOi8w3sHjQ7qnxHcZxyPnFwA9vRjzYla+ZHRdQgBIgvmAUo58fUsfxds7RKGj
w7a2azWGRsdhELoCvIjPjFc+Lc8RfIsTWgpAtFqrbQpxrG3KG7qDbIRZz73uzi7L
xFDnkKqVP3Z8rXmA6cBrsmF2S5K5si7Sj3wZ4IrgSJyoDeCji5W47BSu6/pAtPKF
Q5QD77rfH840/MdoFsSfFOPYTRbl4/+aaIRzzH4eTtkcKEuLwyyrYIHI1iH+UhI2
spmZes/EzA0z/MzgRRn85+coIcpjM7AwsK32QEPEf0P/zaamUIzldSUuBDQLRJvd
7aUr0pBjzkjg8GGtz2QrvXLm3Jjts/pAbgywomvaAw9E+HQqPAsFtf7k3gc4HAL8
T2hiL/Zcc/DJ7h44659HnAZJEmDj2GxIo82U4i8ZV2q8yAFFbFOaEa/Bx6JYDQqa
fhcOvVeLbKz9nlbaXxy/fyLOvgJctQWCGCNxAZbj2TmwAAniK47Fg7pthUrcdNPT
Rh34XQJAf5c1wtG2Z1aTHUHdCaDBIKxnm8/CiJ+w9Gyds00Nq+VF3VmJxxobnIgT
IjSgCQEgPFSGksBzn5Z08pzqPCXE2FwJWhQNYX/vgpVL7/kYOuHcJ0As65mBkuV+
qUVIzm5V2kCj0uk8yj365n30XVWXwUwMmc55Dd4dgqy/FOPieSV+R3sM/rgbutrR
EQnkruLiZYrSbWy80B62tGh8ixkV9uwtnP4MzuNYfCJ7eFjsqsEFH6xdizr6Sp6E
Lv20twKA5WPo0fvhVjuQ79SnsU2pZoI51fvG3UlmDPHRdlHJp96MBHZcBJpFf1DF
9zCE7AIImXmcDlk9bn2GXxvYFAIGdjd2hWqD/ZBh4aaZeq4mzHfn31m51ix4sZ8S
TqywC/jLgQ5RbJFNe6UMcJmAahActzsYUrgpN8qfU1mvLzgteV41B9waimf0zC81
d9JiELGxAKfCipKkNatDKiaqZJmTpU1lRAI+rIqb+D+1jUJY6VxwYJSA0YdoAkEV
+sDTuVXr0f5MafTqGJ2Ial3/6eASbL8nkhVH7UaHe9OAHLrifM8CP9kjfqwCPUxh
4sk+CDR5KiIri0h5REz7SZ5XDMpNtr7WGwZDD8lYqSwr53Z/W4MhF2CMJYhuO4bt
BhsJrT0vaNTjWs0Xqh4vgQsRq0GnLyXKmzobZshJkOkDndwc4phj0EuVyAHmpQfe
GFTjto1NmtGj3j7tiw3ZQIvoUFpB0b8XLalV6g9n0BibH0YXAVYGYIaPuzx4Z0sd
ZLA/4xbKPE0KumrnioNIt4jWe8aYp/luy9kDZUu4Lx8yyHdd2EugCJtAVJvZRsn7
3M/A2zMD2ENIJZHXjxs9j40Y+KTSVp94qxRW1VvqrracfEGTsQxwyLf5AFM/1efb
ZlsHy8boU1ngUk/uBNTq34vSTNUsurZL47lPNBKoXYn5nE8cofJKypga/ye/yS1O
3IV08zjygsUlc0El3ySoZSq58ehpRKLK3z8NKcF8TJJ4pfctnMno8wrkAk/CqE4E
Jwpgejb9hZ0ou4Lh453ht2+UsdDU+yn3/mUoJCCmq9B7g6lq+gUqASJCTowjKqMB
fluaI3jELv6T4kXGXXOcLNsEg6FzIGsWt0IT8nLr9GAZeTg9UQ4FHyiVSxSqNDWQ
n4VuATUeE6WEg/U0cxm4P8LwO6h6u8E8DO45zy2RS1vqX/p9qhCay8B2+fGzqaJp
dYHlETxdCKh8Kk9U7r+Yn0TgqEVP/uD9b2LAntwBeCiQEp1BNMUcqnH54cfDTI7g
QtcSlmYDWmffoBt2zwEghcCQC/pAdKWej6n6hBmOsm4neCaHljFFBIOc31mMPUqr
mcb3CpRBgIBJUURk/lVXAfiOwU7ojznsUKIHRu2qqLmlBJFN2oemnuJn5iquIOzn
QYTy3khCYcSNAWqZ4Eg3BLzZrR2NsmvmmUogGe35lzIWwizVyCzkXU1lCCbxRaDO
W91Ee9Kgu9o7pjClx6FAIqdcxQAYm7CsZDUnr7i3Fk5YJai08qxLYYXbwU6CoQYZ
KAMfo7qQqCoK8h00Tdll4Semp8r3hTPPX9MLkF9wgkgDEsJoaDKKAt7eCaNrD5IT
x8ophIus2pAN4lYuOC7EtjUJQ+s3vNSfx7nsPLxLsvrxiZsWWc27L1ZFSm9h0ycr
C79eDz+W8N1CnXfbbhcJSpo5Ed/EcDJwrOCGVXS5K/EpaPMQHjTkmwOe7fPjEJjw
Kazxicr4dv6lrnzTNalNLlSEk9Yg0KHuU3Mf66ydwk/GEp+ukYMI61DPMaz2EUUA
eRH8si+eF+iZN6gmvNaGo70lzHxg2u55lXaUxieEHzJHgD/619efKSOLWVjLPYVW
YoMA8CPC8pXzP0JkSqo3fn6+YoS7dwlYVGKeTvUDtZyF37l6wwF6opcXzWnf2I4/
wDCz0fAjeozebyI2JqtBFS5NW7+MBRN3WtasVaN464rNej+Iz+f0jwydN0O7eZVn
i/2yZBGK5/qYXZrojZPm3iR+1YrgRNqOjuWezETerW7DPjiOnGTb90x2JxsBvGI3
6LnbkndHKbJsL4pt6kTtS54RmIJQ2X8DxrFgJX1RroMlx/FbEOPDY7j5wyq0VBAL
gBynjM9TNe28O7anSGJxl8mdHv0dlv/KrWQbaYAUyYQzN8o1+uD8r8NOby+CCCQN
TbMmUxQ9ylgXGSnl2jnWHwTKkCdLK8UGOiNn9zWwXbmo4LUYNCVfrzgPM7ZeZLVA
JIhaEjimNLKZP2iEkJDV9NloaPkVomoL//rzbsaOCaPRBBJ7qJKMOL9PF9TvKggh
rEkiXoFZ3vMMES3qFTWQdUTaJBnYvT1r/IgZoZcvk9dvmwjcbuNjAOIxgZKR5XWZ
TQRxnxRwGEEUjxChw7V6X3Y155niSC73/XT9nc85pabfqHtVeE+A66+3lWTkmsad
MNrqucjnFsskBDi4RWE5yCQvRddpruP22xp4SWELrLKLJxZur7y2a6bI8+R2EcGV
Ume8EeGexteAvvuz1FCTf5atXcItV/HS2zaKbGdsSUMk4kbJUGsJ372JhSsPX/Cq
Gu7gRkfV5qjIX0/hUSpRywBwPxDVDZDY049CCdGWrcoJsqi1sOGMtCLRuQ5RZw1O
h18OuwmBhU5URsK3J2KFw7hDfdVABrmlYZpKeMXT5SKgGcIufv0F8djdx9wA7l/s
oMrB5Gh9ovBxFHgnlky6sEDtFiEJ/rW63Zsfqp7EJoHarR/djPnoiEYrAgK1QkNe
qIp09D7Irxu/Wb5IDrQP3+fcRFGS3IYMCKPsZkHrg5txm7XPX7WDj0jj5kQa16Z3
FFucRQ+d9ibS5WXZ9jgYOH7sb7R1IoJ8eA6x9S9ficG8ZL0kRzV/DDbRTVLQvXDR
7DsYyAT1D2jeOwxDbBLmjN3GbLlY1ewEEGrugh0IXPB9NKfky/2aCpZr0eljUyxg
A8M07kN6I9t8qtjDmMO1nxJcnsCXBicHG7Ttiq/JZru8coXLCo+cy9n0Gprei8NW
45r9kBibusqyE/sTcAGfZ0naE+g3Y0gYKJBcAIHLN4ONpVv91AGHNBd+lVBTP5kb
mFYBhJ/m/0iZ0tqtPFkdilCXhZNH0CjzLi1xJbjfyEFSNdw4qQGjfx17BRqu+CrV
XrOAbF7/G8gHzeLf3r9S+Z+Q+07RBrqX72PyhaFL/fzRSJ3jfj5840dw6n+7xcrp
DGn/UjAin6oztVdCvyqV0XWwL5RDXOlShgM0QOtoOLn37Hfp/B4f6CLViogUx+Dd
a4/y3GrOoFN0ISnN4ugYoRzIp5ijLoIl9ojeYpQDt6tk3NQ+xFS7kbvv1UFwMLTD
Auy4S7EDfMcnTeWfdd4hRvXljSZxh9tjFaZ2hj0j8pjIezoEH8i9tBmFJ56Pysll
YlwmDhbJMNa/RMEetnK2ngxkv9pPtdZz9zQVv06xBc9gcReg7quzrejw5wE+Blsa
GeW5IsgZaPbF69cka0BS9MdNX5HD6EmzLvLE2kpiRXp1jdjmS9w2tFt9Id6i9FjA
WrEf2ynMuffjCCUGYBtvmGmmpOFBKLRRlL5TLAfWS9EqNOpkg6NpOuG7vt9BAgdE
kNMjL6JfaaO+ukKrXQmIVw95kGLRWnvwqqAV5vpIW0PqO+/ghBTwIO8oKbL+zatC
bTrpxSIWOAPrWjDctGHnuUSvKvf5+9WFiMW8VMR9ovNj0SAaTt0oBfyaPunowfga
oOObG/8AYrrKyIXcWGQUtlzihe7TsjuCpKy9QKyTN7xzI1wdQk1RS2A2RufqPPHM
NYDY+PVvQ4PxlP8oFazGQNaT0afTum+5aYbTnjj+4N26RDIK2dkUR3jl3zt0tAul
Ovm/mrn6vdWoBaau+MpZG/9HQR1Kt5iGDH2sjPqEjqpa6cWMZPFyMmxGPvuJween
vcGj+45/+QRQ3sQ2f/Z2qvBxbKOhK8mdesQFtO4crYnIRAR6k3bR5/RR55S7hmlg
HfNMyHBHqDspE1J4HsCy/xcsa/RR6auVDrJfbMPBjmThZzlN1lzZUBnUGPmdwoL1
IC257zIlUsEaUOo2EhPlL3eKMySxY7Oz1cpkzhCj9lia2XihJ29jwrWn7x3mNq71
2JxOQ5DmFujLDghdEWY02MvWSlBdPcqaU6XH3J4ALkF719StzqyMOrY5ob7/zw8E
YFB/u9Wwkroq4K1vGSMC5bkr7zqLxl3tkQnipUce3eveGjkTqZXoPDAgEZUCrS6D
274oQS0LjSpj3FNMzt9dzplC1OrpAEYZXGxInWEdgTw6oMPq4NTfQwePhnEQagwC
u/7yBfZS7NtWEwphRgI50HWG1ECGIiVD2O6ngX8WaoPMa2914zAzqgYD17VFlx09
LGlGzBrR0tsi+yBUBCsvLepeucWU2UvZEfjvG8ljFoKWdWYcCMjUmRX9Nclb/zzB
C0yLPxILe6gn5xgKWoevQzT67kFTfZGd3jSxc3cB0xK6CKVkWZD9KDuzH2z6CTfd
kU8YIKsvPDo70BD2mdM8AeGjbcxpuJTiL869OKQJQYtRlenmPo2vRIt2ePyEPjuE
hhD6JI1eZ/R6xtDI4ijAdBCx/e+/VHuaKAVwSYhffvrAV8f15LP5iUy3+KBBJQlr
ET2Io5Y0I+gJeHGHT6TSDwSQk6/DiSoe8YxVw3rfkFFm6sJF+pqJur8ErE2yYfhI
auZZ62oqrKplwi142aWhmQ11L82lACI7AYDdAEp4dy4Jct/u6yHOi2xLY5qbiW8z
8syuDfRMfStejrt1+fGIJsgsNeY0E/ci2z+0+6KVZgF1TmBklTk6GpkVv3bvC+OK
5f2YTlTrlfIvsbe3O0ZxcPmxeeBhY9ubpVKIMBtPDW38jHV5V86sVAyvgOFoYg1F
dklGYy3ZuqAlNvi8abF2zyGob3g0YPjNrguMRqIdDUHkSRYH45RhFAIrPCtSvgq1
G7+1/QxQh5aNqogrlZ5dpE8UgpjB9cgpnLHXD4fPM+Ryj6ya43y42ppI+VAZuJVM
xljqOEUWNuKKZhcDkShn3rrIpF/RTeZ382N+sGVhCgr0xylQM3nWaJNeigbusYHy
c/HMdAtlTd0ri56DBTeDXt8a4Vx2njzUyI3MLdHYvyg1X0L90EeAX2A1xi7bOMIt
2heAE9NKwsHohxevYNWKBeEijqfOJp1LzpS9HLtoWGvOTZgvfry8cLfl5HAMgKyu
ArfEGnY+643EfUn+3nGLwRL97D32TnjDccWffI3AYucaka/OIWDxkBGtAzhCW5HN
+3V/UG6h1/VhtM9Jp30Liu/p1TgryD39AMUyD5+uoFhautDvrBmuMuG+1RGVB9Bv
pr2izMuzLqr/jYwrCrmdyCU03YUt9zgcgzYP00Oaz2gO1oYID5o/HgNhBuMtaZTq
SfCt5SBKzaHI/eHVPJlAOLH0HeQjiVBT3kZUssaRfKUYHaJ/SvHenDgb6ti3XhZ+
/f7S/ZFJ0XNc2twtyoLaX7YLpVT6+nop3Qur1FgGD3NXDConn0M3ke3GW8pOq4MG
CIqvMEc+y9BhpwEcgyYFrHM4Lwm4cKFVKSJFe9ccjEekO2jFj/7BoHBtzBjhdWSs
1IxbBZ7ciCOdxmwOqCWUtZWuCOeDG83XzREOZO+UAGt8akGUPzQfRpaUSrIyTBGE
EYJ1W0s/E4MiqXsFup544kh6H4luzMdqoPmh0uylbUQQ7r+GuA/18144Wu1XRGS5
/pmyg2I76D0kArfvLrHTSnjUntgoq5DQ8ccvVZ7Nw3xOxVLLFXVTCQ0muJk3J+wr
NfNWXCr3b/S+1FKHRIDN9R/8MsNIFKHyBAoerpJD4S2HEY7CiTA230j0aODDQVTq
jCqMXz4JUCjhmxxyGrRu3oiWdOmZnuSfPeqyICOKktzSSHtkegdKrTNcuB8ky166
Od12g4/FaD2c4D9Yj+2bPo4E+pZr79ffj9enBuE3iQICZ5ObCV1jzQUxXPddYOmM
ZMBV6C5MtDzQAiIzhpcbKHuiC02p7tiOZWGXwRec+Bj5q3BJpCe06hcm8j+gFRdR
I5FZAP7k6mIxjyGfNLhdQLDZvc1d8AINeTa+Mitw+xG2YSGKhCll8kjFyTXUhWec
ODQss+j0Rb6hY6WJOHi+nR09ogbmdbA+7Db9lMMjxA8lh88oXmT2OiwMLDWrMn9h
XdPi7iA1MKQ49Pl2M0SzJErr4I6wniksOe0hQKkmC3twkw+FNhnlejDXXAAb4hOh
tVQYWucYi8XjuXRR9yfVVkUmqvpyKjNgAbi8PA36hTj1SGNcIGb7HKb4AFExEVNv
G44yKY00ynqnGNMrG9Zyv/vt4shw69xz0iou/t7hdqP+nNXnZBiSeKJ+Xv/6RUEn
Llyk4y4CVLGdsL8MT6X0Zqqd5Q9HLlEGvW9gpxOS36gHY8JGMtseRt9C6N6iBJCM
j52ES/31kA0lX07Iw9EM4xdhuHrc3kmNaJo1iG+PD3X0jSSBuD/Tf/yuhkzVq8if
BlEajYK3y0EQTpkSF3/owgpBuG44luQgAPfvt9zgEGsFnSLD61dapk9RIj4dgyoy
tjK9rpps4cAXFF4Lx6gQGYI/OdYcrfFkYgRv7Tm0fc6TATsLf/KJ3rjAA81yUMkQ
hglEI5ghaHdP98gy1NXx1W9gY307Rlo2bpk7yW4SF0dtYoAf2tDLoJoRQTRL0h1T
JwEY0TOJIDRBh5ZJQMnwiLiQLZ5EGJ0RY8pVo3+cEEyP0POgtrZqCcUPbAQRppqH
TKcqUFzJ/hibUIQvD3IjJ26yo/Ei1t31LeT6x6vdc9ysLG4AF//VgDimXjD1LJTe
0wTfCSy+Mp3Hqr0DG5p3i8P4aZeH0tXVaqNgkYsdwRIXcY1EBXliVOQjuATX5Qd2
r7OBZy32MD+029ufoi3ecHr8CnGYcWqVdadp+4o3g4/8w3roBP3ErhcnrG1CjEpw
DA5jgRJ6fBBX77D+wyhSoc76NnkaQ3YFDBSGAxu4fsF+iwaX38nxBuEOqI919jq0
4Wgti5h9Q5Cz2VXzfOOBNxmb9m+6/qu5tOY73TgwOcI7Bm3w8Xf6V5vdxgY3SMDi
xneffERtDCpygTHx/Ae4R+7DEhgOMIVkueHDjFvBap73JFetFv548ZF+w9pU/x6q
/1pgiv5mxsEA6JZcNIKoxmxHQWXzs56ROTdXAjiocZxNC88nxPaPpG0Mi4kWRdwA
ejRxqttcsUy3Gc+ip39hxJ5zhKqdImKl09M2AWWT0+z65eXGRNfXt8Sut2r3EI2f
G14GcSAnvG0XUVph7V/j/nvpuJrXnustY9GKIAOsKaNwzgIZXr54fFhwZ1C7nnnP
24XSiXHZqOUCeaCQyK9kahij7Kaqf8TB/ilqSD5jhCU6Zkud5VyjU1UQChinlirT
Wc6nW2h9ogC1Ht4LoCFbQL/R3q1+5L0jAUPjq9218jthAkbDiyjAcW22V93w+TsI
L1dTByPQnjXyZfRonvpNAKC8vMOI688qXw3Ytb0LOMwkSeM6vocz9+tWmaoNJMxl
+N9OmS94iSqvAymIsB7aJg1EdCeJqg22cSxrKfwmBmBpUn+yeCcX2FIq9UJesrMZ
yKmqMqucK1HNgDtzkIHdaaTmkmTx0qgVuz+x1/DndLYZCa58ennvjWI8848Sdbqp
8D1PgA/k6gB9Nsqh1Np9xJVWDZakv45OzGgetyGYMRnSv6jXhvJu5eDI8QoRpKln
8xDgF/IU+hZIH48sT+YROIe9v6OSQm7bwC+siQk3CqDVDXnKbwWZMBtg5ltjRoOW
3yniplF9vR+E3ROfbv+qOGm/PKu6VygAPGbPV+fNb7vqNkpdqRBWVUHXSugvX6oo
rFdUpsATICULVLwGCuQY9AA+LTbqPSvyh5h7i1M3/iA64KjCVbfdDbklFsPTnv+k
lui4n4JmZ5jakM80uLxz+psn2azNDUbsiMLd0rRxchTZofyuQQoIGLN8qL38+bkT
IHsk57+iL6WY7ZA1UieA5WB/996VrFGtmjMrZ68l0+SDziytmHOlUQd/hxNj4jUa
IQdbqF/y1qjx2q6woa6GH7iIOgG99yBKa9J/+M+X9jnqiARblTgQfeh7Im8lsKUQ
DikqzLALc/SM5EtcszY+z9z7RodBuckGn0E8XMKXxZNiUcHDunO0himwV1MjkQVX
IgD++i0BZDmsJXmsQQ49/2LBirHjO0V07qW41EMFrirX39QYQA4zY002esOwaiYO
6p+kn5NX9P1ZQ/Qlyv9ktOtQYsHI1uPzv5IxAbKbowqlSNH/ZRn3uPKHzxP5v+Dm
GOjIa1IjSplf8RPOaAnrhIzoWJEIMArcQ/lHV3Yt3K+NoTeD+POjGuDErNj/juT8
l5DbNGctJq3oEiOcWSpmUKR4EOmfG6/X2mB8Y/M6uUb/Jb7/Q7OA9JbSHhvLiMld
gNEivcGRH3JMFI1BYWH+KAgIclMtS1ID1978qPqZm18Gdl8VwnfxjnMuTjvfwO+Q
Z8MvnloDdvqgplIcIigmyWVMW/qr8eXS6ILgE+RauRkVY1Mn++HRV7LDGhY5ULva
VKZH5FFJ8MfGiz0Db3gcdECdBHMmGfgm+MJUbywm50qJyM6mAm0JVj3aZ7/Mbwa3
6ESZyV2wet4Ts78FKMhii4mr+nuCb+pCqpnrKcZYY9XdtZ/3Ck67EkRGoDSA8LiH
9njR6Vx5FKHyusFBPYz6Iru4zpTha6u4OnBv0Xh4Fyyl+zuLlUY2+aH9NmFiFJPD
U3KdHIt9YSowNTVH0hXiifJtBYKL6w88HmFwroR9+ZDRnyZvkT9b0rFp9juk3L8J
OnWuZIAcruhHsN4OR47XVr7evCaMactYA/ltv2xOAZkqowVmrpp6DopabAET1d4y
/ShVv3Aqzkjc6gl2qox0ryzWFcIFgWNS4eyOsfa2f/DTpGK85YyNvnKO7PZZVnFN
3ZZqqhgZc0pdHZAMbBaMj+iNADPhjP0G1+7RIOLJTyKYRNc7VM56O68rVnsu6D5m
jWJnUsEXAiNQpT+FLEwjpFb8HZZPQUr7OnN2O2Ko6Rpwj67ZpGNzUktHtv4Q4YBS
GsQKs6K4wsM/JPeAMJQJqq6xlj1ownAw9tPQVPIazaVO+1oZu+n0UfcaEwN8m0/+
uOkLqrfRuvlxCSQfKszaJ1Yxn1ohD3SjCebmfk5hT2csbRh6KgGcukMJXgKr9Ozu
BBDcqoPEhb20Tm22xpjOo2885B3w9DFSJGqPOFdIZN8wvMSB5Lfln0l+Lxs2idXV
aNQjs50lYrvNVnrvDiLe073gejC/oqHI7iBWnJ/xwSSm7+JhOhhF3bDH1ZSE45Qr
bSpdr3MWX+7sBVjbrS1JX0K2/3oHeCfea5eWAdR6pb0aJpkXp5G8wMAEJ04nZ1Ih
QC8St3HjaGmeP7nCNG5stHa2WI86QfeqadDsMLQ7NCPtERV41S2Ujc0YZA7JAjzY
PME9ZtvpBQNdTN6KWV50Ox1ZynHchqXlAAGPN+Kbi7Ztu/PQlgUG5D1ykeUyoj74
Po/m39Tc5ZhnEFtFfWtrcz/ENlG2tYTAJyWL46mZCVpJt2/AHkN/T4q6vHtdUJnG
cO3O42ATkrVVDqYiN0XcIc6+Q+NQZ4b4zZUktyHa6rMLOhP2nVZUPwqJNKDq6Sz1
gs9PEsAvMXbkVAKKHNN7bw/H5oA4TnLPG4mI5x3cSyHNGOrmJWQO1S8IIs8qZDE3
elKu56xt7q4ejpR3I9C6cPXvL1mKmDQoa1UVD16jcHr40JnNJ5/d/WgSN98LHzHT
dD7dAqwfgy3yML+5znIUrzQaTIyC9rFkcYhkkhsl/zd+9I/3YFtfH0dsKEfF9x3p
cCErOpxeh0LMQ1U9ORX7oxaFsXH6QlJc37chqAkKaBpZ593XwiPSxMUbygeaNmPq
va8hJveCVzIW/hTmZa7k3JJnI/4GoRSZyNjsx0tBnq5sWP23tAaAIn/8dtinSuZ8
l5c7yaRkZBwSps34icwvSbDbeHuwGlgAjeIHRWElQBy9WMhE7IGQDv25K3SoG4rK
M5nfU4gemKE84QpBdozAWvs1Ayy+aQ1Hql61gCjnwhT1YvpNhCjxHjQk7PPq0gCk
9mNuyvSN/FbFUD1nhdAYikqHIgmtFfHQWjs/kScM5NiXXAW4mhAYDdLhzvAotNDn
VoAwvTGpACMBNDv4Rgb1KhCW17FRjAH15/m/OtuYlM8uZKT1Z99UFtzAxwzRtSIV
7frgQnSgq80h4RoPF7nlDweYWJwlktj+wXTp4n2dMItdgF4BJJdwibJcYi6HL2J1
7l/It9mqwTkskHfyst3tk5/oh0zuLY7wN0/WukE8XHfFAqC+X3+nYD9JHuu37h3q
JCbD7uuVbrXQfyZpCRr7Kc5L6GykrSDAGsI+oL/cTTyBx8ZgtD5tC//XElJA7Hhs
mZvVGt8LFVxlRptTua1I4vp0Vi4wz2iM82bBGBNml148l7B8TCuyTU/47ZZsJFoN
KrtstUEPZy30LueJMHxFLr7jqLiCUlnYStt69oxaw6XwiDt4pC39xjRD3AUpGmLj
T8x6DK9w725UCoXglK2OtVD/vnT27JJAyXpMjV7hA1vPF+iuN65T0D+znaiMSmNm
ygApNZL8JBj5voF4a1AhYIHxtAOhJGeLaF3aJ/uw3PUZSFiNsFzW6hzVPmvnt5cD
u2GGhoT+9V3krp+WJ/ITQauRmeErGcYvWLuTnNUvdRFFHwpQIjWuY/nsKwSJb0KR
oXqEkOdOqXhYGx6arBt0CVYCq+wCWc7YzR4Z7sm8LV0/hpyEKIGbX7A43VLhvE4a
B/YtXCJyjV4F0duXPBP64NnFwWOD3GExDd+hhaUb7cIQzoMszeG/gK3BBRQwqozH
D0vcMM8r5+elHpNFA8IoS+tdEhwmHN5Aj6iBGruhrK94ZPfSf4tMTQSyJxASfLHz
IWdBsNohkfiKQvZwisvaaeMKA0LBXcl/A2KejZ9oCePg9ZleTrEMoHMwiYXmhypp
Nn1VSuQSVFMRFFw6LIDHx7hLv8KYH6AApPUkXW5FeCHa04nG5PLi1NuHwN7PoZMG
wyV/xeOqc5s6Vyr/FH7mBW/2VoiYs6nw18VkXZcLZE12KcdGQujlRJqXh96vyS26
dPwWN0jW7ueXIogICoUTVVrj7p/sP55Z4wgfuqRz357Q10C7/pWUmWUSMlZeX0dK
8skH8GtrPtQTvoYJXFOFuPbw7oST7SLRaVn9Qk8qEBlKDW7FON6Y3oDg5JjJxGoX
NQXnrYdFmgpppkkky59m/j16avyYUdTfUtuBcj9f1OF6/HGYdyLqrq7nG0VxLQJk
Pf7nX6y4WZN6gCAJXzaAoCVG8Ld6DhubtrXJkx51D8AiaBM9+xZ4RN1FruOlNQof
cbTgvcRTSIGh8DKetEhrXc8Zg4LKnWatTKglrnB0iQPmvw/n1UJ9kwpPN6aBilsl
7qEywHBPUxdgPrsOc7zEVTgj3AkhSn4um12nm9GPClMwpPNRq5t0u0r0E3+x1SCx
72voYHMaB1OFBab+1qMi0F+Jm1eXvpRDlWyEVOPt6amtxH8SvFrjqQi+4Lf6mXtw
AR8PIkGr369E2b+YyYaYkibkNu4iL03OiZLOPcr8lOsL+FzB81De3+yt38CXVGf0
U8wQaEIr0nAejTUSNOSeuQ72cF+roUdP+OaqKaG5vPNUGxhiy/LbfBxTeW+VxjO4
5ojY3UjaCabb/SP6wTH0PDuGe4rln7WDXFKLeWXtNY87Ws2fHx14PZgg9y73qBP3
YqyVjMhRwuvKiHEZId+NVBzQnl43wLyo2/Ev23BP9nlJ0Ekv2zfd0O0COfo58n0J
Je+1zsvpLpykAqocxPJnIuHZu4DJcuCmvvS+X8gd3/ZVvkTBElsTwXRYS+gj9NcA
Y5UV8k0VzeIOaAbw1Tijcl3AKezaoYmEaOHM5QwhXIQl5rLvtsj/Ji5vSJm6dro+
FKLIe6Zd7JLjd6Uy+2WSExgCg2iWoTbrJY/RQLrt3lejrlmguEQdGbTcBKnQASS/
EXoleTeIkyvf5JzXz09/KD0T/rGxnOgtjGQ+ZTrgck6hK9jg0lzrwQOtuOYHNzvD
JtBV/3lhIAEf8kNCT3qFtyQSeXPoOEbJTQxQ03cq8hCDVJewlplZRGmH+fQSpvxa
9zb7NO5b5y47OemLf+92luuzmGU8Me4d7K9dIVKM/MThDHZGBTARiK8UHZqMa2sV
77su+6nYf4zajwb8loUrwdbx6zFCBKXWW9OncYCWT+07gZD/dfQmMIoByk9ixyQE
tTg47Vd1IiYOcZiNpn/J9Es2RTmT5eSEzJBkjNXEu4+nxRNFHqifg//F4VfuoMGE
zNMEFFBH5LkTtvUoyF7IufV/AR/mKAQv3Fv577VuUUWz9FMSb6Ch1N9xgn7PEP4c
b7pEkJ25yHZ99JovtO5UL+bwLTbshix+0dOSdmrrMBpSpg2BVNj0sCRs+IC/VlP1
43YaytqWH/oRTw4tqormTp0Nn7g1l2xxmZCHxfQiGbeY2P9uwn29ovWMl0aQRqho
pPhvj0X4vlpALmavbqfDlHlVwaJNZU5mcfGa4LvMG5sLgFLclyaHo/idaIFwJwIU
5Kmg7kCIoKrvNJHCJ43JkkYKrkgzmNgR+zZSTanJ4H0jI1F2nozlbWdsKxhhC+2H
BQBhEcl/sWaOx9tjI2gJDl5T5NRRgfHpKtX8qQrbW73YeZA3HxkBF/JOSS6Ptifv
lNqLNVOkv2BDzysnMt4F8nZs9VScy+rV6ZAe2/1/QZGpz8ZnYnJ5BGrUDkl7TsNw
eVOpQIcsUp3YUClvPZ0i2B8KDJDSCioW+HlouGdMZVzCCyoJzbipUD+6/OqnHfGb
VJFH92hznqQcpp445sZKdPYXHAMh+kTHRr8MJK9wZ129sIQ3mPges8K74JGFDjZA
ZgB61O70xGYsnd1pwoStgcC5Yz4jc0Z188XjPYYgecfjMxRv4wIeS9l2wW6T3p44
VmTCbBGm7QwfSEOhHrIrAJmm8HsY8mhWulWYZs2cfgjES9NV9n+pFvAb9dFz9XVG
+ey3RCnoO80+T/hP6z3Lo/ck5ZlNGFnv1noboHafXzHAtBoQdPQtjeEwm///em4l
9yy3m/tcU+i+H53rECfylJQ3HSmytKjb0RmIxAyPLQFv+MLy4tiE8Et1Uq+2r5oM
IraAClXMhWMb1aU/WjnfTDkhdjxFnL04Ieqb7lBoWaRa3Xl6C47M06R8hThHTSbz
SktNrgr8kygcExfXq1uaiu31zwAYj+7TV7yRnYNOdHni2pZjhnFuUQiUcKdNjlef
/d+FKvVOiHBE1ARl8XEiWro0ODLiasenrEo6GcfclywmbB/sJZZgG1kMuJuyeCO9
AcZ0PiQd6V9RJksLmhx/V+PKacxCSO+Y0xXJ2Qgtu0vhFeQ9EE+DS1xRj2mlCL4v
5qd8NYdOiRetbhud+EIEBlc3j0Y4mMaIgSXHm4YIGhwRUjp1p40l+X1OWpuEJS6a
0NPkBedYB8idcDduyglFJGGFSRjfQCbmzFO6qzfebmcBrgMflVzBDsLGi4XnsbNe
5SSd09GAbfrcaH+XdsKHQjkY9sFmYPhNq7p62WBmz1trlaFgQloim8/oiEf8+gRK
cADNsOlz5xsVkAl/7PKEjsj9QSACyLt9QNohNGprD/QaazzS4dMcqJphF+HSgzfG
RnSIY1+MKdCFH+o3w7T6KBnzDnVmeA4Fv2jEbnVkh47GT7NALaJR2pfKg8vXEz2Q
OI6Gcf2KjBaeaPfzLkVFnUns1siHjCLhjAcq4azQJuH+lvN6+UQYqRuNZTHZku/H
aKQX0aDIw+quECwpoCIgZKTvInataRpwyk14bE5K5yamT+JA+wGXP7aTAxCYzkXt
YsJkF/KyfZZmhzh7izj5qplwcGsKwIG0uEMloE/UUKHXuI5N9KwkhuDD4e+asNM/
QSmTkfru5wXlnwCnW6vXsZ1uA+Iemdq+kCzjf7gyeYTh0G0s/uhUa31U+SaRkxKN
Nc13XO3sgfkoqc1TTURa+W+IvIS/QO4s31Td26q+3PkmADefuwCfWnwxwPf5ejwX
WQgXBOfW0Ey23v7SlTHuXrHnPM2j6mO0RlZNTIcQKtndwvuSthkqRaEM36l2KbVp
A3IWJO3yrnyaItj6iaV9f23eXmEmwzZaIBMx+8HhDZlAtcXSz0YJM6QQ4yWenacY
/t8/aG4SJ4nidDLHhXS5eDT3Cqyex1iagUi77qiMOPNO063c7S2O/6PakuQvy5Tp
/seYbQMIrDlVKuptvH54oxi5gUA7jGNrkLjQaN/fIe1pbt1pR6rd34wlbGsKQbYL
YIHIE7JOLiWdrmsxs7DSshLT89pRtZtoWGEke+D3JzVcwmIPgZ/5msF/IUu6jPe1
NRmGHRqkqbcYYm81dq7zRbCU48O3fm4S+iHB4FKaHENtBhW42mR18xywC6GSDCog
zinJue5YCsE3AcfrCI8MJIy4wmtvsFcFVeBhhvXK+ur9W0VJNDSHa7QF2xQQ0xDL
zq67nKjbSu0wISYZJ9se4d3xTGbUoQ+8aAV+qCTinbdwKMhW3pjSGtoR19Ix2pOJ
NQlGsyK6JVnbcfFCwEpB0zo3dZ3WHhiJtlQxp9Uxior+bWqAANTXno2NUVyR+cN2
A5r6vp/vca/vAPVEfXh3ungmeeBRTa4ezk6AuWcPJulUPWoStz4kpFIziyywM34l
KoAddVmDUGYvKe7Cr7N/yRMoXBp5YVJQm+f7wfRiidROJNeHYlTIARDgK8Jwwgzf
kGqYbk80FysXyKflp6jSL0qrUmVP9kPwRQmXe11ip9WoTSUQSUsj+jIrfUf/wpfb
oxUtQjE2cN25ZT+KueDd3+ODCWKj5VfIvxPjDN6lIBnw830+H5/5pQtTaYZi2A/u
O9u8ZqUcvbHS+v+94hsLKzVuyQdCBBYj/9+v8MEShwMCkz9tufCzc6G7VyQO0MGD
DrHxAN5vrSKNedrUdS2rU2RGheuGQ1KGauvS0sKtJ9E3n7XDArM8XIWblFWtZGrv
/6IWcWT8VtImPWzcq4/pZs6L2R5wPFagGWLD8vthoeLboVJvMemhjWAp1laCt4cV
zJzy7o21yRf5rzVuveyR9qsb7WzuBLT2FZ1e88li7RU171Doa0eJGUSgXb5nyc7C
ToiaX7hMwEdnmgrilqtWSMTeXRVYv2Py4LSG+tdtbCwrgbh6MsOZ3yVYvV7Q2WPx
k6pV0HENuAGa4zC8AaKRyeFoqgMVEyvrRc+4Nf8jpVcCzvy4k4VYJ5N7bahaXwwa
vO0gqOryQw7oZx8xptZvkWs8ikY0VGnKHiczbJWUDkd/AAMxQce5CTPT/ttIfWYH
tegsmegj1+ctpzjF0DDEYB7cnCBvOD7zZHTdaHQF9iCmOj1OTAX8fbwOkboVEnCG
zG2/AGjwqZvEm1vw16JjwbhqwUaufggGL/9UuJ8v5b7aDL9L+1NBpmAYQKf4OQqM
9SWAo/Sp1wCdEzbRxlEZgEz5bXxSVyJcows3fM4UCJTi6BRZLJkRDUbmR8zJTvHR
ObSCuVVoCRf/vj1FnrD13j1vFdcrGLBWB0vgt3UqabkGULLcuu9MTusmOP92G4MO
vbwOCQ/ronymuiEAxH0tcPE2BcQbHuhKMQe03crM1HJCSyvPTHNLyBBTavjORioi
9Paif5m70BEI2qlnmg34nfQEMgVl65zUnayBgy1NTw/umMPVuYST/n5rPgoC4291
ppzIc89KXRmeWyYkuYWAimXxioovxJKBT4xyQS+YCw7Is3oZIuCI0Ij62a8KuaUw
RwMvNuaoBdxW2PXnKieCSHMMPhPGmvPEuGaAD3F5u47niooDQ6xKziBn57LLA8Qs
GTV6zW7/jMY0XEqjGZlOf9U6F5oH7ZLpI88jkEfIS3OdR/9/HZOXQoVe/lMyITNd
sp5WnnV0QIJBCQfXHMPY0VroeALE00ypXEVLlC6KCrpNpZ+7qvdQNpkuB/sWmsaQ
gq1gLmVzNWSoxmH2t4MU0B9qj2Kiy0lJXK1mjj5qYeTl9GVJPIAsL76qCOs0ZxUe
40yknvNykMwtMwB2NLdjxz01cWcTjMYcn9bxv2jGLbb5TgGvnXYt35aZu7i83MTt
E0WCf2YRz33fOt5AUFT60Lyixr3HhzBITLu+07i1YMK3QrFhzy8sbh4AUhAFLp5F
BVMKYFJiDO/pwLo/3LnaYfMgprFxvechGTnQ6BNzTJKFGPhZkfs9AmgFiU06GliN
5cOoIYWAByc5l61OGiAKzLfj64qb0XCKA9XM2ksT57Olr6Y0o6fZw3n63IhoV39W
CLp/gnTUe21dMRPKoLMBNwhuQ6U6Id3X53tR2cJQmsSOXPg5AZIVX7Q1l9QVvHr7
SipT2GuODGW/dZVhSlOjJy02BckBfquGeA/xmRoU3mzN4nsd6Wzhmdq8xMxVGj/H
akCGzVOUQskRkcjnPC4qCY4EpivU7Q8c5mXXYFTy4cWM8Xc8r0Yxc7KodakkPq+j
sBRRpo5S2m/7Hm9+4ws1EZoQbvaIMsnPwUv/aLjx+0kH9jWhZas4zMMhNSPz5K8N
t3VHUFeA6Guw4VVJj9NSR0UmQCzIfedEWoFC3QIZDTIZOXQCqZr8w/i6biD8W0d9
5kfxuTcS636pI0/Z2hW5qODYPmaL1/0A1LJ2MsHMkNWqwyTOMfHChlCGP5yqmwWr
ScgjsBaC1vpKCkovJYBjXciQqYrZShYyXV68z6vb0gkgOzgtsmDk+gHReHHc+dz8
+0fHc1bsh05USFCF4YlTTRvUlPowUXKKZPo7VvF1qVO8WW1MeFSvmeNhWFLZ87nl
KVrMoLU3LVji3ToRS2R8A39ujoc7cRoYKXPkmpX9WcAPH3tqUcs4MPd2jKDciuVs
sEp0cAQs4BZOgQzzRaLMWNtK7IyWpYmcfcUduHrCkpTsdqDve8fOfPnvI+JlcO4w
1IWfDjOPnUXQzr3A1tfMM+0JgrsI6TB+G+sRl6uX40pnIRhvViup2oX4eDEgMkS3
tPTmMcgkgpAyRzZai8HnSzk++fG8fOHdqjO9tP+55ykWTJjffnmEBPPpOM9E1W8Y
PBtxAM8ytKGzbA5X0nsDgTDowUVTS50vAspTUkC3ZMwU3m9DFGyuwP3shGFkgR7+
sm6E+nszbcZJO1Ox/p7uXeWSQu0kq9GSMwA9KTvQ3ng2S8c+NPlxljnlbzVm8bue
XTqZcxGR0Txumx/rvDUD/jb8DugdPyLOG9ej4QsBgP2CfZfFZTZYvQQEK2s1SJcg
HtYyokWNIJOJmEFeX4PYn1xRaZmwIR4G5tpzYKGgh4z5RousEjgy/ZlbiCVYk15B
+/dIOdmebITHIYuU5c7sfYjsTmcavi90Wjp0kYw59B1M6ARE11FJLZxu29gW2yAz
WelQL+LUIER+pMg3NQmnlhbtz1gPSt7XMWDKqvykJuHlDLaYh03tNAwGvsW7HiFQ
gjKKZCT8EQbk9ZISe15igWRj8maxjvq76N49IkwJka6gBI/Azm3/NMV1YtTvd9LW
6a0+hLAqgMxWU2DOquOqTFQRHvCeJ/EISX+8/YY1juiGrO7yapw0YtilnfJBRPje
FScc6LaS2za/ZN4fYA0uHcVP3fGHd2JbOJg/2R68w2JS+7Wgjhz+QzLeLBhJ8Cpx
TPYWpcugDgOgwCPPEvuysKJiKbErI1vcE5LHPufgBwFyLC+OFmku1A6jbRwah9mb
90oCXusqAsOeupDIbAgDEYYwFB+6bcg2PgwZtnrkJCZVaT7W1T7qVwSJteVUFiKD
FmC6H27a+8zOExIFEZcwA2s8VYIpJdd53kydcuxmzth8l7qy/dByvcQvZtNEkep+
DcnBt9WyiK7hzMmYqu6+Z1nqBBF3L1EAbHdjpZwjIUDWJSoLLONdWa0vGQIIovZ4
a087qGgVhVenzZfaYv3Mv8OaMyqHpMqC0n8MRO/jdZMLg2Oqu3At+noAeMwIDMP7
8poQJhDVfGlDz27z1ckKjKnrv4FsdcleR88dsO4SZ+Eer2y747/qVCWYIJ9P/7RK
ubarq8uVxpfPrbxbPNzq9Suhv6oSsvSNbfRaYJ4GFUY3OjixS4WpnmJN7TB31KxS
uI7JwxWITRrIf+L5tdJZQkl/3av1xxlFdHKooQbM2rPQ3HrPGEgYAzv3Wiq9nP+a
6g7Sxnt1lB1UAR4J5f5KM95QfKdEnDVYbNQABXJLXGjslfsHjcopRmtSvNNVMDyh
BnDjcuJUgVmmMmVRYcd51N+G+86TAXefJpULbCena14tvxKcdXwZ3tJGVkGykcMV
yOkcyWkYZSBHgZ9B5zqcwohOYXFDOcl6zgVu6Tnzk6L6s0zEnC6FfKIX0muffJku
NqDGP+V2s4TZxUFOoN+Sm5cGIRgfsX8NYsRR04Ndd6VHSG4/kcKFTpSLbKJn7WLc
VvDLHndVzANCmhnS9D3gYJwzLmh1PRgtESMq9uMuktlZhdnAA313rsz79TbspLUU
gTPj83DBgpRvbvzZvlc4D2DUT3GZa4K0VS2WRqS931eEdllLwcBSgIZfVH2wGfpU
Gge4S3rGrMh/31JtlPDOObHh+SyIKKWqZEHbeU0kLnLQqvtgGzoIh1w7VwCyOtgm
nU5qYSparFTzUax7yfKXuy1MejgQB4i0F3K7OW8bNj6ZHwp3fFjThVGhOZ517kxj
6YRkSIqUmEUj6AVoxSkpzF3gaXAgIPPViVJ2Jnz0p2gY3dLZpO5y5HhSQHhx1xLY
5KrO12MW5vfA+q6bZbTY1RDfXv2C0nttiY5v3qizNjHu1h3TceoE0T40IkoVE2Pj
an4MoWdf1v4wr1NRQukMmxlDTV0MChmeI9ELQ7Env7PiJdyuc7rwvMI9gBu7gSeL
9csnxmD/PACr1+PCwMPBksu+Kf76LNXSvC/5zzRL2SwEFHHD1PXNej+7A88YcRGW
LAr/lNQtQxU5ELFixrQOH8cdgDs/OyNuPx8Nwa+HGrV72JlORHN9SQikkoiYjI+u
merxOfgLZV9kwNBiH2k3O9rsqG9DokcH4IlHOtRpnL2qYQSG1MDP7JY51nAgwIsP
qRjzoLTVKmY+V+xwbvyBa1kHJMTOHTWtr32MbN8JWvybaSRbb3tTZGCPLjYfntJC
zgOaGTr8X16SRkDUTBIVu0mlvozXdHIPmYUPJ6fUpLC7HDPcRbqD4nGFKWBan6hN
/bnBEMGXFudwfp9z4frcQbm2ZDOw1dqbd0txH0+nN6oug3h3QjX0uzKmvo0/wTRw
+Lh/iktmHEAdl3AWuNtI4XE6oJMM0Z3Brx1akiuwDO7A5p8f9zu3BHY9dXzz96pG
UxLIswjCPNzn9ftIcmvxq7ptA6A1q0yb7CgsBaEILymw0VQAjgW/gEbIDMA19Pp3
cQI73b1JtgCxDFh7r7AFu5Ml5BkH+U1P+WQ5dELgDzIc3z3BEAiX5mrhiR1jaIJY
z8JK0C19Doi/hp4+XbZAaHTpwjQHz5JvKYW82YBhfnQAPrD4FD7ppwtPcb9nf9op
miDTPbkAkOrmRXjj/TxS1FEU+XrVXVd112zYkWPdkxxV9fQun49M+4+2wpGlfJ/I
Ouy1BK97YrpIj+2U/XR1HxahP7eUNbO8Eu4yynT42FC7x6CYJ/nDuoXww6Ht6Plw
mQsQ41Ex52nfxcyZu0ZTNky1HVnSQ5HGbOviw+fxVz/6slCawUp+sgTwnWl8K2Qy
HBAxaVYJ5fqyVoV4I3vtm82FOPiDkD1UHuTWgwTP9VcrBWkRhaHsaQpXrwUXtD5i
LOL/9mzLsyU+PufBOnh4Icf9bMkehA2vAUDzvu1uV1kDfIpkT0j0Hn+sqbRQSL0z
7kanDvuIWfo7wwpgvpX3CudDK31x9yGJGBbUyOtI5+UZ6xg9L6KFkAzZ4sTtSlkh
w1teOCYHpwA7a0MIosBCtDs53zHJo4KkJDInKW77mGl3zbYfTuq8nJDQB/xL8q4Q
85bp6R4kkpapJNDUp4/SeraAxHScuFM0fFgUmxhfUrISzwk13tqxZ8o1EKD+lZ+n
y8by90PKc2qndMpMcWBu+LrpDAO2o9yol4Gc8YQl26RkCyjbdGBrAkWM9GL7ZXnd
T9wvoGPjjWPGNBgVduzSMkioxH8D79yFtirtncczdl+VSWx2jGh5bcFhQh83js4+
Jj3sMOhNVmqatW0lbbx0Ez1SVgvCDXjJjVzO09TRkBXLxmHWmG2afudHc4+r4gwy
13DH2KOvJ2B/qzuBQP/p4X+mKuo2yuU97+pEkEIJDNIvQR54gQlGcb62bVjw1DMu
ZoR4asZCCwgs2EmuPC1lyeI4Y8D3umYcsWidPU9CfCS6/QywlLJuv8YKDJy0a67K
hQp3forIXgXL/ftpUeqx8rF61TyZ8dQnFR+rvbb47Y+RSx0AkWosd169N7ZLcbQ1
A4XLH6nqfpcCmla8LuEv10fxrDRb9Ps4txUwSFRGOdhCDm3gswLXVrGCWuS/lt3h
sOudjsPe3C2b6NCgnj3BZ9vVzghdgfNUiRke7sDWawCHvsTtjZ6HXvbFpT0ExbSP
CSE9Sf0ba035NpiuPJxMZfx03DnPSdbun5qMdma/rDBSJQQPR+Dle/jUk17m2D8s
eWdcpRr82xoNpPa7kPohXcCheVqplLf49BWwm5jF+w9tiaxvxbtqOg/Oydy/QPbt
IXxW65y1Y65KjeZixf70H5E1AhGh5Rau7lsyD2j1JY8mfNd6ppAJ1zDdS5DtiuUw
JMG6jrnaYGTuoo4OsQuqZQiM3VjV2aTs46RVN4peC0PatSGcQoaoQDo23gtTqKGf
AEk2BWM/f8vZv7qNJBtxKni4LNAsUjBY4W9pNu+NjR/W6SitmpamP406J1gDTsAL
wpGZLQpRXSRFxAao5qbpFtT/jr72AZLjNJ9T4DfP2L2pRa0dQttdY3Ed0SxmAOkm
6xdqR7KfAnxkJPjx+DjaKNhphOvzdLoQZX91lQEFtU/BiBIaRQbv6YPe2xiupLTt
SBD9jmetOIDtu5AX1iQWhx4T2bcRcRUJ18aW4HnV2u0ESPq6O5SYMMAb9+m+iho+
qE41Gdvx5bEmG4PQ5hgIYAT0r4ddFXw87nloN3Sq3C0ncNWXDcYGISd5rSzcxyyI
H1OwFcksduXhiCjOOEgbB5C7c1wkTEFygbX2dcfLY+q2eglPHP8WcYVYv7q59/ku
Z7zXsYA58hq5rngbMFz48jdh5l4RVnmDxVOPUbtUxksvDCf6sk60Eui9x8IbqS7O
IhnDLiuvSVJoiF0PP02VbRe7zWBjETMiY3cnc1Qoo+lUzE2JDmVFFl7BwCbAO9kw
y2Yr0vLXfgUKvCl1YB/Z2ZipHZ1BNGxYh9R/gMpRquykB0pvM+cC0xzMRTKMP26i
24D+5Pyl+9WytE/xQlt4YKHPdRbiEYrUlEbMXdEHO1qBSRE/DNPx7EPOwmt2IuUh
Z2VkB6ZBJch4spm79oTJyf+pwhSaMNv1Z7RuKgJDmI6xONx3Y6DIqz69tFcpcixP
7PabEGjNhuOZg6Fv3+xr+WpsDDrMt10y0NHr+fAs+exVAPRyZalS4QNZ6lPz4YeK
aT0JPnyXa7qTVH4a0ttC8gASGRKWhTbhST9KrhYIsefZGoYgYvKbMnrRtlmurWrj
lYe1jfMilXBiHrme29Ue7DZZANPfgESfYll4yH7cNiB0YzEJ8b80Kj5rmQQo9lkC
AsEzWIv77zC8hMPBBn/johHmjlHFYtDdYzZV++4oh4kdXQhZesYmX8NOIPzwBOtp
hzD9YPomVjjVLiD125QOgZZSwFyZg8B83epcGc2q43lCjkvN6j2v1FW5N2hglur8
EkpJc54ebEa1rijznEt0LJCJpoCnqKtgZpujqZHiJGZ43KBMtp+kCKuA1cxUaOnm
abJFXn+B4gR0UjPT0tOf2yZbi+plHS9z/doaoi3MTARGiZKlAgXC9DCCTtuLt/ZF
+jHKUCqRXh8JhAIF8CQncrOFmPk4qqibylBjOPn2SkRDPJaejouL+6ypwQl59bzm
Tf3EcoJnRuT7XhusNNFSue0V19WAxcUgYPJpDl6PkDdWXrxgFfQgLwsaC/OBPJ7o
d6iLkNnW0HYHxNhJrH8kSK0n0sJ+QV77Az0FX/zdwUW/7iUKo1b/VQh3e0lW2Zlv
NhWFHeaJc2SXGmvKmYaKLRxsmeF1Y77+lvi148/lCbc86zcvFZX+fml9QOmNn0C+
85eVBlRcaPt9RT4cm8Z0gyq4urudwuP03wLUc8FY07Lbn3jqq2NXg/uTVCKJwVrR
jgX1YiGTwJ3I+rNAPRMOg9FOAafu/TEF5vDYS4s3coWAxerxuB4n9gPEHKTv2EII
Lh7XXV/G5szdhV8jhznxUXu2HTVgO6q5+UuSSR629PfjYpoWnDUDGySGBEvPgjbG
Uu/8FElZ4zaoYoa4IvziYepHFGVm1Oyh+u86tO3Wu0lRWs1PebZR0neagUn8ziHh
LMUCcbkHUNmTUUh19hwk0dPcX/ci4lf1P4zWM1/8/tj8md0yvd0OM+aiIIIqqCe3
O+s425ncsRgqHJrxZmbJf7zOCnpND+W000bqKAoTB1/BcHsrF7dq9NUrLC1q1MXw
GESjVRODXctPf07rCISwOeKe/U6Z7EOPfuXM1AIMFLyXfdY5EYdcvI2fzef773ZM
K31bMTY6R7k5hFl5IdWo95u1WDylDW2CqRxHLhuvBb/Qy6SOJ9wAWdnETt9gox8g
J+eCXW8DqBmgHJdrXeJI1viXPgAGePSpP8sCPcA0WznpJl8f6pb3QrmFTmDD3UHt
OzPV3htQPq/OHPPoY+4Xa6eRGRJM9P11wKw07Hzq4D6yTfOpq+LGxzDqq9qYjXSM
pV1o1DM89bh7fpSqqBTPCQNjuU0EdS0yrX9KDmByq/LSCzJ3e0HkpIlvgaScwmLP
gzLkud6bLGd3x59MxPgvutnuq/ueF+wTUaNajOfrQrjzvYi1KPCibtAeAdrSnV/4
9IXaQWTURJfXf64+HRmJU5UwAol+iu+lZAoPl3a5GqQtljjdk439bUSxvVWGaTMJ
aH+LU6PQy+HgEFX+NT0nOjtnOz0CMrNKOc8zR5dIJxAm0S8nV3x0hwsvEyluc0Hx
Hl5CNc8q+Ao9L9tbG1ML/CaclCAbGZ4i5KVJwC8HJoUL43fCTinTKhEEZ0qSt94b
G4Abg/XSLDAPcQenrY04OyQboZb4yZF0a7ii2gzla1JhV4EEd6/P6MkAZDHM6z/A
H1+RTxGHcP6q8FvX1u0eBFYIXPSI90I7EH09C9kccY9PMdj2b5LlNm7A+ELhij8P
l3m/inVhfxc6xEllVVz/dRqDjSNkHwAzMUPA9E/Cnk7/LIBRys9P+9CD/9eiHBC8
dyaqgrcmjb09tXypZUwK3MTJfJiBemfnHr0XWdoXoNhkBS54p8eH1IJ6wZByxVKP
eETdt5oRLpHAvQe8r+qRpR50eqMUbRgtYpmmGTin2KZiqqzjReycMtn7eBo8ijo9
1nc3K9VXfGdKHD+uqOS6By6v0eDSGk31hg/twkL0FDtgEjTte+MXjj7paco85u6b
anzf9POxJOOmWYM38X0DjQSmuaClujG1dlWFEiJN83QVYdc+5ZC1hBtY9pWtvSTt
pxUMTSDBxrDC7WbfxZNLyyMFRctEEhRgrQosGW1vZiyQ9h2X+ugil6dprJFLlVts
Csr388DzQU5MQK4iovaKlt/15E18A38DxC9uXU/N1Vw0e200NYTD/8cOlRJaxrp8
4q5WfS2wJoOSX52LYDH8XOzauGkxRfEH3VuiMgq++CkKU2z0yuerW3DJju0lONYn
6c+1aHB3zQ6h+81rW3q/CnYppkbRl5MtzHpCObUVw4GTINNgWFbbqkhacR9p74Oi
znovfPZcx15Zl6GNI958fPGVEsOFHw0jMC6Hkbzl6+nXIN4we617zAEpnIczVPSW
dO1yQvK2MqvL/Z2/e7kNH7VLodR1m4EtRE/u8XnC0MkJ7HMWHOfJLnXxAL9SWuZj
4gxv+Q8ei5BMXHlhzW1NPfztwAzZsQOehI6SSjAgQ2SGZRpSDKA+heHeWVaGrbkE
8W4sw3wyCz3w89XHxZ6u+QSUqxBNmCCWYWJMSJHS0atUojtCtRnUEY/u5D8cz5cb
nZyBWVmiZD5KMI1S+TmbE16wqCVAcdkqjzSCUWbQ2x7oyRu2r1KUg58OiIW0aS39
0IKYnGEb+SjrWm66lifRojhVJEQC2gQb6AvGw//83pPcop1dt8FyiFy+XWjGhY2K
+edgQZkF6wk+UtxnQlKve7QkzwtWOefv9QE/QK1HZP0Hy31QN5gaA0fhzypZjRcL
ZQvqkHGQF6ICqCSc4pySohqEBPCGYa1GMLqPebOrlDTJn9AZ1W4Y/Ldt1u2EK4Oi
Dphp7zC8vr0SSR+M6GT1aDDDTnT/23xMl3UvGCMq35IVUST1HjpQfaWKSVf5MWZD
8AeKnpVspmThat4CETCg2iFRVcgjrUuK/jw3wfGmmWKXKEDpk8ydsne0cyhGAina
TbRRixVuUQYpzZ4ruu9+2bEzqtcNd6eGITMflCdRe/sV5pBifwH5FrZPhaCtphJy
kc4Pf7ElnO3/V6jQbN8kDqK2m4Mmog5a/y9b73A6K5BkgLOqIs07Xu6uJUZ/Mrq8
n1zXRXt+uGwiWy563B+cmW3Q2OC1r2iEGqkMfXjbRO+hdBBn7xLQwS0bHFKC1Sec
qwLCnR7VZYmBP0NOEm4enR5ladP+7Y05cKpOb8McOMHqpfsb76p0i+eIubrZ0X/p
lNQdxhItgyDhmpgAtXK8Abh0lo0i8u8ocrrb2WjxCdPaoEM/UeDIVvXhBtLx2lTM
cyvAmK+0kX2ms5IjM60i+uV66f3EqkcGGyCHL+CEAjHEhSo3ef+WbUle0D9DXpPl
AWWHVzJqvdDVR0wU0U6kGGoCcwUrRI++CLlSczA/x395OCRBsk0dDnOpH6tVdTZt
7dbvqajuTcAUI+/ynvTNb2aKS0r+NYQzkEttEaZGz/w6hihbpjWcKRKpJ1/u93Df
ooYEWF3m4l61Jr35uRYSTOdKcR44bVE1LtKtWROWY5u3L3rZDL39y0buQp7PYMho
sw6lQVDHwx9JjVgEZX3vvJg2MhN8oafe13BFsMiu/gBr9O7NH6LxR68Hg7qmjtlI
MMENUTwTK30mPb/s6h5l7mSvKErCyb9I7L55jBdGSORhfsOe8dkKUinGPozvtrcn
TyoGq8VgHUDspwC05JhLApXLJR2QB+Mtv7qnA/d0ZR3eooEaoj1uWApa2iigIV9X
ROf1Ffc+5h0ojFDydKHtpfs6N45VeL9chUXKFi+XG0ZP5H8rbU9EHLOtAYa8QZ29
9qVLw+3McMpjB2t3fH2lkPKYI37EZsKneDnD2wiCPpL7AbuCIMC8X6TkQCHny1ag
bK2RTBVVZKkI48oUQQo+soTCzYL71l7x4GbGf7l440Sl778NAvIT68AblChJSm92
uvsco4XloSxinCZhzTtu4rCFkBu1wP5cXJlFQEkkXgr3yp/cBeBmb6qbBYFUevN3
Lraq2ORZOJ4WhCk/0ilFbEP5Aew62bCTkFZeQvKb/+Ied9RTCM9vR+TMb0g4tr7e
1/7h8h+3XRB5GnEZr4NPtvwNsDonqZEZZFICOkRDwDhilpVeqBTewfO+zi46Yx+q
Q2zxbB+rUI1VBQAqx1/NvEhUE0zWdRiTsRfV1uOPAtPlMdh8yasn2S3+xBCzBeCI
9EWdSJs1L5FFBjO1JwZ40vhszTLZhMYORuipF74Bb+aC1ZyrjM7OMc7dflakL3IC
U7DMOpIQfqcf0kJqZS7vRWGytIAuIBaWzeaC6q829wQMIk3ha60YtYYsOTRKnUe5
eVkiqzMPurkIO/zbfjysEaBLciA1gmOFVXu/8XiqOSLe7FcEym++UBRQ1T8tL0fO
gyt1Y97S3y2VT8wdRWpGn+2vj4V6+ov6XxY13EF23b/3U2J6QXBozSTpV162OYRp
3P0Jf1uu2hz3R/8Zu2JTl64+LN80VTy8G5Mlx32MKc10MqfCovfPFnG2Y/1GNzFG
emYTpv6+lgOSL4V0Nz45m8tF430EpT21rR1TDS4UE5XY9rG5zGs9mB9yxxEE3x6A
NL8Q5wFhM+pNyDWxFcWgucQs3MvKM/WzTgrnrSdvr2/jGTF85GcIve1Kniwc7ApH
cLhgz5dy56mKbi1DOIR3XblV6jBLyGler5W5Rwn2p/JOvtTlXEy7oZ4NyPegWkIH
wf1zrDOKCufj4R4pc1r276eu77aGp2Nq/fQ0ZvCv3SK3c4dyPzZTnYpddVGJvHG3
4BUeNLmnGYsugfuBKcpjTkpkTrY7iiWa/u9a6VF6znTKEW8nPNIEHngSXN84ZF8X
UQL1KZAxcqoW3bj2iWUdVWmnITZGmGu4JdWk8lV85y670EtS3kGmbmG+kBcZapNX
U83h34NQm4dc616dnCI3ymFbBOc70hUqAjZ4xCf2EFFwk2tijJdwS0D8jfoEFEy6
jwcolf+2lIKZ21WNRtYGM7HRKpIz3USrq9ZUKo/9wcblmcfY5PlHBCjUEQZFIyRk
VPTgsx4yWAd0BtkWQPl4SnodpfRnYpCKbsKiUSiy7rCyOPZMwX/p4mB2WPDa5l/w
vS5156gsHuwboh6vpmLCrnXNq15dHVTTz5V+i9Da3ifm3XP9LVOJBBoOGAp0QNYz
9cLKXJuZSIn9YW1vLqI9McPhhl380wlgljTT13sezzQpzgwNnra8IQGGe+S07hSN
/aIoMh3CnCI6YNu7YdIayg7qnhdSGUFIO+FIvEV/VfbiWx9HHvX1TnEjb0QBy3eY
GSx9P1TkXBQ1qe8z6cHC60T16jdf+SQDsghPNLiRGPvteE2pkOWsjFWY2Mt8FQZo
h7sVv6A2qcTnvoo+x2/jIpEQw3xoAWjGmWHD0n5aEqwwytlrwDkerjmv1J8hhD6t
91998fdvymVh8Pv8Jak3i7+9AZNq34uuseuWy+LJyB3V01cW7zdA4HPRkNiVLvo/
dGaCV3ntHMYg4woKKlXN6AricHYgLAYPsgGgk+2oz7Zt6SGo594jn3l7T1R71w9A
T99eZpSFnqhQbkGjA1GWdc6N+WkIDUBZXXktYLjsCYV+zrBbZNTgE3W6nu2aT3sf
6us1s1p8FvVoK19no207CPz15AWxit2GlHepoSpP/CZAxhChWlj/9YFzAbp0ofMJ
ZoUINeEWvWUfd0mwpwvaSp6V3ImV6lYJRfBP63hafO3+S59z2cTf4feivlU+6PNv
C1ipZWuId8dT2Y82yBTL+ku7EGTHKTVt8JAhVAW0E+YiXi7aIh04XBAHvd/t96T3
D6UgtVTZXrYDVjD4NgfJqDnOrVevjpDZmVNE1grgfUbgTTSl/So1memqLQsLmYL+
duknRZpCzk+J/YSyUU1YfJCvqlNUyZgyIMEWj430YZewigFn0SPmuPp5Swc3zzFj
2BYb3dJkQFLK3wiIeETrfVz8YIePjFX9lVlwjVwKg3n4/jQarOCofZvnY2Ue7qX1
6foo+NrNMvlEVNglqi4XmzxHJ/B3JL2oJETKaXhbkZxPJ4aEeeSaxuQoAPASXOKh
hvBrSoHef6hHuuJjbFRjl7x++OrHaCVqLHlgrN2jePh6pWqi6VZexuNA0azcx7PG
MZhkmpCd3fuOlP/hzANzjC9fw8Rrrz5hGdDTcoKlT2JKx/s35DkBTKaMzwD5kyQ5
7cdM5zSaPgPq+cS3EkjpqJe0Iu0d9GNjFPAD6dZN8IZv+SlGCwhqKDqs6WhDxC7D
ODEJPvTHyMfOh+rhd8u0WExl8ybV2Gh9POs6fJEu0jkqjatw5FA4aJCkpTqdgelr
Fe9DaPbXN5UG8dglDiWa5yS/AWh0bjWTiQm5uRQf/u0pCNW+Rq8aR8NzvihfZh5I
N/W0hZdrd7H+jYDnwe1Jw3R5A6IViOgyO3Behgja0/7zzLcSJ9GAOuXalRKcPGSr
MH/NEIX+5ptXz0BwZacBDyENq/IG2NKz2nlCpitgnsa16JZlijBYHNySWnOeF8sP
DEKCQRFWACq53lXIXgXBmf95ItkMO1iBLO+69LspBOJsu+1Mlo4LLLhFPgex4KkR
qALHHp6dOiolbbqt9J3FiZ2Sy7/isNfeQqpyGyKldgAFPajAfzOKHqXHzWBoQ1CR
w539fCYOaJ+SClSm22fRssLE2QOFs0YtvJAIHQheyocVxHlBg3pV6BY1+mOBjsxf
t08xLJyDBZ/WOMq/bs0sp+JH/6XGTOQLewceDjKoT97pPesqJoL2SU2t7cUdo2NL
3bqps7VNWEheIOLvQR4T17Po7HuB9y0SGR/fXFCXfkj7jeBw9JH49nOrf/pua3J/
B8cbVUzhVSpo2BcH3LmWv2by3IY4QQUAPDTXwW8I0lqi7n4eK2ao47w5pNe5QDx9
gJjZkhjOLebQAR2eq6NH31/nrpjpY02WXNdz5WJdWwQX0F5xgcLkcHE+brIGtPIs
9eRBHyqWAsmBnceJNqn7/91/O/23lH15qRboyZYQiBTS8u5VtBe3aT6FCHEqs5qf
hUQftohFV6num97iIpk0HjmQF8tX9dHqarN690A3GoyAQS8zAXY7DynGFmE2q1G2
iR8JDR844ffNk1MxTwn3N6ePTy/BDTw3r/Z24S9giunLvx+6SpwIykWaGgn12xg3
9rtRNhSOvOkW7f400KlIUicvz1zQ4SaWbnHy+rT4OdEKRB29eggug/lgzl4SGz7P
D4YYUsCfwofMrCOU5K/0z0B8Adur3o0h/IEq9ClpUAymrEPemlnHigCbnyS63b06
tjw52+1PHYEjsUmGsVpkD1NnXUXUOVOM/Ff5ZKppMswiSmbY0qgLy00x9LfQur2l
PzmKXDjwP/zBUGhzrETvW3V8KhoDc2ADAUS/MJk5iU5nCKsrOZefl1Ar9tIs2r4V
UriKAEnfLHZ3wYielr+KjcmSDrBQ4ycKFpFORfUKWu8bdirdAzOyDcInxy7vmfC2
fz2k2kY/4YA5Tf0/ESaKY4dQn0bBUM37/9WC3u3JKYiZaIaaX7z9JwpIHUGlNLwj
Vbv2GaIQcAsIjl+6/Rn03DYf9BHhEhQwmf2uQ1X6HA+t4b46K77TbuqtlEP0EkNf
Z2wjkH3T0GBJSxUcy9ww+ocQrD11dVNvyl8Zg8i0gg8v87LRBG+89kGbsi6yR8s5
9FUJaIvRAuh83/ultdufYlD0/i/lauitqb+cy/AnCVD6jGuk1/1T6xM0edZDVIoD
CyUfWlgZfCS8rIuTYBDjrybKp4V1XNGSIKoglfam0gKPaL5rWuTLuyuvq9gS8iyI
jZ3g7vNgUsXl+Zk4tWyZ0MFsT4OCeOCpSCwK8UJ7G5kDAa/w/Q2PlaefC5WJP0F7
Iy8MTnPAF2j44zDPXmYQrHHijk9nI70+OMt/uPTbaGk39nWkB0caETQxw9z0dFA9
Y/tZ5e9lHOD8KueKFdEyt7h9beKXSmY5JQ5BsE/hcbYG+7gPdrJzxzegY9o0dfHP
2sIsEtd0VkXqaBl0PIa4Ls6EfVC0eKmnxff4vzaPfsz4kQ2IkG0GPmwcfAoEHowm
jCX8Ix+gfiAD422r5CcsSg2kq7xWbNaoyV8FVd/LnMNgyY0wrerKU+XPNu/kcDWS
uNwpXtMPBH91tuFhArDMEHvAa+0e285uqMQsmXmT71axRSzj15vFzzuah5HGAF6q
KGdu7oQCelKEuP01M+dxhN4JsbQWIZbo/5KvwFRjN7BtO2Yc2hqShfqReZvnrGpI
9cr0E9Aa3lCQchKCufIzVeGSGqeVG2YfXpH+fuo/1rxHMXKd1FhVAdTsUgEC+rQY
d3pv141BnSn9XrF1vtmTkNENBPnQe7YwbzNCT6OI2SDLPV20xkdUdr8VOLDkkiHH
oRhP2IMzR7hoifu9UCeEHrb69x9f1cFS2qstHuulBWOw8Oqya894T19FK9/xKmMP
jfS3nKdk7nCvzd9gEB6t/GWlJ7pw6BX6PnpxtyVJjBFELhUbTD3NiL7xjlkk7xwz
iFp5KJ4MZiuFj90/TH+Ajxu6C1X3mK7mGm9ehEthWP6jU4axk6QDPXC5BK5u/7HJ
4c43wqg6Z0v8dvY/f+BR07ZsiBONd6WXt6eQmKRGoW5ULyUWzzdFG1u9KA+AarvC
yKDDZ9z38aL6PrRrLyEaqw3s9C88hDxoPBd74eivxxqSaboF6Q1t0tNgNXQumCOG
hwE+Smtpcoqit3C8yL0k8GYornOz8bCb3MLNTwfwW5exlCt9zPl9N/s6X2BFTBzL
3qFKFoDBvTYZe3vk27cyWinc/a9x19SaJAOvFLhxjLar2CR5h5NiemfqnXEFtUhG
hxueWR8O2k82CNNNArbkK8pyTCkBwyHbjO2JfZxO+U2wAl1WW6XZEU7tOpcJVCcp
/5dmVBgG5O0tOxEINJErsQsPRifn6dppYJaAdBerwuRSx38exOSwnnbARIQhHiw1
Lqq+NTFFaitbtgIzOxnCZ30W0aepZDP0AGY/fk2tE+0oLlS0jVGp4nXsmUd5xCBS
oJk18za3Dl2IlLXj6rMrCWifdJy/p29aIiohLPhP8q62w0qmk7LKBLDa+VWyYa56
Xfyb1nrcEwBRv5nw0KdiAGwrjtgK6qIyloBTzc2Rxio1vmHnWkmhaWhywjY2E9Ib
rqK7HYttXsxpvwoJq5Y9nu3Y8elErON4ATfiv4F6GHX9grNa1CLnseAX9+NrwzFn
0uEBDPk68e22ZPox0MGZ7twL8IBc7D869bXh91Q39zE0QzQWKLW5DSuv7GKj7Ln1
+YbEaxk82vb64tpeqjhDfQP4dPqZq0EIGn9YUzedK9vxII4RlK0xF54+BdUQhufp
bhlFS0+uHZ/s7iCfE1uonmziTu9iPs1SlY34C1gpEO9AfVVhkwPiLSEel/sLrqYk
Muyc9NMiRUvX2WI8QFCh/QCECbsGTnKAwDXUWQ3n+j99Sd56XgGbF8JF7g/wqGn8
HXmR3IGBLQcOHG0e3pAf1EDFkASSQsg5Ba4IoI5/ZspJj+sD7A9XhdUKQflSVavO
GzbjQRyonLsmJeulR8Tmt3zU4rGK+MPLL6Nv9pCcInxV3Xqsjr59kkSmx5375iMK
XniWjGgdGCKowzT1IY8PTjfDOS3eUCgzh0zDmkFjkY0oFDg2FLcaNIM8/gcam3+n
V6Ab3Eq4HwWhU8TCO9fsnL6uLD1ISgx5HBClyr91Ib2jAG3NmcckQd/osUixTdYX
Py0ESZB+xGXu0Izknhm1EnAtoclN7l6gUpUg7A0WLI5wbA7vRwA0LXR/osqAabhg
vtS40PiOnn4i8uQZhS1z9CHCsDM474VPt8Mf17cIicYWGF/+DXAWY4LkkFFOrTtW
Hv90ef2ss65Ulbk+emqq1xt7X8COgV2b+fNoEBRh3DjwtsCjRPjp48aG4ziTy4LQ
950smfLlFnmUKKyUcx/OTWtLhVvbI951ZME5epyvjOtTmWsgKa2NrDTwnUKsx3tF
SVemptToRn8sLlP1NI/DVg6LGOI4FNeb8OHuoNNN7NBw8ZuIbCehZCntcvSbbZwV
oCpQvBv2G+fwpBMzvlr4RL02Csu6jyecUfTOa9Ykc7LYkk7JtWujy6emVFbD1Ocn
E/H7PtKtUeVGF1uIcU91k6Oe1omvWuBgaVO52taDfMhbTYLRZcDi9PBK8H5jXu6g
PKjFedTkOXLjBT0wY6ewRSMq68HqUT3O17qxtaw/1kOylsm2STifC9ialwuefdmc
2ddYNEB4kM++YA9PSHgVyXYZ+lL4/xzzdK6P9na+ulrX2bsKWHPafzdnHtMlMj2r
F0v33MVxtDVlP6KDULYvJ9J/D0oqzlENvUiqeuSFlNTEuTEXt5t/65qy5NWiHSai
3Z2+NAWaVztTPooQKH4EWMAVptCPi1UALj4ZBcGavtXi2uNOB44q9gJDm4foaf7k
ag15nG77dUfmYRKKVNPiVaWvzD3PFsROgmvH9zGId4i4fMx2XLd5r+fAzax/qgtt
mMavI/pe21E/R2LdOXLwgSjV3cPIEqDVpB8jhwzSuSjhv/MT0iIzO8+NxpHkHjtj
YB7smJffuvWVnYDPd+uNzDJysk+hPjkabGOca4JzX+8hQVBOXe/Lop4lBhpuYWEs
3tIVl4HW+QtMzHYwEwSd5s8/ISjlgGqATxWTYGdfzbLkx5EDYFFamPQhCTXlEsKq
m2Hvyd02Ejdunpe5Q/XRhc6u/4HLZrNvlc/oVGErgSnuj4j+G4MJcPu147VJ5VL6
6jzNz+Nx7xmFUoFBoqYWWn8jzPXR7xzqNJUEDbL0X+zeKD5pmi6AzCVwwyxG34r6
Ou/YU8ItqsyrooUeBUbWmpxigg6fhVODiMJV3k8D8kCxD+wzj6d6NpjMRCg1oVUA
MnSBJvom7pkkhaStU9BgRURgdNlG/2adqgudMxPB9R2iwdqY4vuAaETvy7zFNfTw
IW83rpSWTxbZz7t2n61/L+mZEauQ/bCU8oU2me8muI8BIlvaLCvgFS8ALu0fHojP
nYwchJSOlYKPC+XYm5LWIG0aQRE+/HGoL6+706xVkmlUmbbDAMTPlY1iPcS+LKFb
2wyiOrmsg6NG0QYPySzodGhj/qnKWA2kOFOae4arubdnWVcRWWyjwepuzxS5N5P3
2jGi9JIWAHVVPHpmBHrXKIL+m6iJj10LKZo6dQuBBWYEaWme/ofZqv9dLeMNKeAA
SyND9nGSBkxxKhUBr+FlhhYnZ1OLnXOcrcNv1mS5dOxQJ0v0sCZMfNJ/pDRuD1GR
qx1RPVsk3LwVJ3J5fFXlJqlDfW5IlifdkKBnrEt67LGXNl6s/bg6mHx66BwUiVCC
m7qxFpcLtP0Mo4OzrfGYiVT72h7JdwsVSKDG2+qyMIWsK/4EghsFOL3i6nptmh1m
FCuV8XTrY8k/WLJskbI2nx2z14XZuiD01bnGJVLCrH7Xd799HBgyEcO2UlDv3MNV
kkIXgfPHOrKyBzPvbiX/F8y2uWP8vUhM6K0ovTfQygSgGQ/r58KdGLtUpbqOEJG2
NkZZk6wBxXAvh0Nt4V/fia21DJyQummjWJSpx0XXSGRkMdoTeahEgS5uT2xnvvn7
KzpFGEztc5lfvihdbhU1/6OkdvI/2z6iPYWYf0qx8iT7we0ZWG22AlclTgAKxrH8
br+iwrP7nriULi/l5hMzjas9Oo4h5XLC1830K+HDA3WV+T+Ad3WlXAtNpDQiMnB/
LPipSXKLNriEmYE2cqIC081UTUml09bwRkZldGeZ+yDvpHhNMK8DOz/BhKTU/Xrz
6uv9D9HsIpOAVVZUBNBK2S6BXWod+ZN7NsFmEW+zMiHDOFVbcVmVQABAMk5W2zHt
L3WgmnUkutxt8UlyYRFolLoADut/yH4daxkSrC/BTulPZ6NNbJ6bk6zcaLfU4pic
yKV9mmUt+lr5HAB1KLnrAJb3NkI+2K+6H7S30kHsWyxgjrYjrYu/z9tQnFF/1UOv
xT/fwqJNXBvCqJonYD/oWdybV/nM4bxHKFMMomGBS7jP8u2HZmVvH/aW/VPMQygA
9brPZeNTmLRQbbP1jiET0avdn9HuL/GSYdNOcHQBx2PVAUV5JniHYElsbQh6zGYj
Abvoi02kF8s0O3uu+mPkIFX4+/tflwDXsBQp8pOFLSAa5MtE4GvYFNNiVdJjhJ6X
KeI3qquFQNTfcG2mv+XDYxC70Hv2PhhCywxSkbjqgnMGFFSfwi/nDUG3DrtvQLAs
8MWoa433Eqim9xFMGbiRM4b1Q1gNOE38R/M3dA6Tszil6uA2uFbvx3AI416T6zan
fIGHuvRDrRN6982GxjNM5au/9xPM3cb7bR7WdjZu4vR6xqEJcc4UubaIyALHxTgk
HDR/B7KP09ILKZlrlaIAU7uzJ7p6lK1PgazhrjWoIMabCn0yFGyib5EMdva3kyQM
EHyeenPoj879RMPhLVqhtYbzXDfaDN+oSI0kTaWcaIE02StKhYASyDAEB0nS7OhZ
CE5aIqrWCQ46UOAm1XcOtzIe/xu+6phEEIjmfJ4ip/VJxQVwyPPNE25+/I1+5Tom
DRtIy/q8wprXR80K7e2gKmTeYnduBawY5cTMyK5F3fojkg4lR71SB21TzMNOjoa+
fNCnX2Q75+wbILdAuyFt4vSRNxlLP6rXnhgzGA9E2yCAzbCB/5TbwrkspOSspae6
HKG70v0srJUBWnMKHVhbyF3SxJsAtNf64IGAnsa3qOfpZlW5kL8cTEWsYLcGbx0Z
H7ldWfON47UNdi5aoAdBlAHVdp5JNUtxyfF7vSfObq7Fv8Qm350eXnNLBeMOKVUC
7gJ7Fj3qhAT7yu3nbLs67zxdfdNhi78lBfWH9qX4pK32DusUzgitt/G8qhbzBHCd
rj1iiivthtrfQathlcf3XNmYGw3fjywunz8f3KdNekrW5xYZGsi64wMlHv6RL5r9
DIDxYoqJiUf3wSTtf+lDBvMfv7dkES09PvmArgX//237+tuWg/zgbVIHed/pYWC3
rmsnKzZOftbv6afscpNwlJklEccAlMcHdLZ3UxcKgoZeWk+qx0UQmMRTXckjj930
lJCoXLZXAbb9ICUAa7T62nCf0f56azVen2sx9gMFz6C7D5hMU+dkSaiT6peorue/
aX2UuyMjDVI6a8iFS7TSVpAIixCcwUcfJ7Y2vjuf0giINXSwHoZxdzVWow+pfsbk
HEcgqOwlDZt8xswmUvQavtHfpULaOZBIJOtitifl8gUt/COyzr20kaNa2uQ9+Fm5
wLVBLrr3O6Nf19jj1inO6Eg1Ho7wEwbELaqWYaJZ3s2kZMLYNf0tBdzbgZqW4u1T
lbHEC2lkwB02JElP43f3/AjDdoSiRKqDJXtuQRWU0VI+YeRBbwIwh4b63PBhTOd6
74pe79e0zSlRkrkWw1Tnoc0jjfgNw66DnRSJGtrCNn9ZNfFCoWgowJhTikprRBiy
VNHrSRo+53RLtuBz/b+3HxWoQWNMMocY9v0LNN9owkcXYBPYODfbIWUWVV8zHkRV
ct2/l9fsxcS2dCb3CaoX8rSM5m7EXyTOo4okiIrEu3gVlMPffyPy5kVsdq0eopU+
oSmX7BkmVN+YdtNbz08gMvH5s4cwoPKdLbMHYAZsmu9FLCibccKH+dUX8FAYHl/Q
Y3KIqP5KUHeFfEBmlShsEbzF2dNAIVNElFuakrBpXg/qRqeV4jddARPykyUMNxzl
yHhAcIrTUlFInMFh5blia8V9FUHpVQ/LzLOQwI/XYCEg3Kcflh3yj/uSE2WmNlsC
oHjb6NTODJWWNvNfKTl3fZzfTe1R9Ei6mK4jiH7o70SpuU2xdp/wEtCMW4x9LXvT
XLB72qIoQhVw+CrcdEU5lS+gFh1bo3YF88zmd+xzQyqykln/GDxF48ZmfNCGm4co
mn7JNM/3vCdtlLm+p609EJhNmptBYsiNsya8Hw3/x54mRxjdk0wRPn8xaADOeThu
+LoZPItcSyaGWg/qV8kN2Q/gWI/URDgIUYtAxTHR0DVZHTlJiyGHcbgkFtJZEi2o
Pid0KhoS3G6l5clXJa4YMlPTTVX5PaAjtI7fTtQM42tPnwXHTY2n2UIN9uou7oXn
1NS5SZ2e58uOIHUzGJrNAm80arGA2M2mowM9ghAbVGkbDIRfbdFkFhk3pnfWBHpt
jrUHfUM5OgT6+PJAjyUjqZZKQMOvUtSfW1RS2dIw/vEMPRk3Q6w8DArkS+G4IIXj
+F2+Y55VUYT4tUlzjg8wkXVT6Xf4evnB1+bZerv++OhRnElosWDIIzeHrnqz1Fjb
61CN1m4EDkCwaboncZJORxE+vMkPZ1TWDr1wNaOp7GKS0QnO26yIOQPK6OxxzQJ4
mEm66GAo9YsMxSVJ7pZOrXwq+jiEHp8DMnYDyyXkTAYhTqkT2Lx0cmyrX5XQm/AT
EL3eaDCSxGhTLisYUQ3GbQvsce2foLVVSgMsEM+XK7uMXsKx26By356XqGprmHfB
J6oLMS/FaJk9KTyD8MgzrahPHr96OKGDHkWg6chWpb+yG+E3fGxTveq/tioqWAuw
We/KzjEq1HRxsdtzXuLCegtMPIbAV6bdpid/MpRw2j+cIUc/oeVNGtwPgKLFM//a
1PEAos0CLDgkFwUeQCh722V13x8JJfYHxGaREXlCu/dA4B2YunxU3A+5vpeXTlw0
pO+bSP/ih80GQGql/eambGVzpz3JGQlKL+JsTBiJtA1VtPYeOEZx+I7tmZiHSFQI
ESe9LbxE1juF4Tz/I79QBhoPsO/WSRPbsLPJ7PECROxoAfrn6QvSACj2cS2wru1A
7Utv2AxnqpG0ns/ybG88LfrnkX3uKWUCCMd2N7Y93tvF9lNS/BPAyHRn2p4tf0Zk
/2o204gdqlsEGpEQminpucpDzp8F8qssXLrqAzfMtR2JezfImaKCpaDiBapnONPe
1cU0VCsNRmrcADjqn7dxQR1Yz516pr+DV9DRiVZ1mr7o2f/i+JGrxoN6Y7IzjfyA
vWPtstJH1C1bfpMqauPrQmhTOEdPlnYPLuy2Hrqkc1uS68NO28WK+OmFUSmH4SJj
bYA1/eP/rV/tx7aSkUknxL3yNjN2j3pe5b399wjTy2eRdIpg9xHG1gRu3nTMG/gY
BXp31vGNAKzQ4U9Y5ktNVqwbv09AoswppwWPhqcUqdU8KHA3uTNq83zn0ksdqnIH
LOiU/eEaN3Wi2gqRQr3RL1VVZnYhNU0baxYeYpJA2RiaWTfUpjc6UPkja4wW141V
vK4t85kq98mB1jK7zA2PYjGF8Pk6slCtMiTvCoHtsKmTZOtvEBuaVdc6vlcqhnWQ
uOfO695USeecHuqofcA4qMVlkLTx2ztXB4ZVpHj+104Ugaa1OAi1c63fxp2iYlqR
PIp5hnrF1gaOZy8nB2+93WvmsburSVarRcPxvR2/mbfN9ioIIsiGJZs5fPHUCHDq
+OkqQkGjqtB7zLWgyVVAl57X6kb3UV5b/+s8dyReKOFYvFSLri1WLnBDX9tbX3bf
i7lYDfatIwUS5KGpKHl+6Pw+1K13pNa+9wNPMLTGPYOgai4TrjUa6B2U1u71s5xQ
tjFTRBD5+pl3z6DrqIAkxKGsfbDBWdr6mIlfDtLUIX5avEpmAVGmM2zBak5DO1Up
z9oX6H6Ud6AftuPApAibWaZ8QUftd3GHHbTGd2DdI2NoZ/HZBm21MJvDzKDWXhL5
aliRiaQtlYhpXxMZ7CO93pcDJG8Fq+2eazhkgi195tLYCivUswJjtP0GoM3Dlcuf
0hr09Tv4DhVd0jgg+6oIxa9QVRGXUrRSjFU7jYoZISNY5yxxu9VDr2vJuLWEQCfe
RPm9hLoNz5XG8H4wtmMcI5RYZiOey3xdZ585zlKGMbnf9bvD3VwEL/ACFHht9hBE
3zsBMLxg6EOHVExHwzgBo3ZTX8QmkN8pkbyE3KcdmunHNktlDcAsdiIXmQKZf/OB
RVvcMJnVChhdTDn492WL1kxeplBrzHdcJgMf+RqpK5OiaZbFj+eqsLZUA0WK/k6e
v0j/Uc9l5oJ55HxdatxRKPfgI8jUFuX02oNyzrkgbFPcqwohdkEDG535J/2JpT6F
K3l2vRLJL7bafC41PJLgu/w2983pNJLem2Frz5xk0vn260qHJXoa/tODCkhbT+wn
wu9ucPVdnnLtO7RmQ9ZoLCkqWF0Gs2XLxEpyDKcDC/vm+gu0yVel/2YAAwZcztq5
BUyTOpg/IJL3zy9MziAv6sMG70m4QHSC9oDHtyabqDQFC/uINtlLMLY73jK1SViC
eodz6wGSTeys7sxj5g3S26pLFedtu3aka/ufD5vbNxG4DDw+w1ps80RxeypZFJ77
Q6wWTBopF0R8CmPBo0Y4vD/BxllbEXfccUn9117kpsmFGoRNGNGGokwKs5FJadCK
UZAoby13BGhkWoRjZYM/ZTOlMMfU7N/e1ckj+Uu5NGB58ruvA6b8br05ljfaY4u+
RrBxje57T+IKE/PSkYBqOUOHNkbO1WdHHG8Hiezl9soCGriNg12CriDT/qRPwyXW
8tv4CXiCHYoJJYZZH4zq3lON6mwX8wJJhiomwWjk3Pse6VaBRJZANGSG7LaNwb6r
HGMRHW54cjAr1Ssb7QOWOANBL6rbTZFgYCmA+kskQ98Wqsd8QoGRzweORtvUdBPw
FdzmXYcx0/yMfvw8Eq1tCY19M+Ndz4tDRjfxOn1ht6mXargvmzwhvoOKZh8hgGDt
afk+8iL8K+XW9t4UqHXH8yrxXLgkjnz6s0Q/SO/Q+sogcMB+ewHjYR3WmWQpqQxU
n68S3wtrADs2okJZBvMs93FhvvLZXh/NMhkOE+rOP9N/mVzWSY1RJWQjEMJbSHdD
06UBVloUcZB1kcDE0A/pH/z5Hmp26Ic1Ftq2Dymnm1Sg5HzKd8tjxZrMt2atOOaB
UigbvPbaZG1ZYIzh4Hb6Q5lJEL+gU4I0P9qmi5ZicjqI4aNBYEFOX9AZ/sK6Xmh7
RpE3aYBh1HrqUcdcyJUf9y93wJrT+gjH2VA0ArDR0qGIdeRNwrQlZ9Yp+kBuglxp
tgJaqF8aGScXkYww+TjkmlcUzhMW+jhtOn36jJwy+tWwzfceC9Ref9xfbaOl2obZ
1bMtozLD6NMB0VgqhdU1a41jHdTItOuOHDPw3YiJ3CdosIm4kUYB7bU8q0pvfA12
7u8iPrFYXs4jIdMbmjGGsE1jXpueo6Myps2flg4F/FwiZj5meXCXyoaMQeBfXN1S
FEziEjkG3o2pQ/zA9WmmEusdmlh3jMFC5jk9NsQOCL4g0Ycwdv67pekXPnE1jKHZ
p1WkQVCIVK0zRUN4gaMHzyBotak0JTePgqcI6NUzcNds4GGWzzIRnsTczHEd+4Q6
IF0rWgTUZpYgl4nXh/xzDHBNkCBL6q3vv81MhhDiGXznfaEWRj42LHb0TL/JUBy7
CnUVepwzxM1rBJmh+B3v3fWl+VThuxUW6p0mjIYKwMfDmDeXSWHTcXZkP066tmwk
iubsJnCxO/SNS4qAJFYNS6lDXI1BZ+dhTEp2kJKhkr65AjNzycnoplhjO+JqAcpK
oHN5+ALXYRmFJvS391dO6R+Xczf2gVlgo8t7N+eyOA5ybH9/gnpFrccUQkBUTUBy
7CWkStvv0MPpeYYSjAYaTk627OkbniTcyIh5j7d1a4RZhtPkFnZKpUMVkTbfyW9p
uM8Km2bK2skregRUS9WcGWugFVuX0eUaEZt1nTxvgoOlvsYhtYGn795uxBRtTb5w
MBhTRArwVfqM93dGMdSmuNH6Q26VR9UzX9pFKnyJyZn+GKnlBySI3K0xoa8Vrdke
jDarY2FKcGXlJ4SbozWvU3ONlnhjGZKnV8RSd9TN1sY1fTLiY7PLp88AWYUxi/A6
rSlWCwRIK7Vo/znxU8R9ljISF9I2PGnmYqOPksosJXFBoHQGiMas4MNb53tNj74U
RuuD8ESEnNQQCWy5gH7mHDx+v9s0mloYGYzhw/oWYaOgBPO8GRZCxKUMu+9VP2RF
twfRJmX220tuwrS/L66DepGM7aN8xScIs5xhM/OfMrLFVafjdnnSUxwfNFClrPsg
SWZMWZhHtU4kY4nhBD2Cn4fPPSCUhNipxchLY+smlUde/v22H3SVyX5DH9K3yJ3y
NKfBPwgHTcEJpk4YngS6XpumfGUruHe3ABhN6niARiVuGvIpmRyLUb/fab9eYsAw
xn4PqBqX4fo28AM+YgVWILaYVsICVU0K1qT+Q+AP3zUZOhF2S1mqu3s5HsjHv24t
V+1o3zjQ6lmlhWT8TZ39Ii8xJ/af3kEGwPKpKMo7or7PM2684tSKnEy2awkfR1jV
UIAFfL/JSSL3m/3sh45dKoDb4GHa3NkEa1soMY0ssTsyxHS7JAe4ZGsGGcxN2hl1
gr5qf6EjONi98DvAlfHA0/+N4RSW8c+tl2DzriHJt6UoR4EsJs0O1smRbNGueINx
VRmfTqiqMPacFJmkVPCmKr6gwNjzpmhl5zj+yUk+LXrxEORETCbB5EAqedn6ubUC
eocPBfz8/DAsQ9xJQlTLEuFdsNldFXvPykgo8ELPT2aIU9jIjlb+mXqM6zUCLa0b
VXE0LbwWskC8O16xL2cZJJlE00VoFBV5guI1t5cz+ecnJ9H+XT4e97OVNkw4apAd
zoMJRxrATFsqRI+PoIJyljC6oy44dKxTuLrEQDfHLalZAHGiwgxf4y1fnfDIxz1o
t+5I3VN22+11mmJvgRtFpg06l9J87JwMh5Zm1oEoIaPB5KNT+FzHVEALmO+1p3FP
KdGdr0LotrAUdijAxR3ZaN7tAKj2B+wSMdX8beUb564ZQKABs1wBfJ+/ntzJJERF
nh7RG/994OsQHbAmG0p5bBqwu9aSBkynrfbifl80ako5z2iKo2hPXbvjkErFnAMd
Eag/iz2ZMeoEN8g0lLk0Ow9r8DDZaq7uBjIH8CTsgRMJ6GZcMMXg3+ngRnoQ2qQi
FL9khFyxzG6XzvHsW/pzLeQ9cbiOMIYKyOPfWYrjrqeT8M9ClanYL0u/ddtC+vta
8uG+ERe0Y59zJTZPG8tBszOXh6U+g69/KhJbcSUPoDnsy10w2Ri/L8Xuh2/9JOaR
+TcTkvPizn1d4yIVGmwKHlyNz5HunX7vANVtAlTToXtCduqd/uYxv2+HoNeowmU7
JA6h6tgBXojBrsGb8zxzFaGEoaXcG95t4xbeFGN0PWpZvbd/o5yKOg1yD526aqIH
9KMK4kcVOaAhkMC54oi4/VX32oHTuBrpDUG1tPK4zXLUTnsklXWouLfpw2tbFFDW
7mVtPeG0zBF9oHb96fldy1afp9omB95lt7EAmcZTcNkh4nIqkCpkerGzwExDBDq2
nw3tF1+9mQxmpj4gsnzJNSbtebtISXruZe1tv6wDkuiNbH2dYxrBmVCveI2jvOqT
tg9r7iPZCibjuB3kVbffo1aRlRn0k8lTtMGIDW3ErSzmBFNMHmc2AamAkg8NCkzO
0LhwTa6whSCA1XLRbRikK6rgeAHZdfwpdmfEF7h1+Vxaup0pDUIkoLFZEv+W+bcI
/g7iK4tc2+p8SFujsTg9aUlOxBDhTu67dY4sw1gxzJknRBxJRHIY3Dq73bxTnuXv
wLBCl7dS2MmujFTTLvn0Y4KqfgOlriuVBygFQioAhXy2TENBoR8DZJk0ZdysGEvu
5BvjNBN4PQMpYPdcKLLafYEMZAiOOisO1CSAHJ+6akTI64Aj9amRkQ7JSz7KQ5NS
uHLFBZYCQJXB+v8zQDla5B9DtqZHlE4xVYvsP8l4rscKKEtHImZOtw66cQ0A/CXT
9hU6DNnxchPY72kmgqRDaKKYYGRWwwc8vJsOTSAaaZITw2/N6LE1WiVIAzKST/Gf
zSNBRUA0EcZWFu5FX99fXrKVMS+SXsIn/UmDMPLB6BwaBK0UqURJVjuae5FkqMG1
vqitqUhxljzMnMUAfBUkZDvUuKoZlf/N13pwJwqpZyKMi4IelylLwAMM7npcliGH
S9DD1FyeGV/jcYfTM2sv8FIxtTAukptnFtbCL11bedKnCSeENnBM0JxePb1HxwZM
yqnJNU7X8UFi4P2vy4F5BSyfZ6YezP5HyKPOTIaONDCbDubMPNslJQbqc14rpWFN
sBafT5fjIO3pUVva+tVbybm2SCLpXRyR+23ihvjvIoQ4ZNfZkTnTb33jShl2nI9b
GX9ifpDQUiYQEOl+1qXhRnBEJAbjJfsC+8rMo9OVpdnxSTpsyHFqXe1rlgU8F5YE
mKraogRvRjOem3lzp3qsivllRvA/o+JHg+zZa3mjtIPJwZP60Ps1gsstQjwmYBUj
EeRrlGNMV1T3/k1KGLbXFJHNwMKLyb7tDD5LRtYD9GGcm4URFeXq99GFwkUO9YTl
zX2B/QUa/mkeB122g50McVJA0E1WEkoiqavMd55ojQPFGol+buTlYgGRZdgdWOH1
5vyiAKWMsH7Dvdrp+h66L5tvz05Bxu6YNt8M4bufabi5hXPe70p3rS5zlb11AZYG
7Bt+hWgXqLYtu0oL9Hsj/jLJDemUyL0PvUmbZjdgaUC93gxYrTmEfZgL7TIDUav/
BirI2JmFeVPhiKw5bpz5sPFImUBY+UoeoV+ySxxim8Ye2mJqVUs8JhCRqkygPlOT
8oxZbobbsUiQtK9eQ+u6sBxTjrVtJI1dLruzo8hmWDptotJNtcjCXpd+4xaGF961
Es9J7eDpmX5vacCHcSyItqbn4PiidS8dNc8ZyR+K3sz5hf/eOqy65SGik/9W5N0d
gLPNc9ZpkEK/SO+YBwoE0fczBeMh6FpZdGvQfoX1CsuBEF/25gWYeu6Hn7841WcB
y6ISGLqT9nH2e1QQzdHG5bonXXiefWAN0MZ8cFPB3iSRg+hFUxilTGlXOw0T56o5
jNNZs+SCsUPG/bQMvsjuJkFjaFKGdIQBkpcCd7h9x3xEtR8OTPcy9owg67A1363K
EAYSkAtFepyvu8tO1OVhDJgs0gCFfMMbZSzqDyC/YkrafW7+wIsKVlxyLjrQFi6y
gQ2wXIBKbJCs9AvVlDi1jrRUjRJ50dqRi84tghihBlrCWDSAGJe7fdQpQmm19O5R
S2UraYKMA1jKTEO3+ekrRM5qL8fTIqaGTKEM9Zi0wHDTCwgUSwjEMLAKcttcJvqQ
OjiQeBaavIQ9pmx057OHSK/8QuWLOl6SQS0Pmf1Vln05GGKdgqcviJkLRKJ+8mZA
blvXuK8XTMFnbxjV27RVB+m5r0dVWooI/DWZeCqxP36iRhyWV/CkMj96I4NCdmXi
i+qwfcAsyZj9AhHYhvVD0V6yjuxx8habjxL/gF2TaaSfi/zmXRSul+4179s2O+bj
buzR9ypmcgy3QTOn1dTDopSjDiFotyfR0Apol88iO6IhKYTVgRaZx5B6eDanSBjB
BypEUryeNHF+tQacIIqSU4JFqTAc+RI3r58pLYKDwcaRGvSdUsYxOhbpVvK+cyMk
TBDZYwJm1Unp5b6D/sKUNWvF3f90ixZ21zs2eT0D9BOa1Gq7mFBkASlde4I0VlF2
U06UknxKKGtPc4nkv3LmwmWXrMcenEciHbz8JGTED4e6dY1JPHNbmF+zvMABSGc+
c+88q3sDWYLGpTESvTgt5e6apJASKxXMuz2B+7MCdYdU4DYft3u8lVUmdyyZJEVD
95x3iSylN7XR0frU7BYF63+WDz09dKATskUIiVm+E6x+GSqvzsVXFShwA+emW/g0
g+LIpnQwKcbppDkVGVTH7vdUTuGU6N4B9xHppyZjMntPV6v3KxelylFfSmtJ7UrI
c1bugG2DjeL664xfHi0s5XRua+GCpk5Hq8EeXNKoOuiMBghwtv21v9GUbDdXt9Lr
hy0V+UxvNYVp5kvJ4x98rD1WfN51nlgZu6XHBLP1mOr96PFjGm6/Us+CHLQxXHPQ
2b31eLnQHAxwlKWnFweyX1dppEe5cK86pxTs+6wyGGNydErHItKJKHdTTJrVEXm6
WiWqvpuagrJEXfGnLDVLeLX3gp+57RCn8b3qyVe8CqnSvpC0GXWM9In6uIxHf0pD
3h+j6qzuFxGz7kWW3i0A6INwL34HE+wsdgcs9RvxS20i78ZYdKLb/+DDcuKRc5lp
eKuyZqkWLFvj75k26IZ/fb9aPYI2MpqFHStBfqQahS7xph1XGNxKZd5wcYjfD4UY
rjU8McelfKSSa6J/9lOqEoWc57czjwBnBuaQlz+NQggbv5hqWCyux5oiTSEpU2sj
kFWsrAYQrGvVYbkqqULOQLDoz0wXYZ1NXkFjMSxq8bL1iM6ow+SIYdHepvd4rube
lZcqFJyLmiaDvssu1uGbDMRZJkbs5TZyTDX1BplQMHbRa9zufp9Tz3iJmMRyvVmb
7Q3iSlha28HCPogqLbs8paFU+JIQSDm+iD7zK9DkwmbA25nUrm6WcGlXsCWWBbbb
ws6fSnGk1dHSZaq+JeEi1FxJM1pE+mfxQYYW2Wk8UwmO0V5xVg7SRO8Ms/0RBAhm
TCRjQLqulj4nQhSUJOL3LigABtOcBwrmsMp247ixEmZeLtfOfnNLm/PX1/O6ydAn
+kNd6F6qAPcFY6BxzfHkQUkwMf4vfdOS5nkKlqfCLdmZCjGfLWCG1uVvW0EL6OjD
4hsIaxOmHa4W+5Up8gWnP5COaD6YU/+wFqrYW38ZWaHqiLDLqZRj4NL9mpanTN0p
iQk/km6OhmzFoLmsSJEENufSH07ExzNtad3vmwxtPhTYnbkCmOmdVmbDdBC8jwfP
Ck0T83u2X8XHtc00U67KfruifEwZouCHRxJ+t0vPfAjB4+S3SSFgrMvnxJYztwOq
PYN1l3KhtHrr9StWqBBm1UOwVVhfxBAbJemdq+EUd6MCk42bNCPUAiUI3bHUHXzn
8fBNWzTWWp3Elq0QjtnDTbTVgXYl4zSXbeRyz2cGz0lnMyRrKr3V74egru6Qmbl6
BmQArwulf5qCUGN2Cj6U9U/bOUj0Fei4iKEa6WUjVCUTEi0MN/8+Cc0/ZF+xQ1FF
9pbohfrtdZLXX668Xyf59jSmDw2YzU7gKHWApNDrZxBdb+V6zIp+AxQ7aQuw8Hpp
DnVXIQdQc8dSpB1+VapCxEFk/7iVqVTadIVwWdcvPgQfe+4/+1kT63YjCwnzMqBy
iF5uxmvTrh3JQrKVyigTtF5E/YqIPVlKS2Wqq0BPeRjNa2zwK3jLzvFvrx3QoAaU
r8v4fnoyqpxV3qe+yDSstFiAD2rQuvC5fyO4Mf5TvQUma0gLPB6wvpR68DaNJwGB
tmB2bhZf23ZkHjhLDdLE0D4TH2qJZwuX2DzL1co/WlugpLcOiweVip1CgkW9w+6E
q9k/6v0XwRZfbE/AQFpX0dWe2H1ED/i1A3qnhq34Irr84PLJM9jNTORhT7r/g52u
HtwYhmFk4xQh0+R4liyWxsP51YJLXzOJeYHKA0sPQJ+C9WI5+9LaIUWrGS50/k9b
py8y3zsASDtu6pLYEzOamGyX5p2tNj7a+dMwoxGKRml/NBDC/5PfhVdynS36vgDz
/BulxBhxi1ExSmAH8EorvgSHdiPoop83VMMkUzrZh+h6G/eZoz22+gMICE2Ro2fU
+B6gCHaxZGTx2Bk3VNqgnxbwEPgPBvCx6X/A4ZzVDk+FzNi8BHegneE4A8Ew1Zlo
95lTre7znTrlzmrSRZpeunvm2WL7rgzBu2Hl7bNqlf0CghwqGbAFo8shlBh12dBc
ceZxPUO6O9h5Cn7ZWmlx2HKN7XoQzddcz7bXfLTDAvg5FuSHLgh7R062uZ1Oa6DT
7cEnNCvpDr5EaxyfeB8FRa09TJSbv/H5IInGi6/gyZ+xHdxaZxozlyTNtRhL2qW7
cnCrqEPchKImBk18e2I3hbEVd+7X/5E9cVxPolgX0wTxAI6MBNS5ogVyqkK9i1y3
m6omm0Yo77fblMgEjPCRjdqpCsa67SIJ6dZt7Y7TbD15am23SJMU0uCiyN404UN2
1D9O5odJ27d6u8mEoDCZL2EK/7G4KypOcvf+YAGdgoC00wGUq2Sub3oBP5JQvo2u
eU1GU8YGrOe5t/ATnM0jZ+zlDGPawE6n+63cFBnZrdJZ7Q8fHSClZxmQabTVCvRT
OkF0w4jjRC4HoWm6YCEQ+uji/Q8iMm2bKbYEk30ZCwvqRgIqlMDJ0SaTTwY1ykyg
8WE/1kaFPD7ET1nx2lAGQ8L4ifFHmpglQgJMffmHrDWoPTfaSFS3l3dpnscbnznB
D5jjG3Tw19gyXF8DH6dujn7nztEExV/7dVbpz8QrKSf7+XDj4qGC5Vw42s3Tz1Dk
PIc8X3rOStYf81dsR2AQNLU5PN4UiM5wtRg2AbAgoJ/Mw6bSk95r3jWI8hoke7zO
X5mab3gIDX1MEbgqt5xlnofgWFirYb1fDGaSSQX59uQ2ow0maoRFHfT9DgBgpmy5
KMDc1nzNJ7dY6W6rND5tXPZOXpNoAhbTMhaY4QE5uEQdStGvdnOp4OZbFXz4K/AK
qb5LaFqpiXfKpcVXoxME8ceOBmmOZn6b1HXHRzf7+L2+Pa6mSB+Nv8SC2FUu3Fr6
fnfcojElp3Kpklu8V1UXH12vwT2MUo5v7tX868hHsofzLwnh+jjWO4SMsX4LePDQ
XPgzuauE9qGugTZzU9SSoKVLm4AMLEWNR5xgzOdRo5iTRm0wU2RHKr3ubCsxht20
g/t4O4pYgckmMp9bozhGUPENcV9ggSy3Gpp9+uHCUCwSK5QxsVV+LtOfCUMVkM7q
b/10F7YeZcWABx0RpvOLCHtmA480UHGu5bGv2vNybbWivK7Z2IvsFdjQLllo+fKd
rA/wrNs9jA9NAAt08sRZS/D9m/nSLpd4Sok4tH/GV5qFMvUt4q4dBwqdDAd/CZ06
Mryy3D1WjY6lPF+/UGDI0+2peX4OG524iUUjRU1Nr+g0LzUFj/aAA00d6Fs3E468
97pyjw7Pb4HjGvH72yv29xWnvUFOqhMygjunfV5xXMX3aOT9GHWHZoOaM+AL8EIi
RLb7JEnkFZMQ6hwoo18ypuQywVqSx5LNeT3L3+mmb+biRKCvVZ6mNopiBn/5lHAj
vCZrkRYwl+8FhalEazOUTZBxsGdl1KZC37V6KSikxM8ouFZRujpkCBJ3NtWoiFZ/
zmij8A+TFjfsIgrxBwdUhhEpbxpDUvM55uNSUqzN3OtJ1mTMJBjO4ScvRIhOWFLX
JMpBYDF2gxqYfSIIdPRGPuz4+sWfeYTevkYLkW0Onlk05vSTqt6XV6zZWCuaX5GP
NMBtwMRxAdGwWDd6tK5DGlkCmEy+jOJtjpwM4Jc8AwuoXEhNnwDPHi9KztUsflB1
8QSTODodTpPRcSXeT6hSIJq9pEfCA+bxW/oeFpU0y6D5ZMH8SM6T4ZZjr1ZvRq8y
S36i0mbDlvRN2dYgRezxnjkc1qMKYf1a9Yy/5QRcVmwcn7DFcWIH9rRGrSIVG+yL
jxvhuno/HXiyj5DMKabtW7ouLPUpvDbrZ9TgG3qAKOQdlvyNdfiSac9zBy2GdAOn
4Y9mvW8mkantJ//BJqej0N4IpnEATRzN9e9vsr/Yrecoj6rKiyzGPcKMC5B/D1CT
I2gXxw17QKEA3ld/FKj1VmHqenNDue47Y7wZm60BMc572Dm9X6IvNpKu34SJOz7r
N1ZUIvtMSY5YPIIo6VZBoeS4PVpDhgVGs/y8/K4oc6Rj9xzv9rX0Bi4mU8qEdvxk
y/DYJyjktjlqVeHJIkojPO8vc2c7Od0sn+XonN0IvUGhlRkh/LYW2nlNTEofpLYS
h8zEYcfk+6QK2O91fHNRF2ReCTJYbnWmkZDkwlQ9lUjU900t8srJOcJoNN6mtk0K
wJ6R/FiBZilRB8QBszRXXqCAqeFWxmMJZGtXpnAl7hf5dElZSy7x8oumUtOA9mQ7
le0Mx4kBRHsIw12MlAt922cSVIwiCvWPZo0hppaFIfutHRVuVRJfLtxOlS8jAQ7E
Gmc7zx/yBXFBNUhiHGtoYLKqy6/+vosW+AlQx+hPiGDUukuzgsz/dm3nM33hm8Ka
vwrNHdCVPhTNjndDlWfyAFSY8uz/RcGxmWQOtvuSoZ6WgkPYQg3g4lAL1U1+2mi3
yLUqbB6uwk3XYFtgFPW1ksiOMVo52W3oRouckej9p0N7TZV9K/Xp6x7oxbhj79ZA
TMWTMg9JLA8vSHuiyZ2SJIy7Spnl/rN6zqWCOqMpz0EkeaRBcXYoGwLPiyiSqEBe
6vF3TQ1aJ3eBcZjQFl3frvh3NR8xlBI2Lh/VVyxlMj93h7dv77HuFrzk3jlJbKgl
Or7EVwxf7SISsSL+hds2A385LdGXHZmvEXCkobFBLILAztTRegmjtU34yTC/TCq/
0rinBCC0K4SliGlwbyPeztN6rg7axKemLQKzeXpQ7PEoLMCR8vd3LfEb4xBVdiFu
MzQJHnHqlCkX//fVE9kzLfMGnmUc9sfI9H4AjWzftdh8yrSsJTKtaMetxy33J4yX
euXV1DXp5TiUZ6whSJ2N7NXYfNWsd+MeSvYC5ZsK1nlx227d85Df3sfQq4TLSjaT
hEP78hgUZlnVL4a6RJ6Awvc3CdcbqQiiKvju4a50SDt0Ino9+35174mu6YE+yQUh
fxikJJrP4L8wkmGPfwJauVVbZ1glIvoYieB4GWPKmjPqaAdM1Yi02MeLxDUo3dmS
q+ddRob5le5xCwFKXCLj8v9cZJ5+8GBBpbWWcv6ejti7P5V0lc6zhOtfLZbnI5IX
tkamzr/7BBU+nWtDyMVEFtRULM/u/NlcgC7BZDw3HPKA/TBpK3RM3DVVjQsJveq0
Skexsgcwc57ta5Uwv7U3Nw8TtcN37ImoHwWJyAV0heWAuCAGQr7HSEcfy1T1KkN4
RMxhkOxBbXvcstOpwRu/PBSCFTmePvjtg/PGhszN3uhgd6EbHJrNWmgXafUIsyEy
mkSCEM0uslplLFyPrnduD6bVxlSWriFrdxkbflJc/pkHBXKie48WhIEgO9ZeAlgY
n4TxIfjekWByAR+4iajYsjL0uYL8B23n7FHbxr38zuToaP+tpAkBCOUNCH/eLsF3
t7CTk8yyVSmPHJDnU9x1HsyJRtfIKTAbL0RG9wJ5efe1sqw0I41o5c5BWsO5jkbo
ywsL2AWzH+s5BPfHxODpaAyVeAyUrovZe/FecQk/291+D4KXyGFRagiP4P3xrWHU
u5A6HyKc9WYPTgwMyPMBjmI1dcMCUd7XPrOa+zmWYisvL7YV236I77buKwp04tOZ
RH3p4lwNyAAPWXtw5MyRGUtXcHq0bOl/d17+C1BwJxfFXrv9n9xcfm87et16YuFW
WlD+UHVJPTeWrwZS2FV346+JKPSER/8d9lSNK0GlS8mhMin8nqHBkOixiHjhMCVw
X0ZyGES0SdRqvRTdpcpd7j/gYTrVyZPi/lmxiq73caSCBZJa/1dvzzFYLGh9DhNn
82IKwaAz5RulNFIw6kmYpKYaFSwZCsl8Od03yO9cc19IWdW+MRUXwGBer6nW5g3G
G3JjU81s0jZErFKKnbhGnkA5L/gVEpWv26RvgzJGnjc3T8hdFYFB23cu+Nc/P/zG
XqoscUmMe5gr5o/fdRljYKCHgseSEU/QSuC5Yja/FKWKG7MPfko69Y3KsmZr7s3L
N0456XiScZN9gt/gCimSPTk58CmNTkomQbSKcKvzD1YIskcOGf2NLLBmMAmU7fMR
aKYnvcm21J+Ho81+whS0Sa5gbEXvlVFKzuPAbhhtttv4HVFtFT6iVZ91BNz/hHKt
GHnwNNtxiiaQsFFOH/uhVx+ckb4CrXrjdYhRNBP8JdKNYPDhnl6FcoSxF4RSsBVb
37XEPmoT7rh2OxLP8X+QtLEMU5gdc3BCyuprqkOFee1ILMXIoaVx0EmeEwoGQxWJ
n9oxGF2xdpzTHKbgB3/z0CGtQ0Rku7pHUAVFb8D6DWrYlvIx3c6t/d2UAMCnn7BG
I8h6MA3voWZGgy+R2ljFhjo6bvJ8IuwQKZndqVqSoSdjs9UKybwN28hIM1qLuZkD
kGCq/2sDO8rv5iKGZhUJl+J8OZxZVpNFJ7xAffEvRBnWkQCxPleETg+mqfLbg+Dg
wUL6Ym5j0OEyK8D0rh6RNSNiNEGHBhTd/POXYTF82SAwQZdPWTAO71etJtetSx/m
YXblOt6ruBwqRy6y9iLwD+ANg7BvPOkezORWT49JqMvpAZ34L8iloLg/2yG1Vm9D
JTZOl/m7fM+lwHsDdIMUCAJ/cAuEuB7m9pvSUJqSWretspRd9nA+IcMKl4ErmWqn
i7uWMqDqEwUDR9nkYproSevtAzlTw6Utw5Sca9bE+cxZi4h/p80xSLDqWVC2xiHH
fLliJn9Qdbv8B4ECvY6wjkvU6iCfFhddYtZ6fp9qiu8RNQY2iGRGw5Vdc4cMWVrR
XCVVz+T8feAkDREbF41Ti6Di28q9kzEpJOGwupyXTrGYlPNagfTDK0UpmXI/oSOC
WWi37fn4+emKm2tgzPLGVTS3HSaTERCC2xKvY/v61AhOKNjcHC7xII/hhFoaet2T
b4f4wTjqnSaYWtGnlbKM+hULp62T+5pyf+KDfDUlRMh2peJpZN6mE3N04R3qSimc
muRWqWRtnebyPJ1wrbYVVw29o8cPty9uK0IecFF2PZLxdfC+LbYWsgOqQDefeDWu
IXP1D1hdKDa7mE8antiGUKYFCx9nmHsBa2GrEc0WHlcdH8GlZQoux36EViiHmLlV
LXqh2OK+k9bcvv+Gr6T42oG67S9gTeiv+hsIbE9YdUa+SHkxeEH4m95R7p2BU1k1
hA+QKCVM8Bg1ZRlkHgXxoDSGdJgXz8IHQT9ju0KQ8hz4yI/1GiQSFD9I+BJc7pK3
Y09A3NTYiryk9ndxNssvjj8mdaVeBuLuZvjnvdlZ6fdEbqfAyGvAW5r6JyHiuqop
32ZANMuF3L6Qa2IMHzjyT8iAsiy/Iz12DY2xZQDNHLWP49ljFFnOT7tbm0REiKky
65/T5tt89BPlKUkKlY52xRmVodKefrwQilTj04bBYt2BLJRyZTqgmiQ/7cPUhVy8
wL0aiQuDxyTQLRhsgJtFTgN58HRZMYoIZtldqK8yhTZbZxajkQ10tT+TiKp4X84+
3U4MXdHQaR57d9DgWXtEdk3dQdMQbFn/iQJBSVfV4LQPm8K4oJy2/THsb1BCv2ha
MH0kKE1ouZLVp5jOXPEliCof42c1ORHBxD41+XHxYOt9dEsaQW10PVT2DHiM6pRk
j1/ojgb//8duz4GqF1Rn+e2u3rXtIvfa7ULhBMSj1KUU+uFlrJl6IRa6qTsCXgdK
2T4keTSct/STGZxfuWapQQqs4Pb8WuVUGb5ePgEaWSuYOA3rdI0iEDRqC+zLpWhk
xCKCgKIOYHyLXTfiM5swT4gsWZcFstWAAm35XH24as6BcGv+QBBEG3ei6mJpsOl7
R+sR0e0za+6PGPpVqsUpC+8NkL2vnC0YYUx4kMqXiqzy7VyjMTWGHpVp7FzxUox3
qABQKzQmHsQ5Lgqj4677jWRhUb8FRGDwP8vccv72WMNxbsICQY9M1VsvP1IhbdIo
aESi3BAZPlqbt9wYqxCBhZruOvhSiBINCpUZa6xEJ4giDm/+t+uMSiRA6sl6yL1p
m4QID4bpl2lRLlcUSW2C4FBae7WSX4XIEOa3Gh0C12Jf7MXVS8SJCKHfW1MMtSML
wPWP2hoYFVfPYzdoO9j6ipzQNCq1zcMCxYb4tvo6Fu+xh5piNpHrtUEIR8Q5mBMl
9trPmow6rLovLFsTK7QiDzpli3y+mHV60s6EPoVFvXjt7od1XAICXGTfXF23ZOE1
xDyqmiijo+agN8/MFec0myD2saow0p5gpV9oI4DwruE8Vf6kE0VTanXh3U/VPxTu
8AymvadgIXLoor0KWwbXRuqXLbgJcOuodL5+MvhUYNB+GKc01HYRwiVAY2Ot2GUb
Kgo7NTvUvcpRRYtNVbUTU06MN34KGp+bqzAq6W8h4uEQ+J9ATcrURWSKBRxH4mCv
lAARspj11EAPi39ZqhaDh1cVRS/ZqoYi8SJiKo0Jgr2A2UwjfJx6YemqFoOa6Oiy
ILUPDiCBvAHyGDsFSmIknMJGuz3gpA+WAhPlq1IfHpttEbZybmZrv5Dg+S54nAnR
QRfFoU+Art+BRCrLOMZbvi5psJ0Tn+AS0TKCa0eHtGK81Bl4a4JiRBr1WxFND3n2
HlzXo4bRESXPzq+XQACG7fCbh9Ag6M4H4s73fNY8CHC8sKR7Ic8hokBWNhjesX0K
V938K3m3pjH70MMBDFLL1qkOFafbhRU14KvDZtbf4BnJtrl9qOPmKZv6xTHWIe2L
pBTjfNJP982QT0c+7Rj25sLNK4qymgmz8tVj1WsozMIctgApQhWlgnfpXNc6IwEI
54rQsO6OvfF9m/X0wsA8CLji8a3swklO5i0skObowJMXeshGGWxBcoUM1OcXRa/X
PrGO9J5Ch2i/UXSMWc1oAMfI177gpy9aYMaS0vWN9uWRwiCnKwny1x/3trLMv/2Q
5MyGw7sDi7KGOmCzGduSMimGxfqEUgSL/xBEjL2H88j0+0y9c0bII9msFZGNVmOA
gTi4Is/anGDx0WOkPp4xKRCE2NWfndNSaFxdMBuAxkheSaRiB9RCvOCIyRMP6cXp
DYeDscrNEEAPjDWao50CWoZdc32kLRoNXdlVleDbSKVMwWWLdFdKyVADHJekTwny
dUmBjbpgMOHhHU+PzmR9kKwD+MzQiUN08T2FkmgUcwl0u10yWSdxUJS3lGjjs3fW
aeoB4x2M4DiLWc5o6r9k2dFHPuSzm0JihWrZiQok0SO+J2cSijSlPfbggk5C9c7s
Guyqu6jue7TedPIzkuDsrvHo6G4WHgT50ZLJ/AKumumLlD54HyKjae7Z+m/xo6DY
Y7C55lli9dXg06RQof0RGPCzXB77Gzgp3swOr7RSrKCOf1x1Qpc1IZbi5caOE9wZ
c834pB3lEIcBG2b33Wkr6gdv1BNQkvxnDoH1FcakPowz2UjW4NUoYHgORpNcp9cz
AlOScyk9yKAtK+5qWo+8ejmLOJbLK4eH/5gGtUwh/iKsgVJox/p1/nBq/g461Yp3
cfwIv/vGONak9jQ6H+6CFSiXfgI5zXqRih7NRW1Plgi959lBa/gG5xFQA24dhGCZ
tONN6HCQ9w90m3Mho4XtKEso/8AB4wDiS5EJdk02b3JX4qtvALKD4R3B8r+3MMDd
PVt9iVcP9ryv/o5nfsIpeKs3cU608UrU8FKwiYqAagSuXJsEBv6coqKwPGbZK32R
J1EHpflU4wJoLHoz8URM7ieJtrQSfFqQzLYk1o5dWNCZmgO8fz416KvGm5NgJl6l
tqF4IBENaeGIeOwJlDJQL50k0cpUWAQqQcxg3WZtYRRtXRaj6kGW3vXW+o1P44MC
8dgd/53ZbbMNYeTeVAwNbsa4O30FE29p6VkeOARQqueRY4HYCTvCfJRaIONQ2spX
HoBP4r8/Qj2AkMTEdKxAGZq335HNmEmN8PtFyCeo3ISgnsA/AeaxsztUQk00Ae7E
tsi6jDLkhzzc9BNQ3XMxZEyVEDUtV4CRpeBFJLjFU4NvhcdLTavUnHY4fAte7Rqf
cc+mKJ0Kz8dMf5fYP9B4pwSisw4csPv572Tlbx7LSTOEfsQUMsAirut+5oiB52em
esKSsuJuj4uagqZYbsdhQ+zDgS//UaQ20GfjvOA1N0keoDJRyTXqTfVIi0c+tXBO
c2Brym26hD659UJ5WZq9HASwQP7tzUUvF2lCUfZP3LR9HGPwCQZa2bwfG792+kPE
5Q45OHF7XlxxDEtNUJB9OT2OhvqQC4QI13VecsH/yh/e/Yt+Q8J6wjVzuo5NFS84
se2nRcO3WASgEKD2UgGu/WJjuFv1/ze98m43mVoZOnMXP8gDlBsM/bJ70f8YWVYJ
5zlzWpuR0m4PiVX4chCpY7TtN72iNaZPiyyeETxZA40+87yEFqURQVrrjrft1lO5
Q1vcSG9q/RdbRalU1hCfTfs44GzPnQnAx4/lX8KsSbHKuZI0R4XaVDsYKyLKcE+W
tXFHh5BXTQT5CoENAkoMFI5tMaTMWyw7OrtUJ2+mqGIP5g08ptI5CWaw/BzuH/Am
XijMG8/CKSOzBRQzP/eefSU10n8HO0p3S/Naxa4Uub4+hgGdFiX9hgML+jsWVAyu
zlSuGsyMqEIF1ltd2Y5QoLi/d4uNzerBcbts/ahBoGV3ECA6ZbfSO09n+1F6Tppq
fi6D8DRW1rsKloAPYzvNliNP19eLnpwHj1NqoKpMxgFQORVHf3Eadt5IE1n7vjnB
rxKG9Di0RCLE0oMZjqflRkcFPyVx268ZkO8Uo7gy3V1ZDhIpSy34SH4u4JprMn/m
3Dz9RuqK1UCkrtdu2B/3b0I4lHr2myS8lvW/38o4CfI8yZtTNqHs93GoVBRKKagU
eb/tcTfTTCkgtvU+Z2wj8BPrEZ+FwIqNHKxBRD1Q9lKACCjF8KX/1AGvMfvsmf7d
GlY6mCwd05Bid3DbN9gxPkT2I7KGuEv/QdtDldushJsYlvEzl4phRNmUOQ3ncf2t
PpCunH/CRSzGxBnDRi8nbDH+BYkbkP2QJvRq6+TUL7u6M2EjiedDxc7P95o2ZAHF
UmjOzTu1PsAJZDzbl3ajyQLgRvKYmxTlFAQnddBzFODjvNMoAwZOk+GaMzJNnsfV
Uh3uvxnzgBMuWQylzDVxf9AkdlFxDhjco4ckL8CJ+fNbCZ122aV+qkdIE/5ZbzeW
T9Pn/0U2zBNv2qQ0pjRHJ+OSOxVuYp0EzkR4wMHPNegpaEM5uFURom22tOzl8RfP
8EmI8h75d+K8Ed8FlO4XiqxuzMeTt6/7NlLUE/lWW3t+SFERvk5VRSSz0qFInJTO
EcUWB9sGo2iLfxNZHiHpW06YqxW8pirzqyBJ2xV0BIdo9PocDzYKdFWDuw61xVzi
AVg/ZRBqyzLqPfNWtTsJNfZ4qDM0Rimb/5ia4IuL4WSQOvWw3NDurcK5wgr0UXkB
/KnOl+OAE4QYPzlvSIAgOw05+fkiYLiiKUxyTXzukzYp5ho2OQIJ7UArnYbVcPw7
YRvGj4Ja874V7DL/zX3XLTV8kknj9xsKje3HMDHwLM9M1J6S+z1CuS/lkr/5F030
7M0HqZU4N4yjJKiK2JArZ75qnb92VGq/+eAeEbKDeBQxINblaucpcwZKxBLt+luB
EdZRBr1cwSTW+FsA9dOEVACR6WqwD+BG8KRXhDmQKc9Qv6Ik8K5cIVg8/vw0Y69d
drnTxtymdiFuwo95cGZVKjFTb8REJhbFcegr6qiRAU0OOb+bKwSCgNj5JsPUfnJ1
IbqlnlB6MP38NAuM3jWs4lF5xlHkTda+PrMr46QT7UVIY5I47+kkqr7OzKNa08YA
7t1ZcgnEn+8UA92dCDLF0pSs4s597GaTHgpQeuec44GzXcOz7e0QqoDxjSbT+AQo
3aj+tB0llW4zqhsBgS/5/0DGJbXLX0jrwKaX0l5mquFSx87caJKLFq/G+rAluh4g
b4rYN/Z7ojfR6UqRnVMdbtZCEgss/+9xpS/2HHpa2L7SiJobgitFWDF0jBq8u6dH
cTfkMN89ylstV2SKV9+3ZUOzFkr1K2G6Q8H3o09fqAHkvMFkyHBrOQ7Hc7kIDIfU
sYvqR7en4869hAOkr6/RN9rQtOoLw/LS8FodsMAySBWLkcyYByka/I9dAdpFGg38
KEx1QGb+aQxo9TQcDKmps+r/bTXmMCQs1+hUFIB8lQqlI1gLHOgM4HTaJ2IhGFXu
AONtByzg1BmqKJml3+D7GZicDVgbdZWpEowcBruNoYlWUDhj/xEjjL/Q0X3ARqz/
Dwer7CzOKJsCw7Tcc86VOPkT1wCzXvgXwzMN3CfMN4Fsi+cvtNPct4Vf+Zh7OB2X
RPqPiqKYCSTV8zF/+rMmb5/FBrZhlLWBw6CdtdxN1P4h4v7qdmUC/wavsEzbBoFe
p7LLbQmeX16OCvwMfDm50ULYUg7jEqDcH3TGjFJsztOMYgN08z2Kmc5Jzg3ydKDs
MkqNsYgoAMbmr/Mb1yMbb3gEk2eJCo+G3sVL/LZoWR/X6Im9r9gk1PbT56dJG+/2
u7rXZMsolLVb0HU4ZpjegmBcTUw6iiLyGCcpYg6EBN8QyC0pOejrfevEa99wVHod
XDP6aDLLskji+OkW80StY0VaXF3WW6swWgfTVCKzUuHg8XkEmk6womI+5UQ61Fqz
C0INr6O4mzokCLN586sjtFM/1/3zOrUwN3vmSVIIZri0PD9rOQOjnJzvFC+jyzF3
wqrpP7KCziIAlGkJjJgUUlClyq8HcB24yKr5PI75Em5md5iQI6j5KvZGNSVowvHo
+2RsYPVKMV4AV9k3TRXI5C1ON127if/YA8oM8WfeHUYOwy4s9cF7cTGjpViSR3x0
fsF58FMvPN6GN69LmAeqO06qOMOryHMD6jXm6nkj4IqY9yks7A3PuLxzjF9r31TM
9joJ45aNT5b00YeMy3oii463rfY6pCfbX+ly05yNvHH7IrGh1X2vkWD8k/7qgIkD
Fc3TN611Qzw8MJEJgIh6OisI50vztkOn66444tIlN/h2YqT/8Vo1xORw1xKLJrza
XWCFPaWIqkiBjDCpgWtYerRwUW36p45CyPIndo/py9Usk5E+xPcQaQ3xM+IKujpW
8uRzbyPBjjFiHefvsgrMcvz5pQE9hRVGEkhspNw3/us8eYcN8QZuuSJL0Jge5EKe
rlP+P7FKvJ5e2JvmgHiJiOwkelKr1Uu6Qja6WrYEeOWHXveY9U03xcfcKQsOiTTw
uVwZ/JldW1rhI4z413cWci9jE6q9ZwqZyEVO31Z8gVxQKmE7czgzTMi3yjsDY7uA
O35bz5dKpgq/1R+Rglb5mHuhY4z+rgrIg8/K2efYRpeFrJgkN0rEp8rCzR89ypjh
16JAtCf6trJLQ27na8HhZxM1m/ok04sqjqlCmKJ+Ae3UYvX6j5dA4UMSeZzwicR9
gl2cREI/giR5I3WPb/YDIE0T5jve0hBYJ1ZnNbUBpSdqfX76mxXKqOxUvCE1oUa9
C9fpG2PA28J4hFjIh8bJXT5sj/WnUL/vMLzrbDgUBQ+epigHq2GxOyIHjTDbbn+2
yjSYrKTIJAe/HYTIJJOcg7X4rS6gIpVwbQhkC6nEbENcD5XcVJ/ygm9g1jkiIczB
AP/2kfsUwWnuRok4qaMssioy0FwAogsTMSAev/aberM5kdPIHM4rW6ZKT4jr9gCj
5PQiZAUowzB3PyneQtPrpusIV6h3Nac2qg6PolQm/+eM4/r+xd5JgNuRX4Nu2Lu9
dqCnI7QqGaZUvd4hKqkznW7a2Kd2k7w1mTRfzlTQftj16+HnnTiROsgoZoewHlZV
Px5NnxalisTot+XRjnDerVWmOkHgwyQSuE3yh3zl9klVj0NkpP5R9f+I1PsnqfWG
nybfyH65vLre6qDL53gb2AwGTHUd1u1KrGBLxZVFr2ULblXmE/d65QxERrWdLG9s
0/2HftKR5LAPNWCBcM5L4hAJ9gOVaL5rgQyHH+nG+3pAtuvoHd8/W9sPGEJcnz3g
CHrKE80Tod6UeSTqs8UPu+w376J943roHYMJgu/Mc7CHQMoD6JEjpGUxb4NQEw/9
//axsxz0w5LNYasPHihjMnD/Mobth+lNeukfDExyL8sy4C1g4dlHCsRRZPt3m+jq
3jtiUgMCgiDwZ9a+gJGFaCNi0SAZaCnkIU7LGtNyzh3nDYJ4ry38NSNeLTuh+jJy
QOc99htpc/+tw1oC6HAGgThOT8aPxcOE7BL/TV6UF1vYyHNIVxP1SmMgyQx2VM6C
UtsE9Jfh/WtnHqBBc7PyvBOIrVxXmzPn0ljPaDnEHaoAWNBz4C6fD4CDn8w/HPEy
o+x55bV4hMPu40nDFP/YA2/qlyqEvdrHS8mFEHPP33vFGSnqr5AldYFv30Q5Pe0Q
cIAjzsODGCrL7F6iTI0J7jljaX3MxN1NWowWyXDn6tjt+9y5z6VUqjv655eVMzgB
hNoMSzAbYIhXGLMvJ+X6v8gNyk/0KqzIDeklb4/chk0qoJGgglSdhwgT3zsdk7/1
x9tMt55yN32LKlcYKkyZ7vd5kC/jN491JOgukdWDIeuNFePKjB76C/qo2Io8DZZp
QLIc77vdO47mU+0R56S7ggrmNo/Y9qQf3HjRpDSDEIZBMPUqgf8J4QBesHBWSiF3
5VUSATtrzdTCk5nRKfKzw1kXwKO3JHTVNHzeTFmIupJ1l3G1G/fJyD80lojWMVwX
o3NSfA9d+qq3LU4GiXi3Q29V/7RAMNMHrf744srblWav4AYkkiNMLCVpNu2o1dkX
lMHfKj/unAMFD+X3qETxorLv/3VmFvNLiFpiEsYWbQuaT7R3jTomSO8Ij602VuGK
88mS7ZkCKujV4XIDAWO+cjY1DSjtsi4Y5gI1mAIyzFPqB/4IC57Wr3G8zlqWXvLp
d6hnEzfaiJJ68dNoawWADH/l/DH21uEmKnuRO3+LfJfBho5dK/86gnRn4BWc2V8N
TKIfTVi7KKIC/Gtd2s/u4HYO0mbep6YWJt/iBLEgR/PdoVZtfUM6gD4/WTUne7li
2MCkvdA77d9WTGOW1Ktw8al5Vw3FRxjRI/Cf4MDqMoSdkukTLzxMoCkZ8iYr3HRx
U8/xxRm2chDoU03TPTQkHt/0Lu6f1UT0et0Q8chpw9TZSI5+dP/H+kxb33COxe/5
R2cnt/fqxl/MEkP+1dOQnBSvyys8lVNTSfvgZKrTJuNhmB3/O6WoCRWgBl8/XP2H
/hwSi9da9q2WPc8SH/uhxaqtNSPWsrcjOS2AyoYiaPbb9dxINWfDuz+s/8KYQwsD
sPWuyXaaTEQlKqKAbqZ3G5sWVSb+0lhkQDDeI4nvbUEuwCe175TXVx0vLULgY4Uy
rNzCVdzxLD2G/DJYfRqM+1PLeeAuexOIfmpYFZiijSbGib3CwweNjclwiqbJc5r4
CeN1W8w4RdpEGhj1yyt077nFPnLKpVzVIaUJhgcsxlBu7QPU7Jq9z+jFlX1UBlbJ
/S25C5fdvDZ67izSAOMqCFLeIPnKLFY/4bOC+M0FI0UueRIqdniM8WWMrF3RPTw5
TMmvu53YlktHARITWJxaJ+rrm0fRYmtD0Gb8JOyBO/m5VUonYT+uqP3iXg/as0Qz
3d+dBFDKUJbYkZpmrSX6PiUZXEB9TT37kGFyXKwO3Jnl5w29L76xRT8r92ZkaoAg
sJ+n4OCpx8xsjQwyjq0lqrWOtbyy8n5/Yh509OTZDLeEkdNMILiCyHn8eXyt8F1N
Iu1iXbk5LI2VH24Og6kpqC093h08FnPTL9803AUv6in9WO/IVegio+yrrIXEqtIl
QS2zcs4ut8NReHP+UmMYKnbvA4xyZZGEJcOXsc/C+1VTsIHtjwZR/H4+ESjmBHj0
RyUEetbXSxyCEGyIucybpa8R6SvXS8557v8tiOdhGd3kWAEZ6UaNqybl1gQ1Vs63
IUrmwwf88CJ7Q59NF2zuVdityM8/g9EW34LKHYaopb7hkOmPJu6Shn1X0syv6ARe
urKB1zSrainK3S8rSYVqNX0x1aKU/p5/ZEIXGdEupYVJjvtMulx3PNI2ORp9UXma
jsktioQfu27q45O1Efcs+SiEVth6AfgvQSGFoTdXGLxgNtHAZLtRPftMydE6SoZz
o5gvfUgrb3MG9dP1NqGi4S3BgvXoF6nc21Lxq0zfk5k9Oip/Zh+ma6Dx/0lBYE59
51cm0Mi6rQDoDVvj/JdRDoizvUOwe+WkUfdOA64W8CdWtHrBDmDATsLmgUGM2Eve
5R+0sMigvjaisg4YxpXXCd5IggFmdmoLV/AV+TCT7GIEYPuA4izwwENM9pgrkwgO
Aai8P8jLc+kWW/nsAs5ebaHs5awCoGwPSB9RaZ9MCWxTyWn45ZEECdLFaj0+6oAi
tf15XilYfc5oFXJrlGS+JBMer4xdTqCbFpFmHFuvqeqyodzMpNLUH2qc8vqWj8xs
Ciy1rPjohy/H0RWp8p/kovSD+mlRBvM81pZjQjDhU7FhRgiY21VApZTNCwzoWDEG
2lpxY6y4dN+7lYu87AHVOkg85kQNf84syrf5mMOINdle7GBeCyy4Pke3kR+buukc
Ofl3YSKCC5xSab6LNtBLvs4wunO0Y8OlOQ2HgSXSXtnQs7M7Ofn8+f+n7q8Xl6xQ
E1P4ooDjjxR/Df4AdDdsSAr0uIflWOJGxJqB/ywIun4hCOffeMQV4g2Uu090na91
ReZbV5OORJeqtksa6Mo2WcyoyWOjWQ0cCghtwC9NGKSUB3r09J9lP4E327zWhOd5
p43BBdGKkVKMHppffl9eeC6vWSQlct1Dc1ltj5IWdbvpUbEbvQeWnJczam0/DcW+
o1HkrF8pm7UKk0HjRwjXj45ux9Tx1VH2Rq6fyfe2oKyAvavkXf/kzCnM+k2/ChRq
KebsO9Hnlt9CUytayfQ1ce3lt2KE8QBSaJL9PCbQsPdeAjmDpUOp/01J0PtyGK/x
1YlHUXNrEL1QnBbwZar3GQx5Ia0UnSoFd4nMNyHWmvN7AB6BNNgot8q8E8nvEKDc
URaHOlkSTY+7a1Gebb4MDftzDUPCT48oaAvFQct4cVGQw0Br9BBrD6iu/8lMDxjt
zJBMnZJee7ROAXVVvXZXQ4A+IG4OutqaGLMIX0WRg2neAcyXa70roA9I5g46qWdi
1m6ImSKTun+2m7t4Ormn2V5CWqaGvhMIJLjBg5ig64/PRKdd3zAJ1Tb9phqdkUB0
RoR3csZDFbDz/A/bhJqBqHMowbWVz62FMJv+V+Oo3W4/l1H1RUcEd353EFIpzLXy
R7gqs20St0GAfT5I8/noP+ZpTelcHzVt3owq0nWqayIxBFqIFCViQ2/VsGehSHb/
hDUxkabNSEmU36aSmspcun5/DHHtPHBnHUJp7CTW6dHDKg03oOaJrSUa3+03qJeN
M7GFHZbM71TQOMFv1cQ6z66IDI7GQKpK+HrtL2OYwluSN7O4b8acLC4iytRw7pST
Jln1x7OsFzghBfGbPEzY2d6HIVPgnDZThtciUc8ifPMrvUX5LOmeSgn4i3r5T6dJ
ZJX2vRZjaoiopzEn9IPOX8z8z4xyYAV37nug3SumBIg77XHUiw3086+w8bMhBofd
zzV+639jCAee3WuUzUt1V2ZY21RF+WZN4U6jbRaBPVWfIJTGrHJ5GY3/rn4MSO7R
BOqYdQQDnpsuqOLa3FpFMACJzI0sjMIJ67ufWBOojA4+ZRLkwCt0HO2OZgC0Snvg
00w+sjkAqiqZ45jMHhjd2PxYs8eCx23ZyTQlAmnZyCIADZOiF1YAu90u5AP5/mgd
6GbY0+weRTBdA3cAzRDVWO0OpgMWwq+izMO1zPaHznpROVb8UQPn2j4d1J2sTQjN
ICZlAg/XMj3bbq/UA44TE7GuEHUU2GEWSOXu2ERgrZnzyMKMZ3Hvmv7WOPVsM7p7
exmRI9dNq8PWuYiN35J/hhuixfeXavaZDuVUeO9wGshD7iHRTHDETBMMheaHjOY/
BMKosFzIbBXGfyazbXzl4fKfc6MOnTpTlwo4cbGYwjB5NDA5ReJvz65V/Qz0rXiQ
meLnX8rDABliMff9h9Wt1wdpVFtxu+JnLS15oH91GQ9adX4APZ/D+a2fe2i34eRN
ILl23xwjXKKkUTaNrkDc3fdjYgXjEpRXIt4bXai0Md/sGF0osEXz3mNEshsNt6Nj
mIFCIW1Dv8+7aELBCe+aBMH+g1Wj5xvxRX65b92LiU6e6Jd2lwmkelW4ii6Ko4zz
jMddNFK+zpvaDoXX3fUGJOUsINKAtp5KbFG7MXb4dCHx31t8jT3qfmW2/fiw89qh
P64keON5WSsmvlspqRE1R8nxQijJh9D5sOTuB+JPk0RXIns8T656bYXThIKenSek
z9m0h42U3glUtKUhFeyffDVNYgA2pbAxFVOW+1TsS/OXJEgDdz5v44ed1TkiGMz4
LnfKwS6Ke92e6WZRZFMO3EAJrwrmkYoBp1xWxwBStUW9oQqRZaIr10duZyQqWAkj
snNu5PgzCW/AxDUnJBi5NdXrIyxuiAy1m06mu6RbRHHBzozDH/VtBR+lvmn9TWUf
TpTpfsBUYLP3HP2Mx462dmsQHQvouGMdKsnKYzg60iNOjgtFq5Krhu2gb/oFTsZn
zHVizgMYfkXyVz7uJtPnSf4pJTrzDDYz/MLrtmNPCfalE5pZ7LllFdAFi9C25gWU
r5qrDOuneIx176yjhI7DvvZyRZXJ1tVI65YR08VrIkwH2dGBq17tYHdnmjnaPK5V
ymEQJmeTlfYrw+gevWKOGCHmvgwjPhxxsrj5fAp5T94O5nnNcH2Y86Mm8ncSVcor
LzKaFKd0Rd4hYUx5IhBSY0P9od9VVLqSDsOqUeX0vJYBI6ADKHRQ9w3kCOLO4H98
UNTFfV3+UbF/CTrH9bogCio/L1SlZSmqncDEmqVEYgmIGVfBpLO3aJqB0yM5dtBL
UDeyYy8HXf2rZB0/bA7IwZML1VQ6Z+Ie4dvZtjTY8ApTQW6JkIl0uJ1SHNe9T+Dl
WrRi73W+JH4eejPosKKwVgeaJ95QpHvmxfQtd3OoGfYNrdlG/wFS9TTN/JQUrZG8
nk0qvpFA7D/7Ei8FVeAiRywtqvkRCSLfTdStZjhy3EYmR9bWbkb8FM2zbd+Vfo3F
pWP/MD/uUAQ7c4A5p5m8HbY7OYEUzHiIVQsLKlzq8545KQMKv+JXEv4EkkfsYRLY
vngPgUEa/yamSXE1iTETUAVQzPmAyLdyH8vdp53FLQjC2YvZh6j8fj+nfpVWFCx+
Nz2ui+NSogfP6Ins5rIQmhkR3frFn/tIkNQVaZIvCbmq9p/vWEluhSpf8Bn/WRlG
DJIwGq2uBbjWV1nv/HDnUD8iO03rPePIqM5JdRy/WqX1JRdSL0fcxLUo8+2VGDDG
XQMzQTt1ZVoSkCOlQ2jxYsEz6cYr4v/vA3hjxxuotDxYmvuhBQa1DfHpC8E/SUIo
AfGGIJE+bs4OeK/ySg9QHltFG4tjqHyD6DJnYY4s3ziOoWsu5GmuxWmFfaoh/V3y
OlSLyLK2lGvyXgMhUVZlOHbXGLfoKSwucnKAnmUAuk8utj2Jtl2DVM2qlRDnvUM0
+8uin7KM2O3131/K7EoFKoHy3Ndsl/+wi5YHbjjDSS2lzl5L10RppsuM07zxVKTI
t42tLe9Vad1o1yTFHFVSEyrM7XkcgreHZcds07c7jXEybOaH2XwxA1QbaTr2OQXd
qKu+47k0GXUlQn+qbSr71g1B8Jgag5SHT6GlYs3nAj3BBhZUun4DqJtdQAD+1UTM
56fuIysqecgKBUenI4zsoxJznzJ6xh/TPdmJs6uqzMMzxxlGJY8LMjHsB+gSSu4I
l6Ab4ZG8sFpwhZO2SXFv3oqz3LHKGxMB8pV8VC5HgosG5ICA11B3BceXcs+yLrSJ
v6atV6vbYO0c2aY5kfYEM5+M25piZxsfj8CioOiUMv/DgL4WKoPOU+w7qI5/4DPu
GvZer+BtxltUzfpV14kycgPI8C4dIjnUT40ZREeRjZDSEkUoUUtQKk2Ljs5XUjaO
AVQkGucyzsjkFJ0pDuaj12lB3O2kuo3KlknocHQXelpvvEL7bvl7vYf43EA0AM24
SxOFkS5YC9jGKXAwHWnsjrM1HuORyq1CW6CvBvb/c/mHdOqLmpfLSdFW5QWzFcCL
7XvmAM6O2dCW/OV+EYUeRxuS2yKaap6XmozJ4ZobqEy9f4vcKV9LdZ6VEpnmgZVi
ydSCp7jbCmJ5rHdtJYa58yoftz6R+NTERsKtuQiOXb9xTY9DduwYPWMWNtwPvxTw
Eny5eNZ/5Y47t7ttEXi7QYD1ovgLayLNEO4RSLuEfXS2b9+cJCyXFxCpFrOioRQl
3IWk4EzFa+K086DjVWSUh143C+Enjla5I5IfIcFRJQgn9paGLmit8J2i1H8nlzgU
A5vZJ6Oq4hONPGSPil/AZ2Z+KE36LqN+rqV1ngUalwzFydCYhPyWlxEl21Z61APZ
NxUHBGUWW2lt8gv6D7nlFTBpwjo3cCZeQ9RjbQO497Lb05BsIQ52UJvyh7vVVVKo
lowOK/xpeIDWWqPpVoqedf7TChR0ZVLXfVM1mCSqx9epSdlyU0j5jSF7hJn0kUlx
DRZX8W6RPALDp7RM5wc6c3EbRDJ8WKwr1vvm5N7LHtFYniPgIXDG+I9Q+Ag2YEe9
546QmNOOFBVFXLeyBPvxJJr4uzWoqV2GrapgjVgbO+3cuPUbVlUAQUfOuuEsYfK6
zU9is1JY3bqGWgVpDKBx+cqHcH9xw0MNBar0txn2uH/7e/CrlaIY4r1W/QxFIm58
VVbWMOy4cVol7ANuP1Zx/oneJwtdNqlpmPG0UBYl2Pguk3HMpdR/11I7uJKSGLbl
8DOARrZ88L5UlEByoZcN1mnRy7lLLrJdPXsgpWPbXZtJ1qaNCd9DvHGb3+/1zGNJ
cnfyEikbxooVWd/9LOnv0ROeq74DHIxbV3BOOn6TGAoIueM0n4F4x/mkmkaf2PDl
Ng/bewYtkPKHWvqoHaw2GgD8WN3cmz7crD0llcTMtIkD/zD15opfsDTs0JpSVJDp
vXXw8nOV0/beatDuU2u3QSKDJcxmuiBGZYjcMk2PEhqoc8pD1I9QY0Z7alOsPUVQ
Mc5ejsWdQ4FnPhJh2rW2Mpxw4eV93YiaGBj1Vd6UC/KW4pugg/2Vx9YtH8WFcC4l
2PrKqt3NAT4rGnyt2UNr/C9n/s834UY7jZjFjPQvfGtiWBpGMJIz3ot62H8i5ipM
SweIDG8wyh3DblhRa883vnf4mEisj7ugmqfZnKWxlD04pLZePfvoIdqLWnDXuotz
4B2OeG1Bj9g/wL5qHPJeTHpgthYeiA8/pyRLr+q2hHmyA4ODUNtRgFqRgk8OEE5j
lstS/07rgvH22kwoi4M8+I9LydWuOwmePqRcJ5wZOhbWjXg1dNU7KzajZAeOC0hb
nbCjGizIjbuX6d0JvwKzfIaNy5yEetaBoP0tv0sXxazK2XvvIEFGblogukOvF54a
yPIM6DcSY7fzP2hcAjdVtqf6cGuAToxIYoQLsM+9cwmOlIRkaUc0m3BCLjwuHwnA
UiGXIc3OslWD1312spsn2oTFvEoNQFx/3qmC45odedzhPGcPzqVbw2OoLRnd6aSt
51NrUDYPLxuqPoM6BgmuUv+CqeLYZFvcUFobKdo1DE8eWmFC3h8kHBuIf4ttZJQV
oThOQwNyTgAbwumOXMKMR4YglgoDLmw+RBgtOzq34w93v0LDoOW1GavBgc+ftF5I
33SeaE+B3NO3Qw4JINP+ScPWg+keRD6LIFp03CdVilnpIFGl0FQA7vXqkJVUatvj
r5h0e+klNj7Xl143tIAG3F/I+M9wnb15P6MFNIBiaMZbGP77+WiYv+9fBd7Qudp7
SeYKWR1ywpH63YeNj+YXjm8v3W3S7k9rKwg9KkDeMqCMW8U5sfKXLRwpKAoa4VvK
Q4cdtez0vCzNFd2bxxsVOPeb7CqJ0EkSs/GTNf2WxGCECm2slmMbAa6qE3eEhMPp
kFHO38+RUaydF7y4uQeg23wrIMDnSe6nTOxXgq3bDuHV9oy1ZGtxuY85tz5PgQux
4mMl5HaLNjTU1RW8srzdc9d9cPTxzuT2RsGY14T656UkKt9hdwFGGHbHxB4ZLy+d
bke1RRENCqHdf8HO/Yb5GSRqXlbAKL8FQHOexKDOSPNTXF87Pj0hVKMzyJQ05RRq
OdaXCIEanb4Re1IKjk76HjG5NOeuKVYMvWsrCWf3NPLpc/v745MZOCjGT9DHHOrc
rWT+y+RtsJuJLOkLbe9Oi9Z6gEOdOdvXP2ZFOPf0gGjBf0t5UYgwS1W0fSyzAYmw
yb3XJQSYsu15YjZZkm3whM86kfp6cbsSDiENFJgc5N9ns+FuRRd41vCvnZqszz+U
/j/ot+YKUKhnCwloqIDdHPBsHwNrITG++tQwVjEltF0pRSecEPqqpNH/I370+NGi
RKZ4yP3nyKBhq3ddyUExbfSqtbJ+BBvjjI8oqDCDrRVKNn0UvTz6HbF2zARGTIBL
HhH+ij7G8ErKv9EtIztIV4X83QnjzcQqFscuJMrbm7qpXTGHfGQ8Oq1jGsHXrgtb
lAVepMlrO0godKL1m1nhK0EpjtXu6KO+mi62JTW6/qy/yKiQ0IrsjtDm7e90ia2O
qcsVrpgr+gemln0NNjIB+sJBnGpe+4AJJ6/VV3Uwd/F1OeCeTwbY6JZvVIhXxeMf
p1+Nac1aSX29u8CpeEtxEqgDPLmhz9Yq7GpkAVsonFSMiUDi7482AG6ENDJTlfK2
p4TU+HIczf1feq4+IDIiAaeca+xTUQiBasbzVF5As3M2mg5JJlmvLyakcDj5mq8j
YIn7Is90h+QMFw4Zbai2VDuJqGQd7I9Hil/LBFuLW8Zh9HhFwqe1BVpSw0GuKvxH
NOIjjWtgN3nVNXKH2L4Bjd0SgoDw8f96nHYne+jbDmaFRR1MYicVKdLGiIGgi1yi
WJwJxqtaM7+bzpRbmzRynWAwrPzUVEm8J82jRF7pRHcSDLf0eX2UJRFp73e0MS8V
oAueDNMacAV3SLzvZQbvzxKy5Jsi7h8NA3ObWWwWSO2z9UvGctmwAhocc2iIluRU
jCsPwJRvz/kOAuOpjUoqwNxK6evcAzMWtUkekUwB/eyE7DF7VwiHngqLw7P5TmCe
qqTvGQsT0vusRCyvrwCsaZOuG897sAjG4X1fEda4Us1rBgrpvmjm7x70F3awrud5
R06hUEnk5aN8hVf6XJqZoVAlqXqqYYO2vwi5XG+P/XUH+/RaVaU7eaH+UxHFX9KJ
z1gKgahcYhDaLrWi9nY1tXPnB55Wjjq91TKO5Bk/DLieDDtqe2EuuarrOjnjuQ/A
FjtI794YtfQA8IEziO28kgoaqO3EC/+MvYJ6scXREIT18lQNHgGIsum/Tii/D9oB
un9HmymssqGhM0USV17NIerQsMt9r63IRlkEHJ/88G9TfYcd5gpepW1OAw8xDqdW
ilYUDH4I0ve5GNjiN8xOi6Cz6l3rsZ1wX5Y7bnHz8xqb74k/womonW32AOjroqkx
MZxUT/GD94AiBeEcpeXXsBJavr5xOsnyuyRoBUG97u9CK+lMHR2UbSGmbn09lpHo
YoNHv3HJ9vQZHswkcj+H4LQ+XT81mgQzGTHU0QQJZ3/AY65aDMOM1xrVTgdfnpeZ
97UWyO00VYzno4gvwWXXle24voXGutYbHbE0HsvF60+sr+WqRRaqF2JmMWuZ43zO
8WnNWZVqelNc+yZ6Es13aQl1XG9+7zbapHBZmcadlSjHezrS7j/7gyYcgtgj5vJc
Pz0ihNrZUAaTH/0WB7FNvgv6lHv/OyFkZ33y48MQO5wdYUpwAep/GarAJ3I98Jwc
cc0JHd+mgCgFI+jOK612BAZHYgy26+SK1yfHj7QsJvpJqkmAZ2L9zGwe6aImVHR3
ZX7O03WATv6h0E6EQPLw7HYS1GH/rlcBkAOGiqXY6l2T12dhhPMTHvdHNNhoJufQ
sT0qSu4gaMPTCOP69unt8xPlOSbCrKwVTxsL3H2DeZeSR+v6Do/mZVAycR5s5C0w
UNWXt0gV0lWv+qOKYtJY5dHMR+ibpvIsZTE4oocqFqLo5setJQFNAjLCY6FuPiU5
RihZiR4Y4vzb3g4jr83HG1LAbdqpI/N/LE22nArFvLZFf8J+OEXYEowTeyEbb6la
MQfQRAnYEWL3J5sSuTEsUvkqhF2Tbl+Bho3v7i4DofiIG6e24c7zzLBlAMku+78h
UDwgz3FJbn0yJAhsIlqJg0hY3xTeNKzyVRWUU34K5nV4Xxel/ScWhqCEhcxwgUR7
TFpdxBMugOJZKLkiJNB/6YN5HMO8s5tImho9N8VTwVD2KKEptCe+4HfWXq8ks4jA
cGmvVO1efRUjZzcTD9OUSYQRx43j9PNJ9whjb7Y7db10h/7NJKmOhXuy24EjkBdt
cLoYML2XWvfdEO+w7LnQ2yHsB2JgrPPpMaIG4q+IA/oxRfvEPgJvHFxAg4uMesEG
L9uaHB9S3inZDoTr7/gdg76hzPFQQQJybFbL0ThsNxbahpU8dTv2YVE4TuXqqZYm
EB1iBq3he/pW78fivQXc36ld07fe1xLQoefrbh8Qd3QmKxWV64QuiaSjI7DDl5A9
fYx9NsJzW7KdnIksSeFpsx5lMwEj5oOGf2pRptpF7HysNUsJcApZj0/eM/LLH6jr
7n2+wdP48Jn49WxyH6ySw8gAX40UTJ1pYFYAAmhK7pPNH0RjcSm5PjTbnOoEJj5K
CS/XLOiT7IoPvuuo1ykBy+gn9WE//s5U8030ZF2gKOr7W6LU+pgHnvPhtOP+h9WB
k2t69uzyZg/LGrLVSE6RxthZP+vMsKUbGjvcxsd4b20/Ytiz0/vPISuupzCllHpV
hGJPPZgQWu+H4oxaQgonEXQvxFgsf1Phunr8UyvvV6d/VYFiXWIpOe/IPEsEu+xq
y0pavRydCiimkrRE2dT7c5F7icSSijCuFPqBmKAQIlp4u5OrJ6aGn+lqJlfR7Vmj
16LAGTZyv/3yPH1HOd4bQgvIzLRmyKMyq/i4POAGx+brNrKa1q0eL/6HmVXWGJCW
KrC2/AhzH/jf5YznBseIe7DcEAUu11loUvaclpvxDDvgI1zilvh902JeyKUVw+ks
EiYoQA38n9FhLo0geyL0FrA3pkYcJ+SYmo5lM4ZzOlSzmLm3gNmfAt7/xBYeDDhU
suIGdH8dAZu07VIq5dI0NNIcz4uJUQw/3MyUPfUvFz+kHe4jvSn0YQEkHdElT3sf
1QhPGDXW77nG+L2jo0F524Z9W+pZNzjnvDBbkeKSHRzYQVfpfKFIAvWehSgyS6gL
fsoCr4yhLmRjaKOpUHA1303e7BzmbFwEH73tR3ZflZjIva1UXEdsE6FebkZN8piC
g0NkjtI/eKhsiQta+hbxRSdt0M1MtifhMsbL/0vf4mrEhXQ/j2+5HxxBmhKopjcu
ToZYz1VtfVCYfaGjs/yN8BWIrSu0Nvh0X4IE4ChkIqbvth+XfvUjiKORkH8kFCcE
Dd2k1vLrpgLFWPBBQpqd9+1OayZxDfJqyFmPDCdmes1CDTXeztZ2RMVwcjGQHdna
ndsijhS63tP8HEbyF1T1lvhPVXuWkjpu0Q1okgSvl1kOmmUIt1ZYWbB+E+/DNdVJ
6mkkK3AHv48U6vMfOSVjGRiSP8p38XGDp5/JJh9VM9vW4Xe4bTQiITY+aeAMxXS8
VvKkcrKpAJ773aXK34o441d4rKTqmg0EjwFwx3JMy9QE8wTDFNCodDO0D9OqFvlM
Nh8ubjvngk2EE1qHzkr5oOwW7m9yhC75lNLxGND8EY0C162GrqMqstPAb5FxTPXU
bh8vYWy9Z/+VP3tpuHFyR7bpncWT0milSD0o7l14gt4P4GU8bWgza1mIH/TBY9xW
rWlMv+MZ24pSy66VN1kxI4VtkOsPq0sEwH/CtHnh6x+czB7u5dMiJY2W2YMJTzNC
RYelyaYW6Hv70M6tIxEcKoIVyTUekjzaLZ52I3h4X87GiEsTHBngvPUGOLTXLJnF
PFAJAZSbvZYIKMiSohK1ACtx1xqZwwEokIczjUPzhb6IZ1tlP2zTTXWs6APc/nfZ
mU9mfuqIwbvyeYN8kM2Ty8n++FRbNjK/lkFIaacvIcSQ58kj6McRr8tajHjSZwYa
OfkWOUYefWBAQ85ja9waLGxhrkzcqjBN3OFRC4H31Z/IL4CWMZtd1ZGOJdxKPVRz
jtyt5VP5GetYvHywdVFehT0q3Sl7E3Yh5D+MJtOBbvrb6UtqOx4r8IE5To1wWM8s
fAqKtU+umsg/yQUULJOGBe7VWTjZtH/JJsm6/OorYM5Reda+udlnNJy4YLDivbwz
q9GNzpDJPWE7tut9rU0rWZ9mgRo+IFJPP/7wG6+izrm9pf0L2Fkgl/L27YBSlZbJ
RDQofk9WM4b7xZoQ3OHVd7ep2sZSv8SflfKMzQKworHMMhZXglHnNruvn3DbaHhs
pt1/D0O9eitKrL8yQcinDYlkpc4Ie2GBV/IW6D5bN/0qxgRIM5vatI3QcztPpMWy
lpT2a51sc338oCKgkAlWl8RARfMwxA9mYaTmMB2r43k4FJ8Xy33o+O73oWSeq1NM
jwUfH3nREGESnZALB+VrQG7vXqMjubiPKp7KQCaqMiWdkKE8Bo8iNa9/fZmHl2Go
CQZo/k28ldQ8C5gN1UjC690nvoWWHu0+YDPyoTTmLcOxLbqtlgTHTibfkuMgcnrp
Oi+pQINo9OAmVSf4jCgIVMVaUiJA0jsE7FoStI3UvACQbEPlBUH5xjrZw6gm1aWA
jLvRm6Cgjc0ZhycnBx55KtPriAE+QMfwXdlKQYIAwg3RWm+jem3WcUZ+jsVgU1hU
S6ndULZmthGOHiWGzn3xsGjq01PL0DlbezvTKPea31nKBP2zQkMkzkYSMgagvbDd
mE3rLWIwMZYLgdG+4T3MMLsSqsCzbHRMsy2LA0PDHIXEmsVRT0hvgAvn+FbbTg28
tJi9VTmFxo94aC4j6uq2BEA+NcifvsPFfah20W3D6tRBo9e4hObkwTxTmbGJjOEy
OzaIPUagvSfUVe6W+ncsNMjJ6IQXz/UF0DUnwqGRTBXMO+Mqi4dYR8ojdYESlgB1
eoD6RgIKtf+WuI5FYKY9uguc4N3Os3kAf/MiiiYFEcAVybDa+i8Vn8fZz9xc3fp1
fEj4pKv9x35VkTQ2ZFON0KtVmJw6t4n5Y95pq7LBTkwUNVn9rMzZJ5rK2O8DixQR
M9giONCqDbx68O23nrK68qMTG8DjO/tDFxBBerc7P+ZbHl3FaHtc4sFoGvH8b9ok
7OHRr/07vzOhXtZrIFU/CSvE7dwsg2bQfQcjVqd321zzHQW9yt3PsTmUw65igWRC
Kq2sDLJRkMs00D7W+HGaFkUXSSMRpPdhfV/pEzv0pRoYHFSWOKujRj26QMd/lRpN
oX/hD2oVHXfGdOZM5EpGNaF5huKX+etyr724jUdN9rUSNGHPo0adEiLK+FKET+MJ
g+mxBsUdSHF5QXnJoqcs4HasTixK4bRG18NjaakcUratTMgnaE1RZID3rSCqRFr+
7dtGuBe8BKYG0d406lfuNIU8APB43ZnIAbBj/pmUlmsNzpLcAXVlA1aZZfTROBzx
HIqbj+/DUW5b2IdWV19em392OCOT04g9+iAmsPF8vQ3n1dTRJv7BAvWKR49nKjN+
w2Ehg6OOx/0K7MC+1RagRdQLN7OqIDcYgNgIvu5kxh7dSJ2slPIptn5Mtx2ovsm9
GVRKFyvC9wymsmtfd5mIlV1QXwtA7OxyCRCMiRDZ7T6CEj8X7UGwZTife3qiThdo
O9L7qdN6PFZMlem+JgywOV4LS+TsRZOc1GOLg1UboQVwjfUJLLZeNQwYzOSW4gI9
F40hM4rq6uj+TmolGxiqvMjKS2rxDiM4LUN4KvUCDr9A7eEGeIvKlcS7va9Z17SF
a1MZjP3cqE9o4Mcvv++UuVdurqCuJl+klqwyPJ/vcxXE2XtruzI7AmdyVvc0ovoi
p01/0Xuc994EbJpBHv75Jr8sRH7yp3TmTekWPX/hHj6eJlL5bOlIDH544gl4foMe
O+z4JdRwJ7dc/thMRF7Qd29jzHUxeB3DqXNmIzq3jqXvdzHQnvr07jWWVY23KCBS
VhCOBbvFmUf38r4Y7qOIG1/GQ1V3uXpeysxERCULSLpxLmFexl2b08ArOPUXvb09
jZtt5TQmCam5qxAwojcsn+uzKtHkzUguFbvrdldcuWvPTBR8VW1Qjp/b6tRIGvy9
icfuKFIIDyuZb/6I5DHuLq1csEuFTiuSuArFqd7NuYIULhhKyC4r6684+Xjb798l
HSH0mv5qzNMO95yhy3QEH1L/9/ywzaYD+uhg5q2DajqXgwCAK+/UOucaTP9pLqrv
sMDuVvaMcRTU2C2nfvyIBAcWDcP0LrPqTQx4u8Iv8yjvhUO3/wKtarMG8N36Rv+3
0tGsgKC4FNoph4LokVnIhl5/3VxD1iTIwoYsI7SLuJAJvWEB+7NRtZlUxHEsU0ct
4FU3YxX1iMKsIwL7fzhsE4ES6ftqkN/1aoaQ1ETTchW4UWt4OgQ//JkXmho3N+Wm
Exg2Ikc7hp6CJ3Aljj7/KR8NRWHX9A+F43ejbsHhH2pfpYyU1Y51LCk20PNu9hvb
MspYnm0Fjr69sbShnJxMhzzzZzz1uLN+I2BBLgfizx8BJsatnmUFPDGhx3F0/RVt
o2WimJ6D7YqI6MaYy/GX056CccmNV8V38DfXHYTKQxX6qk1HE6gG6zGn2V9MI/nJ
32hpy1xRsZGr32Vugsn6KpdqJ0W4TO26Tf3QHA6PgB74Rh2/042fcl8D58nKBDVu
mng1HOOKMjz7IkX+UfOihpzYTXSJIHz/n3YqNE5znrMizvN/iqvutejqpzlND3LW
gVLsnVbWEgyXfFdYL8W9kEU7xFTuJ/1BtetO1qE7IAl1SiepLu5EXQyOPhdol4We
s8x0ocAeqkAygvZIBarSjsiL2XGoj+8CotDP5L14zlxqvgmYXqZBfr/UKYXQ2WOF
ixK5ycHVq1iQDxzEAnY+3G2GZByUew3DZ7aF3TYxhMgh3Y99HYAITCBw3z3bCrMV
8KW++TNaC+1jJmWwWdsEHD4hJYLARN2iGQ/bkSK1905urxcLuQOLKI6SOmzvNpG8
J8b+oKcoJgvFmXcsiH1gRFtwHp4CkGIM1FkPZjsDw6BKnPlvoDMo2TGmq/yoi0I7
WT5+TzHHeUAd8O4GV7dcSXYJl5OOe9SlkT1qN9V5Ffekvuew2LIF8lgEg9jNeA2v
YUj9V41OzLbSSV2GVxhyS87oYAeoGQiYOM5oRXbiwZn0r/ZrdOBPswR/F/oZJU8C
/BBFJ+32dTZi021SQvkqtPEYGBsYot2anCLwRmyterpT7+qrwSC48M6osrjRA5uy
pn3uayqW868Fowd8OCnf4/Q5lqx86+lgBhH2BIz6Lqi8FRZrC09Aig+4r7dqw2ld
Iw1bOJ4+gq8DA//4vlwos6fy9A4DIqVOHBdpCEDu0B0npyS+aRPM44mPNHdd9qDt
iROkEJfjhrlfwSwwnV9BcRSL1xJaxLrqUKfcUkv7bONVLmkfjA1ldmcYyefE7IlU
VlAnEfcIPBHWAi0fFksSQ+ZJCrxDE5JcjjcPVVTPGG6VhKyFCIMkqOWbSdqi2kmO
2WAcVAGSX+VByXyciXkZfckBkybBWHcnDwvSuI7RSspVxQlCOZCWRqjriwHayYkD
HgBje14guysPWqqRvbgcTGhKMthPnvcuygCaoM9+24f16j86HbKQnCpTastzGXDI
lUWAetDKs7z4aCXTzxvlTsvEfYIloYBcWuEMvlol/qMjY1r9Bl5L5Gy8qjz/LuVj
lIbIoeEh0pPp3EyZcAu9umoqnt9qqpBIKKK9fL1DvGmoEbv4a/sI3k6QCShGKJ6I
ywvgCbyfcrV5HAPb1AfQVmWSIpSW0y81KXPpStvAIO8ebVO4Pfm7sRf4eJZqBRR/
J/WULCfPfGpSGeDLHPo+Qn2WvzW8VjiH3ZKx7gblId0etNXbZD8Peragr5AK9lig
ayvY+VSjCEAVj8osA+PVs4ZXdY2pnUaKNcsZnhIeBxA9JnnfKug6vX5R1B+eX5ev
AD4VYHpzn+G3bqDzT4RQwMO9rCePleDolQjFm4KSHb05vARJm15EH+BJm+VEg89u
lz0gYWotKoKQzjgozDHtVHhDo4DYz59Oc/PKZvcAlIpeR0lGta+365XpMzd232XQ
3NVjhaagXxdqksk0VjPDtz4aqvJG8xgar35J3zCI5njquZcVNFWyT1Y5yIOuH4XC
ha+QZInRtROEysNRu5QZuXAsJ00y20//z5oEUwBLL+x+IjuSwKXd+ioXiSOK0HD/
bu0yciuZVn65Ye2qmbYB/s4Crhb/NlGJ+JbvxUFi67iJT6cBN5BhklHKUZOoOgq5
q3t3VG2uHTUTJKJlh5B2f3XILFChjj+AN5HuL96pwEcSFx3wMKTZW/9spKITEMK/
nUz21Yy2YIMmCjeEOJ/FaE65mfmgG3R4W0+zpu8sA5OtY7DStzxyGgTmKF2zM0d9
Mbp1yVDVs4HjsjNM4lO8YsDTPSUav4cQIBZrqRR6OU1C291ctWB0K4zfN6gxMB5r
wO+utYWHVqLh5eNe3whDQTnEdVJytXY5ZUs5UmNvQSNdCsTgCb40ViNKIYUa71/e
1wJHO560YPc5iYv4OgrR6nGZffJxJjOeRj/0N1K+scl4X+w9YAC7/hC6sjsCJfQb
6P7EWfZjyC7dqQ9+zRyeMj3l5mPRxJtJWTiqv1FboA72z9hXsHrplEg+GOxOlinu
aSC0P6XEA6/mcWK7eJlSjmchUWi1+P+xV9nIHopAmNHThyy0E/5mnGXXG8RHFkys
7o7kaDecvySZ+/n14Bcd7qHmbl2A/wspe9WfVPTxU8KBIuMzNag/gtOLP6rgE8BP
CrJko7GqfgNIfM26OVh2Y1T1ArwHZNqqKs5jlGNK4NYm0+/zvjfQ7WHzL1fj1U6r
oFrc6bRx7uMNULLUB410LkkkAJmyylytMOwBqzq4G39bk/YxJOHUH1hfFO8Jqlu3
++JerheP6v1cnx/Lq3YNdRmuO+C5AfDDHignXhwqVuhiteq9XuzaZ3q57Gs6qIys
mDiD7NaZa/8/DX0ROuLYtsFOD3gKPe5gcdOKWRXD5CHK6EU4EFL6B1Gq52GoMZX5
MQRYff9NZILGAQF4idb1+yncs5HJi4s8mk613WxYUcpbIlEYAlZIxrax+bf3GcmC
8aWKFcDJvJjSZ7YjUwks73tJr/n4MqWYLYYDVf7ljrYMSkQwc0M5hxPYh7ee9XzM
KHGUOjMPl+AbswtkkXndBgGueDNDSjehjPy+O4uSxV8wZ1wiZFDp/8bFuqasoSn/
jBnNt3ruCJ5sxe6tQZChRoulJCKb7vSt0ABXzoyP4X94zx673XmmDDYNlceBOxVg
svvTnGu5y9NtS8OmN94pIn+npR/RsnC13sXXVAMyUiyWMmsJ27h4g149+358juen
SPPihgIq7H2Hb10WlF0IAyRwPezCDQHgay0rVyo8XK/3rTlnF6UF50UgBrDb7LRG
xY+JE0naYFAvkftrddlzkPAzt7dUevgkFu1X7eAB3HZHkKuY3iMbyr4e60g4MtFY
gMq4z/ogSySi2FSFL+s4nDb6usg2ZXUrdrX1upTCKmErf/vDib0dN0KYI8BDJ8Dj
7kU4WwTrgrnVW9EQY0JEo1zxyew5grJ1x63/ULHc4Vhoj96fmDxZAnlgjXS62qkq
v3NWlUWZtmxNiLd8lUfQIYKiZDVMI1huES82WwIfJnVGH0wxT/rAzRXpDpjHbIFo
TUfWu2jqSO6kGYaSkn4ptBirIOh54i6L+XZ1rbl0jFTQihSsSXwo3AoqWYaqOg65
y5CZXECsOuJz1fLAviMyR2xMl03TFD3jBAxJNAs08hVyktLUlggHmG3jyQzilYxa
n5Phdxqhz6UnR3hBXjXYLrHGRs9F//SyPRBWzWUMIQNns7r1M2/LVqr7DfSZkCLp
+AdAX2KLhAlk7x/5LkwyIEi25tK1wACBXgBnJVHQBIfxVYxdS7Oh1X4i1MsQDs7F
GRkQK4gViWiA50aAvfaO1v4qIYsX9/afym5ywX3qwGDARfvokMDlew31CgwWqxiw
h6LpirrnMfYN2mSc8ExucFUZFVTUUm6/nNPGAesYXQ64/EiO5a3XscCEZu3Vy3hD
N5EifAf7gCwhK3vGyfMnVjEH/8DvbsBDRew8XVSXTaIuU7sn1a2P51OTa8H7Xx4o
mW4ZvmBVwuLfKyisV+vg55YB/Udy8DlU/wnNYOp6iPBMFGB4Vc84ycQtXP/EyCK7
Am9WgcMrdLX0EcrxW+hpMIs5J+5ks66e1a7FhLIrbj066Pj/IhSwKFi4kuN2QgB5
6uhU8ZfxqCmLXNfUc9HAo//w/xH4vYWfftWvQMFI8INNwH+yrSqExtLKXrGHhtxa
b7r+uvGwD2QJUWdcGMKWN6v2JxkJ5IZt6nkhdGwH2Bpz9BKoI1bHAwaXYJA0/aUy
avyw9XihAlhYIJZrspUiQ3Rgb/WXtlVhzIVDQ+nsdXrqxUvcsSNQ4g6dlKQN06+6
CXSSP3Ry+/+HS6rXNboQs79b0ZOH/neuhXmsslaHuRM9LNn/l+hZaTIrqUWSj//r
FsDdQ5nyD5D3U0+xk/R6SzQqF0jko4FFGAWUrDhZBDp5O3/DamJTiSAaOpoz3n9w
LBBMsh4bC9Gb6GDcufFrjt5ptIGOGtqfP10+yDL3KrPi0Czr6u+zx6BLvItMyg/n
AI8vMIfjbgjzt91iYKLyXEcCCWV2a8WAzFc8iawLiCl6E/+F39aoQ2D3AMJ8ZXVA
DVEpD2lsPJjsyqJ9QsANsrOyvSA3RN+7vHIpKcAWFvVaNlE5gJ+dmblfTw5ONuni
oPLPeCBBVMTfrv7BLj8GbjxK60rGBDLo38ZOTnj+4jirf3YPA6g5fucpqQTGsQ3X
dsqKFOiB+OqAK5MHqpLZneGxTpL3yNlQM9Xg5JdJYS6NfnuVqyzWoH6ebs/bEuBh
G1d3+7gohgMeXRjIXyob9xTy//Fb6OPlUmUJIWi+0/T28p0GgKPw9RhR6NQLQmre
9YMkt6SEe5UVEueWNszvlQuyGDKxiCgw2Q4djb8C+Qp6YQMl0FryGEuhSlKypYns
tGyVwGYaoJSNWD2OcSKS/46QVs4ihrLtKsAHMVD2Zd3PXyWKceZEDiPGtPymI+By
jJGxgGCkmX70sOmcyIe4qUo2inf5qiXe/ghIgEm2boxTKrFf5R+kc4wD99y5ZHZh
C0UAiDmgXFg1vyaYWlwaDD6WZL+UegiIflRa2jx2aWVJ+zVjcLdm892v3xBK+yT3
BdhF3gjs9qOGBQOTTVyq/G6Qwn8uZv0ZUFIh7OG4eDHBqh1U0LZ4jrvvA3R3iDJM
2qnLPrHEeSrnoN2aF9OBksjZJbq+9oCPk8qBILkJ1esthhD6hMWhg7egbyts3M7N
W0T/Ads8U6z5TXPSF8XQctfGf5zLRW839ZY7K0cYZYdXNMMoRHdd2L5MNmuJlmVP
qn8OCVdVCJYYrOIgUVMGxqebYsvLgG3tZGvzE+RXqtWE3j+LkmMn46zH3qZM/P8G
5Ybwft0782DlqHvSEnCX8mP6Ymrwp6GmohIr85b6wgRo9kF8S1KDB1n3R54DfeZA
LsGQv3WxJvh8cJyzC/CigZw/CQJC/QsNhA2r3id4spnTH8YeJ2gQINaB03kVC76f
cYDjJADpISWyzT9b62jzro5KLEjXEQmCPna3TCAm8ZWtEB0ho221rORVgfyvoCDn
dLWif4w7+PpVgTWOC7yPahmIav9TBT9yTIonpnxURrKSe8YNEGRDhiao1FE6eJUC
ZqbIPFwA3N4UweDFQMtuo87sFIXFTQKZAlOUDwBB8c854udDevraj47rXrhZs7is
0euiwIRgLniMMXkvLzkcrO1ELBHxn68gztzKPV8bKpD30yGa9UdUg+lsQ4wklMuJ
yoDMGAwu7IZKBdOzAhdl9yEevYqcchXlPX4uxPQexsIsa6MECkOGxOdn06LboIbc
k55JLNh338Rzdpt/Zgw7lSSXL+dKImlw0l3NaClxv71i/Xz0qTfKVl1d+wNI4gYx
gjM3PjmfDFtj2vBZXFGoYxSr25an+30QTrhkX0eAP2sVbu4CbYYxL4ovpNnCEQMQ
DQzCc+AKXwUlQEyfGW35+ZpsSqlTBHcS7OcPCIi6/mUvLczOLZDtL+/v7k2gRz3z
5AItPVwZZVWwNeYFH061M5TYZk8Qq93TaS/nZNKm8RmcQFLSRc2U0PD008BkjPCv
9KYMYcGBQ8B+XFbtxHq/7FJcsxR3QDxH4KVCxEteOA4Dvqf8YSNeEGzh+IB72I3B
6JGKuIhW6AvmrPrIiZ9JQWYzncr7WQw6sEJfFMnv16qxowTKrAdOEcqHabe9dyoy
eAIZOw9bmAZjrVpRJQfTiPOkdM8cPOyF2/LqASKf6WzxulpqbXO+n8GH/+kDX1Iq
kSDvGzI+PavbsqlBV4Gi5RBF1YtUmtvCrGDzEgeTLQJBOl+gbJ66ta2oEV5HnCQH
Sa8V5tF4+izrpg8zi5U6sRVnq37p9d5SVQFBhDlCpZn3h26cqiyo9IrlKmkMdBkX
XmfChXg7v2XRIgMJKKlqmgMg8Gi9nFEH7o196SMxz4kykTTVNFOdtkaZhRkhiCwd
QohrPTzyw7GQj3O48C2K9wHZN4rSYaEikW+FS/96FhNtgy64Jf7mGiy0o4QGN20G
TbAAPRrImkVQmgVOxg081wkqV0OfKKkt5yO53gnC2OW8R2jiE3uaIWwao9deHnkc
4DgQkCfa7ALcpq76dVtwWOIPfHnH62JcgQ7a49xgffW7u+eyZV44L/oqBSuuniw/
hU6Wwxtft4lzMyvC2WItNXp/kX1riuf1c9CXSC70mOp/yBo09ZZkLy13mPAY/xvR
Wi+0amS30CNPdBXwP+Pfd+w1fNLyx1HyRhljsaT/sl5mp8z5oSuJ+pBVlySB9OGs
eKvKvTbjGNRPdoTpITTXi8voLe19De2J/nIdlirixmWwjy+t5F2IV8/NJlkRjplT
REBTFJG8TUjCF0bJhVAQ5TyR9KHsmOAQCtd2U/Acx5bpCtY/4ax4QSaNNRyyiKfU
Y3GqqMkLZb6NpGPRIQTniOvGZ+NIm2nDNbexvXHnj/G4zMFdyi8eJMChtBO/xSjw
lkhm+W5iq6u3Mym1Tt6jpOGOKzM87fQDEIsTc02AxbzJghvfD+FX0qn1SpMk07GQ
Lok6yQD3bTvjZuIoETIaaWII4ntdKRMtrsFBsnJtDrw8LTjzjT5zBfCZWs8rSVSu
C3sVXF/NrIdK1mo21VT9KP9N/kwLyoKCiHQzBXirV0Ny+Jh9xYCPXoYFAYCKGTgL
vizWOVDbf66nl8xbq3o4+vmZuUPtUQyE6c6qvExXQ6Oj55Mtv9IYqnWBSQcHKLtG
27O34jo8Mt4hoRc0+5fr+So2ylvqh76klF33R2hRlvnt3q4uKEFsuvwR+Sks6X2V
E4sd+pmB4Fzp4gtMlwzwBFMJb8C8DjDIdofgNVru7K2r/YFQy+VGGk2O3/2YfMJP
vh7umHOL+CiFcOLZjMy0ncgE1LqCX5oS+NRSE1Cnprzyc2ayzaef+sW7ft2d2nVW
3qg/KI2cHvjj8YZAOcUmPG22e3gbG/K9ovg7AnUR8lwT74hPcIK4y3XugGf9AH6q
tUJSgIItJtc4X2jL3diQXQrDE8qqnqwYZCJR1sWs4BqFyTUiN79gLaYNNyXqJjtb
zCdA3gqEDQyjW/NyAb0V8vvwrMDmUQVzFCCWK+Y7lDmpyXZTQ0+Srt6hMN0oD0u7
x6/nTVbhjvYJDkQRqjVwgPsnr3LG1Ry+mB5HRswMspYSjr5TmN54ckwBFbVdyByS
V0o72/WmQjd1ceOCcehgIqvzB7e/ZOx2O/s36Nz94HUEw2n9Tkvdn7LfdWVzLy/a
9MzLsOKfqX+r6vqcsLWpHWSiwM7HFzpvdo9yzqXeiVbdF9Ielylg909aS7OLHu8V
1iJr0sr/LZAHCnNsEwsa6Mb75+Dx6Zc5i+eNBRofjZFOFOHxNnEabcfqkzLeVXoJ
JUM28hLLCuXirSSQ2Owwo0nJEO41YZwGYCiTHNu2KwfTCklSX7DmmlcGG6IOJ5pW
PZHx6LPdUwRH9K0jHbZ0pmXKx3772ZgaVH2W6wkY8HZT9dJBjsyjIe4Ho4rWpIQa
EENu3dCDRbsllHj2IJJ39oDyNIZcuPGEKIe7GjjmDsDiG2sGp945K2yAMoLuy+fA
edtkay69bQjL/Q87zVA7mMmmAogB33KS8OvVQVgtXBswX1jWyI02dNlgy78e0UHV
S9WKdZ57pn1TbR7Iy024DJ6tkxy9m+e/KoBKHPueAIt8R8vRoaONC59hhnNLXWlx
WIQmkJLkWgg4K5iY3nGjpSDm+PPHXqrqOm0ndP3TwER+YWqcBWvK6cU+PraUOf9l
Tf0KnZ7FjFnHai2IXjk6aEGp7qiUzgHxJdloP0h+AeJjT9hSGyzzc2xnUE1NzHXs
i31DV5GHJ5BMGdZ88cvhAO5f5ddUHJgvYiJN+kLpQyWmF8Uk8XGTZbP0ALkxwxhd
4PM8ECIQlU5kBFfwjlp0qVU3CEPRhY1ZB32WlQF2VOZBGkRciqll16WYrwfg9HXp
+d7ODBWmlDNLEZIUjlxVqQ9Hd+OmRG3IDtsk7jfbkZNL/UnvibjiNZKmIkuvhbhZ
h5uoic/dzK7qx/yheiYaeM8uYsAtpiQFK3xMT01gwWTt5O6PKiAbBFAqBNmZ8DTA
mRm5Q43CdfZS/jaqNEvk1iw5rRe32I/ZAgc69q7UD35H9nB29E518QpHgpRMRKax
mqWDK8Lr3Cc7kjznY1bnUUOBX8dpFd0BVjZ+sEV0HF3h258rGeBcJCAZzgvrtEmK
sKW+UP57IoYI51LzUOqJNxNqgaNzZ+Kiig1YC16L3tfFYzESwNG7uFK87Vzkon5e
vfbTZx9gvSItEpzCSyJyH9c2tQcL807UQEmq7wjrhkEAhD/g7iBu4pS8P4sZNOvC
d29dxSKQKtaFJ4dLhoymps2D/hYSjCaRG4ufOIbPEQcOYe01thbDCH6JSlUTQ04i
8yHWtMqk7hNa+kgEIslfAVg97YpgtoYgzWR0rdEN5svIJlqlHjoCBj0zElEoFHzQ
DskNbOvadYTkLCdOKkmcxkGI2aiLSIPCOVZes5wFZRx0ssMS0Q9zH5TY+f6WUHTk
ku0cFn6yq310HoKEw2b+M5gcuIfb+nhK6o6/MlrHCuYU4Hqx/YAFMxcMZaGZZcXO
6koMt5g0EuhKcWLEIYPZxSHp7AxBgQ1tGHbNNZ3xgYK0Fn0vM/agMFvw3Hj7QoQ7
7CkenrCFi5x0uQ3+d1WZX1qihkgQuiufKTzLOGCAD74BAi/Cqxal9Op1EGSTnOef
nCdgQ67dQijMJOuRzomInSLtDxXKrp2Kor0YSLK/cIlNB2ueQ6fdDs38eM86/c6U
iwxcEUjFAaVLrCU2rk0qzGGHOzJOsXbJsw3ptXS65rrlpGAszB1b/SnfP933zuu+
sAtiY3Bde+zSZOUP4zHWWGlLXMbBuO6AGsIjcDYMb55xtyzKeeCnlvRe+ixv+Msy
/2oyYqZpzMLjbk8OY5aND5pbpbGc53V+WZP6JMS1GUE1xUbWnc3kiUHD7lf2z2Gk
Eh+HZuIn6OwEzknC0x0Jw3yhnusyq/uSrWp+GEDjEdWa7GvUH0JqXy9abGZ1fPtf
NCEnnbiBmtR23N4Y5gMdGdhi2gh9MnUG90HTx0JKmtqDlNooccXeEk1ZgUwOEs2Q
2/4gEm3/92BuNRYsoL4ABRVYi3OdTd/uk4IEKKTVFBWjh+T86IUCTCys1R4CRiw7
Vyy/RDXsj3YMmuDxcNcD8FgEAGpresboYqr0ekw+ta7LtbDfhBvF49JGwmiyN4C9
c1p4m8WKTpEPkzEjsuYETQL9RlUP0VqSkHrM5+D7YGh7pqVNCxo+Q5PraKdbgm2h
N9IvJugkiUYAJ3zhj7O6qQ6zFFrC2UnV4qh29xBQdGYi7cAKe5Mi9WluqwORnp6V
PpJ5Nr3PP/eihdAvktNxkgFKSsPwjpIO5usqxaM85xWKUh/IIB1L+Y1/7lBkeNu6
65FmC7e3AZHZdZVT/TGTIm2aXw99e5uH+QHPHgzGtWt/itMxAG+F0OvcpXTnlr4e
a3nroxtxBpvgnO19ClYdqqMiLpIEKrs/JLo12IZq0o1+sROLp5UDhYxxvcrAIRHo
giV3mLvIACvmcRlv7PTl9NlAZmLPhoNijdpDa54I08LUt+G9QGP5gcw4wzSyJaaA
fbUf/Nu1wMeYpDH9Oq6vKUFtnAIbY3w4zr90jSQWftViLAmTwfXuUqEh7WhccUJK
M6/T/z7ECe2hBroYOt3scQqSVhVOhLrK3V9MB02LJV7TWQv/QHlq66MQBjbB3JoE
GzKIu8Fuyuw1KD13S2jXdj5aUHZhNhCjCrO1lZjsM/NPx7ASD2Usas+O03CrADwr
C8q7S8MMRDEV3vt7OUAyPDkwouBkLAaOYZZYbJCRrYAEyCIdfw84nb4o8bikFS8J
IA0vzU5SEvbasK8P0cYBWGc8K9Ta0602/pWTH5/bdndP8unLwxkhEwqaHlDzoo/0
lI+nF2OPMJlKW/awvDkaSs/FYTmEwQ5HCjSYQPPVWKQHeTDz4Q+0dSe0kSvwzecN
e1Kz1eAIBSi+LLYZRtQEZYBOuG+an33eZsVeuY/D3P6FCG0CN8ZxJ3l2Gs/4BvKH
UYt/QPg2MsKGNGQqMstleA3GF02CFDV3XUgSoR7Zo/m8Iy3sUz0PNRUUx4drp9Pf
XM4yEb9zDWtIk00La5SVDvRaLhBPA3bFYF5ItAZ8RcRVJcZcbwecd0qHjxJ4UWz1
+ecHSf77K6KnSPfUMi+OIUHJuunl4lOeeMAteyDcIg1NHGJ4snaCPGc/JO2AF9IO
sUb7K4NACRCVnEpm5BNRku5x6G1WpXdCnPGxJZSu2uff/mjUVOa3aNgQ+fH64z/V
cAFex6EapOC9ihGiBdlSYM/vyknYnaWcxm9BvecfgtvRpZjjDq8dIRDYNRzmk6MZ
pLPcFPdnFj+ld7KaqkxtVu+R8R0ITX3Pfo9aUcZOxS93o94akPO74H5FIarIgMNV
UkQ3x56DKaHep+YEAnenS/TUvrHPWat7Y3cqeik/hbbSLbmsVy6II8xc7TYkdIq6
4Pgp7INmMsTH67zfDYKx2/deGK0XJWVsTPmY/DTwLxgFgksba0Ev5SAPZb6QhtyG
INsaJFBmXpI2uQczLUf5Ic/vnNN9S4DVP/177Xaf2/TjPdwMfLGJLTr6YlzGQR6z
x/1Q4X5ZcS5VxTVswLZoXCUAofT9UM+JY8UtEpvDbRx2ycm/W4R4k/5eYoHBgN29
La4mf5EzsJ+IBOxPu3VZ6BzcFi6j5F3IS7CnyrcRmMFQoPJizyYLbpbJEMto4o0+
RuBLDXwS1vlFvGdoRyi0VRPkB2z/KdGuuVe9gN/vtV0OeSRLJc+SXwezpUXYB1GN
aEF67Ml9C94dIyrY/JTWVMjIExUaHv4Bc9wBMWgqmAfFP7x3LZz7eUkEEsOjT6Rv
nE5wKzZ2ldHl/1Dmx1T7dpOVkh0lVfWILOmfBMqTi8XXeSptz9CUCnli1IOw01lB
qo5n30qM1U2tJEKEz9saKbsKb+t3XomT1syqOFmSAIrxpD0TQH7Bpk4RZ24jcStx
zG3cepUxDxKlV82ApMTb3B6Pg3Wy6nRxuQ3W0kG0LgaX2T2Et3bJaRBN6JukUbsM
IspcUMAxythOFZmgHoSdUtC1Y34BrYCzKBB9H/N2iNYMb69FUG3rwO0rRgaWUhDq
PsTQ/xwdPSUWVx1xFG8IQb3fEqmn934Y2Mp1bn+HTVK1+3sOwWJEH6/IE0WpTzr/
vU01wBjLPJuvIxKOM/fCjMeWnOor4mokhzMSJY7nWR9Z2w24HF/5WBHo+jpQMHEk
5RVW8cW76lCi4fdjFKkHd4cuLkPJMsqBcSJw5fx7ok/36B8I4Xp3Pjf10HDSevle
5QPWqBQCcIg4cBTt6fWn1/Yv+0U9uI/zQcNa0VIQskQL3v1UlaaWKKWu06iM3OvM
FgkESRaiZx2ovXuxSYvP1lR8I/omQm4bfjl/uI4nt4PuzqHuftEJCOe6WREPvozS
lmrdOrpgaeAVm7yFgbmGtZHcM91TcHLIxqw/Ge2FQsk7+Y1DesK39djmn50iwx3S
O/B6IlCgcEKmi8+ynfxZ9rc6xgCeRDGbzkbeE93+oyO0PzmQsQUg+UvkxmzIIOun
tVunwqLS+Sfd0kM2uLorQjJyi03pmjmhtLrxNE0Hn3WxJ2oX5kG4o3eQ+Ah1DGsO
yT5OxX9ht8LdBgVDrYg9aKq/WFmX5NEXM0YQQ9sXnGv4wms2RkYs5NgfxLzofXmp
Y3NR3IDwuSfUSlXsHqKCaKquHO1lYccm7xi9FS8lnSQ805HqBn0z2x90TgPwnm99
sbRJELfXe+lY0L62GfxZOj0vCfzTC7gNL2VTwSfceNvkf9xdS8j8e+Z7twcCVH5x
YSoduhsaE2vmymjHLp4KTOZPWL1R0i9FJF9X5zjojymUlCU5nCYDx7aVM+/KJL2D
w4oQmMUG3ueTbB+IvTRdET6aYdUFYPlroHhVro6yUTK1KfobzE27TQC1e2sPcHrh
oiLmRzZ2Ts9mav8qyiKmtjNua8hMpAkrMJ/XJvL6Y/lbzxZn3NgdyatZG4zQ6vPh
Vxj9Eznvy3CyaOi1pkwAQ9n2PncqppR4eNpn4VbXUMRTcw4QIyY78WBtJ2bL/OMe
MfTkJG143+Ik05K98DARalt5NtGxAG8zdsNsVoaC2qJ2T5QqJn5l0QEkGVmYp9s0
CNRfiWwyaaqPW/xtKfV1x0AxzyQ1MvbpWE9wvN6q3+lKJoYawM6xWXFfdpvMCFSe
8oMG8cmrTa4Ea8+EB4nmkIiV31beIvWmPhZf8fdOsAyTvvWMYBdJOvbdXz8j3Z+y
2BwB0I7KIsDPLo+T376nDP+eAYuBs7D6VP9JG50amKWtZiJKRQiZWhfagDWIDh+1
z+P02RN6FAI6jipnFjbCudsSTGHI7H4i6W+RdyZHRKGfgSaHL67pblejwmux9vge
196D93KZDsNvndmpF+0vTW9dDJrOF80KS5uO9Rsf5akoQiStPmSJSVYCwOt1X1mN
71LfslyNq+uuX/WwOVcJUmdk/r5DJ6TZA1mUxuGOv5Wx1CPfVgrTc8sZo5++qFhp
JIhd9Q1ytVSEOU2Rrl+GL0vbXkTAtFqnAfFRaT+oM080e9Xk3CGtiWfQ1M7Thpbu
1wIUTmpsefhvXB45e/leaG0gDOOdEEMiDw8m+XC/8Czh9NTdWuaWdtwCMhAs875I
eFp3Vh4ctl9pkAx6Ka4++wnjXjY0qZ6WwsiqYkPzB49FRcPF+q26Yq3CfLxcSzuH
e2g/TwqUS5SAk2zX7oFmkSfmu8pPWUNBCy4QrFWG40Lesp9aAj6WbQNBXppPWYWg
/Wb1EYoIdIFzf0HViRLlAnRdF/rUY5y4KxiwODVVD+5QtII0+RmsVF4vaEPcQlW3
yqixAaCLqlnKYHLA6GrARIKqwf0PkYZBqkkS6+jT3Vk1ChOHzWjG7uLxlCOzB4uC
4k6976JPx89XSwztVgglalBQWZuaExZrt5+QQR6Npw8L+7IXT0uqQ/9NKL3ufEzU
uxfNz96rUJRoJEYsoWTiNh85XAG0yTHH053W2cc+/EOOfdQm9juz2AQhadF/Expc
Og8x//Z5FGMy3FBOnaE9PaEKKKPehsKVoY8sevmn7RXzBsiGfJQ777XXic6mMCVX
4WnYnh0bMJiXZ8otYuC2p8ApcNV1OwO8YBlkaa5g//lOPEd6IaMZUEO5/DtCtUhF
bJURlEI2kI+4f7Fpb1P2JhwBrIUz/3Rr9BTjxvVUaHBwRb4g8vkl/RoOedWGd2Oo
AB2Mw2LiT3/6A9OVz4HicjwvxesXRyc2t7dAOtIAxw2W46BqU4q1J5BmLhjMH0ys
MxhVqsdAO5aV72gv3GPc+q1Pgsj+/e07WjhHuWBKDUrEQSKS3+ZyFUW381eSRIkl
evIcTsQ4Paq5+SCg+B3QpWX103G+KpLYSxOgz2rEeiavVpFMdCmmGObYVxclxFmf
Fj0JMFGN/wBqEB8WYCAg3WkDp3KpalYNbYB98fGbJWy10oqF5dkVNvZGqHf1oQmm
leIs/x2qPylxjwggAAOgDYm2E1ExtpeYm5VM01wiW7p2JKsqe4YBaFsRAVrY+SX5
IQjVlzI1pChyyOByn7gg1qo5HpbqjmT2oYMUq2Oh0jPAyPK5GZPIiTLA41JF5gsr
B7deW/AXrvSp+m2ucWgtRoOYYxNO+C38uxSIhLkJhazQekqeoXAXtlB36psKbFE/
A4DXJNp4YBEZnawoxiLB+sZ6bKphXyIl9i2tGqO+jdOa0AwDnVjxKHhUDyuAH3yR
+fS5xN4EFxu39sq/ag5PLjdfnsjV5jjnnefy8JlQi2GGb//Oq767/mi9sP+qTZpF
sOp31Ctens6zFluflDqR9O8+wp0pvwiehbQ4l36nkOLSr+XOFMH9f4C6v7e/ukgG
MSBCaPEw4jHLOF1DRp+j2lkBo5/ppHxmPb9oyKvp7uhMveZS1PKvLBfWV57kLK9u
USuFxlqfFnbVusDVkS6FoVWFpgnh4DOwNRXD8u+zAb0CuIGTjdG2wghhYAFB32bx
m/vmKnCNWynieXfg5oBEKMsgsIJrNGz7MMrKPR99dKUd+xP839bDO3QzRTz9DftY
kNHgLvCGa4/yFfTeZpoR8FjmVK0clyqaQgSrWAiYZij/TMTGREF17MdIgMUk6RM4
zeePzQ9PzngrcwT7DagDTFgeDOZmfT6kj2hFE1k5L+xiAP+nwJzyyfsgGzk3GHi8
dSwvlcLEx953MH+LqLQTzTay5yT5XvoVRl7gGbgjKxr0l7gvgVG4QfSWKnHGdccN
Ic0amPlrGGawFWx56qbRJ7apkMbOJ540hnzO4CfV0efDIuK1/RNE+emepOQjZ9mL
eWKWB1hNZ5iQSDeP6M0rvIREEJenhWBYg8kWGU05lH0y+aWaSlYngClFjEVuFP7b
DfWvnDRqv69dgmDQKZY5TQibWPhMseCradSvAYueEWgutFwOL5BvgxUZoFKJ2xd/
zGBlLZyd1XUZBm+zlAT6+L57mFCkk3YhkDfqI8QYmDgtLjQ6+qVIEfyowShoQ+Ei
DWNkue4Hib4/JdnV46vwO2ewJ4aMLlHnd7i6PzFroeWZr7IB+ySyC/AhhizwaxTf
azVzqpFkKG+csxlUiDkPRaW8s9Nl2zqxId30ZsdD90LgANPL46USHI6eZITW13dr
z7XjXFN55y3nRjO4JDXBmcqtnZfI9V6hJIE+TLqYjR6tfR08L2Rf3wDDYBdMQAJG
vmCZ3NEAmsIzfN34M8S5tbVDjX1A9hW1mtAHIfXPhlcCJclNita9dkvbcrU+B6IC
fwi1ApLIRtl8Bnlz4sCXT5ZXYLDCDnkUfArsP/g8mw/yaaWkq2P4pW2RTLt6Uxqa
XtOIMa/iUZfL1aGskFukDSRDSRgJVnx2g5+2h0AnHcsOCxvrWi42pk+u2TVpyGc6
lvSK2cgQEvSSeWdE1uw0opcNjjLhCr/+vLUZQIKxg4K6i8bRpd/noHpCs0tFsuRg
Ru8uOFORNqKNp+rauCfPu0FSoN696U5WCb1cMNG/N935bNGERlvceFCGIoJrqn7x
7nQTLtVtnYzdF/PDAF7RxLNyQpbUJ7ca0y6irGXrw92Wyen8FFsgUdnKBkSgwAZz
+aM+9I5wyZ590saQj0aA6uJG513g3jVMAffCsCjJ7SnXEdPUihX6QkHcecieCQLD
7/yDZRrs550xliWGQlzWnQ9/TNzkf+BTVp9ku5hjJptzn0Ck/thB5WH7DXOwt380
FmiwDUurgFMbzdeBRnppfcY/nJXBTKn3q1/2ymRrRlRSxBKapOKQVAtIKVcWLT4y
i7+4efmjvSvnLvaVeRZ8mOyj/LLpfw+Ey0TSjDeLAt2nP7P+qx4LJVWqHAYp6oPN
6rSgRfjc8w4Wd+KivYzkgtFJ1TJv2BGGBBOwOClN1WxBmj2b3sYbu75p13fnMVZD
0m+Z6W0p+iEGXsFpL7ENVkBRr3Fsjxky81vl2BeL5kA+5wiVzzJtOhLXBuTGxaxi
uCIct+62IKTaE7QBeLN9NnvGt6aIVZC8A93dv9D0Hby4Own7jM7dfQ84K67RnvMX
AIAktygXCVYDqWe/lt+y0ZSiYWVitDnSHEIK5Wyvd6oGTtUSQqORIOURD/m3Tlk+
VPKYZrnx340mIC8dHhe4F56y2FZVSZVz+xSyKK+svKqzYqIUiyT5wlh2C0VEUxtS
OiRU9ml3uwBS1x0lL2LCSyG//sHagFDQn8neTn3lEt1AQvcqeIXBY0i6ye14gFtZ
S1BwKtRiJw/OolzsUv2+mklyOiE2b9Bx2uahkt9qLQBtKV+Y4AlhIqb0xtUodvDC
ZKZiNlowvpmficoqeUJsElm0TIRNYw2PZYE1hlwyuKIlNK24q88pQ7D84vwNLeg0
XuNo+PVKEf7esIR/HVybDVpKAxXInAyfa1ou59ZX3e3wMl17qj48CP6qT5yjO5V1
O4XbJyp3J3RCTun/NzzOq34QjEuw1aZLOsFz/uoT8pbH3d9BBIDqPMZg15ZeVtFv
3CewueRCaCYrgi8xAnK5OwLvEF1W2R3ObTIxRAMtrL92DCDa/1+U2LPhphhPZKuB
ZVcu3cf1RWpW2TO8lbdBdkr67OAd5VB70DJ9Gh5Z61uO+WoqdLy0nrf7RENc7IEJ
Jt4LdZktXmSi7kjKI02OiP5DlnjwwwpmH9bj7aRVlTf0hO+jZk9ZqnHbtO0BOks6
bifMCUMN3tYNmtmomtJ7VqhEpJPYirDV89YTR1Mckv6tvCu49piZ1e2wFY7zVKmg
/Ln0L+agiUzzpSQbSOUfcQ7seyuJHoQXuzQIDai0IzAQY4RgzXBEmCmWykubOogH
erEgLEJ95lzU9ZcrCNlrFa+x2hklZCiZ827HUBMBSIy/k9++/EfK++7SPDnDhNFP
nIfQSUGE/gPnaIaigAufqkuWtG4yprn0NhvyL4Ok+aB1CLnCVFuHncZVCngxdse1
ZDY3KSONUMTTLApUYuI4TeamrLxDQcqtkDg+JH4QM1LQao59iA7ftWpXLkH/uNcJ
vuRqO1tyI2pgT9aCRrMlyz6yZoEPrgksUHkaOtAWR3vvvaVOTJ4t4AmCiDGYyYAn
9IUvca4GAtQoRnw4yYJfYGts7HPlP0DSG/0wqEnLIhKt9E6nQTabrczc31ylpKWK
EwvKk4DLwNs4ixTRfAz/983k+uqki/XnXevdKem//fCWhzVZQt+mLxPycsWdb8rX
ISj277zdX/vjFJTvH9F8hwiKvUERnkSUXR+3x/2uGu4jyo6kgG/ITOrN7o50S7jy
Rx839oSdkQmWOOrLURJX+ag3P8usZAPITJXLSUwlRRklkDuxsw5Skvf2VvUUbPdG
g0zs1TAFv6T+IDDG83QEl3QekByzexZA3GSXCfYrV1GMHXbUj+EYiL/tz5Fsv/B5
s1NiyOTWKRpGvIM5xHmrFpQQBIvGMIYgAoY1wFlA+ACmvZO3T378quPXamu+nKJX
fCXnyQzA3dUNcSRaJbs/w1RscJOx9j4znx+9OmL7vMtg4R6PrJP7HmBzi/IZbgpW
eHYuD09JSYif1aVB8iIJMu6zdLMjbXkYICMzRjm3vvPZ3N+UpeKoLbSMdx+UHlmf
jSGQWdeEW9ftpZUnlZadJB5rd6YjUlMwx2PDdFau136u/SHyVQVvfqaGmZ020KTM
RKspn/wTV+Da5+Gs3gcXHDvfrKjaXnVIS89j0fhYJ6VRuZtMQYIYgWsXbk+1Tnz2
LACakvL1qlCIYZ25MPPXUvt5cRo5wYIcM1MyFouqzCdcuFOgmAMXak+9glXT1/AA
s4nmQl/EHj5G2/keR924ngac6iAGzUC4vYs1SwFasCqo1D6GwuSyIa9woxq0bDFG
WkN0jwQsYTbjQMUYop3vBze5hdYtI3MlI4w6RWyE8bZSVZvTlQAYhWICm9Iic5gD
QRPDJvCsfHWPiVaLAq+7GH5A2RF6qN/sOGTCuGTtBhHDF1JH1PlikkQ9OXg9blya
IyjAfRApnMnAxxSSmq/eADIbvJvf01gs1NzrnGoegxXP8zxUlm+UGIGtkVsHM8Hu
lX5pPjGVCJGJCNk2UDYuqau4FDFOAULyGRAr82F18UpszgkK+Zg+J0sHy6m1EcW9
iOitY7XbZXOlAzRvgMUaq5n4SDwlkGEFwql7GrV3BYA/C9s3hr6JJs/OPhFlw7tQ
mM2PJXnmKa98v+ekmVq+puMQmDa8poU7MQHG/WbicqBSRm6ph13aYfkEQLUVBe2h
iTXRn/kg7UG9fGPBBQVo0CkWhxe5LduGcjg8xYU2aHgG6HVOM9sAu8JXRffX2j9k
ZiX132u0K9ajRQHcXA1aCF8bfQ2lH5yykxD8Gm/4lSWLqoMgzspQ2lNv4Xm8A5h6
q1WmGyfWNniZv4UefOB5i/LWiFNgeWRwEbreV1vNWwCUsQxUNmYepsPf3DLYqvd6
YWKWUdwOLmWxsdhbb6uhPdGGE2v0KgqPZ4WdDNNyJWW18HrqRrmL05mLh+pfO4V0
nC23vBHgW2A1CN7p3nFOIQx/UO+9Sxazo8XpTKKAnp8pvU3DnQKNmi9kFdmVl6iO
qTrhx1S/EcmXex++LIUZlI/sjkF99mjLe091sTsRM/xqaCrWgPfnFe2vGwHw6hyx
ZC30JkDrMSKQuWinxbbzFCZGcXHPaSsdblTY/Zu+IuSe1YZxRSu52+IWNm/1+W1X
zbKbTsG3VWAGZ5YJMIcbDH2iRlTsLXcy1vAFUcdRaz5wlBp1PV2pdCfYeQLWJutF
cw1LGolqx43PqInkDn1ij5ebWp1WLHFfK9lzIM3Nh8OW+uGpu+am14HX4BGyR9Kd
RrsUXLK05QSCfoEdCyNXnJTc/qYJoo0B9NAQ+aTNEze82CnihI4lBOsj7flM+Gs2
EwaGDEZc+dlWRxr1CFCC7umJxruWsJZN98EFbxM3i1MwWfgYhGyhCQ7T9vuoSWWR
Sde1zc45QwQgcP4CbooGmEsLulXP6XtHSDVNXAliToBRyqqvR+5xWzQltkxeswQF
xy7DV4RJQd/X7lU0gQQ6RdwLo89+eBjRi9bJorhfXWetnNUkf6i076jSSE1fQxLv
VsMMYqysYXXNOJLGil2Glt47eaPGlUUcKdWoPcq/aa9JNY1fEF7GdnkOdiogbUJ+
obWL34QreyERoavFiU7OyHAvy0NLYX00iEzcELrzz+R7ud2NMrEyfWMMyrDFgPVc
H+FKSQqkvIJRqR1ug2UbvikZo6aOJ7NtHl6bT01Ryf5nFcWTnxFe8q8GqepdkHRe
4WPfzatSTdXEd+sRSqdCh8BFN1vfrks3s1tPnwBMAi4IP5TvXhPayYk9bxGgH2hZ
8NWw1uLWOgKscGd9Ji05GQ/g2tejeTsSra8EgmGr0OfHiQ+ZwdGFMd2413RWTL0Q
Zj4Za2YnHBM5lHp91Ccbhki5XVLYSyFzo4sguswiLfRfFi54ZtP/PlP2aUlCnRY6
e0qmdv08raYOQlxru0fAaBXNMx1Y+R3yFZI0j3C611TCiOBelMqdeAOkyCQpETL+
yBVFt3JriiNSmzyJy22CSE16w+lJRQ9PzclEk+64kLjHCxtGZdOGmJbfnPPlsZuz
1cKSrLLIyzTbP4+P95Idr8WTqMSw5utiPU7BM6HKGq7EyLiVAoXaBaDjTNinUjYI
ivAVd0hi0ErN8e0R3ivIE6A8CM3Gk5Ej95B4f09z9k5tGQXDjOCO+4O5p2B0CzOK
0s7qgFqTMpxQ3oNjs1R7g5hRSoKT4YIYPqDpyHeBMBHSIBcNmVLF0JTs1tohud5r
rGWeMBWZr/3HaIakJXgqWqFRBtVXxob6wKVKKypvW0p3wIcivTE9RE4iQdIYhjbB
9JGpQwvBSWX8N0VSt/rNkGgR0ZCN/vuHeELOwCNYmsPzH9Tx99CuY8SU5hWZZM9f
OZPKyiHXq3hATzia7jO74fMkk/79qPPOB7Pc/QS08kVD4hc5r56g1rmXH3qtAWH3
1ScXzQM4KDtNWr3mPM0hXOPpBI2+/d6Qk1Pd0EHEjE9OP6scX+ur4V9RNYy+cOnx
jS758QwzRMuPQxn0Ly6Sh7BGT+2s1/F+H/wJVmbOlNRN5oXR8hv8j8x2qAnsIZwY
b6P9A1rZEzwrqxjJP1UGqj9JbwsvnpBVQv8qhkW4tBzYrQGRnYtu1mSFRSlsxnzU
k+mFZwk195VhDru+FUWmeUreXXLEXdFlN18iwy7DQhbWk0KvFidty0elJLIk2yLT
zwZTgFxr3dsoEbuh8LcnVFuCLfq+Knz/MMD7YoPEVYWH9qKALgf/TPGEMqPS5f7Z
XLedDyEpuGhVRYM/d9SsYcSRRDH53R1noc5J03vgzoVp1xeo0pRI+ExneEnJjraj
cLSaDyLvrJO9eFnzl8YBVy0nrDIxScKp7dd2uTgUaQXVIDlDtVqZhHMhZ5bQmlSN
m3KxD3u2EPI2IWW2YQTlyNoq/jYt6D5FhZAFG0KSMqwY/OBmdqMtrWn8DfQcD7yZ
kmHzWBZeMqQK02cnBtUxLik3Cn3DShw5ONHGwu9azb7cihcVK1jhT5SkuNH6hL1g
UUaw5U7nXE2NL3WvN2D3/lI3IKHu1qdUWrXPs/kXvfZ5hHhlKPZAp0AnKPbfwHQy
UfJQTrbcTm6BGLlaoPbp6uDzHMT4ogOI69R8G5eVMhObXEkw985m0MZIlxm7eL9d
BMUssw4hAgYAUW7kXcgRuHqfRgrOTO4SxL+632IdfS191rF38VotC2yXm6rT9E1d
9UY2SYEQ5x4UASoono/3ovnsda3KijFT6+d8ZFSaHSnSn5pM53fnG+4xhaE460w4
CSzBi3QXyZGts4pd2mWFqI64G5zwIwcK4BGDdg1E4YGky9jDGgR95nTd/lEik4p5
fToGC38EtfNDL/DprtItoL4GTAGKceLMYOH59zD1poooOwh9wZdHhbs5c/aAznqE
NCcjhcaTNZDMlkal8PwfmwrNRClwIzJzxCMId1MzSgOp7+G3ZSJESRVeFJcA4lHG
cqs65ykXCrWrpfLEoRSR0FAj2ArAUcJhOIH9oLPYswe9BzCkh+cHuFK3/0MMZWou
hYyI3jcHmFR7ipBhU2NsUteQivOSVCMsBalT5xzG9jGnHZxdioBRE3ERRradvu7V
W2fmhTyhSEeb7RYBotQrWGxqjBU3SHdWfuWNJrn9kzArNevwkwgQr+Q4JezvswwP
yNOUOG7gdlck0jmE0qNmNiRgaTXF721SBAISDU7mlMqIt9sSGuvmZExUI2uNIxAH
5gmXp93eZ3fKksQKBa4GnHP/0DTTwfP5I/L895lXA7se+WaYAQsTE7067gbqsuvV
OIdkf+0MudEGzAaiJ9eirdm/N9ZvBYy8AUnXiSYZAOLoLDtD3BprcZl6Z54EPZfT
xnhVNO46I0g7XVGuHaAa+E7l3yTxZkUSrBViHxwFvMncoozohnoLZfVIGD9rmPZT
gPuAzLHuB8dgt3XBXAh0qHyavBxqagZFXl1Pnrnrxjf0Of8B5nN8W8lX9DjHeZ/V
SG4eLybhXByFpf6GIiyMrcv+WyZjCKaYzygAI9LP10uxVD5wzVz/PrQN/jogFS7N
hPDwb6JW4qAJwzQsWZFKSR8QYKoI3PkFO7qccx3GhPYXDOMEZNRE9xzeF3g8FGQS
GbsR/kDk26/B2YLh/UJy9ufD2G1is/TlZRISW8oFY83gdP+mkvPgii1K/yJ/Al6J
8/EvMR/FEL3wTeMxdOYzK+cBn8O7ZLKS0c2wOkEPlVJl/dy3oy+tuuIm1T4sZfJc
`protect END_PROTECTED
