`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpxk7tyhcSvA7nJNCBEZkOyjNYJyX2gLxr9dNe1tbbB9CrLn8EOFeZfeJtTTQLeS
7k6teZJvTVXkZeRqg6wy/54tGR8ZojvMG5TiUUSPXNXfL9SgLgJpoosFQPYAOxEL
nVuEEvNPSQ5zoyR0xcQucwIPhHxLIZb8GrI0ukSRWCMIEoZahwtUggbvm0QdqpJs
yDeMMh07WQv3zy557BBkeYmQfdEHJ6yA5hsUy28dikyx0R2DJweL+sjgVqrRYpt8
GqNsYRtE7HJPIT0n8zqcq2jOGOOAWuwa8DpJUAqC2zeQbxD/gvGVzRT1a6k9TkcJ
nYhqUJGiXqMO3Ee9RVMYw65SQv/2R7r6Eh1vQOUQccDsqcqhaahHGtzlTA6sXKhV
53gYzQhl5DiJ8dU3Q/fIW6NI8ykQ98LPB7596cQJwYVVM8etW1qViPSssSHRiSyx
rY19ji4qDLB2QqQHD9qzG/d4CegvmcqEOcqhJDOpV9YBz/+11xt1kNwPG1SruWfE
3qg08hyieEf5s8zmoWTc34Lh4H72OGruoJjuM+1NXtSOT2rhiaA0naXjat56EAQ2
kwpPlVF2wyX8c/zIVd2v5qkoM6vy3DUAseCfHAHSWf2iSRW9P72p9VGx46ccuJFl
bK/Y6wGzgAmhkfh3mOcJ7PFW5FnX0O5Feq5w9E+jsHd8wGTvHEwIHPNJ0nPlfznb
Oc5jl8JEmSg0ZOOfhUtP7UIq8pKWOrLJ+kIM8m8MFwulO0YGvOd73CB2BgdrDVFN
5Ap9ZSTSgP63pVpvreNvzo7F7h/8rYdTSTtmfjL61cHAdV89UFFRereby2ylHC8O
3GNNnLXzSOoFZyIdhJaT8XM7IFisQh8G6H+OgcoHqEt3oj9xypLdMQ3g4LkNANyd
o2vSLOaUbtlxyBFK9Vp2EuCfd7U57fjRlKoVd+B5Z5EF7kTHz50OM+foJrxEH3Tq
58rf83Mdi8S0SIA2EmKGXjozWw1OmlClgVIQWDxnqOCnvm3dHCiFLk6M4Y/YqtBo
7/F9eX8U9b0Y4EglzjaA88p49qOKAdwwdPV9suuU1DkPRHauWU45LIQzKhIBSWZR
wVBJmPbNTwssZvZ/kaR2XmXoHJkSUSzcS+D1SdcprMyIqoBbpS8OdmYaAQKRL9sD
53ZpaQEWy3phG2SLDfgEDvpJ2BK2CpzWxjnTF11wKe4DnWDMaWksKt4y5AV1Ad00
ygsM7J2PaMnVogmqCvlXxJTPQL2zoD0jy0SrMZ/VqSI0lJMUJhA+EnQTQUa4j0gm
xQ5rtgXixq18UVpHTtpnjqh1LJDDpFzJwweSYZP5VU4el2P0EzUFmu+Yln6xEmS7
GE1g7abf2hYe93/S3y/R8d1ys0AcM9YLQ3+5F4OWSrz0V8YGcGbHULVMGkecdToE
Qw1nGolJJt1QXMZ1CjfRg/fiYS5FxQjVB6mACUjAGel93HafRu4cYomq8xtkkB+X
FINMatmxmeAVyYFZ51K0CV3We0Q/YbZrJEb8nNCQRL/u0DuyEx/diDQnAUE2YmJE
i0RS6FeOaTvV91t2IvblTzh55DnS5Tei8411hRIHdjAzsZzJZJRiHjavHM4RxDpU
6YaZo2WEv2WBtM7dRfpdQzItrckOl0PR3es/D6idIDSzXg4LALvFQ0uWiVdxdAwV
kzdYNvjrj65XTH//ZzVe4p6kktOzk3fcuDt6E8FsFUMDL3t+YnG9fSeyskMN5iBf
W+Y8JGqPtrzoO16GOyt/V5t3wjw5ZRNcY4Z9EXJwQMPxD1UvkYk5MyKBKRqv00xd
fmoiai1XkGzu8LXJkkG3n5OWFtyNiQXZOXRDY2LzWQchIuJj6Qnd7Ft2Jj96cwTf
smkQxJ1YSYilX5q+NCVJ1xiqsW9uqBuE9y7E/muj+0df6lGFv0mJsnIz+6TwGFjX
kPV5dEcLNOkYvw1/Y/wFUkRaXBsPeX7clW6tPNZij/7HuB3RCEIDOCK9d2lKa442
VxuXHsT/ILv6aJgpL1iHZvSOHKZNo/VKBpvcsSpD8xkcz2dXm94aV//s9Zz03CSE
5YXXNbttqnb2R4YGDDq0n5SGUwwZorYhWr99rmZqL+BCNpWp6bo3rl47zRuHpRKV
YaBHiGnTIplioKQbUbpqwbCFxEBHFXK4fRvIlwWRf/5ViRQTqpldJHiS82rAYLOn
NFRDhcuzz/ukk7T2pUeH7vkjUyTS8BqZ6qKobrX19lvkx2k+K6dgOgWNOsj/ceIK
4AZs1Cs5EPQdmZwLoQbh+aGqeGACAUuMM9xTizz5CjbcvRy+gkYfDAiuUoIPRvrh
mThwrWxgRG4zw1z5z6wgm6D80+XjIn6QZW303AMul1pf6e2ekYk1dVhSVzf3f66b
OYGZX69ws4InC0gLOucsWkhLi93InrY2Fl0quZfvXFSiSh25hfbOO4DY4gPFhSSu
PsMyPqFxK+NlKYE2yURINp8GnUfNiIXzcE3RPX/2YMEdzh5X6YmcyHsBIika535m
N2T6XuZrAQzPd96SHY7rYn227VwTbpW+RBqIA6Tkv6eIyq4FBV4FXUq11LBy1u4e
Sog64VJE3E1SGpzbQB9svC+QqxQk2siPEuBegFPFblI0kK4X4ntEz4gpdMPP+DQX
alW8TtS6zElm3ireNRK2u8vUTUhSNJ42K9g2LrfWxRqpRBRalN1KXsB4RXoN/QLJ
CEztAFklHQA8O2E8T5nxMOzYODPZerWaeHHerT+7HIVXx6F5Y85t68dEwXDyeQAu
YmiF9W9LkKC7z3by29Yutf7iMLVexJSBNJx1J84FyNlBQ39khSbrxM9Kua+hqrJb
Kwx6HZiW4I++6cn51fBozkuEmh0W6p+q/SSh12HNv43ruj91xyrjN7cbuq6A1HXf
dOLww+hJLZLTyAdtmZ8J/GN1BZFDIvlPyXHTzUaBRqqkJ3oGo04LanjIO5Ou+PgZ
6dkmt5v1ztdFqEh0Ed+hXjaO4SHO8eBLfJn8LednwoaXoLeMO3hdeOu2vnAUdI50
pM2LqdVUHV/9yHexHVuDSCosdbiIkBH5N53mKvZ5oebd/p5n7yyZm+z41rAesINZ
QgqaSYsg/nRpkhjoriKEh4XpLClNFw8/5YM09R5uImI/zJGbSYjw6uiCWj4QQjFr
KlPB+6AkXDfgVQ/vpVFeA5yeF6GHiYjcd4M+MdqscMlZojkw6rFhivGaQvJRuK5o
eanYNQ4a0y0YOFIota64hAYCngil/nCwjOnJ3O5/1Vs6CYy9kTz6wnHgCgcVn7wh
hGt5B3nfgwtjPBc7i+t1HBQMezsNA1c4m1InuLLfk69on1W4ccfbScJTUW6gqBYO
EcDuR0z6X/0fP672sGWCLEl6Jv44VqvDMsNrufuah0u0lq1z07zbXNzPpPPxIzFE
GMLOKTFPxpPGzE5+LGFblEYNIMqaX4WofCtEcvjoQhwdBaOacP3GzUGQCp/S3ZBW
KCgtbZW5LU+RLXr8zqnprfyhHtcgKIOXqdZLTGonIe+ZFNI6s27QwcpR5q8Z3sYO
+772rz3SCHqFlLyrTkDqnMYvxMYyWmpWT8KjjIyWqF7xwrfGa7PTGX797QCMR6yD
+eWUfue+TtCs/tb40h+LHSZeP/yX2V/no1UWe39H7y8eWmaLXUzQvroZ+ruOxqNv
RBv3iAwhMSIuJ3Jif6W5Y982166irQR+Q+TXF4USBdE/Yr3JIpPJTRR6d/yQAoTO
Cmh20TIU90h+6W2CyrXiBBezxrOuDBBkndy2wJnkD0j7JgWaLPAOKkTw1S/I6vnI
+9i8vqMtubaNz4AOX8nU/ul0uL/3hMrcda75RjCBklfCUK4+BL+nVL1OF2mUv+Kj
Xr3/b4aMnoPRHeyapdz2C5NlpgGu0PGzdy5qgoaHBnsaEQEHjSryXuu2x7PzZHOX
itnV8H54SNhDMrYihbiDWrJ//rNS/QanFWTzvVBKKBmklkd1ZaDqumI+7H7p6Uj7
40nMN0RVyCNwh4HjyIFONLeN4QmMZBxBlg1BuBRXf0f+t813s+uK63B0kwOWjpCL
8c9tgLRa5wdhZ9DJRf7Gc0zV2dMbEo5z4lH3TzK0YJX/ND5tDH6kSe5T3ExsPl3U
yJeYr108PQTIw5025J1vQ1hedSJ79BFG60x2TOX52J8V8QPprFEIx00oH8wgnxBA
eqeFALEAf6NHC+sCUjvOiPCnLOSXQPnhByldJl+ZgLXTJK9fVR5xQEpWb1PoslEV
ZNIkakLZIyiYRh1FfkzVtin0s4k1qODEUARHB4XnzuB6t0MPzRyQ3KnX8KpFWhfF
9a05+ZaxixUKvn0fw3/goUcbqhBmMevqL2MWzPShexx6wlcdYtLKUyperEs5HV84
poRcyy9GrL9mK7ng/Qfba6Jr5iDNMeMLiIBNsGsn585naiCO4r2TBngBGQ1fQWsB
DVzD1jRy2TpbM/OwUofFZGf4jNBB0NhXl1l+hido3hl+aXo0+XURu9wMvcgxwVnV
8xc/99Ij8Z1mmCPiCmFhVJyfo+hz5p3kb4qN5toUk7zhdvlmweTTFuMNj1YtOf4+
YQUDw3OFYAeJevzudJOjamGFDqJh4D81L0qdURKxKAKhtsoN56w5aR2OjZQZhRNr
99yFGeIAc14W+SFy+u2DOPr6PcIzfYB9zRbrmxOYwVBVSryHjTH835rNB1qr4HqV
jxyNfLS/DFWOO67/3PpSG87Ph6EdPgQxYh+TOn5vIpJpi6CPMem1CiZTobE8kTR8
nmyB9oR5STgQKJIeSEByGGtoU15e1TQryLVLYn46vPTrl0ri+OHlWs2JIpo2pc9U
uE/dKVDt05U8VniOk8PChbkfChJSKn2ypnDxXDeBepcXS0OJVGU9iHI9TjvGQxWx
61OM/eW49va5VcChwsEJ/y0MXmSKISNbKBTBFx3yFsulesHW3/diLQd6YFc3uNJH
UfCHCuM+TNQhEEsDdC1uoYJm5PIChod9YeyevsMkaYgxoYLcoyQI0XNXpnBTg5JM
Fj0/oUPNPsnP6oqMPmrF5NHevwT4jc4rYlJdVJn0mz8ZAQhJf/aYkWvNqURL5I2A
PScCjcUsNWLf3Ue4m4Xr+7Nlvn81BxcHTcvQ4G9MCfCzGduqsimB9QnsdbHBrY89
AamMGZ558x1F4rl+UkAx/Oij+BtIV9oGc0AgoHFNFGzjccUlVreAR9Q5Eicz3iFX
J7KHRKsRiB2URhAC3XAFQo5s5yyOsygVj4eFezUZZB9zySKLmbgOZVK0i262fyWH
m76Jhg59QyUYKb6o4teJFnasl6sJjPcer7RokyxVZA05poXHrWPRAynOYmmX0emY
8a9nGa+06YCia0CSo/R1bS9SUrJOyUXafEBJvJXjDOYyw20P3/m8502XvbjCn4Ft
J+Ud5l6Zitl9RIV6VqGDhITsKMkY1dRgxGqAa6RK6roPtJskwE923XHkiA8OuWwR
SV+PliR5yHI2u9ICQyDCXNIrK74NiXnLlrAAhS1K1z2ktFFvD0Qz3KlDmPjl48I0
Yx7sfTMFT9uPK4hBQRPbNrZ2wlJOeVGgPnt2FMCzllgIGD3ulPWw9rfEuU95D8bY
fB29X5b7PrrKAZphEJ3ZyCMfMnx4uqzDZ0Zuxd2tr3Y791uuXI8FAPQSM0SqXl1Q
ictbhYt3eaXFsiPNvcSy87ZgqV64tSe/KsZQSxv3D8nPOfZ6GnGvArTfjXhqa7tq
Eq5tdy1VQj3r5z5Fz7c2BSrgWPDb2YH0Bp3JXI6vsCq+eQkQbmrmeAloDvl64aq9
RKUqb1pic5YZghDcQyoby8NI3wMxryde9OrL8a70v0pDGLCHVC1vver5yUMrOfEp
jBGguvMr5mhssJ3Z8jH8pn4pXrKq1tY3FGGNUFJihYisAhW4/iH+5nTGoFEFycWE
9Gfnda2vFQoUOqCB7vxTujQutlONKmU6eptSdwppjKEP4zwp+WUQstP1f448M2r2
edYJMkEVQzhHFem18Am5afoyma9l3j5mS5Kbj9KD3TX4w/suTiBqbkXeuwdyNABd
KXNq0l25bYfGo+1rOeEnb/awZPZoJJR5pp0XOvQPsC1FGF+AHH8gP8CRcShUV4lb
I+SjMzsX6WA5mUtjuI5K61P5SBsUwvcreZdvHp0KyS7zc0A3gx/oqqBvsKS0BxYo
KgIOi/64rUOa/lwGAP2EHhlazdmfcLdT0wx9nb3UmicbMAii8+/vJrM7e128GSV2
TM19aavOO88O17lWCfDefqpH+WQ+5HDHEbI8XL2uV7Txrtyxc8qsMWYLQ7yxUQiw
LO6Yzqcl20z7evRkVFJzOvN4tlG82Hdu3XYPL1SAjQTR3UMprFX/SCWyAQyc/czw
lg/kxq1Bdpqxbx5RF5+NMJo8bShyQ1cTiXpraDi7d6dZTO4guZPC7rNXkUzAU+gm
YWSG2KdFqrRmRFSqW2ZPkIwypH7lM2sKlimy/stMU4k5h2PvRBhgpXUhhnuYjqIy
EfBLZRIHb55DvwhatXq/5UjISTgawEK/p8AOyOZdTnGTOsEFYJw9LG1/QfDwAFND
gUtIQM5fT5m8rLDzvr2+gam8QncmwvvMAL8krgtu6X8JJNcea+qA1ap5kP7csRSv
VY58Z2DlmRRFHUD3dj8LCWK1nQFCWG/HEkF6iRzVni4LSNGje6lwow4LheCZ/h+g
Pb46eZ3DAn5fsYk3NFPKhAcotL7LMvhx+znpPTSbtZ4+j6bsP3me4DsYL6Sv7e+h
seBpRvdHoQSYhljpYJ6gTYJ9TYYWA24fiPHONP2CoW03QJJq9rO9IAmi7SbsgXOe
8Rotp2S7t14t3E6WkVxmxdpL/lQ3a+60ATLuKLwkSWU+O1tVHStaP4qmRqZ5cT2d
3IhDsDKNmkhCofFTDuuodfSMTqEmZQvnhxzT3WtAB6YWEc7+XAUC1X9KglCs4h0X
gndw//fJPc64s2pKG+AzHDH67xqPkYlEvUM7S7bHgEffi3NiWoMY+H/MUbnJfzO7
K9MJCd5rr02YdBtYtv/UdFPp6Y8k24eFHrBKwI/wGHnX+wSFpk0+SiPOd5yrYo/U
y59twYOlygNu+C/UioyhzSqIBX12PkZCzk8tRDbL3Ra5tX7yyKj7xeP8BP3cdQiF
W6TM08omlp5whHAGXUl05dO0PNOqJ66/geiM1Q9Nb6tdnUI34Zje2eoEs8ZResM1
jkgSr5+MUChY+rkocxnME/Few4tfiZ988zWLErRxb1vdBG9uH1I/C4PRX77EFKvj
1jJz0Y4aFY2zbnxpj59TU0e06q/zKklbaQ/6MMm/jQhJwWGbl2T1dqZc8U/zY3LK
hz4G8MZJJFZclZR1mCzpmdy45RvCyYkB19PME50EGLw4MIU7y5xD4Amq0W5OhI1E
luuUu+gJUZiH7WDTkxNiWRaE9EP6b+O9IYkZ+prUQZFZhdGyLroQYeFJ6fOv44ar
IqkNmYBRrrHPAdNynX9J4vi7wZoSVTl2BNUH+tQhbpilgodH44yM9pxBXH3k9yvM
a0/n84SgLG+R9oreWtiAnHcqHemmNSFO++W3ZmUmJIEnxqDhf5IEkeHRKyPAQb1A
CaZlZ6YAIo8GSPJJ9v5FrHvOmIIx51A+4MwAi9xaQYhd26pxAXyaVNY34AQjN+Oy
BGhdFaDw782VZ5ssL7Fi9i8xHRBa2DEM9kt/TPBo6Gsk2dfYNiiKOOiUVusw4+Ra
YvjPMncpQkj4KmGkB4+Yv6Jd9j5+RI+3GIZFG8ORQCtZVw4Gu+H/GgxsKnxAlubA
P8hFRcfL1FWh7TFYUi+cY4e7o5ZNXfP59Q69l6/UFyMwXTaObHt54GG9K+e1So1U
B0IsU6fhGfLmQi1FsoKRmaBHHCjWa/shpbqS5sU03cQlSjer/9RpYbX28bth3Ukh
QqZ/URGIiUjVQ6lDOIcJrzkxCjH8P1fp76xTf5L9DP0PKSowuJTE6SO5xU/qt4uH
Xx6vLTPd+YrO8FfBHPq8gG2gZEkh8HOF+RPO5kI1x65cB5Peg+AXCrSx9LZWJgxG
6epJzPsMg+j9c+qNjnJIfRy+Ij3GeHsTO9iZxdTKWbkD1K2gE4LGAJGB0nOoRJEA
HieuzuTbNugl24WWhjot/fulA3QebVPINEclESputxwdHEO3gqukWMY/McUW37HU
9s4x36ju0xWNtXmYxfEC5kFc9bbzFKI6tcGZ5pZA5RGjUxjOvFryzxtSFUCfnX6f
Sf5s32joNsrVfcbYZEDTQAKNA5WucYq9CXXabYKX0Rq9htwyl0kSFKSsgp0uh9jy
OuRsq8i4zlCDg30o4EVWzjosYICJTyRDVEN1woXFotTvsfqAcLTqLdF3pi097P6s
F8CKJglnntqdUrqRWXEIO2Dbh1Gi0PCF9eVz4I5ukK7WXRyAlKTi0RHEPRmjQ0zL
Z4eurTQHDhkg/dGrRKSnEQYSY0pRHlKmMwfzyufmkMktcDdrEbUNZHZAcsfMuZa8
hmIQu5brwlFBkj2UT3aPelK4W+enANfRVn1rcCEzT9ZNUjGjfLYlyQ1njoSI4gxe
69uKYsjOpenGgu44ukwC8gSZRJHm2deQFZ/HVqAD4o26wyeWF3nQAnBLtHu/Flyn
LCv4KKM+R9hHW4A3lIQHOlf4tzlM5YYeUiTuDdc8JfGHrJ+JuHq86S86CGZCJyem
aVKuWzhMiLDhdcp39TIJVqNd3TyJhyAgiWcLezG4JljwcNubvbqu9BaxaBP1KnI6
MDtMLrI8NuS9/llRB1/Eaq1jI4hJ+PW1wC4qfSsMmv3VRfJcySnekK5lqY+/Zsh1
hmvJhhHGuGu8ar697nbPQETm10Vtbp6HcKCY888FgDaxLqSACew/uYne82yTVYhi
owj1B7lxRWIw3D/BawfDwIsRVa0ABsEpwu1O04VeHPa2M4jSqC84r7+ue8kJR0XP
it6gzxSzyJxPYSI4nXFaZsRlB1QWvE75AEUGvquKJqnkbMsVzYKkhyLBoNWWNnrE
fczz6XtYmjOU7ZQQZPBgb3cx8Q70ipK8ssFY+pCv+vugJWSo1FCB1NuXYujKTf92
NxyIBkgwMVXXPytkaou7xzw0rvmbfa0OM5WczllgVdx1bozTu917ySZ06ythF8QB
5h3AAWyZk3duxUGxiUPMP9PdGEUlCFHcqXer+FyUPvcExtiUwtChlOk4M5nticwW
Mfdp+RNN9JofXvVlqEtj+LWGtNlvWYydCMrXhADjPg1Apb3Op3k7XqesESanaFR5
oB2HCy8yozIfXSp7VvMEWGOkgchH5+QSxmUidIjV0anab0C0qjz04JmCaPsG/5Sq
FcGH6UcdAVawJcT+GtLolkKbRi3TAVfSNRRCVBMr+YaAb+LL77KMb6aYVkzgUII2
Axk89anmx08dzBPLmGLftqq20pqDkws4IYJzESiAiGGCf0qQfIImhtgB84aOmfox
koJi6ScGfvCWqJCc3oxr31fTob+kff815S01w0QpskWMh72zNShTTgARRxp2VGMA
RKdJ4TzzZHF+y+0rlyoktCYGzCsasPwB3tK5mwjtCpCMq9umSUM3Rs+AbnTuG7E1
cvD2ZZ4ctgocTNp1HJqiRWcvw/+m0Y/gFmGZQTBbRK8FueNhnZSP5VNWvuBlvKrg
NXujJx/6dGNrJnYvRyWiyFyRthXLVhm22881FYml6r0Tf68KgF+NE/uRmkwyhnHs
mN7+YJ8lsf+JI71bry+ZNFYy56CXE76/y03aVKieECsu3wjVOkKKLVutwf8YXnAp
pftwVIeKVSbGlkUGyvqQ9E+qJZCPijcKl7W0DfroMY3LBXUENSabRsGTBo99s07j
3IRf01QPnXTb+PdP8dxn+dwL+x7ycIityx6pWaahuyItEH721o+T6NtlP/RERtuZ
SfALV2hqqqDdBo4TeSKkgZ47rmGIwoD+MfFdDuzDckIlGIzN3iWwXvi+R4ZIGwzq
pXjkIo18QM7TB6SMkkRI283670W1rSvrd/Fu9o+Pwiwd0yZqJrcp8XpnQ2tDfAbZ
Ho5Q8cd6ZfKh/AYoYWiRzhBsVCDO+O7gO7rOkypZkGUHZGFuWj4VLmiiudRkdRW3
WrsaG7EYkEuby3hYbqaRP7toeyNO0qu7xVX+8FSOXoR4FpwFJDC02TeK8KHr6sy3
lEZL3SV3BpvqxC8kmNOj2lhHOdSKWckqM29DfxUt1kzCamg8yqHVrRiYGE7EJPmF
YdlcEOciNs8739HKDU5b54lJM+aUQMlDet+KJ8pTkxIXYdOb76QbL3z4bt1m+lHN
y4pFU//qc1lFuJKVo6Hvs6SdYR0BiytQPoBjtBxlCZydKCvZCZ6pixY6Vr3chajn
DpLO0Wf0te6/pEw06oS7Xc9I/fT1lca/q+lyavowI9XOUFtwS8yCKlglcY7LSH8z
FG3tGMpcNDmtNnFnDia0myshhBlAsudznmdlILX3FtfjfZRwpc2VH2BlIF77Pfy8
FuanEbdzNkLN4ij76UhdMdWxzEnpCYDeFYZxhUAGDDQllYGtgQq5seA/CvLdaP4D
o5tfuEi0jtngMg9tz8/eC5+WNWEBOXZMLKXp87DKOh/GoL9Sh08cvYSS5rc+xP1j
nRWOl5K2WCkw7f9qWBWGTVnhllhmZEXq6m/EgC7Z1PexOG0cMEKdd7KOK04uCOJo
K/VeHGcjv7vhZMVUZn6rMcfdAokdi3jx+0tlPwSx6dRcQqjtBrYnnaduZJsvMHOa
xg9vcsL1nXgc7hPi2jBkeQvHT186ILeda6J34OUkRNiCAPS12eZClgKUFAfDJ4qI
td46dufWl34yJ7ddsEBqSMl5t618YvITnnKLPX8uotGgFSrArd4JX3j+RsoLssty
S0HBtWcTK7JBAXXHFA9zGWY42DPHReha7CQOtGFAD4nritJiLt4pf2nHTFWiq4Xb
uH9BLhqm9PFR5CoDc2bT5R7PlMTWZ9M9sd/AAGVb5GW5AE3PBNslDSUu3sgYQAnt
ETGZdVOfcTaVqRzhYHMD2DA5pH1L3Q9Eg2Anhf5wIMA/tIEgoTiSPULo/ZictA17
Ct+iuEpwD9WjZiBACLnhASL4qlzvscZgHs3W2vLbfRnWzx5yy3U2NrALJrC9YV6n
FLaVXClTlfJk+0ggHm0TivExo6u83qrAmVgoJs+CIA+gRK6oq0/r+l1kgM1BglM9
2df5TULXE9hddNbbm4EeertmDHhKyg1s5VZkquxu3F0yb6g+WgL26pwIdfOvbWBc
abXR05VHHPvehI8etCgzjC7Idj+NrWwzepww+a0LasdZ1f9KEijTbbXmV78OBsvO
fDfL9wO3/LrN3mtevvnYI+UGTonSUR1lSYOdE9gFrzDTdtJDsjawrMmiF+cAa3Oq
Pf2bJCFPpSTEBKrMsUbYKbjUDvn186qZQ/IX1oWnjHvgtKNexO1rpJ1jJtguG4z4
BF4r+NHJbDtGNYskYDPJsF3Lo/exJtyuDp2yBocuzkG1mqU12kCQ5XnBn9LzOfkj
nKrIFsCL8FQezot4t656B8GfobD84SdZrFVRkLWt9td/sLaYETlaChHxocH4vLwu
lebqLgmlBhEyyg0+EwLAIyrOzX06v4W4gaA39j9jFEMxPR9InYxCgsTr/vAiZG/q
JbBs6xWoUMia0A/NwDHsnTvyP/LjwcKEwoKWetJKolrNak9kbcHKqpGVjlOmUf/I
7ZNrDtf0I6p8PXTf8HbPZyAJMmyH5nCJOrAy1LEzPCjVCaC8UgFT07kKoOZfrvE5
aHdknA1PjD6PbjeURCOmsUQj7r/rWrPd1wYt8Y8WD/9+zsv+f35pQSf6qfBTbAAw
4OS0YsmtLTFGKWXTaMSTjHEdTb3qTXT3AJC20Uo1Fw75IyJppASL86aWywoPVr+8
ml+ABpCRVNSWme/sjpEKxSk+CocK/MDNPzZsw7FVW9gwkrT8EVfwPsfD1dWKnpWe
JKALko5BNJT4Ta5IUM0x+uPsuV1CAGaUKj0SR7vU8on3SwqxcoaP8tcJdKqLvuUH
+VSkpfziqF8YMsN+9fwRS0PuVU4ygXNeWkkZLGDAhBOP2vrbYB2LnOR0AabeFI6B
vcDABbVAdw3atwnMCGgqYj9a+y1F2rdl1bojsyfrZN/Wdc9Y4wCOIwTVvdq8w/DN
8R7K4EnKFzCmI/WIazupiArvg8XSv6HQP6uMY8YabVbsFdUtkcNCVR5yPgjxxKWb
ma++1lADurRdZcySTx3bcDDACfjNcgfeCJTxeD16AlunBSTYJxnIVCGsoxgkw+ai
lU2jAuKVGP2ofzAFiiJZTW+tAsGWNdxRi24nPkvFxfxdbgxUXXVF9YJfqUocv3ZR
Ys6GcGVNnVPkZRnWbOQ83iTxtZfBAWjD+jLMKH3izVI0TPMLxPMRd5UpUlBFnOrj
sy2sBSwKKPVJZHXxE+4d2+lPf6XXaCSXgSsukzvW/2I2lAmCQhFaW9sd1mlJBpBC
3y0vPOWNQ84CFhaGyLqNi/H+VPxKP6Omq5fSq7Ufk97klmKdIdSmqxHfbd1k/PVn
rkvCK7FA9P3Xdl+hacJ2pC/AddAoqa+MDdQlIcCDJnkdCyIn95+4YuQ1E5uEDgYY
VlUoBc3iRjn2smEM+dr5yrQqrsmy1kRcfFGlRJMmcgiERhwh2QliJSeZdTx4C5bW
KrKpofD5DhPojyV/ffsbdW0kEXGrpOKle8N9XwA2nwVPqd5fh8SPCzQiLO1O/Vf6
9RLNNahJ/qR2uddAuW7D6Z3VU4Riuhg+H+Bhvo+Adk0DtKGcLZcPZi4kvWsp6l2o
llSsniEYZdCkpz9VtBfJfSAaWTiBoMlBx10LPbt6+jMetZ9TCUiFpWx/oeoqcGKZ
K3wgVIp/5hAgyIi2oUsbiE2loWbLHboTKpW8fgprHLlVcngqWvjo2FbdsFkeGqaT
myhAf7CXChVeeYn6e075GzSY/5IBL5nfl8euD1/7F+EudjIUbO/azWi7dw3XAFUY
knUxK6lgMct+KEBysGxQeQpDh/rvYPtixeCKbRJp64U6hYz6sE5EcxlU2FGqFQZA
X+zLp391Ue2lLgB3RgtdTShxZ9/Y+SsJmqhazgcmBSY4fc8RDlL5qJRsJbd/ZaAE
3yfYQ3ZnYhGVD2GUUX2QNsvslNEC0t9MGPAt8rBpwvT9hDX5tQVXnYREW0oZq9v4
MDPPuI0pJ8DPGPIdxjgdbUBdX7pC2ZPkE2Fx/N9bmPsi4NqATma1+7DZBH9zzLEN
wkDEu6T27Uxpn4FzjD1vzmHIywh5CaEiICahuSzceAAG9S2g8SmSf9C8geMk4w8J
iHfatYdMbi1J4vJZDX0GWamnPSUVxbceE+qD9v6i1ufKyaDUKIWTUFm8wl5jh5oo
Kqz5DurMcHOtDj5L2DKBiH2gG6XALO0HkhcNyARtu/eCVlHz7YpxayPOuH/LFvM3
iBhUS3wzQgTrqUbG3e0F1rUSiknwUtIDfKbd8vwO8fKFRWi0Shp0tpxdPcqVzVie
EofvqBixaVOkvj1JUcIBJr9FHLtcsoZEAQ0CF9ZGg950Wtg3lfMv0UsNbuX3jTzc
k+CxbZYtWFo61rdbv8D4xjU8O5sgNOqgYw2/n7dqCXHzwFBisH6VtM4fhJjIT9EO
w2dfZPRIv9r6HS2qLzlbPU5rp1p9BrX2GQ75droo6/iegOYpt94WROQ10KKYR6rk
ayS2CsFC0zaTb0vG+YVHfDgyOE+5kDqsSex3NusNoy/R2AlwE7KylV1d627FFDuu
RuRJn9QGwPQ+6sNZw27erGCT3Wv/F2psaNhUZCJesMp/Uz5QAj+u3VnpBToSzbuz
yMf24zAqrnqC/+GQL3pm4i5/NdMBZxGB+D8lUx9PyBXewcy523vdiVe+LLpkuHsT
QB5zRXp8cb/Cv2T7Hb1hfQ2071t6mo+oGaxL9dcy1ZJ/qdQ9ODQfofAiRuagryaY
CGEe6/jEFFrgjC+Oq3eNUgjBUV7h0XbYc/m//qxOIK/w8mE+UiDRRHY9ThWB+fni
oTSiimiKMOytKw6+Ug3e1gxbSdroLF4SfWCdjFkvpb8MzsGOFkragJ9ki31JaVkm
Q9ic2bFfRwEMKnfQ6zyWwRqUbCGCeJFIAR1GNQB6u70jXQHSE6IuEPrH7HUVxn8I
1f2XLCYp64otW+mmqVL+Mn34F4fHLrC8Xk3uC2Py8WcxrhhTPE6ES1E/SCYFramd
PkEHtwUt5ZDAqtBGDCe9g6iXdPvDWF50F/gFMwhW2/jRed1mVC730XuARaBJk/y9
IkC/z0a0n/FzArcnex3g+E8qAfa48LOUcs7mGfjaGnR9SFNjFVlwmdK4jKboECt0
+P0q0XF52Rh6a4emzcPVfCWmJo+SJLEuHfVxNhrC/KKB/e/8EosLPfN6UU1cMqkq
itRcQxvDE73zG6VFbZazKtcrcfBvzng9NnOYD7ufjZWygjPXan9IQ4wtSfst4X9c
r6oVtOzbz3upenTHSyY8+apcaxcm5yycsQ/R+sU3c3Se+2VhwlysWU+LnBrxw7Mu
+0PwOj9u+20YXRTQHCeY/r0fbG4f2sCI9mhg9wlAasMvsq90d4siqNxPgAzPAN1b
BxxNj1/CM+AOT3upAmVStGpS9RJoAs0JoNCkYwuTwdj8gT0sw1JQ98D+myaigd1V
9meNxM0gX2+s0VGPVhLFj/IYg9LKdNPyKci99M3s4655NH9Y8HJEG/fBVA7GROiw
OeazmFmDg3aPo0vRH+uLcxXnFzQlABOP1VgYV6/PSJT/CIj1HimgXQIQJOBpYX5R
MOKS5RtGzN6x2A0GtUflfkXZsFVc/i/ZISbOBgkMLmNZUct+IJhSLhfJwmZAyLKb
DS1BD7qQk+JKSep6Z759edh5iiQK1Jx41ILBVlV563bSwUgen/c0fojTLFIc03e9
bv7fNKvf9aYcIKwndheQGzWJWu0Km6Ik6QP9sNwJvF1SlulHu2N3wVcoNGAERpi+
kE98+f9qx4xwxqYqXl06vyg3nyEmE+77JST5HBbJwXWRdmDs9JlSTdjclnlWirfb
y7RVD+swEmHUVFInFbmdptAx9KSAVLAOCJ74EQ2WlbtwqNnMrNJvPni3y89R805Q
NIzh0MuD0nAdV4QNwacN4gpxynwwSaush2w4QkEMZzxDPTQsD4jQra58iSTppduQ
LvE9w6aeKBQAxDXwrqM9joRkSHf5Qc/eUxbV+mRLvypGS5/plfYDdWl8NArOrCVX
OcXlUw1x9Auu06qFLpkgobr5bE0F4X52LzvTSj7Rwf9ofHCv//D2NSduYibhKPla
ZVJQaqe6KXIUO7Md+VDibe/WXcPGmyvTtYd3RN/qLUtsC3l3UJQTVbAwzScMoX0h
VRkUv9bY1clHtNArIztAzCZ+Sy7QVx1Vc3lBeqddP67yJ05TssfZ+MAZcR9e9K3/
9+VLRFAAQotNbdnfc1AMglcaiAIaeczmuC368w+vmZjSALtwxHYjbiMC6sR+EOTO
R6qi78F4V3s9am0YpiynM0oKTdwFxtsUpcj4ogjTz22tayylNVQ5Tp3r424jaPeu
jdZZtJi6Djjc1XJFdogCrZX7nyzDFjlQZA7cDOMmGr2/ALBBJPIZkRPf2gXliBFu
bCVW/GwmDEdEyDfYNfVIA0VOUSdalAv0D0YfhAc15mbbRjEi0y/uNj8oybd9xqjH
V1qPNLnbdhMjuX+uEGhZ405c0rxBtYHvBhFwr+1kaqzZGnJrcvLlB/LnQtQIaCHL
Allns2wkRgqRqUfUahlD3tjmG0i6ZsNMrVa7cPLz628wX53gmOgGCk2lmWpBflx6
bmpf3KjntkSeN5iwpfWP6jRuPGBOrPejOjjT2jiQx1MBZDsaFUUymG2d8YBtAaau
T4cbGwN3dygUsJgs97pZ3Q3/qKjuntXunSViiyC8YyfUaJDko/VKJyPMw7TG+mLe
KX2LBBRIPHbUo978aVVan9fo7+KfoAL29W8uik0Y/JeZUGXcnNqihALQnfKflbKq
LLYp2u3XHWZY3lqSfX5tfmAclJCoMKYRiUYEQNI5Bmmz0TxM78wm7xDONOL7Ym6x
knChCtU1awJwI3uOMGb62372bPEQMGBL2GUmyFDlb8Ubzy0tzTqEb+PClD6XHV12
yA+6g4zGU111ianw/bavBhqHKBu+on8f/nmhyNkKAvjpGE46Xj3MYNkAIfUrprHE
9CoYTAdiD7xI7aYNApZTaN5pV0gcp1eTDMI564+6GkjWiGYdr6Zjui8Z3LVmSH+a
aPgov1dE3rKyfjwydNTvtzXAnfmc/iRiDG6oI6clKTqKQG8zbCKP9thnz7GAPNsF
mSHOXPDvPaycN7lFIhAg2ANfCuw24ZPLSCKY7830UkxCBm+cTOrAg8RB0P/N3DOb
SYC6WKW/biohK04x+VlGvvWnHeXuYWGCtmw2EESXspwWrQqU7c1xrqtxHRbbdrBZ
7VkEHMj6uWkE+92Os9htNMLHZZ67rOrq/XOeirawEyeOMVMZhGIzii9wy0vjmRtk
TKO9SuX8gB5KNwJnynx1g1pN05Ts1O0oBoQSTqJZgjir26kQc4pYnJ7Dgxq0RKgV
aKBBr5Cs1ZM/tWXIbUak6udZHyXS2D9v1uGqVFvXJ2VrC/b55EcTVxGXVcqNlz1y
lNDoS/z90t07fIRwGppkjY5QlQbnIpIDVtSPF9PwzVHCYkEHpvzgJNma+v7VHtG1
8pVfUqIA5GK6UzZUu2ghy0wahQjxBF3GSLKnEztxO8wiz6SQIsZy6DtNw4MqOajx
KWLujSCok9p5CAa9wb4/jvShr976HTlCCEefan4rFOwQUrUarERBKeC940vcfU+B
7qp7xMrGTFpdCuO7fBqBOH9H5IaMGaBdNGS5aTf7vcmrOxS8oneEsnEGZMNLheod
rpRD9Y6ifrlIKrbWLgmF1ZeSQAavSJcS4se63Er+nXGCo2g/3mSA1WtvfsgYMzWH
T7c3yDC9Jc1vDbZJvanEbW3ArrT3p7bgljZ3RqEe+bYg7eKXtVWIz/VSB+O15q2E
TXfSVzsLFOypi+5/iURSI4U90sMN1MFSqAZyt1ah2EqJ2EBl+/69jeG7n7mom06R
dF2MO3ZcyH9AU6FtFhgp4bo4EBeQCkxYNh3QJKeunK8WCe8N/sjqt1mMRQtC4Cbh
ewi1HW9GtQYW5V1SnzWKyIjFbPxtOuPRWssQFSxAejSp/9gJYpFkaRK1ohG5UI7L
Kzbf8rZ4gXvVpzfdMtNElffhhRv5k7afmh43iBUqkRB3Pke0pyExF+3OrW+5N1tn
QMSInfC7nZFwuKzB8jF81eiAXBB0HZHVfKN7UCFYM27Fx+kW3jniU4L+gNgpAdCs
2ZWyNmbcnPAceDuyYzDmp6A6t5GOTSQ86PpZ766EPjJnBn+YKIYODNh7R6DNLa0u
OqvClDoVADwjIKEJ+RuHOGC4peBe2LVVVqfU2ZOnM6lVHkFpMMwiyCzNstsr5Qkj
UuOzSdfWXZu9jEIPL4nbeQmiziL2+ZvhDkYfeP/psrGJGa3OIhaoLirUOAAcH4X0
APpvkEzMrSxDLSskmSWvkoy5CwKJORjjafquQlw1NinQw9a2EG8y+WVDA6pA2fcV
ktZKGFzSI4u/jKJmcrJBiw6UiGuAOVeh6T5FHOVHiIvPnvwbhPVlzH1yLfHr/DKd
CiswDeYtLZqGF/4Wn04ZJZ8s4vFyMFx+Bbg+Q94gBJDPoWX5313zsWjBri7EgdZH
/JxJQ+HLKGHS+obtsol5llgf7C/VNjrTOogoK+pgtYck/qExRxJ/usfKCIYeIJ50
tfRJwmmdAhgqVeXwRTEI58oTuTOz1IS8+X96RxLZHAUzUYpUHlieeJgGcJ7XSr8e
L9GgADr0uQ/lL4HLTWbG1+IrLGeyQNlRc4FrrYWtMVmQeHVzwVuLu6kek4iqoi/U
G3WyPjxAh/n6691A+z6rmoL4MqdsaT/wd6Fx3sEuY4pAD5HQ3iDLfd0Ts1KKWM8k
eMoWDNJLm24QgOhBqhRA2gLNk74qxHmGY0MVOXYyjUspdOn5iByxvbnomy7b72sa
i7uUtWJs6YreCm1a6Wvc7z571TMH8nryndaa/HsHIRisNU0eDduIj37mbUwJXYRo
ZX2L2RxphYxJNSjD9YE3prfsfOfwNlYHxQjsCu0LCKL1t2kCn27n2cAOdztfH7pn
s1mHDlhlDelv16U314PV6mKrSRWiDxb6Fieh3yulsVwHblxx9k7r2xctEbUpB6Op
vqYiPwYak9ez9aEAMkPBOORltNBAXbXSjX0ayAZQ/rpvXqfKtuSP5z4Nq7dI+bh2
mOx1lvjvpxdDwcwXpXBpCfTwxvtTzOkVBEZB+9O7mP+HuM6i4tviv5IZwNG3RR1O
2s/YqkulXhyU3YszL3eO/gBldd4syxWWUhiklZl+Fgwj+SGGv4cUQV8/Ne3RRg1d
d2WWvKEyTMEEkF2YdDqjP1RSZUHpA9GANZYNxrD91X7Ux/ilQUiyDNv2iO8osrjx
PhOmTClJ1fKEtv7my5vWUtY/p7PWkwPusg9g3lQNOv0nDotLVMhyDyB/eX+AzJ8P
ZMdb+DeZSLJF23IOjHfi1wh8FIOuPmT8P9e3+lkkD+wcXwOhW/rMgh5dUjOLRq3k
UcfGJ79B6d6HG1mHBFa1XhoG413EojObk0Lt3puQxZD76y7tzSyWJ+PjdQc11Lcu
91dw/EBvqZluE3TjlZc5VXcsPWLkjKiHErJVTdeqsvl/ryr1hoIAn/Y3N3jlM5Z3
9LmnRlXy8hCEGKbUlO3sGU11T+tSF28vo67fNmruBXXS/dkIE+ku76Y5f4El/YIx
JtvzhuEeiTt3LahWPfILTVhklISdlhjM4Xo2S0ggUG9JTEIjGrAeekYemSx7bYyg
ooRsBGodOUdbbV+xnTMpeX/7DFONuBetBUdd+gLzXKRgbSrrwyUm9OblrHpT97GH
4nsF+wSG1qEbOs7VdIVwK+UtWZYdj35ev1EAG/EZCoeHU5BgXUATHv+h3TWoLvoZ
vDksEn1ha6jDL1HT3jvtffDOTSV2IljiKJ3nB7+wresKx0oIGjX3havq61G/xIrt
SDqvRMXnHwUybBIPASj9AnCk2ApqhQ3lIDedMFm9C2F4bYOQrVsGZPcWi7NQx4YI
8P1KumLFMZ3M14/CO6NHlqBoxd5MjFa++QWVAzvgPuhGxQMPpzpj/Rdky5BRex3B
GFNMdaaIJqpOlZbgJgeuqr/XMfS2JJ52kztV55oW8W8RbiiiO/aSsRbSl4esTN8G
5XQcQ/0Fa9Fdx3aR2h3m/uDNQG8rWK/EokOk9a+eavpsUzQ1Nm63agR3pZJ7Mom5
f+axg0hy8ApKMT9wnmTKcEC5pWicras5JNNqOmsLbKQr0S9UCj7gcAzyx0/cr7xp
+Ppn8jjVtPou08zsh/JcFMCNNvM5pxP9v+hzCcMTccxZ0wvTNHLoqz6rHwdTEdLS
HmBR5B2tYtPZFVRUo6Ez35WgHrTFQLmfLEkPwOeAHRKhX45vNi9S54zdOFoiKL0R
RgSWfkcsGNtq2SE2+BmAnoBnvOIJHR6T4/Uu5TE2E6/IS1age1M6OV5hKgnf0dY3
52F+GlZyh/9sxbWfPp8CTJNQ3qIKA4Tmuz6wJnO7rpjxu6v8qkY9QK5Wssb4HdRj
qUT60JshFzlzPPFVXS3T0MO7gKCLGqAzkEIrieqFH3hjHyUngGWchM25gL9PQP8P
3GtTiW+eCbYqMbae93DF4kA+qmlsp0oQmLWZ0pHXP8ZJzdWZTyNyM7ti7oCe1Usz
mQ6U7eyDSTvdnG5P/oRVhSkOscwy3tmTEo//tlun++YmllSZqKnm/buWFOOjT2rt
QJiUz0Pc5J7IB11geWz6GuuMZN4HJuoqUg8UNOZeVtnnq4hvGxSqSuaN99c4P+Tz
x2ZY/VSQoSASFM6CCkhzWEqxC5YYvNoJRL8qxDW3iskMD+vay++ucd8YOAq2IQgM
DBISGkktM+M+pxDmRkiT04wriXpRwcqhDwS6uH8s1t8jrv4I/bfYVwxH+xo5SsXN
Hl38PTzC1x0b9ofNaWJ+kTeZAM8JhAcWlnGDJGwY1y4HSczxfl6vl/Rt6hZu4oSI
kdHsitHMairth8Ydijui1Wnolk8s7ov7kue5J2K2etCs0eNhNutg/taTEWSWCbX7
k0EKPZFGzVTduS8tYWhY8rxZqW3UtmapPQy+g286e1tPFSAPZ+luNkf+LxPAZX+w
ERcCIVpDtUtjNTgmrafy5O+GInJwnT5qT/74nbVrSLdKJynSZKflqMZrjHHipWO/
oKf/OOuLf+M/Nf4Ba/+B2wQojgcRZo6FvI3ZVjjqXq7+gwptUKL1rbVIb/u/9vCI
mngMSZmFPgW8Tr+XrTk12BJWGIc5YOlsEIiCLO7ACsH2YmQ/rohk+gjP0U+bZ+x2
sIsmD6qdqAtePSRlVsEz39g72PIskXOsPZxdrxrsmvwfo+EgNbMsUUMVzsOqNfhu
oGWIbxvLqQ3bEdmqetGyKUlwL9kDejo5L3Z9M0u51rX7+cC7wzPD7+ULPmWIDwdb
ff1TIdGyuGjO20XJfL9SV8XT9YMQUUG0zcWgBpGBm0ZObpVv9KUmR54hirtRj2zu
fUMkhz56L4/kdVavvWzrRfJSQUK1d1gquPX0skuA7Xr6rszEaRh6v55ds2v4obRR
NYUbtl15u8fKPwSobktG8z+Zv9dEqpqHhM57x6cgNDMlnEJvu0Vr+9xPhd27TZmQ
a0WxTjxsrQeCLegyl3trKFvTvDOecXG5+JHReijEntebSYOxU9ipljLApGu626o2
JP28VylBAA8mKeR00kpC5PBkshzMAlUQJHI4BavemPnCRgOW+PTZ/Zxj1I4gvKfr
ay1wthPWJRhxKIpI4rvdZfDm1YiUxx5hYwUAcHBRKa75mxx3u7C6aI8OHqdKNF3t
W4I2aGjoW4gVN2j/+meSyig8dyNcjWQdGEbFNduzSnMal9G4qNhqI6fu4uv1SmL2
KD8Vm0TgM/FmqGlDjyvgciimgdGu4OZ2pBdL2MwHxBGDOjjJcYfVNujoelxA0hQe
w/Poc+bqBN6bQ2CcRTBs27TTDIE0DYIv44VsGDcLdwk62F6Hnimx9LpIk6xsGDEu
7Q/eHvXb8mfC4F6GyC+m7LjELrddV1W28/dTpA8aRhse1hKPZwBzH/nzcHaQRhaj
eS3cnvGisG7IIozm/WIZPUxU0DmoiuvmR9JH7ayrj0KkgKeZiev9oZmamsjTittv
XqnmdFPBfkIh1jeo2ECa9p11AIyyxO3kcX0J0qTF/QsBdvdIQz7CRbU+Lewa5ht2
DXE8bvzdoqlXYFezOTYtDgnO5LZ+zsw/z+BxA0crToeMSeRxCUJy2q0Tq8RyxQSK
vgem8xGSFtAT3RXpk+5HYEXLQqE80SWqd5puZvKnrFnYE6UOrCoMaUyWFwYBiedr
boQhI1Rb0ZGSfvZMcuRfzYHtXgtRmf3+C1HL0JpIpCF8QpQoHMz6x7iqxlIdStlV
TUl1f7Lz5qaNt/Rwu8mGgJqaDQo3buFTmT9asz3by2+0ZVkK8HvmKYSMcVKPF4Tm
5kUGLFAShuDMdDHPrbLsJNMUlSFq+unY9YjhVTWKxVmCsZH2b13HZwYvU1hY4DWL
uH15CPW0lJe/jRaLliCgfzx5lnwnbBhZM9LQQghqdDnsI3/dgxt2Dun/oxvc7ov4
f2FJtPUzgLKEl4ktqeI3/BqosqhcetMxx951GreNCUePZjbtcpchprNBiayyjiJ+
pb+6+GjnnwEkvNfzq6qVvFy/4hCpLoeZvoiKNAWg21d9+hW4PtoxdQJAEtwhhYJ/
zPDMK77dMCsL6EM9TFyTvWZKOSf94/Fc/qFKG1dB7o5lqwWELqbtdRIkUMJt1BIF
v1B9ihEGngIl+68KfTeAauOlTbhcPrTDXXqp3M8k+GMyRy41wXmXdOeifP+j0SQ0
F/zQnMt0H/9KDxBMSyWSlYJ1yxLNzcbVEGDm2CRjCkdtyCVg2RVnLmhmoYdqO5PU
jpUQeG/gawIVvwDZhZP5dwAgJTAYsWObo8HBwYoEtJvL/8x9UNWDDGTHjRwhNbAY
wG+feWRuvUhaJp8PQj9KDBIML2A5ZllMzP+yXIQi3WiSXQ9IjsHkD0zVKpevTgmC
4luWH4bdj6mnMFN7ZLgGoSRWfNnpSv9ff1n14swP3S+2LeW8EmRRkmk1iqogAyG7
n+7CxIn91qgGbFCGdqljkqEpP7gaWd6486leNigLe8GvAB/bcCvQYs+6S98TfYXf
4plY8s1BPbkmCq4DOpUV6aCUtnGOlE/HNM0I3WrtSSYHzQNQs+yNKKs+FKDcxmbd
Tye7mNwpQ6qrs5F8nXm8ceiPeF26lpf0pXHOvNxgotxE3sbm3zpf+JHf9R/O8f0M
qXPOQFqjGd/y+PW2fkEpXISUo+aZJ6N2aHLtzsebB7QLBX4jkBru8Nl9zZWtWgVR
npuveSsawlbCFADZG1HKeN4lMqyNUOwDBgToSQgm+arYSlSK4CNEgv/2sOWQl9Ay
ZoxyraTcurwVmhpCQbgqmjJESc3uWnxX9Teyp5WAc34x/b9wY4qFJGf2XuzAwu6r
SQecxRbKFfvaC3v0hJ8NW2AHfTSpQlW0HBweNswL3YflmEEApjg0ynsomCbOvr5h
tXjVWnJbDYylhcpAIUSsb0pjnSwUQHiIv/qJQDZxh76X7i6Oeh3lcxygARVjZzAV
QioZjdJB95CDMf7Cvb1f/hBlDC1Z8Py9J881kcliV/WtYb9ZR7RwSS5gti4jEkPp
8aMPBDJbNNaD61TrG16VR5NbKwsEYL4CdbMyY3PUWUGF3jxFtKHFQ0MrlRmtULbd
cNk4FWJ7F9b/zO1kw7bL+sfYGztms4JKWLKINYNFZXS6DqamGOuQGTF64c62pAyH
N2MNBgYtlcYZyTvIgwbTYZ7S5k8hDztRoqdJ5JyotLv5s74oZbWSzcN45ltMHUcP
0eiDl9BuxGO0y3nAErPL4J4MeX+2RiGG2CEjilCqCEzziTUzgRzd6vN2NqmNq6PI
TWjLAAU1CCGzjo/M2eZlAkfqVJfKr/OdjUfB+0xo8B3cWIzvPr5A7wmEWeqB6O6l
Vxgf0Ba17uiOUzng/CXrf6q9eu7bsR0AGRCfnuHYS20K45xT5IJM1naANqMbllZE
w1HTdZ6tzGv8LxVQp1LBBLtwq7lL0J6YZuWQfz8zJo322inxM5lAwGNcAKR639+e
dUPWzKarHM4yQL9c8oI2O0XnQeK+zeXXU2lBO6cCcKxaPRn0rH5NfKvGkT5N20nd
4rMYpZ9uVzvgBHaOsYMXjEHSr4seub91hxCWlIOtMyyrXqPhkoL/G2oLx3voi2nK
3wvDTrMExcBzHKbYfVQkoFafCGQC2DYkUzPmcxPHyimZW0ml/NjUXsA+KTgIf6ga
oLCwJi9hiHWeuk02d06Ccg03rDxsZ2GyxPqwmoeGyokBDRft6CV/fv5yRVJ77w96
FLftmtGJoF64+clbpmuK0YnycmHNdWv26x/AJLXh7AhYJQ9F+/zdVlef8AIJl4an
/TB0iw1I7iZh1SbhCRyB6JiOw9GR0bPGVMX8mMwbSl3IomOe8y5+T7x8ugeYXnz8
OTl3BpkVNClDy7kCQlfGOxTDiR/m+5HhTedKwLjatpcUr5mPbp1VzREona6/6p46
aVX/3669YPf94fdBmsTa6lrOL2oyS1CaRCEfU3VUZCkJQY/YHo7C3jv328N+ZLD8
P4BhXJgq0R1e87XfHT/S7WjObioQ9rv2YGK2W6nc4LF7lpUiPOvu6O0VrgPdjnyf
Qik8ghXr72/6jYC8KVCTUKsiZ2BxjqsvFwoH4zyVcakvaDiOzM1wr6uO029+D1wy
8hw7gdbc9vs1QtAWRlnQ3WcNzSQYXHpSN6HDXbcKZ1MCkgmGPH9dGRv5FEwdaAXH
nIY5Gh94vcLF7SU2kLjmwAEHZy4Sd0pGbZsJIWzulVCTp07P2Guzs73UR2m54vSa
Lcsx3uNVuegAMLCcnthQhtBCG3iE+INEb3D/ChOsXJqlaONCrbTH87GAfWUibXFd
oal6QIin8G/rQdAYWW9xlxbuRNB2+7QY56cvhBOTOEJ45z8LDGHl9VSyIIRww60V
F8sFHVx8trR0lc2q8WtuxiQTJtz4ilcZ+FxAluaqj8Gk5igbSXt/vYuwnvk77aB/
SmoWC+/Y7XAFQXsAjuDpr0axxKgNhtKBppLF3S2+I1M9mQCrsSDyOofMIr6LWXFj
Nz/eEoAiqdpT48MeN6EbN728lHmY7/pfGKdNDk061m7kALWYaSOAedZ8+MJ/5gwn
357fhRksu6PHlajkDtMXbbQZke+1NWtKCqGrUifnA8Wh4CEkid+C9mWRFIAuYxw9
UqyJvTWvUA3D1Q7YEqqJmsOL4eNXAqIpJguNaB+4bCxNq8KtBfqYHFJSTAnJ/4gi
wgHkw6RqxGtPhJzzClD1GR8TEPKHtSn3K8SOPF0Dj/TLCZYo4VI0CaInaKC7hXJJ
mp7sVyssCW6a30peDe9sdPbJe2SRkXzoiyHtjgmkyfrXuo9PKm+BrIQRyXopSbkJ
PZfnxYbFE2VAimAnhAYgog0QhrLB/rmyoaqTADHGnN7bJ9uLTat4I7Q4jn71y3QZ
OUC/Hy1zXb1J1yivkEqqZPDJpt+C5nPbXU0SiW7RmEN63crKwb4GrmAyTiWFXkR1
ExzXTQfmd094A5DBSP2/M5LgpAG5rrF+2PNZMpy7/E8D45Hi7KUzh4Q2bRD5USEz
mVUDGTUPYN9PGSF98XMR4ZZ769WK+O4ThaWPHmXOAwbM79NFpEBmBkVmdxzeAcY0
Y+T+Q/2ps8Gg3xFfOXx4XJpFw41gtnkexaWap+gkIZoZCRlY21mvsU2Ry2XOAut4
w6kRfomB/2eJX6Df85IDrziwex3BtDJ3Zx/c/8gQo/Fk1WDJ83riPJhuODEPCojp
YQI+jJyz2mfM6ZnVm6yAcH18+QfG8gKUCEO5JlhmCe2UK+X5c5lgPYAmrVrUX6H/
VPN+d71kVoejHKOj3XW1dNnt2hjzapPdcE5Qg95Wtg1VteNHb+ki7fbzjR/KGUIC
stm8rJsDKaC+cZZocC0vEBRqdtgtXAugsx0fKxiTrN4YjEDYRBT+wCf/+js+01KE
Yfax4bN9zWEWLOZf2tcB0dNDHNcuEzn5kJh6kf3tFylolsW6xfQm7GqLrPim22VP
Y6qYXvwhk/nt7lqQdHilm1Vgd/kvzdYL2aVql+z3JG/yXjxyWlcxZ2M5+T11Qab9
eCrvzpH09er9qUytkzqGZvTPKJOo3hUW7zMj2OcqcFlE08PlWse3PN7o8mqSHuve
XofCT+BnZRncTF//C1dFtJsMkNDTaq2VYL/M8vYGju7555hjAeHzM7/TS6mRY4oI
r6P2jt88Kjfwt0KKUl2ekZ2vbUT4cmC8SSIOv0pATIrEPe0HXTb1PLh+wKBTtST/
8r7vsWpKNw49LTqd6dnXVRsS8jRJ+sfJlH+e6GWx03YfUVfJXzEzR57k0mjY4OeW
0zhbzmRhUWxJLTlbT8Vtnpr7NhqcpHQ2dVHeML4ibC5zq2+qj8DfDSDRUsYxQEE+
Tcqerwszi0owPmUwREdZY26pzq/9qgQL4Gh7RBBTccnUwB9Jc2B8sYfT2A1K7nq1
Y31RdGO9hr/EisJQYJjdjPha+kpTHFI2vBM7WAMRRe74DuRJPQ3XBAXoVYLyQtPx
BVm2Nnl6X+hnUtK/xGo75MdKXoIRW8cggNX0OCexTnkC8tvwJLB/EERjtUm5DHf4
aIhjoFsfC5YPROvDNyCQdz28hNZV4Zmz+F9m6KZ6PilRskaCxlANudUY2VsmIhpE
W3XLkjfBLr7HWVU0sH+0B4MH9JRjwcAxYkbfqS74aBT5wXv8aFn0VSbZ+9+99Bu/
jhvMWdBpAqXJWncwM6U0lFzm/qCfm5KrLo0BrBUJLnHMkUyfk3gTxAMb9y/pwe4Z
eD72Sm7n8QhFl3xwJWT4YiD5gnA9mAw1FCaEU1xoynN1zbCzKlvIUJqgi6fshcVr
8si2cTtRW3c1jkgfB+Qr7hTeahvOZXOI1HyZmybPN9Z8uqsRdRG5mlk18e/B/71n
fBlilYGe4gi2KGX+sP0g6TAJjj0kZW1TjhK/CNGQinczzwKeGflxJ7mkwhMLlIE1
lX8+3GPQq9+gTyef01ED62bADbc/5IroNJdvm4MjY2rxFfVWimqkLyu24OHJ80sT
62PGqKBA7W0HH/2BxCe5wKInMBSNPi9LHPqSFYvzhZrovG41r6DPqwrNT182ssGw
36NyxRPm8Cz9DYFJkvQ8O2EkIM26bEimLKLVFbvjTV1R1bDvuG/nQ05f0+skqCpK
kuANBfdp4NF/n/HLiwDfhUiDicE6KV0BaO45AbdYqOupPQtsc3VIQ0GtPt73rYoD
zGtbTWX82dFN91N0yKIDOYBGG8PoGY6ztjC652Acsg0uvOtciy/Qs3NuAZ5b11sW
aC5ySJxOEm4aaBHIlLhG+5ELq9sz1E1ToxD8tnc3iLASK/8YSh1anIfJzLWA9BMh
+5GFB7oOsffm1OPgNjLTvBJmkyGLoNvzX+Tgh5TdQzLaOU3RIMInpVs+RHoaB3d/
yducDKXTum0s3nFuImMbDPFZieSzg8tp/s/KzT0WAuwQLAQ8KGPi1Pc6OdLaDMUJ
a+kwffsTh6YWHHWLkvhCCxG/IQbhggKr/wJVOfM63d9mZGVk0YxJEF+oVIR6wzFK
Ax7N9hw3CVttA0oqZoTTglrISfXT99GvbTY+NAkfLZu+CZ23mT7yzlRXeOCtvnTc
oB9nkSDaGyUQ+v196jk0vxNFcjBmwwaHyDOOTv0Vtltpt3ubvRGOoMTfdf+InjEd
qzupIsVaAru8UuGpd05FEoY1qMw60VAHNa4o90TGhSk0oxxmPbHYn/dTHMGV36nQ
4tBAoBCPODSQuqLu9NQM/kLi9e+5AjS75shUY1k30+9Pm6kwAJVCgnmcn6ccYu7G
IXrEwtcOkn3ozgbGdwKfV1lYpq2VO9cQ8UABREqUdyVG7Qh+O/kC8EBtR+Amn13C
T/afkw2/L+58qGCwI7u7I0GSHBe/vi9KSjgAL/KoRPbtSHNo0FGRKBMwYxE8vpPR
C/GEEsZInS7yiiXwN96dEDgKbATBHXTgSGVRYcVwAkeb8ro4NzuuLZl3/OgGgZom
jrSlPvGAg+gt/9eh7UIh7zhV69zJk9tNMItZsIWKEpAv1iWsyVisGNpUgoNd9rok
w860ub8VBqWONWN4N75Vex2ogop5jHVGEDQn/3yZHk7F/KazFnFrl5VGhP9BUNlv
+D4faY8reHm0vnuv2X9CEanW8guo3qGZVbhDd5RaoX7xbZ7T/xHVwDfDJbYAQkbQ
FM2P1BmSNSkbt0Tseyj9p3jkvRMwJ7pTwJLBU6/raHIzrGbStkWtQ1eeRaoVyBWh
jt9V8FPPRnTAncAjJ0XFjefvFitiLzOf8fS6D/e2E9T8GTwNrvAsOI+hUSRSa6kM
g/NngSw88VtzA9YpZ7OvKLWpOcyB3jZfEG2nW8CsOX5klVPkLuT+FY7iMlkVVmiW
MdyHLIpVDA6V2XNFe8tu0yf9fBl6ruMcHvYt98TSyjmLfqgyAzfXEUPtAJ5lSDJK
Oi4kU3UdbJOgeN8zV7ePW2lZ7nC85kdE14NgTDSjZHQrfXXHD5reiZl9KeZZ6B9y
9y5Tr2pTc04Ej6ZGFVovh0FJcj5GKTMr3Gt5UoL5IAsWML0J5NdCar+T9ojKUK0T
2Xk/Q/BicXwslh1XTmoulmVKY/GNwbhFfPnDI8B5eqT44faznQH10S5BNFlp+cwL
vECee8FkoyqDqdjLpJfHXB8Vy6ho4OIdYtumILMdYjUse1APYxMVqWgpHi5dn3be
SfW7Ux+oSwbF5dIUyF1qKFzLh2jNUEnXeAPak/NU0gPzboBknsYOO+aVxt/N56SN
EIMvdiqTz3UBMUW8/hY3J3XMqDaFmRdpYzj/j0mtR5h/bNDSuL9uCnrPC9Wr+4nk
EHo0jkIs0poVV76qhDA4cMCYfKU/t3A2Fnxa8I2JLW0iG1gLAMqU4bkVmUu4+g2g
Y2cSSmja2Da9y0wtnGH8QsITscU1iln05+bNE/LutlfqOKHp1L10OeTtvenaMIEg
FiWtqWoP6wlbxfihl5+CRjE/VWsgCoY5BamFGRHMdqhU87C8kxmC7ZVYVrq2gOJ3
cmfVQedamVxjIlvD26DehnSLE1+ObGf8SwMbQt0Dc6zR6mv8dvskSGUaTS6RKo/l
uGbka/sl43GONoTQBdyq9AYyefm2puCUSZmUP+Uq51+TZ/7dHI8pW2vIDaqPzo4P
AXfz9DRlc5f6FoevvbaG0xbMAJ9mP9yjU564TGKLLZ3Fpgip9Ns79Ip7GNryTbsz
VJTVKGGqWqUBtzXbGWNDUepVcYcpgWDuAIpqqSMC5/hx0/X+gY3D3sGOGjkZ6HZn
0KpRPuN/V3J2pbU5Hpv1TICxXAlFK8sZ6SUGAZG7GnTS791V/kt/J0KA8sK8BHbl
a2T8VcTp3nI5xqQETupyaPqef0CaYJOzacq0hErtBwPc5U2PW5IermXoqlqRLMci
FFpNQZiAvvYB0x8Qf+YJu8s8ti5rY5tTFK9/Jol1VIMe911WJVw2iOSMiUaTeQ+k
9LtlpSHd+hs4bCn7DjyCOSrysG2ZHzdPApMvesJGx938pBmxqzWP27qN5DRJ3Q4h
LhKPKnDc5QZLLjiCk9f40LlDIB3dKI3/mAEu7nszR2jCEzqJq4mExWQ/uXNBU5+I
OSv4q9nBD4HAFScg3jGz5pvj51BgB50j/jlIZQ3uBvVyPMZ3qBW7yfy38GgyBW4W
/3jok+YWzg2fXmNLMbFbK1WvxlfAvrMXZP+NMXdHBuGL0IGXBGIcl77TyhNCI1GJ
hSOdJysFYjwZBlIDYNIgSy3O18XrTRFYwZ3F6MGIh1P5tSNVqiM3cnGLDgd9kAOG
DhXrL+UzO8QNJRx2jvZbM4SZh+BRPybfjGAz6oWOpOybD1ob6p7VCbqZwFRIekkg
1tVkw+MiX71pvn8f/klSBBg4OgIztF5FwT4/Q9HM4Wo++1mFDpCMPA+eAAXSjyEl
9dazUcVTkjXBmc2s/uo90PqZ7SouOI6vb6Wb6/8EC4jj1021tAfA2q2rFXWEynEO
UtVPl1ygGz5YsJrR13AaDEJK7Bde9IMcYOK7e0av6891MzxtM9fonJRYCXpkeLXz
nkaxfjSdDdlLfmKxnkjK8sEj1mdTkPvXeWemAo+YihSUX0Vw3toakQH/oYx9FgLT
nrDqN7CWk8ZyYSTjKPHx6dz70nzgNniQNOz+JBkK+PLuco//Dj1buYIRe5KKEpff
+q06phunVDmWeVXVs/lFRHVLi3T1YxenwN1xuTmXdWHyESBI2ybvBLfqLw85xb+p
m0JUsb7tCPoWylNIUF70uEP5i06tKb49KDcDxf+Goncy5q/BPC73y51uBcea8pn4
Wz2Qfd+kdBq3nXGaK4lE34Wt/UR8VQYSk1vhv8NLzDXG7Iu6wr7NM89NAPmEIzaC
miFWCvoqFX6Y59q19U0e8CCFPwhMtoa9hWtBJteU7KdZi2qP3fkjTvasChXmeDpw
zKCybOps+Gsnl0Ow7fRn1zqx4W8zwAaEb9Kuj+s27a5P7RFukX+X6x4INfNhFei3
+g+MhoonXAIXn7K5rSt75jLhjNSc5NuMSagjbp/bK+4LmflRc+kONlysw1gr/jAB
NtUqWIR6HvRol/JaYhjQoueA6kV4TV3kSiBNIJgQI3IHwxpI9S9fvY+3tUpfTdss
Y6lgOhrbFCTpYZ8PPEBK8vuKg4vUgwQK7vDcKGvgyxMvTdMYYDqPjYFzqWsEzOZr
FAiuz2ifg0cp7SEcTpxL6CAJ6YoxKEdG4pOyn/AtDfBaM+nmPtuThI2mTzAFGCZ9
wPzX07Cj/jwQUdsDkVVC/PtGXLcs8+iZ+cqF7O+XSA/8W/DXE3g78iNSiaHf1o/m
Xz8tEtwZnVu8D/vwPXizg4/PKUceYJw+qjs9uE5K5wdDBsAQGm2TVKvDhfHxeUkB
NItaqstpSpRKdO0n2SZzRfgiwd3aKH4dPPgWv8FPN8Cjso0GapjPYjOP4kASMN6p
PycSS4mvhQWpiXw2d2p81bYExP00gYoVZoPwFgwTKKUA9qF0Wrv7tqlQpb0amSYP
AZ4e7H8B5iQ234KYA/W6Do5nRGgX0AoRDonPhYlXwMnVtSi7PIhnVwNhQv35X8s4
lYbLt97cD+GwD8IhE2cCfHWHE5ANCGwR/vqv117Lt2qot0hBouWrcRy2qbQHOsX+
2UMblAAiOSqbFLD8H2PgMuNNy72pQonaX8OaIExhLV1zyPb32ZspnI5okUr63cp5
gIKq3SiYWWs1FhbjgCnG9unhyrC9F0eKOo6EYPHfjKlHdqDFdIgEEWk7+aWUAtkr
NVDAkSm4RZJmdCm3r4qvuUeTscm5EybQS10RhzPwOPUr2teyqr/EvjGwD5tGteCd
FlJ6S78CPbpURqJbTxVHWwkMSSqa8LVJk/7Z5cVyjDUahMBikM+9dbAOGxn/TfK8
NIIYokcA/T1sJrtro9vyahwE+m+1DwgsJKUalrWetGnf1T2RPU/fO2y7Xc+BpEFD
ZYxaK3IhHZRG7gzp3+ldCkPLcwXGdoHuRP9yeLeodixi6labspoeX7kX7Er9e5FQ
flpU9qJvBxoqYsKbj5uic671O3m63Eet31I5oPZKLDxuSLVmEZkWoRnfc1yHBMqF
2eJcXeQSK4jFvd0SULMpHghQF9igVkP1iUqvvuXXVHb3m/EMWK0JJHEwNg0cafYl
RfCZz93WmVykZprdTaQkVYP3GECVexPdlyGNIay0cYl2XkxdXTq1WTNXhaEgQ49F
bJnrV8o68DtS9hCLpOAGBHYYAoyplb/WrjPcVtMcTeM6zfaJPpIVao72C2K6y7iy
8tGulvMNsDkkzD9fk6jxw84TrxDmIvTfq/Kh8KBMg8nXO5QUTUxOYunPy4zTbtBI
2Be4/urpFIvA02G3xzaawdTHMbJBWK99G4C410gT+tIR1iza1OpP8Kc0vewE9feV
gT0n6mlgDVf/LQdgcScVx8slQGPxXsEf4Fknx3kJmZFZdEUjfcH18GuHayjZV8bj
7L2ru0mQ4mxf85PiX9np6cFP094nci16JIJmHTvhe/u0W8ZP19gBZeTorfAqjlMz
xdSVjBAM9z/uI2aHxmFi+RZIf+IIhGoI35IMqXAwlY84tjAXi41nIw5hlIZ47eAm
pwwHopHf3AwS48KN1Thjui2aUZJuBRKoneTcplK1q9d66ZreYgk7j5srW/f0zGvi
5nNIO2l0zbSNJGI46CXP7xiftfMwsPMJeW7ru6FTE79TXIbhu9Axs622ChJV0rDs
3quC/bziBvtsSnvqVpUrrscBmOvHhheOIddpi9KnSW+bTcHu5PkpzHfpl4/kxo+u
BmigB9RfSfhNVtu4dIbz0L3ZJN6lHfIBXbbwK7KGeO6jqBoliDdoAyaSVI3udS5S
aAv7xiuAYeM4aPRW0WD7X/m7BA3QoStT3QucnjjLfb26ms1Or0n5gs+Z8OhsC/nB
AtmZxIA45qKNJrgcYNWMRWkiGX11Y+Fea17pfB1uBXe21ytvGmYH+nsQn55HlohN
8iB5b9RXliH8lL8EuoeP7/ynloryD7EaO+5TNojTo5M3GKo3PLQvSDg2dPZvnrpq
htgGRr60WQHB3Yc+c7SlLtQ3K7RGCVAnOJsi45XrU3a5zd8pveoBC6sSTaHhtigE
VU0j0GBgbMlZytAcz95cvRR/r3xps6wfr/E5yNv40AUEttzmp80qXy5vwdP8ncDG
GtLi8Pw6/6j4NxYX6LkXRmBa4seHFeO8helGe54yeDbH9OnmqwjB0X8ee8ZUI7YA
PyNHvC84ZS/i8AS22luKhTY1BRd3wr3aAlK8x94taqc0gVlaZN7ilX7nv6YpguWw
sCksNWe5DDu3FVTZHS6CFjTY3HzLvkBbmst9bwNjDUqE9xB7das2Y3HmjQV2SWjY
0b14vFmz9t4Snu+Y3aVeJxGp+dkAUUeJklPHWhyUCDTnWz6yn6keprM40mOrcxa8
2I0OSGu9X7/jws6XoIsW7xUorMF8/TJnF+RwNg/dnhbmwR0RTEP9/FU0wleZXbui
ibez0hZtSqVmYrWdduTjZcxIecOWVonjUg4H48K8X6XqG7jcCaRypdTX3GxhjzVv
GWzfi6cza/pw/DrQv3tE3qg9bh3r55eBPH1GdkS/dUh0tbIGNwbT1/Wdd91ay9rA
lej6mNXx+cmJ1yFG2j8htk3GoKyC9OZArddjzj04OYwJdw7iqVxMqXEcV31chjsm
FCvQCEVRzJfy7BS1qkB6wHmiKsNehC7Mg/SDsXbZlySfxyFwMV0IXdhK/1KPr7RS
9Sy078efRwkYy2J97plqnm/wrHRLFMlSPDKb2vw0pT8WQ+Aiy8QQ3PmOLtC5pVFs
5cOqYj35Q8g2rk0EKiqswJlTkdJTLLgeS59HzoGtDwiEmsNqmPb9/syOBgZdjECj
2YSgVBZ2YQWvFFUClv7psiJPMMwqEpy3YKgZgovTML7wY0RK+BQMcpcBS2hapwcQ
2pEupkwfK6eu9Lvgy3T1DUnSqPggXIsJ9HBKHG+vQn6Vs9ubinK4TJNo+wXN0mrs
I1PbuyocxlGcWdb+794BVtU0igWVKh52lQzjMBlCql2he4YSNbVIm/fFXGu0J4NI
du/xuLEyAOUrj9XishFdDQW1F/ZbRgNm7WgAN+DL3fQLEk1+YLvme+dboIBmNEY5
eJLijkNh+aRwEk+/cSvtp7JPdyLyhnl0oxGz2cGJoD7swaDCIkV7dPoVAr+RHoLI
dqg0/R2jJWZYZTLLuNK0vzyqF+cLZNDcJImwZosY/+jYBD1NKIxscaxgFXDa4Vco
KMP6sCz/qX6q+lEpg45iXnHVUtDqcXvXE0Ojbz/qU5oLWAAadq4uzqkoC7cAzWWa
C31qePQD7S4t+bHiTdjSsI1JD2zdwJkCDBCPwRReuHbPjTUPYNucLhoThAszviSQ
JlvQmPToNJIM4CIu0m94lOnQ42+6ldDx7rVpsiHm4VNFm1oJQsaF7OLZCtDrgRML
Ak7EV9bxnPi1TXsqTotUPe0P+7OpXoPQdkgChA4/remQ6xUBVY5FnRy5bmN3gCpR
erx1Kg9sbR01AY/us59milKa6motzwskDe4yPrBlZkLlIBIbGWr8ZV2PCUD4DDl8
yZYeoaeuHWcYhGmq7JejlelVeWH9PiCsS905ts8vDnubhL1MKzuX5kaN52TWujcR
6qXj0fsNdsjaJhwUSw8YUA+T874NHJxdct7HC2OZd+WB/RmMiMNZT0GQnxOgZpkV
6oO8MGQVhG2Xeo2uz6jW+yySknY8IQoSFW9S4/RnK8YuMy/fXWdjlI4A8Hkfelup
g8wgq/RVBwDqzdTaV9ejKXDW8FonLeAzXqnqIvPfTJy3sFki3kzuVn1iMvHbt+UC
8Fukg+WbPTUkZ0FRJcpzFtum62Z5Q6P7pNBwfSOBb3gVgeUXd3jOJ+4XCeVgddDa
wQGxUVsxT2prPVY16ZarEvqL7X4G4g3M4jJRATcO2MKytI2j3+0pSt6Qlw9w+r/w
4PNTlbtLXzsBjSbq9ir349lYBsvv55h/XyMueuHNOE3O7TSD5oYDeCM7ts3LCM8g
aWAnKSx5QgsRwLxo9k11NbbfoKBP//wmWZOBjP5bxDDnHbwnyd4vjxkwX1lpqpZ5
IQYmtU/ipCllTBfYooAWRT7ziRrd1x+bZdTs7aKM+XRDgsCWbAj/ZHXqZUZOFQtn
supcmPdXVrFawq9Q1DtPB8T+/Mn0uxJXP7+plI1AeZN5GvRSvnTgAKnY6woYTsVp
xRuAxcv1tE8vjJ78urQhSam7KGmLC1NpTVSY7cFFayXC11pOa/1kHbdiS63jI+eH
s+5XH91fiIk168vxgF5bGoGFf0aMOE6yFfJuUroLy8NWYbFyIyx25DqWjcUKmjYp
icWIKe8x/o79aQLDCub1+4RtjS/FCzoAQrHE2/FZFXjFGZkfN/JM5crhtfr8wKzU
V4/TsqZYJ90k4dfDz7KVebnD15TlxgxTZgyV65ase7g8zWTGymYEN8tAG/Ev94Xf
00+iLg4s4s/MVKBn1VHapGY60AijQE3YcfMaAL4Nk1hMH5TE3x8/15D6Ys0usA1M
2fKwJT7L5DQLo3QpQ6Lss66jBTmsdi5j8OkJL8vil7+xyUNv3XTn8kaZBRvNZZgy
O1IJHzcGK10jWwYUo2j2rYTIFise+sC3DrGpKjqH7LkzE3bCHIgGQLbvsfK5m12u
LqtMRlP2tjP1eumunnIxGNTQGeV43gftdV2Q12XV34bJnhpHxSTnWLhNJgDtCbAH
VHdFNigAAWoYD8y1FjBIi3SzYcRB/TT8VWcvo8rpgs1OohWI9Rtzl6So6KbEELSn
PyHPX6qPLlbzSrfwuzP/htGuq3/zA3At8vNlK+UEFolZTPoqRX3KlyXubNKRSXAE
5Fy4g7OEddHoJiierbFC8v+Q5opA4xGyfjnDQQezi2cgTMuVBm1/ifn4+8oF1ct/
M5gMQfwvz2c3K0HLX9PavnpAvGtdAooXW8TMVkBDbCuxfzP3cgtWmD++GwWqPOLm
paYZ+7xdhg2yKOPq3g9/TQE/5M8HDnQLfx5YHywc3h9Mza609DT5F72p3h36Vq9d
H/go2O3apKDHm9+xVMAj4Ggec+Xlm9YbTGA6VSltDQeBvWcpiSabI52Pnq6+KziU
ikPjO0ghcV2UdVrEEqyRrwLSMBax0qttCTuuFEmRirwEEDnTzpQmolE4rtTC1YNQ
LBYgAEOqjmKb9QouSYrcB0QJNX4Xt8suklKhitM0UocGyMtDKHawTr6vkg7GdZ8H
5LZbnLiw4RFYjBN0T3Pp/xoY+flksB6L6aPGUH/jzovxMzSwuXOJFE9Fv+/KHSiz
wbVE2hpNHpPerRk2i2wtWByZU5nRLSAAetBxz+hgINdlAMNyCmH1eVGB5QFU1qYf
QxGQn5l46uEURXzaUKEjgvCaPKNvRWFoHYkQ1IDumTH+LaKXbuxtTCKA6uUkqwih
/BxIpQ5NO2Q4wiy1Be0k9gihE0LvuhtahKKPVTSsn9IElsqhbiYy0476Vq3IY2Rv
xxupEIHtZtEAHtCtMDwhKVJWejFvbO2xwf5jsRwO+lLZWheS44xAtywuyGbU9l5m
XkUDnjAznJv7Jl2WBYbv077lgqSGfU37Pt/7BIJgvR3oJM9pbj9wW3TVgRaqDyfc
vKlz6kc5G4hhPgtjO4ABVhMa5A+RvTdk+KLcs62ZrAZ/RRvF7EGo3FgICeG2Jirq
f7SBaoNHBsOMhglLUBnRqQU730tlOx02lwW6x1FjJJatA0WV5DN8WUx/X0DnqCkq
ekttl2GoLpQDJmJqWf+O8qVPA8MZ3uPuXd5unsByityN/LAiHCeLt/cXgTR4TP5+
Y1KTCTEV2RDoZpKOsSrMBkpRnX9HI2PRzyBJb54iLOWoG0YGVOg2DMrbZZ+OCA+w
Mh1Q/bL+TGeauMbXH/lcMrM3bT8kLtuBR4aIE4iSWHC9EmpiHOIwGcGHhUJ/xyDo
8yl09QAW5wUMXuuQ4fKXOhBLENiv1IiS7PDs3JEBUamiJD0cRii3HJCKYIZUuU8Y
5ZDZeJF2uS8Z+s1o9uSlvZNPJoPWmtuGTl8620P3Q9OCmlf/xW7sQM0LvngMcN0/
ItDCSg2OX13I+W2S8jFVQXyr7Dtxh1K601bQ8dLrvygWhGw+tFC6MlG/na33ADQ/
iuFtc3uld2NcvM5pLMX/NQ+5oDEOQRPynfeNWKmFqcQxh+uqXG+iCxPbIE5b9H5d
OWJo1ZOYX0Cmpk6mksS7dZ2uRVrpSJa7XKrK44f81yMn+nT4Dmjn70ws7O4z+ANY
GLSG8PCSzQcQvX9faD6vRgfVkT2DffYj18AlALMssi0n2BXlCX/nRbtKaivnrxSB
oyz31uGX9lhQ46avvyxRvYTpNDIm9xQnDSAErHijSDSzIPPX6yyRWT0VGu3BEEGf
yDdGKB7F/8/J+WgDaq/OOH41ScHu96WqUUeJzlqEupHDiHEF3QwJ3lDCRstVDWgd
7E/z96UjdIAHHpxiOlewwbxfJwgley0TrTxBcl1TIW2hg3esDDORKYFXb9e2dy5y
LHifiqMoBAPp9ndkN6s5U7miDYg3mscAOj39eLcBuikAD23SqDBNJSWT2NUzNEZ4
mjHeje5Tox7rxxc4ybj5YKl5HV4JWccJ8DokZAnDqAp69i3X3spXdXQvZ/lHasPJ
w7k0ZDvCDNwhkE2s8hg9Hwzb2JjKFv0Nw9xVpNkIrrHzsNGSYcRtdRXX4zQajLf6
r+U934iLuQ4r11AHt9NWsRwuBhdYraYIdKG6RrJwDmqr2Oy3aMM9g1IXpsj9ZwUq
3cVtwV/TPT+8OeeWLqXrY3oKzp2cb4fgD/kAt9stR+2ewoDw0w4zIaEOUdOKhzJA
Ny+5xUHmJ4JCPrmTjRfO1L2O/leH9yLK1dZpAfermKB2qiYHeQTf07wBpYGsgnWQ
2bAq8pJauyrC0XMYJLyD4KJsK2DdMz69rEmPSIvdqaQE7SCvB261ecuGgD197fzr
cIRje8t4IRVKuEXz9bVqLVvONFdLRDrQJLLKQ7AhBWZJlhWrJr8Jh2xwrjRdGrL2
41vI9DQVUzQRRYRIyrdqi0hnOtk30VolSzbtPW63ce57VOBy7CRXPKBvA4dfLYIZ
6eJyHvZefbuG3zLD/Jz/PIGg/2e2bg+GIgto3Rp/S1LH9ikFpnrR1MElGBeoasBK
tIUr47t9k/zmuRcEd+j+Zw09KeXnI6wGGbD3x/nUuHzqFowASwWTMU5e1aoG6rIy
Tpk5C3EhbJXLm72/Aqis/hkHZkQBJ4jwVCFkmRuYEv8PMqkJZgwhm0EKplO268dA
uf3q4oTpeF5k2JUS5Zp9N6Uyuikomo6hjcI17H56jA8RCOqnNXgme6XgKhENKuQu
Vzzk/VSwV9gASQN3b7emShVp1TGQch0uanpBKrDCIemyAf90WNa1zAkBwiTcifvh
BnH0HETdXv79b/M7Iygm6QoFhsQVl+PAny7lLPJuQEI2ypdfbv29iw9Hb2ZOqwJB
05K9w189CzzwgyLu9LwcKp8xaiKO6dT9hrd8mYysTRtDkVyhOuwWvlKXAYC7fbBS
K+I17cgTAHfA+jVll9vxyzhi/uPQIanctsEWyiv1LdDSt9y5RQZ4lMiSs8Js7qqe
h3wFgiWgcwIBRDMW4dqYcxpFXUrTV30Gky7aLQdL+PFRYU5CsxJlAuN7US24THJ8
ZPllS/wqlh3W/TuJu98zlAFoCuUvY0nqOUxzS1B3ZwDmjrXlPnAKHSNhNefVCXK1
BQBRTh+mvhSbDAAahOx8sayziM9cGDznzinqUCiuyx+otFSd3aRRDp9gL4RX8O9c
H/UDgDK3LREe3uHc2uilbALTHeV/WofkUng8hEK4etezw2UClneUocxRezQ7MbTV
lozIFWpqHTuhRm5xITMCP12dmiZBJiRSMsM/TS2hmi62n+3RolROvNobu3/s8oZw
hal9UfUdSluq9ic04fhnzR2Zqlv9d1+6uQrfr0DZ9Lys9JTKKhKMP2NPGZKsVg7t
MSMkXk7LUDbks4qG3jk6b6fkbcMdUvqjFzZyIo9mLcJJ97qavEd0F/+mnXOHtd7Z
8b1jqwmdgLS1659ra0SYOfC/iEfEpp6O2Euds+V9EMJBYx+Tee1YMFDso34SCdzd
Phe3vzc0EJ0T9zW5fWwkE+9wxLS7/aBF+SqnL0Ee2o94XOtVkpNl+znDuuDaT0+V
laiwebz5c18qExhOWQ/aov5U0z+w88S/xOL6aTL4RIbDi9j8cp/vaAi+0D2rm8oP
F0z53SVeTgtFt2Ud4yI+/PLppSwE1Tl9b6FG1RwLMg9gi5rtheM88Km9S+XX6ZMD
/qGNv9BKNH2CDAlxAXHFfpDOXq25hDzrsvlFAesw1KMH+IVsqfmmzwem50Uy7EMD
XPCRBbwV8LWnqnfFygisYXpSUNeeyybfQqidw/zQwD9NFhFgCOk36alkkldOxp/Y
KhtzXC20S7DkCfq3nUaO+QCFgeIk1De6vFX9q8XjfqloFE/hu3SOatHK/uQw2mgn
UIjNsp0EKpaSKXQrt/cn4eDgNQWFny1yTZi17h5iEy5R7yJEzWUgy3Ym7Y9ddvv7
NKfFq3JYz3g1Td2EqAOcQjI5gIck0xGrMklt0uaWpbjmQOtAnbdnRe43btj//ffB
C0gLG5L0StPte06UQCjFQhukHNNnOrWTnAU+5vrFfs1V44pBC+f0O5V4Oy2MyaSY
Bn3Z4rF/2POP+y6otzl0mOVof+/eooho5T9iGCO8DDHq4o8jIsAyIzGU39DlDhey
vkmmbgvcMQOdm+yfOIX6r2OCqO0kOmUb6ose0KVwlJRKT57vg7JLwroiTf0lBK8Z
m73+5Sn/LxoF3dyPXvzoJzTUg/N0YrSdVXBwtnAwT4u+Bthuo08h8mOcI/lexWof
KiPcQ5YCBpnKa075V8AwWnpvlx6ctucRrEs9hdGPhKYn2m7U4gq8cEBwP+ibWu3l
ktz6F9AJSdzbkVLFsJXw8qtWBjjGqlcrwYEJvkw7Z4igevXl1MG45DF/4Ep+iNSV
uOhnIT4bNW2kD6rsYjRtSetzjWCuxGYOpTUfh6cbUjDAIifBjaxhNjt54KnZuAZj
b5UypoOjqSIpxYC/a/U4sxKyefnW2MRyGV9UfIh3WCDnM6eilO0VCcpws2f20VyL
dG/rgTTTiK/5oPXO4SbV54uWdDaL9xaSwWIpLpiDxlnYcfFnljTzLC3URbmQqMN7
qRqgaRWn01gMG/nBFkDziWCz9t5nVY5FDPiO39VUZsuF2TPLUzLo8a4H1qwjRalV
iE1toW/NnMFmH4rckuSRnZn16ZCmXy83mRE6lJKKtlyGh+04FDYOGPAggyavQpnG
Z+HMO56guo3dS5FfGFLvDaJ7uCdugIdvoGxZLIp65esoSF4q5gCmqqUUqVoJlx/W
AkWf5DJDTCBA8pOZV9YK8Gws1IJ510JhTZNOoQUHMspZkA9Y0PLAhA0vechsJUPV
ZF+9IpumRENohjafZsQukVQKKyzkA17pwdRPxfapc+hPDoRPNFSrpI8VxbgqSa57
4guvNMAp2Z+7iCJBqpGWkTyt0S7hUDLPF5Wlowv9mmWaH2wU/6nkpYJXlV//i6qB
otQ/YktvqOoIbHkLQG37VyFwctjNAlzn+SqcqMlH4UmlQvEL10/3odBF7gDXHgSq
KML4l5rz6xTdrjJyNtuXHj1RV3dM3TNhpEtroqSs/DDrqE940izzzB/Yj8GyHvqN
YO/WHBoEjIUNYD08NRFK+RowskNeL5oKBz95/DQ2arDlhohok7ykQW4DHTLmo2bd
kHGpC4WI1nkop+jQTGqWKhrKhLQnegdw8FRFrEuFnhfa9S6vKBb/zyAMQtDW8gJk
HuCBIGjGf2QKs75L8+bIby8MAc3AiLe0DVXaozhHE0x42zglNcX+iMBUXURBsIH6
96U5M4ZHGu5uiDzAkw+Shl2ZQRxBNXMq099NAqQ+0TCxqXIIQCyi41kiHxJN/m1e
EG8eJgIiydpoTpT6kkHJpJvBGufV2gkoZz96r2lLJ7O9hpYQcn8cPTRGnG+z7FI5
/y7q3fmPQUj+ytg7akubBi9qCFs1koRK4KI6s362Mp5gWnY0CUZi87EsuIHkzai7
mSe7juKFMZTr5Z+xlwXfJA2GXVxY1MAbO9yqarqhPmmpjFqLo/iojbTis7PKAvM5
s76X0+lLpYMorfqgTIoVUumctbh9K97ia2qV37v013IIwQ3cAqbJbFoKcGetGof2
COi2JivUoNpOS43l78l56+uH2XjFz2O+0+fAIjOTCmq4FZ/HXmIP5TWlLWk5je/1
8owBMYboLEUVSAzTrU+Pbp1RJsOi5II3ZygFPsITj4tW4SK1+ved43HDyuuENWrW
2uchzWlkwSxvtfJrA5zZePRRdW32pOToV+v1wj+t7jagcmEnIyqW3GOEaB6miP8W
sdf3i6LVPzU7v2z5dOHkqmM+7Wk5Wml8dutxw0hXSwYRq/rRxlPrhkTyUlJGjgtf
rUVtN/yVwvngkM6zD8+L9kSv57L3M2tjTlk3gBS1YJl4aLrfzPxr8GI7gXTy8DoE
E8z7BUxkm5s37HAiD3QT2wajAFCO/f1P/o9gZ5Obq4+Kpa0URHo7bQB93LAUP1Tu
VYIbp+rIO4I/MF5BB98yJN2rIfnemOf979OG0TutfMvaUumwL9Gdzm2eP84UQ6Zu
CQlgzGb57GlhncswIoLC5HmyUETL0diprL/PcIdqvgGBOfqyD2wGWkMlI/agZH2J
3fO3dBwlBz3R97hJ/Nrj7HnD00W9KugrC1fKD5EEbSNPt8SDw4CyT09yAk6/wqJo
VyaH/34fy4ngx58+PtsuPhs0cqGt1vQUaVQFX/WzH14C+FSP8yp/Pw0KuzOHp1pB
8BTWJ0J1AadMk9omeY5CUVCTN3YPXIYJ2erQB7qqhoeee0E/Yprz0ZUyTKSbksmT
CCxyNkJlX539FadXqjKkrp0R4fg0/9+97U2ImnYWV/JiySUK/+rLTf1idtUn3agt
QnD15QvSMEAZwzCw66EtlzYIWur4WlrKXpgY6u8tHMB5MMQ1d+QQ+OQFEarCL9tA
2LIA9jMzQb0skSF7Ihja4r8HQ9NwET4zS0m/rcVkKLPltKe6+HLxbFpyTt0tCjRn
QRY1u+RI2t4zdPKqA4BpqAcUFzJCQZJta+/ZiYKxmc7T9nBDB/degp2lS0dG0wdB
f9jII23Yd6/uVyv5yhRBQOhpj86d+tmgBfITrlFgjK7UPQ5k4zC+bvcq3+SSQlLh
kivbdTcczocOOHe+w+AdDYk/f+Csq0Q/o7s7inNX5MiCDPypmx8U4mKMyVt2Mi6C
tXT0lGrgbzXsqUtPvw+cLcgHIVh+3a9tc/K8xw6tM+FzCIZCAJf6fszegzFnJPWF
JVkTEYNJhpFFp3/+4A60K5++TDh5ywk/UyjHOA7nrxt6mh/aejA66uAq3upqkjub
28LK9gpvw+Mugx3GgzgFWtXTCINu4vpLiFDUi4cgvUZcwbZy6F2L0AD+JC9kB3HC
1YVNgiiMSUdKDQBg+v+0stKclKKIX8q+OqPBkq5de6f0UAjZzNpmgaVuwAc2O86B
WROWEBoZ3jlSvdGYtMLDZ3LodAgy60u0SEoUXrH5o6YLHhi7Ysx8kwooB0IIQGI2
60IR9ZKDZXRlgjldVEDAKsB7gt+ZO9nSS6PGGi/YLo0hyyxGxr8Mv6zZYU2tnNGt
xt2Z88LOXfOfz/n11D/sy+VefD8RxDsVOeU+D7duYF0xXxRZN4llVEJ34uK4W8fd
pXuUpmWmvtPTc3iZOQ3gIrsvTFpuYYuTTohOjXT5PPnXNN1nHuV2anVWyg3B1IGY
cZfbGK1NgVZ0QtirQD9Q5oPLSjIQjeG8HE2Jo6nWeYTV56dCF9/DPqzFovUGUaPg
fFISMfKjpNqzD+6D1JhZdFWu0pvpGgGSgD+pxCJaNANq+0Y8pcpciHof9gOYqB4I
lkyxi5KBrevUUt58Bkp06PqhnBWdEtM9xciCFsJo1d1w3bs8kZfvyFvEkwoJ0JqG
qTtiGy2nyAQOpNDRE04lYNnrsY4aCGvvSz0UzSbuX7NeXKuTiR4DyOclh7XM2pCV
Uyc4xsthVm+kqwHP+ESsIeyM9eHVcbCwPisHUKOmx4THgomD0gZfmjVwc/zyXQI8
929R8aIR0tU1DROTIol0u/vDnEpdBoNdROtlUETEIbIJS72Ivkwa3zvSgponbvy5
6BbhD1wEgXjfc32S6ijjtE/2xwAk/P7IvuEndqXFzUjURMq5HwiNRT+fREe2YNEF
EyldXK6yA8DC0bq0+C01qA8OmycMa7ByFCjJyw1jzHN+F1mRfT2BnAIHJ8j3OI/8
jUul4IwqAZUCYcpbQagsp5MAgTK035f7cL58XTtxCFi8rgHKo1F7RZiSbWhzLfYU
tWyVN7KF0zWQB5ncIHVBJYxHj9aeIkltJTlTImdUl4cGQny7AsY78q1M6E0LO/2N
M4RYDTUpXp9NJk+NGhQDn6JxSc2zFW+/mB153oWzQw1vMqy3RO2QQV4WcMvk1Ied
dpjihaLlabc84JL6G4eIqGo5eYD8t87hQhVL5hd2vlYZEbCGkN7UwWXftSXxhxE0
Lo1PdlVbDrVc7WZK2hyxoQPoLXs6z3Jwi0rFytE6zbn3vEbrN1cupCFQr7ABfq/n
thiPo0zfwIOGoCXsI1nfNnkp7RI15RPfd94KD+6yVuf595ULUrwefpxJmviqqlhe
h3w8gHg8B1Rc+fRj4p/NH0ezt1eN4yXlF8WYbqkWhGxPkgNMXZ2DaLRn2sZP84+H
k3kPJ1Fgy3rqTcuuBGM2DHF4vctHJE9QNBjpjpP0Q7zsduQriJDc0lyNvvRLPD3s
ZkZCJL39DJp0tAce27a8LZ6LNnIJ3rDGfuWJh00hu6CwXTcXusSu3aJNMsL1/mB6
aWi/f7lAEC48EQHzgMagzraVTYSHy9dqdZlnDFvtBNdJss6puDt44H3UbXKJBHow
dpuUxCt0anJ4QY7rK66Sth1gmrEcqZNQYpRH+n/AJJr/LdIcwtSKk+RBZ7L5FlhE
0vjz1IG+aA7ukRJQ+q1z2lQf7BpfjJhxFH9RNPB7k9pI8nSthXfW1G9maadJ222V
QrPh1ipNMY21yeLkm2wSkskcB+pd8MHQzonSE4RYgtn3eUz+ai0mXjJqaJeMMQyT
ifZKjxUNbAafC7QJlSeGD7M4N08UW8B6bK0hG32KAK9GcD24+UXWSK8n+4XAP8oP
FVCVhnXVNkKla4xNorbgfF1T1dZZk+ulUPITcwtOF79tI4kfsUOBYl8ydft9wNep
U22G+vyBAD1sB5CEHkhm0HtsQzjyyl4Kr+T0x4r7QpP7YH9O8uylCRqSyRqJhOMB
QSarlUsYmeGSV0oJjJ5H7gJoswguIgY6tHjY8uL3WCkt3VrfzmHAaFyhaPsOmfXJ
O0Z9+Lb136khdn257Co2pr3OBNhuvG6YokYEJxlYP/sFwyqJ2Vrl6mV5fOBfLnWc
wu3qPARVV5L8YZK9iMNUIKw20dUcRPDMZyiURwsdlEHkmTQBFdNc3RwsYrb/JO/b
dt6V6RMPpYKQW/eVcvLnRRESM2qLQugpSL9JkRfUFS71qR77tbAX6E9KtmlEKneD
4qSZE11pRpWQ0hs1N7c51brsh0ztCgAfu2MLYaqMDPqrvg93/pLg8+g1OAqDCQ3z
UzIkxLWJAr9ed0jQ+1u9iOvk9l8CnC2S+BGppgia+Q5vcLVVvS5avdp9FOIYHbcj
c8IsX4uFHG6TcsMZOrgpIiRkqzOfg00yRiEFwuNnce93wnFUahO7hPskgbaSTS+e
LrMfkVqP0zXE3Z6gB9f8TPjQn8rYmDRD+RQW8pcQCZBE6NaQ6JdtbaTufDY3wbsH
PlE1246ozWe/v6ucFrjkWW15Pm5lq/SIT0c7aKOcxjucmhXKGMF6qLl3ReqK6k0C
ORREMyGHtkld2b5moIlunezRyVnas4hOc97qweU8ZLFmKoFuRTZTmKLhCysS19Gv
9NiT/rkCoCJt443kopRilIXHJ5ViasUzCQBKnOtlFppxxAZboXP0XcCBSVCBbCZc
FyuYmpKfcvIIZq67m+IV0oNanrvnSkGHYUxuS7mSyGcd/s0l23zdqxZQaiv3wqdQ
/ifeLf7Ixd+Xt0Z9KxZye19dJnkMMAkOFXEILHtzx43j81cb18ItN252ZIA+IB3T
m4QqKHPRRdLh1DLGCcDlih0aPDikF4BtuTiNQcs4t7HVNczlrMq+ARnkRVnsD9du
SwLMnP8MXKNP3tzmzLoiEQBVEztgjgJlF3hS6j9lELGXiZ9c8pX49/x4ayBaHp8E
BNYX/fCKfWYfmTpQJ0GRTG48sDAxFazRNMCo08tmuKHq/fZz6p59DhQ1eTmMeeTz
j7wXi8sqoo4xeSQgQA7U45PQhMzC4pvR9ibPmEp3fOIZi1gy+V8ZJ1P74vCxR5kK
ItxDKwjEF3Ta/BIJRCMgZ4+ih1Zp+Gz+747bd09GdDr+jXOa0ShrDgQrAeBo/20n
QjlL7AynUbk9zb5ru8guBlAYzAlPu2jH9k4ZJBVBXa4FNVmEclmZlM3m6SjDlLom
tJ/QiVaP0/1KUBiWboWozVATxbj0aZ44sqOgE+jKByyuM3+XRYyCv9sMv+RgDmsq
IMQhhaIEr9zjAr00KrDRm5WPi6xc/rE8URvZsRVrVvVK0Xoi1xfGLlcUQKAI+V5C
wzxDzEjfszqfoLEIMuQDaCBqsaq/B2YNDvylgKYg/2Xia7+CPAcIA9b7H1ztmfRF
578nDujTQQA6ewLdeSE8NX59He2QaO8GFAGm8LmyrvfEBDFZOL16juHi0NrflA6A
y0HaJ8KEARqfzAvv7Gn+pd6gaeOWke2x9RCiVJUfKRhEBGhLdrjm1yedKvfh3CQJ
6yyFdHHKf/wTLQt8sZV1sH4SQw70TT1Rv0q8PX+8A2AmPAm/cKcVzu8MRNX/UHBz
Rx0ouGIcnHVhp3ywaxVgL73J3cdQS3sP8IKvKXziBH69+JE6eWPQWrITS+D551CV
2nrpqJiuCPSIVQbPWX+RGTb64PfNqhCrtJDNKkEvPi4ImR4M0/pZ1/RTG1MlDCYY
XJfLV3Ut5YzGkK2n8AtnsIbLyNn5X7cT7R07dixXTF4n+topwGZef+Y2g/3gFw37
7U1SiOd10hUXHwk3XfoZyPW66b3gS8JNOl4OkTTbYkUWwV/A1vVSlexICUQ1K+Kp
nq9PxuNRIHhbswX0883cx8yXKKVKPswCVjh4i2jiszLTlGma66A3sY/ATvf9jK7b
heNYwI0JScy65j3cUqXkRuADxAhe1P+j6WLrW9olIBgl1iZdFNoNoDhuOYE07ltR
HPeu6tsT67uq9LWfMN/yg2CD7VjmqgtQ5KMrXa3KlNAoJXYa6gXTi6bicx1Qbrey
j+VZL4UNTH8ZHpG0XLM1jX8RQlN+6UM1J5dVOLF0MYyb3qeQik1HEMBdt9TbznSj
5FK/zDtDQxMtQlaGmO36nOd6G8ZYUOLhDGG7wE8qFMCDD5OoPbkIVdSKpEwAFMZf
XVg8906K5xj7yjD3BCxgo3BKNx0zJmq759/Ur3T/ugTbDZU7gzSZhfsEEpinQD86
ssLlSt8GOoMhVpU3FeNFKzhRQoQTcR/6e3JwnokJoiluzZ3XvGhdtC5kd9qNjfHy
1qj3V+HEIz37F0SeSR40y037G901kxbM2WsjZ1HPoRqwIbp8hN4hxxn/SFesRnox
eMw6fwzvKs+UCNsoScjcuUi7Sp9UginGkL5odxgOGiUHeZ1I/8eMwR+Qu5ul8JOu
EvalFYeJQ5uwsH94XOK6bZlWmb1qcQvg6Bp38yofb7BDp9cJvjSovk+wM3WyR988
nPODdfG/yNpoJIztJ7pPUynGYtSkPWhX0KNfzypY4ftO2jyadij1Z8c241dsYtaN
Umt7jBIqTCzoNsqigAhBWCfSpBoX9EegW4tVLHqPU0BPcZ1DUCkNRL7/ziMQRe9D
dg4vABflJPjmz0bhCi31l/6/nxPdqnjo6zWFBcLmVu8NBwTVTvWvXNxAoXR29Q7Z
Pv+9W/cnW6gM2yDMjJCS7WcjuV+N3X0aGcbL/uUiQYJeisQ1nhsWI8/mREFtXQvk
lS4kmcZjDEQZHFVsrt7xVgZAlotyzdeREfB7fJAkpRGKqVmI5K8VoL5HkIMR+dVQ
ILSWZ+zj7qTMVlr488oVq48M1zUcVoL0keVEU85Hh9rEtKloLH7Mpiccb/NHJFXm
iXj4sa9+xLgCgVMuxnga5YSDoHLh3QfLVEVqRwlfsqnsf3zCo7sJ0lx1FSoQho3K
k3QL7H+j1KW9kKA/cI658dyvJtjJKbDlLmM2+Ui8ts5Q4hoJySdl5zh6uwVW/8YR
qi5Eqe9SeJWD84f8XXZFgvaU5u3Rybxa3mPYnID+auWiiWIAQBq4sOAj6ifOIOU3
2zJb3bQ7E4fuVx+G0w4h4ADUSSDpIxAeBolhusOad7nPJEb4xf9L05gvmiJS9oEE
/fk6Ehn2rfVrmRp6Iy9eFjSQTG5AsopPaW87+t2QZ6aYQMQDFXajxT13jPBgRUvW
GaZD3W7kO2/JxJH8e6T3TN7TOVhtmBynKROHjhn7ENvdteuBk3ACGptWs4euUs1l
0Q+mlyz2HAKh3gxXxy0Cz+pgftrbTgt479YPu99gh7iJ15voSzPxz3/LyMmwg/AY
CEx62zWmYIcCbFZd2Y8rSllFxtgLyc/yUc9LcXEKsEEpMqMZVGXQtZQ8KsGvB38u
tvdJKRryP4Rx3u0iE58dbWyr2N1MVBvJuIjOWI4HzZ6TC4es2OA4gRdof0r3CY1X
rcGEkGXIBMMgjm7qEQ9rkXGGX3iJoZKi3PEA0OwiUqsdkX7++LKNJvqYvfZ1sXop
C75ulPxRlP97ykeEe8W8+hDrNJds5rpLQgbOv/pD6NTxtJi1fg8lP2RbU2C3/MKI
U1bqkIrOUE1im32/npXHRVgQlhHkQsg5DvhAKwMoQDBiUcDsS4AGQMA33x031QRM
Es8m7x2rEtHjadOsjU5C2O/Mdbg+16D3kDgWSBe4A5MWJ4FYwKkdmQxZyMyDYJ0r
28FiiVL39pipiKFhQzkAY5fRaeZBzwESkLKEX4S4Nneq8qnlnXfYAslEi0nIzSmb
2riOtuAtAzta++I3Gr9KapeHPJrAxgy0UJnioFdXBrJTy4gj65edI5tsTgqrwyL1
ocxmeHPUkY2PZqpAXWSulsHfGXLYo9M+VKjJj7JYhmEfhbPsIgDE3Ui3hFAA7hWD
+ZsRJWL81l62TSACu93UD0wareaSBbxSY/P9IUlk1y9UOpyBOW9GO1PRUTIq8klP
737r9rEi8kWlNn82NQd5Bp/TwFwLr8HwPSNO7VFxEyAZdxejZ86D+yG/sxIu7HK3
5fgH7Dx2c9rSLB8NauG1Wg8wIDZMVSAV2KRAu7b892dLoem23L4pS9vxd1EZlQd3
86lGnQyLXI3U/d53jKdfDBJ2JF6pw7vWmqp9evEVB2mis8Gz9+6PIHytHN+vQuQz
lf4/gZ2iCrhEJSwkpUxD7YaR7OpfKma2Dd6zviAMu/dZV3MoyC44nrRFMF50Z5Ea
ufClynWdkKKIryHg0mPdfs6YkBG9hhx1YaTY/9SWXcRs46RGPq3U4gFsnzE6g1Fz
2Km3zM54AZ1EUo5yBWmPVlRIa4YFPdfuz+zUFh/zWgipHzT+SizTUR/O4k4c0N30
d6DD8VRhiU0YSk5qtuX6XKeEn/HTVF+UHwD3a/o+FI3bYvyZOEtnYSB6Mlj0g/iB
EpgmzmLbxo8ueaB8rMK1NsC9Slmh7thnQ5mSXMeSWkcAXWVIujUfn26P4uSRktWP
bdcEuHLrosrd27Sicj4J1QI/RiInHbEagv4IwbtVg85+rJNyAy/MSrTSDQN2uF4B
t0H2koAKhXqeru94OA+9ZXTkecLn7DriM1qMCuEKmjDMldUk3ScOxM9lpp5ILXE4
pG/4UldaX7igVEVdic6cFS4/uAzIR3u0+P5/1TRxeHQ4qZpsGEKLVj6hpyhXOsur
6FjGGzONGRuG/D50LPcPykZNmr3FB9l3EKwKsoUNFDNCcMD4bbh00XxjOpT0N8D+
xBpXsZIzzScYMM1YoRQefAgS+qZQwJvn/aFAwix2Pt0BlAJKof5HRosqzdMVR8ga
oYDbwNak8S0SoSpIq7ftFevOFK3mhhuLpZIyH+NC2op82Pht+orwlIsSmq303sll
c4a0ltvCb+uIl5m3MYeV72Adv2zp+L7LQBWC2dlzMm8BjmpVNCSXLPLmeFluLcnH
WYgRdiUdNGCivBSw+J03ab8TnbL0grcv9O9plLmIgwtM2hVJCceIZs390O3uSshK
fZ9BQb/P6KASu4SA73kh/D93jepAMLL2A4yfQg3QviOyHZGSaBA93QOELraw+Hpw
VBHfN19VfpgWZTjgGiypYcXAosmofK5GViHklNrg93GLPFTSn+7F207NubDCWp9A
RDrXh+zWjPLKgz7NRz2axLUCNmhW1rQZn6qrq73MXRZndBpGrzreu3fNrHGvmfJs
NmI/JU4mdodYlvycUpQrAFz+qH8RkELLjntmTX1MYpc8edRKG3qz56gtLopZeno6
Hu7b5tfH50t+uY2PvO0UT7wL59W5vSLW5lUt3GU5TvugyiFTTdM16kDiN2OWcb8E
wSYASEt3xFj11Kv6Nd7xIoRcMHoeFZ7k4aE6YlZpD3GSXTBuEZahULAeyOftYWGJ
zngkZC9ZDHCXTLIXBFRAYwAWtWCl5n5Ty71/mRZPfuuWAmS4UUWzoPhiDkKzm8nJ
zwtq7lceop+YZm25KQE5hShc6nURLfoJGAiWRJIdCrPH/5EbSUabI6aK6Ql9KjE3
NMLmM85EIvvYBwCFDGQ6mACC+RjyOFKokBadX4yPjvpF8c7XBiFn5l50IHdGGnQH
oiiEvQpLYSuzLM3cRZ8rRfPJi/uQo7onv/ixR6e7mtad0g0ukQUTow3WKlVpvncc
KRG89u888k1PRUilYOKO2VPe71UZSm4CPxPsdtMnwzKP6viqTUhDwt8QvfiZ/YPq
xsQwSQbCKmis56dgL5R5kkd3th6bNhEZcZ0amCH2UedhenPN2ZZk6kus5U8Qzx91
86bTWB9/9zGyrXt6vQ9kcaOe1jOZqJfMAxdvMNkibISaXljmK1YNcSElB0j7mmgW
CgmJvdtTRUlzxJ9rVvg0UkDbVTgfMYBHa3sKgaiW7TpUgsuCwHRxd1UfBnDB2TgR
Q8OB4bYrZHaRX1POrOkElycnKZ+n15MIHji/5SQ4+CFxjpYcJgzIx/3gW7t+wKA9
R6A3FlKK58lOJo1Qf8ssCJQaO/amjBx8Dxe4pCww7bKCiP65fghxKPnIYrqOspHP
9u2AT0zBSWRqCCdfdCVMpi+Qt7zXwQr9MRaNSG/azbgU84XvXIhl6zxtJVpYth8p
28DP4gwrPlHkRKEDnRyOQGoPUW9EOKsskrTo96zxw8Sk3DNmYz6mhg5v87pCz0SS
mhgXMtREOjsN2dnBbuptgvoHxuSI0BJ2vQeutahPJW9EWLOFnGNbosjGpjlADzUk
VgHUmHSYGXmbqD7FZqmaAbtWaoABvS7eoPkqhTGgCSH4m2GeJWNNEILpUd8blKsp
ZxS/yxaXuljl+XQr9JgE69H6gsZQjB7XMdfCojf+3fd2YFhRynU0P+JU7HJ5OGGb
rNrZvcGd0AuHyE15MaMmP3dACivyB+UAjUFXCUXh/pXPHIirsnZN9ZcG9CWVgh/I
MIXgXXmMpe5qAjl3BNcBZv5rPN3YIh2g2UEBrv8k5T//p2baPB/HynSBjsJ55K5k
rDeSdCAgdn0+XUO5c6ddMAm3us48lYw1URorFqbhA6X3hZu+yQsCsuBXSesyQ3ft
hHknQufaNqhEleyce6nO5UAcKMZFVwukanf3ttazsr7J9hLOBAFH4KIYb0LGUexk
4BpWbveWHbtdlFNc4hq52pG61BbbOO5fYD4O7atwdlclmnmn66SqLG6ihRZXr6CG
fR3SpsJqP5GhXKcWA7DlPt6xjhvvq3E7GP0lF9Y6PW4++U3fR9vmaPphfUpv7xXt
GKDOGmoCFKLnL2hK8yp6hlHvMh7cGbF3Su4hGBUX0Gv/WzJ/fxU+ZTvme16/H2Cj
GhogaK3pEYSDTC1zqtHNvn6RYap8EaNyEW7xLln1QCfkNjWXmwm+fJLPunRQuLtJ
ZZFw+0jBaN9GqO6ewrr1YNzfNjt48mNnJgBt5MSGHb1mtZw8BO8RgEPhQ154+D5X
gmS4pb59ufDrtRjOrOBHtZwZtHyY1052LLjG82xjmno3PhaQVAy/z5qmOgIP7JBi
LXZANk56SI+UH7MnJlGmMGJyUHGV9N9gVdPRBOyideN4NW+NZJThhZ3cRLi4IcVO
Oe72bvQEMYibLu1Uc8ZLgCUITg58tOy0W20C7rlcC3p28+Jj41w7dJNbi3BaeSoy
uXKicE0VM/b7tyf5RjRmsU0LxKOzZfBhyrVCfN7N7QKonioaF+GIzdb8dUcpynaL
I92ApW7tEYgvnjj51Mnxu91BXSUmq3MRkPjFRDx26ukItPFnoSlGBY3l8o1pbu8g
t0y4+z2CNAR+8eGkHBrRJXSQioGf72ro2MWvw8Z/NbutbGPRA0aSLKG9yiTxIubw
ACTy/GiJCHxX+Mvv7tnw39w9Mn2NlON6Jw//hH996cSlirp6/Y+cUmdcwezATAvF
6wk9OVNr3SGGJGDGZnYYWMgVmDyKJRJVyGJbLuOfXYCuwgcMoOkb3JB8JBNF3t/I
oe0nlzHw861qSafDv/1csiSG/0WXek3/hdfA80Gc1zhs1P5wIxQCLoJCK2RD4x69
/WH5DmazCIR8qfv8EOuKwIXJaD2oWgRquBghIeXLzdXnuGifAwNR3An/jB8f5HFb
4prZmDouOVW3rS2fljArxQWXJHzIHmzhBWxDweQ6ozLgQdGI5UdYkbblmxAHzo3A
rgE0d3CtVLIy0imZjtPJEp6wgqLycZdUJ+6GzhaizIFXez4926siXLKi75JxRKTU
OxPNiaedxMOcIHnIxWzzvsstSWdZgY9B/bUuMcEXHr8HVFUkDeSqsb3hI85yAH/3
LRiQ4FVgSGtDCK11zFcft3ClKX4IRXBGwCgZWv44gC+iXIfoEOyMaKlpzYLS9hl4
w+mIvs10e0poXtswEirSDqMnSDh8jR9nwLspNgFMxCredz0tm4KjKdoMjUH+V7p4
MdZ6n1w/wENpT6pQIbzRNsWPNTBjt2BI1i1KMMieHzKSnG6eqOdCPSG74WYWg6rp
srf+ksozW7mTSOeOmxI+DM/S8WbXNV4fYgmRoRC/ecpRyVXtZglsV0RKaoSsvXT8
0d8vTmtlOt8GKq9HRZ8nfw6B0i1u9zMehAwXrr1gxalfiD8K55xQIYTho7etqHnq
bo2KsnN72Uoj34s5gE4Yu4/xSPpSnNygQw/bSHIfJj5omAB4lP5EviVTfi3Rbpam
APxnzUpkYCIl1oGlZ989mrTftQ0FPIif5J/4O06kV0xD2kKU8qxGnhob8nBFU4RQ
DX6csQ8ILn3P7PRRdG8Ah4ZtO5FM+IDJzG6reSZfJDCwPjdpYZluzotzjvvt5NWM
G9CyIJgONs6n5A2huZD/MghFb2xEfEITuWCAmy8JxW0EpEBZq+/ovyJu0Q+k813y
eJdSE7IlaQQqvGCzBD6+X5e7vV5fAPEbLLQ1mBpjcDrbHcuejoDO6VL5TT5Olg9Q
exjMRKlsHsHSz1YPnYzBPlE0JFdhFHbovorxAgn/YJ0+eSjoh4izBbtd+gdWvwAa
hkKA8JaTNFqr/QvuPdWRoxhEtItTa+0K3LTk+EutZquFg1GAZLdUgClRimvLqvOQ
+/o8iGVXASU+BI9uc6jl/SluqY1RxIi4Iv/GM2O0EkwtPGg0vugPRda9irWBxAui
QDZLbbPYhhO9m2THOCSX4Y3ae7APLrWI2uATa7tTc1fW+Ja19+IWk1ngpw+DBjlU
P/NZq1wuL75n+VoDTlMG7+8YRplTpFpRq7Oboh51r0LzgnhxDeuWrKQums29a4jW
lYbrORnptounG2DFhnKkvmpqYhbLb1IdWVDzNeIux3L33q1YrV8/6izVkswpl4a9
Y3c09F2x/ZOQp4dwyw1UXPn3zsEpq2E23BCc5s9Jmsk90jqKzwUAjOwrMI1ukySL
cA48RVvdSkAe0YC20OiNVfMAImsctV6d8vD3HlOm5L0QJ9zHf8a63+i2Q5SNaYUJ
PnK3Ousj2DIFxui+ubOCdnJ3kq2d4ZsPoSnYKWQKRk0758NfBIIJS0YkbaUqR2Ld
/Ntlj96tii8A6SioC829RV8nz93sz7uRw+G0syLBr6Ic5VlXo2e63TeE/X66WayH
dPjc9A/d5FgTmCuYuf9zrXEuL4lE6gKLgUJRgFf35YN2L9Lq5Sw1UK8OtDeO67/P
ltA4QCl+H7hnNEpF2EghXc5LT6k+DsXSd0kfBu+DV4ohqK4x13WVjrCLETzdsb18
g8wn7B6g1ekcA/J7hZiUpbPJE2ZqeQ6noctDY3WQNcbBE0PCHqbNYQ5eQp+gukLm
Xsz9uAaGS5Q7AV6MixhOVT7WK2Pq3LKLvaZrgGnKhqRi8UxsBzebpNiijrBoqCYc
7Q7jRXgVkGc7UWmdahh3v6I2peV+T/muyNz81bprQjZkHaKGSuF1Dsnwo+k12IBF
mKkk4u3WHelB9R0AxuykZI/EgE+qU9XiED8uBb94JIB6yqwFvgLVvk0a/K28EPt+
s6dYalnjsf2V4VvcKcJcKIG8ZJgb80aPYVE8WUFaUvL2JcNirOZUZOB4Vtveickm
JPkzi1gLvkynyXGwYWx0RPhwop3WSuiWbQloN+Wla5gLkNyg+81+vCf8xf8w3x2/
5HEaDu+SXfB7NfjWVNArV//5e8B6JSkiSbU4DtP/a3ofsZNA+sY3IxE397yadIOc
6B2J/3F207q01IuRVrNibdHTM0qX3U8JMlxhOyo6cUbe0lqxrjuPK+Xfz+tIwRdL
eFCD//VrBt2v0rbxXlWhvqguSgknxE2uLVOjJGr65ldAOCvsA0rdXMXK56nHJsjh
qEvtzzNSvtHTiCfY7OSFvWkCaAZvRhFhJKLVWCPqD+8oAu1QjNV9fDMCDAUpvXYU
98SvHsKqbM9PgxjcstiyCtyFE3EDupYHHgQG8pMf6tLrfh+G3T/B+fs+IA6AAOGD
SjxbW1d6eVaDnyBM2X98l+pn26QVBCRQvAyLJI3F+AvH4WX9xMoFcLuVatbVB2po
+alIW3DGFQQpBFjlhWjZIWX7eHF3HJBFXAN8Qof9SSgPyyxBBjc2Kic4OEEpHJNj
ihWC0l59MOTWH/fh1SDc77Ra6oawXJdaKeuO/PKda7MLo9SurOSYqHpI+34mhfGk
N91S32k7plW6cfAVsh8xc31pePxG9MAbXc6OREOhUv4lqJaKaNMtho/uN+jWDD0M
ahBXizUJoM3ywQOMzU3Ns5bZdceM2MUv68eg5xsUadyIbCH7Up5MK7mblE11iGfX
sZV281f6v9nzRIS+S/2Oj2fRC6L3oFojbzG/rgp5JuYsczd/pgw38nq9HCzYm6vX
Stc/iPvYmOIosRCgRpQaZBADMu1bqTUH8a0/f8QFohOYXAdVow+ciX02nPm5xF8e
Y9zKgjpOdMvVauGCkQmNeaam7ytB6VG+YF56D09y//WeXPldzE5aZm9Wwihxn+Fw
uoKSfWhQNTLxhAnaeuNreTz6QWL0keKNe9IRkUgMZvpxW5RnQteInHrtJdA3kVWI
O8ozPMK6qlsBag83FKKotpUUb+0QDcSdUoQp8OdcZbWizVuk/+KTJhq2JbWOccmb
v797UN601Hofu5U2wZkJl/AxggcMS5YTqYwj3Fq8V1kk/sl6crADeVxKsYSl26+T
HGlfNeDKvrsePziN6SIBlaiIglvp1X5BCdIGe74nJps+zWiw1TeHe+N9kfji8M+L
imzIBIE9dfW4VTtUy4UxI5KH9iqWIzrt4nShcGysBSwXnQATqmeA7IQpaO/gjqA3
Md48PF2M5ISw+xmDZZ6PMnNaAMeAjgGg42OBLJEY+3xadtD4OHreOROCX8gORigj
fnLm5O253yKX1JKvR+xNxEmPPHNsd8CgCVuUbS8m+HS47dLWeaOILgrpBvmJoFvw
DwMhNh47v8euC4GNhNpjtZyO0p8ZGPnFcngQBDyCXfMpY5xjTSHmnN6GANTTF/NR
jnBGq4qtFqNBVKdMD+ARMX56F4udx/H/VqW1bom2OZYcfM2ni9t7k0gIOxdGZ1fo
c2pFI4I33p/7UqXGH6nERk3M3lXVNiSwm9rWO3vHlELDREHDBOexp3AgpKeRrHm+
qxlOTqQ1Lxzg5A4ZI2ui0AOhBsegQk6FE/MaPrAt69Ntl/k9INcjHT3dOwZo9D2v
ase6HbIszvbFSSHuWbQQh4JQJumyth0ZlyQtsITbhvrO2sZm9m94zKtk1N7X0kwg
YXhzpjsOXVvWhtyHqRGWto+Gx6CvJZ2Lm1D+zIW53x5BbcSc/GM3vrf3k4KwaUuE
LjMazmJe5aiqnYsrYRqnk0s/2RWj45/ASvLarlijnPVjKE/lrv4CcdnN3IyRySyz
0//h8le1OlAXhNKO7PNhWNAEC2XydYj4QFC5H8C+Qt4XQr/F1gowtQSuka8gG225
K5feaIdT2Q4/0xlPkYFeDhJoYKoybtPrt92OWTvjEtTbze7v/RUPxtq9vsduqsW+
lBX62NCGALM9LfONrewkYJMqjUwhvr3TUVuMY5uDIL4U7ErLZ+Qrg/y6dL5UwCfU
8WcDH7lDZ/uG0TKfh3YhuttHn7TDkN5hVRZ9Z7MnXIyQTOxqevTiwB+hmSyaLTKj
72vK3q2L+NzB8VRSSlEZMfblejT3+brlYVtPbxYUN7gTnmXjjoDZ+nB/MYKqmkax
9gbemjc9jFk8GaLXSCuzm8KmXo0ICEmVV2ERiaX7s+2iCnXD2he1l25wRKNPWvSQ
4pHGJQdeaXWOv1dPNTQlsM5Z6aSeOXthgGV2KICb8adqo7pqhmX9rKtbEzWoxEe9
LCOBeP2MC1DNv4vp6o7tZ4n8Nt3T3+g5xJaQbv+wCfXm3aVjSuzu+O96wdbSkKS0
9kPkOukXa0VZvW7S5rYN+4OvdCJmv6zwdcrQg6kpSzxESEGywnczlg3KPz4V31dW
YUzqa16b4IIV3Ln3z2B7d/+xvde+XeXvJaZTXoAyFTgam4ur1hIg6npPSQMHeM6y
nabNclg9UdSgxFi5m3NqZKjkBEnhZTmOKmQF8dwCFOlOZKtoyAKoTKi6QDsf0lrT
+1N7+2O8wkBIfoAwsVlyihEBNWCv3gkorOqtgfXeEE6H6AhPO3IpYH4NyJV/C3HO
NSTV3UsN7+i6EWehSnJ7dk4af5cPAqtVftJywBiY7boXjW56UzWXzRB1Mz4m8qg4
dikalnOlCN+wBvUk06lG1t7y2FuZaE5XI1ltaiNzqxwqjT0xEvS1B57U/4G6Z32d
2v2WHayHkPkNj/yPcBUZSGqFxmUghpH6KW3AWkfXRYnV8ccGXzlAqT5kTnoSBFkc
oTmucZroegRn3wSa9bU9/Z97CaqulX1kzUD8qu3GZyTqEiYAqnC9S7dUZBm23jrI
Es0B6bPHLsS4JpFKjp4Ee2cLZWE5WczL44kwzJJyaANFnFXQ7V1A6+JU16mNFkx6
7/gvfwL2MUWQO+JZTlormnoDRritLYEsR2NjdAfehoB4B7uq9btijHKdRjnR1cWY
klwQV5ZgxBfVwCKTqa2KTSMn5hnclDyBQka7kkUiCqm8NbtM1tFTCggYdgJYfaR0
9MIlCbs2gcWsdpYthDTrhY6cbG06KKKEprDQgD8ihXk/96hUba40yGVlF4Oi4pkC
j5EKUqXuta+MsRbyg3+a/2dbPLwesgwHsj6n1SWwgXiJ7o8BUphDL5B8YDmLZsCL
oKdlghA0PNJ8/hCmhAxIF7WZR3U5mvCQZ2HIYifJ9uoYy8fgkF2wXADSLIGTOodI
QXgm7q8NDSJ0hVPm357M1Z0tQsywiPrSnuTrjf5hoIOQKVTyseFV2FiWCk2qJeFj
l5z/tzX1Ki5Z1/G9XLl8BdkJMZ1AJSAkljFdslhVIMFMwmmqffIXNQpncr3P41cw
2dnjLZMfv2IajNabqXgF+EUfI0nJrnpNdIx9w0BURxZXu0jQCJEMzeJ8kfiFmZof
KbmLqXQ33hX/5SEsQOrSAG9XdnP1KepLH5lnJJzrWl7+oRF1VRzmAMsuDjhgMkRE
pClPM3pqoHhTcJb1dVsShkFLr8zHzi028TcDnLlZ4T16tdYE/TZL6T2RYA1wa0Ha
aHENj/J/eEXAepXPuQJAHDT2EAEpkZTOpe+vKmG9GooD19FK3nEbXEoWOxOkej3W
eJLC9s2MHJQeBT4mTkSrJzGxHF/Llm0ODCKpG5AM8ycp6BYHTKXPxWoSkn8McmGl
yNmIF/ZpoMKKYkxl+5hYndZbRmhhFKbsUziUv6ieItcvXJEt5yQEyELZdNsFkVGO
FllfNo8eHPzrMjFhG7f81qSzxkjGqeXSePmk8XebvAlkMoYrWUf1BTMP0tp/Vp0i
ZupP1q6CfRU5bVnFEvt6dZfcHv+qOqCej7SYtoYWYO02TBmG3Lf8qiVF+u8elxVo
+/cpQYtpi7pQNQUJgCxhziw7HCtrCWpsSxcl6VtqL/6AV9j0YiHGv7Xcb865QZNO
jm7D1YBT6iPP16SPvx8jgMLQLq8s/DaH8IlEqQxh0DXijXQCKuNGlXIq0GH12Ofy
7flePTVTHk+C7EPSe0qjWO1/0v1K7SFs/TExQwYH4SW2m7MDnHMge4g1KnYvtNB5
fQN+M0fw0iTsbLYE31t+gwidaBDu3PbPZDxLuV1IzgGc3pucBMLbUVtYfUaYuA51
iNi8/CY1lSh6fhTCSa28vP+v3aA4uup02uSmQrjyHGzM837Rxenwv3WhbKGLYnty
VuiRIjeqZXIRR9KtAzMsKx6hVPylEHduLMIwBnq59ekNKDOW9c942TAkLsZAYAVA
atR6j6tPlxPIn9ZCXZnfooqKMof+BOTsLGgjZyxwIsUUHInjxT8pPafgtmCrcytS
4C4GJmO2Q/6dKW3eOwVtYd6RZUimcSEDpvSx1uKlwBpTJR2XrJgUfdTfF9hQC4fL
7YM3vgt6dfAaFwNyPK23B5GW0hiTh0e7ee2QzCAY+ypvfmcO6Y9+9SNPx+Kkajms
P+YlDLXwMHnxWBiEuQTfD2Q/1ywbjEmbnzIC5kA8xeWKZowLS4EWPYyUuMTQADCi
CpE/mKgOXt89cQXjdGzfep/Ehow9iA12rK6d/uuP+l5JkVV64oQp3s6Zp1L19Q/o
sW/8RurOXUJOO+5WKVe0+PaXu3ReJL3tepuQHxWY9J1N9xbiMi/fdP35wIMSG6WY
qz/xN8LOOo4IzsBjQgpAtmX9k3h6UdYy+THx3mXeJtZ+0ZqcxNQvDCKPTeLK0d6t
wvmO8dmmJBcIZNgxbs8pqgQmgzU8+oKfQDkjGJjdAeWoIcbPubD/RxjybxKbSvbv
8MmkQS/BddByx4giT4fTDh9M+FqbeJei4cuJIK2C75rHW4X3k4ta/2uQqwYSNk6y
6KX/mIpDJ5uLxcHG3tsYLKNv0pcaFwwxtQKbKEj0XRkqSwmXQmyOYtlKgFWUF88g
eMnvtW4eqnunOrXienBhA+2VYZAc3fL4ulQxxty9VqyClDSIcXyojjvgsX5mpqzH
VN8Xu/z0VKcg1tLyH6n0sBf4YBfOw+T3rPWP7ccjJDgUeHz1QateptckLxKXeX6k
lmST0wR16tMuor/UWVTjerz5LWV+TMTHvKrrOhwfNrUibWxBtMmQpSRs8M6HkXJb
g5kTZ6ePG8FKNq6/iPlJOaeKqODTlns0BVRHMhmCFF2SC3uv9cZ3018uEXZEp9nD
0Pl4snZ5krpPggQ03hnxzHwmbuC6vOssEL2T+dhDjKxcDf/XO1rOM1CnAIyRp4WJ
2YTyVG/X93GPloil+EHvvHqHWsaKBKEcRZY902HhB0MtPr3VQB/Ih+UzQZPSdqBY
QglN7/WzF9BqIR2tiziqoDvgmr+XV8LMlYmplpD6s4RYgcLpHiot85N35bhulRv6
sUdE8mYqAAOHEYB+EVyMe/WnF2MoxOPfyYWgLxNhX2tsBJnKua1limnNH53T0xBB
5/SWHnxhFGDsjoSxiB76SpLtLRjFJXiUwm3IEpXTAnWRhnT9uJOFXA+Ihenao2Qe
iY7Qy+0lng/dRJGkr08Lta59ckwPb1YcWgnJyjBeaAxI/q65UExytnaHdJL/ieTD
bS+3jbycqEb6w+jEdR3mWb4BoFRkxfqbAMDwg+pIcdF65hzph6rRh7WafGcTP/3x
NlmansHzeMfUbWxaMkxetw66C8lODkh36jVd9cMuyeVUg5I8H7sWm2iICh7kePMk
b/0eZrVgkEIUR24hy2XwBBI8uG2jH4341+663OvKmglB6VyG/mLU9qQO9WmzJCFw
UqrtcDrKAUGr/5k3oU7IuS37eG3uLhVvNfkGq9q4yaZxZtzmWWjyuqkTGJKyUE84
dRyqm3VKttcLFoAECcgMEZQmEZWOoyEgZmt0L0UioiDs4fnIumsEpxLajx818Y8j
zZGsF2BLfPHnQ8LzUUTUV1JN9MUkqkaHRD6zejsZJvxHJ5yaC2g1w8ODB/bJLYzQ
buKx489TumwpyRf2Sg2xdbRWFyjtBuNCHUQqZH0o224+PIBWF2qfNZndNHlPjtnP
GWM5DGpiQjtQm92BLVlr4tl1FLT2lR2R2trbd/i4EQTqyyL0Kftf3qXOd8zkMbUh
XD865g1oSHThr4EY+r1A/7muHiDvKiI5Ae6YCRBY3KDMHEWb+9x/1CK60Jw39tgc
yJB0d34rpOG2hspVuGZvszTsJpMNTmEt0rfOzHMZZkWUY6uDegF0Mu5rxmINqDfr
Hv1OLC3BnXxBXaMGZ+MLRPEkiYuk3PLZ7xTi2Vckhl3kTNv6tQpboIdzmMMee8hE
b0hLXEiaatHfSZXpwfZ18mf2zRV64eUNa9ybyOdkYRff6v2gU3oQHHevzJ/Zcxwh
R9VomhSHiy5UgFaUnwcWkAXHmAkZ2D4kZXzMwJb7p/d03QLzLkWKAknJ8yHtPmn5
5fhWADOphApTSlz6hPVwg/Le8VNKB7G4F8aF1vutfGuTsLH5Ethmlexsig00QWyS
AUowvHfDGvn9CkkoiDTGfKRySkKNSvu/YcMtDHYpPv2dzp3GcwCrxw2kCpxXkEoF
MhyQdN0NxzAVhOzysQB3JCvY7jvcJeyC/QyGMlfuEq5aZqYYx7h1Js/it/xcHK+4
vnmZdREnmOSD4AdKmLDc1VKL83HrvkZqDszv87RKw4FNidfTXTwCbKbWXGTQlPx9
Ha+pgKj/rCgiQluzVIWd2QG4FzWUWcCjdIUpMAzs4yAes55bhtMdi5MaF2crylUu
6JtUb0w+R9Pl/fTgWumTm6bVkiyUkjLwPAoWOwRmjTm/7yH+2LLpzgDHKImi4oIm
yhf78zvThPPRTuvEIIIHurQKXUppiHnKpuWVDwGwGDHQddztXQwA2LY0HZt2OBRo
rR88MUVQtHjcPo5MmuaDIneqbR4hE6NdWodCHgOfrjfDUWgpzmeggNOYwEoJFAWt
wGUXRtK4KY/vQQB+WL2yY2N2kDK/qVzFwYDMjgriZk6C3QRdbdbvvdwkuC/wTKh7
7X5PJttlJ+FNUDFsvuKxC0Q+49DBa5c9RnVFx7FO7H4XKy6cuMaAVoTPeTkuLmlu
NKaPTwDbCtQ0m23O7wthIgspuoG4oiFuMSBK8wgMWdebU0Lr/iM5vzkbfUZeJ6yA
oGJuGJxxBwjrnowJrjYEHF95euiWuxJun/riiVvZ1OmnH4Wc4iz6w4ezKRwCayuK
mLWiDeCOcnr6MQLqyZhqxpfMUaGvuCMk9JZPUdYmhmQQLUt6IckeaZpWNs704Krc
KgcFCDdNIX+1UYBHKXxTiKrYOy2lD8AtQw4n3eJ54evn7qW5vi4N4U5uwudWenne
LbUScldFPalSxHAwbCZxrw2GnxAKvy6sdt+Uy/gm6kcYEz11a6tdqvzD1ov+Vufr
RbafmohkgXvRK1jiSYtLiY0HzXxmHLYSnToUgYsQZXrSFEqSbf/uWBJ6fXtHwyEt
Lep/ylyaNHFBYCV1Hso5cQ0NhUhiYVWgjdOxNEk4HDIg2SujbCHl+Jf8/dGIdF9d
mDUJFODP6AMJftE5DVfxj8djPyU0a6nKLxXALEr9gzudsnm5oAOOlzHX9v3Yrz7x
pTWHHWZGhdSwgEp+d/m8Z1mjnQaJ02US2mmj6DPu7UG0rIV60WAk2BVzLpJYSe92
ytLpaMw1ePMe8LvEzB+rUCFp1A/h3n4GVavYJ8q0XVx80Wy5wRhyWIbp3x5+GWNL
SQIsGyY5EijyjXyJLEwMU+Zcku86hPyn6noEIInrNoVjcIi6KMdtG+P8mJLmniC6
w6oC27vRTt5H1Av8i+PAaA46D1OHKU/BwBUP6WKql9KNKGfDz8GSUp0LqxrLByea
DPaKdzlmV0qspt1+02Mr+kGlPuHKv7v3I6WsKtKqJktHtly3YE+uL2c1g65S6UP7
8RGqDIjyE92bZU4zWfwDyR+3ByppTqg9g94fBKlfxij+37wvn3wAY1JkTkJ0Y9pZ
WM93ywaaAd4VRjWNdF0z0JxHlKXsetAm/0Jp/ezFsEDolNV/0TWQmdB6ObOVKFh3
Z59P2QDXxn0mctMQHNHsPwA/5h16mXRyee2vucx0mlvZoN0st6r0EY1zcO2atyPK
UYBaeiRA8qi5c9htT3vx7hPWwCN1cIiOm+oRFxjjxsxAzSFw0ODXaG7ffUIKF4ES
J4sxwot1F9xqwBVaEjbBJKACq/G3ySm1qjwXdyDtoHVZBB1wF7a1UKxVjgvm41ml
15pKKM4wmrbTVPMrBj6NEUkMphwCluDrIkQPcc7/bDBSHsPX9aFaUIH35byqRC/q
ndh/dY3DG93dfhkUKQuyA9VhjgTgyBZ/YdR0Ctu7kKi0uX+zzJx0ZLPk9RcbXuhg
sFjBgCYhTeb6/qXESzKGLn1KLX8hRbyNBm8zYc5KBW///hBddxGk28iUeHfRp9lu
ddI78ZDPb97VgfVl1Im4apd56dYBMUq3ueJa6lvc9if48T+QRm2xsa3AFefGpt65
BTVtrRJKXE3cB1JiTYySDgJmO1nXPAh0GS19brLg15EC2KALK3CXVJWHXNo8avwx
V7GiE/g/HT40LgNNTsAj7W5YC6GEoFPmLRHDyj4nLL4PBuR+fp4t60cVZPKaw/GO
oq48L4ueD9Mm1BL7EHAfMCZip9PJdg5P37rDH6CimA/lLIdT0Qjl0nV3lb86YGIU
XaItjrERsGgrSDA3L154CDaLVGnBwoElQrWYVRATAPRTsE//UNgWbAJ0z6TfRJhr
MbKdwIzdTOliLyG2ODQ3lyhFYq8wFJtsl6eGhHlIdpXoz3Zx8d+GA2pYu5zpwkm8
7Yuudd8ucOBGmYAHGwuEZlyCf+5h23zjTrBYjUKQq/XG4BlKQiuUaE+fJnoKShcY
XaKoKCVfdXq9Y2wKSfRn0LJlYHAd8gx4rCOPYggjfysBogKI9c4JMbMWXypURdRs
2Vob/DQQDdFXjmBezTugoPLK/4/4OijgQuaycyp2X/NtfVhVPG1Ya1A3v/As0xpp
Jnm99fDCEmeJ8Np7HOnm+Uq1U7WL3egcylSL398K60hBi2HYuYEHIURESuHWvaGX
tWvf8dKb+AuZet+rM/jUNzB60F7Q4LgVAZlnwM20TWYRMszghGPuzGAcndjsv6GH
icdSLiJHf4Ikwv5jczTBebOpjT6lop1CKlBuBySdxIUJtcVMiPTgEHYSvtO+ttyB
taEBGoS198QYGMgNvRx8kY3MaMXqzzqq2FEZwsYqCaGwRN9b3EW0F2BfxShTNnOq
OSB1LLciyOmRpFdekpK0MR0d9HVFLpKTSIr/T3BqNOqFWKmqBkXrMKmq1bFB1aRR
LhrLb/wqLj/P0iJAY9ylCwvXuWdRjNjzSOy2VVMy3E6xWdM/0HvTX3JBgW3O8u6h
E9hFJKG19nHuIWrOQM8xYyMjiOE8oN9j4TSSdaAJTNZSP/xfM4oFOJqdkWgma3Zf
fsWTBjnql6HJh0oERj/TEtDtBaDyursrdeZ490BAvzYXWjx/h7wM6UrdGY3PGgE1
SPa40UETZ3yP8asFQcVVb6EmmJA9r6gHvhEhRdS63TeH8nGDO64p9Q0oJd5JGI1g
xjIUcSqmEjbdTnsNOQl40VM8DFRdNovJNx4Fq0NX8PK+k0CNxJVZQ+76yd3wg3h2
gM63c+LWx5kYLpv1KNmCyIvgDSTVlpkJNxO1FW+YOPyOYvyMjbSk0mION39uDkKT
rXa0L8plKxVqxN6oaKDNVKDic/kid41t/5p4C8lduZeGT7+09g9kda13ZD5w/oru
M3iunuYk0pN3noYUWTmDEiAGiUDbjB2atVL62ZD+XPtxV+7DeqmHmWp2tr5RyVN0
zon/19r1gi6stL6c1ebfn1k2tZLV+VIk37X+nLXBW13pTVL3mt1hUsm62So9NdBM
G7BNWL32pinmbYw0NPEv5Vz90Wfdy5W49V3TJuaWju3dExu1Eaz6/rDWdVw0Zda8
V2zOe5DJF1gH/0eVV8Y/zPRBLtiC0eMO4oj39s2VOD6Tv70SAgQDIQo/RbcOdNGe
0zrMfO1D15x1l0BxyLnaGJyG85qnxTCrFCDYX9G9AeBF5CY+w2oj7tebOsaQtgTY
Xkh69Bwd01hJmRs55bOg+6dmHvJCA/NygPq5MD2cyG4ZGytueYk3tvaqheq7HyXc
0Qfo8vG2MYpPUJr+m1eHgaN9ljZPi93vSwCY0HH5JiTONldCWJdfpFXIA1RAD+Ky
MKuaGcQ/Os+25EY+rO7yLTB1MItrRyYyhtNnF0R8AAHjz/puChEc/qSReb7kil1t
s1RS7Joe+seX7E4BALJKgm3xNeuYxQ1EQs+BuEZllE1q9uw86i9TOI4n7xNd6pJA
XJ7Bs0VS0Z9A8E3P4A9YtqAfvKYFG89c3RnQ+f71tmP6kUzK6ZFv7KpjYwmBBWW3
9d743bvG2ijmgaZalr+yq3SzoFEQG99nGUlDE+T3LobrD3OmYA2+i/1Yymh92OWj
ouWH7ilxK23JdI4lgZ88RjoT68k0ehuk7wS6jcqsSK/OZETxgg3IFZB/4ObuKLXA
JKQws0rSIHiLY0lhzA8V/oOAgjAveFXp/V9CTafTMKh9GDbaG5NKpvQ8LLcI8evQ
iRGAjt1YTcHamYQdtD2bOt5D0MEk8xnhCiGZKjov+Ng+Co3kTizEejHC29uvrhXh
Gi5jYjiPaktTQw1X15vKVV6ASd7DLsfbhdZXKYNxGej/GcUoUDUm38rzWsSQPW4Y
z8bShaeMZeHWvZVMhT6zdGGAUQ3fTxr/sZuEqYtUu433CLK/y92hHVnsSOpv8m2+
5N9DwW1q71RCTSmJtr6MzkDa0OxKpAxwgZ4zZ4uwQ8CfZO0+6RC3jKWWRFjwMBmR
xNQPVFoEWFO6VwtTRCfMzvVykQUfFTbDgbUYuqp9xXtbbFyHRd8jjYf78Jysz9Fp
WeqkpHes8G9VgQ2dcBWu+ZXRVtiCDiyuhYRZg9kGkHe3A6d525zmGRHomnI9641p
J//vtmpXv5z3huUC55BvzXVwYE3EkSkc5NxdDlBM7GLC3SA6FaZSPhnZXI+T2Msk
akfkdtJesCz1YWFtJD5Q1CqeTSnT4filNXszAIDsvP7uN1IQNm19frb1QLOzDFO5
ss/zhC927ztbrNLNAsBlONyHuRccMu1iEeDVo6Xj9GDLBDMv0w46jYiz+WRxVkCp
x1B/Dn7XAhdVIiwRm2yYSHnMhDWxBHFhnyyAisf485ThS5gfW/PR7Zc8W15OvBex
sQhu7tQynbxSXjP1/4OxXLFc+sMy0lotZ47/+CvQ9nUXEIWNMPom2+Dy2tJSJWSE
8SKai6lo7I9EPstQcaXPQo+QgatVXrxErcGypJjqNTFDNTMjEFSZSyJ96ZwoOLUN
q1f91y44CmSnYC7F7JajrosayHKaDL1xo5eOgRgnW2bgg4A6++atDEJ9BfQ3DvsK
Qd1RztQEuigCbvhg0ShRsPUuTqIH43Vt426MGeByfU/vyNIFmDK1/70ma9MyORrA
Xx0f50Aod6z2QPkKjINz+kRkAGYgeYqWe0vcq9QZoq2GOBNOEnp8sScG9RIEV6Vr
nJLUKvdrPaSLRezckxVUX29WBBMau1D9Is1qu6fNcBho4TYNApxJWN1XDl5Yz/3y
6JJj+o7Us8IPLQqk8j9mG72gqDNxEbhYikvvICLx2wzFoBqNTqD0Du32pqWAaWZg
kVIHJCh+37hQQJU0mVQIj5qOPquEHlxn6Nj4dFwSROeMzlZloWMU1dxh1lF49zsK
Ve2rWctNFIb7fJPH7zi7aoGk+dO5SbI2Ct03zFxLjcZTnS1FHiN8yXIHYbJUB6bT
OcfVP45JL6q3f3jCyDRQ1ARKzmNGBOG7PIKVvssCb2aAyuw8N2/+QbYP3F7iphWP
U1UYG0vr4Hmm/WFlqgT7P5yPfNOHAdKljLBLsg/6UNi5W+vvStoubryxZ+fWLqKq
vvSLhAgcDpSMtJKD5RLKpuFytk86Rf92pqDbFIDiuuG7ifkyCf5C3xyqsaBFdnAq
Re0+8nPPGnN+2dKg1bpf6yZ29d5Kv16NAhiV/D230FPIBQPYmzYMynesznGjill2
whQtXpoWSNSc8qF0OS2+rrRgKqlmgIUc0Mra0BH7CLxwSKSD7CkdkMl7uaI3ofxz
p+9tlK5djzxKPO0KixI4sCUTKIHvffwVXJf/4ZzHOTKJfEf5gpQedHtsbkz0Jut2
sB1B9iIfwe06SkysdTry8uti72+U9uXzJvihMzQxFUztymDooDE0EzGUQXWGQb76
8IdiWAQ01m8DrOLXjl74qrI2XMypPuvV09YpKn+9lGTko6wMYHpIXiwCSmPg1J8z
HRLvF7HrELgwrAoiO/6VW9JxtJQQGhfwfgZWH2t7lDJRPymlk3SuKQy7qGhhex4U
fAVMxkRkZzkQapI1ClMBE2xUVYrBIvsl6fcK62vyH4dD2VHWmA2gEn2+1953aoX8
/YIyBJr5GAFzrj+BVSlYwHUhnLp16gIh7SkSsq1SSb6IbGTEXttK+BYJBABstDTq
qakUX8UIteq7P2pn/yPLufT5hyHFL5dV61FI6j6HSR4a7/pijuhlKINtqZ1CtYNV
h9cpdJQgzOHHRty9X5GsD7p5Cgzvv2jE6YjPu6lbJLQLwgsOFfptAwR7a/lfqP2q
95uIn/BG9cYAD4CO8AWWo1MTfQ3Mkd5EHJNvX4YL59O1P12OEsUm3qptzQ68pi/f
snNpINNkLytSsYTIEWqliqWs1qka0RXjjXbN3CBtApn5kDlm/ldUTGNNL6E6toKe
RK9t3ZRxaGRYkxsKQCb4kM0k0bwcLwwSyE4ACYKgTU2GZY+m6qxEPc083kmNT5rY
QnquHgyPdoDnUcHnZZkeIsmDBRLazVjjczetSR20HSBbdhyxvS3nrMf/dkKtgXHO
Nd6jOn/y1d+Vj6vTSx1T1rJuX3Tgja9LUFmCXjJea+JNpBAfGTAjnpagZf3TSyvs
kogmu/Dl/rM6Er6vi1OHNQZvFKlivDHQD2012LpGNQYxE0W8dYJZUmbMfWDdfn/T
ax6GcoYmpblAVMP/cvCGHZkIjd3FF96IOU13l+v98eBpJmPGXD82qTvPjvYw/Y10
4t9RlEwNcGIpsM8wicpySQHeF2l2fNwzE+bnL7BMoDs1gTKDnaLhC2kdcE+Sk6g6
h7TL26y8eWR3NxpewajeM3tCM4+ja4ItZ+mO9+345WYzIEvOV6O7w00Bkd7duFCL
rv7N55Q2wqvEAocsIu4mtQjGrxw3w+FnmdW1dxKletyEJXOH/YQ30FDY2Flv0k5e
WeuIlN0jzi4KJwLI+lFDb/d0OYN27oeoSONkmEOD2x71tBxn3pv3vi/2BKi2FG6H
kSnq5bcxjDsKLhisJmfj335pR1ms9SmFpM5jf+6D2TJtQMNycO9/765Ngxe0Z2xn
LegLRQdeQkC91Fl8SbqfmpbshjsmcXHPYN/4yxzBGRAfvwEKG7T9yJrpK70cMOrd
I8aQ60zzFT7sVTJsn5db+olVGDXGVA6LP8qLtlpYtw7b3vvy5tK9MgE73DL8STGg
ER1JXpWt0iCv13rfvVhs5/lTjyALxbxIygcjbTeuMmexhuA8EQS86W7zVS8KyGkP
ko7VDGecMTAg9j86tzC9Bp8cCIMkR2iRdPc6bHr9NENadS3J4CpyCyppKfe/TV/C
miNVUbbmwVixdfIL99M7GTDsRTHoom94VzzkDyJHNvvjJOulkCViWmmLPVv/WQ2P
GOZmFvDLAYCEPgIWpbYJBMVvoBiPnu84lMPVg8etiKxX3tvpK5Ij5SUrJ16m23VK
UJ6pKjvV3cLYFPqReJ0wYF1hfcbPYMMFJpttxwT1h3lAuZDAalNzeWNvgbzx6Vzb
cNLWwyvwSgA/LbjNGG4wy1cOXgFT5imK1otmmr/r4VY6y91rMnu++iPVDtG+J5Bj
3oV30xaHAb6C5b5yikLAhRm0FOI7FfNCIwMXoFZLKUMzfUsjoIJZU0khQjLweZaX
gxM7nYKLzEPFLuNgXaBiVa60v3aF9GvOYX8mFfz3z1RzT3Wcci3GZyR9KwF4vy8Z
LGaFFvuVbuvhObBb9WtmrtLrP5rKwn1PvUOOJb+JpivWIJab1CVKOz8W1yE8KEV/
kZtmMjJAc4sTJ5cPBk0l4mRtHFPlKUtvLe7CnVXDGrwO+LiV074GBv7b3PJ6DygN
s1vcYdykYMfAyLuow+uN/WKrG3ds+vO6Q1NIGGyf6NlXK2iRh0An1zDpnWBlG6sj
/OrOfGJWpxwFV7+fhODiFD8dA1gZJccZj9VgwLJycBm6fvOhAq/24nxLZ5k/EZiM
vdsoVo1eNwcOB5BhPm3tLWtIXk98wuCTHqzsjfoO9ODl8Dbp0Dp/5UddtmJ1HbfG
uWnUrHS9+nKSWFJ4q+J7dh75fbN0S6GZkJNNYb42EbE6HVHHsfm018fv0jy+NBd7
bQW5tXuYSGFAzlZcpNGMucn3ukZUb3rGBrcU2E6QCfsbl5YWu06CHnW8KPGHF+SJ
/pSpLjKD8taObPCW+FsxRuqPqdoi5dHgBCXxsPjxS1P+gxCaW9ycS0u5P8evp/2n
dSl6mpRl00/OEsDMKoY0jVp47rItKvf9Pu1YyR8vc75ZjTQejccqRXTnOmyR/IFS
Z4/B+zK/vSOT7sRRLCJ9VIECbJfohLsUeqJpVsfj3jqhbyfHXrO1ITnVLe1ePjQi
SdUQyrDGTqxX1NP8MtdiXzdUSOXDX/I+l7K2TV8KyUso4ypehtUKjhysRsNV6GRl
EAr4c/Ii9mc6LI5vhoszH6KoRuMIl537dudUgdcjdZXcVOcTj5XQVralcmgoHq3w
DUvXfYlX2rMS0pDVABl+6NG0xEwcB6FciGURvuJYGWzjAKetGlxzsU8ictl8iAMb
gBV2Xg2KxJ5SVlKNhRXOoVp2mq8LWahryD/LBOiRhmphiKLanCi+wkCAJk8jRihq
BnDFMrAMUzpawbrLOgEYiACdEvZe3qhbcFhYzyNkt6P7mSy1KgDYhSIY3npdBo4L
ZcfFmNabwepV8Fca3TIXXM/IN7C8Aoyvf1IUyChbhH++6aOwbqHf5qrqH0a2OkJ0
PDH07fCT+sxGFeW8lSdbU1leDMVIfXYtNYpdpz8zN7f0k7XkJcToI7ayw4WyMeXm
FfxwmQWan0SoxWN8sHhsfPlKS41nJdHy1w8hJ5FFPgL4UTmgzZIXQdHy8espiwBE
cN2Q8ZppS53h2Ko9dOGBdbAU6p7/NZOWk2f5r/PWmj2/BY7UY4UhZq2yHxEJXZTf
EB1+3mQAm8ZuLYkVS7J1qkKAhyL1EaBpQrWiZwsVWoP207RVuAGDRkcqemIVsLC/
qhmw2OhghtsfendqdIZ+c90kQfEDLM4949izpAUXGwMI7/l3wbcLepbgoTbB98Av
eVYtoyrqj/faGiHOH7N19kCAhEggrwwZwkC47svrJD13SP3ely0vxrCephVEVimj
Y89JfZ8q4ITjR3zbnUSfn76/EOGzp14VxSOfVBQ7bpIttQIfMbRks1oAb+EVZEZR
iPaxTdpVaozfUB0ubl7mo9nIsu/tIIeb/xaRgOQU+Ukm2PbVrA2d8NeFekeUNGyT
1ZjAJtR9NoKTK1aOf89t1YW5LJEHaZIiWq0fVpXk2UB+zC3/zW67E1LxfYIWxssY
3cwPNlWrhRDWuFN/Hv0F+KAzduagd6h29aMKdrtl2THI1l3XQlC0pbh4Omz4CCMT
2Uk9pPJWA+wYfUm7SpYI2Fc+3OZDsFUW8y+pAjbf1oicYmVipjXnVzDCtDnx3M+F
NBDrEjdPp+wxmoy4zQ87M8vjqbvCi6Qzo/1GUbl6Kh9iqRoCcuHqkKCf+hxkk+2y
SfBfh6B8Ulsy9JZP8FvhUXBvpyKis8dkJTEwyhZjK+lQXvl31qLLBn1/0XaieTss
DEahYIVCYjvT/rotGcNGQ32qX2haSOSPkjO5OCth7OeVP8zw//AtBf7ALheNNi3S
Z0acbVcDsidSu6HgtnqWUTQV1aKrgyiqgtlUgBjzOCbN2dDjV/nAhrfius+n2JsQ
4JlfFZPTe+B9tTMG+0d+pMQeVg4IhAqHwRZdwH5NtBh0brKPchFTquBbNGoOfi//
Fh8c63wBTPcobGqWrd2TefvA2y50IfwENQ4AbtV+U/mbjA+csMZolqYsl9qjpSwx
TqMvjqcL0i4iRz/hswts/Nt1/JVZrqQKPTCgaimbQmdyXyOg4OdZrdcRxSbv16gi
TJ8oBH5D9/tP4WlfyZj4kcmaQluxLDsmdmcjIbGY67UiPygW7OEJ43/E2JaXDFq/
3lShOt5z593SRTha0EkrbN+0X+PUB0M/CA4e/bwBTnoMHsiVFI+hoj1xhLj3hhQ+
LvaKJRouvcJcFXkkkgczd7xrWhOSQrMTl1NUhvB1yczGUmtSkttb9UXDi7kvYMlF
2Kaq9HH28/twyqQ1Wcud/hW/xJW0u1JrNjHUMBWKoB/OeFxeWZyQHyEZpDhnLC8P
oA+12Fs+1GRrE5NOmbumqB9KZxGMSOTOBMtLvrsmWbGmCviuDa5cj4WMCgAoxB6V
LxyGcgvnRsAIKCm3pE28hLQsgdDjjSA6C3b/sS7w3lKNdp926tmolh08Yk2DfAx0
PWS0bIvRcb9Uls7M9Z5yRAZbs7cOuAr3Wx9kfa8g0EHqyHtrDovs4phM2m1IN/fu
wyU2V2Hp7uVgC5ZVbN4TIy1k1ul5/aAYYQaaxJfwIYd9UFCQTWY8hYPuGQL4kIaP
/xFc7BHpYjKLcPw85ptBWoz8mR2Hq1XLmQJUUUt/gnOOluIw44ZPNBNIhB+4pl6v
SpyA5uuSiITuwgVOVtdDn5D0GqhWGe7SGmPCJlZmOjtgaFPe9TVL+pyPvBUB1XC6
ZDWkCXqshsqJOqT+Cj5JIf+AWUCrWhFvFvlvwm2/N8DcSHqTReI7YwnemV7T67u0
I//Sor+L3XeHSegcgQIlXd8ZFNt7VXWXsrT8TBaPT0L0D8gGK8ogWdLrbuwrugkB
MP7tMJ2RDQt7/zebrOtQjD0GdPC47Za9/co7GW5+kgdrst2WPxbO5DmykfN0nIoe
p5B0iNLzGTPK0ISS+sosiNRNqCDR+6usB1eLM0/B7MpysrPwaiqzKMo9tdBzubON
g0gH5bTakHy/6BwMSPlAJEx7NcWeN/Lfv+9DbM/RSulS4xP9tIwdq8ptzCi6zWV8
xiSad1ZIP/0oOT+KN0OsOaS9e4WbbWrjhBGrlRtop4jvhTSVEMGUlfssFvKOyHrD
WxvznAx4rwAfswOgsSjsmf1trw9YWN+MnGmyqKdHnWkrf9uMqrA58eQ2tS+GpXHY
W4Fej9csgOrI/8sJ5Hp9eNpr9W1uLIaQoXCnBsz0Zl4bLSE5ukX+V+/lExnucY3P
LhkQImjwupldArXNGhkQs4tVxgSjo7VMoeQbOGJDM4+xFBeClADxBUif1aTcKb59
z8wPVGfiL0pEhQQ8242SLpgYqVhGWUELwDpH1xDnaimEl1skRZ0xBWnPhGknITZj
FJCgnifsf72FP+nvBR2yajmbr+lg5OcAC4Newkira6ziYnNl2YMsW+KHzc0yruNj
rQPYakCZvhFthD+jP5b1iHM/4ynyHE49i0NA1i/b/L1fWDu0bJnY9Kr0ox1Izefx
CC6OBn+UxXIPppBGSxrKRBsGNJF4yCE+ponh8XDh25MXm48S17Uf4xDD3DDcO9qZ
JmGQlh6wCOjgyqvDPEC0rKNhC8JMuKoZG3LarJJNsqcGi48dzie4bTIR5GrKtPkS
7ejWisQu38hHVxJtmh2S7rftl4ZBG/kwVpU41L3XNvJJWTBD7r5SnxGZuDXlVM1m
+8RXj9nwPKxoWXZRqUJxFxC1YQeNVtyL1/TcoA8mWQrDgLp6qA1iNfTyp5YAIW+j
Yi0o7CteXs3O7J4ro3POVrUTYjS2/Cj+MfS+pn68lsD3l5XuBZjk8JI5/AeU3Mli
QH1mgNf4i1g9o7CXyyHgnVk0cIUUwP9l/LcCoCaxcV4wuLvWJpQck5NTrBiRxQjy
VcELK8ZY4kmBhtTLuAbMtCu/XcHYtPu6Wj0BGeHaqgZC6RyP2tEl3ziWIS5zfWHU
UfDnvXc+wR2CyUiTtS+Zjwk3O6dDhqEG84YMzzX0oI6oNhCu7L7HSsa8YSqpSCea
B65hC9jycID2IsUcqmekPy+Fws4Bs7fS4TrO15FpiaNFqOhxe2yufC7Y4S/qwtDd
1MTsG08sKwz7QwVnNTavgJV3shvRixgFEt42b122hwnRoisvlrRZepcmYKMuYLYX
k/CyWLlXQwazXU52Ybi5wzc5bjW5YQn0UmBnXt/PfxoNyX2wymw4oQrPf1htU+l5
yWBNbd4T8mcfeY068WMYabX5sPNWBt4+Qt1P7EPMdOvcl/NrQXu8UPVokZXFOIiV
rxqGwMmNQ092feivYJQmzETxaym/LI/mIN4iCdHC+jNwy13V9MuxPUuPDnmbN1jT
ZgdyKfbSXPfAhAiGJ6dBIXv/meC4/K0rsBQi/fCjInaa7GIBQazvBC0nDc94SG//
d+YZhoqF/8dfkEE2x9EUnqNIXQ6/Yk3NLM6X/Go6A7fVJyddEtJ6EUJJ0uYgFcT+
za8js5qi1g/OxcmtWNYV8e9IpXJEDCyX786djVn5yb57vwMC8XwUvmq6+uwGP4m2
StqofrJ5cHj8WyohjX+OpgKSnUIRKC0YhJCuBn3P1ljlCU/mmEaAh8p+tn46xVmc
oESgy4vU1Q80KU5AuFApYIjVfyo3vi9wRLyZ8FGvivpPX64jfU2DREfvazgruls2
8KMdfKnonh2w4TjviFRdZkVaerIT2AyyoEqZyzN76vM6Kxuq5Sed6q2efUJRjbrK
40UEYn+fs+f3jqtrai0vPVwF7yUtzqcZN2jpn4wqeFEZW9iGJxFFGBgXKRIc2tDf
fjS/hKpq/CDFcmUkQbrmlhiIOU9YQYasceXfYaI21PeCTf1vilm71exObYKm3ybO
umjOuLACfMDZQByrS1JwPdoqTRmoK8KVTKjdS0tDMtS5HHqT+WPyE9+4I9fGLvBz
6FdKaWC6wr2DI+F2YKi0I8rLyPgGmJUbWEv7n3pPjWU8JFvZAIsyo5o4NKX3365n
2a5A70LHN0I44NIl8c1bd5vqRmf9rdZ7M+ov/+i/Y5CHBv4jpPGIUyTXDlvzceR5
ZLkqCrO6L2Gk9HPQThLg4DcCtBIkdlOIGb6QnjGD29v3FLhvhOsLQL7FSkpJQoi2
bEA+GyVmIW4YucjYE2WlI2uKzCmO2j8m8He+8mfGeUV+pDIKSoBlZGDbFplNlir6
KMre5g/+ARnnedck+LqMRWgHPEuSiR7uaR256w28Yu9SHx4SuBvFL0wkgTyYg2YM
+GDLTmVuydklsUeXuLVbW1JCGgsUeCwGMyDCiMxKjJjmnPJAtEX/ieSrnySOyCfC
htbwjdTNs3dbLz+jwIZDgbAFNd8Iyr0bnWT5ZyarKWFgh2CF+4+8InS6yQidx/Im
SP81jQLyAkqvVRuhDi1oiPCcyUh5qR4vZrkaZQNpu6/ou2cJW808EaUytv8Caxls
aufQrumXTxveYgMHN+hEF9o6l5FXzE8yI7mTUpd94+IZ9TdYhPV0/Fr3+8j7o032
YwV5poCVjtYLg3lIQjhnViH9XxHybqc1Kj2A9mnQ5/rRAwcQHV7bsQcb4rIwbv96
R0PMWOGjRSnBYRoQq0uDPs8AM3XRGseb0jzthDz79d39YZObX/BFJCYtfBk/BERm
ldX80EKZQyTYIh2NhoCk3V1sLSfNR9Jk92QiemdzS+41gYs6IrvIZRczzf/enke/
97VaWZUce7USgmIn4Bg4NL9p2l7Yg+hUUwPHbiLwA3fLqhotTb0UIiuywH4mhyfL
Awfhq4GUyu4mwIj1Rr1Gx2KiwvcRTZwdhjq+m51h6jRRzAdAswqcFBnZ+JdrrKGX
jP7ZCjp5sF9NIQgGQcQf/cXzQ+P0pjeAqtJVlU9nHBykcBvnpU7IWJfAaO4kFw6s
ptgx0flZ1i2YNePzJ4SrE3vaZIkCrVcZcP0Dy/JJuRsI+53nOOo1uVpVhf2qgrtY
fuIYoU32DichOlThUQK8Uv9vlxO/DIUFPTscDyB2O/tc8siNBN5u05Yy9zBKVlwu
/MDcoYbU1nZ09fsypT2Oi9obvX2dotJ0lxN7YZQJ3A8C7vE5ekGUmFcPRsEqrooH
M+IMK/X5WhxpV1WOy/6fcAal3QXorqkHAY+KYdxFyrClNpXMiwqnfNWlru1KfEel
r2N8ykl3U+E7xg+BxdIpexJUuc+c77/j2xOJJeQ+S2eOePB7t+h1QBJKan6TDafm
3XbTWxKOM1Uqq+kOcXM0oF3yDhVDT5XXL1GkSRMFSFEE5ylf2kNCfb7SJG1aH12W
JlvlYvY+TjM+968OIjkb6gEioa5V4AYzuk4JvCOtOEzLw9/8FWm5EOSAyhQfAiHS
LnQ2uJG/iLGbNJAVx3UzUrIEb4ippROmk/PjIRuulpVZxctEW/4c3FOeFqIRrxXG
DYf9sLz93USDc3Rr16uBMuPN4/yNbilfZcO9lscpSkortouHdN8GQnYbuSyEWUr+
mMNubXt3kowfoU+suJ17h6bPfnNJatTFWtg38i4ngSoYUWuUVtHhRVmOdBtToXHS
Yz6BGhOA4rxr/00Xw7mNsS5VJjsZSLWXOjTS34bUmF6wY6Vc8lghgQXVJp2TBUqh
qByM9eRQzM71s5RT34AA0A0BacmkMUIvA6wGSOrbUJXm9pIF10CQjAxGpM1MKjjL
CZpZQrCKMIGbLMDIQcHqXTZQIIoG55rsTH8q0fg2H/Lw6l6jYP8MJ0MxEFM4iI21
d1vgpLdeZTQRMb5RA8P9RwZC5QZAzO1LM11e+Iy+rGjfQtRxswkhcA++/aLNJUGP
50APqyW5TCVdZG30C5a/LELkyZNM3wtQ4z4QabOJMgNUBkhJus3ncXZmMWEB06kA
k7EGQFtkzuv/pgi284sOLb8GyAjIsUItsy33rLD+XM6HQgAOueO4PUjs/S2aTZBu
wBoY4VVoj52TAViN5fWETOCsdNVzbVy83UGyL6NBv4ttpiviCBpjvvTF10rOuunq
5ptRh5oQDbQ+eQTy6MmFUq1qO5bomP/T+p9jfWuy1Jc=
`protect END_PROTECTED
