`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7cZvtbeTyzyLFdF5YA5c1rx6BnW5GcZkYw3Jv5Ed918n1XEOLNr8VEGSe5hl/vfU
2se7TQu2VaUWtlgP5maAPE+CnasoAk93G1TyuWj/SZA/qCR3zxu5sW/dhcMxn62a
L/Y2XQxlUEPfmu5XpiGeSiT6s7Mp3MQrs1hz46W3tjmUPVlFsTOw3nCLmw3B3LnJ
Pi9N8UiUF0ei8fRc+8GLL6CrsA05VMGW1nTq5eG8ojeOVBjenMG3qGjPH6oozYJj
hlXSqae3+Z27cuh/tgkqqrNRKYoYfenILH3F5Z2z1KQP1TlkUnF9hCXizylSQpTf
h/CzXduLCH+UAfQFvInFHgpPsa82/b6FkG7SfaJpFzih4Is23OKsdbveJxXeCbGn
t+IR9e+1AzLRu5RIzWUjz1PxPasOnFTsPOXZjQTZ9bNUufwiEUjb2Obi5kee/Eqm
GvhIKQwxm8e8hfOCjMsUrBbutK+6TDinjVxCABBqDV1UpWadaxUElIGu5KHs3LlM
PHBwgKt7XOE20ZJ5mXIRrg==
`protect END_PROTECTED
