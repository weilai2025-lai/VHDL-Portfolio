`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlOygCV3urbbpFuDuarSP/RgbcG2NPb0O0G6RLxW5Mb1IcjEwjGixAeShHfXG5B8
l+PnpkV6vSCWgK4JHTZ8Btt+MU4CJ3J9qKRunynQxHkdKubcEtECv0opVxV7zc9U
GB4AX3V+B0uTsZdy8D0d7IlV2RqxaqpyYGRLZEtjDX0esSfTntivrnca4CxFOHVd
e0ipD0XeFFKFJiGpE7alXte+GUo8KkZJRk4uwffB7gnuPuE1zLRWgnd8u1LaWE6k
JZBEICF0KxEKF6Z55PzkL4aBfhTif/HYWrfhLmVbMhCgOcXhYBp4id3cXwhdv+iC
s8n/RNQmOQFIGeG2s0fmq2CaV4pb/STXlWaT7UJGFujoK/EzXyVM4CfoU0wyWRBC
M7469wNgO+mVlyCApmqMOUsITh63BtdIg7EirP0aIaLWFF7bQcRx+8ghXUI43XJw
YbyIpAM+mJrSaN+AFH8Kdxyg/8Re9eb3A4CrBQUmAJuKz7sK/xO7BqzNFG6fRD58
B0KoCaxN3CS44zUp58d6ubzwpTeiLVp46mDiFPPwK1x/pEcBq5rdHuV/JF5sVdHG
3ukUPjAgl6zcQ7EuYb0YDLqnKGEl5hEWva2IH5WF6GdiHv4qr/NZCYhp+dbi8Mlj
GwpMVcUby4uPigBCoIOJX1a2eb+ti3YDRdIxaMVsDdGehRmDs8ob7SopKoHDRvq3
RwbHZyNWc+WfqzwgGBsusjF20T8zU3FEoa3UVk4zTTpN9k7nx4m/CkwTJ0MULnTs
U0urJQRYuNk+ndW+4fvWXRxikfVUeS2pagqSUlM1ng5pxGqc2M22gUjZPv4tUMLw
ZeUtuFuX/kL/oDKYx8OojGRXcO4/HS5Qmkt5EZeweVryU7XLssugjo5se85g7zuV
qmjWQ40xyuY33z0t+LohGfhuCdqrpRh1BDySkewJJeK3R9eu+BCK+9SibCJ8KruL
WNksODDXdtZOFEhEmbrdD/Q84EuVNducVpL92I+uRi0iYR/+06wGkLnmz386di49
KQ7r2m1AS+s+c8ZrSuprGNhfFFkc5OETHiqXk5cmS+5g17m5mUc4ZDiyvE7l9497
jxs6KCFH5//hB2YofUzESyIjdZyCVnmRCJ3Icom4d5AKnhDWVswb2G42wFUyk14H
jUlUDIHt4ddovp3KYOe6R6ZSPFHiHAIiu1m5L5JkZGB0gfVYDdP4Y8sjWKMz/fkn
BN/cD6MKJXePOJlSgu1M1ggMboOT7cLhZHaCFaLP45nwTP4qzySBLXgul7kmPnlC
nQd7GDf52eyKG5kUXjlcEVEzSQNX2bI7CuuDfEVQtiXp3duBBylslmqHY95Ot+H0
EKPG7G2eJqB58+sg8D1mc9nthGBdjRQoEVDuYCSPbUsuh3Rx75V6bLvs1FvPdFvO
P8cgHaobRvwkbTrJfn953kKOa2Wge/sm5OUFfI3Uye3wlgOnuXGB7lW/PO5Yq9Y2
UUqEnexxFIelulsM1x7zdzop0uaL1OYJAsXWERa7k3cHJcG/2fSRT1glQJOjjjbS
s4S0O0R3EvJcx45KA5W2GtwNpa4PpZPoRZnXjOnssSrP3tkJIFSgFHqaP1MHZRuT
/6bRkOtPioJyhiJX7cGu8uw5FyDo9ERO6K93n3VucXaSOSey0WERa1WvN40QGopS
IF4Odpeuq4bbB3sot2pV3vMhVdng9wy+ZKD4LinCaD88mY0GPR9eth35SAhIjMWt
askZC0MYCLukow3yqx9CHY7WyrFlhrBPwC8Y8CFlHu5+icodQPRT68cr8QLzZS/0
WjoRmQ0CQOxWTu2qZDVyJyLlxvlGxlvabfkAF6MbhbOb/xR5yAyz/0Ceb02wyMFF
KbANbwW/Y8UfQHG/6Zx0vFLH9TNiTgwStKIintemdDZJj1yhhEGKSNh6QHpPwPtr
WQJLkYxZYnPBGRfmVw94/PBPvRCA1aqRifuavxsYhEo61yk5+jGY17lGtz6Xxopi
/5JGfFlmyr8K+/W1P6wWWD1pPQ/ck5KJw9ZWKwxeJDybEbWzue962DLeQ2mIdyIa
wW6rw/MQed7T/GZJbpb4gqw5SVHms/DupBLflVCnkZpx94px1ffOdpa/xAWzEzxw
ivnEPMNSEv+hVs+gFhE/de4CPHUZ1lrbH9IL4RXgu90dc1tG2CN2AEbTPDalP0rp
tf4ZlViFPvuGHpLwQJNQU8KcZohx8OPa1aUHt+As0DVKMWrgWxVcsqm9/X9fH4IL
LhTxIRDw1cvp3m2F9golyzEQrJAULP4dPldFOYhsuzrRb58KpOVgXFflfp9MbMRE
vmj21/NKjdo5uFXLPBlN//wpWdknISht0YF9kbPWiBGWvbWV7KTWLs0ymKwM8KUw
JlBqxgBsp87wCZ6XRv/hjUNrOmFRkq9XCYosnB3bCvasMYgmqI3qvsfp4XCXlETJ
n7ZylHxEvP2hPbFiZ/ygkh3fE/HVF1uEC9a9Jlftg7oWSgL5fgX9egFcbmcOUvPL
/l4wPQVk+iXWDAUc7QUihVOOQLgDX/1rPGyhuJnz4ukV3in462vb8UUNcm0iLpSV
5O6jnz7yVOnIs4NdUEVktKuLrkP6R3wxbnhNIPIMhWwGPUJ+PZiG4Ia8MW8csMUX
+dwfa9xtDqJrXlSwuJwNTYQ7dP00LzLThMxDfrVme3VeoQScNy2bXH+pFiMLlU1C
GANkr3OTWW4anbg31dZ81pY8EtUdZ+t0k/TzDgzT/ZctG9EjILVVud/ELsnOe29e
H/Ja8YLBUbnRsMbneOIRY0oMzatyJ+Jnm5mPGW/dvAa4AXKzQ0HeUG0gseBHtTUS
28iBWeWhjofup2czCYuq6Zji/LmCDl9t7AI6bl++2MPILDESySpgjCFLZ+nDuGRx
mNzarJMgQ7ZpQoFW9ie7TCQqUK9ca0P61n7bowZcIV5dCSpmf+bhmKwCxApJ2qrs
idEcZlMUyftwBDtmuLMuJhUClQw3vKSauc9b+x5CSbArFECBNhNYcr1PBGhfPC5g
X5teNwonlQutafvaCHPHNuPMtgA86sFIq5G+nU9VylsJHj/glXUcybUyopyKoi2+
QAufplBOCd0OpHihGuqkBb8AQy/Q7ZhUZe8DwhiIl4B4Nt5qUy2YtvlWsGSTEFex
ftkSHCRB8o29STqJfFnq6U8s+yolQMYLxmqBqp8SPyiUKjaRjr0nmO/Df7v6Dtsl
jtTuChGA3slBBm7awCJ6t8wcGcX+aGvH13MLa41cQIEagczdZzOJWOk6MxMCy79U
4ufFK+8rkLtf2FiyT+rypC92KhrhcyjG11D9DkSR7WU9ywgUKmmNjPROo4rhLXfK
P2C8FA5lTeABjEWsgmqoGnF1UXiIpfR/A8Wt5bBNSW1daxlMbcH39ctVW5RouwoR
kWwGUv4Nnz8f1UAgFO5wpFMOTCjukUMyUdnwi4t1G/E7l/+y/7en0YCwB8jrz53B
5mHexu/eUEVP/15YXOwj6xgM32FZJ/0MfZNo5YBtRAwrToPMe52LWLEnw14JIuNZ
`protect END_PROTECTED
