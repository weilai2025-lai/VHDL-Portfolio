`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FdkCpmLavBS9R0yri1hCuC0DdGQmXlzhl3eEP/1Hk1jTbCu4S4olfMxhRlzzDqPp
0NiowUkhJsoP64RKy9vNGMC8DPLmpv61AZWtoc8TmTwWm/gJ9R4QYeqGL2bKJYys
v6oYAO0uVjZpDpJCmruR/CR6dlaEfNDdHAI0267SpU5+nWBNGSFKqiod72uK2aPs
GAaCOce8lwle0XWz588mHoFz1dbE5ktH11Njx6JPpJTJ+3qCUgCFDGdvsyYm/4Td
J8hnNywwYX58ioNFNkYqYUoyrkSllfzANT9ATNVNf0thWen3PhpEoXhjGXlP4UkL
Jg7kJ5SuNQstQRfLC8/49WNp8vdNJNdL0wP0owkVgHdxXTfWCQ+MD/iLWg/XaaaH
iQHU30RP8cLcXEmCehIubpsxGC8+s3jlT09iXRUm8LwoyB7plgggHGC6EKytntRp
9370ojmgiZJV0TNMV2UwRtfTJALOIFqj5wLmZtnLqsE=
`protect END_PROTECTED
