`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIH8nKzl1DBgAiE2Aek8o6qRKD2zcAu/fcg+BqiXt1bwngV0dhVZI5eNwgSnZedI
SrFSFrJxlZ9QRi4rRPWxk55Foj2cprWnX4wV67EFlZIKZufEd4uwzXw/w3WpvsJZ
R4l9yhhVwWBnFJQVQvWwUl9qpbXBXRC+saJyAnK5AYCu0XSENy/aJYdn/tHxdIm8
ad9t2pl/hBLYL0NjMRdhGOI1SuIhivIF/job43oXJQQTwBF0psjzny/piPHDCdjN
9oPuzHb/nHmKNW5ulNiCBLY0YfqNaNMZd71Rog6cbTOiNojYq+zuwnTnmQyT3ASP
ruCjVypDes1HNLCFucTbT1W+6TOqsDlZXBlDYbd7oe4nNeoWUopDxnPl3/fomM9y
5ogxWH8jYCc/486yR/A9CwCUnBar9zRmR+XXVq4w0slIZVti2O52fLXho/n2KNX7
bd0vTGZfGi7/uZwWsRafCnbO9YaISB0dIooo6DxYv3SqPAOYMW3LEbQsOsC7hKj3
A16xAjLA7fq7/1921gMxTABlndLTRgNeSV1aI5pf2g9rbzvszZhu+MCSQ6yaT/8s
tIuTCuSxR5g8FKQKif51uJHZ8TB73DBY/H6EEzL/Jy6KO93ZtskFmcp8Nmgqs36w
fci70wVK9WrQwjirc9K9/9FYBN+izOz5BnPhq1uBGKr0tQyTWCDQyRgmxlm+2aJc
xQ9/hlQgYhRgWNY/9Bl/uAIPJ2XCoBWlY3pCjqJ54cMt+dUJriWL0mvzuitHm/ju
y9Re/aBHbuKU/VuWGq2qrj4dP/IvEZIN5GWpzz9WcYt1+lxVkpvDedE3IIDLRb9K
KJpngcbURPJrHB6S5xLIxWkPUek6eXHXSprYFezhm+bngcIP4ML3QVRyXX20buL+
7sb1O5f1/odIgO6FKRgcv6N6ShClRI5dg95bX8UfD241Fw4/lDshnQA3BTDLe/AI
IPgNMBcEGojvV3zfH1RgEbtaJz1n7Thq0krcc5xEaIsA8VAEjZD8kC4UsQGflXPL
MTgym2spbyFRKsTv3BIt2GCMvxHJ8gN3Uak1jT21lnCbADSM9GJ2aQS+AaWBIsU+
cfFzF4A1l8WOhHuSLhOoJJf+NClkaswf7Eaf5uvrVXw/xSqT6Qz+XhII/Ku376a1
tgdYKbVcMhPhLYy27xxQgRufFAzqkP5269eRDeIucxBulMVZEl1onb+v/pgn4qkg
go10QnCDVWofY7eNmfaSqN0rwkK4kK4HdOlBWHT0XWPMQeedtVsGtMj9egLTDPbK
XNYNPOFK98kNnhCEUHffyDWydpbxwEEE+dyghd6UEgcQQ8zbiLodqHfym8AIm3YT
ZKwF1aN8j4jo7ZWF4Nmg8C2q5nVSn9pXjn09GH+KnGNoOXKXLhWgcR1vj/SXvcX6
`protect END_PROTECTED
