`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sTgmK/+aBIIY9H/VBiDxoa2DjYoGWoqEHqfXMPjPomLni9wGhT4tvXWqd4R8Df44
fdgX9AdFET9NUaCbTFFFBdceRAWzGRLvRqLb+t+T7tbLRxST+bUkX6CLLjNrWK7s
qQa6ZdHTJph+prlyw/v8QP/kI8FB61XhCbx0o36zReDP4oaNaHk1jbfqQn+zMtxS
Z+aSnSDsEhF+ijz9BLJj00umyhJ6Jqb834wIqjc4YW+qcvyydXh0kKaf5kuZ3Mk0
HN5zDGZeOplxP2q8VmVzNSRpPCJWSs6z158tsmGm0szGIUvgXFcx2mqEynecc7fs
cdDTtOnVs+vThm2QOejBpMtf3An8ZAIVl+Lxd/m/AppL6wxnvIRDJI13i1aYT8QI
dlPO/Dz+moynVy5tiGB9JZ3BdGXCk+cc7+tqdGadBtQYZfMss0jGILqY1YqONaes
wmGrhMWOxWbXrniCzIIq+Rbzo9zbfPHqRCspPsMPM1Wgk1X8G3UMVtOU0NoMQj/m
OVRrGAh8gY5XQ1inIsExTtPNpmC1FSu0TnmILYnZqQtsrLFG4RR+7dCzkQMbE3YH
MooOSh/2CNk6XntKQiJmGB7cfTDhDCDV7zlPL1SKjEQ7437n5RiUUpPC+GHI0akp
LdQoumOwOU53uIlJEhS2y4zBNQw2mjSeBaQ9PoC+Wd+fAK5SFVNq1fGuERfUaIGQ
MqV4hUYrHmTss2yvmFx6El29Wi9OOZ1+b8keCY+xcjTz8fnWiUJk8XuiyPNcxjXU
w3mMbLoaxN2KQo3zQIowgkhxMB089RYkjRgwqcPWtpxplHo7Ym59TR9KEjVTd7Aj
vzD4yzLxmhLzIjraSJg+lsHZR7jyLi3hxRPOkZv+029pTH952rQRlKnCxvTOwIZ4
TnFNbsKmi1R1MxSsuwAxHUkAmYWVfveWd3x82t6QZ1cD5R83xbWF7psc8YRhYsNL
RpjTtKAuEbTNAEMZwPxt2MeeKrceDCVZEJJ3KkQjvBUnlRDPN3ysXSa9M5tzCKtG
w26Gm06X0SOKeUb1mqedgsGJdEUopVph17uVfJm5AcORoOCgzaCMy6eoIj90b2v2
tmGIpK+VXDBQ8KIHIW3c/ApqS19Yao0oCJrCKOBwVfIgbbeSc5enXCb29Aj4bpqo
17EoBnpv54UwHGU93eYTTUv8uytGdAlK4jP+Sm7xnR16BjCXim8J9dVfXVTfm5oa
mQGI3C8WkpM8yQrnHR7XVzk2EGmT1MwakydzXiCT4cRe138vEKOwPY4qPPZRlk5g
qDONNYPqmr2DbPW6pNZPklHjEjIH9WPQ3qvVYh0uvsju2bhUS8rRTCijOXClguId
rTWZxnX8zOl/9ZJOINj/y33kNX3IsWBrmK/TAVWdNtHfiq4uOJc3BcNEZ6PV2nDW
YqlkksqxJ5478dRV6KZzg0b2QT1YnHWYocfqNhV5LJ2jHypGXkxXben2EMctyt+b
6uRqS1ydLhB4j/WF1tMnijvhKQ2LpybD2HNLiJl7lfgNp/SOn8kZDXu/uPROUh1S
ujFEAYywNP1uPrY8aBwQ6SJKPbWo6+104na6mt/qIm5A53ApRqC5S97nUs8gHexe
WYmFZ2wMa5+WD7/OHHtHQuhWtDUaLGiAVaBgSL1cpGO6KpBvMuNvFIhwcQk9XV5d
wVQiZ+cFFW2KmDFoZgfX21YA0zHsbTaNcpGOALacoPs4rP6tIIa06yYmpgbzjzDh
cf+jjjag0xNOSHTLK4qvB/RhqMkb9/aMOlearO72PZzsM9uA9FLdplppWLwjLciO
bPyAHoSVp8nH+x9et6t7+XLTQu4BAmZDn15y5OsLOJZQbXCVnqu2lPu9XpIrWYqW
gthZhsqJ1nNAGi7f4ngwe0uOvZp/5FGlHin66PEpYG2svNfaz6jowEYHxCLGW1Nn
Waf36dNxRjBHBtS4/KcbpL/xlap2gFoUQKAs5TI+sOUyRz8l+XAsyRkDZMJszQbH
DbBSSAiLY83elb98QWW5ce1ax6uIE5daiUDg1toFQhrIPIfIcxaGtVtWP2oNE+/Q
B8CvpQ+n+sWzaTqL8sVS0ywEtKS/4naT63gRdlw+vN86K4UJhYOLsr00ypr2cDml
kcTh3i6O0Rl9zplfLSFRZbpuhA3WVhLpdJw7GKKaBcroTkIhqv/jIwFAaPFLVmA+
eSrL7ZtJYi9G5aLCa5AT3EyfcysuoX0m8uB696Q0WQUbcDttwiaS5/VypxLWpHJQ
p+NeQuzkccmWAA+cq8kMqOgGKOj01Ux9N4k0AxoTqzOrrWmjksRP6bRTf7/B+5jY
94iACDtiPpB75kiecn47LrE+ZDAcqcSjmXzWo8ZTK9kd+hnIaEWkFngrQjGPv6o8
N5EfCKAZSYSWOmwfkA7whW8S9iBUN1IZ7sf68M/QGFDBxX59Igbm9EYW1d0Q4hE0
xtvD8d2xVNh/WJPNgZgBTSXz4Wbiy2yw5VCe8NcJguCn4QVDrbW+qUFC+y3hBJFZ
xTT2dfOGFKVKvy70HzDfIrQEdR4uhw96cmBEkkeo86+wS2SaIBorGQVfqWVo7TiJ
n8WZTRuhqlONg8co672PmH1BciFecclsKoLJUSWJkONk+0cn2QhtW3aVxooCBhMt
McWfjUb+6AMqaTFj5hu/A80kfDIbdCja1GJW3/0wGkTp/QHlqnv4D0H0uk5AN2Jw
HXaMfa454nCKDJnhqLnK/h0WfNj/Tms08+g3LlwE9Nb3MC5hqs+VueqYU6chUQrW
7nj/mK8hrJf2oRAFGdJoPl/ciVzfJmDTfQ8ap0kXPHY+Y4wKR+lTVL2lh60HWnRa
0D8BfeeQT6rjGcy7AL2FMlCa2ElcC7nMm2fXyJ9jiMddW6ZplqmANGiAgD0/5bON
LL+yxiUQS7m99G7/83P4+ABlD7Swh1z6Mad3wtz/Tmhn93HvXC+pDCOaspQzBEbv
pXfMhLobsv9uZhCUZO9wTZYH+JJ6V0uGATaPAltsSuHqP6vmBLGLl/2Nm+IM5htA
`protect END_PROTECTED
