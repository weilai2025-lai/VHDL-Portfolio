`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAfUw3bAVFQrJSQnIMxpEB28gJ2cwxXUG+xa0ZpAu9T15+9yjypYoAfrHlWcLY21
lEFdsyO90vyP5DX2sQHSNQd4YV3xhQ9aQgexQzreGigsvUQTXJRhJ6DgiTUuCXph
+uXNWxDm+HP5EvLg9MEprpk0hkYF3d0YizoAXiWZEiGp9Mw9ox3iLOiYmaQxSo9y
LcXBTHc2BHAde8fgql9zJhx5jvVbnrWgJQvRExb/91VcIS6G4i68JEeCq44qGemH
bsJbE9gRdJQZR/hS+40KuH6HbIWAOPc+MWWmstCFha5CD2n9iTztb12eVia2asIR
l+SPKLo13k4TGQW74Jr+pSFJv3AlCQIJNS8++vXUjs8/wrz6CFgTa5XJeeoPooLu
+RsEUZ9HjM4VAP9KX+KWMlyVJKjRY8crD51Xif92D6KYz2iFarSzlWGE02YmaQaI
MH0BsI6soHzmd83qqUsoo+hBSJHbcNaf3rFCSvLt9Z/QGWdZKMwU1iXOJDvIpsuG
X+RzZWTbr5RDW2xAq5gk8Twumvy3ByUPjSXkq/InS6BUGIh+vagAUV7DyfleWr8S
aYwVXxOBojvkgfFN3HfPSGkfDPJ2qD0Dj9p0FlZwil+XCnhytZaE4pGYBwlhWFWg
5F1s0FDWU7Aik6onYUkvOD5aufd6M/KDVfyMbqLyOAUSseFbqKzHQlcxdcfar4Y/
QZY1kP5dScHKQoDWFmPsriNf7U1PdDw0BcTQvifM/imravwGtJbt6HftEYqXaGSF
ub3O0XfglOOT7Rt1e1SDI0UaqL0XltRXTsQ+fYoTnA22vkhzjArDqfPy8fptNq8F
9mY2GJ2+Iz9i63RnlkPsBckWQC/ye7tnx+kvKAnOk4N3qjcQAwLMEmxNTZ9bdRSW
pF5VqXkqxgknLF1TvJeEsfY70qEdB4cEVc5Vy36U3e2eUbwRo6axXQ6tbeduUcuB
u4uVRBhg4i4pHgtvaszIIkmQRnOzv79Hezo8apsMJas/tP5n8CJp+z+M8NzcAi8h
d5q2io841+7V/ttyyACDuwcIYZtM/mCygsjAQL7rkmcmxQLvpMy99s0tWl+IAhbU
VScRsW4F1bu34yuc58q38ANHn2/F1tBEKDibuLyY07x2fMX603vbe80uQvzuN6zL
Wh482lR4c5mEX1bK1L7W3/A3QYTiD/hBMVxzNJXZGo81JKn4fxeCIdMICvlNfRvR
9xRjgOxoxWAisWunJEM2rXbXlH/ovmq9VKuGFnOKjGfuC/G5Q2JQcJCecmvYkeZT
7uZroG8ywv71Ls7Y3tRMqg==
`protect END_PROTECTED
