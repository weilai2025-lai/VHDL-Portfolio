`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1QPdm4xIWBUWb3B8HAID1r8PR9qTxGPgGL9a1EK3HFnUViZq0uVa8fVf9cJfTAWn
38ohyTdDH/3XE7T/npmKvFAGeCUDF1sqpL9R1O/ShkOFpU3hPVIOzxmyHfvfuDR8
1AtIi9H0CoTysHEdeDkCyi26Tj3b1JHV51IqdeinJaQxJT8TS0+ywKDMyQabYrKK
LFftvptjBT3cL3BfdZdOL0hiHPRGB/mJZnhqeiT8TzhvK4Kos/8J4IgI4eol+6cO
E6tm8pinz5o3HSutIx3mkgMTOluT4AApcY3GVZoV9ucWVyu/iokhGmR85LMARe6n
jS1SmnkUsFjG12aP+qn2T7/Hn+bZh6DFlmRq0wYy1YYIXr55852718FlyLz+iDQ4
eUHaR1ynAqnNDZf6SGEh8SwWbvh4kCEs/YffjPI5usD0dbg74y4EuuqT9Eb93M1+
LrHjguZexHaAcZYaGAlPmW0LEniGHIrWfUcmaxuNjxc=
`protect END_PROTECTED
