`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qy8GfO/uhNlWKplKOGpg2Cj1vLVe9AaWIXNjmQqKwKufND2oWaM9jjwX6xcgLwHY
1mMoQqspaxyEZmhDuNhoQmStQWe1bXS4GTLSGcoYTd+HGcBZiKMMu4lBG+nSrTbS
2ftsYt78Kx+WLl9dK1cTaPRJgzA/thZIjzK4pQiLL3ot1VNU+UMaAX8BEpE7o2Lu
cWVOEhBXrdc5giAzANERiPAha+mqPiqlgAfgVUIN/5PnTzVmDNVAP03C6MMVNMMI
KoQ1J+DAQQ/LlQfJygUpuZ0wSZA7MrzV+GG8HNvN/YoMiYce/l0vOS4EZpdP3G1q
TZmEBvFEWobuM4QaFux6TPGmYJVvCJa77yoOB6m5kR4Q0e/0Rqa1ss5HCsGlXldM
1R9Iq1yYO4mbLP0b8IkJ65tP5+pckbXpAfpavCprJUChXgkr/9vgrCFZqW/1PXib
v0Ucdm602Y79iUcFP+L/sVT5ff980m6QumEIbRqwaUjXE6a8A+Z8CjhS4QLY37kr
cmGXbD3vKmnLkjqH5CAsgKnMLRFZ0Vrre2xv1kUaNTahxmSO9mVS5FLOVUbm2l3u
2g34YJMz+aCbeHMjwgxEwmsNfF4aO9XY1wIfOQZ9xpTTos5yDV3lsgvLhvuVg9SW
2kmWJwuwvLC8FydrGzn3KGZkTBwIgGgc0EG7tQfjyn9+SAAEcOfX6Mq8iQdRKf2o
u7Znu4QKQ6ck7vJ8snqu4evjBr4TWHupP0UIl0CCWudCSFQZqjMh/69g/PQjlHbG
ZIF+dJ0DMKaoLEmUU9Y1jwiiTvW6cTJACsc42ZxeXYBY3jWpIO49txwaHdnP/9i3
AgQiW/eMcX3Etd0oGTbyEKCNOlU0iggRIXUZ3Qw9zm86LorrJ7/JVM/+c9gVF+ET
19mDonp3xKXI6e06B/ygWE+wbYbpRIHLNIWs6sZHZ5Gv/vQodd/TqXmIFRhGe0eW
Iud8bm3cJWVekIUgtZ7NIaLQ+QLpsOcubatyhuQOc0j52lkVJqa3vGESmdmFihMW
WOqC4LvCnMmqNyLXJphaEb9ACbPMB1lQEASa8lltUsPWrA1egxSOAobAjCytf+kP
D/MmEkyPhIXAs/PyMh+uP19p8Wl+Vd6VZYwKPw0F3WfVS9+t0c0v43YUMfyqiCWs
NUGIbYbkg8iB3HC0rAfbZkHuJJmxZcyOw+C1PqEaUrGFhDxLBHBV2+oeOUZcmgJr
sNoTbMfyxgILocl33hvWTYzSJIgnU9eNNWLRERukGGSZ0vXbBlGetpby1FYPiWqf
VWc7e+/UAU+O3C4FVdMJRibM0gwnIlsqycsWpF/oo9wYY+Cj6cfw2gOWGaDdZUuH
SG+UEpiQqibB615Y+5I1QEDEPlXdcg7nrcR1yHG4uSCuQCzCMwP63qcr0nw+FCjp
XqMtvUdbXz9W9AUdDjJFGwXQoao2Mueb0m6aSFRC9BTUTDP1UmgMfj1SVga7lk9u
SHj8njCFGl0QhaaKTyFpOgC9Hrm7Y0QMsjDyt3mBi+jrYCr+iRiczi6ndp+oHUis
ibpAE70TwUmIEcxVTSJtVu0ySA2fvOSGuLADdYy0DTztuqA8/WWWrx5Euk5ZJ3Iy
czoONTJMk+okfN6Xe2wq9GEF31lLxltMDmLRdW2UjjxtSd9469ovl17lIHfwy05i
npgeBqyeAAdcO+D9YoBk5y1hudrmZSi5kV06S+z4/1YGzGbl3BRo+HdZhyUYHGIo
W2cm10qFQzNp2GNl0XYP4894WWWWz4brlZWucWum8QeUioIdLhxpBn2avOGPLRLH
KrLqQXDrxJmja7BdZPBNy9qFdXwtaF7yr9W54qBhtUCC4QtBo7iwt2uhp7zx5DOa
Czje5jYKjNBkTrX0vgzEgtOljdfg4Qe013VrOaeluebiRCrH/t73WRFJ7FA+lqch
WAQzBHguyT8AQz2T4e+rz6oQRcCkHEz7zW3OpomRjZnUT3SrOhPw7Ns/3IEnHiam
xW/ARkkZ9fJwH581nhauk9Q+Zs5Hk8QYixnNVq75KT7gWwcqc22lbBDCytVN5IIo
jIImnmlVXfEYz4QeGQausA5Zj2x3YzuFTHxNjKvAB4ZQdn6XhdqrRKBdVStEL5rl
UG8CRPYujW8y0xGwm3aTc5LKgNvwvmeFlF8Kzl5GSVZDuXiGITANP5wMmHrqrdLX
zl+REsmEksmOvQ7NcEmgnpweZBnVMzr997ZOmBD785bswBlOiRZ6+SA2fbXchIMd
5ceQBwfsIUyj5uOQNd+GCM3McHtf5fS3Cqdqv2jyWG4pEQ5DUd0qSunl1JfdgxPQ
6x4gz5mX2RoXbH/PIg+b2evprepNEOTXWilqDwnbOz7DLYyc4wjv73OAolwEa4is
nBWUwjWHrao4oUsvN7Z6AaR5xcZkI+bVOrTlj3hXeuKvwokqExSimJ1hxZR8idGR
zx4CCz8y9cDiqbKCJGALmibbB3lmSNeSmMoSHJuW60rt+JOS4/sU50660JL+/bha
o21CpruUM1Hr3mb5KXo00cMZ8w4rgUZPMuhPRpTXUC2IEWwl3ZoyD5LRVZ/E0yIc
9M4iuoGzs7ra/Kv9TGRN6xGNTE3hibDA/9pqhWJOCYVKcCg9Lcsn6RsBtjtP08kn
RKzWdoUt8JdXeso2zLyLbUDsU46oUJXXPSzJsh2gXpLulrkrJziH/ES/cigUZK1l
iawJEx0BZ2tIohgV6GiOzXY9eRQGl6pQy91Dno7nFMWKZzgeBhNonKxVSBcXiyyS
xhMBw+HDRH+qnjhbrofABc/YTSQp3aMzTJKGFpPYGPjQi4HFbFW9GcKcpyieU7R2
8rzGpJFM0uwJVAID1438NWhKrJt4vzlHbP8pQfcnvKvuP1qr3NqCbP/ZItuE9vLU
aQ78BhXAIsmiwkFeBCRxCFyFVLfuOgG4tjgJILb+LGmKOPUCoWa51S9fOByf4Na9
AYOEHoIPVgcylC7x+xWj+jJlY+TijcY54EBBpdaG4EgJg0t/Kd1rnKMNkQcsgcuT
IYWQsj8NNXTYvf4wjDCfKUITt/ATlSoATbJTjIN2p3lFEsG2q6lD7gwJt3MEjapp
K+SY8O+2VnpuIszaIAY+jOxzO/KjtubtNUVxqa7Z29yQ92dTC+9Kbmm/HBw1VXHf
OgzzVrWD3s2bCiYrzyPsO/0cyK9Sqd78uwr5Rqb4Nwn2/ItYS3y326euCz7tQDHA
dzLNZ070a2DXLD+7srjmIHqqGeYJj9toTL2FlSn7/mzf4m+FryPsCF92T/8fy2ab
HDuOAeWob0KnNmtPEqQdqb2r0ykGUGNnk57UIR3Nmj6vE5XfqXqdFnaGQ8XVTuFI
UzYEHbIpFvCFgJVA3FkmADCGmFsuBQKEw+4xF5iGSXygKOANob1ApxZ+JWCXgYoc
xJXl54YcaIbakS9h3KunXmdhPetaETNQEfOztxPGFtTWTUpUqNUJCgUXWW59ldFS
`protect END_PROTECTED
