`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sz6ra9AiaItSEuYz35E2VkYjbduc0zjBlHo8iB9HJziYeuqMlQLY4abv/ARyPZ+L
J+13bPIT8mjhRkS1Tv0CIGOIKks0vID9kN00gsyCm3lmFe4d4f5v7bXYc46GJtI+
0A2TSgVfaAj7Ek4jTbvc8pYkps8yEQWXbkPffXEA77yXV/aBq9Dt7U7p2bIzCHcE
PtovQKo5wFEKglNpdllxUYrFTcwUpLe0+Jrs/mBNkzzr/SD04iGDn/hH4Mvj+JYV
9xsHpJnAI8sUEtCTgQDy+Xep9E9/SxWVLQ4EcCiBHYgHd31lNM3gBkrDiAZqtkAW
wfDFhA0SzsWodChTq5K66qODdV1dj8SlzrzpXXYdtRtQHMtHMebC+cK4uSBNjq+R
rfunyz2/Q7z818rDIs3im6wBEWrLbpgrGSAK9LKPCzcb7NupisQGsim0fHS0WrbK
FastlB4fNmeEe5Iw291jG6fUSuE5LoyknnHPsVQ7987msKN7BJUMxFOOKw0/wWFg
mBbje7H1N8JKHeg6kNvo4nkASnPKOgHHo1QBSveLoSZjMfVhnMPhC+qQnTKJNs3J
4NPZKUrm3izdhMbxaopmQEhxC/DAfHdJtxuY1DI/aa/3cIGGBHqdimOKlUxIQWpW
Ke+LW4VyrTeLn/CwWVnxtwzNwbivQT0kCNgJz2KDZogY6Y1k34EidNcRiHEzvpZm
DanuRgyvqlonRJrESyuZt2nreWUAZ7Xr2BQbiIfvX5QzoC/h6L3aOo7hNonngJUW
Ua1fn+paI1UQTKpi5Jw6wMtZm2tsfu/2IgNFrh+sSoeMTzU+jfy46lDW3u66fASj
A17UWXFS3CofgNbFxlUtbEzCSdAPFkCUhwDe7/x9XCDNYUbSO33Zgby69HKGE48O
rdwANRXVP6vKqs1nYzkNCv3K8I4OIuKl2tI49xfn4Ezn82jBm2YcLfZCSJU3nJ/3
bDUUY+m8DX3ArUuOTPaDmhjx0yif2DdF/hrL8aw08Spev3VXwYoDFO/AvjzX5PD1
buHvsoI049xUpNCaQWJKQDmVaPBjctVz0qNlWYRdvISfheCOi8imMShPNfmhMDvm
RcXQdy7OndvRJtztCRIZsT95hWq0UZNn95yFZx8FXkC1VXqJQ0tk9mAitGHPsrgX
AdJO5Cy74wiYYdU45xkxpOnzDr+zcnvDI9Wc+kn/D6Mo3LRmTl2quZIoaPcBzZyD
sW2nnxJQugsr63IhRynWoNj/D65i+sDaAKRDoNLGYGZb6HYyyLDnNKM46FZKi6xd
n0BtdQULGMGKqcjt+3HMRUP/G0TvuuuB3rmQlTS+t/JbLhkMGkcURKJjOolq1Drw
mwV280dKsnYEY8BsnzqTm2/VHvOHTvZtx155I5VN3Q0Njhgkyx5T3c66xsRHGvL/
MAmdgAZFHxle60ZCJ3gv6jQ1cCwcCCfbIXQxr5KkchvT6xYHhEhzNdbneQ2/rE5d
IhGacOXtEZL6PVGv91uoGD8kKnLILmhWn4BnX8aULof97Q6JwQG+xuL/mhyBGYD2
oyMY1LirQwQXr90IXuC/pZ7nPg5NpdfP8ApJ4vwAPNZlXVGoyhmlbOnmdTnJavfN
6quVKR8T8y4p1ti7O5JZFRUKt5uwk517umjo6XzFsHkjhxDvpG8k8aOOxe49SlgT
SsS3qxAqg0AGzDnLgPvl16av7hsEk1pCDtCfRQEU+I3yHEcqID5ifmmBj+e7S/Ug
PemHd2U6Ae0A2Vc2naLlKfONrXnaiYv78gWysVd3DtI=
`protect END_PROTECTED
