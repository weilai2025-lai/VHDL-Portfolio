`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRhe8vaW2hzAn0gRZ+Pjf2++9HGEL4XTVeygASyh3GyMl7UW2vuse2CW33ZDAZnb
bmz00OcJI/DhAwyOSvU7oGPmWgijYao1wFJ1VbQhDArQYnCdo3DZwBAQ3a55mtK3
Hn6oftmRQDNGXzORYlmrW1f/YhXC7xp5RIX3swTWHSfrMCE2yRQkig9VSevZ8zFw
ByLcJWuKpHPtiEHLWhQbKTlpW17lsvw2OfAeLrQ68SLiya2MBeqfhK0AIsKT3V0z
o9fsE0lz37yG0lUGCf+65FJyx4zs/H7wDFbQnUDtEuHAaeVZe16JMgHWXyLLqfHq
cp5Fquvc3hWqTjZXEveZ5xoEC8Bjam0WF/nPD0pUEr9+Y8IlMV3NeI82yIRKSKl/
0wsy91Hex0Ew9QgcLpfeWJtl/CqPdpg+psTzbCx25iM+UQN+J/PD+ZiEx+29JJ/O
RP+BVMj8GofJYodzveR88ej1gWsApdusdsOEqKpsmMNO7p1Dd+ik0NO5VOoDK3ir
sVIogindB2DrLjoKtnmuPiim9xhqbDr5WrCFJ+/Dw9ATtpRIUK5aBF4+ICTg8dTg
ejKUpyhE7xaZbrBP+W+MTIqBushZJjhbE5YT6eSMreU7jrFQidCQ6Nlf1G/MzU4F
tU3Km+1Y2QKP4T6G6+8jUyfXLB0ImvUicRBAys7IezBObfG8BS3hJ8aSnRitkV7Q
GHqm0TmZqPQr5N21X7e3i+s7xWaGliUKKh5fLFe9Tluu50YWLNq3cAwL6xrFnx5R
SPeXIApS+v/oZrqgr84ubfOtGG9/Uc19eT617ViZEvRKV3nRIlY1HwwFFQHsmqdZ
vH+qI1eZeRkSIcoQ2SrYmSC0U77LSXR719r8sOS0gskYpAohV3pPdSC0bkGObHtb
IVmg0fWQSnoT0rQL+qMThMhuKJfu90vTICpQTaMpzye/uU76DwynKkJ1VKXtWB+U
lc/9yi9HENxCRItTV+mHIi2d1xiq+y6pcn+QTzmwttYBjTPJBE5EVSbgH43d32rC
bfvN7p4Oe01c/ONjElhZZXAtQrOYIYrnFGcDyjntT8HE6M7R/H6AlSj7cKtQTV6L
YztZE6M3yTfydWSz2WfLL8sZsSRmn3ftiDC+N0srUguJ59goLjzuRZSKKmpvplN/
vJPfF5wh+ko2ciG7NSxMj9uOj2JRVO1Vn0Wu9RKRMAtdWQwBmOMALRBiL4lYQB2j
FYlrsul7NMAcEIZcuoSJPITr5UbS53y0NF8Pc0ar8pCiMW4RqsYYLqxeJWTDBxzW
oPW+GYkYFmdX3+uzCGHnnLmlncknCWKH0p0CBYJgvEaP+PnyX8ZFkEfhcDeEo2/P
YbVXameX9+AekA+8EdzbjoXiGjL3f3FzS0/sa9NkdfcpweVWeV5T0h5icHzwNquk
9Xr19Q7fxpycGMv1QqmXDGGQMSNK4xcP9HTorKTLV6OF2uibaKemyhFU1ikMK5By
MwrGzaFjGTS24+XRvxQdYDc7AyqamV/4HNcDUPybKom+k8l5LBiWdnqXbSwS4KV+
IIpZqNiWNh6/ygyWb0c2iz6vi4MhaF+c8w+IIbaljNvTN8kBzU6msJTJPEBKvVfY
SQX2PMaiw7xyI7CECBKpf+qsUphtkdYZGoEXfmHqBRYZ+5ADsMDQv/6gUfttzPQK
5C3oPMNMvR6IVS/8xVnjxdh5ckEq9WoxhtdoHTNDrOiAaTAnDNnzHtUN34mNcMEy
CCkh71IcPFTxJcDUzeX2XGx7LY85PsIemSMlFfM3MlCwdgZYboQ9/aJr9X6qzCXN
+AXptgxCqH009EO3R0sbMlb18uCRjtqwtDoxDeIVxLFhepM0EuW07kr+qln7Qr8i
UbkTTDWMQBqXjnP2sCLrCBHv0xvD4/rDWSZRhmAJ7njQMMsZSrqYffPeieI+0HmZ
HnuKIoFTx14ThByq5tVGBGa8FwnOKgY54qdJZvaGxPOmVpZGF3yDKCqkgIUFpryA
2yek4HX5118TpOJoDnVbFxwxLN+0pzFs6QL4HXFixg/PuuMtRc9GqnOXke1jTRwX
RyCasVN+exOOrBxCduVUC6qPrJEw3vW7gR3XglDc5AIdhl3R+cw2cXHJygTRJ7x2
rnNXxZkH3wKUtiWFk1I5l0nKoY94o0780HV/nR6nklKITNt7gFDKvBWznqq5dRXB
u0O+zH1KJTxfj+jHRSzzwZ2tX8+88mCdof2mB4W2Ct0Ed3czB5NHWaXmbMjowK/v
RhDVvTLc2GijspnrHAClUV08QthoZczinDiZ/HkaswGIGOa4TTgKQPLMYeDdrn7w
+3thSwe4NW6FNhDeonvx7pX3rHmsdcSlJWPfHgxbB00Y+2W7HZWI77fXFA1sO1lJ
gG1KZdTaHOIyJGX4zV4MNtI6VqgVaQ9FSDjwqBbPf5lQwoNeGZ5n+fd2F+N+Kyvp
n4AXoKUj+FghTjItkzZVjlJueb3uKFjfHLqdQn69DpK0fGtAsdHEOKPP5lU3vA2H
Qwja4PDuEhKXTeQUDs9YHmf8VZShlSPRoCT1Vd5oggQcakbXJ0f9/1rYIyTdK9Rd
vyhHjZE/85fu4QBbvA3XTWYpeb5vHYJCnorE0ppDcVaWCEe4uBXS7McSW7qN5cS5
L5epAqXn00rJu3clycYns0xd/9DmoDksbH6ygLDg77kDxSuO1oC18j8GltSQxi7M
92FBW0kfm2F3YBtMoD8vY76rs8YsgOnNFYzE8seumGM08q9fkcn7xNasLmw9oHkK
Fqpf4ai5mUGQbpKi1y14m81L672Vf5SZ2Rf1RK2Pr4U9dCFLGOgoVxw7o8tIm00c
GY41NwTl3YMEy59mJnGJ0lC1MiOEVzwarDa9zwprKXayaSfTJqY1fk7ggDO04k5l
NlsOaE4x6coGBJIg+rlrMn8PFNdrdlIZAFPLlyQjSwGHD9YZANO705nOQ0ilHVyI
tatW5K1yCtZxyQGa0amLvSuPaJlhX3tKuaIpu9dE1BelVMr9FvsEfH0sP850dj9x
mT5zt9s2M5gS1EruEC7nsqALOXyoGNiEs7KotWa1uZnabLUcJuRFLpyeT3XyMpNl
z7mq1MXmhoJE6TSGAinxHE/Uo6LoxMvThat2MQdHQ8jyb1LGKWPiEOR7JgiQvmKx
49yBYMfl7osLKgBsTA4m8bDTEuQTrJElYWn6Qj1tmEEGVWtFSbgcttY1k9rO8Onw
sSkVMRiyz0MZJ6w2ADhdPr/PBolT1ICtkLq6xXbx20RmKI2+JeVUPMTuhfY2B4g3
nJrJzSw6e1cA9enT1FTpBDSk80tqvCDk4J0FPh+olRFSCal1pKOdjg1HPHnoJYK3
bi4acUHgh5Ym7J+FvtUmIQhd4I9QVS21XVEIjer7ol6pPGDltRbh8PWWN2ge0X55
lqDUacQJbEiJgvmL7sSbKw7M4t+jYY7AwE9y+Y50pVOksNjDHmLR7dMlMv+3Ujqo
Jj2tEnsDGfmRSW7bpjRN/NA/GqAK4GvmokE+yblVXk8DJBmDVrr3yA2AVl2L5/Yb
G5OgS7A4yijy5FztjrqucRCNHCQhNLQ10uvVqhjrJ/CZuligujsLl8hV6HlAFRgq
K7DN1BUdkBl3utAUcWHWtmmRZ0sB6ESmagX1+au2YjOGfgMZZHQu5Folhmfwc/o1
RusMPztuikYCS/b6jbLkEGnobRePXYO8892ol6lVO/lyAeKdLZDaiA3UfuYKNyJb
5UBZzrHiHtDIIU355ShxwGibEauRhXVa56r0jBftIjnyWQxACnBIwtqIVWD8wjX+
iq6gJan2qoq48fqOtv5pKeNpRbQB8OMUtUFK9EPvi6JtPVZxCQjpBTw2t7LXldhb
ZQP+T5RDvOVDPe5f/yY3JqWB581/+3WRCgYca7PWzEkNuUHsby+OIWIv/lcGYzA9
wl5SVzd5JkgUF49fx+t7gtAqh3YNf3QqFBleGCEZxQL29jK70z+SgDftLJtM2nmw
FH01LeY/OYbo26/Od+uL+5AkgQkFnLd82jP4rJxbREOCNzqmmOGNy1jjU2dwRcep
WvidxACVJUtbeTOihxqeHg7cWOCYJuByC73jY2N4Zrr3GJx6sPMDbkG8O6lzoPa8
KI+XEEWnCkJSnllgXj+fX1fECLn+lp48AfryRq6gYJ2rrYWoht7bXGX+qcGvecBr
1jz8tmGbadR36RsBL4RbfB+mgQFO+SNKS8cCKGTmDRywzQFljZkwnyrmKWdA/8AW
Sw+I6fXEL5OJOUw/Z+rDHNyuLLTNOJoFqOtNjmERsBEiqggrzBJHpwQdHCmIW7R1
BjuW0xCkOAxDT+DoOyDLonkeLGXNbrWHYWODIK2HIizGKEQ47e2WDJWzFNu3PZee
0md376zV1axJR5pSdbIp4tmXO8dtCvnQjEA0owQ3Gbq3ZREtuTfKaO7yYJnCJrxg
6uuHcAAiq5Y/HtACJdORXdzBl7bJwSe2yWoEJ0HoRxJER2aiojGGug5yiC8LkgMP
IFXCeLI2fFce39VS/GLc+Jb0lP8U0APqNmo0GCeuC+AMNyh9EGyGOdjg7qIw2IBk
KBaajWTka2We9htMqqJj2I1EETC5pxaj9D8ib9r7KsJw4U8z4aa1LDHgPyv2WBHH
Ntl8fvmFjWV4MF2phGBm+293+Pbz0lhh4mROe5FNz1ttZmpkd16A23IrQvYzXxDY
g476muBEvpv0hNo8evVH/4MIri/YqhR9ug8PoIshevqt5CtqtjawOSSCb8SqZdmA
Hvi4LzYY26fOj7nen5t5ZvwO2LgR3k07nzWVbxpYR4ohFZgjH5t3iBgCJN4n4/m/
6Xtd7VSmqdeHT74l0Mw8DEerszmbwu80Owz0+qwroripfcovx3JhbyYCHOCH8vBS
KaGdxSYslsQ5MYROVKc9GZTfqCuRA7SqWfUrOFVt4Ma/afHfsovC3jGmVjSDiP1/
7CZb3RdjsdrTYXda59C635uKs30QGaYG3/ww9sHXWzLCDsJBzfigtkzI8OHTJwVw
LLk6ba3DF/+0qFooiu42x/3LpHBapD5W2p7aVWOVzRCXqw6GPMTjrHfmUCnueJTM
Uq8wkwwjUsc0Se/vIAaUxCs6P6uOKsf4Ukdf4JoelKAJiRt4iFcSlJQFoTij+bAj
fktUUSmzOI5YGCdXRnWpgmlNVRCYInpVpkGhAOqZtaGZB5xzBInd+uyy8eZtXF3b
/RUdZbav0nqgb0WDTzLljk7QZWPbOkqLAoblhW+XZMcz+MaJaS0wXQwRxSP8BMNL
iFZM2d3woAacjmHcqRBMt/B4xCESmwA8f+E8e578KpAMDSpQDiB+6DYUkHcrY9b0
GYMdXL5a9wVqVPS27770tKVerrJf0SI63vq4y7VCqJBDJAB5MKQAGNQ0RzLDwJjE
UemDJN6a28PNTfm+R3TPHz+ILKlvlf9B9pRMY8HiwO/rAet8NN25ZhTLPfuz+wqt
PH2z4dHcGJF0k4qwJENYoLlXuLIKmBsPm6dUF9ZSg6v7iT6F2Ucvy9ZU/ESF/OkK
Qd8hGA8YdaEpPCx/z1rcGLSLN1758q6pvi96Qmus9EUz1qcC3Cji1T7ByQ9xDHT0
aBeHokxFji77Z4BSNM7zwKrD7p/4hVqage0qdkedWA5NGIR48dFYw6ZYzVRYfkMV
sNNBptV6FUpHFhgsbdDm1BNqwtjlLDv8c9pbNbv9praYNFI0/LGxXwWo236YwkyU
EKeCSK8Fu5NBuDTzaaecEfA81fAkHs+yGouhQxxnZkJp7clUtc+WvlnNCzXlenXc
/AGiZn9QcWY/Vm3SYKuNt4zJns0gtG1DvkkeN/jrizOelI5w1DGkWFw8zoE7sv7I
HA4j/F9XpYhmOCdMK+/PvEGCrt/cIM4TDtN4Ad/XetP7f0fF0O7w0/3kOULuaxIX
/qUD9+KFJm86536KJzVNm6pS8sMwH4WsElitTYHolNHSgXVRE+oHGVOwCuTlJGz0
8As6tCO6dne7yzjXs+iYMBe7gfPUgSNuHXmDlBQQbXc1qAX72EeQaB6ZYM7ZYXgX
RmjnFQd0f5bYoHYHrLQgtf2C3N3gvlfEYFVvCvvQX1pKo/r1T4uyPVaabDL6Ae4g
dn1KirdF/A0ZwaB6hGZtn98pSZ8jSu1gZRqs7x9BoTDcX52Aa85W2Aw9VwQ2EEZH
OKx0ekW5GEZzVgEFiFA5s3VvlAL9sd9Eqn791qEJ3F/a3kFEd9hFd8VRw77dJbTA
e8dw772ay0jKJbLUdpoc3u0ElaqL8A7aVluma8l1Y/YhVJaxXOej56LByJ9DqbpJ
ct/4Xm6CpAviBefmakiZFBuM9axxixH1IUARtBYuzo8Hzu/u3xclMEQwsWO1VxTF
7Stl6DT60iLm29F2D6fsiD97PmCw6d3fzWBxQp8VGoa6j9K3yG+t62pAjzvm2VWk
XNTzq8q3Sj0+7XEWdAhf5PWOh3Y1CIZhDRgL+ATi+CSbpHpAAF+ZoMqNMit/VocX
yZALtlMRVsxwvO+AAL5/OB3xQz7hDJDCWFMbgI9kjf7Xp8vsAWcVodEagc4g3tny
dcuj3dH7l9G1FiaMTmh6CrUXOaZfBwU3wAEsF6NnqttXvifV3rSNFdL/d6iG7kZ0
t/dNuypLcvzz53m7T7nXv5SiZzRGdydFqEvbLd1g04Nk3CDgkZIeObb9RYm3cyYJ
MhkqdT13rJwqyDpifCbUuRdry3hnS98tcNuE4w8GpldO8kUzdz+KFks+jdaDMHjE
F9zVAI/aJawxX3Y7P1prOtuLmUsd2bI+IHfbfEY7d2SNEd+DCSYdDRcdlGpoloNc
XWUQ6/YsAMeMjct0x6UjR5jgDYNUhHeKpILmZG06t0x+EtC57uXqNYb6m8S2kmc8
zrUGrlpgvkrfR1ElT37DRHY/QPAb/Eq0E3t3Jh8TjnFCIxyZGSACq7zHShfMaxDR
v8Lm/JBUv5npz3Ssq8CpOfbf2mJ6l9jC/HvU4GxMc1LGEUbziwz7uZw/+sVViKGw
XpicuKUUORT7DN7mhVKFUs6bQJpGrErlKYtP10If02Ft13nTNQzWWhYk4US+EyVU
KHmRLfFr3GMspGqPClblE9ymQgd6dWg42+V6QxlIySk4W1VP5QgYwBG+f5ArT3DQ
v4iy7H/pgxXbwD5Xush/QCuSycG2ggPFVDNWJXwDx26lTRXfuItTO+EXhtt08a0B
jAGhXoZkyfON5ORvFgLoba01lqdf7jY2rNXBId9oFwR9uWcRSrAcysRnYZdcPNW9
6qCoWliQQ54pwA9eaDgTFeEncqQbKVx00hsRzbQuzvxlLyfQ+lmMZyOGCTnWkZ8q
lSVhhzzc4RV8BE0sHz3ziQ==
`protect END_PROTECTED
