`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1l3liqmboIAw71mjK4RONBjpyH7lF8XgpqdcS9gr9y4J7Dpwf/SnYzddAmeQbwee
Kcucvdls8GycRemfjW70U0OpUnDBOJlkciKSt0OJk7CiVHuvyZGoHhRsG7wdPFxC
qqMh2Jl4UhqCEE8BHc1o3SzQgEvcoaggbpa6wqPx8pyum++yHtR/MFL6CdU438P9
yDNTA25iwDEtoTvLb6jSspl+TtivuvxK5IQxvjTt8fVAQ1djsdvkpGgg96sVC9uK
GoUjejKMNAgjAWcAR7BvW7EQwcnLZ8R5l86iGVGKm8sBS6EeXIB3G4XtnsKgxmiB
rLRMthLOje212RF7pW0Hy/FOyG3U5TCTAj+mwFNpDvSd9L+tEr0TKuMUNpP0WTRj
yIzC3WFBHeJ6Em589O+qEzkRHkqlfu43uJ0imHeRvSJvZlQNH/Wfp1A411lQbp/u
Am+Yh6snscJGc8wjJ2vVGMglqzGlbwVuAUWREa58PxbekFX1x7mUazq8VExs/Ppq
Y5eqvlmPFFNSyrtdZmieG4gqulCv+zRzd+DAE9P6kEoYtOWo4sGa/+3hNIj8wkyP
n6ArCqVMA1DfeF+fU3frJNNYtZvZGBBc9WlojYDTa8k+wM3qho2JYqGmeCnYntze
pEUbaPsuZ5l9ujCswnohtC9BW62yGsuq56z0nsh3RPxFaHDupJIlVbwLSClLn4Bc
+nz01dc7iTmJgSDA3wtR9LuB8KIXlLneFa8rBtQ0foAjzGWzd9V6fRZEP5pYhzf1
/gimNkRWOnOfr8sCiN9hjTDCNrpGkN7dhKxQ4/h0nUDwBrGhjj26ofoey/wpkiSl
GfqVVoo4yvLmp+BMSAuLFiuG1J5b+GyJsAgh644xC9br++uJ5vHi4WmObzwXWeP5
x0Vsh1FOnumlaiJOrvHfOcjCE3A2KMunGBeSbYrTnfNx5OJzrjO8VIw6R+DVDQZe
P/1g8triTrEljLoE+JRVjb9lj52eDxseu15UQYu+xtJIZVSC1F+aIGNCVlYfommg
qiZAoKYws54xCfAcsMHUsBkcWKMXbRu7BzAwTdbAY5st6K4UlWXuailyVhxeRwS9
`protect END_PROTECTED
