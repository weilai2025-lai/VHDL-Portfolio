`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWH3Y2qCEUxDbVkSi6VNc2l50Edx05+U9cyVB3hckZz2xebMEE6n7Xf3+RzyJkKK
f7/ou/9MWUQMEk3C46EkpqN1Vc0iqkt2EUi+osMwF4hJhl2G5J4i6zUnXWjn4+47
Mks+YjsMrhzuOFm5bjb2zbqyAxbu8SZcpvcXslrr6+aA4jen0ajW3g80e25vUt4D
W7WU2PdFDTq9UjTOs6/p2V0Pi8MU86CtSKRamD22MMobXIP+0OiYtJY4ZJ9TO14a
LmNvD5174NkWGqt4Y3GQiezOmUrspv+CyX829qFyGHdNpK7pQ3ElxLTaZzBqXiun
iMvO3jHOL/8nNyjOzPI4iT/oqxjXI71FJ4gfkWZyJ2rtqO6zr+dQG19hNWHpiY+I
vxijlLvr8cXtWCLEM5NCxctTa3J9d4jDyU3mxQdpqzbumafvzWFmQgJDGipPzSuS
qFdeffOaaTFmzM7A/DspC3Ow+UrRDFG6dNM01wLe2lG3IbMoPKoH8NLXhYZ0NkxT
YALBhKEBqYr984HhUjyJRzqtQtsnWKqjyaCrzJghvtX6wZzFaV0/uG6P3ZArbSYU
EDny5sHs2KAeczxtobDWjOBPrApHT5QOKTwgQP/a0XVS105tTxOfUvIPZ09nKR7c
RlPuqg6KijDYtoIkWTBwq7uB1RVfFV8YskrFxUbRVz/yuFunysBiXOjBq07ILH52
uzRs8oG6gA/l5peJ3KB2TI2iJqXF04EY075/w0EbjMZd4xR9spr5JCRGYpmje9NF
w/6G9o3fv+RFA3Ia9tHLj7boLlAqMjZO4Tyzoe/OfBZhNzYnJZkSOOi/iKRu8WYU
R5yfFgHBFnlQ2QDqP00NW40Amiq3oJXV8MlwdNOcfnUbUlFBzJX8GIkiecMZKdbq
n+kzapXsp7go03lIF7eWi0ydhM8BV1omb7x0aKrJ4IE4NhhvPFR0+0UASDFGQnua
WOv+avl8WHS3tst4kZFc2WQkBs9S7M28PL7+qWHJBRsVZoFxHjFk0Wv/p2SzPAut
/x2B+uZnOzH0XQ0UmSDUWfIjPFX3Hyx7Mz3WbkdMtT3KWZNpAuNyavESBBydamGd
9LtZeeUwNxaB9n7Tr93aHme2edNU0A21RGovo1H1kbGtsB/Wli2svcB/JBs1mmaq
vErdLPL6lnILn+JZPS2/GiA0plP8c/rS9lG5K3JCuh2FVzV6+jA1sMRdyGpBMxx9
0H4BhFo9PlUrSYgDEMynOHNdKueyo9B2kb97wNWPofCHLZ6HchmVPTJ7VsPj+uzg
VS9dxmpKRFgAF0Z/DkyL8QpoH5KE9bwY10yBQQ2EViK6aKuM7DaxCdruDGACoCA7
zeTPRiwa/dhrsjKZBkjCAihd0ArHHUbB2920mZFMN29n1Bc4lZ7qLJ82cY2+8mea
Z9MZFEGInsKZlGdnGlIqj0+ZDOA6d9nxgcDdONsMMuu1vb4f4Oddvde/oG+0gzjo
nJHw97BaZK5L2BKj3zHwvrHum8cPmBbUYXrwVGr16/cqTD2y6ifamwhC8pbmZY8e
xPHqDNEiAy3IGiLJr7DfGJm9O4a4si7Fs5pKLeOdHFr0We0f72ZLvWohoKbOYzy7
UxvNHhYXJpCrsU1r+mP0uSm7TZeyfGiEtGc6VkSjE6t2NouHs1qAPGgyk3fzyLUU
CHUdirV64TQAH421/3cOWxNdCW2vneKojL0H4YroDN5bse9LL/0jNaXsj0CDyPaS
Xd+Z5IEbGLwjPCdQBimVBwf+B5N7MzYN2ncD/+c3Xz3uBTB+IluVljNktYu4DPOu
yb9LLfeiHk+l1kyJlpBlvh/ap0z6uvHsmzPI5xaAPSwZNoYAzUsZynrDRP76Udqa
ams5vZsVa7CUUFDeXwVWRS84TNG3DeAv8l2jChlF+gayWjpX2OzGS56/juKYCr9L
EAfMW8/nk51zn0mxhBxX5eHTg5rl0NLtfsNRUWlu2+St0HsEO5WAcmnTopsunC9g
g+gxIJvjHef5tO2yMVo9VcNQapQQyJbIJx06soaYyC2PMaAtRMUlvyOangSNIWEd
cCuD3hCZy6IwBQXjXoWnvcBKn1rceKZtBUEdehMGcvmC+0ZEyNiBCkLNSxrhEyo+
imFX8+zLqhBBvG42Iu8PgqRt08y2Ynin6Ns/vz89hELciTjBfO8N00ZH7bDoPIPe
Xx3qwVCXPCH1DpWzbpF2A6WCLU1Ac8u050r2Fdhb8nZ/PVTBlDkSGMr0QkU+prPA
37q1mRlnUuwhdLcbCTyQiLcyEBqHpSTe9jYMT7OF/ibjR3CFUO///4I09gJsaT7u
9gQ+8cZ3CEjfL3En9YIahGgfEvDrQVyrpPFZSe8i1sjdd7w5fIQ3ipH6sH1H9G2z
ppFIcLNnCRAqHS8q1h0d0NJJq1UWTSF2z9ofijzctMahdthe0IN2eNPIY80H8biL
msEedjqsNxcBOxDe0QaRStvElp+ZesfH+3oYly5j3d1M4AXTtkpQAQXENvySFif6
nYE7CjTfgFoQL5/GfdT2pryRW2sfb1ONyXndxmh3qiv0lrPJOd2CXlO1HoXtjXUO
yaNTbZs5U2yucLuSTMvd9AgkqhK+eAIEsA2cXTwNYtUxxkWA0dU28zkp9rWOZyGX
U4v2iMDzJmgI0RuBd79BybhLFBFpdgMGqK/9a4kuHXdDKpQY1mvkdtEHfqtu48e0
5TpnipvApMYZWMukXM842fs3ANSKj0RkD8UAJiUrhQf+55HtI2LZncEFbRW0+pzM
fi5xX+JIuO8/Q1aKoHdphZiPiPKe+3CsKGpukA6OBUcmjQswGwMQdwkdtneJdR4w
LBulwn5fsoxWp4l5dSZZKzZnDV2IdemfRQG8kmolIeiHIysYSSrjkrCOR0RygBD5
vKxVFLEjl1YMqa4f859LOn3eARaFjQidunBUaWpOoILTF/kpPkFCRTmcZ7Ko0xHH
333igOr6ckch8kuRZ6eSj6faQeaDZrjkwoBn2nTEwBkEwgoPnBk0eiFSXIaraQh9
FcJm9axPafN4cmQ55OkwnbIMMBII2YwRj7x3fw1OckGewA7ig4bG3Mm9Jpnl1VLP
Lx0IuGqOvrVsK0r4Y/lLMWKHOTeWWApD3vNhCySKiQLPg9WvuxE8WPXqTjzbwHH4
qo4rRcaZK0CJZDH3bzVrvCE984eIzJA3W04oq15QUarKKCEAhURejjKigLf9AaFk
LZhJNxASTPbufcqPo1UDnSGkwFlfjpLrP/2z1aZ6qVe/K2ktrE4QB8/LUti0COiG
Eu+YDQQjl2TXn9pEqvPxt+VA+UNiSRDK6aiql38OzfPxRYo2znY85/VVoNq73Bac
9EEy9dk9jVHZXdQg/RHHYJp8hXo3DUqC6zTV/0A1hNuCedwVAIP3yw/qHwFUv5HP
/rdeIpR10mNiA6LcnmujmtIy1ntAhesyt+MYQ0Y8+oBYfuNfdAjFls+Gzmg6D2tE
9B7xXEP2N+3jPAR0ffvwax6JADB1cauYShXCXBUv/UqWo0MtrXSJ7KUvf7riPtYt
Zx9lW4IpDauyrk1vgpvi4TPBGWKO1wKA2C6RAj5D3ypN7w5ZI+DqTVNDidhOIAH9
OoKUQmZ93uunNEIIrfvkRtNRtT2PH1hnTu2LW05MqgyWVZdIyz/BJ+cOZhkQgq07
EIuOB5grv8Z0RD9xZG12i0nBA9Q1FGle2QdpQIzzRG6nGOpQeAV239uRsYNEEfrq
pj2k7vhIBeedDJ0Yq78houviPzuWe4drqQ8ZMaFvEZT8T+eEfr6Tk0s0tpatYsBX
Z0pAdd49PpDWeCJdHlcOxAfBZqfGnEp7l/VZZxYQmWJ0UJ8qPSp/VwQjCwYhmwWJ
O6jOELH2zwF4115j0Q8VVwRp82pnTnFZkuMBaOWpcwOh5DrPgkkyUJGG3YWBrv2o
YCuH62hxBTtjd7iUj7iOzLQI8qZVlfqz+4zILrvqyUSGQHEytB0zrcOTWKwXbXd2
`protect END_PROTECTED
