`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAxW9JTMzDUokVajfKiIVkhXn0ixNvg3XXkQQvgER4UmL2/GnAC+lmue8JqvILnX
nfrc3wggFJQubvaSxz0QRFjOd4OwDeg6HqWXR/zvufAuQk9hLdhi0l9KlDifY42h
bPjwPoCMpRTBHI8aQnllKo5dhwKfSH5Hikid9TMZqi4zoJJ/mxZF+yY6fM5AcD55
NpsXp91R8gijJwg0deeOu6o9BuWfKGTwo578GU+6SpSFr4TahZz84yt0qhYzS+Ti
DoKvLEgFyAAN6K3GqQ4mJTeM0ZSAI1ZWgaARLb1nGX2FSNgj/ftNccyFaX3lDcXN
vyxyv8zMFXu3+wT5ZWQhhTnsKqawLY7d/Iof9CAuutz4eKX26YqcwQQxS2aHAmUu
UvcvPdWWK1DFH16OhBoBpOyIL76PpqIrGomLzJCHByn+9mRNXKjKwonIFfiHTKYR
ihljLtSPTDYUOYRqMjFHE/wk3+IsY4XZ4Ai00ApxCm0Ta+rlxwAfLNYLp406cKvF
Zyx3BnLCAXv7TTMQ7PlIO4xOZfB7aSm2DB70diRvvCLa4NgL3sdh1hos1G3aGCfg
Gvbk4V2XuS7w20sna8bsabxhVFR7o9vnrKvaIN30T1IJSQpO9Ate+qOUb7CCjZIl
dMJBcxSgYS8y/KjaPOU29ntd1P2Bto5gb8vwJOyfvBZLWh9Zts/w7jaTtE+wSnc2
ybpgwcxdyyqAmXdJh43r55AfqRkJGy2e5UaihAlEOn0aWLWasEG5RW8K6yIo1BWG
lexJrUPs9Y2nKRca1mg8TXCB7E2c7CBNekNlGgRx6INj+Qmo1ayVm3nAgoxKlU+r
yvUoQD6lvbnYoncTQWm5LdBi7UJ6yTXGAw6d5DqYR7JUGMsEA7O/SKZuaesBbQOY
XHF4nusCVCKS0iHZ7Sh12rx/QnnCtVjtZLpDK0Mj1K1UEHV5E/hji69kQBEuL57p
C3+Jldlpag7XhHxcL4+yx/4nKvI/BbXXzKvra6g2hzbxI4FjI6ZiaBNCuoWnboRu
qs2DyP6DFpbV52AhXlbGNUa3zYXW1/PFOzkCXH6grRD0s6mUQli9YnDpCAccmN/M
a4YnvNkSIwI1VvIXl7jzTKYRGojbp1Tma2zqh7Ry0ZsD/u8kaAiEgQFhR9gMY/lN
l2lJvq9IFOivn/Mm9M4oh3GDC/SQwZdqRDo05v4uugcN7tZHosSgEmfTSLbtUo6D
kmSbYh0QQ4UqtaMC3MyodmksdhQHVOnLg/F00pWHlOy3T2+QdNuLuKRpkK8WJKkj
+Ane+holTbmlY6eP3f2YTNaRtBu2orJ37Ee+7OtRRxFakwFE3a9jBYYRCf96la1K
VBl+PWZUBTTcpvO0MtLZ4Joa5LEtsXWD4kqrjC6y2qA6Bg8qoa0zBhJYs1OSJrji
gteBeIdeSHEqAbKHUg9umvMmGMW0IpJQqxEDigsf0woWGl9PPFNd8NRwc1+65uI0
BepWhin8reWDstAgRVR7FCDvzzfgG7dt1UGfUaLCIKKQSkeMFBCC9gR67zJ5mpw9
8h0tV09gVqTE8pgjooWXP3hjnHl0SbyAdCQ1XB3JImecjzo/2e8qTzHSV01UN+y5
4hNV+7RGxiQnrR4/JT7Z3mmvtGBOKg2BmfQ83l2MvFk3Crm6tnbLGG4k4fMDTusy
atRFkqsmLoERiRJHS/JxxJRF+euTvC6Rp0AeMy4gb8drYkAvEwF50sy/Y2mz40Ob
i5RoU8WF6hHBkyG/1VZKm1/JjTBXO0ceAmvqNtOT+AKEsCbuXeHGlOeQ3oC6ZHo7
EJlj1hMdwSVctvqxloEpApHFuwd0bABIBcvTZNc/JEciypwaEgu/m9E/+bXlPssp
yzFCaOpjJR+TIpJ27phRT0g4FfKWlrvlQM5V/d7a6KmvWLNCdI1asmZbw96eA6wq
AnPaZrCMCLdN7Cu14iFC+ki3COy1YHWbNd/h1ReULcMmYMkQ0CHOItbXonLVOHm7
NB0xvpHMIv17wYpTSNUkb6VlW5vT4sN3PGztgQjHUgeNVY5jl9WHR3kIgzmiPFj+
5slxE5NIwgnvIpg3TNyFcayjXSh0NiBdejgz8c9f6ovstD5hs/c+ZLA9/Yg5nASQ
eWUKyGGNu58uZYQ3S/OSggQtBFwuuj241Oc8od7iq3oTZDsvfu42a2txDE4hy71u
/du4cjwsMqEIXwnsFmkOgchV7VaqR0Kd5nj1izCW61fPvOrp7jwv0RXyHILZgyUQ
sy8MIQQ4u7p6CpPh1ekvbyf7L439w2zbX2x8wxD3IBeFn33YvLDNtLMTacaxsPPH
OPKVY1LsmApRADKu6YBE1857LATI9DeFA9SyqR9jgzLQDduVWm3CLsJ3naLTEjou
CZwMmyi3CUbtgq1gwqcD/fTVc5GDkMg0Jo3nldI/E12P+QnZ/F6RahpCMVxOg292
bFYAwn5b+JHJsIV0TgspHZU5G7PpNQGi43Oa9lkQ01pe38GUqUF06/dxYif/8LW/
DKXwCEPMt7RJ+3Vey+x7j+BDSR/c88v8CYup1+uUNfyahHL4XwwAWmpco8I+vuT3
DqMmesUkIo0yNocmjdCORPL35s1kyt82nAKhDGUlW87TPVA7bIKKKOJJjmjAJSpF
4CWPYtOwoFlY46ryvD5R7E+XL94popQfDqJ/U5G6EyGd6SClFec6Y/9KEjTLQugp
2+qSD0+h+0rm6xQqL8NNIgohwzIW4UwyRT40zWpgbn9kIqhEaxMXJlig+CFbrX9k
pu38uk8+idiMqhWggdXD+DKakD7aihinVcqgj55rw7LvWjcHMu2yKIaa3MzkOWeD
ixr7KMu7m4iN0sxrwBkLhcR9sAC/DvSXMEhsAi6ut5SAobF4BEhLZqdpzHeDHIUa
1FsjzPJseu7xeAJAK1QgULpOSGAZP8dntKd7AvgvFfxtkm+++qKHOyKyKkxW5lsS
+WhHMwuizE6pg+9J8E6nxMu3qkS8rcvp6prWLvVb9W5OQ7s7KyTXg01MvvnvoCMi
cMleuB67w9g0h2rQ2U1Ab61ZsOPLgTqkcDMo3ZlWF+LwPcUrdeN2mtqCGClj5otO
SMCvqQYBRD8x9Xd8O3Y9Fu8eCHsgSWMTgS7zZz+pBmXtUKdLa50/PoCUGH210HI1
HDL0uyY/duxZxr0rFPVQLSR4WqO2rXNhmL1yvO146yPDNUL4th79A36Tbk8p/0OR
6KH4v/nAsaU64NQb8lqkEBNjuL9CUht3ub8OoaT398Gha7w4ozK0lPQGhzfE6Oj8
F1eUnCDXIIlbRb3K0VSujeGFOqvsb3eBAnW0erx1D7MQ2lmwN/Qe12KH0wPztSrq
ecP/7lkzWgXFKVrJP4AEgR1OQv3Ny0T6vVt2KqIszFSgUZ98Zsj05VKuWLI4vjfv
/I8p9Z9kNnP9TMFup52IufB3AGGxK/gLHykDdH4ViL8rr5E4vwwpP+de7X6BBBPz
791f0ro3C6AoziXoMdgwGzMIzmSvVTy5QqeqKrU+KpMJ0pdgaol5/GIpBvDNAj4L
SOD4BZO6hBiOBk0bvMQuW6S0aa30tOxAs7rl49tlwsLEb/cKn3Wp6n+YZDsSOUKb
5OmWItPRK2DWQtFftSyWd+H0Kjz+RMoV9IiH7h8wqaHSt5Ls+b/pLPJj/ZJTonEK
oGRf0bNofjC62CFqD8g5FcXBGVCC4kOOnsPdzwB1A5WbO9cRfkrTFlATepOGXHHp
EMf143wxn3JRP7VoxV2XiQFaG7RQ/F9Pe3NBKve8f7KZxvnHAWAKXKA2g5mZhMeF
GJCyll+x9Ln7B3wPT9PGYQFPetTnY+qe3Z8NtMPfpVKu6RYYrgI0utO3l524I3CD
VLy6Ufsjf2VQe9T7TfZq22aq+NKD3RSkq6iY9V9sUC6rxcXN59W8cdnpj+wEx1w8
9UxCf8TTwhksASI/TMK/kqs1bytby/fDmSQx4HK1cV6Q2vy4H61p3sY6U3ong+Jm
cwC+Tms3cAylqpuznt/Hv1C7fZo4pRjZ6L6+mAziyk2QEaxShT6K1gLO1zuT5+ui
QyHOVp3BPEy49Vuny4Rzl5p/hHC81Ikn2YapobR0hYSX8tFWjImmv5dgZWbbomaK
zvar/tXrY6NcROX/5FGAS+SdddKWuTanUVSMp6drMq03p2TJuKDiJpkIkGsJ8T2e
A6xy/50oRyKBVo6JJVuZELevkdoAoA1Dp+LvZ7+K3Aj620FzDe3r8JK/v7K/Id+h
oNOaTmK7tY+unRJQVdqzPl9kczfsNpxiML4gje5tkYnwrsrptQbZFWcHhnR4YDWv
Yv8e8vBD1LdnJVAjD0Sz4a4aoNIcCBv3OtKCnaxqGYfDAHKtRrQZ0AOyuXmbQPJD
WWFrzN/dCGlstLUGUSm9LhkUfbqJ9NgiuR6uwVEjl8FwR94MFtMc8dlgstwtQJUo
p49kQiY4EGPHblpfLkItNUryV552nG/891y3h0WE3zzW21vVBcMdco7DnpFqLHev
DqbICALBo/bPPU5rarBJjUuzBqjS5mBtydCKtHpdFlk3sRPgSxvSdRfClFV3V4Om
D82EQ0N4WyMQME4IBDOvDIEqGtWzol4rT3XR/RL+fvKPYAS3Eh6yl4Q5nhNG4MpQ
Ynq6tXHkHouY3u7GV49VZLeVK01xx8Du7WIWOVETxFhBr2AtQufANQhwjeDojofy
7syVq2NgXjRy7eXomA+ZFi/PqOr9EIIDzHwGiZ3/H/x7N2jqGHUjTBiSBFK1Mjrx
H64b1y0icfH/YWmJRNP0fH+0Sesi96F01MxJyD6JdcVEotkb18levLr/yriXwcgM
4UO56Q5Nw2o3mwC7mb2YFmdEH81ITwgMLfAGGJU9mfnqOn3A+biZMjDEbB9CsnyU
iT7NKFJCBtB+PCfc8eSckH4SObQmEN+qIxAD7u/CrMWZF/mNvF4Xb2npIUZsil4L
ayJ3lZw5DsAwbEwPEsB41ACdpUQgSt8U0hv345BxPPRbgJi2pxm3nfGJ5Ve9xv3X
Fm7ZvMYa8HPjNpqHEG0e2GXcoqIFQdABlJGDXylZIWAOwPTey3NPmjSsQS/P/mKt
V8np2EZCboLLQZyoyvwwjAjyly+G8GsryrmtKVtr9ibALXlDXgphpYV5RUD2oOLi
y+pez+Ka5L1HjUoLZr0Hblj3Ny4dnyIPenrRt0jmIsmJpkxeqI/9SlnpBtiftWCP
UtexXjfqM3sIDmIVQaH4wHyK4SGGR2PKuB1ySov0R6J7kcPYU4f1udUfm6npKnSJ
b2ud68zOnan4k+rLThdrL69Is8daZoE+uUNflbsg+K+W+K19FegnuLN09WXX4OZt
Q2NfGl6bVhdMKdMBHmMSTcN/P6pcbzA4nixYXmECM6s05xn25q/wb16tC9rI4xYp
yzXU3Ny9Q/LWbpFYc1F5L9aT9OCu9ICcmLbFsz5fTY/OXtDF1kNBIbmNf2ZTzsCp
KKuRB7Bhf6asMhs0SBzKB0sAsVgbcfqdIeRqLqnB01KshF8zjOGDlCb4ZX3jlzk2
1tQaiSHenyZ/fzdvRQXA5gsV/ZIohAQqEu24ARpS2L2HqLhYLCFa0Wtiramew2fK
PYowmZfKLVsPVCv7RkuitDfiAWlN01SopDs3Q+2n+mgWk72r0egXnV2ahwMcvGx8
Mf/w1PI3w8V5lsDxL+SL+6tB6yxxXXOSOA/jCdfvyfZZAjqUrr0kyuFqLaiIw2qI
whdthVdeAUe6/AmqQkARESFzLaZBzJyPFUzayv4g4KL7N/qHW+xOjHBlSI18J/mD
JeDg8GmzlYhDNt5imDOUekTfbs4/8E/OLSKKlkKh9uc=
`protect END_PROTECTED
