`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U80S5Clrc26AdWt6/BFpejsu/pheyH7HRe2aWzF1lET081O+Wb2VruzrQ1CeYkcw
6zAhIgjr4deDfmqmy6yV8c+F9oohSrVTrKPVJxtp7gjOCYDk37t9+GDgWhmsF3tD
ZtTOZxayLuc07hyT2L+8c2l9ysm0NgQfwIli/b1ciove6sL6yIdz9dQJggrIje9e
AJB6Q4G29QrRvqG5o8xEYijH75F4Clmk+JfgzAos/kTzzV0uQNbZDBD0RvsexRL1
y4+1Q9XPkPj2yrEeHI22aJZnSjMXW4vASccbG3rz/U6BKkFklgul+9Ge4RS2xDu6
oIR0h3nBK4QYR8WI3sVt5fW+PtjdDj3PoqqBq+ZvaymJr0hLgAJaIKAh/z3A+GLH
Oyoiaf++Qv7GqrpJ9SkIcpnQ48UTaWMoNwqU5alOn9B1eKGcaxSy+8Wtyxw4bnLW
mSldBssqgM+i9VCXdT0fVQSF6kJD3n0ZRzmkbERjydI9ExNj8gBgLoQ+T/gKsi99
vcEX+avTgoE8+Oatvnp5FlbCV8fwB6l8uAkDrw1Y30LW+v+OIILLBDkfduAHtjdP
It0Wzs2/uo6+58ufUNGTHQndbOp4Js/sIPL5kmIyxH8feu2ucaPa1GeiMgVlpeP6
euacCzYVnNlUn2HsTN5KJcA/PrW/S5Shz+ENs2wJEuXSHUN5sy2rXAMikh14oOBk
+P7yNjVVyPB1GbwYZEI4YjZ0whdfvUlf+FAoIz/OBIbxx0fNNR5ve4iOyHtSh0Fw
8/EdYFRTgdbVSdfR25BXSRbMuJJVP8K4TevZVPxcZvSeY8Lg7hZB+rFd7XY9Qu4v
OYPZwGn2XTzp2/XuIjLtGlhadiY2ejrd8LqScF7kqFQ9vcI4WhENpHWZDqm318pk
VJf8LrV7FCoXQRZPMrTo5WzS5QX0z/yghMgdkEf5jKWohZsOpPDm1rua2VjqkGNW
ieyG63X+iKWyiK/+01/gLjVOTpr8ZEMfp5QwUfePRNMnSmBkiQc+dLzzH651m93z
0/6j4UqVonUAXEuAtZ26cOwpAhVZvUUR+pg/MItLbVQVkR+IKz9fDs2li3uUNYsf
LPSteBxUyTVtzHiBlTyF5UkgP2fk9+Ou09AcGM0H/UzC3w5jUFHOSKkfuH6/PBIn
lnfNDTPaucfcSbLSkOs5075n16yInhsg5oiLJRx/U3x8aRUR4/KR3Om1hGdy7wE8
S66W1UQ/Ua7k97NdsXubCpjXQJYXAZrZEaAaSC06Nw/wYws0wAmcutPMLsKgtpO4
cypQERiOgmprIs+Ihx+JZkNyoxp7nu88rnahds4gRghispe9pd4UZzDilAIIqr22
6TqDjHFPOxy0I2KN+o71DgkDRaPF5lYr9LTn+DSwzSq18Dh1/YsZeRvuT60X2Bit
32LoD6LAJ3/y4+Ip1xmj15sEE8EUxbOu8vQSbQJWLc3vzdPgw3IRJwl4npHzx0dh
NeLx2DEKN9RZcP6eJPDZN3oTRZkzmk8sDUHnYWcuP9+abgtF8zM4VBJRJvJac+zM
Brqzj6678zSoEX9PZ7AkYvZWU8StieXWUcpVRJmKBE4mOtMpobnBcG2G42BYfbbB
InH9w7Zk+qAeNuLQyUPzYZ9mcLjcyIc5SznQVHeaRAEpTt5OUWr/4IwH2U5um+mi
nYK3/8tQsxlqpDZZhGLtJ8I5yK8hXhZpzerPlHfAqlu5zlSNKTUc5QKt5oFyH8QD
pll3Zz9hN2WfTkSYCJX0BeZbC8RV728mtv0+juxw7n9phXqdSHjEdFf02sx6PN7p
/CDNeL/cL/IlUh9kdsUQHwP+Lq9qpcLEyfXJS60vEWGagHs3nG3OWGK707xqMCom
LrGkRkkP0JbQup1Bj4UNVPJs1IgPo6byiVkGV38xuNVXJLyoSVJus786dHKe1zJZ
PfcIia/Ep2CNLu1YW7EySdG65/KmojuolgyKnoPewxT5rOm95Ib59NgsFO3+j1us
Liv0wXB4eciIrMX0n/zJigK/YCeLaFAebGDKjcUOV3mflCxzcwVZhUXqCx2CvdpK
SU7ar62R65EeecyC5HiKYDM7D5gtdZsUxP69FreEyOtIAtYom9qRhzjWMSS5dZwy
1gj5zy0HGmlwBoZS3IOyNiwEOKVAXVZO4wJzgSpdi9JGDwTf7J+jaUxM+Rjsrq/y
8BVUrOuiihSM7Xw4qTEDLPZxiD4Zc1aUx6qFKZ25CwaSPi0QXMFL0a8mgM9PnbG3
5j6QNiS0wIZ1OJxCog8dBhxASrcel2I1qLjA6a0oqrtXHyNtDVrqQsd6rr/xsPAR
uRAFJPHMyR7wx7uJwUkGjzGFUPdv/6z50ghXU6kHlSiYv4CMP/iAsdPizG3gbSoZ
e0IogVMYnAaXLnDcq9dmtb9hh3ATMMMzSSj0UZn9GwoyooxHXW5p3tJGoD7V+2EL
k+BnMRjwIUvE/uKmBeefK0H7q+e/4OVmVd/2RpyXvIjdOJXLFfJNqAubatDJSrLq
pJ3oi2vtOVHp90Fw/LbhfgI59OxDInmufyUVQnHnIxalo1ebXN0I0w1Jcd28mHh4
Yp71XbRE+8OIAbfliTmVTKNKMd1w9d4ZF6Ovzx0gtN8Cy3vIrYxjEdwEoUyc91sP
587jMjT3kxmvl7QQYueB+pHeFWukCGpaGV+gSP0gLUkDDl2v1Hag1juX/OM96B2L
9IgGp0NHELd7pANCoLUm8Ie55kftC/Ae3f6zfhFnFjpChvYhFZLpggyWOinLiy5l
0Nz1Huou6IFuQ0cXvDtoyvfnROZWpgLRB1zYB2Kdi4s8iuh4Za5o34m7PcMw1xie
fMXHcP29qWL4Jn9k7CJ6pQUwGyOPBFr9wPMsyBCvmlQ8yeHqnyKbJr5RaUbzZtde
KGEH7/x35m4oPZ33Drv8/oH4ThjivT/WTytWZGOzVZfCU7WzmpbjQp+f6i6tLNSV
hPp+Amml7urCBdIWaXfUZRaoxusx5jyySkmbFlUMzE+iVEnGoYiatp1TDzgq/v9E
+6lXpBrfa8ABYeN1zK2jHvSQm1+F0Mj48DnovfTU6x7zpfTTLACz4EPBcOHcHl1y
8P8j7OlvVi4pB4HjjQugcgzztRt2icRnmtlKTdI2LwNt79kg7+zghYoBIF3ad0py
JcYCGYFpyrRspoPOggSCdL2ZsYjeOr8UcqNVC9r9NqUDq7ZHFpboP1ryN5AY+SSB
SDxwcVudCLgB60RcvRbdNQGEff3S42dwcopCTn+ccyR8Qza5hJUYoD9O9Dyh6RvL
xMPSd30d3L/1L9QQbB2Q5tWFgapZcE0DaZR0D1BGy7oAXi7CXAtKHeo/mD36pNCr
p+E3noeVKM4pTR0vCKHdmSaH4HAcqggwpj3Y/SUAoHn5iNcJK8ItdPmAMrvY4PGQ
`protect END_PROTECTED
