`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVOiSd3qBbtyyAqq8N3Td/vtUu5L+YrRD0Py6RWKjsVnviIS3yNp57SuKDzCWh12
w9MrTMlxTxIxVCIIpqF8UWa7Y8NoM3XSINn8pC4lz4xN3saPXo+qLTAOMZikPbJB
jgOGFhZe0rQZHbvMMnHD7ILfbHCtdK00YhDR1cQzBShhMFJ95+yFNSXSZSMes7g4
eFJycbdtTJMwitQt3rcqm3ncZwm4I3PlX+dGc8fynNHJl8U47HtUgAn6zAoOmQ91
dLyyYxvpBMPZuTOAQK/SrhL/IkyGQfgkR6/gEj+BeTAQa8nZsntqAlXph2qVADRo
qJnMkmRhUYlNF29Ry4xl+1m2wtvWF1A9v65lM0u56oujfuu2vLWwtYcZUVDt6wJG
Ku4JfWacjv/40VrYt1+s8jBX60P6PpNTAmiZn472DX1Dt/ZIxOY4m1+V4Hak9rgu
WwvTKilbhLqkIsKsoK3nR1peFah24TFVkIN8rv++bvg=
`protect END_PROTECTED
