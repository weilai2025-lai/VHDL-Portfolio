`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMVX8FybuPQnP4D1tegmyf7IWT8j29kz46ecBQAnpD3f6PlzGkNXpYJ70eudWx2I
c3SdcIx1p4VSSsCtOhGfnxBbuhasQtPAV1pMYBIkT7XrAhoXVwxajcVPlm0bE3Bp
QlXAgMib7VoVylHSB+Tm40eyMAnQou7F7nyhFqtY0CvDZUNY6Rpl2NVwhJGOJjHw
i7j4bRER/asCGC40yzVMLo9fDt3eB7QQaw2Kz8kz2B8Of2Vuc+u6N6tX+XevNUsj
MuoMIbyOh1xT22WDeKc+Cu4NQYbVKYCd2YKGB8M5n8VAABPUb7BdOy2vhshQHOTE
OybAOtOlDDgHhFM6AmyjmckdTOKgD9SziLwtNEjKxM/h4Bn5OHaGcEmiekGxmcnl
ehJSXea2AKHCEvPrd8NL5InHZ+NsKZKQqR7SRDLxlbP3TqGeSyTxSqRZCGXnG63J
JlBnLxhAiB8f2QGmuVX25BNuXPx/KbXHUiq27j+/NoM=
`protect END_PROTECTED
