`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmAemBtzkwXuqddm40bDzsa/EFqmmuKFvfstZHdu8NFR36cQeTInXEQNTrD5FDKL
3cqMjXoJaV30nnbVVyL8v9Z0StKp5B+TP25a7mFTkte2wcY2WhBcs4Ost6+hoRQm
n3ehG5MMSujRHRi1nd/uWLgF0XWUpR94VioX6sijedMULbrjlAhfYhSNSBwEHxMh
01QF6tbnipaVTUK/LQ15gaGIzyneE4Ry3I1L3TpeMij7IUeP2NsUJeR1nLT1OffI
LEB87uMglRnwe04S10XY5BMYJuGyIzuf0rnhPUpCVvAni49YQS+XNzKR6271q11/
3bSw0IeqTrUL/3I5VP/PUngHD3pDFjCuq47Dn4LsnoXsfIJo6ixdayzk5xNrtJbI
vya+WuSswL6Niw/H/ToePdyxS73UeIhBmUyjw/kTsxhvmQvKxK2xoh5oHyRtWsd5
Yk+yDhwg8fZrCUwNohH9NVGoGEAYbcjSYaPwC5h3MoLqCO+KwI7GYpiN8LK6u7EM
CUI5ozs2DpLTjOx9rWiazuCZVnGGJ4T0S1kY6huO07n/KZMmDmWtroIxJLqkDaSk
FzUo1lUhxQfak1TcLrCMgExQemuNYeeGBliPT5G2bAT6QVFSQd2tHD7wME+XRLUz
01Q5nAsDIzOaZ6JqgRyPKYICRTdM/AnabrgCuPj1TVPt68lHSFkwZ5tpRoP5kN62
e94BE15VgekpmoQoE4GKcMAdiemL5ebAtzkETodDLGgDsqd4WJrKGnz8NJ7BHNFH
UAokhe4NwL5ms6YuaqQARAYDguEQBzDCcl7EMr+XTXWi0mEC8OXTLI0ar0R+/xCq
ijpoyobX9zBAWw+LhsKmyR3PCM1T1xHMo/mxiIKJ9Ym+4u0DBp5nmtz4UXzlwZrB
Yi5c4LYhK+l8FRCKM1qYATGg8p1hHGY2Dkm7KpyTrMgJM3LFEgFNHKMCdr3CMd4e
eBmilb3cMxeOwFM9VFh8xkA4xB7CbIMIrooZGwg5XfZjRmpglzav8Vx+ubYrn934
SSzryhSyLUce+lbUjciVOD4sbJTISWivhHXYqVFPx9JBt7TgTptzudKnbGSltvo3
bXkluccgrMb7t0MqqNDSl7hmVAeyEDhoVP0rSZEbGSpA5iq8gyfAw3Epbd1JDxnC
xc6YpH3BTBeIo8OY1i6wuUo4CetHOXs1RNINOk2jUouuAVCrhRl8+Dmro8/6uiIn
a3cyVfsEy8BHXOUhY9jSOdLUa9I2URMtnylMmMlbXtqngmV2L6CjlBHTru/HSSKB
FkRwunKa9relwOnCQLBhmZ3O8mYo5AOktXNPz7qrmp2+TPVCIVBKascBETFkR7Wf
o0Sr1U2AXGV/v5Go1GX9FEg/tslVxDOJUGpgb6c2tciw0pl7xwek95+RiB8+WJHo
+8gjFuFPFGdmr9U950P1NzIx4XnZ6cb8sPRw78YppPX0YHFOBd1GpQ9rBMSvZeZR
WzaWImRnu96a/FSE1svbxj6poke0BrBLZaKBGf+AjxsFKe8ZMht+vMAShRXvZmfh
YC2eR+fOZomGTSem8axc0JEAgUhrIU8Hm24zXz863CCUAk0VCflURIIgIB/VI31C
JVq6YkvI58tV6yJNot+Z0F80B+twdEcG43fgaWdilj+w4Z0HDWFISzF4n/z5Bd5s
T38S4kuVJ14FDi38PmYEUzKHjWKa1/S+8FPOljM820owKCZGzdw6AbtQejPFRvVv
9N1RaNnc4nvNreu3rTUXj+dIFMLLpjp9n7KcvE10jfEZC44O7TlRNt/4N+KwxPas
WP9+wLlcQB5fVUf1+rj4cL85TWtgrU8MKA1h2ckp3pAJFFvNSp5FGeduFTx4H3fM
8xBok6jmtCZYid8RT1kUpnqjow9FwOpFsJkI0aJI4HQDZy4d9/33ZjMO3ouhr22p
QL20aVoET7Hgci6xCiu+mqFg+NCNaSCg6RGzUu6TsuH+FJ6VdbJWrJIX0JUqWskX
lz3Jx2fDdH6sfzAbe/q7LV+dv/OV9RAC5O13acyxAsuLW8ml7QrNg1OFpuVbv3bV
5g9dNjSjVJF6C4lTHAUbltpLuUg/QuFRPwFHgToH3A0++rGXbJpUtXHVRAqGk3/z
XLjxeg3qlL6/vsSZ8EvSXLopWz2FHjb+z3UdkuKv+d7VDAXO9kImql7JLzBEsgmg
OWrdfFmh1iJL1lf626Km2LQfEHftYAYp2cBQGOOKrMwi03XK6jMpz5gYJAQ2jXBw
6Jz3I9xE6RZQHYcCJskMJ4cr25KVwUj9vBfKQ5ZvmbWaasIoqDFC9aseRBLKG2P9
Cr2hOWLOzj1dF2D55T68mDEUjgFMmFFQeYyBZ5bZrZ0IhKoYib0yasEQQwRtMv2c
pajh3CBiKCQsb3f9Cg3akPuIjOB7OaaqDaFfAxCzOWCxqSbonsMMvoOV5od+6kuF
ibNK0WLdmmqSTLO3d2BfkdKvy27VZtgFiab1RzydO37kRz2QKrHl7XRwO7mevOcK
FzVJQLi013IPgQNO2YUZl7r9YlKgufAYQJ8efDZbPv5eBz9A+wZma+7FTxLi+viq
07zOtt66MkkmK4xvXYzZBadlCeZ34gKol+zavc70JziAFiSq2bjgGNDYvgvG4IlK
QvBmDC0Axwts4ldE8lT8NX2kcABZRMjieLMNVlKMuOJYe4JRz8GWqUyytXONSh0d
TSp90OIGvTPoPVxI8Sl5ERzoigPa7r+l71T/aReYlizuRRsq5Oz7ahzJiNNUMD3h
vAQqPVRJ4ntoeg+q9Y1hPMLNUpLP9MWTf4RBWn+vsse+yv0K76+a1mJTHpOpciPu
jGWs03+DaiA7oou6iZF8thINIFDOY7jmvEzTuDfWgXxIoAf8cTegscZvAGu6VleM
2GM8Od9+5kpS/HvN9/3xvtOsJZieqtykKhaFz/rjhqooOo5fZ1XFOfLqGKSlHA64
kHAxakDwkC4ak1lbIg8il+1QBe+9OPvSmceodVEySwSOi3vJM5N2CnAJHkbcvmRu
SOdCQ2GKX3rcdlx/lUtVQAIdvEQeIfwdkJmSjFKooOCPmE+XJEhHkVN/adbYyrWM
Qd3slaIHWvwYsvZ3ZdXOKw9KBYDL1OYhxIfniNKT9YAj+lRXNSf0R283CU/DPBRE
FsaKrrXuT2HkEGaWkyIuXdzFnkwBS5T20WvEaFBvetOA4IF0APcuy8C0f8EZDST1
TwqyW/mHHxDZtcnQMJ59Q5HTRgCa8PLvpmLHFrsLUbwxc7lLKW8c0QJTh/IksZ9N
8K1LYpwoGUP1tuQcNaFfXNz1TCzYnmG/8fbVkUihpTnYxGuka3vM1apVkr8ABIs2
kfwcdLI22ek1e/aq+mNPWVIQBlrsvX8ATEOFFbmzo/uudn+vdYJJkNpNx+Gu4pRb
iDfV5u8k+xHTap6pw3T6xCXVVuOLz2BUaPTzSOqYxFeMqwAYIYls+fBLl7TfGhVk
8wjWH37qVLRkCzB6jr43YgFm6bKqm8FqxWb8ript/e8Y3KUYjJfeC+kQeUhgMOzQ
3Y4WGa+RfXCkN2iKcM++0yQ0Kh7pzrk4hZTtn1xUStNqgBGtVjEAWCu422BH/PYh
UJWT4oirCuvj8gq9ZA8RugSFyC9PaMnYe41bvUJuvAkRkMD8Ah/NERsMA9cBgJG7
rPwoX3Dt73Z+GEODMoLwNgA3GZc1Oz/8ndqiyP6ofC2ACZYe87p7hMX/WSGS0zE9
oC3dRS4jaE578VyQcy5wAtGbG+3XUSlVNWLgLmtQKFBiHGvGZmDTXa1CDSehj/Fz
DJrBc9w5YDRtdMAsPAR+lo9OapFFPxrdR8hPkgA6MCZ3G+EpbWccWOhmQepo94kO
92vaO9/4TLNNJ+d5HpKdlQRWg2fRXke9GmaaPCd6pxOTdFDFNwlkqkqZzroeDhI4
IrcbP7TXpeRvLVewjapBfXYcpUDyEd+TaRO/tNSMrYfk7z0l7cxlOU8CR3CnjFYN
KUV9YpB1VryX4m1SNUZxgl0DWvNrlhU+nKn8WNSYY/IJtpmmQ7R2coN4u1HfXg1R
zd84Gs4tAQxwNrAlmzGJh2buU2YMAq6k5ZbEvJ9j1ndZEKocgHPbN6QZryg3CQ9L
m6DPZCmhhfA6Ar684nqvl905V306fShIGcNEIn78Mf446yKSvnfcPkq9jZUUQ1mV
57D1Y5EEjKEOwUe1E7NBOp7N7LlBERNqkvPws1FXw2d/Ogcv+pOfTihJhmWAkH+O
vQ4VbbahCAj3kTmG4vuogyP2bg7HjtmEXX8pcx6hfl0Ze5ImMolAMQQTerBYuKI+
BNyThBvBhSuXP0pAQlpPt/ln5qA9av/2efxPMHR05WyHlmPxlLdHDOruWFNZY8xg
EzIy6g+l9TUiZ5+hzZ5FaYZ9xLsZJx4DmSkgrlIz1a5p1oepAQgBZWHw4Nqy9E2Q
8gxepZYmdw0op6JctPhjjVyFTRcLRcf3XdFdX8qAz/UoYXrbzMHtUqgRxa6wrzmj
uW7ZlSfdahcUZE/lhU8atXkXgbGHSn0s2u2+Pw+w8tMGyq+77RtRyuvHpUVpWX4E
EM6Hvo7geLnVgGeTjyZ6pijhvD6lZExSAV0bSWfhuaD/v9s6ewPUIVomJZkqHOGX
oIbRcr28KP3tpGN4VKCdGA==
`protect END_PROTECTED
