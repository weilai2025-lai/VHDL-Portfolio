`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBU5qy9FH8mZVuLcJiZb8cgKkrRTqjyv6J3x27VCg851xHH+fdKBOWjamWvzKXqB
d0ZhaAA2TXQrnKo4V6blQflFnzMdzoOAOrpgGps4rTz3WnSgl8hyiHVKjZZSyFFD
+1+7i26dICGvl53UzrKhQPZHeweXYrz+XhI3ighMdu4YEdJkKXEZ5juZNViii/E9
MSgNvgzhmce0hUgaKwTk3zD4cvlPEJw42hQsauJrOwyFGt9+J1xCllKkGimyZ/Im
5AiH61Y5rl6OxFrlFlSJOqjz6BypjCWcyHZYkEj+fxSms6evaw5fTw6Vf6mq+SdT
DkFy+uza9sfAPeZT5CcHiCNPti+Eo1vfxjFmmOhAaZUAuwa4e2Ckl05spfsudSfQ
3pZ0agxKK3kpdDLIjvlr8Q4YNVLzbvI4hIJfbZWdIyQO9BW6mH9gefVEvIYTJZ9U
JDS3jCUIeZk4MzQDzwdEzZKRal/r0Jy8NRbcPAl5/AcxhTaDpoquKnjd4TPU8/RR
NglfPQ7Orp0nLOkHh47l9uItj2YyAeyCvYNMqRrzWRrVB6kRbw6NBifD20RolWpy
BYbxlIFKHFBMVhUut5+Tbb/t1N71kFufH9d33B7Ls8oniad3BZnfxPW+iFUlk8vd
ojjIXKvMnX3KqDDuirZ5ZtRIn3jzDWdR9Id7Akn3nPX5sRsBVcTfbPvywIfhpBjI
N248S83yqUctWTq5c3HYmzjwCTO7LsJmcBxjgbH5/LcpMI9PFWNbY8JBFl+HTstM
LWZRx9QdimdvCXde1iHJjYTlzeizvqoDS7FFAJefaXqIzK/jyxz3IQpU7ENKOfKS
iERk8HTn/3HHey1GHnZ8bt8BzWPhobM6VTX9b7/GvWAnG/I5UeUAh1gUcSHLlk1z
2WkdJ/a4V/wKLQl73kej4FAj8P7XQZVf9BmsztvyWCBcPgIjq62Ar2tcLbpZxneB
TSbl0uEilE0ohnAqtY539RCmsEnanSMsvcm0VuzfPJ2kFJN+FOyr6Dk/pOmYgSh8
URzFs1XSvwhfpU3KTo+woTrwQ6ZugVDNjWIL3qWpPgmohl8Uhajy8WOJYZTKuyO8
Brn82reK8Qx1pfhqgWdMZ9qTU3++FZE/gGuJZ7c6+QL3EPBNNBLmoCi5WhPaZi9O
3cvlVxjFQVHivWaooEOlPaC1/5MxfyxDu1DmzsE/mR1YlJKqb1X/5wllqtHS2L06
ek/CIL0fq3WTD+DGzK2TYpFJm27pCPrLyGQUslTmwKtPC0TIaavOGFk8v8BJWLEQ
d29eJ3/2PcOE2yZC5wWHEaQ4G2MqBHoOuKPJ9fuB/QyQo3b3diEb5aPirj0mzQwj
7ItfG92lEWuzeOUWtrj6GxeKvvLD5JKfmq8gOQmPDe8RFv4vqR8WhrWUyyyUHyGe
cl8XU0HNw3Eed99GpsJuQbZlWljVxm7rG88qNIYblnSpKPRvNt1z4Qr4+x2aFewH
6rRa/Bxn9e1z4+H5fe41UaJS/xM6JDzuW+UTMVEi3vsDQYuzaKwajC7yd9x7Qea7
lIefwgCSxAlp2Sj219zFD1T+sbRm60PMVGZ1WfWq/kQ=
`protect END_PROTECTED
