`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5wcLnIep4CiCBKgOYdXS95b4Xyc2KVQwXenIUHzsH73WlQPabHKlVtDBIYLBnKJ
6nUu9jQJK7ScklvcZsfKvh8RBWIWkPBUd1B74LJQHMlG6LpWKZVqZsR3x7fI8Gw4
Olz3Di8p72wxbnmV4EfMsioj0vqNOhzSc0jz7TaRBtXQv7/Nrh7du0nWdJRd/33G
Yp3pDA+k9AAW0zILQA91o2Y8q4l5lfyHDn2qhYuGhcUz+oLVpEK8hIGGLZGBMZcJ
7CrLhht5hE0z7iJRxtPsd1LLfz3HSFQG6AMQ/Hqz2la1xS8tKqMFSy1G2zDKRQ+B
Wq/UuiiI8QnqQrb8HGO2zmn7IFz4+lI0faqiCw2n4HrEUXUQCvkYR1VhBEbM6sAP
A7syym9+J7feSBj1uxnbnCUlooQO5GX5+CaOl2G5PSIuCYovXA2nGPNE2/HJn6O9
9MeHrqkbhL8u8SsddfbDQsHWENniWaGn0aSMF4urCqYGZ82guIQTsG/qcNd7XsrM
syFBj6hgOAn1K8tqJiT/uEbweySKfQFeHA8wjlw0EkgkDfP1KjbB0dGKWPsW/XYA
ObJ8G5GAM0GJonNvAhhGfuOBh6SkfTkL3fVW5oKrvMHADPTaBbg9mnh8OufO4ZeL
AsVj8yA/7tZ+u7PI9rm2kAUX8fxbfnsKxQqVkgsW2oYYNBkddX6lnMX1mK2i07p4
TOuFBTibfGaKFQrq1y2x6Q91ALRnQaqcNLP6zase7l7EkElALCle8DEw37Q+H8aw
j+ZidTSX+WlUhoChoNx3L79qyA1DOT2MwNBGg5rYGVRwRnhQwSM9U3DyHMFQW+fm
9LNW9yQmbAmqL9JboNUztReW/e5X4qOBwQ6wCujYskjCGb1JB19/USEJVrGWo2KY
e5Sr3SrYts+PZMVxGLOT4mBAWs8n4vFtkHRjbxywdylOZ1b+hFAR/us4SIcHZVww
bEb4e+cRCxAFPTmPVSVwJ17GRa1otFJLmXnpj4kgK8RSbsRlRRjpYPVt4h4CzRn/
Vj4pfxdIL3x7Lp8QdkmZ4riJBC9qEGihnXpLPPW4m0HaNGJZIKt4cYWd9eh3LMna
DzzLbumdNlFfc6KxDyRqQjXX7HTMEPxNmhDiM2HDfl768ABXHJ7svv0+8TEeP9se
4ErbHEjm1M4JqKF0SvL31kBeUouf4rlViYaE1Ogac88+rKsx52ctdkG6KDQzN1Lq
dUHC4Vb2YsWs2e2c5nxLtRnOy1KEdQJEU6OrTuRslvai/StXRttNM1KEUl0hxNw7
awLyFKNB8wg2MRJ+3jJUtw9Hw0g/vWcCsl6mfa1CWGbLhuAMitQebR7s/RgB452j
Qk7trJOfmRI4kxWFOEL2+w==
`protect END_PROTECTED
