`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5CAl9Bul1Z6TuFOyIL63J7Oa9KObL6z6LMuRuW149JwqG53Ujyy7ZNVmP/LkClI
6LlMIUI27xsXJlDlAJL2b6HBLtV0k87HoQuLfOjJUmQyREebdkNzeQlKqOeOmmV/
OKsGtNzNrw8D1JHU9IgpfxkIyaDvuciG+nKzRHStV8oGAlNwJvdIMG386IwZJuPh
3D2huoZlimKwc5eAghcvUdCcoExcI/D/50aRhvEqOh2/K7LRgRt49Rz/cJkG5Lvq
5nOeOFMPrUfsTLO7QGXUWFOTmHroVORucXxetBsx13fVkR7uBaDiCSVjoVf+7HbM
1zTBAYURtXBnCx0m1En4/WCuUry8Yu4yfXcjIVLzavcXxRaNDx1t7CSKmxpLl2gw
jdoLGZRlFuZ9i9C84eRcW6KwAYa5wvhEgRP+4/Cw7nq7ESh134lWiH4whU/TZIp7
eIqAO9+sEaZqhexZoW/xCXqGPcdCNnWwXwh1wridXuPOlDdNsX9C9azQikFaQ+xA
G5gZ8Un2sPCxWtel9bKkLRKVgLTLq9LU0H05RlS7RtcJ0qkPu7MM3OAEEfpBFWTK
cFdLcL8gElpZsuQ635bllTYilfPrnS63lPvMNly51JmoWsb7YBx8QIhcV97QEOAe
jJWFHaUSTV0eZ23N/niFMF4UPbMRNYP4A2u4LbL0qfg4w+T5E5yAdUDXLNpSjbFq
ulNwQiHpYgvEz7mS2RquRhRkYzBThc5f16Pw3kFpUpdBm4g8M3vJyxqpG6Fs4AWJ
15YKPjpDo2shMVfqJrwLkxsxh1wqZy0WQ3SYdsTNNWQ=
`protect END_PROTECTED
