`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
638ydQDTShX06NzIbmnTCRG0r+OzN+VmS4MCyYMktE8FKx/vOAATfEZGZpFKsDD2
UxSfeEK996jJg9lRFxI+LSkLuRtSwhlaoVbaJpcoLS9YrQOjMVlaiGvKOdz7eysy
HNy3AnlaKPjCvR/EE0zzieeakXEDFUl7Hc5+1v+VVAYG2r8Rv18tL6hL+U9Sj6bv
9c3HPa/5BM4eFXZs1wQwRws0EbRSer+8xUrokreRxskeZNZVHGKNenab5eIGNEWE
ns3qgcx/p7ycg8HOv2/FmKjkNxeYTC17tdFJxtCq+SDYRKJ4kcFWNs7nCBpdOUyQ
Dg/q4LZRs0a5swqfyykzJTfXBvA88Ck8KTBw0BOFLCQaVDui+fOaEKQLQ0VGP+pK
E5fLKQ6Nb7fSHJQT4UW2UtXU7S0hkKvqXKX26PSD2DH2DxkuMARNGx9QiiKjsqY4
ppZf5l7BORn82pJp6UPBUWeZZy3lTn28TENVRJndQsFmj6xzKAZLPM/3dfjFtFqv
Z2q32C6bET1jI1JMjVQRHycfK6mP18xI++L/44H2wnB2k/8UBJuByA04vBBKi2f8
tK0rzlUvU5GyypW9ScfbIYBGy0YricN30cczSg/E7uTPiZn9yId0Qm3yn5IWyDSI
hoaUODeqWJhIoMogK8gFsw5c7Te/dDlfCOfgbhaU4KotLQ8xawnrIN7enCgoo4H5
Fo2CxfdV02jIPR/JSKI7e6pcpQz5qPj7BElIuK5AULGxY8/SDcKiO7Y996mLnNFr
2b40WKoptXXdvInh3WvBYAOr3J5cIk8MoiK5Z7BOIiUfeZJOOyZeAwX2MilGZt0x
JfOO1w9IePv7YIfnFr492YSyaZTJr8RjwuFljtnxMktbL1bfkZiDasg3PyKbG3wJ
B9PcTiT93dL5g/x0vhh218zvBmXm8N2co+nnhWl8UR29r89wnCoNkGKrOM3iSKMy
yMqqrAmV8WLmz1NKn7Z8onRbiEVLlDSv/Npasu2Ia0vxZhmPjlYgVqwHScswF07r
LNw+NXhGgP4EPYb+aQ8nwJxsjYeDGRrtnP5Wo47ASsA=
`protect END_PROTECTED
