`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5Zdlxx8oFnEP5ykCzV0v+/Gm7t6h4TFo6z/iuepc3rKfBKUuTljiL9TvrYpC2qk
1I5WLWO17wD2UaWmrwAH4NyYtRuRrOdFRSFsxi9UFTkexhWW5XgMa2zUrfGO+bql
MdsRKOS0Rkzqj27CafH0QE1IuHYnnwZpYg52LpgO/1/cTwLNTFLMRH4vb+taIIzo
hsbT44aOUAB/XA6BMrz06OqgGjC4SmQsCbbgKK4X+DUFnmOOAGimMSuPSHSSKD98
+Wjwof6QFkTe4pE8XgXJgbtP8a1NDjGd18Y3v9a18qGcLd9Mw13+YQyeOGIp+Yg2
cLaTGkTw5nI3iwH+NMeEh0tnJ34Y90Kq1WFWIUI53yx++p/2XXD4e1EHj2ax7b5u
K+bCZzti3f3sEAX4J3+dZLNy1gxY/fCh7CEXknSy9XPX9MO5cIZgF2F4qUpND4Xc
KIHJPzAj+Rmfu3Bx7df88iy1Un20awkTqka9zn7L3PlCGY5f0CbmkaFe/hPN/5zm
5+cLi8VXPpCqOOqxRfeQYNw6TgIEyZSLXvJ9Ix7na1s/qIkpOZTMYBjGUW/yrMuO
28R7vecXKoGbw8dtvuxPyv4CCwnF6b5Im62lqRoN4ENTayv6XMyY2MphfV9Oljnw
TGGnGBatUWN6Wf4ZVjoxw8bRlcJTZIQdL/cv9zaC0sv2iNF7BJEvxHZTZJubKR99
uDVpvuLkARbIh35tW37SYRoyd3LjiqjjvYzRKum/Yu9qrZOMGwmnyUc3SojLMKDt
+sP1U9XSwsWcLXGJz3vtMHcp7NBxp7Ot3+0jRcTPRrTmkgwk7Vcn7bLytcdTi6by
I1d7/AYZU5DwbQwWc8sWzGthw4eQFWP/kjK1Zu7J3KUqyY01UA2T+I2Itcrn7UNe
gs7SDG2Fzfv6d6HjZBdqigwV291ffBhpcgG2s9evqCGFaOXyJ3fuRlgOhyBZG++V
+NFvT/sMW9LQXpPXeDUZc/lO2OwPOkXLiVsMTg//uvqBEh5ohafJTpd20rtPLeEt
FbAmalCtAQr1gkeCynBbzQ5HVOVN7rlulqhGT6AxtkFIDTkNpx8r/gco5LZHkzeN
6/0Iu2FzmQ+C0Ml6649puA==
`protect END_PROTECTED
