`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y0t5fxD9JWUVf6vlvfO+lDUAbySeh4/Iz2a8VZpjNXh/6W8Ri+cwaC4Cc0YKQsCd
H+14N7g+AydgPABVvk2TX9RaU3lRubZySS/173eG9Qzkn5dTetb4GxnI4p2FaZvs
dr8Jc3+HnmvFRxbclh+XYLjS2qcaLZjFb8fIfpYtTuGuwESihIZ79E/lWmXmHZfT
`protect END_PROTECTED
