`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
13mntPG1yhhyyPh9kQZN8bkSJ998Q9lFhmT8bOFxweCu1Pl5+zDZu0Rgjs+NgJ4+
kVm6FdVXWcSqBy8TmtB0oQUejJAHLvzfNCEUtPf1/x+paeAn9hwOmyRpDWLpCrne
d50u0rfa16S2OP2BAkIVHtCuo/ca09z0YGLVO7DvhEIGQgPleoj9if0SuVmhZkZU
rXWa2IEXwCkBrguK7vObuOf16abxp2BP+B5SM8FdST4xwbFGcT/VEQXUeVBULn7u
ZYxcFRR38FfaVem9UAGr4UFUyJ0F8Q5n+6MtNrepVL2QbsgFjHQ4YwhedzjDKq+E
mDdUKP5z1OeXY3X2/2gcn4Xx7YQ3Y/sNQG5lR/WHwpfXsT4etidRy6ySbXOSZr0m
SYGYTFx+sDwQXnK9nw5K00nROKE0gqJs4CcitlXmb9oNtbzZttZqbH938I+k3ZNs
Ah/8F7Y7887sRy6OR+x7VWFhOfQXQzlj6oNstVxiVoY2VXKF54Z0vDRU6t+Z88Sr
KAhW+fVDhSRo3L24DCfKRyB94rsUDvMb8yyVIZOF+ADYzTy7WBZBUncuMkNwEu9T
DtILILtO2fR1KQ0L/wZ56YCAYG9c8mVQDF9+YPJ9nsQCnM7NTDlleu3OdR/RNycj
e3p3CWs7nXQWmfq3oC6RlW/AD26Fkq5Zp7b9LvkARc8mYi57uY/SwMpbGFdQFRiy
Hnol2lajGeofm+ZLKc3cdWfCE7+VRdXX0mXA0qWDMK/u6WnmxQ4XsrRgMwtFdIVu
y/f/iP3qCMcpmUoJ57ay+EPPDlwFycNprn9xoxWNB6eovcEUprThfHG88NPT6dWJ
Se6QH+uUldAUZnfS9NX4r8LyPiTv5oTU9mRhnre/dCJRZdJVGjtIFwpi1utxGxtU
ZVU7vSwjDVei07P1mPZho6bEVHrbZA+TNDWtt6/HuT9/gQjB6brjOyP7TlhnO5N3
ytv5va2JbGRyvcammKI6Ef9RTUOk2uIKqejb56yPrbSq0izAuCOzw/cPUhMxwkZK
y3Metd8MNKDVNEAj4jUA3+pnNddTnwZMP0xNnXZPTwlWQczfjVrcbay55XtYY6g1
qZCn9TDcWUnphVa0zs87l6XAb93VireSao7KLHx2Q6gAqKH+Be5uj7M6SqBr4enF
0h44XV4RokC4Kr7v4VYIrx6DwcITmy4GzboOhyVY7ht6qnKceqNk4q3CXdjRTwGF
UZUivCFSYSraaqdQ08cHf9vYDI6p5qh9xgIr6ioJ1jWgIkxrDjxOBNprI4n96xXp
xokO1SEy+jJcO4gzbWYOjJ6w5GWKnUJwqAxbASGuEghLPYd0uKa232qpRVuUp3fI
ErVcHJbhN67imALYe5cbNXOv3VPrwVYsAjRcEwJjxSzyT3Nt1Ax+w6U6Q7ovT9ot
6IsVycJadVI2EykYS3mKPK3gXMzd0HnLuHUveVi56RPPMugUTO+jzDz2oNjnM2HW
/A5ursXT4By4Wu+zp50FMjmjysGbVasx3EZci/9cKxBGtiNXqv0dU6Xwj70/41Gr
XOw6NzJMYTd5Tu4zQ9uPxODNgFiE/GA856ZxyIu1gZL8euxLu7hKrvzpzN9t/3ys
PjctCww3K1uxY/Af9GeB3nKvRXVKjLTXWIk+f5MRCK8RlCaEOAy6nwYjrCxGr/OU
14rG9PCcUmCVxsN8z8ZkJafyk6GHW9r4fVkTSJdK4y+Tj5tSOaTjAwOSYP9tDJX+
mvx8JT659RXDa/4RaztJXeV+l6HTe/qki/Yridcakj0ZAeUSHFvM36oaO7P1Nmuu
3BPrHYusRGhd3RXi4HXiqbbzgjkzhHyVOscv1YKfOBCF3+YAXj78iyCJpS+KbcJE
6TdSyHE7wzVZ81Y7DUnzUBhKnSDcx/r9phIkroTrkO+K2tj4W6MbumWXXaL6tX/V
V8X1WxHlofcieYl5+iivt6YCAzUDZFVaNErkhvm3OsFlREpnAWYZi5ZYYQ3SihjN
7yCdBbJDFF967we1fAQPF8u9K3THRRN9lu6rAbvI+YsMHIuglqNMX5Z2toWZWLVr
3lHoJhoWGbUURsxorZ/dKG1wQElQTaFUiYWdxPDhTr//2pVsKowANwZE2HRPwU4J
crmjlLXsGxKyUq6gRijZkDMprvHol8nR1/1QkU2B7S0vwYx9e+OTKzZwNXiHD892
z7f3SvV9O0St0eNz+zaDjTRHMBUz35mXPbliiiuzKK8cDHUekjx2zqq1fTanEvhr
jMMC8tKXo3uhTG4UL2IRlCZJznen+Yj0RqDfaymqmIlFi2HDdI8qdzl5kl7bKB3/
A8imcNf7VVwlAOngOkYpajoYh9dry37fb7iXoAr5kcCVFoKnxE4EJlAfCyoI4YNK
Te/yh8sXZIArTNvzTLNC/FcmtBH+Yc551PeeXfOl0HNVCQwpm4UNI/7Smdxrs8Qs
lD+BCgJo4pbIiVnPqrfu2jGVN8jjzJEOT9EAKEeBgJaCR5Y79+fayQLpjrN1SvkQ
3P16CzCZI6sn6BAm2QKRggzPvhaSReTR84QWq4h1e6h3W32amovMBfH25Tx4mWph
3JxVBm1HdmPFSCarN6Y2vF51Z7UHNFDujGbjg6DtP759aU4D3rHOg+evmMEWhV8E
37DLlzqAZza/dxmZ5B0HC/e2K+QJ8eg7lC1U5OOpBeOBlcmlu8RudRatIZYtAV3O
npzdobN5lE9D6+f7aw4xrzJtDHBM/yEEsL4mvP03nsQr6Its0EkLRS+tM1b4pEis
4xdRGFW61fhQoazI0kGzDDvTTuocbyhSFOKBNOlM2p8HIsfMpugeiMGZIUgPOY2u
7z1zT5jSTD0+yOp2ZUXkuw99cBmSVvCacZ7MO6heEqW48fH92ftNgzofq/TjlDws
vFRkKVVWKmPwMTc4d0JHzKZwuTEXE51sLdSzyqnKXNQradldPK9qgjIZyL53whPU
MwJ+USgHbnZ/7B5jE40KoDgRBKieuo+jzRiJT6dflN26DbOXuQrVYfjaFOF11PXw
LtdfkKHM8dISXQmWjjrSFVPoD2nxeKPgzrsU8z3HROsV0UTOwFTl2nK8+lNISLGy
2DQjOd94sxOCIdn+qf2kZkgM/VWIbfQHEXEo72d36lDy74VCEZJ2Gyc/joat3Era
DBUOmJ9vuCLqp8r3y9hsKgGbJX1ZkRsuAeLcZeO424LznwosofGnOhk6WTAYhNJC
MUeWt2tPFJ1WrTZKcPgQpcFd/0BtfQRlkNN2OT+bJaRC0sEwQI2psz+rpWG80B16
YKoyY5CL8h97Vu/lb8QM5/SlVKJ+XsRV5/7rOPS7Zc8vPUuVk7uTK3gUntHT2cGh
fU2gKrqVhYNCA3lRL7MVWrhZvoCk7XEnOopgWm1ixVeOc6MCyzaITrwurEC0h6yj
bWY0wUmyd+AFUlmo4O0pUzW4zBNzqBK2KQrb3Uu7tM2iWJgl6HffqH+h6Vza3Emx
gGWlg+oC09owVDap2ZUJQbz59+JB0oqYkLYbl4q+abLcun3OJNx0NXgWyzt0LGwz
R1P9WIHXKVUINJexLAf2oohv9mY6KZARCjvl0eX4BIAj7YnNlsE5y3cQSmV65oaC
OoUXVhYdIXDCnJW1DxOi2JtxBZIG9ILzBhFdKHrriQnOf9Je176i0nl45Cg0FFwQ
FVsnCERSZ1/rkhsejKJjHvbEBLMfSPatNzOTqobbkpUvB6GOgwGS8fevMbmGXEbP
3/b1jb1ThNnK5PeXMqe20PQaV3oWBvm/SXdUKlKyCKoNEtRlphGBcAvoDCglr9rW
8zFA4KjikqvqyDY+8qavxWdEnKm3kfAGo7UJM0dFsBmgT7MJ8CB3np2dBgbtRgyR
1Iqay2SGl4xLztSny0ckuMK/YwouIBBXoWTCAaUUWKslZCbQd4OPaHQJ7/vkmIa9
D0qkVWQF0PnwziwBDnIZYVZ67AzRQGZJ+iH0xLziVhap03O5aEwloLC/06MRE6+W
0pVrXEfhzE3IrwxB3rr6R/QIFzf9MPvmQb4UI7Obbudf0OnLxEfGsdw8jU7/xQQV
eZ+nrF+X1jEmlwtudeaWHbBlqkeXDupc4g4QRJI+ZdMWQVobKMd1wlBZZeXmM7WU
2cmVgWQ7eAhosh6Xx+sFiTuhidpvRt7Aix/J5Vy8PnIcEEIoLcp40JlqISczBhVK
VF2nacQPnalxWJGw5I4kqFR2M+aQmd9H4BH4DXfyBsqiEIhPSDcuXXOZJ+ARgPsq
Xhj8u6whh4u20qz1HVPZfpA6sdUq6gxPWKK00InrG3hsPUegjhnMlKmH7KVzN0ef
0n+jlRXG0RVjmwhoxj7zPzBbYemoezAaD8Cb+nZ/dyso7HUbq7ykg4F0xHvgLoEv
em2ZFRcCd2TGDxqLxe/QzLMbFBFx67QCEvWvWro9og+peOHwDZ8vqgCcFUD8lMuN
NymJNO007u12y81X/89MExCAyfPURdhgehbLtcvWKPuKpZflP9CSIfOm4Cfum0AQ
ChTQwh+SqC9odjNqZjt0zaGeCDKSnDzVfnyDUEwrws97UNJbCh96MNxhol6bWz6X
7XP8n66cuHeNvD8plhd/CKjwgDetKnVyus5uwGAFYte+qw+cmwimtwxRb/unaBBM
wl9NJ6h1SsCWKt5wvucfnsHuttOZPJH3tPeULhQNlVrZcBX04NsHc6nu6j9ZG0zO
bA2fftt1gh+UhBFBd3B09I1Y6NUtX3fHBhhEiVYYbF61Q3XyajRjpRcqgtLBTCQz
AFUEslj3/b24j6XOiLY1qwOUmMM7dO2yQT3XENep8QuQHcRDz/ZjliAmrW8eK/3w
B+r5LXQembS4asu45/x/acBuTRACHXQRtrEZxAc9W9N9/iO+cNh9VSl3KYhRNsa7
3UXKwDVcHkRJeXRRpjkOTFigpPEAytPpCzYm+2mT1uPRwHO/hsO1PcGSeV9Swv1V
ZUKSE7XYjw+V4Qbi3Fft6iCGFG3aVEoLhGWXSH2DBlvb4SjSuADLPuf/Duyj/cen
2W91d+jKfAQOR2p+hZgBT0DSpOg47TRamgwaidHh92UAGy5IA8iqq4sjjZls6kDa
U9s/hBPnD9r55WycYB4EoKDatqhFGuqGZgVeGRYJuRxtKGmKlP/rse1e+d21B6ix
SZmYqvyQiLDH+yCnfPDi2nHc3/EvWIInnG9/pZnlbYACxnjUPyd5gSaavRhRBrcy
CLmyUGbGwE7jiNpcYDm/jF+lEKohAVp9Pg+XrJZSeFULJIFHUNPIN06Tz1pWLtse
8wbziD+Dpb1oWNyW7FpXNSnvEbFB4g8vc1inJJ9aPZ5+Dj6KwK9zb/LkGLWIQfiK
T0bbQSiE/cTdeTxhLOZSuTuTB3AXEWG0FMVtqklQCVXEYTpEewQwY8MoSM0eH2CD
vAqkPnrCFtpnyYW24eUI1c0UNlQeM/50L8+uxvhuT3/0m1feWlHcom5GS//TRT7G
FrKVxzicMT9ZznUfgC5G7sPC3nKWHsImhvx7VEULbcNGqhgYmCc9Yc2D8k2KKZbj
Rl4IrzSuHIuiTfsEh0ZPuHR+GATbXACcCpdfg12v1Oy1ApuG4e+vZkvFJLbSIp/L
c/UusasDmzU+hOyLWvxGbLMQN5+b7pnjQmR/qPnt0XbWxQOTFR6so2wdQbU+K7Fn
C3n3uW6v0lLeU3EV19CCn/14FCzfwAsw6gvDZODOcD7pNtujarI2QyWOUkrfzWoa
2X8YNUv2Z42uGSFjiT6KsKIXyp58OugauVfO82mLTpas9t+T9+VZoqdE+3oPH0s1
A9MTZwPBqT756E8tw3oGadSfg4Hg3DEcwid1h917ceN5LGj39Z06t6DBOkxfW1uJ
3YMiXD0kwmje9QVRsngFCpKbGgwoLu3sKool5adEVSMnn7H1zQGF9UJNaJ6HnieV
tDUahV3CwrbMh2u63hIb/bePVrZtCiaaVYIjRgzxFFzUkToS+Te9iKV4m6EZOVMM
/Lyy0ZexaM4OCkZ/0KDNYCe7EL2iquiyZzGm6ykOWaR7/a9/RenBRzrcSnGN9Ggr
6VPJPSnzpc7t3zyQXZTfTOloiRbWio9TCLrmlf3WKo966iNY33EyB5kW6zKoPG3H
8l/f3fuk+4CPS+mFlBcgkR0tHkdCnT5YDhYDNJeAdZ4PaS5tn5aAIflbtoarkjII
YLhJ0CDYbiMqCkravKcHINXt+LIjGotI3XNNGtKExJT1WIWBCVppT37SlHd/aKVV
zFckA0UL6S9KgziNmWT5kJttfS5cdpo7T60S2WuL+NCM/Nr5mugmOiDygkx05W6a
Z4iUtNlehXTlrhfTFt4oq+aaepvIGYTQx1Ri5nNMLi+mgQxcvtyy+fTF5kct8kfi
6fd4GyIXsyfEbGsP+rxfrKNFsKOcRYEcvb2Wmt8CLX0oVM83gPn0PzMWAe2s2h70
4ejKGa7fOGOq2ZpnRrbj/7wczk3DvKQan69Vkp9eqvJhJjnZq8SpGgkRg5FFnDnP
hth6gmO8goQnpiz5V6m6wowuDduOXI3x73y4lSTOQsXE6F38OMkdLg1bf6RoPopm
piXVP61/apaes2NtXvBXlG+tzlIM450/I0rptEYqWtDnUtPx9FWDXkX7n4v5ydAw
YrbxnaWhkp0T51MO/JkqtsA1RxmYbEwLM0qK2PIjMkQK1qvWdpdxeozgV4L2bYOq
Lv5WhoAfmV2SlS5pyLe/VbhMcsO4qe00RKI2P14lBBtouce5MevEiWtuqeCPn++Y
urKh2GcyF7YgFKNuxgNiufFcqOge8Y6TVl6ZPEXNkGwmtviABsGvZ4q42cPOXfNy
nrOOfP0WiC/sVXLjd506nBCprOd0LDLq3Uqpmeld1lkHfrBCKSyeVNEfsj5XHFYr
riLfsVBfIrsiqH1326tlByIOfFOXYMgRN5n3KiOBs7+2pdAQYKSYIj/NWiG0+9TQ
TiqMX03dGOmfy7DFrubyL+b/cvJFf2RoURHCSFNejx9yjKu2t5ACEYxUGcZH4XBg
9u/y1Mq5TVhJFF6vondxRkSdGLarp1n+JiD8DO2cpbIJGJByroEj7zxbDTW9fzYo
vv9JrADJWnD5yI+fTARcwptqWP37DbHb7ZB3p/zqzpFzob/y4c7TblxLRdkmGG1k
kGEZRwnd3T4oF6rHhunoHCLnM9OokF16Qiurj7KmEa1j3FKhCfL5Q5rvh4yb3dvk
6WPGq4pwdmJajDCBWEMrr/amk8X+R6QEuiyGwr3eMo6Dx+8sNmw8uZaJ512ban9x
qzxYvEBCE19abR36LxiTBDcoAPpkHEMgQxqZT8VdSVHpDGcwO0vpmArH+Z3p50JS
xatrrviDwFmbQZfQy+Rp+A==
`protect END_PROTECTED
