`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08Sd5LibV+V5hbbTeKsjw2nxEQx6as2MBj6+1XnX+lQsdFK/jdzFHtBwrMakBBuM
kQIdhFfgi/uWR9K0vUyqPoaynHzbZe+I4KBvz+lROuqjVBn3cUFVGRWAU6g8VTkR
zg3FeoVt/JkcMfHf0iGshT0WJZyd9rr+TeU25MvqY/Khqidq7cYmx65TguMKZic7
HQ/AoibuE5U7L9CEalEEchVH9Yhgo7S4WNCqUSHL4os9/wT8BenXO+4QhTpoEYyO
kZitzAMPH2pyehrBZv7BG0UOdVNjU0dgvVC+z6W8CNBKw1vV3zAiteWcI3qK6pVP
t3zCCcnRkgOL8AfILMgBjekB8NbvUsR+qPcRy/uGTeXhWKoQX/ds2Oj8AOAzDgPS
KciFv5e1k3ZIopzI79PMl5p7r2VOlXU9CG/cYN5+Vz3XPhjnCi1saPCwmeM8OOaK
z03p5Spwuzc3/5z1/+N3+8TLTAAfiT9RXD9/3MREWfKXDoWrw3LT3g2gLHPW5iL3
r48oaBXbPVYQBOx65Tc1yRuiUIb/t+E6x300nvhsYrgv1UY8yyMoemhbklaW1CWa
EE/KALC0QgF5/YsudtYzAMFSgp8/awvVh2CziOgEhXowWkFYrFK6As4HdpMDoCuY
+1Azu1W3mNRsC3ZzWMZHkdjccaqywowWsTUpQBP/To8CUphaw0pp8QfIdnZMHL4o
j/2H69Yb/jxlq5601aFDPj4mqJtR3GZZEkKxZmrpYDx/Fgci94P+PmorWBgqpkNV
CzqR4DTuX0Vdddy2sRsw5d8JR8ungfs6eIm9XIF3lADRtJABWL3SUUMnwMZAiDAt
kI/DQoBVG0KIdMJw1RD58lGHP07VHa4czhOdrXiFc2A3lJOjbqOtxIC3HKjNLWW4
Tu2+u4z/dTym5p2TiEHgleQhViorWhyuOnYupJGzPTZHBb0QwhMafpW18BeqBt88
/xgt/oR0VwJG1bD1Y/kOi3n2UJB18zw47rC77Jqr5wMQ+5mTOzQj/XHCUX4cjHhx
QMG7v7tJoE+LvG7RGp/0mJbyLe/rnD2+3cyZAtesdxvoXsYpFMur+flmZn3nXe2E
MNz4HODaZhWTZqdrzRoEGipGJGRUmcydX8QoUuO0F5fBeTD9RBNA7lC7B1ItZV5x
Wue2UTWdc4hi1Dests2HH+3wOkj8uTijdTmOjHIm3u9UCQPDRB8UciQjHotZ6nyx
WQhQpRswL5SI1YgCCIZJ8TAqkRW1gNrnWZqb8Gou+5884yF01nih6czaGtWXqb/L
Y3gNFEFdR9mn1GL4eskM8gpeBmEHs4BLEXQIZpjxxmOAq2dnoL6rQy6F55gc6Woh
n/yv5of2OynAHb00DUVX4JyGQNjx0skd13WPetV4i8z32XnQVAIi6lCXb4y2w0HP
QM240D306oBW8ucyWmw+HRi9GwJMuy2aLVVEYErQhAdNXYlALgyfWqK0fjkt7Bmp
ziPc9Z0NI3NnyB1bHeM4J84z2O/J1D5EZDk8Zd6pxJs=
`protect END_PROTECTED
