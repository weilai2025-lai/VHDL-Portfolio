`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrqxlMoEbRbLf3XV+rTGsfJYTDCJU+xSi06ObCU2K92CfU2e9AE/HJ4VnjcVGgDi
FxIgnPVk8SUGuOCaTMxfiJSCxHjtHcMPIxXEvjF+NVZvPLV+AFCQR6TNWGRlZkYt
mWPF9FbdAZ42WLQC9Lh6sG4F0T0W6Ym+KQh0rUVhSmRR7IlOWDliZyKiXXDXx9qb
zwTxr0w24VMXqtc7XHxf3B5XlOHRcqn+a5iT7OO9paMp1eP6XR8R9HGx1gAJpzAd
KiSpk1lwrrpXE6Mw0a3YQ0VlM84Q2DOxNaLyy2Uuf3P3sg4XsJs77TGqE2adG+cu
FqwcFgzxV/CVDX1rjK/Dd/+wzxftzarkvIbpVNJeoTM5ZFSw6vI83b4j1Rg6sy35
iAC0Xb+T6F6RY9u5w0V+Qgab3COmoRK/nwFBzQanJfMkcEmLetfgydeiaWxLjuNi
4b+5x1WL9hm7jLOHXReDTlOjsDbkpPkLMS4Saa3Nxv0Iu3+30xzaZom/j5DeKmm3
Ogu3MKFO25SxvRcaPRoT4RTpo6ufN+8GQ0jWBjmJ1HkalL8AbSN1gnoayGFLKBzB
Nh1qr84MX3sT/2RbdKrDYB5seS24FIdqY7b6/Bo8+MOSc9F/LwQ7R7E1xsP3BW3Y
L7oopcIGrICyB+J3/L23HinhKL1OuOzDkjehVB5RGn2y3C2WoM0c4Lh4Kf8Ghoe2
DzRV1NPsa79ailDeS6c54iGisq1UGDgsyZfXP0iCtq/igSl31UeTq4G5cRCUjdxP
rXHqmyOF/HXtUuk+uDLPt492U7yOc+0/fi6AGPQaJcdPpFoQIZA+bZYKgp4tcqjn
EQAEXSTBRd3fHKHLAYoXd77tazYUr6FNsiOCHDSGdjk0G7HLmUcVKcRb5M+9k/Ef
ptITSiASse7jogapcwhTx+o81/CzLCiaWyHM+L2h/MsJh29SCIsbhSsTebBTUk8I
wzS4f8A67wNm52roCYgfPh3Y2opiDoovnitjMmPlNT/ZNE6zOlLlu79luvx5eFma
kSdhpLafUGPErqnC4U6EEcl7kJ9/Hbp5GcW9Jiyu3ukq+dNqo9ngp0WOETwzVo+r
QuTfW9wrKk+hy8aITZt37f7mC9c7jnK/u/si815/xg1vIOYUU6JOkWLsSAtnK+ql
h0BLmo3EN4yGoUjG/TSaDrUrWlYRM8aDJWVcbKy044TzNhDFeGMkyqz+WTV+kxgo
g7eNgGUPUBixqm/mBx0HToD3N/n9zNMOCdu6FNeBJkRqTOuHMi3t5gVPP02AoiuH
Mq5VV1VvxjuaTjLzXyCb1sr7AF870MIJVFiGDbSdhsgz1Y5AFW17fBV8sWqXNeaY
GpHZO9wVlWNZSPA+w7EnuRwkw3/opE2lbKQ79pXTh/4=
`protect END_PROTECTED
