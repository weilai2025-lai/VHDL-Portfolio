`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFBZivLGj9v+D2lazwb7RAg5G/9vFSyAjYY4P7lKSDf/p+bOpO0xAxiHTMPj4vRz
HwaOUUW7hZhQ6yQxdUVd91JyqGQ9N7//K8aGmMCTWqQsD+eCf98Ytk9mWs08eMgM
N8mG/SCbPWVEYEn30AnyDbU81Vw0FK2hiRHgNTLbRQakGXOozBum4zssQkYXvqLd
TcYhlGnjBHemZ2VLdySHmdGZmKcd7rRWUcu0GQj4/nECOaF+wCtVfXAlQa1LLn1m
P0CO4lc3g4lo5pQhKMC637RZXNPiv7bKzs05/VUz/ouEcGRPdUaWYS00S2/6tKY3
O9wzglRUZoeQ+btz/Pk3z/FLwlknHRfBB2LToXDzBCXuZFKLOwcGmIAV50KDsX1m
Q1Jc3fgTLSEYeEkg90Z6vlAJ8LlgLKtjryD0hfN1u35PxIdg6XTNuJ/K1pPNODXo
3KsDH47LM7Q8F5XLijijgsYW4+PzCeFDEPqlI3B6vzCq4u+d88N5cH5CB9I9EKcZ
kxZ0Eh3g81Il8LyQ+BpyXkKatSKQcITbBqA3M1zR0pbdUp9lpeVklB69iVa4IBO+
Yyf402/zV/z7c1lQpsKrf0oSV/HhwAATAm8H1/GosU+Wea15DL1f6tSybGpNC5uK
mJEUrxE+WOrXvIm0paMbJT3Hu6HM+pQhE4g9sN5RhUi7JWyac8PSHuim6FDieJ9B
022iAhQlaulxod5FY2UTAHaclnvRokDYgsUzNOLomoygusuAQriyisOyC6FXoEuX
yQE5lEVzos+Pey1Kb0Kua6ylyFDHEEmbULYuY577AS2LalzbO/a+PNo6jSbnVtaz
Hyuews5RWxORSHS8dppHjgWpHYucJ5vCuj5oOwc73eTQPxxCF50fs2Q9wPRTbxwp
kFDP7Azx9/Mp03I59vUAbKlYP4UI7fxw/eMeS0R0Oodm6uCokDWEKt75aGB2idxj
E2Fb5GYVf0GTXpIOY9tGpOiPDvm3/CgyYmlPz3d0LwBQeoX0SR6SOuruuJe/nQc1
NLrVExlYYGC5OM3gcIrlTQWbqhpBU93anpGVIn/UxsBMYoN0ZIptVXFlcDP8l3ap
+F8HkRHgXftp2JJfPlBSxkzqcknp73RKkq2WKYv2BY4i/K17RQONocJc/HQlo6ha
Egd8vLpnCbdpUV4Wae6TUarBKWA7IQQa2SDa0lDOkcVZeXS0M6QIK7+RC6SwzZvU
KeWR3FDj/G63dlhGdMQnLUdcIHSAatIjxeitVgMQRtY5g6cOuelJaW9fhSnMivXg
TcJlFbFlDtdleGr6J8CRJl/APNxR0V/UjR+3mF89l+myEhp9TkHY65qlS90TfLwX
hbY3Pqdu+r7tvfocqZvr0m+7Gv3PqTiHtzRQjcvrufKGHnvwpBDEaKwwCVM7J3c2
uc9pGN0YFnmFiHlAVdSxOhcE8j+5a/DuBaPLjTkquA+7IovjfONNfcEJEAJOjaRc
5ucJmzwL2izE2gJfajaNIelEkMsFdRklnGXtTnB8thFmXaTDrGRYaeT80s6R3mkr
4rT0UxKFgqxL54qltJjYuaWJ2lS5qg+6gdDjjOYpjnuebuaUxA457WouUDhTENGi
4zitda23kO4QUA0PxOrxHcvl+Op5rMgochNU3d8bwwsD6zmutm+8CokCs3LI5gPj
UekvZBVlkxodgkkrQf96XvUlapVkDpg5p1HYQl+UnH3MxGFCDV+QIcHVNL3Ns+we
jkFlRrJkKiq91bQIamXp+S7gwjSymeVdXMBNPOUYXJU1FAPJP3mvv/+woQ/Y8mOE
TpdYCxaUOQNeVFKuhhfNz7iBviYmTqzpiiB+ZXITiFKheq4NMLrA1UaBt2Vq3sg2
Xnd9kq+POJL1IXohLnVGYocQHVI1M80cnh7NZElVavFLESXB9p3N/jidlGW3+fIn
f1IZClnYMj3pI8xyk7pB7xgEC6e4x74Sp4PW+hzzq/+pY7Ojah6dIbHyxFPHOK/q
4h5L7RntgXTFh2bNR1OO5H/JJM4qWDCYeMGE82OcSkCVVu2QsW43mfg3vADr2c4Z
n+OBpfok3mBnzGL9CIsB81flTtxDVZ9xzEd3IixFYIR5vMH2hri/c0wR0Sd0UiIy
H2AJEysg0PRcTENhH/UiP9F6og4eyBAAPJNUPITDlBY4Hbfy2wPZt6ll1i+S98kw
zSM1q+GyNFgYy0uLfmcPsAU8ksKHNjGajxHb9wynVAzse1wxMAtpkjlG54zoTqZv
aZP96Yg8mDSXWvSXTYFhkyVKFU/7no49g/yABWVS4AUYGGAvx0uot9kwycZHeR0V
u526Ql8qEe9WKuPy8dBEWplXCKmEHjkHz15zKJ9LF8KUJlmy5XOi07/ArCJaT+A3
Jhx6auDPeYBFymVmZz+QbDygt2Gk3PQ+LNPkpoB6BQrY2a5sYhEzLk9mq+JEkb+D
BSJeJKEKY0AIF0PhW2by0ng4AFRVS1+N0suHDps4NgAyKyQYLhHXFWnyfZg07EMX
8AKk6g3yY5U/VPGDnK2Nh8Em9GlI3VS66817ikhf0Exn1inipzVftZq8JBZ2WcMZ
yIZXtAgEVfOhB3Rygw4kNdt8ao8fJIIxt/vD0xO9xFgcvg/CHqoU7ISDAgn5HtWX
5ZaldU1zVH3iBwUpUiigiUzApz4sNN83L+qnafVzgwT5jwK2sZ/xAjAJp9vPjh+X
O9c0nRfSWF015GgFXQ4DZkI8D9qwrshDubnH3hSj9gireH/oJewe3otFvr0kArfw
xLHptT6NasNmNCyhnKEhecwNkhcaNguic/vg1qnR6PxnG3pg6ErC96sryCsqqe3G
dklxTkhM0ZY19/bpqTzUUizwitUPiXZdqdydeGdCE4JACoTuUW+sL1R9iK0Ot6eK
/Y0MPqZKOo/XnTxOwW6bHYFvFDYpdmHp3ewNrLAyoiooQDtGmYLfy9Kl8diEJ7fW
UExwYXUp3hYL99lJ69sNLGgQifGT0Clq/YF7sfHAQ4v8K+actz0gNs6O6f5fgibN
oZAUf7RMHlaCvxmJTz8eIQVDxgAhXrS41vDB1MU4hZVPrXR5Vg5jKJSBRYPnp0mN
0w8GT+h2xRE2mZfPFBRB+SKgUi+fvH2xqQp5YKsY1X/UeyaKupc5BkSkNhmwshnZ
AVVMJgxPWTwaWIlFBZWaxl6bessMraWTT12JGo4qsNQWK1Z5k4rZgIHPFJM8lMx6
lPfKaTWiMRytixDpQEzq7s+oaaFADB03FXi2aUkaM5juYcDdFSmqd+JOYQDQ6YEZ
oX2uYz1Fnlfazyklub58pRktOmhLmA4lnY3zhmMHUzuO11RfNWCwxQsz1v00CQjL
AxOVBno7uQnIOqNbX1dP0ZtO8Xz/vlcYcR84Jqlz0VUc+QxUj/HIYKt76SGEw/o5
esMu4uVwhajH6Et29/GjRvYMUV0Ukok6W0cEgUYLHmVcBnfzsANHzofoVVLeZLvd
Z2sWjUu/7r//b2UvnzNJO7MPuj6w0WLZnT/VIO2CqNbic8/XEd6V73ct5FrH9DDj
vjziiCKQ6NRO6cUTVZu9J016k2YqXgLjALS2crCUIVedqvMossEhyuktEcZL2yg/
uR6yd6LEenJl/GaEcjdVLYwS67/sL81tLNiH57rIR9lA1r+doqurlriR4+7Czcjo
jnxtX0VTCPzF5CdfF0+x4+uaG1g/hHxvFe4AI36ixXGd8H6zHUFiAdvq+13HRYgi
SlN87EgZiPvZqv7XbvPFqmRjRXTdZ8/3D7LJz7mQ8+fclgAlyPEN5KKR85lCQnFA
CKHwjocHqJgRO/L5Nbhz5hRkSYCpG72fW5htjWcmfyN1uJ485+cEupmupRH5PKrt
nW0+OsqVAZpuyu3IYsIjVAFzLS/GSFoxiGIg8JWbxLZCXbVnyQxFUHbVULF60Rd0
tQYjyAmN3VNORR+65Y4azYXcygD868QZAyovXVNQN6BThsrcRuXb/o7DJCmlpQEu
CuR41v4JjMURzw/10X2YJcyZNmGWVECLAEzIQXlYNKhfFuEyWTO6r+ud6a3C2oDm
KTUEdW0j3eTaVzUcErXzSLxOhf6s5gkeiG8WKNZvqIo2PXMiA9X4Ox3DgAcHdr4T
I4yQaWMb+Q8YcG2OWS4FnLRebIqa9WPhpKr433bzABXPTXZdoqAeZmcMku/MCDpR
vRy925ym5t09BaU+43IG0ncvxiXHg3+/m8v5z8yVPR3uDNNGwN+NQ67K/5eZ6Mcj
VRNC9yRPr+6TL1zuImFF15985dTFI7i3qrMcbW9gvXpeWn4u9wcjUXEQXPV96bqM
Rjzm9tAAmf6v+SS6s6ZIOq1BM4AtRpltJrvJJ6O+cnaB9FfyOTGnEV3wR5J2sfCx
fp1y4FxPxnbLBmFQTI03uhkxMUr5KsKzD1uoxUzap3zdUGi5CSJX7nk+0a4JhQl8
/aAEHoQ+OfNct9SCOxzA3JveIGiLiwiP/WWknIiGkhIUdvFdGPNlHkvJO8/qbIP5
SesfoZ6UD3yOp/emxYDC8tQ6OCAo8eQwOGKD6oTiWddITW37axyJf169CF5+TcuR
Ci60ANmM4lSqEMRQrKVNHmWEvirCkNz332tfln3W1FsXiBd9aDPdw3RdFsGrmuV6
vlv/V3IqDZjXZJD00sJgNMAIMTtN5sgtTKGr9/bBVOEUQPqNHhbXE/+VTKU+7jIU
drRB/BkyBgnmqdrrcU7z3Rf8Ud/Yfj67qGCBvthIu9jCcwQZ4C7OInemOLWvBGXK
132UL1Usuh/XBaQIeIA55T5Kz2XxNWO/UfL0HLI0sR5mU2GnsGDrUVKoJHTdl7de
18xDpZm14xhusOmX9rGcSEz6TZ9+EKgWbb3cUlMfylGQVGckAA6wMjOxi/PJpDf6
yR5lbaxyJjKER7wV6lGZVIOXrqnvzHSpgNcD9LVNmK74jCdd3vpGm6IOK3IPuv55
cxjsM1NxG7xwmT8oLul0jr1wKYROF1/3XvnyNeWOgbc=
`protect END_PROTECTED
