`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmSL6xzlxbi9Vy9mRwXZktxIOaG5uFWSfXOO8l29OMELkR46NgqojfEXjuCYKQc4
+Yh+0pwUpfih8cH8rtd6wJP3HhtXlVdS53DxgWb4TledPqaWyO9QXSZpYlb3mNPy
ILf5uOz/32neVw4a57hyvIWMz39KARv8o4mthXMuvKtGxN9IAkuL7MZGqU8MFl3t
ZzWjSXdl668xPBbnOjV/DOZlrtA9g4lS9yVev6bdZvK955ikk3M2Pw4OSrnbdX/e
tIzs/QCqXY8JbZCFi5P4xRZnMzLt0WdG2vgXcWwPEvs/gXX4iR0iqlwO+Y41Wzp/
rPNDMcPL4ynBL2HFZg2pvB2nGOt4vUqYnYtAQA5BFf2J86LsYTfQVgom4RiADE6z
FXaXOgoiW2lr2rjwFXO2pmFQEstpXMFznz6ckY7B4I0csozHqWowfGUuhoJaP+Qt
bQGIIIqYWlG8F9cR9e0uEKIooJWbFCiAVlNv+JbGfgLdeB1dvSNMQlwp/fcxE8J3
DI/bYxDEQNwMZYuuH9Ux8SKDaRDdFbWhJOWwl1KLO27C5lxteDomUA6iXqmZZuZx
dynEx2C+tEFKSA1bt+SH1/IhSSRT2SJeYlZ9X9Xx52VR7U7UdzNnX5YW/u+V40SD
va3PELMwQceqUQl5dFajNbBDZiVLfjYm0f1TOpt9wE0hbKVyiPVfVgyl2LErQVIt
N+/rjBpEhJx5jx5jUh3DZwBMNmt3MEmGUU9h5Sp3XUFo95To5kyV/QBV1y5YWQaO
HM5qeEaqkE34XpENkOawIu3PTslmww5lA4wwD4iAK0wqBXawFP4RjC07PqBk5g47
I2AA30eMk4mGkQcIFnKD9QSK5bGTtCd0AFxyz7+bA7DzmcmQDEpWvp74/vYx+fh5
QAMNhhBSujEWjvI/SPFkNcrHLwiZFWKKe7CBBih76FAgWggbuQpi3H8v1zfkV/bs
9j/N+vxt1fJTGax9b73bDmDF0qjKmEjLI94Ez4L4qmipeSwMrjeb+errONsliORa
ZnevGHvYd0Jx64rlU9maF++IYcUgEh7nk9QEw+p/9y61R6DGWWSrHXMV4fQyZxA+
C06VIBVNJSz+0Yn7TJXK9n44kA51/s14p/qRu87skLc=
`protect END_PROTECTED
