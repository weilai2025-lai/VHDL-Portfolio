`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOEOawHpkCQB9Ncjy0CsgRjUR2g1HoP70wJfnC4OpYuDa18zV/vSGSvTRm3JiE++
wdZKk7SBKcxY6+V0FYwv69xpaRCuGYRNUoR2m9EaOO2w1wUb3Aj8mnuXHgklF2Ty
NoDYCPCPcZncqgygZsJqvB/gmrcknGrB+ruIRBxu+ggQugxXWNx9ytMUC8CfcbQM
EyxnC3WlwdyuIMCUsfzjytFyIJKsGa5SrIa0WoOXErZNZMH1+7mzebNrigdN9Opg
qOSyEZGmoR9XkkYq2IhSnlDRUh71xP+kuBcCVYANl0fjyjw52J5OZDyLaKkUCtg2
wjJuXGBTBRUtq/qrvcAulhmCuX85zpWN/XTBeyBTnf1IgZXIF/2whyrOv0CrJgfR
bjxCtsa56GxsNqGcUDIwRv4DOB7EVGEkA8M4/GxYqo2ebDD/kzvZY69ebXjo8Qa7
BT+WHgaJBLTpqMk7tL32CAjqjez281cFGDHgojpcZslzFF6Qc+RDqloOnNnypeHw
ZaXpeVg+OmuUhsS/yFK9ak0b2t9Lgdtq38WBdZrUZYB2Ci58XtKQe2CfFu9OytlT
SEsXCxyydkoccz9EFh6MvEivJAUOot6jik3cNUkvDMb+pGkOH4IqpV+al0bket4K
CsgVkMsCDxiniUOYUSZt0t3I7t4H1GeXDIf/WZu7vL612W1uEoz3bFA2ncrg2gwr
ucOHDPNi070Wgdz0jKMeNdfaMfJqYxv2XEdaBwE0f+OfH1BgRMireL7t5+jvZDW9
2e4o7MBN9SfcwxDcKSTJkhDLmlc+Ma5Vhp6Tw4lduljdFeipbNBK56/2AWeaV2ld
XmFHvpAwojrelJIhfz+OR8JoHU/Pmk1Z+nQPPt1zm8Il8rSGgNiQxMhvpWTgXVJS
5v7coWMP/mLHA94U0eOa9vMLSyjRomcB9Co4WN/NDizbBj8r1WQ2gyJtQkFX9F8F
4InWhdV+mTnrUDPhmojMUq00t7E8Mlxqs/w3clUllzWqdVWnhtqnF7IEuTsI8MvL
546mszaKCX6H81clY7BTFOjr3qf6EFkyGXkpeHQDENxpwW2PgqyarTnuTq629582
`protect END_PROTECTED
