`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jNij+LqTWX6Ig/Ldd++bDwTGKoQdquNb6Q4NG7b0XeN5oa/PPVyb8ESK/pb28tgS
bbo42WgyNTaZUVxrw0ATjlTNetjWg9YsaENYOleAqnKo7VtcLa6Hk8tvfkHbuU9Y
ky7WBETfnHz7iS2vbe5Vd9tLc+Zr+irN1kbGe/doT/or5K8GN8cDOp15UJbrhYk+
LIqRcDr4DTTJm/eDWIpsI7YJA4qnI4lAU8p9zSEWC42GAUEPaKJ91xMX+uh1XcCd
28KmEB9Rgrz0CDDDqxoyj3grAihmVLmxM3iJoxznS5EwsSk8O7Ln+jaMJRA/yOYM
WRLE2CSDUqDDoCMNNcyBfDZIU457wcE64Vh2+LDBFCy5VD6nJ1vC6KGUH4ioESWm
wRyH9EuKANIZwd5/NYoBDNN632DKyRTlqnFJcqCRTMYQW6iWkutvLZ34Khc4U1AU
QhMfJ1BftOKLJqf99LboanW1uQZ474EVSS+GMI5v5nI/ViW1xWKwfROj7sionSk5
2BLRmHVBYv31HVivv4W5zU66JxT0F8jd4wKdQHIygm4FAj0+UegzeBDvVhKJEQmm
fX2o6CKFfdf1jzLf//3lsjhMycM5a4tzEtdgBb8AYq7gTziYbdocomr6ro54NOmZ
nofok8h8g5hgruETLRoCPxhi166s/aDGhIRLfmbAqWT7TaDyzap257w6YZlnYVCq
o+EvlZlmqgCmgiLqH0aJz84+Qrj/o8lcEuv3h3EbSYHak0uoqlz27KV01OF8zF3S
ZxLuoKbbVIL6E7JAu6QFFFRNfcv2j5iBBplTXd6YvRbyNFFG7IN6zC/WskgqOd3L
5WM8LQO/SVwInDXj550oxtTcCWvAXzGrXYMCtkzHB3slPReV9Mu8vRVFCxZ8spcz
TzLdNOJJbM025fe+sYFZYVzNEUyka/lKkgMhs2+lsSZm6Hr+BBmVyr3RNd7Q8qqz
CGrXmVIyj3F8cuAcisSocfs6+Nq8J/TJ8ayHr/VUoOLPET/OLe+kANphwT7Yd+qf
dq1dZOAfQPT/dlPc6OW5K09JP5ng3oNtO9mNI+PixEHlc19WV2VCupYP2s/BlRze
4hRpOTs4BtuKkCxb+1Icq+7gIMrY3DHF6LMjTlfMc5Ew2rnNZtOYjokPiy859HeH
2L8nEbAWyex/EzWvIYE61zRCWySoNMarAvGXOQFUdHe8JNEii50reupGs8TCDQtU
zL1MKyHAfErE7DbuXGtd+ZpfG1dvTFwmDN+baHLdLE2AFt3uRQi/UoR7ms9MZNtM
ZwxZS0T6Yj2c9sQgrX0HCeCx+zfv8PtiGdmdG/JsB77HXSoUPvOpFQ4sFMEl5OTp
fGrpCXxgx0UCMBH11Ac4YgwlQNTCikhnqylHHDBGVWdn1PcrKHPK+g3/dZ4/oYfo
HNdjCexsxuvsAZIjNHPlx8s5zc91VeV1/djw4tPfEuOfYQhH7JNE6UkhBzLz+hYf
4LKHorb6w72aKYXdF3yBbkYQkfBeeCDAJgxwOWRNZTnf4WQPVUmPkaUbp4zEIzEd
d1FKkC02pVJb29jMP+p+NDy7mVHZw4PLy2jWxMRdi2FW6KDl4VvyiTorYjGsfFo2
ozl5Enl6g9C3YxhCzSiPbwYUvVLkq8ywFJdsaDbL4JHslfIz2Ey7pjkLTBIYXCcA
U00BaqNDsbmlpnkxzyKTkghHSf/gVQ7F6EW7p8o2kbkgCJORAFOr4okFO0KxBXtB
Ge4D9YjabnnMh2TaJIAkKYxvYu/BYpnvhdOuW+8Lf/bfs4YbovbCeha5AjdvXioI
/PAF7ZT21PTrsCZRXjU9I/QPpZOkkCy85FSL2u17RlE1jb9rdZ2EdBaXjb8adt1d
cOzVjoz8HV+B77vJnQN0gUKpdKXguWK43T75utFapSmF4ZHpXMN2i4sFRa4yrNOM
FokUWwxvkXrvIWGqcli4a5fY6G9usIvIc/eEpZn1AE7sRPI3Gel2B0A5atZD5ZQi
reMvdxoJE7Jz5umQOLSq1zUiaSYywM5Zu9/i6jg+dX0kOvIhmxxInT9HamJ9orkl
TyupWPU3P1QFk6Fm3E87UXB0dMQ5nZebV3M9nE0lURjPjhNqbv4euUlKBe3yY8nt
ZodAit7cyjrXigof4Rec8ajxi+B8zTwh2yPkRosO+1G/e4zABlwrcD4AaT3VLMbW
kwV/y/WBccmcnsXLvcm7K6picSIPhoiPHWXUQhNE7mjdMXrG286OarZwZ0so9z97
wOiwgq304Cv5r7l2F7p6RqyvX+w25Cw8Go8+gFCbRbQ0JTwVpwnra+VK0CPRlzAA
KSfxnA63Em08xg9gAjv7QQLHLZokAhH3jDQ1nkq1pDVqBHYyREgdWpTZoFX+sFCE
8fgewoiJXGiScFyuVzp4MGIy/XakktbjP2L/LzDlFGjn/Wqo6rl5cRg3XxvqsTaO
FbSp34mFhhKGAwJ3XWQUjHAddWajg6AdAi0A35nmPASacM+0zT7TnKR6Ei74rlAy
THrbn4iKuB54T2b0vrT5w1NWoqf3K5KQRFZVQDYeovKBeV6mqZ+a/Czp356cYlP4
tgTzUIInVyYS7/L64faDrgsrTNQpYObUOWL0U+JEdecwjk7jX8yXmDRUygv6pTRP
aIJ70VqQWrA6Ydjew2qszsKVDKA2vr5MGesxRQwm4IiYbF1qgAmsKP4OSdgILMCj
rg88ero6qpR5CBhCaaBTdKFSmP2Le0FTBFBbS1TYeWGKIkEtmY+2e/x/GUp9RrYv
UI0UhWc9KeFxKaXPNkl07sAu3A4zBaKoI35SYaygcimgx7T3hBpdWrLFyWIPuEjM
dEfiepDwIa5MAQnLTsLZMSE1Qe5DE35COwtmCI6dbnJpv5n+hhZ3WPOMnlmaYRw4
XT+MpVijIteAFMViejm79yDTDv9VtIkloM4iomQdprELnMK+txGFQscs0SZLdy0v
6RzLyn8wb6ezvww7/3MrSQrGdJ5x24zkCMGANkNo3Mr/ca+6h+g/4cs3sahWG79m
vTsKKt+/SadUdpQkaJfulRjte1yl3tEnW+ALyYzpnVO3/ywQhEHgbWUSIJvHE6Dj
3e4b7/vaSqy8LtDVlupdVm4wGh7YNcFSUyZVpoSvvooyijSheyO/ypqkXXrNS6k5
yxpu8qLpE5cFD/JXLsy+ozP0qUbEArmvUgSGaBlsNAg9hyzLk4iLQIKBmdysOhNP
jG6gS01iu6UVTfjcnMmYZKQk6W9pYsw3ot0Teu6ZCUJnv83JvOFpegS8Mw7VTmX7
O87ypuf/dljem1tD2CTJzBHkqgz4SWnVmxTlECPKFSMCz0dRZ5D9cXEgpsbmsqU+
GbmvCIgtE3XHZ9eCh2nJ0QizsT6z3eYYABUtzarm6pUpfialkWiARE0ZHAa/MVs2
poQzARjLNNdr/My9PKNlAl2QvcHYziJ1YG/6/g1kydOLFUPIS6Qd9+QfrpAV7k7T
sPAX6LOnqSDyfvopgyEMkft0jVlMeZRKrCq8eTPPmS01ap/6+j7nLnooZMPi9a+r
DMqEpZ8BFdDI1VT5VQAfZvFQGdi1UwralzB+WN8VlpZM9D+lzdJNuj+X2mV00KXf
PM5JHVyOnvX9mov5mtgjMn815Cna7D9Ma8tsSWP0byEP8PjpE6f+uTMoJDy5itKI
Hy5ismDRq3KNOfsDmObapcquIPjbEL70hQKPRLGMF/2dhLlQOWEFrlm/9gp0WqZl
TdogVo7W8YnmNRpwln4Lwd5+6hdNbCwhNe97oCFoSPPvjbyOCy5mulubHKzLnqD/
MJUsueyYKPiE+7JkYnv8nheIDeC5gvjItvMDfwCpaYjm0T5KUvFKTbonIHz8sFNo
y9zoMLA+kAqcgKml+orlKLeDzJF7yVqyqYWHtZNQa6HuYXJYsUG59KckMWQcZxVJ
hve9E1JZPy0GfhilqQMckZ+WzlAiPCtD0rXc2bLMa1P80nj+1cDhOzIJkO2g+pog
/T2StMzKmDVnx7q3A3004CZL4cqUCPKOEs5Oj7Zz1bq4vflKKYDrzxDLT9Yd8RAt
Iox3V7FSGQM48Km8bf9fhDFdmaCmzIv2M8J37Xee/nRwRyyGw9TPYxBZnjLtb4Co
NuvyZ8jfSHuUg/jDu7XQduiQydQahyaYIIU92Eo8z4zLp/9O5n9Ye1UgaSgJVrPP
ki8YuP1fMvzEIlG1MQ4Ma05mk6uphXT1qZT0LXrVV5bFakDPig+4ncRB5s1ZVp37
337r4c7r7i+fskiYCx1RiTtN8ZUULTnJ99k+RneOWk/7RS+eGx1/gSroWvTSietN
gFBavUx1paIB+YZvxmP5d9cs3yROemhyyJt9Z759Lrx8e8/250Xx/zf8seaenpA1
4QTkKvXtGcrqrdjWsifSd2RpAh+JjBK9hmIPxESb/0te7Bmt904mPoz86MxGgMq2
IydkCfyfl4tktHL2Qs29FCTUmRkaJtZad2Xd7sQ6PNTbIxnassEdhLz/1fm2lgHB
WjH8WycX/w1e2ziq+30V7dtYb2muSOKqxZPMIqxKhv2MWDRuTifrDzhqE2EB1tlh
2KAcpfV8gEm08MUQ05aFO/fMHHPuVxlMzinbqNtM9VWXLBuNI1rz+s3NrXeddw+T
yY2ObhY1H2wMQvRVocckYLtunJ/cyAXN7MuzboKoVd5jlkkMlTC6KfVRkYBI7dyW
NNtbVt1pE4LCjREAdG3m0rn5n0nSfxWhzchOQGHoKO0oJE/yMtex/KFVnsVEb5rd
D2kiNYQMijr4sWvdPVbRbe9nZxvvPYz6t0vxwODGoaTtfWwcaNNiWCA84VlAEdYx
JTrD4IFM4UCKPolf6fY0xC6IAaRoiwe5KMEb0Gn73Jo2zKMGc77DAu2dvio7zerf
LseiNw38mIXu6o2GTmAObAA2LeIcvDsxs/sFR+DEToceI8i+22kejw2CzVxJRUzT
rCgEMrvWJTkZ+sHp8FALIrqu648kaEJ0WV6MyM1/p4Kmg+Kn6pXfAVQGNvhZ7/lD
FmkGiM7N8hOyu+5WU51P1vBplwKlY0JpvGM8dPN63cbzOia4qMJysR6BcSAr85n+
4FVYjFVpvQ5vHHlndSpWHImIPy85LHApNYfvDkxgx8dYugjBFst9nyj09vQuKmzq
peqooKIPiGtvFBd9CveF1Me6heEwMACGhC9qY/8W1J1m0v6B9scDskExgoSKZwoc
P9hv7dOL77ciCss5HaeO2/OezysOeIZbRJ06xbyAF7u0kxzHE+LmBkszrVFtcTaS
2JuOdpOaImERsoxWOIGq9nNM4bUAmzQZ2+xXxugmpz8NSaOYE6F+UPAPmSN4z8rt
x4+/TxDxYd20Dv3tSLa7QDuIXR8RgQf1UvCjpppNoYpInVFLxSTnH+4MyfaUC2C1
C0bsmxzsjb2X4hLM18U3/8cqdafTcASZEqXxk2/T/go83/+iQO7m1gSXp6mUZpNa
BclKDyXpDvtNTjtGqE4vlExCF8JrjgeX3WHMMlpnMtVztvTm3S+HF8A0P4+BeY0A
AmB8rtJIHO9HhVscdhLnXDqR1RfG36wH5mz1ZpQP0/9BgRxas4tw8b4kOEICKynK
he4JZr3bsAYrOqcPtKXYAjsFPwu6SXY4eAn9l4aM4RW6/PzIWPwgeC3IciN3YpR7
l/yJUfBkZJuYzygpgMhaHPXhzhoWPRxGkz/KPLfFPXGr20OhtcC4/b02whSf7Lx8
/GzyPISi4c3IrNCKffDbtfbNK4bakfQI+QwoqY+bTX+P9TA10V1v7wYr7ieVlZOm
RQDEkL36ZHnTeuQ6SaaFcMNrLuI5+Jcb9KY5PplwQ5I7RL+6N7Yc3uy4uObxawne
2/r9De5QP8neVBfjGP8Jr+c9vZzlNfFYrLjJmyq1IFEmILtS9yUtHHbRRr15WCH+
3xK73pzLWETw9DmR9i4EvMr4EzA3R/bX92ch7HtEL76JrOUcdj+aH7zT68Mxhdjk
hI3TxuY/R8IWSFiITmS2HUE0bqEERO8B2ea7ylJbBF82l8ArcOweB/G/z7+je6X5
GwKTmF5VL+sLI5XkFBLXfPF+LrZiWB/sGGbhmrSRceaiaCnzXsOhy/GBcKMuCKFe
MW2MR2k0LftI5t7zTUQvncF713a1EhIwHgTP9DydN2lq4bt21B2Z31N5CELLL0Zu
g7YKvdkkgc6V/35of86MVHk+Gp6VmXBPyWv0EKFMxsBRHKqKoDzspou9TBkqUhbt
ojIfkqCZGzkbNov3wOEsx/N9+b75B2qQ2xLq4MVppC25fkRkbSEQwrRh/lUEl+kH
+hGkAUnjjOzNQjhvQZiMIQI+CdMdVDRz6HP0gOFBOPRYyqT93srh9yqNXOjbJYbn
9Vzpn849DqmsKspDLYFgBZkfPzbDQQ/rN8xtBZTzAuMBd+jJY2t4wEeWtRKfUkBY
3npkxCfiyUo5ERggBmPWBTAvv+WpQ0tMSoo1uQ8+QsYt65Ye5td2c9rQYohR1ily
ufbCOMRUhijui+vYGMhucnqLDUVH1UEkn50AYJJJttPmCFSDOL+E3urZ/T39kjEv
XMmrhackPKCTvVklRkhELl3CyoooibwYl0zxbVFe22yMRhB63nbePKTq588nObAF
aC1KvMQhDhlH0qJ9FzNp+HR+fe78DmjSZMSsJOxXur5Njv+Kzfit8Ff772tHVncq
9kIBosmsIS16xk9Il03GB99xqKHQ9i+JsZFQwGZVEGz07Nx1vkcrYzVzgdeehE1u
2XxLFsnGHHiljCGqptsgXXb/+uWf8lHvvcQxjywxKQYVoKsHMIlCQQUtdSHzNST9
d6Dc1lcvKJOJ/kS2M4o2hF2gcu5A2aeanOuzrRmpFioEQCxHC42OEuHCM9Zc26vt
COwyrnX6xavKv2ljGc+QQ4csLQYf1NPHIZqJzDaAZJu6yRqgTOmIsvDfIwTv3Cx3
ryDQOBJcShcP9hnfKOygpuHrYjaD8EPuOPQJcrSe7WUvCAIHQgUa/cTHbbJh0MV+
`protect END_PROTECTED
