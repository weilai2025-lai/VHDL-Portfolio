`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWoNIJ1RTeZ4jE53W9j4U2PCJ01XyioYXzU4QIHywhy2cQyEZsv0+4KPAMFs5y3L
P0ZPeejoiDe/Fk5KuFnv+v4NB1DGy1wrhfkDPZiXG1e3ac985LqETb7lByN92Csl
gj1Gy4m3XbKdh/mWERwvJq2ecNbEOg23nchAw8VvtmJWoHB2C23zgXz7GB5sHXcc
I+3Om/N5OfbCfNrB0b0NZckXxd8Zn3FNtQrAjbpXuo9NxL5bYGUUhjW2pYMV7aCW
AEGF9od902xK4if1kTbDzgFv3kGP3JmaIFJhSVAvJXtIIgEi/k9HQMfPvUA3Q7Y7
c8M8yRNRmpJFsdymdpUw54nJua7T08JNcuufZSxuC6b/f7qIm8SEyeeVwO8FAm0q
wS0hYp4RH75EO8nvK+nNRJ0C0eMrK3HclEzdQDM6nRhauhzGXqkE0drhp6bTSrs+
x8lyrTjzE7UcDQOl4Dqa2o2vwJveir2NJ14j9N8f2GrnKnyiGdksyjsESKOQz3SP
neQo+FbXOkkhR99uUwp0ET5O1Clknn48mCMmZzNE4XEckOLQiQtpJZ+59DY7JSS2
VddGzg0KCdMGsq4PEf8A20UKpUB6LFhvw/15JEO7vGVI2PqkpFFpIwb3rtxdQYIG
Bs+i3L5TiB81oKJTKSpUam/v0IhlIBOWt3tCDEcoQcPMEzuzirNhDTkhyjk9n4BJ
SgxVZ7YWYU4+bEcf618ppIWh4f1p/3/Jvd2PBLm+M12c8g2krSmtqRN5v80FGk7k
AtGLatf0QmeVRKLJSPl2WxjGsstDthwHc8tC1ECYYibmidKNEjhW3yByx7TSnpW2
K/cgWaXAB6RxMnv50SxCtKbMGTCTssUhv5uVHNolHk6O+xLcW/NYjeMSy7GgU1sw
fRu5jmDw8hTTQoXhsw51V8p41Lpvo9XA+cbRJWJ218nlCrTvrFnhp+j6eOi5+7Zm
7iyW1wDASovoYGN7QcWcUOkGf6M4rXFYZujPeRWnQDC0w4RPdec8Lwz7/6f4AFOc
ppQtMR0hc63o+N/WYkUm36m1AocWlyTMptPdKvndmxK02gxUPNCN4WiwKPue20BE
6p2dj92j+Dhw24I84kf3EGNYbDT0c10sm9rxNreyoxhWWNXhcT4AK8tcf5OQy7xD
zJ2tcXqZz4zQ16Kqr1iP/DPXo7gE7XIk0bvNoYWoHJ0e6prVP0tXJR80OTbrFWUr
yznWMJuJJuLP3iLJuhGhLidFObGXOiHCEPTl65WLspUreHRDPPMx5DsRkDVnYQq9
`protect END_PROTECTED
