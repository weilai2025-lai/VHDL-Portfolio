`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YWzlUUZ9pa993HxHHLOzAkMnhZ/xDJPHxglzX7K6Jon+MCBu3Vv6QMzsIKB4QKz
nmDjFObCWAGc+FNXV6CmxC7zW44dMb0PrZjBqsFTrYyXiF8dAyAs1gNeVAQevTjo
+XTvrNOUlBlvWQJ27UiXZEDNWl5LBZsfRtBL1P4+Hz30Ek+dk8GN5Bj2Sar121JI
58mMQmCeqB42eiUZ8nHlAp1+msOHceQO5hfZLihCdLr1F6a4HYwWZUXPHqKC4mRC
hzE3hWJxtbR/JUYJbMCUvZwmQGLPu4hkjz0sYT7uhW6AMZkpMxCODuqwcn8BXHQP
FMYVx00iDRcrZ2qPqVlbhL8UoNX2reENN+xVl854MftH7w+NdCs2Z8jSxdgb2wQv
rJfngV3bcPoSxn5z87E9jJdwmuL5M9Swz/gFRbZfLirU47pn3M1PCBu9+gL7fekN
AQ6XSELFrDB6j85SnBjBmNVdA0vOGdaoFAhkZ7r7eOi8LdQpSeJ6ui5BfXyowsnl
/HiVv/DuZ69iIh3lX6z3GlpnDwjpphFxD0qy1fRlwi5dsGKXHtdnLpSJGHggL529
YIZsT0B69wCFF6+FgREWvzkfG2kbdq1ofHQj1SYYy8o6y7f2D4srHo4fFip/ds+5
qrycalqW9Gx21qsK6PeEBHzcdzurReA2/J+nXn2KphEhgzf69qS6iwRIObYpntuO
ByAS1LJCPnr7s+QL1GCKd9ElW3MSFDGBMSXzF/x8L6rX75gPmwfMqfyXxRXGjCw8
bIsM+tN+BBr5MhbcNw4CXvcwFT2fBZjUaSb3x5uIeIKuV/7JW4ZxGT6kpw+GUoKK
03h6ZFLW0jjILZByJkQhfHMakjKrvesrdELOgy/y9T5upjQREz/IN+9Xo0+wkPp0
qzWEvlnPp+WLpIq23ekC9b9qjTjqM02R0RcAkbKvbMk65vBk2H52DiND1p7q9Ahk
MrKqcz11tT5FBe52rZ5WR5wfsoWfVy8IUnX+UAK+o7SK1lER9GyiKPKXykHm95nV
STr1Pi9K9efo4n015q6cyC0rAWDjRrQGCsv697GUhIu5QO6nsUJRh3qp27/c0lkr
bvJq8gYDHbIwcjcUasaqqN7JIO63+8X3k3uSs7NI5eSmd9w8KJRgXX7188fkO195
`protect END_PROTECTED
