`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6tS4qp6z8Ld4CEbipBlF5va18xKSIVxgs/2vwhUDLMv09lDQnQ6925CpOL40G1e
OCN/uT0H0aOoksS+6bK0YfF1J07vNKVkw6JTbppmWh37dC+/NBhCISaWxUG4Q2os
Bm635rmFubnEDrZUk4ivi1zQ7kX7TpKxe3Mti5Xuy3aq1+uIux3k52kqZJ2y2bJ3
j8WQ5ULH2yg/I5CEudqWGcJo814Uo7c5NFPhWeQZC5sEnNWE3u1yupY+IMiDStk9
g0vGMwxezDpNlxOW8tC422hNpZWX4vc3U0zBwViFbuQs6W37Jq9AzxfYV2QNdtuE
yp/a1m1J8lEYb+Ym4H/1UsZ7otDDHu1viXDvRh24cyi8fsencVRAWNA8xuVgrqCK
xS2AtwOSZBnr+h+SPZiQ71k0RM2DrV8cWwbxR46ijl2i3alAuOA2NfZEH91tqOwX
3rm9mkfbIYXBs2OZJnB+mH9NxxuesMCit5Mu4XHq8ca0q9Gnbybh/31+xoqz9yPn
OYpvwIetI1zEBcK42XaGrR3JHTZNFlCg3EDBr+InH45pAGkCZWT1hlSAyy1L5247
132vffRllhZ+44IWhyWF80bGJE7ybgdJP+rygY9LZ5hM+lo/FPA9mJYQswyKGIBt
2GGKdqWPshrKOQiq0u6qUIoFNNTVTuc0tGjrXy11xAk10SnYC5kjxvxSlPMUbWIS
FRgl/aJOM/6HhfCaPnVy8MwTJv5FYqtPclgU/2cBVmCL5REtuzBXQ2wIBLV4zTqr
/N7Kj7NZBx2w+kWXCTUzafKdaUdRhJtdtNNVpIMRi1ad4a0U4h2LXwMqrDXxuKh7
BIJPlZ2vJYRgLu6McOMc6GFtB633804UOmiry7+D7/pQFa7WYgxdne7aup+jlVpw
m7s8D4n3mUkkvSyYF6DsTKxycKhXXQZ9hzOjsHWbClKURrFCykTfNofoF0Ytu0Ew
8fbqnfHaHGZ9tTVsSpQxAwz6YiNB6UdbwrWixcND3PxjbmEy7vvP+XIgfaAKpwvz
zC6gn+5p/OVVw2zwUxqds6gl5ES/VTO/R87SwaQESmTUWFYv3tB/tHYit2llANsG
BZv2gcVNrS/sGRmv7dBrt1jMp5qBQ/daQIZxJGFatKviznpfg1JpwfT2Q9F/lLkg
pzKeAFfVZFeCODL3NG3nY94EE1sE4/Kd4LbYTD0dVIFtycEaaRL2kXyFQz3Ev+qf
EOLvjHDcEISw+yHX2VXKCWvSxxRajaexrTCEYxCSZiG2aK8HfFbwFsMgUiokZf/p
4tUlzml+LPDUnHgxTNQYyzYhjmDR1EyOwd1hEZRW9X5amyj3kFiZgrc4BfgHUOJS
ymYXTslfLqn9nN+FEQi6/Fk/fqlJdt+U725ZxD1myc/4yYN4aRfTOsbNZi6mK02P
ouKKjvr/LH1Z12WdIkcqjuRp7t2RhiHOzJu4Fh9/TPyRrYUY/VWSEDV5QnO7e2el
9oqZLGF2200ehZb1eLLP5WgZtyvCJhB/4kh8b3kjr6igegFOeZw+Pzf+RDdVDZl3
RFGYyLQhdzzt49Ix6eLJ92yJIKA0RkS9BAExENditonp1TjKP52mjxcvv0y2sUpB
NsvgpDN3CxYmsFZQKXeVg8cH7p4vcmesVyJEcf9XSBuGidPdlJD4ixJN7CloDCP/
81XtK+qvagc+ALwdBA1AN6ISN+19OwYpNjMQXIfZsZ7AjTWsxT/9fqCGuWbi1VOH
HQWWuQEkaKCiuLXEt4oiAXfnf5UOcg+nK+qa6aW6ieYDsYoCeJxQo7b9p8X0rV81
1W7cQYLVuC106OmkNsM7ChfCl4sBGeYdP03sEJ8Nm9oxvUxa5k3SwqAkpDnGUCXs
Rg7uoaW0IMCKlzTMe6CheFkxJeckGFkw/VC9oLDmu3QncSO8xC6zL+gfdw6Un2KM
TODmGcLgtgAtcPtWz9hBHjDR5bURhBy+aa7GtyQm5ltKFGbCg56Nt9urc8JjEKL6
9yWYCY49P1KRlJcRK95ApC1afTOhEFnAOFy+KzYC8eyADilJj1G74aYMk2J2dGek
pDGkUzCJHtH/BZFp3kd+Knt3TOVIOJ4YB9+yC62XqGY09TMHOOu2TIpYb2WXcYeA
X8afJeJMoTn7VFAbr2Spq22lEmn25s0DK+8NtQq14UhihWVin/F/NhtfV5hd+0lA
jpYd27VzvvHnP+iDZx9ZDZjc0upKwZKqIPMWCQkmwMR/I7FMoYK71Yu8ME0JGxkQ
e372UqXCFhVLGt80TRdDd7Y3fqYp/Uq4KrnbS99bP9BemmoUlWzUFRQJzr+XZeYJ
pNN9xWGFqpS57zDjlkOHP0wQvngwQouEgTvTtpi0Agc1JpCeswbURikn06uHoyP0
BsC3NctJUxOOTf9raDSVCFmyTL5ERA45KRmd/ziQ0DB3se4hQPeRG2drXCwNc8pJ
7IuuKR5ekjrxKJaKH10hivIEksTOp/A3f1ijjfrQdcsLGIipOZS+/qF4GEHZOmzf
DaRhHeRbXYUJZscCo/y+my2+LTubV7Tqg1myrdsO/GPpikV0xK6sXjktmljahQgx
RdTF7azgCh5NyOZlJajcDt5Tfo9HLSKBx7fdLSuzQi2/8Hz5gwGL1AvbbmdlPWIz
8Pdwx9NQSy4XbrErkAxhcD1wJnK0p6fxvNuX+c6VpIAvu6Y2ofbkS/DwN8NiJWet
uG9XHThr7pw9PvT9o+sX+Zd6FFCz5Hl+0y6d57SNTfPeLjIbZ4iuvrmAQp0odIC+
OP7s80zE7bUELOcxYxUwbfavdIhZZ4EsKJdP/dzNGB8lrfYF9fIS39LQ1Sgnfus0
lxHNMSgg066AAd5qn+fsSoA94k8UlU2Ru9TFnJA7C/jRpTjDDCApT934b2NztNd3
nDCV7wW16T+PL6HxPd1SokhYwQdXsuUD1CBwu6Peh55Knj66w8WPRi1G2uoApQgs
HgiamIrt6Q1LcchDCLHPOJIbVAi/Cw3+dflj9jLE/Sgg1/FCDmPoY+6ZuNkkteUn
EXY6aHqcKsYm8hwqo65nMUSNYssBOIxS7nTniL+G0VXJW6u8/lSKtseR6O55cynK
UU4ffv75IfuFUN3W0dAvCwcjoshTjPZ9bFueqYO20vdaTpkYtxcOjDJWyG84Nkfj
nkhbZdWcrqbw1a29XhQ7BwfO8/Ky+kPaV+hFXX6jzQFVo+GB9B8dhZQ8LmM2gTIk
+iG0riJavpzdVuQyIFSABjnLXTDo8evyk5gt6LP/ChdJJRWuyJ5E0Wi37lnWJOAj
rW2zHElJdL1qb5f4650qizzRtL7wZK+cnk0rspizIR1Lci+ew0B62+7Dk9n+BwMH
8hKUTl5wpuVQEYPMEP82dwPjdujePj4l3A8QcoFZVOPkpG/iJVS+fejsI/snyLAd
5HhWHlttSXCX9MV/WYIHp/lmx3CdYb87AFVvedqgRRMXKwAzKnggFIUbMbi0/IlU
7jhVANJAUuBNzuvvyf9VXtz53CQ+AdLxsChVsF8BpO2j7XLaKNpJPpL84GIjy1NQ
wMD4BATXFithMpH7sZd5VFoMNBEfTRzZqfYYy5ShvMzg5tzofqN0R4XNwJ7rysEJ
b8kI6W3nqSVyyIgVyCWojRUZFRI52/lfxf7yjQLaMcVLZadTFWbSqOac5e+iXq6S
A/C+WHPCasdD34KsPb1JzqXOrS4Ck5dxEzBhMPxkaG+MVTyM7hWgEQ7KTp2CnneW
Ikc1TZQ9vIrSHHVenPycIjQVYoHIZQYRx/TfazMCL+nsxYV87sNWS1Gp3nL9caiR
tjRXqrO9+Q5mSGRo2HFsLivKUAwqAyW/wIJ8baQY9jMjfqflGDTllhVzH1yLeX7I
mHVzMJRh8ZJEy7KWUFYZOxris2GtaWecO9SSmbS4IkDVDhENk9sovWwbJQftt/Fa
eMHr/U3MUw3ZoiQQr+80e5ITPy2E5sXxi8ijQ/rVIxnpvr+HKbW/wAO7sJlOtkRI
yESncJB4n2fHHDlzgOM8NgyDBJWjsIJpqzSK8cg7j6j6JHQDnTk/olJ9l7TbK/jN
l85QJ2sJxZjVP5OaE4Wo9bHE5900nQ4K3c41OtKJQ5yyJUq/I7K33gmAFu3gbJRa
MsH+JOYMjx1nv3wPL9rbBHOEoPQrjNw+zpZFLICpYE5qNos4xtvMqpNzqZUCDtCg
5WwN8R4xN09DSOOJN8/XLM7G+SrE9v3xhVF01hDYnHl/1ZtPtcCBsugFGC11Yfcr
u2P2q2Naqpjy1AG8JSCcM/dkqEMUe+pEA0bCk6gbAi9oOk3HVmQeBij0d8o9i/Bx
oe+vDxAZ4t15AMphS8rjZJaIxYxijk3lxbKr32Wuv5Au6q71VSXJok3wxJZ+ZPgp
NHal2jSSD2I/RnS0Og3ZihHwH04YwKzFDm4Yas33eJxrafQt0HiiZ4UT+iFvtqPu
ftv3euNPh0wD3zqGvKVWcCTFn8QbQ5CYHchSc92+kLqmBlS/eCeq3FGuVkDKrDFu
EX+wMbcMPIPqEhf9jn7kZEeK1jo+qos+V/1J7tG4NbXVwVYwh28QGCgvneTqrS0E
M6SczkLluvO0XOTfvnXkFEqsLv5yQpTftcIdSgm4/g+YTajZUrgXTsoLw2nVW6lg
8YBHOYmS9AkSfPX8s980hca+nz1obxz5up822u5MMhLOo94srYhz5ZwK4EjgYI9V
tdR7nQMXIzC6jPIKDXVMi+2OcG61mXp5MHj3DSawPYv0QN2EJw5U7sn1ubizEQYP
9EBN7ilwGCGVpwJ8EVecysLftN2ZRVnoSR8qNMG7oCNvxDkZIl568kwqQoBuz62r
BodLK+Eu4tpRIUCQRwr/0N5IPU8S0G6MOBKQbuQiIseEshCe+JAw3gLIDDZAMUos
LEItBrl7UzecskxGdiaaleiABrXNLwOy5UU4xTe/+Qq7pMGTkhWA9cqZNCiwgPDe
t0JenbCRJyxrfF2UZdCdmIeBSiey8rhqdVonzbAyEx2dq1FlyRO4Hgg3EYkcoh9o
nw5/fcfjob7OKBUNuGFmglBZpEhCwlwAaq1NOMmB6n70J+IZtHtV9qadFnYn6v0t
PcykUy319GYgQzx9OlSz7FENMxcUx8pWiRbsA4F4YDDzu+vqjny/uqxjo8taHHre
2+neAxVE2V3mtkgs1qfhwaKVvMoSMN0/Wp43C11AjBBHx+3jsgeP+yzKzrJT5U39
hsehVBz9HFjiDjfAKr9FBqJfdRtcJXUJuhg1s8f9y0F0epYfy5lKl+Wsc/ispgxh
noQadADUMn9e8nm4kzFUJCuqnTAjBgGE+ax4Z3L6yaHW10at9I0fM02K5lsEGdbI
pLrVe75hY96at1cO23YIFwbryAOrNjPe6k0bOtQLXVJfWbd17ghUB7cs5VaBwtPy
pShWMCY+k40cjkKQgCMZEcnlRihbbvfunbaPEEP4xpFfPuWt4mHwH3WMvs+MA2f3
vRUWmjBqbXFN3OVNvLVc7KkNlkC24+4axQt74n9Cp/ZSW6/GepoX8XhMaz5BXCm7
I1SSnaol1+qnMiUvjXWuJHtPsVoc5pneO9m9bspODvucMbYQJCvNfoeWB7/VI/98
NXARGur3UmH0m1SHdBDiXN5485+Cw67bUov45gv24O7VaYrrzx/Quswpz00pmnAa
rJMk7g2/j1ZMN2ILcb0QKqAb5KGcAhmSYS1jZRtiYdIlyVxfCy7z4PnWTFkuUCIU
3owS1jaPCGeQOPk53L2H5wQwEGJlXCjVSXfB+TekWKKueqYCOL7FJSELyVkbBCKz
C8DkTUdNuP7yryB6ifeIs4vVHAX7KeGmZhFduuajiXSODdaRvXcmpInKHXsiegw3
sW0bINQ+4RIqL08f2h1XqXNGr8dm2i9M1o0+YQ9jH6pKdZft4328X6KkXwXSdxW4
s7zMIVkAwhFs4eiF6JxGfChC1lBwmpxrh7QlRiyI75CuL9LiWZJEzEtP+1rK05Nk
0fVbqIQj0PuoWDHhfmf/DI7ELHG3dxwxFJieyyss9WjUbUzI7KksWN1h153DVnZ8
3yQR3H7rc8A+K6BS+qGbuQL9ygQ6LCW6N8o911Tky7PchLaxWuaaZuSpqINYSBqB
i6V7flW+iRbnBG8lqD2F5ErN4azz9gAO9xOHxybDLDTxh7PFiOurNhfmwr+but8r
LkmZsztjJBQ1vbwiTMP8bqTmRiDPfEbpExepTbhVxvMnbfZ8D5660A8EwYEUWAp0
DdKjgpAYCqFwom3YWKQ+8ZjdSijqcdfB61sES9XwjPO0bUfPhdywQDQTjlDqXR3Y
4WSdNaiVm+lOHjj7YbCotBcv9QY+T/DsXZ3wLqTqoYtNX7EcZ9cJtYtyD5C+vwBF
OR/alTTsA5GzHV38RrRmguE4GQnLkUcqQz6w2Oib3yCsivu57nSoYezYtLzXAB5R
//roQu2waOE0qdIgcuKhCe9alIjjmxRNs6HCmzt8Q1JhaYXKOi/OrvofYRinSD/z
eafGwyyMl4lxPwzXghRdXTSBfZz9U87KmEpKzhAAQiPpJOoNQb7DyAt6pkXON9cu
DMdJ4C8ZJLTQ2zN7DNO75fDmLZJiOtzDbFjAiDdRKdZocR47JnP2FHyulCwIqk/L
tPL0u9TSR5o140ABcpjpMlTFgch9pUBSjWXtKCJtFGd8rF/A0lMQXIzX5zzWMRKA
aCt3q083hhfLus5kpw5DxtpleUS+eBeDihKhB/i224WnWjele8STtNzRz6/vdUMF
glmr35RaMG+ZQejeLjhKmGd95XaqpNwMScN6TPvIA9JiKlGdZGh/I8XAi6Wr3Hk6
YdoQedRGqXVj8QeOdpbpJ1KrRF7gz7lnXdQrZBtXwUbLuoTo+VxSEo4JeGnSkwzs
ynPNE610jI/SDDDuR8r+uarqo+cyQp4CkQoR+yASu2AYQyh3REU3ZyLyHBl7TbY0
TfsQYwY245702UUiSGDrBUgVsTkypmnIQDYioW1a6aMso+WLnqQC2OWmm8b5ooqu
bwvAoS4ksJsVTaViYZXE9O3NR8ORNN8AAr4R39RcDnveAsiLY1pj4xokCkmcqoqa
ZLmZWttb62JIxLngNSAiV5vW1ln0Vk+S6JiOpGjzIbfDo2sYV0KNMKWiA9lf2X+O
bCkrEXBhnRhaBYfJfo4HvDcrbf5PqJp74FVahgXfVK9+RxpI01DxTRuXgynMqEd7
10Lk9ebeFDSbPcr1OCUXIg689Alq0B9wXyF4PWI3AoONYB5ZSenKCQpAD+QRzkkS
PJIK49oJrdh/KfWfT5NX3kbhbpnE9mS2c12ZGtMLfdI/C+XtreXDIL3wOce0xK4k
zkgWm/NB17c0ZonLWx3jnTgWoKAZGMsV4/DQmhlkgz09etkTY3HZGmUdgtWge8Hp
AMH7lXdLsKk9RFmNG44mtO0rw5iJDETlRuCmmDsJ0r51I/0Z8ASwesQmp5Q4BFFX
RbmCByqg1oUMKSrIKlATScKd6FkFmZAxdJ7BGRnlxNsXv20IgX58gkvCs1Vl5YTX
UKGLjUUc5uklXFua/8YxeCjZvJGpjx/l69+voLQ2tV+XUxhWbv1bnOoOoMcbKpjY
Y0E/Wuf+XwxkDzZbf6DYXHozvs5F+OTQwa+NXIJ06i2Znr0+KFRD68r6yaJruxJH
qDqLr8bREKfHtnOWcgU++mOmPnIxlaqo0BmuoWNgSU7xj10XFCGT6Nsog8Z+x/VN
p0WKDH6ur+I+JmkQvLhzrzD2ytghmaSlyDZPXtcz3JjXJ9BOxpPiQAkYHkCsCjTL
UqMA1Mr8uPisqJWlNcgM0RKW7u7IOF3Ibha9+Zbp4i3MIczpfDWYoE5GknbS1wIH
LZAiHkUHurMuOJ5H6qMrou9LmlXhiGZvHtddR5SrX+hXUBrx9iqe387eAynSk5g8
4vwFBzYjrUluO8KqdiCm/3GNHgUrcPq/JfuVR2kcNMX7S82icgE9tuIV81pqoYKc
XfVQu1T9EK0pzs+wl8f82fnyXgYAx0rFgxRsUA0Roa6q4070zpzWeuXb2b1UpI21
COAOHkB0xPr3TnbS+FcS0mydUwqmzRqRYy6HFEr8nJuVK4gcE6cLAO8394K3ebQ+
c3YgiHM0FqIzLbQKDIuXRGZVBJ9hpkbbBqC2nsn7VURXbEKKJ1ysk3QVXFoUcb33
2bgGAVOQ8XNavcFPFAhnz1IgnGzu6/afFqT/QdOkNeerTg3G9dAc4vg5G2KaU9/l
KavZ9j24Tyjr2FgoqbwNHB/tShe3f6n4ajbmEj7Z7UKrhAandcmK/MRH+3rNRDEV
WKKohjzz3vXCZRamvaMqcp66/+HwSW1hbeB3OBDSgZArk8qtUQQjt8RD34x1YX//
/xpGp8pirdyneoh24StG6GrPJ8KnHt3oQNxOgahunSq2i1rfavTJ7yy5+MtMVbrZ
wGwcXKxTVOOFKvzw6+Z9GrzD5/8kratFSlO+/ZQcXHZE9DN2qYWDTdQOAkgkPqjc
O0JJemkDYvL6rBS54o8FnkX3LAJkPlBlMhZ1VWRXA7PquvxxLpVccYzvQaRRdhy7
t1214gpP5p6niLJFz7kflZqmHSnPLo57u3dgff+cX3TPoRIle/C1maiioE+3MnKE
9v+yb4wHN4vTVjo5UI+MNw7w9mOJNhG3PLcf04DvYz7oUThUq6qNMajZuQnWyDKI
dJbj4J40yteKtf1vNFkTw7XZh2bpxyBTc2hNbbuzPgMvJAXYk0Pg2tUBPBr96hOC
XF1y0nuPJUFOlXKCtZxj224tRMOh5hkFT6vPw7baEgwqddhNEbq/YChbR4ykMrb9
k07lU8atiu8LAswakDB/jLuEBSsrzoRQVRoWP0wiYHoBnpXJWXhrk1xT4zCLJ+bp
WPYfeUXN0vuuYaaifZpbkEKhuYimQroTKccS5D2PW8eZNnsqqvv1avxOGF0LLIrz
8KjBwPBVsj5RMa1QaR5Yp4rbu+2GXs+ZO7NxDR2FdIt5Z8QxwALxv99V1uSy/zrn
BAocqr5HbKhqfHO57HCeUDvuM9OdJ95zzzoddEsA/FUXJVoR5cOV0m5NzTdiy2pa
AsW782k9tphy9PA0Uwso+AiQTLfPVfvyycwQzt4EP/QLepxHRzidLHLmCy4dPM9z
L20nCUccp5C2Pqx1LQ45HIzlyZjS2j6t58QFjr2eM2G4IMFhMbAwqgF/eaLyMz89
HKqLVKOc8pVTNPHsbwiTaRHV7tExVaaTNExfjBUwd4QtaXrHXKF85bTFbU5Ukpf7
J2B6hll2iOvWLImQH7aMNIclwDo9AkU405rnVQCfv+N40Xnr4T+cKPonX/y43yAJ
A5bQjWMaPsQRfOwekWnGxR1cCQEs1UqALvcBF8xM0U/Uwu44S/98SD2uO2nFGpwM
0y7y54xb/Y2IB3atfyyLUpwvTgZQCIYWmWEzXQYruG6v2IOW1Qygsc9S296DSrae
jIsCskh8fzKBGx7DQ0zA+CG7sY+Hd9Pv8oo8Q6/7faL3r7qQTSwlyYbFL0qiyACI
QU3G5cJ8PGjjF3UBIB+6fnNDIL9Pjt/VD1ny1P8uQE3i0rAYi6dblMDLF2QLNgQW
WWy1GP58I2mrzTNI5ouTk/4i3lP89nL6ppsP4ymIwiom+B16Hy9P+LWyk5b7P/vn
6jAxKJxWVjreMpPw97xc27zv58QMgYqALdf+DSKWTniJOofUx3XOcNcI6ChMU8xs
B6wEt7vwvhcsvIOVkMKfD+qlHH/IVMqwdNSwBN2Ysbw/Op/eZqG98nMtaI+Ez3mf
/I0JHwTb/po7+XMW+sGPILZTyhvZahGD7uuZnqWKPQtKWsomymRW00JMQSKpkwdG
z+5kOQp9iljUa3Bz2trSSUjj9DB9RklHYPJfqR6QBp6M+Haxp7I5N1V13AUlNX32
xx1I1B3XGbM/uP23SaQb4nh1eR2/no0bKyrU6lw4KDZhVIkHuE5FYolxboEWzmyI
TWrXhCLNl2hSBA9H2mwMrFmyGZRvz3d8CS/nVW48LhlPhGIRmfhNDxn/o/6GUDHp
MfrfDfloiwxHhSo6eipjL9ntTIsp0kxzR8iW+SfyrzN4HIxornWtRd9wrPgCPrjX
YFjwifYnP5vOBfD8E131XvYTkcwJxnMZ5eebHlLqHXa4qKHjdLihjO8mhvOyiHpb
oU9K2A90gJF19KoDrlQCesf4Kb0Gv90gNkSduGYPLxGSOpex7svYuPdoAgdHJ/K1
JQnDG3ndFOO2/LqKwMCOfd6mVP8wt88wnvTLRQPIgNnm+fG2Fmoiqny4/BlTqlQ6
iW+xfxvkg9/4qMBvKADYfAAYlbSu1SRgXRI3gWWxenqoafYvRXhLUF3FUxob7TFG
H+Uc/R38/HjIJJjo/mAD3CFa1FTV41kIPlSHgd8zrKiYbqCNmHuOzwbkr7L1SGpg
e01YE8WtvJdZ5bj+w1s2p+z6x9cDupc3AC9uBG41VzugwyM8S8j41en/vIL+wV70
sy5HKDYCKLEqGUOhNRKBDTOemhvBkcG3y8Wiaf9VVOaGqegLB9uW4zGTS/rJ16YP
13f9vXxKiOunG1KLfWnVRdgdr4gOpcNbPyb5ZDaDtaUpbb0vafE5wacgRDXgvGvz
/5iV2/S+GgXo/g2njfwqmUX0JlN0pr6JqfbJS+13IdvRGmUvuNTOLGzPsuCR5y1D
lW4NLvm6yNM0CTSfi5YDboT+ZXX7aZarFgEcsxs2ZspX7zzTlCiDhEAcXm4iKD9Q
WMF/f1wxyHyr7VKKI3U4Pl3G/k8VrGI4xZ1xd0Boq0wRnyADFa8tSL5mCbp7Qvs1
WPbbwN42zQ3GfC5uTPFNOPpEEfGZ7iuF8W99ZgxwKhPZXEjUMBaqt73F0+xmsuIk
dDplR3PqHM9Mwvy0OY4+/fWYCJbjhwO3Q+L7aD1r2LYpu+IgIAsCvH5EvvvrSqmU
`protect END_PROTECTED
