`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MC9ukahTTNO7sngqdJt9KNj4ZZ0aWDezzE8wHaezEUS9MUtJ1LPrmnTu9Kcjr4dz
CNNX08Y5xJyLkFpFOOfAa0GlDKoe6NMOvVSKIEX8WfOYayBWXkOb5S9kOPJ/RRdC
ueJKaNJ1SHW/YebfvRO5VcynWO9tW3tJcmWRDKQo3UOKQuOHHC3vfQdPW2Sjvn12
LPUt2H0b524786DbmtDiD9A2/vs8LVO/ksjJhmibyhukWrKRr+knxJMqXzDxt+mm
P5d+xN3LjePKG04RLuJbSHATKheHZNyyytSdRz76HQpjUKzkR+LAQ7cnP7mZi6zY
KFN7Pesatzjdu+3gpcs0x+4Zf3RfodQdcWBYfHGAoS04AI3RCISnlGPsJbNrgMP4
NHPR3/NNW10roOvCaGBInMUMyb4dc6+ccGGA+ycqi83UgFTY+Z5hLuQA4xXkPMg/
ISRKVfTz07bbA7ZCV6/biy1ANOacGji34Lr5a2wl09JUi/L6adqFEFdQW0PPHoNX
F+O7SUeQfFg0wT3O1iiUyLmtjn2AnV+o70oO56TzqTg=
`protect END_PROTECTED
