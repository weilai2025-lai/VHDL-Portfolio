`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojRfEoD8tHqscwrEG5CqAmq6qY805uknV3K10GLJNeDK00hcWWwUwcKG4NJdGIcr
7wj+UmGFMS9htjlTvgVk/9hLqPP4qHFlTwiYAw95Gf9DYMQDTX1X9CwZIeL9J55d
WcG5JTBLBF45r+GnMo937OIv0gGq6PpU9xxFqwnvIZhgmlILClgARxZ4S9doVLL7
XX9hanWCXuHH++7H4oO8Zfqfskmsmd3/G+C+OOKUcwuxiW7SfXpSQMCB1wqqCvpq
Y34EWVSZqzGpSQEIDszaMVy71d6QjuIwXtxwFYGQ0ZogpTRP/xtx8+dGCqesaydK
V2oVgyVDyarQ0qjXyLWXn9+OlnzpAW7bkTyUZv5/WevVKMkaSvyDGS4dEA1mZ773
CiqzEI00lrNubehSUU6bhQ9T+79CVA6Lmmq2do1hlpyntOhofjbnHONPmmYJIy8l
i7qR+nJjs16UbGYLesLUtSDtZ+NvA4FwRtPEv6K9ng2uOrIwfzmXjywNq3sB0iKj
V3SgDg4UabJHwMVBa8WRAQ==
`protect END_PROTECTED
