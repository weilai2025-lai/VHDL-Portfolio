`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dM84rh70D5/u5Q+BX6+uk3hIMHT69Go11tLvPK1WFlB9pBbNpwAFzHS8JT5bo5j0
KY2TKzd+QifLkprL0lfpsjRWhuLomOe6jdjeG5oNMlAWNhfqyudaBbDqU0a6cVdw
CtrIcoFa23a5La9gFCFFWFdaoyPAq+4iCugH/HI0lxsQbGuSLl8yjet2mJTZrmXz
Z1uuZcr/RCdv1ZZX+ZqZ+uBjH62FQ4jNwpPkU0VsGZc2Nqs3JapYGHxZemDJPPWn
6LMMsZwttEOJ29e1mwOyPNKYmpN1peTRA3PtO90+AnfWkFNA/INBbu6808aHRQs6
3Ei7o2pbnzjTFOfn1OdWamzto3Qk4GDq+FZQMI2atppK3tueIF1mxPtI+pGOti6w
RmcWZs4+csf7jQL1mNfEUuKfllP4WqRwVuiWYYQAV+XE01s28R7ZsMK72PQ/JHbf
lhCdpAUnrShSyQNTPx4Wk7CNybD58yyklkoT6XAAAdeW6bwPfcqinSLU6DV2wU8+
A1kI11JL4z+g43sI+tAMqu9X8k8sVXbr1Pqzkx9ef/yNfjbrr5HJIt1a0iZtE9Rk
HT/SNH75ULcKYVTXyfoJB7go119IFm2aPPnPVdqsNl8MG2CWEiDkC8xW2wm2UafE
MYX/TuFMMwMLcQ5fezstl8KYgeW6X7ntDN6AfT03XoHW47XVJMOZcjZAa/e2/Ip4
F05/lEnKHVNTY8xpEYLTmIXpRjG+VFYf5K7Ur/a6lMxGDyqX2nTxcxyaAyuN9/79
PopNFsPtJdhb/xS/eUKh20kQ5gQMFiq0R2jMEbzVRljqiQvzfVP6NRDTCmFSLo59
tuR6JCCZKG4sEIk3s41luNthj4C4i/mC8miPE4QNCnhA0PztKd/8FNhWBtU8ifig
hTqOu+eX+T1qXuQA3mBSPIRyPA2C6KPcnq/AT2/viv31+5bU7OXFgbSM0ldU0E5l
F/oFG/JZizcj2WMHyf+iqxD8VlrQi83Q5a6lofc8gJb/ZuVxa+Wo9CkPw7e2as4m
z0MlxTDyLWTEqpVzyqgp7KiR6jY/NZcZI4E4cUithVfZRderOaczBFZA/t/OHTyT
aidZutUqnqECDwOUGKpn84MIndg7JA8Q4kzhVnZfRAt/oQk6agS0sXsyeGc/Hcs1
zN7oiRreG3LR2fB6O1z9am7MCNzjPt6FCeSn7nKPNi7hs5sfPNCoRIMwuR+op9u9
Kx3ctfteyZXHSGM4WNv1Vh6WevKB1LCOUQrS4a0srak13atmo6+54Y97Oa4p5RYs
NbiQurHT99szd0GSQMeBe5e0gfR+IjPkSL2mEpmlZiiRojVmMmwSfZgP2mjmWHFY
747BigCH1FrI/ULDysHIZFhewEy4ZFsYtPqTJLJ4hHFBvy256tYxcnb/YUPWIUq7
9kSgWw/vHtq0R+U741xlxWuWiaocE82EsIqyTcnkH7Jxpgs7YtZtrB5wj/LRYX+l
4A+22mENFEZ5g5CWN9d6a30hsEuwUsKiWeKbh6ELXmlhogu+3THxbvYO+Bco+zsP
YdsvPGPT0/6gRI5OYljH5JTjz47nwH6db4gcy3HW/p/oambF2NOZrnKSCkfdVukH
9MeYLlzM+p3FcFG8G5peill9hNqETtpbnmatiAkvSmqmkqliqFMwyEBjt41oux7+
1aT16kd83fLQtivYe6wVGR0BPQSOKtgM5fdig1cmZB1am5PsKMQcfp+igMI0T6zr
bebsWAUMA/WKuZskNthDtb9BOkB+512Pkv+K8k8XVSbTr7zUjYj9qhLw2Vuq1LN5
v8qxiWWrEtHE/Ktchh64dQEgWJIskEQF7xusoPfJeCCfzg3nT8Tm9ugAN56Rb3rA
OIzBc7RQy3Bw1wy1q67RvbF8TeEudc7TeGL++wx97OZm4nDz0SPLJXudHSXMlLEn
HVhpJ4vFpFG4xq65IwVXdJtPNCajcLGSNgF8awz741ddmXUYRbTwDNRFhMakeR7U
pnqZgNXqx8Map3qhqX9M3MdlC9v2FMIld7PC2Ecc4lGwLtWfke4hi/JG8eAhF5P1
M07b0w0PQVq39zxjYcviCrgJaaNHpUQK18rn+VHpIlH39EVxqVgXiIDq3L7qRmaw
fmNC7bLMF1w5WKgMKfdL9+118qeyHT2FcxIjVgrQGTlSYc0lV1uXpbd5JpehYP/n
hIGhVKHDQtPu5WEgTB/8wEhgqJP07mUI8/66Pc384Ia5Irum6cj4TR8PVtO9SdT9
SeI7Qx6CFNr6VEcS9RxJM6sc5V25hpIYm0+PTgzFkFJwPq9XjjgYPbS57Tq4myVN
cAwerPU+sSgHoP0QUoou/A065+MLxJHykFyDeczK1ZhyLrxEgW6F6/TPBht3Pvnu
sW4jHR5MKQPEsL2LyJqdqRze0vjT5Wj28DxIySuSgE2NBiO1u3iVNH166kNIWsVf
qbaYg2oP1XeoO3B95qzejP2NTi3/9hYGvH1I2QztQ/+ZGKi+oM5R06Sc3sJIazCE
YwNL7Z9Cpaf+EwyGJfxhhyMWKg+MF4jVvCantfS+Uzo=
`protect END_PROTECTED
