`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xcvlls6caYzE94YFYj1pb2RRCLswZboMenfezqnOZIIOx4crsDU9l3h0xzmXE6O
konGcbGPjp3lewf5/48KFmNrQFFtOFx835deJmAt+hE4EwtG9ouUW5SrMlA6bMWL
MuuHgyxt6BKb9F+8OcXuVpsGCA5fkHwYrTVQrvaFZQHvR0rM5pfry6TiFVdUH+J0
oQQ73brHs4RqoMx6EWGSRFdpZytwQKClzEFnsSSc7Gw3DBw1vphLUTd0II+PsONs
IDUlaGv6A+ecx/g1OkZuC5rZzn5UedFYcspat6LRvSTWhXyHcaxDVnpS7Mh/WWnK
7vCma8ih1Cwhp30Dk0jYOnAT4PXvGuFMEJku79mQg9EzNc2/5A/BRJ4HXb3HiVe7
OZBpGrlKvwCr1IAV84Hoyy7BPGCPqJ7N//6Pay1ye5NcFCfbByAmDt+Ccs6huCEJ
yikFMJ9n8H7ijzslr1Z+5kXI/7EiQn5HWrRjEp9rwiFO82ORi6Lad1uePfRjAmzs
8Lc6ZSiSFm71QDz8mWLedY6z3AQKO4aYBpTJnfP2f1CnBeFgGz6gkS8hJqm5gjEn
qXT2LXjyEv3ihX0E9NaZ4H7oFi0jnTRgFec6CLQvc7H2QmDaQLkGKmycbG/KC6Zk
08W9omzTO102pfRnc9b+3tA7twDtZ3yvLcB6UlDsbE2dquYgWrg2gb9TqGz1c3+M
5DZkP1IDmfsgnFKterC5D6Ra8QpEumtgcxrWIxF8QCQVz+8wv6bYy5sbUA5x5fWA
kCTfZ1g+3PSol2r4Ss5EhZlxrBVK1wQIwwk5M3JQTh+9a22dODKC2VxD10zFYbJp
`protect END_PROTECTED
