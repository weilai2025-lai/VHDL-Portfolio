`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0H+BrzxWJeYoBKob+3YhVrLFi1ZiLO2xMlT1L5Hkj41vstlcNZ6JjhTRZ6VOIY1f
fYX1RAyi75tO533zo3D7oGuZkccx7lYZdlcKBi/uk3Bk4tnDem/64/GQoGTAnhiE
d5kQL1NfOaNn85q//u2jXJVSDQgr5mIAmiLLlHfCqwYB64qARstVTKXhGlRF5/6N
eeEndhFCgKqvc4P+q2C+vtklImLXod/3q8pdWhBASbVuaQZc/R/UfCoH0v5X/qLN
yP0d+c9FsgU88kYL5iHVgSIMiD9qKMP+/DliDPvvb9JQpii072wWoJQDNK2O4vsL
2eM24im6Hw5gg8L7q25dYMYOZsIIQihsz9Ee08aYfnyxBYy4aAer2dNOJfhxiCxG
xQ20lNJ+rwSeKXiOJ09YsiESBENsI0CGdVAD8/DkNZ0Ru2QD4sNKayJrpuTy4Vk1
Di6uhrdoCvDR4InT7U2LLqW/oKiLTH9cpL83Wmn/1nZlvSNJ4bCjuJWrEe6FF0Kx
/oU7OjJPmF0SEcVnu886bUhmZ+xOVDy0xT2JW9TXLHnd9fvw+E5Lk3DgDyPGFM29
002HILs7KaYGFh6huneCRXh913U1Z3KA+Hcxk8KbXBxVjVpg891r7OH0MyPpjrHZ
rEW/iiGVG2VVP7ooWiDOfwmCUP3oDhCyPh1muGbxxR/7tpsKsHelP7wdNgW2jG3v
D7Mc/sAIS1WTqiErFsB6PABqunSx7XRxWu4HSEUg1IHJ/bhTcZwuHJrY5BqFyUhD
HA/gShsVdF9cuowqVZHTrJU/ZqnYfT1PxkgvW2kIW6+DZwIsZzRN1Btei744CB0Y
RrG7oSqOOntgl86lqhpDo7dGjh3YzWtiM3TY/p8M3kXVoC6RS/hhb1gofbbNoO6N
Gy/aamBbJ9iD/RCjqd4IhZCJ+eHaHw6e7aBMftcO3ny1SwR9s6GgSMaJQt+JNyqz
gdlot28w4BcaJafPYk4+vLq3S/JxQmvypjzEzvq7wgYtG1n3BDTsA0d1/BeLUR3j
BBPK/9YWzDeOek1iNLa9tE4GjrRlF39KDZX+wA9LKPsb9h6lrza2emMQ7NPipt0V
whg53xkHwAOE0IGRqsgmNwK/SC1RVADH0S/Vr5hBqCDFp9w9/7uknZtPocYNCx/v
lUyVnL5QGJqXl8bE+gGpC3VD+mxQ00+dE0ND4QwBwKVx/RJf80mWe6yaKgAhi/9e
xTlDkKJdQIQHr/4qqov7KZAHAKXYFIRET22f8gPVQS3ap9tQZMet6N1y82M15aUQ
8nmPsef7gQF0G6EGs9MyD33HgxNBTVXhd1ZsNmXIm4fwkvKH5ja7YySm0tXO0Nzm
hfAvm6+gxuhH0v1ngW8SKLGGyc+e2Isy0i2aSDP6sRL8zOarMHYw43jxKClK/2ng
nf2tLjCGLZzp0g2BCFo5ZGFhdaLcW51TzvOlR3NL4Ib8jce2y9ZNzjW3JNrazIWf
WoW2TLaQdpWM2uTUsJ1INxFBg+XZ+wJvsLOYg3RsF+KPO/UPESpkM8rn700ytUsv
M96JxjPwVj45wzPxSR78vBT6ORqwroDmxB2I/BXaPw0j8jXi+9JEIT/eK1FAD5PW
28RZ51kxDg2rZEoWhktXDA==
`protect END_PROTECTED
