`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0LoX6FMux6+NqGQZOB8o7hRGlSz0TP/op82nySYIJJRGx8lf0Pp5iaezxBADURP
+0+rv2+AflVe5jaRbvdrWEJHfNNHf16xakKX9Yl+V8Bq4z7VR+BD2/BcQk16aMkU
Kjg3qg9J9PGIddN34QNMu5TzRCyve5rOOtyqrIkJ8Dthy9HmQUfV09eCvhGvqYEr
OBeBGH9U3Qex2iGYtUnCAH6XR59NH69kwpDL6FI3JVGussMpSdBdi7+UY8YJvnnh
rzgO1E1XnjyqvhX/mTGLhA+bRVabHXNqdpMNf+U+8ioqYlDQaPMLTTK4dyt7ktuv
mNv1qCt/1gGSzXwWdSYY+KA+sMnrDYXBzkfkI5W5qe4qXW0CUO17IQ+7ATjA9KuE
T/KfYXjKYhRx5Sqbn60E9lMdv5KrEEaBaUvBunpfjyETRVHN/DtgmvUYVHkZNXDy
OC1I7R4gBh/YPOJq+9UB+ZiT38MNCMREi4aaJOSupfnUauLuxTs2PBD5ZEOvEU2y
h6xqofWDPX4eNYBst1kna3Pofr+sce4KvsKzJoaa/7krC/Op1TBdEvZ/p5qPQ4rj
NMV++5rtZdsuBNJOqwPs0OKarWGScq9CkanmgxU0rt0VnnVrXA8KcNT5CJfB5G1N
CuIxVyINe4tM35XC6pgpj3VXRZNMx+dIZ2eTriQF6XrVRFWCjCvveHMNtW1jfD3I
cY+iKjFMm3aQkK/EmehSbjfe8j442R/OMKWve/Y215LstbVrbTMdgq8PNLn7xLar
IKdXJQ3skHRaVYbi3aEjP12t1yWPhDJ8zdRtj7xSo/mphoFB2jPsHnk1Kb6ymDRQ
Oiov/7+2fjPF/Z8UhKvAlS8jXaHBtWAoGeL7Ih4AkjxiI47RrAo7+q4+8NFxyNSm
0FHxTqMsXItLkvN+El6Ux65QjtuKa26cwUDORLdE0HCgBRNpN2IlhIYr3uzG3Nmh
HCTX3OuW2X/HYbhcupkj32+zUhycG8xlvkyImRWBrF61x+J/jIZIMJcKpj2n79UA
4DWuDbBHuwp0CAc2elsDHbrFp4epNIOIpxnTyEq4Gh4eaABSN7UsmjePBIL93950
jdItyGWvglROD3raIvOWOerUZjP4NhX1s+KzeszNSx5VoNBQt7j2Za5fBPTz88kr
29aijNxgOCiQkZJ4JcicRPqXuIh2vdy9A3WTLnty0pyzUQ0QosqXF0Mrkg2Tz5LU
7Ngdbe2/mMI+gBg22+hN5FE9KeXpl55CgPK9ndAM85Uuxb1Blsj5WlfXPwOzWYO/
hES/5QYkv4w9SfmID8ldycL9NSOnNa2JTK04pby/PD3RC2DvgU7iiP2C9hi3+gAj
8kaQtXTNrqcnByGGfXjVBQdlrQw1sT+vG1xBfKbGd/AGoqJ75GX+3oBkXmXJismF
e+GQCwv88TXkJfqhyOOJIH9FpJAgbHWxYVGynXj7yM2oi0RgSOHVctBhgYLlPha5
IJjU7M1eGDAwRgS+eizo/v9u5bh+vZP1fs9n/gem+YFjriim/myVlfeUXVbrjrOM
S9icEpRfL35bhMBKZhkPAPEJMcda9IEqSeK0XFzwfK7q/mYWtjFTRCuRzYi7Wj0v
naafnNKA6te/OL6cHc1M6VzBFguyZpmbTNd4YvbF8/BpqfnpKcaitG9j69stbjzA
fFD5VnAkTT4DRYT63ImO2FipK52ehDOe6LS1ovdsbSCNGBOW4MVwTbbTYTbfH+y/
bUdDDBQsOyoJFwvyFMa61LRWCGk1U14AZujiE1G+fPjFkoSbkG/HCmo7gVIa3xtt
UyIK4iV7SGGk+tleRHbeDnwQ7gthdJLiXVWC4Zont4AwKzaKkbhBRZk31Xr2YKME
tza1TipBtp+mt1hRlv8A8bBBRIgOZ7GLA7ZXccyBJX+wxfRVpmnvkwmDZe7H/fhN
MXo182xmIaUe/+GQjLEmQMIGN5hkgtU9w+LCuxFUzkkeZy+zPKwlIJJz9fosCfUi
8j/2S/M2X1RK3QeUVEPKAr9o05XMqDEEaNuJ8pffpt3uahUHssnFQhC1r6fwYdO4
fG9bcuzyn4z4il47bXWsOa6rC3SFdjLbltZs+8bxAiZwNlnQHcaDzHxVeAogLG36
f1knNVClUWza7MY6OdFknWO2GQr0bKZYTePtVL9QHfqUtvjNNx++JLguL0GzBbX/
WzJUgSyHP6cFUBMeE2oG5wXF7m2uu4kl4jM1wwj6RPJjKaVi1dtwDJC+y1tH/1gE
Jb0eaBj7tOoHZivqf+hep3WBSwWafpYFO+28JF1io2mqZ5gw32Qx35zcfDlmB8No
XtlSmeP9PnZDXhOsMpKJVyq62NQpzJdc5FltQpete1yNR3L8aVo/NgKjEShgjm4E
WOMVRzGWG3MxST2hYZacj4q/3iFBgcQygyf5lyT7NNLmoy1+W2o7Jawyx4jIqw7b
Q5KAzOQE8+78W9vM4qHSCDMNMO29nT/FhEmLZqVaS4cs5IG/pLCbc5OZF3TjAV6K
sOqECfnyIoZGoFs+HoZcL5b57faQ3p2LAnXwkLdHyhir2HMUT53vRivxVcUExfkr
/CuQ13IIxXN7gGlapGowRc71HgbJHVmBzyHaZ5E2vAS5ulu5KQQ7KnIfn0oA/ZrS
kOK9Xdlk/2o+ZvvvcGCWieAZtY3gOTYHqe07K2Lljjv4AlBn5VX1W8NTdL0RJ7EY
YjpZ1VE+GSTW/Km0+GJxxL5h8+0Pd2qFv+2HjAcB53St1RfGhqsjGUWePvUNEJzx
i1Efrsk9CkNay3STW4+g/K5JX5r5+5f9yUteJcaXQAEAqN9jvrFfZSe+6N9EZv+k
KNlPHbj8Coo7mcsem9I19buctKY70d9qW9wTinP/CLrZiLoV27w31E1tBdF+Mnax
g0DVaaJTU0WxbUUBmtSPTX9MkSJ8fJoPEtCXAPZCqIjxeql3ItCn0tatEh1Fecwj
C452ys9JjbdMAAQNuSF+ZEiCFwX+y+AtZR5AryzLpwu7h1+I4b6HbYb/CtbIIKkm
J/nf7Paa4PES2C7n2ceBOuDyBIeZ79syuqe3dzo72YX6J1m2WkvNcPzS7s/Z9j4K
SBs9GFLjfnfjjlOeNj3CW1ybibpwqXkfloltopR6Ybxbt5t/dwhFPExZzz63Xinw
YJBOib8qmj6pXc+Jf2rhVmNTGMJ08tV4R4ptcwdy94C/5vfhZ9jJZgiqraaco8xV
pP6bD4O3gzTNhoY1y/urh2/CPAOOtHj94/30GXjFHT8STbctc/Ei8alWNlpXb6tM
QQ0Pv00S8Lst/+Xy9mWOmkHMOGAS35iPpGIYJIW8O3f/2lapcnt75ioAUQc4fL/h
SOWRn1YBR0Qy6qTaY1pl9oLogE3Pu6U7pCQdVNIKHNh4q50wddxEieBfgusw8oRL
sXfX92NuGp7Kwuc9y50x8nNt+MsaExHFfWNxOGVXzAv4kMjcebUgUNyZVpgUuq9z
htFhqX590grbZ/cY5nNxDmkr4VKO2ELnkRfUtYxO976+oM79ePUujTpwMY5vPmTF
SN4zDz3Gx753X7lCKEwXS/5pO9kuOPoY6H5DivpkfEBhEFnB7Ao/SlcX3inSk1T8
8jhEseVq6ckocAgm0cvnwG/csZ7fvPUE0Rz5I8XGAwL319dcZnkYC28MIvYQ1fNF
lvdfyssKjLyV9dU9zfIR0qHoQ1SeJPUs/EF//5BpQRf7VeUtbuftHez5H4YwrH1W
GIZU9LtqqyazBsNCGhzEac/+D5QDx97d6XZFJ8cHz5iYO4hecK8cDLgnZAVgrsCt
NnKwOFdMvbJgaes8HWG6JmMst+xIEJ0pHD20Pc5P2Wbh60lzRKISoJcGIT4gMYD7
hVGSISnJhSJNIJMljh2XA62uc4tsyKjIf4ectqJkoTXAGjBHq5HfIMSDzDm23M/5
yOHK+NkCsfhe5iLUS5vbI3q1Z2Hot/8gx1+ep+9iFdiwYtR8h5QcPeIo96iJfDCV
DmL5Bj/P1dFOQCnT5nr24DTW7PROcWm5vYrbIy+XyaX3JiByjZdKaWx6uTSDiZGZ
lHQOEGIBIFsvRW42jJRleM51+Mi8+x6IPvOFy77wYCf3+la6po4gbMBLaq+VeHjf
RmkTgpeVtdupSSibO8VunxmDEnG4Lo2W22S/bWNV2rfIrLJjJEqq3/ZEiO/leWxQ
OmQOPPHbEdIcAI3mTtOnZN56jsApi2l4fb13Lo3LqPDu27RMhgdiZr8TFXywOI1o
pbdsJbQvVyA3t/sH+jhLH+qSVQeHah3Lt2aPE2CBLVY=
`protect END_PROTECTED
