`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQ7i6xzC54eeWWztiGpw4d4zwN1qpfuQCZ51z2rjCwtmjnqU+B8qsw3+wGdzK2R6
f/sjyW4+e6UCauOgSPv8O7IbGA+zgK1Baw5ntDxeY3qFBL00fPHQ8dAEpELW6LXX
PCys7Sw+kDHndo7VRpGV0eKl7ID/dkDT7vGon2xaMImiwneY8NenWRxOs0pesxkh
Xzn6RVQNTiicGISBJHI8u+C2ZLtstnCJ1ZLi+ZO5nboi120hbB7nKtQH2VkxTaCL
lf6JzGvvTMLA8SRWRI2ZO4Mc0CGvylQa7NIw4JOMI+f9wOSQhyiglvFI0aoVqsE/
UAgU8xyyBb9pOnmJynmBqOvdWB5KhXuX2jj5TZQfSD+GEf3TQsgPe8SwXE/3zt1g
v18PZeIsfXFIvtRMvmrIZF9wlyMpyY4OnmHExZzyWMoaMcEUGMBxF0tTBjVKD3sR
wRcwSSkOM4BygSxOXXekOSRYx7ZEk8dzxFsBLGsi9TiKaDqQRkQLZ7u0RzJdeLRQ
l/zTz30Ob3DhNRXm/DHIOYRp07c3NEsmNSRXD3yVHKXyvJTBWPyHjdJBKJTyFjkx
vIeB8X9P8mt8NS9YnmoA1oXGptQLnqhcHfqNJJoGqcyqYAcPbNghWchY2EccGQXk
mA+/Sx412Q40vxWqoeWG/0s7lvsX7aby8N6L1k0iXKBAScGe0vSg+1y4Ohj4TIdd
G/PHt20N6U5gMWcRZ7bt8mPzs/lB4cbBU6TlDVXmodAGZJdI8/Z32f397MFnAoiy
wT0VrLvdiLE+CXgwjZnLQnFcjxFyw3RRHvFT+9axk4nMEX0D5BJOTp/cU95aYHTF
NJI13OTsZOCr0LepEGo7JmUgCx5/XK2vi7ungPdWm00ao005iceDLt2wwEif8MVX
IYoQJMEzRNYEGuj5F3QGgxuKFQhI8mb6ib+2Fts7ECQH0tE27O2dArXxzirg7iQy
YndIuuskb30F1uQTslICAGZaXy0KNd0ulSVXn1xwlT7oB6AkPA3Q7RZVMI5sl+hk
UXmXCuMCGtLEOQFB1DA+x8exokEJQYB0jMnDm9c/h9jA2Zbghpx7EQrjA4wW7Q9u
`protect END_PROTECTED
