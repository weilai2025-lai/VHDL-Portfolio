`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ep/b2EDzYKbCYzumx+vSefD8bRpcqZGIzndnomubpOmxdjZUSC7t9kyG5vjMZWGr
QaifCN1f4Nhdl1SfFxslcpYQ0MK/ZUP7gD5AEawPLYz/0ie6XSUzUF6sSY8aSaZ7
ftxgRfjH434wu9JNHeDUamzV/EVavdbyBWCDyfxBsOwAzmP+3aZg9F2DZhdzgc7L
Tp8FcQphbGx8v17e0RmPMGboH55NBwQKWs1LdEpvG+NwtmqY+0Sq1EQRUoJq5CFP
GTpWhWTzAK7mm1iceTZdI2eDdeUNgxaGQuTiNMlCGqvzqQMeQ/gbccFc3LUPGzBj
Vb4cEq6wP5qDM6aNp7tP3VlOFkTYqU1xp7jp5Q5GeMlQtvCcp4h3Xqmu6vVhIK2U
LfapErEB1warvotlJCyn4hp4ZwvXlZd8p136Mrobh+OIZg+x8udq0FN6ph3ioEmR
swisDv+P8aBxBHxyI/C3edS8wHh+YkOzHJOMj0FEgO6i2dHCCuu6IYI0vOG7R8ZW
LIiYBmFA1Yc30yn6u+qGCE5xXetZWyzxj3dCEw2b7N3c+bCYIbdpzcE7JzbXZrUX
ja73FDM5aGUyDXzHVGqEmc1c1CldOJK4x0fZ2t8L1vk+7goR6hXkGNWcq6VA12HW
nBwLSfvo134UJ78Sv8s45nZel3XWkK52bkcQp3SwswXcH9rIP5MoIRwBx7+vzHI7
tUwTYyvNwL6/SpZk+vfDIFJC2hqi40ss+6I9gWu8vKrxnyTvE1QVXKk0RvbdBbbV
CcUpqNlVySwKk402eJdab3Z/LP/Ursk0ljy3EWcGR4yDTBNaeJw0Zdp1NTUnZz0l
`protect END_PROTECTED
