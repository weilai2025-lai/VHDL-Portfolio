`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYSnM/BSnwhbTKlFf/xl5zOMKkjBcFl9OxOT7kij/F4ntga0zEOSSc5rFWa510XU
R1MVG38VEmrd/g3xWcLsyLraOaAXk+56FWX6qJWvLkyxQ0d02Tw734M55PElbddV
xXVRyfTih0WjCDC7p1d2TiLN7n+//pFxSPHouIb8EyeQ5jYTsuAMi/ddJaLZKSvJ
BcQr0W9W847Arr17wJdkmSN4ZJcjT8FcxJUy7IKwduTucjOK0nK6NT0hZ+CrI8Hs
DAAxinefP/KlL1e59dt/YLNTU3p3LMrPuVIbMPkdayZnfzcalsFgelMuYJdq7WaP
uT/2ziv+wweFsDA4GWt7tD+XKhSbKTXli/EjYXu46meOhmEm4r3auOE+8t0y6End
GLlUHc3WAoIEO6/gxGj1z1BuDK5xa3d2pjqfddSKsp9k1780oFQrzliZjzbCdRV6
QVvV5cU1A8BZ5HnUy3AbR2vY3v7044Ix+y6PaxjlH+UGFMsCiVML4gI77Hh94lzG
E/udR8vWjZrYtplebaqwkhBS+n0ug9s819XLaBWmoXKsRy5UqzZ6dey04RqtN6l0
AmlS1r9ppsWUNtz02Qd8KyDaiaoSK4Aaa5+QT6KBpJBAw0pPXXu0wRt6pSbLQVWk
+8XHnQUT6a+TNXDv7E5AHZdnj0GFHAwnSrV/4e6oj9hAMlHajQ3kjreSdPD88Nxu
iOEjb+i7r7O3SMFmvGBVYj6p17L+KqJjOCL98g3s3zPuq5BHV7eJno1H2PtvodNM
FxCsZIjxxePrmZRa7AmFA1e1oh1HI0QGX8h8gfi1BkhBENkac2EGifd/y27c4/gD
vfcyCudYp6nL7MDFLkC/iFaLk7dETR8ZQTWm1UJoIfusABAAjBz2lWNAB7gYxk84
S7AQ219CLNEnKJCrHSxU1K+BvDo4F1FL004LjHQa76Xs+8CkgjM48tdzZwpzGs/u
X1RGIIxkhpAIuzIPq+4ab/rUznNeGJuvaOYITvW/+e4YyzQ03JMA4LMDWU0IhWcO
ThIat4vB3kryPXB56NS+62+9c60ww2QG2A/C3zgoxv8gEXPxYFqAgSOmyqW3A5hs
jqIgt+SMbbLrGsiNjI0C29ATA5E57c6Cb+LQHA329fMXKV/9ChxNhou1ZhBH/+JT
JdnAxsYJcSLfGtkdvIX7sSviHZ3jwQw8CdZEAe2zwB3WV0zPyCL4rNfXLsIaDqk5
oW3TuhjnNqrjwZZv4XlUKkKXRy8bIYOBT3DZBLc4VXXvEjbktiPZq6WFZKTf/qkp
v3FfvjRvrtfg0t+yO0pxeaRZ1EFk4quL7zwyccVQiOeEB7SSIRQ4YPpJ0C4ZkxZS
+kFIDucB5YR2XEGXxrq2BqiWLj+IoiyUkCGuWTq2wq5xHr8epxPoY3LyIk70Z+vA
uVW3JbfG17EFXj5k96UK5TFuJsyfkJBfMlSEWfqNxCGEvSIVsE1PeZBAV+nPymYI
5/keDIdDxUgXZzjU5QHGAH+sFk/pmpUT8pcPowf9waMV/B0h5lEkpipN3/l7fQjM
4qSbzNoJheQmjRFAlWGhGBw6q8chjUGg7MgMKgu62xJgus4SmALCwc3xI83HHeit
oIhXTOec7x+ij2iFFJ1AVfoxFy+KFZeonGMITn3taf980sMOF/wIks9bBs2E9dFq
YNcBlA1wlfwN1ILt2+WGGkVZ+ZmOCt6/NIM6JTvVC09MMUvztHCMMM6OvbuAwnFV
AHFvqjl+MECBtSwR0W+s0BbBRgldje4Hn+Dswi8KfYu7rtGrD9MRGwo//ngFm2qo
9uv1CDGd+zprhKKDoFNCAT25mRScRuITfa5t+qioFX5RMIILpLyXpGndkKsh84ga
fbkTWcQaLuaGDbG+zdeCgT+OmLTwJzu5JYbIR4emaouIIpHtG0zIkkGJt+9SvE5f
R140GywXxDYy4XVUA2ZivkYrBuL1lJhEozdp5p+AgjnFNn8jvl7L9SQYsDdDiOzT
rXXPfkR21sKQShZAmumFXDmq6CzqB3z4jBm6GM6xt+2tLWTNrHC3+5Loi2MCFYED
cwIsIUvIIbLlN3h8dsf5rt+lzD8RR1Nrjh5kzdURlMMPqpquAOj7T3BUdO48do69
CtruiCjJmQ4Rd2GcbcZDHLhnxFyAtALyLWyXJkrNIZtlv0GgqbzQuK9hTVrgMRuJ
9Tp+ehmafHwmtVv1Z6xBIJ5q5fdAxPMqnREEeb2v/Rs=
`protect END_PROTECTED
