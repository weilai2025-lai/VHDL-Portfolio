`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8r1utyO63imgoyyLqD7oa0kzpOY0bxwHLlKVH0HGl92y5FRh3dvzpv7I6OWPzUk
0cBLjg9Ff6NFtrU1kSHvmQ2r7MuqUWrwlfvuXUlUThVWSYTFb3+HH7emuA3LG/us
+8i6iaUGx8Q1pR4tZNfIpd4JYYUnpxBvbzjBuMuJ6yqUoHLhl+B186AkfghvNdB+
o/2gTRGm+pB6lhGO0AmYH/UAEBphb6GZus4muHk2MEeNSWBJlouFTg/YiPMUiwSb
nwEr1DyK/iNVBy9481bAu2H5U3eZPxBhuOeTbYQBIMmDHasA0GFef3JvpQWIkfqf
lzAZ0uJgYvRfCmwstwM6ErRPoDnTXCdab0Eg2fQqe13zcWzgSmAO7M5iBNZJ6o6O
5zs6RalUs/maarSCSWUOtCoe1C1rJXsX5Iennnqsh23VdclNSb9LcgbTFK0AlLGR
ySXa+p6vWCXkVZy57+WQUSvMFXxqZmmjkBQHlteJYafv0Ci+cWighz3nvVNg2Ei3
VjroTnvERE/G8ZQ4AvUtRmGeNcQdSe/Sb8AXi4MZIyilBFMc4x+pBvfxgiRuFuGi
WN2a1q4Lu0QN7Ryp6hODGpRb8ojQuFYWyDJss3bQqKf7UXR+c4rYPHpvTfHH9gp/
c0/h2iID8nm5luyT0/oSRIkiip6xTtXay+vj6AfUTvPo/0GHp5Pocl4a8yfbLsvq
+GYbHxpGLJ4ZoNiB7cSdP7iL5ekwV487PLtqNKaCnP4xRFCYp/01wIE6bAIvj2xQ
tcx6QkNqSZIA9KIVDFtk3TLyhqXTHUOS+5P0v+kSMpEpGmHlxaQFui5tfbEJpiSS
okXK83DymlwdnAM5kbgVmQIU8FibMRuAkFBjPJwADSK6GhPzqDcmIK1XknLUfgIo
vGRK5ZlQ+AxzXyRBdpgxZBq7npqCArG5onHM1Q6rA8axuoKX3TuSUE9okLDaIBdD
pzDdNxz++f/E1SxPH6Ynt8fkFRbvXh+ln1xxzfAbwoigmTaZkhRc7GkRzWX5PQDA
eL3iPU3UGl1G4jaeLCunMYclglj79muZ79XHzU1eTaayTTsNRWPqwfPo0kh/5rlL
dwsD3+PkhZDovdyr8SZNMXIS+b+GMRNQ+UHI5XFnrDrA2+XLsGh5a1ebpt+tDc7E
BhDYLzYPHIBTcCtHaLr9yXh/N3ejaxAcm2DON62XBIL6RE33pLSc0hHZJrnlR51R
GIkexkS6zgt619Hb8TKGol7JRp3kpmJnbfgcAk5KTi22AM+l7OHSyIk45sCEgSFH
R/bVeJBANXwH9coa2tkcE6ChaHWPjaRAqX2iHQ0g/lM/6Gftwea0F2tlf4usKW6G
ul5bzEGKwex7McG3g2GDESkrH/nY3YFmpOKvrfIVgJ+s7EOgLeJKlBgTBciWtEBj
nioCeZM1u+A6Cvcp43g2G+C8Kia+VCBEIsPmAytmREysxbcTMZ7nsndX9BMtLKbA
jDHAJXSIJJh5KVp4nUU2fbzhgztAAAO86rcbUqDq4PeredKWCGuaYWMlteay27W9
MiGWt9nRRysxUMSRk5uOGQ8gK3esT9lpj9Qg1iEckJ0gZaKNLfH8eN1gKsU6efQ4
44pFqc0ZN5cz+dWpTEgYBY2HdJHJwzfda2QSx70wrFEEHV3O3DzYis7Ixb6msGX2
LEsnOh1fJ8TEjRux+97PJYZ1dkEr/4BYoP47Z8VPmpSpfzJGQJlv6APxk1TQLFXP
RRcmodBWUdsOy74dYy53HgenwDuoVYloG8BjRPuNfRyr+Kg+p5CSHuPTn9sc1WLI
oeh0gRdr+hQLXwdjBtGBW3XRyPGt4NB/fw1bzI4/DflF4cRQcWwVKliF8aVjQAV+
ZYz6BH9N7FOYEFT1DEgrk/+ZOQRWcZmHf1Ffga45VrT0KFD9v7Lda9hirGwqmmG/
Nv6XGLt4TMBcdQKdAN5Z9dFOwwoMUMUh0CnG4fAblyqwzaBuhekL7qB65dEV0LWR
fbo6aMv+IXLwkjMZX3I14KxfLyo9JUSwVVWjpvPWXDSEf862tBgtWTYreVTHf3yX
ERxUIjUv8Yt1twrtIDQJ9hHiR6D0EggnUcY8e6OUr6puRy5A9d97ed3+rFnpK6OA
tIR3fuGH3mO5Xeeo1dYUHYAj7n7FdpeJhjDRuCnVN/4BkL6UEf06iiBap8qHHyNv
4v2SZfugswa7cEMRYP1rnNsUX44UlEEERaaJXwHXHzpRXyN9297NeX15Uo+06UC1
0kMo3ep8AZ20buLxSgihfJUeQUGjZp7ZFG03oB31trZaZH/DQkfpHgROxzgoElgI
xuUlQngGe9BVQRwem/si55bI+jnMxC7cSR3HSXFlRFoV/kMWTWr1Dtotv68afQPh
foGO89BQFWa/CltXboR//sRzlI7rO5NcDnACeDul4QDy4FgueG84jq/VYw+sTZlK
Ds+3mRC+Uu4Ui9ezZP65gZrZ1YETIEexW1U7GJrDSVxOZ9ILas/FKUQEo9FQ+HYs
AZbgYxnSP8wWQTF0srWwtu3JE7gFRma43WjfZ/dRwHjYeYV0jSCNm44eoeNIICMM
CcihaXjVARjvCEry6GPU8EDpTJTaKCD/XYezpefgIUq6Ga4uOWVPkXw1kKIPRI71
ioUmuPOu69KEjd4yan+pGGNPxtiwanJ2HtjpdZ84buQt7XJAhZEsAM0Z1tAZnJyy
+afW2+4HtqOI2ycyl2V1viY73NXS0xn3+AfOecppomKyH0ySfaAFkMHtmgZnGMWA
Q01ZeK1Toj2DzDNOyWhI5HG1n4O8FqYIyMoY2x7Ti04+/yQAutwwMMq1Mjw0HXmN
6R/HM/AuTtXAsoFIW29HAZ+462OOZgiI1LMRmEUFOFo8bvcb8hOK5DB2Y48Bf75x
Hp64TWznFCv9iAOAKSvBvA==
`protect END_PROTECTED
