`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ruZFpIgM6cFcPLZQmu4wK+LYYuZmeRKrMnyDDur74Eix/hxVcwKVqWh/3nQDZuX6
fHPx5CPm+RS2uz2UTzAkjRJmmeqvDf+Rxj4LhJyZpiearmqUOfyq3fY0x2ddUo5O
4+Ma/Y2wvC4mdpx7z6pGnoLWPjyZxtBFu8UHYPT/YHBTBjpjs33BGppVSIJNBVqc
2o3160SZVIYWtKYlx8WqmF2DvZIxLi5c7E7OAAyqtjdItkKpIAwtnOFjs6mU7C+X
s6AsVJqbS5tu5ZqYb/PzNhiSS0cdAAlIN0C3e/8xBCFtud5anXdIKdJHQmUzGYe5
KJCHCewIoUPP5C4GIIyHTjyXKC3bhgcLOq0WAqHmOqW9AL1M7eGsfGQVb5zNiYIY
mNDCVI8ePZx7bJIKxD9eO+xZ/dk+Bsi/hSSuQuNFfqVSKO2bWSbvv87Hx3dSlCPc
F6kldUx3GUpxpgTJsghVfbs4omT2N5dqDyhrEU1xptxw18+WCc/X3CRjV3hWtlkV
7S4wPm4xqOoa/Quq6NYasIelvCq33SXFaNjjZU73WlOFUaMZiTegxOCVfP31euDZ
/m5DQ6eZjJlJ446hSvY0sLnUk0O4NfPA1xGKs+x+b1oeCH04W8FO6rs6IQwtp6TF
IC8Ya7g7rVznkqAW9lQczicq+ZJZizdncbNVgJdrQefH/PJ/4A2/1PHoDUCHcfwQ
VVh0BUjZiV2qxLtx8lNvF9ZEi+jZ/Jul1gJ9FRat47p0nSZv0Tv3IlILKRz+Kg0V
wnIU1P9AaILMYOiYWeXXvqqn8jKghA7ihbbu7pa69oxrwW0fv9SD1mckPxyStAiK
tT5VzVFu7GHOCAmfXShDiHYPpEN/7Ko8rD+1n+KDdnHnz9IYSurlLWmYy1GEOqX1
8G78HcKY4z47fLsCu9leZOZzuh6ghmyXQuvH4SJN7gP1O+t+fA4MPFYHDegJhfS1
txLgItC/3jOIr9uqpkg2i0Jj7KxOLAmYkEJBa2aCAnyo1WDP12taZiTVbk6DGsX0
+LH28/1CrBd0YYFGvmRJ5f+hljMch3BNghOvBwdWgN9RhU67ZOwtTOGuKvbDi8Z6
lxkKTncCznGU7XbF4smMaqiz+6qD2PiFukwByl/dp+ieOCe3usjkdAcaQowHYI/h
hHwxPCDCbJhqdPiIrQSzhbU3nHFG0jmZ8QjukGSJnDx45vS7GTSdx28di/8DwiSu
ePov3bC3xxme2DVwJBXqriy/mxTgWx3Z/CMDN6pHC1S4vNhkEP1VlbkOv9I1Z8xr
TwtRNscr2h5KR/pyCrbqow8twzMGd09B+T5GqAYVzJqLn1DxDxq43xWta/uuxUTC
dp+7DWt7ORUYa/o4+iDY7543hFfQz3xD6me2srvmzypaNZ2trf8Ez1E7Mc5GpDCt
ORxV7niOrL3Uo0CYnF381s6UaT0ezNA1+rpXm3yLnxvZADV65FurrYnWO39GUx6V
LexSJVVHhqQgE2oIf5kKZle131Dd961pEugjaJlRhW4i8gY5gn23C67J2+L7m8pI
VGO1Pnu19w3NFjpNYjico5iKFXdY9SY/gx3IsXxVzE0hXl4xtRzsmvBBysd9n8p9
K3NiaXRUFG5vsChq96FvpWJ1J16ejQZIKzioUQ/HWYHg8Pn9w0AjP1IYK9zQj32v
Q/qPM2HHANA9NAHdFozouzu6psOqDgcbbgLSG6QnF3YGsIdyncpEWrh5PHF2w0JG
pIJKXdPsRRrEBtp1Q+/5S6j2feIiVsXCCABVhs8vmqhgQw8RDrPn3g6O2gwcgJUJ
rsfgjBnC2ay5rvPBlJrutObsA+a+1rPYnfZ7bkH+uTb7zBV+mraNaWLrpf0H5xyT
NrNm2Ge76JGxRG2zwNRQzsyAqrV9dUIlZv8iT++BPC2II+g6U/5qzjT5/DTlL4zZ
sZBFRKOnPllkxliRkPzWusxXlWjcX3nh0VFCIotXu89P+0hPRZrhlWqyzOda09DT
NevMEKfwtUCQVU/gm94K1O0KvrPXUDvCJasjnWMDYq/G8KXbaLt0SAGfvDuckZlK
S4bmfe4tgL4Ocv/+N0ZcoUfu2Hj9oTFHFlNs2L4KnHODRnqKtZmdXr3iS57O+797
8I1Ynbn+wJmYlJ8U+VoOp/LnI0ed/rfuSR+ji0cI2EEke/T89mEkexz8wz86hafS
brdKKlCtmzJGiIBEl65w531r5tGysrflOUKQOjrX77lPxWGu6cwM/9N7imF2FTMF
s84nFC+8H/0jD0OlmzpoVGSM8W/j+8NfQ9vUDhoUNECpUVBi4/TCT44jT4q3K9oO
leGu/SbFLqvo6KQs6Rr2ti0i2dT3C65PIrNmi/KWyuJN1W5VM+/4+vqthvTTZ9RG
+k2x4S7hKxBPHAQ+Spm7eSvbXgQiui/vo61qvizaElqhIh+8lA0wPPWKZYUxFrER
1n8/RO/A9DytwzQlYNctpldtWbtOTAa4wR5EEaHWxjQGVKlokyp9fR6KNw0n3gYw
YBm2q+XgQAkvx7uTFMcCiKhh2n+1i2+gAI2KPKq2X4g1sHAdCI0qG2LvZ0cYGHrm
5cRz6ejhbPaNv/6wxwS8vPPnk2dHX5rJ1+DgxKbp9ihapzKmZ0HjVVnDkKHy0bgM
raCFZ2qVT5iM4vnBDGQmDtMn4hvQdueD9bqVo3RbXMirVUHVjd149ZgKxWotMs4j
zM/1y9/h6XA2A8Yk6aLnzNIHorhPENJS25Eu4O35vGLpMewDQGViQ8Vp7pxuqQTC
jzLH3Zp7VSZBB8yUlYVbWJI/2Nbjm+htOUydI629/ahKDhWpWEgcdgDddCP+as5z
eKpgXvU8cuk3bDL/ncScRlF7pokS51FolciOjZPgz5FMDw7Tscu2V5lWeHa9EJrE
VLqTWCdxTzcW5sJ/DzQW+3sbairdQY88T8GdgHEFfL6CvxE7mBFVADAynUZ2O9Dn
ptN0dBYDxE6Vk8Z8kpDXPmaN+posBf/0LatjuH9QW9a2m22vtSEHJXNWn2p2Xvra
AzLRnTnMkMMrh7gLmx4UPtL2wUdFr06d98J8K6lU1Nyre1QsfE7ccLgWkPJ3Tonw
OdqfCdNA6P/z0qer12YARyJUKoQ+QXc/Rb5Du4iabYEFYAyDaDSNFmS8/xlVHGhh
sZl9L0h0chNaBk6fG2zgK4gS+b+9a5HSC4+4dhVsc5LsW5xRznac5yo4erx1a4P2
MygzTqi6OGd4Dzp2CGH/LLtTj9Ipdgi9D1fahuTg0FqVtJEKxlthrY7IsRx2fg77
9tzysdw1Kc9ycKcNsq7rte6YA8+KxAYgwfKSSA/plstYZZn6q5IJ4qNC5xI3i8jg
/DmPedcElY0yhLOJ/P/u+KFIPtD3MjBNpeokGNkgmveQU6WBuWyk/gtAV0QQo2VR
yN1Xh+eGQ4OQPVDcweTY04dlqA8uozy1Y5LYHjTXhYWGVh7ASFmFCYeIP5Bo4PVz
RDQJrBA3ALT6acSnXehKn87gTnSlQcaF47QC60WCKb9EomhQJ11CJQkdOtZQ4H02
zfpJM17Z4aGxzQxGbR7J8NgYSI3kGpoJ1Q8uBxQL7XFWphF/6VvSfRHwjnMaB+cP
7LinXOxaWT2fTxaZ/EgOEiSTsnHAJ1jQ9a11VXFC1UM1/bIELWVX6moOT/K5Ahiq
INpmSgmtaqugRUO3e5gRBsL2SGNKbyQMACftaUq8gamVTz6Yx0lS5+3TbkiE/fNk
HB2HRYVCQFxerwvGAXNBdfAe8Xip2nzjob41NcqHEaDM7/4dCQEyKBzft24WSQbx
lNvNCtwES4UxvrbklLa/qDJR5rT56DWkI3WUPl66GpEYuKptOpLBSZ0Za+usjV3q
Ulp32qCAKYdSrCj+KFe8EPeysgQEVSvpmPa606mMkk5K3pkaBIgWA7MKD9ilXS08
Sx57dHhHaSOZBO7KKnQW191d/xUS06+TIxIDCQGFopu0kDfyi1SM9d/hjiT4+Byq
MJcYjbQE9LfkzoyCS2KYAszxm3JL2Rj5JV3+NNgjKFcv0x5UJcai6pfybtnXdpFu
E0FRtNNydF5vIkQ/QS1Q1K6yjuxO6QQs4qOZ7kgUkQri0pmolLpspXJP3yxO/g9t
BtfXgAY3d7thDc2gv/MV6om4iEkURbZ/uGbIp+5Aoa6m4kITroMfMlfdPq1fDXKg
1kjJbSA+ZmQ7l8TGw5OpfD8xrDl8/1ymbfVHnrXj/FtgLpxuos/nFuCHqZeUI/+e
CKDmZNsm67ghBOZrdZlvn5vH2S891ky9IQSdIBHtODQBlZPEG2sctyNxKM5fIvGW
oPDVQFk8Mpqeos8SZ8oBqvCMWwqF1TNoPQuef7H/3qYX9DcR5Uvpxd4K9+81ARgt
EEkclVUP9LBd0XSvEYRRaf6O3UCrBZTdEYwFe0fnkcBGtY4ySOl4VLtWphJnX5gQ
E1x7a75LEDoWCYN9/plYRGvFdXWvevE4EtxxXT5IHIgylqis6yg67jm9maUt96ss
I5bncw0Lgi91Mg07h3OZJNBhJZWbNvXVETIDOGfv0d6eQbnyWtDk9u4zNebZhG4n
uM8i9z48KVYWRgOjwH+Ftd1AI84KKln2b3hbbu6EZrORGqxsuXgnGNQo4E+bFvix
yc2FaTj2tPOgkHUP7LDyD5HZ6wIMx4dwGfgvf23U4ETbkGDhJ6vI2MO6ykfv8T6H
vn2oInuyXcm4ox3T9xKy+00icWli1ebaaerCP75if4ZTWUmKLZH1VRIfwP3LxhQu
fB2FzWgfLKmCQy8zTs0VToUIei7I9MDVihfojxHJj9OHUabDQzayLszoQzyDj8Hb
X4MN0WFODX6qPiR5aYs+2uQVENG4iJ/RaocQNDqBwpjXyrk/08vQbsI3qNDLTBzm
nedYl5gBwY0qTvLTDtjBgnDZTjxa/+ZuuSrMAkmomJ0dFzEjQZ1xFQJEXP/dx5fR
CpZr9vVxF3ODQmCywz4peBQOeaoIq7ta5nfAxRRwtNLVBjpBGxmelN1jm4uBgl39
w3sBFef6Dm9CqDTJPrzOHgkQJtWiRgBMkLHVDuIrg1InFUX4hKgEWuKrqwXgCJOz
G1cT7/OnVYrgnL9uLso00TqE2Vf5ghpu6jXKmk0q1g4HZpZLLZr75O/llQt1YziM
lU3/N2qE7QiWhPdMLYUBvbTfWvqAW5AhF6JWFJyuXBqxyZvgzw5Ez4NrZrsXI8sy
hrsrQjigEiVRJM9xkG0AJueu7FuA5NakurHJ5Z0IOGxoZrDFKldrlndAV144LjH6
2OjRwOIsAZFuApN1OrOt9WdEHHqlVI4J1k6Ku3RFfZEwcCPDmKlOhl+jb/2MttD2
aSDVB1i/uD0xoWQ+VA4Zb+k0gm3bM//4xh1z11Xxy2qnKg36NTQlfP6mSKqCAQs+
s9IOUtl5jU8pyh+9jJYSqAW8xaQwAv4DrBfY6UZDCaAeAMGtws7+Ws4zNYC1z9mM
r54hR8dL3JJJLjIdBkoE/z8UsaqVwLEcmEA0LXI+vXsV9KRm6UOrSuIg5bZjhQAT
xWGG1RUl0ciHlJ8YfZfkTC1m7c4dVR6+Ag9kkMttzkTzv3oAGzyAIUw4+KyymT8O
kqmJlyuujnCAt1HE63AnkrIn7yNQ7AZeDxX793X+XxWWEQzlbKKtcU8SdaU/vcd5
Za0IgxrdIgxuuVTyPFxDxuqgl3OQPHJmo/eeM34oCHpkGAyYnMRodO+/iJmSTFso
1EvnTlCDu/bqP2yy754IWp4nl3YhWQ5yTG/4INDKc4DzYb/iMOR+uixjjSgicXw9
jg6XTUuWyOvIlF9wWrkpJjfr9xqDFOpzb78cok83r+ZGTMNEHZdHjmiwPq5sDJTq
R3oL9TqXJzXC2kHYU+kROXFQjOiiGbvguJo5p5kd+iMfGItg6wEB1EAo7Y73lJMR
8uT1WWNs3aClKmaUi+26GQnkDmcMMvI6GXESYahpdNkVPTE+YEJbtEj5+IkBTaKY
DD0WL2KtF6Z1kiLMxVTu1Tq1oR+fXkxMIAqHJTxHY6YziM0NBkiZp3skI4pHQLPi
peNClc1MWw86c2wRJpLKDYaMlYabWPlc2AVZve14X1J1vfy2tw8E63u4Vsmn8eVQ
5tW+G3/aCUDr1jfFg1lh3MW+/Ye+j3KY+ct50A5B1lZRzF8Tq2umqrNGMwnHdM1K
a8v8BaVdDW26jtrm5oSZJF4HyWx+Lgqnc2YA6T8laDoMzEDpVGesAzyBCDH8cZMt
AF5j6C1nOLKkv8lsL7hrXZC0P9VE52YmVSRf1go6FhjMy9Sr9QLz7h3heSYDMrZp
sNs9pkqpBNLXPrTst1HeO6CTvs3h/LV7JP036zmKkxAq5Rrkv+HdsIeS2YSQ/XBq
eYUjfZDYgkPDEx/pwGm8I9BNp0eJZDI/Bpvo0QWQVRcjfavwhv96fbdJjLwkgJ/A
JCRJM2ldgdpOYUsk/6vK244p/5BlZfaB4YMQCRK20kr9S6WUXe2NsKnFmheUoNbt
g98zGV1jsbJeWfIxDU/Tz75U3PHTrT7LOQ9dQExHlwGbVkkrfOAaNvn2chjlN7xt
8XvCNtavG4z6BvjH+HsWfL7vMjd2zvQyDmlG/z11f4bfz95Nl5Zq5lmpejlqF2Tk
HOQgEzPmMydHYDXWP9XIJIh0HgzKPGQb5M6sjCSxvq0ieR31O+870hBiRG4Z0FXf
ftScVSQrWZ7dn5TzheZlKZhOsM0JHUGr0tZRGIUQksInR+BQgoIsZdHDP2FtyktE
AKGHrTPG/PokTDYBRhgZobzFK2xFC6ho6Owd0ev1M0wNee6eKAz5gtG9nJzl1sVQ
Ym2jNAs5ltFEAd8C2lbZVFHlzRrQWHLYydGeQZ9VLwTaHpvDzpKGfsXL9AKVrU2/
nPVKYNA7pUz/a4QyaRcGzw4hxcnHjBIXeDODpEmcS9rxBxdRFxYxv0GrnKJ/UI7t
rlVMCNEDyGRFjY87Ohx3Jl5SYQfMMMunZALqiO7GTmL89xnf5VxQyekkkxB/ERpo
bVO1apQdV1+zIuJqehiu/zeVjrJO0vEtqUdGFJIWUzClov31sbS3kuUcAOnAofvJ
cEV2jxvGYq5elxVhXyuA1YRFZtMNsGG6/2YKwhfEXIj8gvPgOONk2/a3wwNAVsk/
dj8DJjiVp6ZBuCPLgb87Ua3CNI9FZg+v0TzPuhWxHv0kyAybRNWkr/vsPovW5e4D
ypbOudgsIBNULkdW1hSH+K4ExtpjIaOGz0nVjYnsWpSFl5/VdEhpWBfFknqHCW4o
D5YN/7HJ3u+4NYVrC4znI+um3N8Bz4pZgdqgR8Ex0JkNj56T2qXK+bOQWzK4U9yf
ckJ/wtNGWBGXAG8JqLqX87UZuGPDDsU4N1pkmg9d0eS3wNoVqSn6najouceK671O
TMf9jkc/4HR5tP1I3SwrzNxJaEtR4mUsxQp0iRD1a6N/GxpagYzvz1PtVD3RcdAX
9UeCZ6Yg2OtYIAArVR29NSStrqHThLcEfwRj7Ehc9JCy/9layNvpkLCCHVm81cqR
W/6jnYtnQJ5EHtB6BQ0EeTLGj/vyRpLdeOsJJN4c0G4Ty8EtuqOqfjsxIzJ/TFMc
uiBkKOmluOZ+7Btb7crFQzFCYX09cWYN7kVYCIYix/uEfWQL7Oab573lOlqvuiJ4
pj69PzvFh8l2Q0gMqG8lgxWbSInDzyStDL/Nq5+8xexhAoTF/wmtvNwrtouZo/L1
yuXu2Ogj13hMaDwe//7JSE5t08safKm8uh8E74N1TPEHYGk3zUpVO9DYkvZZupOf
esHc6tFsaHDdXRJAyInWsBn3FJSAAjx8ifuNATbKNgS0XbKtMLi2E5UD/QqKMdeP
HzcCS6fFFqBtOaiyjRJg3WHRWiKJPN4if5T6jPqJaUOsaJKzdLx+kG2LTiIllpy0
inKQf+jqUa5/S/stIOAIkUgkuLV3VqYWrQbkXIhZ39V4eESs9l+9sZtPsTsFxgHP
6AYunXHgLAPel8MRG/VxFAbGoZdzk71l+2Uq0gDH9+uqMxZ+Rxuqas6pe6Dp537r
kBbfs7pVwS7Ha1/w+YtrEe6ppngMogAbRvNvP3rU0Rs5vGNhG6bq4gBZLMm4ooPA
UtsHiH/a+I32b1ZOhsgHWsH3yAIH2LPYITRjO5tH33ZzJ93zwthC4GfLmK9/Sn7j
QsQCBq0fILk2nTz5MUL4QMOXwGmCqSvF8tw1V3oa3cUFVgwzXY8lCtgypbDdwo1G
BUPKGW49MuE2nIDZf6vQcLVoZEsY5xnPB/b4lnlwiFBEXClT6ttzbG1T8n48XNVw
rQApM0EIIaVo49XE887c8Yl1Wx+idIv7viY3scrgDmaLqwtAvRJglkXCvlkg3Qzg
15CpSFgBmj1BKm//VF0dxYkAbOTmpJKZPzERg0UkFdKgfhkbSwilDqEQyaRDcOat
nw3fKOPcc3kyE9PrmDOjYrdMBoPhGZLB4GRCwG2Iqzpoptc8KgJMsvsOLa75ipH4
ohbwj6ye2Nz0MgaKCYp88nbEa+pw+nVllMEVVO4oNiqTNgqTaIN/ZpevZiNv2AN3
5/i3fjIvzID5rXIfOpA7d8maiWqOEyVS7UuUl+YsCGJVn2EvQL8kF4PnpgzgaB0o
SKW6MvjN3zQB/yEawK8AxBs/MBT0nnQuTEiz3WcZ7uqt65Tjy5YTzX5MrvHM0I2b
qpN2XVpRpunp7p3BpkbBiu7WaN/y6EufEd1Md+W+F+L8SA5huO1MVGEoDPywRNmi
Lv8bTV4uq6lya74am0tvm2VKoediNErFMj/Q2GSkmA6T+jG1e9mfbtSskqNUuJM+
6LE3Wl+6ArgZmlpcCjYnJXZ07DYo0XYAUdZDeNHjkv99RBG4x5QsVn3GAN/KxQUe
EzM7QhlTErBK2Uu6OQaMiT8coXwPVKbXYTxwlR6wbrrmb0Cm4x92eIXgFD50J315
iM3RWUD2Fzl2wTqV4pb4iJoRVe5Q2eABu+vbfqItWy+53ylgtwAtoIMNPbwUClmj
2U16N6MEcHXONehfZlbfLAKTPMgU8TiNAfvwMwPqslfwBK6WLKrSv5rEfDWpHICq
9t6lOaMvNEPUdaRKvqsukTv85QCnmLQhqkkDDqSKeUkmRwjPwQqvTob5NTUfvoA5
gS1+lMWbCL/09Mn62J22rvh5ae1tzGXlvwie0XundLvJ/tDOcEv649IZSAlwSXtx
QTdrqziTaSCJjGFpAVX++tbTtfhTFkTCEAiBgfU3xrXNtctNJtXZLQkMG3VNVSwq
4dsV7EzwRn4MsW4Pbp8fwuspV+5ZysC0wwDZcfw631XwWeCTjBx3/9MHJWGhWwBW
rMdiecIEPIfYrEwcXzdm+JCiFCAs9Wt90FbpzcCJjl2w1qDaGVk4E7nPu8eOY6mR
kH+hM/Z2NjbkFYKcu3PC1affaCD1Y8n3itV4jUNv7Mf9S6mQnpaK6nnx1d0eih4d
1lugkFh4qv/PeDlfcjqhBVipjT/6b7n8WFIFcFquGf53fpZmg3LVE+DNb6KfbPUx
n1BjMGhA2rb707RkfiwdpSlK7nm7aMJ0qbeX7kr5FvOgoqp49F4N/kyAXucesDmG
ml4W9qGsAmocSuKmODAmVtH8bKkGv3pGF1UAQ3dT+yZj3ssWUN//Pisu7frqy4QB
oLXqFRdvsr40VUYuSH3OgmvTIJYWydEyyNaiJSuZMBvN2ExUnWeyw8d/HuJLnluu
CUhNMvmIZ9CjLthPYEZCkmOXnwgmUHu4SVo5BLzxfixwhlkKagM6s6dLjBgIVfRi
Tenyj96COIRpvLWifYyOojFDw3uYalHn85Lu3zGkZaFurqIZ0HjT1IUBfksYZJFe
7DFWrC83RzRsiX5SPIFaRRQPwjU1q3ZVbmmX8w4QpO1N2zWovF99B6Juz878XMVV
EpXcwVlFKbap/HEf3K7Ooxw22jlunrYMapEZHXLUh+guObf0Prt2FzVcOKev5nu8
GgaK26SKkZxoh+Hu0C5Hl4S27s66iDFIjNDs/rfmQqwNKsZE+HJAbn3ctTTV9J+0
urO8r+TKmxYZcrV3CLV35PdUwSkJ18xGcsYeJMFrZVS8cH4iGf8eC/gApQPZepQO
QHnNk+c+diIuoB0uBWEp4sE7y1jpQyJU9u8tZd/KN3V++lKsiBFLQCHTCGMNy0rF
RQeuJjNKR8VeRVBNHCpNE+8dvVs5xr48gtLwYAvMsatU8jvenhA4L+TTnvCNjrdX
2aakXLzGFl4LvAXtjLGIMUCGbqaCoHFjSz/v8O9fcpV3/7JBsev3uXd9uk349aMU
TA8MsYoAoEPgTU58vAa6i5lqqJtbe82787A9aCTMWJ+8x9dN0JWnWcrIKPAAQK/1
ETw1Z+XJTeNFKZJmn+fAecRWrxMLeiWO9yQoV07Wr6GzCkJr0YJJY5LePFKHJSGU
NzANyCi4m6vkITdnZN3y+z7v1OIzf4UkMCRBvxoRc1hwaOqToxlTms/wIWQTYj+4
x4XfKpVo2VpEfAs5Pvq7Lb0ff896/TzPN1nqADMqY+ZIHcscntydW+AQe+Xx8It8
PtRGaR/WVZpfAENNjfRMhZ7ycodLIuRDJEZZyb1bioC3FTWN5856QU6bAv4xR8Mc
sjK5UhHErOq01xMfJLGGIn08QSeGpttE2odSDKOi7cWobIH28ra3BX+Zh8YD2QWq
cY9Pe9mwlKqF4r0cCUL9iAGBzCeHwtymfknBDKo5qlBBR2t/O+hVHAj03M22Kbm1
kqy8QTwqtWUwCymQBl+bbcK9pWhBWrqn/mwsJtRDuHeE+UgJeYiCWvYIfJ3wsiFl
p8Trlv2GC5p2yAbYZPeQoSYHb66j04SIUFCM/epl39+QXW2t3dRAYEfPFm9qigCC
kLCcHR+Vn85hbnmdfRVaxxNQZnjb2wcV3qnbUPlakiXmZ6FxO9Z06DAVOasls5F6
lxJMwsRSzO/MLTGx1qGUF6xakOvZwuwOvv1CIK13AJ5MA78Z4hAytepfXl+ebsAy
x4fAM4jx/aB/xTqF3Vt7yc66KSi6aQKvRjkrHaSEKIkZT87Rn2eNHuioiTMI3LLx
+jzyhSnogSokB79ycLnfxRfcqSYlt+RJ7d5SyUtOvjykob4749JB7bglJM6TiVzx
VEX9vMoZS8QMX/+TEqn4bBEKZRs/IEVulLRgrA+SbHIMJoshvb63KWU9JFPeVweE
f3INxoVbjYrgpsv58d+Lulm3G5uBcEk9A54ziWHtAiqleYezIqeHbD16mhw935Sz
KR+z64ziYqzpKhIDQkoiDNKHCS9DLMJt43bP//qLt/6x/4kdiBmV5c/i3JMNIMe2
CoJrp/18w2ndrYYuVBMIMGYuRrD7fIZaACblUsY04ungKT/PsyyfxxQxeHrU0AFd
8g1vQKeuna9R7GR7D5fhpcsmaBJJLVwUgNRXF2cAf6F9KYvKu2yfIVI5w0EQoo/J
I6o9reQhukI5bp1dIlLJVCQutjxs9R333cq5B3/6CW7qqeuiEyWKOsB0W/h/bCVk
UxC6ieN9uRa9sQdoGP+oXpsupQzqOAoUzyrWD09VfjVFOAtsDrOPEo/PpzGsikFy
2jBPA2dE0NekORIRYzW/naJ1KUMe2c7GQn9PNh/iA7XdpnuY0uiWFz0V2esZrfTK
V1SCtlZ9Dx4mUBZlO6ibV4c7qFIIrLC0qL/Fh4GrMAyilHPn2zqGRnrhgjmj+wGS
f/gsFtT3k8CT4awXN3DV/DoSA5InX/N2KyLdar7tbsZ/q81CcklSEBz1ml9mpJV7
2AFLjyHHR74LMtnpWG8nJ126CBhjn15YiFr+Cok2mgQ31VdqhRaVlbkmoIxYQ3dZ
2XFWcX32sOUB9oxsWOrRB2JywhXktD++l9I/0LyoY5odRyeol5Go3fefRpeB5Xq7
XZ+6/z+WTmtkqtEFMruNmuUnwuS52rOYMUBgN+cwmjLVwUzIvi+0xiSrTKLVrIDU
4eYweYUQmEjhcr14Hy1wTJ49orn1BHKTgpuonzS2KOTPkZXeXurrTxTPxImubvJP
ddV570AuUeHGXcSDYnSJs8K/y4aHZvIWzRGhdWxVS5K//rKN9UjgJ1H3kjqBRrQ+
e/Xg3dAZcArXLP9ELkJapiuo6ZkjdOMKs/WbL9J0JvZlm3ReK8vDJMg31fuQGJDZ
PMO0VpHO0/by7+9g1rfOR7byPiKn7r6mArR2c+nCdDbBfV4JV+vMhDx0IBnFa3lC
CEkbrJS8/cyV43r9q87Iv5L6DufofaRVMlbzbLD0ESyrL+6NiNE7MRIJRV5X/dmG
x3Z4O0jrNScjp/cOEwNbf+7ESimVdCHDLkLVowYlptVeDIRUbMqO08Kdf/ZEHV0L
u+g4p/LvhM8svtoPJfabYGjDnebQv23ivmL0kiZUXgFgZz7WS0mesG2W+bH27E2v
kXPMggIRk2oKTY7A31pEbBZwrVW6pHoA1UWXrbmYZUnsj1OD9G9vRjbrMYnmRDLD
0VqtxIB/ZtyPBDCEeP8B77Wzh0Pcy7vcjeQqU98EbICdLxyNO1QV4nf0ZUPak7KG
xI4gMB1qj5s20Av5ULrfcL7ZQCweB9Rgkan9J/qMzu9N/WPqte6TlnKSqbQjM1y7
NFt7cTD2RJt0QmgvODaYiRHvkAl3WWI9tqv0/tr1fxlu7SLUY+Qvumfzd4bcls9S
G8eJMmfAGHsft9rWlRJuMbj10Okjs7yz1nbIvDA4kkXY7m7fKN4tDdE+UepDc/ft
CxXX0bT2VQygsVt/lvSKo4wzPaLA4oqjG9WzZeG2cUqt5F8NVcuWY7pVvsZ5wNQ/
wiJekan4frwqoUXDYjkZDQPW7oO0rPnGzZxgw0EXehBJlfcQPGh7dWLHrK3Rcz54
uSEtZB/pN9s1aOkiCBDfZk8qcbXFTyILN77MW6XZuouvw2boy1AymmvMJ+HabRW8
UGcmtRKtkLhl53x70p3Np8miY8iccuhTf3UH0vC0+nucRQ6nVLI0dcJrQgZqHrwB
Jr2NvXwMdK+/LC/EV78yczuiLgGddVakXs+jqPieWEYb7EdUpb9vB7/Qtvxxqqkb
yTNiisImd4aVwAzIbBGHnqhy4214DZei814h6JtYk+1tMlLq2aAuKekxXh2S0Icn
dkxjlnRa7Tw6Px6mPK2og4pDNpqh9GuzIFHUPn6ALdrrwwrmQI861LcWDraz7oHT
58aTMFDjKsdx3FLcss5mFkSbB0OYoRuakKlBsrb7aAtGyHdhEMWavS9cOU9yOJ8H
wopkFFL/iNnP5y5O92d/sO69cbojB+XRKUCiUQLnMt6jAeY7MWuLcZSQtnnTaL0D
vZJapKAWzp2o0SqtGO/Hw/isPkACrGfYIhpf1c1fdAtamXifE9/12UDvc/fxgwIP
zOMkMQ9O5mg2sQE68rwQM9eiRJdhox+5lcs7LkvvAX/rNk1Wub+AL31Ldk4LkrJT
CCsLhyTQOWMZpi6NOHf8+Sg+Y65K4lSvGJb0tAw788gH2HLzTaZdSDOBWdYkiNCO
51QVSdsYP4mrr8N1BE+W6BswhPOQ6YqRmy+QNCiNCUoZwgtOy14jDyGb/OoXf2sU
8AQrf+SdJLyiXUHZ5Olz7wk2whVxPQNnIxTJslIIBh0hhBZtbBBk/8nIxLBe99rb
njOgu0KhQiDuRJ2wt0jeN5nUMHYEO3wzZsuLEEZaEQ5n4cxeI+vVsOd/3v+Z8NKI
Ca6IOE/l9+3sgrFXwsZqDsqJz+kc9gSXqumqJkWqJBbIfOSXWaIbn3vkH6GypK6U
JmothrJCmApfO1YAE+KufjxwEwqiMihPEuqMcefkf5dUhDRbDNY4mYt1wzozjp1Z
TWjbvSLOXlZ+gDitZfDskyaulo2Qdk4d1TYQOO5x9BC8X5IiA3adIuLq/jEWAXwA
HAtAdtETOu0VY6N89Ghh0YGVsqlxHdjs4u0sBUVxudIN+ccTheDN72dsInq0MVOB
pfW16iC0KiRnmaL+5T8jd91AjgQTDA4gmZRA8YQ8oWyY9WIxiiK1wjDFmY4cp9H2
nhNblmGOg2kRBK/8v+Y0hXBKlVbW9g+7zYZvkAJx+txz9val1pYm1CD91rwYd4Dv
ezGqd/g8Ufk2jpfxoHHnaJQ/euN+q9l4nCpQDtWBB8j6oOL5KVDlaz++If8TQic2
xuZMWl96LQCE/ck0eAbATvyUNgp/lznZxWFS9XPw1k9nM1a9cYSwas/DXObAM4tl
WmL5wYCqo2qXqg4qyudKPD4at3TKMx+hqGN45FLawtonqpxrDFS+JPKC9nqPISVD
AMH1dfAKyrUdE9hOY0SkwU0EIfcowuiz7q/fidCp/5acZjdMUOldVZqB39Cx2Tbl
RXb4gbUZUhMJJtAAsfGv3ljiNQ8axkXItus7qak66+tYQqXDK0NufYyDboWwWQhb
HC60l2qKCm8FdxcwJoUJPAkGe7wwm8I5oJdTU2hfSJK3msCePVjBj+/Lz8B42N/X
a0ciDi9pu+hVGxfFP0/lcMTWY9/oHsH+kXEEB3ImyBsu+XnjCw1Wr6xsVriJGa/H
IdhygNN/uka3Q9KpKlIXuGE2HApifEd+U5vZd+NnaYV/BGWWMByZ399Qn/H/Ud0w
JNAu898RwMv74zrCRtHPYfTTiWcl2oBUpFDcBEdNPEfmdYlJbL1VSv0CCvdyjNW3
vSrAL7i/AQkuNiytNaDx9gYxfmyEszNtgTobbLw5j6omrvzXdx41NmhjxwppPczL
UgoVesV6+RZXAguU1g3qrdw1P8cKT1d7IBgagukE5Zf//lQ8wcYRAc/LngxOMcyJ
K8ECsTVzTl9zGZQJdqVIo6UpGaLxn1rXMnoUVkzlVjd3bv73RYqHKMHCR6YMiD7A
NQJADS5xryEpTW0njE7NoNIWFGFqhfD+vHeNZmWdnhlJJb9lnbQeWiA7THj8Jmx2
wcnEm+B6tbX3HGxyewd8mJeW5TBVofg0lU7ua4oEGR2SFPzwC7gFLsmV3X8T/a5e
2ednkpZfYKSeP7OAkHinTlgI2wzlrsZg/Cw8P0hjRA1DATnkHkqMSqN51+Iy1uZB
1mhxHuKAP1dhivz7omCVXvlmPazwN03SaD1n4ZTjAns/xOMZr8aatc2c7dh0uMXF
TUTMx6ichmpw+bszw1hPDh3bY3TgURqSQ0WHmuLxCPbyNKqJtRz9SSe5gO4cTtCm
FWwaoRK4I/qcMEb17YiBQm2mB4W7BiymPKDJZEcBhhU+RPrKhFXE5qXKvAhDZ8Ir
tap0hMyt4emuAyH286cFw3OCZ+VQEQ2hnsV3Bil3nVzG1W6N42fyFU3maKJMkybw
dIggy8Z29bcojUUMX5yF8zoZpzt+x26n7tZ5XHr8O8izYhH8AFy80+Ty2bSgTo9T
iPWCmhTck9B7f4XcD+0q4wRgRl90N5GFMYVAt4eJJc5QUg3EuOk7BekZOwDOJYaL
hqzSsK52TftU2TGv+QHU+mqByk/2TGuOPV05qcpxJgXwASxEAQtldBFKx6lq+xk/
94KEOUlifJlL+fhe6HhEc0234okfOYjrKQuZHjQVW7X1JdEQJWWV43H9ZoPKBc+t
dU5FSKalAkyv8e6clQC4xBnl4q2UbVlJ0QXegoql0O8gxv5sOyjEDguFKhpeQMfY
D8mrfD49h6ow/LgMVECGR9hdkXZoP70CpSR+dvQHA2cRu/6+bYWZETBB0iO22rX7
hnjUAPhRd0Q5QuHH1gRxyoLuSqTFsRXZ+rN6X3LFyNajeDag/IhDZaemaDxKd105
wK8tHJaJLPAh5Cqb8bDiHC3dhZY+tFBc8cJJvmnhi2mNaLOymu4c2ehF9NV0lLhF
boUBibuduf9UdIli/D6wnN0wv3BV9064g9BgoU2MCem5C9KOOz2Pfak2Cehs+CjE
e/WTi7JgSLOrKSOIrTr7L4vL7tgKpIPcey64hL0yqcZuWM+nqFiCjuLhsv0Jp6jy
TgeCUhOiCw33E//09yntzg5QvbL0rNwGllCECpf5Lue/HK1exJ5Z/G0pAYvfkRsk
7ZEDFAxQCidncMEUSNGL9oQ/Py0GLvWpcyer+pTHM783s5wRG1pcz/Cn/XbTkgVy
uX02TqfHCOw3VgHn/KKAaY8CQHNIAHk7VQfdolli0eOh1TqZajQoWju5MknILNYJ
LNr1jBIUOTBS6hZWM0LanHgMyWGViTywlG+DrgVs48Kyc/pPJBgFy+c2c3U7aDwb
FCrvQpZHPvQXYsa+CFaNnZhbeejrYE4Stdj37nmWG+mohhLesEKHQcM7X75YcYWU
aOVrnZwuLp/4WV3ILaQbFz7L599hb6XCoQ7Ry/gfiIhq4DAAJwQykWxJmK63t8cx
aV+eWBYnBYxyi+xfOTIsK1ROITkigKDRiNnUSJ+Tk6ONXRfWaOGn5felweQHOkKT
BzkGPtmflx872jV19IFBAAMzT2eKznHoQuSmNmCrGTANMXpJXIpJ9fj6RbCxnHqF
nDsjAQ9bRsb/epssneaapaVGT+qe/ALa6ggt8AHMYND+AA7QsljTxL7JmBuMX76h
RVO7FJsouFMdFup9jAWp+MCj1P5dFVMN1okworGbfsK0Kkaexh9U/GYcv7e7I8x6
+rWSSIcstZ4k4jTIDD0x3L1Ic/srkAzg9QAPoMsyOeB6/W1yezcBcxA07PMCcv8B
DoFg+3crE8rY4ewY58MP1UT7YhXP9QNEEq0kVBF6ywTTao8deNU3Fv4S59Yy4uwv
0G+f6KKLRzdnFfsqlsh+nJTYvOjsex+7dgk8MFQ0efMQa9MKm5wDEsVBl3JCgz5a
HBonROJLK4RDADQqvCM7SnfPO9glgfsJnxGoywkEDjE41ahASgAkF2OXI6qagiBK
8BiWK6fjLwCGCUSOkUXh2DHDvvB1cC3zLVoCTvITYbatsjubr1Ug8/cvrRbBgbO9
IsDhTFDUEClDLqucxtnrlrXH/IM0JHAjuWf6YL7jtHMda74o2cqB2FxAFqqc29l4
NgdGHG3NStDQhybBt8fplADM0e+jewYokBGS59fNWMnSQ0zboLw9eCbLCs8uhRur
4L5eBjyALzIPzSxdbvZz8XVDgEQ25bPtbvHnulNH/L2/C7xrFa4hj8Eaw9O/rSh2
Cavbi0oJxdqQf2ISyonlST23MbUia9DZ5XWUQ++nv2gXTJzc8kfNVHCdNLK5ykWe
WrLO3OsLInVfjJe2km/ektKRn9Tm0rsQLqbhjUOcg7jF5Gg19PGSW0Uz96yVhh2v
Lm6Us1rKnx7+cp7TRfN8ju7wLFpBL2AHD+VjVlzp91DIlh6PIlndsQHj2B42XFLX
NXDE6LiWEt/K1xOTeSlYMm0pkIz/o/DGwEPTwBAuS9rFTRvYCsGacrpYap9LbQws
zb/HIX2AiqTx5JsQd3My4+nUHph3G5WplU/q7skfGVlYqLxTzxSzhe14ylpzU8wt
a+zBZquO3+9Eyh7la8gxey+57x+0yb+eq7poO/lRuPai2Ufs/N+wJDizPv5UZIVp
DVADrO3EOxGPk+gAiCn28RqbMP19YcfaQxQL4p8Xy3oGj0vjcjHR3z6pcQvNMNur
dQoDReKgwQtjg2Bx2Jzvg7EShNnTCSe3Mzc87tVabYdprXbzPUKNs3XR1dVPSNWn
eTQiLBjLwKvFNY84PH98SYZg+WYhN2yq43qPs4cfqh2iOdKP5UNDWkmn6vwJvx76
I1En258owsMJmdfU++xv3a1MTe/6HAPe6CTCKAWdf6ZUdpXrzfqtGLHHsJpKhq71
Yx25MSlTRum/66tviim49LCuKR6ReekT1DnG9gyMzZjBsz6zdO+ZHuNRgi4A/yG3
1/C3wH4iNdkjS12i9SrOfgjj5AC9mZrIgLoR0boMdBEecz4SwXjADYHWcpPdx+xa
yc95Q+xwaSooZjcuV/k9Pqhvj58Spk2OS9Wuj3f5luAU2fWdlfeXuEGRl+1uITxC
tuYOTCLGuNCrf4h+Chr3W4lVyHqJ06jdy3/llHI4iK1hWRHuuQZihYbXWqH+6dGx
ZKOn+kf2IttzM2wCbu004k7Jw0dScaLxhQ1EUHQd9Tn/GkxUJz2MaSpsPqDi5t1W
vZQ0X0ZNk/udnfWmZo5CTpDMlvAY6uPDzgw8AAkAZPKcHzApQ5gW7Ux0pgGrdxu5
NKEH6OUeYboVBcEDMhfXA3wwXaD43/QDeNHTeVNwJC5U86lYz8u6A7vW+BEJW33/
1TE8YXVB4yGrj5JUsumGXL97vRpA8cSRYP8y0LCzIK0ScncPJTECJKWHPs2VtJcj
DWZvmOU6Aw5kwbc1jD3rHpf/rRaemFl1cv8z7R0vFfAbMQcAFNR4w7tRbLbjVRp/
ghyP/OIiFdBWLGi8uxffy4d8WnSozswC1RsifdeuPKhYjtU+5uKQSV0HZPP1CCgK
IrzNpUOBdR+BSNnNAInbCI3laund3vZVPQxmDFPdns8cbVxWAKE8nEm8cUOqrSmF
zrpIBfJAUgcNpelgyZeh71sKRYA9XoxTJdLgWLKnc4mWeUQvM+mhk2cHk059XAjn
VMxoZysr0VeBq0sQvMlr0YBQZh6Nz0uDxouciuW0i9wRl4vdx8s17wmZh6nIq6xb
WLzS32oZZMU8GboR2jgqtl+nt44Hw2oKsPzIXecplZWvL7YZdZrLMHaiDdmmTt/a
wgOyI24WvmxtFVTV3hcLD17U+yPTskNFnLBoElUxoVS1/ZpEJIxxFTvQBWInQ7eb
b6YMj9EdgkdjFOODABb7y2wsp9Z0xMj84jL0hwP8Omqq5HCTlPPUKYyjlObmdSEQ
4fgv/GZhb4JdylTMDapJK37x/+ke36u/qUml/jo7UD168I7LLZZQLd6BBlRayZcC
vWDHljAxjHq0rnpH9qes0Zpgou4qHjeZYDeh3SAVy+cIjfrYgfpsyAazq4km59dV
hr3pRDtyAH+Y3DFE9VMPaqYF7o3ZawhsraYJwHVNE/UnbJLcBpYI1HTdF3X+fZ3E
JIRdrHa6/Kfy82WZYPpwpal5+huEuGypTxSgWv2+YxZi78pcApoyaw5iYbIIn9hM
1AR5gKWSSs35LvwAXkA8oBJX0nkLZi8b2Nm9mH9HfaU8r3ovPhJMvI4eJ5NvV0Dm
dvTuyA0u5U9C82JG/VmjmDbnJen/nDAitROjfUylia0DpNnqGE9/+v52UZwSoF1p
qd8dYipPqWIcyfMxrcgWbUp5h/euuMbx5GXGNoVfA/uU3AfGGI0OlfN0oMPlwSKo
a9APkvFtbLD9qqfab1oMtm31BYZopXQnb/DaauD+gEEElIm7Z6EH0ERS3YmhEeLH
Kbt/2Vf4tyLAgwvBpYTfSwosMo7EpZ5P4DweQwA3IwY0iomC8ex7Fphh1w6X1zd+
/7+JkGFeyB8pqub/HOFyMVce5e/v+CwfBw2TTiOjQgQY0KP5gwxcCt5AdFipQYTx
qy1YF/4mUJr38MovJStfMD+gvEmWFVZzYY/3ijNlu/ygYCl+tsdAcnivNuxxtxC8
mMJb4tx+hn9O2Boq6A9FLFLDnGj1Vjs+B4c3jB8lcjZi4+lSVmczyRJ0FZoscDYm
3PhnCNBLL2vypazvQjEe9kCxsqLzaorB2ubWZCdaUwVuAJ3SW6mAckH9xewd0QXJ
8cM6J+Be27XiKWJGwHO+kz0nPwur0noGLfLeHpsEJWzz+gyHUCocAvaeDNLl3SVO
xAuDP/tMYds1Mge9LAgV5itRAtU7TKfAC7z3t2Bn/qmE7Kjf3seTxFvE1s+Cobnf
URZdx+M0ia6Yt+BXVPc/gjjGejaxTlVGy6DBoo7SLEXqykQnytmm6lEDIRWJEOPs
6UBCBaWZL/SNmSlONoLknREvbF68IUtx/7l5J4WXVvR3LI1FWWwR9FClKNJOI8iu
UBHmoXbsdA2dpjQqbFQChd1moj+Fr4mHdwFF6vEJznNbkvIkaRYcEEtld0H/15jF
aVnTDYgukcS6rFUi0R4N/PHjI0C5kO6RdvPMKLFSHiQ2Y909mTnB4W+Qf69FKBzQ
rtns0GRVmULZdSZZYVo2YnIQf1jQ2gB1TvW5ylzVPjcl69U+1XxvqiLrxb/C/J4m
Ut5f7pxwnp+aiaAsmFhQokKI27Oqj6tztdHVLGMLkH0BKmE8XkYAhfXNLPB42DDh
1X6Hp9DwzNQsUdBdQ/YlQIuMfwsF4oafO43ZEv9BNb/ur/2AIr3yzVQheUzZ+ps1
WlzwOrbiaP4vsnu5cF+vAzTYKGr7GU63YWVOF1qhDO4MoHvJS/UcesnJraeTRQYx
FSGJpPhESL5lw/jkqIJOzCT0Zx6IQjmxfhxEpQg8Hf9laBKJboSCXPTWHmY/wNdu
vFdIcMlb9V12AemTEluDRtQbxCXP9Ja0BjM7antTCYlBwKEzVFKDy7EzPCWju4Jq
05GuhxnQ0YaPSm0WcAjQqCtRotccPrVeCn1LMcmubESOqWRRAF8l+6KV2J5Dxq7e
UBzdZXk/y0LkHBg5/JEATKR7EnbtJUUimKf4KFuCB/CpcgsUAlbsI7ALzYIwBk2P
DKrrxb90dNEDYWqrsMo4FK21Q2Qwje87kNdQkLphNWNhoDOpHgM+VJMvbiXzLkbA
4t/r7EUR+zFrkUVhKF9YzKd2aMCH39j6jwUAe+9flpbsxT58Ug3gZNf5AuADqkwV
QJuLcLBiNoHmAh8FCvzhqpXEZ/lglGjKYMl1g0iRRGFVCetfJ3SKjVi8k9U/qtKW
13XGidpKRv/KxfZDwdRAPtnrF6sZDtVaM0UWy6gkXjbUDWfAYhUUgDo8syAzrcKZ
g6cJdCrQsNPhA1b4iKtJfD5MjnGIJJXPHWxMs57aQT0kBEgwaOIfjbq5fV3ce34T
a5ZsIyfp+ufW0miDKQepO35m+NjhALBJ2hnPJH5TmjRQcRBdJhsDkMBJJXF8sp++
YC/jWMmOzM67UIc6BHi5GjA0koQuEx8x65NeZ8dGqsTzmKH5fSE41n0lSbYLJABR
YHYqjb6vKD2ftQ1JKgWPRRngtGylRzZzEqbsuB6ywNNXc5O+ji5zfgbjN8a4KONL
7qT9LEqQFA54FzQ95BBnyoMH1jj5Kl5u+tA7FV8PeHeyXob4Z5ey8q89cknn67H1
1DCTfe/M5h/kRdKDUT5cKDCEC2ruqHEvhYvDh9TFUDWnOXzxvkPUZsEQ4UeOkEPL
3ym/sH+/q5J9RDGJaQR+LRgth9qA04HraaWoeTJPODOe2twakFYzBLvK1vDsD2Cz
tp/WXtA18167odIQo02Lm4YLZ69lchq7ns/bkqo4fneNAayO56CkAwCQWZtEamBl
sWQsGvWE/Tw1lBVonQyB0qe7IChaSLFd6tE+dGF5Ol+hd934dxxbL9iu8vVGw0zW
bw/ceXfZrvn+9w3Sn4cOhAIQwLtcGAM6Is/4aumptZJyyDAgXfym6gm8zl29nZrQ
Wz5Et4OTxcK1UEgug1csuOxDcgm58O1k9UQVs+E1qG6+6a4s5lhGUX6b7VXb2fmf
51bfukvLU94mIT57q4EYOvG/myvOcH15vdW41y+53ySz53auAdjmsrnAdGSda7ce
/gsWc7NpDIGZHizFUt/p8VTpYN9CzUN890k3+6NY7v2MPwt20scWRvaG3gvVV4sO
pDFqNZlw/O695u/GMuMRssVAP2yDjy4MxMqzMDSkP7VMR8xohmr3fkzKC+MEwMpO
bBOiMjzewj4uSv357aCnre2j/aW0uwdsRVvF81IM8xStS8hAYHwAiFTRj3W0G4/X
qAflLIXH5EfzkvRRtPIaU40Xu/tWCyvj/PQHo6LuNjupK81v94QDyBwOzwRkPXQT
EhtE1BV2kvzoSoKIrprS8nGVJ0Bm/JQlEK35rAQaz7e5SqTl137vLQvfNWWFZxa4
K+VJwyV1G1FTaofF+RG18R1HS5DlWTcx4l82A03F3ebeSEY9M/7QInp9+CQj/IrR
pTu6rDBc0QhCYPNKy+9xJ/Qroka1+q1awtYbPD33JxSYmTL9B8IvGzzSSbD/10UG
uGAjjGrZSQ/OIlJJL9F4bJLSmh0E1Nj5D1XxWCfgj/DE68Vu97FovV0tOQZe1AaK
Jj62MrnAixdMxFKuhIOA+y+ioWpVW1v30qCB0fn6kDaEtE5EHHqUoSAE0OHk3AZR
jDeo6NNYjIm+iMtfheE/gdlbP5eG+e204Nuxj88zQUpxufe/SNY3tcaocGvBPQZa
bTtUl9EWAA+JvxtYcWM2OQwu4lVfE9aWvN3gg4lJ2DlQKZDNc767071ONjGWloZP
semijqfNlO6CKHVfGuaT/JJ03KbMjmesvZ/VKy6Iher6vJeIjkWXlKXEdJLIQORH
CsfqTxVD61ovK7oZhBl0+V4g+L/ATQpnZcxVFbDpBRNKuNvcObfwczd11nLFu3Bp
NUs/6DWArZ1n5ZFSzsNjBScwxKk5txGJyqTHk31sFTrbFHiboeWwzp9OygRlZGpD
yxehekuJBVN57k1rrin7EkPO1v13bcSODnP0l0AAyz5HK6nAVy9a8kO+4GTDVnx4
K74O9cDhpLwTwqgMheIitGlMyybkoAjB9Mc6lWLP9zKhwmpAn8kquCt/CENN2zJn
xIv2ZCNRQunxTdPjvHen6BaUvdWgSNvNiV51Uae+rBpvsVxVnXjlOxrocqqOqfjI
xdpPFnWP0zXwAzhLGPJ7oCmOoafshtdtUDvRpGY86C65SBxlaU56q9QhEI6sISWc
biK+9goiaUt4HrRmE/pzIPIi/l7A4KxYmaeDQYxBL00PIIwjwH5jmUpXl4rUUuKb
es7uuWfm8ylFdXbt+PUNQK+YSZ9lLUDeEgHWbRt8ZmjSUhsGgC5PKZjboy7qAgg8
sUdetgHIdek0vwC1UH7AnV5Utipne9uCeMD6ZhkiNIDmVxxwAYt4bVrTW9cbz/Su
pwNZzxFzxukfaJdQZss96USrQesz1EgMQnLgQ2YRAqDM9T2CDQLmnzuin62CFMsX
Jml9CBVNiLfsOOUuNT34SnZ6cvw9T/NbIf9ysEvqXbENVf1rBidlpsolLh7ojP63
lm0cHal6YKDTu2lt1Ar2aePWvy557ABM8Zsilt6jelJwxGA1YyPOWYwzQoYT/c8X
ZdI69eC62rEb61pNPNfp+uXrgIxWF7X+f6HnjBtpGwLSKLNSncDiBEBapBy4wokC
jnDPSx21wL78yukFeHHTFNIvKIjLMzgrlUkvyQkgoLrG49qPeT4moYCyo8YbgnO4
VfTfWfLAhax1BtnXkvAzZNh9eNPef+XyvydW3LulX8NtVpfmXWiOD8zwfQadyqUm
DSCwTtvrzCd2nmkY27PCfs3SVmUvqNRXBFqpHWR9HWZ5cLB8BSd269GU/At2Lk1W
bOvFcq86OqHIcrmc5uBMdwcUxSMQ4H1QgGjGawcRTA6aahM0i1ibRqOC/id5SYU4
PCa2lqxuyCoTCgSPJOD/nVeCY15xmD8nmkSoeBgpjH74K2CeFiMMfEpGu9qIVQ2I
Mut/+skCh8NGEN5/FV9Rk39g1RT0zfdTxVX0/JKiOaYbh/jn8aJsPMxXve/CevWT
mH9PIaX4iRjGnapI9TUN4y/o1CLbZXupAnCFH4q+jDJMXEfzwNqx4eEqv8OWWJd5
b+0YMQtCWJx5G4aIwg2n513Hk8a9m2DsBptfkLDJl4lyDf9W/XfRcyYnMp65zJ8Z
jr7cjZMauQrDgJZQLeTLmmUiM+d0r0J3B+ou9v81scdE8CJ7tXvmTeWCXc1GudaW
aD7UCKWPBDlP2Ke8iHI58mX/7Pr8Q+p3FdTdbTfM0GWYqWFSruVfdcrK6xRM5Xx8
siknzGDLBsLMqvQcMOLo1zy86lTB15L/EK8lQ1qEWMzOfy/Qr3ICd4f6SWAZa13w
OH1DAddMC9rfOluwff5hZT+6vb7/+bpq1w+epdZ2sjrFJH1ZVmE96n/LpDCND+dG
9O1BTkikdMXxbWK4e7XQnJaRBxObdwAPop9UGCL/GKHoqfDmyjz9B5FnqlOOLNGe
1DHsmRsE2eWabGPk1YM9SodY3onfcasx36bsFFoGx6peGApGE8Zlccg+l0mU+2nK
MRd/SLGLXIXgIZn3CnfhTWpDcfiZj9FN8DOiBY5t7pUDOfRBgksNIgFCDdDfJD92
JZsr7sm75s3dgFPw7CTvrz9+4wX0VH0uY+tiKoxG8O1oaKWse3IWyUK1bSiVq2GZ
JmTplFcvTTlMr/s4n/Vy4m5/YgczxW+5uPTpMuUeEboZ3VUnr6LWY7Zhx7l76gPR
rB80xtZ8M55pdkSjA5X5r/2rZB1vobtIdBfUvHItZZ/gsvhdNFyvZO7t0Z7AG9AU
USHskiMelhJiIxC0FQCjj6gI54I5X8h2Co9IGuO2AIQd9ec6hzy71/qmH2IzoF/i
UwngbsGBlng9VSAgK2jFP2hgLt4FiUf+bPd835QPYnZTYNitDNeEPLQlA1Cor0Pp
lYTcM/UZrppSfeL/nMiZ+bAy3iUzv9D/YujF9nWac1tqjY8WEx7IUsUeyT4DmixT
qZnkjehGP26sBj7xCeVDpfOMYVYHY5OaEDjEJcafc4QZwqHUn4Mpt6UToeT91zEF
ZybDUC2k23TiSclBMCtKSjj6ZhFEXydEDqBumuHTn+iLdDcMU/RjPQPd6jn+bkOJ
H8gvEiGmD6OpU4sY+2kG69MdSZ16XyEyZqTVx5fqCRobXUEaC2XNE8/JJutt2ZCV
Z6wPbENfKajkJ/U5wR18YAORkWYsSWS3mZqQGK9XrAR+Ysb2fkrwjAphCzlg6nHa
sL7Z8fcC9592Vtz5CbzDcF8vdUuDQxKaarBR1O3XZyXLdyhBOpKPx5/+g787FSuN
6kIJ3hkAFdlqmAkthO4BrT8N3LC9JtR3LfuV3Y8BUmvyv+zrZGR2lmSicKPe+HN3
IXIQwaLIf240F9j8Hy8zrKiKIXqXZL40lqQjhAFjEqfGibzHpgjO6Z74Zd0Pm38Q
wi5qrY0FQYR2jrWriOBHsQVUZr/GCp0UX0Kny7YtW5mtP/EL1AUbBlHnsfZh+PUb
dLVwsga8xlWKOjsY5a+1LQe+DXMvTjxgl14Gwh5diK18ahTwI4rUMfCZv+CQIfcY
VGnrWTW9queo/pbiOG6jRvI9w/KJEBJS4SPbGg34vXfru0hnHSef3RjQHhLqonCs
yTyUT2Mrbs31eX5zWLC329/kIWZVdJx87QKUvZ/XLI4pLqXUUhFXybRin2O/K803
ovANvp97hUnuwX8eThPrKCdsnNAtSWwvPz0hgUT6j39+dIV6ev9Wqi5WkH6Tjp1a
Y75AKgQqq3BtxqAUmp87fXqUMTemQ+G4LVn4O8lBXxwgdsqn0cty14jqWswRlP4M
XrSCkQsxoO48ZIe7SUuImbQUnJgb0MEwQN7OBtjAsardOQom9Fl+jgLmOMQF9vUg
2/uXQVe7Scv1LeRa455ebiLBb8FV2QokCaV13oBntUoJ9shOH9w9ZGpae6m98XrY
kxmsM8+E8GuWkZg5odnfM2OvyXOKcOweMzlrdzRMEvKGb6gRqQWRIwYGpRHtbuL3
VD1+uvpN5BCE6PVVmvk1LetURuu6Tfa0bhAKH1k0S88ncvnLVBFLJc3fhW3WdoUX
ncYbTwncAK81d7ah4rT4GOfUKdUM8dRwC5MTjb/vh/ejssJWLZPxfKTP+8VIhXBm
P0QOuM9xg0ePDNFvtk0sLno9YV0hSUNL+GY6B0zSmpPYR1tfZfqvD0+bD1aETXbu
W8kEUk2EUi14gmf6GLoLmMTmE//mQV9Au/eEekoeKORTfpanrJCBO3aGDcQGQJ6Q
rv6TXm2voI3K4GtOp4m9fpzLBwgzDQWeV+2fUCqlzgvgzzQNl9+Q7UlgtGGhnmL3
6RfBp4BB8rtMjRkVIu94NQ8TtSijJanGI89d2a85+dP5zpX9TaaiimHNH9GWzodf
IJ+HtsH+nIxPJlSgzqGCgsfldpq2RCP9pw/6fZLGQvTeHZSJWEzslCrXtfD/j0W1
YtLajzzhmeTGueSKttA7xzAglawoZiQJfoSk3HzggeMv7zQM358oJxe2Yt9W3Hfc
VlowZZaIqg/8Z+tjDs7QJtxOAxbCZLMoB03iN8iCo3JbBndjF6IsUUWCKsuOTyVs
1zzzI7extw8Uw7PqbUdqd4uhZhIhCatPuZHisAzcpXnGeIOtnPTt0Cmw9UtlqhLJ
8Q0ZJnjLBqCM+nCVhI/tfLuthLH6tKXWrq34Ypu550mCpGfEvK4Bfd4WX+c8CSY8
ll8vwVUvXP5Fzuhi6gJm6/q3NvergTSd8fXySEcncsLmZBlNWhaaxTdL13OZFP+P
0lOpNNRLF8ODl+tXXuCC4HlDdsciSL7NyEXcuj2/fmm1yL6N4P0qso1QcucbKaUS
KZ7uvSkxrYHpMb034lS2CbT2nM/Rz1nPCwT9Di8tMFnwROUhDTnegpgxKrmPjeW7
0FhJD/L5T+mmnek2TzjhZvY9fvK6mEAQ91i+j2pDaQ78TN9hFcu4U6sZuqr4cfJf
BltQrsH6xninP+dzJewbEvuDv9fGFbV+wl9te9aPUo+Szbmm40CPezQ1MvcUb6vZ
qVG/SzBTGjEkHukpVXu2cLWrpBs+Sx052084HR5kkhMvJrR0bzAQl3fACgoBZhtm
abn0ITNY5Tu1yCFST48mw2kJgcvyiP8bfdSDyclSp4L2h+zsiXU9UByIlJCoKaz8
T+qmFCudNNO92yNPd9EssKraAWplWMZgnK8cz1Pc9O7fZjNfKySuNPXKm3SMxyZP
AP1D718ihkD1NSVveE4H7QXk3H1dog8io1x8kEjWztC5V3sCkly/qFdn5OrMCCYt
QRiuXMm4jEYzX0GI6pGxTbqSNpHKcJqlmzVoVbhy4XQlOUZalN3v5dNslnN4Jn2n
BN4CrV/L+omGoI2ZpSQQns1IFJ2zPUZJ75IpeMglKGUhXqxt0OnJ8GE4ewZT9p1j
KzAj9MbunVxXUp6UDdTQwumT/EQeD28x0b0G2lZXo+b1kS41+DZD6lCeBELCT0KR
+5P+KdFSaUkUybq3zRqPndxji1/kujYtkVCSrgQzYcoXBAaEFR9VovrXZNZR9/Mo
/Uq3B9+ZIDwik9sQoKNyFgUAQJar3iZMT7nj6Y/GuN5mzO4OGe/4AcESArE6ZhoL
IoFKkZw/5CKxnaw1sBXQaWOIcJH5LlqJbRbw/Sy/d2wbz3u+HJ2nQTJisDPRTxK9
vigCHy93FGQNqwuCkqoGAWIWONrG+YHzTGL3AoyUciHjDOlXEL6OrgMGY/1Qe+Gv
y7j0vUDYhmqf+dNBQ7JfPjJjw8t1u05FO8gk0rUPospZ1pxqIrc1rzX1mxMWXzSX
fWcAhSBiTieSw61HAFH7gmjcY4rAeL+ibDEV8XbwVcj+NiNJN7sZ7aGnNWGyG1yU
H3m+FIIFkTIKXBlC4oFy4pN1ygDUJMBBkNv/cHoKVLgBgPQ53URD8LKg9W7dzlRB
EK/2dtOvmTBNFn+qA7QO3GNXI6arzUz8yJFG2aGOn4YW8VRgT3IafWI2FRpJHsin
DljKGUr04k+G4UgDVY+KNj53fM9MK4cP4llmWvQC5JX/Yx6nAdu5+Xd9hYTqOR5C
HjNGuxPrdYiVZbYzDJWNMXs63RGbskvjrOyGMh2f3UGvZtpOhynHudySTMa7cX6H
Ay7Uq5t6E8B+lSGIyyJsN7f63n9mEv5nKBREbxjGwtQtyMsluHoOCE73X9Tll339
uMdqqQuLz9GH+lwHPFoF3C4tZ+eVX/rqXUMdtHLZUbl4ZpwFAhnZdWiGU4nEkDs1
qI4A/LUna3xxmlBMow2b2MK6neDXDDMAZLMfDQlajjgOAKvhn8UkYllJWtyQeTXA
iFcvZ2n5WdirG8PqhKLueiH6MTGj/EszhdKSxRSmxwTsdj4XS71v5s2dS4nAAK4E
/XCFrhBffzeUXa4IdlqMArOR9yqwKEh6nw9uuJ8xsTUFt7KiYQifz2RlMJXL2vk8
6evDd0oIfnuk0WqWgc7b0CZ2UzkVJB++Ok+ywWh88sec3/CGzkfvd1kgW/bdFGVg
fryvuF46iwlgW26ZjX1zv/Sn2Az6x8LkGM7gkO+lrTKjDkysMMnaj4NvfOOyWPU/
MH3Qq+Pka4o0cfIhh/FQrZYPlXMfMmymHPz9/P4D7bGIG8G9a61PdEzrALg3NTvL
nWvK6KCO9fU6T1YpAFog0aElkNXEu4O9fBe04Drtw82U6UrjvJiHRJPU/cjeWWKM
9qgHWr3nJpXasBYKj894JAb94Y3/Cgpxp4ezwViI0vkdNR3BJdqf9PHXhIds51nh
qbwnyuX2yCgdVJECFwPkLAUp6zcndbrqSnUvIHQBPPI/mlRAu+IYyqnSA6jVfm3l
b3TnF4Q71nWaj6Cqh4s/8UCaO1IAyJ41Pjd2DhE6vdLclOlwA/SMPtIf4nc1QOka
JF2JKTMx6kgwmMlECyJao//97taommSg5ds/ZQZq3YEng74pdxYZhjM8gFcWF8ZI
nbboTHZYYxoHA1THpgOgNgChWM4GK0ysROmrA1sprkDGmyGR/SXfXLlVDRAQPZ4j
hqoyDtz5jYC0XFNuRTA2UzXERBj51Pqzdh8mKOP9S8dPkvZ0wM2DMeqRg4lKmzA2
7Q9sb83+OUKJ4nhG3qNSny0B3xMS3naB7jFJMwYytfMfASO1pVXXlsxckA5kQb5j
ACMBP/BuWcsySG7nHEKQtNKqVdEH32Gv6trZx7X5r8iL0DVCXbvs15zZ5mebEVQK
YbpnYKXiBRHs6RCzgUsU++cneIRZifWG2xPl+Sc9ZNOOU+SEj3QQyLuHOmNQH8QX
Uj8F/I/dNi56izKLIGYLSUlEBFXtHFkWjPxew1Dkat0RhaoZ4+mKj+hV9CnDf/7f
4wjyOU2Lb0jgQkonQoyWsto0ZmlDsZy8/kM1XLMiTvCPHLp+GF2b/NvT/pouF11P
BcWVEYBxieQhDtie2lsLb7KMKI30mYE+zdiPQ5FwujezvWnUKJ7Sq3XxSk3MVlnV
dS1QtBBPaNhrJUfFQmI9T5G/+mBJPxgAGwVXk2FoiBkv7nZhDC9YnASZ6gbkXqB9
p3v0VWZvt1cv9m6MbnuV6GrC0ZhH4Qt2iD23sOvh3yaU1qTnKIRUsuqZSXwU9LbH
zn0C8GOTHow7R1v7Ak7V2aHnXmbCxekOzjNX2BsDrVgz6V3d0D6I7K6deov0egOU
VTAm36BiKkQRbC0KXW//ZuIvZvhWtszoOA1C6yzQh5Rl3dge/Z+L+Yj27O5SUPgv
0PhlJa772CA91hUsuARweYDYxMhDO0Djy5g5ktevCkoz0YpoCkbwoLZs0zM7Bn0e
DZJk3BqBQj4wCsRB+p7A8zo4Ue4dSlDeLHPbArQZIGZWX4FCfk9FZ9VidwrrAUEo
HMumCE6aGrXxvvFEXn2lZgmC6EOL4AmsGgz7Ft2ja/LF9mdox8+xv61V4wwJD4Qx
k7XJV0aT87TSzbqlH8rIvsALk6vDgyU6lWlkNmK6moKvkiwWUYSr8QGCdqh95RTE
3QW2vFC1XB/dq8+xZJh+Z4wfC7jLNjcUWpLoypUAc7wcK+UJk8twA5dWJtFN+FVJ
flCDQJcERSQgww/balFvgFfTw4Ukf0c7KB75Tw+YgtZob72KRGsXTs6jE5vn3o7X
Ge6A0CC1fKwxGxmAMSaLtFiyyOi6Cm1cdAJJhDfbuscQUIjUfGcSh17MbIQyRLFj
S+oSte9HX2C+zZ9zXmGxT2oXnBP/TbAolpQKS50PWRcZV90uhu/3Kbs7cPEqjWb6
b+DI/00yGS6pP9U+oat9tjhy0YPkXD0qIQkMLokrQW1v3n6mPzZzsHMLy5adoMuy
HtyVLqLP4gjlVaZ21Y+R35NyH8n6ziYFRg9fv80mqt39uqrhXXCsG4QW+vFnM75g
JfqvXezanMIWQq+fdvNVCKvB/BY8eSSRyKStwqc+l1jFwyobS7UCDD+UvSA9lyid
Y42PsEdKSezJHJsovkcEZ7qABgp4Wlb6HT7ygrNvoCKLqYLOs7uwpVLI/nBVKv0c
2u9KyA3PgLYBsKuJpap+fsBmFlcxfWIWzc9zgfWAsWvgu1EVvFizxyKmwkX+l1LC
/WkszA+Ln2tNA24NYGQiJL2wJEDtVmVe/WE1wDvkPjecQPTgjE9AKnAo998KfyoU
7z+cdDUL6hTrqxITbedAbZZECKD0eDcYiGosDaFXlf3Y9ET6OwLlKMSZbsUsxgXO
gEZDet3ppaiKEFZLglKCAO9HxjzOvwHR3icJlE8nxRwUWhrgWtK113y7HYaWl/RV
1umNUSAt11ewVN5r1cmC1sL3DewwB9tIV4ftJ2YcN/1QAiVpFh5T5Vvr9fQ8vsBu
avXMvW7HJL6Mxla8QQF/Da7HVRfOOfyxjEa0SQ6DAEcbQ2DP5UqQmdiXsk1GIwvR
mMpMPB1996DXbwEUu5hx772RPtzDnFqNmjtPWYDOl2HicRQAOPRtMaUroppFj6Ci
kNi/OM8q0Jj3O/BVfDnYW1ZDQftWNBC4rnvGRaGrw3yatm0166QMIMsvIbnvBB0n
69ZOmD+lCgEVq3vND9RDVVTjdOwbb/r834tJf1VIXFZHRcaJgzJHEfx+P0bsEMwN
cL4th8LcMOcVrNpNNKA8i4Qw3emgsN6za/PaaMDG0ufGd9jv4BUwTkA+YywxdeSL
XGmsFnp5SDsZrx20o5+tnLna77RdujvXjBL251WJJIWor51Ac3fkz5FHP2Qit8Aw
KqCT2QRprSjqoET0akmG/4DjSzdAU9e/UnI6g7BkIL26GEEZ2q97PFEBFSKd8K40
krSBvf9aln0J6NI/nTI9227BbPphbjGfWOh+snC6pf98UDTczE3yppeJi3GyJaOv
6aBzKP0k5dR6s6rdaQdiJUCaVCLsSRnIwMAwdJ1vO+eNdcGWqwXBb4GVCPGJCN1t
BMGogHWMbmrRXX18iqxqfUv9BWBQ6+JbeVNPL4EZnjCG+dp5+Ra3ZnX0ggnQrATl
5O3Iz1vrzyasoB9W5dOuMJK91wNbeD133PHkfvcAt9d83H2n8HHUcqf1kHbZsegZ
oD2mfCxuMk643ZdnfQDIZkcOy6l4o29Ivta8v6PQMP6FSCjxhEQUEo91C0oPhOvC
YHzNi4wTEPr2CAnFjnvT4n0ZS8X8Zb2wTLnJccstWxFfDGO9EZ5tVFfpW0MFrF95
sIyHMRhCkwliSosGEIBY2WEIWOtQq+B2bFXL7biieuNcQ+Wfxga+TinuJrvFB8Ks
aeNFFt8eci8NBIIW1HarPcPa8g0zHoL9DXYUyc6rI0w1LkcAFF49h+iP1d20IHYA
13J9azx/RWf4BlErGstmuwKiRBleWRECCaZWz3LKVwhGxquRoIHe7ZnvEPH9k+0s
tCIYAmAG4bb8XJ4NfSZImoQznE0eMIFhGlCR6TzMF8MvKJ37TegZ5AWLlK87Ma7l
O3/mKOMdP2IxgglllTXg3cRXJq1eJXvFJpJOFvvlCixPOusUfHQmLfoQtiF1wI9W
lofljjNcwucl0z5rJlaLhYprnSNBkhQHfTR7fMLmLhEcYQVf6hoECLw3tn22b9b3
GjQ6Q8MiKDzQ4+nwt4qakyJzJYJBzTCy5Akg3ungjT4MZxt7Kr0K59KcLR+Yv2/o
BQOwuiWUVkYUuJ/rmqyFdzkfzbNTv9h1G3SDm71XG2k8tE+sk8PAAM5Rkx6tiGLX
q3l8yBsdCrMDui2Sp/eabZ0bmmylALxZWPkSeFG2hfkS4STrTkqJMcpPKYOrFr0G
3xEOZIfWCwLD1mHR2KAN4wBiKwhnEZ+h7KnF18QQpM98FP2w+GVEHX+XIRi5gH1b
Hp8gk+kbmrsYWbyIZw+GSRVrlvQB75sbTwQo2taeTOTn2YJr6sVVE8nEkNWPrOhR
HQH0b+oprGlVNc/FUuIxDYIAMJi4AClM2p9PWTtrtdUp1VwOvD4JJyRRsJwe+xfJ
mUaS7wWQNQpza0ph5P9137SaoLTAldFTB/koowy8Bh4WDrmeXLyW2H9Sg3upXkjM
dHuokg4OlF5NfBZJ2bpOXwI0+cQXCpDnWqHOg4xsdGXW26jeWJYmtoXFyI5dJODK
MbE6vaPH/ACViMe3B/olmiwF0Sz/fo4Og+yp34bvT1H2FAdLOWWIRkUwDGviYetF
MdYc7Isn6uOUzgbGHuKB2UnLYZUPmlGq8GgwfWmPhTuWLF+Q0lsfhlxmBj64VcJy
vJ0oGI68Bj80WNYQbq0+8gwBFoM21G0ewPPAnLR2TUQZ7DVsnS5aG/NuO/B9B9rM
bbQ+BUyxo07x3Hi+zdT4pjECYqDFYkWPalXnCA6e5GxVBnfSWZfp5ds9ld8k36eK
ap3DY15ZK/fWrAQfIkf068FMF99sWfGClBvze72cSZxQ1WIwF31kEm0gH+s6sJ30
9sg9wQUa0xMWwoc9f1Ze3NwgyGmkTREsXrBjD4tPHIdCDZLbla5IhHsrEG6MJ88J
EecmaGyl3LpXiT1XZYa1CwK1LNp9YzODN0ekN0LbHbjEPrUUY6+xnCvsz/JFvNTe
9KcJrcY2jmXzBfXbJzHJ9uY4ablCwYWDjdiQOGJSBAFvY5Uk2fb39KkFwuD+3Lpy
gKqwgOH1q8wFJI14+pdmrIKyyN/hq6IMzXL/b7crESBQPDPrL1fmm18MzfPI3zo1
B4tHkSFvKuLH/8m70qplPI8bshpthwO06bTruWcAGJo/bMOyUGJPW4wvxUg/G1B+
Tn0J98byJSSThSnIanXfW9Za9dkJYyYbB3griFhRDZ4PwCb8VMBGYeuIHx8bJREg
H5x+KeaH5bEMcQYqHKqFPNMjO/XmflZkzCyoyMB258H+2vC39GYVH6XeXJ/XsOmP
n8JTFttrX6hqEGXWavJJwmzMeiTj/Iwy9TVhCPId6uh31p5cTOABd4sFmgCAaodg
FogtLS8bD7SnOHIy+a8KZ0ZP5L7ABBW/07kNJgE/2xm2mL7Ly4jhcxZyrLDnjHsR
fdbLSNezyo1ccdNsySHLzM/PKo5ugOO/1h8e+AHu0LiUqGiLlPqbVhDsf3KVkoff
HcA3dQ3n+Ru1J/V3PE8r6PnN4VspD0jYq0r1/R+C088oQGQqTXH2qrmP2hy633gs
bWfKplzPB6TC+BntYqdCNVbD8+qadnZq8DxwOt5H8sD8dF28U22H8E9iq8athPfB
giBE9Hrdqbes6dhXRIZgb11GaXlaQf7c50cRx16/QCBxv+Lx5Iv5oQRFCFN8EgjS
1mee2hRO0cxOYwHmzN2NpQRjV0hXOetZyvzfjmlzkkxRp6IPefCH6Tqed4Psolyo
E5VEJJyIXDqWuUpuBnkKAUR36o4reCLj1r5wGLHYhvYB2xZzQm5IZr+2mucECCLA
tC0gnwlR7X2Q1fwMlK1S1A/9kZTfiChQVZWCQ1RdXBHmz5AthsDC7X6ouwwuFJfA
MBX5xSjmS3DlMjnMkU/68dzLtLr0aEvBS7AlViQBgSpPcNWzYZsCluMuAMZwyw0L
xaYJpcoaBytEAEuG9N52MaeE9CRiwKqmXBU1Oi6sBthdqR6rKbEffyMs2lO+sDLd
U/d8pWkv2hycVsEPR63m0EV5lpfPCJt6o9OjKxWeo46EEanXN6dNIGiyuhsy+s/h
1hOULCPu3R5Cw8CvwFwkvbkCEdqvugzPQy3KHsC61gXNV0QHPEJ2MF35SR1BpeX+
kqnwwYswLfcQsGvmv49s0DpoSLFFm8JswVmzIOTZuI6e+2Si82QLBo3kTlFEGKRW
pS6VB5Rk5V1hpVndaocqQU6xZHuYqVqTXUuV9VXxt4mv5M+5MZXsCvAFjPngE/wG
snoIoodBXMupTOeElSw2pThdchfxlD8KiDsi7evSh33HrEETzncE2/vrk+VztRHO
YN03gn1UgKl5axmYIF9SSd9LKXYrrMBle+WHdI5e1Zy5pHYVO6Ka2BkXCvEkiZYD
5c1qUv3iTINkYGqO1q6g/caRQQddrgmWG8xk/xS7459a50xAdSCP9LHQ8zy6bJTQ
Qho+WusbL8uy8pfoZ+JYzJ/NfaUuPKIG5iay2z9xxgR8r2zKwbQabtNmYlq6oTpC
2Zt/eKYV/D0QB4xfgqpYGIDRW4t8Yj7r4IpYBLAgVtoFBZe6Tfk+EeEBqSTKK5lw
temzIw2oX4FUA3JljazuTLXnRHHhE+Gf7pIKZYieVD7QJhtwDtSyEzayag5Iky6z
xHA0HsDyvhjKhNxWL1ofULXus8Noz3/CKkyafrM8fe/pASPxJDQZ5GFZAyF/S+u5
ix1RtXDas0u+X819Fip3cr4VUsilyzyOcqFt1mwwMk26AYI1JK1gqxcyhbmGXlF+
wduD8H3hpobs47ji5byuYFlg3Og5KFcGEE9WocEob7RPFgmkEakvzk1kS5S96JQ+
9f+6qDO2OkizgQ8R6v0/sUjKTZOqbeAdIy4RjkjmQerYSmAiItfN/q30WxGl51vH
Ey+sC+4LYyAs/RwoZBhgeiy1LQ5qPmorkw2P2XsyKGNAGYzQCJyZS5Q0LV9n3fLL
nP7P5ntn/lJ8LRyNfE9K4F/cUG/7dwMmJeUv/+rNBi6A+Y1JphZeutwLEnTDgoT0
62Ew9WgmV2s4F2ieibgItgbZcUsYjcXlVxQMBoKenl5IYOk2Jl3idb4eGH2rRSag
ixeo4ys9GJLit0AUQfN9iSRzvMe8D7JJi/LOxldHRxO2qfVl7vgXWzalRyqAS+OJ
1dTcnfaSvuVguR3owIQ+Jmz1vmYKettj3zZGReikMVNUg80oF5KiZ27hZtODSbWl
vIhFEF0knJvXTSimeuU3hBmZrufZvpeVPOlpoiGXbvdlMYzH80WBgnESfs1QWFWU
rVFdR+vyB8IoU1CH43X8BGgBfNWgcFsYIF+P22L2TGH93+TrBqXAz5uI78gqRjkY
y2FVo1l7IyIztes8r3XLYvFWuzPbsAAmaNAfXj0c2U3rD3k6F4Xy20IWGdsIhHKG
+qyDK/TQ8+106QTazg8iqRfBWSD/WJ2sKQeZ6bjxMUxI78VYK1dfk00Jt4BZj6jl
cbEsQa5/U53v7ahs3wZd4jPYwIbArGL8c+6iiz84LV4KG0lvvn0uu1SPoHd9cSdU
6MepcXWNFlvzchI8p3tZoMA5I2ncKcMrrn2AFrh76QR+QwwtsRmwrrOScqkL7Ynf
NS3vQyNhnGjXX+CQNid06xtOa7apa4ga2tiXLGJOu4Ca+GP2agCsSBeUiuYMGWPy
cVaNpLGplWfYc23ewkNZbmITvO8wxoydrd1xEwrA3va1ph/iLk6bdsyQT3ygOmx2
oxW1kuIOdB4L6a2sCy1qJphjNjPA8/fPoUSoBcTkF0oHnUsKCfxxggmfN46vlk1e
bqq27NDPNH0n3rZGHi4YWui3h1cGpul+3CMwsqK+egbTf+0xbRMromaSYDzTDI3X
h/t+qrALIBUddo5qHSwX0dOIwJ6lGvRWnjH5iWcBHOdVDoxLA/MMHsMQQKVFMm0U
Ssa3pOrKqvuDkOSl8RjryBnV3fRzyMPfMRatA932LTD262J4OMfhl2YJFabDXJ29
Y5dEl3l13U9w0aPA/+6u+zTPAIdjTMPi+AASgpePyv7huvYetgUUNF/EiLcMiDP7
W3TOso5xcAX+Bc4lVSsN2iyWBE5pYGZ/bdM/k6JXGMgZqMMaBUfMJNfh0tMoCqbB
fWAB0eAdWp0CVN/FVQsKn3lQzxj/Kc5anHL8rW/MedTmvlvt2kQPG0YQ8n8qtZvj
m6GUTeFiPzMvAJItJPQ8V4vTk/P6Ujuip5kgeIfzjNNJpQhH9yooIPEEYVkThpS4
hcB4fAiPRgbuComxl3ZPhShGFAkbtkq1nKn+7nJVm/WYMiqrzgN/3FaSPVnOLvqC
/ROLNzhIukgxN5UkdpP6KJm1Fu1PeRdNvyoWn0WCOMNgOTLXyF38gMKH/2cJukxL
2UoLKmjvNyAWBEVRU8cmCv+Azxm2Diwwdf6rjSmwYlytwc5tLmNp95/k9oXaV6m8
9urJzZ+nch/kt7Eh7DRBElitS/28UPfYo0MScHaRFLvKAv/VmeXpvIPo/h3ZaWgI
Phbmv5wqowDcOmm+RjaRGuABp8Pv/P1POG12Ky6N/YxIhDR3nKsMjtt0RdjQbtP3
AZ5MRF7MKSi4QDiyU/PMO4dgSZtYeV9c7RRuI9+Bz4+IQ1YYpuwQ+GBqHqsiG50H
nMbt/MaRcAldbn32dYNlpNZY4DkfXdZEYYYu0W0puYPOdK/ayuTYjlEgxvSxwLgb
FdXukjtJEiPqYN4GamHYNtCImZdkw+e7/n2mBUl8KlzM8tPesl87UL/2WtvaC9gq
0r/IIwpwZjnR+f3Nfp983hKkCSUGMLn9uKKRK5ES8VQUe5BEc0e2o3ZqcZZ8VH+U
0PRtOPFE8WdKvv5J76Jmzzs6nDWJ1wFNyDCMl9vz0jLNP5sqS0ECN9vy31RgaoMw
7sQFNEK6XKyKDAKhypP9BxoFkDyvUBbjTd1wcOjd+s+H2mJhqjCslxjtQEn8oGfH
daz8VKn678pj7/KrfCE30VWR3W4sX7XfmddhKuGoZd2WBvn9CK0jazsp4v+bzmfk
CpsahkA9srqyGvxn6H5awk+jGHKHbPDe0zOGVawOifkZjXFMxCeewMzbvTpm5qTl
uP9iAvVNfdqEbtP6Xxe2uidnsOC9cZKXS4si/dyITEtblL3x35bBbh4YcqwR2xg4
THkOrvorunDgeJqvQTI5TkmQBFVTrF4soqD/NVGbJj4imPCW1lsIJBZl75bg2quP
cpgG3ccv+xXVSaaqaEMEubnAE2Ap93IfPLE3nKyyUo+Z1HWr+HxrW4o8hvvemj6l
AY6sywiCVYacsYcu202Sb6vh5R0s2BJblxzqYHwu+U3AyequHE8IyI5cpwVjyKVA
fL8a9P6DjkZHYb/S8ZqwUo5SjyqdoThuQZTuVgdlIIOi5JFSESrmIHilYycFL2cb
fSEOPQWlGZHK7URwIO0yJ1jHPBCKfVBUzKNKsBEAb8IK5BUvQdsdtFixKsBSa8BF
TRW9qUHFQmw5rKRa6m8rjBQWzyfdXUAK84tTSPoXLzwDLoOydLCYbnWKMRu5QsAQ
eTYUjFUqNIDpIWbrfpSvR98+AMHK/+EPHtbQbkgaLCBQsresIQgv7RAtYZnTxgVO
dIiuY0EoUxy6pKc0jOPJYoy9sjlzqZbpUGYP7RWV0GHK9NYf4/lN8/z8atYShSwU
2p+wASXseeW+RSVN71+RwKolr65FZnku9w/R4YrWHx4VU6aZ0e/3jx8d+FwYRqO9
xUjwWx3VOZf8xBMc5GlzRk9QPP4fAS9GtqUwKaLdAPjHaBT9QRXiZzRqFInadoQv
oMHCMzH4yHWkIlS8YdzCUnL6tzpoUPoYlI/DgPOXiydZuzIRvHeVsj8QQK7I3rti
97EVGJtV0yXxsYvU14vliCafakowXziiIMjNU4J9e5D4cUJI3E+5fYgWP/CFBLtZ
fD/Baz6D+yqq+JBj+jHvQlhhJJabVYNSuzpBpRzu+1lRMtzuu1v1DhI67ABZSp/t
TT8qLFqkCw26Ur8V1S+vZqHM24CqXVvsp/II8/jDvtNmMzSCtDTOEV/SIRgSedHk
Xe4/WIITe8F3BBPexJpud+AdTVN1jnU4LGYL5ppq/AY0M1UTA/0lLCZz2wsVt+HS
39SI0BVjihnQikZlptolu3Xs775EtyDdHM2wMWfau66WCEZWYpuQGJ6TKHJ5hetL
1MGrsNCISw8+KV7Co5B+o6LvJgxalPArbzqh8hbdv3Za/GAC4uyaZXiGPtOVAdGK
8qjGM78Iw8HFbmm350e4d2j5cE8JrFOPujPTFerTnx9vyANyEDyhH7lYSriFo4FN
c1wu1ftCZjPGMzmwalDZ8L/q+q5tOiBvS49SYwMYj5srwQAaAn4Fk7c6AuXbgkNt
UP1bxkHS2KE9GgjguQ6W5dpVSW7S/QuQw0M/cTkNzVixUZpg3Q+vFmcmuVP1+gJ9
z8tZHU3Zx/DiQX92sRT0xXB64QFmbQeka9cqLnOPLwT5/QwTTtaRKMyqZ0l96HvA
ap54/yYeni7QkDR/OvBTUgHq9eIEEZvb4RGEXOdnqcaNl7AgBT+rF/HrqVueUPoX
wGG5QTVpKFf/0W+WjfJKDbgI2cVSwvubgJwE5z/rsrGvMJt2JyIPUSWJc/1Wtt9S
VgWJoxB0af0/JiVUHcrf6dxNYmKntSNkdMaRjsztRVklurT09xvB15oWh8feeITh
Sm2GAzecFGwtaU9FU2X6jSKtYpNiHY+Ratwjmxwx0BXiANMRlnqM6344TFzb1yD0
HUR85RLvOjulF7EIY8+0i6DPVBpzxzmQl3CH5ERMXgOUUwuu8ee/Fwf7VWlTH81e
QjVVdb7xKvOp4cFXT8xVKRc1JtgxzKB4KfehovEZXommmRvMpIbaMGoNoMYKsu3C
9Z/xiNqSJxpJkx5FrY+gTY2ErW3kTrwNIjo5FPFf/2wv7LouYQIPdIo9gcg5T9r4
+dpxCbJHEiLq+5W3+ItDk3cR4ZDQM1uZv9ha/WA75wX6cRt8GOwaKP+5dUpNaaRv
xObQDgZ8SanA2PLgtQA8grpk1T+wbZh5MNCGrd3cOG1JkCl5lvTlVMzv86/Azbf8
BSPdt2Rxclyi4oiK+spJgrfVPi80qI4AGQqBgT7O2f/hxm0XyJMJ4Qp8Pu+FHQTe
QUd2HyrVmZBvChxDJ7bay1RpVsAoKV4LzKBYCCOxZi8WresVt38EQcyxrgERPzji
huBxO4fkcEzOkCfZEiVCeX9ggzyzYTgRImJhZ3DdTaIwOb8JTl/K6gknXK0NHfR6
v4AYkkpcqtp+ClksNNeVeUw+n5eC+Pbzkh9McntE/s00oD2afQ5g7yiMaRxMLser
KsWkqo0z0Isvm1bA/iAtKixPc87tbKdC+a3FxewS3ic7r4XNBHyFzaQmjVQk7GpC
+6wLxVGmoXpzzrSrm7183UtNY6cRSJ/iM8LkIzekGpmW99R96dTm/C0E+IvC6KCu
AtHYuXNNNRNUAaudRhyLkeABt8JrPCit7QKvuzepOIF1gE3XYd+WaETpRnzY22dq
nM6ZZ1K/72mAZJ0xzlEggNLx9g3oErg+QJ7a5PWAJNrnkwM+4PgiYK/QMCiUgaim
Gd3LKwy1J8PwgN+55Coj06TOStyrlCo/LtdWNkG0dOBcqsK2e4oPNFmVsEhgxNd/
TEAcvLqkxhgG1ujzjk8SLgXOtCEgRPsJ3kS5J72yhUVeVo0kBcilkjr8T0FRjx2I
r1fBXhxQpfx8oLM3Gv76NJ7+ES5o4mqQVhlbREqxTAasyaIyyvVQXun8JDL47ogX
cj/k9tLEtRecgblJVlMjoJxfnnkXVmxckUiw8/ee0bQHKxzF/TtFSzxlwBDRXUYA
FieFLbN3Q990uGPof5d02eqYOjLImIVc5cxT+w8YKOUvqHk5djfMMfuS09pmulqE
8mN1LplU3tgqgf0Hz/OFpm9R1/0Hv31lC5A5Al11JZ5DU2/yoIZHZlqUyyxonfhc
1bcY27pe6s+MxQEeh69Uvo5nVwNrm4hu9zbejwBBSZEkVRlNTsZeiHeXYN0t+tvJ
NxfEu+dca+Twg21oqLuO1zfKbv5VW5bM4DA1GegaxxuCHDYdvUdrPTlIdHBp2gqK
7SrQHZgwHr6heOprXn3Cib0n36IZFcQ0fjqX1CW/UQzM42fhaiEFSjBgVertoUC1
nARJsRMHt3V9WKXF8fMl1d+TDCS4/fTBmz0E068cAOMc0xKb28gk+bzm8CjwwMlQ
keipmPFFx2PykwhoMy1By04Ns5tMDHySu60Pm+7YQK99Lb1HsIzzFTvdGgAJq0xr
d63FCIxNliIq6H0IA4YwVUEwRdGWlxliP+1SVifKxS5WvzRPr4kvLFeA99rvLB0f
GqbLsL2zddCoGM3notO+hB34OaQ3UjJ2y1762rRpZwY6MFqGQDEcq5Qmze6AUSxj
otkiSRGhR4CdSYHZ/9O3xgTUsOelUtagKm12pKIgO5/SXz/t8l4YsSSNnEtZaaaq
W7M8NsZl+sAbhJUfmLvUFpPvWBSL+QPCLTmbQSPEB27o5Kr1vSupN5+xl2CamEAJ
3ZkkR5B6bVS9Wh5LfP/fMo+HR2RegxyJLO0tZDjbHGCVyNaCvUiWhC7L0jpZO+k0
dUv+NoZqusNhyGugkLDYcy5BKddATZ97RGFeW88+s8RV5XYgpcKfclYMmvlLf0BQ
o8HSOZNAvsNatIc7sBRh1NuXyb/LiSvnUpnwZnZiVfJoL0tqyIw+3Lh0jNLBT6Ck
muZE57KCa83s13fCIV498oF1sMOLgVvfk4jTzGGxy9nivjLccBkVn/dLCnHueeQd
k7h71WMrkylbIbgh4nrXq3q2MSg168Z4/L77LK9yOAg5eUx8AhUlSMLNxmmgjioG
Ut8bcxbdaJWF+pE03Fl73/+wI2ELWRJYPLlFhcjGx6Tt8l1GvqX7Cb5bWw7nkAKu
thrbo/iToI6IHbaYb9z6J7suS880qNel0v9wlhD1bkv8UFXjGH5CcXpEHHIhHDsQ
syGrxFqV1kslLdGF5FHMzHsVg5aWPDwGROHMBjMvVet5YGb6wP9mS9k4N+8G+Vf+
+qZN2W1KIHPMJpGUY7fDpxIo0NHXGMlq14w3AxO6/V1rC9opU1WrdtcivgsUWdCE
cZj+qEMoJcI/CpmjzpMVlwcG6fx43y3VJwC1UzHpT+Z5iTwsxXXGe0LZ/bl9mlZy
jpuM/lBWfSEcEP1rus7mQzFR62Oy8ujDJIIIwsULhjP8A0wJ4FxtcH9cBTHg3uQj
mA1/2yvVxQ9GF/uheTtj98tIon3gF4+GgWbRrIQHAqZzm1vrc5p4v2YETGq2wLxe
pz1fXjNmLRs2rq7UiVEy4f556nYuUCEaWKPYZuvTpGizeu3lR8AcRCmERzC180Ur
JPIOmll5WuWM0/KPuf1yFzcwYmN5KCKaWIfWEipbpBGU5Tp9TNVBqKEJqZ5t0Aa2
OQZz1hQZ4iWBeRlc2WHv8VCS3gmxjqWdFqFvoAtjbBMklek4WwEg4UIJ5pniZfD2
sbmKfZh2TPwzmmlBuqEvLtZIUa9dyw1Z0FJu4tWsTosqfmsTshAGXITNISaH3GPZ
PdsDNSSgbe6BPaM1aQ2zCsYfRWBagfSeW4BrKS8t0BWjyfjcTgNfIK/KsNQS9x8r
yHoRQshp2mssmDXjSQ1Z0pCaAPqgZTgwdAbYeGkOS8serlLdz4VpHRyeOpGjSTsj
76kixhTxM+GGUYAlw2vJHKwiMzL6H+d2E7HHQiRxUR7iivhnPGdTawV7toV99CTj
loshWGm4lqObeacxumbXYiUkO8ho9Hdq60BuXy0+HCRGRuhhxg4YDT5DdFu8c5sj
4WZVoSpM1cRSvtKrgcvC90JcT4vVI3pBrQhKRn8Xg6GHzyDpqiKuvqVfknpDVHoL
7yZVE6pv67BTDR1Ybb4QdjV3oLKGVzk6JSICkPyr3jqSt8VpQ4Tliz10eOj9t2ex
uMKdNCL+PcHeN78z07EcVPf7ibyAItAo+Vf+GzsrwLNl270efiIDjEIlp92+Aev6
ZiBQGj+10KNBupwfJnqZIvQA/UUe9YBxigm0JiTw6fBR2P+rte1yoXBqWrrWvkem
rmzjPjCYk+wr0A0cd5JvDgGbmIMUJzzZ9T8gKDmFVxd873b/9qjg4q6FqUVHxk9L
DpqcrviMQn9kve9wlM49pF2oro2DZ/kaCWVjHjtPfSrHs7L7MdYQpyK35YMm3BaR
9IqnCQjLv6wtoU7l9/i9wO1iWrxvxfiNZw7ZVSz6UlYBlD8ToujN7XYDAJnhQEWe
NASO4nL+YWgjH4FBkXJFSLYVcsI43iS2pnP4jKu2M9EQ3801/T+YMoDdWHbRezAA
B8iI5cSS1940cPYKLWFGYyJxceROLNNWk8XviS2zjGFG9ZcqQEa21Wdil1nIzvHE
C085+I8J9dSjjipWE3T8I/FWQQ+vsN/zN/TlgwOaiB0pKNDkt6gEuORJ5vUmHhgU
9VSs5h7gLAyxBT74YONLZiQGkrW/tkRzb0iQ7djSLS4c9Zl3xVvMSnIDS1P4qp0m
1QYjgu5bztLZIMiKCj8tkyGmD7fIb2cERudPnjbKxlQhkesSqNTXfFY78PPsgRok
3fD4PaHSM9Gf7AAi+qvlOOVUIIp3furOs6DLTR7mBtHDy/tw4fJjI4OGZ+mhH2se
vjVQHFk0Ldi+biFR43IMRhNwtNIleILZ+E4VE/LDDw7gDl4PxybennyUwf9Q2a2S
18vr3ELBOh413iG2RHj4s3OePlOEjqvk4OiwL/7o5YxWgOh7wY/Njcf4CL4GI+28
DaYZbZ/6CFHmP8sqacpk3NPJdcIexWsLOZfC6VaFS2golxrxeTJ+aNyo8v4xiv4/
TBEJTICC4c3C5CpiQ0SAz1/3wowMFS8HgJIciekoemQvZT5EV3XG6TV4PhQWvziQ
aWr7XHKiUokTvdZxFr+bNqNeCXWkUZo2oF8962H35BKZnN5Upw5YsaEVpVPuLGZy
2hlCe56ApyUv6lS/MAO8ERk+JQTHnMKZGJMuCdeEVMMxvgQZq4ZvJxC2EmhcIGRQ
e8/ire1EyCnTeNj1RSuplctPQxbKc5wOulunMDmIodf22qr/iTkW3dxZYMfItRKo
OgFjbPWofOxukhu/5pdKyOtD5fwfnxeRxxfgczPwKCq2ibVazLYL0ayxqwYkwrwJ
OFFfgUBxUf5fxm/1AZrk13W+bmwNa6+u34SeCL/y9qcutSYs/bqt5TleCb0fc3tO
gNoTiIf6HB1Qb7U6/1U3EwcFgnHhSKRUqOS6vLDO+REJaTmOKq2NLON5LfnpXaqf
quvYOAlYZi/ExTzj0KBchaWMGQZ/bzKxAspeBj2YLCDvOHP2Wm0+JFCWDkHm3wjs
NrnwJ6eRJstXs9wQ0IBdwtkGGjv331OkNHW1XdED8Dp1qfksPsB5/22sXAXQ8F8m
5GenFs1ZjbFWgfYujxsvzqHLXM8xnKu1r1HSXcqFDYJG0CyFbJQ6C0ZypEf89Fbd
Um47AMIBxpfKwSQ0i5q//5PSgopH445oeAvtppFpGHqNCB9w4kK6bXrdiMeH+33U
HsZ36rPVTSQhFZEkjYfL8nep9tL//npR9yj5WvoIonYKZM858wRgA8aBxPzsP0SO
INIqvyb+W2XayGCBNlhoEqILFZ1NSZFXC+cJTAatO5uGOyrIByRyxaAlDlBWwNeG
2iWyeZq5Z1lPEA1SnkwPIUFBEiMv7T6/orS1XbAKg58k0gbWdGopeBmA+OR9nkAu
0bXM2cPOcHMY1/PM3DQnHiMsexIZQRgQhAlf4jwout4UwRQsf2QaSPoWIN85iPyB
vj46iUYF5HnmwMazRvHgtkBDWCdPC2z29YQ+vHcYrPCUYaX0Sa80WG0Z1R4EVLj1
2MBWSn5HVa3kzQjIfvwWX/eT9EWs8RIi6EZSN6UZV19IOWQypwJPc3hKJsYqtVTJ
WWV1WpaA+r/QXlfysBXpsFeV061uD+lzYjYG1XLHQh9PIleb760uh55UtjBj4eUe
NJ3rjHFH7WcpFQf1qt95W4ulWP9EtEtWoDQnkkRYwUTt65xRBLcy3ogmtltPpDCv
PWZCEI5WrgHWc0BROA6+krrau4ebuQRc5UDQYe5l8qEkboTHzSWYrDIwnUy1IBsq
FCITHEsDLykUEiHFxOWMcs4RZy5OGiuPu2gDIo2lJ+M43KvXZ7eo96DuDdJLBCcp
b4l4fgIH+ioB3gRowQrXn5YJ8ARWziDF89sRVqk6kumQwJLZmPPO54d/l6J6kuBw
XBb+GZf8wgQ3jufBpsT33Ip0Fy53Ad93ebfhb1k8sqfoV7zwDkx4q6O2VzWt+rOY
8Ce4BZxmNvWxt7+on4OITx9ONiEwsrO496U704zCuLGQ0P342LWtdGX4cgG0WfAa
Atmu6az+s0tVGiPCSCDaJ0wbH2ZXwIkBjlW6r9am+3hAkylDNSQr6066tUJbHYGG
De4TluIdkiL3bGNoHZH+5EWmugVAN4V75qjuoXkF2tPbzorG3JKNozU/sDTJaXBF
ItV7+L8jEkjBO1vGruuwOaXA52ZlFuhBbaw3F10wNklfg8JKo4Qc3HYuHAcLL5U4
pmfW0OFUSVek5y6v/KpEmDyRKf+Ce+8mQkwP34346gJfhuZZ/t8dOkuVfqnTyxoE
c46eTnGirOcHnbSP7UYGlLxtF3irVqE4Va5yFV4JqqbfOef4lms+i9qPeFwXDlKu
fYf6bi6GQBTZ11Nl+GKDsrBsisJpLww8nmO+6HXLSr5pcln5+vzFj9ilVd3/X9v4
ZgxCRaC3DLcIZ19ibKfBZb7ZF5twqFu4Jw4/NEQDy7VZraoX5piPsQ6m0CrWIJKm
XK7dOzzR1PBZbZIOymWWVqbIaGUs46jpJlopS1cxSyWYL0acW5BxeNvNbwPeIux/
d+4xfmirNR1FJPzgRM3Ndzsie60WZfdwXFfLc2GR0x9Mvvq2irm7GkayCFOSh7gX
ZdiFN1TxyxNkoTQ+3jEDKJxWVWnrBfeI25EyBQBOAevyh/Hv4OdvGzOYObYc3pT4
cOz2aP1Wn9L8HZVGuYcy8QNY4a7iQ80k4MwxnUWaLVSohDWZ/k0ZZnAOywHRh2af
trB/hV2YW07BnJtM4tEBxdVeW5ytcsgjxLXTFDKmsvwZqK/sJOzlZf3BQWKZxq3r
insGzdHdhDDZ5hR3ZYbMsHW9R9lMtoAUOM2dRo7J21f2zOn//1DFVV4ScJdwySGg
qrhAqAJLKDa6JBVuT+FfzcDDmRfJLc7MmFSCGnBBMBxaAaGJJunD7NtwdJcK7dZy
/wTPMW0lDO5ZSJCd3HXwZuCu9vWOwV6KRwxITfxbNIqI10bVC1adjnjOC9VEb7Gs
Z3/YOWdkAb74nixxpa2Lbp2N68ZabyTzus3muZ7+WLBj4wFNhZd8UbyyiooSHA7V
PLKreeRO/FtY3WvaOV2wt0A/++jRcCzMRSbzZ6RiaEWtu22Q8ATqmDrk4MQBgMd7
zPaI8/vQlG9vIsQ59jlfRAhsK/pPRg4Q2e0reSAT+4Uipfye+G8uqd+DYFlJbmDP
2DyJjdjWjL8GnGoG3jk+ygSzdNXOB5BvgbsBrA/Yi4DWREhXC4hC6b85TTaAP/17
YXIybOCuOUNJZHsCxrlYrEOUcRK2wpxa7+/4YQL0JkV5U+GrrzwyF2b5RhWQchvj
4ZNVF/McXcXU/pCSjoc8ncQyeH77gE2xQL+mZNmUDk9/MivQYoGFqazPsw9sW4wi
xFMNwpxGuZVYToU5lSUg9vz8i7RjOomCl5F4gsHd8s9JGvCCjgDhIAnS4P7pIxo5
mOQFRbQynnYobCG2dMwyqerNVOl8INNmLcVLk/yKW+dQSI/T4Y5C4Ep8jvUT2VI+
Cc4nKSlM/hgs71BV7ueZydTVsSgbgV8wFSEBN1pv7f1Maa1nRwK8p302wvJZfNs4
84Cpa9+xx38HKx3LXyXl/YuoxDtBA6zQSi6qZ0Mk1qaaql2mHeaXeD2asuMwFNVM
p6/xhhJ+cBHrgs16AZ3JM5vtXFkMLqH8mhoEEivJLMTqFdGiWJuCfDsVu421YUlX
wgpABmz9CsYYh9xqK5kMgeOKX80ng79MbP0XTMyUaSkMoC7XX+0uL7t6r7ASQVph
1T6zWnfdfSd2ntOUSdQw7z3tX14ouKaLzX8+kWl//iHN8cd9Ll6a0M7gVbsdJg2i
sDKQt0jTQFR7ru4JQvnKXtW6NitXIB7zl3Xij7XvyjHq6kafhk9h4EWlotZwdCHh
YAuQvjax8pMOLLVQ4bqHocoDzC+gYBKhoNj5dE5CGODDKCQPRO1nvrRrWMHIWbMT
P7IBjSyTI4EPq+AlP6uAYy8Ry6NYeBMWla0VymCUbKrUTNlQaoCZP6HIN5jRd8nj
Z8JnvQ7JoOqoyJkoo8QKBmZu15aB5U7p1MZ+wORBt9GAxIk04kQNScHMf/NQ087G
ROaB2PtiIlXNZizO3PN5PCmD6uMk6pVQNBAsbtPTt2CeYP4jCXhWRo8gwP0hubd/
YmklIlXHbeImbsmHuJPJNm2UDWh5VpQdZz57jlKy2Dn2jFs+lnc42Ese8kEE54TG
E/yU00jRBdaaR1riNJq4n5OOFv5h7Ekisfad2PgYFhwtcCgbDAYQvtk37O96YlwD
7tyTHTVLUwhcH7yzSPoqrVpK9n9gXUXaei9dEVL7DnFrFh2am2v12Q5r8hWC8aPG
9I0jAievFqHR7wumFVTYE+SArpu40uk1DE+B+tqWeEdz4BnazeSXoyje2h9pfy86
N4pF+q5yvR490AMphtb8RS0gUvi5SAk2VcF/Nu5W0C3rp4PJhXQnUCm9IVR94nR8
eS3DO7UmKU91pXh50NO4hZDn9QG8+cbLPtp6B7oLLIdM0N7EbcmHYSlspodfd2Dh
v0foz8R/ySgvuRz774vJ7quqPiqhLkLisCr38pcpHhTMfrV55WCYbq+tL9lnwGQO
uXkzBEcsbzaoANvJiJNadt+YDt+reYTX/VP9rCOYPAJ/gYq7tDzxMdQ/1tVQbvAy
FOhbjRmP1Db4COnbswNCb9AnBdF/jDQ9OgU5YeazJAJRq84zO29KeuNW0YrgFu0Q
D4G+q2gTICuXQ74ybBhLlL5XWVQ+2VKQWIJQ7WJWdY1xektJdzcuGOCopKDc0fOu
H6mhmRMlLIdHIGODpJTvCWbgNZ8COly6tog49OrPXVsUuhEDo5Usd6I5NyIqSf03
/aplQGC8GexTHyepDZt+ptijnPFdicgeRJfxCJru590JjFAHaR13bOwM8o2ruWJY
9t+qndq2ZXdEo/thPzvzn6n6k8VOAMR0bDZzX0+lhF1Ps+3uaSoc+q4jpiu4MQWb
Sg5EhhkB6L0x+qYTKfBZgjtddE4+/gjuT2fnzY6Pm9G5V0pbx0I63rQib/AlM/T5
g2Kst4Xi83EFog6UE+Lj0cAdKxLClVQ6wHHXSlNhW0yBoxz40bXVG2zBOXUumi7J
2xK5O5JenAuQ/wFfjHx+uSO+INcUILYsqh0qAnfRbzpSJOj27oJ9W9X3vHNuFaBJ
v7IITaR7BBEZPKZ7VGyYo3PeotqHh98da11o2Ocv/REy8Whf09KosTT4axPZY4NI
lOC6UlaP+Fe8lVqAyhj8KPy6IQgEGLoqeFR3fP+EVut6yVx95RjECVDWAVJvkJqS
fAlOXXINLEx8jbZFUqog7I6i7hrvhyvr2q79QmYygusqvlb1+vAl00Gzm9DQ1cVx
J91jWg/s85PBfhZ/4F4IA3tRthN5FukYI3Je7P/PYdAd/u2OHGnoacnueogesESw
xQocfz6nl+bmQtOOTSLRgzdSe0CbPl5VT3mMKHobDQHpNxYxIvO1kArq45WhS1Qg
HkzwO57F/K2uFKnCcYunmU10Ne43BMcBzDbcOEJUlmypeg42p8EQp6CUCcfH90xw
mp97DH+udObhjH2cYrzxwmUkQr8FlqwgG0DP996/3d+cRj8tfh2KpRq8sMT4gXZ8
zBxGH+Dl50XYBpSAwfkHxK6049NKIP3m/oY0j5naE3y2+zx/+hzJCQtLFJYYoF7Y
WFaU0KKicOD08ZZj2R5fUdK17FKHpJhQTEdLI80z1pVgtUUEvr2uhWJeYXrylNpL
j9z4wHT22lPm4E388yKfBWWTLK6WcY9t6HRZLowagMiuYpD3kU8ApLE0Mi7b1tJV
cv7EO70KSu7jqksSAN+t2s1SLo2L2zKX46gLW7iDrlo97lq2evEEt/0VRQf4GVce
F12CM4PAcAkGGfKL7sc2qexES9FdZphvb6WXTeMZAfCL4OZU4IZ4rvuVYwoWGq4x
6eEP2xra4l3tFU0kBlhRjSVtyxT6X1FxBcKp4uduDd/31jPK9004fWqZ8ODgZyvP
W3bcfTzN4NI7LBtRQj0QAi/qMgnFyCqnyllvrEsvXwbed7vqB+jh2DyI62Uas/cz
S0fQCj6GDHhtPkEtYLYq+v7kWlU79NEkT7NZnoDUF41pX3jX4uM9mowRYLHjaHcH
VQaYwiYxn3M73IGBxdqAiEqAC90ahKDcluoGLpyoe6iRI8pNbByLtxSSPmaHFB9M
1soCRkzce2/+NTF9E/0HyTYU+y+WHkAqeZDJrw3x3H4G4Gh9fMdmMvC20n2Du6UT
ls8mSwNd4e1eFeVvK16p2TLuhmOWKRyyVnU2wvf61f7MPrCGvue6R5jg2aL3/Jq5
/LWnBZKJyim9umggeIocVd8foTzVHsa5+v0nNvY9EiAk7cy545ZDVkgm/DdwdokJ
PoNhpYLH2nuhrRW5IiG9dP6NVezrp5p0LtL5V1InLXH/LRC+rl7vr3UbHZjdiXdY
/8mX0E3rbXditxq6K9FZZNZQggw8kn4fh3Ctb3/Hv8yJJ5SZbHHL9FlYuANZwrh6
udodGjG4bS+Qp1IGcz4llQ2xhgXWEM0dNe1+3q45bslgJqe/Ua+QDGrUCORFe7K3
QkN5ya2jV1s0mFdHmpYUPH4F91g/GTEJI3H1HTHnJDUBBTYsfY+J2wCw9lq3xDb2
17mwrVnMZ+vRGB84Qfu9DCkFGC25uJ1GYx0mUvwbJgSzUiEGu3x8eSU4lr8gBFIN
fyfD6tawGfny/hUhdrDKz3cfZS4BKnK7OQKEdlFW039Cygo6N5bintGM1FCY6PMx
dJLNKExkqHJwKMKI60ietyDNtX7mryMuRzmWpHhq4QB+VfXF3daghF32nTztWFfB
oUCsQgaVFIXXYUVbXC+1sdLHBieT+U7ufLzCXUR1EEQu5NR5QMIlR5oTaa/OpkCQ
+YkY1REx1RpZcU920sCRFCp6UQc8kkStOyVLpKj70/ptLjKkUHxFmwVAl5zV5upA
dpYEv6KsJRawNo6f3GQ+5JGYfZAa8tTBAPg3vIc8qm9AaCm/z38EdqlfvGTFGJMa
7+z4xCGRquTuhyqfdlNvZlm5IYbmLMqKsJOVTf4AnTSRD/wHI+9Z16h5VojjKShL
mOzjIZSEAXGA8Le58q26l5JZLl0yFx97yuYU+cLj9KvTFN7dhxoVjmGzui/45PO+
acmZ2JQlMbslSk9D4dHSfDXhMABbWXBADQRXY6rRFrdgOCDRu5o5Q1alS4o67ohV
6mnVmY7PCUVpZzj5Rie5UZY+9z2lLDMrDQm2aUPjJBUB8sWP+ZANUlrPkGlkZnXL
Kqy/8UFZDHnufXqJJrRi0CFLHeZcIHnW47X+9GISyPGwNYLrGKXqjVUv/v5a5qDA
LpBZ3jIX92ceZG1UkpbmYsgfvJQYufTPE8sxs1N69HIieVIDQo0JLyvqQBiJhya7
5yqhsFjp2W9AYoBg2KhQ3nMpXVy51RSWH+M1Q+LfGssIMrn4kUEiPyaRXoj9sYmv
w+8eka0OH+xyrJa58w473m3k+oF5ZnP5D2BOoVqfaed7bbCDrfBcTPGOjz8r9Bnu
8vNYIrp+PRhBXDmdHkvtDlqbLnRhtuUfss5XXcWSEUU930IOC1U1etK+FZwZemsQ
T/8uATbB9KPDMZWMQNdVU13rZ4994grOXReFqc/Ank9AVQ4T22kLaRq+LBSUk1c0
ojnwskDr0sxrlRK7OS7UIiXChiAXV9tdG77TRlpQpacYf5AKQhBKIK2NRhL4lHkv
v4A9ZmuW4Ku8bI9t/ZE7SE8JVk7tjHiWn+lCY5cvhAriFHtS8dvHYBejQc7rvCR2
4A/HOmrFPC1V/SYSzydgbtm+dsYIpKohiTV0XtuVWEqb46DLNlSfwyBA0+Kl7DSd
6MhDQJmdGu4/FFu4e1mlgEWDtNJkuEjq0PZVWDnr2r3kdb0YP+QvCzfx3ZJXYcxj
elNtJGtZPtKxkRxXNswUVkkEFj9DdZK0wrDBODqILHDbOl8eB6+mBj/lWyp2oyP8
hwNkxDTFx6ewc6stAJItowfVnlj5pcy0Qg4rhzV9AbA8qdGkeJBhcdJqOSQl7YKs
tjqF3ZJtBEeX00eMfnbtihR5nBSa0ZFwzosfF3FLJMj5ACpgil2rDDp94Qo7yx6t
yIBxMhkHkYwX2lm9Pwok9oCEf9fcTy5p0kH/7GdP6v8Zg0grACoAA8nbsw2Nrowu
CvvzFwXZ64wDe0kauiUzudwi7QsIm3tWaj4tWr2MytEZa5V/i1aD1UUOqVse42Vg
OIV83C3/xDd3JwQJipK/Nx/pnhypLZQ7swXwbTgMgTCuzA6tuhJx6krRPAymryvM
buHDtO7Dq7cTy+MGTTLY1PUJYt4T7jhmLzqQuKY4xWJ4bXhhCHWv74TDhs2kzszT
N+m438TwzSE7xIcmBMdyHS/OFy7nJ3lu89hI65vbirjUP7V3FFEAnLu18cZqNiEI
EPSZ6p5FHTG5L978xhSfMK9Oluzekl3XNgeSHkj45WejEFiNlm16JgwlRD+npfwm
kL+AMP2I7oRBeB7qrhjJVG8U/hoZoJ3gJ1sqL2dZpnLnsxgx/Vt/RSILiayMu0JQ
hd3eEMs/61Aru9bVIc4CRuySjhI56OAo0t7ZQsJETPQfYoK7/0OIEivBmb6jSrAp
wpgfYJwV3k+LomxJvZqMgBHxmU7NuXFr3MJhdKyzESOqYLEMTSJWh+0l7vhWuu/w
V+WaqE9GtTr0QYYMF9MI0E688+lvRp43cN8W/k5Mn/j4RigKftUrUukZDQB8ZqVv
xboLch3ol2DOnUN6Ns6FsNsvAfyPMD84KnxI8UlOru3PiOSYK0YREwfo6VIMOO/r
uPCZZy0jSKN0KZBBRd3yI7Ds+FeQLC9C54z0vnAu9W6llIkbUbF8DfU+MnoNYkLH
qqd5r8nXJMoJz3ESuuD9IZg5XGnXGfBiAhcC9WiG0v9IXh9PxklRtbeq7k6NAf76
z0BGgz+6jTdg9T7D79z2W2vC1wiI8BSD7U7pBo9qdMjqKyLk1Y6UhMFvWNzM1hNj
P2vtbIXc7fulwvQ+ZspVef8KG2hMvIyNUFCXluOy68pSKpOdCzINRu8poSRijTdr
5nMRyDiUm7Pa9vQjln0/jF2QhFxQ0aKkV96Dv/jfhLQbbrZqgNmayJ1agFAiOt/E
Vj+kZ9bjNs5cPha8tfIAfpWAir/TVByWo3V3aomx1jSWVMhv3tRWZj7F2TVNJcmE
fX+KNix17z+GOYMxh007AdH5RFV2OsNMgz2EYVVFCw6/GSYWWMQNY2AQnR+Iz5wM
vqZtsgWakd27vcaGzQNz2n0/Gb2MMSph0NDFkKbq85Rm+uChxhrvelqR//a2Mgxg
7LQNSl+eWrsvf6oH2ewKZcIFMwY4UXjVHdz9dI19TT+7o/BZeepylD+KO4F/2zsr
FYjMto/hvCT4s5uuFJVxbMPnsdRuKBU02emx118mAx769ud19fRmYTmzxWAMh8G7
gZ+l71j+r8EayTgf2Nbb88bcCuv38EDsxudWT3TMhR2nkyy4PvEq8WK2k9glWViP
czc9obAY/bq18gsHGZy82zDOVpzC7iK8D7d5Vs/9CbmIA8GYUlhDJxzjrELxZWhF
/ZtIuzcntiLK/TPJqlnWEDAfatHKWEZ4Fr+Yp2ivbilfAoWkT0UFE8aUZhvLs5zy
mT9cpyDNHlcmPUVLMtXtHMlqIODBu1dHjtxUldbaM7ASmut1+hmiaJillzjV1cDE
eB6T5hVXEsp1SprF5N3cUEhLGtnH6wUB8xxi/aRSLwrL0XcvQ4aiCXvV2sLySZJp
dYkszJjDJW8of36akqYaTdbkUWEWvSqwtajG8TkXajMWmQ+AWWgS6+S6A4deViNO
RikJiR8yIf5LKepQj3/zbiRLtu10Njz7KetcBzaTvYbIw9x3CV5WIBwnEhH7x0XZ
kHP0Wo5LYnxIvRyI94baV0RLNZs828rQ7xZm76ohAOwgoCRxE/l1wvrXzLcOrzb+
hAPfrXKI5D8vFEzfVwmHrWy6fSf13nOCEarLhAKMuwAcGF9EQtWaJdVK0nrN6Q3t
WyKxkYonRO3DPwB1e3gXBjiJfDnUB4C9ZqsnM7JTzOoya+230oRvdFZsu2DqiECb
uJOoC25RLiLhNbegUr56PnLfHQAPOgmhleOU1te696Cucg7MgGYUreyYVHpxyint
R0utgxfgy3dZfzuqiTBpMfKlRg99ggpbcp6hfUQmfXATf74glAzAUq+8ocylG51J
rT08DlK5rXtmitirekGGtwygpciMvfemswuoDW4H5P0W7jBAbfgkgv/6jGpem5Dm
JY6XgH80DyFEINEqkwths6LGw0TU/wtsadp81e+wqdscnP3/9Y0w2Clis5hWQ39V
b9W+xcvrESR3SwR3WZLdeLRxFZZMBXMKAYgnXQjlf31fimM36Zho2Tme9CoD1YMQ
Fa6WFZzK7bn/gJUUOr0aTUmAbKhZOsxEpwuaF5CwZ+WT0uvHURpFdqqFL+Z/DFm1
jXkS/DqDrYWgZEFH7ZEubO7OmtWaEIwOaYyhcTf+sv20aZLR2vT8Xg8Ihsue9gWL
+2iDiVgie4BjIDajqS4bL3h1V/KiA29BvGGKMR6VJsjN1T9RkO29TjORfoP42OSV
FL4qzB2meNKPAREGDW+nVaZbGCwCBLVgYETed22Zm7vuzZbsrEFLuDiyRFhS03Ot
19eRvIxdWZ6dJOyVCRhruJbtGQi3BHPtsMyt+H+3G8o14vifuQbDWJIaFDc7PkZd
upw5A2v8wD/6lOr9RQ+7wDzMDfzNCxI+iN5nBCPGz8C+82kRfi8uLCPmNZmWDski
boMNxaRg+z/7yfcPTmKijimd9SQJZ89CxJKaJaknmKw+rTJ5ezS6csoAi7YXDIwJ
xZ/WNGrR0Mn87yvwzCqjLY2R4moo0s6gspi41jzreeiXw5zUWv6F7WjEruZ8o49E
vGDJYobvVAc1FLwVWA9oADTj9VRsIKlzJQ+zTgPBXOwoGF4WH6oilP4b6rvlmaEg
Lvrbo644E3TRLJohDEZXOMJ9P4xnJ7Ns2ZFOYxyXIYnOqgc2BpiUwMy9f4rhmTOz
741CslH5qEbrFw3XAs9NR7meoAT2eFZLoYh7emBtx/+DZwVo9OAdvPnvxhvayex+
vX8y8aG0snJxWEQ5CV2lj1xqg30Yyh+SWaPbZL+7EQgqBcTf5T7aAqZCvLsNpq/k
5Jkj2xx6KJvC2T4dRF+7C+7r/wC/arUcObLtd+GcOtaHnM25HubghdJEH4zA0L7D
HOuk+GLxGpklUG0Q6Iw+DgYqAFMWBfLu2G20fGlAHw89RXgSxHjVVqUBocSWlVxz
/cWcSwcGFsQA9+glAQq0w4BpM4eLHocuanDX4Nc/8F1hvOUumM4/DNPCxKBsw1vL
tpTPdLrTyaBPREDWaINpd7g/aWS6zvthtuBZ832PKW0/TsaJCG2wEAksTbDHeoHa
7ffDeD1d70lA+es8Uxjlu33zz4USBcUhgmR//NX7Kh1fPCTW3p+Y1C2Gj6tsf/sf
nRbuY4xEMYZy5y7Sxp4vGuwJ2qcWUu1fJJX3mC3loSiEz5P5s4gPFPW8k2MqebZg
VteQ8ZRckzd4wQbu9VnUTv/NJZmQxTPZWn7ZvrGIyHTxTeL0JhPey0WQIiH6KU+t
RyIi6ePw8rUDmmxY14rdTSNq2Oo6XBqMVRqs6u2HFJzP7xu4cBz8vqTZRTZsfJaW
OKf9uDFG4auL3fIz7pqK3q/FMyLeMs0x5FplBqNlJ1nJASCY00o9OtyQ0NDRXrHr
5WJlHf7waHRhhXyjVUdIMnIXE3So0PKLcu+Z8g2VyYyIpIAOr9NANz7johTj0CNg
QKbHbv8/RpVP+V2ZVbjBevWq8vAy40oo8cMo12MVKyVyyFtXqXAjUmzqrzRJpDJT
FIc7uGgk8IoKgXkc7mrY5GsBLm7mTceO/AoYtq4qGE5WArurLIC5+j1gTn1bTmPW
kMRMlu65Q4whh0M4zHTmWxqWHJP3lZITG1xq8ymHvrNWjeqY+mIqDjUNOrFDUjVk
fn12toZ7V6Lv+oYlS0pCSYLou6rSNuUAr+7U22Zpkc7rMp7tV6truNVWVnbop/0P
KD9SzCZBehsMoofeN5jPoDPqeYCtDRyf+aochRMUNbLPx868DarkZDwRKZF7gOg2
7uWltAnj7OHJ932kG7pcj6oAWhHjjkTDNx9pEROdT2rOJ2oZfdKPggGmSRz8SGDM
c7wW3FJfm//20YYiJOEyilTxEsdg4mhVahYgOFo3IraG5cqZGO45cccgarYxmHhU
5hKYu+jVNDTv4uqYhA74j72yHJfzuB7tjiHOalBgU2bca05I8cBnVMtFnFTNUBVQ
41NGHqrKqcmh93s4dVi7CMpx2hX2smx0TVe0MB6OYG22JCcxMmiQVEPJKT7+to5I
x8MzZES31sPfQHcy1rxWVPIoXe69FovPb7v+E9RID9k3XB6KIREzc0ae1hwmnMAD
XVJr2uvj600SE2N7cc6oa4mBKX4ji4MmFcc5AlCYlShrkoDVuJ9Tp0Cbf75e09tr
xoMYlS5PeNJCgr0E/+veV3O4ZW5oots67TXoFc519AM8H+f9bDVu4kGGHGf7JLUR
EpaN9IN5uJ17fpvyoyVE/2YL886+svQjdQ0FyQaIMc38ESH997RUp/+tAMp0TnQv
Qhs1KUyuAxrXrxXZtZK9IroK554DTYyZ3v2QknymEN9CyR1HltqC53FUg0iPnSZc
21VeQpdbZsAKPUEGMun4EtRnluj0plc/icsQDXwYDNk+ZgKmQ9llaCK0zqyFFuLp
a9JpuHCu4nkATK5ge9zD8QkWlycdZ1tGPsDLeaBGaaNgPuedHPp6MivPeEpVpv/K
EpmpMsEFh9VIsrQu5ynCSmWlLEDViaKwQknr1x+iMsNFGbrbxmDRTj+dpIyudF/t
m47uJLpNjxd5EqrJbFNYPZKMVQ+cuZDY1N19/5ZQGpSaaZh48C5Jd9EGjNLbj8jp
eWwK+oK/p5nAztMRZSq6s/3vWeURfvpzzbytGYoan528eMYqVq2HyZo4Q5V7SrUh
tyv5WXnzI3EZNLU5z65TMEzIu8fB/pDEA2VlGiZu5N1neQMlya+YXUFgBcFmqu5E
85OmQWLjxGdc7NWo7JfdnKhNof425oOxgDkT6/RNHTaOkNVRxFqGcciJXS9EirhB
OXokZLv7Zn8LcCPTtaxPxSkpw4eEh4SqApVEa5HKG55S0BSIwb1YkAMz1gHZ4sL+
tFBKr5TU0G6slsOZEnB4BOJXgzEB375RIWFTNonQRtcnyrTVZynf/8cBF7IyGVT6
jVzuC9GzB7H2do5GBGWiz2Ly5fUSs78DjjgNlf1qDZOhNJobPJbia7skeXqaVFTc
pubE4KDHMBRNh47gymlHwFfPifk+9QRQ43l3QAvpJAjysSJ0sxCSEz/QBxZMUHkp
nlNa7WGgB9F5tPGVzieK+AHhuHOFXGpnkFMvd8gmQ9uhyuGM6FUvM6ZTH7OA3Nua
TNJF/+Elf5T7i7bJYgbNBw3i8QXH6rN1tSUqhBQJhjpBq0yxIbz9AzzF63LWpNid
T5EU/HDfpHx7x1BH6XBYUG5S2NuO3AAxlPBALWMrLnXMoYW7z3ZjI7syYuYk++Cv
QAgewroexeuINltvRg2rN2eVWuAxwHuOueBtrnEG80zhRJDmKCAemhvT3X7fHPbw
eQu34scJEMK2OBXNwvkuLIIRnMevwSrBecOYkI701dU7DYPqCPOdcds92DlHbVuk
bgyme2TJYk4SdSEcZA9vx6QfDRMD62qoe0NMR5tjQI07Jyq/7c2eJ6/sOn3GVRCN
GS21j++x7Vw7J57J89myNus0nour4xOEDR4mx/fOIfw92nX1ObTuLNITucKE1rr9
75suAcHgkkPdSTYEHEAYuSIjAvJF0uEET/zrhrUnX9SfEm8nY3E/LqGUS+XuCGZ7
fJbyxWjAvRw0ZJcU+2K3EccsNpA17N3DCtlW3pli+co0Fkm4hh5W5BEjJzlUBFvm
K3ueVVo0iTc6TmVj7x3sLwxwySn1ONJLAyVckcruRteKh9vqtpaAkKKHBp1Q5DJs
pQQhtfQJnBnNcESiUqbb020hfymtuM1VWsLBM821iWHnvp0otxTdcUpzUCWubn2Q
3xs/47PZMOgnX2JqJZizL0Olw06IxeF4eG3MbYivkwlMtOPGHH70D/8iBU3Rk23d
mfPvbKLxJEShRU7sxhUztcaBZBwcoTlyQ7WIF/C8ROqhyoRdaFwqgKa8G4slug+V
6Vq+64ED7mlXWqvNpcEudS8VpSMY3ubeAQmQUNN1mPHqjAN8aSHvhcQh/Ul/JTXK
zKMk9+0qvDlvfNccSmbHYipmBr6G2jhBl4anYu4NsFn1mjWCf/p7LXhVoi4y0oR5
IVvIWplagC/EtjWrhguicw22DF4V3zdoqJpjixvmp0doD1Gb+gFItKs/xCgqXGrm
eDXxfTXJdxpNOqoUPU02ld87jDVfFVVYuNyEehnASFW2nHdSmtcv6AQ0qE2+28Wx
px5ONlkjhheWvoN2vYOTttTUiuLN1k9lcZHKY03CwmspJgeZmgHudxorGNSw5J/V
fak4T3zKB734S1LAb6TmnMzFKoeuRE5LvISbBK5/e1TZh0XEvUo7wzrsFQXD6AuY
/w6MJDCRNc21Euy55cCSZAGLVhu6ZoRcmCWhhj8v+gMUP2mMZrXRrAaye6hJUDRK
VuFrD7mY++1qqgO+aXIgiWLr0yrzJqy1s9PeTHT/JoxvBbsTk6p+p1JKdK5nFbO0
SrdaFFUx66MtFvAS71kpAPPCTxlFzcKa9WWsYHgkHDa8UI01++O4RGbrvtxbdZCr
jYngUc3TbV9AHw5hJFexCcRi2UcUIYRp7Nm+fd+CshJnNb0EQxan9ODx+pBRQzVy
oNLDM9mfHd8/4WpNehTC2vCNJgnRickNkwq9nJ55L9wsgV6H49KtXqJMqJzJCl3W
wMQAfNZV2DWEA3a9CaFoe8/hNpHb6HMgU2iVizUXrvTSMRq4Hu8sR0X9ZcjlKZI6
Q4ajM69sLoahdarQPtfSCj08EnZLSV+ZscZ3znO1feHmsdxf+pN9hMGt3gbmALDN
YNP6ZsHf4/n0qmDL3SGTAOEr53Ww9mmBvRINxdoVRvHOVVzZ9zFFyU1C9wuCUYdI
VoSd6TpTFCLboAeg66CembBYjYwxcNm0GZOHfWSmT57NKr/C3hg+rBH3jFdpLznL
biCBOMVef4FbxVq23uBZP1P0yuerrPzmk9yoOztj6Sf3zUjc+z6CF66xgqrVUPDC
Ojoc9kDyEUzL82kwZGmLuR4nNMtKEURABiX8AmAyPTxnihWN59XLi5nVX1+N4Gqg
Ajz3as36JMt2AshRR4aMoCiwgUZt+KGDxfFTVSwCucD780fBTibvbdqLpNCKgPfI
4dctJsLnc+hem6s8RtQS8VWTUUI6dIOZmcqTvL3iqTuzMXwAjSV+1F4QGe+w5TIr
rS4dOqTFyIshe+ilQZymZ2Y4FGNvSNI07opdD8yzF/Jo7EUjlgcV6fxhbLUaRGH3
UajjKbEPgHpquU06w1su3dBCncVPvW6oYQqtcLMwqPWuU1VjBbzdo+3YapoSk8TL
IkKGXQG6+q81FYH5l8y2cHtZFOdi33XJAqlDbtzanuHVBbRUjz0BT7JkdRxiNIFy
v5QyBX48OM7jOq/TKrxZ+lzkhFvh8YepHFDa7irlGQ5dPpnazTOMEZMLyLuXUcXb
tOb32rmlXhJ0taJqeP3RgXDX5Ceb53bwWa5XPJa1SLbI1/OkNfkohT++n4bE7mg6
HP+aoOv9I16hmLFrmWgdBue7mwhoxfed3gfUhxMaS0mt7t68T6YWdBduXJQsEIdr
osDNKYJ3RBQyl4zTuDRAJQto3ZjqCeaoP61k3G97iry1qnhxrF8OWev2YVVEunzd
ve5Dka6ws/VqbdNPf50QMLh24zx2vqKdYVTFPJ05KbLJRnfeTcKE/Wz1SQ6KNZvK
o0wYIFp6jqUV9ElSfZqkOZ81/slHNPdBPz46gfocixi07rwnfr/Y+scksXTkeVN2
twtsPeVfexVlCtCAM0uz/aXQjQGA6OhvcWocDuaJ8th9tpzwZ5HUqEhMbw5+oM8p
c61c67iVY7IErMNlH9BvzfIcDmxsAH/fAxMccWjhzsCQQLlNxu2e6RPRKohu8iiq
Kr1orL7wpRcYHh6Cej3jLiqUB/FZV9NoZtDGTXhC9iSTWQ8JcNQGp2H6qUz7cVTA
mjwnyw05VrEGgn4CoyaywdiJ5j3zV1rWhxYEh/JiF/TwapUmQgd2qsXeopBC6BuC
3zFptQIHNi8IC6s2vwk9F1hQCxis7trvk7lg25qJadgNagk5sc1x8tLoDE8GuaUp
XTfmBjkCT1qz55JVc/vWzkKHAvMGKBsDVlA+BYaSnktQPcPkRYYZAfpX4pHhO8ka
BjYvTEsufBXNs26JRZAXymqnwVT9dgTCCqNbW5YmQ4CR+RbCw5VHeFO9ptJTKPsc
byhTeQKz3GKfkaNX3T2XpgLLECN2gZGxL12iSgyg0W2OLAQgtgm6rYEeLtAMhM8q
IW7HBKGwRCXfiuIOYoEq+SKs3ivu2NUXmF7z/h8zWF+W2wZngIq7WtqXFFeAdEIg
/b9WsQlbETkeh7OvxM5CFv+zRm1NhGS1ivFL3sClc/ZlBta+zangPhc+A9iPsms+
H3K6JxxXP10B/nmyBa5HdPcJ7IyrV/GGCewYrax46nxLlHQHBQMWY9GdlE2l3IEP
2b6V43+xgHKxHAdym/+8mejftlrv71LrxhF3XiLE1uOQ40a5YVYOzJkIFvheiEmg
25sCGQWOYf035Y6iX32mQt1obtRXugyZRIVL6lp4L1rv9b16L53J321roNd+ckSO
aXmXpyAXt4ixn90XAwIiCC6N/bC3NCd5qdwNujC7NBv0C2EsivfWjNvDjUINkWJ3
kzgq4lYLKooNFPxu3jSGREDHH6qHnoVghwxaZrIRg5bidoskNiJE6f4g6OZuJl2r
78k7bSObK1MQSVnRiBOjlZhhA3D1GvjHDHIe54l43jk/cNRcCsC8L7xHcmcIekpy
Kl3Zn9WKe8LE+N/1mkJf3JO4KGaijXG1GI019CkJ9uxnpvqnM0Ch3O4+Dqf1bQ4W
Yt8h4q0d80OlALcGjL6gMEiS+iJuo5uZ4ybIKIeBmpGYmDRA+5zzRb05A5G8U+Sj
7LZAstnagVBXZAiKz+gAM39fjPi1lrUNHjazxAayv6nhX9zvE65UbptkGF1QRxS3
dambzQ/mlraxwix3LpLy5eTWJn6V7ZYJjpRnvzvPcbZbOzx0xhqRgIbEOp7igCjH
VQBi42PR0dVJ6akyQh6LmGzHW/kYP/R2nM3pFOVRvVZdZ9cjbuuXmzneTSeY2CcK
RUnqHnLc2F9jro3PfJDmuHda/eHXD0EDi68uTPIoCOnuquEGPnLd/2TPr7ZE72le
MtbE5ah4f5+GmALIrBmg1K2zeIl6lpJYeWubAvc4kZyppIpuoXBx++AuZEzgOEye
6xJpyhy3WFENVza4tXGtxkyDkVy7eDU/NNRnicZE8WJm6S9kWRYJQthWLV+kV00e
9I0RSDzvUQBlwJ82VU3KFnh77z+5CjRnvmyuSTleGXbIL3BP/2ulStd0EtDDVvxx
LGvUQ4ah9xZNohRa3jqVsmBdZwl2t94A3K2IYusWxVus6/Eh1R7HORLmL/VJV1sl
NRF66QO9yw9l/aHLws5C5EoPOCKVxu5kFMAHi4LSA8z/qgJ8NuyRWIrBoOsjFLBL
FYs9uTDJ5/asqILaeAT7HMviBPDKsdmpgzVpgKhPpa7kP/zNX4GSkPPLD5Qk6wXK
TGF4evPK92FI5aeeLr493nl+4zZvJwWpXLV1TLBlepId4HhocU7sGTKvz6y+NngW
oP+mpj+CHCb9lXOJziD9/JMMgB7/1yWQTyykBoa3FDxCYOZk189vwrjPkPpo0YfL
OvoOiLf6W0bT981Y4suCc6TRYnY8N/q9PsigMDNFcYLJSf54j7GhgCR4XpCOggfH
cIR7bMUm+AKq1g0Xw54hAR8f43Cgr7J6u7cFZZazLs9F0jjinEMOLVfrTYQRrINN
O9MdqC6OtsniIoDFIvXqI8zpbu3vgjZ9y8DjET1qt6/qqes/pcxnXfF5uQx15jKl
zmT+bHGdMgEeVW3SojDyJg0XD6DO36YTD4GR6FjiI2KrYMe7quTQ74PPDasr3tZD
Rurz2bGSOsSH8/lxA8Yif2jxCx2W+HdL8N/bIn5kyuW1cGg2Sco600j6Oz85knjx
OBP6lrFjdvTTcHV1u43DMiFimWn5hX6fTM9ZFM2yZEwznb7NAIIYNV8m+L/7f4ke
LKQGZvfVFvncv+I6TkBoLN2lOOZGC6+bEGEbajWuszwa4BBOslYu0r2Z3sy1/MUa
/b4Fb6c2WVxwyqnLV/xWLeidGjUMhXi5YdR0NEljB9sLIAvTjFemqyWI9TnuloYT
2QYMdIWRTTe/xcBgrj20olnWFIw6sysEfeJ9pLOFuLyCJWn8VpTSXz+slE3/oOvl
9eDmKFinabSDttzcnaZV4iCt78vFWFDlmYuwhP0ee5kaw5NHsKnNJtVCnJSHVJRU
snhMzSmpe6fJIRwhUkP0bzGhyWKBXvM5r0YbkgBHQOAzb3kNUTPNY10p5etGweBy
Jb8E2HenLTh8P2f5BtOdtf5d+KJKHZhr0wxHWruwMz/Zp/FNbdH2pre9I02nTb64
G0wEPZTNEZHU8T7SUQiyyUTqmmjTYJs44ecu7UR9lVGaGu1kPSqYeIGHEIOKrCRs
t4sCLmSdzM1u1hJRJwj8aNcUytYOPjweaA/n/5qRDCYRSiQNba4Q6Va0pF1OCHIp
U0ge4a0Vd+tN+WldDpyFFAMYlcYwIeLPQmVLkqFp5fA/RRtKkrDmPCm/iKr2ovO/
BfDfsynG8ZpLMLyXBAq63AlpJhwYQ6CMAXeWaa2NudXKFJVZ6BSgqd62iW98NiL8
y6R2O0bSb8xY0JTWv0pO4DhkfkjnT6DZo/NVAvPS+Qu+WJ5me83fALP3DRuvEc2l
6lZk0chYf5ZkV5MaGyiBZxEroqy/Dar6MO0ozwiNeK6Gf31l/yWyI3fibSY9DoQM
pxrxKBHQgHXxt+DteXNjstb1VRIYK1dFGb8cgqApi6KvKDoV9gYIfwVvwiDnIJX1
E17PdR4naWHNTRXc0JigEjwHj/k41vGlXchAmoXG49z2bPNQ24OLcmxOMoYjg6v9
rnjkGp/0nfrPC/5Ey/8Uqk1pD4wvcAODPkXd69lcpjLFWuJjNGU2a5ZdjsmslDi3
veIm3/ymC+0jZCWSsk0g0eyz0GriZz4+oxFOz4B2HO9fZU6fs5IugUtBCOQpWtSD
NLAR8wNsFV+xNPAAvobXg70RUuOtap/mB0WVUHnasGTYKSlRvvRfh4ZB3JMFaaSX
MZAj7ETnhdiH9nZUEHFm/RIicVsymae6Fgn6G0KWwJvb/oq2i8t6PzpFzT4dZQ6P
2guUTIID/P6VGowFPcVFdKgvGZagaPmDJXKbjS9dhjpgu4si4T8mOeZpukm+/eOb
q0/g+fZAez9Nu1H1CprjbLmp/AVs43aYeEjRa9zCFadBPrpOJbwIHWIwHb1Crd5J
OkeUYRjzYpQ1qhsPT5JvUoArKnor8QYTloq2ELHvkhBWHutyJoRfOPGh5fLRCGof
c24II6nSKfMPnVLCG50wrmoioZD4NaciuQYO9o3NLoWoZuxYxrchIVXSJt+0oirB
zZPo8tb9xn9gmvN/xU6AIruxsz/L7cssbSQOrfrgXrOO+AciBbuHQey1RKV7/Hmy
LWEyG8YWky+xSnI5torzHXhKnlsCe0nGmd9OO0/ilk4ywQ/K1E18lZ+Kx0fQJzT7
vcfJGiNqUDiU9BoPgVLiEsr9XR7lPks4SuFOjRIqyhFY7KDxKl+LCbVSt/xtePIY
+TmCfIi7OdF91dYBfuAoRZdklXCCHcQgfVxpXku/Weq58ZXeRhlv21YQAEIc5vAd
gHvph+/yFJH0qn/2n+tD0FieyiO8vELGrKsRW/Jhy7h2E4uFCgLxzzamkBjbkMak
M5NF3pLF077sjw5o0+hOUCr9HjO8umnaSzQYyc0lHbk0bgX3o9wChPx7bxuQKc3K
uzxcV08jf+uNORFgF+FGJNWxv473UFpwDoc4iU7UIf7T5BNtU5MkPUSc0kLi1yRl
Hy1J15Ia57qWf0o83t9xFg+N8kHxpyLeTNEnOHCTYREJDKPV83gTuobAkis2H/xK
qsBfALHwat7JMvx/sXYsNkAeVRUhtArIh59WY974WuhIfOc+GGizoZ8bq/stlaKD
ZFOuFvw1wu52VFENRPF7CNDLE3XIVH3O2rvfbWXVuqAt8+Ubvs2Yz4xI5n38LAhn
Rp3qPdMCFIIvGQyT1AQCKpe+jxFDbRn+Y9+SV4zHZIO0181tpoi2aDHygQQzADqu
DYm1u2yVm9SdqLwOxbk07L6nq27igIZsSMxsuvkhKSvGbLATJv6Adrz7xleESSIG
X/4fycdy6wcWNEIRKQJHZ1o1tWq3E2rpqNkD+ER1wFVkc1A3Z+gxbFMg8AsnZEs6
2dl7LdqVvZ8XSWC+k/NCvEfX5aKVtCPLYGls6zLw7YC+fqiBDvmkn+h4rLB+KjFT
CapmiLdJDlaDPEoPV4UB3hM7Y0ffxROK1euhb66GArdJWYgHVMDS8OQyP7EPjM6P
ozw0yR47iIWwUIT+4Xgfzjz5gX6nj6OdNyTrtz6v8VTFNponFvoENMBK5K/20wZe
Rgpv7Hd7juzlEcfoKkhg76QfZ/4HdeZP023NPi/rN0IhcS3o6MZ56Pn3eGPonAz3
OW9c7t+QIxvE9QOT+VO4IDDTZUqx9ENzbXUefZjzurgq3osF6OkiLMVTIC6oy2zk
+Gy4Z8WiscMOKmiasLFrjIb8U45Jp2WOK0PzHG62Zus29Whwm5DKZvLhsZpmQLkV
MY/O+o/FFmBqlW3DD0ezGvwBi3xOZwij2X9QXASWjxBZHIjZ749q6n6K1TcfIyv4
SjwwqMdU/WLhWjlBfCrhjhunPXPl6uLUqdwFG0/lTfhpqUk5Erbgjrk7VMoHqE8p
9p/1UqjY9yTvo0Tm3xEwLgLmQPKOxrcT32asDz3HKfAHGspyzS+DFm3dlRSZj03n
fc5uVpz61uutt/oJgSI9sQAsIQmB2x0mgjzR4Y1U6KG/J+TkvG5pw/2UwT8hqzoa
mIBU8Zbr4PLtE/go4U+BP+n8z21OHKgsJQLo8XEjEHU5hKwBLVyWyVh0jjMTWlJu
1DT9xHCYUc9pNu2xWU6NVlMye1QMazVRKNo4KIEYQQGLaSzZuBpgy00G+SctKvjT
o+I58xtc2IKqiIRa7cMX52VrWoMx3L8ijmrpup3dgj2x8URypKrapRkmKt+MOtED
CjPaRpG7MTMqY770hYHIrVeTnyk/pacX3BlDYjvXICEGn81xiXKVW7Aj+QkTNVCu
NK40U49vlErHvvNC59PDc847ESJ0Bc3fXyEzv8f31+ERtlu5E2avQeDzIFKva2eq
4UBws/2sIDNcq5A4Hr584GlhhQidpfbqC4mdIe4Akipmb0WSX24bwNbsy5PDCdH9
vXwhTz5vF24AM929Z2+2UWSboAQ38/GQJMPo9O+mlqy1FrdbvgxxXSTyNTuMDpsg
13QvWSFWP9jr97m5TSh05ifP/aA9fEkIe8dkJPb7f95k4nc9xTPtQADKzjazIu5X
FNv2xeRO1OAYGaBzHeSSw/XFtwBLwE1C8CPlGPL5bDbimpxUZiOOF7FdgdjnwmSI
iqgq/RM+6/+rU8k7ILonTs5sZ7AOfc9vFx96JUFBFoOsUNaj683VThnp1VQRPnND
eJ4mdpmBs59OWNqVup73PxHKEWwuYmZrCiosaRPj+U2H/n9Ri3XZrJCkpWnZkhRo
WunKCA9/kpH4mXcdkIVudzKcjOKlbZTEsSABPO8O1LrO/U8r5vByMimgMeKFeqwl
+hFbDAmW+4GRsbae+yLqSkIuMEfX6r8u0IoutpSy794FZmSLnqn+Ki4J9q7z0+qh
bxYOpequtKcsSjtCO6e8NBpDvJuW36N7gmKi4mcOsoaHmMuyCaNVtWr4HPw5BGBr
R20+AM4rL1KxiMd9A0p/06EUMyBBS6SHvKy+mP8N+dWOmZuBJrSfKWzbfBrHhQH1
JrfUZR/4xWS6ngvwuAp5vPw2cHXlb9E7vowvTAtsgqXn8mE2T/33lUfarhaXtgr8
1ekqKY1cez2g6fOxm5Jcm4QllfE7xn1WLt3snpX+g0w4ZVFGwzbxeRjecyoeiYk3
iU1HT7RkQLcc20Ett+QHXz1MT57hNhdK3f7nSem4iwD0z2P6C95Na33F4t/hPlWV
EUzD5fW+NLHRN2kW56Dxxk2wd65FW4rLbBE4QIpHLuUfDfjU93j0sUJ41vp1Blxc
/ITxvHlvxsPEjFgrcMe6YMK7MrPDmi+E4dME1SDY+ArwWbVi8yj1+oNybFswctdh
BAP/gRAQ0T09HEhP7AG/8geYzk/7K7QHF/3ps9Y1NS9SkKeN1LZy0+FaI4bF3eZG
uZlxfrpM6Z05On8eSRQKrXZ5p409uZ//Zk+PSbw0a3rVi4PROxFiul9Sxz2HWOAi
cYORCC8yh/5eE4yjrttMEW/2r5FYWfB1hBklwHeT+QeVmCA2Le4fMKluGUI1plbn
S+whteblUAWpZ9H1mR+wB6ULnaR8cI2ne3uJkRPd6Gy/bWiKqMZC3jsyNXJ8oQ4w
wWuTXfSdkX6mPuJF2H1R/FtiFe9K+3V4LcLaqNCAqlZ9n2Cu957RuuOzeeGsrlD/
cJRLA8AeGhlKUdpya/Ky4+wbuBRMkKG5Pxl+AvtjKg47fiNq2ROFeclt+mw+UXck
qJvibzH7aM7o9W1d7L5j3jJdbadNEs4sWvgajfbJB/LaA8ecSMhCS6pa5tFcpK9v
BA0CvMxxGXizOXH3F51d5s/cSEuiblWkOI/YyOVY80VPO2nOik7WAIIeKD8kNsiR
F8voEr0cyjR2vAlQPR0Gb2KsPov/N79cNLIxBXxJmjWfbA5Q2LSwe9/kVM8eSsiZ
HihHKMeDWmFAX9vR4vqQ78gTkp7SHCXdTSzaDkVmGXvwlmylc9Y0XObEbrDxvybp
/+fSNMDJmRGa5OHgFsZNaCBqSbrI+OdFEju79ihWF5LyMbgrROAfR7vjPBKGKuGe
KS75BKpyrR4+yrTXpBpzHfD2/v6r/2BPfUR2EmnuO0+ve3R5h8Bj5mFVobJ6/OFN
mcJzLCtne5kMk3toaMNxUGquTJUGU2nefpaoWXF1dt4RG4rX/p37esNn0ytNl09B
d09cDL7hL8QoH/vK4eZZY0xW/WII6Pk7fQb1sT8QFUkgut+suF5ycs+lY63n+UBr
6a4zrpSmAWpEgV1DgEiItlehPG6dphrf1/EwM5kOXAHzRNflE9eegVDyBjkiFUaZ
gTKenphiyJJDbHhA8c8CuuaEdXzsQ12bAO8GIudXIF2sZVS4p6ghiikEDmB+PBXL
PPgQa6Az8cPw1ILbejb42u6XvOUjgOBaqkCsgJKVDfl/aKa7isOkhXzQEnEdpH+Q
w940b8i0IZiT2f5mNyDf5caKza1ONN/LbGdJPoYGdjYZGMVeiI0oYfbLmfa7arGQ
1J1eXeNjF56Xh0cgWiK7EkdxpxhigQrElwa7MvYfwuIZpRT/Iz1RjaDQWlpJ+8V1
P9BSZ4p158m2b53hZmyfPq6u04IlvAGYioF5qmU4rYoh/VJxpj8bjhLsX+Rg/3Ec
5xPxczg7ZBqxQYCF8mgi7WMBawLtBkCE5kQwLpXgzES3+tTkllkEyFaYbml8GaqH
OoFMQHWS6UWbjv2ZsKuWk58bUBcSvOdglMAGvOCPbDjaHC+uax4pwUClviRCUC9B
VmiIo/rjOkEZCqvaAfsJw87bkPL3Ma884fVLmWqY3gAtW3qm0zP/7lwD0rqRuK3T
g3umfN3hRfP7G0/FV+/X3BFAuUyMjiKqze39c5Q2JUX93/5UkSpPAeTTbu4M01Ow
fDQ1+as/RA/af51J3u5V1OugsGrgL8ClQcZEjoAmudtBCv9HEsJlV9SQcdT0I+2E
HpcEti7s9x/yoVx+dsWVRt1VzbU/T7kF8aQ+XjED3w+66EHC9hCI/3aWa+zQKFkn
kWx+lInPHp/hjzyStGKzugOW+jTk1BkA6MqYAhUtp8eASaUkmU/FL2L0huww9rNK
U1AbOJ5jfYu9V/9QabUrl9B4XefmxLYMcJZT5Q6rSuk/ZpYpkZa/PTElMrwIwkrq
juhtcxUsbOzb/cd7jwgfYExfz5kjlwn7AdSzKPzqKCfSY3Qo0FhDEYtvmrs/oQGB
SKouzhHv7JigHHyI4yz1UFzB7NSY6DwW7FM8X5WUd9i533X1WOHBGNXhgGdf240s
H7oRrHK9XmCd99HYmQpPM8q9fTHVLyWkpHzEMf74bsM1bvWTw13KwhWEh4bD988H
qAyUZ7zvzP8KiaoqKCpKuwmecDgQh4lbGUnzwx8WyokbBu9iq7W3hJMIp7m7QkOZ
4HDeAno8mmFQk1p5Lg+RIPhLghsNSSpikbkhNm9yOt91FKlvzVvN18B/uF4KNunD
ERL+0B6RWIzIPExfmAkU9PkXS6MbeSYFtGUQHN/DnwquCiXcVFb5Tj4slkIgboZ/
P55a4ZGUxc3jP1I2tbIExuhWLO+vSxKdFS5F18YyKEWoljczBAeqR5qtr/4fYHln
e/vrJeOAgteFbwuGORDDr7zKGCbYpnoN5vE+d3OH6rln2O7QIXZ9oyXq3Fs1Cs2O
o5IC83XSKBy31fOzvkjApye3msDNIicoUfNxeQdpm06ExZ7WC2v53DATEn7/uxw0
IjStpa5o3XdFLaELjUPBA3SykepHiPV8W7SZacXWGgpXeN46PceRQrTqCWilpHMJ
W6u4JK/ehmhf6/a6h6Dpe8qJLX3pyHR9ZHe/atCdqcB+72fzP/OInIje4tlc1xwf
DIF4NcFOekpT58sKw9rpqaGginpZGefDYc90oybqdQv/8o1vFxbxESJUISrN6lIH
l8oRryYc1xqNOE+10jvCuxk1lM5uJZJZsbHardXhoiUy9F4xKyaTpTouBs8b0dU/
s+Wei0J9BjqmE1KR6mi40/Jr/GSTh5uCZm15OeIWN6MDWqoVaEwHASXz6kv44RpC
/jNRexVHGmjkIlpIou5nH0mp5t7KqProMrc/tiGYwGIHh2giOcffqrHaSANfxUhd
MyWvhmp8BYykro/ZnepZkiGoqoV6QUc9Kx2UhQWOpl86aC651vKjIU8pQP7Vm0RA
cysrPJB2CE469OBDHYBHDFh8L1/sDn4N+vw1uJwrnlW0pGCt8aWHmB4lOBEGgLOW
0ODBqtcKon109H6nU3koc/qKkcvts1DX6FM9axc8lgcdDqsXJSjkKdqZ9HJ7hrBB
sIaFD7V0lf2c8nz34FuGr4gYCn/SMKvUShEdfH/5fLTUCqIzcTFbldRoMski75t1
RX27CSURk3ieVwZLm4fh5C0ckQBkhHaThAypv2zHzMlfMTV8r5G7fTjBm+YLOWWN
cAI8MN53PzWpiOsYNdVWsjrireHUxidBaxJNZMii39hs5DPMsce48VIUBO8THc6A
PZt8NmWl4p4PaWdTWRI/fA3R70iwZ+c1xJu2Zg97DKTlMk2BhtNPC4CMFoKTMeIb
2zDUEXXKMehy4kv79e0MDih5hFYo2bGQ54YH+HgK2KElrBUS0gFukLOtt/7Q1Dvc
jsPtHUZGmkNcAjX4h62nKHBWV6XF5pmBTGoy0QgHrbKPhRCvDaY0+2ptMTCESfA+
aUJOuDXt+xQrYDTkkJs9REqUWxkl3rG7FVHGPMUnM+mMOL8mjH8nsEvMSLrcYW4R
52yeuPrCSwmPo6lslMUF2i8/TWHTc15aeYosWTIM/1JSnBXM9Y+xPWDnHojPsR7B
1f0Q5gtoONywSj6gjmQjpfDZOD1ljlY7QBumVG7JoZbKfulVSQtCgzM+6Vg3AsKD
8o/OK9QfQ/aexKmt7FkyBOde4bGjWMiusFxAAqOuDIV06ZbHArfwyPFw83pP5Y4c
o3ia8yeDvxwOj+x5mW7j3GDLFLu2BHMUVnrTti+4kCPX869Ch5w1S2vdfV5Tdr6J
n56bDbZTvyFJgCUS9ITlBmRh/Y2oVPSJ9ehh+AqGyPsJpXTQz/jqNM7KEJpmbPV5
kimZ7UygKNSRyt3PVT2TYHUBoUP4BsWYkcHceyp/HVaDVbee9E8ftsNTNMvZZoHY
gImsZ7owJmNKFKgtCrkbMug1U3Cvjt4FMy+EAjTDahISdrdECRIPP0vBpoKpxX7S
ulLTPXh3edDPHShIISE17FOojwL1FIkMgn+TRyOJDDWOo/wI3x+v1DjKvyQ0KgHk
OEvT14WdpEb1/SGlYrU7BuN/bp2z6NXgLSEr2sUCIB0qVsu5sDVedhXaOlIL9sEr
SgtjJeC5kMoFzSYlNZFDI7s6GsTLLtAt9KVtVV7/5oaxYB+minKNxJSxrZ9Jjo5+
C1cfF1YDKTSje9G1GMe1xWXlO4fuEmaDsUaUD1AaEQlBkZVEuOfg5OPZwMtsxSDy
1ZpxTH5RGy47LAAdSdgcELb08Z6vDzTNy/g5OzbavRBtAw2HoOiTRXCO+GUgTJHU
PIW2zTIo0+0y1lbtfxN2Xzkg0KJbuwXlL9YBm540pGrvVMKfzHU17u+RVKTStk7C
q4xlNBSAzgOjcAZ4MjBpOJP3mpzLDyYCOzwXvH5wV63m7D6ud2Tlc4Wmf2Z/SXF7
5u+EiRGzvSIyjs/o9hNYQFeiaIQkd7lk3Tw/tWnmSEMWSEirADdc/3os+80SAnQL
JlQydrkkABoNZ/GoLDBp6lOBiO0Tjo9cKyVNLAq6+VJ+CTTa8JNREjFXla62xjpz
3LMUlNhKSIjp8aH7P7HUOvs64aiyrXLCIke9MDiIIAVKxL8wWE8B9zjam4JtlCAF
nWjF9JQdLA+oUs5HiKeRs1OohRFwi+0658/BfbDWpLl+zEuuaN9/kR8Re2FZLvnu
k6VxN0pOslahNbfLge9QPCIrj3Co0cNXdbRn/V2eRzUE+dVZgSXQvcg/1fso24vd
zviGuaA0tWktr9Ac9CHCOdG+2penIyz9Zm8q6BZJjT9N0tHd7z+oam1LukDMwW0o
mD5KrxvwMGMzLydTjiqsXjgxJmQNT4bXgnEuAW2D6ZA7cdSrf/tqCJBNj04Grp4R
vCOsZ+hPvgxGy8gSUDbrbxUH49fsXtwE18sh5BkIQYMqAAaFhQYCToT4aC3O7RIk
rwOn24mXK1zZIfXj7h5dFG/gwqbX768+o66WkBuQV9M24bW62+0phOqxxVM1LsHb
RTut1pAk3YLk5H/3xS7vs1A8BPVUfChB5R5vmjohqfAo6zRe3cZMruvgvNNAf8fg
uZCRpYApGUlbgJuw7OIwyYtEcRqmDlCKe4i0NRdb5mkr8zqsAfskILOKYeUTdJdA
d5zTBbDddzv7DbIEZDbuPOT6k5Y55RxebsafDVcf2I3E269TEkkxdkdE+XvAm7oE
H28vfKFrwVWhPXLyQ8cq54J+nF2H68XrSBwnhWZ2c1S/5mg7FZ29YvEF9G0uB+TR
ueRIpWIxhXY2VFBpqSGG/tqUuc2Eo8BudDlYCc/8o4VhqH+exHuZK39sDz3wbZK5
LIq9g4UMIE3TS0gMWxfTSg1Tp7EgWmglcmFjtNsaZNiiTNRlaNx0lTdb06ZtGk95
bqI5u6tjNDs9FMhACGUeB8qJ+0+86ICqH6SojLFAv9d8RtvqbGBePJeXw2mcU8Me
SCM2P5f4QzjO8AeXDaTvLRfFtSJLp0wb52Hc+9SDhmRcbBftYU7gTHlp1SPrdmm+
Rkmvzmf65SRacY3dm/0vPuKTqZF9p36BSqxzIhWTo0kv/PeaPcC41EcGUYsiEr/l
1qC5J6xX9990PFyg7pO+G8DrTMeWp7nS/SAbFFIOKKASwXeNWJNIDIdwFj12dyUL
8UspDlKJkTR2zPEUdet3upF5T7uzvIZA7QDi7JFRRnV0dXAZf9JPKlQZK7DdTfwQ
+9+p+mHq7OYlW5csCe2wO5hqIk/16mA9e/pnAcNYNfN+naPphxK1qJLpaJU3Ynr/
8aKVS7zRWI2SzOXb1nPOEU6Dv9AtaGW6Q4vLf/5QBh3gg4Tf7kpPc9Vnfqmo7rN1
ej3OBa4FCYPAw7irTI6nvYxoag5C2o6DQyvf6aWzmu9PwEkRtwlEDCBGJn0oKVtN
pDw9trD0MgXM01Iu+MjvqBhR9byRM/YfMFhvqDLTg+8hjHB9H3PcihN8zCSBeWyG
mglrORJqXh+Bi28FRFSHtKmXWGPqb0ohhYbKkcvYxaRvt21GsmLjxzmikRXDB5Ys
hiZ4iPxwGvyfrx180yRI0eDbLDH7bTvJBQTYk39du9ZBmIz8DjjM7k7yljgWrCRn
+TD1F2sZdNl4Xy/Bda1ap9UG1I8kcqflhYBi6m30Fk8dl/I8g4TzUMYoprS48WWy
6Ffv0grC/N5pcyzStGZ2il1AXHAq7GPigaF3TH8acQn3d6JDJIuLOR7xlfZExPBY
KpIGCQjAJJHWA1T1sT0N74Z06TYqTwzjePSJEH1N2LcqEtHNOX0OP+vnl9yPfGwE
BXLM/3aHfBi95R/dMH0U20io0jp7SQrl3V4pWRsPztCD/SrsKPVgWWfoc2jcJX83
qSV5cKqzaBSpgZxtmg/q9ABMEZKSNWPLOsA10uyHWGP5RpEeeVP2U89O0XrsQ1e5
9mepA1YM0WTHp/FeBJu1lXFYxYH8l3af+4vw1NTi/O0cbdyKbh11cERbnsdMhs/U
PApYUvgCR8qL0NZE2CSier58wLRN8Q0PiQU0Ko5fAbCkLfJrxNffg7/FqY6h/VvI
a9xbZAaGkuvuQ4LkAFrcUj7Nutt6+22Udlp1ltjAqF9n7PiJ+m1R3J7y+R3Wf1od
u9BNH5wbWh64n+RXqLZHa366ORO8DW1ZbWKKv+q8Gvl8e7Kd68lGBgHwLoGmsti4
N4fMIBWqS9RWbYq479wXwWokwMMSOHLWC4KO+KA02gYu4raMT5/I5weda0xiHHux
OSEaQq0SewJwApO04RM9i5G6utgAo3gGzEcojqoIQr8d8kn5abtMad6KGoeqI15h
lKIQDzVJjgY5llj4yxK5H40OqYiu0nFR2vm5oC5iqOiDOl02vba4cfSh8bxG3exj
8X5DQXGoPxDkWj5U2g/635txFovbcpeV8+XR/+7EdNrtSsbpx/ABB8Y8nVMU1xSl
xa2sE3ML8lOyV5CJ/jFLC6X4uf5YOhedetmHv4xsFfiIo5UKttGfOJ+QY+HifxOQ
wqQtFX6rydEZY5WpGaUTVUlGZWmogrNKusV+8+YOSoQ6Lg4Nz10Aa2nohFFA+1C0
fmw1mJafellZumC4i+iC/6rZJjCflaJzHp6mu7XF+PuyrEI69CovtkwrH9uL+ICR
2UDe9NmKlPT3YrnaPQzjG3l8jcEj8C4H7IYOKGPPbk8gWsS/iVzZuADHfnoKT+i8
yZ12Ou4UczgfmP8VDEBU0XgLSTNnyx7g0x2ObeJcE9stV1Tdb+qqOF24t4SMsqci
1U144dng6YEAwPL2m4SzeYnoeEMg2jqoJxpqHuXC69mbos9TYtoG3SaCjB/PuwFH
dknvHmJVoRMgUVqU+6QA6t+jbK+NC9G9MvXgaw80oLJX3DdM2nRGoWK+lA4SBCIi
S6GUaa6261zijryWtHmue4q5cDZnGPoL8f0Y8m2y4q00NT3wIXZw0RWKB1u1gzKu
p3Bb+HS1EJWQRLiReGmioaefe1+eEbpPOoFoX3EVrkbAu+N//ztnDnG8lmX6o+NK
1zTqGiMIoBdLOvoIv4Q59HJzCNQdAO0t32GxHxqkMcUh8PfiH3eIffGN00DV6/bq
SI5R+NDmoQXnqzzunRugmKIPKLWE/r24xGEXyEHmXBr34nrmMi8W2SXyxl9v0QrW
PcjqOf3/3bKCu9g1K0v5353b30n/3rQSBycJYuTtbEaEu2+wG49cWnXstJB+vLbs
q2GH4v40Vo/HDqZWFI9/vuA7lrRxchO/gOChIkyUn3s/Zw769vlcePypOAqBBKV8
EXzsenHLiphIV+eQmA8IVy7UArpmynRJ2RyLaPJx0RMeCPOnT1jONpl4QnOzhwNz
G6goK6dVpA1eqFP08zpNOCBHzqQpT16B6fV3R+EahGuNBoNEd13psr5ZRMkGu0So
/mMB6EZT96sl0z9oGORq2hQcjUb+cO1SpFDCtK/fHM3BY/R2LFRZnAQsy/WL9J1a
D/geq6SSj9PDU1BML4ETh3s/CoSvFn5hixheTWRZ0nVdNTzzB5YjpuM4b3BPj7iv
3i7lcA4/Yvw+MOwQAeU+WSY4Fmi3q5jXTAYn3eESi3GnUyuiTGqLSDEkZs7bPcs1
zpjm7QRPq5cUlYaXVZ2yxkTPLhFdofHY8FiNozzvVV/XWfslsrnukKdXRW5Rl4ry
EMCEGulxd4UjLwjLSGH1J9nI06y22rVOSHiW29KxvhwMwhch+thCb3lEt5NvQadU
B8amEDlG8LVcM9WclDExo38oESzA1cl35TJv68LDzqrzazUcokGskYxJWe6VBOFC
49UJF6avIwO6vOcCvlXUIvDETqVJHVLk+VBfF4L57X5vX6mEKUcCVSPl+gPSxHys
yLR0S5ZGDEhvWXQREfdMmyTODzCopnk3FzDocjyCQvCER5LRZZf/rx9FtrYCqqiQ
6yvfPujVmYVSaYsZktgoYNkeG71WK/mZX60Mv3D6wjPa8vIAuX5fnKSwV8Etg4vJ
GX82fwAf74bRf6sDQTKs9DUeXmLy1fATUp4hiumhWR6e66WvdzICnHaN1I/kEMtj
tDrQEJye1BB1pk6EgEvnti7QnscBXGH71tqz9O2Lbl2QikeCH+WcNTDFl/LVaGWy
FwRbCGt0quKR2FcpJB7ls4nSQD2fTepkSwjy2hE+CkS+o9h3kKJxkeHg/q+572rT
RBjAFbJxfkzBJW/uTo9tJ0zPywNh+ZxnbH/0T83/zNoaLWY9tpDVDq0RLhZ7dhLb
5R5W1MXWy02fkD8de/KY+3hJW8k5Xn87OWvEwsSzqxPeipzxhd0PCa12Y8QyfvJT
mQxCGJMVeZISYW7HoyLtHe/W6cNBrzjc98Am/6Ivtm/4VFRejaUY8WgRgDUhmZLP
HkW4vbp8fwmajJL3Wcxf4QAqZD8AcAXcLuOceibehXGI9gv+ETxau3ufT8Evtfd5
l1Jcvc/Z/ggJY84gHEwv808E91C4iIfhVj7WbRocvW1OZBBV25120uSRvJuLs5wl
E3/sRPhBKngjzsa5h6Xvkj/T4iod3YWKuwl2VDV6z0G0B8nPqjYgY4U/zh4RYIgR
ZqlaQoWGXSdq+pr8mzIhEXAHuIhZedT1UftI7G4mciiMMVmnNCZtyE6uGwtGJcr9
Dz8Wjtx9tcuVR5r1V66Dh5SBsuH4wn1zT7ybuweNYU/vyC/PqmndRr3r7cxHJUMC
aQIoMwuRHxu9C/1g/UcUgaANNiEyrGrL60jAMZBMVN7sKSU9PeUPLOtN3ejR0i6k
Jvdy+Nrs0v6WJsMZvfQ2SLE+a9xGNFSjajwDRxiicxf+WphgJzXyMdVtP3pXg112
OQYU48UJBGfMQIgSK/TbuiCR+OuH1reDf530wSeHAeS0WJz4zFBnu+2HKQhpW5nj
jxB4SU7/U3/R3eGXTeTW7Mu6lTRQjwXyWN+Q9J6pEhrYKe6YTG558W2WqPfxouhB
h3/Cc6SY64GJAsUmMNB5S6OJncrmx7gc4A/a2rhGt10naprHB/ryZPeDC3y76PeM
sLcZ3V/MAuhV6izHQKEEG4gIELyH+pIxwER5ylsc9B8+2KTJstxdxUgKtIdYYcXi
m5T1L83deC+HZ0cDniyX58fbmJkENKrWGSaFQQCeYRtS34JYcGKtAy/U98yqpdSz
GT9j1R5kw9E0LhGK1i87lJS1ZfGDMC8aCnZ8wNZusHTXzM5v0QvJ7xgmzbN+fXcA
dlutWQGAemVM0+mCHEASf6LOFLBgbWCWT64VTzZpCLv9bFo2QafLzjY6koNcgX3N
Lf6/zqQu10qCw6Nw8QtaGHemeqlpdZMR6DePmxwv3CNjofU+1KKELQq7graiZ/0r
4cJLLdGsExWXK7rqtALQQk3RDToCks2/l9Z9xrSs/hvj0L0FJY/TAjv7kxuiwWcU
pmcTQ7DN5CvkVyGGaBNFt+Uzfw8tr1d2LCypUl5etWDBj+CyziyMDKonZ3nJUA9A
Um3auXmJ0QPV2oL+lQc04yUNh8aMi+1K0FOAvt2yLVsSZLSywcPbHrnIXkkgy7Q+
a1T3sotL21kDexvSuz9ztihmRijWQHHK0xaHLY8be9svHk9MFIfQsJUiSIHx1WOP
fDzdrwJ+EHhdgFigvNZz2whFTuyDD0ye3OgOopeMODWJYF8VTCsR5lx75uty9brn
Q5eSa2JX7hAjMDkuyeWXUen0Bry+O6FRUQyoze3M8mlcYbnWJckZBLIc2qUoHU3d
lLLToyaLhXsyLFYrNscFXo2wLNj4q0YMvKUza/C4eVg4/zgor8tG5co0UM8CMLOJ
nXLoQ+V13zZh+alXOv0ghQIAE1D9DBmv9N3OoiCU3D1Q/L6TUQV6K0vQ5/B/9NDj
Iqba4wvW4lGMcQpbMrJF4yLuMxPCeakZQ1T6aE8glo+EzrIAQ3hKSi4Kmh58NbVL
Vif9xaff+hOV6hw6e4FTkz8nw9eiC4uWjNjFQxnu29oOvYwWoXb1pe8/il2/S/3L
cU6jfSjlO8tmH8WNojWtZ5+rEeuRhZf579PPZgNS0Cc102nyDVjBV6137K0NgZ0U
kLK5E35iPzT6O2qqkBuXsZmJSi09ajlR3zfe8RFHzxSq2y4twjG0a+JuWpeOjx5j
Y/ge84Zkkq92DlAQS02diWCsbVnoIjhuya2mTCsNtkwvKSn6HRTzFV6UAfEQh9hg
j7YNH5G0CpDFdYElAW63YDbrh8ZFLkhgQDSdFRV/5w0J0g20H2QoKSoBmI3w4fOT
TlOmRLvUEp7cyGEXHN1bIHLyuVzQzOIqkvtfFbI3oBpQMteutrD7jOHLycZ246ll
ZdRArMSzUazhk4UWIRV/8tNDpqS9mCScZh/k1X553eRy33Txkev0T57shvj8z2Ti
I4uCAjM1Wzl7msfUQnmas9VJbRBsuyzChBjVxQSaEuy3U7gutrLSCj4qo8mgI9OX
PcmTjqNK8E2ObCHZt6nLCAw8/es4usmoobiiiP8PQsySmUivyZo/UDRL8N6zKBCt
wM6VsqxkIsELmZPnbFbdiQT9QG/x6QnQH1YWLUxH8tjXz9sZg/D+9S+KomP/67WN
y1x6L1jSJg+Sdcysbqh8HZtgKim3FOw1PcniUPM+ElLCUqrOxYUO8omzwx/r3Gb/
Cwx19NOpzn9fm0Xkb+ii+5/0z1GNiiBqaDQR4IF/m0F/RsfPRrE90e1w4zBu0Lgz
v8knGtsY4S0zjxXaiQXA2pGiw7CLDN9NicXdMRbbtgsc/JtItaWFQzfiuE2p+ZM/
sEeHipsp3hBqbjfff+wkJYS/2LQqz5Uah5RL67PQU5m6oW3elETdqx0nMKm4cZCG
7pAkWI9OXc1y12M1FbwkbxcJdXioi5J9hex/uSORLEjRUoVwWoB3oi7nuHd9ulwj
Fy14i3+DbC9JlV8nYlUBtOW1Fy7RPxM1xclNkrEujw2zXPiLT+1fV0f33mFxd6h/
vdSsgQ8q7iLFboe34omY/V09GgN0U82qYM9k2GwHDwEWJoHNKrMzqyGYLHcG3jWE
znfbJwlq//rcgJ9/9DM9UjVnDCDbCIyafRbeg78xAl7feVn594FPuls8I2a6PoDn
oGZmiNjhWlnUv/wC3uXVOxCcFip0NqQHrhxC3NRQkv3gwf9zw73m/R7r7CGDJoHA
eNMSbXYl/fQpIduVRBPFSpUlGhSr9j8h8WtNbTKuT5GZihf6/YO3qSkGTfDlK/y/
he1HOep81OCz1SGc7boTlpj4zS1ckikSki7YRKfqu63i0YZRh8xOB4u4P9+W4eTh
irxdQyoSIcc908g1JICk/L1TZFmWFyP07RFjYTowEORPyeeeJBhYwXEg8RTOP1x0
Sp5l0O7RaiBdqh4wISjuAJGpWRE3mz8APhwH/Xpmc1spWO/LE00CP3LfHRbcL+7V
Gd1+wat68GMOX6eamzpGwpKU8pCLa69PURNd1MzAru1FySEAFSBE2GXuA/QB1Ogs
ls/zu+CIrGGZK6nKdbryfyAFAdjR6wHQEJoScgvZAdHu0U41Kwy9FaKOoWWvQLzo
oaYvTc2SAoCgjyixpVMo/LH5aWtn8l0CA03vzPIcp4mskUzWkp7fHEKHWzjH152A
AjE6bcxZkZodRZpklR+YmNlY4/pdfA0bOOLgQ5BDxRXtOnCzvo2ErPhnQhCm4aDm
g8P9kSIWona6AoK6+/LIjF3o3cdjqswOKVomPA4GmZ5bITw5wD9CyFGc6o2FQrUg
GYHwcxaBX8U/ImVVBbNuWEcpGPMCeW3TFe/e9pDXvDeVP6DmUmqi4g9UrEjzFCSJ
RfeQb/WI2XjrILMEhTYRRqFUbofpimtsKwL2kyBINkI0NunC6BxxXsfc+UbOfHGt
snL0yZhS+TFqAeYht7wof7OfM8lA9Ytf23rkUvRTCDRMqxaGuPUrgcUn95shwpXW
RvRri0C5ItuKn+5NNJlZhtVXW5rXgNZ28xOARsbsobTNVEu0gh94tZFOY1yKgFvV
gaTzVD+Lk919/SfLcXrKrzlK8tye3JMIkqwZW/8qSLU674nqb6K9WPUCKlQtoZzJ
2vQZCC9Ba+jn7WjcEF/Ql7EEav27jezBpbGY83WcS/XeOCwFvpmugwWxDNBuh4Qx
CE84oCJZX1pfGXGUHz+/paZ9w1urCdwif3FSArHZAp3lf8SYnjwPZAxrPhCKch4q
NQ7naxn62SY2tlJUcgvUrEbU3Izak4bTlZWqhX0R4JkbVpCSWMYzGMtBmIDU0by5
ax38wpgKtKURmwbu/SHHToyWdNvkunIr+o0FS1F+fHD50q3l4vhhqi8sVsb3MlMF
y7MMi82CATAR1yb5PsNd2xsynH/I6ZAjhDDCj7im4Jw11Knr1zyDzcFIljY9vJDK
zXLRtv68gvKNdyXVTBVpbnCDY9iouYxpBN3DdFJyzwmL5UnYQSkaRrFzJ2x703Z5
rbCY4N2iV3VfEQ/VOGHbkjJkdr+oVg/Krvg8KNgv44SK2TbOMqzwUhqh56+y/u9u
v4h5Z3iGKok0bmgBFyXFCq6R624LxLClC5HBRW9YJuygJC7vVJ6qbrazTn59tDs/
byh+RYhrLWGdNKJs+0Vr03rI1HCAzGwe3qvt3KangVLDX7W1RunYrVkITxNaljrk
Kvm9QARBo458RV1eVdqMpV5xLkOg3ttak0h70/D56StAMfgnVtwSDrVldQTKz/d4
RGwXCto/YkOoQZITw9bnX5My1KJrDp15rH/CUNwPOAEFBkOMiQN2YN90isTcaLyr
Tpj3cT4/UAnmhu+n7xZWKdAoOMoHsfG8IzkV/UN6sseftUxPFLe95OBU7tvttNYm
/+xMfB8I6W+O6GwHDtLuAuG7ifFlwfe8Zpc9sl+6HE4KZm1u9QGIX25ocZnROQvS
Ptw5BnNjbKriiDJvWwkRQUAiPG3glHxD6ACHHZnkA/qYN1xmY/z8Lua9vDA4kg/t
O4lna4r+tUJjnuD1o6RAyLraHjT1fnvsTPNkI8IWxGTT7bMODVfYLRPanYbTokka
VYvI0KPdivybsmwo35bcnOCIB4zzY+Tm7ST3WphlHeIoNi6BgNuMZ368ljnaGIUK
DQGuU+ECXWEEui6pM7/I/YukBCQNOKQlRAZtoVaj4iYXKRZwpYwFgHYnMiwPoBhd
xh5rGrjq6LP6KJjxVXNevqYn0tggmO3/3IKergFE5abOR5Hy/FqT3RdaAH43vUT9
EXNEk0bBFUGwEr4yCCzIbhPSvUfeU3vBXxi1EKbfFdxZHGLKeUCBJ6ZvV8vksc3t
JkAifIFw8cHh7rRCG5C76x1F0gXIQOg1BYt9syTHKKbOCCLPR+3+fmc3qMOSzqCB
pmKDLag5D63NBfA6/8JhhSS20HVAZMOecYiYcCDOhyXtMfKc1q/a2U6Vzr1pnfs9
TB3e3JFeDGdGTc/zlyefpAoKG2qSciRO7aOfsHD//6UbLjNm5bV1zzxwvXjIvqR5
jZh99o51VobGhepD4yyW9CxE9z0jfRdnSbxSHKrbOHZnqLuxAK4xIMXkx8BbcNzX
cwkCCvPkJ8GnA6T2UfXNoWPQiGpVq+QeEmIxyoO+qD6rBFV3Quq3cIGT6PlbKmmB
26cIYTv7cPHqfOcPNrxJKf0TF+guORE6t4FTq+QmyzVRt5+UXzu2IaFlzcerlXd0
XpPp/AGPFNyHOPbfqaE7qRSXW+nw39dUyZwWXzEA9KiQ2S5O/0OiMZqwfh3st/xV
i3UXz1/g2jy/MHfzw2usQd3mQdZC/OY0zV3Pqli59TpYpSfb5J+BtZxCO5j6I8tM
TEfKMFBU3gePcbChMaNKv//DJ1AyrjkhPlhs79rfHtl71VhIpA8SX03EwbdkRjPK
bqRRtwauAnQmUJbHQ+4/oX9Za9Dzs2TG2I2YB7Nem4HMcDVnV3sjScWQfqKL5jYN
ETQfstI6sgS6drxqUakywvIBCPkpUcrXd1Jo5qqeGlrLooHUp1hQLIOZ1rhT5q7V
4BJ4kB7YocFXmsgKj1TOTVYGWfJ7d1dIli5tnfSjKXEmXAzpPealNRPOYvdbDq6W
4ulddOm1bCQDY39rUfYIXz5PHt76aJsZSVuqv+T5lc68Y9ozKlI8F8SS+/gx6EeW
MEDA8z81X46ANnIN4vymZB8Sm/iukHIxaaBiFofMrmdmza+G7nUPTXP7rSFSKfga
E/iJxrEmwrfFr/DYgkHe/S5ULZjKnELx4f9vdFTtDvj8dknoVfHvPX44u9VpFvCu
TH3ZsCjQstSJsTDULQAJ4kTwOwkbCNDgb/vY/SNaYl1hn6tYu/GYgCIgpwoaHcXH
1/ECChKcrVAxMsvYCWhW2JK8gWeHOwa5n7/5RtAzl8xpIwas7IvhixSlhQ9RhaPj
UcVeUAGnC8agq9bQIxsgm0g6sYLDYlRyTtP4cv7WRyQ5FSdDz/fu0BAAkNNMG5vB
tUaIVJH1ErrMUjVegy5kIgQGq5/m8a81PyZJe4X8ss26V1aNJON/8Ln3xmSeHXg7
4ddGj/Hzhj9u0RHSxnkzkle/yavWlbVkk0fy06wiNhlHC8s5TL3fNFKbEYBnZRtw
JQlO9fm5fui3NLUxKCjOtS+03HLgSYa+Bwhg342JuW6GSiGbiCldSKLGl4pZptBJ
wD1o+om9G/asyGs2kDz07/91B4Uo+aN23FR9VdLO/yAUPVAJe+DNlaeA+dGZWyLk
frKxlq8PhHZj84AyGFQ84VWvUhr6AO/IT7hnnJfLXNDY3ofjDgF4kIC+YOEBmBp3
wkTPeAjscP7J27Pvxt/toEjAbvpZyNn99qPpPQ36dLRGLdFF+CUKDPJc/tXLdgrj
fhgT/DlXapi75RI5eyvwTXAjTV3rjv7YYaeRh8oCG5TV//gDvBSp+IhPP53sChYq
RMs7771IxTn55ZGm36VOtkdd7Ctxc7AQMoHedtFsO8oEMVJwi+3YobiPfXa5zCS3
tV4cvACubJ+44LISUBslGSOPRNGovHf3D+RlGXhzO5k4IDG14FbqVTfHVep9Pcaz
MyhjuCdXH15C5ib0Dpm8J1Kmlg9JckP0SHuJCxdkGPpcdJRXxqqFqJvNNCBjDqvK
wdWkb6mXew+mRv8IoqfQHJcSvKn1nDESQStmWZvq0S3h+KK5q22MTXfoWPIWp9QN
VgkBpIy4L03D5tl0zRoWJ8LlTY1lpS6VLeWfhjKjP3/f5DbUnFB6iwr9FUb8jG+w
6yM00aoD142NVozQ61EiOg6YaklU23seQ8EIMgdj8rIcRU7R1NcHttr396qT/78p
GuSuHEHG5fsD79aKvLd6lNa86W/UAgic/ilYwz197GbBilc3ADdWLaXAmeUuMCI3
PVm6KJpLoQRHAu3EvGSMHih1YhA6PbgcA4ieJVu/By3vo2Vjf4r28E4A9neuHmtC
cVLBJExqAuDd6l7jRnew2OWSTt6dgpTIY00ZY6zF5o9KCrEUHcDu55QdGSh6ws7F
UaA8+AQHazKghCdxXirOXvOetCmWXAF410BL1SjTCquGjUAEyhUWdWRMev0xIuGj
+tAsYGpeKhbwDOUIiG19RyPPfp16+EI9fsF4UBy9Qj+j+I6SjIWN8xHq9rKJ+Y+9
tv2+7FKkvoMbnYjGLEpwDOHVpDDHDfjhRdikLkbEGPqLK2y7SB0KzHvugz8u9aB8
I/S/WpjmJaQAq3r0EdmcE24dOf49gA7XCgmRDMOsHsiF0bff1It664pz4yk73tpB
uKCI5UFWos/NrancJCCUIK4UeW40/wYv2t/GNRBx6cq7mqBICmMGm/2IhNbuaPhD
EBmg7b7aXBqIBU0rNqSY01451hKJNK7k/UFksG3R14anbl63HQXkH09DmfcgYWuw
4YxKoJF6UghQ6wXewh9IdC8ZYcHzesiBfmhjOlYl7A1mc8xiAjRtC8Psew95OaQq
wZEVO/HgGLXw09uj8pyU4CJ3MbOhctLqcbQZQJaybrJxh4bP2xjdv6LmElXrISfe
UH3lTv/c7WAQV9G5q5c6xfkwhfUtLG2WnVtxNW5ygyVMhQX1FUuwKlovCEDVAQu4
DaK0KpNuGZHChGkOijjDc+GPq4Pw4eVyZ+2+REL0udb7ybo9CRs0SpzPLT753Y3U
Mj+c/E7VItwXETCdlUQFVRqB2/e2P4BmaI+4OBaYpkOlDoWAVFVVgnGE9d9I8WR7
geLdIwD7p1Wog72xBGyOTWH72UYIzO2KsVbhSQAxFrXOmu2cD1P5ycaKQNlOqT3j
csHAatIvXNqDjKL5W3f3n5ANOmUlshwbuEDAbkVhniilWHMGHNd3t6YBgUUhuLQ5
OSr/VeK8eDK8wPb5TZ/pKVOrKDhZOH3B5O+FHdjEIB2+rYTWfta5MpfdI6xtgp7y
xU8zdTyfjtTjK1LQQwMMA7JTxYHbJ8COlbr/yDK6KW8NhBl+aH5p5TA13YbtKLBT
JOu+AGz9/JIu3AWHe/c9vOf28Z6Q3YP3u30ZQk4YP+3syP0b2Z/EPaT53gUOM/hf
9bLaP9zedXAaBq8ucgDYy+QEFPOH8ghThSERCWzk+UQ43PeJvZMntcEFvHBjMppm
s7ttQKgav1sciN2DwDIlg4rxzVA16ISyx6T7OdVL9H2BCTv3ySJhPX7e682NQCW4
gSK5/daDD8I85+YOi0nlA1zXCHt7N8OpX/foRwnH2nu0gonRnPybDQz5IpbuBGzt
OeZyhpVsMt0yO6bZA4SJNBUfGuRIqbeCcn31HG6yLl1DWoPsLUZ9EO2Ohv4/6OoH
CIRCcexPVP6aU6y7IGdrarCR7ngMqIneLxinkhlaWW6aUu4pk2Pzddoz4pj2zJ6j
YiNB+R1CdkEEaNJJNEjOM20ZuaBhq3kK7xY1XnHVbTlZmk4OLJdy29oMupTryGUs
KrbkmBc5JJeZPWq8bMFKJITgT6YXfJ0D9EDd1BI3PzbtlDWQe9xe3jUp0sJY4AK5
6KR+HolCBPRnkkJtoPsVlNwvcX7ghaTxaq8bDgXQ6wIjELv4lyPVYjeYpT5nR2LI
l9+CO4U6iXuUiYTj7n4rbyb9t91GI4ZqvigtvSsEmZQf/QpAp8CjBAMCdX9sCxl2
w1vuHAx2GJ8ef00e4BdKhAlotb4MqkQOtGdUrcvt3BTBWG9+C4l16BYtx1FjgZ3t
AoIXqmk5sp1HXkhjjmzQkBg9IkN4x38lW9Kr/S+cyeCRWhNJv1YFmzA3IElPC+lc
4Ewh4oXih+aXisl6UtmyQONZpZkJ1jndjr7cGxhTaq3dqCpJ5PiC3d7ko1YmkQSC
zgyv2wWmSKY/QYhr6/a2hevNT1ernPR3rDBXJgTfmySSiLp3oL+dL2YtaaWmlylB
Pgf4pRAH/zB8K7SOoKSQNMP/kOSMl8zqNCooV31K9aGs5r84iW4N72TYnjwnHi5l
PtRVC4rWAofdIcagT7xDax0UOSBlDOxiserv1TVUgiAZCsuWg0Cp2NXqu3TWQAYl
doA5KuLnvxkG7LKgfWeywC7SEMBNrN/XbJOXuWw15X7Pasu/wpkqg3B+ozA/vX4E
EjFNE/YSxQOCmuAWaJQKAnVInu2wfAhYuEBtvVRjczUh9uQxDh09vFyfGH2m+Fbj
7CP+o3JFy73IoJ+dMst7WpVTH0sriWSD9tWxp3moZcAvFSRYumQXFOR76vLBVAHH
zdu5k2XOB9Ez7RN89r5PTcYZK3q+2MwLq4ZIHkuccoKWjyBbg1Lbxiz3DAmKuhuV
+beK4t6GJfIyvQgXvn72oVrvTZfQO22on7wjwlmWFDZMLsG8j+Zpx06Kk0qI+CI8
aFa67XtvsT1+eebfzJXQ5AvEoNzDxvwguSHrC/xdxDogwJNZmXF86s7jKWgMiJDo
h4BzywHClnnnx6auNuiFu4C67kk+J4mwvECz56PeQxDIi6Uhj84FLQSH/OKLYHJs
cWquYnAvtgCEYH5oc3YSr3gaD52TP0xlTFZ48ZZKPILdAOhFlbG27QV4l6OmWrhS
c27LpngOf7ThGFH/Qm/+EOhzomFEu5tREZckfQuDY96dgmPg87TaYxeeVoVb8he6
WTplWF/Lqt0orhpCtMRy5+i/MPtxQl29LPxSIsvxOr5SR9bxwo72ACUgIgFGd/Dt
9hGrQr5lUnyWUAuHb7mLAgEivUtMLpLU4dFvCHWAaeiYhII2gg7UTudGyQUPxzcC
RnDRjvUTADU2SR9uA6e0ZLuEFBz7GTkULLfnTml4sfk4213b0NB47wGTnYkCtV8f
5kK5MF/CfA7MNw+yHOMt6PItbPefTRQG9Uv4rzCG4RZ8wlrXyJfsZhiPThruhws8
l4NrjVyyEqxxGoDAlkVUysDeFvC2Pp7cuhbhatb4FE2Vr5sYzvqZuc5wo3chwW0f
lBHdbMmLP5etIZu9gPWgeCBB25Y7ggpGzlQAO73/W0SZgHhqpFpSbpn6V07ejasq
YJk0D1RV9Kp3jFslIN0bNg11dhZCCj5XLOcjC5eBMe73b/jZbGgBW0x6dLhywrX/
thUz8GxeVtSKz4Jr62AapHd5+DwZgcpBxsGSiNFeHpq/+7nvZbjszbA3lHqvx4cj
zkLRyyKpr70MGH1B+4huFgJZSKXW6RSjfPqKUJji+VLAy4+kVUMRewTOKRXUWUeH
Fi7zUB9ql6O02PUPxBx4cyZKejFJ9WLyoDsR85JThq/WxT9YP2/P4q15WLPmABt7
SkxnwnlSCxSlX0gtHvP8Qtdzwl8B4ktHY8NdBjNA/8q9im+CN5YTG5ved4CrWJcA
1f+k7frRb4JikOJsY9mWSv8CnkoI6OHFyI4AxIfgla/ktMjKFuVTnRPR0vl+K0IN
wjxSdKhzln1CTGsamBRMkNtSDNfPKHXox4+Zjds7apl5XRTan/WMniw70CXiJXfa
4cpKUdcqNA339ZFxbawSH2mGcfDfhR0m6dN5x2UcqbUvMqadcOohVgkVHXOtKumb
fzbqQYk5rOLkieoIVzyHvit8oC0B+pWSqm71Y/d5W0QZoc2bceUS8JidcB79rqqo
WDJpSrZaVSu5cYUde7zN2wYR3x0BAod36r6Hq+P+0dEZfAIdMLaVhHCpXV+TWj/3
Zz3kR5msV/51yfzEM5FdhfYAKeP0ZSAFqNAn2pfXcekScmZpp68jpZInjSO6zgAk
LvQwev65UcHFEdNgq0/JaTcUWfwSWcnf0EhFC/e+Qe87pLFkidve917n/YX0T0TA
3UKOaa4GH333HHJgbhXvwRoPiBKhy91BqFJtQ+hISEnV3iKaMOjDVsKba6CfV43/
WFHdwzbl8/stHFNsJOgxvFT6EJXqYcu1x3ppxbP3jOR0Md0C7EIuKWeOLkm24c7V
HQKTornhhzSYzfnYWr3iwbMG80j380LrK8qIoghbkGt7s2YK2Z6uDrMm20Cl0MZf
QjdcOGx3dPajlED1TgW4AV81Hdd0JfJPiApt2otftQL2Zr38BH2ygYqu16Sglj+w
D/tPfCgXSEzkvdiujzymfWx8u6D126INPvjAe9uYP8N+jfNcY+W7T/i8ZG+KJb60
0SyikqIPG+/xPRqdcEuJshJeIM5KWbS6fqpZ+HuzVU2nFkYtnJAXYrTaGTw4VIhO
1v1RZdIGZKqSMspXmuHH8q0ebtQLUtAIfRGL6gvmn0GwA2Becs2AHoozhqgIrr8s
JMdU4jawsqaCfA2sjSZ1LlAhVE9uXQz37aLL3OLhWehdNsa63uHpWhqOeG2TzGlu
DIquQNQRTzKbtB+TvDdK/lJQmwULEMe3vyGLR/il+Ur/05mM6l2zuq5Wgivj2DlO
XtanG4heqB2hmM1W+GcBeVtq98Yi4CAp7WC9t5uHYpyd+oxGOHFDMwaGYesPpOmb
K0d3rrRVRvoMKecLx1kOPz9sByF5oChWk5Ttmz6xn/+KuDbeChCbnb6+v5NTSvSu
eWkleLSEepsacaQHA0r+zLePxOyLwDgkprGXUq/Cn1DzmXCObUsSo30PBNiEkF5Q
ioeUQEP9XR4dG2PGGNTnFgM7ZCgzzjXXYWHYfDF2CmCNmE15izILYG4ds2SLod0W
5Xst1+qTFoaDYLB1TiOyYwFu7UNF2PuOy+XCVqmLVVFWN26h/Fb+nm0M3668KUg/
85R64/amGI2aLre7aWQt8ajPPDR7urAPlV/qpGo/VZr/EXNsWO1XjYGev3vZFOe+
VXbFXjxZ/nlw1hN/jq5MmQKmJJKW1vspzBOeWHce7iPDKiXwPg8vha+3hiV3hDIw
VPQ7pnhpEQLcVFejnSzW3205sWXXOCLs6FAHb+B+0JSK1SxvP2ELdwez9pC8g5Ct
Kdk/DN9F0h1cZ1eLaaIpBQIap28ug86NHydL7dxuhIB+X96b1lw+tW0ZuIpHOEdJ
6S7hkI4DEdpxNWh5xUV7jC1sJ9o7e8y/YbGtFdHb9y1w77gC0kEdG2ESiWAA86K5
pdhUdI5vZPiW/AJdw13p5Y0Nvl6wxleLuQFeh4y4FvMIoA0efFdYqzYNAKcVr0Nb
61zVorT0FwkHR5+EK/gxFUDgLMtU7cuKaDNFGqQnb3StbBV6a1PDEb4QLiXXnXBW
wfQ38cB6kl8FHqhg5MNc7NN+YxfWsEgqjJi3Kp/nAFCpynJ3lNAI53s+xuoxceDA
biWBBFURqKlT/lNOQ9L2v2wtOVeKxfMmWla+au3Tv6xzympqOsy5uOQgUEI5k42Q
yiZ3/hj5gbm8KLgdes1IxEbxh+PD2ymIz9fSIuIvRLhmDS2sNGfWP9Q+9psKwY8O
mKZB+Qmq3SU3lMLAyAKsEOw+l2NKZOfC4lGTQ0f5QgammPYBThn0Q4g0M+q6O8WW
din7+9TESKEzhN7ATfLeBJxu95Hq9wBbrCkReKVYLh1811Ig9CqO5knCtQwpILMx
PRaUb/zEGJTvy00QKNnrsA6VuJ0sJhNDokqmq7y+KNt55pkjfR9eftRWOflDOWhy
Ig47FRNYvNyuUdBUii02/LR8GrmOAewj+4RPV1oQVj82B4MmqU13aSWE3jOw1LAl
zqbg7B1C8fPhVhue+wzjP1+69JhS+WYJ+HZB7cvPSSbGrWBjNVcwTZD/38TVRosf
p9eGQ2jUiIhoEtcovvTIIe3EDLLVnbp1ezgAvLlRluBXT0yBPwHIFsjjRL0CBkXc
9rYKVKWefIBHR9nuWL1RrCpbpXpYYGevKWo+dN6fVTTLblGtWs+BGjNHPifiCyaV
xw8RnlSfhgL3DdSi5byJAnosK8cuOuVmFFQKG3UnYyW+qYCcVjJoOjS5CzEyQWBi
7gXFNeDwDS6WpoF3CBolmbKl1/hncUqZf7Vsyl8FRMXGO3Rz80vT/DPEeM17cDFy
C6kfr3BmkpdXWDD7jfz3LTjHGOXOnu3omY6giOjwfWJ2+5TCR0fDjoz/m27GtVz0
oRpDRi8arKQmILzCza1iVa6QuJswwr2rDm6OOf+4rrjlzIXtqxAJ/TdwCEEYJzTs
Rk79VuEGLwvM1WHOKWB0VkdZJCOIpMI0aOWt5pjSImkRihLhfkbOyurd+XBDYFPi
QRKczDZGsO+dmGxHLW5+IoC+A/ssmn6fZzc2R+i2ehyPViQ9nFcWxSfadSzH50G2
JgnIQO27wKm58N5y3PpBpDhVCgg/iXdezpRgJsipUzVWqOtSnaurtFqR6Adx7woy
uEH9iLdkE3v50t++vkSZYa3MhMBameGJkB0XYgiiA95Yh3d2sMRLJfLX8wYRKgTH
VcosMwgFXhtkZ8QwjsIAFOffIAZW9ftgbbTqW6sg9jukQYIO/5r4BVg06/7sVpUr
u4w6d6TtXb5KiCbC5wk2l2GLIW/3Qz7f46r5pyxSE9NlAdq3ZH+ztwyqDzC4uzfh
/5CWJ9Xlewt0UWQRFJa6XPmpKgZ8x+41xe5gpzf40mjBPR0cvf0DBHV5R6iq1SaO
nPTHZ1v4dQKwIPCHs9ZMCncX4djsEr+bdzWC+0h5a7xuf5855rhbEJYEOOl1aPZ+
r2h3X4Su+X0yjDcDZqux2dLMkxAG2nFrJyHk+Oc+lYoS1bLLEHfYaWxPXsP8UY5l
y4XfxNMansSYtvXvIKLxvrlrHAs0zSgwxxY3xsJK/g1K/jk6PAOb4GSKS7BnX6kq
m7/iylJOaIoJqzfvgrXXDQDZ41F+gatKZfvwc0Ejv7LNCsPplHtTsQT9rysjX7pg
ugOiKIGMIsReR49kP2ncfBL4H9jhX0T6P7Fc3YEqT8OwxoLXFjXwKKeQzYiWZxBo
6hYmQHU0m43PGrFwLg0Zlb6ZFxOWyCONK60CPRwo521esbJ+OysGRyjjnq1FbHIk
NXsmLWLoLKkGrHrOaWXa1YSSF8SoOKlLw3qGcwPnv27f3APXjzDKDRsVnN53b4EK
w2TqhKIV6+5OTMsEA8taq2SDb8ROfoHX8OjTf6ldivck7+uQFj+8NPBPY/qHPIgc
/pc4DNHZoemDoaFrDfdGbgZ/pbkuMPwOr0YW3P0K7YURp08zEguATp32fYUeiLJ3
A5W+nE1QA57dhaCNW1ytZBghPIneE5oYX/K3QLaXA9mW9nEBl9QAPJP/QwWWCElt
G4YEkUv5t0KI0ZnSNU/vyLAI8h0m6OvtkpBwOcjnnOa8iMfV+2pgEolcScOxJ0Ur
25DxCkxN1noXSOXgNHoNCGVlXSwc37hF8TZY+MzFOUnGTMBXKKs24n092CYN60Mw
h3IYC4cBRnsTHVSTs0apiWSHecJY5lmNF0FN/s8LhXogchWsV264xiyUSQGIePHj
c+VY1wahcy4x47SNh5GPNFw2jnVsxLzVzDAem2gaPrCUEdJyeqJ7MXOgTbwUzebn
i2QETGPyGMC6RHYsjPxyNk1JLT0E1+IxtdYs001RKWb7PPPA9mHtJG5+/IEpMi3f
evHVgLiD//OdYjeAHGJPUa1sRRS76E6dQsSWUSkE/za3T0cu6LaILuVawx0p8TCc
W/MD4btFzoglMZ+cW7CbQ+VZOt39gasLPCHdlvNxtbRMAHeLYvU7LxBwjC2Qk4xT
k6JviAkOON3PFxG9R0dklwzgeH8bqFQrMsufOlTPKz1kpaATbXZX90Zxbe0synK0
yS9XAtgcZgDTFtKc24W713h3h65LuQJA0yzgZ0CTbdDTYqk+975XxVDRZ+IMlzjk
O516TDku1sixKl2tlZ/48NmJ+CLKw6xCIlzFaqkl3jei/suXxXFTsJNbQT7uGOdy
+1L9ruAAsyYKQa0d/i82iug/gIrNpcDGbNYDTpKA06rzsNDeZYornP88EcWHoZfd
NenIxyA5nrknYsATijzzkzVciGJshfIRWjYqnb+XTJnvbgOLgPqsvDfPv0VizUMj
NGpt1/SroAgs051KcHDbK2xWB7XQwpwM8WPc6a0eLT7YChYOPMGoe6v3kSs3ZE0y
IushIRAbVACG+UbHBvwnMi99VfItpl1LK4KY0RX2KLy6rFsOiihGVg69X8CAohyx
h1YXx1q+OMG3jbtK2XKKQBFc13fAqRGEp9K1vXZ0b06hG2UM0SAdvj64n6kSpHBh
xXpT+fUibUIZnuxN9KnvSdxjXpIPrE/D/DrupvtKFgKaGleipIEnsrnJjZJ4KzLe
WbqzB0fPhRU7Ob1vwPRcqRwImzvjbGY/iIXVAp10zdKhorQdXXpIUQvnlhuWx3Kg
CuRV1BmfRmF/Hsn5KfZB3Xo1kWXqx2Mdk+DCNDcg2YT5K+ZO3tIen8kZ0iSiPtQM
ksuFjzQVAcsbAab5lUiLnWzF7TZOvnkQk0odyD3nwCzlbE6iSUOdyxZmoESDKOWO
knfd4e09lgsGf8lqpKWBaVxs+qZE8AAzm+Wt/UQFosEt+LBpdfjXY02fhAAmkqam
dOK1HzipdlJYtn02Q4x6eJiDaSdbQqbRIJ5olI5WTL+hj37CMVvlhZ0i8GtRUBV2
qltcR3HJIbxZwGQOcQJgVDxDgESQ9/SMUgAqMQwgjTTBIrSrYdJk5Qtt2mxMUv9X
vtG9i2rwvAUFDIk5YmzqAJpPPQz1YJT1QM8cIA4q0EXuNeCpK8t+JLimZmql6KKB
CoOdHZZ1UZUIRPY3fcIBE4teCCb2iSh1veEZmJHSpenRwIydrqO7d+YCgN1oyRsQ
uqlukDLhWH7d9yph06rea9U9NuqSjDC391CSZxzRf5bbAxkkI2M/kU3VCPmzSkhq
bO7hjCXoa+TtuA49kMTtMsCn8coCIWz0/PXfi63vkUbl/3ecJmF76ttnrqeOHDn+
JfPbCJxX9agg7E5l+/WKAbUZJM12j9g4TwqWE1XYQmpV2erZl4MT5y0MQdy2uTm2
h51LnTN3KOpCFX+46mVI+iwb9BkoDrfXDiwu49/9IjJ6hfFQ3OppsYoLpHEdRhDz
ncHQv9PLOvFWRil5rjd4suP78nuxvZpyGvdU4JJe79FTJm2N9B7BRwI9AfO6Bmna
VHs6H4AhA5KGthfqMxkkwLtgM+SRb/HIaytyXqyawJZTRg1i2IRMQKx5TRs90WGl
5NqcCbjOSB2nhyhoFAZ6QodGsj7heDDMYyMtgBvJCjy9WSi+jQ0/8r6qnBAIQl6X
ulTFB3KhCDTKkgxT/Zwa3tcR7/2UuQvg3uqK7Ph/iEz3f79lFO5WUifB+FOjWScP
XVeIYzx3EgaLi0kIyX8OaM7OyAtvZoNtT4pl/yzbq1coB8PTc5wKKHhI4rJRrtHs
jnryz0472nlKSFItGCsaY+htJZd5b44nhRTsvLG8FnIzcihoTMSXj5SpeUkBblM5
RCXAvo6WZmj/XhPFuG3UVCysWra3qWLqo748i2zlY98CdtJAoLHIqSmvL7PLytPo
yHjw7+4v8NMfLhuVuHj3UnHGlr75w/vBxgNXUVsDmHVIQduwzYARE++lRyhpoWEq
i5W4fbbGjE+yYFMl9jZ0Kl0chMT3HmC1mtsnxSOrXuDzIWtLuIS7fG4dNXKPtptq
YsLGIoFAlbj4mFvbsE5Kc0ejPxRDJo+oW2odg5zOseQ7UPg9X/JbmuG7kdJZ4p03
zSgBAoCvLSs6ok3/6qUqCi8fh90gLtUalnQ6W0LPq1mgIzs9m6CtGOAYaiSgQxWJ
aoVMTX4CywUUzDoi6WuID5w/Xx6IvSvtQAOFY0GzEk7hQksOhXRN5RoqmkwqThTD
pmZUK44rICaRjibMBY852hXKmKYQGp9Baf1gwcDY9MgKLpHFWC4bd0C55sOQ75K9
KR71j86UjJ2tM35roJhjiitEa5x4NlbUsI20ZN9ygNM3anpEqPylYol+Ko9jUhnb
IB4rbOXh4TmguE9XTOwfp584+6Ni3bBUTKiI0hsRS2p8iN0cXs3lUoPflxlyh3q6
z8pgoIsQNIlI1XM5sAsalLbk2f+H37FptjS5crCCJo8IdVIvJJIepUaW7NkZUcdB
5ScGLquusvf1fA7v7IPoDFUgQQE8O/GEyK0mPxJLtKCLLlnXMnV8djeeuJZbDQti
e0Ytr5+AOgNZF8z1ELxKe1Rau9SCIQn1Od9GkG1Fsy0VhLlac9FD9WO0YPjTVw/P
fZsR9HzX750aLkp27zSCahoPSW19S8eJUdnbSkH2xvmX2nbuzxpJo6sL4yEVSNWt
WuVrhG0Ib/rX3eU3e28IIb/7UHQtTgrIiipWTGMtud/S5euIjtn8BrK6q5ogRDIB
TpVhFUN6l0JmqQTFQvcu9XP6+hocHFaLUYb08N4LC9a2jqXSs3i6i+rrtYqsg6br
XqQid6rC6XlRo7h7nRa82RE+1ZDGIafVXn6NGm/UFK0BkTDPmz4VNwWvBzDGvv9o
DFMHjN0YV+UV0eu3WLKPgy7BCppTdNnZzq1V/BcOdlkaveBNNUZZah7lIo+Fm3GO
hcov6gCcrOuWH0wPNQC4HQouMtRpUnfXkNYuZQPVYZFmLc4ASmucX5NLNH6ogmz8
d0Arn966qW6V3UnmblYGijMbu6AgPzP9sohitsB0MntQcW7xRCxdZ4PVBJ4E+dVc
hdswpoROFhSLsDMdQkBcP/Hf/GIWWHkRmNlqaddzX74mHsCsf6ckWJ3pVI0iKlDa
f+j32NTkJes6740BFISYU2+PfikZOoWGPQkKMWbpl5tIPpJ4CwivmfRhqTX0xFed
hecAX9Z8c/TMrqz79Bu3oT+m/pqQDWxVccQM7w0Ydq9HVUCb4F/+1wkxwwmo0R8s
D3deWjyCmwkjIzaslt98+4o//Bf78EnNJdyvxVzDAax0hdyY43j5dG8S0Yz2Xbrp
DSJzI6GYM+jlJfCeAJj1rPBFHP8CZghCkwnm3nLaHsIzNkpEMt5pNYGGr0VCltlI
2yG2VCNgKfwXNJoS+2chFosYsoajmtT7KMkQS9a2pnY6A1tYzVugul9yi+/9BXcq
eEzLHckHomaQbPvX8ztKdBwcFG4dG32nx3P9lLz6JFveruqOZj6BJUAVTRigsikA
zEHi9iNElSo6NEI26kahx3VV5t6b7ItnfsDd/6CL3sIIhxRKsVICFsmmwEMfi6b0
ETCDSSNp8WkdcmeqkmU5hL/fMdoKIjXfwJcKLpmIGiezBuP7jPzMeDFhlflIK1Rr
Xvm+HcqawQ4vRmh5poVuxGtq4mUtTQBNXInPEUTvxSsSnJTTA5hBNpSmsVm3Q+x1
qu2h5P13Dd57beybK3o0cwD7k00GdtOiwxhV9CwzwR59nqqM0kPKT3D2PrumgaKt
x3KMKHa7L5wBSauh8bxKOU+smR1rM72xGeDXdWQOaoQkO1L3YdKIS/S1ddNcvTAT
1Y43LQxwoaMCB6mX4g8+OnRZn1uzH7DDehcmTOOlv8Cya9AtszelvwDa7XVSp3J0
pOC3hIAWGIjfA9AfIxLUvtl7Z5Y5e6VGVoYZW8YDxSEGcyHoAUwCGeh3o8ppxGWj
2AiEMEVzr0f8qGzn/Y9rgZTi5rbikgPleRILZoqLUFxjfe0JRsrDJzWEPjFDXv3v
35e+Cc2nVVt35ks5UojNQbLIO6rAb157HrVo8Lv6EQaYVKddBxXqQ9Ek8mhLoJEU
tXyUlQOTzBTN6aBMQRweWwYeN/01EnLPTKKjlfTRHWY/j/LhXnPXOIeD7ZCW1Kxn
pAoAOdslJnzN/KWTrgiRTDMDhW4ZCM6uBxKwslT0VS7zQI8b4Lxu/GAOsoKz8Rk+
w16ZFcDHrNzvyin8D/wiAl5TwATa9inhBNidO1GdhkF19LZC5Wb3eJMedbEAVe8j
trRyVlkwgH7ooi2hwq/2Q+vCMo8w1MuYTZB2Tyrl4U2jaPzvUEEnBbAWO+OKrrDb
O4E+9qMxLEvkWjn5OqxARhhxcAqsS4FsHmqquUGEP3xd60d/hpIS+eL1a9CAHyvc
6RTahlaNZ0KFkXjaBEaVAk9aGsYZArVPyBySGnjNGi6QgjDIjIe3eYa5COopY7Ma
dhDXrv72OvDHBpPRjCoFrZ0fRYiw9bftDdjWawOBJWY8Muh3eWbVoJft4xrbIsm7
U38YEL0V33T74lQHmOsPli2SsDFTyXiJkjkKGm0PLOWoPlNL5lpl6hqQExg2GUF2
SDWpKbMqBdYRBTDKq3lJkc0zgUt/gRVX7qlu6Sc0rH0Lfi/OhfhR95ZjBMblXb+C
SbHzKsWIpy7HjDvsn9gat020kB4nR10i4S+0HsQZPbkKrXxxVBqHcsCgZtul+mqt
UV3uunfs2zHeuBLgwtFLHe5dQ2TPJ8kVrQd07h8xoBdXS4QTKovS87kR4Eu6NIsP
ZzXqS18FsSBhekLvkKzHBx3XIRbp5ct9hairOjK5qos051nyoZLpYxzHap+amgUq
yXDCA9CWchqH0n14N46xClUqYGryI0OLYYFAkmA3itBiks0wY6z1sutGNXsdjhu5
FZ6k2UhIh3ZepWluGge0SyR6tJ8TnBpw5rOnhCk35iX40Tmh+8E8uvfSgvyhV0pu
fqB47lHH+3gtc19bnFMomRQGa0H56TkkdEaXxtGp9E72gEWBuzSaUNDqqWeVbbLS
tFl2RutahnHsptrcTlDgnrBwoIACPytA/VjxSa+EuyOH5ZXDsfzdBC3UAswIBto+
c60+FoIcpHYM65fBpRbjFywlpyK0eNE7dCmia2DGhPlGgE2ceDL+fAe0rKeOR7Wa
WBG1l3Af5dcnp/N5xeMccsjYXZyBktpeew2l6a+HlrrJgAxWyqntBuqaPZiTX2Bd
O0wd1z4jmO9UY0EMQZdER6b88iuYsRxgIoAQQPNzkdICjR9RliPie7OQmP1SKG97
TfRjzACadbF+g+G2WI00CTA/4h9pazc3vmJOsaRrBOOesyRwx4GV7WebRvjY4OEy
At9Jk+P7DTHSFstbC0cSLdXORiaOlk6azcNUw7GONlNPaffePtA/i86wFEWo1hBY
Psefwp9fXkN2HancOxN/gh/HHFEY5VA1aCtdpcsISIiExietR9sAp5cBAd7cMSxC
WZuveaJf+pGHlH9Vg4YeOWZzNdDuCJoJEhj99TGuqdM5C4MzFR9IQOD/CPxumM3m
/eTRFA85ESrbO8l0NDDHBvD77wh+oyIckBEVqGFdqTDkZnjwYxGpQpaum9pTVOTh
s9Mnx1tcmjSWiWdy3NStjlwQFblQDnFJdWJRoDJyCcQG4Cg6g+ypyG2rKOtanNSd
hR7dNGhVAuCqaVCMWWHokE8fye+xxdc52PsqYl3Xq1iqIQ6rwOguzxZCPF29QfrD
iYJ2SxC07YNY6rHBMc2hthePiptOgphzzT7uERvXj1ugAIwtwGbp+bFHa8r3G3eY
nNm3ElAi00nwtkFltLJutCW1EHzN8D9ER0jmmR9FF3BvwGxE4GMqXRHdzZKEbiWj
jAaar2EilJSKl/xJr+v6ne5F5EOBKb/vwk7LSt4GyRzg8sUu7S48r9b+vgstuma3
D/SFEKUuUJxmMuN0knx3vqT62EiNQfOlKOXHgH3woT3HJzOIVZar0nvdua5RCWoy
XIea+w6QiDgpZ/VNCppna5flnL0vu7EivM5+IMmVPE0nhp+MEyExvJUWHO7qqgFj
U343ipKVYX+LOPEO/a8wPn9uatu5J5KHEvuPiM9dzm0voy/3Cp17NIBsvd8C75ky
xhYvrbCWWNgVqoL3/6m32ik/84tSfCgfrXAbDQyJ8aeDZdEmgsJqJ1kWd3c8CNE7
a6kZuBaWkZRowPpbUf/jJw68ZxSYd4obJhHi33MwCm5FJJEYWEi+gSt0UtLzi4pW
AxKwqpE+3OpXz6lyXCuejz6Y+ZQJ7ufjNq5qgkpIGEWGniJ0nghHouGWc9U7ou8i
bDSXT9paSmyPo7pVEFKYSLesWrBQHU+Np0I+ug1t1qNt+lONO35+ej3KfzhrX4lj
`protect END_PROTECTED
