`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRCM4zAPKH8X06/zozOtv7SiNrw/0jgftzZDNNv9aOi6xZfrVd4xfwzDdE6xHkpi
ff8uN3hVE9A4a2vqtqlNXW87nzRgZP/owTEA0L3RcnatJhtKbJrqJ8fxdIE/Cn+y
IAbCtxoNe1D1nJfFAXDlXapuU+9szl/81Zxauk20cvC9lwNFFwm060bXHbBs3yev
VI5Bw3pxQS9tLkeHd1BwxagC7LrMLt0l55cmsCBuqnE7Cu5ZGw5j7XK96SaW19Xn
DDTLeAaTXFCkTndvxlaKAnRtkSfXI4mTJrkrffktu+un1j0n87+XqD2ZtfGELlyX
izeG/gKesI6W8+cu2rK4c4T5kKfwmE7Tz/nHaP/4D+zvtO8hK9rjOZqqzN+HCb0Q
EbMPeBeCJ1i3zye8RMOXHYuy3WfbmxyPCfdjD9gBnYokwXnvzVkWpR0ExwmmUfTk
SrqlWYVFpUG8tuW0PD4oKf1V+CjxR9tjPDKosOfnw6aXkW4ANNS8vZTP8kEi7lvp
c+5TUFzwgv6UA+HfMBgTjTJ4QGncfyCs5SR4PgxCwl/HKW41qzrNQhB7KLRUpdJU
3mbVdQ0UY6eOaOTcz7TLhgObXJ8s97H7xcBqDy9BW+izJzLjDEU0hBzgYu4kHAPP
UE2JycI0NiYm5vSbU8WbA/vi2mB7hCGDeTIp7s9Q48N4dUvybl+IWBwY7k6upPtt
WB5DMl4eVd0FT/SPTAksefcgjPla070/udhRMVeAuA8L7wO8pVaGmd1mfnt4HGgI
xMxV635OscoBKPaZnbNEA6bWnpkX/MKgsPjxDtphgOTlllV2LbZ6LFVwuIS1s8CX
sqdXklhSWdsIkSiw2bsnAg5qolcjhNiKsGSYytQnKHt3v5FfccvOXTOeXng8klh1
eupLZ95ZeiHue8h5i/xCh0f4EASr675pj44LR+suStPVr6zpmX/OVB03hqUKXwKi
7lwM7i58BfOmOPkmn93tfBFqcEjW+DzN12VwoBYjvvvZXdzlPt0RQO99doE/a0Ir
c4NXlAbJISHKSZZcL8aVj7Ah4X4hn4WU+CE37U1EwuFaksuKD0FvaPIloQUIdoQa
XkaBiEbw/YkBf5Lxd/Mz+bD4sGgjczBTxnFpy1Br0Ox7zKYjOU3t7SH12CnDgQ2i
NklTVEhCmpii+p6akX/hOZfmfp8GhYbvv4fKaXFCQ9UOX6dHnFtegfHVlNcGZHzV
ZYLwO6gYjwQs383pkIPUoGXxxl7iz/9qmsEVMVA4HzDTLNAo3xKk40+GUxG//aTE
QRWjyLx2EH0Hrf0SR3COfipfsrB5gsOvtRWcoWlhSlM1DSgZS4S/14npr9/+FrbZ
UQ29pacqy27gdoHCvwzZmnUXEFgXGUuo4hfy0EAtiS8jbAMcyeOJYte5JeGCvzpU
cdolBwfrFGX2kWNI+t7F1BtEG7STVGIS33jyUBWDGiyH6uqNU9qZLaPyAAfMuiVc
lWDEFTUzmFChNUq5iQ56r2au4m2qZ/Org2TYzsF6BZeFNLswR5ZWxOaPNyrLv2Oy
Ip0RjO6o47nNxF4mjb8brJdCF4rGOvljQE0IpEYf/Px7dpg+vYWMoc1ryLUCIyq3
wEJM78B0rpu/PqLiIno+NMr5Uj/Xgq8L4ocCl2mzmKbkFEMEYMieDv3jBLaaMqi4
5e2qN38uJx4QvK1zYuQe1RlMljRKvXN4geiSPDQX4s/ryoo/YQ28XrGx+verhZQc
laxRcBiJMKMhKNUE+6G+a85UbtWsRUZ66yaHi+Q/bdMCrVKdezKZ2K5UB1YZxPGu
DwpSw5c6CFdF+Cgy0ycLeYX8yQzETDDNSZuIXtMfzLDfJUNcd3DppHVTSv8OWwAh
2JKtZk6H36IA7t9rD/9etqVTS1wb7xweeEiYOI69mNZmCrjcgx3aUjtDqfO7y6rg
xKJXxnpDS5SibeavXrU+4ZVs2gLPReuDN0mFdU8WL7NaP7Y1bEKC+ARfdJgW3WJ6
BcKHaLSW0qTZiA+EJmdGvlF0de0Pyl4I4ZHEilXgZSx/UhYvKjj6CCLLH/hwtT3e
cvNUkarUa+u1JbsLXfuewFaXUkRWrSGQZUHlYAy4wH875t9364g/VWePocyrBG39
G/LN+TGtLYdLNRPkBF+QDFG0unV443GTT8txpIohNqnZ+XpjGBM9PqvJPnD/Ok2s
9n7JlAmMbBt7tmU5nBYOGbT13JvbxQ4ELot/WKPGOKB72AoQqJFwD31VAzpOAv/m
BvFGgBQDRGZhEiDyOINbGyjtlfEcPdS79WufoPBjNt+zhSIf5YMxcmjLQOdgU/AN
/vd6xh1605/+VnWPlH9B+bUxVK8NpJ+B5nsqmkvDkQDRncNlAPvmdRae+ouzEoVP
4Ww/aDrxXIBpGCJkUiAJqeE9u3wgxXJ6fdYEN6YFLGq5vGArudc7AgUgU3A7q5oL
4sTLOH9DiHZca3NI/KsDi+HBrj/mbKJZNIsNADBAIHp3MboIYXDEijBWm9eIqRmX
HhB3AImN+SUrORyf2oBQYOTdSvpBO4BNV62pX/9kOPsO9PbIz84MG09rcjDVUYx1
BsHPgs/fMQC5sskfhzVJ/GmsQdkmr44mMuGYcBODdPJtMFloSCTvdNRZHhOsGMO+
groZ+R9vgsBUzXabcJ4v4gJus18KpgIuz8tbamIzAeC3R0wcIFPsiZQ037MKyZWU
oh82y/bXBkkwd/HuuJKjiyCLTF+IWXYdwgSIP2+DfXv2+LbeVs/TxRuyH/0SRyWr
ngBTlwjn/1A8uZUGQCnOakArL5vVV5QE9bzlWNFTmaCS9PcnvzGr8YMnn2jPKGs4
Fqod3a8TV1IVaBLQK6GT47oFFVNz6Uooyex30p4nZTGaAEUkTgxpHWVhu6a6ip19
ffMZxoY6Tx0are1sQOzKBJ34WQdGmixRMy3LrHHg/L555Pn5pUnlFqlPZ0umTsMj
U0pZZ2QY0s8KtrFMpEISPcVszbk9YoCaSIYN11gaLUoGdvhfgfvP4LZGASXHd0Ov
U5z+v27Ju4Y08VOa7pIXG2Z8MH543grwNdIwknnzsSOntnLVy2sg1PsPEnmSE5vw
UK5Jpk/upzSyCIm3tsy0vGLs/psumTF3L9s7BsDxl1us4k/yqaWwEFTrmpIl+pn9
X+GpSt8/hBSHLWPpTMRe6QVrA6xzkGHNLZ1GWCqmavBt8h3osO8uYWMGX4PzQpJH
mhcJyZHTGpeg40BnozkKUQiFMD+/5Xhe+tIpNBMQjxZrcrmLa4aTgVTCZHD8SscC
685XEYpIqxfdNtrcZzrBnmQVEqLn5qCc/JHB2OSHMcQm5Yv7i2H/8309IrG3Ysd7
cZqlqofSwgCm0VBPD11zcDEHqayz+SinMbbM3ih5MvIfuamFIwkb8kgcze2+gifN
RyM0BdoMetvmTJNN1vAAr/B59jsUGMfJpaozyzweQoQ86oViGLisek8reHqozM1t
THs2f3s/d2K1R4AET0PXuecTNsYyz7ncCdMVKdOqlKnNCn+8hUI8cowNzw9Ue+JD
mfaKKeDNc17PT6PniWhvsFG6ztjm1QzZpOHHX5wwzI3743bFKhI8CZmyXyQw9C4O
oZ0Dsz+nXwQVKH7fM1yzp5DI7M2a3ARLxvuRTIhkZ565jHz3zDyhczO2hFlTBhyr
8OnW54/vd+rZ2pJ8xGojCBJHWe4HM73dMWet0TsYLgyXFLb/iZMQTvpMX/fJlQP1
ei6YIBZ+og8zUdsoeKOr70SCBliBOF5leVwNybYgz8jjOTjywSo10I1bkBwXFRIK
pHjEmcygK0NLkUzl6jCBpp1YmTk5/stuEzz492qsRrlMUG6EkM6WVkkBb23mF/lc
v/ghheldsv6dhY5SYWcORuCmPamXK0lNleOEX/I+Q/eJrzZWw6aFC0MmlmQ63oIk
8VeDRmAWeQy9wGX0y1k146OCfKopimVXZMDD0yNw/zM4WKq3RIek/xwVc2akPgFr
BpFc3BjlWWSP/TZ/AD5OOaZ9HfPG3Dxybs5HNQCPTcTSX4xxcdE340koCxTGkny8
mVjyoc9qrXBvZz/SyyarQZHQIALKDar4DYQAY7xYW2lkJ/m324tGhdMFkXFMAmJf
9dmcOP4F7SEv3PwDMinrjTtVIb+KE+VyszvOqWZcEuUslPnrvYDN7Z4Zi8zaRoLF
ljCUPLDnV2x9heovk17/VFOXqQ86pGJcLRj7t0fhSXufqB2quilTwZN1Mi0tzsGV
ywRJog3kT9qL/RrodGANYTj+e3K+CcLGKTqRXseFupLEc97+QUXgIWDa4I/ddoPl
LQf3EppK7ItIGf3MbAxVbGd/FhkEMZ1mU+0TnenriOpB5d4NL+ai3gvw7slDvbwp
RaQavG8bX9OyDH5lVDj/R/4fOycsjlgCWvaSzVDB6qf5JEFTgzReghUSBxTFWONJ
2SoDqaDAG51ORlfPxjG2TwbP3oNu+pePTOfdN6mgyihTBfL7qFCcA2ia7bOJ/10s
S5D3T71aN6iIIxZEuFNdhO1XLyHJ0SJG38qiUij0rV9PsNHXrZY2fNm9dnLkrxRe
ipXzFIJtiHb2zGIM0eCAj5WavN71aZDTPeoUtsrNQmanfNyX4csxJTDVZINkbjaA
`protect END_PROTECTED
