`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+1aPQ5W5euqSQ3+Y5LfUSUtIcC9Qy9Qs5hCb6886N++7qy+AKFPOKG3wiX/4SCe
eU8xi4zrQKmkcWF/tM8K/YrJX4N/XKcNaXN5m43dh4bGAY6Lpox3KeXMKu/WuG/p
hFrRaByetduZ7xvUqcv1otg5hhk+rAMLhiNucGzsXysJLmZR4NPMCWNBXZ5bcMe1
+NfbpITit/n8cd9VW2/q5Vzc0zrqzAflELIGAVq26xarFbg+7FQr5RedvqhukB9X
k18Fzhm/o5rT/KtbZR0KJHj++SGc9D7UkISaXhxp+zZANtRuaDsCizdb6v1SSiCh
ChtiZaeqRJwjdlEoKbzRaYgm5ZTx09St9kWYSG3kDR+fgqQrf1NgBkmH09TIUEPB
a0CNviFX9DVkS9T0DgFfCCMTrVIfSNnvel2ugym3ixc0sxOExCXdVcLdQRgPUP3i
WW9HKJ0ifiAbQsiylJvs7z4lNdRs/PaVF9KizmnED8Vq1v0gKxy03f8ofncNZowD
zj5YAPMsP0Yrwqwvp5SDWBMBQr6lkVTimEBU1bwrltjlAMRWqL+0cUOHbnnnM4zh
VBuMD7k1str73x/dmYQA9/fBoS0KkYQRrqdDz/A5eunx+buNRBey3R1+0V8sp9DV
X8of5F7aJgHKPKZ66XhvOuuEOfEF3C+pLyctN4ppc/pSkd/QLqaLjjh2chiWrcPy
jonTMxshszvEafuJGVfl15X6PZbcFMJjNDXH2nuxtXKnkf5vSzE/Fqb/Gr88QH45
Y2vFFjAMHc/52HlOHy05xGIDnum/LHBKirPIjF3AtIXqIrDtoWFB+LulUtOoHJxt
itz9W2khgkk2RQ22SBsrhh6dMItHM38n5DAoQYAyrUhqpjGyjm5yBYQL9mYxLaVZ
3Kx+RHUM8AB1yWWMwkf/9TsYiWd/FSG6hjrki+Eddmoq4Dh8QnCzG76vpPKcuogS
ojBFyXE0bCbLZu2KlZ2Tw2Nl/SMWwQg5huuDazpZA1RLbpnU3vMooj5uty/ED3tE
/ypcwf+7UpNvR13fpMDIevH0OkJIdvXRc1pJbZFJrYAnPDtUrds73U9ZcFZHYyu4
6+Nxk/x8jL93+Xsr4AFRm8MLuIq2/qirkOYjy+yhUDmw/iLM6sSXohZPx4kyvYgT
WmuK7xmKt/oNEZqxagwnrnzZ42bdJMwk3y36KLd/urRlc/zxyflSL6fFT9pqsvWC
ujZZSe+Y5W5bHYegn3ujKWbzkGprHAKEFgS/JI0S1U051CYM46TFBZB54UNmS/Fe
lfUcJ6uQVzFNVx0jNGBQ9qQxHu0B2s5ThjcNcfKbIM2uh5ZdkcuMEU+nb6kRN+Zl
2tJLCpeXtsM6Q9iMRwYW5TpsMj3e48+tRQO3YUmlisNIVg78PRs+vLCXBhdT/Cwt
Vlo9qFUBppzZzgxHrUcpmTUotC26MjISEXmaIOTkp0ASAqsVCRXQ+Jb3CJ6x/h2R
MDXPTxo1c54tdInf+e9lUAHtyhx/JzjdhEKoj+3HGzDfJ5Hp4O2RdHmNuGdtUD01
mDfWu+TjrHTK2PqEHAIWF6L+o6D1AqmJ/bhCHK2ZYr4Zlm2GBdAtiZ97umjdXHIx
gwGBXoBOT0P2bFH3vsmPLBf5u8V7ZFI4iw0ANZAvGJtRCI11LMh0V9o9EkFyrrPx
37fIuUEnMTVW+bvQ9P6ri1k6eoSFxu5tPAwQRHMzWTmYby21GFcpCDkx50ePwMi1
FJYly27bmfYtlU0KG2T51zsLbTGtLQ7uJZ6QzwkDBQBTFvM5f4GJpx5kQo2HqVLn
K+FifHcoYrcU5GaiJy+rzogR/M5Sr/Hmiu1m4dHe8t5eIuMYi+SHvQ2UjIIe7d+0
z6I1hNZ8u0VJnPz9zFKHTODzX9yrpwGQYKcNw2eRGhVtVJOdYusxFI7QCiV86dB1
oeg/gwevdx1i+j3CTN1AuLDdRv1n0pHrooWYeH3ZnKCd7Vl5gzuwl6MRkh4AbPpf
JHcCB0ahViEiddt91uHPYQx5taau9IO84/e5+IdZOVVDp6HFnKVTEIpHCdTv/Tay
V4a3+LNM+cygQfpRqXyDqnT4t+xfZgekWhmIMRN9yxkNDv4kt2lKc4MoQ0MKFeXb
9bkckEoBH+nr2gw3r3gSKZ8PYuOP8ILxYEFGdD8+Plxu0ojXs1leu56DpNAJw8IB
Bo41oEw17RE46YqcYZCOzMWRcY8TRn4445yVc2la/LKz0NxzEfk+4AerW9xYhgBK
Rjjqussm0NDonxZQECwnGfF6+3KozU+5NBpEihetUnpMlR8mJhPnWSyjeAfMyltv
6u4urvL37WwKW4lztkD1/0O5UeFSD/Mm609LQWKETwb4Zoa+R4sV0+qR+u8GyoGY
6+aRgIWo7wTzlZgzI13enaNN0zD4Cpqa3es4j7IzLNLUsYA+gi83YDhC74mw8aEx
GVIZEew88OkuRibxUBheyuYrkSzJuzBDmt33koUUTJjPRLuWhYU0FVpliUyohDGl
hTZCWTFTHjy7OwW/lUbWGEGyyZzfFLwMyIRUgD1FzKKpMrw15ARpje/I7HP8EsK4
XPg4c+4IUNoNK9Sxpi7fy1KgcAflttDLXr0K2StctomT6niANLKeLDcz4JmftTO+
9ANgwasYckbuWSXGAGDYaTwxL7iiqOnxy9SdIcLkhx3qeKDpCdyKxVQgKr1iRN4S
TPh7V2gAkeq0gZtqFmW94k9MlrbWZ+34cgxGUCN8OLPnAwsDuJx8BAl1nSDRuUOd
XN0aL0Z36VPKjq65AuqKVhB+0criD5XQgs87mRAiElbvdbC3yyijVPmsqE4zIPY2
pnOeGw3VsFctA0UGRKHVhfI6jJzXWa4MxL01ZrHiCv4hOOoA7ez7cGQuyc13o1LI
JOkL2dQzciLWuLx38swoyvGqlgNcFpotrvM5AZS1GOo4sOsoQXhtrAyWm9sJgyYs
SmusqkcJJj4kgaNEM6Cih9Sdz0pO9pFChKsURDmFjD7wgcB+tEtkM0bw3MCYSiSJ
3AfevbA5/ruaZbVftrcRNX2vVNHxK0L3WbB1IGHCz2F2U7lbCKgjCiCLP+lPXA+n
qNpRlCGLB8ae0QnhCD9lRNOEbNyc9gMWUvthlfL325YVfY7rj4rsk9jKi7OOE1Y6
DBgISOTBCDfRQmvETcwg+BQEnWsdcrqSblUkSOIUtopWyVxvH15AJtEgNnDOE3eC
AYUeX8CD+VV3wO9BIrS+SkLoIWOt35FCmxGdKRdXOdCEg931vIbQyxBatQCPAM/C
s1hsCep/krM5NFCLP4soeBka+XksXMQV7TbPLoQvggU955ydWu8BT2II58p71xWp
gXLlSFLdBz8utxA/TX2etsN0z4Fi6nDIJYLadpjgWcoL1xNCec25dr9eBhrFFbCY
ovBpi2jE0y4a+ehHfo6504oEobyQgyz4bRJL9JLY+tr43oSSU6yjed1NY84B3X5K
H41Bmrx6/7L0qbyHyVj3VLp7NMh4RFTS29USNoj+1nmGcB49Zi+1WcvdXZW5sQoA
Ef76sCrQBPjVrVvQnZBjJuUjQEEeWSCOPiQxZp9pSvhOHSV2Ui9vgPGhVY2iHgDu
A+DLl5vX404jRbNpf9m1T48sjjUenreclbXA74GxOcBlyT4oKJdt3RpXubKh24S0
I7AFJkVXGy09zDzIZT7LgpDh74OiF85dhx5IUW9ExW6v2/HShPB2dfQ7C5A8gfxd
YZhgvl1t8R2EHRnepXZzYSXzYPn0q2/vKbxnXfjsYjIjVbuQOZ1rH6rRnZJJet1l
qzNmwbWxr3PFofjvkQlGehHNh79rs/PN4dHmo5W024XSFKXf7QFG2Pe9ESQvIne+
oVEME/towrGl49qSQ+nPJ0mYa4dqpz5Y8eh2SyKLsGVjnVUNlWHCwgivk9MPW2dq
aR3luJmJQjAeWdnsVCuDCWWk/zbhLZs5YNpk3HSEBLa9bZnB0DstNqorYFdtnvVh
vnFEwSWlvb3GDhliVAlfv0wm9aSNMH5dVsSRBSay9XH1n60C2oJvv7QkqHbzJdln
ZfphpHoPOK4UU0/wmF/Uqf7nk2HLGVT9yhnfGSi5xoryUVdTXGXnuPcpAjQbmBoA
6UysrPdtTfPtYgpKVNgShyHjtJqiZ1tMH8FGOlSxcOgpNdtaLfU8S0Ew+Yo7OmZ2
apxnjwQU95d4v/NDTxKi1HQBoaNl7WsAoX7P5r/S9KKuXOJGJWgVjLGSm6a+e9ZZ
EmVV+W3ZxOmRO/OYqjZmbUMqXU3HfUrKP7vIt3zfPyQRSgUEXuBhSVrqIY/DJmoP
Wg4kfU/exjPs8Yyw5EAP8qynx+rSqKeMxY72RiaZkZM24sipmTwglmF5nT2CLCo5
b3yNuntcGBxm/3TSBCWjdBuIgy1FARW+omWqQI3Q2jzgjjoJYVAqUCbHizNnVyCA
0P4uIQWxEMqink7DlDkueLWxLa1UtaVHDPygyAoSKUq9oLs/OHcvLzt57CmXn+tl
PsmpVfJJqRFWrdE8Tf59EXh4WHqSCAJOjUYrH/L3AVFQY5E0UW1jlCOxd00BxRPx
It8JnlVHlmEVpJwG9+i7PkTNSm3Eq3ieDstlHho3LOGE8zTmd3Ij3SaylFGsdd1l
yoGGgZ3XA0yu1r2USywfFM03t+6XcRQ9Tk7+tURlauRwxYqyee+GI0u6MWubAVSJ
JEf63fg2VexYE7jb8oNKZFwWEUExLXd0Mfd2qvS+OzmPUt+aZqF3GBSku/T98/m0
7Q/u51zRsRui4XuZbLkddUhSGUFgr8+N2MtOmp0lLFeEyrIRnIKbRhfhVevjXPtm
gdWKcQNoyhuSOE3V8erykNykFrw6Ng9pRetf1D32tbgHre0W0kcKPQ2DPQVNITYn
hywtI3Yp+C3SPN+VRi+3bEHeG5OKoB+5accYZZQgBBNDWW6JsRvKK3u04cNtjhkp
W9KFRMI1ZcNNbW3cYW6CU2ZGkDKC+50XCtcD2SmUIsJZD0VgPJXYFHJYLmGNY7BN
Idgvf3qcajmAJlhinFXr4jIyUE+FD5Uo/eE5cS/0I3odnxjgGoL02afG0bQsL9wO
pk+99OvnLHFOTQtjx9+a8tOXnHlWYpwYpi+ku6CL4N0VMBefW2wVh7LBkLo0furV
O2y8Q9rKf0m1gChBbQ+NhWs3a9TaCdkD8ufrEKl4HE7jlcdaDBVa8MuG4bevc2cJ
rSOUYuuS09PGxiOCoF/+ecuzkHt4pA1+l1HGNgQdvUO0ELzXIqGs80WEkfGulp4d
0BfsiSWdDYFo4jT4HAHvl12pErqNr2R/XHAbmSa1qjE2loiwoYqvZirJy+hGOfAG
1Gs9/ixR9CEiE/Jyp9LhRimExf0OxdMLjQVcwrkUNHzBIqwZWN9eS9pWTwd9MlEt
jrBEcy8ZFMDiPX06F6r2sjeCXRBXgvE8B6xWj/fT3xDSij4a/BSViL/BQtL7bi45
hGSmyrCkG7P7u8/0jfseH7ATXtN1s+HbOuG5INKjnELBLDzhToICliZ+rCsAVHbf
RNnh7AexWkJJ0qzAgnEaYshrCmJvnHxbLfhDNrPGYAHDs5LhPHe6c/yedFSY/xBh
e3rsFetPFCjCu8IekgyaW10r1+/UStzhXUa5EBw96KCf8mp56VfxQUGO5tWhta6i
aLl/6EQ3QK3DbPbiGFPm+vbOxGCdwLrOFjbMmAuEQcdQgQ8ORAhGy/xLbhwYHtDn
4r9RMf+Kv0Cq5AY4c4PTifwb6VPrheIEUurz7/8zkNbuDgAiaV+HZqNsNGnhj+mE
RSqJEchmpHslsMcYak6dviQLNJ8jLvaiTOL8fF0Rdgb8dEmxK3xjSh1xdBV8CPxm
zAlAF++LUuZwDoovfQz0UPNPNhaRBAqDWOCa5N7MtLAXRwTVABc6Py8p0ZIWxoBI
c9ToZq1zcOuRGCULa1sxFW/FYnYY7ridg965V4UGQdQya4Tq3icrSqyYBH/mxDMe
Loow52Gckst566nff+FedndWkHsIjEGyHHya5w9ZBuidZ1xrE3/X/ga79n21uPhl
PNZRx2chHvzPlUQgBYx9CdOuiPPOJMET9ihTPjL30Ou3CJzblbyv6BdvS8hVW1HJ
HdP41Be4/XECmLovKVUgNuzz2vMJVvVByfvCn8w8m9oWpm4eo24PiG3S0GXp6iAR
xemJTKm2z0gHbpHEZzFiW1hwVYgQ9zKHVCPmAovTgtvowIGVpABfns2reRsYQOHC
vtJPZTW+lktBZr6rxoGN2f1p+tOpRWQD9Mv+XzBQkwVNipsT874nqxUGBQIrihsZ
+fXuHb1DvPvjvFJmxFd6jGjO6LsxrHWvgNyFTeckT0c3cEPnDdPahcvaYoafL16O
9TT1Sda8uYNAli/XfoOM+cProvALOqIQ1N/pyI1xR9I/ta8gQGvMQ2aEG+eUmtSo
lcua9UVrXMwyMWGXPFidY+/ldhC/hrjBjx7MnjKZVUWW67CWxUEYfGyWJNHTstXo
dA9JdyCszor0EpkGw7vgmR2nSAaOzZU5auALqLesB2MmXNEcjgPApbs99ZoDnqji
UGLRtEG/n1NHpwxEotfUrvIL5YszUpodSyn6qF2/M8GRoGYpJtWEjsHCkPttIFuW
AUi2DjmBV45GP06ftMZj+KCapys1yLPrNIZSNlUOhAe13e+6PDek6dErcPAuqZ5i
1Da0otVs44Ltq7LkHWYXMOndfJj2U7E1Zjchq7tgHvzD0f6dEXjOmUsPs++QcSzG
TPLjOTpip1/aZ66EyWnYwiS3ZAwfBCPGCEJ9OuI94CI50Ol9aswMvUV1psyqhqhc
aaQ95VarWwCfNfl+HFlSgTHyca13vlLdK5dhyflaCdhRiKc7JADmHEPVgXEesgRv
0nAkQkibieymTSP29f+PXpIVp/SxUnu0Jt3OaNL7XCHxSpubuc/I8lVO1xStCR4U
ObmxmMEkg96YJAUVEqXJC3PbMKS0yUeWtiHB/3Bzkh/w/hqQRVgVGePWb7+LSd7W
UMLZNX0O7WQgzUwSao6ipdwaBVo1wTZtDJBr5icj9Qtebz6Nxr3w+aW8PsiVBvC4
3H/Tfhf/QhzToqPult1FV4YyzHheoJn0YyRqAHEoX0A/bBdXprOMzF2g8mAWkBA5
yLp4Btuvc9VAOlM6al04KflSfn1l/JaK6YOSuwKCELlNgC1tPV9zNej6EichhdZX
R1B5wJhKrzmIDMwVbGUkmOpFU/5z52WfCSLhNddjm1U7uzEABin8Mn9JGUcDNDpg
2aYDJTmtjzr/g+6njl6HYp3zZYmWPK6rQI/jKoXb1gv0BV/ajuvv3vkb4ya39ekm
slr1CsgGDVRh2R+OVQFOj5nk4V6d63D2mfOHIRJle2gmEeaU/8eJFiWUB9hoYtAr
HZ91QTNrm75Hc0Z/HLP8SFJTBw1aRV2sed77oWxexwKAe/IuzfG5xkGENghvmgr8
UAjpfWU/5XItQfA87e5VdsLav6m5m+T1RMfI1CUwzZbHG5lZnU+DKklZgf0Haelq
Jm38EELarOzYweH4qawxerEZs65ZfWhjqw8HP+CSn+/cByXBrw2QTAr+RWFqPwlo
l5oZpKMz7W3Cfp0eJoNn9cNV6KbE3vPgLwu4CKM7HAGJBtDW100owRWg6eEkytNB
fm6ZQikSjjCrpaqEGWB4OKp4ZdBlJoqvaywZhnrgW2r13UfXuIx6ZrLnRH0Uiz+a
umQ9OWK2sZr7/WLollKcXSFGk51kkNX+6Su/Or5oFo8lXa6oS70cyPR0Ax2vaLv0
m+XV/nlilYboZe2DfMfcBjGNraSK2eOxUEFPWgGK4wBUiA6KuW//UrlDjL44yT67
Eht3g1NicbDLz7tmCQKSZ1Uj7WA2jBRfFW+gnccOZ+bGHENL/2/8tq+lkloF2zqD
LBQETxvxnT1MxlQcqe7aVSQiGawDiTGod7atyKtL9osRgqqmSLcJQ/OiC5QunXK+
aiG4NBvvkvHVOpUZwWEG+3G7wSB/0NCUPyZPuSdiEroUy+pLIhboUGNjdD3jsPfS
PdNGXccjSQCaiJqUO4o9+12f0OH0Ad1iyPRi5S7kSNKrfskwz1WRSRnm9Yzg4E7C
PW+3m1FoyJvtbWFm+RWJT2S0Dz2HU/FsPYMpqS6pcN2TTF8o6EsYM1IhP/XUfuJi
92mH7ftOKeeDlsNNU6AwIaYooArq7sYARdUAdevj+G7FcdShYMJ+gXnHXAqO/iuY
3wfptf79dJSYUvbp8XhlTr1CAy+m3YFuy8lyPji30HQaqSsnAdj3Acq3dzkx+ghN
yGdkyPO4ySZkCFcyYvzx+2qVHlRyv6PlRVprVidq9/9/17ExOtngVzMwfXNYuwa6
aNR0asOK4DzcwtDcMU/lZk0KpkHm5TbLJJk2j1vYR02HNhVMrOGamk7cUoUuGg+V
4Yo87HuV0r4hF6TP/Wmry7E9fDbbW+/4j77vDnP1+vsztbJkYWXD0xM4jhmLrjXW
YQ1CdJhgGL56Fn3NmB88N1MuzM/QTDkeAZ3KwpUuN9VfmYxvFR4htFoPUAadGPsi
zHvRzcTdBN1SlVw1xG2HEGfnmOAPEj+jy4khyDQRtuyTUOzOqUkJahS4E1AhqotX
aqWtvfWGgo/dDjnz9tH+D7a4bexWBSkZtPS7iNgqzIkajn1MLwk/66W0izENXqeX
9OE4sfIMMjuQsVVO8zKFPrODk7sZy5gEbFRVTQXu9ShbXeivjEkVbbvkZmE0M/0n
XsHnJZRIz5loM5jVDClkyk7OO1puHiK+fAiI2mMKluQd5BKSt6VGjzleJ7O756Hd
tSkm+OHnTOg0yeI9S7JVHW+RPX5+8WkOsGz8HUFXoX7monDe3qzP/dIb1kyBnVl2
O06mvCnaBowfqDhrsEHqaXwE+UUadrAaN5s9sYU8pCaOp41l8CFcOQi42Br+/F2s
6R+Lr7xKYBeANWCP/zdxgR//ZLaAIScxTBkja7w9LJu+vcPw1BezmQvfexI2CqCq
VZX/feZGpZmdIzHlV+Z+F5Ox9SJwNwC3foDrsXfnJabP+FpAzv+sQxsgkD3YpbkB
7aFiGaRF8VhiSQw8yNIQ7BbQmwSaAx53Z7amrE1vNR1S0Vz651fexdALQz3G6ios
vSYRopGYb62dxb5vewW81NmcK84UUDhS1CI78WvXtnh+OoEwNdxZw5I0jjdugycF
QfE62wxUzPCTK1WAi2fSdcL2lR+rUn1JoMLvKTz+i2dqMIeYGMeMOdntG5ChmoFH
3TzrMYOF7FFOnb37mqSEf534IeqloKSHrA49TUj74pDbUn2IRo4lsdr/P8vSAIZn
62Db2EmdQ/EDDW6vz7o2K2W1vr7al+TjpSxAi8Lhe4eEATb6lCsX93lPCGi2V4d7
yIsh0c1DCoIBLmaijK660tNfQPR22dsRjm2l4uJjMADzTBfHNMa7M0zsRJQcxSRm
+HABXYb8UmGtkTEukXnOz/2HlDVV0COGDzSqB7cLkG+MCWBFFsHhjnE59QZ7cLPA
vTYHUanVSfUXq2/Qox0faFMslAjCDbl4cqULtaro3Z5q18AD5q2iG0khQQ4psmqi
lTVlKNui7KCbS/4ztHixeK9N4vyTSzjB8KIGA7VejgzBrpwJPwaO3m1joLnJey6h
tNlBzN4VZla0nFf1gGX5MvxJdYnaAZ49KDggNaWeVdQP2kioQdr8h02r+nd6AukY
rXYNmYB+KRradOUDF05Wej84qwUvRECdlB3NJcOzolnwMt65JoPxG6rdbk66kbJp
kCyEXY6MSCm7+FxWlSE/la1I9z2fl55bUeWVgwSQ98uRZtteOaUnAKHrz+I0R2Hi
YFa0uAw0RbMF88zPiny8+pPIoAJ/6l9EW4apBTm4xaXbyNu8zeGE6TVL/16mgyPN
yDw7jPKows8agwXnjDE145HdxQK7+J4RF5jSv58grtoMiCiFi5ZaeaaVKXpSTJ0q
XYrQMvy3C5bRT2fG2VvT+EgaOwf1CAZDGIg9EBK2EHpT/NwpDT0GQsqaUElgbKJ6
oAt5lzRudDqYZTyjgiHl3N/+fn5tZuUtJ8NSirOKBu2eChlLb1ByaFEuokBSwjn+
5NMPo6jzH12UoijsRTB9MST2amSkXi89vCiMWdeMfx/G72XhymcRpCSJ0YZDAbt+
P84Dah5hSYIdge0DkUtGn7Yji5Ojiw0bIx5CiZJzBZgvDS5sRHakkcn/MNRlqUCA
YSKBK4mok5IwcoHQDlQFu/1Y+2crZj7UUprHBfZbkrx5Gf+hEVbP8rePmnEcCZ8x
BZurCyPoZZbWFekJAYZjBmbxIFUl/4lBppADcVtGkcsGXdBv8x1iyo1iWyau/OhN
8a8HUv4Xfhbc4B7/X77HEYqNmXqNXIFFdwdsXBoDjbZAfPmzQXVlkS9ZLxP7rQ3V
4szroB3ifL5pSSwy3YwPItaNKnrDvbJAfJ9EtbF9lQHZWxK1BZ7fK3BD4741bOiV
eWTSHs06I93HBzm4XTfhS8SIQMlPIQMjFxIF6snQvwmVwX0grXszc29uJ+nvzioT
KcGTOdkWEuPmpxm+3/6OGl/Fxjgpk77PRuZm5fmiu+bUtVROJeK6dLmbBA/nAnul
LbtGPeqdebBel+mwESkjx1BjnXgVwNKWFuxjc64cnd2w7/wiHFO7s+mvXb2yzoxi
Fyd31s4uUF1C4Tw7qAoll381bAtu9OlQZYgWFxCDN33VOSCo9kC3tTJzuH0MGEk8
FVCT4q72+1UPT48NKcKrq16dEFcYyEbNEdM2eHnSrREW42V8NwAdxw1Y7FDp5gtJ
Vj7SaqmdTc3z5Apg3acCeq9ezA0dOf2dTzspP5bN9Qoffdcm3v1pZ2yZLexKFMNx
QyfmS55z+90NTwtenIUF4tYLMV1AwSHZmJViAYnobTYuvdtrTQmEIh/3rFn+SSx4
n9gOADUVsL6e+vVM8WPJhYi6dV9KhEY+6g1ZEMdKPLX9F3DIu3MM+EezIfK9/7uT
qBo0mGaTjNPbKuu+z7PwkvVxTZdkw36UiefDUSFtAH9RU/EzSzPOXl1O6iQuq6em
C3FAWjzsMF0LFtQxbOHryIVhPkdPco7JSxfH8KRZSdtyYplqwnbGf/AARtHanaDG
EYdPvs+AX0y6xmE1lJLh1SFpJ0RyrNXcMoVsAFcpuQaRF+CdioiUz4I1ggUuX85Q
H1XkNC1JFqWlzQe3BCr5hlr9mvmSIVXccF9ElToEZleNdaa7AitJmZyJ7rE17nn/
cisvYJCB7ADsFTCH8Azm3Uxdz7ReibHRwc3QofpfPPCKAC3934fZb+HXpXvRxh2I
fwXyl0fG4UOA4NHesL/+5SH+yfNmrJsBGhM/KM/8OJ8URQhlht2hKEPnAJ8o84rA
RLV2vK8F6bRRZM/bcRKkxbZfhHTA1ARdKFxctlkXSEpUwTwl6b7CZsFE9znfRoH8
LJ4TM8zIdcNY813/dOSQ4x74m1iunhJnv8CeL/qviDZms3aoTfJ7v0r9p00Q2pq+
/oG1ZdCZDl8CXKdTRK6x1faObzJDjGOJxMq6zKoZ0XLABjDT6PxMdq6qrwq7UJLu
XT7vhFbgs1yMJ2gJQj8uSdIVH6EqCkczbD1oI+wt8y7S2Okg2ypcChdHPNQQqc7S
BzI3O1wudMr/dzWuJ4PR9Jw/ngW8pDn+QTxdYR3sJlHvQzIxcdLJL71JOE1uQ/Lb
JtnzVsMmksB+S6DzfEguOKYtsC/7ZAa1pJVsCoeYQHxL8a4Josu4ovn9/fpqVOV9
gsMWhrCGZAdAXzy+UWX6FSN7lt5pywA3GGszmQsYrCz9wl4E9KHAVYIW2DVcflrO
0kCZXn1xKmK1SqF2FVOuFSvYL5gsGtyytiiIgI3lwALuqKodcvnx039Bf3zXf3Dh
PmFqcl+zvCZWDQt0hH8ARGrz/PZdJgiEhnvNxOCSYozYIQZe4hqbfSN7HRPfCIsa
vV5SlrqgFNupPnCgLYhExhin6+nMAwLfjHvoMPf5pRn3VCDm39nXwdiXMf8pfpMI
kt3gDesfUt4+jiBNJS1AXigyNzlT8d1A4kNzgTEoplj/LEn1UPVO4gzXUo+DZkeP
R1+jWt2vwS7/OkAgXqZtAGF/fOsBc4cMHUVa9wohr8fHPEOuiOI3tGzLYYenaQ9Q
5SDFPrFORdi9JBurUed/QCnFHW5MyJZNrKFBy0EogPyGvMwIvZlvc3RyIRJYnGZw
Ad2Yya6qmJTfQOkCAHEqSUHiOQZ4//AJqeNkew8cEKf865tGgS7uyDbjo+9PE/M9
oqo9RruCa3yhhSdbBq36sV0jSUzhKuai2ZSveqgHaQlW2NdwsBSnu/3fiOXLE626
ATIl9rkjYTyaUIjGmZtdOtiYajFbpbe9PMWl+EWm5LxLihFNp0DZyXJ91sb2Wlpd
rKFeD8zGxMPwRVAnc3ptNu5gx+URtaCrp1bD9GeugCJmpWmhwvtpxXKOWRj/4yT+
LtgjlQ/Ns/lCddCGmXaaSqK4LXeKelK918QnzzwxbOM73+K1sz5p+iF2q1Aqu+L9
gUR9cde5LGae9jehZFixGz8hR8bDcroOlF0Uk44xUyw=
`protect END_PROTECTED
