`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJz+JEdIJi0BolTMmyhThQwgGqykJoBtSokbZ3N92gGT6mIV69wNnNZnhSCOvYBZ
gAhTHp2viXqMm7zYojFbBk+J7kIpXOTszPzD7bRNc1BPYPFmK97QoSu1qPTeyskH
Ddh1hkEAbThO6e3sAmanQSjzfKA88PuZu9xCEB5wBB+3WvIR7HnCZXxnXyGwDFqD
sKvm1rJNvc3XJGUBsdRdCojGlWgFHgc3fFAhWmS+PVSb8pCdYwnsEC0PAwv5j1Sh
a+uBM23G8rxpTl+EQ+G2/zvqK+XTAiKiqzVxrTt3YzmxZ+YGhIozcWJkA07Gj1AV
o0DeKKloQLYTAD56fhDcotuld6scycJtBHuj6ufsypobL8C/sKdysPvVH4cK2Vea
QeX3UHaKKFj8XwHe3/V28G9GCAedxvQctO657PJ4GJnNXdls5p31Gjv/nfsfNUId
lRLUqEaDQlYrApo8Vc4zq0l6R3gNRYDKYs33cxoNAebLvq3xa48Xr5fJrth23WNo
+DaFmB9ijJgyMBDkt+kDmAciCIGVLibWsJK3+vpGjEScn/5KIs4HFJJNQuWVf0D7
thVdvHjR6uLSqAkitHr6zd3sRiSRfE3hTQ82L45UhURWEN3h7iePm1Fm+IY+OWmF
E2V5zpj5csCRPvcT+h5J/XQkpefFFL83+q0i3Qfc7Jelji0eVDoGUoi2THhzbtxG
/VSfTAN3DhUo/tZ9cCnJxXB38vbI7lMq2qywWHZQy2dK9GyP6TMfToC7BCZaYqHT
IfNw8u0eD4pPQNXlYE5UtcwcFzZWYFj7YRP4H/UiiRN7s4bDCTSw7SpOYOtMzQY5
8rjQQk1s90BawsbLlDPqrEuJ6JTm00gnyN2u7kWqxxXhznEAQv3RZzfkXow2VH6C
mu6SdIyu6rAISJ2EheBNLF0fLZLuDnv9LddcxneDG9pEIiAbPrSe5nkkAwJFQUI6
6HtSuVacODofYY8GYG6lTeuQ8MNcYFzMgtMvBuvH+CDHvzhoaBBcDhx99AwERobR
L8HsVf+kOZyQiJJEC4Yz7opsRUTajGUugtOsP/O8EUXHdMhn1mJ/zcZqzpYOhXJF
pXJBPjJMKQfLXWbSZj78evI7lOmEkXqmCB4XnHOSpUjrteiHc4ffyQeRLRROw3za
hLxy8Q6gCD+f9SX8xikGWQEOMA9w2SJRCCI71KXoZhOP6STwmjJMNgPTV11c5LyV
bXZwuCohfqvCqTEboRmEv2DqkgeWB8u9v1RniRyKdQypwVt1dBtodvFQjrLgYwh7
Pu73DLkbyMzBTotpR4tjpPfqGusIQVf5ByrtUyMYV8it7T1lea0hqpF7XDeFQVsd
171IDTyn0Bazz0qFexDFic5K4SrGOFzD4jYpDbisXmCCQ/A6pd0e+hPGe6802Xmu
OZznXuv4e6v8CmtCvZGAyfRO2Aih0wQJVHMUKuOP0/ccnFeelnuvTq7CjGzVcwt4
9EoFepaJ/K194E3iE+D4/Bw4WpZ8bLxVPiRYs80RhfrEqsO1bEwZCCQ9wXw3c/Nh
WGyN4QAn85zCesbozRXsg90OeNA6AObjq47iLSohAR00RPalPMS76ASvj0YhwkH1
Qbillti+Ngmyl9G5W9bzOaiZ6R/4gxfs9FKIkrB+0nXB+3fb/g4JPoauXnxKvmv+
B2SOgG9IAuc3Vp7tZChGOpyvRTpefixKfnNs5dhJF6HwSsT/LRyW0B3y5UcqXq+a
fhgopywMZaUA4RpOLkKS4FfdmaCg6Fi5VIhgNfjNFK9ISrdG8j3UAyyONYvGGc6b
GI60bR6YmVJDevlUWIXal5YM9Y7/UqtgVoV0qfjXCGzhrEOcmZkjIPvsBP7BFfzF
hbkzEh2ifLw0UCDp8Km3sW2e+nkXOOKdZy1RpQdTKjIBBDLB7o1RtOOqAm6i64Ne
gfDqfJ1wNkJ0NzOhh7QzN/UmSu9qhR02xphUvZ8Cqfi8+zkBBQMux3q/UA20byyI
hS58j9ioAi1MY6Y7By9oII1WpjkoVQMrRNYxsC3k6q2FkYsskQ42Dx97MzgSPlSP
60MDkxv6BnMOm7ZtXeSQvpgciMal378rf5ixTflWRIzz31w4caM9A8XB3q0Qa98j
98Am9rMstlQgLU8XlbyNd7IfGlpupllX72ws+c79UmhzFtwp2X6Z1IuditIHbwBw
o/ZAnB6nIawTbo9ClsMIXyC0Rz172Xn5sOGkUzWMKmLHJcpwAMSBPVQwcpq92riO
qrNtttL6fR/Ws/oZycGOGT6ugw9/cgTncOtXov4zQJz+UijblT79I8DbnAI9A1/D
Sut9KEF+EJ9okdAwgHWIjB6MCkY9MZh+GE+1J2ZMMXFv3yIJtGDOO15C+lPQ/cVg
M8NRUWOEtgZWdvzjFOBhwNby2+QG7BezB0bb3VfweuTJGQkczIkzFaiYc5HSl/S/
3UNnpUxjR5RChRo3BOQs1aibJyFA6WzZIcTigjamrIeCYhYiGsMYDCYodTi5oaah
3AVyKePD+5ndms6Rs8NS9fMuqdwyXmv7bRWokvsdbRLpdBQuGzv8Gjq1o5bm6INW
vg/1eu10RjLJ+JGmQSj/zfNVemuLFVinbhdbs/nwONmzt9hBgOxC3AytirpFKCSH
T5a4nuPnLjOCLUJ9cqB2XHQCf7OGAwJ/M4ODXBxWQpQsBooRnTUM9wBZNKp5qTMI
23y39YM7llCZTGEfKdwSe0wWd7dU3Xa4osdFZmPMR/Rdildq0oKGCvCUOjg9ie/1
yFDfX2UgpMvcPnsxbuWTV8Ct1E/9sZtUhLiSpInOy/vGebx00hpjjjKwJ7eDd96v
4CzzmbA3bcuv5NLAf7LM5Vd1rwxvhxNo0dwSDfaxyJkoPED4rCDXclu3U19LVATy
2+yIU0mQ7WCjAkTez1m+4bV2mUtgkftsjNQiY3AT2OXmuQbwHz73kTXOkV4TMdcb
ioAtatvr114zuNM5X+0A1lb4p625VC4Lqe7OlusxV59Q44diUyQIsCqUV31Z6x8B
Vt44j+gOgU54YxCoLcAyme6vdmdCtwU0rFtL9SERGNo6vH9tR5mx8zY5fnz3eczB
3OhKaGtXB31VKSb/w4dN10n1hFMeqK9ZlIaZfXW1tk7SF5p5FMicFha9bg/DRT3v
SpK9y0OWTnw2w5uW/9uFFZTs900PYhXwSgF5VdAMYsdBn0cB/Df1cmB1MUh7/Ubr
mh53RPET1N9+Atu3ECsrL6xcb0y9n6IiyD6bUoz4D2hQlHFOY4BAtWwP65FXXjc4
AsMjl464nawCXa90lycFm+NIbd7A1CTFxQQl4hNv/iP3UxY6FKAuawNS0+rSsdpa
xKH91/ktZ3ynDsSz0oNttg7SopPN+n2NUGXXnxUknnFkrPtfC3RXYG5goo0V4Xhv
fCDFyiCTajFaD48lu+G/yxJDdwjZWcq+vkjucM+5dCNnP+7VxVGW9XOvRDNp6is6
K0hZ4WkOvqCTanhtDD8pHiFaOHiAS6H1dkF5EoDhLsfbiUc2EHK/0H/Q9P2Cg858
7bqjpLmtYymLN5fEbMXIQhUf7c6Gelvumhi8BRR27fsKFhj3wgOcCtHpU7BF6d6n
2YfGASyNkUSo6sjxrnqoJUhaYv7cqGvjXWDrAuapym7eouDeMVQC7Cn53gQMSSbd
OL6ClPYggos7UZ5MEQA60F4pS3Gpu+8hkUsixLYCdJ2gOx9LyDH6TAY7aj1N5wvz
GK6C6uY8i9zoaHRD9jjXRLOlVGgHWCIvelC5YTMaxGYX7iR41XLvg7QEMiwRQmzy
p5aUEYZDVuyM/ntroOnLqa9nowMAzUz0HizJY1TbUerAL6S1r4r7XWyqvo/m+CHX
BNj+bO2QFSLOEPdqo2XaJfB6wVxssvBgCRl6W6p6vvjgtLquOdGnO662SHQzsYFv
8FgH4EhUokir4qgzk/qKSZCFPAatfqgu1W/vtjTsVFdvuHXX3QH502PA+R2z+IFB
BIuL49lnArpucwTdlnm8BSM1IyYz3pwBJ2WVuJFW2YmBnUc7et9Xh3zPXCxCvVd0
ucKWuwFcpfNZjHa3BRNpbXECZDlVqkLwdjO8PBsOYbXS7+tfBiP9u1kN7W72xotP
84gYS89XQk+XhemZH/2JkA/Uyc5hBiY6OIyyygoaeHD+ubt7jCyuUmjhGH9tAwXV
PMgFy0vjU8LvtTp+7IReDtpCQaE5hFOcTatmSaSfuh1pvmTf9roHhzvo9nSAtCXD
rNeQ8zuDAdDDdR8rBUuyhBqyHHnjh1hpbG6zU2P8QI01DJbcTh3QTA7BI5XlIBGs
cN8uqgcoM2qfUc1RqEmmxu7+rLxyfadOVXCvByyCrIlcDisovNPnr5fs6gPzv1dh
vO5/yzfvC7zX2Sp5Dm94bzr8pQVMWIw5B1DnUYTyeC+rQBA4472ibOGxK4XoOMLW
aWUlfP7oXqIrYfzjn3gqV3XGTn0rKb5Gy/p9tjJHulN+Mhqw6ELNmTSIAkxz9D+L
BPxCge8r3Dfg3/JYB3Fw+TdGDNYNptD0OdOLwDPJ4g/I87GS0/2NyFEOkilyolLX
MqWAiKQfHnwSIKmsN8Fe7AmmTgmrSOaW55rld+aLj2Uhf/160g7WlpCLZ6ClDr+R
cHm9BMuuZpi2dUtqA1iq57aDbmbc8ATZM6sXfM+REnN/ta8x+UGxysC2kReYEdc4
g05K/0kLSEfdHMID7k/2tUWDU34wfLeD1bm/dCJImrApUsDp3bRg4FolEObrh6au
zQ2DLazLhKoOrTJ+BgZgBzkIER+6gSLQLj6I4A14C7IjZffg4Nsc6YUafU3GFMk6
yYe96oTtPIjLI4GjKQQjAQGgNJCen9uPhn/UVzEGjF6xwC1pcv7G7qbI2YhOCj46
luS1iVy/y3tMqFkgApJSZarOH4uYIbDvUp7WCjNDwM/RWsHULs4nMktr5wq1XB2R
9GeZPIp9M6aiUjfVaP4HenR+tuzyVn+QaX662bcuC9e1Gu7Cm2w20NarY+6wSDey
stczNGvIxSkDr+Hrk7A1OwqKK29+B9WLhUHDvq+jwLhZjkJvFl3OqFRzgx4n8zBx
3p4bRYkbMVxB5BQTzaGkrs6+R/EKBhJoYtNHN6X1a1aCks3h02NoPesnoBf+T+AO
dTiSE3ezUxYHgvG9Ep62rEgwHL8xcEURo6G577eCgRzvMHEo39Z3OrsxcDdj2K1F
MU1Tuy4esjAaViHxraaP5n3vdKM/A3lD24ZYQjmAYhuDdwCMDHaL0wNbRSsGuQC7
GL2OLee8uQuOiyZxX4TRxfv+ntcdY2J3WAAA+7T26+UBgUt7q2ZBs2uG3q6SV2oF
zfuTsbRsuFe0nQPTA6TCvRabE/M/lX8clU47D4asnj2eR7WUTQWiRrQg52o8Oj1F
H+FpOU2MeT5YxiOnMbgNlRdd4dWkb2uXA/iABfyI0KRsfoH8WFVor6z/2VMt8DrS
cz8ohZS2ot6MEuWTzADeNIl3Ha0UC1kJ6Op7Un+QxQ9B9CngRQv/GOJbWZgATI8T
QW0AZ2MnIpPMIYWReVvVRZDp/qz7LdLFsFGAxHyoL2Dm3vfFjvrgCLTeWP7cixiu
mksEG7AeWS+Ew+06hJJgr6cbqdrLNQ0wZGM7EMla4gds/yHrcTEtakpP14aqBi2g
HAIL4MSuLORs6Rf3EqXV1XfIZn9ADGGFVMQrhCtRP6Yn0VHQ4zO4PoiZqXG/LKnc
CtY6MrJhQaYxV0mcy+3PsPpWfDLu4jDTpJ3mClPBlps4A0s31Z14IeUfgegY0eQ9
dpL8HAl6IF83u0BmKn/6Dm/gN+HYynB49nEWbS+I0F5K40MvHpwiQViXs+HGxHcs
WYfmVprtGc0+iSlXcnmC/V3cW8ynePrGr4XOA8sEvjTt4bveV5YLmNf6p/Eht7RO
I9JXsKb0snx3o4LJU7xX8bzZqHfdVwJipdsaGzfbmBBOdKlQbHi9P0AbZ1Ayq375
iB/2Uyl+e0CeYjbrSJ1zgCTPBiehfS2YS/azjs7CiAnAak/ugwRsE13e/EXjvyK7
kDNEX02TTfhUpZEJSVekq63M95n0rIqeJTlBau+tjg8t6tMVeHNcVb0TVIuyrcfE
uooim+nRdLRsYR9UoVBGSJmwXqH1OehawX6DdohILeeI8XOfH/JBrvlYGJlj6Tzv
sFgU0R8SdM/8t+8RFY1WR021omAIbblDyhnsyLVJwbzcWvaQlOC1H1W8JzRA4IDR
Rd+78l+0oxJ+WpXN9BF4PAerApfdbeaP+wnp6nCvQvz0MRuda82uvVF6yRNmgld1
k33J5VS29sKLyhaeqXGhizXcrgFatCsd2VrqC3e0zsFsdg2HDWE/ph+8dDzhcpyh
d9I7Mxu0Y8tnujZu+vA1D7X4nUukScxxbBb+vPHWtq0AYcAsUy3Nbt5Vrv7SSXV7
7fJF+zwAEFzm9JhrZVfCIcWK4AAS4rnOMydwost72zRztOTPD3B+YoD7WBRaTII3
t2ofEesKf66L6HENxZbsgndBWg+b+LYg0oZJiyjzuv9RlFkfDyX4yXjby3wE9J9V
2yZnn/4KhnM4io7jfVqTQvxs4wvggF9wUaEe8KFBcMdhMK/FuifU54ue9SaET2NF
72REn1UIYTA20UGpH0DlZ89XJl0wq595rfk0uMMtv6loDTDKenmWUcQldFiYtGVS
xp2h6vs36co+CVmMrTU6XWP5pf6FxJTMX+HLlmB2gh0K5ARKdd5/gH9RJ77m5xfA
NkawtK3ayCPCudajTpTL7zD117eUpFJvhskc1oF0zHqvXWV8CHBtufLxqcOCkpVN
8IJnJ4Y2OKlz1W8XsoJMSW68Fk2Sn1pfIMvzaqyaNE3O/Qu31I0arb0IT5at1GJB
vC+JsQHcDSv91Kvw0kdWN9UAwCseuRwA09oLp7cHrEABJRuKhD4sBFF0eJals6z2
+4+QPFWAZH3bR+5CDmnK7rXJtXAYdeazbx5IWsVLuaVTwjh2UwLAfhGC/Et8TYM9
pvXYBF1+BsRXuVUGpQG6IqqKgMdhlx9sB7tmsttWBRucVlOf+LNnYIt5QsEE30Dl
ZfZcYFR/EYg1CxB93vZp7rqQJzsv/hVUAlUMEL2ZzOlfkcRnCxFtKr545wodBuCb
Oa1PzL7dm6K4CqT96grtg6AZQeSJxZ8W6De+06M1/IpTk2AC7h1jCabJEjrDppAc
BOHEi6tajtXmLVKAGj86Y5fYTDd6zqzwDYRw3jNaqrae1MW6zJm1eO92e81v1e7N
KYdC5szxAWfILdrc0d5+JPuArTOXGD/kp7YhLkQmMi7M4hApBQvEERm7ECV3pdEi
K7KC5JHIYkmRH0/3KJIlT7PBH3KMadGzuQ11Ewo+FIkFiXq9y9ZFERxsKLSH9pG/
ez0WEN7uO4j8ry9qXT8ya9B2G8B/sL00D8j40alHq/f8VnmBLyoT11+8QAa/FJfI
su9iuEEjouHwsQPpWrLF6/Peoog8xhkGo7BFWwgj7bXluPxouAHm/+cu+8Whm1MF
gVLoprzyKyPejLCG2TqOWuBKlNywX3r0WTpkWB2L7ktoG03AQvRZA4q21kP46y+g
0CgECBCA3oI58zUl5iZKAmrHEyfzAA4HWck4Jp57qipQscS9wLmvtp6y5dUBXSz7
yS0EC6fjX0TRxafqs+lt18IZNp+37WpdklFLCRD2UNh615rd7h4FwoPc6/Ol6eX6
3HS4cS43UdLO1MVIacltUUfk++LCjO13bZvA5gwKEGbO/Rd5OfHNKvFCZGjnOp9d
QnZX1uC8cDKML/Uu/OLR7RZaJwGTsPNtLYPBUBqPYVW7cjogtFJdVwA9wyV2IeNE
h/MNVN0LOQ1K4AOVhiOYC5h4bpqhV0Bkjo9AudsIe8sV9xN2R5AaSkPvT4kc8Ce8
RMn0Vat8TK0fqaJIzeMmaCsJkPLGtXIkCb51BaNo+fFAXSyYKkrRrT8fTKDgRZOy
sDCoAadrGcoGCeu/1gcugV95fMPVPbg6hJEof/sR0kfOmWsXSP7TA2J3kuZfTg7w
A2+stEu41Zxpjy7QqVaxB9AiExSbBRaXJksbCeaFPYvtdPq1W4z8aMTF3WH4lrG3
t9qAGIol97LQnn29a+y5jE1KcJFWrJXOTULSKnKJskU/K/59aUKy88tnBPpg+Qgp
7UcgZKT8hJ8A7HrcZXhH55/zXwEyUnW87ac1uqhWs7z3B18/kQ/wqa2F1H3EQYw7
MUNVn1AU3EPFz7SpA/eJ6RToSl94JGukcNhV+E63BMg2DxV2eG3A6Dn6f2KxXuio
SBa9exrx5xFVZ48MGjSqOCjMgOuDNqQAs8fzIrJxm7XvGrUdFeTCaAlpgYaT68KJ
LPlp2r5L1KFp7ka9qenAgYxPn6egNzRef8d/JzUMdSC/53LohPNlMQMN8lZNOiL9
jdAyoBaupMKFJdaUfZIsVn97l80/eeCMQz1Prd3ELVdhqHVM5grvfozpZvMT/OYR
EHSkgQEVKIansSYYagzYuGJ+7c2Ka6AORrOOzjiIx1oLGw/IRtqFIX2terbMadWl
VUh7BeQOTMlZIWUhs/26iFoGs//tKrltj+Bs7g22l96c5VIpSHcHl0NdmHrdEe2V
1IinFyGZFwIkOvMqf4YA59BxfloxhdlLZvLJBUH+A9isYp43DrVVHO6uIymO2h+D
5kwHabxdjvId1rTnzS3i354d0OEE8q3b1qcQs79YufFlX6OSS2PSXthJh5UvZIey
+PG9+TT5o/DG40v3uE0KwZ0nhExryXHtTm2SwG4nEPvY3wo+J4FbP2P/oVqml5Jq
5Crr5Ll7FqErTQoaul6Ag08ohzJ3ad4bq1VdBKpS5zIjuqDbNthFdXNU7iXhS7Xt
EHmhO8Z5mNMjnxK4nD124yMncwzn6ApUXeSkuPPlSGwhOac+5pX62iscH3llg425
JvvEitGas7jmU6JqmYPJBpy0NRcfXSyMwepqPIVNxD18LM4Hph3RjY1LUk7JMdXR
yI5mnoOxHpt/7ABIe8YNoerHX5KDboy2LtqvqtvmuZj5sN3SxfQYP5ZsQcZ7ePUB
HynFfaChKiY+hkBFICguJ5b1FsHstqWDtU4wFanITgfjMw1c0aNEYNBpKWpZbW2f
BDbOQZNp6i+FqWGMzwrYn+76LEu6OsLRze1r1SJ+KNHieOLRFE4bBUXw6EpOr5CJ
+RlxhkbsKOir2c7zXQjUWhbs0IEYg2L0yUTgYy7gQ0OO8v/sB2a3vYF11Dmf86tz
8FSY9b5eZQvyqRDADUvREpdmZ7P6SybysQByCeT170uPN3k/g29FSddTqwNSuJUq
MtoYkA4hu0k1EI3fRlw4O++MEGAu8vEW9lVM7kxL0AS8ViUuX481MWOgcrZ/sUGk
eN6EYA+2AIPxbEFnf6SwswJkaW1FPN27FpDBx07w9ehKixrbWFY5K3MSLtgHDEha
XXj4KGbLOoZ2uFE7LyE5sqKzAOJr5Ywli/Mvi5cQbmhfvKV0Zllxo0/An7+nin7T
rX/6yyijt0d9vGJrwRJrIBUu7DgLm6uvqUpf50uOee0SA5VArQWmwFTmKR2u1L2h
NFjH9q5Rlfh2xMxnUDeDI07zTiSgrix0u/kwktfnT7wvsuZhovK4ZuVIkktaTQpz
KBxoCQTVm2DecH3zs+1zDPurt2aYutt1Q2PZ0CokKioeSy+wL16sH5vLT6PT9w+h
6zRhDBVmrRg+yy7z4bjB+5sPkqHxOvHtvU7G5aPYY0+JoRXZm7110pBhdoLzyC7T
1Qptg5lW1nTdaezB18pWK0L2qOz75gN21ZdI3BXJfcOJb5l+G/E2ctgZ5u6PCvjy
5OsHgNA9oBAiL/u1WShns3wFYHQLKgWxJvNv/bR6ATneNdqYNk955IuX4JZ2bytJ
oqK496bMdZtyYwVyFjDjlVAf5QCZUO+LWleWBFVY2Ol1DctTwuGGu0qeje8HbSSY
9/govqYQTooYF6E0jlPvkaKUiDYlb1rnDCP6Hi43q5/ZISoo+piOCdoI32kHM04A
LRi9TBtGI9Zy63AJQF/yVZMDD7GXav7u7TsqdTFnOYjS9208ruBDxdWjgNPOY6/B
UcXZeAVC0kIFAmJuFZSZq4X/9QqBeRjZ/B+BWyp/JVxlO6J+oXresDY4cCIL+Qx/
OyGRORb/PNZM1bHjoov1+o8Fzq92VIvOiKbG1rUTfkJ6bjto6bEKTChaPmk+eAC2
H49n9t5EXGjN78klk4tu630bOPUQ3ZgnWtBd+GfStWF835HybH0Q3WY92gH3Z5WH
xAQ8LlaRzlon3efEGzvDI1/OCHUurZYxwE89TjtV8Gz6YdkDTxDx5VnjF+q1x2oj
ClCCfgFY3DBit1DTPnuuvt7e65pVUv/4MpaotkAWj4st/4P4JHteAKIRyUTNl294
w2OuMhBd4M4yRIuke9hdCJdl3uoDdzc+bEDoMgjl3ZBqHy7RnpJGPe8YmvuXBGls
NPXbxCMH3KbCS1miDhhCs/LVcRGpmC1UUmfOYNFHiNaNVM4jYzqtKSuH0WAWi16O
0OygnCGw5ukvINMr7jmDAjHb/nubavPtYWvQvGEOgNEp33++tPUOWtGPLoOWxiC8
SQo4ALFvHyXEY8FcXuhksHQBoH/Sk+0T1oELFv0jliRqL6Ftt9WK5DhNkbxWOpEg
Ldd3/MNypERfObD11cus9ClXeRxdJZcnlPo+m95NnmvQlf8g3EK4fot+RhQItSxM
Vdf8xEqwC6TxDj8w8W9uspcdFd87tNROSGnQR0bmCIiCOH7ld30ORI7gHyJMNywk
eJ9Bbjx47AIVZ4F61a2kxmhDh9el+/fW5HEWix878c3gddzqYNct1VB7GQQXFIdb
rKNQDVxeYIj7K9B+CqftafD/MNrylFPpsT1et+NSXTlT6k/jzYb/GcZ4lyl/Icjq
i7NS3OBSHhc96LjyncaxTrlSsN+7BioW0paNQXpgjnpooXFq+gFkIjt0+GMehDt5
KE7Pk+UOF083g3ChboTy+HhQvZ0KLSOFKngbNAp7j8iSdhcjkqTS9ap68UAg8pRn
GaRs/3lZbnNR/S+E9WrsJ+LxZN2WfuStGL047ww7BY+DAIRuR+ljZ0Ro3c7xswyt
xBYLOJX9yNkUFpq+w/KSsugVy+H5ulYMszDAoh9cyoeRvXQJt/8FMOytEY6XiBCy
KdBZOizsz5abGDeZwBeGcD1t/6UWsaAphCvEy32vlnGiqNxLUNA9SvkPPWlQgnTo
I33iGu3M+Rz1kt2dRpg1ZkR8EQ0Q3DUOgoNjUtjGzVqeWV0vC76LY8Czu+I08gqv
Owsx08z5ldPStheeHr6D54BYBT54jFRAb4CXcW6zmvw2Fd3s6uKzCrX3azDSDt8+
SskrGoapoJzjt5x3/1QGkBSMt8OPMJhXuyuERt2manlEkSfQY7LigkDIryQoPql5
fBljeGGJtj59b0uvQ4NsN2UAFViF+9c5QPXB1OQ2fp7DBKdsLWCgQnpYx/TutTpa
Hlr5y6/OuOZy2r0SnjwwiXBx8JmpmJlpCdbn0i3D1jOgXuqYzUj8AM9r4IVW1cTV
io6Zk3ZOT26Fqg0p2f2XAzXBcATSzdkEXspJxEF/MCk5d1WU2ms9xsJxLtlKg+h5
c3xFbKnqUCAJ/d7fOPgW0TxKXt9Y9ESm5kQ+GvVbnbQ+78TRgT7HQPPlXGQjSOfc
Fcvd+yf0posYTYaJPP5IiOT0/vgQ5nt9Z1sLoPsQZuRRyGRUwuovJHMP2Rr1iGRH
0DIophzE5vvvdplPKxNaNcxJx6WkDKs9akIYe2UsbJCo4FXXBypJBrS1JA/TkrVA
05EDGZR7QYwE8Katoif6h26hqH/Nrsa7/48i8eVoBKhmE6tQlBEoxUGfujM1tF5m
UUeO6D2Q2VJs2yhaYNcMJKTJTBbZJUmLTxYNi5g77z14knxIGjIyMByf3RjFbdtj
W5oHr7x65xALnwzsWqvZBQYS/V11p91TXXMhNd+rG9p1c/5A30LZpSO15Hwo8sfr
SK76i2F8RKYcVcDS0bbIlX927AYl68UtGX2l2Q87FfaQ3SF7I9FAtJl+b4TW41n3
0gp+UPwNubejubscG2TYMcyY8bAZ0lzJP47jJ/aMGKvLMvlQVIapL3jYajrHE6al
G8Vf8ajxRLUsYD5b/7QeDwh0SVHxNh+Y6iCrRx7YZfmN4tmdQ4o0RKfOfv2REOah
wSc9yN0zKvITr4RXC8s4wRkJEWacHfYvLg2w1zJkuKj7FiiWxgSiAUoTYtuDUj/E
zLXKW6aQjRhDnZTa4SInBkh78l/yWPbPOEmtlAAOU7AtB8sEX33A8LoA0jrK95ck
Yqw2zOm5HMdXLXd0Dh36lQRK9LjpWDJU8E+jB9tcgBs9AaQlu17EeG6v8sfr8IXA
VP2Hr3hSqUhSJhkSaVCVEW6tPfhyeMcsH0n5GZbT182/ENU5h8qhrThZFLvKwk36
dMb+TZSlNItLD+1nRzes6nuY6LO8nJS/icem58a9zAY3d5OkPd0hjaEOkyHjhlB+
Cp4hvmwyDNgDwOt3hwhuhcYP2hpqUc2TGeIQLdnaOs+dApAxeadTq7qjIxytZrMU
LHBwd6KfzlOSEi+iwhOPTEyz9/wHI7DXm7divDICYKPUim7i8FyCSrPw+okUBO+a
fYiWq7I5eae4qSIYUAQQXgTYXphABQba5oBPW3HXpeBB2afCSvmWbBxy6PjZiRyE
5egQD7Mb/13jWwymiUqszyEDdTtrOOKHeLaVagHG/dqfPo8HppNLMNuP831PVj1l
ZiM1gSrKvNEHqSQDlNbX6eumJQiTz1y8MHD2ouaOrszfZfmk2NAFAKe+6Grm7QVI
EbGq6GcaW11yA5dmMuuwldgKVafNHPPcVKO85ABM4hNIlPES1v2bko/W+8HWVba1
9afP0REKy5T462N95LcyxKW0Yx3fkdn0V5+YQq952meSqcY5kv3+svNw4EJIYkFi
ZGfUKEsbLXO5u6G8xQc3F+/BcXjRbPAJma+RVcvcPmZ5JoLzq8WMUxztZ/aZWe6x
v/83eNSN/Ztwpo+d10P+YEArR072kiBjjE1guijP0bcuIlYDFeWP4bsEHTCqwkFr
a4Q80/QqrXP82Dgmv4YggILr+5pUGu4gSfs+NV21/2+1Zu6Td7PBtkUejoNYd7Ir
xkbgPg4fqdZaak8zT8dPcr1a1eeqYCKB/rmQd/3jUt57XBNRQtlhkK3LVv1gTBi8
7jDGI+zDfcGLTXpmmfHzEyx9pafZ2EGZiyXfIav1lYsKEG1J60Knm9mipnqXQYia
XMxUWVAfTKNtRiy/OiRkyfHMpjgJAEDiC/d6IDxqW1iP4rpTMDvLthln7A2i5inZ
3mlcjqWQI6B/mRXNLprRi0EP3dXahWiDrVGLLoaCB9ZV2MYl4t2CBlcrM8MPjUJY
M7PvnkBRVqMFeVoG4z139I7XVY7rRY1B8HiNqDPrGPILNMghBxJqXwXfIsu0FgYU
SN956HNhBWTiPlfcbqTKUTjP6VDpffVw5ce0gljiVt49ILU20UAybBzuZAVCx1xu
RbkET945SVqDTfhMINraur5wirZD6lR2uTmEIqgIiWuP/ezZrZ7sOff7StUdK16W
/snDtsmsk7ikwam3Q1Jh7BGJpIQuf1VzyngUzTa2oFsZdyqwgNkb/jv7dM+EpTcU
dN+HVVDXMWGwfJn/URFHuQVchHL/Jr+sr8k1yGx9HXtyg6jdmFotkUttOT43dAvE
+V0AQHljrw+Ywhf799jsb0XX1Bky0E1rK+Zbj1HLDkT9tNtMYg5NazYoNp5EmbdS
aZUsve7ATenZTq/e2BHXIDM8iyD3Is+QGhy8EVfu5AT4dKp2ZdZJVIHYqH2BEOUb
A5LGS1YYAbkdT1r5fDw1C9mEboji6m5SELqdrqtChHn/Dzs0Iei33FtRP6DbL0Jd
apD5mZUJGkcbljPL57WKXLREs5jn1cV51a7EquypQsj/zR8A5DoFEV1IhaCi1Bvv
qepNuOjMACSs0g/gPhjGQXY3RYQjZsX3xF37ie5RSkuiRr7ZI4NYXbCXxFLMnzvP
kK98cnq43VoX9AtydSz4/nMW/cv12C+1Xpcfo4YmntTbBnfPMqxjrbxH14/y/KJO
Q7ygnBgS+ToJcl88jSOJcrS9i/iCX/1gY9MyKf3fv+Ne6sbvYoFfvWw5DzsQt9DJ
87EfDWKCMYnlLD7gsb8hcnyHNjUGoCqHYa32vb+SuF48e2yG05ESVZxlALs0R2/o
T95PrzlfroPKwVjfw7t3IDsKdt5CdOphzvKgjbFOnrgcn+SeYDDzVGKm1ZwB2HB/
cC446C3PStypyKOBugShCbYgecuz9iKz1kMllwjXKeMXPulRcpExNeSHcQ5tmDCj
ozYVLmJlbfsHVLLzXXUAVRIoT6CRmy0aKZipVi273Um5xi1MH2hlfdHgkxQELsUJ
dXKMXxje/1buKJyz+ME2CD5XnB50vDtkiBI7rMfiYy5pyUFd5xoezd0ZBanGXBhK
SOUp8Dr7UMhjkjFGuwQfXpewD3hCNJkecjFNgi0yJl7JkcbpudsJVOEafeAHw0M7
/n1rruGhmwwZeAEj3O1J020hEzE5JTKdHVibpqPMZUVoibIeDW/Wjt1AzIV+II70
XmaTqG9AVU0pp2nPQQ7b6gsX1ITmDFh6mSnZC3ecHfjnXS9r5aly7K/6W9F57Xsl
C5lby8CI3uWN7OB9KXMq+SvOYUfhHoJ1WEn8qOLsyk5FJL1V9tQSvymuM5/G9sKo
h6V4naiF5oyvCaKMk02tFODn7aqx7LgJ6Cdxd/Hcq18UOCjljwvA1dqyxP+B9cFi
+0uCi+9eILZUytb6rTkwGYTxeZdotaO0s0df9EZVP0iTwlNevwriUIY7dwYlNebe
7i8EgMvSdfpjaf3UDi8hNNx/XkQIgMaVJVlprXkF8z1padI3+fMYhJ6yZrxEc9Mr
Q+7qimE33mjPcBHpnci2Tv317foJXQlXcApmFLwDREQNwdUTP9luALkjABIw6awK
eaXKIii/FYQGg7vHj8pe7VAcmWPVKLxgNuGvTzn9O0FSkJUJgmhas5JHfq0GTw+4
SVcan3Geoe1pQOav+7kK8WlXPfo8SLtz5A9mQv15AghX0b8BItUNdLYEWSJxv8HV
edanakyB7jr6x9uXeoQnwhkbyl89F49r1I9e1UBlvB1F76fDomcE8fpe5C/MJoTu
Xxj56WhwyqqnEQTmq59dafhAKWQHl0tMoyB1HwGI8VTCJln+xUMR6Kb6excfHGtU
+rotBqmv0VDE43zh/nEQqAKyx0X7hCp+HyfbhlN5kV6+XJ0D/EXa9OyXhSCD3hDi
I3727TY9ghTfTDSlHuoXz2SklOCl00zbuInqB5aZqNisL4QAz+psnlf/Dyx+wEOI
/gRFt0n2fF5t7HwGWAmh8rwyMt0eg1s7AWKFAItyShop7RhlRW4eJK+IXfhf1hyl
Sy4tPrLP6413uREAcJp1eUI/DIzyN8E+GL11gnpQa+nJuAf/1u/Y/JU6u+M469EP
rqzXv6IwAJu0O/MG4K3DuZZgJM059eFH+dtyBO9GHttsRZy3PLW14//BVPmJDjOC
WMXNVhzlsTAVRmL6qrblCVWyWS4p/FxjDIoOalFLPpP+4b9KS+q5XWsi3baRWB/R
vCC6hN6G1pdOEMF8nRPg6sGSq30dBiBJiHLISnMIdnV1qNu9Qz3mTZjek4q3dtAT
PYW/2SbIFdT6QTHSWc8tci9f/6mBgj1YEfBmL/I4s3UK4r0fAzi5fd+Ht7UYPaBf
qsL/tBKzlb7zX+gFU0TWO0DnpkEjN6EQjvN8WscaAcpLt6nGDYEMKTSYs+CjegBn
s239QVf3+Or4ICEnaQYJvrEMwVMUGGVRATys7wM09VzGyPJBVi6FSk0Byg7rygMM
en6Rs8ElSJToA2WSEwSeljXC7FQHlYjKZJj2JMvfsYzlmTgAC6YXWatrmXIKb5Op
HGJOjrdrgrKwIrObVH3G8w2zGLBMWPxkY0xvITPcI4/xfh9EGo/ZydGws2VuBBhA
r+KQFHzmY1To60ZaV91Ru020fGqrn1lmllj9VtM2caSiu4C/8nk4nsr7M7a/CTb0
iIhD5hVzg4TDoWqvQXpuVQZjh18uU9O/R6hn3QyFYRxWPrtNQHnDhA2RNa3VnlzA
VNM1DfZ6ooClautRUPHUrEmks5nCM1/mK7FzxCVPEeK5l9sizwPzMGBcnSTEgece
2D3ZN0rimXmNwpIFjxx/EoP2bAaPMmDhWcpeD3arp1IjNdhEOC8w4pPaEeWnp0Cc
1EXLBpxAT2+dPhFWU9GZ7b0a2nfqiTdcbs461udcZBwC+pDRxWPfV96MOlJAvg4A
5kJAXMflJ1wBEVQA+LQ6oYkuItOe+HxybMvSB9x52BniZK3V539O35WPHaMOPnei
u807Nnp2NQOYPn8PeTzLIKQ8ZQ4W2d4HmCrhd/ZVrE7a6ces3G+HhzwLoCMxZJ/z
6RUeQvLohmLavx8VTrVhiQVIShOwKBMTfMNQfowvzy4UNZmiO+0MmRicNPdAUypb
crCMVkbgBlRoN0hP0FXmoWUJdzSPgF4AwPbcuj54AShzXM5J9sYauYzhU2Zr6/Ge
MbBHNaKO/uIDjt5YYODcGb/4MQ5RguD34cLTNi9dtl+ez+ZbOx6nTSfpfo/Kn91q
tpYOJYGVfhjermqntTc8nIu7K4ipt6E+CaLTpi7s4h/RxpN/WPG8NDHJWerO4pth
iTKFLR8l7VxQ/oawrQlZ+Z+PCblQYI7mvWXmKU0/hYNNOdGKF51yMlm/Cd4AgrzD
gGH7US0/poyWiBzBcCx4HUcrftW/YVuCQXZ5/wNZXHmUMlMup0a7tT3O0aGBhbU9
f9a4nBSgE+4D2K/NKblmeVWbjZZxR/6BtEPazXjxS+xcJ5YbziLfGMNbZSeod5Q6
EBoilRDsMdjoOUtryXZTVnVmDtEXjc7UlW7lRvbdDbLbUvqAGjeYT2gO0bmpmUqk
anbdDb6J/N3K012/nLSdNXGq4kGlNsxOVov7PACe2wV2V93O68HtkN0GMTDGWM2D
KkB92inYbgLrkYkwNCTJlAbjE4FIHEtbCoBkYu0sphx7x+9ufcM4NaNZtPZKP7G4
XmlQ0DZVUo8FHvxupPed7ZXNKeWU89gcCxzb+yoPt91339tzG7yoO6tg2eKPOOyx
lKZLv7TUBxq63Dz+zVcSXMEQKfd30ACPXy/scFNQaHZS8kSQa2Wyrjg5GRNQrt3j
HSbGKdbJIJwWEC8XZu6VbhOKLcyTQXPrCgkRPBmHNKVyQ2h5ZQ39RsiQQcSqdEtL
QWZbpwra+i5llZkdLhrNmiis4U8ByS0oFX6gXCz0MvBTlTKsHK8QXA9ACxvAoZAP
K77HhQZ81aAeXwKRc8pNACAlJk5w2kvYJsrWbgJRKRQBRTPbfGTDCzmMFOWnHkzE
l+6f+ofaf2KBpuWgbhgqxi5vuocdUGgRHDM4HkMN+CMrrXCcUCHSMGjRgqIu8E6F
7K+OCP4Kk4p/MfAsoEhcJTn8e7TJpwxub6JkcqfPPbg/WnDowE7Fe4gNqDZgyMPT
OHf/jdNvHnvI+ObxiDHI/e6ewesHfzMSXMgcy7O1PexIUVu6GDTWoPzQrZ+PEM+7
u5ignjzaAGoPyH0r8Fu02NzalxuzOylawnaPgVZjOkrDGAFPImJfuxPfPZ3LXMsN
HS3y9xcjvxh+CvnEtGsAXkTn7wixqcRQnvsiSFzoS1KUsyK1M03il4vlA6RcNlkZ
X9RwRdkC8aea62+RvJjsEIxh3Dvml1/G/7E8oiWusO6DiVXgz/ZwSorYOL6fhN+9
MB5X8iqeX/0cAI8c+2D8ljkfLVrkK3J6BnA78+nfaAFkOzft0+xJYWY4gfnZII6k
wJZ7uf9ds5JsK7x8EfJcZ0zVRbf23SqJj9PVOKo49IcKpRUDmEwskTtQnyK5Xkkn
9icRe4uINuuUvya7uwk8mzPc1pqccbGh+FXR6hEkmBvxfgPUul3mfjmFv7AIBbRc
/jEs2J3lTdffDDfF7SroXPsYMRe4iTNN1LY6bugW1U8pVfphveXNdxfh9XMs/RI9
rleI1L1NWPfpRPtemxqCKU+1Gjg9iJED/OnWOL+cCpNp9orLjFOCqFKGGkYma+RJ
xfcFNWYiOy/SQ2Ava5FaYtMXZvdJEHgxK8G+w0WvEdZeZ3ELN+/ogC8LHydcm+xl
2SpBPJiirPUnw+8t0H4131WaZIxYVoSCZMtfmUUUokaLryBCi9kJYlYG7g6fMk/U
G7WanlCCwwiM8S5u5AVqUC1aVTGiltcKQad97Ue/gOb4evpxApJrSQW9hDPoco5p
OBPD4BPOCWcv3+orih9fLt+WV1TeptqyQvgYvjVvQ0VwukXCkiFE2Ujcv2BQg4IU
/fkRrBcUx2YavWRdUDxQ3aMQZn9A32xtJTIE0Q68WPCRfhyVPV5sywajDdpLd5ad
TaXA7Fsc227cqdb7YtQgSfBG6HlsTZrDvWcFrJJS9yY6thw/IT5Cl7zqh5LqqZyl
ApJ34nWNf38btJd/oa5GXrUULVchDUFwH+e5SejnZJpGPrl9/bEGnMc4AJWmBrTp
jT5hH+qg1RARwwKE0c7xxaSd07ex6kAYprM+moNALbBCermMGhRiN7QAQdtBpepG
Z6ewlq5ErqADOpF6wwrpZsWmviBGg1pFSrBICqxVXst+juN9DLNd0HWGr4eIhZhR
lK8RDngaYSPm0i6UCJkwF9ZrFOQ3Oaey47hdxTOG6it6fasYN5el6GXO8ZvXliem
47qvWAAOTX8b0H+XpODrU/awkTJ3VWIholpryKSceykUHhgpUzGLIt73EReUVk6L
1AWQTNbeOcZ+4hbsxolqd4+FfPs9o59PMruF4AdGGC7pcogakWva4SF7YiyQVhHm
F1vS6C3/7e11Z6piQW+hHFNOPv7dQpzyjXgCcuhwxHqtt7wNHsxkZlKPJIGq/yWm
9wzGJB5r4MYCtrU4nGXqUeCo633Y3If4xRZrUb41YHJYnDxfG/PMDKFaBVis5DX9
R2BMofCdpddqhcIfxnNcSacUNCxf8Wwd8xXwm2Zn2Qk/2pQqWvgFxbU0qNUUQbK8
SU8Deu7BdvTItpaMdR2h4la1S9WANVAByGN/zHqPRMt4/OvGftwkA5kl97GCU5C8
JsIZCg1tws0Lq7voOGV0E01qacHu91z1VSJNeJtNK9M5ML7kSjsYZ4knG2cuGve8
MHZH5S+jvPEkpQDKowoPWn6qbLQzvXrt44mC5Gak2oiPrUQ7+VvqvGV8GOzwxORg
4gGO0OeIm1PHBStIE3eNlTnTaMCicMuDcAWXI5aSSzKvlaKn9uyMgylNKGtpXq7G
b2W6CbvrZnNkh85P9ES+B4OFXxUyWsyHCkupz3my6PVNVzfBtf5PO/6xTxUs/q9M
7JfTvqORKoOTODZPb7DiopxLqQd1br+CEitWdTiOT9WncLoN+gGys6jdfbvAKXjO
yUGrLJ3RlK/su/PSQoZKUEFDm5Ue7QT3h2C2gUjJOTVDLn7khkS2tJJ84lTqIneB
qH4gQE8E2hRQqYPB42xOoa13hbl7u/XQZ7zsOQJM5sKeMohr5O9ZgDrkvrkn0xeV
xqTySVFYoOOyzbVlERii9i5NaL0jwKQRMDG6v+ixv+mxzrriTKBMSalecmND6hKy
5DVwjI8YrFsV4zw/ZKyGUIFdaLPq89vGYUj4jf1IZDSOMwzUDKA5J9pA9anACVnG
vMyEiNLufa6d1ncCIsP7RafgyLmmyGnAOB6bdyTRljWSe/XIUU6edmLAvZDXeO3P
nKPONJMgXI2BLIkqtZ7isoMKsB6E9uYimI6SPfx4gk9UW+8F/shK1MO07I1drFc2
BdSmO3agx0DR14plouKZLOmM1mGw0dD75PxaDtP/e6dvvXNq8FB5O3dYlHzJ2g4K
NWzPjcv5RbBNZ/FKwhtl4/fcoJti3V49z5Uv0tMlrqLOZ55KNdG1zZcchhbFqYGp
HkIJORpxJT/I4asJdFKCl3j4sw/DueLToDRRaR3xoVDeblDQspzEC95yPC7Yh+jf
zgR90OTBHzMHV7w4+UfX+baEV8/Hyq46FtDVe5cUcneIhd6ng6U9GHnGzDq5pZrl
vlI5ht0IUN1Hjt8jVSFGPSttTRU9Lid+p995mQqMAGHah5r5nTKUl37c0wJA1b0C
ZJaxVJds38PDa+T8TIazVrfYSZzsMDI6EiWpazMHCJd6mawT/2CIrNPGrie2Y6Rx
tOnCiChSMLChuGCA00Sx9zC3MjFoSBQdWR5ylNXVGwKKeYV/DGNuNIxvghHeJ4+A
TxK95QzZuQLuNpgBqZJQ+GM3B61Put33OyntWmKq7TmErgA6YdD89vw46EI6ozow
o06UY16ZGBKXtlbXn7600GXL4GFFMGISYAAHxRCWdcUtix4y6w4hELt8Ci51KJfq
TkAdQlYu/9CzxhpeT2VeFWPkii+Ynw2MOyTnco1zn7TDYUGfWyoR9mpEGH4LmtHy
4N1xpIKKAVJjFZKFn+GbYEQXr445w58Kc5dPFIAWi7FAjAEufvKxa9NbnWosTYNN
cYCLdh8HS52SUt1+2ER7MTwW5InU6e2gQdbM5hwpUvPMjLOkBEKSXHifHWAn7QRB
2HI3mG3rLru8bBWQ9R4As5+jsjXC04oi6xI9jxwPwGejap4drQWu5YwJuik4WR2b
k2ZmEw97hvNoE2w1Ujvu9JgACU3MvB3PAnn0D5cFXbsRiKbBpbZpvAuqDFiCAw5c
pSS8taqNpRVS22/q5UMfa1sW4u8x93L0Fq9X8m6p77jsc0fxFuBsFVxu0Y8r2UYU
YmrAkUQrSXFnSdgnNUzy76aqc/xBj7Z/AYdjjYqG2pDJ7x/jdNd06lJUqNG5QW7g
kZ3jEfWHU3NCQPaYTIG5y6bdgDSPgaiL3xFf6wkRs/QxhPrdjAh3EhDq83nO6dWi
BEkm6611kiD+pkXjQZBfDP3QVE4K3ljAxWvRSREqpf8Z+d0GyFpwQ3Vs/Q7symTG
KCLV0aFmzJs9Gl/lbj2pKPEak0on29zyGXwcvT+xFgckLffZALJc123G2s4VhSuX
UNu32rgimh18i4Qi/W/09UBjslhKmzST+WIHG6wTpEveTXCZIYWhx8/7kYtRqPfg
wumqJyQAZmW0QyGahrWhiEprkwbfVAfb+oolbABpMrzDl39s+puYU1+/YUrm6Q2K
yBhXVPgpj4x3DjGh6WPtGu+DChHvlMcqz5zuqzf7eUujFES2r/hXd5NMepScUkDB
3ztKsu+jgFm7klzHXZ2nY6mTCD8LXfRodJL+xczVfCRyZRkpmBig29aB66x6/ppK
sjBQngC8nSRwzlIExZe2Wcoiuwhp0OkUtT6mcnxjzO/9UtgTLKKJvq3s2ev27nDu
CzoIBYH1Ja3G+XaObygXjIIYaRwkPRNE3xO7rrUUAaOSTFt1DJIzWCQBzMCFv3dH
tNPAOuTv1oJrMPZPSD44pemb1S+0RjyZ6fmYram2gTIowPVFbFSi5mcNhSiY7nOa
bdZdQad3XebZTfqfOYlTU2xvGyg0fYByOTmel81YKjRkDcnoDFQs7vXuFgS45zxI
tGfUOLdT7xK7OKJEr+WtSQQ1ioy4GbuLqO87w3vRZ8NME21QC+uAFxmhGUk5zEM6
Dw6hKr4yw7yX/KtqbSLuexu3gqWvA/+U+ZZ0RuqOUh8k24iP29CzuKtmH1P/CWrV
9XuJnHk2UzxwEYtbiv3h9FQwEStrjupIXq07vvYh7C4kskT0yuZBW1BiCd8mViWk
NHXBtlMF5+rNGn24hagEEYCL/NvF6grhzlNK4MULTea/s31On9bqe5/lyvXdoY/Y
ns3kygrJVEMhO7kEnThV1rNeQXFQFsVx0LvNxdsji6ptBzKAv217zSoMj6uOnhiP
o67F+VXnuxrMuSyVVIa3B6sakrqNsloMG4lLk1jMJ6xvENxC/gplZ7h8zlKe+4fO
3lCjiD5uLbDGhU+AY60ZddAEvI6GeJO7qOKp3IXBS37lp8Z2BE4jWlLn7HGFTS8k
l9ZYoCEEovFVEC2F29StzO0zFYjHKZsUBgs3ZNNFnPixZHyA9N2kKsIqXdfCvyF1
DXpxvOOSiSViImqo2uRY6Oh4Ip0RuQbm1h3EEDyDcNyzrsHetBcGCTE5B2uNGNqd
klKymEJLFQUcPCiyKWdRiMfUZndc5KdfOThKfB73iPlRlbyo+n+BJtfP2QPVH4WQ
bijiyToZ7VBLkMFkj+NECl3y2ntQ5rHyT+YuBEyQHSS0OiXKNa/JBxKnaG3rmsxC
ebXkciu76Pxv2DiHqALECOZGoBaIG/awXG4KyzmBXSgsovy/dEPlPCtg+p1uEpgZ
SNV2H55dx5SWS61A5uLJ5MrOtQ9oWomJODTXoP3+Li/31Lq9V4b1clv8kOrM6MDi
7mA0NngDm6WgLgRXlgcCmqSaRjOLhyPoGlV2NXkAP21mH0Mp5PGu2DEpODLnlYyJ
5AuK3U3COKlhAFeyTuT0vKUBYtvcq5YIPhUcDYCWM37pdEG1ME50Bqkaiibj4xFO
qMoTUepe2B6s1qtA0MY3RvlsrTwuWcYKKJf95qkIZgFT2xxJ6kIy5SOwo0XAo1Hj
AQx1bXKC8FMcBGDhIyn1qmW3dVSTLU4EFvqD4RtND7Di+FHUwSZcr1KN98QqDQqr
MSjA2/MpubOEIs6BYFw8OEeTm1q4RuF+L2AJ0DCMncAqEaRyrfYKTfxyNpAIlTyo
s4GzYJVX4E7e5kDeTH42avyO7pJTF0QleCggJKVzn5OUFl/TsF/yB0CLIbBSC0Os
MNItbFkR7FrnXp89pLiPzw9guMXhJalI799QKQKrzSOmApoJ5g9I2OnTcC6bRdHH
j5u/Ly35XanqU5beWiQ8qyhDsCMgwwAUrBKgoDMA2AyuNPJlBxWrJQCRQ25BAfgg
zg4r1HFSy99Qlay5km5N4wOGJ0QVc2IhFZPLdnnHdCv3H9i85ivEHwnY7KVBHAE8
l9Yq9wlQSDUq52SwY6EW86gyraw14w+HAol0U0mir8JaoA3AL1NZOMzcCV16H2+d
eNK5hJJ0yeTFG/PbiRzshjU26YXdTyZH3sHVkqC1cvlMTUj78vFD78PTqlmzfton
hvM8gMNbVWmjBPzYMebBPCADz11OQimOYX2iwxO2iom1cS5749zRtqZ8tKqq/hx2
jN6iJ/qjgJqCtk458f15MyvBahIUcjHX1liGlOho+BB0qvKRCQ4sCpUWcD8gy27c
q1S4tBG7oM1Fl9Cc0SvMvd2Tk1vYTFtcKmgbSFR+zuavShlQc64+Ygs5UJd1ZANU
NYZHujWZGsM131GxI5/gBMSO3jIjB9MtiCKR6pumVHqDGXj3olXyEQZzIPOdL2Zd
ibCR5EMABCgg3mrYANEHmil5YMkwdWhrdXZCKFonbuH+/e+fo31LZAJGhUsHWrG3
HV3UoVCm0N//T0cV160zW+oNeeNgiilltHdoYEhhWrvSFzfFBHCKe9WeVNpml8E9
hyB+FiQcRDDqknBBqKjonzlcBU9mSGeB43vCW2MgaL9MCBP0AQ/jp9WcUzT2Xq8j
7cNxRqc9b5sgxRjvJ2P2BJ6m5lWbkSjur9lRkP1CXH9JqSx01WQaI3/WRCBSc3PR
f60WKOcOkLnRKPqXMGMRvzDlStaj3nfwY7QCmJ69Uif6ZuXQSyuAtp6mEdI/WfHS
ZnPMDiU705FKeUXjDAQv855ibgoOOGjjfblZntetR+cpzod7Meg8/d3/yMdzX/20
nMh6gIVGQDGMyHaHvcM3pAUft+nCGO3BxhvW+oMt2LI7K9Xoin+/DiERoI3gaghd
A8ec7y/7GmFxRdufXKkinl+iYL76ilH3UvHRzzo2PfaI9bDcIRNmYJMWBEX3xZ3M
2jhZxMD4mpZ+mxexR8iLqv8GxCGgLuOkTlWF1egnC4L033TWjUyG04NC7t9oUc5D
q8zRsubFBNrtpmLpyDH3MaBSbIX8J+bFilH48A6qBdof5OGdcn6MbEFWf9ycdYgc
BACPdvIqIdkhWy6yeJPkp6fToNvZ2TD8gNA2Y3vJ37vlrCTI88PAnJ2baY8dreIi
6vn9yXwuYtUlT7Yno18UWcnR5f+uvgwP1TUn+T/zW/3FfmtMWgQcnCNkLGz2iyZU
L0sDL6fRPSzWmi1+OBgFKROouKiFFmlrEX3RUoEhxMP98RRiCc0yhysAMnV/FJbD
VuPXIj/AFiUQGJy+w+nXZ6KDuBrKbc8i2O1oQrhXFVLHp/TGBsgm1TCKprxU5+/U
l8CklL6F/OW9+e9biW0vKCnx7VyVkqYsBPjRjIpk4FQb3aIeXv2il4nHiHIC71/M
u7JGrB1tXumAy1d1VMCD5TDrpWtoO8pLj98PNKNaIIGxlRvjuWjKqUgQEdTtXxGB
QVUfref7XBdFwJB0aCtuMPFjJ2ym5WH+iz9CzeTURf4iWSv1Q5dlk3RXIgx8KDdB
+eiAH3XF4/fnLefAasbBWGccUdifUNRVEleDOyxsRZV2hEZpUxMDyCHeHLIGQyK9
0N3a/ZE6Uzkx1Ia2PQCNQjesontt2CMLrYvzV/S+x0mxyhk23BR3czqG9EY5A68u
XBMeFjn9mac15iLOqabeb4UOc0z+8G/xil3JukAa7g9qlYb9zgZWCibXTDn7Vo8B
QTpZfFK599BIqwWomTkRjmuAT5KKsuxBBDloUKmFYtWjaBig8x/GQvlaE2pbO04g
95rEFJvWiGMv3WsBENPbN3X6NR7V/diWdQkpGnY4nJPKJGI/MkDOyoNbNnn9gBV8
9SxHj4rHrow3coynvAJheFFxa3pyXWp8WOOXi3l8U3HBU31yqjHGF9MdXkzFn0qI
yTftnOEXpaCLhiVQgHAXZBpJ35OrLBTotiPbghML1xU/b1Fyp1Lv5VZW6O4jDldK
N3oKNCRida3kZ+yYbOS1rbRjJJS0Mu7aBxI59R4WSF4rK2veX1dj3FWgsNI8gQ15
JE9ImefnvbsSEtCfnGOdo9snd3pcn2brHHPyEvKiEsj2XMjfCu6hQnNOynaUG5JM
a46D6vA+Oe+EZE2woNs8E4fnZEugrTQW5EOT9PrtGOXQdc8BWLmdHZ7cEEPzu7wN
gbSTxkcPZ2sFg5bRIw373HV3mk2wEUUkcfUOrd9Q/4YSeUkTZtIlm9qHh4koJiKL
wECF7pahi8lirwqUx0Smcf55N4Rs+XJcUhtjxjZn8vL7nricOE3T9bMo8adYu914
wPiZK5nMIzbCBmgyHFKBS9WNzXEsFgKqLrmwY9+zwtfxoCCf/1FF6wNuxuLdyI/l
cwCxP9GpzzV1pXV/zDKFxdBsyChtk8iHIDqnNOp26n1FBmTIjRnaN4FO1MZrNbcv
oaEwEaDoFjWqTLLuqVK1/KknV43mCRMTEchXheaXAg7Niq7hhwh14drGwsjddJXp
6DrBxZZAt+ULHFsoASuv0iwmiMjvx+iyGbQizZvpYBJDrl6biyxj79Lc83n9QBEL
ZV1Kz/Tu0MOH5WGNJzQ/1lCnpkHqFuV/c8v2jUPGnKU5WDnNv6GDdqL8NNyUMvsl
T7RU3KYwAecz4y62bj/4orj5qVW1YTxYkF/KARp6SAC3SXOb8Jw5ZFfxs0p5t2vH
Z6qGF+DYZpsmE2g3uH2+cHZjnLM2CgD1lT4Cd1GFrSV0Wr1YPgHYx+hjo6Ux3shu
rkG81Vfr7MOHmW3u0sTerYP/tXuyROMkgonwsXjUnP7bs4aFQlli1Yl+w2oGAYi7
AtebFXstgX37mJ+W8VPKojhWXzguT4v75gIY2tTtRhBKM6xX7etQoQ/PZXZ7nrjS
biz9byjVJK+6U721GemNjqxATv5WPKwsMav+9OBNhfa93DyV/6KqI7/UZGPronoP
Hx4nLmjrnjbexJuWnQjmGYPvYAd8X7etfR/ecNDb38X6JJbuDPBST7hTRaI2cK3f
lyQ2yO07mTxDKHSPZqBBcVkDW5U81Dcl0maXia7J6D0lURFhEYaWsih9IH5pcNAL
gylxAckRfqwu34wZoeH9CR6dP1/hzc2dKKplOwJUfaRCjkTsws62jjshlecRhL8G
aZl/LDwG0g13LtVM9UUX3FhFlz+4zNsK+xcQB9eoKL/aBOop9S6HIXa8164eBwG6
FNniT5SDHubgDPiAY1j1Kcyr/lP7QAVZy48ebvcUr+w3fIVbfdL1OBHX33hqntOI
Hg4pCfEVW+m3fbZaUPJafvkM1QGjRl/Qbejqpi6RpoSwCkIfKh6Z+Ui8tWmxUuDC
BoUPj9j0PqFKaNh1QhgrRI1C5L6tLvH3IaxMmlNoB6/v1xIKqO6RmhjABVsJWMGF
rw3uWoe0L4TF4sdHdWyz4ZDVb0Gkg7p9nbLBMyq798jJW8m9kBgFkrQ5KeoMlJMq
SHlxCfxXrzl85Yg5jHoKHnBWN9+S/rZYOhA8GmGCNnMxhvA2RP/bYWA0GsxAVvT8
XWXYFrIYNcj1OCbJ0ao89yZ/4bkASryMaPIS1Yv60cz+KT9l026/B8UfGMXy25ub
KS/KTLyHUBMbNwzyvPi0QLVEqE85eURUrSkeJ5gG/T2vwKYxQntgko0DQ5dpFHLc
CBD/rrAn41f0vBmAuMciCjcnRBbV0vak8AcRT0sVBnQqb6zxObHuiceZsP2p+UqA
7Num5T5B8+VxOeOz8xeNiInVmFHctgeKvVsldB7fGrC0+TxWHZjWgf4uPGfIhEIN
lNeULqUIXqKm2OFlKHwv/VPH0JaOGGeTbM2ffiEmRBIYpNlp3cHm3idQBKCy2XkL
nU5m/sQnF5wUBt+0JAKsBU0LV59izw46cHnwhAIh2iCmiqjV8YDiDgB60TYdfGA3
D+LeFhEu/MgdG+Rc8mJ2xxFzMlRf2ftJs2AieCxxFzokUyt6jixGgehed+QKTo7l
RPpwphxYhC2ZL5yLinXj5YC3ausUcZvvNZ/cqNhO7bHSWEs/s9oWrsudw81Fhys1
76GSrDp7ni6TRqHeoiIs+7WwIn4A0WoDGHnpDo1SYLc85gj02hZUUmPs9K67N0+A
AtoFy61gQzzpDK5DoP2MqPASqmyTC1zYhBKIz2xz4QyVUTzx3Cib7y6NPehvxJqs
uERgU0QsaorMeMRkcFc5D5sneuVGy6Hh3qmHGQ78KU25/vq7bwnn4Yym0oVsvlvn
lRyqsftkUlF5vMe/auOOjNQq4bIME87NgJ4Xma5FqF7m0auBr/0E7ctMXjnE3ke0
bVfUQGGCdbzAQfXXIlTJZ3VQ3aMbu7BkHskMDoxHk3OXBBCPlWCg7eo3c5wUpU/D
F0DWqakodXSGzA4iKuGtuquCS8kXeT2PtujNBYPyil3+2M5EpNDbHrCLl6yo4vp5
pf2xniFdMn+KRRAurV1rPkVjfuYjyXYGwwfbHIczLR40+qlWe9zRBcHUEZYvxLR/
2oTmunaW+o3L0PUbl9ONC55mbhLUE5Hk2W88pX16zX7hjgtuARi3JPB95cnvr64n
exuaCZbJ9gYKqrDy+47m1KLCNUk+j1AQMzjc/kSlVLoybtKVrw26lyqmL/6JfG68
g8v8hRZfBNLhlNkdK4TsFXefrH8xueHaN7PAX9QG18NnF43sRqYlz6IwHomNqm/e
SK+47xciHW0eLt9knuw3qMLK4fGfF1xwyv0Ki0hcwR7ciHQC1UhUpws26IBwDInF
mnbhnVSGroUqdVbQ/NxSJfORifggSTJYx+hxtSjmY7GEdwH+Q2Fn/tgAJJlU/V+i
wXMhfFNHhaw5UJz7WnchnpNUuT3KwtQVHN1+0tT67p2/mXsGtrNsIBp2AW1MD3un
WZHamPxBDxCilqyLlnab5ifZeippzoALCiw2Kv5va0iGY+5nf1VXoMnotRdmiQJC
sEqkIjtxDPDEYCfjsC72IlOfjBwcWYefUqU3jW5rgi3JDGMK8Xc9vcH2Wcnm9DX3
XEkekfUTpx6b0Yf+yUQy5ViYq8kgHua+KZbn76eF3imTMqB4StYM5CYl5ItuKRdG
xvQPJERo9aQ1udia7hYfy91pcK3maskbn8wk9j3+ufp/ISYnidSptGdW2r+AgnKh
SENd1ni2NH3GY6N67aet6/K66lB3qber1HGwYFcMEix2dWxMWx1RVKQWWwEaTVC/
gfp+JT4GqGqa4XR50vpvwv3G18gpAgynZls8oeRFxB3Kyg9q4SIw7grz6PtBtExD
dQso3tzNTPrxklx6QQbgYDwUox7myRAJJirPhSUVq9JqIHqMVxJ7can0BNGqByI+
it+ilu1OaeXhSYgY+CnUscz+WkKD0XgArebIzPLvDKoqVggLjCvylgvI1uJf7WEq
GgTuAmjeNmvEeWqGJiB9qS7z8XYT6Y7w5T7Y0GdSRr20lT2A/m0WBjqV8e4SuO4Y
zTY2wmqjdvQRBawLP8Cn+BGyPo+5BeZKQ2SeAkkMbZaARWOevS7ZIJ7l0bd6Rk5c
PyG8AvcSM4s+S+pQupwtkhuLPHccBITvddQbEjZNVM+6GOYA7OlLjCioa5OT2z14
YAf1HhaAfS9RQReIYjyuKqji8sjlEeBxf3qebIBi7zvETHXCF6n68tYOPFQ269az
wMndcg6qtowg4O5ZGQq0OcTL+5yEMh45AUeHzOjg7dz8V6SqVrIzqMwroE1/YIYH
yufQq3FeuTvpbNnWTRCaR/LnEGakgsFdURWRcEeH9loA96sc3d4SmYu4JMH70IYu
GzSpMmjpj7nlVg7heTbwbbhduMYmdNb+f/ejbX1y2UBDj+biFWco8mWYTLBQMVrJ
MeZ9xfj2QWAj2vpkIf898JlUBd/Nrf+2dMUcSXQbNHQ4+sCT2qA1cOelMsyeEEf6
iDjbbk8424dj+iIod2viB4dpx91AksNzeudd+yxb9IWkbp9JVUY6Efmh/mRewv3Q
M4cOwEI3SdpzT2AKjSQMjiCnz/X7iM9XupaiLYFGA65vvExTttKjer3kUXKQTVI0
OG/+m1pU4cWPUanjTwXvpNoI11V47OGKW5CyX0Z4JV80ASsNswChjtE7yZVI20Oe
NkaluPHg7TIoudPEW7zod8pZwVMrWgBoTBNziLxeVfCrGZK0/4tRIcjiFK6Je+dE
Oln4lLSAsTY5rVXDxVoMErVgjbWcCVtU6MWg00e3F7BnWRaTIdPCdO7eytejij6g
/Ith1S/VhmsgKsYX5tuEi0u7GvBl5vhLKY6vWuzH0zmnbpM33kU6BALJZC25qdfo
3Tzy4y1Z9dKp/mfpF7BdE7+rq0yvJoL7eSef5poBE4kRmN7wIP95L/LFyLEBdAiZ
JgU0nomdTAsBfEs0Jm84f0Z4qjF82m2Eyojkr+sCpe6mVA38ao3gvzTehm28284r
5zeF03tHBJV+zpgVX2oAt486fAiOiLeivdUg5b2NtPjMZWGP7piNsJVTdgdnv4hv
RUHZl6jX4c6RMK/J3MVxSsNqGitkuA3CNQa/E5XEjzxFdb1wJzkUhRD0B8CngmTU
9M9H3M2F8DhSk95vaNHnu2m3mqeDRefWJptRScz5SQeqrMGfsjWkRfdQCOfl9DJr
clTQ05l2SzexZ0vfWqdwdrH0zy/QJ030LPL0aciCj9jRduuQp6SQZI8G35ixqe2G
4hLeOMzgpnH9tGXzZ2QU5Rj0qdhZv0+Bn2wD6SX8VSMJGIKIm9IOXIXQRGpN5TaZ
VrdTq+VR6PCFG1BRTuIq9bBtRqYiY+dGOA+n9LfCpLiFi+TxOYjxnMvbxdVPGU3y
KnSYx3Gsf78au53wy/A2BT7c/MgIkvxoaJxwCVzDLe4gLek4S0CoVQEW/QevqvKX
GCCz+2OqwmAH5I868ZagRIq+xqe71y2jEgYF50oCDcEW066FOkoMScy9oZvAJPcl
GMx29FnX1B14vBmzG7+60ZEt0P4P7WQJ5YoWO2NMfpRPf6utC5DgNjNdT0cjg6Sf
+gm8rrR/2HPATJ5MCm2pmvZK5YgBGB9okVjJ8bPYePehJYajESlL+evw12Jtnr4H
Z+4a7ocErhdhIrRkhkREhUr8QlV9kt+xgsRm5geApgXOWdzEhfPLBDAixTQon4ce
k6GMVg0yEVa2lQT+0uZPQ5n0q4AcLCLAsoJbcJYcmsyTZ3uZq93WEfyYRImd2cM+
uHd8PDuu03eRyPf7/d3/AWdic8cOfhY2+ToebeWjg1vg6/ZWSqIohK5N4B420zJv
cOluwiTpXDdR+bM7zOiJV3NkKRDLCDOHiWwYMfvK5H/QLtlQBVJ7HF6G/Rftj9en
CD6JuwS2rCfm/oogUFWHq996t7qR58rQ+U8zd09POn/y7n5M97hbjGRmHBAQPsC7
Kbdux+yagq6lGua1UuOaEwRBvSiYeQG88catoo24ib2vbqG18ymnMRAJS0MBXlkX
jizeAHfZ+AW9Qd6Xao/2pHIox5E/RYk3jcf6nGoT0O/3SYbtV064Mx3w3NuCgQl7
16FvF6xxjDokZED3Xh12y5yIszTAaFaB7Ih60HnYIfn7BkQrlPuJqZgCIY0Yss6o
XFfXGzPWUbsddmoJok7PQWELVxcv4AzwbgYocLmOLawin/kuC8VR6nxWNRQLCsGx
6qvqUhUUgg5wLBiWyDxViAwK+H7WMiN8qXtHBXgRcOm6UTOGwhKy1KsJCfVEFlN4
/C01rme/ebRPLultmE3XdFNiyPGxWXC9OQ6eqO/xtQW8/Ec7klHi/4kUSvFverIM
o3DNBfZBNl91SJQnsNwgVNjiTN7dxIZBPUU0mHVCCLZQEN80WTb7AosgGSETf8Rv
4610xyqsdMPlzX16lEQirFjmY4g6pASGrbAhBAIvDr66+BxLdfxFytTcdSFjWf5D
5BbndNaZlmcvQZruvJs/L8cd/rB2wLUaqywbtBrvDWGNMf4YSyKhsZ7Wrq6XMH8j
Fd4CIfRUrwYmvq8F5WppjWt1sPMvMtFY++wWnk7mIMRKddYYtVA0+JL3NF2euzYR
VzzDSx1eylwORpuP/MA1JAnRPs/Asa+SzB7o/k8Y22X5J3MXuPE4s9LPENkwx7I9
LepOfRV2QUEC32v5QXP7VrEMKVQD4VvXwqtDpA7wzM7oG/TABXHYdQDmuo7pIRUr
cRtnJZH+AjIgHjXF3Ahcr98sQRP21N/7QIw3oeqSb709+6aR3Gfidc6Ou3yvdLVv
+LwEO711Hx5bSaMNsmPcx6CChk/jFjIqMm7Lqx3sHnsqJncTLztiPZxing8A6IY/
/qPAHQRKiCRDVv085nHHgmxq2Ejo1JOoU0rPAzCYnMQ9mA4KE2s035aCuIfxejEp
cW27JOkAgUaMxr8NeGmZR2OCIBa0rfb/iKYUXJuDQJNmRh76qp/dFUtuD+9FN2dj
QBGWBg+tWqYnngviwu2ut146NmtiozP6r8oKhsssxRuAFVFiQNP+Z0HN5cpvECnz
yIx0sImCnXgtNADU0Ty9szm672AsoJzTUopJzYAemJOiBnL3Nen7psARbsUnGFFY
JtRVGUkrkZ0BceTeyDer5XWgIVnTMK1vwAVTMQx4BAvdW6N0mPIEOAa7owYP0nAQ
p7CbEVlufiJrxOir4Mm/X13M5fBWAXshMaarlgAGofO5a0/Ch5vhW/4O+fDnRrXD
dWMkeI9jSdUXlVkM3jsHunYeoXVY+CO5I1Rs4gPWlPf9yNjKewMZIudLzW3WBpIk
KrUGn74KyUGVBMEv7Tfa/4lo+5eiQ6SOLuS3BS/fY2pHuzcuisqn4vXySKCW2y+t
cTxGdHao6CQ19xcoI0u2oSs2qv66AA3MhJcCcOuz47gsx+sC3apTyKpmn1ZaNqAC
uP976JDUGPOlHpcM7sJkEithswYOOVBOEzwpN8rwzfp3gTmi2bepIP9sQDanjY/x
RuMw0b2Dbexlt5WlixNiPXhbD6HQzWDPu2L2uJt0a3AwbsBz8CLQQRHyNFskXEzf
qVA0Um8XIuaEmTo4fNt8c0QIM574aCP1A22ni0YopTidQnNstvrsY0ONpq59bYdd
JK14WpksAp/6j/YRaxzDrJQvBOnTKvNjnvZoDPvkceLEQ5QlZsRt1RVVv1sQD3Q8
ZGII/ZHIDeBIAcstw8ezRfNCIbQhJPiA/tUgzIthEmHtgnjMp65flyKDOcFSy9Np
Krk5qTRgKKYco674yoJJ8MQiM4BjHxaPltAMb6Hkc6Lkge0MeJgavoweIAx2yt8N
w0IpkxOA6kCgPjLcOo77oF9TTNvCGJdvTly61lb6CTTuncXztsdkIX83ReLXJMxB
7J60WWV+FpqF2Z9TIeDvzWEP50yET1ZyeXIZAWhOxbvF0QRFcOFp7s2EsunTPEfh
OggrUX9uLhYdf/4OR0N1FH9kV1fZGHLFwvh05navcTx2xeo95lJmbKmw+q6P1XhW
DzLTF6XnIVr1f3KRAh1OgPoYlnQeA45Xt2Glz81MqCmnJM3R3CH7ueii91JOz01D
Az4sz/vOdocmTyHEg0NhQ37e6Ci1UUW6C8V0NF8s+24Rlv71Mu0OeiOsPlvDy6MJ
sWzW/f54RIc+brP0KaElFoB+21/rvwH5/ASzb0G9vh89lDobHTmKURRTGLIc/BXi
Z/zu1Qtd7fX4OjDPyn7WsU1AzeP5mCEZsMyoW6HmgewXHVbqticA8Y2u7bwSL3Rb
X8QmylCZqfYVcLhIruzBwK4aPUo9WW+kVloEKbHXiljpmus8umuLLE8qG0hSjQzk
M671dh588ueIZ5LfD3WxwTp3573Q960vKjTF0V2VHfly5N2fcyDJoUrIuKrYWqJ3
j/W298KPGIjzDKd1DeTM6M/dd+DdXOnBFEljMCvKyiHTx0R5+vnsQ3ghZKuRuvUk
US1U7cXWnhN1dVLrO/hYkUXXQSt72Tjytm9luk8NObAf+3rsYUmJRRVC1gGITAwB
oOet5oaOJfrqvYJ8maUT22p9VQKzk69jw9Oeu8F1mjEwr7mIDM+0BeDxSXtco3Ds
KnGNM/P35iqFY2DS9Y/CXxYBRhAjTydemQU5UWOxBw2Ul3uaJPr34xoTaJ1cO0GI
HsJ+Zie2zEU78O5Pm8aYNjZlpXHLVXrhonflbFuFnTiF2bsRX16Mpk7WYF2lr7LJ
meFM5kIC4XOqdI2aija0IAkTxRR+Lf1trt1oU9sO6/pQ+MSOwrcShQUVZJAHSQ+J
vNsO67pZxAPDbzNjq0CvNZb3UydAN/46YJ2o+O+LU7zuW9fneeCJ9KHKHx1W03Of
ObXlsIKytnT2u/0Bwgpu/AzdSWzWSmH3KqPc0Uv7WysysEZqU/ykbPvb1rQnoCSZ
XUE2cILBCKSrw+fyIcpumk6nfU8lDDU4nGrVxm0X6apbAMknlMDk4dNgJW65rN9j
hPBkBAKfRG9lNUkNPiVwtTpHKcwlkFGOCSG7vw0pz48GUdMjLe+WlD89rMGKdu1V
iehVh6D6X0WAYPSFKBAigXxSgJaFNq9a5sx3nr92XzmHD7VnTKN79rEMaFPDXSfH
uN4ziE06nWKPU5MXuVKFEd+vuY21VgnC1jtR88kSfxBhWGNC+pFnFojlq3q8YBRR
SLvE6JwLo+2qTlcyRZdFL5WTZ+OGUUOPdPTvGVn6DmC4jzevLHTcEXszqukjm0Dr
rBv7wBPvYCEOreQ0U4DwhZUDRaFhgRlq9SeKVGU61e//ZjhVUTgKHCGEn/hrT+Gk
pSseim7m0OnzOQFsY4U31ztXBeKc1uDD53ODfDwLa2eI52A+zkRMj1jMPIpnDQQz
uGNHelW6/YEbne2LetxC5nn1XatnsDyaP1osXHHn6YvOecyMZsInBNOp0Oti+2xj
vEQ7/BKHp97aIWWFZA32It2mI1/K+HH3xEg406azWnIpDMnRgBugw/rzdY7/iU1R
PdTVvN4pQoHTp+66q2RAeaA3NKNmWMEugwipUfHvWVxq8fmYrJiEJbJry4fshC1Y
DTQPzavvDxErtv6WgT8cKBwIhzjVqRI8vqrfbPVn4LdLvsBxJxn679dp1R+LmSYY
SLDCTaLJ+OmUBN2xEsaEzrXvtvPCXpEXR0eRjLv0POv8T7if2++8sX+NhZO62Bzp
sVN0AtwswFOK8kwEP29WaCAfHAqnxkX6YWR2Zoi2jhktVtSSXnFt8KalLXGmC0x4
KTNogQiO30i2DrRSxXpNV5KFgvMsN7YfgSkmPvQTMzdPU86cNYmSfkAKtprL7KD4
vJkpYQdlZ8azJ0QGBO1cOn+Ir6BojRsRhvnBTxYUifBdHkZSIBNRBxtxA++DNZ+T
syk40W4oL7UARPs0o+YOzwclM4t72sDI0AMRmnubaBBDN5ViVn8NklfZiMp6OPmr
aVlJqOMiOxnIHykW+VwxxRp/EV4BauC9aeulEHJhRCqJX0g9D+xvKEPnI0DZGK35
dl2zALUJeSLg6HpIIvwB2O905MYMGiDlS6lPCf2XmQm2LAi4+OMHZ/9w6zkFfbhQ
OX9pbTab5QI3Sks6cUW96sRFsZc44STyIUbiaumCIZnI6AvgL4W3Erv+VnfuHvrE
ukA9RCy2tPctbQerqeaf1AudgTfCVWuT7YiPcMeW388X6DdFloZRStB5DKJERBBz
tJIw1CCcvNh4zyCJxW0WGFKNGW8omtapOzeQO+RwQztl1xR0rfgSmrNpVz0zr6bW
DvLxEVmB89h3FcNP4foaYYEQkh7jfnDOdRESXrSLClCXyvkQKkox+9QfY1tYbkzn
549IZ8LVB5X9yA8Np3aYC0lzFuzFxhnXZnbDu6BnD/SzXaK6WLke07gaLkjmKjKi
muJiZftjV/xdTJKnmMpbPeL6FGMT+ztxN8ghQ5GYuuuVkgdnfzq0kYPLsyG/mEPh
xbhWQRA+Pvm/h2wMM8eXHC5hGrKV5Jn9AemMtWxBbK7HUX0XJyWL2SxAWHkIDDC3
f/NVh3oQ6IqiNKynrdnFLYNXT4sftYYdJfDRMmzxRY/2U/hj/3+yxfweRYPOUMIO
qx9QwOaVhdWHbAYY6FBKaYrB8RINLVOpemjJrSesJwbBUV3Bgft3XcsuaLZDEtoy
xpPIgulQUvn08p8ONPTr4ZaL3wFAxXZe/vqPKcu5aZ1xba/3NF8yMO5NUaG0dOZz
V2Pd7rhJeLqa/PUvcbPw1gsPOg0/SU1AS/IRe06NsKXvdn3saUvImS7+0ptpSfcR
4c8mQBtR/gfte/5MIC5+GM+ri0NjTPUZI0v8ZhHyAtNsxdVgyLdMpL74tgpfuyD6
rXN0YUkxuXZlTNYFf8gp7UIg6keZbCR95Cu/8vxkA5+K7m0fF03h8LFxKiw0QPwU
GK62A8paUpq91qPr2QBH5UIcrMgN/L/fboQ2624jy0HLUcNfxrKEUa2RDEsOAWbv
tfb1qC8tPM9sZbnc4fFQxTxmAlfQnJtR6MikQV6rWRAVqY2jVbZf49VZWiaZbGwe
qftW5/BpYPqiOrdaXqi32IDAVVZQKECYDgDyv7rrDgAO1+pswBmc7LkWdLX/YsbT
j1yvqCRGROqq00H+SjTR+/oXuJvn2cHPpjzwI2AWXjrVoODzjQvw3Wm+36LT2kFF
TJL0U0GH0SgwA46Iz86DGBEQE0dArC9pIp1GHSijxgwEQK1Oa5MDU/r4fsoqt5jm
0dw93R7ttk+mvWKuqAePkgqjdopLZyomfGws+5fx/6UJsLeRZ5AY9nZeo9lU3vBf
u7vV2LjFZK82f4MeHdUCtVcjqN2yvUbh1+B6niJosFDuzzNdX2OhrccaUV5PyEee
WyakEFld4FcBHeneLG1QNkV1D8/0UJbgMbgqBZzCSusJWKcPqM1Z+BQ9B8syWRe4
h7KUFRPeep907CLO+Af3yC8Jtk1gQ9xamEw4zxBpYfvKu829YC0RQl6EXmKhu0zW
uG71cI9wffGRnwygtoxwwPT/RfQq7WN3yiokPGtPd6PM/8YKj969ws0R1W1pf0GU
TGrEKvzadDG02O/K8H5nmo6LPDq3TWH+FernJHH1+pwzmV6YTsthf60yRCwzpRZc
0lk61RDY4orKphS/IapwOwgf22UsI/C+t4It2lDG8aS9pSQX+df5wkSdpQS81KaD
QyLysAeisxs1Fpn8QZbZsCqEI64Lo7itR1CcSJDUpiUUS//97WayS4CDSynGJ9Jh
7QB9i3HtrimMlZCDi+My1slQMOSmdBicHIZM/7yLlY1S+Sh/oFpR6IgSsR3/kP/R
LCjRYV7EJ/vo3J78RDPxW5nIQ/RtQX5/HVTVXtptqmffuLZQqf/HTwZImTZ4i7dR
dFEMzVqGegZ6LOt5pZwyLqv1OLS2Y7GpN2G2yeZq5GhrpTCsGIpFoEXXogba9A+6
R8XFl2bfj5BnNh+wkkKh40/BmgohwPqe3k/pMtuqC0KdUByj181bEX4/7jR18ieq
MBDDmUW+w3rl3unJOH/rxe2FvpNQBmoK5W8THD850X4yvau9IIwtgkiqqB2KwT2/
rk31j4hjyF1hGFbbkI9JV2NNqX0Huc+BZMtzZ6iQODllIsDCDp3JkVgk9r3k0+oJ
s2hjSpXrKFEtAsclx8H6CQpM72zFA4MvuOwUgbiTiGtAW8o5fqy+OD9hIOavVM9A
Z1D/Ssib1W7F6mhVgiRAZVtHV363n0U4Uwo48qMhrL5njG09E82MKLAsVcT6vm8x
Mhw8zzo9COepruN21e/EUh1e58TFHjIzw7mjXMmYcdf6KkqUj07o71yn17fpdSiv
D6fp/uF8BTbECmtyg0kfDcG0n+WOAG/VxCHfe2LPOPIz116JpaPbxa1N4M8rN87x
lpGC+M1H6YH7osJMDYQ51XXA6SAkAGLuBoIQzniWO8Ker9vgv5hCC+gqxSTnjVGT
JmVW/UXAHpEGnlAhYIXuJ+wGMrSVpx6xqKsafl42t/CNTUS3N5Ba0zF8dh1GTEvq
ESiQdFZzygMnIU42I3Z1dLmXYh1CDQZ1imMjbfklQq0qKp7UjdKXc8tK4mOCkRAa
nYNWKNL86UbqJfNbXTXANSpWlCSWJGddhRsUm4yPw4x5bbVURSVvfbMu0rchnsO8
WVOTDrfD1xRgPhU9zSlYxJX4EU7ecnl2iJAmXP1A/hWEfOqilHyfzbo443AobPR/
8XQUHv38PxnygTWI/XzExSZGjeYyiegW+E4Ey/+/Vpcux4NbigwLJmO+y7M0fXEu
n3nYlk9kfPQXNFa0XIa2VR000D/WXll6VfXcO87dAzU+rg5zFTqNgjezrjK71rXV
5fop5PDTNCzc+OqxrMKldmZD8bvAsM7PWyBvqikfySg35qU4UMlSD2yZQP9WVpKH
Y1D3DOsrLL6HoCdOT0HhZ6HkSMpLTOWS4AuuIb6q6RyeB0pGg1brQrB2brCVgvIX
s2A2Bi3AMI5GLs4H0UpdbGWb7AssoEt1r28k3Gi4hJEzASnYpbqko2Z2fHHnoAJK
tjPZT8m4CQQ4C+9R1OphdCfyozw6XJDDWBT4BMCBDwcjJ3b582brFghmEDa8bKmZ
lYZVgTPS6nYCMFOxyo2FCE+p5cgalwepEcb6deWqUTLoS3eH3Es63iYdmW+cJAs+
ZGJRCMwyMUx1rhUqoauu5JYT3eTreDxz82poas6mDf5PRWWrXNrP6iXZ12srvFQ9
GJGu5qaYdPlnFkts58vUiT8N3Fs6ddQZvf6DD1iqrERbQF/etmvmUOUP+Az93CJh
Z2MJTb9hVCyJpMN6wufMEORVvIvlHWL4opsl9qNeaqQg9c0IAAvIJQq0h8L1+9I+
EeMPddH8SlJYGrQB+Hcx2xZCUiwWFJW3y9OoDjUL6wVbfn5GRYOBcPwAk983sJEZ
ZvpGdGaSq5AFpUkOsYxOtLswf0w4oxH80JRcl4tTAVJhfChypTv1sNr5NPWjaYJ0
Q1pXP9mUExWWLbJ4cdcM//wz6jq3jHkrV6wBVKUUD9c119xw62U3uN1kNxzCzyLE
W3LVFnwB61wA29LJpKMlSNk77D25VJvH6nBW9NJ+ZF+CZO/6a6Y+eiqChUUZew+Y
3F39CqdeGknxVh8ZaAjypcy8mEQHVpz5zGFicLgNizvP76F4iprW7qpMxEVpuwpt
1eqEek/2w0Q8mSBYIdjKgF60D67I2GbEiD5f/uM7V7U+yW43nmJPYL7O9hnjoRwR
hTr+RNoSP8NIMj59I4pN2Qw2GbeS2JFVw1oEqQekK9Su7h5Rqf4elCLfX3fH7mYy
LI2Y+jMU1HTeGRAK79zt244XH8zz9CJ5bXA3tagqcxIEWDSEKduWR9zsZdWMH7E+
HjJhp1riDtjzL8ti01RlN18HwKzuwdu/NoYKLSM+QOvLbgZJBxkxZJEmJXAjtftW
rr13a1x1zLozM4htozFgs9dwn5pvj86mXX3P6Ix56mtpPOW+jr5vj5CcAEYshqRy
puyw/ZbAhV14f3DoxJmFDF7rg2dMkmsCcNhHCaRrZI2tg/N4NlwRNtg5vBfp9SDf
AEa+RiGgkUnfAGLX5mLLzT4RKkQ1osRcjPpj6nCNGVkcoEhjemqKrMxftX0oIQpr
B7dM5Sa4myNoGuZk+jkxUjJtBFQ84qan92bAC9EXccG8BDdu9kD2n7mKFuooF7jt
Q15is0Ywx7P+HzNGkOnuFHRFZDq/7PhrbP7PAyg5kWTv5K5D380By7aNHWsoI6+i
2/ViiqEsHibYmJ0Q3aVQPfImyTJsbJdHF/Z2WK4DGk4UbXmvGXpwiY7gk9kMcfak
boKE6Xn9EQYdZNpNSigg66MJTb7+UFkj7s+AJ/9fxi8e32HGAidlfxEy08uMe4aG
KDCncPFK8+IbU5zzeyz3KvO+7thnEdxnecOrcmKBkAJIP0pFvWrDQFJlEv1sw7A3
JduKWFiS0AX3X0UvwVEiswafJ5JLXv1o8UMTgLqCznsufx4ospwejLd2W5tTWemx
BUVfO5a7+BHNIWx7ZqIyKmFp6b+f4G2w9IUBoun7tAV1Oqf4fnq5oi0ABOL24e+g
YaCZciqZ0BnI4oKeIFEzIm/CMW5QlKorfrl4lcjYYFqftFq5qbzZITh/OF0hO7Uw
AN6CN3cBL1lkbE/FKC4lqvGhFSvgtq6+AwRAcQa+9Qq0nwUJYXvK470nP+pQU3hc
kdavU6rfBcAhcRT7ugeHTmugwsIEaj9Iam8A/MjD7voSmt7GPW3YS4GhqvuaDq/9
a5rsTXOr6MfU9y/Jmd4YsFo7Bnp6gKQcicAVEI8Gto3ikcUKm+RJYJ8jLVo10Loi
0oqpzh93n0oNNFAfNTGRpqQduaDgufYTYQXHj/R8wYWXvM+lI5Y7edy300pCadkv
0yO0ZWPGUJwCWiFmCnrKsdzsaQSyNf9JhM1Rn+InwX6UuUoXm4hN7A9J+hOnrmYw
+lZdppLPdEfVmc80n8pYOT2KbqR8n1lJISww9B9KnkIszjs9GTP4hj4qLqjTeK+W
aQXsF6KqD4gZ1/QpdWwAG8Hl3PQziLSO15c3zR1YP/1Y2UGq5xLzX6SPqbX/tOZ2
MdRSCfJzqz5hbViOiyxhI9KCrPeoeWW8EOJxRuMWiIeL1iVsZI9XwQ82R6NNucIK
wuHbIZEkpU16AXR1iDyWW7uWNS+2+7ur0mN1iXUj9hMU6YB31veRVzSEK4oNeSn4
`protect END_PROTECTED
