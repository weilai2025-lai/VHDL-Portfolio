`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnNBJF5t9A0i6R7s+QTHH/RabzKU2Y2JGifcurgDH5iyFubaiDt6s7Hiki+WMQ7c
wzYl7yLnZB8g34oTYSoq5s7eKZEmOyjBmcd+wM/B1Bw716dIScv6sq+MoOc7un+y
yp/s441oQSSyVtez4e7O667IEZjfrIgIhRnFkv1+y82Wpnd2RrnxtRot1Lfx76IJ
eXgER0nP0IAuPioyt/nbNm+pOEhGEk+SpoEkhfJmX8SvJ0J6A/6jfJ25vAsjijVn
KisIXZ+QMNDIjRrKDOwPSGmzfXHdCU36/z+Lt4bcawhtjP5v2Zk0TkB4HBXtD+Ss
+1pWIXQOOH6VL3TcPn6Thi8xT4idiFxgdW9xtsgSjEoex6cZxESGjAUNmXtwOppl
6St8/F/IKKn+NtzKPhXoGBMSLJA3UteP2nrVg4EzyHn+ySo1sjDcD5/zM6pXDukp
jQYXlID+jE0/ylwSm/Vl/SDmIyDo99/xDqSkWdhWpbtf1JGNZ4uFVIqoXQSidLYO
QOkpGvQIZxtGizCcWwmajv65ekIv5zWFhIXft4UCKy6jgNfhCcH/MB6+XqV8lTwT
L5FmSIE37v0C4d8XswB+3Qh7BsvtJvED5SKVYYfwRySRK93aN4I9qMfSrxywIjfN
wHvhAORjYmX0rtgLy+vffNckcuRmXQCIVebXtmbFHjW/HbwCgiJkPe0D1EYKF4wk
EsVTg1AEtFXEBQslKwyVzDabu6FAmmRBljV4TROYPGZ+mFIK83hXTl4E9ACZVL01
J19QTaYPhLJchi843cvVU++t4BFzxs1kPA5c6FaD+pxvNREKBYC1VjU9I3aWJ6F2
Ex0ytxUfCRRcooq+dXYj/a4VzNOatVugbycC69I66Gou655fC69AqiGq18qwMJhv
TpZHC5EfnOKceX0TJ2PQs1FPHwyQ3W0ZBd8oBUJnDFN/8VWWSWBb6YM/OX7vfyPy
/0vQweVNyRJTnMaAfBhibB9WblAqmFBir9ER7L46LThGZTgR1G1ZUVH7HXWH/ZpN
pgWKnhRKsxXFWIMf2DHP88XDqXXjWwCGKY/cSygFP+O5CHP8weXCosdaeYXF1TEN
GMImm064ju2Nm4nNYnnlSmLwnPZqIT//GbWWDH30Mn2zqIJWMDeWMwDIqNOqt4zj
g0ZN1Djapaxv30x8aLw4FXNeyBqo+zhdX6spzQFW+UyiU1HgZppqW+s1X9q35cPg
/AhBG2X9LyJrPyMhf8UrR7SpaR8VtKF1MLsfCMHtbwXvl4jjD9vtlm1EOeC72+r+
7XYpia+Z7P4jznS2CGnRSBboHfwwPRJsTklLt5hN18lQ0aWzKez/MHql4GKZeii9
yDSz2COnRi3bTsBeWVCv7bEmQ9TUibRE3WC5bv6ziQGkKo+HUzWweMGCXOV/TalF
S/U2JsCdVobdygJZB6CCO/9U8ZIg7MQYNJ6aZxnJXZloo+uWg8qFloRI5P6VwVLH
kU1HI0NDrJ2RVrNTOjTcblVfohN4Q5sAnQ4gbw6leeiHd6BKfUi2r1/sdaKg1not
aL4FNfJ44EAS5+nKcvvT35Vjqv7K2u3hPtvLfjEl4z+0kFyh29ilSGnXQIpmC0zG
ULXb1cAn1Eem5xeq6Scu6R3a8mKGnHOImKAkIG+VnGOV7JTx3SMJDqIungOPfGSt
4niKNBn6HRvElgtUljKTy2kIIDO8N3GDnB7B0oB5g6Z8EaGLPgZAaW0HHuCDtSUA
GvxqJg6CZwjZQWiAdETL10F0yPnJ3pAIdRHaTT9cAjiGQYKgA1PmNWSFb1m0z/jh
mRJWUJVsqJ1lTpY2e99qv8iU042+RQBw7hOjcctdduQvSm5s/gnmy+fwJGOcRrYc
W5q8ZUe8ilDnyHIkeGIZ5Sykwha+UfcVpUbsScxyqLTi4WkeLWKeKIFxD7EORbhG
kuUSBVuFRyf8ESJv33w/zg==
`protect END_PROTECTED
