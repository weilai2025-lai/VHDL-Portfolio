`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HD73eRY70FQ2B+CX2yfFUi8/G2Ys96buUZwC3kdUszHxCbo44KfRPw42e9Qvg5ts
XGH5yrNM71WPMgk0d0lRajK1vRRhP3ZiMEOtNDPMFPLhymWuwhaU0/C4DxcWk+MA
wqGh2NgOuzTfDBwR9mdEvS5iognF4Citbe+qsbsaXkpllsfxUXK1smbrI4E3SuwR
uncfOF2mVVRcrn/OruV6ybRPg9EHilIxwju0HtRdskIkIbtL2CkWzZVtA2tZQLMt
a80j6JuPMwTJRUu/R1Q/mXMoL6sdIMNrIAkGth0EKVrW6VVuU/f8JRmj0AorQBNM
S3NfhhyqK2JrU7YhsCd4d5jKitEu8l2qPjqzbjzli+Gw7pNY0HspwmaEfMXEl7c9
zRHd2rmI+NHUQ5P4T4JZEMfM1NGmx94eVHAB5X6r6xk7UOQgECPHdEBaxf1ZQJY6
qPfmg1yK+WOEe1oMfVw81OCAPTEyoJQOCj4g0RbJMkd0ytwwgqAolpDvrS1HnsQp
qKMxS+8SdITwqEmGIsvmIe8PaciXSQ90ZpcCBbQBrI34Wz2XahtIHrBhyJ/WiXwX
Hk41pQ4Rj7sSU0c7MSEDJDkIbp2zVtGxXAWej8/u9ljo0TS6fxH/xXGA+ylikVNf
/5MssOH7b2pe+4dUEwN45C7OOQbzjiJDEDY2bwVBX4VmQTa1cusiZFZQcApz+82Z
E8N7TD9zMLhKvMMxk5kErLgjAt0Mc2rWbdTehGASVAWFHXPvT1WEzNHVoC5XvuMW
OF5gmMsnNxGn8XZWPxpoUezMY1p3BH/+BWph8yHi124EykcTHXAn3hU4fULWucc/
jPAnYQvE04422fuTCMxS7ZL0olNaz/YW5XDy0OfKomFHUPgfPUMAjqEoM1AFu2J5
5GuSvIms9j9NlcsI5IUIP7ZawsyYX2QIawcf0t5t2FZYIPRjS+1oR4zbambuRMV1
lenDNXoudw2knST8X/36XI5tenFRGVKx1UnqmYCVXW7PFCSqGzIJ0ra51UwtAqzy
ShoO7vbs2JZ5KbckWPjxMDINQltIygyl9yTam3nggfA7of3rTzWroqIDwFe/NlAB
Ul+2AzhUZ2wb6ROKn3tkmffAMgDRfrRzqs9Qo6dco0p72Oibk3MqP9QHJ0TMvBO6
Wfj9HqPIpNVT886ZWlpBy0V7qRHjAN7VgfvpiH0rw00lUO06095VSx6amsgsJbm6
GQ/RbtBi1CJZiJ1t7oC7AT2U343fRUfxJlatqRwrWqsqDK9qBZw3Dzgv8o1j/AW9
aGWv6VXWSlf94J3AOXs2mz8IDh/+LNsz/P704cwZfyxM5U45F1UNbf9uWNjsvtDn
lBBpX4Dbf7wyrIOC4QaKv/JFcxr4Atptil+MWIFxjNds+fIsv+EaRVmsWirTzcks
m/VRvbEqT0bmE9VSOd/1bHhCgqfdzrWP/piQXvWAByPSEb8YFEAE0Tq0UMI7bu43
YjCnzBI2CV/7lmJVBZV+4TnabKnBRMIYvP8F3/KjiOCp9Z2LYlSQaRVAIYDSMaoQ
P3Ll+Lij3vjI9n13o/N4dXs761JugabxNeNsS1D0PZvzJ0JWlhZVYqkHcauezQHg
F4CQ9grxURLZrQaXxaEjTuRyPPZRQ1bB303l0HJt1LFUzUdpQwqpxlkkkb6m8aaa
x5rTOgSJEsoQ1UxnNTUO3tDEM0hx0t9/Cmja3qE2+ym5PNMQCb6Gh7uGbchxRbxa
FeKIJb2EV+HYUVgw/5or3xi7XNx60WFb/dtkOS392d/sU7S74n8uyQF94DC13Ebx
epS1rNvulDF1Be2hAEL9kw2jwCJYkQG13mYO7jtTENTyMGxX3bdFFT4sMXvGcPMm
8jP7VPPS/EFURjlbYEZdWPTbM2o1yR81NfVdHlNVPFP/Udqro01F5FdakeDoINLp
weEMU0ykbF3qHcxxIvm34eo0GHeLyTsBQK44zw3PDAql3NT4fcBJuEsNGEFI77uz
Caf/J1ua/8szKSofguCW/5w1cPZjHLArZvD1OYPIlKjKxqM61KgMvZLhrbbXObPM
LXMXsLDHVS4Cbg8sJNOBjs1y+AayWAfxnGwpjhwQphH+83FjRpBzxqZCNbu78HDw
bEo356fxJNTtj76F4azCpLPwTTchJthup3PZYnUXda9uM+iCfvNWNAtQmBBtUFlZ
MEYUjIrRjpgDDTxsSl5KvnG6e1l6PmxHg3LeTcY03QhUNs2SzOgMZOsFu/K2K8pg
cPYUlRp4E68D8VyZlWK5ulHuWALeSgYLdzvoFA1qfPND4jonXXjgtSzheArP2rYw
fKMsougaP5tXtHaZZ1Rz40KoQ+Okvf0I0501bLDO8otUg0XSf+EGPVf4OjMq75Lu
6JYrNmpeKyVfWU2hDenLzzmZYo9+ZucjKvXg1tgKh37PXZF/gz31wgTZ1jXg68IT
VQch3UV2eMob4X8eC/oUTOo2rbhGz9bMGrOhKw/mgPu3+4uBF/xRfBnsToco+d4n
PQQgj34E3XM3SYLrkdaas99hI6QeOtvjeA8W8F7Abacpb3q7+yGDV5+PIaQrwIB6
IV446RMR0d64EXMMWuixtOoHMGQ2AjGegp0e9N5P2zEuuAoGKuVHgUuuM8sk8CLu
Rn5n0YFDTPYLAisIRuD5QhdB3rdvHzn3w6WL9QtAOCi9W7r+GkAxfd/5TzPHmSb4
gyW3VvSZwqdPZbQI1Qb6dQCIAyX494ndtoTDqKNYODm7LLDVqJvGos2mQsr/PvwA
K1o/wEhz2m1Y1nf8JwMWVDvJkIu+T+ZUYGdBh2/vOXneRxy52yYnFQjuMNW9HgY7
r/xLGs+qJfMA4LtACV68XXQ3Q4Ixttgqsftz4Elgq1wP5v9ZX1FqqzuKXvrrtdWX
KnPTD/oQby0QBZKU6Bh6msap8fmjDopZG2hF8a1ECm1qvTj6V0gJkmErlQRB7vf0
ZABHdInFRxAf2ZpsK7LD8DUyTedPegrdr2cTTj8IUhO3Lm7tWHbsjt8LCqLV+m2J
GspjON11FUrBBJ7tcPVbtuMyLsZdZFMpiNu+cmBtkkTXr/PTAxniS7LoR6hLcbqv
w1Nb+xpLG25vKJsXahLDIXZK21BNgtz/QnuPp8i+3aGpmcsK0Ee0aERfYLqszY8Y
e2X2b0cDXqnfUl+/i3OzSNhe4QeDGty87aBAy/YTNL66C1RbNYgchJ9AMWRDgLFS
14/aIrsExa0D/0xlqbP4BFnJ+JBIB7Q5LSzWawaN3FYZhebiIPMt1MHyY7Z4GPTk
Y3la4ZxiitxOP6stC4BmB42wmkAHUJEUxA2v6HqiG9lUj7bqrj1fWTZBmv3IHhfD
NemP4uY9v2ck7rHMEO24OiULQd47oyswE9evLPN4eJJs/isI17/YYGdLQ9zGBWll
qLN/7vWhGs9ZWqFLLKxhWmY79//g8SZB4mDOguUTBtXyJuAH5XHX80H8qvvJj76g
ihZrqEdYfbw8a/+OsmLQ3xaAkIhftQBQUZsdoEvcNb0jsu97cvOC0HBqM+k/D0s9
`protect END_PROTECTED
