`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/R8pCMb4orYSYPkVf8dsYwsXojhLcm7NVTVor5imfmtEj91FOacZ/zz8Cq6KLnLq
lZbJ0sYpC0x3sB9kcFqVb6dP5UYY2PduejGhOpxxBkXcn0fKSBzMIwzFZsCcaM3y
y445cV6uab8NXICQ5umhQI4B6NaCMk3p+9bogzvVwEpIohtFcZ/h8vlGCzRa+XPe
UmqBwo+DYozyoeZZKpizjMKvcumK9Wu1amBSW2UoThwD3Jo3gKlyd1Uxqo/C8I8w
NDRnYMnXwPOBC0/WqVu5OqV2hFbYpVP/OxNJa/G1+1KUuYEti2X0tQRjxJrvKp2L
pWxseL8HNNrVzMjm/u58H+56YKjd4q73JPkFiqIFydgxTKsyGFq9btge3Zgqdy5j
rpQiYFjyr3Hrqoo2Cak42Qucdhbe1lVkCJlrm4gW0nzMx0otLVgWkDaFjdI1AF7X
egVlDhNwf0z9jD/1D74vwv6u6TRMrLsbi8xpNrX36qWJms0jU0Q203ngTYWpd1bx
uIuKrHb+LIxEjpSH+1g39AhXjinyq0Di1cxCZj3Czc0vfUEq/Wn1DrHdFEeU7Pp4
6Bke0qVwRepQK2eRkb/2ogVCHHx3Z4JVjkg4ww9IunVRY5FaQbGgT5iKL6hdeNcN
8g2HTzTAxEtM/zmId9ny/uN/iRs1eHOhe13Ye8bbGl6vNt+3qbXkLlpbSCaLiTUR
jYvGlY8pu523XMKv9HSLpi1Bq28B4BfcLbG4AbUeOT0ViL0WiwdwHbMUuRqPQaiA
5iGkobHZO8aIlnzwFnQ9uW8K38IZzazu80u0tlzh8ALQqq3EQ05N+5tEjifrUM3M
/JaO5su3zHy051XeiVIAEOjkx47qspFxCfRDEtLhv9561VFUxdldyM31n3l4tY9V
SPM8UJQPf0tNzjYPeJeEfpx1aYOTB6w3aeYfLEG7D33Kgg2kEZjo3KHfm/PVME1A
ReRdxAsQ2sZ8PkwhVBfU/1/hCPYHGildXbe0TeFEykktQqo3NVUqiqHjG2orQP0C
E3PeQBRUJo2HVgRyMOC+9f1pnqsEBjLN4JyqZd6flsEvWRt96bl/iYb+xbG3jqQ8
3J4poAL0jqE80pSoVMC7JoPXdRg40ZjfmJ5iX3vzJc6j5gHHqbLeWIENaQiotDRO
10dPHivxp7MCa3HmP05NzsANDKEMaXg0K8zYJk1NocNDvDtVkMh8HZy9GUO0WCy7
V5wDf8psEQ6NrkEGxsPNvAgJopQCyWZz445CY7bwBKrf6Xd4aJYQt90T46U0AJwg
jYtWkQ1OXW5JTFkO84n/kePIM8Om+7WxjVnIohjEsCiBkjkd4Jyput7UFWQLZ5iL
lEcQ5EdQWij+sNv/NdzP6vlfYK53viVZ0HKmimfNSIdZmM4T+3/pANDsdDqtHSZd
b4fnCHHwycuxV7xFglK5ZR74kvey54/3gL9vb6MtQPxICw+3j1uPXffEkjfDJPFF
hSuXdKtFpEqe5FNSUI0MZ4pqcOVNH29r/F1FdXmWY0YfBXT563o+RjalpIo4nuAD
x2Rz+b01NJWH7z0zeBOdKJcWgpX0Pg0Pm+jmkb5sqXVT5FUkKDgz8L73s9KODHTl
ns0Su4KFuhN0lCl0NLOVIrGsJIy0Qv/9T8F6T0W16h+xqdGd81H8hV+y5kSpzl+x
t+tPX/AWFsYk40LTmmCAt2pd+1Ymq6RC5qdYqDYk3i+Zom313J4gFHQSLi1jqxz/
5KQCaq2WYgqhQHNj+oCUGWnTPv+8kwFtBlli1sJthg28wac8t5fq5cfARX2csSwR
ANZ2J0UunlyIgpYxg4LXfwZUCV/byBpmxLIw7TonavobQl5x4fbflAfUEaDN85ru
mvfKIoYC/xQk8qwUuw38e8ybLIWGnZ+sqBUn4kcgE21Eyr/WfVLub0V3fLvEvtBj
NBN8GNwFGHgPlj0z8OhXaeu7NBqTPrbczjQkZD+5mrNcx3men+syOndIVSjMU5Ft
nvm/RxrDQ1zJ7QThADXDhA0kAnuHOJMZ+bYil2EUb+8EffJZMg+hzHRKUrujotm+
9wXbRpxZ4qL4CdL0ZesaLbQSIakrGWnuK3LK/Smgo7kLwyX+xK3mPgHjGudNcxFX
588SZMN5/CWmIptlRHNsRSkGVVFBOPcNkm0Lg0AKyeQ2axVCQ6LaliYnHCca2K9z
kniyn6x79pHdBeoZjBgMc98gwOQygBA5fSyPZMaFvbgBdWP58IZ7PzgM5HVIpf+w
Zqfw9C+y2lSNHZ46w8oNNb/fJvkDdMbNCkGqU7C4HqK20g6fCvcrrREEo03uHfQI
rm25Zyfi6nAXz8pNR09Jx70oysVhbnqJq6dGd/F5+wFHwvVQR4xVdNfBYmOrvhiC
FVF1w6/ig54uZ0FIOgqrxFcet+XY52WuMLmZDB/ONYieqV1TaNRj5iONeVtPBNqh
NdMLCRH/jxYNhXsTJfSe/z9lIDV1oeW7LgQFx2dxo46VeYN+CjW5wyXBiQlHMXer
Q91RgzhtrhxXmaZdrzxlsGk2v6aaXjEtV0ogVaMAw6O3T8LKPbcRzQRkezBpScHb
TSwxDPakl6I3Ez4swMk5xCPHzIMkdOcuGpr5REM3nuFF0ep1rhWn/Bzmdl21wmXV
L5Ya3mlUTCxL9LrrKInQshGUp7yV535H1vhHSpIYo9T4ohPTFrz1qHNAOepv+zVM
DCWE0TyXMLHDQEb20oqcalLvZ6Kc05kNYbS9adwTcie67/3IEY/lg7okxyyS4loA
hTW6Yc42T2vqUivb+fC8u7amvKPtTNyRIfuIqQn5YWeflFrZt5WYMSG1YaBuQweU
SB1eM0iJCTCMnaImBsGOrQxGI08O8MahITjD46ovFDk8On0BnripWlwmbtFTW6/B
/LFSox62bHfxvZVpkUYEkq2wJoc0Ly0Y/Sfi1AW2RNmPtZ3HjXVRNNUG0mgt7ot4
4KUPiy2wnsrctQjBNk3+KZDyzxT5h561jYiU/IbBLvFkmSUcGuNe/67Em6q4SKqj
HDn6sM7xYlWTkSoVjMD535ZEiK0XFe41q8+T3gn5P+VZOZ88X5ycruMby2EyrkzQ
wNJEKFUhKWTuYu9010giIvijY6LzRT1KzcNkSjwE+VuDtxPj9oezFALunJLt+/Sq
xYAihtTKB8xT/Tr6+io9TduldcTyCXXbkDdERXeBp8q1rtq0hT9d9xDBjmbBk45n
4cA8IW+IaO2F6aK2MpKKKVdSrmBiPU92US8QIiEZrwsi8uZ5gHLpf2+FGUkRmBTy
pWZKhP5ZzS0A44VJSHpMltMk9Eo8FNOHZpRCv00R+8qu2LuXU0VNkWnKX5XaJFBd
5IKUmvR5Qd2/E66gypszqqLADbVm33gxEo0D8P2oD6DH3ZS3EB5T8M5WiluvddnG
IOw7pR1I14+l3pxoA9j5M5BJsSrBuu7e2nk4TN9CZQMdlCSMRYnsqpvLJMke2eMO
FkOGFOp4KTve658hzxQGDUw0SjBPYaQOgISpEfojIICl2PITn47UeRIhNSoBXBzG
fBjuiYi6vnfDhjxlY5P59FQ64cYJbDqNwR2TNmFFZ3Ze1Bv6XnQkXqNqTzyrR8nY
1tSmcV31Ke3HVeQ2u3pxsx7k99glHFUxBifU2RFXAjEcXtEvXX7EBNg+kSXYVhuw
6c/1s+RX1BcjfVztuwvYshU/qYztFf6kDdAzPjQqPJgJSzOnrkhe+u1pRtlNEO9b
ZgsqrJh05WxmIqKjaBJreRVuSBAeTv5QAZ+pfYDVmwYRgpIWcI3iY7tb/eMeW+gN
M7n0+TwY4VxUor7+RuV7FOQwRTAJHyl2TBTPAl06axABhm1jGeJimKlk+ephibcB
sPevceTrDR2nXeVVfuCHLF8Pm+JW/Svfku8xaPkoyWJcM6MzA0tmX+ImEmQCUi35
r1wqW3+BQv361acN42iOzHVdYeXtzZ0LadjHuTCM5qG30B/hph/MZXiiZZI5gE8q
jZeAIu+tSvMtGXbSlWKQfZJJeuJvx2IytJBgmp2SRnYD+no687617SxRdzkDNWbg
EpuvZjKB3OaK1FHeWp/CA2MsJn921e9sX9s3cfQYeyFjWkssq++g+uHHBtkqnwgK
p0SWvi0S1XwqApmzso/BQf41dxFo5EDhZ9d++0X/l8Uie7vvzqzqUHxOr/I/rq0O
A7Usd0ULM5zmMEEiYV43kj/UwKAUBjaVGs3Ug05qS290D7xVcRFHbzTJnJbWajzQ
TnOitXiSbSHpN3zMV12QrYMU+0nvHjy5CmTcyWFE3Ms0mw61i6HxQVsKkrUXYkDj
/0YBFbrkdXyJXrK32xH87O1VyTsETK6d7y2Ap93nLGoyu9PvDoXsrECE/gJniz8B
Zw9V0xpf1du4EUYp0sZbxk2b/kwPeYKZQBO7gaD0Jyc3Pms6JrTb0sryr+6FM+Jv
h2gkMoNwQLNE6mATzpFY9lhlDUUojQKDFVxvIxYnSy3ZMUq0sSzEhnqPWLh7IYdd
bC4zkE2cIn5j8gN0CLyA3fUyeqwOSrJbtFbsMH2/ExVeIzLAqi8grbKpzacOaE5u
Dfo5LOEkFocUZBlsFNeO6HLWhpBp82xs64sy+Y4vrrNJttsTeOPZQsc3I2/c3U/V
23vyyvc7ZYAmRtfwDIu+wM2zLrKU7yO+fPneYq+ayvn9GqK3psB0A43UiDsyeBA6
5RLhQl4gCaYIkF9iAXICiYGBNiUv35f1Ba4t8woT6wC9nOeFfvU+s4hSaO9RSFQh
uqmD9MPe4RI+bBY5DSoZVzwZvXa2H/z/pTd0tecuf0X76BYaFrIcjOcRL8zbFsyj
cZHih52czfcnMctVI+ReGEftw1pBs8oZLSrYm+CsQ3XSzHQBOfwOVl2KEx4W9RKR
AOweRjcSnkWuZ/+T3GgrwBoIAyQ41Gbd8Izh9SYgGeoFRVgqNWoLM/Rt012PYkqw
pJmK33hjyJ+q7uuFU8Ixb/GukDIwHpG/JN/sGxg5a9D5JfSgPeCTNPopKwgo6q+9
tQe2ESJh0lS4OTJLJ/hvVmpFUggeRlpSPMICdPD/qsPZSb0sTb5ZWXU0EabHHYn/
v8+XTd2UKakMVX9uY1asqh/mStuZduMtvSNOm7KT5GZY3zWrvZuMxUMA8Hxq+3ax
+2+PPiwNXlbQ/8lqG+mTov3cpoEW8HPU/H4rc5itQJw+plD/J0XXh9hzAyqgj3aP
kDAGC3OPx0VqD2pq4mgUgGa7gMgIVimFwSh1HDJzvbp/eKmgPdT4x9pdAXpP3Qzn
o93iTXBPizrP+tvw8bHGx2RrI+IDYOfYoU0zKFtya5bZt7sp8Ta6EBC+kXIU4U2O
8AK7hFRAVNWhzE+HtYNaxC30YPLeHRb/EEJvRCHDgshod7WGOPR98n/4lXHtYGFE
ostEvrlMw6jIDOzSeTjirSbIqE5DdxI2kFNc5hipQzbvlDp6iK2m+g759vkUdf/v
L9dv8SssISp8xGYu4D+at6/44LScMAEdfCrfj3grVBqjLxKvgX4oVLYPIZQ8UiPs
0hSykfnSGEcB4Glnsw1MghKLQ12gB6YyvpsI6J6bmHsgBapL8VEpKB8PQ1rqJN/n
ViTgun1Cpcso9/BZHJ93ieqEPUHlC78cjJJwe+P7ueXOcr6Dmd5gPijnkVcYpJMI
jSieMIotySnCRxjE4e8v5VXb537zyiCB/wWAi127No0yrLSVT38XPz0CehXBtNpu
pyU/F+6WI0ATHtoRZsbvc9qJJVgSUK+Zr8GvgPHeca188eEfsCZ96L3d+yWV7mDx
8bPs6zARHjtAzIuW6TX8MqA3OL4GnkCvbw5BBgymbobNKzC5jDSVLa/q9JXmszfN
OT8rgXKqsWVFMCJvnpBZShSrjg58Pqbmwviw9oRVZjc0s1pDPsv98LGh47OykCX6
DLO6ILO864iuU8SYdaVzer/LJAn7LLPx6jZhXkKDrPr5LPzXFB726gInU7jJa018
ZbkLfHnOHrAcBBRDEBm6ggCLxgWYJvPcSJCfWGq679do7iLnsTInxzt4jZHeMt3+
CDUoILFe09QsY8pfjAPeiaWd2RXvQRVmUdCIAeMquHw8wLhW3d4pJaCfd5FI0K24
VC0bFjyeYG5gSATi2EOzG3w14WEf0gZhQI0NkYARHxhw4mIoCWmZVddrd6a8EFL3
tIrqkfFTzD1kYB2vJR7weTg1iI7di36B/Hh3mja16Xc0XzT/LtgItFXyoTGtlb2w
LPK858u/ZntEB11MavItAxreAxsGcZZLzOKeC5scIvOi4a++zuzODmMHN/HOe9JG
M7LmeEEVlfHuITjF1NoqqP2i62FjrEOxNl4ERAQwQOzNlR4bxh+tVlAoceR1RkpH
ACi3nqpRA/Ef04wmXs22Wxwsmq3lgT9ph1rjGpZxIkEV+1MOh6kZTGnvfTzwhfcq
qr5BZ6gDhpQ88WZ4gAq36yRis4CUND7QgyLxpH/w0rVI3Z9eNd99SLX/zWx+nh0i
i+Ct1UwBbVNSVBsgPSuh/sYHtPRcGPrfERKn8Iwrgtq60t9YTqxSh2G5W6+MPlqb
lpVVPBcAnFSLZ2/yZqvLcOUYMvIhH0o0I3MCp8O2Uqf0/x5oubAyLPq/Y1/Rqxt4
0jAisjj6tC8CZYp5xUvO00iytP0KD6wD2JW5Tov1EBiEcwTXrJJo2rfSwFvzLEcv
p96IR2PcBKxrSzuRN3B8PCXdIK7rI2AbRCszpuY4N0L+gFhsi+S2mzgNafj0bZaF
rWeRfQsQW/OYuDerx6M+a+OAXMaCki7m7mBcOOaAJXo=
`protect END_PROTECTED
