`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2QiWexra3bVBwlC0vdlrdo+EwxcWV2bm6P8ukzcVOyZGqiQVNYKnuwpsygon01O
R3P/hZIvphvLql4v1KsHAnJdC+luEgJL62WtWUnxWkVvYy6dezeplSu5BtR5Ve8P
RRcb48O+rnpt3txgL1m24XT2mS2IRlcxMQPyIerZOJRiFm5jblge/Y2gMFlAYmUy
gOD1NNy6XcKhDtNKmDCqLN7xLV0zOKQRsq837ZqblfGy4cJHKmZ8Bj5F+87EnExQ
RGeVkJXVNF+vXCI/HArvTBIOyYE9HOkmsRczz3l9WUENMuwF/i34fDGoRF7gpRUe
2MGUVDC4MBhgbXkEsybjoGx3gqBryfIYoWNlx4j4PhkTcWDkxd6qh39MJ+RJSV4u
hP5r2n/UF/+Me6O96wx1qCxEmzPEt4XRrubXKH/D6ERtD++8n7xRmEYCt+cKwpyw
lfAEiDFHRh2UMxGgGiy1zgLoSX9uyWC96J5UCz3ASeEwRAhIQxonYqMDQjhjNKAO
oNQIgVv3O6F7n2ozP4gSsA==
`protect END_PROTECTED
