`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYEMYrYT+lm6gGviBOHdieFsPUgTpJpxendkwZsSBgbm6XqwlUc/x9CKDcQ4WtbF
ns5pJ04nRIFOtiW3eFIiOvu5z1sWFlpfwWXHxptr4MGwZUptJWVInXvdS9UIeyV4
JlUCrDIY1Vud+BEtK9IwLS2eKe88vjUDsFLHDseshwU4CsmdrSuh5oPK+BtQWGUY
n4Y3rrpEUounztAwv3Ge0ZK+DXKnAj4twLpvrjhAgNhnDupQ6ZcmjSHEBM50Vlpa
8/dL+zodD4xlqrDcHrkaWEtdbLRlB/ZUOnLaQNAB31TqOl8utod5oLEKomTr2OST
P8dW66baS5qoigF2uwzZ/snO5fjUVlKgeByxo42Y2rb57Wq/tX2jBooNZojsPzVR
cgoTSdZ4eXspnJeAlR8lw0/Glvvpq/Szg94BRFVTMOXM9YPwKDFSKq33W4QtTcXJ
hkiysRzQ9kWdL5lBI+539+LblElKPvU/VSeo6PWqgDOnbmu/keWtLbcMeLA33QJI
aJ5YLght/TKzYcw/Wd6q2ECTutf7nNk3iviJhEYcnouxNYi79zXDQ0H/Qxy9WmjD
n+va9WaRNfjl98P4CkP6bp2kDOaPtIl+B3W60ih99LfiokzQb95/Eh68HnIuQyF1
DSskjCj5DqLwLDdWVzlpKQ/F9vFx7ycDIRS80PY4KKAD4M0wLgyhyu96AR084+Bj
3F57lzxsqGw+up3VfxNBMFvrNf2BgySo9heFEwRfOIzlcrNu1ezqHtNdfQR/878h
uKktw3aoBVmXdiC0KjhulgY3rFeV2tHlIpqdXdiEFmaMsiaZYwxEiAWCyUC8oHez
ZJC96JzhvMnBaAC76i/nbqQrV+ZX0T9egomswElDK6smcrc2ziW7EZE9gA/3qO6P
W9CmJwh9RWwtkYhEqJ2Ag1bq3IJKb5jKBCNysk3edVBr9jtCyWF9N5+T1fz9zbX9
dw0EsHV9pJSEOfl+aadOcTOGT13WFPDDbuwQREyg3I+tC/DVAElT73g/nsEmL7kk
s3I0b/eRSldr+MDps96ZDZJ3WKVkVpDWrJPCMV3suXBkgOIuxMEuxgs6ru89PKDp
Yh+/I2BvCbtxzZkEELw4eEFFlVUqGnsA9MAzcu8Fj9IqFg9zfySLls9uI3s+pv4f
RExm4DDAf1rezM15Ys65X6RlejktbgkmLDdhdiR7rryikAcrgDBeAgw94qITOT7X
Y4cC285ZoWLYCmtzEFD22S97KXYTIvTcWM2IPTH5rEN0QBgY6WkdUodVsuOoid6G
4WahdZJtXUOnyIfNEovliIgvEwssYu/kixQ2ssvsx0ljZ5qP1f9llSsGJQcQH8bU
704Fw6Iwtn7x/hixuc/oOyZm//Ukq1m4y8opLBXMh2ErQXACaoGfe2Q0CvOCBqs4
olV7kCsmTfeXXgwi8Dqi3CH3mgPJfuL7i9mmPEzsqb8mp70H+hzVkJDrUfdZJbjj
eXeUub8mbJQ0e3Fc9oeT6QU5w/FTrlX2t8p9LHwPcNsMI65Sw2Kq8ZJ9HWY9STkC
6nkUn6tBxoaHkxXDL+uVmq+oQB2YjWaMMLWAoQSHmQwc3e6COWzU8KOG9sXYtRs+
2wfFaPB3+dGmSjFeM4uet5/+LaUWfHhb/p3etzXNq2gmRgfIGKQAc9T405mOjfu1
3EdGubZ5nGh55x1ajyaHPR2mIuEfF2x6513HDPaKPGVCv7vY9GMbSrO2KPdm9da+
3FrD2h1zRMj1uMbZPnQ8hqIoPoRUqWegolgpeDrz+cyLW1MnZyCgQvlL4KcsRAax
WZwhYZbVYxGwFWYg8st/6g==
`protect END_PROTECTED
