`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h13aU6k5j03INs8Qngal0Mnpln5/zPQtiHYBsCAGsw4l/odBRYyMW4NQjOP0mE06
IFMxw2rPKlrxP9kOcfrRANDwu7TuwyFIdxKK3cXjRwryF+bIja5rAyxSrLI+RRsG
5qHeMDR24VttEfBB6aDXH2P71IMt0LikZ5Y4Oh7xNA/2+ba0uMueacEzKjjkMu+l
pe9i/C9EUCBZJ/sgVWwtw7Mf0m4XMc+pkM+THrH+90VtBcy3MT0bhs3gcgVJmw42
eoj2IpPDewR1lqCdDcAWO4XRyrUy5VC9xXkKClggPG0s0B/Hh/wRlHzV4azdRT2m
PIMRAv9J9NeWtnpbsVOu2CH9Z2VhFGJDxd/OFcqJsl+ejJyaoD+4VzB9VKksK4Zf
C7V82ROj7hpo+tJH6HLLJNr5dBHlE134c6b2ZpBTGoOut86ENx2rmMOqcWYjascG
1SEwCSLQshufk4q0WnabO6U8M53jIscOuu453mI7CcWbSgWN3sc+TjMFGerxXGCm
kj4v8/ESClIdMoW+zmKPwFnTjQ0CKM5ruVQ2t/pByDVkCnbSiAIngxhuUW3JV/JZ
yHswTeKdv0ZfTujuHQT9chCEl10V0+QgkJjhroZb6kRklBDui6nMLUrlkw//sNDp
a2nsx+rSPALV/EW6Gsnk9tAb9DL10NQpyRg3Nolomp0S9WXB+sgxbv6B/6OWAsVA
Lw3sR+hg71SW2jyRV85XeVXivXQi397yGs2OamdaoQAIvt3SN1PZQoaUqseMxH2F
TmnOLGRVHDXYvx8S75nzQ+suZS8xVJG/d8q7dSi4Vg39ZyPbuTGLidcGBku+f66U
7eUh3BGguW+AoyDgT55gJj17W1WUveXGjFX2BjpWvchA+h2M24NjD0hNj4j0SLBv
jMdRBCrNxmTbROuIBmjmREobY45Ox3VfqJUR7uhKOzHj3K7AW4sAH9NCusNTdqk9
U0R9ICtiL1tSXwyE6m7MAyBnviDNgWi5pXoZChukPg0/xE1SN7LiRHbY0kURvCVo
KNVlCGYokPjYjF/3MHRZtswk7+rvbWOQEiTb+UIrjEnfYQY6Y0r0u28vwXw4x9v8
cR86N0jrwxV2dLyEXLYjNyEhqJjPOlAgLKr1HmnW0VLG7d/K4UlDNzRgcp6yzAbR
hlcmcODlgh50oEjDylwrdpSrp1rIiXdrS6VK1hBikO6IGkIlnbMAJkFcq3/oPwvs
1nXseFzMgq348/7dTjUQLDxhsrkoQgSpZ6CtnMqqZvyrz1V3+y+zwgTct6E0GkCk
nfe/Z1noqt8VeqVHA4zaY70LWwtsyrtJFKX1yvaKltJ7/EMYV2GWZW0uoEiK9mjw
Q2mEcd5yWwybKCiYlsVq/LXxejGoz2eK8Y1ugFCU3VOMBQpdz0eihWI/50MMzA6N
TEAVoyVlYOS6Mvh7TnVgqlyqHrXRGQLCXfwNxu++so+L5u2Q9EHcGdVP1ZklTnB5
BLus1C4xDLA7hXvZNEy1qLC7WjHtZ55bnsyX723iWi3+rDRfc85zfLEI7480KG9a
8vLaAhYkKFJQ5su71H+/h3BFcP7uwTY/47p/g/NdUY1kdkZ2FPFi9riRpZ+SoBbD
6cEK6XkmWO/tJyu/pYamM6qsjXMPZQQYcH6qmEPRliERpDkQ+39r2CzH1Af//F/4
2SQxNB8KzUKtOjeFnj1/bI/O/2pjq3NhWMTjBORitWKP24rApiqKG5smz71xzcqS
4YVUJThxkRcvy1mIajL85vgBYdcX67JXEXuW9ATLwUr/ps0qEDu2C4J54FIza8Fe
PT43/RdiZpuvXRqUpQeBP0o20ONX9N5jDV4kvpbPKNyFChAh45fuWX7vipz92U5w
bCeRnXCdvLGe/cmWR1osRDGWJhxMx7Ceaip7awsw+coqTmlKBWt1UWM6og03C97i
OPuPYwPb6EzQ7QTbcOxYtWNAtr+C04GqR8MBCU7u3MvX+8QrCTNhDYrAjo02BhDn
Uz7K/C2nX53WXrI4QXvT6IzTLVrgKgRznNzMhV2eC0eFrveevvqG34QAxUr/4YMQ
QD+7999+tsxGVLA6SQ6PgZNmntJ1FNGhzD1Ydx5JWGodN/GblGrman3Wz7+EmkbP
VYm1FH5JuFstrZ2S7qVRCdIrvoUQKdLikbn6Fc02rOeIWV9UtieChoku6My3CXsi
nqzLWKPKQKC+dN/6iUQsUlrJVcs3JkStjHr/9Dzi8UzOshkJkmANT6+oRy6tm7Mq
/hYC6UbCEWZ31XsuQRRvtTWA6QlguAF3Rsx4+4fPVFOJaGr1VBeb0pZjMsWpwBXG
PJOryJ/5zZyqQO0LPcjpF8Eyv0SKRSS/nnV0xLYvKL1m9Et/VK8ky+cCQHb08J7N
+/5TpyvSoycNHQRtLnk9L6N1PG5Nz+UJNWMB5D8szyaUGu1aKaULFqidKs6XcGTJ
/bkeVhEdqSu3B95NYitLl3mE+V/iVTJWVi2OBR7s4u1vjMeUEbVF+78VLbOPhHX1
Tq+9uZGqSp7aH8LOkMxiuZRI3H7UjCKyyaKFH5zuXgoxjpj2mBiR4uAt2FrF5+YN
eKL1Op2d3rWHvw2QzlEdLC1PxCO+UI5u9j0pmdIT65geXhu9QnkLchaZ++3bjy39
hha6S7QJhd5sB1jHPIVZF550bXIwq4MFusdT07XB18+BxWrlVk/s/KyZlN+HJ/5p
GL+VaTUueeb4lr8VGpPwi6i3cN/Y2WxKhY8gY5dBxjkbcH2m0Ey65yFU8G8LsKhC
jRFBfGIovdhTkGP97B4QgPfjZd7h5bhtcpKx/cR6Klw+WMVPTBGFLChonXUSfFBJ
dnHVD+OSl3e8RsTBpT46l7l+3zh5WboDafj+3fFDwYhL6JMG6T//vKry3+z6QwQ2
KfAn+9LKqVy5VcXMOX+8hHSgs6kac9abBbEI2wMax0BPl2qABHUvIZgRcmQwybmh
okm0jc4ufq3wwYQSp4lHylUr8xAaGcN/06ym18G4rNCF23Zbbc/6Ub5224s+XD/V
GhnrE8j9Fy+nGFfMSG8w09hNYPC6Qcln/Y55+zCrpzMPkl6tfLj06obdXVJqjghE
zRD9b26ID78OkAGBq2pkLuXERlyaHV4vqgJEKWjPedA8OGPKD01T4xO4NK2+wS9R
OthMgn+Bz3QFsT2dLQQEAXu/Sx6hTmbKmleCb56/gk2n54F29LquYFtA10cPoC3k
idVBs45Efr4UyF7jv/K1qCzAzb2rB/JBF/+y6TqjPsEbzvMhVwqLEElULCnf+mQX
kSsuhqVYcIAnKxW5Upn4/eHk9SfVe1aoKW9VI4boO+GUlzLFqvqVhZk9MmWLkDd5
1h8kWgyeNQvBPaAVmhACjU+XIf2AAtUSKJMgT/xiaVXKMR8xnd8xTSwZKRF6QG4I
65u8hUrEUTKWIltUkPYjO8u1cLP9YWbgsPcig5JOACi0EiXnn5RXVgVNbDOZopHJ
GV+/E01QjIdrKz2SM4oj9tVlQg7liMikA7tfwX60J4seqt04OVIFGpZGZLXjsfn6
V0b5sKiL3VUmxTu8IUNTQIwo+dyYHq7HMmmLCD8a61fIpH1THthcEw+mnWtP+lgU
tlZyg+swCkj+t8n7Nww0VNkqZeBNbA7OPiDkELacdm0JnOOv9uufoJGgSyTwtqmV
IUNYUEIjnXmbWguvaiVq+cDTROBYV9vidqgQ+PEEclRY8sNm9LHmG1rcVYiW8M9L
XzhDGSn6AdqQBQnE38EHMk1pg9k9PLcCmj7Xv99EX3m4fzm4moLf2c/BV7DBJlvQ
yN3bdnu295hddKMvUcOzE36Kt03fx5C3hSor0nbbmt/xZor361Wkwu258GV9O95V
ghfTzpzFn+1FxaMhkw22YAXjG1AaFkzPnTSU7rsfhpLvxdeqkO58JH7iQhXn8Bi4
pjSBgFtniif1ZizQOfMLPOYf77aCCWbbnwfbfhXsQRLjXVjqWS8YQ6MVFJW2ciw9
swTcW76O6EG3Vq/T+yYBNviBJa+/p6SQW0UtT7jh5xrUGKKnroj+YvEYWQPtS/9o
D9i5oVn+Ds6jhfrFVVlSt11hBHyg2sLoBFDM6kUxcZH4npHCSuYkcYjS+NoaW7/R
tBfJKKHgd6Ug9yW4aSM7Fn7WkVOXj2sAN1si51mCMyFi/YcoO4YxBypdTkyr6ukl
kY6Irr4QATFHV7BJOEhXyY63BIDvxsSckX9t9cNXJoISjFCtGhrQHqtomdDklv9/
EL/Gy/pGAsS/5vxUk2u3eKbB6U3JrZHW/TKe3WG0u2VuUgbIWMAYKo2kBeMdsIdh
/2R4iLWd5xN009tEukeWTvR0EhX7yKhrIEiTOZO93tLXCvgmzrEOTTb79TzdcRVQ
28LlhJeMaDL9X3TJtWXaXKrEuIvme9f/lWfKXjpzHXqpc2cz3kx6QZOV65ehUP1K
I0ktsbCSlQ0LznO+oIFxn9n0TAFuNUKItUcUj0eAh/F9+hHywAOY8154CBvCaWzO
oEKPa06R7yB+6UUv+8EOX8Fv3213zTqtwPD4bsoynaSUpYAme3xM873j2AndlaTs
GQOjzOh8jlafA/woMkZ/L/+Wg5m6mtdtUVru+i+Gt+HGRYE5UNg6+rllJb+XKH6P
Sny6RIPzFKKwPsM+G4zE1I8zkyk8TRRcDcceQRdArG5yTx2H4h0i7HqtZGQEGaHR
PRSTO+6FnEJYkXEZPSNbpDA+EHpYO0BfC+enSfjxG8hVNsOzWLl7ohMaulvMw4np
T9rFFwHOvEu8fMzB8tygO8oGfPDPPnCEeKi9CH8b1FgwQSqFQsn3rUIscJnELhYT
`protect END_PROTECTED
