`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7LvySyOhzKdEe4yCTDihh5cQpngpQDxZTGyGjbVPjSUDsDo9Mhi2Lrmpn8VzGHo
a4/OddMDNiKSJsSIFh9/HMJfqtysQuBnplSsTWtX58BzO2tUeVwpTN5OHGBnJZg7
sI+MRLWLMEd2hNAOJ74XbRKSNIPmnjw5QzU67jn3RrgdG6id81Modukpd0Klipup
llwSuq77tXhHjn7fbR7jh0KedE95zpoN17MfNC+NGth8nn9aIVlJL5S71FNYFxc7
fdSUOC1NH1X6z6JhZls3x6zvfkizWI7fnk8bV9wpVM9q72fv2iSeMce+pb54LZEV
g/s8DJHCeMwOxpLWPobtGXEEUAuf/hIo5xD6CKdSSMDzLYtwqPJJqQmt7erZ4ARQ
N3zVUqsbcpjR80jlhUQ7mqvtV/1T+5hIj8gJMFW0VGCmGnogjpRM49slhbi9GZW8
3DKr/Nk5e/TzO7f0skYzztYaf+MJSzQqFhi99kYEnM3DgJRbegb/B5+pXhjRN1d1
ouhGZqT6245vhLlz32fiyni1MtEHmE+OcJTwYEKkeuSPWghzR0WXro4ypVcXt7O+
V8yw/A69eGwaK1+mpKCAgnP1Ma7tuC90qugn90UdQmbFdFYVYhyGMNy1g1O1Gfqq
LKnQSEe3qoTYAdMvUreaXhWerldrM6H62LEfNY/K3nPQZtznts1T8ciMaR/HLovw
Cw5p0xUisRyNsngqAjdDJwUXhohOL7WEwVq5BsVFPWOh3O0d7+Mo1laup1X88U9z
r1zj+V845O23lGF4yKxrqkepRX6cJZ75919hNximKwG6NmuamNMZ9cbSJZ5tUne8
`protect END_PROTECTED
