`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SFzZG9JohXflQ7w1ci8XlIROuNZkJSczRin5Bp0KWpiLMeFejbUXcbHwT+7Nbk1m
8e84Ko/XoZ908aPTUy6P4vFoqQippYan26qjMYT6iKS6uoD3RGeb6uCKjJSpK76a
seGK+t8QwIRLUEjjPVV0gaDKXGA0esvO2fmYT7UEZm7be90N/g24UF+CMMZ/wzAi
MoOwS25B/LwRjTCAGG9OnYeQdB/KzrXBqM/+hTp8cCNYDO9FALSBtSOeVEr61+WF
LaI4IHJRbphSZEcKYxD3amiKBtCH2jNhx2JnDRCGwURHmiOlhcFzjTiI8cDKWgks
VH+BWG462N+nAgugD02AwUePT3dpeTsvtBUnLeygYTze9O+xS20fd5up7TjQslS6
cfmKHXwfCUH1vww7Xccuh9uaEM6EVt6tVdmnVP/V1XgS/q35SM/2BYxEfhXPZBey
LvoSPVYysz1G0Wq9z+7Gxuc5wgNUzAgeQXhtg9S/NPYpeiYwGgJagQhkVuQXe8xK
jAvWCoDMcghUQpovYCOei5PhQIFyoUn714u09w6O8sCLTiJnIJSqBvC0cqQfE6Fr
FmacjLULVz/PX93C0mDro6rfWbP8FVeW9idqrCpIqOHcotba7fjHhAeGjcEGq9Zi
EeCz8Lf0JXw8x7PqzZnVpBJ4SMnOMWEifF/VDFXG4bP6XsxzgOgD61h5WdMLK11u
EvMkUTFw6fA4GzHDH0NPdcAtEViER3hB0WumPUpj1b5ny5jh0Zle0FVkmZiy3FK8
jJXYNy52yArzPIELpCAK0AxvtfTTKLihxzFAufKmFs7l9H2NytItEUH/HlOQRua2
UQRVTS5Dm2b/2qbA2U4S3uFPBnRskGEi3iO7zZVpvFc3KKkHxEU1kcwTFX4DZ2k2
OKvbMJGaTY3jYnq2JQ8j3PhPr2o4kVYvgsNnIIVkiQbL8hY9iIv4YFAuIvJY0Pmc
pmKDf3UD9X7B/W2i5aghduL0oyMs26ztYFL3r1ET5dKy/M3VBK45QuarjgEBx8YB
u7RF0L8KEHrM3YGDWh5/tKpNZ1QQv1dAbcv5z+HNfyd8gN2UPFVME7HbJHYOeJP4
xaaa75BuJZstTYek6tns+HN4IYBpHeNs6+BgPHAHfUZdnZZsQQ7m82gMDhQLdMj8
`protect END_PROTECTED
