`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cGsJ7D3+jLJRk6lU6GsgdlAc2VuoZxRi7xD0U/jl84E4PnQChntz/manPkxBnw5b
7IbGF0OJ+5CYUX6kGCMGJAN7yu/6pkyCPQUktZ2CvujnIoDB19AgjL/DNhP17CQ0
o7XqtjubJddv822jzAWpS2SoYGX7M7C/AHOoLq40N42mq74L159E8iNmnobbMI33
kNl+DR2IfBp7ciTrCXL90eFkZdLQVsmPRv0/taxae+dRpD8DmgecVdHqWaoZpfQ5
f03Oa2XJIIxLrBlZR/RZXhCocJFByZ1cXpXkW/KUjAjhaQtDe8t04LTqT50635pP
cRkqW7HpYPACy4vIDIOwvRMNIOKmIa/r1Q1tNqEY+04NdTi6dRVDhcfBh6a6uFn1
NN9+YDJ1MavTJUCh60obJOH71rIAkG8W7ioeWnvtXrJACnWajTDP4SxvOBAHtPVI
XQvTEoVR3og1bnOXkkrgk4ZNLHoYaD36leMXBJdXcXxjyhoV07ohnmjRgfY8zTGO
XwWIgHxCPInIrjdaT9KHzzRIH5zdzVjL3kL6na0dJfciBxlOju98dm5DgPgl9mFZ
okSrNYs18txAqlArXVT9znbABJminU5iPuaCAIIxJPGoP0SBbYG6vrDf66SvdLpG
yj8OYCp7+KfB6rZZZCcskUCbAYama3BKe8piVLaeInu5sl1nPOq63kgprHGTqBX2
Q1bRqM9TgOzAwfqPQdG+jASnM1mj7WBvCecL/D/KzzsEe3YDCHUD4PDgWtW36dAV
V4OgMIGFhVpREUEJT9lJIqagd5flQEO/02ciplF6vLI4nEx+uFSkb44Hk6Hm2/H+
fOlDlpso32lPb72eKjtsnu9YMI53o+zl/yyH/DbTQVeZJDb6t6u8RcAFqdYZzar2
3gX2f/13qAIifYXmXVgNCmIQNm9lU8efzUiP2x88XMfEVhfwdm8JyPVZassQ3ogo
An3fPZ8GhPNzajtarc+p8Zos59uQyDAytuS9bz/idy3pWeHewetoY7duPV/fdBal
KMTWJe1QbUSWWL2nPBNt5EA0r1deQ8M4DinxAzzhSL8Nm+CjpFCl8DjMZpUZ4gjL
nUFayJsRsv7NAQwQcbn6B0wIRE2FmBzcjEWn2SBXrE8=
`protect END_PROTECTED
