`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byfsL1kMHW+VUSzul5L4zrd43baEr2RPp7Z8dDgtHBca004ev2VqwCr09v0u4ek4
hdmwp4K+SBt63wuNplUr1DPYX9dVZfwBevFzlEY9fdqVe3h1Y/GQpRgdaDpvfHzV
zGa8+q0tDr7Cj66H7WTirZoOcta8WVC60tTQZ3Yjww8Ec/igV35VnAr+aSNODAWW
/G0B6XIwiFgBp58hEC9Kemwhqo7AunaPHndKSuCvEX1066ydqe0sDa8fIcOWEM2o
AMVkSxz/Nx/VpjADvauEd2EV0uRG0WMwIpLrtsKCAQjl++fjexDRZSbfextW+TEo
tD5+f3YACn54N1DpDWBAQungFdKQjaqmf9UQqPRafkZssl6YX+jv5Q4Ncfs6ZBpi
/lvj4wZyJ3T74yKDe6GaO2ZdcKAAqAo6JwkYxpVzSRBhCtV9ZyWyp8BPaOpIqJej
qh7QWuP7vdNusNXaKhbil3p7gyeHji1jA6B6/UYlrPoHsoxekshEOASMstDe/7nC
qF4c0iB+4FRgV+MbbqS8nJcuKrDMPM3vLA8RKX0LVFzE9hCTkpT/1OWdanXNHcke
Sx8DuYEb8JWDvIsuy1khwL67uzqiIw2ppAg4rSjNmAm1rR51BCy1RKapU/4yyPfg
kB+wUhfwXvQznKJ0qjqZFPu1f+WehpeIYAX7GhJJyYGRrCR+ssCHel7ALhVL6VYJ
`protect END_PROTECTED
