`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSGyrZ8sWXq3Wmxw3KPYTfN9OOz4eHinGtlHocgHJnadiUQrHNmDiQG4R1zN1b4o
YwKNIyYfJuAO8/AdTdkDF9JS6ObeKjC9EUBdhGhZC3NGOK6c7nH/dxGQx4BNVx4h
H1r1i1BD6gRH+fq7qJp77fxOFDKLfU2USto+xM/fGgw=
`protect END_PROTECTED
