`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6grpUQsCQGeMmxvO6Mm6TA9d+rhLXkQKdlPiFBSGTa+IWfEXLWIGPGKaSBdiKvR
lkqv2yrwQcfxcE+LXxrIm9MPUfUG6lltVGkLGvPHRkVR1ytW9DLXWhNjJxk4g19A
IZF2w8x0rV8nuUvqztAO0Hc5RrdmVUDDp+RRH3FgWFL9uDAF/WSS66NWWtb33/sB
eRt6GIbpJy6YRv+AARj2ldFsvdyfWt9WmvFLab8e8pDUiq80owjriiuO3fo1Hjdg
jK/sl0XaPgkbsi1QGdKlSfwe58w5Bc0yYkLRazQH7SHsPV+ysH4iNCaBrhoORIP+
dx3glLCvnkGuB5JPnXR5Bn8tC3Q03gaHsgQLKK7rDBb0Vs9tRJuRCIVGIm6Me2An
wTx24QxSRqLqC8vmDWow5kuBLKHhmmYESwynLEElsZfczl/gFPJi7rVx30djx934
OHr0+H33nNO4Mr71sPLKpAUGzKs/XnE1PEExZ10j4wksVxGAWz2zIjwjaGxh/ugH
FLE24Ekhn29xNcJQd2dlTlmOuHtIAFVmyuZkh3Hzl4BlMV1UJkqHoqoDj2+C19U3
reEdHNmT+xqPKRNjjJAR3bdliEAsJekMeUTDQt+oL497M0zElbvDEDRwd2Aw7JXn
TpEEIYi8Nbf2gE21pCvKU7h+C0O8ogqnsOPw4GjSCwueBdOsMm+EUlwgT+7M/xRJ
yuci6wIAT/d8GmP7RV4ePbbGI5NqbGiuskFHe2A3E6/tQhbcmWM14KxNWAxO0D3e
GGQ9dju/+UYk0FMSHvIoqW39yndckYOz/kDEtBB4JxQzStJOmI8PG2y3pMzHzrQV
cG2aCP7iVHT0zv2ZRGDo+TnifAYo4CPB4qaU6X174XWYTSVr5QNsOn6zeY8FcE4x
E44bJbSsiGgSPtgVxVHUDDluYMQWIOPp1IAuJ9d8PlCX+yfZVZn/N7XY69kDCUmR
mV50V+eufnY6sxqHfRiUuFuyaTcLBnLcSddG+r8PZOmDQWDxprKXJpcMdwBI8N/0
81hMyek/1zLAlhpMhxZyy3MpYjXCI3h4P1OeSQ//Kxs5t/BV3SvEwAWVrRKH0OME
nkbFcYrP8Pih1J3sGJ7diaaHNPGnLSiK/fVV7zdJ60Ex5FNM7+IW6DaEpcP6aBoI
Ym0PpTMBtKU4bs9fEF+S+G+0lFxbBEM+e1tob9ekvPQA809vH0IxSQPcuGLKjdIp
7DVpck3FBjcgmRCvRsDsmtzIox+Hq8os7vz+kxmMJz+dMlDk0AzDdt6TmpQx+IvQ
T8kjRBjXjGdl3nsDS+1FnLPPES79YbRjFUeEqm6G2RBbM43CbR/HvQWrkCuCbunk
D6T2osd0vAwDPXsKmFETJaCmVTQZWv24TEr1+yqiSv2UjA5KsS5NRH4wUIDz2dr3
1NGqMHln+WixVq0KJUUwbPcmOFrGXIigiQ9b0160cNPLT0HbRl/TF9zojh+lvvOb
qCOLP/JEkrhlhGZb2ovamregxAw6DRR84Lt/bUetK8siA+n/YfCJQ2QAjXDR4LAM
jX3hrgAIoZ6IFMcoU+EuAnPsYAjOGasz15dDcnbBuVTZaMO8tRYtxv8atCaGYEK0
nXXzJqnUYjYftCyV9ByGKcZHTd45aKccIjEFT61Zg5k4sLt4ZbJw7Z2fbCpL9DUl
Qx0+Ys6AcM2XXpEY9THeTaBMQeB9ggHtey9JUyzc//smokKvbc3AzhTKkapll1R3
IxfjizKIMRjpP6IWgjpS68UjuiKlNCy0hD7DT1EfJiWW1FqkmKiAzyoqpI0ZTKG7
8IYj1x5DPOD9hSa62I4/vyMRauAqYtHIsBfmKHwTrHH8+ce/1gPvr5aVjew+SpcS
7Jami72nt6Vh/Tjr7++7Nke1bmQfvZOzuOmzd4c4nZSkroaxaEOg1F5HkQdCRTzu
RDZH/RD5Ws3ROH+Tj2Q8HqSwAVJnl3wumh8PnuHHJXF4hQKeKiE48Pi3CSkXZask
qPuZ7qEaPvqw+LsZpSn7HaRYA9eBHrt7mNxGoW/G/GOL2GF8DxA0qddaJRArgzNF
2z9HsD3x/oIqxFh5b3CEKLk/8fa0zQHouIanHksrc07wtOyDVKORrCAxSrRMaQ8j
yWc2trDXQHfGAqgFTSCTwnsGJRW1U3ZR2t9YzSFCHGsjyoKEuq1fnK9xHd7krQYn
reC4RmcN9/h0+o28OKZYUe6atT6pbtJK41HRUO8zLcDEtlJotdTjVzgJuEOUZZgV
87wgottqt0KkksTwDG6yrrENsBIJ337LbxcoAnNXICLXsZL7fYrtX6Rkkvqkn+Fn
6YvU3KQwlKzvlYOz2fWYhx1pM5Y+wl2l8dNmHUyGURVOBUdTpqF6UBN6jZzcsHIX
XYNwGTlsdkHMOAnTTvvESfeNiEy8yoLrIB8zVK+rFD8+tt+US+P7H1BpOT6yn+2k
wgRrywGK/SAjMAe2xpwceNBskCvMw2b+veS60krmZcVsbFtlxzSYg+Hkd3RmFPuN
cLBAWW7v9KJZH266nBMvkbeH6iiKm2mjOGpqBS1BMA6Kn7AUh0vFOQmW2QIBLWGf
0Y1ZHY0F+PtL1OyrxbSAC9MjiFz1LUOmerydFTn53h8xoCGY4YBmf5iTaLFESB9W
Goemt6VWaqaCSvDnTqBStD31LD3tH/Zf6rRoDpWgjx3V/yk9VZbMmJZzaYw7MMuw
Iead5gALEqIRlMN9jKc1MwyJOKoQYvdt7ddksymFtAoqqWijj1F0C8s5UQqlBn0W
/zFpX3BwpmlMGC2htKVToh9ujrTpV77KK8pZHsY9C1Yo/rfbtsxnZHUfTvcA4kiv
nzmXlmy5nF5LzleTQZyIHGuRX6ZLukZRpiYz2vmic2IGFmoM2AXpImYLJUg4NSiq
vwXUaNkRmlhUeWtqqwrW2GmdQHN1pl1yO4j/M8J37uzrYxKm96vN4oIHeN8SGO9L
bRNEicuN9LNw9L3E3LwmPJD6nV0vY7Mp6ZrwHkV+Cj6ZzBHlO9w0BCzHKKAC/r4F
teVmzUF7OkOZ9mCpqGT/KeEJhyh6pZKev0h5jXdGdRti5rWhU2PQ+3oqTMjMTiCt
wn955GFIKekhdg/2E+wbas6hK+zDpExYrnotdBALbWB3KkDg5pCegvpSSaJphanw
OCk9qi5nVIKVscLDyYUtjlZ2KBfPcqlElULxKv3ZvlgqdcOWpKPUzXzdAJDv2qx4
yGKZDogGQuNnF5dN8v7vS8I8NMTMgR0NyTJ39fyZaSKHLmjdt7gJFkxJQUv1Oh48
W5nOLYZ/whJoB5jhWCJPaxFw5e1QOApiERt1R6fG4fLbzn/mHlD7K6mtw0bKSz11
YxgWo4LMb+l0FLV+29pC8sbFjzt9xyEUTMMxVP1qjTpDDJSAxzVueF55friT3LPb
/gG04qoKbxQlaPwKbsVTv2/YkwM6VPtRbPD2ljyO+5C+AKGAh84BdT8a4HcXSOWQ
C5EPFcwJpi/GhPOQAT8v2RJB4y3opoYHg3WDAoSqf5feYSPj3SlNbAeHQ0JLqxoO
3hlgIYrUsduAXY+M5muHo86c9Xx8N1k8RXGGGSKmcI46oRp4kKkbXPhEWUoEkBUj
3vXJLsum7Q3kWgT4Fziqt6YT/lxyJFvloH/3zfEFOYngZMBpRrq1PPcO6kqVhi0s
hIWXlwotsurnrq7FPpwSJF8L4tIjc+8SYcjIa76YwQrJkXwHRdyoCzyaaq4YyIWR
TIC9rG+qoHT+KZe8XvfoPEZALx5kdyJ4ELFLtY+2qDfowQCuqxeGC3GCmkx0lxwl
cMseeMQHGL3cyb9onfVNNbBl4Kp28ldKoqdsQQqWBTE1qT7c9/7FAypeKVEQJR6u
6OiJ/WArGBhnwOwwCQPJl0BP6RYIYN7weSiv3NgJNPM3epnm30yAcidZJMW2RPag
BLAm3mwMU7Dcvt21c282LDKbsVE+QCtCl6uvQn739fR9BfOwStcxfMjI2sCVf1AR
1ov1gYqx1d7Qm7ulSZ0rCalBEueZmvCx5OPcm8QMm7HF3HReq/OhDO3zfA3LRgXU
Ws5X9knTQokZiIvfNxk6V9/u0ceqkHSsIDgXyEMYRJYySzTIBMINJ4NlXYxcHPCH
Ji+y8lP+89ObnwpMzevETFLeVrTztv0OPMSqXkZ1bPH5rJkrhclypXvAHcpUAHOE
tYVOgrGlz/jO2JrB1shMD/3+FdVWMqCDonN0R4ai9L1B2gtIzRhJSZuD2eSUFSjT
34A1aRSDbB1JSLWUkJ529zMcb7WMLwznSv3JiaJ/Qqubs99tjFGObNQwWgn5eHql
KWqjwt0isxgj3OcXKpU20+VQA/FIglkyfINYZGcKb8QvWpjRtQmcgy4teGwgyE33
jgF/TVTxWo/nqQoBpsDn+Pkoz3bgPai40k3sM8FekISfxTjxX8i8HqSNHMH+nQXV
tSVVOgbvELm/Monn2m8YZOadu/DM35jedq2nPdm0B8I29IJYevYg2l5qqm6aGDaj
zWJUFJSiaXoiyvDayWn4JhOOp5smjPqDcYyngbqtf+CIZSJrLCy1IA/obfmARc8Z
YGhuvFya0NebAtEgSSRfUaKv/E8lUkk5KjaknklAu5Rg996rZ3iUijkul1qh6o4c
eLN0a2RSA5IRx0KBmac9Wbnp46EvVAHKlaLCDvKi2RBsnhY3g3wncSU2/0R7fCVy
5mdsScoBb+2HjgaatX9TPmqPbA51D9Vt6oFGdm82Sg84i84VjiH7s+prlJVt1Jc6
DEoU4BGHjeb1j+0oK7ieE9f8cynOYNq9WlRXmFk5AUmjfgxW1TE/Hjl52Dbb/Ex+
cXsz2UlxJyOhdZ5ywemoQ4IKmdS3U3Yb+mUvne7J4NTeL4bt2kPo1s0qUPdnYEmy
hI989hzjvD9ZZW7Qu1r24wXYWw8CUxvhYb3CenzS4zCqiRwbjy4niLqQOFD5+V4t
2q+6sN1XRzvzjiXciMWvWLPre03+IIqG1kBoa3cv2/WK+647fUAt5hvIroYqsXwS
hEro8Qjgsv6pMLxjmnZipapZ1YxIG4qBOJ2cw3o1eGnYIQj5zbOeHHiIp98bWCAt
HhdptXiyUwwLFLyMSnKibKg9/ZevVzpOn+8MHSh8N9uXQq/f2Q58e6UMKCH4xFRo
P0ZoBhUjlD5Sslyob3monHzH+Z9lIdhpCZg7b+orqfiIItkAX6IcEdnL/mJZrwF9
N9He7N5RmA63EyCrgOdwYRnLCmUohL/BsEjUDsa1ATnODo9bMHpZWR9OetZ0W/+r
8Li4Jna5heAKMVXv9FI3Om7fkh2xOJKPcsbovbZOdEr7uYXO0vDJQCyytGgxdkVv
e/1012EzGNFIE/xjPk0eLOFCx52xHC8miy2vFoBJGhiXZ1aD11IFpffw9QJxq5KP
AkFyh8D37mu0F0RDqN3i06xU73Z+jx1hBDd9TLqUscmGTBr9rz9tgxnRw3x+5eqz
hW+2vdnLLViL+Y3ueg/1INlyZo+su7Udh2Cb1TQ233YHyR+v7FLaH+i8bw+ROjBY
I52pkPKMFRETfWPAWzbNJ2IgwUSlwvEbVUSqcZUYXlRiDTEM7i2XSxp7+yRLVrwJ
lL9UZ6qJhcrmlxUXkavaJXPjsM8dnjq94+yYOV20bqvUU4cF4GXuwuLSD7UKeKd9
Qh45gX4gyIsUSeAT11Mdnf9PdTlBMGlA3s9LcMjT/oAiNl7Eqy2r1Opax96ZBXuQ
EoNj9JroGb57gEuowLn+L4spWPHt/1sZas0XcK1XskOgj6Qh4KKsKOshILCTSPgA
HHqvQgAwoHO/lzLPOdCdhx6rkMkdsUfEr6T1FzBvG8xFirea3ftoqSbFmzJiQW12
nALdmXnkEpKnZlrb/UQqvbZfR/+nAIssvao4zNmXLpcm1GGwY2zJ4FiPq+jtOMiB
xixkgavAJRnTrOHdpWjBEvxfga0DcI+H2Op/3S60kyGnNz3X+6kAo9RHjuzdMRmL
DijlXS4FRYJZWk9wh4wkypMJrhfdXfyv+dyT6kEuTMIWQTqRBozMDj7KxsatuTDl
SYZGgD442RaG1wQRvoSaPfW56cPxS/xe7wrcwMqWZowrxFnXXzQhlLP8G97IygPX
sdB/XhBlN7udCzLkxNHd6YpTAcSTAGMxXE9vqkhHcxty0HTTt90PdVAZnHPs0DhM
bqQZIIrzNTAPORilYrSi5Os9mhoZf2PdKGlOBUwp2labk+D1nbw4gYQbQAf/xwCp
6uevSVYCW6l3K91mjkgtY1UNFbgcoDOdYxA3W8BwubVH3CLLD5GL6faMOOqKierW
7ZRjTMNhGUKkI/9CHmjxHjZuTPDTAs33tp2gKh2l2t5fJt6xdBTzKPTk+FQSVaie
I2ZY1gf36Qcr1mnw1y58YrOwaru0j/djamZyVlZQZ+Ontb1CEWcsKYsc41X++cV+
kjDvvmqsAMuwx1sb+vf6ra6Cdv1v5Im+AKxz0Aj89G8YIxR1l/IYnL3ALblrvX9B
GyGjBWgu5NLlit+HhyCsz3umUe0WyUiwfkyyTj5i69Q6c8DKjl0Y8TwCd3j2GLZ4
HYwmUDF/bVoMYKIRG/Phr/d8y/awMrowNo4w1YhABXIYKAkzauVC5BgqHdPuAV1C
fmOEags2D6Ie1St30/NgcfavTqWBlMDKcrLaw6p4NBKGxHFa5S6GBbqIlHbw0JAZ
aknXYoaWyywpe3ONmrMRxE2HsQiMBl2G2OIe0kolqF67zE00VCxbNqAbKoA22Z40
H4C7+TOdzqHRM7+IGmEW0fX1npBLUGOf9NhhpgxziBkmolgkYdJPqWIVRZ1VUE1o
KcKyIM/vaM0dLywdA5WAKTDWHAWI4dT2piQPvGojj5ADX8RMmznpHQy+6jOSbxV1
QDPLLJKtfV0zdpyNTPDoZiX5fQKzKK6E3s+Ln9Phf/xJdjwvBi2FmkMCDNr1DL98
E2F+M15YxJ6RPVGk4/YO93HQGbCztmc59vE+eOY/OJuIpqGEFHZ6RXspSW61pWXn
xLmKmDIf3JhiwYC0lu4wQeC06vfNQRgG5nvg/sL042rA9+t7gKaSyLwY655tNwlA
e3PFy4wMVeK4ACL+jKAnGroW3Z+bOgwSCv2xaJO6CTXp82yS4T+o5/QOL0paiiWV
HytJVXchTRdlx7lbD/jAz7KNxnytWP1MDmrIlgjRDW1VHAPYQUCG//1c9VVN8hX9
qICGsNm9IjdV1+y5+6HTrtNQDRFWSJvwUsrPMu7mb1rnARo0DxWMzzdVnCs/Togb
onipjrgahpI24IUsrNlyJ+rlMguiPuAvw4Kf9ymOfFGpRvTE/XdHLUpj9/seaoP1
QM3aavR4krJjdzpK3sQxGxQfywE/19Rfed2p16og3Un6JEm6uhz6jhPWN4neAF8X
Lq8nyONU41Ngg0a77fMwpBf+tHxnwK29bXKoa5KJIQCmNVvRPgZNH/9a1vJoOVt7
esOuWMO3KACFeWLwytRwQGeB1aEa9gZv5ip/iCE8MFGmxyUyxV8vzfYhx5kBDod2
Gq08yQ8F6sDwEpbwMSRJC9thpsgStTB+QjgsyTPv1UjzHfE2NzZgcqJA9bK5Msew
QaAo9diS0y20iFl7RWXIJVjeyW+qCEpeOf9XsGcfHVdnxkg5tuf9/ZnRRjRT6N5/
8iiRlJoiPTYtz2o/Kr4xDvo/v8VKvj9PFiYpCBxPIzqaESKH2cwze7e8DwewNUE2
qK8o7qDICR5PtnJyDFiUjBaHsGh8kLY+/gAH4zraXZYawjG4skDyyu1imWT2atem
TF3s4eOlAoOjLCBrVKH0bDf/2N2V9IS/JnDL1vN5gfrB0F38mgUreWN6l/hdqXdM
qv0ATUKPI8MKzGmuUsJ6mybOzIqCG/fk4nw34aNWeaFKJsah1prmdEi3bNBuOh12
XUeD9MDBjLoOT8zMKDtePiCcFE6tHwhBo/SllhwlZmPycTxUvqQm0ubQCXO5KzM1
I3eol29UReMBM+9zlzGA4604JgtHwr6iqmPRgw362YZwcvVgXMfJUp22Lm6Otf6W
x8Gp9rCuOBcSi4mYGHP4jpdkUupNOiKn+tdOConhp0BzFepD4StAGDowNyCELa/l
1nWXFrqf0soaiwTXacHMi6it0/Bkij0fEngxdgVSlXzW2QGtCSR408PerSwEbO8q
1Mly4pyJtScjW6PoKrUBhCD1tjjgWsuaAwBy9H6rT3Kdc/ds/06g6wHOo2e8B+pK
9pPnuFN32rbuSpapjeFO+joO5JH9HX2Ea98XkPAsDZqJWzYY1xys3PzPS6/xzeZ7
1wrfSwmFBwb0DPpuN4pq6+LXptQNSu8kSj9L4ReXSqg5cawP3BOkpyum7GBDufDS
oi2T5xx1m08DEYdtSpy+/ILJdMgxhOWI6GuY7q0SqC7Vn2yNnFqzbSSXDSlL4cIo
KgNxg7m5DInhH7qeE6OP9psXquVDXY5wwWuKwQKZ8+YPEC1eCnTN7Cj/LddBTKhH
Gr6DrAywnxs/g/ov0LwJDICit8H+xWxndr2WSNCXcad3aoehHSf02x+n7PjPy5z2
t2x/3Lq8gofluSw38jkzPAlXn0/AtLJPPifZkwOQqKbysA9+/imscp74nIqxd05t
ee34ridVptAp3vo8ShdqOXLCKD8UlfUhMO61gyXGjimsx3CR/wpKU9qCbpFfiDuJ
n3BAry5nTHhvbwQQLYC9mZCfzuGkpYALykXqAcNx5zstPC5MLhk+HWDGqXCoII0E
ccY4d8dGMl0IY7oJ6tzVc8dcQJdargM0M0DYbJP0lF3KuNKOmVuIriMBgJNS+0/Z
qZeaYNlD4e0AvPktpEHTOQ12gaYxeMWaJtJSAE/UNXcv2zI+0HHv5R3A2koxgK+N
9f5Xrqs4dV66Rd0IlG1a1dob1bn9e1Af/2WONgWkn5QdgaK6DeNlRkNit3E/H9la
29eyDO68OpSen5sQb4Y1/AlwBcuYCOjnmqzX5OMah5bS6Q//F8RGEyxqaKqImJSP
O+ltId7DERasg8yHGH0k1RqLSKHKVF1XdISv/zXZgKZ2TVxi/aovpQuqT9v7RnH1
qa5r+BvdTIKB8FYPkH0HUymqpdC4PtBX8GYuDj0o3RBrmljAnln/V3U1C1mBJBPt
fEPp3lMjgl6FxMrAiCiQzaPr94thPNHAtMufDnMfYn6PhhdsTYDH9O2IyiFddRPz
MQYJxwo8YfIeFtTYOvWmzp2Ez4zqHHtDVgUSst+UVxXTYz+GiqS9Ar7QEfxTayfh
Yo41GEavORCq2pO8n8tfLjYu4rknp6n8Vc4tKMdjuY3Af69lKeE6MZ11ziP8N0aB
fZGCao0Irbj9LP7+oueoIGrGMLWCJs+OzCmF5LleC5i+/FmHTrtZPHCeUyTYnmBh
R2LUzs9x5ZRnPmRh0Krbp3O1nRCGNfAoyak6cDSBfYHaf6cD5xseaIBihI0Jiz5N
XgR9glYw9OhgUKfWdgbseg1FEOYrLt32/+7pNC2KRZWOO7pUIkTJGDIURBkl6WO0
5Q4w2/NKs2bAvV/Nd7wne8qAW5NEnwCevBAg/2/iWIhA1nHJI32tE9BjQoYqUpqS
tZxN11xrthv4mTSQ6tMpmc95J0/ClPaQ6E67mQ+lsiM8hZPWoCp97KH6BT/XMxBL
HCx0w8RIOViHSJRpRC4DbCKELKTdUlyH8YAzsXWQGBRvHruQvQWqS0ionpuD44TO
gV6/ciKy8v87eH9rfh1ASVoI01eMq1Apo6tJNtyk0uNrGLf6V/MGQvkY5tykB/+t
VP//jK5yaJ5qAAH970koJbRNFvt1OxMoaR+/Il1hf7L86GyDQ2yy32G6f2be/SQe
caXgFrqH+Ilh7lkI8rvzizQ/9fem0SUdicjW7hYetRpR15tgvRCd3WI4jr80csAi
9b2QM/wvrNoeWhTGt2AYgjKTSdODOYyhL5Mzc5XoXeoiA+cFZqweVpMNLW9iua+e
eLdxjTtx/reOQFgOMoEDQZrOCVM3kU/Q1RNWeQkl6p+PEacuXwPupm53yTir/L6l
0QCFajmz3WcHmjsF3tInowMHsub/bLCumqDtL7J1q9g1N39DYxPMZJFodYVjFKoL
6Npp0/p8DKNUeFbNjrjSZ4dc2qnwsrmsaqwJuMC0H9FC2rXS/D+vP5DRRmSak/yr
TIA82eAap1eCsBL9WQyWWfAfmJWJEAslVIWIy/vuz1hMQicV1vpEkUwmKMdQo2Rp
L0O0J5OEQRZCfK+cidDJ1gvuKzfeheUwSa6AfCot3jiZK0bTtXj3ihukUQGqKbMK
zGPnKXc4ijSPrbJF8EHC6oYYK7iXK8e4CsinJPXtkvAe2hqxkHcY+wD8pYhxxUNs
XejiZ9tk14fCoW3dLZY+z3J7vbq/fZPc2GljOHa4MvVZI4f+5rkXUVVhqDnIhYds
9+eiwDBqKMd3cMJsoWKXI0KmsPvb0hJE4OHDtlIUsmdV9AFZwTE/kQE6+G9u3dgw
VLgO3KSbNtKh7UynYZb0Hmknf/Y13BCUFiX8NQG4/gJCyFMhQX09peIE5ao4rJg7
HgPi+CB9MQExmhQe8Wn4Fs0CuBg2CxFunJuN8PdbvYuT6Q/OY5Z6U3CZJJwU9vn5
mNwL4Kwr1GmnrSP46iNKJveg+7oxhM6Kvg8Qd5N25f66ymHbPCriEN7c/kAs7L7G
CeYoOYSCXURpSDR9SgY0sCDNvNK3sPOCqnj1qmxiRWJzo5KgxYCplZyC3LLz+TkQ
AVU75VUpFSt7GONr1XixiD3xIfshSUs1Gfm961jjXakeCgv3nz8Xysc0JqM7i2Xu
I2mLCeKTWWHWKiWAuvd6ZURaKyUFULN/qJuP/hguNNSptonwg1jyKma756dq9N9t
GFIUSWJqyUnniX9TQqPOMHh3QzMMFuAtuvPdQOzoj/ek8NSCbgaLwuJOTgTMj06+
V7VIo+j6P9b2xd2CiMdcXSD4SRtIteo3AMOD8LQvaCdH6omr3dwP6VtbYHxo+8JU
QUOxNR5vdtuzq3VP7LYHQ0uGWagXrRcxGDYurpSwugEe/0+Dz1uUOhrKUZqDcBHm
SFP9T6OVr9MzisdvSgsqvoqP5E644vtPIt8IQ2kF7calLFoz5BKjXqEM5U0RNOc7
LzDylMXsQCD4xgieelXicijdVpcu9wYA8pW983ZotQCj16p2u3JlbU9Zs1ySW2uN
2/q1lU5EISvuFtFnx6PYnb+2kmM60mANYA7PDsj6AT+8ZgjNFwIJaTBxR7WhcLuv
zPXbW9k7UbEUszpwXv1v0ZAS+9x74pW3Rq0GcF56p3vIX3TLMU8jtUMMZZCha13G
GTMksVM95qq22gFd8MNCJmP3NSXs4je9zlpVvuyLOkeaTGY/21hw67DqCVzX33Je
HpAgwXnp6lCbG34VJvorpHazsOJzZWq8cN4vy/xt3jk29WQfn/3OeqaAVc4kEPuQ
re6UpI4tjqc49He0XteNUzLl6ZIeFNGLplioJkg3fES3+/GR9lV78OQVegMTJJxJ
GqfdLIc3Ma56PesYDQ0uzYDawbqIbHrhaWzs3evFfha6bBeYcKvX65N3INO0E8O7
6HDfp11mDj0x1/L+uVQrKWR4ckR1Ln0+mXoOxn/XixuxEkZA006/e0hh56ljidL5
Y3gTWatlheuL7RRKx9Yo0RW3s58OIqvPQXpIbj6caVanVkarWsQuqKT4TDwPs0qk
ia/mAwbePhMTgunXMX4Bb2lLUDArBgNPKpDE8l5SKw8MAaGruVisy0uvxORAGU0Z
+VovaqGAhSvVgSFqP/g67uJUatFII103mMpkNrbBvGpPFZSduKun3FGvw6hfiIKE
QEJoWn69qER3PBINaDwKPqXqU6Yf46+uE1s8xGNz9a44KMM9r+5nMry3aqvMQeZi
1AswOg3OWwFXgUwBIzWr54O0kcpJSBKEChYiYTwnBNaEvj0dlfm8Hy2o8Bu9QMvF
xviw/bIIVt1BQU07kocen0S10hJ56/TYWtDtZZ5Db7tIl+PgHsez8JbVVOCua3hK
sfihpHq6CIvE6pAg2mjVydef2g9/eP6/AJ6MAMVCk8X+a1JVioFXbc8hjMoOVNR1
2+TXrSoIG0goujr8wZiEnTaV7NPyKHeLpCK74pjasD3tuk9EVXxM5Xrt/J/NLnsc
k8y47HxA8gTKwR/8XOpJ4aNxMFL6mqCPDCcC2A4s+fsHN5057Z7KIN5oCKjNLnTB
GQnnoneXOvaE82OU5RATJ1sQgJD5xs9W4+MqB/4No0NnbBLGYLne9IdcVa0kmqKZ
ojNGSzrMJK1Fu3vn98rbAs4hy6T3+D7REEHcaCikFKqgRvoDJ187hm6X3AoHft/t
QccDWA02i1b75TzWErhL69XWGebUaawplPUAfmfAdJdZTCWuJ24XCoZkAKbzONsf
5psoebay/XJMFF33AOj6/bBk7HSFPmsGI7wvcNO+9ldQDFgUaCQPPdrxqllzN5qk
DUitYRXAXnludsgJkW1n5boomrDIM7Msr9lHvW7zu2xhbH2pOxJcJGws/v7EsrSo
Z3xv6oRCR9cHASPKovxohYHMWl1J+prrkoreW0VVFflrj7kVQkZgJ55QMM4VlA36
inko7vWrqBkiAlgbnD+DgjE6y/4SsEIJsWHd0XRUe917X8kFBnEpRL5WgYrVhzW2
piJyS4f1R15E+gVxhx5Sf3ROTkGtn5R3FbxB7cN5B+Kz2SoE7ikG3033LwVvSvji
Jh3sTRhNh+GUbeAkqsD8+TENJkaPcqqqmv4Do6UuKXchg3UPhK6baL1nbgfgDUxY
D0L+JFdt5X+OYHw57KF1dbWvfMmOdPr+GyRQJgthf307/tNv5NHPWhC3sCLYTK7r
msp8Oge/wW30oan9Je2SQUlrFx2UyvDiHB5IGrLUVueNw1c2z+9sDQnE7ShVmqpd
0ZOr2LRxkPfXa/mvxoFd9qgJRkjCF1LHjPdQN0QrT4oL7A3lSEEubo/zDWYCEFF9
1XwmrlFg946cOp1XNJE8Lgv+3/8gMn+Z4poDYu3i4MTuz1bFh3OBmFODvjbrgVwO
okeIx50XMJss7HJQlim6RVf1+kWrLVEuwojTfQRovztLZHfNtYk1pmKDC2da9mYk
9EgglHjqr1E/4iM0+EzWmlI4dcWYLHh4dg9gArRlsdcs5/HgbuRRmom7PAz33076
9VquPmrFtA2t80kMAoaghn0bNquYh7UIwFAbZguHQ+L/p3XrOHn8m3ynw56AELYe
pSUvBDBk7zUa/2FySfWTYaxrCpPOTPOOwmQ3pB410g4NMShb7lPUw06Bw8sw/q6g
k2xe2uR3vVopxP4EJMu9Pzd8ukSYOQCgKNkCuVZSyq7WWGzNQwbA+InxAzDDDeTm
SOVYjPfd1ONxByPxrqxbGYSxO19EgmTYYWH3w9Tpst2HdLUxoCswlYtKhKswr0P+
EFytbqmm1PzQP6eOhxIMiZ0SOctAEjbqe9JxU2CsNu/ZsQRvgR3ZfvZU4z0m5Yk6
xYJz5e67u1cHnq/tZVsFrVbmC54uEXxZ5ItfuHGANjSBxvyds4fD233kIcwmXijQ
kT4xQgWkegJqx6RHz1cGolz+M2O9Z2arF4DBbZ78UOI2aN9vKz/+xWQlnpL0phm4
zkE/882f0MNo83GYotQDHCHTO94TfB9lcxgG4pbraFgceHGAMyHzD+3F3CsltTje
V/DSQBrbNasl835PtpLMVYkWaQbqBfrna3+t6zj7lSfOjS8I2PYJPVBShvD5o1Mb
XT6RxLTozKFN6HBcImNzQH22eFP5UNt1nnLhm9yYfqSH65naLmBnYTMRBL0/UNJI
E6gsnAy+4PrOHwHGuhhcjl0xMYhNrxCqhl/3uicoezO5ceVt6uIQCRBLNX5DO0kp
n/sk6NKUz0tyhqCvxeGkjvDhgmuYbL8KCyAoxd7OQQ2yrEwVlaoN5eC2vRmxOHKt
ebrqK2ugqCXA2BCYrfYT3765z2TkwtTTzlw+RNZ9OpdhKNTfYkmNS1eC6TMmg9Kd
oslZd60YQ/9SrpBV0ez9Z/HiV+SyMYKx8LPJdKOV5GI1pj+mLsW1sHy7EAnYKpS7
ke36dmaOa8vHGPw22aq1xOInm2Dm5ZoAr1avA6N+H3tzIcrScswiKeSskd+0CugK
Nfhc4Du8tU119bvA1dAJeg6Na7bhNNfcEL9xzmOsdksciOb0vmidqXrBHzvwiY26
dPBma//93NF6K5PtPdNv2r+deO0V9vrgqWMVU4hLHGDlPHTADy6+TJdDADF26eiY
ANmtc4d+Sv8HkCT6CcO3sGLi6FneHP0rPOcgjKlarxSn2v+yHDysv7xZK6LT/OY+
P4ar00wbpIBHQ39X1dwM2EEkzMmvm5vjDfMEMNJg2FpXxloc/rCm5KLYNomT+BsG
sa5Dn5eO+DOy+QCIEkOP4KRPDySWIJUcXPWUrjyMHdpT5NHGjrSk37dkamDXKwGa
c2XwCJEdbhM9chE5DXb/1DrDcCbAUihLClk2rlgwOuWyOoiCO34ipXrTuVONbwGc
XOwH+QxRr/fNmlyNQuVm7V3i11N0d/bfpA1b3nbMYvjJvrAbbrctcGMNu6DXgliO
hwZXK/yrgNG0OZPJozcGsHjYno2K/4VOI6Xbnz3knaRnzt+Rr/ROrG3wTv+jkxb3
x/19Nhd6MiQ9cZTHaxHuDn/dIHbOkHafnLGMjWvSmBUD4lIMqglNm07N6IPPizt5
BQQmfrlGWF+YyBfEovWZt28OVjvEzwZNKbx4XUkao7F0LqVg8TPhsY66goyuhG6z
A0Hsy90tonjt6d16fwc+8qooEsTrN1jxqcwXF3RbxwqiumnX9I8zj43a5LAcqQPT
qqOENawEP2CLZKGozIpnNzc/xon+OgDWFx6sCcNSgepCvt/Ut5BJn92rVt7Sr7HM
qb+v2MIsX1BzgGG75XJdQBX1MmRl7lNSAUjkCoWoF9gjxKoKLeN+pCB7kd57/Vsu
BBiCzuWJAW7jGtJmt03+mfXx7CCVZXf9GZ8Q1obYCFJYka37DXbshwW77oUun7xi
qGo2myaQzhARNPggnOEnmvRflrBz7ay5+qKZD2aj0mU48SIaYjF3NnhybK1GfQhO
aNvzazpebq3JPLXVb54UMDUV2aQYXRf8mh+6yRAniK9/ujKXYAE3FbJl0IOxM2nk
3e/ijIlwxNJvvEPQY9pvPMIhCP4jag62KUcuz2qCFjsxsfVmU0yJUQxV3nyBb+G9
B61BfxYzBa1bOwM4iNHOc1nHolaVazYShV1ApggYHpNNJJgreJDbXU5zxNPmNhh1
A8FJHVGjO9Py8SlCL3D6Zu1tUmfcP2xcwdKNdFaYMHsK6zP1F3rxRh/iEWKzWTY5
hAzgiAw3FIN30iodQK+lUdnaCtpiatYW+m5fwFaePBOL0LPaycSuA+wnSAKMXYWo
yO42e/XP91BpI7GOwIdM+Tm5CyfWVDSZsDcqjhvtrKIA4/YWaqyzMNPuW0uXRFMf
Ek2z4v0tipDVrgaa/bZY8MMkkbDqKEvmIqT9dVQA0HKXEg7L+ch0rlvLk7Z0ASzu
OZBe+h759JNAoqkXe3ldSMuzkd+o9DX0BVXZz24KuquM8fqOdPuySzP3i2Ft9sKK
HNjJtqEiwWWktBAWancRJ8e4KpZtPk3Hjitk9imdCslwZhUx4i6Krdk80JMmSI4o
eUAuCFQrKr7wPhJQ+zfxKVcZX0cnI/31BEiSz9EIXDYt843eApoRzpQxJ5NAWJFp
5C+/jV9MmAx6Rl1ZNUa3QI8U8VgH1kPfBfBuZ/ytGSsKxsz4v4LbalDUhaet4OIM
Qi/5UQwxIq79uQ54v433NDD77Uzb+FHqxTPfcRUX4HNxzS5J2AahsJmxEld9OSMY
Fh//scOdrhm7j94c7jm9MeXtToZbwHy+aZhi38tDa0ogyOz20hI6xiW1p5kKpwIY
NEuAWtaBi2OLFkZDEJPNew6JlwsERr52aJanCVselCJqgMPcDwmBQ1h/1DB5wBQQ
WJQEB9C1efy9zs57P7a1TEt2O76i1luuYEVKy3k+bDmc4jQmo4D199ufRbae2XL2
uVQxInVawxpihpsQNTpONU9NqaO4b0HQAfzvVufhjDxoVkoylD40EGfgIivqCZ6Z
RclTIsD1mlG3IPef0Q+Pi02kYRBXtxLidIW3/AjzlUQKzh3iF3b+maOUAM20I/TI
Ls4ZupjATUrd7GAc+vKIlmOU1/U2DH2JDRia3srVg1uUsrcvjcOkgzLG7RPNIcvc
j9F2XO1NZ/NSH83d4kwJq64YMcY9+D3h3GfGDfluiIrNtbdA4Il+vuG1f9QVjr5e
b1i8cD/9y9+rbosc1H3uiGniLvSHr6kRWfAUTGt5at+T5qx2Ea/PA+VTSfDY2TS+
Lt5tBfx7bmw7Wa8AZAR8WCBwkcf4NC6anHTcedUgkxLfpg1Q2vBvdsU+8Dp63GNA
tKPNQKtTmqK/wRJY2tbCAaOP8lFg1gaTd+T9NoddC2pIKXwD5cJuZ9lmjdojmz95
KXuKR1hIyzd6czyN3DFaY7ledHz3uBJcMstWL3W0/AoO+d02f2d/ooqf4cKiYjLf
XqFhHJAyq7hvU3u/kXM3g5eHwuV8EBfup1lQrw4RVOKr65q1BSxYNRBn6u3q3OsB
zxflhIseJNOXuRF9ahc5nssMXKIX83Xkzjkn57+OgAvc/K3jaz2kZCjf5knOmEde
ojrgZKXreVSDSYrdaNfzxzVxwaroHXPQWrEyMQb2Aym1mJLaBMfNKfQHie0IFXA6
EmKHA77xizuHe+ZNOu9JrLJBKPG8OKbqqfOTZmO47OOIr2YTQvH+zXeWJxxG9/6B
t3k+HSKlRepilIaXQNKIHktCexE6mKfoXYTngbo0zZ1a3T87adt3J43CZnqctArr
rWzbQLCZ0cvddz6edfO5vQbR3BGsGIf6gERx/4jG2L8dlBaV17exwyNjMS24sB+W
x9UJfKj5tYDoUiFS//UX+icbbde48kZ1WA8+2PzpwBtwD5mAylXl1q64hdVdKU67
IApPQQPGaqmzBe7OKH4u7C9gXRCR9dijmKPdGKiLZB3rXbV191KXMIZLPOZE+OEY
uTIQX5JHn4lZ0Td8/rZW3c3kYCEFUInBa0H/NHvkoAkptExOgVNDIESOsdmYnlR0
Z31Nf0K/ETOccqfsRUP0+ybQMBjPi23DFcUOpwKd8zFR5Nj0eAwNIAzI0o8chXeD
wH9dzSLxftBtgzswDsqm6Z9M+fx5JFWVVTj/mLcy+K5D/1B5JXpCyyZg/WQosQy6
CIUEpN9nN1CidAz1Zgi4SHRgXmMBJEveUBTtJuXB7ENVMEe7KsHGB2xUWjLjn0y/
ZKPQCDX9nawtQ8yXSacyJB+HQn2pZ0xD1x4iKUaG1tbdr6DU5eGhSO2almRX2w7F
zaHfXKq7fhnHthvdqo51slkJJxhZNaxLax0Cre7kIQ9o/g7M4qwjqNBCr5SpTdhM
hRJzzldGy11GLPo+RWfotFUkW+7+Y8NSaank6L9hhdTq1GgZB4cz9GKZTFunVsSc
+xzOC5dzU2MG0f3cmzWzaEmk315ZGhUMhz8FK24Zww7r6EfTQlL7HJwnyEApI1En
tz9wdoTdOr8MxwkqmHUHhVSQOqsyl7KgW/WP6uSryizZqOFhsUxgnjbOcqDlUpiQ
F7cx3xpCZBb8nVbYlCuhxXcOEDUk81oQCPThN4Wi7d/OZvfGlY883fubaRvdmA9s
4AogDfs/HJzLbL2MgOXTIHi9soTYcWBc5WyqD2UiAZNl6MUQRZDDThcoEV/v3xX2
GrGmlg1YXmrmCCl5nRfVJa4kABJg3Uoy+WjmeKz4C1WCWXrCMfcZItAICsbeKZYH
CeCdghHPmIvU1Ue6UrTh0a6cFAeAThDZyXCWHiCrCvoVip6PVIHdxS+8n9zxUGdY
UgphRRvIoWBjtlv79vh8qHPs2eBb4McG24BCm0qlJLWGPdbplm1M9ZMaDuSpZz+3
EEglojc2L80ZunYBhD/2NA72ArOAoKc/KseP1CBiRWKEtIXtxfxLF+VsBdbgOE9u
ZbEkYKoRsrECSgGcDFEKy+0OKxlF8zBgM+F2EGUJqEd/lmc5KPJrpEH+lEYkzgZA
QsLijTTlBf2XCI+ZFIkT/HB1I9TZsmShxqjN+8K7Ti/tfYOnw+Y5h/heR93EcWoE
KQPRJ/UuiV1NZEh97YcLj2D9F0eoUIcf15HXNxSI189xqKidx5UFU3EKBN1Qmuu6
LO4rQOLwUzVWZENBhkhTmU7/95yjfwUl1aJZUe0gZ1ZWSHGBZGH7Da1JNBvCfRGy
B+PievnDywPrASn+G5VWCTSbwQRML9TyNvBpZcieOshAbB5XeVqOLY49g1Kred3l
je+DscYOoM+wGis7rYX8pGLUMdLOkaQWD5pAhvQDRycBJx0Q5TrO3QEt4ZjM6i3a
kiSH3+O6lwMQU/gtb6l/yFqKDOemoOTFujTcKET8AwoCSyjl/pRYyCujxGdta+Oc
ecACogoAn5kntPMhftDtOUrwP87Uz2ygE9/Ax9s6LGl56TE+NFHvA7NMpLsi1RxU
zh2imLWcZSvfPJiLRq3R4/G7QLU2D7/hx9nnWb/zza+eHnp2HQH6JhEylSKozu/e
xyrlFqCVNN1796cN/WvdxcemdbNS0tCzFvRnYdtfPubebzoqml/TrYQ97oxgFgDS
hSMsyFb5mTG2EppS9fPy1S7J7KSn4F3nrTqqfc70ckdMYQ1n60M6vEWCPbhaTYqC
2wbafOIDPjuL/bzuguDRF3bCGN3mySaI3RPxbVeYsj36DBTVGsXMAfiaLG03g8MU
7uKSH2WaX2eKPaCCzIDleyekHZk0v6mKAY7IGa/UT5UfyWJGeCIv1r3s0vnnxUub
fgm4/Z4atY+tU2et1yeACyfh0ZiFejbRWhpxWqj0lZH941iNEbU7lfYbk0H13uzE
MKfyUM3ONJTDKOWDoJH/3zUODYNtwJg4KR1oDki53RpzO7rUYtuJLASOTJ+Q7HGw
9VAHSfRbt6Y8Gw4moG/MI2c2CoLIbG49z2XiQOEbI0wc5E96/T8XBFc2oHDwrVo+
uKC68NEoiAd2SsB3VD2Zv36WC0MyCUDCs8IY39Bg+VbVaWx0673mHlD6UGa/v3dk
Zq4p+YFaWC/Ysa7DXE89mu+2Dn1tNBLhqHvSpj3WCnu06MF/0/TtIPyTLXcIilPx
RyXRUhhjbk/Eo/dKduPWCDZdQSkzGoMWi477INp5om0COF1+9VJE6DHEEJ94b7CL
/fSjpVkRBVaAmEfLUDQKrVGZR/K3Wophw6nnmWi8iRp71p+Cj87g0qmdwsqjYbCj
ytUlyXPHyYbor6eVvATN729knydN3aov3zSQLBGsmMn9UhZlYt6Y7ION/D4DiRnB
3K0oEMfErKVzrHJUp9tD9DOha9fl5VeTg1P6Y/N2pIS7Kema0FrRsYCpzNYl3Yrx
iO8OOO4ocDnnWcLJi7Y7Gl6T7F/KtltdOQDhnq6AbD76/uXOSmgKWIKLxwXPZBKM
rEOhl5zchQanqKlCuVAxJvJ1AxvMml2WUUyGDk0f+kjUDtzSPjxwv7AEpNixva/V
xqn8u1Km99nG3ZYi45zCZIrYLkSRXKwHPE2xZz7rZX/N90UN3JPpOUGTg7eLWNYH
l4KagdvVDBUStO4Jg9mj2cgWej6KhQcfiDtJ8ywFNUJG7Hf3yQ5BOT+RgiDArd6z
/owIy4tj6g/nDUaFD4PjMHI9pMdNEOKuRWOxd1/QfkehkPdqyMnPxEprJqefX9A3
4pVuVs/ycsSoAFxo4h8Mq1Yhr9o04Ll66MHLqbvEQqF6vWYrbw0DN2qReFcr2aDF
yuX7u/xp2+p/SAR4MpVmQnl0dqMw5gTG2p+bnthNQ7fXCLLzNoYg0o5iFbL/F3GN
/HdhqnrDs+oNQCpZnjNyZd2/t9MOTJF3+OoG9ohrFSIRaaslyrvwhue0d1wCxi4W
Ea+tfmmy35KFvnCHMOfvbFPmmfVZFpTde/3NPI1SUSft1g1nHqb2TNe3y+KdD2mm
9/c9r+i2EZRxsX5089CpB2jZLPPUFW3D2njlXnX+KEiy1B67hYLlqeDnX4hx8+4Z
5Bi+tstqxD3VowpJ6PZCBCWD9V4NmoiWsGqiepEbBC/6jyQvl9SoHfQEn4nR1A6D
q6+0+IDNrVkRB/aS+zWb1ccUekzPeIvAb4JqgqcKSJrOq0v306JhpHCb5hkNdXOx
N8qkm4M273jiNIraSlb2LPRwM5CjfBxlnxSWt8TbfTp7zTp5Caz3IIu4jA0iYfp4
T3DaOOYwMVgJ+vxB35c4PyyxO1j0bYc8DwgqDzkXHOw0jIJ9zg/9KBif4M50evHw
sg6hLO3LPf25qQiL7ohEvY60m2B2gutbgPibE2bunl1cU1FNG/nRzE060pGQ8ejL
nA4cytcaAw+DuhRrZy0Yx0SKyK3f9shmZAwt3j1D9BbwiJEfJWbGdvP9cCPzIvkd
8MeH6WAjSpq9/BhOK5qNhfwqUApG6s8t7UNrLBJYo8jx+FdBOSiHC80nXBo50C5t
1SFE61/TJerjpvtxl5bZoWz+cL9JvHWQS8NTHnJ89HAdMIq/wvhI0+IWdJoCO4IK
qnTsUSb4hEFCZug2+F/8HRTHlVn05a82bGjJF7llIbXky2nkyE/lj7333u7PiEua
5sd5TuoBmwTA5OzRZbo5YVnhK/Lu+YnbQebg2WJmIfCLYJOmZOmW/8nehGJtq8Eq
+7Fo2Vl4b6vbHniYa6PJJLTELyBgxlRVWb4nT0Bxbra7fd4N+dUs+qBbCey6v5g3
OYHziTWU1IxqeQEB+8E02Ys4BGbMB0GeR6ccKtV6tHpuQMNI/OPHSjnNDFIw26Nt
82NAfTNhCaWtBu48Ip/M4+OTqYanQZV9TVAtG4xFQ5TgUsTc5V9azSwhxkF40LwH
xWkP+23yZ+og63Jh47LhUKy/HYFnfuFigtxfRJxgANl4aDxni4/K6gaUpHD+1kVV
3qKuq/zSp4OQSidl76oUVHEho4hihou0wsho1DYPcWDhbbz/DIKF75+Xp8xpDePU
on863ZdCxK4clkUkdIfjwyEHRytQ8L9k9fHOx046emyUINQYSXzTPlP2u1GMB/S3
iObJoridXqROhOueFCgPGfP8EnpTSRHHcYJzkXxrPC4ozH/k8GlGQzO57aXrSGHW
7thC5SY5tUuqkzuBeFT3mxFSQs6rswoWRB0QI1EtFqcZ/GsQcFIUOLVc2gpvlYRZ
VMgZsVjzNkmNQD69ZL+Ho5Q7Q79ynpXP30O3MlBK0XEQClJO2vf/mjIpAcwnE9dw
QTuYTpym3Nc7tvWv3z8p5AsI+dZkUPbT3PaDDo81U0ftiPwt3MQUabruY3A7cMvv
miYeJFm3b+NW6EryTO+77j7UsqzL3d1rOPXjwOz9zfhqUvo40YO5PEcHJcWouTlR
/sk++HyZy7cSbfvlBhECPCYSfpYYYAqu1gAEYMHgDkURyWS/G4tN1DKU63TlEBA2
ArUbssf+JLJ6N56Jt7H7YvdPioMpZ1yREhi3dcQ91TP8tYWotr9VmeS6TU019TqL
o2WgbHkcfOii9jRW+H59zVwORGdl+P+2Qzk7sFfa3TvTGGf6T9WlilOGcqkYhKbX
C/sDanFsYwp6rN4815jtr+eOKxpg/xduqW2OCfOdJ2/EEQgq1KdNU9sZ+ngYdSl9
JJeOCBwg4DJ/u+iNQ+4bnxavrJmv7b5fdQj57E9JwNnO8aQE53VeFZ/zKQCb2dcA
KGyhqBLlbXKqz5iIl9MxYJ/y6N5PxSsszNTZfAiacMJ+kudbNEHGSHrIBmWhgkez
JFGHxQAOu8Qjputh/ymA+5dSv2Kn3LTW1VCuTUnsTBWOUqZ0ezBZiFkS/FoECOpz
ostG1K6L6h7ysGbMtMLRM14lSDBRL6/Ori/Vnoi50sftCK0e71p7GLKzJyqlRWaV
fhj77mJtrCzfSwu1ZSQD5ZADXuz5yo7JC42JVfElwcp/IPRT+4tkh2HmzFll3YIU
DBYL300q/I91tqCIpiFaPvwBu4jwkOV/Ci63C0tgSRwzkLGh1u8ib5KXOv2nQh+h
k4ttwu07qTMGJDnbCcd8WodqG7B4fdlSSfQPE5YCkX6U2OwnCJOTmrrTR5YRuXZ4
+a4P9H6YlvEc8O58cUiMp3TcPkX27zOJg0pa4t2qGJX8XQOksVsCBAgcFjx0geQd
9M03G6MjcJrqZKiYlcmaEUA+0iFkc5dkHVhRLvEzQ2iiUWw7S8kxD/BgYPbbFcLR
+19vBjQpQeQkGFaKC4vjHeFB3z7bfLNqaFHjxitsappTgPRAO0fjXvz2o5v0K5q8
icss2NnXIp/dfBwiwOHktb9f5ksmynKjTusbKmxrHoyEcRfvC7sPQLKDaVapH19/
hb7WgH9YMtK0k+ER5y0NZfcDLkDp96lHZ6dNewOp45m3kMPGAPynzhwiSmNB5/6i
10IRFcl6a2vkB/+c77YSDqBfSLOi2zzHNEtxLhrtsg1RcDb/txctUjVs8C8p1wVn
N5AS7WAvz4MqR3Di3tCpnOI1eXz2I/HvxBQ/mYFd955311VQPG9t2ECgHqhH4wl7
INb+NJQQOkuxMTlaLmcjgSR8ah0AGGVS6iBtlkW8VpHX27Ft6K4yvJq/fQwCt15H
BSORfbWLgKyUn/1KP3vh/5nQlux6sWXXsrzpvW7oldXR3HUi7CW3tzHg1nQ8Uysa
po1eclhnjnvUN4flgaWHmNIuFVsihW5KQvS/OxIudoJR1g9TAvrVFPb/SpnMJRPW
7D0+Y60p4ro+NuGxOeFxVh6lDN1Infkxx8r5aUCvS0fdLH6ALBQJZCgATyNz65Eq
vXsamgWKyonFJq78JIGueBMwtbB6gPEhOfE1erjszQhtb2nwy08Ah8WG2FWkwvKg
fQd910l9Sl8rEeNqIvTZNBRw8iuQJP1QDB5K0XffH0/bZlKyW6SrkltCLwxfjfax
MX7xMRKJ+HBaA2SGz70EhIN/uLcv6jzPidwyjgVcZDR0m2EHGwxS5iTqtyiPxWJI
alBE8nsQtyLqtsu+rjDPSpitRk0HbfL7uYsJGnslfwI0Uxn0EouBVcYpV/iubuX1
I7pb2AeFVk2BqCHIubYppnfaWy9ngUtZnQLnah8OvUuFOyfVDPEdbv726Hq3Brme
D5/qrTEDct2a3JMcl0FEaUdIP3s9TmgGuL3ahJxdB6GLFSqemCHpLKJkI7OluP9y
xL2oCfHTZKu62G3mizW6MojG7rIkXuZpX953RSrsrMyeX5OAaxi/cP7nOM80U7Mw
wA0ZYjHv8SP4wgHg644JODQhHTjS4nuurSnL1vqYN6qtY3iH46t1agfhilDzMPnJ
Bb3y1HANm6yV9rWQMTQlA0WY6HFnHyT3kWggQNWFiobtA8oWKZkfXtufvXrkQHeN
yfFbwWkkcyDaOdgSMJeoQ74DrffMWiDWCiODM4dFxJL3bns1ZwPZfK2ts/Pp0B7G
NCQXkSFBBhNNFC8BRS5yYLRW83JmwXLa7562rzMYMLS0F4V44ph1m9Xh+SPxi2RK
fCLvrUalZrwK766OCH8vCJoSPAw0OA3M69nzmwnBeTbGRe9QtMQY5ozDuQygcwSC
2Um3ilP3YmiW0l5unPAzoR/40Xddx2VOIKwQDoRarhwVIoLQ5jAOYFd9/KqayRoI
ehZ9teP7GudhMpvAy2XIjN0NLTm0N1o2mMtDlp3Rd8hybxyxdqFUDTxX7QXiO7Bq
Qnn1FCa3DnIHkUIUVCTMbXXLWK9xqi+EkThIuKXI/7zGr8KbRJ1hfVDjsChkgQDu
lUiyT2Px8aOs9bBY5zvJJquD5G8gqAslZDAoQid5FkpM7rnagEJU+X18CWa5wD1E
stiAyZ6C9yuLIxuA5gyZ4lSZNe6HIKtDYoHJkpm4qJ07GJIKpMmeDMZ7l6Pl8MPS
D5rz/YHVMrQ88ik+3kXcJm+5v6snTXjzPnRuIypjIua/xGXqT894DoAxbmauQRQ+
DMWNkaQXTxgGq3qbMr4XgnOZBDT4hf0ryYsW0fUY8uliriI0/7vJqJPBQCLcVHYa
ELLxy/O4ESVtxviIKmQIxDszAIKm6B46dssEAdYYukMbbEVaAxOlaKn177GDCIgX
fnLynes/NY8ZzgBwRb7kGhfJ4c04WO4J1YA35qH6ZcKCLL7rfm/PYEe2+XyKVgaX
lCDcRhMKRCr6TKjSRGviZtaFy6BrB5dykFrTDbOyCWTx1lJU3y83y8dnOM3Aoql8
Ztmbq3vIi0KKWh2WXpcie24S9t93HWeipxfCT/4xah5kDSTvOoCFtHRfOuZxFhxY
XImj31ezvpk+wNXRp+Y7M1jgEdFlrBPt755G54TNYGj//TSqN+apqJhCXxO4eHG0
9bCkEwzlBa4dmQI+6P5zThzU5SrzIlBcpY33Nk461jMe3OwmXDYWVNZexmlFGZHs
FIHWwAZ31knZFtI8DC8dTxL7X/9YY8jr4Flk1jGuTZ565FUjqX2uf9EkIuQRxQ4O
bn5E1CGhTTgIZeZkM79qxaaK+L4AEHHz/gGzeA9qnnOM8Z+v4j9o3M1FXBhcTEoP
rgH8Cmu2ivt1Y+qylPre8bkZA2E7eFpRCACC3b/TI5aJItareJWBagWY34RVueI5
ci4eL709g1qiz2oqZQjJm83llWue7Ay9LpvziFEdtJWyVJ4Ij3uNJQf4jRaF4Emx
cIih8VEArD8yd0GoK0hG7Z7jUQKczXJipqOhjGZ0yDzE71hWi7ZomGEjDvY1AFsO
FCunGRC5x+FIaPuBEk6Q7hWbB08xKH1lTP3QplrSl5obHRIxm/+qxFrvd+hIQWCV
3O9ZZPsDYlGVZ2l4E+aTHZXl/1/A5NAoFqwRoa2ZGbioxKzBSble7iYGYrFDicb1
W25D7+/9JQbwAbv/YYq/pXKRtW4YixXgsQ8scVpcpr1pZcVFeyoUHGbilZ6jTsTR
euZ6d1fCy1V76MeBshEa6mYQ3bLTS8szHJwnT1dcWjOF2k9YcN2WIGjobJb/ZutL
5ObnWJuGi6nBrp811cO6pcod5xw+1Io9NtIbH5hlf+SgfOLrRZbIcRRMidNC0uAj
SqbTLFKL2NmNIEr/xoCsS/bs7dRsC5K2DDXcmBBbzZVd6tF09xZ9aTTcOWwm9ESK
HAUaWOty42a0O5eRsNCbdWPtoSREao4vTORGitbI/veA//75KHgEnKdUaenJD6nG
XRiVF4kVLrsEu8jfbGx9dK6bwuz4xi2l+JPiIzSgRYyGzRZ0XhCv8EU8tvOFk9La
F6fsnH8l/AK8jz6idippv+SnU1Aj0EqQwAVs3uoWTX7+1lV2JgdZT4+7k4pAe1cF
5C4gTYQAz0wjH9T13tpkey2tklMIcTBXNr5n5WVG7ToJKs3Zw23N/hBsShilLA40
guw+nUnstiz9F32C+d5daofKzgmXZYPN4q3yVIMM5NECtGEYO3vvg/QMkN2l1DEQ
Egn30rL+ItqXgTl+LUFqwBlfo0MyYvoV1vbUZeF6yTz+T96jGyMnpFAMkk+0Gni2
0j1hzIgy+t9mNZKtkzs/9ONWAEgbzwl1knujq880K0friaDDrdXGqPoiEHVqUPBS
gf/wtzXsQj9WXpCyNPzbDNTeJSQD4+pRQsQrxV+mGNY0WuO6sq1r3vXZSkoYByY9
eDAxhaUuDNxhLZweqqwcFC8bAOsp7faGi7NNO2cffqdDJ+PcWDKQcVa7kJ623xSR
Zd1clU2vaj37Lz3X2jKwlKY75RU5w4dKZrv09HhzvAuctPtqGldN+FgQYhwr0sxx
6qwgN2jxN9Sip+CELzltuBUiAm6GfrruIuWpL1lKuRoMN03HUPlXmiFoeauNHjOH
Q3IbIsq3XSQL3glSjLyrFRv+K/5mR2l4tMdPLWakRPCKJXFoLKNvGHSX8Kg7oIgo
D+FkYMYFoeLuEarTP21owxwHLKTjOmBWW+AezvyJpYZSaleA2B8fVpyROlQ3YgGU
JfcnJx0zAalyAEucWLTqChDef5dYAQ672uIVl6rOg07OhNPEZykBYv47Pytg5xMA
61VeCKEPfFhm6n+axVMfWoHc9NOXFh7FDJsajI2+Yk+CJGaDZLPnPfXgl1RfrQJH
Svd85yps2Swg0T6zjkGQBsU/67U5moxYWFGmbkA7h8fyuPTNySBevmiTST1ABHVg
fQSHMC0uwoaJ6cMwdzvFTbKlqUGbDYwMABfWQqQrG5pmiZfJNCYbTTrzZZT3NCjn
+GMq0jwrTAcAllNhektbefd3xep8qrSjvv6xORVbW7xmC50jTEAxgXIGZleZDuZk
MiFrX46gw7gjk8l+sXyWQY38ZzrE7Y6pF4+pAOlrJu4+aCYHPu2WuhPck2Tiz+F/
AXFTwD2yfOz+dv1I6harYEHvl9bYUvYWUAQq00QFkwgg03kagiFaKwwAdFm0oZKn
TtR8rlpI4noRF43dytWNaWFVWHVCj0tnd9rz1QZV0M+kwVxwWxHltb55qo1rcGgC
lAEPUK4dGNPOUURfyh0K2BPYlsTmiWgtiwk65f5Eju1/H/an57RHt2mVxDITHOkk
yBo4OPLTaOhe79D8Oyh4N9d19S0yrTdiN7VjBosNZ1oVG4m87x60qJ9DSL+ttN9t
P0Hh1hXczeOG4KOMGR+YaA948JTnK+TeJ+K+adRkerWHDggc6GZbUTsefkeGqaCI
cptNIlde6DWqZaGP+BRZnCQcekKM4vJuJYxhZGdcF3OEtz8t5GHIah0dFAuNkY5h
8cBZ/kxxMkddOvDhOwv5WsR07OAS0QFlWEuJKwWcGOZpEmObZjqfqaAaW/qq17SX
suJuPWiJ/Ml6LK8RM4HevP8MtnMbXa1gkyJlINj2+p0Rq9Q/KuyP8iuC2vu69PmV
rkYGQLMHf+bKkVWj+tw/DPmV9W/YmjVdRA+UjcxMwgRRRDNaT2cHU2FiwpOYr92R
p92N7dBfXYOTcRebDCPj4Y1j2/O//w7trZ/w+Se40lOXatU794lMBmYlU2VZ7vzo
rHZWc6kts89K6R5fxB9vExBwWpI/C0RMvn8eh5xQwjuYyeC1Vz+GSSiIk0P/klsd
EiZZFTo2i4+j4zoZTMgxQygykwKG0ahndq8+TNWEek6YrgBL4rrqnj72npnRkXRn
Pr91aapbSGcYPAnSoygI5klZ/6EOdZSj7mewxKI+cuTaFoXhAhEEunQdJu+hYOPn
bBRfIkDde0ASTOrZe5l/FbOQFAyZ32oKG+A0M4cDrihiB6ulymnydWzhNTL8bwfa
kASOo/QZLkpnmqlBGsdQ2u8oITLdrxIpeICjdPWLu5zLhvf/f5RGqEcSc3ndlT1z
DgWbXwpHq6rYHd6BGssvJHpWNZ6ekthg+kPg+Bb8OZEBYqv+5FViLr0RNpvifU+a
LHChA/xZajQjLu0oSSAtsF91Li5yDvubHExhRiLxXuKIyhgv3Ts7VxnX0zd5CdGf
LxxkQWtTtvmBQ0T5TRXutAYxRoVpeJf50K7LtmueriagRu48zrFVRkPJ/Wf83GXT
0QVFCS/iWRN7C9WIJjlmbp9sAdIRCLRv5STsMpFJSciybVus+PGn2xNklQpIV6XD
2fDq/MgjnVbDlZeCA3ZmNHn6TqPsTIxOk5sBKPrimq9wZjcatlOshan13etKjAD0
HOS093qgynF9nGmWZflNeB0tK+2r/AegGclkzjCa6UPXqTmbNOxQQY8QT3ook6tY
q9HWBU9lNRzZcdKrKHtBB6zmJlfrRNWJF2vcvwlG5sDhaoG5+wWNEfi5haRk/tWs
9UZG2rCtoWKKx6c5Uj2B7RV5JbP5jmUNWWSUAe2gSNOv3U/VzYLOfQ4rq0XRQT0s
yQsRVZwmbHaiCxsTLRBEnZoeCzr+nz68vUNWVjVyFXsEpvG/ZhlupLV/VYVBebWP
fECfSDxMvQ0nm5QDCZ/T0QUQB4Niv3hZWJi8TprflTUGg9h7KQtL/fTLuorg9c/4
7FMuxdpWyk2e7nFIeMHmCbEGt08QZ5gQA7wba7DroahrO0eYmnYOWeYl5a40nrB4
r6kI9f2SGlQz3Odo+6C0/wauJDXa0bp8ik+wD5JPbd3syr+MM2FUmwPzmyENAf/e
qlEib1ygui812tglYJjTfT4Ko+RYs9y8uGOziqKqhoEhpJjrZw0i5DLddJRTuoUm
yNwwXux0SWwfh6ldrwkfnSOkukyR98M/nxZZl5qZeJifIe4apqQwOsuxVB5wShE4
x4R2rjZ9ipG6zGll+/aonLXfLP/7Qfyad/oI7Br4BIITSliD0uu+atdNa43k8y+2
C7cXD2Zq76gIlr2TqyhqGOpiS3AZRSrBlrvUPYea6UFl4/OPtQGtde038VZJgpEX
M5nu1D6jn3IBwtjNp8KAgauVzDApgZdv9tX1ZM+AoYCdJOBdS2od9RV0RYsrX6jW
WYn7ldYgo1r6mHB0yVEtmGaX7b7VU+mfpuj0OsvaUd/H9Knj1qGJY/hh6VflndVH
skOQg0dy9NdjirdZtNsqwZn7jvO/J1B6pWM4+CK5oY4LZzZmPhMEOu4T3twDXf5L
48sLYD0PYJeaBu5HEVIY8OeeaARBrhd6SY8hM+0xQBs9E1tmZ2XnyN2icDogORr3
JV7dtJCmhL88iX0d+O7ezQ1bU+PI5VZ7voyQE+x2lI6PplI6SctxjKn8oseS4s9z
912qEFmfilYaAhhLHxuVkVK29D2pXVXj6o6j1L2Mj0Q4NkZ2oezMXuCcgPiTjkUS
vvmeu/MYKtz8smwfSge0kVZcdnEJS0WEbbRDjEXNJAr2DM0n09pr+LxaR7rRxa8k
lY4o3eQyLT3U2qYyZvBdP9fz7BEpmcP4YsDUCjwy2KT1iynLy7SJIoF2rA9JbZNf
rGIBIhWxHY8v/TZqAtI4FNxmUGw01ZI+N0lfI/zj7/zukQLHI7gy+VVp6WKc/52K
/OS9/jhJUoP9vHouw2gTRjqVpiY1Wd2B4Z7J0yBs6iTZV92OAaqrzhR3q0csIerL
mamYN9s2Grf8vIYm5kj4uWxJiuz+fy7Nw5Fwnu9EmPs9iC1FdwJBhhbO9c2JoT7o
8IIGoh6JILLYPwE3jiOfH/Du6TEqQH6kSxCEc7utkCgxo//1scR1FRSM1jyB3AhI
+S4PxdvTb+qW2/+DYHV6Nfu70mcKYR3rxEy2UTtN1sF6OtNdu2daRsXy7fL98nxJ
V3l3LpUJ+v/KVFD4AGrS85Bn0Y+RWOOyphdaEBZNUytdf+383ffcgDOVsvusTVcM
H+6jLOi0MQuhJJidCN0Lr0SyUh8sjtxARbKga+v1Be3mlBvG5aPnudyJH5jor3iB
fNf5YCfPIHKiSLvRPwe7Je17Y6RkR7YhTnSjOHGzdISNJE60oqqAcBeQEB1cKTMM
PoABlAxistPMvJd9px6an6jtuRSRpZyqmXzun4gD79myVaGsXLxU7cBnegOOlR8h
BM5I+gMu5wICef3y5cqxb2U+hwnHTsmr6AGeEvCvF7JCcZkUYEgeXwULE2+AOMkt
cmWCfBqTet83A6BsqG3bkVXQdyp9J3s45S2idjqekf24lH+16q6/wzVb7Knmideb
m0CWs8WYxdwHRG4ZMqXwqTXLcIld6tzALt4GXpKdzQp+rQYKW6HxZ5v7qYooeYhP
0aVlkEGEY1sE+8N3o641umhZmYrbiYAZT0lC+4wQLNy8SVCwAsMESbKGyfy8TuS8
YnQzdzrNt0fEytoXmS8zFK8ZzhubYeXG7m3D9O2q8IEaoLBlcU9YmvOqDrydAxom
0nJVJjwyIGdbl2W7QtNxo7LuX/fSv/5NV1+lNSfbmOxSYTBJwPJZCzvVlBoMYKM+
SqUfUx3uZsh3+9cGQeU+ZNBDD+Ecz5lqk2qDWnIZIzIa1M1P0lEsultwvkzB6sbD
soCuHre5pobWAErPTUXsuAE12Wxxu+6UzZlrSTnA6N2dmvXgKovREfvZt3WIFn2n
4kb37++mvS2Lw2QumUVkGSYfY56R76I1fsXpCafCMod8o4wNug3G7YtkUw4nIv/V
bdnJ/Jo9F9n0SnGjJzJAB5v8+3OXVP4gKthi+AdOh/HMWE+9wwb9fdDy+w/zHGRl
9RxRm08bGr2ZDj56VX96kBvoaGZEA19lK5/iEjrsSdNv1/19PeWAps7hxk40B47/
ahohYOeB0hc/mCvLyCC2AF2kgzTdUCvTBC7kENjmG7Ay3SdCgVU+5wyCe1ZOrsxt
j7qPcZpkTbQKZg+JEXxr+fhKE1+FYw9ZN7O5mzpqx4emBoXllxBb3nMPE6UlaQ3M
+tsC+HxVZMJJ0hkEZ+epcCn15w3MWkOerwMbACS6IuYvnodBx260Vp/b68iq9xck
udDug+wyakNGSqOWoPr7abSMc2zOI+p2QCJ0DTq438hJl1mA/zduQ+iob6XK+NMv
9DPcL/cMT7YcemAd++wLYhhq6X2/HZlXd4j9GlHHK4nfx9av/7EjYpXiRg+gcrcf
yeM+jGXJ184y/asweQLs8GamwzxN9vj6nI3IuMTPeZQ0xPWt6CmIFQWuhWSgFVBz
iKnhKZRhefpPhjuO17APf/cUZ2UBUUrZomYCO68ukPaqpT8nYzvH6XZaMBAXa2V2
oan7SRbpk8Q+lcONIuUvCEJFkQSgQuXOvTGdYQKyHajwwWm5uFLPAXHXRsUl+zSe
3mKbdq4y5XmeZL2Ga5wRWUB6pDJhW+faermD+hnFy5z66p+UleUPBbHlRBEFNFe/
RLxqW+kRk03Ra/98/SbVENTv24piV4B7Tt35C4C9f45n3dXIpLZ2CbCGRxcg6lmR
9PzrmLRLVJbLcLJVldeHYXrYjJxLxyGjqDokzPRZOWW76VqtY2v9hILEKrp1ZEOj
vbCWmK3X/mtASyuF0l3l35a5x7Od8CgI31179NTGBkPDtyMMu57WHgidJrs8QaaZ
JJ5OQ2OoTvO8LLftaWY9iw6sgCxYxFXZH4i6NsoWdQuPV1IgFNAzExqsh6VGbN/F
uHEnVoD371qgod+iQjJgtwtsgnZ1Uo9y2T7TkcZvSsOFskFuux9FWcqnN2WwP/j0
FJiYlk1vKN3BdFWOwVNRjmK6xLkTqVBXqzNwfAwYKxkll+PB10UOEMtzBDaYi/Ne
hy9X2Q6HyCqcHI5hAxDUJMOTdVOHnRjZivgxi8GgV++M/3ek49QOd0SxvgGSzk+t
qgzg7xHv/Xdjz2U05dtXJ6/EKhogXsGG8J4ztB1473p7bjMu8siNtTULU5nFo3VK
9fGURFj42zgKtPSXNqrp3KrmGuXJu/PoWNPG05PlJCNU1ZJTPZSGehPWUkVKLMAC
Xeg7jV7+IOlH5pL7f9TAUQcfi2yiuVKA+pcgiNSzC4HxfmgI4kr0mtfAGFhSCymz
9B5uvaMKxbuNCGXTl2hk9THe1oqobdBTAu4dwiP2FDuTRiRiEi/i2X/I/nTO9Ahm
zCoWh+kLJK3XH7hlMvo49AvpCM0X5ooHAMPXXEkz+6a9qODqK7gB9ftmeH3nyJNA
azR/R4zXzUZjNH455oqS1jF3zgPFJEHlutB9HSWc46l3wGgd5j3w2Bib9gQwPUvq
8jf/bIzeodSR7ercbDgdUiqnIHDQ9zvhTZVaG2ceV6SgHjczVe9PhplZGB9uSg3c
l9zRTROec2rQbpxCLnPi56yUWoOT1EoMl7ab2tAT9w7rDiCA046ZOJNEjmnwTKcf
LXdYmj0is/75/RN5MQpxd4pi991FXma/QkzSQoCITlSXnf4YMMhSe9vjKs5QIcI1
eMMNjhunSYcgsNPmqLh02ToNVJg3hzCFcQ31L5JxriXfydR/JaXn27yX41vWmyZe
CD5BIYxlmCjA649SuSTNqCN3treqJjXlgBq+XOrMTF+LEerp9x7qnn3eH4FRUXIF
Ug5TkzYKkLw4GvkKjh0OPhxlldz6WWcF7+2POtBdF9SrvO1alYz+GGUsUdPRXuXP
vLg8ikTS+tT7I7R4r1K/FHXHpcccozLAz3OssyBuGtJtzCV5QuzmV4NDtEK8kYEM
7mtTpUz8hGg6LAX3apHmCYj8tb68sKbmroshRF4qcideUofJVg5rLrQU8ZPrWl/m
gxHn76h2IwTn6d6LCDC9mPBcq+rRscJDATyj8IfaHd/DKGa74O/ZacPnFEaoIo+G
FfZnPS9EolY6fAF47r7ZExGPaNl8JzJXItytyl4Fyk6RTcba4dH25vwVxlNkshj0
LEGQ37i4ednFqiAR1wx0RBP75oPwxgqVskKGw2nPHZ1S6E34WlGPW9Bq9pSv9xEh
Dxe51GjOOEYk6TtBwHX9wrskdZEjcbPyr0FYByBURxxETauh0a8RXvutnQiz48bN
asVFqb7CYlPBzZxJDlp4YORffIKhM8D48t3PO6qNdVTdnhaZy5miQU5IJIfyR74+
gWvuKF2ds58O6sH/NMcpMW+lelU/CAZqg7FaXXfB3lhjotQTNKGmpeSq1dwjSBjG
A6gnJ6v2y3mXH3iXSayWPYPCfIk7DVg1hBPIy4GPMxEhPqyoPjo0AP6gAeTyO96g
R11uTdgCNdpWZp0wJcjbIvlyqJGWXItiTOSHgG62lW1V9w0y/ELIJdw1uEdTummw
YQ+IMP22MoEdvDiEJBQyVXQ8CMYME7ObExrYthOWmIS7IQZwluF0UeTgXlS63fqp
Gb6LnVGS6nC6BkVKaiv33+vTdabXeIW97qU+2B+Pg+B1ZC/OnUhoweytbCA/nLHS
7we+aJa75KYZ2tPoJoGj8XtSmUiLjYGNa25SRC7WQdXrkxKmOueNxBndD1Zxk5jr
SVDbZxzYovueJRPLlhAgAGauCWcgZrzZTZklubcvAHnaYnFTk3LMZAmsl6bmcnZt
UBOy0Jfih1YpVyLNgFA101aEBL39prNfJtTVKC54sS8pXsunZWsxz3VfqKkwBuGP
bLdbZEP6u7XvfMn38WwVa+/iB/KWG17pNk8oAbxDWAwJVAQWUWp/mG46jQaAnuPg
LIDH46pvm+p8JAv/Q2jjHE3LaLk6JUusoM8UNTsJfe7D6k0qEXsNVN9g7QWCQQHY
FjcOw5PwA6VitsosL0Onlj66mOeVEvAZUUvruJYmalhc54Y6+LvU8sFIeg2OcDSk
Tkg60ys+jLdoAzxPWFPCUkxgR9GN38+XEM8jXHRXY/A1jtzntjO709wUTPG68z/g
HluFbn4puntkS3hSt0WTxmNT12hQc1lmQHaArDVXM+KsOFhYB3M7jJPpctzsOnlG
iCQrW0J0m04njAphNtbSPkykewRz28MiFbmgIf8Ty3BCmTFfL0WYnsDS6/8oo33b
y7WXDqQJwHpfWresdmtMUpps3U7MfqUjJupAdjv07crlncF0RBgsG8ghUXwjMm+s
xQhieGXnMlfixaMCOc8Rz4gE608rd6N8DjFBFYb0cV0+e2p46E8XRHTeChYXeXVl
MhaI1Xs9fjoDhAyWmJ8K/vFM6yr/XJE9LdQ8UeY2560Bh5yaLvVgTbjA8OoJZ1Q4
4u3C4oytkySRTl9wT+uKQUxXLfIyQA0Z33R7kR6I8ioUOVstmdZvcsvqIst3SKFR
LZ/7k+TIwZQLj5aCewCOpFHWrhfvZ9Qa6zg/0K1QRZjRrLjpSChuw6OTK83NanFK
uogz+E6EiHKvgnAKi0U94XDsmCtyarRU+DKwyYX0poiCdqDvnNzSvgEes1244rEY
K8wU9ymONV4FR6KvRRa6rr5rnWyYiUAlpNFUa1k2WDCrGu8QCicIykgchVlLqnjy
J73gToNkyzE6MDb5zSQ4xg9oCMVKm8Dppt94zGkX5TOxRvj0QoXqvMP1JuApjOL3
/lGe056QKYLONqewWy/0cwMWnb5embogmxf+u7BE1ausbS4GpYjEDRggRn2ml85/
kkPGOVclsNPTVveLsPhQdZYVjGf51/K5Bw09esWRAwLk5FxjrpX0t1Ue1zRwXhNh
T/N0tJ48bwr+rovhXP3yA/MHGFjlbWF+y3zKNN3fvwwn0XVB8ZIS/BeOJLANo7Lz
mYch06KaqiLXVpRRj5nIDComl1Al4HEHQn9Up7g184PxN8m6/xyTvxpKLJLHP1PL
f0e8ED20nngNW4Qkgz6DdimanGWpfsUYzhkrK6JLOfXd+gLt3a8ypI9+N2sjor3W
u79hQZGBhiGHxV5DzBNXIfrnlMpRRQ7rgwWXj9mRBR5mDX3aY9KxdL9gUTiKHlAl
vjOb52zj9XbRmuUt+eSOXorpHozfWWugrujMZ5q1NIhZpvcaoqpXGU0Dxz7FrsFR
2OAPi1+SzRt/K4f5gWXDF+P+0BvGF7PLL2SF82IZZjBH7lp0PdjvaKPyMpCwwAeU
qOHCompKz/AxeqEsd/lkkkmNMPTgGgm1kutJQCWwZLb3zDOwk6Alf3oiy7SJt7ha
YdyPlD3reuSZ6wA855IOXFf65Y+EvWu4KYvwX0QBvB20NANomPTRBtTyimriJX9p
ZleuOML4nkWgs0JlDuwEfJ46ywpBrEyOichY76wX26zUR5Xy4kqrUA7q7wAy1XnE
RtsRTIqLmXfvfsgSHgfehBl0bUj+veP9lkgjlV8Nzf+CeSvZzFqIOFg+1RvZV2AN
CPpozis9MN3gQiYMlnNVkFDElV4nGvrfS9BYKtd0/WqtpogvBfdlDcGoWo13Cnzw
uoYI1aC4x3NXvTTSUfvRDsc0Fm44uX0Xev45QTAwFRlDbMIgxv8ekZ9VgdvCWzXx
eHyK4HRyeHiAe8iACsPPgtJ2f407wR94lbwzU4cn7DMqhlzorOrJ5qFZadKzWkd2
XApi1IbC9RbpJ5k4hZdnYBhoYWaqrKZ9y8e3csVIr2p1dYjFkp9fMx0tPqwmDoqr
TFMragEoIzf4UgEqxyAM/deWdDNdhCj2WePeOL37eYdZk7Pu2GXJg45aPSqyrY5/
IlG6XlTurBSZ25Bcrmx4TkCYE/E4S8DWnTttEuwnWiTl5dI1ebhi0VzH74MthTN2
rsW4DwruI1ZxVGyJqToUUdJgtq8LUvN97qgkjo1OjiWSLW8unvgZSIZ1pIDgLAo1
YdWVkVdfcCNNML3/DRDUM4VchSlPAFvYt7/uHpG7DMX3AFf+im29tkZQa8DlRIFG
AGFBRbmCOSTFTOax6mID3QkLaRVlDHWWvAlo9pathupdE8vUJWwtsCKopXMuFEi0
ZA46+trxJLE2UtVtZd59w276GhtmCS0jrFFVkBVPJKHZ63x+gmV3YqN8fsCVZvdm
6Ba0QZu/0DIsPUjvdOb3vNN1Qgn1/5xLs8L/8dBUIpyPXAg8IOyvnsNzjNA74VSs
2KgWKu40PFv4oqj0AzYuTvnaKTpJtKXNEw1u8vD6IZMQHVZPGdcTHcYy0Ijx7Aze
2cuYo7wHCa7GD7ZCCvT4vB670CK6m3esWwq1LS/zagrSvyt101jrIocVR0M/ffnX
ptANe2ZbATtqIT+bCaadNZc+2IgRt2Zy6YRqn5KQLK5nepLZ3emqVN5MOKQqRXox
PzpygEqCfwAXOH3cRgP3fh7fQgbq0Ayj0UhNYv3MBnyypgGAlg556AN6cotkpjPm
GWn0YjL1cCaMtsq1s1TBLCcKE0WOP/W74uO0OUu/D4OD0kkgV3ZqSA93pTzR8wNa
CdxXVzsddAOO0EToM6UDlc6mwzGQOifjGZoqiuqM/Nr23psnEHcBpaxn8bBY6CEs
m2pWElXFTqvWbVT00cI62VYQD8FkAXeaURFBELR8nNjXKixRX4QtFNS/mvyy8LC+
ezFT7LSRoo0eRw0205wjal0ZpPrcDO6FOBkPQ145D8I++SZkP82MmOscEWAajC51
1Stn6YKyceRpxHRgVDCRwkG/b8SJyqlT1RbuhpUtmNaqzUJWrnTSRaHXtKlnPlZA
yriwX5sfQ1IVfVF7gFbTed1Bi8sezpqaQunCF/KtpdQBzxayafGYQogwygI648sc
2vpq2DKEI0qPYld1umYMkvHEnz6aam/htvdCP1Q25YLQFfY+D3ep54DtCPDKvaAJ
zv4bBE+0N1tIEpheYo6jCIa+25sx5WSB6aVMg9NMd2zfCPlZkpyvany+Y6vsmtIh
R9qiuRqA6qrjMrHfojNUKlbjRh831YFsyGHIMP+QUBUrPZYkTIpugly00EDfmwsr
U4kPY5QtBmI8K76LsybJXptXCZT3XM557sqlltG8akGQuNNsLao/d/syzmA27uH1
tX+Nff5zAj5kQlk34bl+w2OOQoK6iJa+6IrkVQmYnusTfbe4wN88JSqMixwM8oIs
1XcWZvG+1yW9wVcUY4LePtrdv6R0vy/oyGQQW9m9XgxUUj4/E1ERC3cuJtSmyDfZ
FJPhljD8xbw8Kesi+iiz8aZVq7VQ5PjYRm/9s5uZEpN8Nd5qQmIS0a9eTDtAyKTB
zgDtmLpHMEiX+RZNudVQW85xCywl5m4BN21XtAl5HUYDaYQjl91yZPIPYOD4wmKw
m1AjcwrJ1iUWny80O6zkycT4jwIkGQl9GPDj+RmIoPDSij2mFmc5HEPXpaxiY4x1
cjOlkxnk6wUdHXxbuja7qE05HjF0DE5t7WNhMEru1HugQifIq6HYOpTf6Al1moIo
tVKt8wz5yw7Qhl5eCarWHVTiWNenEGdzIYLffr5ecN1h/VjPPi6tyPKJUz3tzNQQ
dk7H7z3C9DTFf3ejqmWsL318OpM//LXWJjlklwmEomkbA4tvPYpF/870w6/s+ATK
tcO0cQQFkzHn5j46KCVC2a9jTEyZWnNV3/+xqoRYnPfXjYtLl8zikWHqiyr1cS2w
/GKmFnnlM20Xb7tdtX5O8SYYdmH31LmIu8cV6MCeyezKR08c8CjzKQZypz4PcM2j
z/FoZ1mzvCsoKGhy+hL+BaRK5qMsegi97uCPB8tlHNcRNZNwCYzUU/YTtVOh3HIX
/AX0AwlSJucRYnw35Khy2oD5syjZvk/7i5AWBRVZY1TtzciXqLk6coxH5URruRrp
MsS2lH5fWuMlHePw7CsK+YgMcx76H4HGc+4AWXwmh8rUo5MqT1f0VKFOwcwHL+m9
sonWDxqvKWPqavX3X1I7ozFZP8ToLnnBi4Jvlf5nyNnKBH4lnTrQX/HMNTfDdy1A
ikYdzE+bBcHb22wx6nnMZpHp1VRLsp4/dS7jW6F8iE/v+93QJAu06O9y2rWvhVDc
c9NNSay/tclVJqMJFgt21/yq4In+hV+izn8PkIxVqQm/ecvHwa5KmeRE7LeUrWsN
ppQOdN2Q75HFwqzFoRij0Kiw3WIVFSZXndxJtOF/fniQQ2IKhXTijHOULUznKa8/
1/Cpd1F4Y5xOhNkt0q3qmkNo3EFwQzjnr22KyAwYCTQ+/HglOVKV4PTeZioLbfeP
ddY7FwrZvDAysOifsjCu648ghi/1zx0ZpeudfTLdlZBe3wuEOE4MMbEC7YnufPJU
akDc8lgneVnmkRWqwEpHAHF4SEndkqbTsg0WLvSmPDVmd1IcBGJ4eHefGe2i+3jb
B9PgRC1NQIyIWiTj+KHVaaH/sSIih+cM9QZRxHsFQf3dE9fA4/193fw60vHcJroj
GHBLl0GfZ65bNb4SVxFd823K9KVB00R+cvlHi6nE8HKTMZ8vX6qTcp6cs35k1k4Q
mKBia4lpdrwlcgVz41m8SUjwA+nUJcSHlT2kPmqVf9peK6nd7BoHOE6E++FpP2qR
BdCVWBrR950lZkZ4sIsH++V5FRxob1MDBVVwNHYcHO0Pj7V9+tRk5Sq3tmQ0WCMa
psK3xfe4pTY+3nhsSUuSAAdssxsmZDn7WilgT2OgaLR+1CFP3Q/Sfa39gzkhxtCi
s7JhEaeQYLpa06Bj+llnTqm+l2Q8pBcAECWUBrohpKreCfTbo/aw6152tPjlrV1R
n4PXFkOe5P/XocX0g5uYpZubKX96R1DFNGu/h39dnbt9pKTFiKrVm8Rm53/wSBXP
dBemKjTREa+Q7JhPjfnoI3VnrrOpKqpMA/LbIDmpAM2HyOvqyNMw0b8VTY6JVJSz
cDfrdha7rw24tdSNFUOGtbS871MjyX5MyZStQz+gwaUfsQEPkPlu1Fmc+L1ALlNT
nGpJC6ieGVNoHCgODsumFMUOIngZa0ltXGr2SCCEwn2XMjhCqJzzql+3hoJVqira
weZGTEo9QOWu857vUvxNtBR+H1oyykZkhd+o/2E4GhgsVbZHv9BNQP4gGGhECDnJ
OB0OcVw3DAbKBj+EqJ/5XXYOX43XyYcWrMQwT9gruJIvfFnLyj4L89xHmGKoVQKD
iZemncIfS9MehwZpxtTHKUcBNN4LfK8bvalVLAM814SywyCFF+Tt7AmwxnVPjuSY
cSIay4+U7mSkoa8Nwak00YclGgyYA2cQkdk+Xo29kV5PZHsqsbTwsfzJEaq1qo3F
WCtiT5DrfpbwfxDwfskf5XuqVH6v1P4agMC5mrj1KB3Jp7G0X5hPePG/4uu0Gt6M
AU0kUltetEJQ/0j7RCo9rQK14slsRIbe4axq7oHJCeaHFyiO8ce7lZrvCanjNEKv
9qLzFNpAJyy/qn7ll1imHhpcIheaH9sslLytmhtXtxXsgiTyW1Cdk/BcRzIZRiTI
rkrh7gLlX8d0fLaInjxVyG2RBGCHMRTdH4w1C3g5epUudGwIvmopfy1qHlLWuITb
8u2RlJzU5pYIIw6s3m+ZtvxWrpJ/c2sYb35P4cHa3LNWX2T6wztRG4pgZnm7P7Uf
RzP4dgpeyYeCmenSE8tNPhdn6dniSTWVy+0NzES6+rQC6Ij45QnqUyIv+cgxHoeE
ZEcfhUaONsuDdKjsnWum4+4GpnuaSL4qj9uvVIBKtipbwhhFtkQSXlitTw5MizIF
++sdH65vATy1Ih2/n1Sx+JaST0sQ//U4yI6eN8BSO7iGytEjwyI4DiK1Z4uIyh0f
zteL1o4X9Cau9qg1OJpoQVR29PXdslCtTfm+cGfCCQOO1gSpy7OKUn6YT11ttTlf
rU6lK9gkDQQEiJ17ljUdu6sZ7ecvIMk3CiZYCsTZNRk94gSPdG+fmnTPIfu+ieCU
Gena1klycFWeTqAKPH5j3scLQm0xiRK4yvf3OBU+gE1rI3V6iq06lWOA9jus+KbX
+ennypvr9N2YsH3B6gF0iFSjkY3vYXnmZU5et/GwCQ5JbcKFfgMBDVevFZe8rC96
e1OR6zpp85BfDKc9Kgzp3OZ0OuB427rsrJQ9BHXbONt50S1jRvbrSO//ivA0ZZ57
XD2h0vLxAYdugB6hysKna3yThE0CfzPcWRlmhQEGI0+czh4krCTIMZdHOIWNoCGz
+OaJTyF/K7h/rC9zc3/6IZqNE5sYrMYerL50o/D18MTw2TXgk4+Hio2IBp9Bh2En
JnUzqfcfGWptym2fGkxR8GnzOOqTvRrZNvGhfP85wzvgJcOwJewSJh9rCLJdiEE1
rsw8fzopJH3HBeNvj8u35X73vQLpx/j3JK4udwi81rrth/xyiBZUYTFJMPXTnJFi
bGN83d6vLptLAiEJSOJvBGnvTEcv0Zh+/od2Hc1rJj4x9behhhb8kvcLnFKrsOSy
WEQrPYZ60/jKYfw8r8vE2gmahGf3a060TM2msxXfhEXOEl7934NkA3WOb3Ysv44J
`protect END_PROTECTED
