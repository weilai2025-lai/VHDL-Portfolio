`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7n5TjQZ60NWHSL9hLsxmCIeB6Gt+l3gFPW1h2RSDUsHEBmveW+bJ5g9aNtRUmqn
IWONXmsfSJGoSRltv52gUH8SkK0lXl6VovcM2kfeMDMZu603CL0lANG/yB9dB1WH
15hrNLPNPuh2uGSp4iokqpO4+d5WeoV09XKoaeIzjnaPyp2vdM6oSTPaT14hy2Zt
KTYSZKX/MLgaUGSQchoNRCZLY85ClkfaACKPbsYh6RKk0DMYjy+4YLItEDPWFsX5
Ybknod48W2VAg60aTsrNGfwm1ySe89GyxQO8db+VLPV+tWg4NpMLcCZlTm0VJ5C9
1LwQ8+4dR3RNSzVlodDPVdns4DrmHcBA/t65gdb2UINrTYd1b93dX7apD5H4KgGB
QoEPa9PdnD/tGIi0doUMXevC31ZR75cCGadcUb4UH+UsIzS+qpQVdV0QpBjJ0WzZ
zZinHND3yLntRELGh4d4oycDmSgpjBsfsMAeDsl7HyOkVjZZHj7VhL0jFJgKkU87
3mAlQ401ejtLtzGy93jllODNINI+7dNg7C50FMs7wMMp3Ya0caCrZ21aDdjtcRsp
FBQjZuzu/6hZlFD63eQ4p2sLlxTtbu/4Apqda9bOEX/3FYBVfy8PiAm1Pasiy3dp
2c0e2z/01Qv6yISm2Bh6n1ZTOdFGJGuR1zN2aNXQSHliMRDXadKe8GCcnGlwC1Q7
vVG+bNW3MJAziTflYi4RjrDuT9lLzhn5wxyjW3CGWTg+xjets2QejUCGFaCooC3y
FH7RmukUzOj2u6LR0+FLxiudqvENZSJF0A1j6789tc8yd4Q+jn2dKLRCvPToLQgW
umr4Z0DL5FdkXeW5zonv6Tbs53MIvFJVghoagDRQG/uLrDCAoom5WTf6u35P6xwa
LC9CfBeikVKaJ75bGvEzu4GomYjtEaYXm+oaET27wRH6IMPWkIt41O2au4sp3Yqr
IOCet6YRxmHESZMn57R6tIBlkHUvd4uak1INYzUJAzgVsGzCdqRnoOwBxAtxD7Xp
dCRAfMW2AQ2yV5TaeqVbKW8iVUx7Z/FvfYAAD8oqAGHQU/Mp2qP1D4gwTuhh//IE
idifJ1VVAuXOi8usinuEuopoZqARZT683TOjHtkjBU1HLoR0YLqpsMnBGGMpUdVy
JpZm6ARct2HL87JqLtbr9ZAnW7JTQNpduqGu+kYHXAMmBsb8QRPO1xSuPWZ8z23Y
NT3/40qpYYyCB71p2u6xVsTooe80gfuh+ErxDxkuASpzAj95Hqd8G2kNkGwax8KD
lzPJu6IZC5QLvh6ZotkDDGfCjj4Caf7yFusjhWDg1e1KQSKjNGSLEEvIenYmVsFm
KKj/3+J4O7mYt3O2k9mdbryBZSZmq9xLC2LhxbahAgR6OVQYOlry/hv1O1h8efUI
2RSSKrM8WWpaWoilZp2Pb/SARNWVkNWjBERm2qQAvUMrbe762HkCqwdaYyd3u38i
zimp8c4bR3d4+D443kDfKc7uqOd202aH1daDbX8juoeNAEVEgjRjI4pfU/5VAji3
/Z4bZFyqdB+n9y/yb6oheg==
`protect END_PROTECTED
