`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/fjabmyJBxOJVk/PprcO6oELAQWSR6dV3YyIBp8nYR7PvoelUqVx906MOE3xvJE
JwISCbNNHvp5qwQjToH3fNGfmsqk9MhehIlt1a/HMzxlVaKM5oJ8ZuCgoTDJ8D3G
AFA7/pS8wlyKP7DRe8zzP7yuN138c8zvtyNvvGR8seAdiD5zvvNYfJ1PykJslMtg
Igd0pE5yvfGAfzYEdTXN2tgi/tC+e+YdA8XQIithAR65IIepuvjup6zjN0kPgogO
2flLMDZEsYsE0lVwTgUMq2QVsfDxdZHkgJwE9u/Bs0j8O7hbQJPijkVWaM6ugG3I
90ORkKsb1t98+KJGsmjoAdHBIC6eglhlh/I5Mm02vFNbcJRa5NCAl7IG0cvKbygy
BvIzCwfqqmEYXJqai7VofNEG316G3Cx0TJx/RnlhS7aKCbg7E8srFT+vyJYlHTlq
L+V6+enGyQcj6bWTQQCIVsprRPqLhfOueV+58I2RnXOkzuleiSz38+PxoRsaHGoS
p4wD8t7gK9qDfkFC1AQw/SyA4wi1xuTG3SAfLZjx2RyI0AL498l7mHwdfsmCnfGT
RXVppwmysWhwONvDkHSRNIMf4BLxpiwo7GkqahGdcjGcsBLa2aoo3dvajN4Ylq+4
ZBii2gSsCqaXTd3wTm6u91y/c0d0H1kaXqFcWwWyIMmi0f6/y52A9wRPDszoO647
J//8ZhfbxjDCbAy+9gTo3n6dgzcFmEKwbLUr4qz+ZFUhx6zd9W5WCNN1w0rFVph7
j0m08L+qHD++J+px89DO1MiFLY7+P2EflKPz9rv7AMQk0urhbboColGh9MSXVgAT
7rB1PSne4MrgalNtt8nwKccbXcUHscZIwZo7naaxM3gf8kdG28lCCUDDNqE1pooT
4m97s0X8aPYkjmRO6D0T/HBdkClu4g90rTZyQC1gO0Duq5ausjYog5Midr/fX73p
Ruc7mRr9ph6EHklRuCfmm342b1JDu2ROqp3JaJobNCxITwNCbVX3gnU1QBhVJO7+
tI9KF9qXlAxi2Vu18wSHFpOFEqnszW37DcPtoMnziUbxhTZ6wsWzhn/CvjxkLema
rGT+QFoDjUTfUGAbU6R0UvmGT82FpubzvFU4arV3uyqLMmOrCdxg/HVhGl/0YBb1
OM+qPXbreK414lv0IlIkBLQ9fFm5evbZ3au2B3qYy3+/ufecQIa8JChGdEsLhDOx
CwsBdbfiH27+DVkUNXwdPVPx+WtH1UiNlHa8VkuiRCAmJtzDA2BYPtFti123NTxq
TgzPOtJhuCLLPuSpJSyH4S2nWyJIqNIFoA6EpDhisU5K6HSVW0fVK9P73/RpjR3m
7V7REGkjsVVA/kP4xFh6HSbdBYU21+kRwSDf43OTVUT/pkl6zEJ3JHuftLIYffqF
MjS3SrsT/3obyWN7+/7Knf3L4A+GGDPCMFtF9kZbrE+Ojr/qN96ZkBvGzieNWqmp
Mf/fCItKqpMs0vCB5jlGr/sXu+cmJybgaz9lTJxqh8LI/2n/RS+lShdfQMrN5z6X
oMw1idKpqpmcjfwOKod3BJycv+rs+C0PNTSJJHwE23Ix73eQNQZJiMr81y6Ya5R/
t2s3jKsZWGHikeVAuixfSSwVtb4a/kHxVnOmmVBmg6FckHIRvARYCUxSrwxR7xpf
D2pXaBWwmv6ah7GF+ElE9JWerm/iGNzdTOKMb8xyN3LBsOtl3emmQauuZf2uc6H2
et4IVhFtzIa5FztqBW3ev/kKHW4gfCiOSZmyvK2q8mnXvqb0wUd4V2/Blr8lmcqM
bSu62eV5bvlsJEOfHZ+6HRW+y4GAjUffszgoBoPL2gxBRu5sDc3X5cHAXhTmulgO
DBcBDe/yoJhW0WzWFHDNWQoRdDqzmsIQm7DNqMTPU63DUbcuXuW6lUdOE5ZHacil
+Ef8gziyACr0UadJRFH7B/xM+ksJcSNCZ8ycPYdkxjlg1CzDwIoaC9Ckm+2ai1iD
`protect END_PROTECTED
