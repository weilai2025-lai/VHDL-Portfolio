`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gc3nvx2p8MK86t22v6P/bNvdFr1uOs46f6XwzGnnndL3A2R5PahhfSo/ubgwMI9
OAyoaZk4cujLtOsxcqc6A7iMplESuvxe49GAKJj/hvhXYpWM9Fc0ba0FR0ItJbxD
FjgZf6lsLEh4q8y8yHDfnl+HBnVd8VyGdbt7akSQK0AkeO9Qo7lO4S6pWKWFBgBU
Wna3BxYSAsL2BHvkWAtaVUw1iiwzOO3x2ufH0fPrwDk66Bg9pXSmzbAXWT49SrbA
C6yU4/6wlCuCU8oNfEBI2AWY/X8CHicT4kqqM7vglcT5bxnzPwu2KpJI9HSfOBBT
GJtu2hQL9w9yjo8AC+Kx2k6WmGzOiUi7j0PiJaqecbuO0D3RRTyaBH6OLNKlJH7c
/SlWHkOjNZ5jULLWkya8prDbixXRV2twbFyoLk/SgLN6YBfCupRKguhaY4toTc6m
SO+eBVGv+vJYtU9d86/dI2/74ht0Etnd51w0HaKragLHxDHe+ZWngWGKkhJQWHci
buPHTQv0osDf1N2ApxkfnNltXXfcg1iY3Az742Kr7R/36nsYYV16njJ/ukBNJUt7
oZRZ5bseLdzvY+S2JQvg+nH/1OG45uYd6yUghUxO9Zw/ZRJySCGDYwKFUhfU/1Av
6IBL1Q2lpBDIs12Nai3HTBc+muH9WTz5ALtw1K99LCz6xIzKZqs8h6gXIMiMggG5
hdsXnY0c/ad8gYN8wAxhZ4Yb2lJiwEC+PrAGFSfMJF70vF97hWZLDmrsGTGM4BTd
azrwGPKBEXsQ8TUm6aX3M0bEygMGBZhSCEWGpE9QEk+7taKkl+uEfVRVwPswl5lw
VVLdx//hiwlXhqtrGBfmffVUSHREX3iXOyfUnm/fvv8=
`protect END_PROTECTED
