`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Se7fJVUHOVger5wt9zxIuMLb/9DHVz7zNwqV2cpju9WLbqJmHIzKQgntBZSR9u3N
owJ9gnfeyI2CqB5UwAO+z6nNgnLT7elo/hZB9Lm3lq06U+FwIaBkyr4MuozKmpQ2
f+rroz47YwMZdrIRG4B1EtkfeVLvKqg3bczEqtJvfvyXluqjsyHVq2NUAk04YzKt
ZT31wpQqjBjGDzqCKe0NbWHciF6PjnsEr/tjAdsrtbBPzgKPf1uPFT8JX2TW1jKq
ihUwTFdQSvsK9ft2YtU3wjlifsQ8FyzNTdVMSfALW7Oy256sJjZojXOtb1kuJKB5
G4J53KHZAjJy8HDvIY3j1uiJQyOq3kjae66T3IcWZdRxJ4w4zrVGs1PL02vzqdmd
blfLioqfEzHnQeqOzaIT1vuUjQuSJJmbtJ60pu/A7trcKw10EGtcbx+yMZy5usNN
3eq+g3NWqCnC2/ukgyWXHFfW8lHT1g5ZulceOShJqIvaOT5BB8JZHCGhX0VGuLf/
1Xop7XM4j1EhodtelceA2Q==
`protect END_PROTECTED
