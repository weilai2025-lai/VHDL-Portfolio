`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VL2911JV7LTvGb9uHLDtUrhru+oHXk3WGMayiP3VWb44FANRHQqFX8HiGLlXLxuo
+OwXKZ+zOMkWNy5CF6q101mtvC0jDvMIZI3kl3OEXrfv6VtbfkmyjiYN085ErGM5
VPg6IxZ+N3QyrLOPSmiLcJ9EmUazXl0rmR5A59NQQsQdrdv4hfNYF3ckIHcGQ1Sh
Mv7BmjC1fM3FfzibbwUDq+iZjwxtK+V2UPnmgevLWQHo83WkYZusQaij2vgQ1D7A
z34urx7bFaFAu+2zpBiVCYAsDZpWQZooOcFzKgLHymTg9f6NNm75tAU/xXp1ciNH
+CS/dfybRaLqvRQowoIyOD1+aKG0cs2zsvIpaNa/yilJz67bE4JsD/LQGLAqwh9z
76Zcp8THBJLyVqH0drWAJqH7rjeV7Rl7blwU0kznIbi9phUlyw/o/LHjY/mrxQSJ
vlStgPDllPNt+VtI7TRUukjDV5rRgJQmKlCTV1UKv9sKhSGMNDXQ+20wycIKM635
kwuZxJHzuqnxbwiNvt6YL1IlzbV8rRsdRKu4r05d2V4KpP7t0Tuvst8VRHpvAGw4
ih//6Fb01DUt2nZQIQVyGCRNgaAhGYLuFXtiuPcrXc4gTdkwZg/M7TVPa6MI71N+
Yu0DTkAqtlJ6K+CA2kuCd068rcf8ocjihlzCFqYl8IK+muI5Aj6MedB+g8OKCnty
SezfXFNdrEbUuuYJBYVntA0aS7LHpoe1EP0MiXoqh6oIa6qke/PlZHpZwskIF07h
Jl0r/ARh1lH6cEYWvF78ZZu+o+5i2g6qv7Qabk+w06QfWK82yXvOIgWgKGj5ocDn
wOgKx3MBEyFrWOBm5F2OoGzFTzgcxf89TXbOPsmF9kYS14cgl0VNlVoKth3N+1m7
U+8gHV4UGBIM9LNiSD3R6QFpgpPdRakfoEXdi3+/lH6+wHY2POJH56RrFcBPzguD
WvmgrQkFVsARQJj7oSbEYznBCvZwHRzn34HpKS32lj8s5eGxoliFtPu2WYreeBBF
jeglxyO8vi5HIwH87Y2TBMKQcqi/sUSZmXAocJ7jaLjySKK7f/zYwWJHGiUPe+wW
+7ihX3xj7npKNkAubh+kzCgUQtP0bOIJMQ78rLZy+FZSDMqQfaGQAOyRMFh3wzIc
5piXSGXlu2gJ870tU3nzv2UF93VBZ26tOmEo+22myrlu50kcIRfkLtqIlW6mEjKG
rQuaNpXldnUWJvSa85sKKz0slIJuq7Gc7xKCzXMQn/LBf6WYJ8z1I8efpnsdcYPt
F32rn7ffuIm1XQbM9TGBt7OZRtDH5qcMNulC4zpeFkR74+I1BnOOvQrrNTf4RDAX
wq0hpl5/6ZfkMR64jJuSzv9jP+NDz/t9ZEC39LTbCif4MX4NNs7LprsHdn0T0i2o
gtPJ6xOqBOzUhNKfzmnqx5Z7fERkEKJK00KzzQEZzH77RKsHUtBEKzaRkfNmvgT9
hDwyxzTcLKqlFa6pqwHMM8Ud+tQGlA56xB8q6KCSTRTxDUPjwycT1o7SWiq2cRMm
L/RSGcGQO2LM1UULlg+d7ZzOnaKDSD87aOb6LrN4F22I59mp1e2BKfaryBivkqFP
IZ8T578OZ+xPcm4iL34MKsuaCeONtIwWXGXG4PX0iFl5LTK4C1QCD7JEO4nOnKZr
gAEJsbWhidiRyqcapolIBtqqzdWESUS0f8egfBEfmCIDCV2HYcEsy47XwZeOH2KO
UcF8wb5pav8lCaBryqvZjV5GLp1nniSr9IDsEQBKYW9wkxGZyfnrybE8mGV5+s9X
+Fr2K55I5bYZAJtzxmAMbwMOIU6GDnO2KFq6hbck76bTO94fgNfUiiCy9EOFr69W
Xca6PlCc9BZgCu+PB/no2YwbkB9aaL+jND+I2kGI1w80DRTtWh/CSPfl+qxDbTl8
XE86x7Vf32wQyU+JUpntzdadsSBWMyEswgeqcHm+dPgugXS4P5LNj9X4fQXkglz9
7PVs2mofqbN2q8kPCpEl+pYngm48RZCZh4Rp7ZBfCGcwZCyqDfxqe1BrdvuWXM+7
pVXBX+RHgeNCXsvwycHrTD9nk7mP1bufjhwOXLPI3z/mKwSZRgcHoeWgzv2U8jA3
6Fbi7/+0+38L6pWthCdtWS2xCLYrLNMj2KXQTzLEb/iOFOAIkzHLjFAEGmP/SLAj
0Ta/Xi5BakhOgbw4WC3d0SvffmZ1wVfxUwk/5rDgiQbiHVQRv2dC98DQHgk7vsC8
QKtx+5EVBRwbZZJ97f1FqTtiO5+Ko/Fuv2HvQG2a8t1FhyUjm7eVQ25whUT9aF3t
wxX6jZPDHSFVfRaCOxNQtI9uU2l17kewXtaisHqTiIbWWXUyBeQTsFz9Z+JpED56
8XzGet12D16gGdPDFbXcvSBO8gGXPV0ub7Ajlo5vbXmftCR9lr7cUFmRhWAuUAZN
R3OBOUI8dRMKaaPUnOUYVlwtPI/ruxUy1HBwPxYEX23UIJ19TgL+ZLnh/0iMvCJJ
sh8fctEg2+NiIQgA10b2Bk8Wzk2EOCgEzqnoDnP0PuU2Jy5tl0os8tDMd/PuwqEp
aOJ6WsqYtj89yEKENJEeN8QepQTKU5STisiZGPRzvwTIk7sH26x/OHs+sNxDKUqC
gKSRZ80Hhoufq7a9IPjeSCYXvpErjCbWyyJKoVHsXZM2tcXs3yd5YGpBWXxbR+Jd
tOrprIT1vz8QhsfyurAmR28AZBLowQEhOYZ2agKGDyYOqScvFuOTrwcCS01t6JXz
Sn8R0uJxttfNCYdgY0F8vsrF+P3BZ9eZP8TlggANrRKcvgjvFXeB/otTAHNebXTt
hSu+mITPfWaG6fUfIbwiuocE14BLw2t79QpIfgbp0o7zQI2ai0Sccxpp3uNWgjCL
w0UYv2H5cmXrleq8cMDFIEt1ftwq4DD4EiSYDMwv9wgMuKFwv/guT7vTKKbqesk0
NOhFSyLq1lY9ydB5RAhMtGN6d7pV73xwkWqwgWUpXRVK7Eg+sI1Hca3KoDHRpx03
zF2yDD+77VNTe72LjzUymLA/aV9d9scO0Woso0hs36mDUQU1WUGhRvlJwRKwuem3
WCEIzc8Wkv3V6BbZc18rDr7QgRuPhRsxLd+kVykEU4UlsDPNVUdlBQeUE3IBkGSt
fRBC8DwaxAfMgNmFbl2wxbCj1lK/Ffgyy1XWbQwYeyphhpoHdCsRPZIWfNSuDqVB
by71W8HYC/T7JFkmRtFv3VE2U2mCqx7bBBrj7zeKg1cKa3oYzrqtwz22Cg2CAoEy
pX34ee/ZUj42hu6P1EDn9WA/HXgXQxYU/FUzS/FzBuZoO2zDIBRZhWC/3Z3/Vnla
DIcafUpBkn4ySI4Xb4JnQuYuQKWu5cUMhE5gAU3pRNWXx1La8Ajdife/TBHgZKnj
DRSi6b3s3wwBlw4QgTXKCTXOn3fkxxfD13LIX5K2RugttKIPgfWN7sDl+w8bQzua
g6Soxq/Od64B/opn6uMHzOObAItKWt/Ij35HFaR7P3eUoPxweaEOBuWhfWe7dlDO
Xxd0G08MLig9RFacs1m/jIkebFuHSbbacubhgbH2zVYQyY1rGVx6BqRzswB7qXd2
PLwvhXe3YmGPYSoxdWOh1e2HTUCTP+k1g9w99fa+BmBwOaVPZxsHVYf++ocLFJ/f
OJAqelVAM2hD6tdAik0AlXls3oQql84TJmlt8JQWeEgVQPVmeM6bRCkhCqhzZKsW
tJLpmRIND2WiLLeLFUMfhumQ0YUbiwDUtChzz0WxOdXgptWalUzs+mN72xZYRu5z
UL0XtXWV384k/uRX0xhhO+XOxo55bZx+5+lzGHdGrFhgHETR6qI4Gpmx8geKvnCR
ZqrTqIPjJkHk3mAKgURFOm9VxfnEALAvsCirYD8mXbL6knvieAjiz/mg5/HL7fJn
4viDlfjWG2JA2WpOioWNFOZabu/dy7e5L8k1gGhsJwnK9R2k7PyL7s/QNXWdWGsf
9QzUXacO7Q3T9cPtKrytMfu9kNliY5PNARsM9tRGJyMwf2Cv7KVcKaVbWGquwon/
G3D8V/KjqIBF/Mt9m8Zz98XRSRHzfJy8X0mtvAfwDrYXq+CH+NpFz5uKCctcX/Tr
ydtaqYjGHpdrwk9zstPVVlll9m1KOp2AenHArMjPelQ1vl/pDHF0+xPTFLEC1Whs
H7flqAGiLUuB43lzvuHN+4WBAzoqz6u+hVZx1GO3NosfE6VkKfjlq7Y0/BHj5EoD
AUJxxLL7tXhM87uMTWi7cu/XCaybLKItSZhmPGy+FgGL4KbA47QlH6E13ns7vmqN
YG1bvvs5u6ygq55S5tzNaG0ieAbLRHyStZyys/2dGaqUEHvkXxjJJPWamoRphycv
WignhDMIfOICrEvBLyV8NhGKtU5lBFo05JaF0U0r8xe+RHc4eDJecmhzmFAxmg6e
C4MsOyyLCS3vTwa3KIpqL8OzrAfuN13rimlke7liM7X3lpj4Q/+pwjm5fHBaQoRG
D4qrHnNcxJ8WlK2Q/EFF2bGfzTvA4Mit1W3V9F09/4ZaclMcl4Z7grMpXAYucwzg
aFLAMB526GGIr7g7TG/yEEVd4wpGwUummFYCGnHqibQOezMOYKhCBB4dI9xkTD6j
/npMm9G22snH8xkBTDvTVJ0Eusuu4xtXl1Ronx+70xNYJE2f0TxmgJIHcLWI0yn/
GZm2W5tqmNfiSubg4q83qVFluC4zP9U1W9CEC75YTFHN2I+K3D8+QjilbLx1T/qv
xohGmfqAYwJDnmefG2JDIcjSWgkgFKCDUC2i0zUTOYc+wSQDToW4p+S2+4dgJ1bI
4G+hENRlyxrDQN5/JD/7am6ApOV3DDdNWxHFLLBK1yUkkU/JK+4blPAo9fk/fyLZ
ksEkP2OiUf7OtwIPYzjrf0DEQ93qgvAkWOQsJugtWfhbI0DThOepNVJ6gKPXELhH
IGPeQKb7lM7cyT0IoXC8tKpRcCY1txtaQVDHFpCOoK8n8/s7trZtaJbF1zZUlUex
wGP+fU0Vwc33/N2I4n1VwnykDCP2GwJ8xSV0buj0hR/7eRsslBA2nHbfiHQ3r6ve
Z+3Z/7010s3ztICL5HHPRacwXI/wr0eSYCHx92eB/jlBTZads+CfeZAztZooBN0a
UxbgqGEetUonXqM4lpHDyS6agFm5vjv7Qu8DSNFI9FPSGB7Q1n1iGsHCl0Npv7On
MtTJ6ZgSJqQvVmz5cJSTWk/OEsv4V/UqS5+MXSrnKXkiH42+FAilp11dTsvA8wDa
r3vvxoM2dv5zYJf8u4lWYxfcMXUR+ndmlgyoI/aKezQEAl3Dz0TStJMtc4ND7v5N
bufEjXANZpdZ86Irdx+UqZQ+DQQxyZ8bBlzs4TWGMIU3M5clIufdQ+xsnd5gaC7b
+wlYa8jHMFQVMyaa7fxqayJNROlMdJse2DYjzf21nQ+li/zsjlt0YqvgaR1WSC/V
SvW8Rz0qmSTm92BvsvrC6Gd+RwnpgxSGYMhautFHToWoF5uJKyyVPgWUyqx8zj33
mMb2HqFRD5scTXZOQwZXtvNoKQutGGIqb0PlSD9gRo4ziqrH6yjyJ28ZVcP80WwL
PgEn2kWATSRZBh+owMHrRlE8Xg3mytf2OB6R+ASnbOIIjyy8HFPOSQlkz7MJQn4S
CG5MAGbbOSG+9GVLrnTOi6ZfFdMKOaqDfnOIO50i/L/ARI1Sa8Br1SWpicHeL5aJ
JSsPo84hu98nSkIpXL8PVrGIg0S6fsDTjds5JV1kHkaep2hOoCLn+QzX3UTzct5J
Z4r5JOJezww2hDU8+XzdB9Qpcl5RsdzMrCG0Tp4xJJ/tnwwSMj75XuwdXUzrdv5d
xiEUvnbTyj9NpdZf8v4CY1LV2LyvF9OZ2hutksQJDdUqbjgeZBIvqkZjkhJsZH9B
63EdeV7TvOVJolzoT2I38urif4UV1RWZ8E8hUiD23qB+GfHWiiM0zugf/G6MFKKR
Vqar01hROchV+rhjbgZDZkjIwvXFmZCNPddd4ix+mdQnHK907qB7I03c+MbFGx9Y
Vf/K0fVs3EdwIxh/q6j190I3wuUwppuHou7nfSzjk8lpHoCDu6lx613OjdkFaaQI
NZRnJxhZiRAB0eU5m77Z1OD2rIGMPFgnow3IZkAG1ka1YO+PKK3QREDR4FOi7uoC
+3wCGi7B5Sk6kcUvReoZJaxIXeks+3dgbbFpUjRSwiXknCITpVjuhz3QdDGfkkm/
+gtflp5uw2CVHsKxTWqxhX3p25DIQXakjsRPtlaGI/8/0CPsOJvjdsHVmKl2Lh4E
0NRuD5LvLI0c11pXHn9wVSqSw5ImQ9SLlXOFDwzoMGAX5KgsIzUtWclHgJKrRsYi
qeRndL1zRRVVmaHYJQe1mjJN56ttslmLpPo+Ql978um2EPhisWb25qBsIVspSXTW
gbXVMlQUXbPOCn5i5eh2w0b9ZKRrDgPlfyNGxzFYGSxqkMENGlvRRHG1EoUKfm3d
ToKBqtrSXFPnmQcudnp1KxpvytAAyNEff1wHQBdwNd+xKv9rxJjZdkwTICJywuK2
0uqIAFLZi3jXp0DO45nf+gcN8qUQ5MJsd1UPY4rr4+Gf86ZXKE5KsO0AFZ4sPvzl
TqCfy6i5lbi485KUlM2Em2yUBY4QeqW8x+pLqAKcS/HIRYx6PbzqiP9AQ2p+7zpV
LfrF6TZumAwBfC4aSXchU5CykeU/wP+TgZhlnGNay43kK03m637TfBmOClMUB4nW
sYq5UXQQfJ+VmXPukjil2RSkLbg409xtehbIq1SrBRD86l2FN6L0B4CWGtcl3aDz
Z1YtOkq7F9kgA5+SRclw9mCheohRS5XcN/djxviMWFDxbQK/Su6PyxwuIrZNDA7p
Qcazeqx30WeXR3Z9FT4/TPJmUm1K33T4pLmQ79Hc6dSLYkoU+awaCjvfUv3Tdj53
cBj1TJPtsmiAtwY3k6H9wHcr2uTqBtKb5vt32VLFT+LOyVaGexKpiNQSUYxRSrxL
RCO0UUsyFx6pK8NMulkFTqE6IdrBqiVLEuVNHlzbvfd51W4rXaZ86fucQy77TfCR
AelxRbXRzDJbQ+EMJa5a3umVvCuUse2nfX2nzA74Phgm0z9ZByAqKBSXPsrH4FGl
usnUiT+/Kj16idL9HIZWBDQm9G7Gq4nDhyCMfGqRWDgK8eTXRCw85RfFZxvJFl1v
AJUOV2ZCHjZWg4FP0RguQ7N6Y3aUMmGfIpg+HnDlRjlg2n0tzgn1MvZDZdC8+/yO
jR12QZmRonNl48uFvI1jkm/GK3gnAS+SaHrMJGzU3kHKcy/1g2qdHnxDBlYFHO0X
ggMVUFO8O2qJWNNcdFAFh/mj5lIAQaa8eOdYcg7p1ynoJEzuBgNydGipsddIghlf
DNTr1/MQUx1ar5yQocIsiy58Bw7lG5UQH7nrF9cScw5ZFe9ZH8W6hP62+aH6G1Fz
6TLGvfHwDI9Jm9ur+0IOxP/wpSXgMQ97unob/mzMRd6VkF1HPsS8VRFjJnp5mPmb
/9ZiFEZo1kQ4BbwdvCk7IYuWlZFr8QtZjKr34wRM5Mn/H4zZIU+ZhIF0A4sIlQTh
i4Z23jCwGLZJJZS/6aXAc616Rcg2po1AgW95bCG4z5/3EnvpKPSVyf+ZAAf914Yi
p8TAGsxE8YSRKW9dbXMvqIJ63LXiRe+QfwcgDVSxvdHUmIQbdN33e08ZjoruEvkv
SFhzBWbxGEV1WhJJD5+2BHRrFrFPmJDqCihQRhtoDazxKe5vft3c4zjgBqZBxwG0
D5KRiZyXQfMzenoII2iAnA==
`protect END_PROTECTED
