`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Beie0s45hRj9XSXhNXa75ms5FWza3IcLdxNdJzJSwROKanfTvMuJE+sKwFmfufnI
Wz9fEDYxs3zgOknUjazQNecLwQRBudy9jBOeYKPrQ6siidGDozkixhekj8byUAwi
ND6q5MOjbedNQ28+rluGBIDnH/BvpNBe2D4OSZetrynfCUiQNeWDOR77tqnw7D9a
b5XcfT788MTs/Txq/6GX8bilfxDODOFEbcXuv58KUANLjRaAHdguO6fHJJ8mW5Aa
1B2Uk3T3yu+ADQDTmSdu0+AOA9Cvi+BsuRW6YtyvgonP73BvfFFN9K5oEzy28dMK
D4DbqhrS0Oe4hkPzbHRCCvVej8HclVCO6fusxTQE3hKTYBKSX5BdrnWsmaeWo/e6
SCjEX23DGFLSrAlMCtu8XWqkKgGgSaUzqFlZfSWZLBP3yrUafsyFPPxtRvn4Wkxm
dolr7ZCo0L6dSsMEi0d+WDt9iTZkN8J1X3tWiFO+r9LRL+NImEuT1Au/zR0Rh7BI
MkN2EZKPC29hl+Bv/5f5uZCApV7tvsmqL7NgMnWnfk3/XCVgLcKl9jPxCy9pUUZK
/X22MMbSbp/qBefUMfXOXnYAH/edeo3A3C4wNiYg/SlU0JCpIne214nFd/Xbw6D+
j0x6MNp4IZUlepaaH+Zq98T+pq0ZOGnPrqpttFkle6Lss8LelqXQFEaZ7G2IvQ0Y
nvmwXYHJ3GuYKwcOwflBP/si8ntYS8eYYMOITgGqYbi/ndcGUTS4QmNfGq9705Ad
ZOdN7dwkLsRLMYiWfh45vKgNPfaKghbiqFHvidFWDsI3x5R3q+XVLZZuOemHViz/
AOPDTsv1NtzzFgbYao5EJatK+yJraIYZh0mGdCkUtYclf0I7S41dv+YxR+0bsY0r
kFEexd85uI4j/EkLz2YY4+kewVD3FaYU7lrE747GX4WTsfX/IGCShs3GXunZ/Lrg
+vKHp+9VEb78gZA/JGz+Kkh4lV3GF9ysUprb/WGsE3nEVDMhfracHwNYAwbFE0Jl
jZ7CknG1BnF2Kh0FQMA514XrsAn2LWhvj7pM2MrReX5gG0tUl/4ki6J4E1fpKUyj
68cmchmYWclhUVI7vYFSdCxmmci6SkF1QeurDh0m6UJ++qwrCF51Hdn221neSsR1
VieMhh5vrza7Rwr2D50n6y8MZIpug574In6uRuAa3RpdzJWr/5tM31YetyAzHA9y
9vCA9DlhCvtPW5XMrUkkyYQLtLx0D3s/nm+uDKZ2k2Gh/d+UPZUP5TbMn1kr44fc
MSwINpzj5e/1iyFh8xxaHoyKoxdLGlXvkc6lTYuR+yakML5qFn5sdLIHRIXz+OYa
i3+UfC0CHecdmkCTJPyO57l5qx2hDvRYi/NbrNaWakxxBqixvb7y4elg0i3r8X72
8UB+T5zeokRIKJ4mmkRypGKDlPY2O92cRa0GjgMYIUc4G7l5N/wreyiFkRCjIrux
vygSbCOe8AVvUDX8Iu8+lEwHGu+CA9DHhz1nqXepjGAunTDgALUS+kZytxY7uD9T
l9SU4eZAg4Ac3CRXGXcJq+2Q7bIeSqbSaUXDA2oV10JMGLKbG2zRDOjK3Dr3tfUX
B+ZvPXbeeSkCVjX9g1NsiBpEVo/kXwBKMznArbzwquB4qyYK8MVIX1srjXq20qrC
5e17pWGuqGYI5xUAlxHuLTfE5Ns4Jpwwqg1a+/LyBK+T7AHED1ireHA3b63g5saS
Rfis85beKEJ679OBThkdxGK8XTccvMoM9RoazyZjQWOy9LXZPLBWAhJYSzwmn/3r
iKZ6yADhqH4+ci0Knis4d6numQcME9cVIFNsHLFLzcALgh7zk6hnTm7YelQ1QDAK
JupfIlWRCJWOBKO9yEo3pWAF4TB6FgnUviQaqI+NShtrSmOQsgWAyVS9N45fPQFc
bKVxpqccLuI3NwHCa+DwOebl8gowH6GzXUG6abO3IxpWkOWfiYmalTsx4rKkOL63
peSXHkxofvd8o4XsogfL+iqZmIppgDO1o5E6woTwJqo3+ohiiqcLseCNXpFort3a
NnijyDrF+qSQpVkg5Qzz7nicY4I8x4g1t5qvCxIyt+dR6yO+108ksL9s3nAdBFtk
79MiU49Zy5KKozElDPESM5FDvfASmIFMA/Q92eNpuLsYMozvdz8fbz5X8ckJeP+I
cOHTWaaS0p/4RnPZajAg+/M37H88p2BSN0EUl/+OFSzo+BQycpQk4WRx4uBGitJU
T2wBchEOtQixp7Y8KfDih9GG3KCESbWNV1kO9iXjv+3GEMbTWn7b2ViKLs7Zxw67
T1OkfZ234TMsQug509SDZ0T7CacZjyHC05QaaaL/4AhZUxbdv7ysnKRYZlRHQeOJ
g5Mjjy1DGKzBa1fmbhhL14SkT3Wdwt+1Bq+Ovxkt3gSTdk4eEK+j3Sft5MgRKZHD
95bpEYm6WU3B6rm8q0CQdWLMILBwRCtLz8aJov77aQ56CHuJoM8pe7r4u3GiYqKx
nuutc5BY4fma3U2vKxbWDVXJ/Cdp6PFIEoZp84NRwVLCJGmeadUrVgfPDG9jY8yG
FzZXm4IXZn16DpNq0Z44fIhNHvH7MfSVbA0jADOAbV8g0cOIQA6IgaoLkAF0s2A/
9qKczFOcHDakoBT4JOZU/TaIjInCYG/fT+B5eJxVSijiGjSOrb0PAcZc2AwO8OcO
+ieoIrp1IM+XZzKcrAOo6RmV9YM1UoDa16u+n5zi4kkzSXXXqcY56n6YajogJKOf
ej7sAx8Nkhfflj2ZVQ+QgB2UND97RLdJD6up7E6Yxb6eQhVl5NhF16qJfADfckNf
DzCI8v8NVWDyIdQFol4iuVQhaEBjKSK5SuQqeDfeTEpusFNMeBHar1k2ApRLM1Wf
mgifQ9WURKkbyK0jWtwZ3QtriBSrLee8Tt6YtkqWzg4nHXP4hMhkYUB8/50RGtZu
fmxRNJbxY+eR15LIMusTikZrHXEm0iX+3czExWMb0cwTh+VBL6tnW5s1zfhXKEOU
I3pR+/OJZxIt5UbtsUQFSVnW3WFsrBgDO5WEWLFk9xQGZcoV6v1X86Jz9jod1HFE
zM+7aIiV8Kjt4jSD8cha1JhUgaQvZtSRB2InOkqe7sIeUU+IAa55yy4q5Wwnnehu
0tZ8b2xqp4wupmW0O/ai6VUIUoScVcFWzGTGIgGY7ddM0AXnnrIJs5p7jrWzzCBR
07WiDyyromK6u7Idy7/ezvOGLYWds6u+2hhpy3shVTFiBD4d092b2VGOZ5nMXZRh
nGFh1Fv28WHmMN8ZRNJVHaHCHHTg9teaSXWyDbePGXNkb8lwhGUPMBEsvuJfPruF
pUHHu8I+0zYB7B3hyWNTjJkbHt935jahD/HPfjKLsoRSTVASk/QOSY7OXyQjByWM
4sKV4/q1XyXlloQHTJ3Cr2xhh+jXxt7dJXtYz5qgl0f+gsajXNkuVVYk3XDwTNEo
Y5w5GAQ0w464zNHzSlxOm5fEZBwARx3q6L308hhq+C1Z4LjYeJwmP4WdX8KPr0Oo
m3oDs0WWhtdqam0y4Mk5o1wSiU742rX0Mr6SsJ9NqUioEsq5t5LzaNCXYxYxqYot
LJZKlHhdXh9KqVruq7Y0EoZ/s4FVnkQQYJJY0GRXLRkXTJlENVL6TvIQlN0CEoE1
pQzf4NWDNsU8/Yk1u7vrw9VbVsngiEfqUo2ATaPDxDLdoVKLh+ZfvCXL2i0Ovopt
N7Lir3pgrq7Sip9Tro7RmHBd7YJc2kTPvYiE3TncdUrR6oE/X/J7PU9yCXp1EGUs
AkuGy4fVG/lXD4vR35pLrKE2qKOfkHrG4yqowYni1JdOicpnTHsGsaLiyhyStOYf
TauUeHOQOb/agcsQqeTB1iBOuX8eGlCYOcQCsZpvFs9YTWbw6Ijs1Y0PXbkeWTb3
prY2sIY+k7qyvpHyk5YrY12dal0GW4ZN0M/r6kHHupFKx/le+erJry5L31MW9fYM
jm2JgzPEQoiZQ8c12lEIm0DzQlnvhHD5X/YZBUbCzMUjDdRYtfQK5lhMbA3Is2B6
jJn4JUqIVrJR9tW42qaibTT1w5Q6nbUYjX3KTJXsOsDIXuVxg6bQwL8olUp4DsfU
ApzXuGOjNdgibBxTRQeG5m4mWvtWTYDZ+Vcmoy75Q2OyRJCSR886LD5QlFFAhPZc
0NaVfxRqoU6rwPV4sFHOOpZsJcBY9N6v2SYARcNZ5RKz5IFlUgWwFsNoRMGp7l+v
sBqOiC01do4NH89zez9D4oP3z37h9ehaogxnaK84hkT5cRyAgGsRz3/CcEK9LnB/
xNsUKUE+uzgXmhrEAErXz7bCL3MIRcuZEbzGhumBAZIDN8zcADtQ2oTmhlEHW/Ff
P048PH36h4w/GhZBxh1teRF2EHAeX4c+2IzErd9Zzkl6c3BXleFock4Wqb/CMlH7
1Pt5iLG7vjOhpHMyy1TTtqmQ6nJmbKLwhjephdI3mHWoJwyb+p52HPgmXkDvPvU+
Crbrevv6iVbJ45kBbWJUqn041sj53ytYcDC1KFzd8fBs87erg6wwB2J6C12B5E3Z
KQ7mVxS3sowJm7TUU+L+LkWcXCz9ZxAg0xAWlnLlPVNjvzhxCBzAIG3R/d9ZRMJH
wWaMoa8VkWfCP/r01FSkpdT8TASEOgy6YBiyPxYf2xWBCJ+O2aFK0ubr8ZGojEqY
NcYJho5h1Lq2rrJBJHUhvo6A+u2DnxihRD+vUhmodEGZwcYQ+HH5xtEv2yx0xPAZ
nRJQn1/unxZm3GmTy7kfcI8IwojgRzBBU7I8CERp/o64tI4EYKjdGIFrzxiIXnE3
ofjVgt0iXgTBvV7rF540Lg7fjWUq1+wQKcBzotiagJEBJdgA4WQmDxdvTU6h0K7m
0jFoIfuxO+3ADVMPx8FRX1D7g/ocpzxlCNY8W0ILVu+vx+m08cmz9Brim0aME9eL
zzNf8G+SpqNpfIyvYJ+TcJ70BjtDnEtkFdNzFDKcMrvt5TQ5VTkX/TLgesT/3olB
yx6SU6r/wMe8f+guCi6yIF9R4bDYWGCJYF+m1iqmH16EkLUd2/jMt/qLSSmf9vsS
8YnHrjOcNwuvspMPxb4Nh6cX3/2EiUroXB0Y7aZkfZljA1jA04nK5RNX5ESHfaFb
sd6JW/0itDZO5B+lA55nBXMjMIJFMQUi1fDaDeWJkV9HoH5eNue6TgW1GxFoB75K
nbAeMTh41Y+XV30Dy/M0KikxHS0+5ofgrRqdH8TBSCcDhOmf00KYC948rT8qfOdR
GHDuSdm8DnKCxFf1J8ZHRKz/XQoVNeXfxx7Ps2lX1WSK+ZpropBhBd0UNG8lmXrv
NhfjpLggs/deed6NOUQHRZAw3fKyF37rmkPss3+Ew15Vhhn/c4SzXBYoBiEImPVv
fO+N6tNMK+Y1XIckSebd5jsIkNp8ynkH34IzuDSS9LADhb5t6bCLFLfMkE5B4dMx
1J3eANdaAOnz7O//Mx2X4E65aRwCDrSE6sM99wLuQOELQMTKBml5vH7Y6dZKi9r5
mkHvdAZFd7DrEDMqbXCYvQJ6XKspVxU0FodFyZXOo5I5Iu/BzfHGyWaj0IKvzfxm
XMTmiAXOueTI6ZHOArHIgCwRwMpJ8Dx+vV5C+QJ5oeq4WRUvZhxR2Nw+MUhkmDNZ
Xl+okpcVdRVaGYzjRlY0AozBiFUoNg3hOWekdSu3GrRtQbKcKOSt583se2AqDUrO
hVTFDY6FbZFt2hDLf76vkjjF41w7ZEHsfmcQamJNdcB1MtQf/hulBsVMxizDA8H4
02Quu4jW4m0HmYGIoyYk7iOmMJtHvO4B8Z2TpWEw0Ta+4aAG0cYemeB7ckx8/fpT
SqfQnxP950RqZUAAuiwi3Wqy04EWlUH8jX6JKr8kEu1TeuiLjwQqHReDvYVM3ZXD
0ESZVXDl1xM4qywX54hI1XWs4d+gqoQcrlBQm0X7X15jZ5iZkqi+b9BcoTPB+KEz
/tflUUB5rxGFZF/h10BwcUfnW6ErXN15MsoofAFol0QXmxIrd7mRnkHCJd8Vkmyj
ojbLs8hfllK8R7JRm3BxjqZc6+EfbG6ID933IHf2wISMMkLc/Wfx44Vt/uqBi0b5
E3ATaS9Sgdkqycsmj8Jlzv/Xz+I0EseSo4CwD2N9JGUDuoardcITYbZi0hjg+2xK
ujBBojw1pVkO/qCaSoYQ1NGQ5qKvBQHs+LjPzqqY+Pe+Un5Up8btmO8PsYFWiwBl
5RHhqxCNU78IWkeHrXfeXdrSEjNeO5Q8BVtZW+caD8B/1NzSrWt943hJqqK1D6uR
HrAnXP7ogXEWcfWj7UYTYELyeLVpa5CgCGtd98I4f0oQx4dw6e9vgwvEIp11f72T
64kZGCwynIJRP1dNeCVIaaBj0MDx4EqnAkglomknl2brfVzQskgcpiws/NS5b3GO
7WzMGIK2YaRn0QQBOYx1Qqapq9nshTCS8E+Eh6pyH/V8NkRQZ7/Pi3QU+KWsmEfZ
NGe1yhQtfOdlKsw1zfKFYCbgLAnS0eSxteeeAZs63yWTVCLPmTt/j4kwxw1lhSbf
6EuAlVTOAOaeUOTDjFHGW7R3dKDO0qCJAqqPfbW3yvQXtsd7ZjAJSFgIfMZvvErl
Wxa1snZv8TbEpDUhkuD1p9sUofeWmrSiYd+pzal1A6yghebDT5tleeKwA7dWN7k8
ZjJmo5yY8cdK+YmkNhg9IJmoFqgBHkxUuJzjsRl8WAes4lDugumY4MDQcPEf+JJu
4g3cbgBgOvNv/O00KlGJYtx5XebEq/NwReSAHbjYP/fcVXfgGsCmn0snl7n4h3aM
xe7rd/G08SqLflSDv5g075jWlox8VMwh2xswPSeMTdkhE+eRvUxEVUAGRvtU2mcS
pxUyqzSVfFPoKcKZOOtUeD+Km1OAug7QRSZV+2EL9BAUd1pzH6kEqxQJBYcRhlWP
negjFxW9K1+Pg+4H8xXx5XLpP50HmrtiiuI++zSZthNtUe9zg6i4naQqsOFzSpMD
uZxrevTDbfuHKTY9aYDG9CdkZaMhejGLvxda/Sjg1L5Crp7qeJMkX3rzf198zd5I
/2eyUPncSUWTMH2Ab3pwaqcJBcR4olNVybpIPucIQjXNMP601+utbbjIFBThv7VK
62tG1s0lNua+how6B38EY0fvbh7TbupvZaev91xJ+aimpo/j/ZD/ef4tHc8MS2QW
kSwWNoq0a06+dzo2Gf9H32cbpPWG6SYUS9amb123viFr/D9rT/iMvFKuH+b/nyCg
q+rUBJp6OISmqEmHq4JgPOGaZZjHOSwxOCW6Anx+qlGlljoqz/Cl2Jbef+pHLdjz
3Z5JZvfTLBB9ExTI6/qU9w==
`protect END_PROTECTED
