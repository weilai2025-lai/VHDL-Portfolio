`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2DN4NvgcZf6aet7B4+OyxyRK8RxInKx8IjjCjQr7a2VbOn7hxab79YEi5kMwMGJ
D3O0D1cDaMHN2ujicWJMbf6y3Si6J/eOxQQAxVTHN1+LibaYrIuFG+iEas/K9BlC
EfcntiLYUuCskzG3HJ5GMo4MFwgs64gDWyCBYPt+ovG5hXwIC5pIJ0ZD+tLVJ1LI
3CnCSsSIiuSGEod18ZoPK4oxriTFvDiomI9gsJKGrAiiMaJZVXT0FbujMExBpoI4
qOAUAih5wCrBeMh5WDJQCUQMTWqoidl5eoA/mtmUWon+Y9lf1kYb87jiMKe6HpeG
qQ7LyeahLaGQgeBB38UzJ4Uqia70oOet94BvuDh9HtaISjCc+TzGQIrL0piNQlgs
pJ9FXvkj/HRmPLHyULedzuX24njrdQKrxVqZnBB5UdBBvGArCXUqp3bXMAKwdkdL
73ronPmxf/aHmjVDsOhMr8px+1lUIux/3daCaWpxbFL2oyXDSQF7wu3MSYSKovZt
Do309jyvotwrzQ3iIn9iWmOEDQMuhM4R4DG0ofpUv0JSRCZlzdrxPnOwdyBtEWO7
GBlbym5bAy9A8/3hbgkibgrd+SXoGWkRbsumehkNsIk=
`protect END_PROTECTED
