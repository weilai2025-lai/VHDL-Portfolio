`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l00MDWXfz2PuQkz0vaAjWwotA1XtHr2sH6YDnQUhnzZJQ8eKV8Dqld7MYBXio4uZ
tmEuPrJJDjk6vHi8lH2VM7KNjLnVcGNcYMZdeZXr+UqlNkb4cLgDxypKjDDkCYzb
QcSL2tTvRL/aa4ETwFJP9+qBlUQe14BNt42XdfMIbtDIYrqv1CUIBQK9S8qfDjFO
MadtouP6sKbO8MaPKcogIsob1kgaHFhrl8zsc33CxovN4x2WLaAL6zxKjQVYfubg
JZhnEHBSTCQycDdAna5Fgg6k1h0h9SwYIfYq5pUoG/XZERaQ8BkxVCcJonRYl9Vq
fznvBLNfTfw6Sb2xaJv6xqzlqXOXMDsnEMhYWvyMjXFN/d4fXkkUvuxHZ1MxBIzG
bc4lKGIb9EqDhg7+tijCxDkd+u+9urtORHz5U4Q8wphvxavDaq64xibkKwFwQ8yN
aQ2OYKfYizuA5t45JAppB7Mw8yDfI6m/1JWet5dR/ZrhYf5Dgd6NqJn6M6xW//8q
S6LV0+4fgaT4p8r/VLVcFN0B9c/hUO6TN+3KBNRmndZ1q983yL1V/7Uf2ZU9p7DZ
Inc0X3teWlxzgW3nHEia68nltdxMKWabUtHkq8jL1qHfL6iklUPg2y/Z0nL3gZpc
zt+HZ+fW2COJHeehz4inD6zGuyHvzD36x/Uly0UYbwEMSuRcvVmf6R6krbHunTuU
0Aw5BgQr3751/HDeNt1brNl1ZrZBVHhRg1QSz2QKdb4w9ekxF5uTthT2OW+hz8pd
n73U9x0uVhx3v6HRRMQyp31UYjubtUJ/+w1qPWirsb7suyaq41e3elNkY+XJbEgl
AjpxJhFo4IbK+4f+x1sw02h51tl2c+uB+97hsmuLc+3+qwObC2IOmSU3w9gSMqLx
jCWVqC2sSdp+p+G8n4TSI/w8OVDID3zwK2aPaICB4XuylPsqqn3ZzY3Ds+dlCABz
H/zHwHqjG++0S5DWMEEXxMUgEoINq7b4bgHlzXfOESnjY+XXO8nNqOLMBG+MwGkN
Hmu9vwVMG5ptuVAYGJD+SkPx3Xt/xhZOTESKuHttU3Ka23QYKMBWAeXT2CBnz3ln
h9a8U2Pm+vNCgCMqU0mAbyRO2mGIqkmXffZJ54Msz9CAbhbBAxElsw6OMHO9nL/z
AGAdSfbUPyOJYKOQiKvJaTRHrtSG6XACiDYZBVPvrRc8uwHX6kSAvcxQrU1CLreI
0PJ/RLqPC8dwDY5u734q16jI0IxopbFUzzpxPutHWyUYbx68Rs3uhnH1+iraQk2B
`protect END_PROTECTED
