`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lcmswy8XKaZgGWTGB3iZuIEAbi1Q1QqsLQNxlgjbj1O5XROrZJ+FHjclwPNqjX9
hRdc/E73bEvAWg8XE2vzibscr50ZaPAi3g3puuGHf99NFssNMynxX4VRnV5AZnJV
PBvFZ8xraTG/S2Qol0LjdcVLlSimQyUhH3259v4+TzBeJX2lpKmzaaNcJvoMnVZe
CEbfKxkcXW9cNjh17ELiWh8zQaxp86d0lELI/+YuIDL1gMWgPz+tWoGlY10260gL
6Zju/HlU0LPl3GCWyA7dttqDJdm/3GUH0m24KjHLeYml3+4+IfZRCqJxRgZL72jv
U6wQhWA42nF6mxIzAdONb4tPw+kdMQLDw8QMXXPvj2x13bRLEXaWAXbux91077Fa
vzf2rNzG5+LxNzfelbILYZE7WfHp6Q5lvKISN8Fa7JGKDtwaVmLXg5SetKchHfoO
da1D6EXkPEhXO3MudY8AdQ2sAfFI+esGrH72ghS2i7WSs+Pc2z4nGOngWmhFiahW
wSayJdYh0hZWBXLODfMecrzVNC0gecv9xF5HmDbtWbSjU+pnj0Ma+rjq1BHcQp4Q
v4a6HK8F+VUmn2DGfn3t27BiKQrSvhTP3wQ8bOifYcGA+rKv/MhuxLyD3Q6Z6ZL9
z3glUCtVHAftdXyzSuPmIjJ2rYFnD3zzvvrZrLgLsaXm/t8e7XqpTkoFE1c5NUVA
sdaHDJiO3xeLGPzpMEzMZOdxt223E5a3spe2nO3dVxrPeEsCW2iNCxaVBHzlvqEF
JvdZ3yR0sERxcT5ji9U5oKBYGOD1GcFMY98kh63JRKz7RNXe5cdfa/lziBo+xi0L
vDxYoXeIPPvTRWSJCEoKZhGoMynxzHBLks1JfkZ0JBZVvnDN/pWXqZU9ZiUdWi5A
5EfUZwtcLtuUHKX+C+3uWlmQjRLw3f2EkAzH6i6fr7ZW8gtQRYoBmW3QYDmhiaAc
EHcCuy9XogEA+Sla3C4a4Ln2jvaWB/JSdpQhBCpQ6lPAnnWJuzG9ry2lD4ZJ0Err
eAtgDO75kT8gk67AxD8a5j6a8b+ObQzJjUCbUGVtnVG52It+gu3bBk8si4Rcpxv8
B5zBeCgx4WB3pSp7WSHCTKqHSTDeO7UxgXtO0lvQxu4saqvSsIHm5oszhimpBwuw
p2yoxpxSKKCtm7BSED0/QKeLhej73DoZ3w0LTOuynjH3WMPlbFjP0qDWvathvcrU
s5EnuRQbw7a+fMFCPolC6wK/7mRPg396FzfCfiZ0onXDjIrS5JNKmq/J4+cIu1Lc
XuK5FJUw/8gvxQQE/y3SVwhNIb0cIVV6RBFliRx6cSS2fkTkm9g7Yb+ZGWjbhxuy
nNxi3wdN7/0KdRnotvxAt800+j34HllYNN71nbs/avdxxrE//xEuLZMZ+macxlUU
eB98zl6/Zl89kXkOsocOERW9Hg4GGPzGNFoDPUi4MY71LvPcW+UZj9kXlPhQbWE/
6mNUh91MlBxhrY/3LyorR7EPgw+2CZ5DPFme8pFU+n7pTKALe6XHBFnqOnlrJBih
x7/IVdDZtg/cEKbuab/qzJ1p8NWYRAXBT87FMyDZbEMBMuadHYRIpYv1D7UY8mc0
sFz2q1eUohTDMTtV9VIalKrkLFao1dkMjsXIUocEyMIA30D5OfuH7jgBDIaStPQ9
/3Xout7raDSaCKOFnGTdj3f3/mQJP03zgnLy+nDvBXW7rgtSmqjwv8orcGrDQt2h
vOJwhkMLpJL+KekwOrK0PnyM78rJRDlEh2MlMbumpvGsxqdRif963+mEWeJd9kWO
KQ+MjrDY0QSNiSQYtbBdfjO2cD0JLCBRaHJ38X3HWm34ZS6mnHYt30pcc9Isjib7
cVDoiurOAEresTEWRUt3304jq5Yh5pcJzwHIVQZOkNZVdY2tet65sdEhzY6BYjWy
t1SZ2d058lvbHZXkBtIo8+o7sWkLJ/UKfwD3S49iGNyJz7HSbYn54aoFt69Bki8T
i36OErmBr2O+CmS+3pjsEghdc2LEFyNF55TbEST4mPyKpZEKmNqc4DhOXE2GUCRI
LZe2NzpkHWhx3UmkvLzDRK8Fkrzcthik05Zo0LkTbp00IrXAweReehodyFYBlxmz
5QKtbvT0+sePkkk0pywkMJqHUV8duRcUj61uJzo55o4iVUFMSfzVRZsQGwa3JZ3n
dex9ZWNLJ3xXxaZsZxkRYX4yQHu6oXug7q1XG6UW1HMFgLYxSvqrvGiI9gx223f8
bwFJ4QyulP1SEuh98fs/kJu2XsGiv0WBA0WZ90h1kE7SByBrI2kGlpafZ/j6VAvN
fYwWz28aooRa0eAzL2lCqInRuYjUZeMF9qDKXzqkZXF+rcBE6RJe8XMGneJc/KN6
b8wBFaonu1f8UFX38fWzBlCESJPASryPhNYkp3XwY3kOIKt7iWi1TfBt0335cMMM
vPEXXnkeOnNqIvRc8jMpm0Qu/p0zEl6Tsy4OORNfDSMaUfA0PmgQe98+xZYDD20R
BE6b6mMOMpj6gF8oKnobkRNRAbGVMZRjTUs3MIQDumDg13jgbRGoMYTGw1UbwepP
po6kC6ir2+1HbfbqBvliDWKb0YCkz2D5n7m2hobyiFFuW1Ng+Nbqn+6ZAXXm4fJ/
jxcLB0Q5nXweiGthEAscvluSCLsP+IQysx6uTzY67X14FoZ/cmCsgW3gdyYVBQit
3Yxh+4bB8rc6LbIpSDCW/ybzd2+Tbj3qTE/8KTDEHsYLjmQu5uQ/FKa6/f3kTatQ
dnBJ59aOjeRpLVPUxy9Y+tuZN3l3FZ5IOqFDI/AGU1qMhujvdZLUzLbHGcMx0eff
+SxD8t73rmMlCAJWn11xUQmi4bhxAsFUAblz9DxfndxT8diIWxL5r/qJB2z1sE4+
vwvgqbasm5bZj/JU34xYmPPj3XqlJvgLbR/Wj0JknDSDvAzh4wNfMChonm3GcgK3
qVe12bRp1ZA6dOsBe/CMy2ppq3swKPOkjHVBGpEYapQJZOTGzhnHbezCGOA7ypkn
dt/fWxRejGuuloWjvjGBaFXM+JLrAAMQHQj4l7DE/ALOO03hp75ESyIMbAt1kHlL
mKMU8UrSX/uN71kSH4NAYT7os7MS0JjQD0pzqdZEY55AjOvvL+hPIISMLygmXtAZ
jUh9OGbU2pFwSLKx2iPbMVxqOV0T970yicOHyah9cJ19D4ifqR8iNbDJOL+76ql8
Gu3+UZRNTkCRzVngE5GBGsYnhBGa9lp7jlbG99zLxKefLQJb9GoaAU4wqcMitYLI
9fwKIpldpuzuoqZpO8WqxNyKzuQC0Ez0iy8yopyqvnhaMjGcVl/t5Y81m0RrS3gg
3F15Pjfa5k1gnGRc1qBUMr8CLm/yon6JB2ALv/NX/gj0HhrPiu2ax/fsiT/F5RvV
dQNH7iAnKw7Q3I9S8rO+zbLfWGXBV9eW0NlxYRzuOHFvcjwL+8VVXlnRxxHT0sc/
5dY0c2Oi3VhLJXTH7HoFFcLNud5xnFV95dOGPAidCiqEAaR2SfFuni/9oigrxsil
KjHUJ2T8RPF0c9bJ8KHH+z7gX2ljrI7c+xI0ddTNYPUp4nIQA7rnsEr/6uKc+TfJ
4lHzLBQq4ocd2o0ViWQ1I69s9FhBIE4dc/Hs0ndCUbGWsr5dmajyMub6jymdn+ut
M1P/xA70Duwb3lYh2rGf34l8H8Oqw3N5dHTPJu+Sqq52d7Eu3v2VVo/IQJXbMjXh
1Lxk4RicigWKzJHdJohpe/uQX6LFxsj14y8Qd2DjOwAqMW4iuu1CwmXvw4jkXNWQ
SoRzJo7e/G4a4yDzr/hrY362xF+7xK6Pru0rHFg1zWj04rmMv9FLYdwk/XHh+Q1G
mHetmPWq0FThZZGwTmNJc65M1gJu756kzNpFOW9FRJArEYBhV2VesTfrXO/OKKoW
4w9Hv7FelchkoKKrHH+p86BbeDwa26FFq0PkXvDt8opjUTj6gVHLz9ElA+54ITsW
ynDrxVUikRsy35unHXu0LKkqb0XBf96T5bYsxwbA2qJpGxe+wjbo8cCKAzI1NbBn
8qqGQVPdhIJ2uUVgo7NMeZ3TCwE1S1oTAT/pIx1zVaM4nJvDCSXSrdcQjh5LEyec
rHKXcdhkAkbIcl35FMeVaaN45MTSgUNl7F16btyVglfYG2cAfvklLjlBUBj2/fAB
xglQKqkeLLVYH9lL4QsCYcGE4uP9AwQcymZHWvOFWfysauYqHL7oJS7p99Ht7sI2
tb1nSr5sxK2SFYwjNsRfCOtUo/o7rYq/FnX226u1jcdOFIjIxjeXM3Tpkmc+kMyH
ysO8VeRy8rp22Tfr4gKx1EZlIcFk5iBhHVwC9LDwIfUmiA3dEbE9ZYr2I5Kjsn8U
f0Q31att3jnk/Mob6pzej/XCCSKMPEoEjqB3+jCLK0w=
`protect END_PROTECTED
