`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSruORE+sGiyjoxE600igo2G9cCnvqnGm+F01V5YzmnvR8QFDBwjGGoX0iB3knQu
gXn1CJ3jeYQxo030Bd5/3JpKdY0kmyqXZ+jpj0RTtfq3RVSUhA9Uq7yy/c7tUmXa
vrO/CNyckwfj8JHR2/EHs3PMAOtEpEkrhzatl+iCeJ4XAsg/THPW1+3N5G/QdpXE
u8w2IEPuq8giAm8pcPc+J0D/apdILUuQ0Yvn04drO9sjco7h8aVqvBoWvv4/wMia
N1SvHFf5BxYUIOAwecatZGt13bZPGo7luJCC101lo5lWcWAaUYiHWqR6LknbzLzD
KB4vTQbewENY8AM0cBVCYORPW73zTLsAF5+8bOTjT615NMOeruo7uHto29F6Ppc+
8UnB313mNyuIDp0u1z3sCy82LLfVj/ZxOivpojthi1yXz5PaHJqBBxr40JMlcGj5
Srkm5YHqTmE7PCSWkPXCaYmFfVoZ8hRQJ2ZtNIYtd7t9+BdNXBUIMTKzCa6Flg0y
VTKVp+RwYNVMDm+AM2AUAeTUU77wg7ese+nVH1mqCL/mSRUx8TRwa4U1xRz3VJ3J
HNC2Oj1F1S32qMsj2jG3gOcH9ToP6N8W6/wskH1dYkzIVwN2z8qiyRRVFDBVqAHD
rZwGV6F89Z36LtzkJsWW7Nl8t91S15NwdbaDtK619v1gT4D5E1jp+1waKizuJ6IJ
hTcAFO5g8azru2ezQKQrzXNGuFd+Nk04/IbAITPbX47z+uMg4del8ej8llSQcnLo
g8eiKWOUIZH3N8fUvidb+N9sgMH0BzMU6xGEGipXqnUEXaYdAV711KLD4qbUOiRO
QobqxI1w+M3H7mGXwpBkmRl6C61hLvqcx+XAp0TM1l3Vzhmzw/PUy2QVfEbO+CPo
RPm5gPKMSd+kMIZCnNYWq81VtABI3DFg8Ro58xKL27eykx709q6uWGsoe1vD7WYk
Br+zVC8O4xitDj2ss3JviBC5kqyy5S9qMdhuI9oENZKg5rspt12qzZzgvAy2NiPB
qCSMwif3hrof3c/0OLa4HSIo5+01Lp0H1vkh0xb6Riy/nwGB6YH5RZIqvnqzJt4u
XTk3d1xCrt0ykyg12wsLzJ0DY8LDqJCgIyZuOSBLioCVk1ZmEAzqTo4m/MYoaoiO
E2Ep6Vu0Y00bnpfoaf9cjJEaZJc70pu+te5PouZ3ZphNItK6XCuf6a11zBbPt92x
bvJP92hMoSrPdJVouqXmuQYJSdEdAHzrzVRrxFjHTUugoaZohjV64fTHTmQ2gl/5
ihcVCtj3P5gUqun3mb62CQOUu9ERPLeBRUPqBo66G8SjcKsTOYeTvFmQlxRgiw2y
JVcUwL8Cy9pQ+K8KFxSxJaM1saKRMjEiEd4FPeeXzF684wnU9D/ld7+asU8ts1Rt
EXXm5oFvMXDykB9q62/K/6t+AU+nwhmeQ9oYGcPG7cED4oI2Vdhj4zfVDPoMsaDR
nLCHs4xrgdDZPaD2G8N/wwMw9/6jjycj9FNvtFoAZ81cGkqS1k9PZ0TdpH8m05FE
INAoMX0TR2+Ie23nEiUoZgTcicZ0Zdm2Ur1WYqECRMbmSJZd2vdzbS5d8nQCsaA/
KUsamwtvOYDZJwG9esUDIme/q/f5nBtXb55zpZAjR1jegLhy4R8dbiai4HC3oi9l
ME2Tw2MWFv80t9s17c8088y2b8QAYmlP0G2GF9vm94J7PLvYNGUvDMSRcrjg3iXr
Rzza6KA6OpEumYa5JFty3PEevWE5paTIlSdSUpUKXr5PzH8tSTfVTzH41qHFdk1s
Lz/hY1yHaxMrykQM5lTNV14lh10sXYURGywWELt+TUQyumvtw7u4kgbKR4exs2di
IeZqYroPX1SD3Ok8Yo39eS5RFY2UlihwKhIyYjF2kZ9Nijhb19Rf1USEYVEsxMim
qJPYSIBaI5Y2l1vwv50GAF2jp7gKqTJWaGW1O9JfysawCN35bUBN2dyUQrIJ8sGW
X/yahBZ+uareqQR2eFdgGVaB7C57kGrKGrDgbrqAva+6Pcf9LbRzahqHuIoiAgqo
t5AZHsd0UvHbwMpqnDjQbjkxMbkEFCcIcCn79x51fAD6g/+kdsZYXvDZLTSSt961
5Ex2hmOLP2Ny3+cHlhFLPTWFE+dcB0Z32JDnMh9ac904xcT8rYQTzCaxqswfjnsz
l2uXQcIVcZbbzSvJm2dyq7ipTXkJZKAN3G21n3+aqrJKUTAAMlsuSEbxhuHajf+0
WfTHsQktxaRXMc5pVg5gY7qWBwdNDx3JHjQ02zgy2Nb8LK4aZFr1OX3OisMuA1Z7
M4pEdoUGR/iFiTSBKP/KRbG+vdr5MZ0gK2A3YEUnzUXNJNdkfR/7PMdhTYiJKYGu
eqM6Acr43qlv3P7Eqbr0ZsXHZU/KcOyuzeuK0LxET3NiUZ9zjTj9EwdvG723vRiI
XmCXl3YgNC3jtJ2Mo+ZTbzfF6IX60VK0yOGuZuOHfRakEEVryiJwmviJ+qn9vnbH
IWKSFarD6IAVCP//cqdvlYjyWuGHvSYFRPmBOxUiSIAuV0ZFrvb8DRhtfVzfEeks
GzVyDGF/qPk8iqJVO+OZbirITYGiZhHKKflyER6oe9narkMaB/Huhwvis/YxL+rg
Cg38p8/X5YrYuLhYbdxgLghySOJMduRnox9IHS4kxBqL/sBrOrkRyIbrYXTtjmXG
fLB5GKTd9nNp1a85FQFpr6CG/eZezbDdwKhyxdSzuslwHk4qI8spgPP8dWAABbqO
yhHtCylKLxUHHNSFQqiSF9EcKoLf1sdOITXYzV4KuFDTGCJ3br8rA0B6i5i92vCl
uC8DUxH7M4/IYbybC9cGHeA+wbcNedoxPbr+6HE5IeZtdlo8mn/qS1run6tOGoLY
yKj6XKL6UcHu+UmMG/QinFOOF7ZHpvDyyL1XXX3l6Yqud3V0MLxIHkARL9KaBa/7
b2kw+mSUFzF+rwNvPX6B7R2nt23Jsm/tWOXdYUT15zaPpo+r4M6bgdNoMZ69HlQd
zmPGoms/e4aOjR9OKnWON6XMV2lDQJQBYEg1vI9hlI4lVRVraUC/IBSbJpJAdmkM
Ng1MG7Vvtwg4X/8ceUJarj5WgR/GXHab8yneuAWMzwfU6QZ34BXeXOJfDVyhtWeG
Y0kh9L311HLsthX1iRfJK0fc3ScyaHgyu9w7BIfUCmHnOX0Sa+8KPL5qzmeZSmAh
yIO7Q//DEIP9tMEVeaYi/M+Jv0EYQcXVEHAoRUBFYt3t7D38req8xSt3UO49hKj8
0dcx0DuL8aondYXdUCe9hsVWo0R+SkhZgs+Qd4KosYZlC/z9G5EisooqYa1HHuPt
Zfg6gKP3ZEkLBCs9eFWPLGK5Ab9cQJE27LjeMQOKjGsojPzwWdZB6x69Qd7Bx34S
H6PcyjMdAXdj78lOKz7JrWMgwm4DMDvS5C/PyxE7mKREBu/1KwMNaoDH7/teDdmO
91VoVPcGObNRst3wv50IuHkwlIJFMpLxT6P3JImHsj6gnuRnsqfEywchRXr1WLva
Yuj5ZLLkHD14+67PVS9aZhgCXFtwMeqo/Ndemk15Ne8k2G31rsk7YdzR43sVhATz
3ojtEzOAuPLC2h3PfoVjt9yAxzFzRQ7pY1PgWUkDhZLnbdQxTb8FrEGZENUfOBbu
b494+CO1cPpyzfboyoJV+4dHsjzMcqjWgYtJ9UA80zEeaLNBIMoZ3EwWVOuIvLby
pxoBUs/DviomkBQtUnevKoH1qIPi1+Ld64C85/sV5f4mQKy1z2u7uxoYSwYzRpd8
x3nzv3tkRlozYnb/x6S2o17TW5/mZsjDlNeEt6JMEQ8AiB198MWGJ64aqELSA+Ys
JonIg+E3jyEhPUxB/fJflReQYUo5Q3IVK9gzrqW7iRG6MIuewbd9sdmq0Xj8ogXp
Mgpk/G5lNOQaT8aYlIrgaRRAfY6LK/kSS/lfQSZ9Y+UEIo0PGyDp+gG8y495EJ1X
/QauNnHGs3zHvTg6zeYBx+6GbbcqREdqrJNrhG61dHK721xz6erxbiw9ysjW6an+
k3W3yor/BNol1aeqqqG82BVi81oxv0Pg3nFNU5CAv/I=
`protect END_PROTECTED
