`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5FFX5XT2b9Lr60bCFRzaU8mhuNX+qH7htusGq2A04OhvHKAX5AtnaEUs3axujJ6T
2uNk9ieAIDtTZ7+MFjsLRA16mp+eyFwaHJ7e4SCTPWIs4gdC/8Icl7KImt0r7N9M
SMLKjyfUCjBdcoclNpm0YQw7UXjaUAlOcvjpbHP17caC30IIinnep/sXRiVVpP2H
Yrt3YvnUGWMvOcSOQWnoy3z0T5Hofi9x5uDsaAmsw2dt1Xf2+/MFuiANnfY/UJYV
PD8sGHzNMhjeBA2I+X3F4A7rk+nilsN5pnDyDUP2LvW3FuL1U//UUZPdSJoUVqt1
Q3f/bF0kcFxT54vGkHZTxguA327BB27jrt63OK5SZejXALLGY2ujLYiWVHb5NR/w
3ZSy+ZXdKl/QxwIwJLjyB8G3kp6YKxZlPkCIPT22uYo4CastIgIQ736Max1Iwxn3
NUMyTYBdqM9GEGKaob+7FGDO4hr2+A8QBy8lUnr874lkmftqUGeaCL+P+UyX/6sw
t/tVcSDAQtZR0dBv20EXzmk2E8vQAxLtoUScn8pAWh7Nid7kwAcfYYft4hsZWQ6o
c3d9Th+7FEZSUq5I5v6OAEt/ETmSSjuLO2p39YQ3v78DhkvVK9mXn6VGE3XgVT2P
oCmVZTTEcJJ39aqeulY5hXUvkGeeXW1gYJn14NXA5oc5TTQkb4duw18TJuJWDTXt
b9XyHMUjD+/EvOed+V69tdYH1pHu5uQ2pRePvXeJfe0=
`protect END_PROTECTED
