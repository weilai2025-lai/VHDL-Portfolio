`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZmSey6t1hezVpV+p8K++35wL61gH7spcdMs1pWZpzRYd71AujMAPtfx0Y9W6r6DC
6jxjtSs6lcaZBsKIxibvpmlY2wy0Gv71TJ15N73PdP2wrnbcFGFTSJ7YxcwfSTLb
PwF+//D/mvLcGvnDyP8OkgAlqdKG1o8cpAi9g1d4AMJmSoxJKWax4S2Vw3quMZsY
DY0AWg0W0H51tsU0Lu4nYSOsPEYkalIlHKTkA4WOWsFnaYXoNvafTdmiYMn5TSKT
Xm2DBd3DmAXziVhf3gOtTVo+9H26xOUO09esIDRwhfLAX/h55Qww755IXwYz2TzB
8I0mic4zoXQ4j3jCvqMmw/kmjbGafWrXq5CvylmVd0W3oJggjh1JBRRiWMW4/F7V
D2qhZNViPjC+seYdmsR2y9yaKYjYREbTeW0rrbZ476khM8D8PmLlT0jB5y0M5OGC
gXhk+GuNSPJdyxMvzNUhv+BlVAZhGTZYAYJ5pOA4W5d8bTfcxkNla1gXjiyJ/xdF
ZJL+1X4hTpZsZxvmaREcATxL4wPTAJB7hHmNxiNXa/IwrO4SlGqokPFj6kpsUO69
5QlZ8QlGnVA6686SlvFElGKkWIGlIcEU4fkILXIPO5iHblGJReVVwxt/rYKKIpyP
DjLjxWwvTqc8Os5HlAq9WhNzbXfrsHhlVD5VKTdSCSDF1dRTk4FxrAYoYZIQqtFr
7MmpaINzyI4W05dfgHBcr1QugYi9DbQbYo6Mw983aEG6XYcyW2ozgyC/OR1hSiO6
+qBryg+U1KkxL2xctD3QKtPUJ3yK6ZFjy7DwMrIOI9DnwpaXAwdxaEixqtp3Hezn
k/HxAlXxt6kNc6mtjopjD/xAC0r0HXl7QUuuZTBa+jn/5tRm5ES3/NemsqLC/5hD
lZZeQrX9pi/yFRbB9T+2xGHBo7Prz3yjpSqgfOtCo00p1uzSHzUSK3RgPUZdtJxN
ZTdDcA/6tz0qGzogqbE4CmfZc6hPXy8/vRUrAdk9f/4cJoI1HO+vvOEvHOKbl6Se
9qd6liQKEPmoreiSJ0P8AyJkgyC4XGgIhvHuDkPweJazR32Iq63fxzSpDSCm6oTe
Sl4+0abRjVRQiW6CKWvXW1GJFphe9eyIOyDb2JHdUyzbfjGqPdjJkwV3428Y8i1M
0lHYJrLxRyVMclkdMif9cJQXIcLFPs9RO44npUxdgmKuB9NNH7AkqYF7Nz+bAqP0
v3DthPHGmiJXX1UZH/LqpzJA0QTL3Vto9tQTqoNo0U2c52rwr6J6LpmGyvLa4x9w
P/FC3qh8zNyP3AoE3xCKa8t/RJmmqZeRRiHkReMYvhzpZJitDLtKDhEZEPqba6cI
Rp3ezRsp9qd5uKI3ZNZREChOC5GylGam35I1l3i789qvW1Mb8oqSdv+Id5vTtsSq
enAiBulV0bvLlmsLZ/JsgL5DU0f66h3eq3rfeZNspiKV9AO0KPvp0lepr9HCrt5I
990EwxaGKNeIoQFyJfNowaLsgDh10XKBgLMycrCflqqdUPpLGewevqugH7Dja13o
`protect END_PROTECTED
