`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GO9FuprCQZO9XD1oWbmh3kMlm5MB75xqHDZBwRwT5mXSrn0HtMux4eXd+4UNFsgs
gzajpxnp9z/fm/Lr8esFKU0SLuyugSRhz0rI6B4If9Yauer8QKpo4z6hMcR53HEp
ZBJUToRduozL08+TX9mTwjPXQd3/V6qVof6KHcmbd8s0oVVE6IIYew4LhGACwz25
3pBt9r97YwFb+HYwU1i1LyFnQqWlHRGWND8o8teAbow1aj7H0uqU2JMNRk5xtZ+G
Y7jNZzPgwBa5hZP5w4wE26j+xhJrkLz9pEb/rngPHppIphs9/PRB5xuouhpzvXUG
NruzJeEc1VIVciy3rSGBtHLB89vtW3le5VPqpMPitMXlSSOEzxiyTk2d/n8ia6OQ
+Rxj9B2DVeJ35a3u4rVwzHpsmu1tBYBaQlaAxOOTNqY68bzL4AKY9u449DxZFlqk
hOB9hD/6ZBbgS0O5pWLXRxyNBJhARpZDMvW3szsKiDzznByrToUSpoHrtahgNeLo
oJWN/9LSrKIl1sN+86GA+cA2a4PieXKK30FAZgH5BIWQ/fupA10ryVV4kY4hIT2w
mvhN9/dkoeOXY7vH9/vqLVCGrZKGno/CCfd0SsT+sGTNgWhkGHyhQo+BrBZm48RA
iCMb5EdlK3Kex+gNxnDO9QGmMNkdqyxOcr5gdZdDQFWpf1ZJWOxzOeQ90BUJQaYM
hW//TyKIBD1ImOxO+Mwa18FQtG6QrBe235IIIb0XE+I8k6jwC9wgfgFMIyFxOqM5
`protect END_PROTECTED
