`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R36kqFLrM8EZ9YoerJGtsFZLPF/2yXyj+rQi2vNxdzShr9mIEy29wLI6zoWMKnLG
G9GjOQaMTIl0pmMF5xdKeHkFXI6ozbQiLkqAvkGs27p/ZNEjOV+1UShBmHUIhy0x
gW3LyszKs1EQfH4N+sEaaR6zeKDmbuiRe4bm8UQ3w6+1VaKJer+77x9cBSpc2UYs
i3nEOuhwn4h+RBsuEvWUijbz1hqbVRgBcZkVPGtvkU1cupXuZxLP5kcQAF6M1Pql
FB7DnKT6E+rmqO4lHnLAQGEymL7Ccn+/AR/G0WF9yLYWBnOSYpFeiYQuv7+ZId3R
nhchxyK6WOtJuKQ7nWWZWzBk2uxU98XOH7z3QFHHIAHFO/NMBscoUZtGUCI4fZmL
+FXZmUy7uxI4iczy+zDb9UXnJK8Cw69xb8TRTYKzxBvHWwOEKU99jYVhR/+UBlAN
XbkW5wi/ojqdzRFbUjVzBR28dRz4DdLc9edBqf+TFSuUBR5minndApRLK1T3Lfj1
tqO7cm0oAxm1mpb+SUrowNwTiPmG23B2FcpzJBP7Wn8FbGM9CV1q9qy2zLisevNn
LmRGv9653Y2yL9R0hDout3RFjo6RWfi3ROW8uD0nfJTRIHKuhuN523PjuaMw3Ifa
15BjUEZIRF67tq6+A44/tDpEtoRK/chnATiReoHvpQVFp/LZchsvpXpIN89FfYf4
EFjCHclFPuzHXjTAQIXZyVQssqKXV0ijE0qYpJk3g5CQUBsBHyapaFaZx2LmSzxk
hZYAExJY1doOzez30Eini/By22+G/Frtg013fIsp2/E8iNbU5NskpJGfWnnwl12e
jbtGpPJu2NHGeYh6FTYjPA==
`protect END_PROTECTED
