`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXk/rCT8NS+3cEX+qsSdyQjK42fytqOAgawLqHM82RkrY2R3ATL1vh1fWaGV9W1r
96BV0xVH8tkd8ZPLqjXDhgdkvSm8uMGsX8yz+HgIztf8hHPsdHMpKP1CozeNscQS
LYQZp5I5WgMi7FEYkQ/h2hgBrvLG9Ex0LEKwO9Kq9pHUa2G/Mrw6+D/xki2a5se0
EnH9zY4T45Fq8R6fzqkDOB6c7ujH/x6vqQiwmwRt9acsXiOCWpiqFWa/jZrlBbbK
QqsrMPe5R6FsSBvXlltOWxENFzNTNEIc63uV3WVmZrtVrnyhbohQN+XVNxAXoxYv
FRjQ05J9nIHhj50QQAnVF2XvZb+0DUs0PBbJMkeXtrTsXzIyj7ohto1izTJMdHdD
q5vZSyvcN4C0StXXN+lBbY0iWpC2om4RjViy5Q+ZhJpor7+eBEFsjFu/D67yUgOr
v1GFR0YcdlOhYS5otKF5OlRldTRJo+X9Sk7vtJjDg/gHsV010rWOPmH6WNGQbA1n
FuWN70s0b+ijqmwqlkL8FgQtikHBmv8gooLXLIILyg8=
`protect END_PROTECTED
