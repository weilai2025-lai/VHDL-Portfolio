`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vd3LQmPNl0sFLEATnkJGzmGo24WY4WDd8VWSOIw0aIf1hy6a38M0Yv+a9NRKhLEt
N89KjS4CrVu0D5ve3fR3HmDng+E6TKVoEUijBlR1yhH/78pnzlKB+4ZK/ZSKVCUM
M/H4cL/lmDAErs/Lph6s4wmjS3iddsIDiFSpj0twvrEKsS6fFfy6OIgo+BOACurT
6QlbPWV8xjDTRMTvHfkBXsG39vZlAqK4hKmSt8LkmiJAdZzQ1Xu5ZjVqG+4+Gn1a
cY/+WsAbUvzl3aKz07rk6lAZInXmEIZElgiwnmu2Nix1rEgb6HtDsrzKUJvC7ufu
NV+K6wH56rBCRJ2yIgwLfLglsvT2D4zoWsZJChE0b2vViKPhPKjTcsQmaFU/1cxR
TZK3qQQPq3BXLDgZ5e19KsSS9wVkFJi4mqbiXrREvuIK1/6dk2cKv7WXbv5EmJt0
xfHU9tq3ny5jzqqXniS8XC6SLcGNoKGw2vGcUhj+HcYh4RhAqiuIQLgS/kq9anhG
UhGDfwNdKx1N+LEBde0XcZy6n3YaXzigMckXuO7lXjsJ1yJ4QxNGu3HXKEQXLny+
8QLvCXEk3/759E0DhBEXETaUqhlEmqVZ23rT0SXN9P5IM2KHN1LWTdTC7d7RCIPG
NJsnvjtRnpmzb+bggt4jA5OMpGh9ZItq0mYiIgIFjC04dmnVHtPOehe1b0bysJvI
VtN1JrGZ6MU7wtII1IEtjTlDNwU5dppT1+2BiTLyrNw4hbgKz5k84CzwesjxlYkY
IN5SQMKJ9uTHtNzVeUo13WWQ3xr9Sb49neS7/OXNkGnpgp33thDg32ZRWpHEhSSH
i6vQQxYTKd+WGvYrkdzOTJ8HORGNagKt8WSU0HjHBA0C8NnVtgcgrZy7bPgtiTuR
pA733DfBLOoN+IWXhKwU129tehBPAeMA7LnhJhpfiPerM1ZrDbGvUAzrh+I62PZf
E6QLmPGjXYp1v7AX+BF3IsSM/zniMaubRS5LD3u08Fgfi1Bcw2WDLQiByasgDbxM
hBCZBdulS/OQHYzOlLIMQUJPjBQ1OY79omVJCUinA6rD9b+vugW1D8rjtSuuAZ5U
Q5vgOoiIfjAp1fqSiyR9NcOwb2UMpAMevf19bEgPfNwhV8/2quA0al687IhxQsz1
geGUfY+GvC67tXCHkNGPt2r5BJCtqhVMZECccFo/PR8RnzVyz7hnuTnpTaH5+VIi
iHL/OIP9ru+LkNBTCIPDRqTcqUTFgb0dm/vgmG4vuZsyvFXWwLDnruuY7OhneZle
rpZ+k1o5dEhOWYFWEnm8lMRnsmrKpE14tFkCjOWBwXeeO/siETyjhlYQO7IKMSSA
xj6WL0ay42n2AepUzcGVr3A+Z+r+Ze9SU9K3OY1kouAypeQbvg7RX8l61KboO7Qk
NGAws/jIyZP7+/Yrs85KOmrJ5WA9vU/e7RNGscNzb4v+MPWTiDHHYTjt7KD6lmDZ
RpS8nk99iIOkKbZDU2G3DpsoXcD6QtRwO2dGydIWNezoPrPtDx4EodYO/Z7/89tr
PSIw5YIfKHLxxYH6hz38qIr4//e0pPlZGuw8r4RxqDjzDfwfSRlCICXZvCksYkZE
S9bAAaPUagf7zobUx38Mbc+PlSH2pjD+mx2Pu+eMIMN09xU8WeDcWYnCeD3HPxZb
He3au/MEwqact51zfITyPqnqWTNSRfaT3VAOSKUR05g6IYXmQtxPB19TtCP2sZYW
c0cXYOjEr8QE83zmBxQ8RDf0pgOVmg0lBxvUAMS7/NpfYQYWbWPn4239Y0JJbASP
11dl8OjihWFJ8X4Br6IPjooktNwIhYDT2qFNPOt1qt2huUex4gFB4g8zb7RuST/J
tiP0TAECaFSzw28PHOsGPnPgWQ+mnQ4HsdrxRjkpCJaywy2bzUwjEexrsuB9Revq
ikqSKPOuGugGsS15kowR1dtQUmm1jy1T2Dr1wl+sFtB1/ih+Iaa4FOPjp/lgyUxd
ovro5R6x/We//D0bUPPBaf/psLTBfzO9nF3TVdc+VIfqwH6Wke27acp30vaKWTJt
rLLuVanJjEW15MUVb2TAm0rty8wpjyXECUhS9dkrcNE/nIDj4Eb+5Dl+L9l/6qIp
kRiTQjpcn6bHwzAWPlR32YWirXkNgUwn6hHnVax9jFfql7+JOvD4ix+1LZq8JFTz
uQ+L9gF+NNAQ1hf/8cdify+RaPEBSuVkTZsK/KEAf+Ftvt5bXjBQyZ7q4tR+TE/9
DLWdgYyVoXVDknkre+P3x7TskE4miMY/RKPNyzm1MptbqhcoVUkt6pmkJiZVzlaq
E2L0xIlvDrMA18nhjR3v+m17MUHLfS5qX4vh2MS5hOBYqxr46lLaXN2wSEYd0sW5
OExohUAm49egrQ4H0AUDc55LPRFmHJBid/Qffc5fomPTPL2MLhVj7snBtXEJR5WU
dsA0k98ojN+pGV5ajkWI1pbwMX1GSAXC2k+R2fJj24eyl9xcs3DYHb2JvgSSzcL8
N69eFHgvBcJ1dZZW3DIG98fRdO1Uuvkct+z1yKulldyhgmHvTvJ1Us/odqEN7v1n
++MwuGAWlZsfaQut7oPIM9FJwKtgy0ll4kt7Jo/woi3evp66pAR3hAGJCUoQYu9Y
+nHIowajO6Dluv4SkwWnk1KGbBk3WbOSxFKXoFECFtZdT/ifGImzzEx+qSII1W45
dFEMpDzg6nPIQEBGy2mQq5b/6n4ozsqetoyGw6ZaAueb1dqvom/40E+CXvFD10SV
aM0kElnnj/M55s4sC62VKOD7XlTS45RLYTateFFRjqCbxom8tlvBY1434mpXbJKH
7N/4tkwHYtCeYTXMHDQzjSms68qidbaJvy9Wn2X+53iEV+FYANG38MQrwbrYtW5b
kKDx9OPq7FVjOLqqoR68+fiTn3WA40JoIm+Sr8qyAww=
`protect END_PROTECTED
