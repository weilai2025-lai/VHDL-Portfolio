`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fu/9KTlxPZB9fledeFmVszyuE7ySc81mK0Qd5EFEtsah0PmYMIMaL/aNSBMBY9pn
MXbtV69MfVBaeLUrOv35yPnUsILN7BqmPLR+I0m18PQie2FS9aydd3JkGHyeaMcj
j6pjU9dliFkrnsrJIJb7VUo/vz4UAqgh6IYGqYBBLiXgNgbGwBuadwhpvAAyhzf7
1QIKglOR2uThU7b/7Ojw6G6PAYRg0v3GsyZosDaQpRNkNRJRSqwxGy51YLowfk4/
ntcvmzbk8eruFF2ZOLLoggeQuM1FB9MblSs5bQPGr2jW3BvAhw9ti8uydhJcs5b2
fVUJ0LabhBjGqehfqj+M74/MQ0nmEv1LX7gh7umJ2hUo3srg4kXi00yQpDIvJku9
HmPT4PmnfBgAvi83YsOd+fpLkmffCAKoQojjBLzmr/5BHqwnKHtdaohDb7CVHXlS
X2Il1eS0OMcQEM/Mz2N67LThz3++NwYniBbN+9huIEXnvfijYNA4y49ulPfYXs92
rCr63k6WX2/JI0U50KgrUO67eKhxDjEg7J2sOxUr73EcE0oCvLPnPYiX4Uj05m0u
5RCg4Nu2/kdezv3Cz5SwqMaji2mbUVhcLzOk3xoE1QMIOzKfcgAm/xRwF5bA+FHx
fZzYG9pNadJUVDzDkCDiI3qvCRp52lH6z2fbmFJkPCnG+ltlMz0bZLauexjh0OrB
jjBEI4y8GVGC+AEPMvIb2ILGga3+FcXTipmy4HYVKnU2KF6gEvkGnvQxH+e1RJLx
9TdSO9UaaqOvn7vZDsgZY3gkN7uIyLzI8v/sVgiOyGoG6TEoTgKF8/qxFZyFjDtW
/ZUFZEVsTJVeOGp+IuqEwVQ58RMSOI4dIMT931lj6VOrq4mJfHCylJqg5tK57GI+
CR0qjN7ySevOy7slzSn7AMO2t7bWyNE/aC5ax22egGRM5IHJypAklwRtCx7U0sXs
ZcXZ0Zv4fFtC3pBZTe9NnDr9EhmPDZB4GC+Gqz5qMIli2IDlWuc89z9/fyuLnqtz
yTBvuqQszX5RF9F9csmtjKmWqSLRuyrV2w2ArrEjM6VIQk7rcwDUlpPgfBkOzt6h
IMOqBVkRfh8aqb1Yjf2AXPB8PEO+6sci2nKTqJ20TLXg6+CsEXjwm9MzOsWqNFER
rxZeaHM8WRRv4om18dix/5beZrX7s9VSlYR5TbJlvg15P8ytcCpYe0LYPsHvPrgn
5eRXaQcTXae8Cwdan3KMUinPvgVUiFZqnti2Ta8fxDHIx0cDgZmRWDcKwdc2ba+2
BkveOFhvEB52v6rfs6F6L5galmZAbVANECtIxHod0ulEkb79pDl0Gp25nKRkv+e0
s368Qpo8TJlLZ9YzeWHM+yFsUq/9d1bk2pzLV+BE+kSNkjRi1IOG/U+uUcPDsxXK
TdVfxwMti+NLGJikXG6Pr9PfheqzEetcZbTlRGQIaYwhoOM2dq8BF56dFZDXKjDB
hJEU9Dqlq9OEHIvtO+zkdAOhFJLE5bDnCFpXdw5PxEsnl4IL13VJ0wwjXvJPecfJ
/pGbLq+ngBVt5sN69EDQ0zK7BvcpTS/jP22UK8mrfNAb6nrMwFMtx/aymis3efFs
BPwwOWbjdfD6IXWyhmYHRehxS6EKWSA69CqIHGcxOsI=
`protect END_PROTECTED
