`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JEvANeW3wxtXAApQG3+6Yksi7/tAP5ePIbMHywu/rwsNve2vPOo76gPi1Qm8sOb0
DmbibGH1JF9jAadFG8+nNuY7PeeExaOfo0+XV19qSpcps22TaOEu0JigIXo/bPOZ
mqvVzU+vT0RMk/qW4hz9bInGNYgXB2ff9XbLV7HnYRZ7P/krWpjYh8mf4+RmTTdp
glmCQcg5MhtNwSNKBykkSdM2/+doc1msBOW6dlu2oxO4VmPUJVzylDXo7piip2B7
fG7fL1AFtYV043LvmkhrtsXssrh7WjE2MTHR+DXwvd1BaBesy/xddvzSBEIxk2y/
H1IcJAqK9iQNE2nt5yA+ulS9/G+c3WdP1GSaNIsQSv+0pBoagA6FwBeaLSrJhzN4
VdVpugpmFl/YI/l2qthJ7t9g0eRYU7PFPZy2wu5dCvy1cYk9T+LrMuHM0Z+G9mZU
E/7LR8gKor4kjr6iti5d12t5BNLntNhUDiSaUW2IOep7ZA6JpC06OXywuvvmFPM7
sNn27kPVWplX7ChrQx8WLl/lH8OyHPofnL3gPIAINyP/YQ0zS6eg5RLu/SaKM+dP
1tSQtuvHkZfr4FELjkOobArdtCfDCkRtSbkwufbTTxFAUk/KWdlpREQhP0s1UTTi
4raoiFxbTOyT0O96ZIAdzE8db4bvb5q8epqdvGr664pHpNT9mTqqkz9YmMaJ5Jbz
Hp2eWlGtB243Whn9szWR27/Nms4ANAOIdWc5Ljox5Jq9gx6GhPBXNs2B6epYEKmf
CmXXzlUcFwjpEOo6rznzq431lihgCvNvPliZJrujm+yva5BtCWWgUs0nE5Lur0hF
VPiv9URY7KfauMAYKbq+8XRHWC65XtZQaH8s60ESkU3qjXK+zsoKmVqBFF9joA79
EorW7WDpYNosuxycmFMdn4pBGODuqf/Bq30uHpLb9tdc+An6ax/JaHmT4MLRCb73
pufBKOIpB8Gk9MvnKcOk/xsHIqQJJB83piIIUKj+M5JhUBogsa0F+V5XL2WNzsLf
patzq7aCO5n9sC04zXU/Xok3NVyA0YXzEKwVHGyPvY2Pw0c+nTeMBOeRHIki52TX
gCPkVn0SMNWSWA85kzQbwa1dSTlBUrmMOuGKmuM3RKIh5oavoR3tZF6nd9ooZ/cb
uscOASSeB40tqTCtqQGTtKN0dkNjldBUEMieG8pIIz6OzUDDMVGQZCe+XOGLG3tT
6EycZnCjKI5MPlOBZYpstNs9USc3JzzZuBrc/Q/7dtlsc0Q7vw9Ko7HtkwsyncIX
73BEjh5FR918zJ7HOzcFQphNl5QRv+MaovXG0vvmFJNxun2U+RWG3KnVE1ibbSpz
kOOqdwnKcaBby4M2U/byiSc9dOsZvg/Y2r1XeHuONseX/hNbPPU0NcAB0iJSvPvh
4NRP4W1rvcsEQZngHmfv5HFDXLCp0s6n2T/9c3HUcUYvQjIMaeUakOAVGyWOSSWQ
6J2nOXW5otaQLpGb6p1ijDxrieh4MHyTBR0uRtdhJmjOU5y1IwLEwqFvZQZ2LDFB
t/gsDz/joRPGFXERGVcYNk4rbompCMaano39zMnPv8VfsrUWQ4V8HgzZtXys8bHW
/+nwf9ax6zfhI7xsZMqphC+xDJEGcFuR5fGy/oyQrZ9a037HJryvdCHpYTdQ5Pkk
jnH8uDpxIkaMLVUb520Fpib6NNIvlH1pTeah8Yh3/PlT5sT/N0wGS35G8dVfBxJG
esS65JTFJhMKpM7I/C3XPQ==
`protect END_PROTECTED
