`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/z7aHUKqf+HERy2m46ErijNeb0AqQW6KureMZhUaIJeA7TQfK8GkE62ej8jPAqGR
5ju0k1zOUJxE5IGH9rmekv73Gd1Q6HzslLKTYwj3wOf74fBEQKsFJznQZmcDBz3O
1dk9cd7Ay+sxc0jaKP43DXs4Yuoa+Kl0smUu/A8poLsFkWxUCWVkH7UXZAQrZ2Mj
ubUZNoUv0H2kjwymthc4Ha3QZR7VLnTJ9j25Iy2lpiOnDAP5NU1Yo1JeQnPX/Inp
+mE91xoHDSHFwWGAtdX1u3w/+p12Z7ecxi48WBdVy9T00md65nzACJFa2rOLGJ4c
KNcbLeuS0pgiWcVhBZpxa1rIDEfW5ix+4rhK1e9/4482D8+SBwspBBpANdzlnso/
51OA1u7Qf+FSUEjMmlZz8mqrNWFj94svDICs0P+fXBtqT/BcXh490q5G+lkPPXaP
ckjGkf7KeCyzHZUH+FsYGRwHzpY1WBz3EdUJHZRyUL526dKlgdO34sEqMZhpkd/f
IWeBzb+47P5WiZwTEb4JJnOOgqKRRWhK4b8WBmusmTimUoPkQQdBPe45ze8/i+Rp
uVa44BFsvY31agZu3uGsVeepn0y7QDcPnWxIQfsCVclgWH0q1e+oA84810oU7T5X
wWjswjhfWu9Ep4nY/cAS2M4QdqoSv6W2naopxxqtavPREAoAxB9qGPGhKq1nlfRl
+3fNHPEutbUiOywuhgppaeVOp7mRpCg3xDsM6WrF6Eq0YPLKeKWENwWPVdjj7KCd
H/FzUnZsNTityjBGBAj53dnZyhQWu8S3wpgJ0dZdY2PP+8M7vMUeDYRNGKAf67QG
LZ9NJqZnFVZFwQbDlntegIDPnV6se5hqBbs4HHsV1pi/8DjBkvFOZXEBU3e0lp7a
5FhBO/NduBM+Skdnd+tqFwjOXWOujIXJhh93HO24VbJGqWwhZmjIMnzzoYIjT6ib
TJMqve8WJN3IdI4Yt9OmN2bvS3pajM+AgJhqtUi2b9PXZkiCpjmUsu2fPqBC2e7X
i7VM3mAjy9LpVf4lxq/YaFOt5mx+xWgMqaX17Cse/hpiZEatHExvHXbz6SofGkCu
9LuDpoXMu3mvyNg8rZGhIpInfGiPr12tz658NvVJEaaJoPVHWO11ur1krXRf6m0Z
AsVcZ9NleqyFxo9YRJCyGlwI2irzTc8weAH6QkSGNDloeWf1dL+js4MjGUagN0NU
eHdOF7tJO3HNzeo4+UJHk1buGwyOmAgccV2L9KEE3cEP8pZIe+ErWCawfMidTKkr
A0+es/lArIZnajNN6fpdVY7i6Ddo9sgIWANFpIZFXpIg+pytSHKWGhA38r0ouhHP
ZbF5LBrvuxFLvKsljHhX9G/ObB63N3oeyxnxzwfqqRJZlF+M8B4A8INBdt+IkvTs
Qjl38tSc6zyRehRkOy/SHIkE5z5GeFVI3zSNVClcK9k=
`protect END_PROTECTED
