`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFjHYNzdWZhsIDvUXuWLYNvrdz6nqHlFbMMn7h8fRhtooPQAE4D6o1q/X0PI6noY
fNaPz4qXrMEyjfoU6xxwcCJ31Qi4cWByFiJgwCO2nISQMaXP/IjgCGCUqjFNBOB6
/3BfWZOFbcfJprlMoL5a/UmVe8uyzeyozTcPaYfLH2C6/p+XVmZSBAbeUzVioP8k
rtXuDoQJNpPfBJ6Zz1ZhI9wiYMc9psseOrNAcUE6wmy20sciHbOjmmUVIB7Pn6bb
3KuWGzAYkzkSFbhpZj9Su6nRecmg25Z89XTn0oKMAlinCnjzkFp3EON/j8SttNdL
wkh5o6PoG0HBOAGcVF8EuNMD9aesNHz9WiG2z3rodtRKIER5kREA7LYpleFsqzgM
Rc5KTtVGCndSq8PJ42JXE94UtvapUL/wT5iYZv0gasEpU1+vLdAipx49dM1YXwIw
PDq5grLHESAul360j5grgUCdRFr8G8NaJ6cFIuVKUrRRj1VVxVHXpKliQIAG+ncc
QrD1wrXmsa9LPy6759G5PloWiXc7wQdq+iSxmgEozPY7LxYet7ant7kHJ/0Xelgy
JmKkwaq4CRnjmvmz0KOlouQPwRa9Vm2o9WFtptxIhLEqx86i6v1NnuSp1jUIqGqe
LFATPEHBuq2KUcJ4TbbZUA+mPOWLqYK8Ozw/XyJ+fmAA8xesSHZTmZwGEBoo1s/p
wx/cIjfQQU91+Bqa0lUBmLKajW+nkga5x7i1leumBVR+bHhggQNthClnx+LiRUtp
TP1CDLiRp4rGKKZuc6bW/MMajEeXorGlKs0zHx1A7Sval/mSt22VZIOGiAHL18HK
QyKmgYVf+iZsy8H5prAZPapp1veYaxn/DU6r7RCNEGMLELERmrFGAVZ91Sa195jP
NUMrzpqgOeSJvWNo3D4/9W+Ov14yA9FZy44BwS1CLTVwS0kqIBwp8mBVDJWjlDlw
cBX/INoboDlZP2MwYTtPimO9ZPpbBD9fMncGHtdl0heJzMBZUUT3XyMX9kpoU8YP
Utm/bjEFz2jEOzcNmTjVD40C7mA4uGL59hXenRmk1CG+hU1WKvWh0sqr6TIyTmO+
+A+QxUT2kt/bvPLD+ER+96p8RkJzEk7whs5CU/P06GlLNkRMhuVRLPqmvzyVeMM/
lKoFhZlyZZXBqEkpBKqvqNj1Vq1LunTImMSTcvZv41rAvGzY4g08yIwU+0HkBTm8
Le7RrRaSQyXDmMLt4aS9ZQE7B48yR1kxSCSsJxahmq7rbAoniE6Yd4oszABIUyBe
h2pfRzs+3iNm8sptppgaYSg4p5jvrWGqBhJms62YdV5p9C9hf5Tb5elMl8ITKoEq
sHUMgsVKPHrcQmy+6s8E2SNAU+WsOAX0OEGWHdBWDcLolQpYJl9w+p31KItTGGyi
uiT8sv3Lpxdq81+IpRY1yDoql8ACyNYBh1bA7/dcaMJbsBGu7tkhrFBfPBfx+W5T
HozNNGJijJ+1ri1w5cG7eC6uP61M50EqosqXtefVm7tXTdtGOUibXBhtIL3ZaaU3
ovupKnyuMBqnPrAE84RHm5Z2BUOXmIYZ9gDAmCc+6cdAKbpxlP/kAG6iGtoD3Nxu
gNaomfuQNB3rwgPSPLgfgcYkF8agOK3mLko17xya2DGx0YtR+Yx/GKxsL46TtwR2
h4ODr3BW+I8/y0LU5CahzEQZqPw0yTT6EY2xGlw8zLOcsYK9IPH/C9CO5SLMA1kc
RLLGhxM1tykdXn1/ISJ/VPtONifwetelDdp3Su4vjYWqjQ5/8mc5sF7szEfRMnqJ
7xzkT8rVMinoVkWY9THlyBYlmrgKtpwwYcaDSUkgHhSktxJ2WJAbpr49+XAXlOmw
HxxtT9R7XsikuHbYmrWdKS0G+guP/o3h6R7V8jd26ok04sW/B3mDSlNXXSUEDTED
FlPPqW90NE5hYI32ywj1P9CfmsWrL3Sj7C4Jpw5MI6gFkVfYNWIHWtuY/tDlzjrI
QeOpKby1HYlaZv5QOJS209RDZ4tn0R7rF1Rhth/JVlHZJOX+uruaqMPwLNbmjXmv
2QblpzAfV/ilVqFYLsP8ZcQDQ2pjpJg1+tCG1yXDZ1zEmMZttB5xC62qLQOPQ1sL
F92L+ihMK1qgcMyNjspD9B5qx94MvAtQwEmsDmOboicbk9ho2nHZVuXQrF/04Ixw
ooaHXLSZYCHexypZLlOtkc9lT4H56Wq0opnyWO6a0xD1dfOCOp+Wb/hMhFJDIZ4U
WEcv97gFexosZXt6hRPptJr9WP5flVmBBb2wqzsXQDLFfgehnitwUPsjwrr5NCUM
ikcMX47jjY//hTCyeFx8Ya8hrB9AmnIlEmkOG+d1OkgJ44s6ufpzGGDCO5WJwES9
EIaM57US+hdF0EkbFiNbCg==
`protect END_PROTECTED
