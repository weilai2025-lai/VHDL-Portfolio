`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fo5Wu2mdIMFwTdHp9iayAH1/ZnxGEx9Zku7KFm+SibF586zeV/5Ti+Niev8VJsS
YyBCt5f2PN0+t+OZQtO10eDJGSiPRh2B2hHfPiag72g50XdZl1GIq9tyympzL0UO
yYJStvGT3ERcNfIBR632gfHerVsu6MR7YewrgHdnCIXmmJG5mktDNffjcwI3JkzO
XcrZcQwcHEHGxTGNS2Eo0Eebb+CkLcjh4X45zs2Koqz85R9KhOQ1/7P60YzTYrTk
GDxZgZcyxvp+T8voyi8afBNscjKIpcpRlrVFV8d9yj9e0lTdKTeYyYSYDhboryXf
npkyVvEVaJ3k1SCZh/+v/xUltM/BTGDpH4MuV/yW8/O/N6hH9rRwGYYDQnUc2AJe
iUm2+oNixzsUzvpbujYm6ggFHkpcv1N5/xiPETghpbh+h1AtydwxBthHbldMUPXG
HjXib6TDe77b/BDI1HiqlqlLMVzHcijt0amIbKaylPiSCMsgqfSjzF8mr3V7Yk4b
JMj7BKdb0WPjxpjKwGlI4Q1rhozu6f/gj1YEEk/gte5GUmrEKA8w9RKBebJZFnAS
QDALMLk3JBCQe5f0w5mA2s97vFjrdFNBeHJNpFuv1CrWqc0ZQqz+HmxqEMvAcS+v
QLEgyFlHCnGuJTK8TZW3qRvD2d2/CQz4r8Ki6vFJu5VJLSzNdeBdZOG4I3BBYwuO
TSPgpxlcLR5+UM4AZwtyhMxXXl+9eOrl2Zhu9a4JKTuD3/YULw+dFwYo94KXDxIf
1EJj2T6nPI7dgkeWZKvv2RegILzqUr0oMJk4/I1LPdOqKx7tBuvD5M9Dw94BGzEm
fnSJnmeUp5L0Kj5EG82YlXIUurXWigmqxKQ+digjLTYu13huyW2RfdluXc9npNVQ
LxZJujq4hoNhOSkddqZ5z9FUQcZOhjoYwM94BBlfgGSClK8S+jJAZ3n1/dYUuuyP
0d+m/FZiYJEt1S30h8q1Dsk1FMkZOY+l3nQvx8UnLGYu815kouYoZXXVsi9xqdtj
FsmjaSLs0SULbfFbjZOFA7Aev9U0HwU2/QBXB7ChcEvdzGHGU6zOon8h09EfPqcD
/TGXFteo7oasNFo9q00DA/EavDZidIYJFlK9rhUphfh7zalE647o/sR3xdKx06w0
bEmCyj45SEa1HGnhTsZDIPfzebwEA0vc7F7y9xcXVBM0/+K6bsXS3wgzJyn/ttIz
dWDDmKxgxAi0ZF22E4oziVWUvbHA7UxuBDT+Jsjuajm8YXnaHYpd4IGa5UGnxAhG
oDucq4rvyUgDdAxXNF9E02pYFPEXuzFsHcgZRF3AJH7zrTqT8jXJ+K5fd94ynrdF
+2MCMfqYR9qVuVRNz+w9zj1ga6l/jXA1xlhLeVO/fP06KMPDhYp6xqkS/vCDc6+h
OSbnO4aAwmcomiPQZeB/IKrLMvdObPGD7ENMdxz69A9bKIgQ5NtDiV1E260jMyoQ
DuJW4Epe4yk52re+dHMtIqFLh3U4NGQWReF5Vibx858ijaTCN+u0J699tSCdJi68
k9FG59dmMffvNnCJa2TFbNZrgTMwYuxqSZW1hbfcPZsNVN/77miEyGtRz5TGG1H8
tjXAnkVmp2c+/kewFaD2AEn/5KL1v2czL5HNDWgEhfWyRCFR7WDNkq9fmEDB5/ba
0jYeqdUqJ5XQFnVypzPKKOjXbRe2v4W4jjm273HY4W0fDKXVKOscmIv35O80Cwqq
tRMdxoWbEjktnQ0yurfP5M/Yv2H0jO+M8/OtpM3ccIMaokfYj7W8HB/pN/hNMrQC
9mf6y0QfBFtcNV7jUgO5NbLLm3WDxZpzidnS3oMwyt8K4+x+HiDQtoH7FR1guGCg
w7vqelFVlaSEbpW/lmG4IPylwM3PRcmCZSB81ViC9hkUizR5YcNNuNnI+WXM0YJY
lhiTshQbWajnXn2rEHcAJIhL5NpFVM/Jd5R0X1plnjdI12tOLcBLARAy189MNafs
sj6OMSwCaZY9rEgj4cnkopYgW5aojcXYT3QWu6p41rnDl7xHHZ+quuuSlPKjgQgo
+CVql8uhAAUWPYX5O6sqsVW+W1hezrj+fjZB7pH3nvYDKmlnWxAAPeNls2E3ff8Y
9u/GNEpeHqSbXq4TQT172DikEBpOAuyj7e9oj1ptKDB9LpxppMdCXVG9Bilr461d
XPIMTmNhaNb34tJwCUBV5BYcA+xX+PRaVmyybL/uV+J3tIdImi5S71VJu6YtsXSt
YKCQIc+Dt7OQaJnfpXFb9ONj0kjrsL/GAsG12tIUB0RsIgSOua/kprz+LYgOsZ5e
xgUHOU5aDOKVAxEa2NWiMl/mB5X8Qhk0oKndGuOAJMQULttzHEFMdqhTeggeP6Js
8eCdDx0affFTfeG8z+o0v2/Pda0MqGlXIz3gbNTZ5H3fzjlb5q0jyfQF+HHNo1xH
vR3XXetXgn6FSh6pXfBM1fGdRHOR68UIgobu/ZPAquOy011s3F62gNToPEdm/7Xl
fV7kF1RNIJyXgSeofG8cy1SVjMC+P8/6wKr6tbgvFvA2L+rdAbWvWvUcyAYYcpOo
LPCfq4j68jmUqrtYciLJ8hK68BkIQbn9NC5QEhIQbZ9Ca6mD/rJx9xhIuVA2Arqi
HiXSmzK53FYjwu3Wg9Qz+NHCxnUaJFXDiK4Jag2MYEtoS2U8kHiCZZoMv5QY6BNc
ZnxkKgR6oSzZzuFbTlWJ8dICyLpSA+91+g4l86WNCtRzPLFmf3KXhhI6yWu36Yse
yt6IRvs6GVu3dsTOiqynEVJglG9GB022R4L+s4SF2Z34g+GzataIeXUQR3xw6WuX
TqkEzsQLP/iYM3IsjeZ0Cd7a1WHw3iXz/N39uL37nD8dXXxaDuGUA66gqrbuqeyI
b7VZNraJj3+paA5n1nxhD/CuVlY5zQYHV/spY4UXRlRbnt/3kQs25wUtiH1yc2Fv
wT4TD3TP5Lyv3+U3BPAe5/d8A59wetatUfxMOccJtURFSyDvkem961R5YWQe7AXs
5+TOoHgl1ksJOepGY6ckYvPSwWlK0gs6bvl+qpAD5yypfwdp3WXwJuoofKaDUW12
Qjht3ey8W+UGpFRlvVgno7Qe1C+0PdLzcZKd5naNnb18qyJpjAVESTEtj4JKasrE
gRxZcVpB8I25gqK8gsar75Zuuy9pLOwg9oKKjonIMrar0k8xCzGd1YhqClT+ooIR
J5nb3IrCZ2LMwHZ/V4VY3WBA4zl+m6ZQlTV6OXsuIOKIJ/Ke6jdj/z0tWJAd1PKO
QBPRjvULy/UKWHCR3mqeQFw1aLnJkoG5jyCu71X6bFC3S0lVra0VkOvl9f39XH5b
XtQTmsNT7fvI6RmYt7gbIHwROA2J32u2D+QM4I2JO3GQfrWnWyX2fZcTvEanYPUA
rZr0AMCCxOybR3zwkwRmFx7pNdJtCa1Spx2IPek/veDc5jd/BBZX6WzuXhn5SsoE
9Dpxzhq9AvtpzuZCQopFLYyYaDkuOP2KNsrF3PtITH9Rkk+XsDj/cudIXgimLlEu
4uG27VMLLMvVN6Eheds26/4JwcedHsVoxCRdtXHpeLzuO7G8iCFiUi9DlfdkOIyC
9dSg7oVbUrX2gW15hvMCd7hcml8cBWx6Mfpv2mlqo56ffYcPOVLvH/FnT15hQ8Lk
5gD8FGzCwmfmyN5GPEnmZe5Ry361STHyZEytBUu6jLGdc2J9BJLpg3nQ9srwipv1
vAV16cwPs7tlmifimbAGq1sbjfzj+RnMTJPNdMB8UuwCbYqen9Co5J9Q8SJ/eNpU
+saOosxkgFkL0IzyCrl0sx/M4cAACHdyewYO+WJYKIB2nkXvPBxKYXOfaLhN5d5K
UNVAHPWhUKWPEkZV+Zaal+vn5+eY5k4MnXKSHCs1aZPKJswNGlle0YTfvjz1b84H
4jySqkC5oiq1tJFQlzJ2IshZh8lHDKTdrlMs1cBI5eIp4ixFs6iQE81GDDRQNO7b
qF3+Al6835lMnGbv6F+4LFgRqoEo/kfSVL9NNdGXbuKnSctAvfCJR7pVvtDh4YLY
/LXZlHVDekAg3fEevccXcKNWqc6xXhNixDyoizjpP6pvGjSAGdEhBW7rEyRcRrFM
ltlP1WYbru7QbIXF8UqRxqpnx/IMkW2gWnbPLsejc4b/GIViacrfTvN0ZBEvW7Sy
04JYcsmUgjwE/bzFrBLEzj69qIMGLN1/6vWh3CBUfnS+PFZGdAk1STcI+6JcK2an
eHynXNNTnqmj4g/PS3789BHBzhU9wzU/yPEpy5epr99iMZ1qa7sA0nfY1ehSrji1
V4+57p80v/L5PIazbDu9LII+JhSKCyLNDaCm3IYLzjuB8XuPM16H3LLltdNl+qPt
7tByFADn85eWG0jztsVFwXq4be9jW7pRGuoLE30RT2XvcowYWgY0Xd3f4hvDCYTf
btg+VSLzINsr3AfpZCYYDU/xiwDpOwcDbL9U3Wt+xgud1s70izgV8GdcWVHq7m5G
wB8TzshKs+6ptupvsQXJY1lklN6U8wZeauB68PmAeK22pcH0d2dyrh6qHqErpUAx
FFzdWqZf/lS3Z0y3OPUcI/FnvXwLTh+n0JJvUDNvVQpKBeyavpOZeDUqUqHGBEjy
RHedEsfNZ5uo0pUQrShzReE1Qkp8M8KYX52C9yMNtGf2h53RF88UBfPOt1iJTDrS
U/gNuaAijkhUHjJX+VEaRcPEl36phFgGxw0KQ/KI5KZ56xQw8mjbLUb60MJSMdhe
z5Jj5zq85ne9wTcqQlhqSMsMtq3RS76YHb5OXty4n2PQ6Bu5dvLWK6+XEfLlrai4
HpEE2AdKhdh/jcSUzznkM30bvXAXGsLT947eFrke+2sDVGSi3r9orub0bnTgp5zZ
Iri1zrg8zyc48o6UrbnUODTN6sYoUhZazyWv50wUkC7u4SfI0EctmmlGkaKHD9WA
g+yBV1VZDSdmxrYJxXjpX10UWCkxkr7JhVbx+XUbv3XG+P26Z466dzpkDJJXqNvX
PBxO8blQjtC16MJGKZEHJ1IRmv0QfqOOCNDyJfttnj690XGw43/mW7P7PGoITsfI
jU6HGIN+FhtsPWSSN6g63bAiJXIIR3oflYxyVqUBpxM/+rp3U8DpEcKD3CevxvoY
o+BsH1QysN4kyhyZO0qEe57JR83f+w+25JO1ZmuZjCm6C+fGSSSlW9f3drgy1LUk
I/aUg88JwSjm7u7wop4UvgYL0Ur02Tp2Q43RQLcVA8XntMGN5CeUjXvRkc5wOX75
3wKkUJIDM0ZWpYAlihN7BsgItpHKWfpUHVQy4upMiCcJiD7/e8TKQjHPMWq4edhy
P6f9kyE+xQwTivJpScc+/SO7Odm7UmIBvtNPj2DlbzZU/PPiaJHb/TGbl91YTe5x
vtWQOaTYNa7jbxL9aKR23Gdp+me2xmMO6VfQ9vOfyqi/ZDIhE4fQaY0S4hzJRUpr
I1onJJePvfK7Sud42woTq39rzUiWHxpLqJsx2oGi2KjuAFumDA2zq7V+iYnZzkDK
l/VZockE4RheIbZ+GMAMqBznyT9P7Q/uloSPRq15TBNweMfSQ2j7y7Mh3Ww1t6Dl
DjvATE7XilimndvoMGFcCbL9srW1aZaxv+g+BdOjm63FUia52Pq2VoKrvuoSKZx9
IJqfLjMq1zqNc68YsOX/lw==
`protect END_PROTECTED
