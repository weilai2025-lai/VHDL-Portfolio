`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/L2wCNNFFQhERUYHkSjaOJj4dOCEi56f8vkPFp8YM8XEy326x55WkgL6pRs/PRkL
DWXNc2BP+TAuzgcykDdAkqV3BnUsjn9QxLsVA+r/I9JULHi+2QVWWTVWH8d7zcw6
FX+9mtxLcbGzX4+gxKkaAotPARoiJBj99NGK9yFb9iK+TMBfUqbnIl7tbeD7lQoI
gIHrn8Q5Rin8qPtXUCBC5WvjyiiFjrZWF54WyMC+KPUqplwBsoHidaQSg1a9ETZ/
X5zSxmqbxduSyLdLWbnmwJHT4Js6ZR79kEQEA/xt0Mj5/4dGfvZ6TSFAUf7EmRjw
riTk9MxsUM45wadIdBuo2HVlFz3lV9sO7qRPb36+KMdzW41rsxr3wmRaapkcoDWb
HL3WXEwVE6taAXBEjR3D5gPqPQY4niLPexYhTdPaY4rn6zGVx7iLn65ocqfKewTQ
WxpVnqptrYQ3ZHI3N6WsWJcrI86H/gp5rQGJqw6lYHpyQZ+uC/PbsaE3P/lY8n9Z
nFa3lEmEgkITS44N+KXUzgdyEwB7yXGF+jXwpwkXdsYcdPwYULkeMHmyJ5b6XjMZ
7GiuIbdRJC/iflH6Y2sxDdcVqot7QWktzHBOXTsV2SnIMbkP1kN9wetH+fo3Sn66
sX8aLKMQ1AtLyaS3z/DcuPAKnX7CcmGVeAzWHv+eWN2LZ+QkFHesT8mLgKGCb9Nm
hZiioiHrHJ47VQwn8FT9vraFp/3sqqlpo0SWjT79tN77vKxIX/ixlpOAw2GVZy6F
5cvLfb5mpAp6sgKs5hZdSbx48cOGjluP65VLSGyD+Kzlc/dtoEs1PO1tabDOlAwz
qx2/icLxXJuOrooCwPnKLRmnCEaLKFspt7hcGlF314AWPdcHUEERwegltOhlGr4q
5sskIwM5nVJoH/DcbI3Q7Ut4Nt1F5FX/Xg5I7e8PwicAx6Jjgdk6M7kBWHpQNLCs
lsX96pjyUK6fdlK0IUNKbNI6ZfckHhjF9sUvyW897uf5u4leQpuR7C7ui3hqMzwx
ZaVVDJ6x3ZIlKRNhX/sH15UQyYFuxmy1dusbKDfo2IVgyLEU9dRpa8T38RY6J/sE
gRfuI9uG9mR7PjFylnYxfabKorVdajPu9AMpvGKyGquEGugugO3koAottyibyFpj
U6P1/8DBTVcjDx0pjWYshmi0/NmuN+0JfwCma3z+A04qYzgfolTlXh5847Oyn1o6
2XLqdh535y3CZCxRFsFEfdjaOXpMnJdtaldWKo966ll0StMXEQDC4X1nUn1iOvMS
e2Y5Jx+rx6RpoU2ytCitDmCTgqGD+O3Ql1BknKKERZBa4VNSnMrl3wJPncIvNmKb
33KpQPfjQQLCCnjyyb9dK2Im++BEjL713NFPNhY85lifAc5qfw+F0mtQk1aCAlbW
3m563qadAd58bVpnner7plND29ETAi1CRsuUaUm44y4egKns52mnsviDXlU9Xi3p
h3J4H9KkDqUVHyCivQdnF6+LHwfQE3sTXUPPSAZzdzQ=
`protect END_PROTECTED
