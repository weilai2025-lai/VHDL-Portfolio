`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axNrOlobRSvvjaH6E1thQLbW4SYtV/VPKZxm3SwDoayrAJozORXwSV9H1dZ6NvU1
gWobMZgEVHHjNUmZtqaQ3f2SvXOiVoGMvtG9FydfUx5RmMn3sv/OGTo7PDXM5+C/
EN9SNfL+jc2SUKyPYgvPEiYMS5IBp+u4kGq/9aFrFfXYv+0uyjuY/x//0LRVm3IW
ZxF/0aw9gNmq2CmppstcEfDq5fDxawH2E/rOaNxJ8NsmBQGVdoAYlyDVhvjviMuP
V/tmSv4GG4YYatGGDiNvrzUJirvRuagN9S7Fl+xwDNHv5wI0DGkz5BKsdkXWgOIq
yjsaUz5UgdsG+N2QgK3S1ddZrFc9KT0iJ3MeNPl36XAtyDgLIXNmQDh1WQ7+tj7V
FCSGmvgoFQiz1gehDRKTxlcTUHKYBpeBmMjYx37fO9mGPUarrKub1NQt9V4rGTNL
0AqwoOoZtPsNIn/UqAxIIZZVSJsnJelWLiQN6P9aR9+x55tdFt9QdshRG2MAOt/k
zMelnRWeauK2jxFJ0Y1nfYeBXkUPdZg6piulZgDctGxrFOZIv0shquNM3d7LOljE
wKo73kiIz864et4xHa+MBcJbvW84327HyIQnRlFLB+KGqY2aBq8/xu3cf2X+T5vl
/G+OQL0qBEsSlUyFaNREdARXK6W3IivHrB5oDwSSgrmseMzM9ZPmuVEhbw2Fw+OQ
1yQTX74nIcFUlwma8nKmdkpBGzjr5FaUc64avYdVqUL8thYKXh/a60bzYAKCmOek
zQoFoU5IZQbQqcxAMo5Z3reTHbCQEqoVW7xl/AH4OwXSGB05i/cyeCmrPERGWc3T
uMBND0aqmb48isy9pz4nKb7PkRM11ffNvJw5WowJXPrLPlOGy6Q+8+NcFYvHaDZJ
mm0yDGkCCT6TyzfjhFVKXv3y2y0Y9TVHebRfhx59T6dvZOuWc0735XKySfFDg9rR
sS1Ch4y5eeGL0yAo3ekbpEWfBnfphtE55KAU28f97gvXz5SEvJkgEkkb9axMHIYS
c19xidzLz3UzY3DctkxjvidMziLwUGU2jnQ+UhjsBzB2hen+5aESAbVTHLEzFng6
rEtno//Zgfhc/Kv8TELp2ZkJPNWjPYUNrG87UG9/vVf9OeSz8VnLZQtR5mnLJoFo
gFWm9t3xR5Uo2LsrD22LM+8nEqneeJMWePzpsKTQbtBvz8VJt/ZTFEnGeu9hRaPD
igYCUwu3ltlq2DnxcRvPWxtDxAiDKXUP1w7yr4TNebm+1zaOzSGtkStTVx0JMEqi
lJZZ/XGoX3McTuAt2dvBF1nxmBSbGNUaaCpDNKCDE6nsG1RrBZFm3SwrKGD8bZZb
jyuPOtW4YP+hYyMMCzEvgLvfgrZYyvVTpO7ZJ1wHB0xBIiRpZoFETDg73/Bgolee
UoOuD5IWYnVBLd8TzmFTn0iWsPjKU1IFG8/uk/RiW444NYe+Y7tL3LVGylb9BnH+
vaeEF9ztktMi/3TkFjDnov/af4ixrfcbUMjV4ANsYiTNH6Y6SVubtMqS6JIFWzIX
3W4G+rrWA2rmgzUGmY1N43ifZirhOsLaaLRBkFDAz0NBaeikpjOvrce/Vjj0SfbF
NONKEXgS4zkot2O0kVBBilXeXBMwVUp80m5AzJ3iq5Mpu8toQ4KeJIaStCnhVMzQ
bklhhZFXB4ALMsv84lbwc6OCJkq3OX4U8xOH2obv+0eZ39Ewzcu4qR8QpyLxskcj
jMJBNnIzne5cif38m+OcekavQw8BWFHlBSda+4mXFsSxcTCnq+h6zVJH9QFN9U5L
K+o0ivBIQUboGiFh+50zHCaR6h6rgS6YgBhPajdtHflkqgax10+0v6YZuqQCi6R+
r79ATww4oT5pgnv0gsQp8ugnbBLcjwNQnQAV/Ow/o1OkLhJCmdl/odREurgBMu5n
q8FqBNDvBmNUpuImvUe5Gg2bxqoErAoEnOYkqJ2dW3JNPfBi6I305g9CSVM19zxq
ioBas3D7q+Nk9NlsRKTD90gyel79tuX7NIE5r/y/xP7oib5pqXlpl/TNHZjrZnxq
ZNa2BYDNNZvqeY+SZ2qmt1uia/dB6PBId8nY51jlT0AeJDBurDdnblmpuljCzcdq
1U2SO7jyAKIwyd3vEB9egtI8bUWoUdXY+SFlY515SHA9Qcs9GBfW+PpUjtguB7U8
jL8AUKXr/RFLSdRKBryUaG0C9y6MO5LF7s4VBzgrFEoP3HQhpxchqAt8ncQ5NJ+8
vCRVwV5myto2GO5ILD/cLELf93nQCvgXS/Y7dErmWmgDdwAOf7orP1u1fCzW1fa6
2r6yt9xG9eoqqoZJwFRgj0mzxyl4YfJ9hjt5tHa7peLLNReOr32oCSh3lew0BUSu
q7GxxJKqvi9FScPtfGtxUZncPGDYUsFKTlaJZDw0mQfegRuYRlfePO6EzpOXa2m+
LvH1yUKyquB4MqGwVyWMTcvawiO0PgVLOCyrp+BviGneL+Ap2v8KCUzovI7g/MWT
B05lF8ec1uOCGcjnatjzC8m5ItAUFwPpyccv3np/iifzJ3Ptny09LkYDRTdhXexS
XOWXo5NN770bKMNYScVyDFMwQxxD++c+IwpsbXgbG8TJHaRdSZ7Q/x/MlM8bpWqF
FBxEn9RUf/sTLBX830sHt2CdEkXeVhYZtdONxIoLa1Evwfi86IEr38QdrbMD+Kbe
cR7PLQqfhRMH8UFvt97zGeFB1/Oki27fu6UE4jxmRxgvR9+jhChP7cD6TSKvo0AC
pBqjmDWXvVuDGBUmlCkPOB5Q5bOzBRk/Z7mLK7IrZE3OcUDyYwcjxP55jQuesm1u
dICBn68c0qsrySR3o7HVkMbVVwtglOS+qaKyedESrtACkpjdlArxXNpfPMdm51TI
ViZgJBwxXt2Jfggf6TN7eoDOce8BBxjyvvqZ03VBo3iua/cdHb/fGKwaCEv89Kfo
WL7+CzmxXG86aYCG+HwsVnUNL36fj8SUV9GSF8kcz5wnfb32N+R4MlrfdfHgpoo2
Ms9vGn/mDDq+O7rImRNBzesifc2j6oDd73uI4r7w04OVj8pfOqew8p5aaspyoFHe
67G9voTlEN2Z1tKomXa21+YqObvJINJkp/5mnL7K3RWmNaR6Wbh71gqeLxTbbT+c
hAD/5CZITTElViy4ghIVikVlPR01ufEpwgSCiulQZXNOjYb1uJdH7ccudD3mrBI6
SjX1dP3F+uhyUrrtBWWEzimx2RuNRCb3SaSucYMqBez5jlWfswCvVSxBTMoncHDT
2DejuE848F9Vuy5+zUrkSnm04q4U2Oa+rGEWMzbZqUKD2IiF5WPChcNCsHFGcPTu
`protect END_PROTECTED
