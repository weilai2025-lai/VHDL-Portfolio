`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k2KvHPKGK4TSu9VCEAS/jXQJwAZyBgtH6XUzVOu3On5m7A9h0yYcdInjwf7ER3kt
F6xKbnlAH7qXVqXxksq69Kl8hhrmI8kH8PTg9frpEtqQ1tGnEHRP8NR8b1xpizX4
+Hh5LOahmc6b24QPnWnlY1Ynwb3VkwzCQ//Jev/G4IN5mwoTRohZQcONBFzZGp8k
wxMAd+E9qp/kLVV3NrlP4+tiA69xq6QQBwtgJVZhCPxSniWSNxtveOav1Y4aAN7T
knrY5Nu0iZMtvXZxPEME3TSEqwjYjaqHd2HUOkizzkynkajfv7ILiuCjXfKvhoZ2
U2VGfjZpuogAP1X38wzx6xTYP24ZRoIU51vcK10nP+4YkTcj/sOqDr7Ng58BpQXx
R38eFmiYGR7tBTBuy3kL2FFAUKJQQCmf1dyiSpYkVC4p/mPGsomaOnJKl9ftxBPo
1X9lqhfPhNZk5JNRDftOZOyAAF7OgSnO6Ulvt+jJOYMk+gK4qOzYI4Ibywb4MBY7
xDnJa3QcaNZOW09JvJHXHV6tHqvE4446uDSOWKxf2u1gk6ShtZn1TD/L2AkxeDU/
IkMf4+oclLnI+8AY1Sq9++zuVJt8fCasOQ8GNAxKqx6/+5c37YT1CDS5Fp1FdwnJ
k2oWvSmW+W/yDSMY8fXd0nn49JdT7mLld4468aaoOOiqJmhqNPh+6oZWf5nr2MaZ
eDjqE5x7cW6ZwzKM6b4kxnLI8VsxPQXHO4TNyYueBhQ1IoG7Q3PTydR4LfgMTupf
eeR/jpzSEUc16SbjCl5l9QsnfPTXlb5/Cuq1qyUVSuEC/HVRm2S9ixAcDbbR4qXY
JzrP+2gY47PQjbeJD9+wYtw9Mu7QtSHKgaVtawk6nbac+X3nuL0Q60RB5o9l/QgG
jwvnKuxtVBGjnyO31DQ36IZWuCkFtfgTnq8jVV6E6eBnGpDGuZkMLsRHxU1fHNWD
Yu6S0t+7rIncd2Bzb8bYaL7KDTRMPoMcUTcylWH88yjbnGuxolEwfue0ytR57WVV
XBQYTKWaWxQ19CeBdjsicRMsEZrVwBtzGQSNQcUX58P695HDnMw8r2FSbp2SbXAZ
l3mAijIXgU9Vbo/RqlhXZpb876U30rMbL3X66MGfk6TkfPMyJXZGNGdarrof4mHx
8kJIdrJtweeNOvQb+SOp3hSushGGDTIEj2MYWMSmyt3pU52KiGm82FzUQmKPvU+o
H3Zo/56Jcx+bYuupWLvnMRaHPGthv/VTarBbNtV628dDznk4kFIlAOJpCR/Y102t
Ox8T2mbN3w49HTK/fHqu0dqf0hGOJBHbzBvkh6s08DR4VOp/OpoZJIABmgIiJpVo
BPKC2o/RnLzRnxy2T6lEF1iKsX3Yr1BJNFP20IzFIztif+7Z47eMV8qafWBxynVU
4pMjoFKGP+PnluGkPbZoXGwTZqM63XUy+XYmGTri2IvRx3pUQkaLgWFWSppXKHrj
CPuVX31OMcuADHDVsG/97r/b6ndJQ7jgPnkUPtVG4YEeygOpOlO4nkjNxjQ2rjO2
8H0TnqpF2Sa1hk1HtJmaKC8iwVtqv4XUeX5Fvu/TjUaFepRVpAiwb91PFTrj3je6
oEPfGuA9vRnkKybvvu+LyMoZVtuSYTIDpOoDmfvo1YskMsZtXrnRRKApkgcFcdhE
U56/desUpTobA/dkOAvE873IiuNgyY7KYlrCTDUWxhMgYm/RqxDZDeyl6EkwfkjK
edRCaahdv//yCeOXA2qLcLt0hODfVZ/gjO14kAqEv3YjT3Wam1VlTNALYwJUr0ZF
lX1kCAS5Lu3u/Emhicxmnk+LKl7AC90kvem3v6jLc3sXLDQFkv17LPElC1GTyY4w
vXz0dXM4yrexzVvzqmUQDGvSibWVz4cFuTq3G/4w0BwsDEWZQDftk04YLQnMVI5v
+Fd0tClVqkRqwR6EamLPdfACxGAqokSgWNWaSwX6xe2Nyocd/uipGxMpZPh/oA/w
RZav/QbjLsovCXlLUDSK2D4WEJZt1J+zNtbiyqhlWBpjfZH6nVUTsqCrzL1dNyFY
qfOzTunwCHIl64rLnoYFi48Pgc2Dcdn5LMwn7Q97bbrOxsBagJGKV5pPZYJHCyJA
pfQHLp6iQsnKIAy83atBf3NQZ+qFtdDlNqJQqSUUS9khJypK8WL0d6YeEXnUPhXg
SYollC3f2vyaQu+mslJarZrFsv4LexFgFZwverbJWbTQOolwcljS+AjsiAdK01+o
mWXmqupAkwC72Ambu7c50F4MyE5mgYLwHL6vJvDJpfDTZaHwdXtPEyAYgR84LbNB
yxWyk4Q4UhYHDd2TiPctgy5x8z87vqzpgvo4q0xcN8a953Gws4zSMrOtFT426eQH
xnRrxxLRWcY5yo11M8LqdFV7Kj4kIzcejTEZxXC4apXMheP32oH9PZonw7GWfBnd
PXEKeo0+k3Plx/O2ZIey6p+JBPge/cz/xTx6d0JtuxqRdjJpqCGi2vEn0aTItRJn
okb12V9on5Wl/XrzDP/a3zNlYMXOeNxnlC45oKzmiu1kOEpMweqgF1i/o4i1BzYQ
qezq0kJGcpMDp6nlo/JwRDHzwxmIkCkBSB2wFpYchnAFMWZYj0dVX39Tna8me/0P
ymrYYBCW64eeqwgax/ONHivKTyUIFFVNY2B4BmPmxb0=
`protect END_PROTECTED
