`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rg+xk6NosI01ucWG9QH7uSbUvrlQmDYcRQ0L1w4TlxOyGZZ64OJZIYwYneKWsHlY
QLfH4UuqpnqbPSSBUfdFXNXmGn5VoQFZQNXqBCeTD7he1bpIQ2AbnUQDfa14z040
vcNpGGNb4HaqNPO/pwpRv2BQLnYYdI++FXCH/q89ccH0OFG0pResnumAxi15RJdq
W5g68Oq9izB8ottRiM0FiWqRLagxmeKcj22fWelWrKHO7hGbgWKY48e0vgWanQOr
prnq7+R5hUKFBe07/vlks2St0DsNFgg/IrFk6dpuCkfN8s0LBz3Z8L+5rH+Q1nvR
MNLAh9h9uc5p9LsitMc+CZLAA3xRjsqkOImilJETwLkydLTpdxE7Pk4A3PuerMGB
oPDhdASmoKok4+GwhodkOdxST4XtA3zCd2XLp0pDXRDMKDppHSOWP6WxQLp5n4lv
TznuaKvTdfQKEhhIJnuS3WhZPC+9lh4yqB0rLu8hj+4SZ5S/OBMlfaamWFS6wqVR
+FwQJakWz/UMr4WWErf+WtvvhnfQ1LWJGIVlJuhkGVfKbhUuQ0/1AaTIfdbplT+t
5R5jdQO9ft3DPYvhWSQiW5KDsTgL4C0Ey5O+Y2egrbQhvo5z43c0/n6dwT1zLHV5
2LtJi7AyGHQoEZkDO5tQgdRjeLMVooZ8ER8zONZ1E675Kk5jcrxAngfxIAT77c1J
O0wDEWCd8OD3KBefa68M3TK2nmheykP8CJqi2sXeLGy+5R5nNMJZh4FxQOyscYRa
cIaCmhA6/3CajVhlELOhD2hOhNN3ZRrcOAnZTpJN8ChWIhenTrrrLI08qXwB2tKl
wN0Mfxc9O+uXifssYRIWjEWRjHoKRVoYKk7u6epho8Wf5mt0+jmY40IJlrMqrFus
yP3K5o5+7ayq7mK3K3k2LQmXVz3o0FVb4BAhvLzp60M=
`protect END_PROTECTED
