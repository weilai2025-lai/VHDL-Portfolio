`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6X6d8iv6h/TD+t8TOqyq89VktI3dMalWfJXkdfLxAYVN6BzCxomAcpwN5XXmvJJo
qLf2akYbqZaeiIeg6ENr+yNL6bngq+R8P5rNWDfJrY5R7jeGAtHOC654d6lgQB/a
f/F9Iw6y42XNcnFLu+KQZhIHPdDDDj2WIrkgjT8ACAvJwNhq5gjH22sIMpfxJ3CW
bZ0MCebKorpbCbDzJFI5YA2mVsCMiHFtetWgug6hApQGKMnDU8XG/R7qPrPQGClm
SSK1dbneLJ2x1zSXTfwzLQw/uygLZOJV4FvxnqU5NhuVXJNlL7pgJ3Sx23nCpjd2
4OBtcgLDhr9Kj8VttddVI0WDjQQsmYLlcG5tvamiZxR7X/bFwBEAfjzmY3mkugFs
uQVMEfbMSopudfjBeP0rgLazIxxfsRdfKVo4UPqJuPGwId4u0mpfuRo8jR2yBlaQ
novhLFkJjXzPMlRSzcdgOTHdNUy7Guf7gm6FGLfuwzacSG+5bOsMrI0wvFlQ2lTm
iv1ncQynNJ93l8fYwjfUjyB11wlQIRrsc8s50nVzc5Hp1eR4nhzaCGYbz35De9Vf
/HW4T3iN0VHxHupfNYlIh75APJkWnAP63wN47uG4/OWWHNOh3jw5Cd4qK1D1V9RX
om7h/9DJm6ptxkVTFBbY5OnpFsNIwMzDyZvGhx2aaHjQ785sjr5AtxlZOj7DY/WA
j0xR/DGIyMorbxBQCPAkjGfwnniEvmdhwSWmgojz5xBXUZIKV1x7+PY3IRHMbUuD
TYeckQC5fHgk/rsKxK78YR64AzQ8ZRWhoXQKeJrAvjRE5VDerCiuapx3ffnTKjvg
7pQuNnoNlb8YfTvIRaHawuwFvWjbjU1Q3HeoJqiWAelIs2/H85zTkxU0IKydSNfx
aPXHKaOWqANJnvzva1RU6dnHY+vVHZrkhWaeu1QgkfZ0/uRmVUrGjsio3QIwETIE
dS+xX0HH6bV1tFgjEQNujvY+UQMqbcbRlzz71PqGXY9oRom1ag22BPIyN28cUTYL
o4l48wD36an01RlDkjmDr4yX3J50wQqjCv+H4Cbo1/8cwTCSUMRxGhskUcKn1EGb
krCJykHi7IyRx/2gx/09eW2FUPv8oi0X9oP43PJsWF8grecVPgnR899Csp9W/jC8
5bsWcz2DPLDs+pBv/wB/J7oFoOiqB5Emr01ETDcKG+y55XGkyTrWX/jUN3KR0teM
VTvroasgnP4C0yovrNQ9TFcesBjcLM9Jb1pT9FlRbytO/e6Vzh7laP6htrRACPYK
E9+r9r0hVTCXfDBCcGDseVbUZh9vav8UnRdU8domgsJu24QxwaFpD4vfVhf2ruTr
A++4hPaPXBLOWISP2Y/OW21DFgy5/hditFp56MIsUfqWEo7lUg6ev6QXGAtSyB3V
pyu2GN3Oj+5ptAoNsZZm8GuJq+hr2UTUYP4RfABFjH+7qtL34Ko7bagQvF+xvXgU
uD4II7RbAdn0SglwMFS8HCInwUL2mqwUwXUerXmHROaMrjXZyG35KVPvdQulglv/
ob0dZaRnBh86y/DGk90xNM9R9NhAe3Ym1GeXuwwkxtAuKScsdxhAoc3hAWD+MEkr
PeutHusTX5J4n2l8ZB4weaMdLpeM/rHKwQngCfrLjoEMXuRtEAX1x1VGjBRHdE3Y
GbVnb51TQoNLYeG9nsw82OV5Vv915xSV+JkX30vwmlcZ4HzSRJKWfbYVL7Asqw6Q
kf7WtCrmfZpBD3WtgDVO+zYNIv9/vKOjRByg8U4ADViKwbaT0s7xcG0Y7hmpOp6I
9G+OxNf6JztgurNI5G6XtHxXYLfV3j/h3GDQH+dSalZ7+wwZqfRCyC6Ka+70ZHms
jcOg5dRF0YktCUibo2DkiZqG0dfJesX6udcsT90dpuFyB9jIOzCV1mSup38Ft+PK
qcIfzWB3Em5bVjsrHzTFUT2RbUhOuEubxAnvuvKX9LQiDjpWfJpHhodsfBGpb4st
itB24cN9oCk2w7iT2SSHuK/frEj3QvG2fwXa7ag6PBXTQoxFBya0TdiGXJAzZmo6
rorTClUXC0c9MQp/zL+t/uqj5NWS9JlzV/gIc/hMK13oRlrMNmwqgQsnx4n+7fXn
FMQyAldV6HlivQWkI0FcnkKO9W9VpjjEaOaBX9qP32hhZmLE2vfELds0f0Fv9nMJ
eOvchNokqVDRx+1IVvt5UqEfYyt9++uB71Hf0B7QnUFCKoR8DNJbr6ngfuS1gGGV
bW9Z4+uvhrIcdd950XSZDMFCpKY6a7zi+4OiEAVF9b5dFCtThZfC7hPD++0xzqT5
zZsfTxcu22WhG/Vw1xngBQ3acpUKZSz7HwcAmAaC6L7HwSRx1Ou/htOhPr9p26zB
JyZceedQikFo0he0/ITIPv+Of97pNwys7QFgHqsf+hP8v2/R8dQD728R3j6xT9g4
EtcyVNBXmNl5FvP3SqOLsrIg0jRWCIVX6gTVaeDRQHTepesY3fTIKmnp2n5l3Cax
wEwd3nmQdYXkP0YU1WXFxYNgnO+fn0PzktcvLpogus8L5O7vJ+AH/xvon//x5d+i
PUWUlJzKqf/nkl7+JL09iXK6PXqmrZNlr8L+gd9g3tz3x1fSw3miqyFAMUtFDQnT
RpUtaA1wmFCUM6lrhv80GrMFxqiv0cWIj7Yz1YfSllU7bor3pYyacFs8pSKklTyW
HC2lWxUfvNfokJuetH7it8euShnx5lRqM7gLCBJVPB5BHHqElHFqOURU0Mdnswk0
D6VHxvMKJSCNVL1ZQvTpM6d4n5DvkVXXsYX0K4DhluO2OTACClkKH7tLnS8e6cnL
60sr7XEtEJicPgVGSIINmGDxw0KUPeq415bz9F4PtHzFQoNyXYxflH54BJTXrV5x
ssOZ7X+VQZ1Q+h1EqVtw63NAoNOXWZPRRf2UJ7v207Bz0OvQQ91/OzioZJ/oy9kn
p4vjmtA6uzORHMfCTk5LEQM9fCYpq+JEdlz22s8RL8vm2MV5ZC0vOmEk/T91+vvK
qKkqUL7vxyzpR/5C7afkBtyIgBvlAqgedWXJi5b9rpYmWFssNf7M9DkZ2UB9gyqa
G9uoPOvvJPaO/rIe5g9rKBFxtW8lE9oVkEXH2rujAOODBMszZjGYXl9rW2XrTsmq
zE4RMw2x7eff7Tqq+WtQSLxxItMIGUmvRawvp4yXahWMX6gLaHMra7YREr8wztrI
xu6GNtWlb907XrGXW3KwqZetbQ2GWJz2uSjZ+9ydyAxPXKE8X4RYM3oD0Lv1kn0q
jWj4c9bQ9wIV1lAkZZNNS0LCMe+TB1d0JOFzIW+lnaQWMIg4KXfAh+6hYSLZvWY7
suR0YIDNZWrhXH39L9pXLI19n4kEyvlrBZcZ7fK2mZmu5QQUz64702I9S74XbU5g
ZZu6pKLfL/edxBxP6nDFJhiSIwqSPSGsEjtT1hRF/0Rd7c/A6XTCpCDgNBZLveDL
IfJLU7CWVWKLO6Snxh5Wmdf2AB7/2wL2TItwwT5d2lffR3fSJNpWetxe/siKqpXs
Uk1TNEOnII4nGMCis6SnIJ5neoua18LkjrmIs2m6DruAyZk5cljHR2EEW6XIgbvW
5tlpKQZfVZHOhLIPuO59ixfN5Z4DwgrPTTk7sjYkHepBHn0fdPEIj7c3DpPEe1sb
aDKISoncrDXHrRfbsi+7FXYyrCTrNVYT3SnxC1JtRMFKdXzx2wbpw90sKWuDq2lC
zcTHKRl/3E5OtIzAiRdXIseqJEmapVw2xSvrthD0pwVcMre0VxX6P2hGpC05UviY
kkiEgh46l/xIybvXOgbTiCU3IMcPOxhkuDjhhtkc7XbTRhluauZtWYclw6WlHMca
Pllv9G8843b1o+OeDoyQiZ3xzNQKbyevcm8g+9yOv2cZnOAAlwSOnqMp+c2g9+11
yRavqm1UAtzBJKcPTeafZcGjIcce6McnDaElV0EbhD+L5N83BL6EYcq/JglXjfPS
smABfW9fHrI0l8XSgwsAz3blxzWDJKJRD+y3cmy02Z6gmGET9ghXySl9k4hV5K/h
wRY4WzqX43DRlzgP1KFG8pbkPFNh4krJ/AkU88qcpz4SA7DIGtCCLG6GC6zX1sbY
jazXx6owLWQI8SkP66OZ0SLXLd6Si3zGY4J6+PnKRwEaHOXxJRFZbF+cjMHeVjGm
LA3AFOAEWl5WDn2Gdug+iZPNOuC9NxVfzqDympifgFUXcjMrcw/hEs4Vmo750fkn
Di8cuLp8s0hcQI5cQfXFxSCIYrOuvthXyfW9IdtWX3KexaT+to8+gMCS4Pw/VJW0
1ex0rh5qGaSGmS3jP1/D+vMrBDe2yWKfy9dClZ1EN7wbX9LVM6yVaoB06BP2k2EP
z2ytp19nFpY7qb6s8jRYS/JzfPtZRXbcLaZ5aQhB00AuOK0TkpIe3WbbpaFJ5JDA
Q68YXaHziviqT/lZVXa8hmC1KdGxu2HYbFyIbo+6qixbRp1uSAu8J5WROS8GItEv
i0hpdYwf1Qm1jHTisVxfGoZRYfod0i+VKOcDowh8Ol0Vs1104E+56bzhF6FaNr5w
tEVDavx/Q6A3tZSjh2lSV9tqRcLrZ3+y3JxanN3NwUrpjE+0UE4jU3e4ocubxMf0
T8O+tjAZLTx0V2w5cDDXJrTbCUT8ZGPoQKZIrsI9Ub+mgvmtEx0rucvxzsZvPYRp
Qt/1eLQ1/vKoGi+t2NGhYbd7zSwayGZOH4EnzjLZplcxggng1IQD9RquPt4IDBVQ
ghr7sV/LAs/YVHiEqA0ePwJCZOovV697UA1l4EodKi+0W/zAJmPPPMJVAG07nhEk
96c59CLShiqR2yoGxGrQciUja729iel5hpGJc27AubcqSA++1y35Bfhcftxfx1FY
DPHWhPfewa+HbSzem6HGlGnAiVO7aZgJyXHWiSp6q0t2spLypLssohWKt1njX79u
ZDpHOZiawhS+Gozsh2n8GwlJvkakGv/E2Fn5WI6hzmc1ux0ev6Vrt7IlVSwAOdYI
ejlSP4VbxdCGSI3poUar2YTfThrLQRRNOihvq2kkEh94Ti2AnUA3pts2KoppbPQ8
tI2TTOUJXw1kxScplBKA3AIofXx9cRtQ1XYtCLc4AWnzb+1mtWIY5g0c4qKmG2xV
ylSOiX8cY1p5zMZO8b8Ee+1VlNqYucqCu9S4CgeeQWjGZ7d9ZYpWa03ySr/IGXWP
WkH0XalgH1o3zAB4jLyAXlfmv012885/qv7y5AhzHLLu3uLY9lfub5tm4anfUmnL
gYklJXRhdpBYtILtuyHdKyaDDnOzzxDmc7Kofgu5x3Hb0kYLWL1ZiQwtEwlWC3Iz
/Q3pTowGOMyDfEegpvD/YPLX0Ww1wREJ0/e2e6hfY0vjszh32BL7TJ8cIqKSfIHh
jmzphqQ9I7zszhvS66neGuTYXHLGUwD/DUYgqww4iWhFXXe8L3L16UJxGh7YS2jF
8a4az5ejoBNYMeonuTCjGmfym+1FFQdTCX5LCJzjSBYj6pTJLVWbxdNsZ51e6pEY
RQZk4thDHt1/B4l5CV9YF/Or7O4cj/Z+3C8wjaHO8tFQCQTgdQmvsSIfQOVVO60v
z0Kdpl4DU8NO7MQJaDnQpFXpJCXiam3oSIRdLiYlVwI82ROsmUWNIqglfgIFh5NK
5z+sNoXd1wwgu1vBUaYZPFbprQF0Nh0sj7WukkFKr5XRHoGsFEj4KRhngvJeLETH
pIT/1w+1z2yT3GFH8/UYfOlN617ha0MO2cQ9IuHG54Hxg3CFjdcMCXNVPsHdGZoy
wSKYAw5YxM8WIB1BB7U6Y9HpT+IFIQsR8bFK/c9FFcZUzXX1jE+m+TK3uuIPOnLy
L/FgemeUJAkNCVXRRy2bOHJev+MRqNSyD4qtoj656cl/g/BO6HjbzrTNEe44r7Z/
Ble5ipmiK4qZk179H9XDbkKqTxLQuNhQlgmDbCDzDz9yeV1A0so67tVP7qRhNnDr
cLleNwvop2qJiT5Fe8aWvuCiCjhLjcWQM9qpe3meqwBjq3PRtMXUhZmkc9waoGC/
+EL+InpSTz+FUnLjlJEUQ3wNufBpHZ2aiAMyrZ0xy95EXLK56nbhZqOvR3xqQfiq
65yIwe2licAbEJnd64e7y0BJRM2AwwDj03jT2dUrWsgW41RcSDYSAOpoSTX+QDGy
nnH08yedNcETFCAefvdpUOhSzBSXtpDNeQpRcRVK6horn+QOUYDLU8bceNpFdL7R
S4mXXF0BDbq+M54/cM+mwGXfDD3xJ7/vYa47XsnCQjJHwc3zCjlDTUad4RKWjcN+
HsL+famxap3nI24PDDsr7FB2DlQKcqeP10vAIuY3ooH4APO8uP4Ep6IbmZOr0mRN
iMHa2vUL1xDL64BS4PtgAx+3rRV6U0PihX4So+oGlt4K5MLDkqDwtTOeXEsG99gy
DBEorkCrjQg9qtEafIyPmvAeGVPlf5gam2elmaqOxGaUZxlqZXuWpV4rMKQRxnqm
NS8y0cCB/K4xffcS7eNyABhNO3KIgZb9VTZ8Ae/BVBr6OrfmHnPmphprAxIJ+xW+
fWhtcz4TkpFqHv7vbjJCK/I/EaAU5GCkWj6SZiDMx1JPH3RCt7rJzPx1RMJNqlRt
vZiV+LSx89F6vJJxop/S7uztQ0+9fLioIdHsXcOPPdcVGJOYa3sHxH7NM3xVcMh2
mMfRPSYDMuyHOABTRy4UJ/kk0CbbSOgxOogR1UMGYXrYR6dPYhS166LDhwRnw9i3
OjpFGdgxxwwVerH3L21GhaayW8RXx0AAWDokwwbkJ8KcNcxdO4OdrYsuRcEy1ea5
kBRNe12/TIy/2XGNpo+tWHYnBrWYesSgi28UoUT1s/43sQscz6ntKbiqBkeQ3el3
h8MXI/DE61IlZlUakppUxOUmFoIEQv0CscUOMca2kco9bQCY/ZMAG4hbknibMwK9
xqWbjV2P5Bkuu4AzzevMb8MxdgKhbtP+Yin2vZVRN87wAkpkx7UTbsmevYpQSsc9
YxLjXzA2JGnvxehWlQWEQzwTxuN1wcW3ryDbAEA3O2+B42dOwSlVkyfJN1mh6Wwt
JX48JEe/U8dv6dO0U9w7Z+rt8zmzU7bEhcDXSIA0s7kcexIYVFx7pRPZnnf4ro21
Fad1mLou4HBtKLu7nxkNg7YYfCwRGOeztkwNO2QSXKnWnPXhS9LfC8Ee2E7XdWCH
MxqfTb30nehSQxaV7s2O6Sf3w1Rl8hPA2tM2/Tl+d69LDWV4IEa89cWvzITxn/gW
IS158uKz5+d6JBjuqN6lBwvCDiJf2bs+0UHvlqO9jbx8v5gZW9iz6DPSdVGi7Pnc
SF5shOCY+YtU/VaJwkzU7ekoE/49pOlEbvR8aboMKf5sDrLfCNcTQmLEWACovjWM
p2pB12haDTu/D+Ez53Wbqi25qCkjxvUzJrNX93vPIaTtGVKq8Ay1rub7Iu0zCHtv
JaTMmcXfyU+9dfznyvPjScZFzbk8Pm0sRjULfvSIVyexE7VnCsYj0NYHcYG++gpz
fPBL/RQTIHKNSy5PCOhSv81alr7+mhyHq/HstMFBLEm678wjoK8PoDsExhkPsIXx
Dx2VgvLwhT6PJm9rYdvTegVIaMNy75I7jOQkaHoknmTbh3RyBCicdR+iLmTLnbut
8e5/6DFrzX4jt41DBy0h/zA/Pw/JOTyNmY33U4e+tR7iEBZZoGJZYL9rrJOQ739g
4cqomEwhFq0tBHfVFGBGnfy2iuM5XQzrm0K11Gs+7qC+6NEh51wxaz3lBwwXP8me
SkAibGUsZN+rbRFQ6Ym9Zaa6Jcdfe7tPwzyVkUbBc8Pt9ssqLN1PrIM4JYdejUAp
/DqyL7f5PoacieAwVU4QSR+cc6ntdTeAF7FpEBJNdKs/tzZLHH7K0KSA25l58O1b
F8+UGVw72BxRqN5MzPyq8YBLvBOU0Txb+RR5SPxtmmHZRs/fXwSg2K+hOa2l98n7
B4fwQzE67pLA1nhNMt0KHaW2QIrkS0X7Bap0/JPHQjbX0g+PWjhgiT3A89e9IUSI
cpkY+PcDvsnGz3z7Nui9p0FebZPLR5vjpKwgebjy7gNjoUTyUnAYBi11zmdbgHy4
6mDW022IRw+rZZYio213pmt/bGos3CwQrWD8Ex5vYquEZS0B6oid0rTFZQkYUviO
DuvhaP8NdWKajr0Mxu9Kxt7nFhfyf4U2ZPdptR7aOzXF8nqmGL125TXTQdjQgo0a
5PWqPsCLwe3jBZDLj9e31bq7g0b6mlGV8mqDyzftkUOaJNY26PV5SYyModBm8Bsb
PuIVXVJ1hU7UVNQDavN+DzA8Cf7Kn5SDM08K/J1meTO1cWu5AEYeiuV7O8VX73O5
dBSNkkFUg6SzRbFl0AJPCM4VP8F8l4qbCiLMltjpa5k9d4YMxVadV9DpNs9qu5dd
3AAswSngX+YVOrXb2EUKn659wmOrzZ2HASDxe6rbVb3qEVaJ6vQHtSzQ4rq0tmUG
gaS3Aw+8MNp43h94QaWCs2cntOLS5wzqzF5Hlt3CmF5zZlDytzfvCM4ZGvIwz1sc
95YYkTXEpwr0zGuIC+iLfLiIu6L2qKEj3SaNmMsvoBaswYvHmu7zqzL5voKUvxXQ
wIjLgU6rSY+aDVghrpGBO3WIo5qxdTG4ywjmEmx9Pgp9y1FGozZ4h4UEKIIQMfvU
nHECERIDbCGujCDCuUyIRMFMg3JCYK4scz0mkaqAiS3QWuvjtl89Kq+cBlaXQO+T
awQ52jux15rImTz8+efq7e+xsPqvU9JvWHR8+96xeNBeRfp45mouko+MS3gCxneE
mCl2iAuFuL4HXNQBU/8qqdtT5I9SHXhsA/uWQnjyqntPnnenQMN76PWNdC4PhTxd
qECU1DJ3fXy/YdWz5dtApV2fq6wbaYIYP3w7Hi3VjjIAwwRFBiiHdrPP0preiezb
GJjKThkg+VmmxDJC1DcUPfR5FhI+QXzpL34YWysYJ8WlhNNWn7jhmATpmf0UBSTm
Yi2aXenQ8Jls4kYyhiyXIb7ovcodjN6DiEKqby1Wg5riErR5enHTRpRBOSCjEX6V
TlfTvgeKousgdxgeBVu9SUbhH/zA7GYg6YWy3yZhZ32bL5idpe7hkvUd3VRPbFLZ
Rx7wOVnzMmvXlwG+uBDXP5BSSXth08bZBrZsQkSAcr/APoS5NFa7ShxUTn9yLiXa
ssuDNWAzddoaXRywW6+GD/2xPKa6Dhjgkudnq53Yge3J1iQdqDuT9JifDldM5Loy
k4xDAXIKkhe4ElXxfSbEMFAbVovohWAFoHq5WEhGhk1JsA1VqKaIdgg7y5orD8Z6
yK4Pq625Ee3eJBpSEhA4KkXplhS1vlQVt6oSyCKq8tyw0hIqzF9NlmIAxelY2I0e
Rrfv1twwFkJgNMOgmLEXpq4NfvOGgva+E3PoYWHrw7hWKt1y+Vk9rjUFERLf5d86
G3D407cKOK0fdWlqIlbCWfOhXvD0CWtzh2pnure+33rXHvpI1P5f/pHA/vOfIRGP
`protect END_PROTECTED
