`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vW+7KQTd3h8wdjf+7BoRJO7Dt8LKajr6TVldq/k4wCt1l1tiTI6F8EibiYIbnOsm
Ljd2ZiFD4zX8abrW38kDcXk7/5wD85KZTdZRDz56wg0BEy8la7NIPHSA24apH1JE
rpSR1CQKR+pHO5xAE1EllEHI3Xttshq7LqIztlpU0beXX9i20kMA1OXe2Kil+qgX
Pqj0QS3/1VVC2nY9f/vzCvWJZpaaIQpaP5zu1CG77xlXvxa677qEdRawNAt0kyTU
YoR4N1zrwGen08UG+GCw3wVOJjBM9ZZ8evU6DSRnle4hxV440UrGW+AFC4ETSmRK
da+z3Ilevrkxu/HUME8UkZEOEc8XKppXVpEd7uDAKD+QOAO/aQG5ZjCm3lzKupq2
jwEaIZAY6ZV6LuaAl95mS5raaSwkkTIN4CcZFA0KFLNglABlnPub/5hV+SodCXGO
wTQ8E39ukzkcT9rezLDQsAxyywVh5qIs5PDNLtoxW+cB2foFu7dJ4iJhoy4f52Wz
j7aq0zNByc7II+q+zooj50u0MPnkoPPXxJ2VS8GBDHzZkPAu2Idhh6QR+7Kgh/At
fphVqynRbfpuu219ZUDMCb1Oa5i7yeDdcgrhslMtkIspUUy7fQL0X6B1wCXplleQ
kxvFgGAVjhXuRF/SGoLNctPF8tmViSUQN18hg6nQsCXnpSFJaQXI6hG+eQonnGM6
c4aG6XmovEJk8+cWqu9d4/4TWgxyiZeEAWcaG+cjj/y2s5qoqxPJ5Bax2O5yF7L/
jCuZSeKn1wczsDQn0dDIqlZ05qfwF4BgaDalgDMGoMBWw8adZ0UzJ+ZJQmNaSvSX
7knpaYQoajjaISv9a/6Om87anQm3EeQEc5q3Du4rNBr4jtgwQyzFjC3AuA+LoAfb
bBBwptpiDcXt8TBjirdq14YU7wF0bdg8c6RKc67ihGImuC2ZyD2h0W4ZmxweUMoc
LtcO39VBm7E1DevPdGg8pRsSS9nFUIB94JWaURcjDurVmab3XofGQqach4xh9XeX
zmYlMIs4syptSKmqJQqPnwwwe6GI4/Vb6EFQb/CQN9ljElar36NDDBXXSAzfwi/n
AaGd6R6HpMAX5pIKWUISystWvzY5+KnG2SeU/Rq3r8elsgMk24FDx1PKwF+JbLNn
0rrT2U2DX3tVSmo7Ut9Febd/5U6JSdfkHZNqdx+hmatSqzmZtlSgiEGLGLKM01lI
/kvZLXxPqmSAGXe2PLrm+uwI3H2h6llWsRBttuQviSAPIHXsSexj6ZgahO1XYZop
lQicnRYU7W47ZcInO3CBkG8Tdbv37CCZmlZsnuIFEyfh9KCVtNhVGOUFRlgAkn5C
Ah5hWUfMttBgXTFbTF041UfGqVrOv6HsZoxUrDYbHWcR35+VzzOCC1n0TOm8QUGi
Xzk68zO12+A4LHHW4apwQsqr+e97kjJCLt/KQQj2QS1g2ReENbFaq9mPICM6OULm
NPrfxet+6cM+lD6PGqA8ansBGH0UVa6VCmI4B0/52ON3GDeLVL03G+AKvh9Fskiq
NeTSl01p/tKjr2Xl9rTkZWijAQoYKA4EI/e9DJcX0Yo6ff6MjYVz5eWzN7+i5yPL
5SZLxFEYyfDzSndFP550CVSRRMnXi6GX8cA5a5BJUT25sZtgnSyiB/IUPdcTGTLM
4vGCDXCq0i1FRcfrw27VK0yCOQXveM+mK0Hfulwd21AcTrxn+Se37dA5pWWgLkPD
W8koUQMOqOB8gTfN7FUZNNRijIDizU3E49l+wSpmpI92RtzW/dy5WD1goGhMQ8hp
8aZCrmBk/YAAfboir8QMwKkxYzZ6UNNID1MpjsO6LkjRnHBWF4g/rdH71kTxmfrh
pS7AynDhrg0KxpYworoenRYfji6ResapX55MCg/+6UiFeB0D8feXx9uuuhJG9RYW
9Gw2+i3Sh7h5Qsru1slmxcUiY4pK7kjVIeBHpONrH2NAYVpoMhdcfl6u1zbQ5D9m
qIjL/6SGtCNy8YUeG2U6TdW7DrZOrXo8AM/7rYA0c8qLadLSlg3Hh/vHnoQBeDok
oXva3Ubs6qLQ63Nhggg/DZ+QnOmPGAkasuxpLtMf3MAk136+n+yuWLVs8TGboD/l
BJwxj5Hvk1SKLEotiOfQfw4fZeyqocphEu+TKSJWfTg864cfQXcmqGALptcv714K
iEg83JiulbYyJG3sR2JRX7bmM3RiaCjKoCNfgv+Lrm2HdSChLIh6UOzmwJykzFVp
s5/SwquYVMrVGUlkyKlnlOhulyeR4I5izCEEieiIgxR1GCEnyJ24r8lTGyVgR02d
rKCZrDYmIBAQFzC5SE9w7XpayLNlOfosqZrl3oiJ9hsVIEUIQq5KpRl6T/2M2W1i
C8ZbplNQ5sxBcWymr95z7eOZ6uHs4tmKf7wxdlTCLukgPGDh2Ef5QvBWToAIqjk3
U6amrlU1e+JdKRL6xKauSEiYCSKKI3d0J6Kho5i4rGVyKuRa6VlApeDtLOmV205G
34aSC34UECRZ+lvPX4qF52auRPzrEgq1+qZjOKmYAKuE32EAKev7561UYoSMGBEX
qOD/PdzuS2Xb7dmHCmZliiM/JwVaGrhuHCd6QQERfatqXMg77XulXAi9j0QGCcvt
5hoM09DQYaJ65ZZYQ1RrpH3t3JTVUE3X7drWmyFzBf9Bv1CaESlHsk0U+HMo709h
4BjjbOwk4oCCSGvdYJkzHscO9vdpf8ZBhtkuKVSJW0ELNH0OZIs9NIZ0K4EEChi6
9na5aqM+9Vddj11aVpVvy8g6gQvy8CqhzUkLauwsHlHsZmSus1BydTIOWpORj81P
q9rhkfYZcTNgxlRRA0ziQdKv0f4X0N4MuUVHSuv0EDByF7Vhhg/Yb+1UQ9GQ3iz1
kgkM9p+I8eADkBzyyKsLm3EeJCXkZG7k8ZZzwbpGnaEYKFx/+6iBw8S+lRFFP63t
qP/0/xEgyIO2Y9ZanJa9Z3jSQLPlMKlAU2Ge5Md+IiXDavv8nMou1JpILgMB7UuF
SNOz0LyYeb3GOXiMaJcx/DAnWN3CMBF1MWfOpYsyBnfruyar+zFfx4V8D2NNZ04P
fsWiUfDv02Rxi+XO/DJ3VnZTGwsG5m6o/4QQ1nPCcJZbGZeRbhtS4GmbxAl2yzYj
hxSi1deFWNe3qy+vA47Vy7o0XuTT8OO8fhLw75H1Kz55pMR24AFnW6bO2eyu0OOr
MXZ2A9yqH0dVFpncomxFI2aM2bijPgqyhFidpqB+8V6+klex5ZP18/849E0n0cEV
WtTibkFCC596D//2hIJ2jFDQ4TfAxFw5FHRQLdTsP5dzFbOdmJPI0+HDOeCQc3kl
tPNCYmhA/ruNCZRC7qf0yD8xWqkcMl6vPSX6RCJXocKqTMSLH6+fRD8xhXDBh9KL
1Wzmrc2hmtoMH1Q7NSFqoS8cBnMh25Zt5HOKKZ7vWQx7u6r8yy4beDyIG/4KmKPy
OBITqB+Ani9VoMTP0RSELeZ8WJk3tnW/cPl/4ENzoqkpS+Y0do62iz0QnpZd4n5/
7MgnI6XKmv5vUkIOGzEuqHHcNpOfDN3m+qq9RAF3UTV3KiPNHFE+qsdNowmpcESv
0cw5ZPO90lFymYZjE4e42MYSJmjLjg8pHl8xr0iraIqs0mO9b35tzkVgh8IFtFd+
rFg4+oFdbkkd4NPUN5O9NMhdJk7a4BtYL2fvp3XvqHRoB5wXZLXv2x2zP9kG7ozE
fvA4r4j8livs7HF9VgXrfViUFcR3nU+7eA15H4dW+qRhfUToYYki3bVoycuUbVR5
eCEL8Mn5KaG9S3DbD9NjJx5qMcASPp1/6EDVI/4r3vJ05GYXDybb6Q5bbWt5pjwY
9CdLwHXpo+QKsKA/Q7iEe8tCtPVBgzYP7bIqs3WTT0L/5rFWs5Y3Uf8RhpQVK9fc
c23BIYObdQBBXqqmtFgGV/vOTYL57Y96A09w8mCJS5czv6CHeKJ8blWXhCsVs9+p
/MExGgC9cJVIBYde/ZXm8UyJZAY8HAHN9SMhskpx3l5euIBcPunTSDR7+gDDyngD
v3Yft6zjpZVbiBT8IB/s+MnGgdy7KZVtM7hnAM4VLZoPHInGWhy/4SPxKq9Nd0pS
hcHdxr0XnRM0932HVQfw3RBH5L+0/EBL0URTh+UJbHhYt7zJvC9GJ1I+BAMVGONt
C2bZ+yJTza5h6TXrP3PfY0ncih8+aufA26ul2AvRhRyXgOR6JZMUS1X+vByq1j/4
buVkC/1T8TEM9jGVFxqayS5uaFT/Us61YidCYUUT6OiyP6m93qFQwX0YvWsPMqOm
/mzTmcFGkkntSU5qo8D0QFWnYMlehJMRRFiVWhdm2kkqL6c7R3jyMsaBPYE9hoj6
thPxXPLJCKZXnbaGnL93GQsK3qWUUg2o3Pfs/tlWYb6AT3MhgTT/iKk6RCPgkuKc
xWxCQvfdVEduRjJVqplZS6jIbTcP3dGb90c4H7adDY8AL6MiMDtPtSmghV/Z0zoK
gdGj6/1jBRNhrT+JrnBk8BEczHOkbCR4RuYOZtZZQuV5ZpGv47/Jc8W/itnHvM8H
SVYS8lW4Ez5BRU6Bm6jm8pP5UkGKpYqGWZE+UR+TJKgsBzAFZaWX2O8MCoEZ0XbN
K05BOOqNWFRCpgC8VYenrgkRLqRVroXNm1OgpsX5cYjMHniJH36secIJBntvfAcY
2Hjw/glsRzCze+L3zF8no6ojc0pI5zpKCAaIw9c3tdTEQRJFQGgoIDiMmC8/9yXS
52TfGsRs4DmZjpHl0MiKnYwoo33hkA42OmvznwvayeEzU2rTnhoMk7mfKpcNCpd8
Hu1Qnho253K0qKcf6hT240WTzDS6IyBjY/vfqz8sAdc0zv6VmHvZJOd2bpRyz0Y0
4p/jxEjNRtvRHaCeQvd0Xt70cR1DZm+Ohbvynce+6ecdkbpp5voraNg827cyvdhB
ct9snx9CMpsimvyG/LaqUpVF3lmbl471O4rALKygDj6MyHoB1+uhjI/XgVlAF3cu
c1uUb89ec1oRb0XZb7QmK6DxxPOxWlG46zA68f9TMIWwNTmp4bHx+gWfiT9RaSDV
DWD9afM5QZZnF3lI/+wqI3RWKLJcTR8eTMX93n7O8+L4MVNGj+w2rbUtSVylW6W5
HoAWTH3IkPs0DtiTxjwEQlKV8u3J7qt3SwvVv6aAxCycJTOGDe2iwfUQu4AB5rVf
3enqUMo/VVRAo5fcp5afgUYwwjsLIbn+1So/A1XrOdfKBlV41ftb6AFmk+Vnc+Nz
IXULL2NazpMwg2C7mfuJba+Rnx1A8kiPPEp8+du3Md1fe1wcuj2YsylQS/oNN6z/
7v6InvMtt95tkTLyzmsGuVBfOVwyQ4pmDPn7BNHm4ChpDKtjfUC3aV3vd6Te9+f4
KOiiXOEcHeZVi9hnJS7gaa1aVnPmaDnVUiiiRcK/UiASAB0elpByf/bhpNiVyeWp
GUe9Tg910RywwvP0EMl+V4XrNtnIDdymZF2HmOq4YdbC/UY3XCU45XuUBqkj6rzA
jD12BUMeFuiNQRXpYVDkJ83Nh7TFVnCu9kAqwUOGHPWFaBgNkFwI+0FszryzTCsf
beYsKTcF8trcwc9X3TMXmwetx1DiY6pbADbMVqLz0m6fx/SMgvKWAfaLR79fWSfj
nYchs1cHFTYT8WBqp9R7MrzfkcoNgN//yAVrIsodHGUfIfqiv232uERqBuCciN1X
7qAPJ5U7spM8xAKHb73yHthsqZ9o1kyb8sbqKnKBWTJpm2c1vkrdFVDi4PicmFGi
Oz5lU3RgWo2sJcb4V1rbb/5Gl8tM6QGSsGZykTxjvkwSTcUcRdx4xMcvYkemLvgQ
9ru2Xk25bjwsh2DfSJlur+rSh6hVmVF2fQVhkKwKRCxcwk7dkxyO9PrUcbzs1ujG
9S0f2URLE7UXmo9B8k986Kxn+ZjbAvjrIU3T+GIM1cL+m2+2DorEjB7BzMII1l4J
ON3Brf8p8CJYHsYHqJ/jbjrHnrVbolszD1kFqRN2Q87RgSm2vNi7ho8ThuNy9Vfy
uevCH0qqYupL8cvAhZtcnb3SnPG7C13TipQo3TjIJ5pnvFUQemJUZvmW8yL246HM
cgSDr5o4NqkGpQK82QtPf1cVpJLPMmzU72HDMXvUg9thk4CRWZC2jRrctAgNQNqg
IUNIPI53v0XDvy5o6sgGo5DGp+BDA5/cexmM3hyBn2lX4wC9DmbGvJYKAOkrPdBz
K0CeQ7OOAT0KTtzizLAQ3VgvvvyfX0gOdoSPErGVQh7eiwinTzPqBxtranLvCvot
ulIEv3Zeda/jAH6Gqcl1u+Nw4JnX6xFZofOGTodKd/PyZHAR5XbhfV3XaKFHpgH2
X2svNhoo0uBCRHHWa4K3r+E1D2SbJFJO/AYW5U0UYRJOqyOYJKh/k75b0Y8QYVq+
rrhV7z1RD/ZtWEVsWuGzgWAvvqT+QETqK1bLiPtVmRs92jfwQkW778QXSnzZCfig
0IIMKUvmlxCCTSW0RYgD7PW5b+3fxAjiY4+d8qcW0yGSoouF8uIZ6EZilYK1Jorq
B74gQMDB9mF1kNxpnCGVE4l9QQw0MbsMIkkRM3yP1hC3amUbHJfcPZbQhpwq6ncP
z12HYXlgj1/MvtL//D6SYjJsfgiUgoBG38JpmBiuuT3zIdB80hVD3YaV91877Bue
wwNkwED5dxifbR5QPAxq2HUVb5BmGJXNVdQQvkjCHP2IMA2uEyiske387TX9vBvF
wcrmLYuqQJYswFtKH7PCEWVHjv1PBJ8oy2vsewT6tz8yagSuzNiPoeGfBZFkY3Cl
HQpIDiXzofPBe80Knm7aAWTgZdwScorpbCEdJgMLC0tnaqHg4kwFAn68DXTcBtZ2
fvqdAOPNRPLsuZJKmLj4iZWEwhdCDBRRH4Hv3nLIQqr7x5tNdR/XWA2Fhqk5VHNR
6pRjbZyU2K44MP8HWO8lWHS9IuDMmbCNx9yXREYCymmEe5IqnEBA6oC+1o/sDdYy
58VXYEc5SZ6/XpjW+3rSwQmYqIy11CERfEc+66beGs4tmdu4DeVu5WTNM8DE3isq
kizJd42ecks/TIzwXTez1wauHdOJ7DPfiT5GpjW50oy/mQ4sCnX6wk6Wp5TO/WAR
xsJz1meTBQrhidhREU6jbaySDHffePfEZDwdrSSWR/vqWO1sXMAwkhbCNDU3MJbA
AipebDMgM1pXI/HBzZet/pnnAFpfzQ8KPpYEwu/01VfQfDJkLuUjG4QzX41Zkw6m
IMw8JMpshF62PkXGCMtlLrauo6F0euM3nHu3sK0mEX1WvRxfU2c457zWnQb9jjhb
vSZQc1KYPt+M+h8tNpDYcdjAUkAXV4E3fWqC1BoLY/apPs7QzYPrzpkkKolM+Vpu
9VHDdg7H7nLfQsB6cg8W95kV6g2bFDLYD/7agv/QgCWpHiHHYv5hbqct4cgtVJqK
l8ENnctJyuYhELP87JG6A0g5wA7/032bLgx0qu5oSZmJr8KdzoAb+Qef5akGRwCC
B6TxD3H0uJ3QAk3Np3CTBNz4sISClL3l8tijVVQoMKKQxTh6ETU5SSAwAtiVX9H2
3ThT68GjdXcO0b/m/K97QCNt0FglAjMgf+11X3fqJ/e9wsd+HsOABG/IziNdsvLn
Yk62HW5G2UdDYLTRke8rCfUnNxiN8xMdR+ZR2TTfXzYAU0smK5FZvIhNqpzWiJI6
QAcKoLqnlfZN3mbfJKIqTpAQ7vVrttuqSEz1fCIN6PEGrmQZ4j7bSs9BRbAIS4Vs
BdaiPnpYZhM4PnheDqFjta4QpIYzDVspB+wEaiSxy+dqcyG/hYHBsxpg3+AgZbQy
ZRXb7SH9XX7Ecyep2w8cKrSy77WJvPxZ4vM3pG5Fv8igrfu2AWuLvBnysLEfedrt
pEwVK6WlSuSEEn5rS0brNlCjARQljJmi4gH48p+qD/8f/+AAxpzIe6Dx+tL2CcQp
/+/TSqDQ+G/TYuCK0qqVfzxKxcTG/ojVSm5kZGOOolmQtEtXe7POd2H5q2xvrCU0
ZBhuBolfhxlILUpIUrjxA65DJC2Tk7yHsg6h5bf1OuILKwFSQnTppjOXP96xYS9j
fKgkTKOcBtXOA9IMWVxvbul9OsdFpA7eNb7gjh7vTBw1AZdY1lBjwhpBQ3z2mKut
brKRyR+fTSN2ZrUSfJxdBd1SAImU5S3f9Pm4JtUAfPV0NxTM71eHBfGacpRYciAo
KjAjFm/KMM8EbaRaC1NBksF6C8gDX9/JhCIoTTXJMhjQh+sSMFSo+ZL0/Oyuo/LO
hJU0LnsXwxJhzSVUD1k4jEmdt67gHcqEDHRvRpI0GKAZW5vG2DNXgOle3CFoVsLm
lT5lCRoQsNvSA96YBxrprLAo0kinhuhm63eO771iJJ9PDSGSiWMlXrkjqmXAnIbl
bimqK8cAL/TpSMPg56usClAEZ/wv/2tV+ABIASK+q1VPx2FdB1TYrI7EAWeqIlqC
z4wgnYn/okZuXThdlNWPCBMhZ0dkGSSU1kbtI/vGbrrxOeam4T2qxuqeFTp+4S+N
cQA4Uez76WCPK0/Qkt3zzObRr1YH7cgAxp6rF3SpFWTW96WJMbL+OQIxh08vMgBF
3Wwx7AafxIPS7vTij3S3T52/aGxdE6KdzG/DaU5wu/dNZgjSwmorTr+JrdRTpZoc
NQdcYWPni7piHcXh5CCl1UCAdv+78suBIO3+F7lOfy05lx+E13Ry4F7A51h47sGI
50w+9E0/rVcYABItb5lU/peXck4W0BulfkU2rI1DKPgIdE593EGQmurL0+UpX3HW
A+8j6/TqR3CpSRn2cSxRA69m8xjY5toks0SayVBfTDyvk9Wh8eCMv3Vhi2J30nkS
yZeu8kMgg6R1zdz8UUXboPUNtNyiEVY03icD7hSctqEN09UEfB93vW4s10RI2uz/
omMPfzN01oeM4AuQqT6tYBV4C2wUhUSWh3A4NSEOdC7956Km3H9xQHMD6Ekb/QjK
zhW+dV1AqiSep20BGtqZ4k7x4H8eB1bFOhIXp6dpz+IduEHOir54mPjT+Bc8GEEa
GPBqgzccMuNGQk9d6/0TMfChqshx8IfnDybOjijyzQNt/dJ0ulcJCOmbbSL1zlU9
QeDZTAm1XqU9/AupOc7PHWzJmXUK9c5mglynpi9Ggj46mmePzi7Tsak9AE9nNdwj
aP7oretUkkezIf78CXQv8ovcDmTEii1LsJb02ZCOhMqWBCG3IpQAjoYCRjyRAkM7
mk1wisxbpkTLcLjMW9ZM6KEkJJWFHKXFIHKtu8VZskPELdwjbp5n1gzscMFUckif
3IKOMty4dfpPBio7yT9hPsBzdi6VOWjG0OZ/V6HNme2BIU2TWoBVI2EaGHaZiYAV
jRu6ZmIBMNU1zMJgIRk/CfH02U+eOwLssREziZqqeiRzmn8a/+VcWMF5pi0SU23L
AiYbdKZBeCCqmn4XC6E8IKGQfHHZkCti4GfIvugEo5zKfxht8x/x+5cKjIq9PrX1
922mxO/wjxksA52scWVqdCAN6gtXjpERLZixhvhP48Z0lMpivmeOJ5hsBee3aSmU
dS6S0Gb2DufPNo7f4EjrlIG5/MtS2c0HuKpl2QVxAqT2DY45BGHP9DDLF+D3EB13
/YgK3ZCjNTJ5ueybSn+i30OkrlgtNe7+dzchlLedGjKwBIVl2qN56a4bbu8x9yEX
42asEhbpWurvhMDcQoZtQNOiyl6v1yovXnOwt7+kmUlyoV7e8ZeMT6LnBlUCgG1W
JLFm+9oQXmfA5WbEncuARMv8jP1067QBR/3x3yk0D/7YswVBoumi8tmKQxJm/2cS
1B8jTT7oNBXVVKLVouuk9JsIpn+wqIOPt8kbrYGN4i39xV2o7kelA6RYeIelLlJw
K2tUvsA/+E5ONFMV/XoMsGHuoqM41Y2R4qHMCg0hs815ELi+QqCoN+A+Por11w6r
a7wbEfMYG0pu+l0mP/u8m9d2DeFlA1R6Rnrv0cyHASOQoFKQnCt3uHPPru/aYcIG
K8asWC+1iBF42/eUGuIrktVchDTR2kf46eafyXSYUY82gExvRuijeM3lEIsrsXFT
MyVBZEX0CcSgLGTPQadDAnXqpAJySWuRGP4HCqTuJ35Q2tX3opRp2+Jaaft5t9Us
CNjKIKjg2gY2EZOtDOO3yEdEgL+6M/498XCLOmVkZluCPbfFxRzAtjuUR1Mv6DAZ
EqImVvz7tvfh+9yM1ac2II4fC2+019PD/P4yK149qLPLlVhPckawHjuA5cU9QFBZ
o0P0LN3rze7gkf15fAJbafs1NsTeE0+2lM8FpZZsjCDM5guxSpioErKsiqWzcWYA
WPMSk8X2sQYRbROwO2cksJJ2c/KIRUmD6M05s/G2kCM5sxrU3jK388lHFNN/DWM0
dW388jdR1684sFRcCUqockQbbiD80ic0IxLEWhEoB977FgA5svizEU9M2+QaoUJN
zjpKcuMb9nPac/io+8ckpo31lJhnneDgi3z7s5BaU09OCo+5PuCIO+QGG6tdw8rJ
HbwPbgSf6DCR9XPwYRRKctQaAzo3Eszda37O8Dq0srK0CpRNLDPXsP2E2FMvumPm
+oPE7ILEqatRWAcvB7/KjIC8ayyeEAyEiz5GGX5/ItA/uUIb3+qyJXe1icnpLfqh
XGv2oFz+XroJ6Psy0pi/DWvlvNlZ8TXwxGFHeQvd3eraiuX0Lgm8uFEqcE8RzWiU
qhH8n8XfdvGXIwdT7ZfXY18Lt3WjLtB2eM0gGbYAjLDGJcj3WCDIJVmZ/l5RrKqZ
5aacPbvr0yKZ69UDp5g8uYVbqOeKPMPIFT4Jvo0LPfbdGGMEjsqvtdUDJSHNYope
dDUFYZiukYCQvOYj3baaLuVHVZ7IMdaatZ5tLrxjmN/OXA+U8qjshquSF11Oi4NG
Snc82qogoyvtT3P2ArOzNFQs75V4GLjd6ugv2I/N/DtHXJ7NU1tN7zzlB6J5KTJ3
2GPdiWnG3INp3cQSYpQz0cge3qKtOU5RJ3Z+GvY9nXpExC59cf5XqEblOrSpa0Ea
74iomcnyB1UH1YcjxgH6gy82xA+7CSuvb/mqDx/q79zPRFaJCZCyCOhwkXojez5C
jsN1nxsVMnJXlKOW8XZpoui+H7oFPnKMMpGikMAwwTh4oBzUncmtMSevanHMOpDD
CGw85UG5zzH6B70us/LSM3Qzh0mqFz4AUrA5ODPa/QUYFwiBTnaXrOWG5fX6uF7S
+oOSKJLXnEqlQzBEvbYsQPbHMCAgRwhoor3d2ZKngkGqSZTFVRuWfFxKq7RTu95o
Q+XnQa3MW7NLX4G0831CRYBLB2oZZRqIW8fDuwoNijQJhf6oFGRjm7CZBelhD31K
4c/IxaCbJ84j1/iHTBV9u1LbA5MyplJoAEk/RSwVrGVGXWhM7JTWgwO3QikxjLrI
4KDY7XVSCga7ozAb24B9jZ+ZUG5CHHYh+zPErVL42hPgDt4CGBBOzW7itxQ8B+sS
wSN+zPHRtAX/yMYh2yXnyFLyB3uKjg0Z8kIqCRnADiLiIE8V3WlMWyn60Aolvn7Q
YSa/nvDETDoYhCuDTNBxTWTp2NthUK17F6Tfp0UPToYwljLT53zG/2VmSL1lZfro
YpTk1i6QkvwQFEv7ywJ/2mV5InuBP2G1+1tLtvHUjtfJ+87gpwakst5hmVQEDKiv
QnjkwXdB5ttQN+8lydvhnERxQeDSUkNhSeYs+JfckqMTg7UvsDQK0pnMViezxWbl
IVXJbt8NUgGKcC0OxVlkxi/7vKtdF+IIIsweptgrkKjt0V4X6ujjRxfQ4uPuGJP9
a5VIHiRqu2dvnD2L4tnijXHANeMGnGR9xy5zzQwJdsBVMIxGkczcDD3V/ZVgvXMU
JBfE8spcjvjkPSBjJbj0zveln8gf0VvhmiIvQejV0Xs1r+Uy3AylfdLCSh+XYNF0
9AFSpglhm90d1IiWKQAt3wpwKdBzqfNUoUCcFaQBAzvu1ACpDvvZGsMf31xlnvPt
1MUiSEmp+qfkMrgKjqjfftdbwVp1jVEoj8nRbeHp6FshNEvllX2SfQjehvKTSpmd
VHbeOaR61ru/W5Q9ooBfgEvurazHXf/X9MI05TgIhl0YYlRdGiegcAS3ufsMlFxT
kRfVGDDJ/oGvvuNDl4ZaNIEF9obpw0dre9vntKSlQt0mEuU9gJQCgo1L5n+ivPF6
MkwFkCyckJW4uUNqmAycTHC8IXC3ao+lsI7ng2D2VXwYHkNFQKaheDYxAZ8GkVBB
gUx4eJ80MfykLpZfYjzP/S3LX3wonsQeNckytEL/ZWbHf52qvbdmNGnNSd+GVRa8
j4saMj99PEGEKs83EcTLBNdKbiUeWpAI/koJ8a4jE2G2+aCkOg1kD4mguh2cxUvF
NUdAjPVFmGeBI0Gb1gxdHsczk7Gr5vsHF+sINU+ah08IaK8YcZJX/mzAqwDedh01
ahR2xxt+bkYE2ZDVxPjfJgYQFIlnnaxSGnf71ue4XbjPjm0iet/ESeQWDKPydovV
7ad+bo6odKCSw+O/bcYc6w==
`protect END_PROTECTED
