`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZK4wJitoMWcZNNr4nFiS7YCDt+6RDQrh0QomC+XtMcurB2LsSDheFc32KM76+9uZ
YVmTTNzAhGlnlBrlEUNGDa/vcR0Un6m5uBsoSTT6qhO8rrDJ12K4QDo+EGTpeZcc
IR+u1vgF8yDeotIa+mpM8yuWeRRW0sra5mLVsTf4e+SeRrnKu2s+NlDogNInl4fw
nnAHdij4t2qdXZGMyTY0bUFLGMdn6++YHHDLBjx2rvuIPygyaF3U8Q8vNkhUqiMQ
fDyhzJUa07OtTArpZpqvfbD2rYVTGcfPkRzmT/WMB5Ere54ms8wGNDARWIe3ob+V
p8i2MmlSCcOs1neKXnIHuinQ85Oyvk3UJhRa+AeHrNKiRWGCKFNmewDRZ/y18+cs
mb0P6ByrhXNp+S2k8Ce4OH1+pkpTYZVjn1dJ5gVH2fdiaGfPtp9/oh4YQVKDr+11
jDpbj+Xf0g1fZ5l+s9/n0MvuMyv6w5IvaUSkWxNWeQMnTbmwf/+LFXqA4JFsIuTW
RcDvC92K3VI57W/fB59HclxEsznPySpPOp5G+XUR9BgwA2sfUAb0zdKHm0MuQvS8
yfanbAH5ZfV0215kdc22KUDasi8jC6LUdpHIY5YsbFtOwufIDMJbWfg0bCXIDHSG
5eCMtbNvSzzWPzPfqQj91F04SA4XWbKzDzpJz6mdVHUEyl59A/4v4bieuemDvruY
Plv+K7MwFzmc6VIhKfhfP5Up6gkbJBNwAFjaAA9fh0X0K/a9+ZrSD7TClVqgAPrp
FGjubr3YggvfT18t0l5wxyFb0UysW1T3gN/z/Wr8bQjcN9otGNVO0kZWOJPITHDt
sF7D3zIBQRnymOHHno5MIhQluPcTorQbR1qv1q6Jl0bSccOoZDhNh/wrygqcuhsW
IrEOlvW4CQfflFwwE4vYFWSom7jw8spu3gQWtZ6JH7w8sIEt5hJQijdXKaaYEJW+
qG+fH3rFn2mT73aVj1wFXM9FnzdKt09IOLGC+fR8JM0So8MMIgvyr/m0WATJBzPt
oNLEo3AZp7XwB84edAbTTo7d6ShmreZytDl8KzCsc1OCk9siEcPfktsK5+3/7kyc
6J0xBvQOa5DnZPloJ/vUoA39yaQJ1VjmYKXhgHd4zSr/yetYuGwwN2DUQdVLe91Y
V2gOu6GWtYzSiA7jyoE6eimH6xuxF+pktwl45ldhz1DhkAXjSyH7ARWGtzo8DX3Z
3CmxxTewPoCvHEoKLE65l1xqYCY/F43Nu7BQWYmDPGsa02YyRv0cgxayoUdxBSuH
Kcg7Du3dubxKI3yFwxcsOomleQhDVJXmgS0POUt/ruNS9vlx8Xa9xL+sJBl8DObQ
3adND4nHaWbBtkSGdsfuvm7vU060/Z092cl2tYmDY1S8HzTqBiTj3RbCelSlWifU
JZC9EAMbnTJ1b04Xk7/v2fb9DHIZUWwVxB13bVqySqx/zGCR+r/iGBmYPIPvb9Z3
acroOh0WKG75dhHtYv5jfEsS/RCzccirGBQdG4RFw4QVy96JbblNqs/OSkVaP3/K
kLxtX7VYICZqUf+vpPvkjfKFWnZxKntAbkta12uMXnfNTAIrRpeiJnC14P+FbEtr
kXXfpX5ttNzltY/suxaTb9SU0wfTd1l/TijFnH67nhREv0Nu5FX4C1kjx4Qud1HO
BNoYEb7aYtaYqQQnfFlGWUhr49y1Q/V28yXMUxapX/TBwU8HgrlyLzgN6KRMh7ll
Vsvj0F0ZrKgVY+j/1zxw+DoSI9kDfk5tlRu0b/YLQEzvyRcK6d+tbxR359OWRACO
PaWKXYHu+JbBSBbEexPASmwC2Klce86pjfAvPrSinAbm9qjWZdPtPbY3e47KeIfD
UU8Zcz8NzaDw3c8nN1+pWiOM9Rj2l5Dhsd8OC6Qgx+EhZqRqTSLEfqPMxLWbBtzQ
QgDn+HBiRqhAdprG6Ji5+4EvnGPEFUH041eox9g/+q3YtY1IPgz1Zpd3i2YpYqp3
0HnraB6zu3XnUJTUsiTbrBABuhgo8FG+3blhATNOg67pA/wAOpnoTslkIqcrV17Z
eCNFMEKqmwmI2YiDgj7VNlPoNsBmC6vUpe8X+oIExrH/QNybiPFv4d/0EnKhHUFI
31pP57foef/CtUd8Zn8XPR0orO/41FHZxSQuo4damNfPCQORMA98J3gigoz+Nymj
F1XkfKpugv9vQOZkOvvy8/4RT5haR1Om1eZ0pib94a7bSSVRTxMaZdFvuYnGiYau
fX83kiKjAZcrpclZkbXk8TvLEaoMEPc3AnoAElSkBq7o0cyrE2itWU/8rqXalIR4
s7Bcr88b1tMwgMJHbqVEIGjnmxs0/8Ca+Y2XJVu1RtGTd4vJ3KV9+76MVgAyiy23
fwL6XV/F3rpd2sbDCKYhKcxy+0Lh6FbB8I6I1oauxRByvS44JskV7FV6+B1mCKmO
RMv0EYnvfhSI8Sxn3BOJJr4MXHrH+h3vBjXoUzc2ArCe0WIFfi5bHihi0Wh0LnYA
G8gokqTbgBoWmeqXqi3MhRmXM6c6RCLtgWuwO1F50VNmkk2UoILzyQwe2TVkzX+l
cRxQeUNoMs9iJ5/NbRQdv7Mvq2ko5+7xYEo60u5tMgzVNGXpDOKkylwhBe3Hcd/o
87n0QVo8283e7zBDB24npAgNSjuuLDiSNSupMHi4SQEnJwzG3ojfLmusoPy/QGtr
Md47BB4dlXchoIYj5PJQu/JjeExOjvM7HNXzX0BaiuQr3ODsmpSfmh45RlfPkK7o
O8nDECwG8Pr/Q/gmMY4CSH656GgV9yv+g3XfGMs150s6sFe+/h5ZKPeGtWVF40kZ
EMv6jox1npc25gk31FII48lwjrGhQHWsg9Uuhumv7WQcrc2mZm+1gqMh1bFD8LLC
fZRAT3H+Fbo3fdZQu+/ZibfA+Diganjxx+FSFYXo5mKEQ61/BVit6n5xbVCGrjZ0
gu+t74EL97JpczCiWQnAnvMXXKmRKvjJlrXpWtqmjufeFNJJW6tfnjGKNASXxZWs
zjG6KEcyLhIFArXfLEp3yjPwPvPIbcjSeINXtvNk6/tofbvAh9Ii5/Kx2wqlaE5O
qo4pRdSCMbzeQY1+zut+a25fZurjeWMC14wfVuKnkcxsYYUlZHdZnhJqbCKaP6Rn
jKiMpyEJDH6SLn/eiaXre7heUpvBSHh0hDrYdAc8sajNUneNTHvBq6a6j2QrSTTE
tosdEEV1K6Pu7h0a1kyLGsAnCqPv80z+gpB9Jshh3xrh990Y2LHg56Yf/PrEpvk/
Sl9hD9/GHm0FHTfqMv/kpRl1+4BQ/F65QCxpdAtcOLNVO0Fo1daaBjF5TaPzEqaY
8MRLnPMvGgtxotz+bvod3pstUJHERrtOFXgflON/1Gq/WWhaP2qR8+BxmtnIn4VJ
`protect END_PROTECTED
