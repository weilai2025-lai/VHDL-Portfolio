`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JbPt1c98vPl94mT4GngHdldc3RURhoHkRs052U33zXlGBp4y3mg7+0uICbY3mEb
4L3tZLEJXmOngoo2S24DA2qPY0M1PP5ALFTTKE1TtM6ZEqVbZaDzWLf9Np/AsGn3
mw/a6yUPC4HyoReywxqrG8wVt7mTswucwdZcPyXpEju6Dk4gnwhq05G8kjq4ibY9
cKIfe8hoyFqwjdcnETc4xqUyFbzmCEl0FIpsvAiT2ek1890Cc6KBMwqCdXz3KC90
BGJp90B01F60nxWdczYaJ8TczwqMQr2l79y8hJjFF47WEo/iJpFSwHxtl4+II1Ho
UJYL+gDWdZ8ArLxC5q5ml5S7ZeEO/aycx1DJ6N/m00AtM/AuJE94zNoh1WGwz/SL
QLE4u5ZtqnyyBBKitncnv6mIuYvuVb5iIGgWf3H/DI0w8v3tQU28NyeqzpDqkKZ7
ZjTtNFVFhLl0TOmUHCwvExeqeYgtDJ/pUVpJjO+LqcmiDTjLmatoSSThEPh3q5Oz
lpDmUrLJzP9CzH3Avq4nLVxOCr4xRwn4NBP4idvzX1eLwd8qePCvVYW7hjilLRwH
bFOmrIHZ1KyoiNAKNdCgs/qSTgODkmNCFVpNjI6+MV02erQwKCjqCOy4swm6qN4F
OtB7HN5su/sCXV82kadrlYWBz2RQWu7GgBlviqgQC6ic147NJdeyzXpRy/ODa0ui
c3onvZ/3YmFXDgcoiXgL+hRsO7zUBklofdqL/tE2GcPwn0wCLVHd9mG15XL8wKan
YepRm7VYPX/dT3nxlU743OTNDL3QKFblV76SEITwZw62dBSsIK3zn5HiwcDaOXx0
YNhx+M7SWAySdL22MG9C5K+Gk3HfD0Q1TnX2YLi22yVjeLBQpCBsgqpOB0/H0L0c
1iKEUaGWdJEv6rxdJcPLisSZkmJ7DxRkXLWESwMse07S4/7WJAY5nRgEY17NzaWw
jmaR+GbjJGRum9VlURc1OJC4mn8xHYx6L0uUMNydxE56+pkI/ocddV4Y8P58Odwn
8B0IMgYzfvxWfkwxlE1ofH5Sx2Gmp60+DDDPzFXmHsWFsLRmwXyAG1U8yZgnQK8p
kO/wOw2WxVyDUyiwfnYztoE7HwEVL/paO0U9Y/ddBL7vIp9onM7/cvWarJSmEZLL
GR1dR4DiNtxPwVo1pQHp2rZvsh/l2VSEI4XZiyXxf7PUa4pn/Z9kNwllYKPE5n2n
qm0KEQLLlQxp49IlatIFklGEA8yav4fETcyCPG18DZSW7vlhC6qV1EBYRsukocgp
paDA7gmIthUahR2ukCTPsBO9XyAr5dfrheb+dfNcMa/qEyF/5r8Zy/oj01EhqN0B
twLfTb2CyeW6wayFwhSTGMo/IcA3HOKgnN8LMY1PEMEe7vHBZ+bgKjHXO3uCsCLT
UOrTxztE/7xlGGMBtj4iDB656zhP3IiqCbqD/mrXi+bysP3QhpgJIOQEfMH/3Rd/
5Bw8ii6aXu2wBuAjgwqrdp6CUA7q3hUGRuALJ7oyQEExVZ8z8PhUDvibN3G+ubDb
/koSKyTKZzj+rIoZ3MAP4EoGcAx+T6h1Q/3ci2XKIvj+J38ZnEFJ4hcBzUzX5rc+
mYT2XvzB11FhnnydKrCi63xZ3EPpt5H42qF4jzxmfRJa/eMyZ/RvIF4xWUw7qFMH
RFm1fVEPPQx78lfLaa35LP1jdtcVCiyP2ApWVH69w9A+bTflghaSgddg2UpJDrIW
5JyZPOsO/02Ry4HwIlzlqe4KhX9GCB2HDsSydBvtIYFjityRM+s7Hh/MLFjOvAfZ
aX6QrDo3+HbqPCuJR4hghjsUuLjUkvWz0M65cZ0GtKMV9v8Mzk6n43hJ4MzJj7/2
cyXZoF3FDjqLXiUq4g1ZzBALtxPB2vvHDbNZePi+dHvlcfeGtSS3nd/ABc/MS483
tpd8nvIotN7I6Ag0yrBZM8eC7qY+3g5MOwQVMv79l4o1rduuR1glebmfqLMnW9tr
HWzcSyIHqpg1yKakLAj9klkePbqnvVZgfCPwxd7zLJCXs+Xy+XBuaNXfgboQ7/Eb
zuPzdBj4migXtt3kCSfcRXhvWEQ3akZI+P5uDiLOjrylDnhHe0KxYHO7MkROYZtV
PgByDQAEfdANatSHchiO82q/xk6Cm/MN8smScbhTMnRfPhSCgnzGlUKw8+52eCCa
c0F2r/JJlJVtFIrxChWh73Uh+nZgNaocmRgn1yOXfAFz81FTyKAQlL4/PbpNFaTz
sLgBkRvlU1o8lhkUbbPpY+AzLUdnTmc0nDoGJMhyp/wUMbbYjWHp2hLg1yt+OsVc
2AB0aa6KkImXOCX97YthFDdnoyX3meS5u+pbX8e1qu3pYEJp05utk09llXiEGnJu
b35BTawU+rV5sxQhKuL0U9vEuETzfYXVajL9zWBeTry7A6ddMpA/bkEVWNyPPmV0
heFmcBXYec5t6gHI2ucd77VNHsjWScU4L6ijYFzkEgU9oYBJNu99AYaImDif/IBd
ZIuNDsAvaMyvw6qEm65ei8Vdzl4esEurDQrZq/uYB6H3OzJ6oBqxbXGXCNRSfjCc
g8cHtyNmWFaLwpOycralEBpNaDNTuwTrqeyHNHSW00RG/KbexZSh7kUNZoIFWYQy
ceVZCMl8IMlzC4KL9dF1WpecZMh8YJQEAWYmshOmt1B2Hs89v3AZrv6HlNtlCFpw
AkbK3452Z2K6HTeDXB+5fG1ezq4lcVbYqmfm8odhqcfM/IaIDGDoycNgejJqj4jk
Juz/5p+iGHGs+QcZTFJALlEvu2DAdDNzFrtujCOtRxfHgQZ2V3ygWlYaAwDawVp7
yR1YCyqo2IDrsqnDEQkjpgwIoAm1QeEqswOUMjG3Lbasl8UYArxP6YWhyjimn929
cyMb6wI9YP/XKyJE6hWIMnMWkdGSB/mAhc2vMV8v3QZqIyVFJgvGchNy85RKLJ7I
WxUKW4IULLZ6FYBnB5n6ZXHgmfB162ECltluU3lR+3PN3NL8NaM9hQtX/At2PbJh
K/aIUYDn1hoXnQV6sBanaubeFmEMFTyNE13MSlLNxn9ZObCsWrhbfUz+Smn7iXPQ
DxTATyHJoG+M31o6Y0yOe9OJI9PwEcNhFwvJEgLvU+uTUVrfHLKu7uNQyVZKUFiC
mAcnpqSEbww0a9LVWUiWCdpX9Rxg8XJgHwWjHQNxUxuJxVevxWs9jztFXXjrgVEp
zh15s73q6CpGKQX0eOYNwoHSFfJwBEwsWYAs4Lh5nyYM+9t3tI2HZcDUGUDOC/AH
U0oSR7PbMHwFKEDfLjIxh+tu3CHJiuxCXOfkhkToiJYVUVzZdVXeqx9Ul8onJvaB
ibDOmVM402KJmzM3q4lzpnbMTYTeyC5qCSrKfgIHHWCV9uHH+y0XyOHdvdPUaz4i
gr/b4dCiZDoBYQAmOEqh6pj+W0Ey5MiCWBD0qVH9E83MtcWbiHvATysmhL/OVS6P
yF2RcMAz/AhasGo6g8IqjHCeA0mypuLnW92OIlOqKYyUfBbfZ5qmdM+J6CN732W4
Cld5syz6ZjYwPqjoUdJvuN6VrCegYOZpLIMRhnbD507NbKSzPPvEzie8hpBeciBM
rKTOozxpVucZD3DwsaMrmAPk5W4KME2n3mBaG5MDBc8Vz4bwrxAIxV1B0nF+SiSb
OxpkhAsc9faxszbh+QqiwMRBZGnguwoBBxGk8KYlwwfv0n9fb1GvvTfowoda3tCB
61+J5dGt0wQXBbYD15FK2xzhS92UbKf03jGccVJgpEIp/DiOjoRjjXzgj8eZlRos
8+rZw8na7KPPBiqIT69Lou0e7D08W638uel8KOddAMH/zrExe+aJjGVrjrjH1oBb
PhlYoo3s9cm2XrxT309F+/Ww8DJjjlCOGsB/RrlpPSjSbpwAmx6VEFf7wB4F2MbK
FHJA8VJVleoMKzk6y4L7sS5ANLbP2Mi68voFyha/ph34iZ7g0OqJ4Jqzi8lqIZOi
GdXtJ9dcbn0PrSrFFxUGIQor9AhSwO7b4QhYx9gl5I8LUEO0ax2nXbDNH0+fdTJ7
/zjuWb+x/QAYZQiyPwdQAeGBUTL0vGeUF+hEvGxHbI+UY+C09J1eG2YBRomwg3sX
UH9CdENzJ0zarrIsTVWmWwSPGFYpDAmTCFCC+xfugqo3Y9oj+AZh4LyIfOKcjzUn
NgDJBUmebYNLSsOA9BV5v/7H3KAVaFxaneM2J5KdnbKlkiw08CtpoS8hw/zoDaoK
e+AcGaii8uui6NU8TJRhQGdpOsOMyg8Qhf2RrM7yF+tDLiMZP40r7nyc9fouxzHD
LCzziQ73LoEzSCssz8lDn2UvlExzAVsmRSGQmyYYRt8soQvICNfiW25JTOGpctFZ
JIt2FZ3FXsGKsT9RuePEazVb9abQZfno46b20PCCDKWL/lDfqc25XV6J7BNv4irk
iQZKZpSA/c6wmt1t9JWqr4eL1qCvYwveOamwM4QD+oh6qU2jleCnY5tBw0udrZJA
iZVSVVp/QjQ8IN9V5iTyHNNRa5CjxDJwe+mSH7j7GBes4Iw3XlBQfRcZhlrqo3lb
4BO3KAzeXs6OUeDGvvgYN5TjvbMvvpnbuPdOOtmgolwczmxRNoG0AstC5Hym29fz
0Io2cLTukBxGgBFE5F850eF3hiz0aQSXDOuRENEeDeKoTXojVSwb0sz0wBiTbTIr
Xgkxfjr29j1nqxj7YbJRjGtnP6norYkSKDeMEditRBhIJ0u4tXn/JMAArTUAS3o2
998OVDypYRYcu3Tu7cM7G4f4Y+ZUzut7VTmKSAdKlHnOf4vsTjens99+2BKB6PVc
chCZkgAHmvRwHyf7wRAGM3eTb27n6wRMa9YuXFLmA4KmK6LHKkU3GKMgY40X+rIv
zBFTHAFjRw9eyKWnCksBex2g84GfYT2Ub3skbIEdelndDh6sQK2ZdZ+W+Y0W+cBB
dNuDiDV9+yXP4fzF5zUERF/JGXKdcRwsYtx4PAx/J1FNtjHSLhC2xnqr76ZAcc+Z
zBkzJdekusneskN9VzkWXUDt1bJ1LAMoVTWwfVzr6bPkqsDbskVCQzqLxkUJRfBc
PbMTf6yakRZEMF5pyNVEGJv4usK/Ty2f83LznKzBxhwmMxkRFj0/7S+cydxQZCJW
KFNyk5CA7tcyOA1mTvXZjaiqJ9dNNFEr802ix7ukdryR96peSRc4qaL1fztV1yvs
ltdTWrj9jIoRGkbi/xCQ7cSoXIlcYHC3gdP6bY4RSeliugHtc/ryA0G4DhmYSYgW
DxQUcsHhaPYzX2p4HTBFMjayFGS9rWhOzQVSiFLcSu8aiAuvjnJvi+PqgnUy4kQj
KpQirOmviC28zHARKExVDvBZlPlKYHjCKiUeoPesAoL5rkrahIP27nh3vyt/+62W
1z8B4XX46mF3lp+1IKBn44BtjcQk0Q5ON2G3qL01a+I9Xh67hPLC2d0O5orohXDk
iCNoOB2KhUyLHF+V8Nl2I97/XecCisH0Y39Ky7IQzI9SIC46zATSyQseZS4Bjx5d
XaEWoh7+tkXb0D6HDg9qRXyiL5TVnSlE3w3LV6hpU0aTNQV5kQal5Zt0CDLFzxfd
5ASqD/4XZgePVTTnVibWYtXrwexjfaP9Dq9FTKfhJ/V6bGE1kO3RDZ6Nl8+QFGQ2
NW6CvxLjEXlzyn7enUIVJ5bWgAMa0CSbGmgsDv8xbpb56g9/0j6MmkArBlEGQG3K
UbpQQ6W4UpkH3a0FHFzquUDBeC2wuOqnRd6t/hTxT/tvBs7ocQfjgfdL0aDzhbzl
2+8xnVxX43hHC/xM7CUTI+rOe6XKMC0r/reG+76pHRp5u428O0ksUvS6ozra7yCQ
Pf0jcRF/ApUSLb5W+aOsKmzz0RrXWjklzaso9WrfUyK18B62p+dZufjSD0E5dg51
5CfE/k9TkR6L0YXwxu2aYuIEI/wSopyhCV7Q1u9V1J8/VSYRNoLx2OpY/YnjDAHU
ReHzqt97FrDhn7Kw2/z9KkEEeEJ4kHQaADPo6LH1ft3V7znaSgSy0fnPmjGSzD8s
wmChJDoTmIiv9tSqcdMeEWjT/l3dAVNowLyKxuCyJpbtHGCeXan2p4NFLXl7rJQW
lbRbZoesAwtNm7dwHxeDBBsnXSFD5UjNv4vMIM6WTuBEDKoesUZOW3Rv7FMEkhUX
BTab/IoC/oKNbZR711UmSqSZ9JCPrbZu00VGoqOgeUH/WMCe93CsgjMEBTs/sm6o
k5hvz426FjExoZnAS5W0nNqiDePRbO0H6eVcgO8sA3JjrAP7gtzEg5/c9GyM8YaC
agU0904crFp81REdGbU8vLYZpxHBpDGRa56bnxj89q4m3+FF2sGb9gjlgytWBwGc
xCm3iz0y2I6TAqmOJ6Ts1pnvnViFigm3auQNHt1HJ65cTG18vDhaP2Eaq5JxpVdP
4PLa0hWA/sA1zngZd/GWSxpdGSE4iBNibMFgn4fuLWL5rKFZ9RhQ3sTb3B0e1rUW
mJLEzim/sh704EJvRLf3jFCBoYCImggDtM1dLKtG6O/uI9xdLdQRaMdGpkF6YfFK
gsXSJACRp7zi8KgZ/tSCtX11NBglm4T06k1aZPM30YulYTtVYmGSQm6NAcQSAnyH
5FARzkQsgf5ateRAiLGnzlGNmOmva8QwFCMLWeZQr7QPpDgZFSVG5wEjINGVe6jZ
pjYWRBDpIrL4sRlCqkRawsF4MEI9kuWtvcPRYZvKMg6LuelcWkz1dFDSEAReQlOZ
McR0mbEhbf3EqzuRaFku1ebm5uZ6ssw/OsWIz3QMPIf5XpRsj+ErOzTaOSg59Q44
NRw/S3pQCvveJ2cFcomgIo4WE3Zk702C7C/H71NDjZ118B5+BbjebbCT8yBIYB1v
LnGukOXizgGBZrSYmI6GuzMXpOYolINpjs0+Nvq3HTjB1SetbsQwiTSf89Lkjqon
38e0qqeMoG8ZCGNc8XOI25Ku4soCnu/fr/vbJbcHZIp/8O8aak5Wrs5QWZUvqByW
xCbZEJAKMNY5C64z6x1H200ZhLE3dzyo8vjpamDgwjmBkzcEkAcIUh3jSpOvKxkq
QYM8kTWDeZJeNcKUmiMCRwHffFtQrcBECwND+q2tki5OVErEtGKMBh38AX26Rs+e
7gVArlp4UHveH3CqeyfxEDy/ucD/fsNn8utn72aQB5RC9YjPQGQdiNx+2jO9L4LZ
UR9febdx/eZq+k/Drm7iGj3tWIOckwYJ6ZCzulO7hFa8DlDzDcaGcOVK32unzbXS
4VH7C4mjweoliA6O6aj1ueDb2hwy5BYjSCLDlovDzjKiHn0Pjj5/JKNI51DtSoNh
hv95HGLJyUg78vuPGN+XJm+YezzDX56eSLXuNX8IlMm4l/LGTP45K9Wk3kEKQqHr
c5RZTdYu7y3wGdEVHiFqn6gcS/WswzEGlP2vrr4V6aMgaxSx+Xr12mhJp2klvCIG
IFLMYwnE3uHGkQNNFO9YsWceLM3ibMm0M86wz/u7VnXxontqAzkNdGh3AwUKBhDA
Fr9Sp3MFFHWI/sknxU7roTOv2OFMxikmYDls+02McbPv3rOfpmFaWKx6AOuRS3o/
QA2XOhk7Skc8rRQlYm7bsjwxYQ1lnH5/c/hgHpaR7wmfXLJPykrfTi95ahpaQq1K
FqlLhnpTKXtmnmwo9/GitbhpRFcOIsxWicxQ1dhJAvm85c/Pn7K9Rr0utv2DfEUe
WSrXpE6aRJpwb83/rhZQjThHiYUShiC+TOGL7lSjOxrIbWAjxNUWXQFkOaMB3W28
TYnjhLK5QOZFi0G8C6V+OnPXziVSWqrjjRgsi1PxvnzzRLA6Lw24oEgVQ64xmgu8
Nf5WO+dGHvjgjKsjs+r/wQDjaR3gtzZvKeNAhdWzBGQlOFkKvNdk1XtOohGtvu/7
3z9LIcOOZMKG2exHrSBVoiHgdVZvW0vYwuVAWLMPo/Z2niXZ4aUMcp7kRWMDiwR6
abzE+HcU0fBv30rEh8ZjEaNfn5HoxUC6xw4CG2wAvIM8aJvuGkvdSriAyo9yIsxe
Fd6VvFAhwE9JGIGB/UUe2q9GctU1CXzHN7f5iFn/u9cjk6Ae/uu8U1b+IP0tPwOF
vRiU24qAfJh/J34gTAptwmAL8Lg6i7441HdebqtX9Daqg4pxCig3BvNPE+U4ayLv
cwk2BV1hCTHMMgvO3kmbY7juLQIvFIHpRa1Q4sqG53OlZpUkocUApe9sDZdFBaJT
FqNDnn+VCgVDxY456w505OD6gfaXUSDA19BbnqGn72lEeB+Eh8CSeSYCVTROVwGp
jNYGgsE/ED2g8GmTcyr1d4vBuqeb4ZkxREPSbhe2oP/0I73QUurCY+zfvqooR3u6
uYu5CYFgbQVekIkCoiR6q9eLEiv5sw1QejtVeIIu6lETBVFWRuY0EFEl2RDjKf0E
1xxKT6J8I8pULnRDjVBiIb9V0Dk5XJ51n9sK/FvUc92/7yLNAyEW31NrGkVljGks
IZ8qmbAv7yaezaJ9UhlPgOgw91uhbUTWz96nniaiw7t79m3WV1f71/EVrf3tKDln
eEHQQrWLgFMzQJMx4A05MxHrejnYbLlshYn+83K83KkDamogm0FJcCUJI9SrmbNe
Kr4as2Y90sjB5JzAJZNvmoYG+j/0omyJxw8VC6P49QXZRK1Skg9MqSGRK3oLmBq9
M2+AQHqsSaznF5IHMJO642CjtCsdrbJOKZUz5SsYyuMWyFThmy2UgKTEv5NEc/fe
rD/wh6+LiEfudqXEXgYJmsr+aX2SI5CZZPvo5Va4uY5iSJRruEaS3dgwM8vR2tXk
Pe+5OH6UJ203f800fHVPB0s53PVKu6Dy9Lcl+HG0oMhtG7G713uReYMVH14sTfkV
PTGAUwUfxg/RsX4PN2lxALHnEvuRut3sctEpyV7joKlikc+rYMHoponqkNuZD+RK
9+4AHWTer9ox3GV2plET1AHzEUy8cJ4aM98j525WdYoOx1xlLLjZcyOZD7u/rntF
7rMJ6fUzTscJnCXT/cfNCp7SsxxkiQ6wzoJjmHyiK/KsSbEpJYMS9Nkxcr04NTCx
zsJR6RfaD/X8IojIDujF8hLsKhQb4QWCcu5fTwZ2Xj5VMH60+pcUqoiT6D+BhFtG
iDRyJyHTISYAWjiLEVE/DjuAbI0KoZsa1vKx1cmoXY0wOVOvYwd9fDfaLxoI0EoY
aM8PVgZlMi2vaFRM1xpNGSYBAewD84/nuEC8ol1Oiot+ZU1lQ6zx8gmXNIa/bHY7
h9Jh70u5qC+WzRC8ctqcL9Ku3OIVE+iqoP+ZUzPFM/L3A0szgAKIsoY8dZjPIcxT
/giBxfo2XPGfdi4FZU+gRpN3OE3x4cak62wkSKghMq9BerXJ0x4jprYe6lmHeSP0
Z6pFQOoiBBA3kqCym4YV2EuMdi8OJ9SycP3R/M0GLOSHJa6AnnbGav2wWS9JcZPb
17teR6ULJI4AQrscoSMYIUK7UTATH2HRiD1rx3V0cAJOa2G9MomJPXfy2DfqB1Uw
/SrC6RUIqY5gtm6m68HqHAbZauO0iPWVw1F/eWxqZoqK8C+G1KoE0NBx2q2+pLkA
gAQsIJAI2cS6ImA0MmbtN3gYFAgfHuL78f9TSezbh7h/tgldJccedHOTtiXHssuj
3rbAYc3PUXLeGSrGs2HaITbEuYxXuWINY6JSjTKuKot2yYsfBpQtUKPs7VAaBbcX
UOIXq7cpCb8Q2EzlCm1gdMPTHUySbue/ma3Dvx6QwD/Y277hmvvXSYOIVkKH74uo
sfr7squJifb2tQcDlBph/s+ELrJwnnAwlUXA7i162Yx1rxoTb8KeF/oF72z3HpwK
98rxP37z9Q/J16DXgRme7n+Wf9iW4oUjkP5OaRlWHI3X+tUp+Te0EQkDsP1/4MVo
KrAQht7QJyZcuxWqed7ODH3koeUy1wA4YQJF0wqGrH5Oz/X8PUbQC6EIKY4eIzZM
qzwnciFCmq4MBX4aSGF/xRTSzLpCVnq/KJMppgdUAG8klLgChf9iy4oFZTNCynY1
I0/3o6Y/boH2L5XqnO32mH0fk2qYNRvegHm7uSpTjEf98tSyBmzG+zJHWS8ZLgYK
qkWU2MaW8+zBTW2fI0sN2UZSeX71ZHQXFSfus4+EZ82RCtwOMLq1o/HR2e0o31zY
z9yJaREIx4JKv133UAKrWQ9z/mXmGafJe1FgXJ5cShkVofb5ddirWfKGFT2htchb
3/F5b45J+k+VO4Wd+takMsyIUPAfwVXOZneJDj34yids/Fr7SbM+g5/BKJmecD2j
y/vDb7ctz8e8Zl9DCEPQnAUoRN/U3zFqO6GlJt8gqylCrt4TBYU919vcNdohn6DG
B4voF5fN1YzDZzLzSYuXUcHjHp9fA5DSj7idrcJy1EXzYYMzJcY8aGMiBFoL4r1c
5KWRV73BrkZ/0NvJM3n19lNlOjqu8Uv5g6M1cEyp6qQgEnJx2NsjT44Pw4RLBdpQ
9m5e93XQPIL8V+r7dJos2NUl1QwW/gbzVoFnZ8IIq9MGwj9SiokhdUtK3AFp2ryk
3RZtKLP0/sFQyJzXJC0YwQfAi3aS1uhZ6WDdQAFbrSAzXYTQPcqmYz0dYmaWmxl+
cIFVhPQrtkhQz9p7fRXSUkTtdPgMmF+9x+6F+0r/ZZ9Nx3MTH/Ter+B9ZtxGPoNu
XmP8EL2TdlOkySn0KhHOdKohQxg3kg8VZ4r7aefoxCYI9qR0CS3HTU1iquf4ECp3
+aUQG4O5WB3pqoLOrmuEykOWOhCkMskvEE9aJUimt4nhgQJGD7BolGvlQY3Ya/+I
tx7HC/8c/J6Kq5O9jCwBMBn8grcQdtlVH11eDIdo16JrM7rIuX+C82jya3pUar9P
igHwGsjFzUbuky5YgvbO2stz3/8SVXXESVC1PMtN/i3UQC03belnao126UKlSD4P
RDIvBy89fapybxJDBK3rRX1sayaLDWFfrqLfMz1gqXum5OQcvPyyawJ+JD9R4UBn
xXPzb474wGWTEGcuy3gzsINi9zYR157yoSEXJc4Z0Wax5x1T+rk5oU+FCYy6zl2f
Tf/1TzbQXg6tMrk6cGRcSrynvhRSQBydlbMUj/FdpzcmCOjF4S886nGS3sXTJGby
r29q9krdfv7hVvii8RcauVLOGmt7HqssKK6PXHn5SwbkvuLrrqzaaRYMgfMCuUrX
9SGdMYAcJvSi+kZiUfjZsbhxfblrDvxmZIMaSVO0NlAWpmmJ/iy97q+hy9ZpoUxw
6DbtaLziMdlJm8+pdMuXDX9doaYwi5tklRDQGuQsdIVi8lyCQ+RowXeQOdix/Q+x
KS27dkuVdYDDxiwRfhiGXYlokIVF45rBqLe4ud+MNrewCJrhS3epCmjGUQ7fF6Xr
mpTolgKjly4EFeT3Gd6Ga1vBeT2OuLNgeq37OefSOkfB9AfyX3JpctzEzPw70P+r
RnrmAp1gDxhy8dRU1ZsN5NHI1xzp+s4hXizd32Jjm7FyI8MDS/faRdNvx/Mi/p6p
IyXjzAALHaJSMsTOgvfJ0cPYi9f9xlMfn+UXLENrAiiBKi3Pspda+v408nHc+Tq8
UWVMxbSYcECcLBmPc8V4CjJqosEbTqKJfDL7XIdbO/zAqkS/jraVvVQQeFOHNOIs
VENY4UrDmEZQo4lgrxMB5nPR6uVFOhyAbyjf0SokE14Opk1WDpW75eW1H0FV6qde
TzRnm/KFjki7JpEn0WQilHgtg8cFu9kSWrHXJgvln/OH18PsggBc3wOdWSyqcK6R
8JQkH1jd1alC98tiEWNAb4tPGJnAd8LNv5GPr73EcXbHupP2JuQERb2JhT2wvDaE
Sjc5DDktO2tVLGds2qQ2eSZPJfRBp+t/LzHfkMj+TZnJslRPTTYVSaSVvslj5a1p
90H9HwMYurci6QGgWHV8gh51uR9hZpfy11JMmO8NBeOur/ZvmHVR2vlD5F7CFYfn
wltA/tvBKxNvAHObuqc8SG4Bd0jvV2dbg3m7yZvQhAITmo6NP44Rz1ASdvD77/Sy
Uxp5WwemATWeyVaTYFWc6JsBhzah4Wor+1bo3PJR9hgkwQOGipF48rBSPuLQHpHy
T2cLZWeUhfZ19UfmR5e/SVzIG8+j9tX1+nEH+j2mCYiWMy85seVUSXKPYO4DKXgS
uCE69mNNdTaEwIcJT3gMms/ieWBVOun9alFcI6PllC4y21mYptpWyugOANAwc13F
DHdtpQjJFXFQsLEoqVt7Y+x/2bbhD8Ec7K/2ImsIC6M6Q3g8lUlKDimGRvssGEAM
t0rZZwcZQ7C9/EZ/jOinpEfnVNlAxNt8ZfZQS9BN8DAie+U7A1aG1odScvjAV6xW
cXKlC9O8pitOK75nRJfnR9p8YkBei4NZoV47WFoVq6C7+3N66P6szij4UCN0Tg92
n3zQQ1YOsMLBIhJygCRlqwkLuZ2H2otYDLEpaM5B3vPxyo/e9vOMGk7at2Tc5iPy
froCDOSNwDGZMpzeyYPcXoSE3ycKkL+rZ6UjGDnFOP/Gu6y/KyyGA2xzS7f3SmKl
36VkkjFz5LhmKJlLR5fAyHEguY0lq2ZfUTyammV4wPU=
`protect END_PROTECTED
