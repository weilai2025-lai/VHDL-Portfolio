`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
geSG74H/yd/keTrQGi2NRuU4rdOM85i82fxl1InZkCISQiKGQKf5YwG4T7j0QIDf
fSx/b4p1UODqWesEjF9gCF3pcUHTj9xikiJCIkaqBMXy2Kck8R0kbf4LcIkpDAIS
3y0L7WjF39F5QY56HgYE2R8PDaLesZcVRSsAhf5e+8EfljDVftRrB1/SY7fCO7n1
D1eDfKaA3/wrYQVbUGNVUCKsiyFhqiJs57rIj3njTcJzh+CE/mSRVs5HCWawQEGj
mCeY29kzmEb8+a9n/SP4xSQkK5iIp38VSJkAox0BAOEl4udaF18RUY1Ogu05s3oU
vK6yyvDVNrrn0eijis/zvLBPpAJKjXXNsXVAiehdJv9isswasd+CCur7ZBVI5jiR
eoxfMCkXtWTfNTUE+nxXLyOMeJFuvogFCMX/LTSKI8lzTh3sZhPk016gFl40WWqr
jp/Kgjj7z8b7SicygtQ57Yr/ZdKonK9TeV5aOmAYSw74WlZ/GchB/fHhjGb94iqp
UXxYhH7b1PtcVGCJ2ZpC5Xn2LovlFKrJAtFhMjMwSVAQ/gn4BWyrRq5QZhU2Y9rY
zGwnwTsCNCBT1GLQpSnmZWKaEIqrllrt/8zO9ezsW23mBFzq3XzCwYPVBxWkD0bJ
cNNa4L0C74J0NQVLjcfaz4eeZnS0xalFKpBgJeCzReHzVeCR1GoFOwLC8m37849s
V/5/6RKtNxhgjRkjwsDM2BR6SMg/gC8IyU3SyWGBgrI+enjt4WjTSlN67XbZrtsS
eTfItYD7z4sv4Z7UwcvFa2lvaUzQS6fUQFDX1Gp5qr+vDK8OrzesI/zsCb0w/Niv
KsjWv10+/7eAyti1OjEX+5oreNDejtOaqkV+cXnFZOfLhofHmuiwi6bJNjxoT2xY
fpJLU9h0X0lUpz0F628SuOUWF9akFYkqkViN4YRNmx/kRUx/Qgkdzm1lwWrxmMqS
XdepF120XR5KQzL+Lhc1JX7ULXfp1M5iH013CkeJb3d+ZCIws6lJgBwzzcsW74nP
Bc2ST9nhRXp62kRx0NBTe+gJjJOnLFE7AO9cjHw2pNPbFlLJ1sdlLHxCNngVtTkk
3S5vk6nlnUt8d+Vv74zEOb7TS4b73qwTO1ddHPx4N+e9fHwgJ9tx2tTjtNvaV1bL
8ez6v3VC/LPpu7/y/zOcDVRVQLu/FAs7YQNOrsLoHK9RHklQCeVL9h9LrXtblTek
Jdm0xZc/7pbboqjgz250yxoKAxenNg7pgTTtoddJwotpwnvswwWgkvrImjzv4iQP
b0c5diQFukjPcBaa8ugWKmrD+7GEIflxy9RyylytYSnYAERQJWK7r3P5C0M2ML4F
/LnFWIjoD58Rk2V7qwEtJYZquPafzUHzV3MyG78C2IyiBj8ao1thk9TMbLBljYKM
NgTUcm4rb1CtfWGjReanfCd7hSAp3vpd/u66YYWrDwF7AWQRhgzDZsbBIhxNYUZq
rRQO3J8hGyOcOMeuOLtxGxq0hBZpQhlH7xiEEyLPXizCLXw5kn862kPoPddEKme6
TD5x6dx99PhjYqwo06r9sxOPZPK60j9cUMTxyKjJpF+imvklBnHMHCE46T859PUq
80aoveZ4wbjZT6HtCLGMmEWOHlRqM0dylPMDvsIQcICs6FqiMhYFDvlaz6KsG4NB
r1ddgp5fx34IHVDKRVnmIg7S0IDgrX4w3rkhhMwZwF/ZeQsAyTQjretu45FuAzR6
1IaF+RnHjwgedbANeC1tiyfzv4wpUitcQidvTwcYe49mPE+UhvMsuWVfNxYeV0XA
JlJqfqAhmlL7sezixTyaPjwMw20XwuiAP1QAJlujBMKT9ghCv15qIQk1IQtdRNV2
CyYnIf6EfmuzQiVrCoXa6ordpKZs4W5wq0SpxwTzdEMV2gdbjJKhZxQLsOJZZOiB
vQu7gPDGH/4g4vhIBYtQlUd1ixuVh/GaM1QOuV+oyxF9lSkyVrMJkZUsnBm7/LFR
i9CsbCoqk+NnP8lbt/Lf/su+rjUGaOVuNCQeC2UnPp4pXhlOILbRQws8P57vzSij
DRdyghtnr0K+FM2kFZ7e/kPKxVI+djMsAllL7hZ+MMyv/soV04jvE15LcVNGlqAo
FpWK/a/lelt4bPhEKTdHkDNx7d4JVl58b2pu2aORHZfZydwbjkG3cM9pZoI3ApZk
ZZYeCAnQguUaf0wSVqh9Fz0bhP2OrT2F34lM7BQEj5JobWnGhkYHGK2PxMV+nwZV
AEYZ8GG3FLpL8H+VdizSR/ANY+YDk7y858FCUUIJI7TaTkUcN8K8NYrfTwSw271S
u8IysOFf6cU7oxLYMZbIPnE+sM33LqAIOGzFQMgAlamGD+0DGnb49/PUsTWWqDd6
E9e2xaAD66G8+p+CiyqLsy3aG6yuNrP1ppXbbbewYSGSUBx4QXgfj5Ar5wf1Crgw
7SoUW24wOlQKpIqHDJhJJD1pWBNyiVkVapAn2JtETcknO4fODUwQNoVG6n7n/aAN
LrGgvdYpeQwFvSwNDIqX2bgZAT3qxah9lcTuv3BngmWeT+TZLsWYiRyMKblNC+Sp
LReV9UPUkxNdRc/BcG4Hog8keOo5hRhE+yIjTe4V1dTldyQb4JodgOzzp1rC9Ct+
VVJ+cBMP+eXmAyMrvLO+rsILUDcFpUAVa/uivGDnAEBZbe2WWSCUKM8aneIdDyqQ
WQA/0zr+0lQxOwxSUfThpFetylqY18IPXUmrJy3TCVa1eUG55SbCRI8rp03sn+14
BFUeLs/BwDd/TLgeqOfjcWXexLPaIDJYeYieHoMMMaWm3uECe0PaxkB4aR0TihQ8
mHHDCXqZPP7p2ppCuGx8jl75Azl19p7IzcBOmoNachkTpMpjpIpLF5UuYRFmddK/
I66qRIR4WBKakCCC2yM5CDafsIWAfqFMG9RpCqg7GC/ceCkVnooTZyIuzuZaNe+d
Qarq1gRP0YGFuT7lHnUs/ZKKNJK/JrVZux5jwqwqECptw3qQynPeifiowaRqp8GU
yMHRQIGWodeRRAMlVs8/U9AXCSJliDcYKN4fAp9aEkfBVHNuIjyYYeWH5YmprVE7
0/QYLXf67njq0JgBa52GJ6XoW5to4xcePVhkLMkc8Pw46QqUOWBlZ7k5fkcMIPmf
UpZLCfv8U2GQjTnuyIuheUA9NgymqNCCK0oQBFB5VrhUPKvuhptUSICKTAb/1Jlz
DudGoggCDi81YxNj0bRF0rUvVpaofnjeirvo6jb9++/D0BrsPdhJsyPFlQa3SDK8
rjbJW8o9kSbCdlzvxVhCtaP4PaNl4UKch8YJ22B676nBDDGHrssHDQDpPQMHR+YP
bqeibqJsMQqc/12TOdIndN3Jj9NwRR3Jg91sEloT/trQ3cud5Hj0XiTEW8S9eqc0
gwfOnkxyB1lXUX/K006zE8FUtkyYYr/n6NAOhwD0xIE0XW3ipYsW7w7aC2f7Mwzw
2dnG+Y3MvvwwDsF4s0dKLvP92xiEF//USiW3mQeR6coQqbstgvipZ7e9TcCzMVoy
R04lB1WYOg/1Jatpg+4jcR7YGi3iMudz0Rn7j2yRq5Ki4LUTKL0CoV+W1XiCjyur
2rpqOUdWkidB1A4dH0lDXistpqo84JbCOeO6/buqcIKVzaLt7WMZDnRYFsVMkjB5
6pcdTWVz7pES5+rKHr1tmx0hYtFZ5eaT3SZBpGQnx8f+GSNwCWJo4KyRdIfN0J77
lPbF7k+m1zPAlarvBXF3gL9LBnMnrptAu4henWv7QtTbT5rfOfzZiHb7hQU9V7Ga
hKgIIqXYELfpTAQX0QqX0UHMiCCFyez3jQXP2TnoQh4k8CmTdafN7S/Pks3tXXY4
TSG1CJQojBYMZNtcwUvF/y7T0gTJrF/e23v52iLQiiBAEyIgwE+53hF6fjXDDtjY
mcke9TEeNIiL4UNgd4My9ZVuCW4JB3ToHrToeQ1Md2tgEfv79E+T0BQLL0hmR8wU
d3GizMFjBWqMtQQjMcdbR77apQAjBsjm7qKV8u+nQLc7S4nWqsZPDMPM8Og8Es+Y
AblavbHaVunlhxoVRonJns7t5M4/5s1LHIOcyxdpPH3WPOeHYqyAYChKMA0udfzL
Vtsi59HJ7MvdzQHRFPDgB1s9XGJn0FHI72i9DHdJfgCSs2hUIda45YkqUfbxemxR
pUzDNrVhm5noiySVEfIwazAwJo1i41P1Dm+HyV58uAfRdFBPwrm19Vg3iuOlaMeQ
HRUFhImLeuaQ7ycXxo8WBIUd3as5DA76BUl54es067w1f2529qnNZ4XaAzZUe3LN
DSMDTakk1PdpSFl1G7BwQL5ZlyxbeDpenvA85VLUIpbfPnTPD6LgkhippJ8+X9zU
6vT33n2Ktu79b+nK0D1oI0RxUGgtN/1k5ofYEsUOa8s=
`protect END_PROTECTED
