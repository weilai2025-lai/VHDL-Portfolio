`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8axyZTumXhw1BcuNTypNUeVdw96DRVH2ZTL+Iign72NnOg1zisBqgH3/3KBzxM9j
Q83E7yaVyKCFqk1W1ctslV8xVArBoseb7r/nIbKWSlJOERVLgUtDooqjzj2azFCp
Bh5OvvBXnJRPnUimA27WusPWsaFi7knEp7LwqFwdls8eKimwN0taC3bwao6oeom+
UNDXRi7ooV5tVzRPYEgNqPLLAgQ0XaJTqYqJni8cj3LxEVGhUv8RtPpCHurJ9Vor
Oyh6Rtjg+IagLQrh02jxpz6+6AKGZcJfhpaO4HdX4HW1FVpYk69OlbcOVlCtv1+U
RBKT9glmCoaBTwXNd2abt7iTC1XrdHRmfRnYKhxT/B58jEdTWIo6yvaW/Agz0QE6
UMWnOBCQuHPguw1DVRuu1H8No+ztznydef4lzfd2NDpXFnyDd9SKJvT4Lff/o0Tf
t2dD+Y2xJPxnHbNfCHW2TTJsS0CVzRAmv0JFC9smnjM54eWq+Z5KJQaL2C5gJ8Es
bXEIviCdqJ3xMPSZ4NdyWRQZBGlTr4ucyD1xdIZGtls4oPfV2fSTfEIDXrtwDGFf
2bOqOYRBi/TxxfCEV8MxzKBuImkrTGFJCNAEfhq5FDJuWA9m5g0ve+OR6SrJMFcQ
SCZ6Mu2BCtt8rcJf9nrJnZqRjh7BamdN+X3i7FLYSzT1Ok4s+fWoE74BTN0h8Hl3
IpWnOfD1Ag9/ONQINznd1PpA/qWo79bZdCWYdmXyEwzuy87weBzMZ6TzWWEWqyO2
wUhX9dg+W+HXkaQaSZ7m/T7MkAHKW/10wMxKLOwBNGzA1LXiQCSegcZ67g0uKZpA
KSrWhZp3kMcxUt3UEgWcuZZsgskl8vtXmKI9/RIW77VZIJ7OYqhXK3rtxrLzobby
7qqQ5mmTPGMy9/0YQvGs/FxRmQYPTYEpkVov52tofYuGIrtl+z3Cd9/8gVSDZZ9d
hXVztGpJom+2/HhvhNhwoLs1BEC3U7dTazBzUMSIs6AYj/OSJ9pAK1e8MtmKc4wo
p8dU74VnPm6eY35jcUV4e9H+mwljp4iplDtycaGy6e27UZ2UGnIOpUhKHH/+Jl+Q
bJ/cqmu/KAqML9OpI6KY3uSuxVuAIZTH0gl6SqSICFQH4+Bz+ChaKxf+uQcPkjIz
YP+8ogL/sDeFbf4PpBDlGB8CJVpUNLP564X993i9afEWAl4zeK0UXWeg4xKQMtzg
bC5tb12EHl30Q+Kz8YGXsvkAHQHUpSfG8Ie3K8fBViOyDEDZBnLrPnHksBG3pAxY
uYi2M9BdNyS64kZYqjCQ6VVAsxHNKpzZyK3gKOQMhjMK1pF+05rDOl+nt4GSTXyC
EoELIMTx9AAsL0zG+GweRmPNtoLnsNVCxbMCSSgHtPW1/0d4vJL7zxhsjnQJlDab
Lwc0UOfsMqyLQWts3gkE3YExaDC4BT6gCwGUt6ibPWZ0+cZOmReSYXnPGmmMEbad
brBZ9DiboTIMquNJUrdd5uQiWHFxB2f26nKxD9IXJk18T0sMde/nzXmNF1BC5KHz
MvINCJ9HAlz5HO1BVEf5rcQ5TnMPrRxYR3EX0CHJppSehMW7XKWcOyaGmxYk5TDf
sxDHReFLRAFk7Bnn/xLwAiKBo4wtsRv8ZcY4/FY3TV2ew8KYOWSPPfdbAkvWEYqI
oXjxUS3vfQqGLT8/ADPjg8plWVRLUg02W1z0CnoNnI+22KCRbc8uifDyhcQJo/Ry
JRLBWOnTVbOvD5tDvXzdqd69bfCA/b9oGXunjCJZCHB2PL2rRJx+9bXOZqeKIUeq
qSI1eaEn0kztKI+P8Y3imO/Bo/WaGoJs79XjP+tEmcwKiZx55ixODBGhek3d2mJZ
2b5L4YdZs5Orr4Rc2posizV/z09pnnvGA5uDV7MJkMC8xz7HU0kE5/X3GNpUmGWa
ijrNzWytT2Zbtc6RMKNhIYZ1B4XSm5xyxwXNvgNlAM/KWdDWz8Asz/8xsgcref8i
5P9U8mkDeTCRLAY0iCN5qxNZ/aK1ntqmg/W6HjiIzMJIT00hC+KNRrXp4E6IJxgx
SJw5icRLclJ395GPIvPkghALaWXaPnB2kKuYyFUWG1zNbcO3mN1IdyuWJGqGc6yE
9FFVpeg1d/iKJxdOEMRJp3ZPMnnobxR1y19C9cJkpBGzGCC5LhEE9XM+MUxnz52L
SiikUsJDkylfWxGiLldapU2ZZhnq0+1PIq7Qr6mcUkBuxxjDJKf8Q/XDci3pFr4Y
rOfJVpYvuvcrW/+2hYFI3F0gtaMD8TbBFLD0zyS9mop+hdjU04euTbceq8UUM3bJ
7ImMpuZlOLSOFF8jfIzXuB9w6L1n4HeJU8ZW/K7OARlPVI2qO5Zg3pSWiN74f/Lm
qBROz3JTGbANrmkyY5uamVQzkjNnecRa5g6uQy0nJkHmEoCY8G8f8zLLEY3a0+oU
NNwGATG6VVA9/FBuXsiykM/FtjzpT84iZjsITnpVIeBA90bUkw0qt4z6WVc8mYlO
IO0d3SYZwxY5C2kuBH2cH+S+GBVFxrZLT5pHA2AtSAaj31zfoJncLNIZP5JhE/f3
KqN4LOBPxiPO37lH+5G/OTeJIORxrR71e6Ly5Gj6x7E47ykX4SLYxKGd33uNQrFv
WHe7jpPTu7esa+qE+KW06xXevTSItN6S5+K0ZHPo4rVNI92cB7cxAQBGnzcsLVVg
OP4r8OhNpdcyvFWvlnfL3iBG4dz4/ZGhah+k5QulJwM31gPT9QwZUXvgGtSKGfvk
Lv3EaWd66W0GgYkf13ef1gA83dbGtzbPA/ZJLoDwyevMtm5aUpDZjXkKCVhHK1Z8
wPd0+i2hSZ2Wt7fO5/fGxl+jF6c3ftrMWQeSPiWOYhjjJwB9TMXXTnfKJbP0x+4k
Y/s9LtFjS8L3NOhMhQtRrfXY1i2mFl63gZBcnrcn+D8VyO/ilR7c9SzdOI3UOhnW
R4uRdwPmAHX9P5ZIMPeSz+wIX2EKci49Q0SqkKk1fO0=
`protect END_PROTECTED
