`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbD0PeTB8eqsPt+y4gHihlcRCZQKQMcnphz0vdgrwCovxbWXJ1wDdM3udgCuAynz
t1P5yDj9ZQB+XF6kOsyICQtWYhVZ/apkAUHwbQMiKLJmQBCKOngXFEFXv+xM1lpR
iqtGyFSaUbaN4w41kairQYEr6ocX7g4Fs/20n6b5yqkn5wK5KAjXItyIGcl9iXYq
AllcZJj19WRLT7c9/Xvx16KE6mKExZZ942Nhk9ol446f+PH2oOIHg2Hgj4X99WKF
dZ303/MT4oe0cHONzBZ1VQ1/WjPLeHwOf/muhWo8+ux3Jx/lTazi4BNtr4HBHyUj
m5QO5momUvn6PPkXZWVrBYeM3tLqmhvYygeFDsHAV4bPPaT6M6tXwkyCQGNluE+l
gjFRvW6Yu2Hv3TCjGQhlKSciV7wrh6Z1oqyX0G80j76W6kF40o4RSilY4d+xlFh5
BlMY3VKI/AmJRQbm6CHBpKsOnJwZrnkYxM75HfUQ9waBtiDU5MXN6LC6YxqWBx9a
Oe4tVmNRGsxQgQ2MqB724S+e53Cx+WJ8SXpyzemEajm5f7P4fvmbF7v+pEynkylY
yovaUP8ZaHqgleIa1BX02Q2DxogF0q0QXvyX/jGc3P7DLkQ/ZIwNcvtMtOobVrW1
33x8kVXjtV4CYlijH2HqjFi+Y5AxJarY1s+bgK4ek1OTu3v2E5FIoGpiPuRhRjz/
uPbErK6gxrEteendWryD6Ek5zoZzVOArzitgCiolq6p5ZgWtKuVF/WG+2x8nqlXS
/QaR+HG14Ezft+aYn77oXwndva4AV0ELCGnw56mmbK8Qys/aeNyOKb7Vdp5ppwE0
iVUpjCkF1wZ5kUJkgmlQQKyoUAemCLbG5R8pqo34gPlbqSrg3BYQTyN8Ul6R4H9n
MGKB+C2T65/VVP8ogb/1Wip68WiaFwD7EmpY3MvnzKaxnysvFsPgPCrGqCKKeVHY
1Z9pGz10+xQX8i3g7SGA/J0VJDaz8c8DJUpejrf8YVNde9xW0+wWpErM6XmEJwdF
cGog++dGpMx1f7i+oOr5dEm4taTWONUsbQay1VuhpCEg0scWmWBH/qzSxVqrzBvU
+Wv9JRyuLg8p7TG9rs7OxK/AgfFegQ4LMi/zQxYSaPElTX6+v09AHveaCWh0hYha
UhDgSXLHWjD1mMjc6Kjch4ilNI7Ere2WrqUOsUgfeo4zj0D5nunGBwxll4AM1952
Hb6sMovUAXIQdlKFCBJU6Twt1h/dHaPTKn4MpiwYhY/6P8x4JOaGSgnJeGMTTzsH
82pY4y3vEMvd7VYBt3wvVt3qyvRm9r0pkcd9scbpPobaffO1P03fzC4yZSN7YVxF
YovJ5lybQUxT6oVApa2M2XRXZMHsd5KBshBiV84L7NmpaEstWUXkM2qXYj7gnyqD
4LTg1GVLsE0E0jCQzJHpRvd97HurUty91UZvhOEvLyakNBTI+rb5+OvBKa1CgKgV
IOTLTUNHFepL7GVJKffkH9FGI70QcSKhR2yolV+He4y2qLw04KYOGZhkliCd4ZQS
GH29Q8Lo42nyc2k2iSvVQcvxKBCdBHptOyhwDa5PPBNPhCbeK7k4O5RSN9sEUahc
kqSXc4M33roVOXBHlQVKrnVa6SH5yjxoBF6a0IJSAZ3f6T99oK9Ag8HgdTa+gCA+
lGh0xYKdWeNCap+ZnOfQLdsHFL4y81HwrsiWjEBlNNSx4CnJFvtiJLhzTs+yWCyG
ZDx54VgL01otvA4rMwIe+2s7Dgv0oux/iMKQAJ5sVDiSNnBMQ9u4kNvMK0bz9KhI
q4TMuvSzgalC4x/g/4s3hsFSEpFDgjz/5+kRD87o+jUuT9W2EhCHW+alI72vd0N3
6KblsOG4/61v4RvbHfulFT7H0JkN2dnfsrw902nNMPohe0RghODK9F6KJHA96hqZ
SK2Q813MTOROyPB+3866AhTyiPD+kCGbIkH8g4entHl2/C4vQctC+mBWHXSMVaMM
1zfGBWpPv+2FXQoVdY/2A9l4xqNHmvM5NJNpfjsG2zZKdqmPILbkU7BXzSSM2MOG
oIYxzUWdhCYHtGlISqC8nUtsf6LdMCGfFXyYzYgdldrJGG0T7y0LPTjUlOQBfs5E
W6foDH/G+zigFEC0jX1ZC2qDRuUqN0xSemPIEzNgMuAJP7HtMcvp3zAPX38vLYMG
xYboPKukWzjLXCS5Hd5Rw409GE+Si7Htw2cmAk4Yt1pA0/uL+4YEdfm3SeCdt1eK
NnJCMMj4lERyLkQr5j4RQ2DjEjFvTEfJrw96j2h9ugz+Oks9pv/AdlFa4hToZGzK
o81zRv2j77rQ9YMxYS0h1lPblqYqBYe9N2THv4MD/mKghCF4DCUrIandC/eHwhi9
FkpHMTvDIu9PBakJ711FmXZ9d5BvtagnCqrutGrZ1H0NJTGG0dlMi5e/suGOqNFm
760oZxronw8epowbVl1+vctOKktZtxQQUIipfrFhyf+TFZ+4kXbYl/6xKcCfQfyt
A5o6celBAcvpLnulBuMEhPHLd/Y4bOQ7LeMJIAZKIYIvsaoqycOkxkwZL3rGFA5k
6MmO38GEeTxF8+XMJFWO+MxhN7+8wZbll+UKyLYrCYz5zcl/e79qrTU6SuuxM0Df
V9kOfoJVs8lp4Ew1AYATQv2rSfqtkT/XOE/uip2YNgtjxwT6RpR7vSptCLuwT0t3
TksF2mnwPd1hujK7EBUytPt2VXJJJfWjJu75hMvDmN/lB8ASa2sCV50hry2b4FZe
sQRWQzcSG4B2n6ImZAdz1HOc1n/qjppDI+Ys8HuUUo6WFMnBz8S33k9PXI07l4cL
XU0D1vU5qduk10Z5tFA56stEaq2hMo3Md4p4YVY+zz7O47SI7PNYw89FbvsAQ/AV
frg96V0UzhHgBd2cHUIAHcL/W612r/X7+Sq1bWmcVRs/prE8gmnDPM2mXPQNTRXs
KXL5o0DqfVDI3Da4oTQbTnbFyfgoxYaXxVl/iWPyraF9RQ90WOIx0FUKJoiQVZhh
cV5HlAfJf8xUVxZZuBC0mE8FXdqQ1Z1ZAc57FAAw34KOPY151Fh0V9JL2wjjfA5Z
2BQNe4549yluDRyrg3tlwJMY3+ZanYzG1/s9HRz4l5VDdsN0TlkE1+B9J6/NxTTL
o5dwu24auMTWY3Vgh3uK0oTAGpOl0jD4C+Fh/z9jhTTCj0j3eWX77NERq48r+447
mTJIbQHyXvGysp6fbNOqhrjvOvmNTmOatZqG7peNUErHpE/l8DW4GW3sRzDxurwP
P6molyOqJBPm/po/pTCyfrh7JvP60HocfTIwcVqVgqC8xeGCDQSDQN/uLjkt39ta
ZowfvoKmEf5fTudZjXOX3rw+ao39y9azYjdGPG0jppDdoIPLSE9tdVi+TQGoTt9L
k52A5jfoDLTXQftNtpLIKjE994BD80pPWybNz3AvHIO9xY8fDu5YdRSk9NuMXVub
wKWkm5G7e1Fi5FkJp6vgSYyWRazySnWGj9fym8a71IsC3PPibpjfPDc1NO+pYt/3
P//bB68XLXaUaBf7N48j8PRi7Sg+ZVVpGXy68r48PiSYrgupIUWLhwViDwzfZrm6
+EsTHPZ+NYPyr1YhRRybrdhKwfLl5XuiVOGFpe7I4UvMZztHcDtcCuFcNjSLe9r3
Ei1ZBkpUPpf3LJYi23aXBKJCVLERMZ5kfI1tAZVCCwjU8SbdwoEkgYlK6WArE96+
eeXQR9Bbc7LXuJaMPudQ8McqHM+ECUnBmX+d/GYNzDeij/h0gVQncunnEfdlFP81
UscCTCrwbyEJqjamNdhEiTkTFOtgrr1ntd5ptkTvNeQBJZusCPG28E1IMurLFoA6
wgU2APNFKXyM0lEuc6Df048IGLCwsJrqz1ziGPXfFHkiDSwANiaqlrI64IBi5y7U
FEW1eoBhezRZ+RyTtdB6yaOsIBCIhYr8EclZH7N/U/PZQ+lS/sb1MTVcxmyQVMaR
XLsMcQlCqEP3dnBOM81V13BtfqASuAteXRoZrytzGhhRmz89xXaHS7190wSbr0u0
Ln7B8pUrhf1eFVmOhSxF8vNfiTZdsdGVjXL/iG+wzzRYO1QJz0AgWqQ3RhsVw4+k
VqX5fMfem3xYU1OQIa/vKYIS4zua+8KExJvXSmhSVLjbF/WZLzP4N8KQdws1Al16
Hi8FxKC+W6OQJJ9Fri7ZJkaOdCUA4Tdq//0sw0TtGBKhkSIoumUSFcWU2knxY0Te
21lEV25NlVL7At2PZ+xyMbGigazY/WumMo3zib0AHFpW1VgIFmxYrkrQoCqvjF6b
vnxVDRc21QSz03uO4kUOJGqs8hDlF5s9ioJPZJ1/aGjL5UraegC5h9JGD6Eqw82t
PQA08vPZ9VPPxetUcM0eJDu8LiPxpycJJWWp3lkqDwE8lPo36yRGipoybGe+8vBf
u6UjBBtJ2Jo3hi5Er0UrOOx/ZEFON/cOCIQeWTg2qjJnFut0EMcqmHlLPcHduLJu
7MYKU4Kz9YGajynPkS9slIjyDSrKxyfBfcyl1WY9xNmK1Qyd8fTN9/KyhMBR/h0+
9z0al6FpImkQKnQ6105OYbboSmVbAZDEvfEhtgMZ4odZ+GOQihUyn1FE7kAXgJd5
pO5Ly2n3mbj3zjIUjrhsGzikl+UR6onoRcuVPf8xOKm3uXAk/pj4pFSd9y7pWgDw
Y6mtCAfp4yBqG5CSjt1eLSW1AaL9R94YH5IsjyFdbLP6H4gHV5ggMZcz2EW5IXqC
Ngoe8F+KoPTRhj8yA5avG4CmolHko/XFh9LpF26zEh7madq49TJp4l//e8lRK8qp
g8EeT5suVBGJ3pp+HOtCKhl0DpSPjpCnBTNwbYkOrbuWnx2GW18S3JrvQcXvWJyz
ScgnN5H+rvWN96H9MaR9l12glNxYusjq/fVC42OtgxgwoOaPjCu/MCNN3acnjZrn
uDgN80GClIzjhAlDftEUF+QouqN3YDr1isxQ9TI7w6/dPnE44dEaFgFiULkxGfaL
Y8LoZnhiUP27ZBtBOWRrXE5/GKAS+IZlxyiBe2kzRjW938r3zkjGAnjJe70mBnYB
1e2BBFSI4fR3HX4aVLm15UxTebNbFZzi7SerS5FJS87R93DYBNK6NVoqfTgXFtO4
BYjBcjcjjC/6YYRDLAuUyGUCh4e1UnhA26Bu2D6X22Jnu9y0Y08Do0WLvWAupuVe
YCyIJSGI7bxSdA2FKwkmUvkmSSPlvNA9FGPnU3TASSQzY+u3D1G/H6y3R6gTUb0B
20nOf16SJebwOrLZVsNZsV1zOpsu0zl9b3OKRLnMFl20nfg9m7BLj4uVDh9tdt0P
1JfQFocZWscfDUFvkGCLSMfoU6JLZkaYnbpIt2T+hBuElAQZFrmqH/fUfv0KXn94
+T9xzTa5Kjx8Wr1Jja4iU0BSqgQqGA3ktEuTJHC89tW6BM7xF1KiInhZAEtx285V
p/WH4FScMXd3QgGYvOJ0tEhp6NvvdxwtXhoSXNFzRBmNKZzMkRIe9MtlaEfn93p0
Hsu2DclfeqQHTh5V6W/ElrfSkbpIXiw2Aha5axJ/n8V9n5HDotpG9WMVSjFnWW4k
SS4g54X4HvqZxGSLleM6JuFJ2vyiXAMv51PI2mrG3f5nQNyRo9FeGRDw3vhxLAq/
VrcCWw8VR34SANrexd7ztVyB4acQlpl0vXtfTpAwje/FW8xYmzkq9BIPQ+AjzIzS
3oHlYtJmJGIbNVnvZ5qlUncSZdfGNLwyshVT6vVR0somg3pEZYc36bIDroaj/OkZ
jnRtpJasaES2N89wl2H5vAMmJ/mLvqDqOV2mVLApPgFZxGDPzj4roRGNyuHRdod4
9OuJRmP4SHqk1q61sIJJBvoBME6cmA2a5JZscIinx4G7AR/pMTctSddQVsvIT0PC
lN+3QsMXArWoI3CtPPbQhDhTbWnGKwAro+NiZ1BEeWesBhX9S6+glm7NQEGiLqY8
epsv3G4nExAd/SqZpR1hMBLz7D4X55NlFHJ7YUXmBhWdaFuLay+9GB3VAmBBQkLH
gjgZ1zZr9jKv4K8yVUsY4fbVSjQXyZmqIxdgnDQSC+4Q0Fy3LHJ/bLzH6oQ7LLfe
baiL/VpZUsKQWa6bxDXB0AUqZSdZax8ZCThYeO6Hx9xJ5dT0E8zKoGJ8RH9Pgikg
Vk9c+y+KaPUVa5DO+8MIuUPPuuhauuNA+kteX7XlcJi0oeASCOH3NsE9CFAdPu7b
KgRiLNx9NETgI3N/p3PM1TvnFh8/4WinnQRNsLtV00BtsfzydPpA615QPM4XobOU
Sy4kgk0JWcLpyU2FHaptzyYEKvq4a7BNK0L1PIlfCH3l8IBvsjA04sW7fduez0oE
Dxm/af0UJIk+ehg9jj6BxU5eDsXX5AivLkq1rCrAhSUBo+sGj1P4M8x23PMkTbNN
Rw21kr/zfMbJweL/Xkr9ho45tWnA8Az/mvUvcq3WwwCgPWsa0SNA3UJqzVGnh1bs
+KCw2wB5hOC0r39IkDtTTHrlivxODb1IxiDe0x0mtjnV4eNFjGeNOoWMXsYlVwo8
UPCh8QIqRoG/auiCJLkLEngsxrAotfH6HQxDMl6HNjD/k5CGYcymcW48cD4KmgVN
QuvnWMGJZfMsyQAsXR3YzvYzrvtzVvBIvf+O8/Lm8zt6Es4iD7iyfGQ4n71hfQlo
N0kWZxuqeRH+cTgoWy2gHS6P/5WXlUK+m8v/7TsUFhZg2rD/k1sT9z5RNeif6Ook
A/SycNZvfS445fSd6AFGVIyoXVfgMpdAr97kajUHE9xx00aRUzYO/z0+cz0Tt0NN
6Cht6RrP/p9pHRlNSXH/9TNKR0czJG1RFcjO5rWTR9x/+retBjPAmEY11RfmbaUy
C1i7HxEIdbEDl0zNHKJqooL1DlgxicBc0ea1SNWmzsTci8iWQnwhD90TTMxl20FX
Dp/GbmXsINDs6j0tkdH5p5O9YlRK5Au/kqXUM+wg0HOQi0B6+9kluJLeD0qEaVjR
ttLgH8WFFFfQnEqo17RC/oKsdGT4uqiOop8SMy1jBonoGUF1Sp76q/US+gE0d0el
uq5vlQpLrpGuDOhbeDvj/V4lYTYzGXo91KnzXPTfjA5cxwGin5fXfh80IT/8Fs0d
NEVV3pmwPqWF59aAwnDfHO4X6uSdltQ5kSnM1Ra8/KbdHrCfGQiKf8tkGaXJAuPk
+icyqRgWNWyrqBEd43LMmXq234DaTRGxbNvaVPAmJbMr69dVKFYzG4srArCSmZPc
PQDqmEpTtZI+aj/obN5TF8vmWKZulaD4Wx0xq7wGJAYr0mJtQ6EAKVIPaVPE1cNF
Nlf+xdi4Rz8ZI/9n1VZ5oqrh0lz7sEItPM6bim7uHb5rka140n6A0E6dAi44geji
zjphaT7w3RdtvYs5cs+u2w2gYrCl9nnukKPgLqDKq25pSklMrBZ6c+3M+WwqSzqI
PCc9uvGNFViH5ygTiLLiXukJ783bYzEGsntxGqjAZfAYxA7RlJHxddcJWBf10l7s
Q6HDFBPkgi1Ij3wjZ05+CKJx9vvkuaizFEx2vpKwwPmNoytxtIuMo9Nf8Deo83ug
h4wgtw3Wr6Mi0mkvQkaANWoKJuTUGTQhKQBAeJ5PePAWQOxYqWL96chf3K9QMTfJ
7b/jtSmk/NXCyGlXVL3XXTXZtkGuZ+DYSqns3iLUxFhRMqk+v2yVISEg66B2Mmnx
J2PrHSa8dROtD7VzPVUoxehKjb8+ZaMYjvQqfZ8SQurWMQrb7sFgEnlVTnFc8jD8
3ycammx5jJh2eoAZ3Scq5IDUfSWIGzJlCDVzn3+eVN9omAkgoR8rJ5FugWiJV8AT
wALzpNtiifk9l7+Pdqa9ElemcOkpOtVG/6zMUzm8BnHkHb676SrYoYY/j6ecU/jp
Iz4mu3+aFfIAtrEmY2p+/CuFWlGsLl4iAhnLPXN8H93LcM+32QFZSFiIqrdQHH+o
Bri4mwy+U2mrKjLli/mZwYRkT6C2DUSRcO0Z0YHdbAeNVJ02rwwl6qmnjUYo79NL
+tYB2PBBGgcYUUh8qblUDqfCRY0eNRuoGAo8wiC36R4JZQHlCZgiBGcpX9WAX7Xl
wT+3VyF0ezDVA2BZtCnTMF05RqPeacHB/i7jwkXNeB6W2Vj+5brQX6LlUe/aZ+kt
wQjro5BwpoxSl14kZNa7Q/gmgN5HVf7TG0gZhGH/mANsYPlcZ/ZMWxz4lXqG0Obd
cPmBkQSEYZUKIieL3bCBI1EeRK7xf6F1caAE0RAzP2tWn9Mvs0j4whRgEswPbY5d
YiuXs1+7jbRAk9fYcXLWYJsweDFHZNBSZMyvPDF7yxELRCWWUaCFqBmtdBos9x9q
leKLkoXfaHAbV+Swx4P6OcZiStN53hW6lskw7FBU9u8zKGzzHpd4tmSCd8Ele+jg
6NckElHNRiZPjpGfm/yt9zGKZ0b4oQH2c27tmD9Su2Tp6SZxEn/VH0oSwYc84c8o
2vTcAPySlM+fvhKEBP27CZhfiM536pn+MFizezCyPnQhdL22/r1sGqR3FW+NJqg3
o9IZgObLjJNCAXWxHOwRqNuD4IHcrSqC6fsA1j8oDLwl1VowjDPJzkb/flPqZHgR
oI0jYfyeNEq3NUXQ8BrXycC8mizpcmzT6XLPPgHCgL0LTvUYHO2Y4c7FDcEYYvQP
AnU6OM/XBHbsfQgqb/G1JVcMTwc9o7sY0erd9OdCUT0RL41cyIV9RT+w1rr0orKg
sXeyaekUh4hE9NhLRWaGOsybNlPbXOv8AyazKQPO6CMsAAeqff5PTQV9YWU0ZBnJ
R0Voo3jzISsR5rSry0AyE4WKMkubxPhPhnMhHGBXV4FiO/tXZlVVjlbusgNkyHV0
aLug6L3Kf8bbpTJLqMYuko/EDfuq2YHUNwKVqIHazBhHgufGcB1on8vkTUnm60Rj
gUtKDncyvveElyyc5ci3mK3mW9FbHjerqF1h1GYUGJHVe3KMDwZ4o7lLmt5Tl0JL
HR6WJNeSjY1Y9iZkeeaMXai6zTdowB+rWH0VAZs/Xo3L8NheaXzf7lKbtcqno1M+
N41i0SvawuhMSAidkbv5InVsqiUpI++dSNdtQL/EYU0ggpott8/eiQrGb/gLUkSb
k7nKqyV6y3yVtm4K0RNHeku4i1osTfBfO9Wcgz7oA9fMmUEPjySq1+blDNEOq+Go
tJ83Apad/v5PDUDMwyCiF6HNeY/wHBos2+nH9Th38j3/u2Ve69n9TeZbLYVemE2X
T6vV0Attv/KoaC1wrx1hsQAHz9sLo1Ml1ztXyXzk6HWCkyeVSHX1QwkuUFf37ewn
EgTe3xPXnhS6O5DzNyNfhc21HYH73X8YjnNMjc+AxBhbO/ITaruZIborhEcxSHP5
8oidwQLiNs21O2xn4/iwC0iIBrRok5YRhPJ3pwAc+gmBgRA7wIF7LgrHH/z6M2R1
cGs9lKf02HXk1Dr1UAGcPwNWMnESZCgjik8bfopKvN0Bl0S/lGVyhqzjQMlLLoce
RN9CQbKPkbfl2H7WmMB4H1Rl5+DlW1dF0cfaUHOqiNaUOA6iK1P/5YCZyb94QRu+
F2MGAtxDz7JNvh3NITj4Fh+u91Fk9XZ62bHpbXlgoDMGm5JoeX98yRU19SsfnOdY
zWu6vjPA/TXV9SBUezjNdgSR+PpZyjUekJwaevJUFS411wgpysg96VWSMv+Pd1N/
rY5iWROoED96SfcfG2hYIToecToh9BCVwaYUjC99TsVpW/iBxj1e/4+YiNDM7bTz
Dbi+WLCi0clarGMX2eH033ovl69CqoT0W01IVIZ0KZPIjb24uvRq4w5NVoZeLdXn
jrq90R0QWmAohxmC21oKcX1Cr6tN6Yxw8s4eGUlHJA5idZXiKMunALSK6sUCv016
qand/GCQXDySJqI8T7lJ6wxaxvbZQpJu9xG6kvPhim+GrOhkvdmomZaz+fcFA29u
qE7EzCBjcjAtTLVoVSQdD3CtvmSf7rl0nlAWEDjFE+wHyGG+gMNr2gkSqL5JYmIi
pe0LxYE+vP3HISaBs95OvD+Juv9zuRMZV7kSieaOySdC3bLfYxwX8TwCogfGZNC1
ZpPJI04iMBalv5f7V9WZ1ogTwHVE0rYp6tKKcBEGcGlwa/IytYoPhTi9lNSk12ng
S365oyGrW5Iv1D4gVQhpOlZz//A/8rw1fbTUQMM3b/8gwVKJ1M/+K/8PUxI62Y27
Kf8tnvi/kK3h8pyukqvBxJH6MU3NRMinrtCSFTSpJKN6oK0yT+NyoWbBudXPGl9W
bHU5AF9nO1MN4p4CxoL9oz3/+oGUUJGVkyEG00I7vxzhyr0/iKiNEPlLuHhLsP7b
IJ6aaBSPsQmYkuCQn3l+oRUek+a9FmUSkP8pBGZsccv3rdq5DBw3kLI9uxcp6LYi
Y86JsDVx7OcDF3tu4Ps4xDkGDIOnWN9ft2rQwCsNzTE00j1yACpmGvdstGV8XuR6
xADMVWiS44NTo3vBu4YUOGpBki+vamDzSX4uqWoU20AgEzRKu+ji0ZwU4nm/ezFp
/FEzE6POrstDlEGoGvLQntb26hP/EHzeXf0QrbjEUujn7ial45lKplcR6uh971LS
lqeNIz2ruLIS3UYH5ZMoeIU0fLuJQifrshI8UXPpGB4iGSlhttmqBmFN73rTbTgF
DTQir9afcxFSbA6hewr5/190b6i5LxztfG6Mt4MSITnzPhqTTCVx3aqzN9L+e+/j
SvsUcmKS8FAIQZ2y8TARps1HVR1VddnJ9tIB62poWxsUDwY+8tGFVjcLuK+UTU9V
rnM7lW2ZgUx/231kQTWU4g2l5hj1WEEkMvLFo51egFy6arH8ubhcA66WlRa6y8ha
4E3c4wCKyH58NWR7RylGs+ZEu0rxDEpOsxanwBVvbYAkfMG2af9VqAkPZiy0BtcX
xWH3+RYRvIWVyPQB7LI+6zmh9+7mnOLppgvoMyGZdmWy29hYXKLCvxCLlXXUot6P
b8xpBFInHdeGVuZrdxvVfjm7zxBgkDsLrEpdtW4FxrzviWKCsNmkS80g+FzjojkM
E7yPat0AKhAKoiOvRAFlKHsc4FMtbu6Ey/OmM7lwbceDLGNOTA7AE4/mw3LD/Mbq
00rNYTUW/JD3QPMBm3dtk/jh2souAvLy0lRa70x8OpGRzHswaWaSsZPS60H1lfeX
cR3xibhHKvYQuJ/ttrAKltaB6PUPPG95Bt3KAkqqv47XurbvnaZ8ENNGNQgXWsRt
rtkWdYd6wqx9fq+mFaRZ2/a+/V8AeYTbM72sRjdDnYahMjrKj0YuvO14/axp5+Ni
z/lcZH3jniQpQY5V437PCw/ozKOl7QfzdobD3nt1FqMvj6ZPdMMkEAvTraiBwTuA
7CFkBoODP5xHmfLt109Buz4QTrbzzkwsPuKgSzMdusRyoVozO+dOkER06JYnEh4M
Tn142o+ppCyRVG5RPqvgeO3Lhks32qVpRmxgqxkYFZMEX3jT47EJmoOqlk1KRSMA
E6UzrXDNfs+Cnh43Uyeb8wZxpxYaQ93Tw9ZAXkkvMeWNkiOrnuPEcZe7bKq0N9Oj
Ef3rDo9xedFJqGWrACLNnWIit8vmRUx6q9fazdYCG5VMGiShXuwjSXBHX0q0nCb1
LxNscyckWpzobM9//5C88v2+FAt16yABObeBrUeDDH20cxTTFlyDuO3iaXESZP0L
p6pAmXDmNwzyiOzPTF/QEJ8HpxroYZsYNT2jMXL8faZxX5CyKkwkfiKn3kyT+vNS
XaP88zciv/+0RB/Pkr0Z8GzSRIVM4kfbz1dENI0ZezYGWjt2OBJvUVks80j5bEJI
2W+z5wIWxn2kxArHK9IWUvgTS0/fJ4enm0VeGMkFA0ej02tIh3uqfux7mPACjfvD
fslGPizOvmikiVz8ju/+4HqeUUPZVu9tYKLvRihk1f6dvejHOFQe4bwQXJUsRgLi
gHUbR/I0F44MzlEIU0kp5AZ23DtxwNfsHx9qI4s2flomLtrQxgxq6wl1QXNOEumz
prDn/nCBeknZ701w+KkvkXvi69JxopUIE63qi2jkpJ+MkMvAovKHYu3xW2sLlXyj
okcJGUzrwDKEp1Yf7Kh/IleiIEwH2sub14nAjZ1m52BlVy42RpnzUCW967hZUPYr
rNUa2Rn68rPSQYbQAwKfB+i0SA3MzZ2TgLkVIO84bl4Tx2t8Dqd9hXU0VPnKlQbI
d0N6tfcv32mpmVTEgsDnih7UyEZ7/qbuDXDlO/wxfvomYwgHGV0iJYtbp51Hupgh
DTq6Xsup4+EV9SpvWr6Ldh9cTA4PGpsbEw4QhmaRCoe+t6S0Vu1/+QH+9q7x013Q
T2rbADeCQkYIgjBjx55jnpadbJ8I7ptEGrIWn3QWyxzm6qPjkhoI3Z8ggV1so1Uk
VoXVpW4GicB2AGLjZlAtLvF89Z6nhtQoe/hJU6FEUIzrzvZAdYOX3au1zoODeWtj
oywSiTBpjXph3swpyBlzCxjxpdNj0d0OH+YwqN0IgN9KWYkC/hbEibZonPZSEpub
gKMdl0IB9DQ+EFAAjBgRW6hZ8QHBc9iSJ52u878viCdmDhL57eMtrqizcOoYgUg1
ZYpdYG4rSPP0gBXQoDESCBRFWPHekAjK3NYQgSqfOawkfSQlOWRPm3vEFp75SHIJ
SnJJIyVrorYp0Bfpn5iZihreODM/JNPDBnuWg/K3EiZ5fbOHJBKy5wX2GSDDegL8
YO/vGUgX4D55vOmcKeP6wzEG/oJoympBtPmiR9gCUj3rG6Z4yVMfEcNT3PUyglT0
B2cNVnQMp83c6HQyc/bXl3ek++022h9SbWalRSrHsA3BUTurduNdR+IFc33flldM
ql4q0Rbz7nJ4FdLFDXaLXBTxXAK/nsC7yZmAZLI+Hs0ahAcLrkQuOM9XRVdampC8
XO1XWEy5CHvApd4SijKzDc6kPDkjcWU4eYY8ko5j/Cz3MAJsaL6jCk1tl+F1+y50
qkhzUDUJqGsqRMrs8C02ewKmdBHxPrvzdpnpJnGaPsIm45zIYVeMUjYfEBX6Ti6t
z4a1VHoY7jj5/mpxD2TAXgF0N/1oPAajGC768XDoZ7vA9vxPPnQpgjz3TpF0zF5E
sauuaxpGz3m9RIEa1ShulkLPMZ/1P1dGwKGueZZsTsjXiDE6iWQNcYYBzBitkCfa
K5aMO+VSb6xakJlDXqCGt4s9N2EMvySlwKYGGCULIpc5amJiJX1QO4gVSn8N67xH
0+xGUFJSbZcYZMOs/YRC8Lj/steOUC3fyMUJWgvvBSgQmDmu3fGJ1z3D1px8WnHn
Yp5SgtYhXduOWxg/zCEAa82NLdg4qekBDPx0CsX2Cwh9gPN/OVYy60fFj7Jf6QbN
`protect END_PROTECTED
