`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GyefIzoDUlpAstmBshi3bITnxNO8F9nDJOPBHQDSP4S23/tpeSOL9F2I5nlw9RfC
CFqKNCEANGWb8OnlXYdsiUxOUEsOIuTeAvXMNzzUUaa+T48UyGkcYw6uQC88MW//
iclJ3H4WEDWkNOFTGplili+XobWxWfuHzMUWZGH7rIf8XSZ1vmrOO90vqpzDzfog
68BCQPEScfQWfhSOYvgojjepakrBj6UIQIC78RUe1yV00/TZJuSY4ONW+sWPzd9F
S0tCqf+HpA7V7OqF4gvqIdFH/g+U3td2Zkom9Dz9SBSq+iOpHzhndPUZjThdrok2
xspWDNcjFJUEXYmQ/vhd0bJPERFEndMj4iPY71Tj6EFb2DLtw5mQbs3Te1uKoo66
IopPLLRPMioCzwOIN583jNCK0shd7umZ+vefL2VaL/dmEf/zaJMWt3IhWqarfHXv
YYjxNHbuvloHGLY5kQbyMw1VcqV9vrw55BJncvZVYdN+OU5g8WZEg8uZyV4+y/AW
54ZS+igTbHCywf8mCKuzRDHt7xTHkKet6u2z+ZDaViX0IIl4iZZu615vO10h7LVX
Ziji1KCJQ+C73Q6QVLx+jUF1GkJBGAKhVY1tktKXS39JGQjCeLUkMsNJgVWHIEVN
GOkkG0c1igs1P7gOcLsMoYHnF4iBLTZ8jbiRkwYPkXOmftrr8jiqQTdO45F95gEg
PyC5rKWU3NIsjqIaDWtQE+fKafy9houGj/ndxOpymovfxPKHk/ZXEWr6gw1t/6xj
VkiOWvK5fuGwUFGxn8XlGkeqaAQjqjJ5zAZGeVjaiU/ZKCW9m1HTNQ9BCedMP1iL
CEAIZgjPqP3DW1JwPfYM5BPV4X2LafPeHTgZ0Cmfe5Ge3BvsbahCH13z3lCHLDkd
Fhwv7R8vU7KgGzd/1pPDsD5aY7fmUSEsl/p6mjoaT1kAERSz0zf2jXa40ZKrkZT/
UTTBfCJCBlEBe1gAYVnFNn2214gGaMFFu6rdaHQa8LqpBn81vTQtxMgh3/RzCKa9
2EoWlyUFedP7rFR0bh8Qbe2/M5z1UOmlZw7eTCCrraHH+D88hEDREB+sx/iJLELP
0wzUyCVU9UeUExCDJM9rj8Y0gYX4L5i2S8BlmQ7NAA32XEte1pNunFUzCXCyt6mk
lheHM5PF56yZ59DaryBimc/esjl2kzIZEiNkDY+BRQ3Q3KEEEofzECXMU+WD6WhZ
xVL4YCh1NvxKcsUF/jMe/xRMYmqmaUdN2+K5SIDpT16dkeYUOQMSsGXbYHiF35Gb
kizixViC2gbYszc9ac7snIjykgIOu7pnBmRVYCLMGlELZO1vLjt2b+/fCZ2esQIS
TGXtgqO663xTLojCJaq2a11e/XYx0lVOrZPTCOmsUHMw8xhBeT6Iz8QlCPRIObYf
siipetu/sWP1ScZ+u0QNQLYou21TA8UfgHsONcwS0eI4pqHkG11ClTvM3T6hhjH5
SreaCabc7m8xBsjtZ/KjO8NBNwpLjIR/I3RiO/sTFlKx5HU+9+S80dxEO677AuPX
3vwUnZixgl73v81rPV3kk1gypfpzSGPCQ8VuXHZmNwXwsDRnJZtX5GcM8Cnk9moF
rLsPiT+WS17uyiODM6bDsumpDryiPg6en5M7KXpSZgjxBFD7su6aMPAEisS5zygD
cRWpKJoLPWyX64flev3Osfg0A+j1SlMT9anV334lxjs1pB2YauKnIn7wHpxsL06Z
54aDGEvHN4p5wpNiPmRcUjsJqLyujdB9FS9NLvHNOURNq7X/lvQ0E2j/QN8hHFTE
pLnVg8MneTijRnoH8JRgTkWbcBzjvtyOyEvl9u07HYTnct8EcDcWPmaNvT39Se/B
5bTy7CdtLla37ZRck37lcJSvQz6GI6c18+nAwFQeWyL2+QS+3rCHMSKPzZepVsR5
K/XYV7cwC1v+xxihTt/QLQVdcO94IeDbug38D8ItLL5QANsaGzOlWUadSiKzt/GR
Kzbe+sVEVJimDDaIru6YlbvCPZWSClHaPt9BDWQ0gljV0j04Rn8huf9YaVsKnQsr
`protect END_PROTECTED
