`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efykrc1IMUNqCl7UvqmkgZD0CYiQSk5SXdtUElfzTUesPkCGoTZia9w5z68iLU+j
+54kkz2s/g5GukAmb+Z8PoD4sY64C2eHPDDX32himSgrIgkOfpOT8iCE5kxF109J
59Ng4KrIIwwPA0nO4VyI92vsfCS4DKAwAtzit7JRi10QGczruA5t/Hv0LzVoP/db
`protect END_PROTECTED
