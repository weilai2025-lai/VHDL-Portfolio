`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Dxwpn5TsbaGdMbQxfAP5579XpbsZF6Tk8m5jek/DEdiWC9nhDLyqKI3vOGVfG8y
QITynbCcxcF2iZhaFLMidPhY2zpfPVh2PqtKBzhMSaNdZjL02eGn3u6RQSma/Zmm
ZqI4JHFVZ8qPf7dm1f1Sx+UMimMNwc8mn3dSscUsf4dzpK53lyzZAvHHIIxc4iN2
fCncDr2Yl99FlZHZMiQctUWauCEYtKG9sR0Zn1qJVDLt3CxHTUXqr2/I318mfcBI
cacbPLfgd0zrRXy6j5IAK0ug9O1i4QDYYyWjXrHRZRzDB2JY2t/cGeJ7f8ob+Ycb
oqmYwUnJab57iUW42WuPssHeYPGhNSlc6UH3j7n3vRxT1wSjk28BcX8hSzH9vXIJ
1yenRHWX+E6SSNEa20i2uVh2f0K0dalKG9hGNHTunGO2eAfMfsA7ohwihnvtso0S
og9WEEs4nUTeuC1x9j9rpeFMumPEUThCS+Jrco4qRU3M/XiKYMvgbSvgncKxJtwV
UxPsZOCaIigKBEb8g3HX874Bq5dGnvnOKbmjktaOVa/C5K121WymGIFiMEtNGfA1
TOB4GXh7y4/VhpBMqEyXbag9H3WWZfVWCKntbo66zbB889olkCQBS2VJ6p0XXZw8
GWy3dTWFOmaSGCfP8GSm5O8RGSm2v3+imQkPEZJibuRtZXDSWd0tE5foonTlTYV/
Dp71tyZm9uYR9NpZ/Id0RF+leCyUL9ixEeC3ZlbOLweJ3H7AkWSORhbVwc0bn/Oe
uCjB08RWfsXNvEkv2lyG0ehKnqIVO08suURPuXtooeQMHfHhPus/Hw8tiAxqnJ/y
oD0gYsnynuojF01cPWa28O4CAYHabDAnw5VwuUyZd25Wlr/3sfvks0Fh4E972Lu3
wMbsNYZwiACpn+obVtMvXZfh6fCVzS+WRoqmfrI4UqwWrWav0pRa3sE3YIQ4z9Bl
CX/6fjEhjvnFA91Eu+Y0hJD90t7JhO8WNvBdo5QJ20Pd2f0mIPu5BX146fQJIlY2
Fc8XvZOVKShJ5n1v8FvXvmuQUZ4hkT5XqhvmI5wubIX7588vHwyrvNlriZ2a37Hf
SizI4de6gQ+sP2gUZcEF7e2FolNtgsZVn9iE1gXxEAkXRjxz6/OY+OPLo+jHV1Ze
z0OOh4UzkdDcgDu5b75MREs3grE8NnqigQ9IJkXiemOPdjfZgLN0eFNEctRVcCTP
OLrAwpO+C5kx3bUU7K5kWdjpr3wJcYGdlU2a7rT30nyzfYtrU9kBwbx7gR9+rirQ
W4RKmcaedHkdyD40JSFNhBiP98oJnopjAD7hB+J0mu1lT2aQLROlUujm93ccHYcc
V2Ias9RJ1IkBGzy39q53tKet95wOrySmFb7ycQ+HpvJn8bg3FMzsfAZ77BiMQwg3
FUOD0SKkZEl/wU8L26aCT1NHnHSnVRAOPjCVJ7RCw+M5Va/MEE2n1o/kiJQfKJ6+
aE6i10YoSJGN2jaMEdllfbUjJ+6mB/M3yPr8pnVY+Edz6LUvWBziz6Ulje9EQvtj
zuOr54OQSAvgpFPTcj5A6zqREFEgPpWgxIiLJ1n5JgVuW4JTPKJba9fPT5/UqPTo
WCtDw86zk0O9rY8DRLWl9yPFcHbN0/aeUKzQ69CqdNH0BXePhcuxJLcZXXoYAqqS
7K6fVcfl4A1Wocxcdk7Q49n7glQYlCC+rCdCTCeiUELUax6ZanLvTJc8FohBbw4t
`protect END_PROTECTED
