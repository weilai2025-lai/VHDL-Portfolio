`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbvbLxZyPeBM8rNXXCihjzBml6ylAUVaSCPA9anTjZaQomOidx8zVeBHNstGdlfZ
QfGNwt+kWmXZr1fG5g7YajHcMkmiCV4EsTMeqEeOKpY+RCKmCHVig5nSxK6lNxzt
kauabLQaMYU6WqNTaZ9Z4xrfMVFcnLFbVbNgXBt6SdLLoEtTtdtriC4b6xsAsdBI
w7qkLyuTqqFu/2mwQOjXmnrkEvsVMQeSej4igipT7f/dXm6sWh0g3ja1PopndWpf
KQ8X2CC9GoBrrlj2Q1YqrYLPbhvci/rgbqIEh/hKJfMxY7olxKN8OjpZV2J1SbX2
Tw6cVJQcFsqjnQAAlhUi1C57fwoi+WI3ZiF1Q5I/18F2Bx/hzSGsnLvWdV4MxUkz
YK/sEm5fwTFK0UNi5OWLfgFa6uQNZYpaek1NlI5HTIC/Xt+D5qrwNB3TU5p2OtDD
M2OZzGqIPvT6VuZgPQmzB5fUmbDTtklZREKhQIx1E6Zu6w6IHFv3dxBxEOxqB6Gf
p0Hm5MzA6Fu1c1+9ZhCfmFRFh4pql/9+9Yvy69Uuhrs9r0zqSgmphYhTFn6UFN1k
sNgoLdp556iSc5XZ5ermuGlRVmDv4VgLFr+u4uTpIDggGRbAGKN/c2QX4+FHe9IO
Kxx4GBoVrqbzY8yPgK0F4AJny8Qs+cii2pgIoCy1N33QzuyiVIfxc22k0Lk/71xK
CpNQVH37yufQgYbo4pP4Gdjd3XYJ26VBq9v9rU6FDVKqxWJkFzxdzv/3ifRy3Sku
nAj1N+2yxkQDXelbBqpe5sgLlf3pGdLGCtTR3CoBUhjn5CTT9xfu0wauT/mmeMBw
vSJ1L852h/y5tBeEisXTMerFEsabM9tAjm8Vn6o4+R0DiooPQTjX05FgExF7oC15
PX6vEcHP0MX6MF3gg0v8Y68fFS5/U42CJqVp1uRsnoL6QnzpX0Z9eaH8xCWQRaSA
aus6MJ2SxQuoyIQVEjYUICXzJgcwf61oMu5UH/GVnSzPTB/RYa0yj89zLWN81YMM
vDREJP/UQEgn5M8sfp84TsGmYezJKXpQPAxYVqlmiLF2eNgSX4FySNaLJUJQTYZJ
7OW6Kr4kljhYoIms91A0Myq4etLUGr9TN/dQ67yhPGV6WLQ8SoN675W50unPeg3S
HUb28Pcs8cvkTCEWJBhAUNGzC1auc9/TDG8kJzOeoNRFZkkO8zky4eqJqbIm2gqB
2oASRueztRJ//Lh9bW4k3e9FECB+o5V63vyerzQSke1hZZhgcD66AQVzArO8yn8E
qAfUh5OpmVgdcurwS0iyOQF0W04dHVBsTQiVztpy9JbGXOf7hxbOzcY80wQck+9f
VVqH/zG9DwKZp3RI4RfpA2zoUpkdfPj6lfOr+7wAnbSUi6Zc9Nl9c/CNdoyZQmPA
sgcFP4mjR7WBvAhl7/mnd+i9j5cGYXM/VsSMPbhbRPZtD7k7YB8xj9a/MFgMX2WZ
rkWDBpgv/2prOE9OBidbwfa0C1i6nLAFIlP5Owa+X48havEKwKNgKE/qW9IW0Dxs
0PHcfSlH0OEN/znx0pM44rkCr3HivFQaR2t8g5mqdAroK7sT9Rtph83AN70144aM
2el+bCgoxDrjtxIHkfiW7sUJkUyr9ADXQWBsxOLpPWmjhqy7dcREzWqBYsIQM+Po
6cGXAOz/vfvroM7K0AngmCY9PtwyWpw+SZ7H3sBu7isJBklUwg4Qh5ECVBeYWn8t
yZYJB9DDVvN2POTgwIOemmtppipureCzonRADSJ76RWjn+k4lBKWPFSMetlB1hsa
f37njWmyHgFkGjGM9fALkUgzTdaCRJE1veARW/KzVKZ7EmBty6pw9v8x10wysva5
wYZ/sWPGEQKIMtkVM1cnDT0UZr1xtwKD3OYCdg3pXFcJdLhKg9CR7aMTHt/9rIZK
gDFhUjQlTO7xaU8iAefeq/lQ5qGbKIWPrIweJLIF52px6v0lc9TI8MKajjLok14q
W8kBcfkVjMalNZflqCoy/jWgx2BjhnByMZbDWIyxFHwiU7epKpR35mAUYLsbijhW
8c3oK0y5CGVfPrdLbt+ZBPTkSFs3sHQbpZp/mfaOplhY1twdo50Q+405u6UqTEnx
JBxD/iCrkXxQmouPuPAiRdK2kpBoAZ2MDT+ksi+cW7xtcwTzpMQMRleOB9Iw7p/E
GkBu7F1TQBbofoZihNWNslYQLxmM+j8rOqYJvxlosoBpNKDFdORIxPbjJl4FustJ
VJsAsZ6vvERQ7/KV5QFrktwOWZG4/7vVgmRb2EyicWpG6xsgDE49IvoFnFF/ugjT
QywZqe6sLEfO6ULFHIqJ+HAmCCwEgsqKqgVAnumjIGIX49YpkYY4l+Tu1iw6auTP
o+IDd147Dz+tpXV5WP0bMCWr+p/zLsuff/2El4TF8BgTbNW4B7zaeqN0I3qJEJrV
VssH0gL4G31Bf9Vd0/X/HCbRXBr6L5W/map0logrIEA0irNrl72nvkjmNNOE6N/C
CSEKR/SUYnt8g5vowWxEdstLUsdWmritJfw6puT46EAnYJcjYQEajS+igXZpf3td
jB3seRL53v6GHML7uinvuiO9+m1ETVBi3ND/UemxEshBIFNIKTK9YCVN56nfARCO
/oTfmjOBBMlr8Nx+atXoAr3DpkntBZLn+Tiq+QuvRLpU7LcKOdQIdt5f6N6+3so7
mozwpuMQzXhZu7SYZiR564RX/6ibxb7wQpk64lIlGMQ/gp5Jn4DfSYibgxdopCtz
BG26gsOgjVJFEqoqHywDaWdFpTNWy7gR3YFTNH3sUWWZxqO8txvpM8ajLrX+li94
mUhb34kM2deJ4T78FvNMl47altqYGY+Nyr+ejlnWXO6eJnsrn63Qw7HFxaTqAZI3
LiVhah0ajBEKb4UhmtwhyLAQLh2UA/LfylEU4jvmUvREHWr8wHWeLJA2CPbpWfUl
4a+JnSDTHlet6qNbncbsNFUOU7HkeqAJlJ/7npI/DXQ6r+iQAWPTRD+0cVT2AAsq
Pp/4BZe1jodQ2IHo7pPc9ZNADjlLZl7bTJY1RH1ZoOItn90CC0mpY0X0hq1qV3o2
bSDET59nPQk9zFP60FgX7TceWHnVSObKnln5hL5FDWl4Me6B9G1+xHH0o2a+NQB1
8Fqjfeu6G7WiU/LtMFJ1MfK39BcOpq8vlQ8OgxDzODjJCPBOcJeTy0UAmmaX280L
mfVeptnHGw0RzkvCtiPx43/H9xCG+arG61hiWqmnX+sqAywrIQuPA8yhTyEpzX6h
VLSvfCQJvZLFnY6z+lN9W1g00TuYqWmcV8K6felwsf3cfqZfkWdCLA4AoTiwZqII
Cet/8iX8oZZclxkfCp3AoC1sgF5mk0An0x2cUKOddyHv60goIZSMmcj8lKwX7opR
yaBWOwmUH0HsL4XGUVuNLuCuegE3ziXlv4m1J1cu/WHr2GI1F7efzgKf7sb1V2I0
Rws2hkDNev681TucgfL6H4zNpjGhGpBdqtZ4B9EYduqYcAV9IhLXljz7hd6Ch0yJ
3ipIhIOvzHDRwt/OlWemSSc8wXxVgbSxZ+wZWEXqtMaQKHX38wwlfD+xBaXn1sY8
PonxhLzFC90mTdqbLRP7l7ML7s3k+cdNqjhd5G5pp6jDJ5iCm8OGAPbitTPD2nmM
n/1DX3tV71SS4AtM1c3qeAvyxTgOkUw/DtOMLnao14XAHINcKpgklL/VQXc/St1C
n7CJYVXQLUqaJ9Gv5b02zZVOb4yzB3bv2TCLfIHT2Kp+Rgq03cbd0kjEkCQ0qsyu
V1RrwZBUukoR3Ui6qYl/knRGLPkU1B0PgynyisTBgmWFgEcvcY8XGxut2i8m7P0b
G6NJBL38tiX8DiFm9yxJk0/lFT8aGv/g79FC2MObYQiX/YGrVLI1u7L9m1fncJHr
0foXJlTLGQhblkZapkxvtbSdowlpLZOntKzOh43SaoYBwGds1XiyT058V3lu1rBq
P0BkVr54b3MJ2W34r/IMgyGGLHRDVK8y11wpQU9dCmi7YfcWY20I/juiMUewpT9D
dmtIb+yH0L8IuUd58WEdyjh+pcP1qdWhgIcVnnXRS7CtxPnDpXcXTGyKB4fhMqAj
BMBDgsVZZ+vI0VVi/e4LDSjyOXkjLk18KfowQFT0prAAIrf9hUOaPW1knCJ9H8a6
RkUmJld1bd+jw+CehvRfbjuBat9y3D+Er116WEnbcUS0/jyaTNXoLdPiySfEc7LH
UPTujeHy7xKlHT2TKlNmyfUNSp4So4vYq8ugyHk298BMeXm47Hq0o0EWXy+zHsRr
uUrejg+Kbv26QnupjehIZyEVaR/V/VXKxID1P4z1ZXNUjWu/vJPs97cjjsEB1wTR
M741ThdT70z1w5MXgZLvuboix0zGEGRE9WoxXsdf4GVvXTweE/nQvXlyOLoKYwZJ
9AP/7kNG1bOQLRm0eYXwYV8T0ihZHK9CbJb537uSMGgJaRLgYf1Q9/flL20T/ouc
2HJcprsuyTWmWc3pC45YfK3fcTOFMmOL45tj/nUhCMkuTTYB6QYGD3O4INs26gXY
3niFMadmL/K2fPy6TQgvnlcdi//cIyjU0631XydbA5nWdGR+SoS3z2gG/6627+kV
BGcivc1/PUZBxqKIGDh5tKgsDglo9UbCFJ3k/7ssLG/wcmutTB1lgW4se+uW+wgb
4+Dv2Nm7QX0mbAqE5HbKZ/FqUOHT+l8Hhg8kv6Zmv9UYv3hPkLTG+GPu14nSswiu
8a/JAnlWzvBnLIIoUPHK+gHZHtJ5pkY1wIacAAziwOVuWGlOC9htu3WtlOgN2qiu
+xwgTL9illmJoDzyVvXBFL8tTKfegqeu/WC8RvoVuZH2eRnNLEGHVVlTNSZZYiEM
8UHXj1wwSdIwhFWKvrlEe8Vy3JG/V0rIl2RrAH1yO+NHH+QIfp8rxRthAyjnhZMx
knJl/iIBUpPvPm8rOqWB5Kxpl/S6auI2dgP3LAJC6AeZFe48fqjZgPqTWMFAzUvk
7IDmLoL1Fbm6zHzZALKqQQIx/L8cPHXQak/euIZxnf54d1GSpYpbh+otcScERrF4
Q1rc2QXHVxQ5cSGGXSNzHAutdPLkWXRofhI/1q2a0BilzA3jJuUGUughuqbiFA/D
MajxdTfqze3bPs2bHeQfnUIxb+UxQkQRuY8z2eZDH2Pk9CnTiqo4heLYp7+CNGvY
PTOHuhUVR4r0ykNnP84HcqvQe84AC3AEX2D5gwpuIShObxigk0DhYFzvKBpnovaz
CoprH34thLOg6AfH/aGV6TsiLBWaY+OSWEjkC/nU4rgPR86aL4jmDeQ2eepBdmIY
PmSJ3yvY3qzicv4F+E7u3vhwOgR2NinP8/irKDmbosGwkJIdGIgIU2OjRXvsiDHS
vzPXBB3QQc9U6e8bag+wXMi/mJptwEc8zkACAlBe4fAZW09wB+ta5FgKUjpydq9r
YoWAXWd1cbuBUctoWcSAaMMNATgwR5KmKi+FFgrkeveXLM+NK2M3vGKUmhCIaSXz
LCeVCeeIIpW5sWWr9HMbI2m9jXJmUmd0JsAidaebgTOZFQ3XRKgytxbK3rZ6nyYR
H4CYS7WbxhusoFYXD9FMcYYuZQIWOwhb3hFqEGVzWVBfojGo94LFV+T5wLaGpEdn
mVfdyLi02G9fBkiPlc38Y20sC8I1L4x9NJ1L7pQsm5Pr9k3+bk6QIN+RcXABSGbH
DuDgF20QSIGAzn9PTyFswH0EOBsc0BxSN7iiVzu9MI1IvBuudnhjHMJ1Y+qzopsM
5JWNa4aksRJTAilrlsaCr3G0OFzzyBDJExsT1U8UfiVAVLXO3sW7f5QIOIKOvPLI
zfeXhxBPltnMNcI6Fg5HZmOZBhyzO6V9PKwt7SJP5x8oqsMMAjR414kHEdK6OUyg
HfH+jzRodYbECb7q65yiL3t8sTHUe8lyQfwpnIGCyx/1dTNwqvyoZ994IVY6hDrh
GtjRshgpjGlgWb8CnfwAaKJGQhAuQJxifDwYYRCHjlx2d2juPZ7FXZOpU9bNtWUP
KEpunmV3RcUAOzjHV2DWwX5jR8/Pt0rnsGsAmWrEnfBjjaoZGEEWbSNSNrojy4Xq
D5jwYInd+rQR3h31G8xbcWZ5xe5jPEUXRxY2Cd4T1FYL34Be0sHK05EVpzM1pLvV
HtXzJrfoNvw2l+kBEZXOxYnBmAbDKbD0D9fd5fR27dVMQ2oq2WGzCrI72L9MAYT/
ZUu/+PPekKC2s7yAyVZHQ2Zjk+yyADn43P2J+D9fM/vB6Fb4ZgUIxcBlyhUj3Jzk
zGGqwyUaJkcGVBuPjHfpz1MV5tOuUOncchsZLlcCI2ue1XPSL0lj0J8ayQxGXjTE
YCYasSYa5/GhWXIpUKtLH2oCkWuHNyKPUZVlznG0R8Maj3g6DOGALRqyS/QYM4BY
yLdFaZHtZR5xThoLp+pr2cnKJPOMfS59kPvmqxUowMpv40p/vlcSzHkejtGeNjgg
JVgZi5AE0sxUtmWJcxjYdmY7hkpwV+bpyCmeCSMUJKS0ZKSx7Mb3vwhmTWuVY1pD
qbstaIvJ73G2As6gZO029o8e82HyXePlXOyYDkSVaULhVXOym8cMu0ZX++EsXIAd
Hc92seIdaUIomjXl0rzJVz0Jwu+UH0ONUy8RylrVc29Kzyn685pskgf34J+h3rCo
mbQe6+VFk9m31uheFlK0s7wvVm0RNKEkAPzroAq0EfFkRbvjRVBuo0+omBqqZ0Ui
wBmozfkplmAO0fhdhFwTlfrFD1MXTCwZTKjtkBo1pkGf5vIUQxAOFoJ+QMA7C2ab
fguOjxCFv4nYTacvxiGC619Qfl9CZUtTqh5giBea8u1G++219RAD8P1bsOK4yIoD
Jo0PtWwepnFHb9FJshb79e/R7T+8nu/ZZdCqMXHweF0w/ErGcMeeWRID6Ei+coH0
R9on/gHNf2B8eYPfguY0Ag66TVXBYinu1LTh2VkWUhRtSni3lZlIYPLXUqLZ4LWA
JDCoTDAUJQ5sazPP2TBLw3+lOnCCtvDBoVu4Q6lT6aWZESiK0OGld9za5K1UmugP
zwnFzojkGEKvP4IKSBm6VaQoWhzzpn84pff9YFrCKufXH5yNrJsYxsUN/c2v9bVO
FndeLJrvRTYVWVT83/LeFUbUx3l5zhFGcR9pCudS+Ikkw+sJZwF0QAXaA4nErfTt
XTBDZMAP2bpLrrWbfq6udUhqRp0AjUQA1z5B8u7E8tLnl6C+5neCHXBuFNNY3GWA
maTpM4yG0Yz2dl2qd27LEC9a7wvL2CrOOI9aCxaf8BbZn/2Y0P+UpT83dtBKrBac
aiWBYOWLwgp0c/LitUsoUlTQU14E8Nw3+GoCPNJbHuqXxH7qZpKimc7a35nwb+VX
6dHoXb5WZDrnzc+KDSWfSOq2YXX0GBsXBC8De5a4JjedzH7FdEjGJ9lApWlPboX3
OV/BzxPmw/hLNMAVBHLOXL9gBryaHoWagog+GkGSdsmrSGquu8Ru192W7v6OKjJD
5Re8DVkfn4CHYpHDs9faXYEizRIucXoAuq+1YI+/K14ul23xEhNv2dyczV0/ayoK
xJe/NzQjwgFrLpK3u9iPvEsI5yPAiwfuZArgqPiF2cOIawWrVM4htcAlAAyHeS2E
X5NN1V2fwCPUbWpmzC+MvciFntoC4r+TyJZo98mIoidhKMc7v/wslQuHhrZ/UKHT
GO1F9lGqFjq4O2UTTsMnfJoAjwFSL8xFKoCdwoFejCKMrmC0cqssd5O3haWZJ+DW
wdFlPEob6gE5D+wnzCpRkQKx5GTEh2e/RHcQa+MA17ARMcj7iKndM+v5okM1DFxx
bdgiBvle6wwtOQJYol1Tqsmkjso9zVq7lGsG2ELqQhwiL3AdrjK0Kqt8pWxFuui/
N1Y95e99FEdpIlh9KdQSqJw8/c0ZGNXhKMLGtYvxMi43nVQKSDLTpAqt1J8K8vKt
XSMuPgwyp/MPd9CWQoIohfmGJ3+lVNot+o6mWvIo2rlmwV1tooLrccMmR3mVSoLJ
AYkvg9JWRUmYwJKHMyZLc0MuCWu7m4eKagYxuFdTid/9ooPj6w12455YsR/fVENT
LAFNy1zBehIinI5gAkEA35Hz8U6e5gq6P28vSBfFrDcvQg95feirX+dC5PieaZgx
kXuoRUeEtPZ5B7WyBmWIprGrT1G+zX1Dj2mvgExcd3fuuv37IiZOblJO8j8RKaq7
3Zck/SnEXewGjxIdduuS1zFJZviLqlOfxYdImKBXskZZjPvh/rE5vn8jUHSENOHC
m7IRDKvuPOysd721pKe1exe4kniQeQUAhskjUWIhAeyQSIGCmZH1l6GcnTSx0Ksm
9kwSEEqulfLnFgMqaD6b3Ysu2Qowj6MTSD0wkukm/bG4gRiRecNP87QCQp3trlrm
Wjh6DOr98qDdH0ncWvU4O8FqzActtiIzreKntewRxTJbH2E8fptyJod8qHT6QBtJ
E8x3/KXFUcpR6EBObiRvkWvEGmgKtE/JYimWRI76pzyblETFePLgTsvUuQs7BC0S
UcxtGZXgrhoceflJIIDk9sJNTXGmrgfFFxxmbwbf/S7e6DzS6z3XRhyz38L40PwC
YewLhubHnBWH2DTYt6S7lmMySkZ2hWNLdds+k+ZLlJnhTMXLk5T2e5MH67SMOK24
YnNI1fxDn3tGeisaptaZLz2UjJ7os135T/QZVbM8ZoOsXosy5hZvuOYxGifZAc3X
ndSBcLnfjiMUJv8Z82gcIdLWhN3HITqaJLDY5d9DxD+qn9tWkZEkZaF0FW9+yDs6
7NVn2e1CYQGwq8iJ08PICvVpPpGPweQwN95GHoGptKk43sD6hILqeLR39bCLEJ2s
RWwYYmt1He0TIh5eFc/nKdxS5zEKzeb+3xFZaYVRmR5TOVoR9XekcIX2CWZNRg/C
PuHZIZfiAQps4+ObrZ2LlyMyDhaBgYHfOhR1xZOehoZ/CEgyDZdloNq2gZQH5jXs
I55+vt+AbatjUvzcP+6Ds8wEf3xFy6fAFS/47rH2OpFmEqFqeYu9QG1FbSKxrvI3
o2tvXj3/B8ZiMqtZNPf128jFohaKoov68slWuCbYNEvyNXl2GHBaIWGjPOkCHenB
eiV36bXNt42yziyL/psVOqsMpTRzFaGYjVpBKbRwunsahHL/vn3xrTO7CP3EiTZh
b2KQKlJk+jTEFqOmaxLzohfjWN+8zl6aMlLHF25PCiT6xY7pxyiKPKN8UOYK/kHX
wc+vvgx5LPBTtu61hmw44/DAddzmRy7GiAC8yzY8udMjNJWvU/vfdJ0KOrpoL4rZ
orGetkNhbbB751nlITD0+Ohw94tuZonst8xcZBCDndIJan/I2JAAfabeacIRjGYV
qCkNyOz0bv5Xczy0diW3aeRBxSfqM3OTB71ITQHPv6O4P7V3oXVM17dXHUR1cTKF
hO1Ko+omPQqlmieXiwoM3OWh5jtyCpr1i3R47kOoscD8ZTBpZAd0Xa1n3ez0eRaB
37hhZenLH4FbTcJojs7q1cjJ9Yd4O+oQ+AB1rzFjkBiep/7SYNhwZD5ZoY7kUtAa
DqVHVQWC/wZDqKY1pC8Jmx5pIYzS3pBNURaxQWwLOjntF7hUIzEngl359kygPkfL
ZGzdNvJXF1ah41JB/3pcO/lKQ76nPQu/xNYq1OXm86E2S6lvFEuaYIHswiDrnTvr
Sslb6t2lqOdfjz0cliyqX5UmE55kVkcz4ouArChzHC3M1N9KIAp31i+hRw7PcHEY
QD+1p7pmNECYLMVhw+zS9vWvLC7siNwnUQo5UbVmhhfpFheZdV6va6aMRPpj29wg
+Zi9d4/cR3OrouNXvkxu/iWQH2otGoHhdp/zjTrDBiWBGI7XFy0EC/2S6wBHmdVG
eg8Dw5Rl01oJpPVPOKmIb5vRNxx2cBOnIplr8Avq0JZzJDF7O4mxZPzJmq19RTY7
Y9zvwUlfg1pR+1fc7yES5BOy+oeTsBiXKnlTCQxWXi5KL1ittZ1Yp1gWYI3KfIJk
s1SVYozIZLq+gBfkqmR46OfTWEX/3NP+Mf+3euXRvnH2yxIhVpbKeAuWAy5VG6WD
59/L8LlZclwbT7eYuS12VlyxlDPbydWvuxa/z9PZrdf/Aj2P5Bfb3lIamS6dJvOt
9OHksnrIJV6n2gpLXuBXVZ7d7o+687iaREm+1H3GSAhw4DAXZ0KlfwLl/Qlo59qy
y74U5XYyoVemVgLUMXfTQV5Ts3A2+dj8KWYgzEGvo77EJ9f3YXsgJbmcGsosnhxw
yngohExI/RJkmfCEXrEWJ+pTrRiqrdfCWx+dID5jwCWq07Ug5UAnTDLdE4KFgc6T
tvWhuOZdzKiK7AdxGhubdmGBkE0Tf4kzdz1wOgEL/2BgYXCqzAn+8LGFxFBdNKMJ
nFZBjJHlQmc32makmuJkMASSPltDE4dIgYH8UblsMbPg8ePuvsVYcZZM3wxn0iD8
9Fxl83ByQmZiodH67PCJuCR0wIphumA0LslkIfKGCSsm2RSma6lFO0s78tWHJYcK
2EGdvA3oya69xDWbtO7Dnf7m7t83pAgP1ot5X8d7O45tOUmCW28kmXadmQ7W/Qwv
nRNUDKoEa8K5nWv8U5YUIXZsKJiqivTp6RgurnGEg6Ad7P7JEfVCIQj88rBkQxf/
h/5HQySRImdo2IKUrogS67/MSRxgTU7Az9AiYjdnD6zlUI/oBYH5v+TBGLmIwyfF
6Btu6MMZln15jhkZpxMcYMc0AALJc3YCDTFEF0XqyGq71IKRtovlpwTeUeGK1Gni
+kRL9Ug2A8ItThKfAqXwZNH+J6lXQ08I9465URcbqqzUw+iJUp3Xko2Vk7KBcezT
5aOgzoQ2tdsyb9UsbMvfKzZ6t+/0wSNKsRXxD7C8ACg71bb1fBxrZv2KjQy6quk5
hdM2FCBJ03rXnr25J4NdEK/9Zs0YtX+QX4hM1ScOXAASisSXgLctCDctle1XMjjo
zqB3ZdBlHMaNgOBRl5rxW6y4gOvWRNQOzrdFiAJGhYXTDGS9KLPUK1EvIdOQgbLF
937WqAbx6fAZUTw3cgc2L3536RCHpGEnRimFDOJJiL4clBcdNlm3HrwDOHiX6DiD
+E0UaPF2KfitLux8mQOOzuYxuqcaDVzhxAkIj70fPJ/BFRMEjiptUL+z5STFeB2j
7JRZ47MwjIWrT7JROaLEwh5UVfljctiFvNdItKrBqbqLF0WqwxK2uwAfIRu5C5m0
zUQFdE+HlcYImHOlCYrT39+8t0uimCi29c3vH/dgK4sQANQ9b+EPqR1gMq8x+/dK
+x46NoSKuEuTQBQdwMwK3LOkvbTAQdK43jRAtb8xVZGKV2bz1YtGBwealSLzRTX1
HCtoSPL57QIaNA4Ty9FWzyZ1iKu/3Jd5x8Z5nPAbRvBrtJAfryWNOqDZsWmFWcCh
M8S7Aig89ICCmjzHSykcr6EnMecHiNtwR0SxMdQeLeorbnYfrIDH/Ea+JPa6EwZd
GGF+GkJUfCzoHfweRwELcxQxo0H2XSUKOv5IT3D3/gOVqo+cEskPYp+QpRvgkzTO
aCw/lTj2S4ThAl8VIsNSKbNZVKV59xOzztiEq0KD7U9iGkW8jCpMdkBRiXkohKFD
8ZjaAVv1tZ1FICNRZtyobW5jrqAncL3lAji27RjSbR9Xs2TSfZgYpyfK9MUg1DEZ
5yczycM/WKNooiX1XLTbSiyGBGeF5qTKkD8GBQs2lPc+BDv7AEQ9mf4kUvU5b4Tl
pD1gL61O1tAkzHjwI9mQ6+wK44ATlcnBKY1NOWBpzyxG67q6GS2V6AwEmzqvVQqZ
sAncaZx2egAdoB1KtlWqrIypz1Qnj4uYOoFzohCjCgSSYnERcmvH8Wa2B61xhEuB
pLowSGvQ6A2pHgTJNGOELonQJqEjNiZeLFORbLLLwY0mJaYCJtlHXj0niQkO/S/I
8de+HYYIRj+0zZuhWrdRoIaaou2oeCpI9bCtoKSuThewhArSEHiOLCRbIFR99lSS
P08BbUVoMt+fq8w7YDMmq1XSIo4fINoda1JFE/RwAvD7vZRrxGHD7KoEfk666QbQ
QWtn8FH3Og4VnOKFq5W9vNhILqpxGnFCvhZg7QVdpddT1j5XK3LRU8Z5Zt1m0my2
+3vafg45zNC1bC8Km8JWkyVRvuZf6i03NZwNx+bZMavgv96V/o5AX92+OgUVkEiM
V5pE3n5IOAiQ3ga9uz6ZDVLkY8HBMoSEmuMeKxuA1lmCEGz2cOi6r5Nx/ziqrdCm
WASmab9drRek/p8b78rJwNVC+cnYu0VqserIhacY2kIefEDD6CWdYoYmq1sKsLfy
6O/p848w+SpGhqHrWn/fDQ+L8ojaqkxUNyiss+B0+hf1lxfzQ5LSDR5iD4oX0fgP
zg4qi8733jVbAuwD3wpa9cMN4Ummvr2QMn4WW00ePuapp011X0wQGlHGcpkopI8z
YcLymgNWbGbGYVxtBTNCRa1dZWKWZD2I2Jow4g5/g6GubIeZG+03LrNXiSuyaGCU
hn4f/HrQ0TxS9rFqJ3Rp8WB9EdTAom8LMXGV0DxVMehL53YHjZCQHcNY4rpIIbHO
gy0b6wwgsWsk+k8tRlwRngy3v6WlGwnqXsOhhiWL5JjeGklOEIghzs1r+/8B0lCU
I9QN9SEimd3RSJjFBxTPbgplvqwfwyk8jHWGDiWQEPNvrR3FZOA1LaNYEhceMIS0
sFfBFLIN0kP0FjkAdc0ihmMLTss630VHChnwb4amFixkBcUh48fDATyuJ/grVs2+
huer452SkkaQQH0APff6rH+uTzXw8IXkmxvq1D5mk2I0qj34gbRwt/lji2f6VEKu
Unl8DJWs7aeGN4s6OHpaQPBMQKs3CVHqUR3xvW22Su0Z1B39GEh98BLUNPHyQn7q
fNHKTNdXKKf2aWqOYK9/iMLDVMg48+z2mJFDPJZkSZMVMTkQajkTj3+L04HluARE
o0Cu2neyZtuuyrDUs9/+X1qrBzck9U6Dp6edl/bwJ4bsMAXI1jPnjZ3hZ8igAzJa
zMM4PR9vbok9icinkNPKy+foMHZQq7AO8G2j38z8/nu1yhjQMNoW1smcLEu1oAkz
+INNIn2wZry/dus2SKYe+wgiOt/QhQqkniN76fmEWBokp2WJpLEvnksfG640d6WM
f9ERHnofMOuk1NQCv1iZnj8ru6/eIL7lwOKRxx8QihgyDU45zRHXguLsogp58N7l
XNWB0zX5yQQczaC5PxzuQ8OUwLP8RclpwPsOLv2rtduIXf+dtRjxNGAhz2fCMVAD
G6xqAcdyFE+QJ8VC/FDp4GaPIXiWB25rAiydO/jXKr7tRklgErnZ0WGrVaO0RfUj
p6/4ehPEgA7tKSIOjs6tP23usPmw40dnSQqCs+256sHTvDZ1KEJfwq+gK0Kf+Uzv
zhiKWY6QH30eAKA4jTRfJoMqGqk2I6ahIl8GcWYxzZeDCTh0XtQxv7h3/z8wAWpf
Szbfurer4727ky0NxCTE3f494wOPkWUYZy/zokg8FGVDm4aYzEUdZh2Hf3pnLLP8
lk/Wnn2UoUV6eD579N34zEh/KnFOf9JJlSsYd9IpRCvIXdyZc2Xh5YbE3WAPL18n
Zpgf+JMhF45fmqww5ciQXB1Opxbig2puIcJRDJ2abfgT4c8AYdahu8/pMuP6BpFA
oKW39o21QLvcfScToWufneIyI5+UuK6ZffCP5+DY0Yz3vOp6n3qutoxPVmuE2Oo+
AlHQnOGPADjjGYnStj3oPLodssPWdPu51EVc9dr4AMTn+HYTapQlL4Plg/asJFhK
rxsq9B7x6eOGnqTCXkeoWwijOt4TRzHWrUiU+IBDg65Fsx0b35KH9FGI3jzqiDzg
4aDx8VAt3kmVq6MJzIdr3+I+Z8vYekospfXU42GmkSznadH9P5QfNv0HcMu0AZ4I
GVUCh0rfQpEmHQS5ZFmkqV/AK6ztet32KcFUoil3wvk7nEbJxUQ07GVqTytlBPvf
oytsa/eYlNt9ByDp3g0WHFnoGdTrtlRmppKSeHdkOOzbin0XZvNMP7UR8tgGJxR2
0bpcfdZVnB1u0hVSJPC1d0pdRMd3lquqgpyimpjy3pGO9HQJdyV9oRgZXCyzLjZT
TwRaY+dzQKAPbLe7CNFUagFgxitINYdFrBdgNTocqvPJIooFUo8WVIZM2hCTgMAJ
wi8Z57Uj0oKwmzv54Xy20+IjDDjL6bxKmRtbbrHNlQwjR2J68hUi6FyYdr6W/Vf6
BIq92DqTAzGALWLS5wIW+EJybjaILrEbIrsJvxPNPnehYqUc819Rj7pLPZSima7F
sR6oqwqkLygrbLV/oJiq1FJ2zowf825AhuFCWtnxMbDiwVQCQL2FBLwOQuQUd/80
BQI4/XVsLVL0Z1oYYUyqkG3TT+xeWr8onlUFbZEtBO0kxxSfLcUIiJM4/BG9m5+o
77NFTzyDyY3OTVwtywgcSvopshtTSoJRvC+FLSKLz9H1iz+UEAR4wq0kIUthwksa
PuIjpP4yLAp5WpO7uhXCM1RZ19tF9IrCvoV/00oCVUTYoQyhOTSjdHMYddgmjuqx
uC0uz+6/JdjqbYF8Zm3yESZqIVbvv/8vTj4L59wJaJVyhkm4zegnZYot25u34tO/
XN6+ilBhgiGJFDidnGCKxFQ6n86HwNl9KDAkVKq6UPLYqXW7qiv3sRRIxgiL7mMw
5eCwMJ2uleyArNAD1ZYm58vsT1OaCS8Dai7XJYx1Sqy5sd8ehNnn673RbDLDOjCf
9J2UhHeBppJwnT+wiCvmzPGH/JfTfMcaBP1B7zaairmKn71e23HrY0w0UnA4Zjpn
FsDIL2luyy8DXodvRPALEHeGoo1IEIRbmWh0ViJurrN6Uf8w+nc7t8QWXLpkFmc7
ILZSLUWIfilVyudP66t3FAFjKs++BgembgcU0ATBzFXiFdTxCM1KvpNj9vKgCdX5
PBa0jaFDuoXR6rPcW2JBI3SmZkl42D2wFwdpBglzcL3beMjYCioypuNad2ua3xaI
aoG6z3p80KC4d7/sHD9ULx8PVb78Rc+dZH9d9dhDf3y4XAY1XIeKYRpa2bpTgCfO
uZxmKyOff0ft/o/6W9tFV4NVRsaBVB4UGyhG1KPQCPXniOosIGcqbGQTVqU/dEjM
6rC4bF9mUTQKf7Y3TPUPNNjL0KyMEat+IP3h+VofrrZxm17jJB8p/n7IkhnGE24H
jH3Bz8+tLBohsd4EXQK6H/9QmQp5mhM5tLFuCiMphw1biUtdaENCVTo/e2f9Fr68
kA/xOCD0UlMEkEhAN34Qj5yMd5V18n6E3Hm5HqszvtmleqPhdYc0TqhfNtzF3nvi
Fl7jbh03338G61eSZViYSlFAvQ+9BE+J5lfFcLWLC4ImGVcqH3F3K2ZUPAnKHkhh
DtlZfznTgd8YWceOgmB+6yDR4XDejyVONktgNuUyLQQU8pBhSokKTEwSYJ2JJCvZ
97+vf6O87X4NIC+k/+W5Z+PCSqsYmM2ZUinDiUhZbB5ufAzW8Gwf2wKjNgJKJ4s8
6jP1ET9M6Y6Ysf/A9hYsNyMOERvsXEKHxJrCMHSKpQ/tovf+2Ra43YOtk5xKszH/
rZDElz28K/+yJsV2uGyLtbBPMB8HbWLxNUX4Tag3S0bWfm1DNY6e9rhGVVApv08D
3M9uL+ZKEPGrg6a+ERcRgCLKFfTR7LDaPAkrDPaiQ3sAefFmMnK85yuez+oOoBKP
R5X0P8r/K/yXBZGp7nitvHG/ezD8zMKQT74ukPhQlNaU3J37jdo6Cpym/28AFPAQ
PkGB2/Abqmf4kObxCVKIc6lDTbBF80TzaiODB2ozU8wdrdbQRCeaUuKUlnNCq7iH
NsZvn5RmFGM20vThmx7sbpk8BmASW3wK0kNq8iQoEETOZoecfkanxhYQ611oF5sv
L6bWgRJBoPOMnUOC+eYLgbo2Kav5jCrOm1I9uUlU48JyVFMP91DHetVAj+HIVNs0
/qe1BTWQ8vAdwo50PH4Dmmu+kPCKixpym7foP0WTZ0JJgEfaNlEvlLvUr81Y4XoA
GYU0xx01UqKw0IFoz9kxLS50R1rAoqKZdsQSJJFFNWBflnz/msf11bFfBEIaoDEM
NmiopxThrsHpZLKnCEL/qFqIBu8SPUtGB4GTE/cZBimEHLGrNRocEq1g7C3Z4kdG
LefR+PS85CMxUyHOY/DtAp84mC2ov+UdeMczqBaJm60Pq9q3ownw8pyjiY+hI+de
EGaS2iKY4XFenSJf3R1byHpnUHUx5GA4iKhK1IZbN8ahULwJUVjtQq1z2/HHxIzB
w277UCi7xczwJJfvIZaIit35Jetr/msMRsPcTDJwqKmSfIVB7zLq6wB1/Lkviny1
VLGxaHqAX8ibBfJBMQFFwLacubnltfB6yiwb5CWT6rs7iRoUdZcAHW7hIjmvVEX5
2qAuKXQ4F4mhRYr7CdNc9oz6firu0IappzVE0mFagEWc9/rN8c+Sps0vCpA9BBf0
iZTVVQxP/48SaGwqlTFbv65IBqayV3/iqvU29vAgT+Afd193+J8Bl2xVJcK5uZrY
JX8mYABf+kg7O82cbhLfggnYkBPKHjmYwPh2MD60O0F3v7gdx38f0FHmWZoG06ix
Y46Sog9ZCL/wcT/d6RoTCv1CQj4HuDcb/8BARtMTtD+byQmhSVoFpA+/fH05bG1X
7de+3wVtuM0Qm8XKcf4U+laW9dQwzSBQnvOobi2s+yZ+5HFeUZQb9jIQYGgqPn4y
xuOui0rdweOZgJP9a9mDOBkVkYm2PHHZJozWQZ/JO2NB0J70mORzTrrqG3hho369
+xnrxIfteekFFxe9toWFdcXgTIAx13/mNvoj5HxF+sVnNeYlGZDEKU6qmxX7eEkt
SKhyX2wYrGugbZHFTmFxsnZPyKOsZCj4j2mszcZuPsVEdyX0SA4afO4B6sjsw4JX
uJvYNyGsGIQl8Gkj48G+ZlGAReceg/6afrupmn25hQVxXsBI4GqVw1bjNtfx3Pe6
W1pd07AEJhJf94z0jaWFTyuHyN4pXFxMm7Asq8kbjIwJJyZrMkh88A+M7qSCffA9
iQSJwCs+HaKrdH7GrTRHoS6/O1BkNOq2oIFK3XmmQVkP3fCS5ZiJVg5YcdxCDxJj
H0ZDnWRKnbSyR/GiblOMlnz4CeNOT/ZEOBw4EIPpvTRAfeke3xIABSptXkQI894u
v4tHjgDetkbaE75lDkppTMWGgy7O60WT1aw+hxpqPRGaDO44rCqxLX8CSlE7NJ6r
xaw5NEW4CZYQ5UwwGdwvVDuLiiq+p+eMlTr3dXc+LnAI4AVTVTeQkNNUozUpJesx
hmzUTzGQNY+0b7VDSui5FkmgqoG5ORIHKi3t3hI3UmYszdGCTgxhaUpox+NqDwN6
bQ7dwNNg7B0BKou0H6x1lZ35+mozWV+m48TtwMk0M+vaxvi+n62sQWARTuaYAJWj
YCDWqnsRx2Vra8tRpU/M1OSob29KyVYyzBiPGLyvSvztsWYVMyFGaOsV5gvgdCge
og1XpSw0JTp1saIX+ctK0dNtk8k9ahFBIINMzcy+UdODuNURyFeJATA5oFTupHLC
myYaT3JvEWOwAhf6LeVhTr+sPUj6ZJzueWLFZ3xCRePHtU8Rj2hSfyB9t7lLoId3
xRDpIxbh42iBqGqtLPMMy5h+ZmqQocX1nSFdI8qrZ0d3EZ6xIs7GkN+uw1vk6AaX
JkLAOcXbGpNCS5eDjqy+SBkau129Ylp9RFqO6qAaZK6Yna1+eGP0OrWd4IOQtPam
ADIqoay6ThirazB6sqamsBeFlbdGmrXkCpXs1ACTO/2Go8vtQH/2sZaZSMQIbxG0
H5DZgpuxGB8MF3TQhWxKw6LCo5RKjYhuFCiLdAGaiD7anDjp1OGnC8uiWL9L+SF/
01kBV3qElltF1G0T6+mLIFtMzg4qh+FP+NkHPL13M0pTIoDj03NlE93wLgjGgP4p
9BeJ3+1xW5bWCz8pqoeJfM1SKqOC8mbyh7HYXtGLrZ4dDCX/6fE28GrDz8iB8iYp
ypfv562ta6H4SFWUqYR+54w3OgblJ8FwRBfiZHYxQHjpGzGHKqwtfCaBkxKBg5Rc
uCd+tnCGl/aPL52XQPoN9GqOHYnf/rRh3Ofksj2MinJtjZ01cuTa5sz8PRj7moqI
kZv/oPdlXdEPRPsusTyZ6x89tjgxrO70xSOyGRoSSDDeK/bGExqcc4AhaoeCuaYL
88ZgvQRZg0iWHSGZouyE2A7qsXnX4oOhpT8jXNHSTgsh0TGZA9TO22xezU4ysX9b
8VHW7fkwshCrKJ0150tm835UD3elWP4L6YRvKdimlQeh6dUUWUj3KlA49qCSiVVZ
DUcM/C4lU3DcauAhbnH5T1a7A9ygKe89z9QfbG0iT7K23mBST40IkWfwPtEKa4o7
UsVNroI0/8pxgeQ7g9KnV7rdYOmNGwoPf8gy9giLYmbD2OQy4HbiUjn4gyucSM4w
qacBEUmjeHacfOhiIyl6w5Yz9bieU4XQtlRhxYTDvf5RC5IXmszVjm6xUCbUoQZF
AY+zLlbaarLMYBAFqd3yPMGkfJ0hFe10nUcYn6hlavCAbbsc6IR1SWP+0tFQRx1B
YZkp/JgpcSBh2FmNiiHgHiQBd1Qk6l6fUGyB7KyuYjUEiXlFJdWtL1Oth5FsZyoZ
TQOUr7TQf7PZgFfTiug0Dm1RxHdMhqI6iGGs+15lUuBRewZK/ntD2DTewH9HyWDt
IYjBvbvl8Ya4jHnZ+JLrULH1e8EzmCOKPpec7PcdHnH2e+KIdpTnbr8gBl3qcQVo
hAaAl2w+rTdhpMFcA+SmLN8g2UzWgjveC8RBGdn9jCq1j+brAMBntgl3fOUP879h
i0m2sq9PMZqnvd+7Iyo0GkW+wjwsEBHaq0s05qgIeDSDW0ruG4+ah5kgtYtaIPWK
8gODCwuYB/Wf8eYFe/G/V45bHJkY82b7HF0YHYP5FkGqkSaxUHgziak+No/eGC8D
uIR08lH3thjgKBQtfcdKd9XoD25a6Iv3LFw5HsZAwqqa2hhXXP0b5/6eDHVpGhoB
Ab90TR9ElSiUElXXstv7PN8/qIJ5c7spkEOu6TvTHq6ur4wPkVCi2EBEQ1CEzBD4
HpHLRwo3ep7UcVWN4w4a4CwnWlFvi/SE4uoHYHsZNlZrUwNMWSZac5mp0KaN84/l
oRSrr5RkfKutTyA7pWbvZY3VXVcgchmO4kRQgHYgT69ZyjeyC+Dm/jMC8ZnwfSuT
vnC0h/kn4QLVLGYuMDsJNa9wTb1bPOHAzTZluN9IkyV8JV3H/hpXCi4IukoiJcTS
4J3harfSS7MNKDY/61Ai84PWKgCwaG3dqbYtAvND22vX5bCwDQRf+yi7gpLhwAyi
WoHXFtubgEanopDd0kbrz+IXrSkp2Qw6GjbjZV8EurD5rIbfEWaNJaShuPIQv5qg
N4dW6FYmYj0h/AMUyUjBIo6Osnqckg5+zogZOO3vgJb3lFugu4fZWuiTKnXvg+Jc
GdDOZ2Du1h7YXQHrg7ZX/MQvgpXTaI1pKJFgySp5s7GlrEZWhoI54UwierZdFOiA
tLfGs8S6MZv5Z7joy3hsFxL5fczi3031JtdzlrStGMPpIsf9BhHr5YA+ZavKFMG0
YON5AOcRVFlfZthFRWDVxPKVjHOgvM7UDgg5gRjIIjZdM24Wt7HPbeSc+R+Ypnaa
Otg2YXvw3wUPiFeJp3liM61hY67I5Bc6QvUKl48LFG/azuAGEKRd/a++IY9/z/ho
Oed+7C0igxGpU+rYR0ZnY5ZMf52RsV//uPv2qqFfQs7mBSEkKQOFZjOj62WJexmZ
YRQbwCGS72DsIxt9iAYDUor2ql2hBWQWDfUllR05rev8+VyryeTkHpGYqZ26azci
3bX77YigXR3DKdP8LcJs5eH9gOIJ8xaboDRUbutrGsf0BVIUe8ihetWGJrj/FyZe
dufx38/CgSzmK57J1BiiWg8dAmrllfqBqlnDIXWBpOOqblLUpCVEJhNdLOIhbA/N
Z8A27uMdHXWYtqXPQ8N5J3Wg2TM7fjztHyPdXdMYbIsmtuJbJzfq2Evw6a7uw0xl
I4lkht6xi2VRKo618EB5HATX6yFxNeUWhBJuO/voHz7XpgEt6DgI2aQJ6He8p22n
bJcUCWB7z5/p/lEskBBjWwKzNV5yG6leaWKsa5r7JvkNapb1cO8g8y3QPrF0RdhF
UNJj2MUa7Q+PKEBuRMU+Km/R33Uli0K45uftLDpmkIev5t9rR5V3n0ajAVzmL4mR
xHyvmJXXYvcARSwlkPIu7WWBsIblmpakKoxQ/tx+weV7uegUIkcP+8vQWJ9z06I7
CYvApzBaP8FMRTb+OV+zmnJCiyO2eV4tu0+Bvq+xydcUCHOy0y+7O5dJ2JQicZI1
tEXkAJUN2C1bVJNrizrgOF6VmweW8esP48mCIgoxmljhiZaRByujCrTajUEHDQbp
MpcsXnMogRPwPfafAQElZH+8kjsap3WfyWt306OBvKZVUK3MwIyl5Kbl9F4/W7iA
kPDEacZFtm/QH7bLu4uTPIt80kM4z71yL9RmnTzJ70xtWXRYYBaPT77JSalDiEtk
UPO/yJ207c3L3yIvFfJ5M9hAn04SbLPqZCVHMJNi5lm3FcR3OesE/qTY23j/mbzq
VZbfhD7mK4G/KYn9J2SX0kgVS0FAdCInAIJm+Q4Au1bmasKVD1BjqX8vnQrndwrd
GayxkKTBTK+nTY/Lm21HAW86IUyNaffUdf+njuocHtKeJ9A2XSLHqltNBFht84aR
wvhY8BCn8Wb1R+fW2kv2W+742QcXOOKiPhxYmbAhXIr4sApUydeYmKxUEdHlkJ16
JfpGL3xanELHCwMtzwJhhZI5Yd30HjcqOtcRIxGZW9Hte/8AlMc9VCCnbj63GoxP
y9o4vWBsuFRUJnOwgoKTIINLwfr6itWevm+h9/FZg6FUrufkjglFU7S8+uCqkH44
+Kul1GA6ez456E5NJBkHysEI2O60sWSXi85weOF5wtyWRpjlvIcbdlhKexNlwfD6
byOYjKzNuQMJXEMpkt2vd08CDXxUFW99FXN1ZILWMc4vi1vH3a9Isq1TBTS+5FJn
vqkTkA7QF1N3KxHpAzwjOu7CjUoQxG67bn+H+/vnavw4LHm8Gdr8z/ipSbgK63C8
d9e/uTdtS72sUNDiiUp7BqWThh78W/BqZ6rtP//b3CxNW+RoSVeMPDINTmSoC2rW
XML6UyUPVIW2/yZ7G/8l7gls4tWasl1IirILr+6rMEVRucvRR1wC7mgW6mIV2N+G
1qVT62txEKjcq5XP0r5x167dMSaG0FNomw0m0YQVDJnAgITUM9AxNZu8lvccKhJa
L+zdyeo1x16jQ8enwDngB3tsaY8D/7Uxlj3LLpkJtdc/nd9auFuRAfe0g1heR6UE
lpCm+U98+CPhQfe3IwpgjcNtMZXv7WVAF0GjwOFSqVA0SYCY7lFppYNbZ+RFQLZo
bRni7RCYheRP9x1yrS6sKvcZoqGQpyqqL42DKq6rK7qMwgkqPNWmZVEiWEtej2iW
iY3w1a9jPncIu2o107pkgHu4SOpf1rYEz3p8Jf14yMQNApT23DrKmpwFnUWEfwtM
hVFd64MP31qPoDp+bsL98goL2TFAL7fWxU0yuzzYieq8uQjQ3eePtwgnMOos1Ghi
G17qs42IULdkTte2sVFZ6jPIyu4YuC2v4BNox1ZJ3apR40LMtGTpsNAKzyE2Ux5y
22lcrZFznNpCAz9qDweFL7+iZSuSIB10Q6HKaGIMMLsXA+w1jXJtIM4x+Apxe/RQ
DPKfYOoHEWOpMyiietJUxpewXu1kjd1y7NBbLZEWWG7LHtOzutHDFsvCHC9z1NvD
OYfEfJmMs3ZvXZqbETDefe3qKSqEqg45VoYsa/Cg+2ZANsF6p3N8Bw5PAXgH2D+1
Sx0wmvZEuL4LvUKeaVRTGh/Wq60pJbrss7KDBU+QSqzoUlX8g6ahNZLwLV0SIdE8
OqSEOTOz6uEawxWsmPfp9OwYhyA2FRn0VjmLrCZkYXjZjANcbmwXWyUU/sjDiZZd
KWSPci51AjLacQiZDLWg5Rz9AHVuEI56GolfACizLhgbw438ZLgywCqrPggbu6XC
fe4z688L5+GIaMc1TPkRjT62W4uQA9xByjC0kYlX0GRcy1aSzaUWEilM5Dw2f3V7
dY3eLx+G8+CoyY5S8o6raIKdV/U28lto/o4Vsei03FcSf6QFVx99zW8IqsiI/rc3
BWv3hhiynNlU8PC3TGY4XSCz0jxbGDM8TC43lqa2Mknb8FL+OfD3lqGVNodkDcF/
jG3uiheiDhHjHDJXufHrL+I43Sc4JH3n0MuGpUBaxjSC272y9HyGTzJY9NBgz0ER
VieHDdAZq6oOK79RS1i45UQAHUsW+lYlXArh608AWP3JHCsewRmhhwz/hTDrdDG6
Q1qsNtfhKRgLzw57+vBgGDL5lURwLLrN3Revyb/5PGaeb+amODBEQS5cxLClsY4t
o3HiG9nh4mxQvikUClsJxk9JkowxdJMpO2cIMqvfqpK+uYm9jAgbiKg3JW5ddYOP
OlvDLMfO4fKaBR9yElv02H12S4VKCmzNv/tyHZL5W5c4TmsX/lnZ8jqjXbebAGVd
amrGBqHsq/2yWaPRdG9M9q3Rk9hk271lHPEaZhaGtBiKmodlPXwpMt1a9Op5/DMS
NmVbv0UQJy9b5JYAWqmd3YLjp7Bwk3kEhc9aTAewBOEXza5H2Z61jCC4LQJei0lk
N+gx7/q5k4r47jU2Co5OOPLyFwGFgxhvrVVSNq/zWJeCWulBmq0KooXzOI+ztUmq
cKfEXnciW3060ntCgwbTi5VGbnQTPuG0oRoC5nWyWrjuFyb/Xrv7W0A5JjLPBEKV
rv1u642GQVY7JpzHIrjr0cQTT4r2lofhozMMqrj9PgVOHqXtjRUvBzZmUvr0a6hi
62hg6VIkKPpBxJyJc8kaZCmbd/f9yhgMMyOUjZPKsrATGWXCjGE8X5dAXUisIDkn
m+jCUicVGCySVvOw8BB6j55Yy21Zc3JsMSzBSE4P3DW8XfKfdA8DnYQztISTSWJi
XxsTWo2GLB25/sFE2ZFt/S0Xj2/HpTA5OxhcGB8UTq1iQd6GSDPasfzEPCLM38q7
9HW1aYWJKXJWGBcl3xItc5ie7ibA23BF32SVpi/Jjf/Jb+HO37WJxqfy+g9d/C/p
i64z5e4kmfM1fBAXRx8knT6DymTzCVElqZDlkQE/+gBFRv+TacUmWQHhUNUb6MBC
Fcz5zxXxnK0rsGOGKJAH1TUiSUumkUZxtdZE/9lN7/IH5gUSG5LifEq0d9Yzy2PE
jmSZxvBDlmfuTehecgUhsP3NnMtaoyhaMIYqSZvyCv1nAaKHPujDjBzGk7zLp3i2
2jYQeQdQCOo1kbZl35uP7NR7VsGJSDvJ8lzWuAUUSTlor3AkfW9eeAybdbZuIO9k
lFWjUOpwn/Uw9ZS338m2jcTNeAIRBU9v0TUdBz3BmrN7jiCaxZUs3c3AaFG0jrsU
XuUKvJDgYQ/hi2VvfZSE6aVZDEVO9Mcm2CmBnUBzLoAPDKI1QV4HEB6QJAuF1ovl
qcDmfcbP8T2YBYlV2qw1W319bvB2DgbEYLbeupX2tbjTFgOh2eqhMRmPyJgYUrS3
56Pj0KDSoMaJi8eW9HnbJD8FCqMVQQXuyQCILCMh3k4a06toKcndJJoESbeAkkVj
kP1sJAiA4mZgy03S9zt6VNAMha/89SZ/FkEnfjVx7icLE9F679nSOAq2MB4Zy+8m
pL0jc27y+Z6jcriALJzZV1jAlpjUz1vdna43drgZ6wMOpsox3VVpxtVhAPwADGO0
kGk71E6mjyzi68SNdhbumSwQTuodKYz8Jxm/gKFRlTuTv9R+d2OlchvvwgLeDiex
yEBY17AJy0HzVBemhyk9k8toV8PrpT4eS7P4Tv108GfoXG6MdnMn4YvZjGz+pT8T
UXqYYbcXi1qHrl2K7OGRHo1i9EFHxe3ApmZCnQfwGV7J+yCk93OArVrSOP+F655Z
uXq9riwNmhJ3ouHkKP9kdNTRFkKBOcvhmK5Bm7XzZSjmG0bKvSYsAcKYb+cg4dHA
YLSueX/fq5uL/YLCuGFjSMLKZtMxtl28EZ22adSif+8neOpTwGsfXBK6exAyI8vv
9mpt9zjhCauF8h55zeSF5ik80fsCXzXp4Ky/sXyalEf/quV2c9nCrlXm6CXtE6BE
00X/ygEE03ezDDOuca46br69FQP/0pBt7nfMrqogNmlFfBPdjRSJ55JQTDqAFnFL
wyUPwM2z0dZjnlUfxikyIM4cA75pVLmTAgpL5hxQ5eI9JjACzTorcJCPjh7wFo1p
+oDPur31tubRsybyBaXUkdNmIy+cklkiQVAH1ptebFp8YR5HBCf/1nc+asN4l6O+
1gmBDK25/NgpphJCtaBjoxh+4oZTRzrKuapIfCZ5zN5RrOl7zmx4+PfbOr/2wGLY
EAO+Gxr9rzY52bbql8on3IdAXOHiZy3ciB60M2DNOUyr1uOIp/mWEFEus/Izk+qV
8bQYWwuw+Es/+0kuqEIV3HxmVw6FdRSB8kXa+gaFnserbN9hRKSXSQG4ixMC2dnW
8Jp5e+7U/4kS3U5heTlmErsg45Xw6kIPgS77wdXbV8ji0U6d4gXeZFkHKrDsj4tB
80OiLY+xFJNQAxqoJjEaKLiRrt+kXyWRMTEQIjiyPiLZbksGzL3mKTxziLE0+XCT
Z9Ian1m1NfX3SYecfKZNcTdr/MmV8JoyE9lWp6OLdcD58BaZO28hIhevrQsMEn6g
VqmfeJQBVaKY6jPqs+p86iUMGhHWpcrBpu+X64V/2d4oYu5sZQMGkDGummRy6i2z
88ox/1JOc2P2gtroE7a7dNS+tETI/w51ZvVqz/R3FlssLC/pBUha8Uw4FyRytx66
KIUHpapsM2nSv+tmzQZXtTz/sfbmcB7HNQaDzIgfnUiLghUFlitztPVjAsYOujLe
/84zGtlw0BU2OjbsynLo49Hz0lZQUtGa+H8xtnhGnH1Uj4UeDXkSo/nywGs0vY7B
DbWOhZWp+g50ce9HdWGqHcAlpy0/2Kor7d7yhtG2mN3ETy8bJKM4JrIeIFJ6bhAW
EawzdwDta6Hf40QdvG+EVx3IBt9df7oCXbedMZAsh2LZMu2UIJDoFhJ/1ZEj/w9B
aNRJe5EPNrSPUU6xFanrMXLio51KY5zLZgyzTqugR2oQ0z/h72P/WL2ijjqiS/Hd
qdeoJIwMulfbbcEd1SxStzz6i5csPyAreGwmPrSq/BxBaRxA2TP8X+6QFj+6vt/g
CTIQPxqPpPaJsLWqne3nWN8lGjG6OBka+aRLzXtiN4QAQTRnqSxLTu1A7d7qI0Bk
uYYRjGioRlXecml1G7TA8CcwEi40OOHmj9ETiWF90wNGl5nQrPZT7sFzxdGxgqr8
THV/M01GPM+p4vpOBZDsIMoIl2dfqWD23LewMro4q+6uFS7QSA6HNZp9QbvVLfR+
GqfAwcY7mHGbH48WswG++3mGbpjPM1LnhvxocDKzOCD9x5PeahpwM+oBsKDtWq8s
45xCspqzCWhTmDv5YRcm+KxMi2qDt0J4jYmv2bLiuILoHWRSYXtdYOhGW2rqCjgc
+7Y+sXEB+lKAWCunxeQydlj4fLNrqWPx4L3w3xIMGbx0rM3wxLesrmc+T8l+aYQE
xx0VY4O9pODT7dRr872beLmQy2mALEixAbcIkJrmrN1xTWICJIm/K+zrv8vAC0HU
BRta7ONjej4sdIvahBjKoSQTYpmItUEZ2u8AtgcUcGlvjxQ9aUCwY3KO+LA2PK13
TpM5x65BHg08EF2Y4cV5JxPpdIRfRYmccSwqpyf8k/6AfdEI03HLOgFYs7iYYGZW
gjirONnSm7IRt3+5chiErZoWAlthviYJJnJfwsexHztGiP3S2egZEDJ7DF7SCHNB
VMMdWwXSTZ9KX8mZOPZT1cDm76/f3+vPIUFjH/d0mbQ/vXkOa076aXgPAYozS2t6
3+2isNETx37gIrVAaVzW+CDfNpUV5xt1gHuaqN3muQdiierREL9SSnhTEsoueiak
wELyvLRooavJgmgMxMTzFM81om5ld+1v1pRSU6nKWYBVjmuDmvcRla5oNlKcKawJ
AaWslRS/bF5DZ0P/UB0TA5zLkQLlihCI0RSaa4Jd18OcIAnCu5BKyET7AsWbK9jJ
YFTl6lWqnbPL9lFa8mxQRMq0fuShDrsE9knTTCzaTeWIRt93SC+M0Ij2Rn65t4xO
1OYmj8Qj7Q6AOnJMFsTk9GjT3g1HAWkT5NCefeFkJXPdMJA41JL39nKeTV9KubK8
kVhkjon9EWYJRJnow3qf9MG4HBqcXBbXwsXe8aly0hEl98i4wZn/Qs4bDvSVo8O2
DEOOhe5KeveJdvYogtS8AqM7n2cdl4LpAhOsP62K6ObAe85FCBUm7m3UNHWW7gu7
NqTbavj8Qq04uHmKeZF54/uzifsMX8PUJoJweEl+MQrE5fbvCbcHBzsHQz1Bc/+7
3sWTb3ZQW7U4UK4CutJVhgxPCf+Rvnpyjpu54vSz8/F9il+z9WyVAO2CsdPQf5Sc
o7ykXAanYYAwpM898XTOcfFy6gsWPfBvPpJOWCC4goPnLlgnVDdYy3fsh4V08jNE
zzlM8NqBvsjZWjFV3tURq5b78BrSOT3EO7krJoH/WMzGClGkAOurmfQ2yC9ydeuT
f9f119/wq8zvkVxwJDQ1woq38en3zuUDhWuO1i4a7ZUmCzmxfwi7A3q+wTbEW/ZM
D5Il5r2CrDgZXv19JToZ/XATacqwF453mLVkUF4BHO67cez1+qYcjukddoxGmB2e
4VOEzXSBJ0k9mgjAjoSAhR0l+syYuWiEPnYZ5KgxjXFWkt9Hp6jogKcNgZr/mpMy
Qb6R+b1bRvILJpwltF7/nBhKjSa5W+XfJjpQCQVm9LF8DUCsxnp0GtMahgDNff2o
+ixou3JuKvzZ10t2ViUr0yLY3YyLXV1EdmAunroHgYXy1DweZMjXGGoVpDFoQgXn
CESYH34bn1TdYAoyk+wDJrHQ5UB8FHRFbxznkF8mng9H1YyBppTzOGUok9mNr18g
7KD8zKJhOimYiAy8j95R8kwcPQVa3MCVgUzDy//cvecR/YRF+RnGWqyDGtiggC92
RIYCmxwfONj06KuDxYLYJCBxSJofNAadpo4Skr077Vlib0WDNQKmK4sZJYxNO4RW
iVwV1HQzCzFa/uafxWwA2OTH9521vEr9R+xRmuUMFHlubm5YCP5wV+bWCngp+6XT
tzT7QYuDJ3UPGvyYO8Q74ds7wp8498Fnr2rbWi/W4PvdPUDT2Qn3hojuXx6f2iVS
EUtptDX5A1+06a5WG18yi/ZxgkjJEMM+MfxW0En01N5EGEujxZkW3V7EbKXf3JxX
zX98NrHm6xRYXrtSOgCgdvEON2buqxUn6korSDJp0rUuXU9RF3bno1CTxGpoy5GA
lJxL+OoCpADMgHLl6Zgo2WKotsVEFrwif4NRsCaDeQ7ExDOSeOW7N+3TCl+zf2PN
Eb70ADKAyN4CwclI493DPr/Icd6DmLgM0I+Iz4hp9MK/TJz+oL/2uNMepph9EM7c
wazbaNkYlF/u6cSZ1CX0uQwUT6XgZ8d3DSgaFBrTLrvQdxwE1sufvYqBcbNTsrPV
PxHgRQp4yrw5oDaNOzrNz4FTeluflU7iKIEg91yCwz0C21rBd2TsHtj7T2EKk/9t
+oozkc2mfx43Z3NIac5/wqp6CyQBscrevODSSUMF7JHXTGzgcSCyFJd5xYD3hBn6
h3gWx6NQT5dzRoP8b4oz9bQcTDFdPk7rlT4zrTi5EMcIMyT3Y9gJoxTvvPoUVr/D
cP6zdtlmlwX4WMlDckXwOgi4tdPOhE8soQtUOEkAfyWe08wLBdotHjqZMgZapJ/d
x87dK7Q+NpmFf15RhHff496B8+gOBlLsr9K99OdYGGPh9oTS4wItyKoruYsqBmUh
jHkJklKA5j/AxjA4jI0fJQjW7COJScmWAcYd7WGfD81aaRdtcxP1wS76Pg6F8gLc
r9N1k5RCcjSR6dH18xSDsYbSuz6iO1WTLrsWDE90jT8dgFYe17LEqyLQRvtlBsvh
7T+YF8meXLwqiTf1npSEkh+bE0n+bnXKzGoGcVfIcMd0i5twVmkK00zLfbk9yhvI
5Yfow795GaLGNliV1En0Xt8gI2CywPsbDhF4J8d170GlzwEqtkU3SDrH9m4JYr+o
8fUgBKdb37CH45sWXFkqwy3hC39etmDZ5fXzyQQzbO6xQpU4eSrxFMLyxqrhH6Yd
ob6DJ1a/oRLeg/XzWnnVw25xt/AgHhj6o5Xec2XaI6fa+VEMiy3OKz8BBZ+CkRab
pCqRHwwzbUysEV1LFcVYa9brzWLfbPH/ZT++U6bxPJIlgURIeH3jSM7aoMwWV00X
aub4BKDcVsizPHlZqhWM4UwHxn2vJttFoc/RwrZviysotgCwObZkIdi6ISpyPuZh
1M2i0g6GiWq3z+Mrxs7lZH2YM3sEnpBogYrGy4vnK5G7hgE++bgU7PpgVQrZlQuu
qayqs6BPu0jlaPo5/ncZcSIM6iz8zygQ7iYWmdg9fKYZCrP3s0/9EdLkYTxm6hQi
oTFBHfkMvTDwfzq5YAKqfYQzPif6TTTEEggx53ICSVtAXTteShJuKKO+r0gM3hB3
vWeljGHdShXiWKEtshBV0D6QmUIQBzxINH09RBuJaRfwrG+EW8Cc0dfr0oJveFN4
Ot2lxnomd5uG9q0zn3Fx4oJIUZc/+RTNiby6pKPuLSychOJFPcidbNquztVKtLW/
0F7iLncIAXUyL70bqFjKIdSzUSWB+R7+t2usQq1uky7LdokGAkekEXRmq+qARNKv
0nV0XQxliiZf0zIiKkqie2A4SjbfMG5DGEBMKsWT1mo3efdpIAhK2BAmhpaA+xau
YNc894UZAOezwUBYaeKPqQPZHpu6Wk/0sjKhwloqTifTX9vTXywLpTx5VejaU+BT
+9jRBxBFdZVItBbLdMUy6UTxZmWJI8oTjISFxvmxn+2VIa9mFm8Lc5+NesL/2Vd0
7h5CQmSvuhX3KN6AuXNHRlYHdbRTt5ETa0pdlerTB8Vy60uGO1JIU2H6ztZ1WzSc
Y+8H4wwSBuVXV4UXjycI8EQXbsOx3Bo2GSipO2yhL8aAsZOrPe4bBmlfHcIkEhVZ
IA3nyM46n7fAc6Nn9OWUw+rl2CDx0tGeZIqNqZnsmQkXhbKWq+4wNPMSs+PdMo2e
NEF/dluIfrmGyDeg/TihYSLcfzZMlsD3utt8dNgFvbAPMcvVai2IkTQVRx5hxv1W
JykECglP1srbh16AmmyDyA6oCzbs5HMvT5MvXFHo2PQXc5N1iDtID/xR6AHJzilB
/YR2IvNiaei8348gHjP97t4qOeL1cUs6BdK/lqfkI4vzjQXm+UV2rg+H+yzyxOv1
PQ+i5+Zocs+wEDcuyeRhoSjiYmI0Khzuf5btOr6t6X8M+0qvFKedvBPD96LITPZG
eq6BYMSdDmBN7dhpCKh5Kp5Q1BAJEKaQ5N4Z6hJPt44+Q7gfTZRwELiDRJTTlaGu
koc3N/W52fESg5onAgTM7EvowGenZNC35FOXbDefdClrhbTuimyuAdudPvd74H/E
wWAaScN5mQJII+K/JZWgUi8KWMUxNGD5RIS1HS8+/3g7wkbpAZHB2I1vS2+e3TpM
nGm860PT5qbTBVpGpSMLEYhAIuI6GA+0CXQgmNfwGk3FX+5LWRvfOI5dBP4cpPmI
ximDHWjUCusSby6YItoqHNo29S1CqRXo6vdZd7CmxrzZO756pILlSleZstxNq6JE
vfY84WuaWMP9K6Nj8/PW8h6vxFT53klLfL3h8EKaCenajUkrZ+iA4OC4jaJgdTXL
D50+2CQMit1Iy3Fik/TL/y04GQGu+H58ZKfgxTwYuw9VEVj0XQ3OxNIU4+N7Cwnb
0OjvQtNY/hp/JdZsy2vhm8CvBl0RsQizbwitQIN5/yXoQ8hR/4w4of5wcl4btdxZ
1Q48yAI2iAMIGC8IEkGk4wDOSb2QizfYf/irDge03rimJeVn9NLz1lmWCVFmScL5
ewourpAD/EMImulXuCqzHFmRXTbh/Cla4OLhaCLppw17EZ61zN/7zSh0bEXNAEcH
ug8PwHPUjkT++2/AEmeTUulD/iAMiEYZHNU8GwULBGpPFPUqwyUXn6XQslPd9H2o
cZoOI5wuFx7ZK5vT7o5zjaJotpITEuU9GCWIvsNKSAo1F10X6U2OkJnXDRLDzIEU
QZ/YtMk42H6s9REzpFTnxHw8YigxsfXijgsd0QRSLwiNGVEaxLsxbIYXhvBN0wl6
UeXIU5XigACeGMgmepPTswOtZz234WDEUlQoDEwq19Ch39Lfz9pAAwfjV7fD1GNi
Z0IIMWJaLLLCJXeQjtIi2rj4vW3r4FxJYGg03uLccY1fFs+pyeziGEnebOIhPYq4
tmpqOqLwKRJgcUgQwAKisyxEOvy9ZMe1j/gtM8wE9ZbjodzrqVH8bp+c6s1AXghO
BUqO0m47z8VRSmKwqJGsZ7c/LeILItM33zcXyOLyLX6zQFTZTFEXJdOrdGc7KeHD
ArBp5DM/VDyiVnrXe11gCDAEESeDD9zWUkiDaodugPZjj+NrpJjQ5HFqfK1BgmsC
sp4P5n/I7I+tH33M9DXDB9sGMbk8qO+PjcywR6xoWZLRQPJ+AGkUgSZqCkU8zHM1
tI28e/bP3Xxv9GO+nHbNILnaLSkFdgwy79CL0klwoaKReR24U8gaLeRBKDe+zjhV
jZWHMf4/WrxVgqG+rHd/X/oFJ+lH4oeCAZV4PaNv+R4DJ4+rDLyxEnhGwJXmhBKF
dtW6E/ewvW3fxLWM2U7OPhYApiCgyIRKjZ97XirG8+zKyS6pKJMIUGHuDT87Sj7D
QeIg/oVf9d3hj++wFDRaQv+PROjvEZLo1e8U9JElYsOnE5ogzeo81KYI6DpevZJO
8WWWGeKGBe5wfKj4o53RuejI7g4N+AlaW7Pw50LN6FyxxU0QI5B51NwKQk0zHSdG
KifpdWTiH7f2DRsd+91Y3O/w0XE25B30l2X3r7W7Vv9+SbeyfpnzL5OkUI8IaR/u
GbXRr8oC2pSGrEk6ItkytMCftE1BnJ+ex192L9MSxSyrnXkf+hFLwS++nKRMZExJ
+bkrNma9jLgCIjEeRrqZwSZZB4WEzUEj8EKKzT9MSO+r+VsmvAFlfXyrhyj17a5l
3xrNCbm/Yw9QIWSdeEvUlzfJtGsuDCcVW1P5AYFlzPdBKiobiMK73cb3tYj68l75
+IEs9XzkwIH0hH1JsRrV4G60Pn0ZE+VLA/fPkxYalzkxq/HLLoCAbQDpAzsRPW/z
RpfvIHMD7aX+oMgrP+NK4cuYhx8YHHiWdnwfBWteGpJ8Vphc30MUdJYjze62EgJf
J5spn6PIFxgYK5HqqEQcSZSNSLtIzSjEd9WYFDD16mzesF/um70jJheXANVMKWcU
5i/oP40C+tVuL4lJZx5MtsjYESTLYlyVyfqNxmztsxUlEc7l9B/SGFqK/4dMrA+k
VJqhRV73Zi8NT1qVjoD8MG1uKDmbtC+kh+LO4GMKibWEE5Eh6716NrkjZT+FAHHp
peQce1Wwz/P8xYu2qGS2v9h40SKUhKSmYjj/NgkXYvHyzHz0/o1QZIZC70UIzLnQ
HeC1FRjj1Jpt+buSCF4cmC2oChRDlQiAOVBdTx3YmiQ1yLIBq66iKN7KnoDKKjj6
NXsL4rNScJmkIa4nEEZGfHj0GakGwCVyxQElCVd8Y7l7VShUlqRu4MJHKJDxHsCa
LGF7+n05tY7jA7ekP+GmCqGo2Q2CjrqGU4Dc35dnSow6kVTOZWWehUvnUBdPmFTW
n7rVifX70+Nxk4Jo3/sChuau5jGjRsZyakCZgWeg5BAT1vlbbkYDsoVLAIL5NUAP
rEdIovhAzzlYlS3G9XGRhGUEwOxZ2xlzdoZR33HXkBLftj5zkLXzuioNSa1h3NlK
ATa1Mlc3iDsJXNNKSNOzictc37wlw/1bItdPSlS8ykcmWPDavyZc/I6N4It34Gfx
XSOnMPIXjAqjw2fS2FHu9KGZjrd6WpLYymZ2SdpnzESYnFfQKuoZuwj/tlrvA04O
fUnioiiLpPffma/kjUp0XfkHe1eD6HoXimoxHcwhEGoGAloguPKdSKhwYo8ojeP3
pYzhhAERtAnS3Kp5Los9C2GAyIe2l8xI37oWFjxtwDuuPOFhJqgBSo78btoJGhg7
Q3eTW9fBnqVdOyCq8EzMfGNDLx4RMk5CxhXODbXrZ4RxtkbTX8Gc3wh4tO6/ez4k
DG8pvZnhNl5hlFOUi1QiIgeXGRizjW8RMLFY7pLsMe0yCNqTB0pFfW2rSt4Il+kO
Iys6+4CjfCJiU4NVHETqWpqu37rnnTQvNek2boMdDpE7rnxbvoQ9OS9xOgnfiLBz
Ple+bhk2syee0wgGJc2jMlKC6hOSoBbkyCUEZyHJekNoR5KwDMlv4boTv1T7C9Id
n/0Wg9G855vB3tX0yxTwDYVu4uLsJUmtmJzR7CcgPWIejbVO+zE45+8nN1ybmgMH
HhQjnPTEMx8h2f+1QmVQXxmcXusKNrMJkLVCiCfHTREZrBvB/t9cA7sOBZneETWI
/+E2+D/3l6c5ueDiecjTwMicYLlhgtyJnzpVZfqIwrjtpRfOXgKcu7jACpuh0muk
UT7hvJEd9sRAkUBzEhPtA+N7SDIcCWsLpdpxx41PYMB02zDcs8wgqzaJ9PjHRpU8
7BbUHqQtbMW+9ocjqlvmVTL3LGSvUPi/rqn7Vke7oQNh0jEZRG1CDHsr7DFz+2Xu
/jF0D2nVqnMV6bkjgP3rfGuJB2TTVEcNTlAO4wm3nYJFSxZiXC/guO5zrjSNJ4ba
Ah88o/PRWv+MXUJCfZ9Bi9VPagJvHhTmTFo5f29euYEKi1IYlqRgaolL3EjhBN6U
Zlz1OHOp1gruOJ38X35Vw3XMPVIlsiWEK3EiRVEu9QpIkkccv6xa6XOdvQBjq+i0
smxRC9/ukxfhE23DVFQK70WHpfeBcnSRofqVKb1uhQ0Jb9PT8ZLU7yiz8JosZeM2
iuOh++N64wEUBVyo34xdhJ61NCEHVI+Fv0Dfo1fJzd4PTNJYcEJoQc3+stUiEV3r
8/8POHXJb+e00tChUxcc8n+nZmi1+G6eT1ruOZ6VwvPtzsUk3dTnH6greGscriYX
QUYg03JHAHI6yMsTqtJzCMO7Z5SlsKrMxlwLzeTuJ3MFVDRlunYLfDTc0u8wbDfK
w5DGcFSGfDvtD3F8psFc7jZO9WacEVZ+vO35TttPOurEMt4QMnDEK4FcBlaZk+s9
p8B8s5a6z1GoRhU1YWqDWABZpgxd9zw2WeoCDBpDFhaX6cYsCOu5kt8wdFjalhzN
vDAFYMb6adCJZTujdyARSw99ptykyq0tEp1rksz8uME1coTV+telWM2UmMLlBvs6
FSY7qQdG+2A61ukNBCr2ZzsKMu+IcnmfSaejED9NN5LcZrYfY8ttSna4ermiTyFo
E4INdFegGjMqQFEzfDolLZu4QDr2XtvmxFJL08NQYVYfgA0AU7TqxPw/vYnE9T5t
+t5Sll9uTK6fP8ZksIeRnqbheK6PnoeqxFxberpjp00ktN/g3zG/0Tm0DY/fj/Z5
OYjBvDHsfmS51zRGsZbRjx1gIeqmG/TDBwJ2kaOWXLIIsc5jrYCZjpVO4GrOBPtO
18zYuWxSew67rZk+z3CYzoLyAgmJx/zUIz04mduD8h/8HSAW5X5AAUUeLtiQvctz
/lcOruG/lMee4M8CbV4fOPpwr2qHxTvLZLqymaRg8QAOeUtJcbF1zvXtIewjpkut
xGLsf8LaMNPFXtFlAisE5fO1KF3gVtUK7rPnLODqko22Boz69CeBS4XzlCyATagV
BNAchnr/JeSNfLQ5LpGfcD/1q/n2GKKpWpg8mqna8lJBjdSIkgzH84NqlNpnZRUI
y0RLwwkRZEnYhwuDk9DlujqdCJCJqZ+yVt+cAbNMpFvERjB6LYzzAtY0ZmfGR5xE
XH626ETQcfwHD/9oIyS/W76BQZoNZtwha4PsckV776IjgkZwX0z8PzAKX+dRV4i+
0XV7SUqOi0STXbTYBCCn9wyIvHbUtcNp08HIzn1kjBtNxsHREoYVFjvFuPDglatJ
Bq0gBpoYeLWtK2ENK3cqIhFQM3ui6SG1qSSXv46+CQHD52fJGKCosfwv+RgYj/5f
IBmm6TlEYMP2qrD1WYqGjyyv2lGRa1+ATeCShzvVYAjQDHMQabk6n6vz1Ml9MVhk
vIcda2PBtgjwGyJJKaODjFfMBf913lOzHtxmn2JsO7WbFFgNRzNgoiXLHSEJh+EN
PxixFvEsuP6i5EHBwABJR4gKtviConhR449PwZq7hGKY3ZJ3H56NqRv3Xm/zjF0W
+STyv0FSlwYdq2lZGE6tEkHoBK+8S4cP8TnA8VUZ/xKTXXBe3d6CEtooRim+3lkf
CB2ZaNOyw/c0aldpELkN+yC06Xf1q2HC+Hh70avbXclrAmSYupVGMre8Hws2cxPK
NWV0NWUMg7stH68l7fFpzvTYbXjsBsQ+zkwvJ9+sapodADa7ROD8t7saqn2kJb59
inSGagdgDq+ZwXBIYkvfPJa+LuG+kcGo9oLASA9Xx3wRjuCKNC2FtTrOMUi0EeRT
olYQwYTds6/+NAJ2Il8flBUs+zW5AHLggRE13sTLVhZhuexDZgkZFN+pef74LZ69
HX01LJXTitomGKyjEsROIg4gLR5INEzcJ0/b8BrnbS4bf8z5WmUdATL2XEfg8imu
7oGaHPASbEQWQYUgEpVe5Xx7Puo86uSy0W0MJfzWF7b9IFPciLiSRZTRwuHwP/RX
IOADbA7IXgY4/T875UY6glaQNUhUnlgwkFZPczkHXEieb9p7kfi+zGa7xOnMRLxD
NrJLXHZQy6Vn/jRYgTC4dhpT6cOVJxuxBam8yZh33dMhJVNIifQ1G3Y2GMu45/FE
+LKPjRDD3Aib76ysn2GXB7TFPopRfAjX8ZtFJOXcbovEAxpApt/AmgRY3+V+OPiG
C3xDEPXg1vng+evMM368n2m+NwduGLFwBEXxX9bJYKvROscOBaBr7lFahJIwTyTK
O3gCHZnpYxawSEYlRYzo/bttiQ/sPcqlan2ojiIOySyb+vr4GkP693PFyD80qF01
eshrtfZo+VZsR8iWHHYPFP5LSsHcDeWa9AlwL2x47TumPmOZXv+Mr3I9nUkGLrYD
KSNRrD/IMf9JtLLnNGn96FDRnjJiN6m/Lnv6RnI5v14Dma4CQ1Od6q3JtVS0LgKS
r73RiMnhkCOPCXVgAUqAPWhDtVOgqYS2Lrpb319Joi8k8/HZpcmU9Jhf9ID6xIV5
5Or/DdCwNzF0v3X1DogMPh0FcmBmrT4Mqb++DG/O4Xn/ibvfobw7Xw2Dbv8tzx1f
YwH6SHvb0TqzvwvjVcvVVdOpxwWAoyqPQ73l7WcNqkeChTjfmkLnOMuT3HtJO5Pm
o6iCjx4JtFCcVBih+dncKX/ElcbLq4Th7PYjd1O3BcXtC5kz2veytTPDVUCPHi9Z
waoCPIT1BpN60+uGxE4SRMWNFNVqMjAfTGg9pZ1/zX2k4x4qYdcsvYmomlB+mcGL
CeqNclJPMYCYBgXKF7I7pxu3Wiw+ZGjk4jOukKnb6tX4nNaQ465e9078t8gxFB1T
O+JnGvYJs7IogB1mvQEemvX6qMyhyBHGTDKjUsE/uZanFMJzOSsSdvSYc9YuUyJw
2Pji6CmrCCC0Kajs1a+7zL1veOfoM+T61+cm6+aJL4pgO3C6VtLSnYSDDmXj+buT
tct8nPKPE49cVuKVWm1vnlIfF2r49yX50GsnYsZEuveJbhmeGjLdWbT8pnYZdNTP
hKI74yZj/8Fc6cI5ehXYDhVNU0ccXj4q+OavDnkXxGVh65laDHFc/uPrCbmPLMyX
X9fK6IrI2a8//HrTKRWaTtcXokM2llM4XOarh/pf3Yg3hpaQvP983XysBccrBiQL
A+oBWcKS+Bsmg0t1HhYCUsfVHX/mVrWliWnOghptmu5/7hgFF1QQpnQvjiCTJnem
qUmuPPBVc1kjPEzHeqqOat7tJUWloV4gGWGB/NGPeRjt6FWI3W1b4L6393J0sNkE
CvW5dfG7NHD+oR6YFPhfenxooGEry3fm4heygWkvAYQuIB9NrZey4JPSHsyUPYga
VITzHkn8Ch7SXND77Yuue4z2lpV+SeI1HARiIFaY3G3oBAu0GEzu9smqX+kFtcb2
hedJiaMAH7wDbsGsKVt2ciqM7jjVlMLVNPXV1lNT8aTcJmOrJYwVGCJt5NfwaC2w
wejGsMTRO8e1qd8v94w+QKGtik4yWy9Sc8ic/8VvcIF16tAYggXuh2QsNS60LTC2
JL9ykOcKtj/WI1Jcnu5a1uKP7DXjS0eTA7Q/igngmJ2bfxA/N9SIPM3bfiY2Oynw
+64aIDfwn5wGDidI+7h2wRj2dVObk+WHIxhKZdoQSscFedfUlIDt0mQcVwESp38F
t9VJEi5CGwfME2Zyas33Iak3bJaV+FVnB0uDytKiTyYgcXMdm1zutLGwypf45hi9
JUhtHBS2t/phb5fEsrang4CHMPf0LpmsXcQseIFtl1eHepIHd3OH8o0VB3uLUSuk
P9bZq1W8KqIeNGbRqtbPPScQ0XbVdTW7/vUPdd8iYyS9TOeIs18uHcF65xX6ajiD
BDqIy6JsVG5GdZLFOGMEdYvgXzHZ6hr3AOvt4lCOsFz9Z0ASdMI50PeSEZyJIvcf
Dlrmnc9XsSwDDcij4/rWJabB94xSFQmzhL0DJt7+9B/1UPenk594NqK+7G95wuvU
qHWNDYkvFeZIcz1B7sKimx5eI3mSKw21cVvMK8YobETL1IA55e4FW8qTcBTeD71l
RRrKxn8YdscK/kcE5WiCR8//vzqdsro13ftx3QRmdkPUQewkSTToW4pRqZN+JqEj
pqiqr9JwAkBnZFHBJIgk1mfjH3f/Hf2eYNVRXxXWRQNFQBI0VK1O6RZndTHXyCeM
UPT4gEOA9aA3pbu0RBzRGa2m77qO0J74rZzBfJ+pG7notOdjnndOeySiKR1uFZIG
uSk/BQ3IFQgPchsq0KlyjnusfQr93knRVo5chpnWE9MZgoEGV/6brSTG9JYEuV58
8sXmurbQtVnBvXrhd/fR4Xh758fbzokM7PmRp4gELGKWWogWwbyt4eYteBCqyaXX
7AWw4GjQhKb1lpkYdP45gfvsffwHRhfjH8q/i57BfXBcXIfLj9kRYsxLqJPegNx6
Gw/jPvOvBx8G7CykWomP9qHeu+BucF0040hubgPByJ9XtTW0+fBHugeFogQGQIri
MlfQzJQLs4VSKftV7O5NeSr0gfzHPsHQ19yL/jxPA957Ng6D/LwTMhVc4ts/UUUL
j8Ht0q26bAInbyqTVAPX/wrYIrG9xmBtMm8DpzMRnaH6Q74nWoBH6VsEm9mvumK4
S2op7sTXTU5hy9lnUxam7Dy4s5V+H8oe+/NKNxYrsBlBmLiV99oazPOr5ymWbduP
+s8qPVxVIxsDiRhv9vJfmLwkLp4RyaNuHJmKe/v9NMqzkPacHdyIS6q5tmACM+5f
IvrkufIMRKjytnDdjNMcqBwP036jLQxoJ3RBJ8DcRDuCWkPxZYh8l+ZZGBjjNt4A
7eX9T5kuFuXT4DVPuBrbW4N+Andmgqu0nMKLdE+QLr8H93CjlXtPH7eoEBEeg2Jr
yPfymqp44MYwZew7UJVpkzp9nRddHhDrVuMOjPickCaU/+ypkU3IH0O7DEwnfuKg
Jjeq4LMhTRfrJhBX3AcvLg3caYBYqclDmdFMmET3HxTNdukguX/pOC6VU0yUZBmo
+uEAo5QZu7MbO34/iNG1pdFuthpcjHDZj7oKTwdUOUx8XvNhwUTkSi6DC/VYUnmi
K2y9NEtHHm8VPd/sAIBkYUz3Rdng5QHdlb38OXNQKV8xklzmGqycH8M/qo/bAfyf
RULOgsvvOEiyEsvWGzShgkmipvi606aRGCAnrdpyGVu2iLrqX4NRB6+Cysk7WPzr
L1qlfoPB+A+dzqgjdN27/1KypP++vzp9S6JWYdhgHGhGZmXI1p+9w5ylJ3d0cReY
T4IwxyI+B8gGBagR09A4JyEWzlqoYWq86azWX/E4GmYiY56z9GwssTyf2MvUfLtq
F77Ab90M2eccG91tIujpLtc0T85KJIo9Ishx2Vg83w99uAC1LP+ZXcMmnLayIkJv
1H87X+3D71QTkBk56ts4l7qx418Hm9aDEL664UZa+QDpdTSIKMIiXFCKzE+ZPKfy
Sebd3DpNKchA9BPz/zoaOv1b5wqPoGGWwWIWueI7tI7qVbHn4gG4gBQAR/6Hg1VZ
f7KYL1bEpnsTrz/zaBMPGcuy0KQXFzY81NUn405drGoLvA2kTr3p3E/oETBHtD4b
aFm5ixVczUokZ8rc+rjVTYdOsARCiups/lm/35EOKYxnNd7fX4tfT4R4+qoMHT4S
NKd7uHPwJXo4i6GI+skZRiMLpgx8CIf7wGO+xvDQLho8UxzBa6im8n4OT3ppQ24E
jK0lIdP330PD9r30+qpqKi5q45a1TAMDJ0+wGL/xVMNXFPn9I+2BERUUEJ/to91C
Q8LK3Ae7hC/vaL8TYIys40kJ8wBHY7Gb7tN/HbYVPuH1tRQ62WuL/MYla0sCgjBt
vEYqYbZrlNLukwr++dLTox7CLoI0e5hE2L6GjzQW74Zw+B+5XYlW11xX8xV94hnv
jjAd91++pwfG+D4bjWRgVpI6Jfyx7AReQchnSZ4DeMd4jS0FnYSQ2IYIfPZ+YUup
lueNQ7E9b6cyVthbYwvJ5rn0Mvrtfod8ZweB5WDGyRw272CZ33rZcJNS/flq5YPE
0NCO2T/qx3xt1EiX+IvUkswe1DIzzkTXNjDT9Dup3su61VzyFTLFRu0Ccc4Om0vF
Vl7hh2szhtXCwpsj8bv2kOpC6er2E8vDlCk/J7qx840bhWu89lUDYxIu5TphRHIq
lNEmUFej7mVcDU18ErM36kjTuGunuw0WIRmStEJKI1hc//PYVY+ZR23Lmq64H3g2
NVrwJW08er5NuDwHC+ezUbZIkBRPQFXwpVYZC64yxJ7eDJZMaXyNiXRE+nmwRYID
HwjvMhiiCoTgDxFpG2A90ru9VE/WPkPZNabO0njFIUuLJizgk9sx7MdSQKChvVqa
vQr5EjHIA4+cA2PeNJCEzRGEU9WdXApmSIHBa56O2qbqrmDK/MYhQBgX7q3lAG8S
68ZpCcZSYI43FEReB9tnB1SSGcz1SBybVZVU2pTveVvTJWzve6hlDQMn77v6OAOL
QcKCpO4ORk9YUgBkTXFCvlXh8riRFQtyLvXMWwzIkgRTjbczgtKsgKRHr+FoHTvH
Ct5xUUNi055A7Hc3mdivujhEcVTzWUwqe8q3AB39/rGA0NFGpQkskgMcyRUFSbWW
`protect END_PROTECTED
