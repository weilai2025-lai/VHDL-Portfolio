`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8K9A1IyYOihnfpLv6rJM+0zyCBQzQayLvW6fYH0ofCi1fP5jvoKybLs+YjMlOad
9M1SOmmu/yyHkz4byLx4C1BzU7sE3TJLuedlnPJR9u63gJb5vonegi1Lak3sJxke
OIBJHzRCpFCfJCrGUINHyvacce0UfOkpfj3cjZA6u+qbWp4Nx20laxyGVWEMeYqE
J5JFq3CCxVHT2e8AOZfVRwaY8txJQnfOVNjJt6Z2pUONsPwar3ugof8gNafj+kbI
Ge6wZ33UMPbOGSEl5HnVurnjqshdqT6OozTpdDM5nnV4otfIcgumgp+ZlsQCrmiT
/z7vbiY0xgQ0bnhyzF6PBeILvPnIl9knj2NA7HA5RtUaMoB1tJoShe6nhzUzZtQO
R+/6HKBWTqE3mPl3RP/O0W7IkVHAv/nBxqmoYDDPP34CSljsq97EZRAo1KRmxcAi
hboyU2k/i3KP37e5qLeTs0mBUae4pDzWGTRh7LitVaMk1QxAwZQOO6g83DScHfNe
+CO2WG9ycwhXlIQToqiu7Isyk3DD3sw327zkj4taKr6VvVCWvF1p0D+8znxx2XjB
Qh7DBsucK9MCk9ir1d2ybQP8kPXt0Z7hl4ZyyjbgQQQgNY0RG9D5JtnC3CzjDdBZ
NLScOgVTw74RRptege5NiWMOW/3f5jQ6hkVBYrEHGq+Mfe/e1uIMjaCpocF1iuvH
rBPEuMx9tdTyUnlc3C6QmCQF09j6zuYOhN+g1EwA+0UXild6d0Cw+oVMr2wY37Kr
6cFtP0pTMNkD7XeDBccKftH6RVl7P8jpucw46LvNzCW5CpR3i3qZuEA9cP27oYvE
aeDL3/JrrRGE1ckC8OW3Xm3Mzd1bsjaVwlyVNpi4rig1K9Sm1kkKLDlY+Pb91uGH
`protect END_PROTECTED
