`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TrCj2QHfEAIkc6Ol55H+CtpqkECKh9xUfQ3iucytTxisheckpMD6CmD0GTwg3rvP
vvqABB+JPS9rBqfBRfzkW8tGpa10X03fWEYD7pa11rchukPDMX09LiAxfgSKEvxY
QHC5EuU032Yq5vW65Jn1RmRQGOpUSQp73Fb3bWWqvxNpU6RlEEyxOJp8xoM/9qSz
Bd9XNtPGL687FcfdtJImFNok5FLwP9gT37bp5pHQJxhQ+RF7zL2sA1COzmZwv38v
E7L6cWVvb9Aju7Ks23zlS+JF3RO1o5LovwER0oaAUK1VkvPIv/BOBF4t3Z6otHeU
xFpAUOdnjqn3ZasH8nOSysw+42psPpAx2myiUNdOnYdj6dfSv/Xia9C4WBPfWdPt
BQ0yXc6uEqGWWVXvdGb+flFflytVW9ucs4ZzArrAPrzaTl6FAF7RExBoCcSaHzF1
F8mtgSiFaElys2dPh581KTQyNurFZptsG23o24dDS4fwvixSU8QbIU+7GDWwcrQT
q3J0hRLh/NYWrPOUIebm3UKfcNm3IdtbsUd4fSwnqVLpnkqedQeTXP/ROLPD/bvN
fStmQGSLncGQBBLhlf7y3jvLQgTR4GVODgCtU7ANTHa/wIKt5cKl84mWIiYseRZL
x3BGGXWOCFTolswoAqSmVlC62bsQBPxcavCjxzd/7jpm2Yw7D2jmVHssfeepSISc
nJSSZiD3goYzj0I3UWLqPhKH3jw1h4pD3KvzBhxXaIZCc71H8hIcNen9ELpzbAcS
cUmWzHNkxiRGWN0BGSDzI/9NxhJvlsWSmeIO4l/9Ik696ckSnKdvRaHyhNSZVRSV
zk6lYg9ePxICzaSYDhH0s5I0wrXuphmMtRC5bTG36OlSUMGiAg7r01H/G/HgtSrS
qvtNCfJLfLuHZPm9UfC8/goVRXZABg6bg523ToqCBBzkNxdyXpRJ75S7JL8MA84u
/kK2LMs3zhcHK6RSLUTcoiIrW40iAQ/fqnFZaMYx7H9ZEwslNpK9+yinz06cIA3T
w3w0rZG+BM3G3u5PNAGY595q+Y1HKTgf1QYBnRT5CACH3JV9TluAGRdoqKenMBBQ
6FU4vovbGSFdpuaMBMHtOxG+Iy4PhFac5gEb2kzZKmCNG12jic+8KGvKYUTF+ii+
5pDdkuUcwbOdXQAtNwMTCziFisNR7JmcaVlElozSG6qrC6ujc1vl+PJNZT6YKktW
pyvHDCJ/eA7kynHHonFy2OvQppL4RiNu9otpLAd9Ym9W/P5EpoWQR5gZO75TIva0
YnIl4QIE6IE619L3aZTZhpdPwhxFsvwtBkcxG4eaBvU2A5AGUo2wzSIqaTJ2/SqD
8VpAN381soz/OJxSffpPvO4ckIw2Yje5wGLoq6+ca+suAeCURdT4nh5XP1kRA38+
l5YfjkeLpMFdnu39Gem2sS5WT8k/FRuNxwXt59Q0/EBgyvNPWpAwedR/O0mVGwWA
jtv0JUnzSBFDp1DLHHqMCQ69Ggw758yh3cXKGWielihFIVdvYSFPaSuzgiIU06Da
tbsfXLkSH7DLzvvr9lnkU4xhqg8IDUpHK77WCiEAA86qq0DQjMdFENz0XUcfoqfq
p08RfZ03FbGrcyz8WvORaYzHRz9dg+sbJD9lrz5EZmRf6MCwp6DXf79skG2phPGM
suDeIlbVhmjrr3dGuplrkAFx7Ocfwo4jOfefFOD39kWQzmHm0bJtQpxiToZfg0ph
UesOvhj6nltCxljgF0hV9CtFUhqQ5OQ5GedySEZe8vojkIqu/aL1enRv+ElZB8LU
91IoZoWIAICN19bSossglX14L16w1SwQ89NL7Mq2iAvdyvTQXnswC9AEvDbyYMNe
srP45qzzfFOWfBe3suuv9XOMonZw2ff1xkWqBmpj9Ie8BMTlydPebjv5u7bCo1jy
ayDL6CwU/i2vcCSSmrrdAio2tzB1SxvyYJnExp+TbjcEYLk6fqLOk7+s33gqcg12
+dcyIaEL6vy59fmBG+XrxE/6c1GvTg/xiQpbM/vsoVWesyIAuqJSAH2BTXWHNPyW
a1R07ZiIyBwrVz6OobWCn0MNGzKK1hZCFXWNXGg1nEjo9xhUVUkoxSnxb5f0FnBh
RL640Ymjfu+ieSENKnYkc2sDsH06UWFDV/tJjcCgs9CeYaqD+ikRhsyjcoR8NTbV
Dx4nNBOLbLPPTrwmgGDQa6ChdV+HOeRNQPtijhxTwCNaaMG7MU88oaDJkmM0Z35V
R3IqzHA24LOU5oyW8WO/dZiJyOuPnJAgVhBPwSnbNuAD5YuBgmaCeZH1lfTCMLUD
6Txrig8aUHGcAKcrh6OBMPyg9LqZ1OOedY1eCMoMA9VuddeHDmBvtOpSxuwJnKaJ
auTNAOGnnxStb2boZb0/RQ==
`protect END_PROTECTED
