`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P6H4UCN+v8k+xMeKTAVEPJjIUvbtsNa8NvRNs5UbCK8/9GnierPOOu4LntQaR8Dq
3q65YO0M0PgFGiTTHBOMZ6jplWbWnR0I+X+k4WNOXR5iUeHJgUJF2XgFAzyhq4M9
luIBPTVbrrOggX1A+d2WT549zWHSDlHf/BX6VrOctRkFGymYcgP984XxBk9ujA0K
JKnTx7lKbxhHdgc98UIHMZVBFl9NFp44JjyodYCwfAtE0eTSDA5hTFw5Oi4kvauU
phM0h037sPDmbH0IfgVYzjEhOMUmIIk60kZmvwmE+91NFixh4ITT6RsED4fn40Z6
rGRzZR2cLq3lozo1hmygLvSyrSj/922LCGXTv51fS525KeZhRM5uE9aUr7I0sfzR
muv4WIIgY56I76cf7OaAPyx20nyRqKe6Ue7+7oZEY2GYrrGCtPblwd709Y7fCEjm
`protect END_PROTECTED
