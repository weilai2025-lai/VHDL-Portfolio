`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6NmlYdAdTB2u+LWOYTck3eJuxOb2JDF89F5DgrFP5yr0PN1ovsH54sv3sDy4PgR
hFmPZs6nZ4Cjw4AgjBHUxW2PIDsmsQhJHg2UMogMKgI97NA6dQdl9Pw62tvGTqvK
2ODSQWAtYKOgsLbIaLnJRR9tdXXp+1Q7uc0RLyYCXrrKaiz8Qy4u5HhTx1aF93KW
djqVEWWarCBrEHE8KqdOTKPcotc92Vx9MDTwyV1k/If9ZEVT3dCxPvgmAB3PDqTQ
kmr9YJOsUgSmnT/UxPtoDblEvUY1HQe676I1LWlOpq5teP/I01UD4AQgcerdpqq+
8ptZ+e0sSxqeVvCKpxiZsODnfWY4fZuYt4E/CTtyNNyQiI126T5YqX8dKnCmohDk
mOP7NRK3pNATgIo1Dk5Nb38KZaqzPROTqt7l1nnKHJET6ZGwT2knjMN2OBZVjE6R
sWQrEfPR/1eAH4RnaxHOK/FQcYhzB9OAu3euaYlYxJoNjx2puqUbkkAfsToNRxpt
/QmNtfpSDD2HT4BYyZsK/VKlWlEWM37n+XScTw5+smE6Mvct4/8c+mR+nDKmrOsx
dHusSD0FjRAVhuhBV5p3QA==
`protect END_PROTECTED
