`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjYHKPl1rQUZKR5JzhK2BnMYv6JuQcB4v0Dgua8GEj4aJ8spD2PcypUobo9KIluF
CK4adkp3bB6u7PE6jNWixmLu7z6pzhxVT3tNCisrwZBF3B3yrZj6K+Lc/FAfRorV
Acktvi5psPZo0oOcxhVN8CIi0bYdxA6Q38IkCtTvekqrsors2L0GsY5yeMirg7AT
1wnh9oUXD5iY8zJNvDQQC1lzArnurWV2z3wKYsd7MPPTboNRZsEjMevD6K16Nc3r
lQRDjHryUje0F2Rk+HoSnd3zgXb/XPTFL7GeBt8OtvUntudhcb330E51qClg2jzb
7RFtTdJ9KapVDRuIvzxoBjf/9TLgG4am4K8Cau2rYJKWYcx85hrDsJbe0bcCa11W
923Tyd1chIUci8YT94JdLZuaNQmj3cI0VZYkOSseTPC8Scm3FAgAbpfd/k8pbfND
c498ps2WFdlud65zlGB2TAy/vgnoIwp88nShtNx8Jev4XehFpsbM83rwrolMWyNg
0vRd8UGWzFi+52AJVe0pjGpcpuMZKGh/ePQf1y09A8iteMbqC07hkoYZ7xgrSlHH
B893YlS8r2cJMcs08G0H0MqpyvSyfSNV7nKTE6wbyR5tlmt4YBrCGSwB/sOiQ24T
t0lqtQeYMeSKB9l5v1PzaDec1/H9n4Qxi9Q5nk0o4+zvu3KMN+MeIkcPP7FFetk+
ZCPZLbmjCOhrYd6rUu31R6ikQPZNn4w6yZbMc6P0g4NWqFtgU7TvCrlZfBdmcuxW
Ir8X+rCK8z0ENYLRMtTSzlO8/Q6xY4/F0NtEbBfCVJ1KlmCMuaRo+LNGlocYjHlL
Vs8WOEQz3SjfkqsUTZQHUXkaTeN21ScUv4v+lKwZ2Hxyw28MepIgrR2Sjtje27X0
R2JSz6iw/izBzeIWysL+de/b68tvUdlz6UR2wJalIfWc7vchCWMdZesWxAPROHiv
LBWB3rgvBuAoCaVXLghwKY5Ki42USl3YvAEbOgiLCCdILRnmz4EGkat2QTqJcALI
2XWikU4E1COQZtNLbRowLDdqNzgh+te0ulxQM8aSUKpN6+jThKeXL8G4NKTJExvT
j8zjD3FYg6US9JL9LL5aTEph2BqOR0LrirTRW0qanch2k59dwd6a0v1/FH7fVFMW
rhnqfhYUs/Cb/4ohU1nBUYy7rZTPVLWSxrPba9PlmgjbYYd2AKGQbBU+HYjb7ea4
C5rCl7CAJAvqzPutDlQYhvnE3CVBk+Tet/SD3pOsFLfKdV63FRe0TMA0baNe0jhc
W4/VZSJd7CBdZE0OAHgSfeJ2qpfQab84uDW5iljqrLI58WWmYoOBMZzFf5pC0JC1
nvCamkICc8fh4HREL2I5O/PDURfPDLk9uUhzsstuAdTFihkS1AmIiwrVr51oBQTx
oHfl4MFAMWKN3ys3E+XXNNYktkPzwZMRNLCUevcDzVy+OSXiZPogfrfnBZbvm8Iy
ion34DLkgtZ+cT3rfb7NYg9ov4JrGZ23Ehzj7VOgZVDI4wTcZ2/Kk4DUf5oOFEy2
/ptOINDbY70pwpZXS6McpP2OKcSXMjlFwx4clbP+HF+2f6ZENiIZhlQ30FkKWpjE
yn9pnWj9mrCfnOKK7KfGT75KW21bWmiVmA5w2V5bADAbZ2+9I9/CNNI5Muwr6r3S
y0B/4bGH2zNmvcHzEDoaXcdlTOODUy7Sto2dj3zrf1/DsN5D3CP5fqxXDwwKQ+t1
jTPVJqnraXXSmUJ2SjcfdbjwBIREb0K4npsEbJE5I/x9d1PhfWBJKqySd8EntgHW
7NXy3yc0BvkWlnxxyQOkdzUKuSBsvhConEEpp6M6WSrFWkZklIb0j2Npfi0FpAk2
g3m2y/fqUErTTqXJDM6pfD+/urZLF/WyF+LoBxT1ld8wkm/6F3p+XecbRr8uQBlV
8NAOiGQhWzgThHmGy06th5ARIXLxYJtdhRuHHOIHRmhzPuzBjCaFGbXbqzYESKpC
Q9UJTDwzZofecNYYPydqPzNWAI1sYztyLgzZWFN3pOGAILxTUThAOo3Wij6tOTpI
5Bk0oL+miFXyQYMUT/Gebrl2b4x6qHBdi/pnCGsOf7oSyjhKFkZjdVleaiYcIFa/
fRuK+T1Sf4tCDYjGQR9zgJsZUKAl6XFRuDOdI3eYkHDKZjhwrbSN2xKDG2lXWq1s
o1fAVTKrmOaxxe8Ysu3SsoZB3YBndaTeUuimngUvCppQOJmg/3EgVpHW87e0kGk3
eEHTRYo1jNnKAioNF4PocoI7/AwjaeEp4m+ibBYq5HvG5+ddQHkW/+YCeiH9xwnS
jtIbjpP0JjvP4PIzOwyIVtzV0Kq7i9U6aQb6HKK6PKIDQZ6fd3LYgKgjuDodRayU
iH/QHMw3X0BZsWhUWdPlGz5/hFhoSlcpQf28sQl/gDKHeUIELcxK7kzCZ+UKP5xT
/Zf/IgjfyaBAegiGJtZQPpC/ROxIU8GWHRjLIvZha+iKwJ56w/2Zi2LxmGUWj3hY
pbbM7rmgzWIgBNjkaGk/mhFBFzH6e29JtY8u93teCHmq1E+ER6Bte2lf/ene/mbN
FAtpK6a7ITZ7ThEy70PfQTvKoQp9uaF8BsDKFYRe/Es1ficrm8B85rvZ4w+mF7jw
EUoHJreoPefADruqDxaG5SnJeJUyyH2ORod8wJvX1mL3uoiTxtiduXtEv51LYe+m
5MFF4L+ZQs+HQnvHUDUJJrl5781knlz0kTORWYX/L1vDM5m8ry6Vg5S7hTlnblpH
kyscOdxxLABGCGEMlCqyrMvjDDUtKwxQVaZIvbIaX1eUYWwd3dDzLw2KRtvLLcs+
SxuRYazqKSQ2SI4/JyrN1RsMQVsiKqUBgIZe60Scjk4W/UY0vkqPaisXPFrCq/qo
YfF2ODRlEJfefWv5z6VtgqnJ+oHuvh15AnCyxmoGXjTDMm5fV5ke6DtbeQPBIPEf
JRSM1zyX4S3+JjCYl/e/DSmyYVjMw6eSUCWjWr//XYEVnIfxCY1J3EuIZgCqI5CI
qw0pFtYd0Rp8LvuGgHTeqBcCWihcl5ZLov4vJbsh2p1DoaZJCmvndXw2HyI2t3Og
MGBwWg4GiLHSbiB+bjqGZuBtZmf4LksNXALlh2pW8sEVQpCPZHtTqwkzEaQJB1u+
2+rDiWvBZCA3ruxb5JMevuKv7+3fcWDRSwdyiJ/gLYayMepdlNtvp2Kg1EHJAyOE
27+ZVkub0R9REsb1PFfMPdB7kFsFPWLG8sx+MVNrPf6dp85Xdl+2BoZxHHSNr2sa
FeyDb4HZzXrIgirgZLPJfGfJNjPjnO62QOFl5BGEMDhM2SBvy26G+lg2aOgazTn6
GmOYzICVmLVhWj2me0Cd6KGkwnrG5dqQuy5m8LDwbxASYEz+zubRG6nVNDMwqvLr
d9bCMdeZT/dZzGqhmI2Ciws3puFsSirRPjkwRqSV3+MJmz9HsNKk0LFfeHGsEqvi
DKxc0blm3vaYGdeVYDD9KXW2MiQ+stkKUV9h8sF7y9QIvViABwliPviYA2dqpqRm
G+lzGRfpuycBqbWY5QWosasoX0c5MSxMvh9/aZkvPvzm89UAjJut/1U7F/zKvPNe
zZ8rniG3BsQTFPoYiglYeQQlbO0ECpdMqwl8EKbHwO/a+cC372mD8h0uV9pPJaet
ayUch9Ot1OxOLkv1zXr3isyR+vw4Y0pH6TThR27MKh7ZTY2rOlHdAq640KBtnnno
MMyxfeEs/NGnJLupkiF9t1D5dTY2Izgp0FNOxG4/PW8KOMhmopWjNfJwN/wHFdgw
nvX/Zz5taNNu1sgXfuEIt1lrTtE3MYWS58g/hsqzX1Dhjf/6Hup1IKwskPV+maqJ
ZtzC35FsaOSIJThXm8O6l+esNNhUkBuGWtMV9TDVYCrxq2l53KPwj5Kjs7H+DPl5
ikEkww5XKsqJqesiI0M2Y958GPCD/+JlJnTX05HAV28qK517tgtmqmFZPU1HnrDy
VkTCtosoMCKo1XC46kfOJ9/ovCHyZ/NWaM9zd7obT9gWGliWRrvVsj9pRzaTDQSz
gzYwSUah+cfs7kITB47YjacGSE3zTCJmwgdczS2/jMjVqHD2n3TTMc48HkMu35VX
dOcHYtztczjkfboFNgs5OVqVB3xB5d3BI+Xb8AZfs12vOuu0lkfb4T5PVGuW9wH4
cF0PdOSz87hRfW/tVT7OIeNSEnk0HeHuHSEgNxxSCF8Q3NdfL13VJCkvtXQUDwsq
kLS+AfOahI6eqry4rRA3/hF1FnUahVcTa77aU0n5VPxNSbO0vYxR9YCSeOE56lO0
lh1bf7OERoo9eRxMVf0qJBXItIdJLdsW57GlDGiVaGtI6MdZI0WQbzDXDi7STdfg
bW02LLrTl4WJwC9puOlo+d9Z+aEe8daSNb+iXCKiCW1zpDKVrUHGsQvHnES9k/1E
RonUppkJxUwlY/xSmdlP5ui77w+K6N/YmWgJT8VAbiC4bf0F+rIkHpeysPY6ktuD
OiP+Si/FpSzw1XGBCCzHuUVi59czk3TJtRccYlaT5cIPKmCbFk2v24cxrjsnGlPI
lYX1nBltp+He5VLt2O0c0Vu52XTbXqfMftubg1vL/xWV+cXt5QfTkKC8XT8V+dWZ
hnOtz87eBtkWYR0P0J1EfF88Fhk7OrbbfUgAU31iIx5ZmpNqgvWS7SB7wZJFvIGM
dDG5YtPrA+ft7v897HqAhNnw4WlDzfMKZgv92dvtKp1l0I9ROlQHt1R/1ke3BFrY
6VqX8fN+paUyMSEJ2VOua4p6W13q22iSlvf7BoYvAv0q/JG6+sRhAAU7RqhsyTkU
8s21dgW7U5DlUdiwQ4PxZd9zdLq+XWLMMkp9xej0+4Em6qM/3G3fM/rdccD8GOBJ
o6p2mYJ9TxKTmpYcjggkwjLy7cmlPk4Nv4pyRW0d9U0AGbfkd6RxtA02PrjvOOzh
TNq9Er/7gZZp09NlVOzt920GyWHsB3EMmUVx5ENRdGbY9AmenZ8Ng73NrABgeLEZ
ULBv+a+ralMCgeDF1NRbVsIpG0L+o9t1c4d0iWUnUeSfOAy8Hor5MQrQ3DxL8UXX
FqEh51Xox2FQXxAtX9r0KkQQlE0s9m+6RNY16fyampiZ3SjpaylBp47B0V8rV4wi
fHtCx5xyAArb1TBxbB0mpK7iUhM8GBeEtIARcFhzgGLMwmiMWRdny+1fBzyDeyzW
JowsHRXJt72iUvOT8ACw/9pe/XmEuy2SJ1489s8DNoEvu5mOrMAYzPpY1kqpBzWK
CVfjWucY/fmrg2o579AcWrOgsMW79b8aovEHn3J6ArAyVZhzMOgug7e9rReo4slF
EwtPt5O+nOmWCV2gvpkXqdTsOua7v5SlcCW+j9v7VefXNMmX2HFRuIoNB/26Sh12
DmKuztk9qNrTsE3UCerKUpfKvN2G+XGCUJH/qk5AxeZ3ieSaedB151L4OktC67F8
xWe3gqBCb8tydzAXfBSQc2Kxpm3fMVszloaFlNIy9tpgZMH+u+B9myTzk4iqN5oy
XtMf8Q6FuTunn+I4eSQmYpQYCaU5S4/SHum6md3DH5/8FuWqKlzMXRviFe0JUmJh
9Q+TTWZkDS4OREYMluOEQPb9rJIv+BAp2XRjz8HC8dIFIinQAoi0JfyhyIr22zsI
kAX+aKc5tKW9XSm7tXxE+PxB3SA505mV8m/ihk+OegRXDCtivvZXFxspe/ReJnPL
8uMYZfRNjOkvyDc2MdCU+OpR7tI23inyAu0tcDjOoHOBAtdeus/7jo4Ir2+Idaob
1ddFU4EavfIpNiiSXi6n41VFDLA0uGjJg1YJXtXhRLsqOvX19Uo8LVump4sLf2YZ
OLINEY3lPDPi8C8OPKo9cven1+ni8WZqb2EBktJZrvlmpKI2TiZTAYRcKNhEjeeA
mHh4o1LZpfkpo/7KRAmbbMrP0d4I0DUgVC5R9DKMyrmSNhEaERDzKJM3a5Rzxrpm
GVU+U+sRwM2t3yKAaZeQNKPrMHKoLfxh6vfNpOU6C39Y2RRnM0uPOdrP1e+Bj7RG
+i5shO+RwIaAP/JEfG0MeZBTAjZRrgDhrPO4OetmU8fEwifL6+2dSyGEuEqzj+oG
qPsZfKqT7xJGOFX5LnoAL1duDqvVUsMaQCPUC1qpk90xTCtztMkZcDQuiXeqJoZr
HhnUB1JuBSs/KgATTuZPtEiP5eGzxr8I0fH6d92cnTMr4JJ5Xlm1G5scnyuZ5nOI
I0MSRs15DqZtFelO8nCdV8AJjfKF9tt2Q25g70jvJ3YjrMLhUFmnEzbZo3TcZbE7
z0oabbTczkgVaEsNN8DXG82uw1bSxaFeCkAYYULJ+rTvLQle4d+liq/IFbMpuM7t
KZAvaXdKEmCSJ9p4feV2fPmmEc3xpLVhFm5w511b+4x4lKAcstNxrx5/qCvhoeIC
/K3RJxc3cj2d9bc/ZwnhEuMBX4oJ/fuKLsMCTm19MlkIvLw3+3Kv+DN114xndg1Y
hEE5kcolYMuL//j5ashCQA6jFSHttehKQXfpo610A7kfYgQ+oCpLhDiqx6gH3EJN
I5dE8wAJDHM2rUiFJZyhJktQzQPAnQf8JX3shEphSAyHPGc4F+OGSRgE63rqvckS
fhX2Zurtjzd4sSVCSz2ryTTcBJv+9XV6abm+MTVyfraOoRtCi2k+QyUu2Wp5Ge2f
hNcmTKwYKbpJTt2FsR5qOgTD5EfU7ZMzcEgHUz/mfPoU945r54W0V5qHurQrAbUV
9kdDtm21km8g742VTgtfXJ8cHONpakGMJvDJiTLDKZI=
`protect END_PROTECTED
