`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KemYGkjtAfOjnmip3kNmv0XV2hihOEziIYp3rB9XZKPy1B8e1z8oqx9GvPI9X7L
ki5wnAvmjgbBLu2cSFAJbpHuA2F8iVTFByJYYPH9QomUuWZzg40p/h+/MtIvSryx
12UCJ8uURiPfhblJvMtLRGB9OJQV4JpZKtEZrbizV5396vYd6OGhrHKfdrjLyK+n
DqLFfFW0cORlisCXjc1+CMJDM/Qxko1rl7qT6ngCg8O/RnvqD3ooa7N2V/Os4eu9
nweWq9UxPcSM+O1EH3wFczFMzYDAXDJY9SLj66csMYWzDRhI76Ul4bjK1L3TStxl
UpE0JnPJfMFi1M0YwjKgElkaSRQSH9DfzExZpMyiDBhutXuDXuo/6xIwGQ/jc+HS
`protect END_PROTECTED
