`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+U7Dw2DHOrQDTtFPoz87qjrlZ+Irauuv/KON4WMuZh5LTfB3CjJOyI4VFCOsM9Z
xW8CYevICdRTzAvjTkZLqdgARTgT8Y7L2X4LXZFQiVMFz4exViwHeUwwaNGrUtFR
Avdp3ZN5W36vQODb6SKWhr45rtWMN+30A+oqFFvexHEy8sDIpuF7lbPc3/XgMx3e
1ELZCx9GFiO6rptfGe8EZN2YBqe4XOCpTkU3aS3f7M4gGmZMq8IKk8rM4sk3HGE2
y1osOEUA5vMXFG+fdF4ZXRQVly0+VTZmpnauzsbVVHswHGWsQmbcZhcZlDRoQ3/r
kV4hMj4BS54WRl6B8MZqAD4nVxQ7MbOGLriSyyFvl2mUr33aJtntUZjQHHvReQZ/
NaIBPDAY3+4MFpxAVr+uetVeQrvGSEiUB1qXKwQvyS0+ilyynXd+lGOBt+S4NorF
M4Qee7ak0mMKEpMnJflCamNCWtpgOr7XlTDVvJpHsBr+BNrb0YnB2eCV7sp0oKPv
v/hXucAbWzoP0aySXJnTUuN95jiDyEtWpx55JsCtgvlehExxyTPoPCQGcJXOe6Wq
9PXAejsm3V8zVETDWYSdK24u9IsJD0yARHMzb9bH/61dXiPjqP1DgiB5nrmCXUgU
EJVaV11Cl5c9SHNNhp6tnBLiea7SgOmQF1dCBH9NgueVePMFL+htlCt2PwWDVy99
6vCAenuqqrjX7vhKYbNmA+JT78D4a1BW8F7v5eZ8VoKSQXc66b0zHra1bqLP9Tzr
IBhhDF4+ZiBqOt7btlmVWxVrWN+i4rGr/gqNIw0XmFtbAuawMUnwoX41muf6Dj9F
9T98hgmNYoyilLGAO+sWel0/mqG5ExNylBsetHq0EotV5F6tCyQ/MjsaqpZLK8oh
xeYV1g7+Xn6iFc+AJndlkilzZiBKw7TmjxEWpBaKc9Ejwk/HchzJn9AZwBRDo09W
pcas1yBp1I0hYbDsLhOSEhEK439Y9iEyRkZSj6ycUkGeAbNtukI74ETG+8KPCymR
7GXLERUOceGYhR9iwyLCfh/sFZxH2m7/ahOQFUR/+6RZuFiUPvHX0dkmycN8UKcp
C/KQ0lIV/NH/0NVTlWG+4ZhymyUBs7PakUSruJOeKZB3AuIJ7/7CfGEtGrZTd/V0
OP8Ru4GH1VSPDPQBIFml14UnSVvBlUFVTE12U1M4b8ZRAxexC8X5HD+n+/YuBvCt
A6uSVjqs2otNlUPmO5dSVIXQI41qA8RHAgvTZZDhtYIgRml5tRKMNFqU1gRCJhD0
lQai3HpchOYUj+CtQWxUOeClCGmkU5kqN/P27RELb5EaztF/kR9FjHp15K/edMJ1
SlaWmUK3291ZddmnPpmWdm85xahd+a9Q6MNM6zLC/MOiJ/BawJLJYTmD4JdsZh+e
AVcBPn4xYE76wEQ4G3N0crZTB9pQMx2faG4Zrdgv+8CXotMOoXiM4hEqVC4w3Ohe
BXhCSgop5bab4nJ9DFN7EaMSv0jMYmNEDImud8i83NDfjYDtc31CvfiV+d0BffEn
nQpqR5KgvVZxaNO54u6kX09Nht39IvMOc/pm3bT6O9m7og447nDd/AmVPL6l8lSp
m8uhsSiWXLoZhQCztvWaeKIeCIj3sOdxa5MQhfqcoAAPA1l/sH23ZBcmp4L/E748
1uPRIB1eAiLPAsvH+QgeV+UHMvIppluXwKf15C5Xxwv+0jZDsthS9/XhTitLqTCH
QKdYOnoCi9NmI97HHoxMzLdwqQiTLH1y0iaBLassDZmARCIUHx6/AHdMsVDZWFHk
R7SoiGLwkgID3Nt0XbRvaw==
`protect END_PROTECTED
