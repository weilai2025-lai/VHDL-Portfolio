`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LswSmcQ3VuYXWY0zg40qxiF24twSZ/XMjm7XGAjUctlWXnogq/M8FPFl71CIew5
npmjcMLFYAHYdFgLlThqzq8K3LcQPBzS1/+ZmTCuYJcLGcPVEU5u2w2xBd+fb5Pj
7C+fHb9mchrj4GJA06xcn+dKC9Wzm+5FLq+D8x6/OhN46ARxbhwPeXLi9vIqwPwX
1eoAGXL2eDUyja5KMdDiiUW9vS4W9Kyv75GerMe/YQIeS25ujk0jF3x1p6D3XHjk
8emSaWm6iSdwvONoril/8yD21kCMizAYhRK4t2gUO/slYyvsggg/EjPdTlTKP80D
Teng7kn1u2DaBG6+oiVMgLAkFu7yD1Abk8BdaWe+ANbiSwbGvcOr9D4/GXQuD59i
AVEOFD8MM83gIlQNClS90RHLGnYhdRe5HUUe0+bVXHIEhRE88MLe5XIP85uot11h
w8xFcgMWhPBVzSlrSecrVq69URDN9TnC5l6ieFCZQen5igaNhJ4l1K0m0b9OWNRh
6cP3o95n0MAGB2Aj8DkdEBRdHFLVxd5R5eu9fTUGi5uz5ckSwpFGTxdkGUydv0DG
fbdUcPYK9U1YiECiYWyPXTWjekhFpFm13E/rqa7pwt43vd+kjb2ZkZkGPtAwl0Ib
ZjZoCzHBfO4R3QBDTTuQ1KvhQalIZDGGHfyQ+AUBr0N1wi6OM+vEb1oEC60olouB
oKYDKfeUdGglrnDKE0uR+xw/iDscOWioEgghiyyXXJHUqdSqJHNqwEZQGOhtEWgr
+OgwW3TH7svPlwk6PCfeUSYpHOvzMRr3/p/eAmYwrsy5x43llqqWyBuVkOs/+ACj
NjiMjmKiqgDYyfgHaI/eRq6nepoqPrNYvKdqXSv4Y3CZpA3Y7idsIufOwbznlQ6Q
e8vW8iUlAidTiA0HZrNGivQIOD424Lc6U8pKw7KSaTcmjbs24tvmocWifgHAlMDR
LOKOqq5n5JdPWxbYDwkyHW/RLZBuAMKbjG4dfyVCYrRCvwKul0tx2hSam7lZ4qjp
7+kViF48bOUbAxFj2NBBLgcpDN/gxU7YeW5U7a6hUXA/cFnzi6nNWtEzDoj624jy
+uInMxATyMOsTMdnqJD9iNGmU16OyJOFHXJpx/3GLhtrSK9bpoC3PWPsJcrmJmXE
KFgXlaCAr77MLKxMIP3xdTByTQaBSVM/ThbWfgTVicE7xf7oUJLaE7uqOs9Ljh0E
UpP1spKHJHWQrpt6I87PBQfrG0g4iwGuJthQASVv6Kz8hT10z4fLXyoWAZCgxY72
Z7GYBr1PRu+p+F+SATPHW1QtdSAR1TY4q+ojS9Q041iWW4SoS4WQaL/vIayHMZHV
hf7B75y3UdbENb3psVqHQieJClAE6v3FyEoHOcMQh7TveJvhHj234Tk1KxsUoOVR
Ia3NJfuVPQGYYnZDWcUBCKUqXQwRTDkej6mDjEcai2xi7havDYEpewO4iRqJnzol
vX3J5lmrJkGLb9WrRafYmqbrDs/+xEJBeizLj/m69hxYUbS6OfF48KQ5XvmZ0mR+
IQku+Molp8dFhBtYoOOHqg==
`protect END_PROTECTED
