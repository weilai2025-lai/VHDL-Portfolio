`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIDupETQDGcqgsM/ozdc5gwsGHn57VWN1mj7nmrSoX4SUP3eQp233nquYLFhC0Gl
py5gfrNbLW9yQq24FfPJvXXnVyc1i8f5pHRFH8b8xcnfhwY80rAWZ38sTsR0LdZM
X5TaOy1yd51y7O5nare+rGKehgBK3xGU/gEU6SOVfZjYHTLHlIO633CPAD5BV7d8
YcN3hIfsguYCymurqk2k62f06dFFEFQyzUxecj4N1MoP5YemXXWphVd8/yZvMqlq
SdqV+zhBAiq2QCykG/6ESCSWgFlF0RyK3HdyzTv1irHSFWPijOg4nFEFb1ZcxOXM
QvIpaKlg7iKY++jNfQpMf6IjjUTEunk9gqiH+aLxyx5JuPNi09H5gHpH/8XlIIS7
kXu+bJRN8LMYS0YdjCM8dS+jXp9CXyjTAqVMAWfmRp0KwqlN4Eb1UD8bHveS/YBm
aFk7dV3Xg7SPET2Nwq2UoFFp990kJJCxeLAasVIw75HMToEcHHFp75Zzi1lULBvd
PhOz3epCyPSojyCOu0cfuWqMMtFYnqTUN7V/0hOg2N+xBZZ+8k53uN7Q431+mVKV
NpR8X8KCA7CmVr9TYYiDZQte0yZ3XIe07APXDLc6tTkG9WLxrKu+ICASUbYBZBOu
I/ms4NGWkn/KZiQ9twjy4bjFEH+8S6C2V6QWoASgyjokgRIktzH2N2LGpCt1q0/y
MF98Dhz/OtwkKFKOfzXbHGgsa3Db/chzgWo3BuqYI6N6dz2izy3tJogX2XaywcI6
onC2kGjt+LiZOw4fdmDUnX7cC83Ie729jja2kSGY1Bdd/GN2zCpg6e0aKwUg2a1H
Hm+u7PfFO8wvJljhsO7nGUo8kZuG5g/KM+GzUsOonD5nJDjguLNxCQS2UuyU6/Id
1ZuTJN0ONuhOrY93z/6Sw2hhHjWEJG8EgihYVM8ip2sy9aCnoXVBPGq2UK2HzVe7
iKZDpMInoQFgQBaju9HF3yfPtHaBzt5NnWlM9zP+3PCJOUJrPhVPWSDJXoRNdOm6
gyga/yIF7wwAoQWGZ/kr2C/c5ofLx9of8OQAOdw4TpXNZlE86GG59M2Xfa6V4Kx/
ZdHs/6ZgGaVdreiAI0Ylr2QbYPQTgYPvFyTb1CyzJNfB0dVF8ZQJBhWwkOeE/oT0
pG3Ysim5IvvpXeEzR7qefMMAPWM5gbuQ1cvP1ATq5fWOl5yVuj+tPvnw1gfqmnFW
7K+dOCVwzuCSGXDLEyD8NUwc/5L5hqHoHbL4v7nPhmhw7ODMR7YZNmTMgXWN0cv1
NBhw5vJTjuyaaT2KBeXOxIRMtm3m1k0ZyZ3vqH6Juw0en0oeqq4qtjCDB318o3tp
LJNpBs0jGln9Ebs5m8TGKpBXgd2MbME8UTvvIVhYw17OcOWKxrpiDmk54tD1F8/E
PRrKUNHKWBWcBlBSbXtroy3+2GFCsU6ziYQrzhwExdhsxwODNsB45HLv+xKEdoio
QyGRi+eari/JP/PHg7y3gxaErJ7/qlkYl5chHAbL/E+12ZMhjF3z1RKWyPi3xCcD
Wkodh+22mnPe5nVb8g7/Q2zXLVzxu7byzZ3q3M9saV6nLcNt94mbnbPUCSN9a1ix
N7svhTeOdgLGjSeI/JPg+/Uj7tk2Wo1+Ajj75oMelV+in68qFL9Im/BDN/yksfvR
dX54aNF9Nu2NVImpCcDtwz9nyeHqYPeSZHU8567cnmSWScWV+ysFBCerNtdlqyN8
zSVl7Iqbm18xPxk13WVdDvf/wEDtG/MKpLXSENDCN5AxkwfoCzN/8l88vZn8xsba
6G6UM33CJDZ1MLhWdCTDS7p7y5OVHKjeXdippMIlBBGA/F0r6GrolV7e0WeUa3c1
ndtGCmyW4qOMetzlXahmmRRzrJf/ag4iq6RwBzNS7NKCHyKf9cRVKHZ+n2BzS9pD
y8yA7x2JnWg9yc+CCSbHAFxgALn/l2vON3PwUCoqAATWislskJ5GSe7OTGCorn5o
9kVnFFYvtp9r5E5sAT+Ue3kgcvkS6fSBqtVUZQbIpTi1ZFeFBCGCgWWPQyeCQ1eE
3wWcjOjCxFbMYdQfIJqw87/Vz5Q0KXZLn2jyzJi5K5/ZS8AO/fpVOFFHymwfc3n2
n/aaqBH62ax5Ti8tMYDnnd6ky/L4ugjte+yagRzJmr05BoPw67YXCkVn7P2QmCKP
7ZpQn4gHAomhXZVdLxap4IwJtj4OD6pbBWe/ZT7W9DtfC4a/UsMQuDOQVoR28nhp
fYQUd0q8w4zbv8cjpNWjzPI91e4ovqB6jN3u6TUxUak1NHKQUREtzgClgCNZlN4c
4e2HoruqJTe+FlZM/qzaSxnYv/48ry9uFDScLt5oXBugLRtb/xwjvxSMOqcG78RW
t+tmVVjit94v2i0+z2PZxknWo3K2sogmaCtGWc7iXHN5E0o1alnoZpZRLdlRu9mV
Z66oncrxdaZbMaXw/apRUTpmdU7+jIcT07M45BDfcZzLLq2A6liMki797VV2X1eG
iiHWc7V7+kEOn9xaOmc6dWCCb1qH/pqdnTkBrXOlWO0s4z8oFwSqhoApAsNnw2kr
7eNeBFBhep1B7g9wi5RV7fFCAY4IFKOzWRu0TPeO1A43461guErZ8l+tlOBbK5W6
PiYAYe49PV/JUe2cHyLjvdJQVjSGHdCUzZ0+UZIBNi0jbk7u9AhzRZoZUggEJijf
INjNV4Dw5lscoOG7GK2czq9tkgBrO6VEXxt1D5k8Y0tqsRtdaaBaU/39Zd0dl3Xy
LULbsuEZearHfU1HachPMVrTx/AAGCyFja+QmsbY/Q2le4M3up4wbhv3ZEQAVYAj
tZYL5aqK+0xH6PVfKQgpEDbILBI3etFFCaiBB1cL3sG4FWGkTCBo/S7X0kTJxbVo
O4v2peZZmORYDU+FPcuy8iWboYZcxGXkVevMCYg57NLTXMesyQJaKyomLcpqJpLT
wsh4PiVDTz8G0vHa4HjKDq6lBgdiuQN6A/X70YFq25eP5ibfEleQMdQCO6SnSkKH
2SKCESm01nlC8leg2O6aFSonoyXAG39VogRDaDwTTv+valf/2dDMltDLtzQjKLd0
opufO6D7QmWKf5FQxAL2O+7IMg/sXJkw9t9lDQbOl5JI1kqkgzzqoR/kYZ7Wbs6c
PrgV2SfnQnYslfKGTMEICfyZhkPhAVIxG5+jWq9o2u3iAa6zxzvyDBQCTUI56abl
E1P8+NkVH3QAkFPw0nZesM1wnjvy39nfYIHEysguFZpHIa6YFZ5GsFUW/OBK9wYL
ntKrU2L77HcEQoXlVh+U9ZMxrpR8LX8tXiB30T/SdHL6aXjsnFicPq1UfA0ngUj2
zsUaju53cTcPUhM9zbSm33e+v3k1gvqqP0fBtfF7qf6hQmkuWZTHGC1eMritjHlz
dz4f6fMWh0gj7519E4Jfc+UZO4khaXhif9wBtqEixJ5cYcbeVEJe8a18Gf3n7ffq
m+H8r2hUTyQm+geQErfrme11N3FUtzQah0gQ4lZZqDRE+oZsZCuWu3HC1U1oWai1
iQaOr/CiUJAFaxXSp0VAn99zJphmYz0FCJ/jsia0V0n76FCoxmgxybRz3KeTZVkn
fHFHWQxHT9xuoIUgACcNJErLlocXELhWMAA1vs6Zkdwu6YR0Yu4VO15xMGRZ3c5B
jC20yhY2GSD4EArF1CHziZf6in08FxxPPK7AADRRoN55NqSWMh6vEk0zSq+LZfKn
kNPSePrKO7+aDRUBIGxxxehOQpqTsrxagUYurWg/VHR7fbArbPOrTPAUl6jf5s2U
W/byGNMxyUCpPc9n7JM1G1/aZiv8uvTuNA9MPjY8rbhck61f7ATFU9TK96mKnV31
6xdBmVG680P9tdcORamuxeKmocrtGZ5IUi51aYjiPP8xZ9LzVZFhwRXQAyU+QmOh
oixfI84GTnTDCN6lVpU2pFt8qH8KHYQq5rEJ0qkKoxpJQKoDOh18gMjpjMgi4UgA
lvoNGUaVRrsNdMXwRCD1802XP+Wa9EnONz5yGZmkckPSIMR9BHRiSEa89n6YBGFj
qf0EsqM7jXaYX3gt9ULD9g==
`protect END_PROTECTED
