`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzLbISjX2NGdqRFdMPI8g+sJDAmFMBtraV7hoyXxl8ypShY8SyUILeqn0//v9NsR
nSkbEmnCEmpdI2fnH7xQwSzIKT7+b5Vn01hZHjiUT8lHeMKkHI8xwfu8z8UMs74O
Pr2FG3kN2TsVrZNVR8hVdfz3sKiMB3XZMmIkU+n7LZTGAlc8+9PRLp++7sY9kXbr
weitZgp4K304FbiWArvWKjSW97U8//wqp18bbl174+J/heuzREDudgjY59jecW8L
fO+J93OdpZkZ2f7oajKNwhHruZV5SzgwH8ZmSQkfEGg1xtw17sABXOiV7ZSpZZqX
5Jc8Uyo8Env0V+S6ac97FxXfqJTR5X5EGCKx6XWsuzbY1eERyGXBWs/ZaF7Cm4xK
uD+Pij28ai7FMs2/tJZwzCct3x0NGGFxd+SqS99CWbBiqV4oDcZnZHhNG2WBhAlO
zBJUFIHw5FjJ80H+/xuYhTTt+JGb9fws21xfq821zbUQ/2zPi5ZgA9vIa0RxgkDD
yj9PsZ4qtRAZThAiFpXtQqdBWmmq+77DsGPYxRqOmhAkXHpghd1hwxWrsPtdtDvd
7OaNqQxeANPM9K8uzgP24zYFrf5ZhD1kGLviIaWsrEf2N4PxpMBa/23DBlw4/0zl
s+xYH3KVKgQ7WlPgcnBeVMvvOJnU+qbO2rFpYbB7PAsFClatLpG+4fIsqgty0CY2
XBFJo886+Ysh3+YkBPsvM/hH5cqU9DL+hbkIAeaeA2E/fG1hy/WCQARZdpWGTy5Q
hmdcGOPDJyZ8MU7vDCpzlmjYjikh4cCYMAY8MDRvYjzgQ9DEEyV7PVzWKgAc4zbk
WNwjneAL7SN8bPP8IrH29a89NP9E1sPvV348PujvXQSL+p7bMuRAItX19W8FjvKu
`protect END_PROTECTED
