`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kf6dKieMNzvms3R3qtq9SO+FJgek1W4V/exKlXsa8S9BGziYXNntcwRKqcH+jj+G
kvT1vP9nQvOhyTaMHT7nUI9CaFHtNLWXcIkU1hxZ9o+tRHZpJl76FrXbI5UnzGyW
+BmeaLICBpjF+CMlZfdzhZCONKDA6sxxTgxNzElHYJHuQkXAqH1xHPbipqe1iNBX
D44aTkMPPDDNFqLw5w3KkMbUGfqGL4/YKb6OhgIVj3NBxwxGNitW5kPj0jxtL+ef
01FXKDkvho6DJ5q2kK0St5MvcO282OKsx9cbHV7qEPx9PaB1lVMa7pmFo6Pg7IMG
ILkq0s7EHo/UteSSZpF5B51rQvrytZMfNovvrhZhQ8UTihS8KgJzopEeXcWcRc1o
KOrJcee5/YJAMXDzipDx7R3tTArw0AzNltLV2qSdImxC3ISKVzglkU3IUJQI6iGC
jjQhDtJCpIFGul8FF3SwUWI8bf9yUbP6LP1CMhqMTdLjfOWVr8i0b0NFIsKoREwm
+dsVBeaUVIdISJ9jLEUfW9N20EBsjBxYmoUr83YSG/sH8GGNYeVHo8YVEFujhtdN
RToBNRUXMcqqTzDVlotlO2THGgDWn+ehR70b878PYKn038vytaxJlZn2uoF3bYfI
1+MzFd1PZ3BtT0jfmvISGXHyffnUfzer/YguKkArp7t7fAomAGNZ3NtpxrvcG7lq
1Ud+A+AOqKDzio0Tfgoi9tgXhwuYrteeQYK9lsUmG//GLVZP799U2P1zEwIfexpY
QHBEU2lS7GdCs9x+w8fxROEvA3I2rC0cV2KiBxTYNi0DM2wCleS7ZFv0yH7Ewk6S
PPmVpbggD0tvUM/YvtV2vo7Y8HD+Hxl2E8rnjN4mx6RolAgqvXRoxl8ejY0oeyaE
E4KPhohPu5Iga/vS3DjePxYl1uZ7SZERW14I/5VzuLRc4uihsDYYnpvh/6W9kUmH
vVpiKBP5/ewOJxrUoDZfj1KZyU+Z83prmPpuVxJorfdPFZaeLucoadU26b5fSLAB
WTLEbS3BbLGwbSUwqpd75Oo8pOwso+fPgTZ6dinWqJLnx/hFJ65m57ta0dO+uha3
CI1fJi9g/X6kX0S/hEA1Fa4URx+IlF9hQg02qhDM85Wh7XaB6imWJ3CZ/1gzQEqo
dZ9vUs3IS4JSOCzRd7/prDo6qqPOnoAJQL0WmO5uUGWhyJEK5zHzQuH+9p+aiXrS
u7f+jffCn6PjRSpGrNMuQ/GBEd8DTwqagij3BZBTeeVhzGsBO8BMUi9m/ro2PPAu
RUI9kI8l55p9OAbUsu5isaSvBLrVHk7xJIdYStCBc1c2/p/6246rKr1PQ4b9vDan
eJAtYIKfxopPMnaQWnTRknkqPLq16cKxD4amjwQu1AyXmJdgdvV6wq/DTORWC9xp
tKScRsABL/XgzxnQ8OfgMY6982lGwgr6WRgW/VQtOg6JeT0/YIhDDfgnnEhd09hn
`protect END_PROTECTED
