`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Id7pYP90QNVQUBk/f0j95PIK5BkwUlEE0SspHYQvfkIWOw29/H3gbxVmTVFulUvC
EQZ07v6ru3sqMuTOzHrPYhnf0LBCwBSzoA0Lq1lo82XsgTdoE4sl+86EBmF1b4Pl
VQkFMDrnDqjGOawIWAI/8lXv4p61kaiGmxJU+Sb8EuxJ23yetGCVp5fN9nvKhQzl
0sV0H0MkQNEtsDf7YqsxJxukq4LW31DS67DhJXamMGWT8qxB+FaL6PSG0dySSJ15
x10Nl1a516lP5gh8YL0g3GnIRtWg+XUnLOejDa6uVklGPxZpXBtZSJoiEA/24MDT
Cp81Z7KdypK2rqGt4KJkH7o7qY62H2RMcPBM0q00SeTyElIplwlxwVSXp9/aZO4b
1uPWhjwunPN2wSrFxCqrxlK7tI0+3U41jf1bdKzh5d+QPFWKsTt4F2gMDnZ+IAFo
ByzOynuxJ+3QithNbaaMMHJHtjt3QsTngiE03mCg/Gfkmf3xXl2YpF/BNHJltP36
jgBV2EJqz5lp0L+SVIQU6QodznqM9r2XhTR0bpXUwkwKIuXSB8YZWgnlWEKIrJSQ
YtBvLp8+mxE8DXXYYlgcjmFylLUCNh+hK1OadP6xXCiuSbHfdXXUOzLpmA0C+FjD
4FZ580vPzPpX5PKQhCgUGUnprUQnW5Wc/NxdguyIl1LZcXQ7RGKCYaTtrkY81ZfR
HvavYq7hxsps/GAjKvvPUrWMzDiyJs5juChjAEm7tkJ2WcDh7QkEtdobwv1zD418
xVsXwZJP4qYTdX2xzivSBoQ9HGE1uuQo6G0++KRGldKu3rYHYM6XcLi/H6nO9DEj
rsMa2cdXdXirXX5IzsnrC67lBJqceR9Sci0u8RVkwzVV0WuITqQUC6ACmXbGO4K5
JlkZrbX2faV1pLLKZSx3nU4l/m7+sPfChcucIhQV1jzRPA36oF1NL64OLGGIRFCv
59tlXV7UWNyQBdk8YuScn5ruFQo6THbc8z5R1SpmmOK4Tkl/okStyVIbWcb9Xyy4
NTXmdezdvx9n4kbCh2HxMukj+bEYSsYwXK7Wp4DzIzYVrTzexsArJuUTsxaHwMTf
Smp96eoT53sh6jvXCUI98os40/E9NAzUl4SsP4hbT3PmTjJ7gwDZksLLjlcKPt6J
Idf06Cv+8LmereoHn3P81jcvLWOg7BOMd7LzJFIwz7/8eS0Xy5+E5vIJa6oWk5A0
LTemzSJfJaTsB7GtbeXTp0joSstoQuR7qknn0nVTwJg8iniFYYgVaoJZ93neYbuD
msi2Gmi+bPrLMg1OHu/wI4rLJUcuY4C+rtQeVaYGPwjdtx4m0QLT833pBg1RH9Kt
qvst4fySLIFWgYHwpmSLPXSWZWkZ84aNFQRSCYjt+NFuCvGYu3eBKAQOlry8Nszi
gskFsf8q9oGqAkYyUMPat+X/kK8ujs62q6fxRFwrO5ONoP+InhtQj2+a8K5PHq6w
haJoiFXNfaBI3JXZ27rlIHm1dWs5mulI1wYUI2neiWuVwEtkLGyrjMeZFNdXzVgK
8WJLFlbpPOIsy0yznyJNUv8HmVz3BcfBC13OGVNbrDInnmkLPv3KsWC+rfF9O62D
0+wNRTMSDIRjyi+8xmV1Ya2QyztZL7Hpnn5SaoAGna8=
`protect END_PROTECTED
