`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tfh6w4lXo1+NsObZlNbdc3GVpsQIQpBxe+Ml7MNI1mNR41IMoNnmcDaHNP675Bm5
pxDu98kDXDpGsalZ4DUYHEMnotp1RzoT2X4mB6i3Mm55Sq5oQC99NDyqcd3gtVnY
hUtN00Z8yjAHRqUYOcb+7KBja1pPFR00Ncqs5qbNBS3DrP1JS5x+hpScsv52ffE0
0VgYwvS+PhdM6BVSceQ4FDu4hsBeFZvLNiRwrkjnXJeojeMUzfCLLVIhwLqIVwJb
FRL45fLMScQLu8y1CJ07EfQnvGrtN0JMvogFlFYt/H3jnpW/UcuZBGZLoear9FOp
wOHyh0iellJBUT0MEOjwIESfd/d3Zkq1Tgl7whJ0votzw1E3RcxNl/PQ+Ylz664w
R54n7wGyAdoHOzPag0ZRJhf4hySAedk8xViFvfTfTE1PLC2Un8m3qv75Qhs0Ma2J
XNAXhwvRUrrrQJOCGx9/Ads+VGT7pN1O7V/n1nt8FRK3CrY15B6KK2Kmkkc4yOJ2
OOEZj7Zw+RXd3J9Gaph0S3z548fL0pKvYlzw2Cz2z0RHsNxRq2NM081bw7xeObMK
4M4LmY2EIT5WxmARatzWGqLUuqdOfoueiD6CTyvLZtkM+X/JSe4bpthziNmlmVhu
TRXbTcVKCbTh4QZmso2nt//JVYNUeCu+/ZEViVtTm7vyvNoHcXZ8ts65cUWz8fkt
dvXjAkhGA8VifrFI9RRIavVewb3HBrctJkScqXv7RmlSGPQlZPuYpP0hFSekT5JV
+XKlBAg9Q4Rf1TUJ8vyrIfyc918Wl+uzOApl1e0nVKSMjKbiikPbvbqLJzZt7XAq
V7GDih1truncecXQ6qw9Tu2Lz/4pPy4kXNoimQk+pwZwBC8BqmW88ySdi5kGZbAp
X1lxS+vg1KksXykef42O7NU28jLUklkB41bUPs4JS8UwtacUiaEf6GrBRUkFXjGU
48vicxkZJLO7W+DUnWwvMshh5HivYBh6JNlEHn0nu38fFnU1PmmoQVYxZnIN6sqc
qX190RakJquUbmMmNZvQsSu9bfUEqcxaFGyoCOxFpgSBJhvBnYb38uHs1sMKh9td
ijUYuFt7eBO6o5iJmQvc4KOsn7iol20B5sTnoUnFqzgyRtSEMbwcHibv5xtCNkdb
T22o4rlAhF6+4bErwznPsd/16EwxIxJEJHkpvgv6xHFwleqJF3U8K8Ozy64pBdkR
igmykWh1IqmMJlcwc1UUJz3gyNa2RPkfGVUM6JOuCvMmw8Cgm3bMm+8ISQ8UxmoQ
`protect END_PROTECTED
