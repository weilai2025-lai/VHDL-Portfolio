`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
phAdtwwfIv/P4akA9L0GRdnVzC3YTCCv1OSgZrv5D3ho4kfHSxWO6GLU6bIT449K
5CJpPbLOzaN6VjglrKmbz9Xq3of/s9kzfzdckVtBzAUdtdw7pIKR8q6nWdh0kWG9
ekrOozB+KmY6XveHiOSScALJDdXGR++KwcGtI7rIApOIJP8bBKpQCumscKcQ3Y8p
ScaXz3trabPCfhcoP1jhg8MlpJf8JLWGzcj9ZoAjdjo/ckShQ2AV41T1qS0cOtyt
IdGS88lSE9BKMhgcYz6lcw3Av33vsLceo2CBsoT4W09NAz754BN/xXCRx40SLgco
q5xdTDpAOo4z7GQAO7rP1aH03m79wyIXfR1mnGc2D+AtErc+Uto84EFxHZ9tUfqq
aWK0VvOeNTlNe0k7auddfW4UmJnEK/cwkXqFsL+cahXcEcVmLi19McHmxyJA2vFk
YtyR/pCV/skv9RoqaxxvHRBbKyKaETaAkFRpKW+aaNcSvr9ysAR4g+kCn1utPjmB
0f9PAbeh8FU0aD9kKzCUVg==
`protect END_PROTECTED
