`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
znS6kjBsA/jfiO6v5uG1TaJ7zxOKHXPewu+gvZ5zoZ/dSSgbcAsSqvAj6mb+6/JV
h1Nn1wF9z37V5v22wk2ioVsn7xgjxs/wan3npZ3b33kwpHuJfxNYYF0RQH5STu83
zXoAWijXUgVNAzimTbhbU08bGx8rNhEp9jhS+e9pn2cnBrvP0UvUgQ5/3o6L0sGG
atjwMIo1L2mTMGN2dZeCAMoNdZphX/x3h6zVL+1F0tL6s0+otWtVTWfsmnfwNcQm
P+GRj/YCwU0/xE1IbZKuLw==
`protect END_PROTECTED
