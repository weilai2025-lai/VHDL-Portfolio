`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AIlulRqq+hufHdOgVYubVWcBab0FGyPROLARnVMtEA+gGqja9A+fmzKAm2qm7Za
F8Cqykzho5BH+jIGydfTyDO47emRENKNw6OikKlX+pEww0U9tSlfN7ZRAMSkCyoE
4svarsN8lfUpi7kePmfIRZW2WU3Rt2TIHdlgN4SuiUSxJXReHUi4r1oZVg4zcfzY
0p78pTXJP05l/CQJ8SDkw4iYITG1ZG2yP/5s37LRrKG3BNQf3zEZ3I78VhRtnTyy
prHLwvY1KrBFOpLkpLsVmXoCjTMDg0vGiwmxJexzi99il0nfkb50s7RuyWUciyu6
Ojgq+YDeB4oXO95C4CybOcpsbc8NWzhgnRsS/NncIm0N+ipTezozwUHMZYFBj1EI
SeCuiCv09v4u5mSQ1wzajAnC58nrzjU7x8CBdx0E0+/rTd8F2CbYSggKzQq47lgm
QQc7UmaK4CsAVcXN8JaPqSaQVFD+guvF2FUtxzVf0lQR/Z/rQpv6SK1tL/bT7QKo
+AhshHxJ7i4fsX+X0kgekaQSnNgq9ua4Mx08U4glv9uddNhFftcQcrs8nD0dKEz3
HCG6XRP60NWKLELKqtZj0Bqy3mmZ8TGo3YIUaOAOQFT7yTHIaPFNuhvXNYOEvNmc
`protect END_PROTECTED
