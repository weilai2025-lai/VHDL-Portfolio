`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hq/FPyTkH50BbkajUJE2KG4q1P0r7Wcp6geIg94XeNVCxTmHQvMYiiwHexY+dMx7
Vt+dWjctE4CZAficOM28yQMFZxJZHZeg5yAEITzrbSydLLulHYGuXftTlKHNRx5/
dsZeP9y0BtiVSDYpvlwWUG/6g/xozAwQ40vpu57dBE8G8X8A0ePj+k7ZPmh3zg65
c2zdHaHW/VLpeSUv9NUZc8tF/T+lBQo/NzlUAjgklhX98t86ZzNj4G1is776TYJ3
Z0jX1JRoXS4Hjb/WBr9Zzb3tfYglOof7w7a+IX1VWCtL9Xr2LvTCpy+zIm6v9t/H
oeozUTGDTxkxDx5BENwPoUrDVADL9UQMyc1C4Ljh3HZlrmKwAlmJO3ArVbP8JOtH
6ZwnreXndRfBkSo7kY59f8v3OqA0lrNtQtjKLJZqg97b4fNhEC8FahlK5JTphj6g
ZfIW6e7Kc2zJxxxctt/n6I73aYnAUxWoK0iBV/cjEKms8Hl4Cn7rtOQIWqYM0yPm
EePYt+GCIG58aHa80Sc3hphgZ8ShHZ/Gn96taFtsbkZixIaniAUHfMcS+rzRtIC6
rzvzVXnTBaGqszCFJQZFWTCS/i9sd9PJxdJNSYFtjIZEQN7LNajmDMkPLGwKgjFD
G4FKIZhfzNa7Zg7a7YKE5p/9VNrKlMQOq0tff033pkTUR7gjX6QfUcXMpKulv5Gb
iS33jDrLioP7vrBuHofwt8jVa6a/1G4YzwgIIxoLcMOCqAEleF7YqvjoWW/cj9oS
HUBKmgVvRVIPJ1nP/nrGNjMvon3FHPE/pz1udsVVAoiyctWSThWUtUPCcA7Tc+un
DCmxfEpBeoKaFnNcOLgGfmxeCh4+NomqNQlilvPASMATKa3SSxNtMjox/XEiJ5Bi
vvpX3tM1rNthyerjdvmJwwyD3b/3i9he6pl8ABoc/md28yBEQbaYmlfj3KDDVsth
0OvJipatuRyhVtl2E7NaywrWtAbNr8oFB6yswtS7+qquUzqF6OWU5xZh8SKfyCjW
GhCYL3BB4lUEfw3voKU+IgrtG/7bGae21k+SnWZStkuSoKS/WZgZ6fbsm/QjxROE
Kv/BDMGvPbq62JtoqzCzE1z1UYeMEBNA1LoGJLVuTnSACsqRnU1GwuNbKyVvZUGV
C8+Nid5wPyfpTYgoBGggDfrtPUpRpvjg/LGJC6UoU3JnBxi+E/CcbXolLgrGH1TR
Lsi8lCDZKUPXTCr1CCVTNl1h3oYID+hOkq4of0XXZk1ztc/i/8IvcFJw2Rr6pdmN
ebSnrnYlamD4f77lSKYgiTxyWb82l5d4x4iZITv9+KuJtd7IqMqxvPagbtSFfHYf
UzyiE4lMXMEN2j1tWjylWJEzkWzO0y/BDrq2GMsr2BQR+Js4U36dEUhMAU5hhZLL
maFuOxEL66Y/p1iWaOn2/4LdBl+CG/hGhHMZ/4VtJUixWsO0iCutHguDL6kC94FB
YIiSPUUNvcREM5BvqQm6C0LHW/QAoj86UzQZmlUArVLiHGsPq4GZU8sdtJzqOLJJ
B+Yh7HRqe95S3egCHW2mO7m5zzGh3s5qgmEoH6V0PCcv6+8/9w4u3mmVosf/Py6J
OMo/vYmOMLhPJ4aq2i7s1CqjDN9/Cw7toWraUra8DTkWoJbneBe/RlUO3k45TyTp
Kv6WOR5pPhHz8rECxo7DBl0I1wYjznxMj5fNlM8twm30Q0lBxFHOY+FEcRrvCZio
gTm4VZMTMPgGr37eAZ2DU0BC4yPVYueaDkPLdv8w2BaexmNmOKVWutzZ/GABubTT
YGSK4Xo+gvKk7gTzoy9u7Ps2MzvIC9cie8eorCn+1s67StxH8UyjaWG6Ut8HZ566
MtBEFLNHLD+tj6TGgxyIFdkjT7OAODqxBb7oJO62yDoFvJPSVC8yJzJBR2txnIAt
fMt24E6NxvCQ+VcsjFQrq0juWHyXccsed+tqh3mcjc5v8nZMTS2j72p1uxdvIT2i
4iUwpvaY1aGpVlmSJBrS0ZDkydVJk4EsT7WxTYI9dGg83vIKhnnxKnqCv1X8d0DI
qe2oFBs7cRnIKtvP15j9WydC85z1WqtnOGJO4eOtqsxupDZqs7obICeNYyLGwWfJ
Fy3Gz7BfPk9a7SGSYA2kX8vgoH9owve1TZDFBaAvqTS6R2Ko3HWKGhxSeXs2MLtN
mifaFPPLX5DZbDwT7AIQ2nUGzVz3UBU2SoYh6qykNUMaq3NQI0ZHX0p4WIDz0b19
tg3gijBAkRF+foKC4mYAea9e9hFRlj8LghaMlZUWPPk9CmmhqjW2ecZzhtqwANzB
IBAzHcotvo0wpuzfMaMFy6xEChT0RR9kggMo42fnmh9mqcax4v9xT/lDFbGvaidN
qtipOLQGkhK24tVPQEbCWX3oqoD9xzVB0qBDi8CX7KM1VMvKoIGaITaLjx4OgpUC
Ri0Wi/VYeRLgCgl2YO9orqTu1MG0GtbQ/EU+qYFFUHOOHUubMpi4AdDRtMJ2vcP3
3z1oT2sFyGubXoM9Uc2mDPxvnxIaULVkEeRUGJIRpxxZ85qruTFBk3CKSAtFOwTp
Nj+d6BEEguLM3pjwI4T0QYe82h7ifk3T7Mu74cUwzgH7m7pI0q0GutGJDsNewhFL
oHxGd6bERSPa7Cc+59MZZ20P0xQH7H+q2l34I4ZFGMyUdUOY3SmN22gglwCsVZP8
F+5NlSMNjMUAKIO87RaeOcjeQ6ys2Hkf3EW77x6FwYzF7XQgIgycrg17qYd+V4qn
tLMohvgAfIEId0vcJl8S8vDn5I8wwuFDiXdUETmBziq+1EqSYfM12PdZndf5U3ja
BH1b9LseWLcZI+VX8SVvFU4fHEXiXbFu2/E+0zBwoBIGq3PAaT/CamoIFnGTzXPH
6ud38MLLFYtT8d6vq95K/R6dHjkWfc4Mc2A+uoh+ljHlKBq3+rLZ5Vu0GPfH22jR
C107jmLMITuJPas2jRjzVKelW5ueZZQpDo8AZEVf2eOiHIQJkMFksS672zJ//0YT
S9bVs0gKLOEIuPVp5JX0j5hLoxo34J/mVp6F5XXFjdbY9wVtMYj5Q/kmAg6lfqrh
VsBWjCTY35zEzS3oOiAUlycrGle30PhMHP6KZcw2NOB98Em0dGNf7BBIpMHCGouX
zT30rpGHXWSnuMsX4mauAHgKM2uXmlpSLfJdRt2wegloocBFsdh2wkfP5hzidIBK
g84VmnGGxTTYImlIqc3+Ua/Qj0jodHWPbNTGMCPZS8znfTeqHkhBdUrSxGEZVZwN
JAyRx1e3dBBRf6nQwz/Q2fqntO4libmYmYtpSabDv87cY/yurHXcb+Cf1Lf9LTeb
IUOf8XVrf3xAdCXMHFnSft1HxEzP77WA6ON4cE0u69GDIdBHQg+QQ0x5cJRvSVNn
++cA8qiGv1Devx1drx4OxFFUlOrRnSKk4LcD/K9Ggab+Gw5OnmX1YZxdR5v96k8k
OAPKEU15V4mPwIoYj6rKvFnDl9cZrSvGT/VL+3GMoA8UEaJQOkhTP9wjNPYSgeyD
XXaftlwUZ2+YiwDtoPFXTPs1ivD4e6+v6bzs6uwuY2d3ZUmN8Jc++iLvVGAEabyj
9qvQpM0ORmFpp0/cDdxOxTUvu1iDVEnkuXTP6gCmpfAIzBzwW+hg2m7oFzTL8mcB
Vf/wwQJGRQa2clRVbq//CE9O51Jf2wsirvo7K2asDgoTmYg9p1El09dx8ErBq0yp
q4yKqtJhXZjF5Bct0NwG4rDHTzJq0VUvr7fi4BfQpRNgjIDcUJ8sBVfbOqA3HjQy
g44AjI4amOTiksUn/WAn7S93+VR5GSctC3rW2B9ySw+okz11lEvmS/i9MZOr9t6B
tRfPAXO4GkFhUHgnp3d+3PcpGCPubpFnkazSViTml26wuhxq2c7B583TN5rT2Zr3
x0QdzP1n7DEkPCEGxTxYVi7Hw09HFNSAF2+Gt7p7uNzmoEE1WBpqKlVPmxVQmFXq
8UTlIFl2H2oECZgftgtgFgngBtmfmgz0Pw3y4UL2SF6egjFONKJi8ElEffaUxYgb
P0NHCxrD+C5FBxi/7RTaiNvtslHm8wz/F+Bbmo7TamRrB37xRUgmSbMaXMnI1JPi
sdAZpn6bg3wPywjo7QGEaGfvYdadM5eSfd3kaB3f04QAPTtTUnxfLTDp+/3UI6tk
oJeIRfMHOL6GNZf99Z3SchiraotCoC+KQN4aQA7+KMQT7VDC0RhyZhdbq9vHPGG5
9sPoutm9dmOqBmY5RTaxEyCBbi5nXFmJpeek+SKj2AXaetoFDY6U25fe1Tgbbbz4
AEW3HSRUSH2wS2ZobGxPXtaCEeiXRR1qyckyw6/SuxSUJ+6Z6luWzxEehVd5wLo7
RIsSijClO86bPPp40Esa6J6dXagSWlY4sqSd+QMljf7eXybIv/XVXVkHcSnKFtiD
r30C1VcATMHW68dvlwzMtx0wGQpuqu06yi65ESfM6vdD8QWXJrFSAapT6tloa97J
KB2iLe+LGKVq88yBgX59Tct4J5WDqiiBRg2tNE+TVBUEJlceTck2RsSoDS2FC4IV
K9JXdvo7XabrIhQzrIv9GNievuGC8rcg0bbFqOd3xojlOtt6xlS4o0EiyWkzcgRE
M9X1hL0qiCDYWdOrd9OFwvli5DzFXd9XFFm6opITixc6R8crAsPu4V2o0odGf8gR
HCPliYODLuE++J4yN89H9kZWPFSgbobrluWMAGn/u7pJr4vPGHrHkDDzuzGfQMqf
6kRsvoobvURsx5SlkQcRuUBvepuWCicpCY+W2wHlgrNPS2RjhcYOYr+ubYSrVMlr
rwcFy39/dRMI2PoC6kQ2KfOrBRzkjQwHJeolIfmsuORUcY81lP7tKqaXPA0/6un8
dkCosgNk3GmSkwZYfywkKAyYKkvuFn4QOIAC6B+NC0zgxGkMl3hAkWbCbP7b+3dJ
8C56aGmPG3j3hzt7OSheGF9cc90K4QgBhHxAsYVs3w4R9vTzrKAawUxIOQq2Hxw4
zfJ8LxLKeqoEtobhobu3Y6ssYk6fZd1+2I7AIlfMbsIv8GXsb2sglpWQ3OgbWNZD
6fp6dziDfN0+hi+Ba+K3oLFlhU7Hs1L5YgaY3sTapwFuooxejzwo7dPk6cpbeTDW
KANNDqohKMTFAgdSt5TFQ6BRE0s+sNA8zlbmYBZGomOzzeurGR4cHr9ZAn3HN56Z
d/B3BzaiwiYFJ28BHEzoVck4gj5dDM/QoW854LVyZ24XkxIylUMtZpX17VcoeQGc
sGxQFg8fEH39nXYzuGV5yJkguw3uV4SdDBeYgyyUuTDb795cVImbqEeEsqRoKTDY
A41/Cz1lUocR6eWNgY3o9oQXBuB3EABp0S8U8Vkyc6AYDKjvKXxWlGrs++UnvJRi
wpntHBmg0ZJ5BEHjzjGZEx2fk69iU6tsHr/7nb/+fVp27je29rL5IjzYJeGjYyyW
LX2+4tZzrz/sAQOWnUPbEhLCTLngog7+O0BaPKzemPOmStHpSP887lrxU/27TjPT
Ney+PPY5EeB7r3V4qd1GPmTluqdGxLYpmLd7IKQixn4=
`protect END_PROTECTED
