`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
akixqfSWgEuKuAtjm3tPFox3Uw+7aPzM8tmSXtSBH4qdygOKdJ5585qiZkgB8c+m
ZzHV7KSWN+T1zEsJyjLIHyH091fxa6zQL+N9I4wAJ2CU4kym7EbWtzgwqYS68Q+x
WOW/3NQRbMvPqWM/ffoZGSbleFzu4cen2qUAHj30U9EaAJjpoU/XWez815RTSj48
l0bhUcolFcdWdoDTaRXaimJ0lrWXE4mpG0KrqOE/TOz6Co82XZn41dEze2qXF4Lb
YkwZ04A1x2Le6b42TcbkGUWiiHHv/S/qCnP8DFaDZ7utFr3+LyDd4c8aBDB9ptFF
Ekg9rBDHV8fIq3wa/k+7hCxOhllm2shrGShXUCP32/A4lbqDS96n04ebSAqvZeCN
rdtCoKDauGm23MmwAX104P0RP4Z+cxuwt6cieVlFkUcJVJuUlchsByv7NBPcHnJ+
tI9+bZJoiuVHi9x/AWA8YiAg+2BxFukTZJ+5DsNb3DsWX+2MLeu9D7A7fj9jyW3D
5RyP3+hCph4k2jFfY4IQ3vOgL45IhKiPqwgAp5g1N2zhwBWG3H9EbEIRYFI59kgv
2zX1VX9Of+pjz5TNa2QN3VqWnrGwpxwHLrB6awaG930xrew5Qsfbv71eXB74Sktc
VHX2AvQN1Uj0H805d+lANJtrWlYgqBtTsZsGJX3IiOm4Ae4wzFUP4PbD9gd5CnpW
lXwrykrnBeM6Arg2tf3dS8gVHKfRUVYnDl9Tt0jJZigT9zYuQc0QTrLbSRQV2URe
7gMxDhPFTAGfT65mVyIRzcrr67p64bCRddh6MsS2m8GkUjN6oNUfi3qxifFcPT1L
TVOfAaidz/WMi8kK9AUGtnZgOXwjjihv2Wp65hvthBQ=
`protect END_PROTECTED
