`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXeI36jAV6RP8VYl7GCf9Flm/opjryf8fB9o0f8trKmxk8uZMsWB0bFH7lNbIVh9
CBCkedeLMCoUQIw6+UdE9FihIT8uorBUA1POUudJRToFW+Pl4nkK+Dm/Dj413T2w
3kxAbM50SBexnQ7KMwIXYcJ9fRGzTmjpVZOEji50UapuJCcD7IB+S9D5vjK3Fw03
2xswSaxkDh7js3Eh9aJ4m7aj67fYSINQC3ICFzmqw6q9giClyPq6Ym22oCLYBSBF
sRkmZ85saQ1udEMa/9jNadPPVOj49yDgIl3E5yhZgJ7RVVBiFGk/wFj7Q6K5v+O5
47ua+fZ+rk6QX8+twdhPKL/TYbM+1tBxRU3tOCo3Av5BJ395bfC8Dw/rgcphmsbs
`protect END_PROTECTED
