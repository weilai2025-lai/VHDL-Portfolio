`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hW97oTyANgPa3/vumvIFDo4h//fQ8FMa6WpPKR0MN+0FoxllJeW79P49UAh6u90o
FiVk0qkg5m4SiwUK28BiOvqzvE0I1meIOw8QowknW01C84sefpxVM7Z+lqVXuYqw
jKOAA4ngtRe5va8kHzXce6HToVqIoFfkJu/QBKDtN9PgsZVxbkoaGv6acWFPswUE
JtKN6EFQjbeF4wtr7QcQJJC6pBSGFJ09zQVx3hpZHfWmlLmXHUTtNjBGpWsU4xTO
xqcD8s5n+mh9PG2XKk93XvU+w0MTsmjSMQrN5q8wBKCAoSGCiC6x1gNeFZNxhE55
YQGxDeUfg3nwPPWqRg+SG3BNy3ayhI/kKC1MThW3099tda5BX0nTZhx2FjKSZRRa
DN4HFMULJHScb9l/yOMbUGwMjdgK32Mamz3+UnNyMmm5mUsPC+ULWG/D36XMJCcZ
xmPbcqjEjlW5ghSqHUh73d1u5ERkWyQ3cJO/5ToO4tKgojJRk1YUG8QB8dOJoEHM
jGsFMyy/oMhfWwpxazWwUlAJ1EXb6CTruIMOPMFiHkgiPtCE7xqwkIpGj0Stx5rd
tYja3XqeCoqGtYY9VW0TSAzjMr+cqUdWtscirU4FTs8aps3keMlWcNgPY0thv9sL
WhxrnBB2afJ86uq43yNUD/wC/4IeuteOLYyHYm8lbeTyGikR3Zb2zRoLfzaWhiE8
R3sNCs1HNjCWN1khVCbA9CH0GuwbvV5/xhzVVve1qaPsmj/cd5PZvtZWBrSU40hq
QVgGijJsOGeY928OtIFs5Rq5Dk2vjdJWDQ+CG90JIyPEyBtKntzVIMr2cKIzNN52
Tj640HtTR0sdOnYg+oWq9F2Y7FFE5EFYw+RyhH4T0vSaReESJqFZ7jRi8QPkn7jD
fOuMQivxOc9gAWudw76eUNUEzLP/tqWnMexFYELR61TT0443QoXDi3S4QQSa9Mfp
vcKDzwFal6EfsK8COfjEkfCyNgoRiClabfmp6YRk7YlxxatZFoT3gWBNLSjiFIar
SLBnz8uXzb8E2DL4l7OH88ITEa0wn3Rr6BPvK80Ahiwc3Hf3mwp9Lhs0vm8t6hYF
BVh4p7m5DCTxmmCVe4V5SMX6bV6dhho6/O230y8EXSCdE/DD5YUdG3gtK0bfnJTk
YYzxe+Lxn9yLjSdYjeuoI8BMuB1berDi9+y2yVTwwvQFtpX0q5QeVe+PytXCl5tn
GP9l5hM9+55pvmC+QW/XXD1+9QFMYZEgbyt373wQEUTzctM/SeTaPN0zSpqHzR+V
2VM/3TULtYwWeN6E5UIH2l9GRWvhH5WVmkXgDBnq71aLcUFhN0Vc35wXGFh6Zur2
p6oYXoqSoZU4Qecmt6WG4+J8J9xoTdNXd/w5tskGxcqbxTp0aigtNKhDuJTe8dji
8CLoKF+k/VRgmdWm79QHtXsWN+3zqfQ8oW3dXWJco+y+nJB2IdAJAbSWj3rd+AD7
scvPVHu0beYuiOms/5CeP9ca3nZhcNaqkkbGdJvGsP6fUDilu7ENWIQhXn9j2wHh
BXO7usAXGzfZij+8oYpPAsqesE/FIH/jZFfP5l+24AALWmvh1HUMeK8QtGW7Jsjg
MFS06Jau1Ysnsr/xsich+NQ5CneUdDfqXySOlx5apheLbiFPqkH3jSxYW8crLbvE
GYiR+oZnSFbmxZqCfY/8FIg9bKky+tHjAxhe5Y+yXnwNd8/5q5aZwjj/e5fdImK+
t7eLTf34kOX7uEo8jtiUfj9jGDjspXzOVq/bxqujlpX0F7EaXEhlDgh6tvqwzVYb
sbewi7kz4E7DguEjftW/kzn6KJ0p3Ygz/cZ/PwOUyYsvftJ3HyjiSDaH0Iof2IBp
koalRnjrZWrlcpXEZOWXKWG5bfUg0eeaud6F5e2GKiSmati+nIm3mtfAkTI36NNI
2Thip0Rjpt+zRRZnu0jAgWesArrHtcy8u7hyFIUVWDrFkYXDAyx89SS2C6BiG0Ix
dNbKqMrN0WDCAaUHR5gIsvWhrwmkFr3ximIppo82PqAGwyxDkbCwryyxY7XMqO1B
w1VxEGGdE/OkzE6eXzGckiRdnmyLEXEBKJVJEyWGneu7NY0mKFiNZwYVjYESy58L
ae4w1ksiZ9eypA741/3KE3VfT6qId8QgZekwq2PDj3AKO1RXcoEnUv59So3Ap62f
txoo3dRK68i4g3yd/n8XdhxP4xolAHpqoZClrOP9f60AuZWSshTfiOx6pfzNHCCr
Bxv6n1ZNugnbCFrfh7J1MqQiA1aHkbX5OlKrI1g1tR3TuhEmmY7TG5HhD9qTwuR0
4pCfLgI2DUSbUWIKEvTdAy4hayFJfd0+5caajMD2vaZCqVBAC13urwKPzQ1R6cis
5YrubbG+SjISgw2Eukf2kxQXEK65La72WoyGej5j89vFAT0H13swU1ERYow6F8ds
ga8AjSyvL8jUadbrM/H1AaicQHfMbQnEeeR0VaYuBCcgMbnlG5gSFk6Aj5k7QAiV
W8ncTEZ4dfsEL2rfHmGyE5IPGJNe9Sj6TbZ9WF6+75ZZ5sbzs34eQr5Oj6gEkSoM
pjpFpEjIK6isTns2E8t5kKXJnoYz0enPVCkS1biMR4A3J5R3zby3rJKkdXvMupxW
j0fTXHPWdy6DO6H2FXle3Sc9iMB5WoT0t7CUcXBfTvAsjX1jra2Pi595I9XSQAho
B02sckSNynU9tng1Q+v/30Rt/S3feynnpIFgN/rtgB7rgsfCLIZxEtpBg8zRO32U
Xy45YfrOpZTRbmeOdp0i41A47AHG6u2gwcwfE+c5QoC6Fj7gfATHJVX+x/V9x4hy
fuNk1Rbx21ygkUs9VspyBwIQCmHrvlnRlDsdnveierpa21SJn/zAbnBGzIW7+aun
5IjCRDgPxSLKsqEYlQfAR1DiyHZjiEATUQohp80c16L8tms7eutyoFLSF3Is8SYt
vSnfwX/COK5I73lc7sYJK+ggNgBeviMGA/58Oqh00jsVAW4EsLD2PpTMW2i9EdLq
hBWTa1y+bZgB2uYndI1rhvHWCKOm8Nvm6jauQVymtdq7tO8rQpaZjkDCpkek9hzs
UKXGz7GhG77rpPos9fouaFfp/+kdTLMF/f+uxNS2UOnwf13U2D/AAE+NlEPrhSVC
dL6xxPEOZTVO9RJNx65hM6kV16ny+JYK/XtekctTuhKMGTEcetVwFGHibQjFXT79
+ee+U1/J98D0nuzIzmcYt6hc3F4DTXpdyyb17Y+l7rGs+e3AlINwofp/g0PfokR3
J78VkH3obyizjm3qaUtBqgFn/frzR5aHROasGSDfTpNU/XHS2dyI0oWoPf4IDXdy
a1SNyRS/D46pPz/TMOpOXQQKL9MInLa6QGz2KBtx4wa5C8CbA9veL5nkiHdYwIKb
9MxUHfnUQ/JUrTKbeWe0G2tnEXwweLfDL8djri8KV9JyKn/FfNrIro2/aOoSQUYv
RfOYSq3ptuKty7c/W8+Lp6xLp6o5WZk2KSS9wS7TPxeUQI124GS4MBaUwADPE0ZZ
XzWybqDZylMMYcizgUgbOh1+WDXLauJnKSB0wG8weVblnZ3b6/Cw19acT6oY6ybK
1LLDqt/rlC5Jbet0Mx3i4H1Ta/1czBPS3BEQqPQZGsPvkaOAci0AF8r8Unyn0jQG
89x7xKG4oboZbiQRuLXcM7YIY4m6OoKsZU8TbZ9bRBGsoV7lGHYkVcnWCTbvhOrb
sC0Noc30m6lnBFvAmBKaUIpoq1kzDZw6BNaVBxPPnW+40FjGV3BQ8f5XnJFo2Vpa
ronPfz9ZG//FBIcW4mJtQeOYkg4iPKlu2dFsN5N6njerG5GjRoNC/0Vd0Xa99eLq
sd+8sbQ7zs8/y8VB7qic6Rs7L5BRkyeZpu6wWvLz+sD5XKA0xxT4svEi8CXqJsQE
qsYyjLpqGfVXs1TbKwhrKw57uH74VF/YWlSJ+YSIl4BHEWZx0MyeLoolUUQF4MOS
KpJm0RIOBhsFXqWMbOBqvLm/mTWG4Qt1igvTLD1grPs6Z8ecGRkVA1amEPOkZDDu
O0OYKpZkWIOjFbTnt9ipbcmhs+Jguz+7/YgoMteLYNMh6u7Yiq8u7Wp3q0XbBVRH
y2B1lloQjeeFvY9Zd/6GEY1DUHfCvCwdHpLKWiYN9LVSYJjYd9f9/LEub1wUR8nO
TJT71gDKAdxDZvj84ZfKAJvjmfxOBxkpcwSCkKW/x2MrMicjOeYfYNVeXAGr9/5P
mOt9/tQU3kHFmrLm4+isqZB0vXfJB0B7FZscZLStVDiAUE0jC44QUwZVT2tm1n4o
AdzwFq2RaI/uVEsvQx4Kq045dlGVU9mfk8Bd2zpjwChjn9dnFKQ58L67zoJ9WDAl
b+CwucN+A6ZnaPHlbJuxvSeFRDUCdWcIzJKNrLJiB1AgqG72NOtZGxz4kpl29bmL
RBLAhxlfvbl6VfxywEZruYp6bcjXAszGh31GtG46H8zhQMpqpPu43GfGEO20qZa3
50xKz+wx9qt40Jdv6qPawnjDR9WoYIg4ec7hSifWz0FZJlW3wtGmkX6WitENmfBp
/A+JH1RsHJQRRtpBYVSDJhSIm8ehjxWkIesMMZ8rLTVPBcRpA2hpiEpOlyYb6gxW
sGM9cM8SQiEG2MDHVpR7j3/BEHyqShxhs2v6N9zN5s20ClGVecYg0ArItJhfO4Ed
y/DYVslzSiKJ1Sfu8DK82b8Lz0XNHokztcSXeRqI/vmAvGh6iZkdOnwzlNYlx32h
Ucf/gqSCSP0Dcwg6ZSOcXDfIpzPBOVyS5ekSsZof8SId/D6TX+jsp1T1kaIoyiSX
nfdRXco0LR91BHUOwaqyI+RUWNEgTOcXMf8iMKwZBb2O9lIWNtt1Xy7arNVBC5q+
OW5f46/95kqk5EJxZwi2L6JG962H82tQlzgzaq31xmq6kDGzz9eWUrv91Z71sG5J
HnBLY6wlrczks66rOThpgCw0CVAb9pkBwPhC9t0Z3Hrr1Jk3wcv93p0D76hKgLKh
kj4AHqSABeUsaSq0UkYZu+hOZEdQnCT2zhQZU2WAtuFCB7FLGY5rCMb1sLAP58QE
13SEeSAEP4JLbzj2Hx6j5/xmY1UQW0TDLUxf22PMuujv2EpasW/GLwHN6IAf+wqI
oVQaWxzMVGAvMuhVTPbQ/IubiErXLZj5AtHV1vhG0F0yfB4f8f9IVVxoUoy8HAx2
gxioTx1vL6gS7G+JTH7qR4y2C+NaF6aEjwHSqULJlVzAcS5I8DNoDwBfLHxOVCOq
LfcJBP6FPHG8MTFv+mOdbMmeVWODl+rOPJ0weI7slYFTjRatjOBTjE6apA4fIf9B
rs/gT72GY99+fDvcZaPzl2iV3nYSuGwQwP9BlA02Py2TqH1Ka3gJogfHhGGeZHVN
gvyiDRX18987+rlS85tmqnXz2x8aTJeJZWNgyrFyiYXw62b/OA9wtWzFv8k50Au4
XsYR+ZHKrAx6EF1PVpPYWo23Md3SEhbEEKZLqN9YTkj6cbIWf1fSAOFwJl8UPs8u
0zhMJk63GrWupQvRje8pC6cCNFFHkOOeV8sz9wLAU3Yp4bWJ0piAHXaIWv5NdgsE
PHS5vaOzwJ8b/2ZMG/jnAKVPsQB1PTOML3JxxdlobifmZWoGD7/1mQ+EDk42/jET
sjVgo2uZqeaggomhWIoDRR+NfrAarQyT8rnVA1ETVw11WtKsfRVPAj66PVJRV5v/
GH5hyG2oAI3I7X4ze43rF3KlK4UY1+8PhjWYq8S/q7GASUb+Hj8qdvGMC5lje6f7
xKzMj+LouVVGbSZQH/7p+ZTVYG15eY/Hp3Snd6X1c6GP+gLjdRGEZMK/SVawUhmj
bOaqxpMtZuNEZeZHM96Zhq4MNcveAriZYmidZJyeZBe5qeKXj5cC6nTk41ctwrP9
aKm29oSS7kSqm14SAVa0X8g21351QV7wUhPHE2/gireqEeX7T3+qsBQzCTfXwJZ7
NgDgKlMqn324rCwnHFx/TLhAW80ChRG+9ELur6Sv/qUCXfK5geWHH//vXW876Lks
3ZlQNOgX3IbbweL2w2WAL4yHuoVw17DIJYiRcXPgiA8vmsBs/axmk+hNq2R7ATKk
B6Apji5/lFHKDzc1OuqCe2pj7ho2m7MEM5K9nCACVliGPnmZpPALTn2gBou8kxeB
3kJNAunqxcku7yRZCvayHLIH9JYNld+Rr3o6q7VrPZPuXtXm7rXHttEYEyzqTNGY
A2F+PxaVhqgWG60w08pltC7boYuJK9vZ40et8CP0IsFL9zG3k+c57VB4DYGydQNp
5vAAKRxWN+TKwzjhEzoCHSW7zAN4IxiZHG7IDYPTEh4LyVs/NVuFqfcPTd45IyQJ
tItkGlySAYyvpAm0amCqRw0RNOgp9Q8o8yNBmhyz2MHHj782Z7P6w5j8HLFp1SAN
aORIJHpEVlcfod0Qod9EXZ3QNxUKQVze0u/jitScg83VWiVGRDpu1VuLi8PDpufo
e1BIST6f30FWsSp3nPrriJFecVjfzDgNr/Mb4rY2ZTXiqLs6jHSZZuY1xNq+S6Ai
CSgUa7a4oDM8l49qt5qi2VpyZYCVIv/mOLQL6rjpGpZUZgHccGAkP5XNlDIffbcl
fmLs6G2gg2dm5mUJn0M1kOf2zGFf4DMWZMFO7YWI7YolPn/WQStUZAhbofgLEpu8
SI9+/Am+eVeST4XwKy7CtExL89KgxMyImyIWKqx36PtFOft2fLhpt356z+txw+f1
qkHZKDslaNcaEBQo/18t6JnhJsPSHaIs6uzo36jfYQ3W3nJeX/y6LIOqqkkJaOoY
pbGQkIXRiZBucWbm6uMcS87ev/IUqYbVI93GyuWYlrsK+IhkDD+3R+DIDto9bL8u
x0qg/rVqHZHPQ76wnV8XYesilPVrkv8Fa9k+7CHhHWFjfwpZNKe530NCfJzvrm+8
iOuvJX4QknZeuoQJRNc10sOzq588Xh3QEctYB0FTCro7Rfh+JeSlGeR3L+2BNSsr
p9ehokFF0vFhOS/9r2v91Q4cHmtN/ETUEcAfBgOcVlMDUTIkJTewkWjU4YC8ojEM
er0V2CNfME8ue8k7jZWVOIl3tIDTVzunUFMe1Y6ev4gJpdPVqYQnvM+3j8qstHxA
tIiE8aEn9FA8eisZSU785HFbV64GA5MNNclG7NdoKDdmHUI5I6rI6IcA2beKPNyL
f4Afo2ivLSUBYLfnbEa64mJBll5rEZWlxwe+5m+AHZJWEts/yRDiKagUtexcOruF
gGj/HCZw9ZUSO+KYji3wUGQPRKbCRbCh4D/WkNc61Ogc0BljbCSSPEL5H3UIEZ9W
IohnH3E+2tcxVrP26kIXTnEVykNhSHwz0cMxfLzyTskkbv0s70SDCfD7g1ysh88D
jdyoRSW9eBbVZ4JiTNlj0NG8vmjAALG+somnPIrOk8eiqq02hqoJQRNBe7NM8M8f
AoPMkXQaOpQlCV/UzLxqSWtAIaS9/6i3wclmIaAIeG7a9zxMW4T2ZGCK1dtPBuib
XM7cJftA5LW3qxuvY9tsCOSAOOJQefAXOEFKOE4gl8zEBVI7AB3RkpB27TjvjFnm
4BzAYpECgJYGiGn9fivG1XN79EeB/c/AIzG1N0IRlQQ2SVdX0sLSj2jEr6+43upJ
Onrg3MMGPQnvJYjJ42Q4WZ4lUnRPF7L7YgdGTjkyhpiF79MEizCbveavTQSHQrQV
BNaG0amPQDKEny6yP7ioUAhLQU2nPg8oTuLQwf4O2rDnS37AVGQoobps2Gg8QGaM
H9+6sIGKYIVa5WIKRRAOQ/uYU5WY1GQ0l4te3MlQNApLXjVImcTQxTR8lkxevArV
fyAXXpQupEDOGVl3PEQ55CCrRshh9qad9Okov0drA1a8GZRiCMQ2AcCjj9RCyqnZ
c6dPKJRKR2xmcf42mcyyh6QI4MSzETtvT0D4DKBMjVMt2KqqryliaxuzJ186O0CO
rK2t5aBc8+CGprQdPxfgdMuEZdqRQANx7oDPDZcqM2IIvfnNG+XDn5Qo7gnqnB7C
Z8EY7HkIa3pH0hWs8O7yqDNVwACYJt1P2lL+VzxdYaVaRugCG4a0FHHx+dUuVK1W
S5MJt/8W/H/iSiLa30gMxnLw68XAFL5zCLQJRAGzrCCqy9imnFAKibAGIfnEoi5N
Ek/XUzBTPo5+R1PNhZ+4ZuG0pOBUe6foCEgoh/Ly4+SIp8D5R9ZFhxlSVXrXDAnF
wZiModaHDd2KhPGWVHSAqHkfvUkR6xEmy24gAFrqEAXOAvDqWF8qHzTJAkxryjbB
TpZ/aGxrcaPRMEnWkWXVmlPe+1PBdcc8YIaxgaPZQB9tkAIt+SJkxfV2sscwiZJE
anlVsz/8fPbt+gf9TnKCuDH7e6h6WP2gD2pq/caFpXY/eCEhaRyAim5Pi5Bs1Ad8
Rgb+y5Nqkpf4N6fUEgMWkhIe9T2WcHipR5MI/iDfSSDERgsggKuYuL37BcyGi+Ef
XltodT5RPlU0vV4D7M+MA3abSKrLNduZfqaablR598TY6RHblf6GkRBc4SSN9gnd
nl9Y4GcRo2RWPJJzyRtLAWv5clLMVAraQYDY26iEy+FbXWYryVeLuKkTcNUtxF28
9fs8EnE7qWqy8TwwcM5q3qfmK0VeCg2oogG14Gl+Ma/AysYhKmqC/68XXFpZJgX8
pg5NtzisTb2E8FxWaQXaBaPOesf/iNz7cUBumJ+YGkf0WqeibTQiLikKBeZIeJNe
oPbhCuXxOBL2bm7cuR74WbtEzYyUitt7bqPVlkQRA7/BVhpUMRk9NJWgh1p3kEF4
CjGMmYFaCaB3u6r4wrm4sb+MSRVGYofzswNfP464i+sFg1btg9GJtlywKbRrz8aI
CBBiL9d9IAABZ+gEN+biz6LgMZlSQsJ2HC0lvgVxoPWL3KLa3Xs6YWmCqDbyugol
sBJlzvesV9fxRo5qtwJYU8I8r3UeRFL2X+gnmkqz5evJwsuABJW7ZPVcwJmUw6qU
hy8Q6eFhJy3x/yPc7gqEBjZBCITeyVW76RCBVAzLwPLLW8+/smTXBJ9YOZKqd3EL
qYTdT6QMWwc6GcLRUNFU9UTPpjjyssrbHpZQSdtAOiCMsSsH+Y4ALM9qxjjBMevF
9KyIjbfUvgsqH+fUef3hKW7Kzr9WF5uZcKOnt2vxOGSGs9Sg3aePk6kVWi1V88vs
uLvga6KwVfMsLFsrKLx1q7vkuKL0Hu/YnveGmz4nThheBf251qiRP7On0Qf2m5vE
HuuVIjLM3y9VNlUUsgwvm3o9jgxVdjg0NjR7OSidGPThVJAun8LUneymH0Wq4/Ew
Jc/cZKES9FvIatRPCALyigPb+wizAo6aWbG3XW2HJWd8qXubWAVlT7g4dn4dYyxt
7AMbPtqMZj3wbPlkJxUPH5GomvbNNbB/YM3k5RG7O6qqUCsLxAMzb5kzn3tr8o9i
Ts68F1L9uOtvFzYtwI0+4Rt2RzwX0/b1Lzl/gjzaDvPy/4VuhF85ctztP6nQZmer
ezWxNfPWOjVRdpwdHtEEMiZ4nkQbcjJvuACCNKNf70P4RD84U5J9AlYWB8FUTwkj
NpykMCcBHryFYlOkEzhqjVAz5VaRg6htyXKw37wNGrG13XNxlB/3SULD7mopMnIm
hibrVObnsVwBR+UEYJktJOq6YOEGwehyYSEbwr4sR1G7/9RmEHxNCNx8509XvbtR
LLGCscCEJRUuFoYvHq04Z1eCENHweS9UEKUIHKa5MU3ct6LslKS5cjRZ/ZCu8ezc
OcPB8gTRsMXzToa3uQ+HVhxf/3lBEOxU8pEjfPjSTw4RpUoJ8s3/tHQeCOeKJTtX
BbtWOBsJFtGMQacoqkyiOlf1FHxpRNlERF6353raxRDf9CDub4HfajGD639yfpga
0yu/m3WS8g+xNZLHEANwHmBilif/jFhWIWa9ooo6KMBwNGS0Fh0+Z5400mJQVJGO
Lq05mwOO9m7pvllTIlXj1nLppovHyWW7ssIffzlosfyOYYk8UGtYIpYgZHqO+wcK
qsadVZxNZ2re64Q0wJs+xcV/2Ij2WC1kfBtzCN6eLJVVgiECGmujXbOa1Jf+1W3a
/+7lyf6R9FqvtFycX05RVZaeSYEsc2ySqC3XZGzoGtju/2mnR9XK19KYMM6VkPeY
CcpsOKSENK5Nkl93jwV1LsOKuh6NgIpyGcmRDt5EB/3w252kxMJeBSmEa/n7FtLC
qmFdKg9JDpkPWY29aiaR4LK+F3sdkI80l85uBGigK9gOT7zVzqF53V5CeOt3Z0b4
phleiaFaRWkPFDNiquL8UKpRCmqzvBn0FmJNfyr2xqSQCyAI6LwQVz/VTAPhXnLX
sxz51v963x9+8+ttriYL7K8KSBPfqZ9HpalgJU5PJJx/51ogu50CAD9sDX4oZo8N
DyfJW/Ll6s+htbPma+y+5Cmqn5LkncDvqqWBJUXAJXt2YACfRXt4s/wafMxuzgve
Zhy3qbnKuVrvvm3g7mH/4W/z+qXVAULZHf6XayKhGuhXs1IPRnrPWFtSaEP+Y4cn
yrTsbs5LIrwYk66rKOkJsBXS81v1eFDENf6hN+tyIDggqzMKH5HBOvvc/4LZXdg/
vyBIwXHM+Ip5zReazUsYE32rLTq0YCLky6dRMYGQTEzSDt0IsbhJRWR6N7oupvrZ
bM51e8sUan9HP6SXR+ptbeWp7UZR2jjHbFj5lMLc0GyacCjM6lTHdf9ZQR9WEi4i
HJxOYLJvPXnkmzFoE6AHqOLc2O4IV5Pu5XztAY5cY4NJ5i5ZqMoCeBpk167wypXA
XCPm2IX7PCIy7Erly0nsR1OMU4CF7otYlBPjt/LfwH5tiOfsYHJm1AHNT637lxQ1
TUNMyHtek6dPZHXMOHdPjHgcDXNTv2n9XJYUna8a8ipBeGp73+Wx+BZoffBEZ2sJ
goDw4fKuHQPyw5AJw8tRnphBmZW4ruN5TrxNDLqXS4FtzgkziLesHoK5sZp4dnJD
JjzfzWnYGzlBjcbVlu8fPIOr5Od3Bv0A/fwTHYIS3h9gOs/vtM2mLiw97NfcOJH7
s/Lr3nBH1Vw4eSigSfgAOdxYdRcw0BeB9QFOcu3p9sKzqOd77GlyNQFu37wU6nKV
pnrFJRCBE6IhupFxEvhb54dDpNnMtviD7kxlWR35OBpddP1IuubtqJd2Ko2836yk
bTytMvyCuwDoR6hzmKAkS8drxFV6mkWdiI9CL6fl8p9s9lwg7svbEOicdmBcScCi
TPB4fnDUmvIvD+NdDseyGYMSHSI4lVL/Vt0UJze8gSbolL1fnZt/qWSHWLrs6TES
Sw0x540b2DeK14AQN8Azk94E6ysqNE4BR7XQzOLjPNMg+IFBRTibxggQLmqp8FXf
Ko4oVuM3b26TWoi2Uv3MvNVFsZuxl9Z6tgzD5MHicY1XzoIINrCbbwGJGgxgLLHa
pPooEIQ0Oto5r9Z/eOZBC0jcmq5xKb9N3jisrJf/KqmzA1HHee2P8MHRC2fLdBmh
v3zwvOjDu4XIGxhOolW9ZWYIBU7UZBukmzv1cw3SEByzEnZJRyPZe+1Ujo93snDR
EQIx1UFuRHWMNmpu0dwOVhl20AZn6cwedDMZG/q4kAbVD8Z8hn466lOx03MOKr8s
3FUbdDWRx77hGdXNHWkw5NW/NwDExOm3VUf/s/ozHkYp8Mi2WeZecfoTu5Y8kF7/
9/pQvqqGtDiXzE0fYqeWUGAPUJ0AMfpcodX82mnxNfKuJhRKLZmvwyUzbLF1quCG
9fKadTWyG0JWLgov1oXvvUOCQmPWoHQh0YooO5ThZpecUgjd8LQOOnOtBFkueWnR
dP3MPRDKd+9DHuXA9krFHpuJiP3X9DcHAlGceBeSM0AuQjgGZBJl5gZQxYCnj2S8
7NGzM91avQ6CeYifLOs6Zx1XsZ8BAP2ZvkiwA2UpeC77iK3nG6QzN88hl89bMqzv
a/qpbPBPwho96+TGvQJDj6Rns/laBzMgMW06tqsZfw1h2gr8WtMfZYOdubrpyLa5
CSdlfIz0RztACoWcvvPE9JCh8J9WKnLHHB2kCyzzou3UGO1xyBnb7I8V7TRsf/Vg
+wgxEwjQV+0/vEswhpSBmANfovATfutxw5joLWvQXWGNk+JYfok9YzCUJekpGAOo
HIqLg9pCfY28eRvIkUyGSVCJf2zhdo4Hs7imXFN2IiSm+7/9a+6MxCLFRLOuZrNB
DjHnJ+efsCWUTQ7mO9yMB93e1RuqgxmUFwhtkhhGSHQz5976QqpO1/TzCsqmFIcz
GCer/rqbRid88oar9tSIddTvrJLtni97DimGN1c/XeWUn2odjDxuKEr4EXLHkx2+
MF86SL4OUiRf+IwRwyaSBdFFdyye//EHcyf2sqkwLSRNPT+tJpvOffU7T33EZ37B
HKyynb50n9/y6Qd7C/FJkoudDqdTP3FtuFKYqnN6KKz4f+zq0bo0f9PDeAHZmYNB
JQ6jTbKd+jIta32skrwKecKO0HbBsc6S+eCuKhu7QUh5UCCupXy2MUo6ht9MRTK7
bG+FScJsqAdpb7d7oYkAKBWBdu3hcqIL+0qHmRcabFvOuLTMvp+QNYEog2pY3XAn
aFbBavQhC/t9h7WE01CyLEmcUeEezCmp4yknuGaYQchcVNLwzdzLZsOYmleFzcKN
oR1ZERe9CSGy6prLH+7FOcMCKyf/FdtTQ/lP+54h75Hi9AA1ZR2NkVUvJnA6xaAy
iUl4cBLXBVVi3TGLEYcRrTUhUPGSyfrzFns83wjTdD33OEAX2Pra4Wcfi0KCZ1T8
H254fEWidpHPf7ofIuejj8IR89LvQhIYrY7SeZtk9CgxyaBThpNOsXQ/1fyDELcB
YE5TRBeqhb0xUK04vy5+T3bRL4Y8ResT2a4KcApiA60+TPR7mWYHG5w/v085wqol
53Hb5DYlJdhizLAOc4hglYbHUxQUidxbKCsydYJAqzQMzhuQlGsbF57c/xUPS5MS
moo1kF7iACDQFPqnX+lICdens7L74wJ9/qjP/DJfe8e34btb0rHz+Dmagdx+G2po
rbsU41Xa7bAMZj22En8UhYxA5j+zPSxydvYT52Y1gQgQkTMnr0LrV4CnnK5L2SfD
Xq3kaAThsL+HtJRnhKindIvC0geSvJPRKIUkWrT/R6l54l4xEb0W8riXXT+sINxG
R3nJ/uILSo4/4sbTuDm/Yx3OOE2AP6KoFVsfq7OrxBTaRRAccRof5H6eY/ECT7w5
vSbZsiLuwec7A3/j+1zq2gwoLlS3H9gjbVvuEKlfkHK/WAfTH59zQcUYEqExxldU
dxC6jipky7x8wYlEmjSuFOlrQUeNyhGBQpX4kzjEACE=
`protect END_PROTECTED
