`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uee5/QIGmAl3e0xoZ03Lwze7PKstnBs6nX2mjtDQlbEABlIProkm7K2/hwCgzg8o
udDVZOsLEJglZVe0wtAJrfR73l/vjUIkXiF4Ze0cs59sUQHoL/nmt/JdXM3Kqnwp
8ADfpKpfPXp2Hpm4P5jkSEOJlOPIF1Z7Gq6KiCmBZmqXNRNx6kA7VZi4sv3AKMYR
GQWv0e2LsVcdxkXZZO0UpCEzLlt2tfP80iINa923lhUzvrF4kk/AyMhmAcyVrEWE
+xd2sF3IbTd7m41IRk2F+HMLk7zUc5w8NT4TSk8IveTTisY+vhuf2r0LB+c3uJer
UaZ3/nrQB/NtkOw5hlvQeqTfY4FpD9SQ6jFLJnn187bTeJlidSvNRwsoQnrdOHzJ
xjF7o7VJjsAoc8eXE5o8nVPa0HxirFP8YTk427nQ/fy2ucqYyxDm2+3UWso94nlD
Pw3lLQR2Ga97txBDmqGnPa+I37TXzkxc0w+4x+4YkqIR/OXbNuULlKFKFrnj3vdf
h/PQIAFepiI1PR3/JVerckbJzoT/D/uTMAQ/fpOJgKByuaXdB5Rr6JKOgzjKDUKq
CC6ifh41J18957Cdx8BwA4x3WCeaISAqxd1MBfp4A3KpRXuvqvBFuDaimOPNb4OD
iAFoiW7s7q0TnQVYvPJE30AoHBXeX1zzT0kzd+z68kW6XJl+QDWDu6vH473xVv4B
ydWzCyuh+Lrcc9m2WRzg7+BcBtl1zjUDEy6bo19kwCJNTr0I7GDhrnE4hiONQgzK
11eGGjMFe9smfV74Lwp7HLphR+5lsMTqXjKpxWaGdRrYkXMc7SNOGFhqDv2lkpqb
d5t3Y04SBb+RhcWFqLjA7FuEwNJFavmc3qLrc84vyYnt2ttTpE/J1odp/6MnDdUh
14eI721vyMLdZ9GAKYmlpEjELokSv9rtM7NmtqR7edc39j6EltOg839oLycYRsR1
+eAWL5bviY/cShIgvRMJhfQHeFtKYO/1b+uv2Hy25zKc3KB1Y/uUrrCKM4xilMhR
Nz/IWNTg8gxjB4mzZ0CQHN7NaetV3jpv9kwdPLR+TuaXaWyL5Ob6HK+NvYlumvLb
cdfv1NyifIOl58EaCy+foFlMub7bOJQ32kUOjBxnCnFbM/To6aBlZ/pmCEKTe/0Z
xLcN1eHDMA1XKyqa+TeIpl6KMdw6zVxOS9BfBVtbIbkyilHC93ImPotA/IA5ZFxo
6Oo3vTbeW8Ju9v7gNVM4nes16bjRXVi9Fg4gq7cbId287O2CxcaGFzwmR8kg9kn1
Aa8sGYaTiF9bMmfO1o+AMIG4OQbJuEFGcqb1CDoDz5dFEPyUPcI+6//DQbssS4Bw
fBtrDeT8t/l32ipu3aOoevWPoCMtSgqxhQw9YrU+cM92mqkT+qETTdZIEDas9fgl
NAE5NP0KdlO8KJ0SzpnKcC5J/r+Wvp/EPUrfKumN1saBxI/kJ3HMUOTRRhHgXZD9
OKnAa6L+nx64qX5P/VJlc8AiVPvnSKY0sIGfGAihc0ZiFIC6zaoBSArjCL/nKP+E
BL0jAWEhN6uwg9N7S2FzsLzqiaFNp5YqAOJJqXGYmwRcQGzTiN/PGLgXsEipl3gP
L33UBkY70dStc9yS+KsAvKrSsIkQyaj+OzkJuCTamsJ7nESoWUhwGGiI6lEOfq5u
QRpJT4P7+wvQx4rbi8NJtecBk4SFS6HI11g48BxR2cQw33CiDOuSN6rMw8fpxn+Z
pAS4MJj3TZT2EOrYznUkdHpOeqnL72kzK73SizH/gCP6p/Y/oRm69AX2OlOtaeF/
s93WLacGSdDXi/Wv+99TFoAFbrVIZhkTw+2OqFidr2hBMAht2wEUrzckqEn3Usva
7B1PBPI1YyXpv0nLXc7rrJr5teF4Lkp48KMfn3WDIdPaZZJGNOeNDc0q5HkF58mt
/DQq7rP8VrVgQdwC4fRuNdM+eDHkoNdtHMh/MQtvKj1+8gtwIOPPqc00Em/DzEpR
mNOvJn5Qh3yhuSrU7oabm9Oq+bb/h/lJ3uUD29XC5Ofrs9nQTk0aXnQ3O4qmi6Un
XkbIj7anJU2yC3CKbCgO3UZV3HQFjyLCoQTpnBZuHuLaqFNscTLFc7a+mBirp8wv
hZd4I9C8zFhVTD4e+EyH9DiXRokcn0jaU+zy9dctIbORJInjtlovfdOenRXzdZWJ
grpidEOAmeo74vXz3bbUday3DMzsr4M322WSdfD50uSqlXWNWnXI+lSlo+O2eReM
pGGQoPMo+zj/0a0tExX9a65Xof8Jzozh0Sy8mXM1fViv0ADLYcMjbfjJCgxKZZTD
60RxWoT9Kg+HQfIak1AoMPjzSHQlgx5RGeQ9nJXr10IAEUiCKq8A7X2TqK0PgEXt
G8okYQYPZQKgjRGhz6CI1hCTnUCg8ws4mvYKkbMHRg562cmWywiMjyLfgqWrHWvq
HJuFUV2JDW23MWTISK6iIl/8L/ggUHHGmRXQCvET8mB7oZFKdDfhWsputl7itIAw
WJHhs8EO9WD8h6koCvayHklgXXNaRkByCjvQIfJSgJhrwFD0cgrRuZwi7mwc2Xjr
s51MgsBKC+2LyDsApYzOwn1J2gBZkgAzL86+NrvQH8chhbN91nu56PLBG0dmfprG
CgvGkhrTSQhBz/xZbOJZh5kreXMp4uR4nWDPUeDvcB1EdLWIsjVLCNmfcLRmTL2z
FlvReUh1dxmnzSgCw1FaHcuFn/dOg0bu60NVQc/DJYn+NHZxL8V9sjKNmzWOiLWe
9N7PkKURCIKoiJOQbbJXmvlzVi3//1l56Kh7SWWc/J0UZwVe4L2YEn+3XjlVfeLF
RJbUyc/9YI8NKKR6xvpxaz6h9+z4c83B6XNcAXjw72Vu6EnzMU/Gh+LzaNRW8ACs
88EEq4wQT7uEXpqMXGJP/cSWN/TF5tP447BE4iGdrSVe5rKUYSZAyUw/Cn9pjMNp
irqWb/a/mYa5+BI4DuesP1wRR0np9kIPcF3H0INs0lHZFecj0HCyZaZNjQRnvz9A
N8R6PKPurYIJ2ATNUae+Clui/bbK+c+hhHpNai/LdiT3gUMjrmQyfUI1BYJI8E/Y
2VSe6ncPqW24B+wOQk1CzHTPniaF/I5qXqmxhq6/rmzWQGRE+8o2nYFbi0SGjOzi
K4zxmb8ESMH98OExHbI2pvFrAsZLxbMd3q+7Y7b0ClvxONpVpP31OuXlz9iI22Kl
emGhXKINJ6GZjYkRKcHxTiSxQreawjfezPkTiiMJC1cWZGsreSsfY6Jo/rDb4qVc
EBpgwcB8ZZOeblzzrBjfEhmEoFE/G2q4+J4SWggE/d6bR3sRFkSdbJBg97Yc37N4
deIL8ZAPPvzy+lDNhwCOD/15im9G/+JItMVkCRf4sllOqjg8jMySmGdWozXko8B2
6WZtPuV1EuWGajIXvehECQYkCezge/RQyPKy3xXq9J8TY2+mOOyaTTPcgd8cMt/a
q9feuDJbDZsCrHzV74/wetJnW++ZwxDRZzzxQPoLYPq83aLG7FAVwl/DKx+KeOAV
9plp9brrvn7uecD9RV6pSDSPqja1VVzX/y5AEygqa4TTjxs+Bu6QPPneXAx1lyFs
1NeVyYkKSPhFvbWgB6epjwZl4mRl3R9kS/d00dUpxPPGoXj1rHqmeaNbxZQR998Z
RWDYucfEQFiyzTNYy3NKDf0sl70/yy4mX//twS//vc+JVmjBHOyAvQ7kQ+ghxUb/
AQwG2duCIAP6rZCnW0cYZEj+K/hovGcZTCTrtm3Mya1apq5xgr3gc0g6hbubqRYh
JsA9rH33mFXXJ4SNmHkTl6uUcsBq2Ep6s6HhxP4jC3HlU2ymLLS93BYI2Y8VpYjm
kbahuLfNXVfuDWUeBA7m45HD1LCQwQL5XN6cZpUfhguJe8kmjTUaZPphJ+L/KRE8
almRqyCF09sitB8HMJ/ZLk4LqL6ynF0JFl/5sCb9Ut98AOPaOSJhz8yUnjgMZ9DU
yuuorb4dIFQgurTztjnTwA3+4+yMEC8YfwmWEh81ILoRy3gS8pXH2mRczgP2ODTu
8tW5nszbQTAp9gFrkr8BX9QMyeov/SzcvT9UbHW6o2EAXpmqbidu9p918TRUKRNo
Ak3l/X92jrjspzlVuXmXQhsoPc7bR5aONqRI0zjVxus35J8+6CKVwA0ecezcgD7Z
9BwooD1/hpBRe+tEofVWdIxU+LwOAtgY6Y3Eo3eeL6Tgt6tq2dgzsr7RjFO65swg
b9RovYob3bz0hzjrTdTGXQdmioK3+FrD/bdKQRiXXtTX0SddLdGVMsEXOGja75AP
dEcXT5vQ6DRj5iWLVLPfHABFRrQ+gIzJITOgtvTHqq2SGuJDuRiQ434CPTUaQWA5
i3FhzNgxjGRstZLmTlpx9F2rFkIRJ2UmO+CYVu7U+lmEzCvxmXK3PiAY2JKUZYe8
Sl6AQuM6+HetzTxTrmE1rbFC1S8kOO3uz2AdJnN9hBM95gXZ5htIzoZD0hX/oceq
nUegM5gwN6NE7RZDFHTWPKq6EMD8UwVsK/bQfrJDILhrQh3DNwlkr6zEneQslaBu
wMgMTtNIF0GnObVmaHii0lJlwQkXVuP7dllPPQejo6vWt9LrX87OU6VyN8tKQjwp
hbcstTXRkr573ps4Oftom/XoLRuOSf9rPI2B+kqJ1tOQzsW9ntJewBh50WCh3uZr
7SxEFU8t0nh9MHpD8b8lP+FuK9on4JT8/O9sn7/HyR1hvMEgIy/JDM7CKjcI7uQp
gT6FWNYCetKFtbCZtcD7d6OUcRh9oRD6gWAP1OyGcf/MikCh60EweOXmAgA4/CCG
pH3xlnNYVA1QKKGsy4XrC8Ai+n52JlR/hpBlloe/05ESBDDd8RkOTBNENn3FlGl/
ItGaRO6a4ZwY02l6fjga8XCvjkPj5weIQFdoSEWcB4Us0EuzOCu3SOHqDRcdxyUY
J0dA0Oz452d/jBMKI0Nnld8uGal9xeI1SZsjtRWpR2khb7lRhbPfriRJsVhGKL0S
`protect END_PROTECTED
