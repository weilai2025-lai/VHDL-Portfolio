`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OZb/mFXGI+0Owp8IBTkTKek/evX/oZQAgbisw+fdKKT67cAjE1rhToGMikLRPON
Qhk9rBUTaSDGPuOu3OMaCetkWywCU51x5wmzRoZVABrMBzWIlbDw1j/quoAIuHAW
rE/DpAZwWiAJ6nAk6yKFbbexSWuAgCAKvcMtISyUzmh1S7nSMZm6oxEkzbUoXlyt
FSo+yWp7Qvq54w/APQ4gHb1pLnVDphB8Qzyqk+nGSxMDj5whZ8UaWTn2HM0AueiZ
c+KYjOE2wY8RPQ5dlLYN6DMbrUHaKyuLsJcQ/VL/2lIcKAUTaeUhRmNFdswEnNVr
Df4fZICVd5qHu9SLj546nqrV3Z+7qbeIfl6DKnn8HRqF9NeDFNc2MxHM21tHmJGY
p1xUcLfASmxKtOV12dCahCzuMNtQ7FD41Fg2gAGUqtESvJrTwVDYvriJtN/Lh+TG
it+2+IK7cGCccs5H+LRNt95ZhFDfIDDzNvJ7Ux0tTUu34CL99Jbs0wA7yrRv4Spi
PInl+aICOySi/yDlPDPCMQaPoOKZYXchbmpgnJR2bXxxE1ygH25ALPzD+pgUFM+J
lD19bAZq+/KttAQDvBW0xQg7HXnJZlTUYxZzeeGVf4K4TtZ/1y9bdWSA8J24Mjmw
6ahW4usxtsjSs1oGpCs1FYifIvLOM8yG7Dq4J+HUhcSg5c0txZFvV07L5d0OCkoC
H3xNe+G6UoiMqIhMJiqg4ZMwEEqCYQHOaIhI7ozoKkc4A3x/epOe+B7O64mBdnzG
dslHLAB3zbJ0HHeGgAGivlUiqHl1rLQElROFMDNRnu9xs/enxUeoVl1eZNz7nqCE
2p0hGPuYD7hB78Vw0kCuOgGTkaOR67RJ9a02ZDWHyU+UoCAuGVPuZc1fEwHHRNOB
qdp+KmSmQ+jszL7DwX4SMC6inRw4J5i+xTZ+fqcFYQ5M/oGA+FGkuKTmVLmDGw6n
ZI3ljLgE3NHKqY4LhbQokacYqdTqYbc+n8oyt5UOgObwACt8FgaIogNDmyYM3sdx
UAfppazwUQZrjR5gNRpKA+MCTB5PLehH0IVP5OmpPumgXymrXNecNqt+B8lvxVP5
V0qxPg4UH/uhmuVXD9r8+1UcPjnWaKiND0/gDBvH5yxQp3n1qYJgPfz/61+H50fg
jElslnqjXZ42tbB37lQjsodaK1w57lqMLrdrp7iPDd0cRwsjAJoKelT1aWxU8QZo
CBWUgDi23BA5I3f9yGjn7Lz3g73gXph5P0Vo8NjQvkP7xRziu7RC9xAdQ9G5IMA3
XfBRJsX2Sy9q3gIbcJiJl8BoFwKa6mcEYwPkLPFeNPctC/g30XjlLqTYYp50Z+52
63L9j9aBYeH8Huo04PQjAmrVoAaUkIdKWDwSdFuI18gPkCbIh2e6XS8JYe4Uhvbr
9QqzJV+oyEWReHPV2Y2Ytjg7O7vPK1IHjSyHL6Ku8OpnOnfhdfZMwZoLABGM7IaH
QdZldrBkwkZUouNxT9mlDfx33TofSRs35WeaiVwn7DAW36u245ex29p/xLqf9UZZ
yxPt3eESIQFq4joj3H5BzCiLJfdG+YJ+ba4JGDq3avO3eVmQhQ2mN/bQB4VoauU9
dipwd6J8glJlFOA8XVQSWku8+DH7nBAeMnR61sh3wyCaVJZvSLYq06XqWHtg993E
zN4kxHcxp1phlhfDwQ9yLlisjZ+GAJKaJMAw4iKc+lljHQ0LIhkVXe+TAK5o+RMT
jTY+GY8nEDgSyv3k4GFrWwNV4i7QV3bFgsXTfgN8li22xvoUK82AA5JlL14E1x6u
bYZl1GJw75PoSGTleAL5JTceaP9d02BOeIKRqfv7Rmdf/nwxz1gWx8+619tLn6se
4xbV2nXxRlOEbuGrV+swm36FUKgSpzfM0CSppkNCddewxRQAg2je2GWA7Le8JbEQ
AiX2X6VbddCbQApVWIEPufdq0iyDHZJvAnLKtQpB39yfCs0Zqg0ml67eClJ+hRRT
FSFlIMuIHhDK0va0gNz7PglxmPCwJHLMU292G3BvgKNWn8GVnRzYouUBl/M+VsJT
uO+MRu34b5K8gi7OpkZBqaW4sQ4K9Rl0uQTWK/+lbt9evIjTi9/9TfcfdHVVSWc3
ktysIdVcmlGsweIfsYdGv3v9FxVjTHHJQjn9eNvfhrev/O4mjTURqX9gWZXhs/M0
ZuTVkIbU02h6SdT0W8mzz7RYy4N3UP01qe8nMb6SlU0HHf5X230TjYjf028haX57
j9+nBIxKz/1WeAlyiSQ614VpbSGVyH2piPCiQqrPPY49y6F2p+j55h87JuWUxsYm
C5sP4FTPpFkDZL9qe0WmiY8xrGJjjzvRo2TvjsKakA8NJ/+OWqQy26NRO1z93KKW
WYComhFkuNjgpDyGjc/VhsoktRso0GxhNFvqq0aII/oyUCbICf7b11sIpxrVkWYm
paCGxDhg5ptlVvp6wCHQTKSaZu2gMwX/oAGbhvMbBLb2S5sujqOmqQDH6s8L9Cq0
AvHLlHtMbnLoGiPQGJ5yjJxEOvChS1Xdj9k6PyKAKMU=
`protect END_PROTECTED
