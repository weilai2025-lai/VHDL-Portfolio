`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQuuvSwL10YvIOD54++Gy5WbZbTjPV6fWE260jVTsERQ0SbJaVNenyRGi70f5Jc/
/9BTtmetQilYQ+vNHqfJh3Brjgm3OyCwHWlmmZrAJnki89OwgVUWhmTRaqFUbm2N
AZ+NT/FzK58jmw5Rt6EaXsl9iikyeUick4/V5215tgpITlTaPugkCa6a0N2pyXTo
dyu6eGcVb32K5GbcOwewY3mWbb+FELsi0OdB/OSu/bKGtLsZfsMHvDIvyq+JjBrs
rZyGIluD0SWJx6NQ2VbVI3mG3Shocdw5mUF2TdMXcK2YYhzNaAV3iSjloUXkm4aP
wtpkdmwLb7XhK9XBxmM4SEIQuodvLWGXm+GNiZonB5U95/PB1r9RaO5RIXmxWwo9
jyjrtS3aNsfZGWZnDkjlQAz72bErSmjzZD32XgwSN1zs8sCSkt2jvh6QaHTPelAU
cw+sT911OHL6IwU7zpJ44z8LuNCwMtK/uJXfRlCdDt6mswM1pgUNoPq79cnPntDy
vjNAylk9ERpIi7piVdRyzi6UqMyFQjmtJpoJcutpQ5wUoIANC8IS0+ZwMzzTyMRG
8eE+GAMdtiK+LbW+YJjSqX9+wsU1WqFPUzti5P5BGr6V+Xu+xi3SKeBAy5MPq+xi
7EipSPqmkKxcxw9J6YJ+R1hJgXXBoh2YDo8q1YQKz9nKoS6gRbw8wI4mO77/+JbD
Mp2D79Gf7C75weiYF/VnADP+rg4GhYxV/BlyILOCJnNI+Ft5MxQENGYlS4+S7Olq
CVRIGIps+v7WODqSkmJV63W2PkJevnQ0uAWhwFIMm/rIOZENnL1P+JHN88mSY9PZ
iNy9rU9SETU6Q1XfspufhqcsWy8X4dAw4x08Y3GbnDyku7QedJ1N74R+i26jaiiq
UMKnFTo024IJOV3tOUkn6sww1EdhpNxXlZs+dAuxXrnTh1fJLkQ0jnteBpA6nMwr
2foqD1RJiTGpmt5w6bs3r5RsO9ubYMHBB8dEDTCB3+CTOizLBmV5QyA/AOxrLL5i
L6Eg0AK7kJAsohaiCvVB3iH6fUD5gxB+lUrrPrEBRV3T4mfDqZtLtmcFhRKwvnDN
YCiqrupqmO3klytgQ3kw66qGTdU7nyxZ1ro1BScL6kznunuAEugaoPmutH7OGbIG
9hEebimCsH57RcZQFvZsOXnPUkS2yRckzBv2EbnFjHJ7PWxekl3rNmxE5BoQ+8vT
+FsYqv+PK3G6eDgJq+crznf2du6dzD4Gx+Pk8mrIAz1XQv6QU6gSJEp4KK8CaiXH
L2VAV6IISIHxDfYwvz6glE3ijU+fBaTEs4vg+QQiL+K+8IwSQregYvUzMW+QHjYv
QivJUgWuKxub4zcdMp4G38aTj3TkO6/a5iABjOUPEzc2wenn3g/UvcVNYKeGOd0M
EIKrNcLgei6RvCdX6aTY5fTVYYI6ciujz6NyW1a9DP1QmBUuWUMRvIdfnIiDrQn9
6yaLmuaim3FaEV/uXRNUL5yjZyEife3sqKczqxJghaAwwAYEMN3xHODLJdYqpen3
esgszejRvvDut5UrUURVvuwGzDQ6eUo5BQzopl+v0xOhPHDSnn1jQxCy1Vb1ueip
7OraUmUn0PBIZM+pqw3AJdLWhweF6NuNUl7OaDHeOF5VatAJSXjgZUDW4WfDlobh
FuH0uYh6HxPXg95dH8Jo3hG1KNjAQRbMWeg2XELeGoclVQ+RQ+Za/Cv7xJw2gyuH
xdpW18I2/pCDAIWNNCnuoKwTbAzDDquOCLSg8/wA4kuLtntC5U7J9fx35nE/FnQc
eXNl/v6kE5bmcYlbZdSHxPnyBb7dtjPOyPOQglxbv1b3POjcOyjHqvy8OrQT4BVQ
cVscyhpXOTXoAwuPPuKFd6uRiS38CmA3TPZiQhpPAm+JH8K1UFyrmzG4lxYkalO+
YxMQp5sBkqEeImPmohpgkhknmnjA61j0Ln+G9BsrM5Ve53AI1Yg5rUcXnxWgU/EV
1VlgFKrpCz91vp9sPKRy/XrxdzehcBpS3dxOgC6QAcg4fN2Rr4Hco68Cv99R7vXP
S3E/UNTip6MgIpheOZ/+NnPyrZEAzbSfXunZVMDr599c+cgNRhBEmq2XS7w+T71u
CSBYGmQ14UKRW5pFU1b4lmALcLAm4nJvA2kPBbIOisp56Ju5PHBBIaFubCNIA1vH
dr9AqRGquRDuNyr4TP2QAgw+83BjX+wnZeXf1qTLMp25ugT87boINhYAI9f2Cmd2
GhIN/Xzjc4JPLVc97SNZn9IjUPmzsXTaBJXhUC0Pus0OSndKJ8LsamlrXJxB4dCk
dj0Z2VvYivtbhN2L4vBEzg==
`protect END_PROTECTED
