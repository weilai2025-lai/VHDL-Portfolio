`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uprZTi507nWlEBJ44qbmMn/Ou34XdQcRCSH2W32BYXAiUlATlUDgEsOY3J6uqMwF
oybwO5bxdKjcw5xMiT/olTAVg0oGbLgC3gKJb+OVSkuJV3leiz0YdmWBdLjwqeqr
1/jVCRy8UPL7TfXdVBYfe1/WzfuSsHI7WH0ePk2cBfQxnA4HefCiqAB2gKVCFFTH
WJF7yBm5bBiARbQC16YkvhlTsSlM26bYCYCrRKYXsVGPKE1cJVGmcJkhK0Xk6YRs
9FMqcLgoAWOSyeDPNwLQwjYtCpuIUbyjtkTOucXhEIvuoGfDoHSTV0aK7wrhFEtP
Dy0rQKIPVajLstgvd+3w7/h29Q1izDktg0h9hq3pTn1K1J8ZgNgs5N1EPjNVVtnS
LACoXDv7IcEkhni/uhwqpuy15NENPm6s/18YuW40d5ar4qCs2iMXG74WYjcaxAIA
HQRK1uljhv2+cpIdQck8lQ1L5TfoLJUsr4qwQ/SesbBXkp9P6r93W6+3lFprPEgO
01myL+pZBKCdzGxD5C4M9eiAbo2YaAmHONuFbbNmawiSOxMeeHC5eBmMeOzwp63k
4lN/UcXaEEi+L9mAkTlZy1uaxlUK009e05ZFnrGin5WrREcI8GbICnV1cxO5bLWn
NhzX2wgUmpv8hCTUwRDxOW9kFztBxYFT3G9NJY26F1fnjs+3uVZQiyfuJMPJ4t9o
gjL8wUHxpSxAjeZLVQJ94SDv/x+WVi98+2jUh6kB7qvbz4b4IKadtoOJNi54qRil
2L3/g62kYWz1z/mhzWyeJgN0KxkxfNJYpjUB59wHoFF/LcqmvBOc9+bjzvnTAX3/
W7ByqjS4/o1/sUTPszgY6c1726PyC6tumdc5tDjtMMN3VGY6U3WyGq12PEipljRV
UVoQJnyX0p+sfgl/WkEoGh46RBP6XbwJ5qhivT/NNeAo9o3/k3kPa/aTnb/BEIxB
4kwdEqvk87SQbefvX6FMWsiFChuOwCJXBreiRfyCITT70uuY1faraBdNJ/rHNFor
09W+ghYYgI3pD8Va8EejZyPvty6PUtDorejYilKmUM37N7LAmzJKAHsDnBJAmlVq
MJxnohSDVaq3bUSH7MO/3ie+zvFYTCrDRphuY0YcIMOkplGon9VjbST3WC2Q4C2G
NnARZHAPe69Jf5tv6BDMfv/1NCBLUv2ZFE2/QafO/u3SdZfVd6SF+D5TDarlPJ+n
KDNnkfwz3zdz5qBsLgtreKdBcCFEONPGYr+PEShK7rqfmEPIstqC+w6CQ8F3dWwl
LwRoNZpN7TKCqe3O+d0SfNPUQ9v61mTcO94szsMw5ofoeunQywdPjI9K9FERi9lv
9FXN7TMIXhbkkTetDX2GaQF03cCNa21/RNmDimf+2DxVPsDrdWG1CN7oFzF8xLtO
CJVDMl5n2UoBamL3gdUWgzfM6Xiuob8tcwhubbJHWHR9Xp3rh1wANEqbCfRvJPro
l0DvtvWnpfpEA6CB0BDlz+Xo4PlLpmM857PScDK0mqg=
`protect END_PROTECTED
