`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tb/e/VPNlNyOM5RKRvadTNJ7O6G1qcd0OEur2+EyyYunjbymUmBex3bLUW0/SL+n
cymoKysP6QpfwjeShWOwUiQlH4Zcgle8fZii3kFRxTscqA9I3r60vKDUyDIhdwVz
828ONKgNJFby6OMXhgjsrMxeApgblkREfDARhbqWO4AvuttTXPm8PYXBXARvNJH8
C/uid8ylVFftw8OmJJLeT4n3ioGlTuzbFhH6VHBHZySTB46GvtEp7Vr6Fa4rRaco
Rz7P59kJPrkgBImKSfOZAVfAPq/nNwbCaJOMtf8SDcMSHiFxj5Ma5vuYdh4SPrdh
DFSSdoePqztuKe3LTkaju/aNDbY7h5HxOFKOTs1KzsLm9n2YgXPO8KXmwCYGJBtQ
UuC0fA65BDclN5ZUoOfbbR++ZZwSZ6JKGN1GCslSYPdrPRDBDNFlxJBhp+omXE4f
h3ahzeim71BcyYdXxFItPXsX/KYJ95q4g5njsgVWAUz8VCp/OSHF/Utp7CgOAjBR
TUdG5EoYFilNPbuFVtq1Jnxl8ZxAAuCfuh5359uQJ8UPCe0N3k8gw/biTfrNSUIm
nurokusjgHBpHdbhKBclfHPWzznsVXGVHoswmb/aafBQqT7a/qWp3TgeHxZbv71t
Lebo9VzncXIOPPCk5YTxvVKcs2HMRmzuMu3/GXAdwHXDW3TCy+J22lF5vt7PhBlz
PSajlfQ3nqubowPGFYB4fvgNL2Aa4bBhpuglifUUgIvk/1fp+EIEf4iVGfGHfhPL
U7H6ThWJgYLYf/SEdMqfSkuxf3KPMss//N5p3xPEVdXiOaesUbpEV+esGBmY7p9i
OufoYD8hR3eJhRi/40zxx9vSpdYx0d+VQIOzIZOvqA20v8SYSRhyMMZgBJHgoRWv
d1kTrkYF+MPXTbBfS6F+jMtDhGcbzKLc4wwhK43sSCeIMMQ/GHGbEJesQiwXVd09
NP3Q7iC6evR0VOwmSqzbiIPTjJtNzsnnM0KPs4Iv0O74GQoUKKA7DOe1Imv/2c2B
flZEeLTpG8tw3Ab0fmL+SveVc6nFNGdeYau3tjOib0Juw5S6yzZd8zwtxQBiXwJB
OgFfdj4ugc0VzkHLMaOIov/VF0NQYZMOy1IbztfkGXyguPZJY0u/zuommZ8nE2Ll
U+tq8FDK4Y/nTdVbQUln4p1AUgwdz7OcWVjj0PAaVTyXQmqkbD4Kb9rUQFQXd6CI
ynMy/1THTsfj3Jc1bKaiWlKVhL2Sk6w73DLk3uESnoIJ6ml65A/dlG1bEFGGRFRd
Zx02t8vPb+/68XBXLtkJloYHR0iT7bvf4gn8pgqww/nTSk6EPhhinsJHL4DMFEmo
Dm9UoAmhvPzW/v8N/oVTPrpUgc09znTeCSj2xcfvoQiYHwMp+N1RkNciGc7G9kjs
o0ZXbBHdMPOij95JLm6Uvr7IqNUd8XwL0DN1uWfV7M/qMyqiwq5KN33tzf1intrY
`protect END_PROTECTED
