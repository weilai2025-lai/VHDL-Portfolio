`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vlAM52OC1K0oVodkt/DGvUVQPxK3Xcm2CdCH6YFDwzR3mmnewhJM4Zo81SRjobEg
fapBxO/8U7wVnlquc7uGQ+1A5PpspIswdYdZIrFWFg1/+m/8ahtg5t+Qex1MrOMw
Ev2WHFDmvTuCTSx+xwvFOhdVAnIOEUnydUvqvJKODklY6wNWK6RG4ddyAVRjwjyl
7nI+yPp2O229NsfV41pmMye2img0l1hcKwNf1UrlAdQsPYzE4/2+Q7nMdi7tOYq/
qRFvRAzxf/dWTwOf3UiAnmU3sUUv9R972rmpcTr84oxQukGE0EYTbctm+MFgc5TP
MI17L59dQlY65uRVyN9TreMLleZZFKHwk4DAlrO2LQuCnFWy2+OLEOA6pbRHFNLX
tCCE04WsvHM7VR9FccNXvOvn+J7SFqVCOG/QN3C4eJ9vtUrQhx0bbyEILmnKcnUe
mxdYafNxUyxte871BwvPUDXnEdk+Ih19n0sAfHWw1rLSMy5xHA/Yvp6WOws9XVyU
LnYPqB0oS8BoixmKNlD8azO3nrao4UtykkCUZtVf1byxr/iM2xMsiYS6+kNfF7qr
9Ig+oovH00SYeTavJRk8Xum5IyAeQ82X+KP17ykoP5m+DxIoz/bxTYaPwfU4aKNj
1t5weZoiecPM7v6QfmIBddWdBqCj+w2WeQSycxxY3OYfzX83Q7v5i2ibWdpIhtP5
ovi1ihdlHGor6roXDZsX5tmdjwBfcH123DPSRZM/aSejJTXj26VVuybeV78Ojaw7
acRzQUALM7BtfcFQARJm/r/q1sBuqZjEZ2kEUD8g9rJQo8c87/WGEdqRpR8fhhyj
+aq5YHWSNfNx5lliCzUE2+JCc35Mq1FN611wZITzLvvnyh/lqM04gnlUAHf/xdtx
JTm8dXsYqFK193LNgnCCJOuWs0VDVmU9dNzeFvhuFTeG/7d0dID7gAYpSGX/avNd
+/okt+xepm6Ngr6uPjooB5FulF0gWuJlotC7J+4WQEy1yJ3lFFvP/3/DRMIFGMCW
Un2fj7AL2IroXYmVUiJj267G8/Jt6dE1ZDAe5SakmHAq5hh5bZ+Xib6qghuGqVEe
TfWCrSbzjJpWBOh79f082Q==
`protect END_PROTECTED
