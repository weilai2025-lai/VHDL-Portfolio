`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yf/yUOIexSewh5JD3kaozZ73fGJWF1MHcxL4WFbyi93hArmtCOpKDTFSWlGm40BK
lGmIv76eOGtBCqp4z6qkeyb7uCNoloNkkO0iUjm1U8yxsxYF2/TXPejBBGcQMQ9b
G38dFPow8T3uDsi6WVuZ6E7trMnG+McPiZsxBFw6vms4L1jv/fDur7e5QDzxfa0g
twy6PcnqX9ll1xfILYUVjNVptNS71h8V/lGDNh5oIo54eYk5ESbf/kMK3GjMdaFs
MgEjmH6P1eOMAb8Nn0Oq2Q6X96F3VrRx3eJoCzj32Pz+13tNMGDWMBzgGbJzvOeR
3A5aDKTSEZz1Yj3ixwfBiEiQQLuNRs9YZkP5SlUvMWTOaR5AH+E0ix1WAcxGCkdq
y8NbYEj2JOa6TtV+pyOmV/huvLId3Dxt23Or7Z1a0dVblkQ+AuTs2XbMxzPAhlqe
orydJYq1M3CXp+tRMlHByuVt8+fXmven5aSZFl/B8EJlTz/aKLV8r/41+2w/lFCm
hi/E/9hwdFJKLuJj+qSTJDPx9rqxWsvRlqKzt0ZF3N6uV6WZA05e2+dYBl1JnxyR
d2OjC8Fxu8Xmcmw5FRK13BHF8whqLIiJbadWUyTuC0LXcUaSB+/FYrktwLVYcoAa
S1Gp0ZWkRFEEpdAGT0G119Lt1nhELgTyPeWrjr/Sh3l+xrsZYp/yFumPcXq4qPnK
X7VXYQ9Ceygrzncu3qkzKwBuGF6BrSahBTEVxyvXelxeqwGYUGX+ZJPKG4zTIPEg
JOK6eJVbKKxnJBM3NR8W75n4n2o/l8gMiI/LiTZgrj7avTR0gERSRwASW/MG/NzY
rB0t4hLMXeitW2AZzVS42yGQBVDZydxDo1dnwWGR+M936r67eiHRKkttgTCV2A6V
5UNGCEVOHaLsWahlNy4QmdcMuNo7BB1shOd7qxs2M3ieS5EoMFNyJ8oOPmYeh8b6
4z28q68OMlRNYYwl3gLHFpFFFg/xuklxeke4dOUetBcEI4besBXTR3VP/znjuRsX
YVTDYwsNbqk6XpTATEKkKIRcg0Na6UaiynrEu7xvAGxgUnQsm4a0Lsx4Z5up8h58
jIHukqjwsls44+uWfQ1W077FhWiTmfTKbQPcRS2EPwe2Aek+odQ2EfJwJ12/AIw4
Aa6WDdrC6WO/rRWTYdaoTKM0fEZ4p6YBqiXocijCz3TElpF0UZwstNebGitv/q9u
wPlarFHi1AE+n8bYjxFEgU/UdxJ6bue8uR/dTx4Hm8N9R05tUYt/B1AODvv4A2Sw
`protect END_PROTECTED
