`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cvxTYDskKkK2F2pt0RKQL7fnBMPnNpPSOSoAh/M6fJkQ9DC3S1kLaP7yYpiK5Dl
iLOW25y92IqNFSTEQAHTldzLpSrkXayG+EgyTPV1mKJs9glaabGKOzgyw9xgesYW
sg6q6xdK3z0taLlZVYH6sCcxeOFZDQeryuorhiQR4MD0QrkKxxyrxNGlr/xxfao2
aj002GYcwR8ZshJM4BI4CCSGFBt5NkC4ElyHeeSmKzkJcq0ajWb7GXDYnjsP9mKt
r5sLF8G/+pnTg+6U1KkAedBRkWXou8qc+nUsnO5612Cp62jFMjT8D1CrgNWjIoA2
yOw66TaY151AcHybYhiRdqK4+L7RbO+D2kSNmvQIrfl0AwJOFSwRibxPvdswE+cz
+na17a4PUjZjVHa4+PjHyW3u6T4wRa/0L6Dg2+ryrS1f3TTsbXENPSn67CNlBbSY
fQQwxTLfI883gIDsgImwEPzXbUyQrbdUbGKhARzYxjTOwFK4BiTu/o7QBl9gv8p5
JzZVHwNgkbEnA13eXcM06BPljpLbg7JCR1t1AiGdP41Yy71ymoc2FJ9omvEAB2Ts
GgJTCY5XkngZ4QKRwMF9gtyr0OQKabWLhzgKF2Jn0biCJgAXnXspqP4Zojdr7Bqb
f8XJKkbw37+Lc60MV35I9xT9K/qSOVMlCDnIg2lILVldODVHPDXPno3DtGA3eKeB
HpI8enRlWqte572Bhni6KMTeaY38j8U6Pu5z9qSCZNW4N0SVQ7hyEv7OqgYgsVuZ
xXHbkmIXvciY3Ksqp40aOE8qIhaSPbq81ZAYWlXuYsJDZKMdCWkWl2lhpM/yyVtL
njs9LKGRZbTi2ztTSNmz1Ixd8s2e7/UydLfcdK2809lj2lpLdXZWhxLaNvDK+GcN
4kQmicBSKgURBlepprp+8WpZFn08jNnr/fZttxtA8T4g87KCNd/c3bLLb1BHrog6
RqMJNLlFtZ7XZ7LxWdwgYBuc9botw6GR3cvpwXJ9tl1p40wGYGiOXt5i2BUXm5eC
R3nlOgdNxdq7ndhhjtF1bwrYwgCYrF0SG0fESqHbMkgSu8nZseDUbAQmjQrVVuSA
B6T+46I3vONmleZUFaXHkHrVcTmY9Q+Di80IhUa1qvfT9IaBmtsn70EbC20eEc7l
hmjRhtatArwg8ClUCkROcwNlf8AO6QmWbyjy/FwaEsPT+jNXXiJni7QtNqMwb7fX
t9VwNuAMeYwYlWoPAVwcOvasvXMfDGjLFXFtWFNoHfFUOifPSJl2WelCG8TPAQ1l
JiYv26m+NTN5GBrKuekHCUDN89EN7yDDUwCXvJaq6wwRC7W6x4JCqTjUktCCy8q7
PdTQ5kZZGnL4HfR7o2xS/IR8zhXDfw5NwQnumiM7UMi7iiXxmRhaIFD0NxOfDJTk
LOiUSdv/0Q9myPj8FUdZcsMK0rPCzNyJogasXnwz8UnYkH5ngwL1Q7OB5xq9423y
pkZVSSFrTEEniwbgXKTEQ4jJLurv/xJHJTR0BAY5Efv5/au/dMsRk1hkeQZz7FOr
xVk9S4pBd0DNOVu8TxlOsGZBCmM6RWEW/2ksofuhmY/1zLbJ3EgOMDKurwVJwIGA
lcGota5u7lVk5YSq6/W94Pa0C/RXuZPHYayS0KXfaDzODvCJEnxmZYD4MSmJxR4Q
fOWoKiO8BYIh6xtG/II99WoG+CtdWAPgR1lcS/I+6JZK8+psf00sDUb5WEvd5AWT
mCcxfNNtHYfoEs1xwnSCY0Lnof8Roe6k91FiEBhP+GmhOIawQaEWgiJ1/5btbnVI
GohOzdFYWk2ba8D5H/DAhi153iRnvpv5kVqtmxeBWNQm1fnHs7FQ2GRHfrgc1Mt5
xk+T5U/rNKh6sJ9Aei73YGBTT4oMlm7mClZ9hogyLvwStSWVyn6VAArYPWIrpXtI
7VlcQouJVd8KQduGeMnc1hZKSr+IThWXEm5e02wpO5r1lCx+ZMqicwUsa/BnWz6n
Ffjipmlo2d1MsRjHhlVPjLuS2zCimx+PP68JCqFIIrgfrR1GWZ2DnUGeAqzQPU8i
qrsGSkz9TJ0vizjrd4xOeuFhreBDwC/2k9UsdfXlMWOUMk4EUJ/odX9CQMorbUxu
ykskzHcf/apyFH/tnOCwqMXGDfowF3pTt1SzkAxk13gcoeDsw91X3GMw/JbO8U4b
77E15wW9o0vHdkjFPCn1CpeRN9rLtuivlP/W7coq9pUqIlmXSwHaPr88MYF3x5Mw
vT00IfntdhIWT3AkIkUxbzkxtvVobH2oZwIsAdmlJ671fX2/tRX/Okw+8szxhA3K
I7t/gMLf02yHuZogY+LDJTVbLXdum94q2EfD9AUNvfHS7odNdK+R4smo7hizRr8L
sbrFrQAURPhCTu8t8kSBWDw1lGIH8ctOgJc+X7HpjufJHDU1v4tzIwB56xkJrs3H
d0kMdp0SFa3TqxJCb7tEYlG03BbmQLuW8cSfDQp1wsiS7sKguK/aF4id8Tx76JhY
ketScMI0sBe1TRFpCMJgRn2Z5HHviTaByC4+gEss1UhZItC6z3o/tBf+gn54dFAe
86IMZJzf9w9EfU66hFgLgCM6zaYX+j2c9gyHlAt5qdsyMsQtV3alEHs9LvkwIZyw
yhc9K/aRg55fC26QNAf0NOf9OGnINMXy/bPY/avHtE5tICJhyTun2sth+3v30AER
9zITxjuxvc46i0gv9F8Gi1mEY8qEqDQ6h7y/ja+pLSOlJ/IMgmi8paG/Xw/8kyFq
cBpiHv15eUopWD86juR624p5b7hRlUUbdXHlugwYqvqqisIHEbCuy7uYEqp1UjIg
eB24ShZU6qqSQpCHNtLLGCdpByQlVXwW4JGrHHS2QCJmDutt+hvkMPOZDGEZncZN
VhBSp/c5aUSc9SKuqIJeVRwBD+PDZaP+6voahYkQ/pc5HcuQPWIRhpJsOkZOkgTd
2nEMLj194NZBVVvitfFmb/h9wnKWzJ8gNMnJ8IY4qrltxQCBqghCWd8ndoYlGan3
fERgzeg1O+8PiWvrVyX2OZa0cJMulWg/qS9ojd1KDLcQoTiBZBEe8c+FHMxFzPkH
3+mWN9AZ5k//PRAAT00JfiTPFF+NhGvUlKdTjDgSxwDSvbWBHnIaqVUFbO+9EyBS
s/sNl6v7dqQQtmoxymG1q25jB4H0lTn8JSo7dyDv+byPP5w7JCbA1z4qlZbMG0Go
MqwXTnCNS5SHe/EsUWisklRg1YCUE3JJDNtUGQANmWOup98yxvPdeQTC5n1HCe1P
UyiWTprRe3+p/rvAEBgPXjiKYq8V34XaI4qWg+gFXXG3YQVyruK2A8zp1bmQl8DQ
HuvI1VTjCjup9UTnUFIJtI4Ocp/O6OclrshUv9ZHwCOWVbOgRuwFEjzNx0ctcI5m
sYZl6pXcZ0MHbyPRD3ZXMU0j71mKb3dyfDUggo9LhGt0Ln3rSJjnvuQeeU3CQlf9
StDYpqNvxNW0/5bJ2RZU0ZsxPhQNTY+D1f39l5ra1Q4pQqo1CglS6vc4DvXLFCRF
yg6nL1SYdAWtRvTL4Zh4FR6w359lZ4qkbFDaJ9rCX5/TPhTW+ocwwarmXQQHmyV2
xdPyLckdfg88QGT+rxPQ2KdAyig1cfhkWqItZRl9XtBdCx+hB5GLC0AO/BGrZvwZ
gbr9EM+iy6854cx3czLCPmSl0KAjfR8a5dbHrZ92vQ4ntw48bc23Djs/bKuLqIvQ
jmfHKcT42NUV3FTknSAfeYSaTS84x22cs2ypEtW0q+Wt59ZnPf8bZ4KLLRJTEoQi
JbxhGcjGxVmM0bX19V/6/rMSbSP11+1fP4cwrSQododSEDsMman/S3bTeKGNZEZW
b27bAlu3eor2YC99xt9iBw/W9xNpCdcpALYKNe1sMt5BOPSLToAIPyKWt/Lk0F/6
U00CgQ9uhKO8KKWBIDaVJYEDCGHeS22rfQm7C+DguAEOq0myzkXRx4WVpls50oXD
TmFO7qoCT1rEX0AdEw+wbRMbY9MU+5nggoCzuWCCeHGi0X+lt4zVcfhrn2UFWoQZ
tG+1w6326t70cnUYgCvjaBb+5n7aQ6tf7NwEfJZeK1IObfwDB4kTFNw92gGTz+Hg
ZMqUmH0zisTG7VKcAmaL6hrbs2Cx0z+VTIllem0lX53ffjA1J30nXGB+TtBuIeIU
13bCWyGgTz4r9heLqpS9dLBvYjkPNN0PgcbfpJVYyaqvCrS+JfkEirbFaPeUQc0H
y3cRAkDxELx5CRGkc2arJfrtvlUyeFLTmkwmxrwCjy3tW3hKygCI1ElljEp4LcPF
wWtrIwV9i3TNuOZiPl9QZ9KLxtFR1AD9YVPLHCZanMKQi2gdaJhFmWDyUtB0/aqH
Uuame3tNzLzeMq4yHafS2n9QPfUq9GmQZWBfjHr59C5y/i4Us7TQx5FSVSpIgz+r
uhnNHKAPMO2VoIKzG9ZFVS3iM/wb+UeXEOpoO1l9gY0mzSOFk8NRKIaDY2LMIw1e
lU00r6xqFJkqZAMujPVpSyapcKAeVYqTAjnQZIjQqhMs5ZRfGnfQBdyNp/tXceLE
zZAHp4BQlhAsMQoHtFGKe5gh6aGp7tMrR1Wy8f0wHf4dKgcThqTp2n/Pug7V/zl7
qjRfI0WTXhdNirhZ6LO2P/qrlUme7yQ71/ZFiAtMny9wZ76mRx4NrWn/BHsHwXlT
VRHKvmvBTNByvzJyrC1YtMXQUIJIbfnGqCa1qS0AMnRRKjCM3R2tcA+sXvLfbd/D
azQUJLXXtaApHzUOOaYHwWDyvow9pVrx7Oa8EYnV2kWiXQazY9huU/Cr9/H0LHad
qVM9CJkm/cahY21bxRC80KP3tve9K4mzlv6jqmxhwmgIafAuJq6YXl9H/PKVEe1w
xmlz5yvwer4QbO94bEXx8qRGlE0B8Aip0S+qZRNmTDSXVUkEsaCVEsNvkWZ6wz6j
NsTDkxJqLzmAbikr9YC3/FoJ0hnjV9ltuoSUyVlBE5C3kHKfAjF5k8THq5AwpNvI
/QUZagaECyUspafszTjdOXuU1+vFlibXPZHvBNLd71g88A5Os7Y40iPTWwzFNNbu
+q5g/dAEvKv7O2ZlZ01MtPE4n7JzksnhZcw2LIEN2TIouXIS2bmhYDr11o9pl9AK
vj7/PEXXdF7UMOckpaZ6UqS6SuvkOBkKcvgneZ2cZvlq3DbSyl7v76uRPtam73Q7
TQrvMlsebIf5jL1NQem11TL89WOP4kkMfRQEEC3hf4vELfMDLZbL/ohTc3Xu7vBH
tc7Tp4sQLWsdBX6MkOTxzR0ZWQDAZ4xtmpjmQiPKK741QTgZ6pArv5j13F8bL6VC
8N20OvFWwlLWOp9gROTTM3CG38yG0tnpzh6cPgaPugGjD/1dx9KK3gqzl7cfYLL7
xe0HqVpUluG3/ovPyTrrP4W9cdja8HcbreRtduGf7eruW0MAd0VjkuSha0Kid/ZG
GyyTCsN4aX1hyyo3P/rlZ1/KTxANI0i6DODI0Wa/H2+zqwtxN2hCUS94zSarRSee
KVPZX3wr8+FWZe4Pbuk4LUHl86MaoTStzuIPPzBNttF9OIHHidDEyahkQYntAk7O
lDtQv1L2qgRjbN0rhS0AlrdfDWsQqf+uwQrTqCa5fj18wN3ix4d8gux2x/oOF1z6
GA4kCfydfPZwubXt83v+xGldak4mCAE80+JsS8joTJKdPY/tGMc9mbDjlj03NFtm
7eWH6174aQPZu9Yg23rrIVuiBBzPtGgRyzb2t4iBYy1UpaP6geD5RpBJulpKIqb4
3UvVJmf3+l0qKdKFcffsF0NMDYddwaxevbd/kEDxs0uIZ6938RhX6TVxCHK+2SeB
9u2eUjRZ6VXJb/GezXYd3mM77vNnk4KaCEe3XxNEg1IPSRtOegtojPXclG28fafu
aTAB5c/lfF7jXVBaub049aQULw1SHeJD67SM55u3lhM8ylc4wG0Hb4rG4+/AAGC4
XlFX9xL9ClwmEJtqxeken+yzyK8+pCVHNN0c8wLCPOA=
`protect END_PROTECTED
