`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eacKOGlnkLs/z0QTgnTmqFRH+7mO9groRN+HpIkZMzHcP1P9x87LzP4NlUldiLo7
VZd8IfG+Kr2RiNZl6v4iq/pgSDo2HL+tw/STnKoEqYbQZnxEEkW7LfKgfEtfP5OW
VDz7ocJlNhbuALQ82cpu3hPyF2MxCacvzYKi61iOH5AcT1kaS/dBeHBOvwCOv0Dg
2A4JHm0a8B1b+PwcbZSgqW8cX3Poxkx2po1/akOMEpbLQQJIv+WNAZ6oerPnozpc
xY+jYIGTgvuqr6iYiJMqh4/x+Tz1PgWU2CNlYTTcjl4hTxJwY21Vq8djP3j8/LNX
5h39vT5OcRGRFPIKf1MfA6Vf8rTsAJNT+vCqaDbxq+gRgVaTV4u0gTDIa3B5bUi2
WaY+T0GLrECFNmTkydF/TS8vt4ays08xIx9vDfbHA1Qz1hu4bvxnlmTMqqEWf3hG
9HY1BkUdsHp1DActdYKEZIEelNYdrosk5UIfPmPjqPYwA8pSee862OWG7mBqNF8f
vEy83gDCPkUnoYsuRH9J+whOH0mbRRne+NgWf3zXCq86GlvPemAm7C6p4Mfnxiwq
Q1jMQX0TQzPzUjtBVQdoM7iMnEnHypRPshWohsaD4QnzQzLxPhjCuZGFvSraOEo5
jZXmuALGF5m7hMePyRdHPik7DDfkrBFxR2KdX/zlgVlKXC9vg1yqcsRJLNEQz//m
i6qEwI2VW2C7xO8dEQfX6+hgisI9YsdSHwcyhwLdtoJrQZquyMjabglyCOIG8bol
zG5ZLFjLNGqfOLd7j8jPAW3yM71cFCSDekf726CrR7LVu+LJe9dWAvjjX70FcJng
FS9DFZbYmtQWsdIORGG/199/V1WMIl0DppLVUlsBkez4CjJGoMeg+CPcYonfSx1Y
Eo7DNPttboYA9ChrrHiN2gINPKyD4K41y+IGS4Nk6DFOJQzfSUElITidFq8jiFkO
M0/tufGHdu/J+3IWJjZPRPb99reW87pA6X7Yeg03Y8yUGEebP1bxTUp47X0QFwGp
wCvV4pDvt6H7vEe+FKrhjg==
`protect END_PROTECTED
