`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PeUk+8RxfoGdGDr3k6O/FEBgvmwFBQPSdjSg14CT8/YfIQYbPk3SBmD+T6R5vV5n
o88ywzCuyrPWOdkSoRgwG10UpIcr5mjF1Is69lt02yDTEhPXGeI705LAtGkrfrUf
mD/0ySzuPit2n6RSqrIB5mMc91tG5DBIxFa+0WhppJYoyqOtdgH2l1ZlaQ0y+Ok4
OslNV0J9TaYYS2LXWeAS/6g+sIwhVh1Cim+Y66XpSNorkQhja54ih3nymkVmaGh5
ULb+WKmfjUnFZuwPLpGo3PG7sXaNHhc4idYAwGGF4xv8/51nVvTGbCoSBEnKYqNp
Cz0VoNFkb1d8RAizHblDE6kB37giBM+1Y0UMq4NroehYdzuI7iafgad0OmUEJmhW
V1CSvbePSdOscU2GdRdNzQpTBAml0JbCqoauqB14qJegz/JfX823lg8pj3K0rgYM
I8Jo6qbxmLrBMi1Nyv55VWnqu5mYBG8ofP4V3GZIpKKlekO8kJfd9+GoiRxJ7I/u
C7hEc3oeV3wrD66F/AEQPcv9t1gSzVWsNE/3of3jotf8ScunCUSp3QBw6qH7biab
`protect END_PROTECTED
