`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8CHyGvqgfzeOPnCvFtXHudXZfTlNOrBw7w0TBHDYiaQSb9QuvpS2g88XPrCZCJ/
A3k0Uk4uRidodVPCcTChrPz67cCx6pFdXyUTJKYM8B0AUJ9M8rUfAwiabhe/MYSW
c4/XpMR9I0D6bvx+MA4ZP33NZYNIvUKR8TKPhpwXwtsmOpdS0F1O0AQ+M1qb5Aw7
2nsqg93EXgXljLzFOrJ6sGF+gvkmQeBwoef8QsCr+fJthK92ye4uuuB/o1tW3VTo
2hoJC1SC3IOGl+/6mrOy7ZEdGR1oGj+YUaLgujYzTkzYcVqnp5Xo/pBSz6Tq39WN
R7kUabYYyBSXAKQ5GGi6kmH4neYH5pGCWilW/fx2vN9XsxZGYPLXNfj3neA67oWu
C63gaAegrQj1Fmvcgm/PBqsKxJ7TziyR0FlxEfJzo8hUteAgj/wU3aEurmupcQyS
J4OysM1xk4TyRoLInMxEIIlY68nD8YLOWP1//ESTe1BOprTUJ5QT19x65ULlW4E4
EgenQkLU+oIwwi2hSallilYWA3INg4CBYUcCURCudEHYca1HNSvkZyoS4DnxQli2
5jr/hF733/9D3AAvkhCGFUOnn3FwcZ23AjIQUsPgs89DgLNp3qQFKgngLXwDQOIA
M4duSMSgsaIf+0/Z2FthLvg9sopYNuvuIdapmrt+gehmbf8G2D9jcU0/v0dRkfmQ
l08pYDzdmO3BX34lGZiDi/F31kGjmq8cJxIpdvBK5RNlMmpo4Pjw76lJsgj9zMdt
lSVTRs8r9vrzo4LrCndcDrzBcYrkDP9A2JDxFvl72lYD6m5mE77LGPxzfT78Mhrp
Qi95CvZnU5nYYYyv9ncH//OX2LLMlTQ9uUo34ULoFoHutk10TBSubzjdCW22GWha
Vv+rB5yHh1H/sq2aGa4qQuVfPSzTvLLoQpj8ZDLWxlYQfnMPt6ISkA66d6qixr49
75YwDqbLp41X2ILTAHhA9ln3cY5iZO4B5qSNHprfTN9VhH7ljsgWxJAJ3pQy8PFK
5nSiUy8vPCu7PtwSZxgJlXyoRZKNcFOrdGYuCg1Nrragdua4QgE0r1brqSGsquL4
uWxZ7GsYryMm+b7sapD4SuvwEk5dp4a7V5X16o5/1pOqTbkT27bTtES1ObcF3ciB
3XhwHlclJGANbxrmoDlOHK9DxXhDVJt7+y+RnlmRiMdldb1wWBz74sv5piG7bEj+
uzEtZnR0Zjg76UFSF5Ngl4qX/eCMRQWjsw0Y61TIYQNFYJQdGe7b5OeelwsBcrJE
k0C0F104EhVabheZZ7gxzToB4E+wsNtBO5Rp86uORAaDHqBtaxRo8wyrHtRF8d1X
bJQyj5Dq8AqRF3BLgZIO2qibceRKXe1nTsbG55ZvaS7b6LZrxtlmqhtltpc2NbQi
WPbD3MCtuRY/dkzN7aqegNuYun/C3VzUk4ueTMGOUZzRObMTrknM4zgAomj77r3A
abtJwoD7YP3cztrCCPQocWNL/nhTAMaL8yaRv8A66JPigbOH67XtEJCISiNpYFok
7YE02nfBxfuoXztNNpSXW0WCQs16sjqDD4X4Jvky94jqwg0ZXGCSdQnLSnrNNK1/
yRmK58vTJZbJqbXOjzmKq7s0ioAVvJ9WKahseFH01m7vQa0I6Qq60eZENYMpgm2H
6+Ox8OuJaYSNepM5dBv2TkDZs0zc/2htsQgabn36YsXNFHofa4z7J5yPzs6ph4fW
vYin8IbsJW/bcOHvnOJfEp/Tq4PqnB36ofVmczlEEJ+L/ZKCqp+fe83M7xggsxBq
JAbVo/z6Dp1VOZ2BdCagVSrTXG94MpMUq/AVeZ495/i0putldMqGjJOPRZw2RuQF
kC0mebZ4FKlFHtYm4E850oeShiT8OE/vxKRzHU0B2ESzj4DOF0uxtukoD0uwfFCm
/+R8M1ypLAzxXO3Vij/8ZkhPKnJvlyo6/FeLN/0KRfs9atnCXdvuEvjj8YkHi57S
CxD0+Avw+yK4hooG2SuIln7IPTv9y5qOhIRjiMB4RtFmuDgOEJOs1Jcsv/023zo3
J7shcRKd8N8iRHDvDsAK5G8iP5iepNt6S4dNBm/ywUDhKbKgwNouy7F+IiTbDNBu
fIClaI2xB6ibsynYucJcA6KWGy/6DLuTM+RuxX9PPFNIVtBFiRfNLCfwuk4PAE2X
Yo/lW0Ae+AulQwitzKB5R+yZFoaCaQcXq+6lshM++F4wY8Uxiqzxh27wTf2n6IE9
L4v4VesoJ2YD8eMUsia7NFLDDfdBmKkoN0/tCLB57zqTBsSVS7eJPCpYfy53vkdC
EVpdAWpZyLZM5HVl0e8HOra74W5qIQc0Lzr1icLLlNpK6LA62KGsBaq3F0WJnZJ/
c6TgcV2Tw4pEvdAGvu/Ju8g9g+Flzyl11pUDMdg20wiqtI12/w0qfoZwxHbpJUJ7
BoMOvVO/uV7I79bEtEa7h1icnIb0COBp5RoLa0xrHavW6GZ3nkcb+VnfXD+mi52Y
nRXSuut9lZcZZoTrll9NsiLYSuPznwF0DnNEYrZ53QQzeVp96+7M1HZhLeM7uOPB
d7aaDQDPbfro6P5ztXO1fGhb9Br6YfoT+T8xINKMzmDtd4LP5LeN4CdF9kmndgRu
AEgMmP8nBy6IHNnDI8SCejPKH9qvc/X0xjgHbkXEp3riYSghIN6Iek4y9c7AdbiY
0hQUx56qlSNVUmyHIGSdFNzRs3u3AJ4693XoC/msDi+9jYTnhiS4vpMxr5siqb+1
4+c2CVRfDbrufKQ6X0MBwGkZnBRKJLWOcOGJ17n9IKUT4h6HqkJMS9mA/LrnkNPm
K4w4BxbTkzSKvwsUl6+FduKTmQOSjANdgC3xmuZUAIA=
`protect END_PROTECTED
