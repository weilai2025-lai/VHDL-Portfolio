`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkSNtXKcCWlsggj9OzStdxdWwnv7gt/juOmj9mCQQxNFNWrRG0KAgByxAT3XJkLZ
B2bY83g3ceZZZD2wSXmxipGpFlHoOdtYssTNTRgPGZoMEipryIL6D2d9islGhIq9
Q94BdUuGCd9VWzwy1cdnjbFfOoGCXtQ3cUv3cW/uvRBnGrm71endhEEZ6E4mDf9O
xx0bxbgUoZwzut0Z8xWbjM/QITgdtwco/PuH2+WROTr0wUfCYFVut23PpEnNcfX2
SedN1mck03I7p0J+fH/rDKoqIVeXFDSNW6h/bEWKm15ZXSJrW7kQ49dcazdVzY1x
I8iBwI+3UVUvMWPT7+WveR2wN4IhW0xDlY8sovhjL2dw0V7UIGt8O9KjoqXBehLZ
iTnZLX5NFdl8uKC3egSrWNRVD72Y/hmSojf9ndZTesAe3Fo3ogcYCfzeMQk7vA+c
+FJfmhJzkktvO47LrDoNz1BAAoz0ocAHbad2Gjwg2s86V3VvWWVvHrdKDLv48KxT
IijJDfMbqRSCMRs/Yol1HbZ/WOW3h1hqGxErKhfNH2Q1fIeBOL1bmQ9YDWC4f6sC
gQM6K7ao54U6a4IXD/2vrc3iP2DVAbNwOWULJxhYmH0=
`protect END_PROTECTED
