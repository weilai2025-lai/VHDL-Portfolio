`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YWOClQgN51IaHmwlUq6i4L1MOaR/ZiRina8HJ6uxE+jO2fezc1RKJD+xH8f9nvvr
C58Nq9x8+oWwXhnvSgMCRaz0W+vbrOXG0ajDgN/wvlss6sr95bSIvXBx7DkoY615
37uhnVPRswEIwe0jQY0ZFpSS8Leg/ZtjcyLKluXxPAX0jGzBuqYyDhTUJQDcbbQE
SCc0VVGShHyGzHGmoDNl9YElRRQEy2VLs1K5GEJ61LTATLEhNGmwjOGmxQgEMTdm
vtEsXU1LtO4XP265bYDqp6dSfKU5Wq+7OyjzeSh8MFqjXttAYcyR1IqSv3/qrani
ohz3ESaQ57++zoRWGmpaM38sfmdkejn37WGFE3rXtfteieh9MXimMMEHvPdV47Uv
fF6sz6ph45COeACk2ef7Vs1rTFO0XWChZMqU3iRIg3HKHmXOr+PiDT7lAbzJTKd4
t3nzAwD4e6c17/xA6PaFnNPouFoFkdF+4UMYx84HcZTVy4P1OnlpsTknh20QhlU1
f3+2RB7n0n/hw68BfCMoB9tuHwo+YcyuBzPLC/Qietz5XkwGV04aTeRiKv0ERL0W
ORa4mbcNz7RAOv9PoiWTGQpGetX39dOLrcmaD9sX07TjYmvaiIozP4jtf6o5K6gZ
ZrQtF0hV7TbeHdFywfPUimueyNhvcElWPmQZW0EWcGjy7+09Pr0gitmOUskhVxa5
Yh9IDSkYnAb4r/DRcxOv22xIymFX4NTP3JzoMh8xehIe8y4bklaMcMi/r6VVUTM5
BFtg4BghssjgFvpdH0f8440/DNzJlLYpf1kqeEZsEukoTkSGu9V2Pm07R5+wuVsZ
poBhp6gwKnG4cGgnu8wKQGFPeY2Tu+dmV5wJot6629Y+wED/2s8d8NR5PvpSBc49
aJ45Se03McAmgRBnVf5xtvNWHA/I1NfXFrPfVShst5pyl4jWLpityoQPPdRcKLS4
E3dTnq8eYlgyZoZXV5kDMz2I688oDX66KlACNRmFcpZnVid1y4QK3VPpSLUio9E0
px+WI8DI5SWJP0e6I1rwhDS37r6UaqpE2Yl62fzTSLMWGy5vhYodcDe5XuprX7G5
T+VYmyP+AphWtWFpPdG/ArzniyfuW5iC5d6IomQFjRlhLMByflIw9r1AfeC7IWck
at7BPlQ1pcJizPzzlUNiNDeNN2FhudnTNZW7Um7xqWxpq7sV96xaqyH4NQgoS8X3
RDKlHfwdRAuvnljBvpc5amBO6rtLatJ+FqNQN+JUuQ/qb7s+/PRSR06PJJizV4yb
r/5d1roGgY5OZ7+8NNpxjg93Es0abnQdT/wKzUW7S2w0ZkxlEnOKbGxStkr4kH7h
QBh3/g/3IS2s7v4fOYBrfM7NFz1HyDoxuGpkAN2moZyhz2r9EmbYU/gAimvJssZs
DdU+vmzxU+tkSLoE515HJrp06Fo2240XZSS4hqKLutbWFq9cNWFB4CWFedc8GwZU
gnjr2IbE2EsAqjKzCCH63XhxBd5P+asflEBlQI7qtAF7jRPvYfKv4MXgGvRG8uBk
dwxQFcnibWmQOPG8X+wGy+09u7y3+BQoOxgRyRXrQNC47KixNi6MLEqSSKPys7tg
dXHiVk6xWa3ZqCVXiO8rS31/12xegiQ24ro8tU5Xb2noiaDXz339zgSz1Tml3cY5
Q1mpp+3AwtI5aDL3J+bbWQXM5aunIfFflAj24uVj4rGpQwRDuNro8oakLhaHdUPg
K+Lhbm8OEn2k3rCr3XlhTiJGbGiEw2VUZ0gYsL4zUGhS4M0oOtnPy17iWyCBpP2J
rd7LA2HZxWsWksJCP98vu5W+uRSwz9iti9MRCQ4oRvRImy81jAE4tOo/Lj7Pu6m8
DmrFKzWyQHA+TJ4HxsJEhnxTC0aitvWyxtwklSKAlUYJ2AtgbDqpL698fLJutfhV
FFFXw9oTCxKsj1XRJGtbOj0S2ZtZMbEqduhNgRarQlQZ0qfiqM2ECydddAvq8EQW
q20tAHwqvZHJ5BOVsPUlJpm4p+xxsIPFPFQ+ygvjokQtA6rgFe880ZTSkfXNdyOU
U4rbkO1viY9syZWYe0WcsNdmweD8hiGXy/4i/WGHVeD4MlaVOiG8Gsim0ahv5IYn
tKdkfpNtSXkVMpwkgMPGnB5iMYUQrl+8fOWhBx8vpcdMoGBo3yVjJceMXdPg8ZHh
0vYVBCf0caMTuChyv0wiyOAjFaSShbqcNgUaVs+yrUbe31smBnuAGZXDOD2VzCt3
eNkhIBWWnjud9FV52kVAXTTecvB/hgidKBk9qJGwSBDpdbJd6RQJFJor/2yRh8iT
HK9rYRe9gOkIu0+hn+kl/Y7YjCZyWqfU7J1TuMOl60DYB6iI9OIv6PG2ZYoVoWyi
aUpyze1NPqsIyT2v6PLa+enHhjYNLFIJY6YhxD8pLhKYrPK0PXem0qRx1L2FO5dk
Rb4EDgznR2ne3GeuH2Du5SMpavhuNdf1lil9fiWEew7zZW9HT8XzPtzo+0q5qoNu
0yq94KUtZl72WL452SLpyq8S5DU3n5T4vqGa6EuI9UsD0LHZYt9Yv5qceD7CWina
slae2oSpRMb0/pEsWyW4+AHJfRSfoYSgSuiH35bKdJhChneX3DzuiStGKOiHwxEA
IT5D2lz6+vGe9a3NXp0QPPwEDdtPDEt13ITuqkVuLgsq1b5zoZrK6m8RrweJhigD
KT5L9Lk+iundLWUV8EXIbAoJVSxp69e3JFds6hjaj7TRXQXOfaAMkd3QFbNL2Kim
il7IColIZiG/LZ+RlumaXc+wUjo4tRyNXToFSPTLJ0dGMcasfUptBrq1xyNqaTPV
PRwuMUdIrtrydRxhpV+Euqai5zzGborgWDDhDi6uJEL9Zb9Cf34qcRA0mhGFOPro
DUvoNYJOvuY24lDDZqSve5P3zXlujxK2vh1h7JNQwNw=
`protect END_PROTECTED
