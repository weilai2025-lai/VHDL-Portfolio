`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LX202dlDbAaEOZ3Y7UxNqg6eFcZS6CVB9ou84zcRRajSB7B9fy+wsGuOSAvCLzgg
PGGR9CrM2QeRNzEdWbezwsZE0SG4xKjhQzzIMiLl/V3yKx0wlfUZHcSItYszYOHT
gM2IgffTbb1A7SJBoDGlbOKqqh/T7+fueeqK+MFfFmbiX08cEaQAExSsBEMxDoi0
Y9x5bxdR/srhZeJOfE3icult6VwA/GMw24ABqxaSf1eDwWE8g/bYCh2+t/I6jmXv
ssIsq8Fqk1gE3eK2xi877JqUqIQ+kk53YJXa6KAjbzLoOBcAlhaVLzKH53ypCEy0
OemX+85vpKPqKwxudM4e0CWf7nvLfXQcmt+rRzUC+Mw84H3Ij3gk6PPTxv/vdfK0
h4TJ8ySeGbi564Te7ALOcdjb9v/yu3AS6xCIKMbqv35NQGTyR9JfTfK1ANFSeE2F
LD9h0ClsCGPddKo6Op+2kZOQNpbJdynJ3OuY01lv/wh1HBrwRqdU4YRVMnhqKcPN
rFb5tMzLOIGAsIBl7Y58zACs2Ls7E5EXBmtVNEuQaCaLVMTLLeFWGXEKGwaA8txO
JqxsOwgK1EcFHGmJY1RJjuZXkrvDZoo+YcYUUcYsuEYfPmxt+qkVfGnm9AZetl6c
CriIg03JYceI0zubwwbjMvvM0CgBAkqchbZRqAEjKb2GrC+ZOgPIg/tcL8PNHq/Z
EPUBoFJgxB5EkyTrwFM8/oKQ+2Bwz+UBYO+zc16MCWh9QdgvktIqWOKPUI8sn9iT
k7K+TB3fpsUaVOZ22Ny2Mje9Lac27cHYtZore2fV6oeGABM3j2zmwKqKCMuCxmUG
EzYbx/k+c0KNUv8+qciO74VFWliehZwTPkJAl6vrFjXrQbwBOR9iX+sJnerCpKd4
cWSdZaIPAJtEyYa4MlD7NLS771gYNWog+MKTrvISXYxhpa6F85KRlNMoadPTw7SU
d5QFLj7YQWVdA38GpY5cZGP9fv36ulbcGG8tY/bAH+7F+DWPSUB6Qm7JqQlOgrgv
AxlYrRJoozHFRkKkCbQMVjJXJUkogz5coNc7RF1RcL8DJk/fHOFDNhELqOvi5cvN
9CT+tAnnqReSBc6J7uJmYGjOm4w8xKIwX87Kxf9eAf5/0189K0OFCZA9tW7J8d9f
mteKvokB7I9DzN8SYO9hzKyxTiFtC9MpLByeV7QrvgR8TQzRoiaOVYWVUsNeiInf
8gVw2VRNQyecoY7ZKcXrHI0GS/k/Z9/GV90+NeFNjF8R/zbm8hViTxt4f71EiEAt
`protect END_PROTECTED
