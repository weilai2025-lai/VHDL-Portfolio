`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcmlVOzI4CzD6wl6AY+a+PMoadK5yQVID8Hz8rRnj76kRNDD4B2tB4OmgiqzuKkK
wluK3LgZwRL2hVWnMDfD0MWdID+3kRQWrB6YTogUngu/ap5OmD/0mzfHiTKWoiOz
okATMUHps6M8szQCQnpxSpTDR9Q7c36qFSqNJXp7TkaoUbygVz0ja1XvHlN5CcAK
2tFdHkc2Az8Fo1MtOiYyxkHe/9ACR3LBk4eX/j5dCKi7fPxp6C6qERfCUOF0oLIt
/Y42qumwmgvkUF9YFlIT86VkLi9Js2/ANj6/UfKwV6Rc+btkP6Uul0/iKc3F7NKO
sqvoRPOSr/p8xRHeJZP5tJGZQvxhLBpzCOL/krvg51eFFXmuZJEjP5M5UBs+Cfk0
WS5mLzNhkigBqSJ60XbDI/gVMxJWkEH6uJbXGAFDO+KlFfES2z1J4WBByGzhvAnS
JUaqwcvL1wILCKUVOpvODdKiTcLsavU7saomg7c3Z/wVeDKc3hdRZChi47mjhuvy
1aeUTCIAl5DJvBgE6lx6rdJfCozMjwsG3+njqm4CedEXK+XgGBSKHixMy8ElOE/8
tOH81C7edQbWSzQWmAibmUfyZueX5YQOpigmUIb2JLvpifkWSxvcJXpZquSCkuu2
/wG7XVS8cZLQjFeZUxHDv79QOsClCFPiDYGVDDSBdWh78x4sEoe80j2E3tPQYCQn
`protect END_PROTECTED
