`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnK5tpNgQLjmryXPu+QsbG3MCR6cECo8KZJHClm1PmcDNeNKRQUdxApzKHWQGyU9
E7bvB2u617atfx/zbJAGhnG5NnGHo/MH/y1P0TZFhDbiAG/Jbc5pFhbJR4S28gZo
zEvtzs0eFsFDYs5EUtLxDmfWtVjrrwn3xiXLY81dNVVcSLVap64zdX//jqIBINxz
6SAvMss708ou6jbHb6FFCj1fXplGGDppniGP8ceSXfBm7g0gY0P4xSVXYsbUuXDb
/EIo/15+atHSpqyhNaXTviscrcFs2byL3tsH9wJhN1vVOa7rd96Hnaz5XoZFLiFV
Vwcv6wQGkerD/WkkTSBWGP8rok/hqXbpu0UDZ3yPF1Qs2d78u0frR8FqAc09Z8u+
5uDQF+0zT02PkSvf2JU0CyDLvB9J5rhaJ/tdYLJ28a5vLEjGXx4EwCC8S3CZBNE+
pbjfGlgEOFjJrn31gC/tn+89tKGLmJ7FBWvfuAKdycA=
`protect END_PROTECTED
