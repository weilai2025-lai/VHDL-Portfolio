`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUz9U2k/TkStAXN3M5JsBthYD8c/PtkomZz8AHS6+HCB+BEyz5woj2MTs2AHPWaU
lYzoeZll5lCJUqbg+FCawrELYtXC482gkIxWjHQb05X8FxS5D+aESy53cX8gNDGY
XwYFLxEmNxmCngLpBfW6sVVvoLY1ZfzpaBnKZHWWQOhtbgSMewhcABVhYnkkPQ2w
WS3xlgO3dRGnt633e0RN/V7qjLTrg3M1H32z0zVVdrQ5JUXYDasrFrd75HTWG5iz
kRiwYqaezuhVe2SMjeDNlsCRi0isGp7w2ZZKUylbmEiHuitCH229Z7SO+QUxqBQ5
4xFTDgK04xrFBHDKkpYsD4DKNEMyi16sB/gK0oc7gLIKsJp47Mkw2dKdxZNWc/yO
jNDPVU2/WWwfK9Ijf+3POSnWHyYjF/tuBLbEfjVrhuvuXV2aBKz5+92H1k73ABlj
YWXl7iHhgZG1wF54DNHKxACbVbNs+h52E4ejynEmHt28xdqUcReOAfN2DcouL1iM
U7ncm/GA43MxMDBo9pApiPmR7tcZwNAwKgCMz7P+XY/xcnyh0RlKS2vVCEsIkVfw
7sIJT1mjPnruAGhJLcmolfzTTUxYQTSdRS94+wtmKucWVpRtt97dBoEHwy9Czcqc
DFPfp4tfl3TVA/sdqc/FiKEo5Czh6Z61OHqFAQaqlKy/RZI68nz0nS+3KM/CsRSY
wbbmHdCsc8zUHumwmsuNgvYCMnAG0i5eb7GDtMweMUUw++HAfWi7Fd6aYQqlYXXt
8fFbsOjCRVuawgGO4JFM+jiF3KLzxrIg1XxvcXYQeCJaY/BuEui0iz/Q21LF+0/m
TTlLp3bdWdhP5KOnhhuJ4hZc5koABYQwVapPuzjef6hf2fGTpOAFvc8teqjbAIfH
RkXCUdXe8NeeosK1StWQZDyL6cnAiEx1ojk+SX7TQ/NjSDoDhdnmQwbtXLyiDdIz
MwtPzvzw3/gizdY9+zPkK8jIc832cYdi/ISpmr4hF6XqoUCP6V6wyhFo+so+ilLv
DucDg0uyYyGZY6yEO4eEWU5pRmynOGnAhyCequcKIHKjQnqSRErLO0Dmps7sw4Gt
UD3Id4HUFHWa7gW+J7DbTRTsL4DKfy9RORE3oV6m7hlMX35QOLFOoE9lR4zB4gtY
ybL6dUOcQrRIGXBEIwZZG4TW+fBFQZb/3Wo5T3CvAEzrgus8ksaXv3u6EemRXCf9
Pu7OaVha/7pEEHkuv7h+Dfz414OJXhCVT+3tAXDf5znrkLoRUYO7VrhWF+t4pAZw
axXyz1lC4vdUwnQhNeOr/sGMx+jMZIoAq4pp1Mrx9OoS6vZmWXe7mtc6tQnplg86
qgTgAQYZ+2ggrw7/mXSr3nyQKY+5Pgx99VK7s2AKDo5oQWxixsukrqyti4M5DCzb
e6h/iWZxC5BbwyQbdv+uzZUbLhIgHboI49Q3zc8ZqUvErXA9/miRY8ZNlV289D0z
9GkEILm3qHrBHd/tEKnOBQ==
`protect END_PROTECTED
