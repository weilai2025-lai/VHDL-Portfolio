`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSDxCpfBZzWRUC+aHJPJJvlHhZ6z3GFmq5PKXUygmHynUuTNE/oYX//ZfulKUOc/
a4HlNgjBqZTV5rhSeBp1xccYtacLyeW5ZW8060rP6A0uxWVSuJRTw0RxQjRlPSQx
jSkPSD6UKZWbnLMMRlkhoMxAv9+tF6bg5/xIOw1xnGHVzj2slRhF3LNmeVvoipek
xFtZAYnXsVLkf/S6Qg6mx5SSuUsOB9Uj3cH1b0hF5Fyf9rjvM1RXcaScLOaHxSdf
2NDTNG9wXyq/Qaw6m0VgS6oV6NHW9Xw9lejXyVrzxH9SJAj7y5zT+4yVWcF3B9zk
R0oNA0EQKHbgoIDpn5h0yzkrRllekVQSYk2uhx3soYsQxkd6RnF9lKN5Pwr8is3a
uW+6YPurE/TThGHQxT65MPMr7WzFzKQ6EopeE8Mciirr7YOnIr6F90pSapmrfwUC
AHOXz2S2i6fcBI/YlBlJZRQRkWkp3mwvRoRR+VWor+eO2zEKVIHxSpPYbzJMXFEu
nt94lqYFPf7HMBHCx8Dj0MpjzwKdFpSl8XDY4tA4JIV9yUEggTu6AdHHJI5ynCjP
s5XEOhxujWu93PX+QhyQsQ7+f/vi+IteB3xwod0EfVqA7P3PgPDwzgV0Jkn2DQX6
LVLYg+G2hcap6FDU6yHqsdxe4lgobXW/Y1UsfAas2InC5piI+eOBq3Uyt/JA8PHm
zp0eQj9kxC98oMUEb7hloQUuiZWf47ttfn5MMfYkuf7QTIswHe8nsbCrWSEGdd1r
bM4SfEDHqpPDgOgYfoVud1Ot0RYNBu5EpeOmX2NEWHFHvbc2Bf1HcHsrrcyz4v3r
xd5FkhVpCiF/YdDlRdHvVGrBHdeFRuKHaXjKfNU/XWCfiKGWrbOyZtB+o6Av8aTD
+QozMr9ZhBonGVbw3xD0vy/Ab68/QjNgYxzP7xwsni86rkjujKNVmTpwQ+gRK5BC
F+65gMjx4DbgzbhAjTliDwwA9dXn35SWxJGOk9yBuvcMyNCESoI7cUPBziim5Upd
wE7urkN6gDjgDojR2ny/2k3foHgpkhmvq/RUvAHS5QJQaxFnT+wVzwoR/5FcB2ML
OqBJvWruyUaJRh6FBnjdsrayY2VQSPJ6jKI3q+2kL1rsm8K+2X4+MCgRu29GEz+R
d+w8BkCO610eypOYCX125TuXN0C/t+38xzTI3e0qFpC84PC1l979os5PX15m8WUy
fBkhzRxulanEBHXCXeqbma5SMEoJtkFYLc4cJdeyDMuwVA43rugmEuK5IiYpVcpw
rdGF6c2qkXLBvUm+67pND7Ok0YXCJNUXsPJ42277LskrQTVSHpxeRAc3f/A9KFGT
aKK3hoOuiRdmNostm4k+NaAovWx6RVR2ZQVVE13YuPCY+sYCcdhtWcszWe/36Dfq
Q5672YSBAd3ewqBv1x1uDN/yphNWEWPX7wHiv7zDSR96jgFk8XvC4Tx4tloFeyA1
r4+LGChRnHakvjviQCRK2VetOn4s11D3/Xk/KZspClZjINqR0ZFEvpQr5KCxFGbY
5EtOYVbci2lhPxsCCKcV5KcNN6yUBqv+aq+ZmD2pc2n37XZvnpCDAKUvEPVE+rdi
HoFd/zfpY2lcVAq3USjHr1zM0aDkMoII7JOTZB1/L/94ZS/U3p0TvA2uHjYJ+GQK
sBkiXIawFrR0lfasBm7+RxwjfsOLQUcNKh0LXWRyddzen/It8kudijAlrIz1WlC/
plLAQtAbBH6zdMNrdF0suabNMmBWgE+q0D28M+MM9BKpIOkHPfCLnqs8U3E9BbTY
ofpmE4ND5vGu0pXH2SCu1hQxITBLtuefEgLCZhihF1xqv/R7SuTc0kUeS7nkPFwC
Vw6G2y/iqy4wtq3ugtRFvxaBtlvR3/wC3DGQ2MBJWVQWAD2cIsQWxqzS9VSN2eqt
a+K1lKfEOTskyKrUX29rHqJ7sINIcMotIE2o1sw7a1NGkn8c/7JzKyOarU6DNDh9
QRUOz167bNUJW6+SQxVikgTmO88R7PT31pGkaahDCkw9RS+sSXNaHXx1nl51zz6+
OGBb1ag9f+l+5erv25h8VWPvXrZYYdsAXJi8ZB+zqvDFJowmiLij2gEqrT22qixk
7aFQqexpNsgRFOsZslIx3Dd7CcDJNOkaZXcCF7Zvt/q6bO4zVbkq3YZZEiNfFFY3
2LoshurCr9HRrrHLSPuBeOyO228EqD12gZaioSIaZdOGBTPVdUVLtBKVRuviyO1N
JQs/bIkX3L3CH+u23gFIuSMxezx17q5YhOqfFLwM5G2bubqU9AmoXpvbIw8vGj4M
GfcOFFD+s2qsxnPJYmvhkF55I15+Fsqgg7mAyGATfW2lYaRXnIcsM+tCaJoSaNvR
kwZdMeRN38H0pqXTZaQsnZWLM0XjEFeJ78OJX6sRdgl4LDNes0ORpbQ5IBxdKybX
r4d38B8aVoVf2pNIOXykPiLdy5sZq9Wyd81XdxgpvNTS4HWENDqmvYJBqZD2Ya2Q
I9CQ+Es6A49cpwdSXYw+03HUiwNZ8AXZGi5nuFUbmPzxJiNHAUHBOBpdTm4oAijg
ziKOYjpZSfHYwsPX6mv/0b+E9mDAvOFu4LBfntYDgvfKI+bz9xsE3bdCUvgvSBrh
U+WyIDUWxGmlK+n00r/7ZgHzegqztw79mUbYaUpGmvsGZMYvOd2PzS9AfjsUC6LU
izlnSsIE0DOSTuRo8fQa+g==
`protect END_PROTECTED
