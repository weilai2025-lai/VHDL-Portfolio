`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U91bDiyJ1z0Uv2tswB9Q+D3Fp42Ac7lHDDwM2am46F/t1IQc5JKLFscFDlTf8H9U
sbULPanJMPALGkYc5eGXx7NjoAaJF742Fcz+kPV4YL8NkeHmNXdRqxKAYMg8vsuQ
hyYHwlzV6y2wJhucJrTkAYC/VT7ZAMeEH1qELESdYp1oI6CRhIoQpfe9FaJa2qqd
0LqDxE2eVUP240ts7+MT1zN22X59RzOPVXp79Em0V5h1a2lWmb2soQUU10zFrvjH
aZ1iMAAWxNjknNMgz58BlNRGyxHrmGKgZ65RPO7pilq1mo9FwzV9AZAQXFADmyfu
Klvsxnq0bPqWAsIktKLwYaMCY59Hsx427KYfIbgq7HMjMGUK7cp3MCTRR8bTXi32
QkWduy4Fc3nBByvU+fqh2CFdc4zgSsdavnY/lcivVEsDpGQiBt4oRKWFs3HtTkso
pKEJpzU0K8V2gi4f7+b9wgJIwDMoaMZEgTSELf7svlRkELggCHGiFVzEWjsqI1Kc
tBYEmtzLqBWiFlCUX7RbwtKv+4rFZqN+8SWETNjTskVLej/pp5AawV3hj/t4RvJD
EtfbhwavUVCnHY/yqM28rohlh0XYumd831EEcvO4uY3XzE6JM18fykXZYOO3UUd4
3RHfI0GiIY3PEGbXC3YTVmBCkjCD71OiGRR4t550AVvrHUfuOqc1OoI7zI1rIi/z
yYaTPQOhILpGR53phx2/zBkih/mo4IaexlbfalXkSs4cf5EEa05AhTKaGsqurn8v
prjj/gw1249wEIy0NZeB0m1FwYhxl24X7yumdA3pIfdjJ5/iJ9EaK1PuyPBIuFuR
9T+OKJcsvpCb/CjC5TgHY6GXiuPXZE/FpcDdZRq0FPNqK+4oD+wQDaCswHbBwgGn
f4df9g4wPXW7zpB/Vck140KsTeEWqRH4mh94EnhbEbuhArDU1w/vmNEnL7UxcPIq
MiQb6X845S8I2c0Eoxn2z3bb6HJsIs4GXIQxdgguV3Q7PhY/AoDPcLGUqWskfV/u
Qjn28WeIuJOpIngQPcLpzPno2NKjftvCMZTH8I2YpnvRpwxy+z3GwTknWYpNx6Fk
FkkBvhyQz4OTwsGvwij9eumgBWEXTlT38raPwLDqzSB8oRc9EnzKCehgma2PgoAa
Bw8AVo7XuphplT8zf7IHzDuCR2bKECbCbXD4VFVdcwdp9o+cxzKnf/QuAqvk76DK
M4TZThiGuoaR28j5da/+1s0oj9Ersa+J52NIQ0eoT/vLk+bqOlSu2zz8PQdGgrZf
Yc2zdbVGNNu3vdnxPipuufftu+Hp7INMriCSpZY6bUER/N81vOQd9UU8wFE/GEHH
Y8NB45RVY97RlgMNX5FxI7AEnjpEjGw3926jLLXD4bvQuKwbY6qVgdhfO4H1qDqz
v+kgupnyISCgdG5Z36hAC/GqbEsikNGrf23uplMUYqkzQfwo4SqmWo5NLgq1igfb
AmDE+LhYbFx+9rrl1Ga/7CgJLWibjMEeG3UD06js8bE=
`protect END_PROTECTED
