`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zdpk90yvs5e5gtlpxw96LXBfX3HfK0mQXv+rNUgvWq50mEmCZaiBA7LzbgSSAwq
s51/Ba+HvfLEthAHujZzU5OGtIZMwjittugNeDed9O2deqlx/6tbmZrWA+kHOBTN
oTQy9pufn3Uf6EJVF+h6fw0ElxMRlXdd3MTTd1l8gOYa28Fj9kyWNtMSDZqYXEC1
TjMUpyWlCfERPcv4kKnseXdBI/1yz6PODoOl1iYm+g6wew5Y9Yk2jEPpVUcDr9mc
nX/QndXaqvy7tDGFjsxMHJ6bPLcK3NhJipfu5htlTbZ+LfremZsFmuD/QN4k5k+0
nAPgXSUAY+Rcnevfxp6ma004kEY559uYLFMmrPyo8bLvovSOoF9UHTFMsKggnRzD
cqsCANyQN3qJU79exUibyjRs/SCOgIkR/CN0jS0cI6TK4RgdnegZgyloTsBgC8oC
vgfYYsAWgWQhbl/oBSkPXj9D5doen8PNguG3x9DPYFgffA5pqdspRGcCuFev9HCl
9yWX0XmozJnY1u1HM18PUULXYfkAtOahoECbIwrABhYRWuGvf8UhMUBJnzF4//+p
cMLdXlsm9SBZsltBZOB1CJ4lFk+FFKk93+Wjb60lMhmF5gW3H45DcpVL1cUpaCMy
GDLubG40pdvw8V1w4/NHLdobatu5SHynaGDTomHfj31gVYNSw83LNvu6l/UXKp7Q
5g51Pu65kRnhxPb0eM6wxMOuwmPTjoT+A0etuC+OMF+eJQ69JyIS51QVnGI1HJ3c
4IUWSiHSe+RikwBPrSD9h9udfLquc4JxwQ2OTYkx3cIpBfvCJp3MbirXLrkW9Dpx
EP9vmH2tWG2Htujiu5fzH/StWik8OcTgpZi4TXXJi9kqkOuhR+QbCrm7p2rzLpaV
QYkA3hy655dKKAFlq6UMqL4OOeGWhQI+XjyY3HiQMZNWSFB0O8KEXhiuqqSxhucP
/8hhhl8fKt2yH8honPlV++UEHkIA/C9i+9XhxaX5Qo8B9RaKwqZkyyfPFIOYdWyq
y5X417K2MVO/8qO4T/MKQRQg8+5didj64o4WqStl9nehqBC0Q01YZ+o6zld355ZW
YBulvqEp1FueL7RNfiY8VQAxf7dtNv6patP3MSRQwaPR5X6MSEpEaEDA3SCSTbA9
TKXS9hWUidKP8RisO/EyQkVsbp40n1DCOGwuzt7RhMFxyRyfwq/PtR78172ridvX
K6cRrHW2APfIy/2C5ZwGSYQ9v3Od6a1HAct61vfblbEfYEvXYImAsdH93FWOV/zl
JsylpXQJClVQanTdx6JHfgmQeSgvSlEDuwGD2e+5jMJtow5NC4/OtXMsjDKBoWrK
s+GcmhUGzeMhE8SbnEP/8g==
`protect END_PROTECTED
