`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nB4z3iursnhXXica0jsfXpE3pO3f3dIg58r6/v3XPW9bUdhacZ36YYrNHN//m1+m
6JqC9892KPUDztZQjBQzq/q3KUuAkYHL4/iXW5LrFZIkqkJQq+JFTuqdgQC0viZF
f4vfrTz9vTtFopu2XesU9N4CiTS499kJ5576pyz7TV/2kv8YCY70RlsDm0VSoJaz
pETdj/maD/iCG+X7i6y2RxH6pF0URUJvb57hjZkoxzdYWLOqmpffTENgWhJR0XFp
vYCK5bRe5wvG99UJLcplmtoQGVNj+cRxZsLtsFWECOcgSO7GBqDulD5dPt5HuwbN
3xkG/SDWoUL4Jn6iLQsFG4BSmzmpWTe7hxSp+25hCWZ04lI9e/ZptIrHisKS7zAO
3iUpFxBWLQ6UV4G4eysMZFc+qsAT/VpxbbLUol016Z+HBiv/kWKUvmIGHySBFyEh
RmVshr+Tcl6KHQUv3KpO6chaJ43LQWI62mNhdPQfn/O0d0AA6UTy3UD/F4d13RsA
BBJ7OHJJB+ECUCNXW5sx/vrrfCbgwyElVThWvwlxpLmIejYExGwPiS9Z9jZC2W15
sEwpWFsY3bAsDIFZ0Myi10C7XEUblBnvXyI7Zog2oMM3y79iWMiZBMTHl52v08GI
i2tTZd6KKdSisD0uvBVXF+iaxjVBjOV+yVzCy0qHih7eO1j6YPR7PjLDOO67reCh
/mdVImdEyBpULcRDx664z+8uII8GTk5e3Fag/O70O3+GUkg16hvdBoaZXH1eA2xZ
1/8zZjhhX+rTRwU6USveWNwyDI6aPjNFzVYyazEu7hdp+2cTLrLN7SouStzJ3frq
gdHiTZyi+cd6DcRbqK/bsCTnEMtqElBAEZW9SdnAI1B6T8cs1C4eKi9uMGM+LzNa
Kn0q1UBVk8Y9MvRE2+dFTgvwUUYtVa+vbHavA/lKTszzXGK4taDJKwV08jyK5q9Q
JmKS58zk9kfQvveU+QsbHnHnb+RPF4mvLkA8uMWOWaaGHpvB1UmS8Q1Mv+8P9th4
yKedYuzy3hTjCH22j/wEnf/7F5vLZBVHl29+cNw9xT1mP2kr8LY9/haFr1MZcZlX
JXkRSXWsBIHKqwlmqJ+78btXf5PwHuSwrDEEcYGfU/Zm7EdjFzMel4j1LaGgmT+u
3HZBOvwRA5RhzWp1fIkZjVfTH0Ow+gyV3zXpx1Nuvd5M/ltRE5/NPjRXiIHO9fHM
CQu087QeqJO8zmAWn70Kr+jFxOSuAqEs47mXUq9JVtGVdfm6XTLZWXYLhPRYmzwq
N8S7mCPjm42FIvcYKoxqR+XG/z9WTll7hjNm4/xTaSOGcp5TxGpSOio9VehukXZ8
F7q/YzohBg/kUIYhNHo97nFhstG1TdjbqlDP3jWmI+/enriB7itFQ4jvh/CFF9mU
d+1zEbllKRlbhv2cN+USMJzUCayLo7mvXS23Sqk6ynhKFAN7GmjIEUY69LqowLnJ
6c0v4ucGGmReR/GgyHQ26eSh3+7Rwhxujtvt14KSVHqbol/yePnqtWdKbXDn2gz+
7hX9+1ot0kmTihAuEoOldy2jVF78BfoD58nHlN3GDZrJPYad7MAsm7agz+lFQ6yB
IStofd0JDRmw79r75aQwufAwswGz/yfV2S/eotTGQNMVqGJ/xVwfMzMLbCJseO84
eFR/9PR+wDmMR28SqKZKAz+t5hqq43GkWVGBu3FBA7d7uJk82FTv9f6ObABAdgK+
A9YRWS9ydIe/MCaF6U8cB0XORNid9+xCW8Vkwlnt1O6c8o2nvaeyuON1BDdZR377
mgBOeb4Wfam1EJW6zSfsCAFWoArj90RPHEAH9WMYf+SRUoMiNtGidKZbcUCWHqyT
eXVBMp8pTUzrkzhFQnf4aiGw0ZC2/Y91qYPp+ZcAOXQCMqsfrlGUTHMV+XvQQ3CP
yyT2gon6Bqgj9tF1D3CBOyEeyCQAZPM+xu5lUoGlfzSYkFfrPkJ7ecrPLrw3D5QB
Of+D/jKA49ye4CBfiGQ6Ohj69BSOZNFQQq2EbJG6UtUjldqMNZpcX6NPvT7hcAhu
5xyuPs8hBXbXZnYLFDSGwsVKefZEhtLHIYVwBIZm+rADHYJJ0+ud7EZOLjNSVfsp
olVLu7dRJVL0E1y6vv+SiRPcgBrbVW+1vjLNIcO/14Fnq2dT5QhxQeEr9IG83gyO
l5LoXi9Jw/ELytzNVUxy+TXQt2IKgouHY5QCyV2DlF5Wu6Aesn4m/4Iz1+8GJco5
YhL8TdRsHK+6qVPxIX7J0CW2M3f9Wwuffy0SoVn2f38pcd/51hBECEH+kcz/n0YJ
GMNHahaFI5qQ3Mm7/hwfh17l1WPZgupMpkOgRDi0NgWuDGVH3HDDMPjmaC8vkyhZ
RXAntSrp8PL8vfzM03m55P+a9isezZFLDFI4wkFLead6PHB1CWPFtEXzSIQ7b5Qd
nrNCm5t3iB000ld7+p/bansSTYZYUK9VmmYANL+gpmFmh/6Z3OxxbN8klzixK19K
X83+nX+QmpU4chTj5VSVIyZGywpP3kb/XBneEG46vGBApcSbVyLQpA6jotewo36D
YAUxXnM9/6UOv80yF7LGSBlagjt4WT1XWoKG07yT8cAWgwRc4gEtjDrvkTHLvDm9
ZF+zudiyXpsBTBgjLXb6o73zEA/b8vY+OmMd/ahdChIjY07VjaFI0dDw1ApruKQU
agIkhNceWRC2/mHMFlsK8Lz97DIJmarGSq1aVPKLXuCgTTG6/S5aDfK+cEmff5Tj
qmrumXOxlBpa14ZnDUbyADkmjh+bO6+onGjkS+ZDNWfP5tFLeQxlWIGHs/1Npb8d
Qzs+7r1A7yLBY/DqA/d7SZ60eZ9OMKoJSlOLbaPtd7Z5Ni77+uINxcL8rHc7kihM
IxYoQmbUevWZcRY/ypYD1eCrHUPHJ7JEBnIrskggCweVW7SvOVKUbsI2D2tBeYH1
+aCqTqd63P9Ic+U4++Znq/I9jMKQo3jARN0+Eo7fSj+J2M6rFU+FD9K6ZmTnjjmK
G8MmNY3jEi2Cg52kdQyxQNfLOrNCVe3IcUshH6kN1nP/VRwGq0tHb7CUCZoODEPp
2THUihpYrd2g+CRGNTqiO9x+aeSkrvw92KeNcAyrrKlm0xcj4Cw5nE3W1/DB31WC
49jbIEoxseNRD6o9uV4bflfv4CVjwQSuEQSFwACOzCK8JwXdrEJA80tTSNCNNCHu
Gs8zY1RGV5UgKfDZfsYuTxOzlrm6cQO04nIA3KhZTMAaG3tanWMzeMkMn74bMrtq
SF2ELbxyph4w7ryxI2lfqdKzMgdvGWha+Sf1EvUG/MWbtlVuoJ0K7frszGjgg48n
9NF1u37dHypYi2R6/sz79+zEn6lmtW9/ManSIjhA7hdNl2gr7uaf0F4f385tUiRq
HK7NfiGTLXWAlOKmQnIzhk+NaMczPxYnF9zqMUO54IOs0uYqRpaEMJMpGhvs1ZXF
JjDIpws2TtO3UGQo1hL/a/AJ9VLRV3rIgU/pDSq90LJ/hAvkOt0yJSh0m8U/hWUq
F61cjaWoaLNlZyWdU4hyGeht2UJEtJh4ZZg5SfeXp90VCe8S+zixeuxI2h2yR41W
aWJbqDhoB9y8x/BBZadhEKykuubN4lqX2rP2i07KDzKAYvxZXKcJCkrHtePNXnO0
9rmF2plnHfbCMHL+rgjTUOV0C0NYTSpeoBAIxXrff3Qto3mfucPz6Ven3O+bN4cd
w5lqxxsWqmvn0VrnL5wtmMIC/aL9OSVbxHz+hvrea888h8ZGOYE/WBaKclOT7CWo
wXR05KbYa5CAtsee/OEnwX6U/nffQzmzIYPZe+keZyE/FJv0a1E05eJS41Cccg91
iMLm2DDJXzVGqyG/3+lB8Xit9lsBr+FxOY8bDrxzypgOKEqnWGDk7ObLTiU/0WA1
2Szmkg0K8rw7DOhwOY6PgkWhEe5f55Ykawi3nu5NFHtmBCSvuVfCV7SSYZsoeXOu
bC00C/BlGRutlGT8HR6CV7D7NePgzisqpvDf+GrUaZwDQCKghhUktv0/SkaVHVrF
9knq3RqNh2ApxTypLP0X4udu7OcZbCfc0R4tcmQ6uhU9UjJ7bvZiO61KI3TbrTlX
EQSkqjKDAmqeaamjLIXN7mWGqsYjxM00XGYygPF/A8ANefTQIvjMqb/HvbDLiTxw
PBZ85Vv0p77XkJ1YDYoi33sbyBXPbBZyxmljTrc/motArSrW+P9qskG57LROUBlH
SfHEsyzY7cDFMRUdUgBKSPowFt5kPotYe5UHbUFLiuuUku2TPU9ZQsEKz3ZPv4cp
oET6ybkmHarMSHlHWMOOGDcJ6iJVtj074fA3wfvB5MlS0EeHZtkoqgoc/kpfwIZ/
i3AxvQNNGlOTgIOV2s406RBAYTrgB3boUMVsbor/HfBIvKxLAupq3aSAWX2cqJmh
TdQJg+u4fob75yOzfQwGuxWlZPbXDTkn71G5rgog0JR1pX01ZEb5bfxtAkQu9C1H
1NMJpqj4l0gBDIWKCGeQhdRqaXusiZw7FjseTy/wlOjQHA3ovfQeGnZ5ur803kq4
fC1U/pj/d6IwKPRX/1M7LEd81OO7voTRsaJYduUcAtWyL8XD3864ylgfFwTdsMiC
fu/epi6iyYqXePQpsXBwSOCUxKycjecc20N/CLSdWfi8ReL+tlg0w5FtMD+y4eDU
o+VB5okBAxriHfMzOOlFMU1532+9/IuQaMBRgvaj7UwMtxsxhEiX50+c4hYJbPnM
UL2XR1kYQkj7pkNnIJGPT+573SwYwOzx+BMYOskZl4/LkK2xwkPQEvOZZlARC+UA
wUakb+H9tRCOyY295uQVdgoD8EiL+NB8/Ed992KlujdgDsKUNFeJ0zI85KD2vhWL
gMyd9rtHf8VtK2KG8xYLsFBTVzHozydiVYPwRtbMtH33AocpxjUkThmkODw6Dtdi
AvzANcVzb6rr+vATPV93C3lePuysESOAIgpqwygKT5/7srsSi3wvy3GJfS6Y5buU
AzoiCgiaRl+sh8/JC3v71ZyVRT0NLRew+HKVOlofKlZEOaKLjJr64F5LGsiE4Qzk
2/V1GmVpoV4J6pm6WjF08zFMnMQ1TCouvQqUK6vspNUs3uTRzaIpKj/mJPs22hJh
4A5kJp7zJp4xWJZkBxjihRsc8T4oi4bvIFR6pq+lrZvcF2yGtURWcFEBAa8MFmVH
LOigYCr2KEp3s14BxguV8zZePrNZsT3Pqk6fHA+d4VY58lHl91AvMQWa8GkagAdG
zrgTvOi1t4ekg+h0kRrxN5RwE8zNg7e5ehrIh4RKVxhWMlxFH8k1BXYwrjXxRWHj
8uD29R/wTsh11G+Q+03nEQCj6qGSg07BO/oiDgvGlWIOIDRy7SNE3rJ8on2Qc3r7
g3q63qtj6GFb/3S/K0Wk4bLBMQbUBlLuJebFHOQX+heiG5IR9gBRBwLt/m1pGGdL
8AHVdc98bs4cyccOJha12Zulz0RyXtcT1hbDTfPGZv06+U+4vVDAB68N9WxRFs06
KQPUXoPXdJhxWkRqfiergzyEbki6hSJneZwEYpthkcwS1fIBNzbITVq4gDefkGHd
EfjkUWljpbmTA3mL1i14kMA23u48G9NHdeXgpo7Csq24AkXe14/bC2C+LXKwvHEs
gnZ7glxqIt4KCfgdI6J2K0MUAzqReftaxgGMsDkttgrHnsrdvY+im4RUS3htUm0s
p7WG+lUWwuSFynmWw50gJe2wEHyNrGrMcMp6ty5WoZ+ovhFV8kzEK5Isvfc1KVRd
UPGT0gqNz38ILOjpz1Hb1E/oNyQDMXCKaNEES+4ulnXxIOT/BwHOlXT+Hd2PO9Rb
WMLr3xZPWDYdtiTXg4EhPSPJ2CJ5pk0LE1ViqMUO7iPZUtvVFGSyR55iTxk/ElUG
FrusAGlTZMfwqMzkHp6W9KGck1i/QfHZy8ws+fB+cqWkUeu1h6epbJizjLH08uZj
v+USnM9wwRQqjHuIYBHC0Pooc0xIhmL9dIiIBIgwsXGnTO1KxcK5rDvUSgdn4bXo
PHu1l9KYjhK6Y9Y6m7c1JphNjgRy0VRp2RGqSpbxgaE2leWYK+Hor9h4DT/I1SQx
Y68XkhAV/ZAc/UCndKApNziDt+ieccK3jbdluTPl58fGJDkpYbCHmhJEWerjX4ln
3Uef86chrS+cBWgU2hDbCGt4+65B3gO0JQMK8rWTpruATk7ySNqjGFZHC5nXgsrK
OROEOLfJSGKySQVloROoIM/9mzBe+LMPd2SaikSqjsnoKLA07bwtOs25NaukifjX
AuH2w5J4TyJ6jaWdY1f9N8Lte+Zm12iIdYRJsyLe4UTPAb25d/xQGDGj8E2OvXfH
218bZOMzxnNIqiLc1TbsSKkS6baVEGKPcYadQvNmQACr61i2lMT6cQqdwgqQtU6F
GgIkI/xZ3zIz6EJ93WUqDfHeHS4mpWYoYsrfavaR6uFOexxh2DIkDx7Mr+ZHZuRg
uVXRdcnZWZZEPLkgJCvtQQWzR7HthTaJ99RtYv7r08koaEjmOuqJhr3wTpR/BZOh
LHD3n1fzZ7fFgvKZrbDNNcEdNlnE2C6f5wCC8DOiiCNs8Xn1KTyZgZROhwaIMGCp
VU8LAnN+8O6FPe9uLp8/XXrwsbJuvh4NaQGN3/fhAaaToLVAUmY2hFiWieKvA+je
1b90cBqlssx+1pmceVATT65cr3d+eBb8jVymgIr7GHa/Pf/RFRsLzVN6P/DBScXg
6nVpeBG4NUhgDwtpWl1cB44qftbFNuZi73JMmM6rp4kdCn8DIwWlqRSIef8rS3Zs
M+nTKMPpyJVM4eMnHomX7YcYg6FlK8ZhN2qQEyC48Rh+SuH6tU6WVgSCPZOO9Hz5
RnLP3QggV5cbA4Cqy0OA52OHk4VQWECg+fNOODg3SZI+NbaX9N6TeZlzqVgOlXK+
kFiyXW5IW/GyeqpUfwo9scYrYn0KN1/hvIb/qTbahFUq8DlEqyy+yK22Fs+Rsy72
kCPYlDFjfktio+TLV80fF+zfTtC38y+eBfesSPxncpzgHhy+4Z7iS2N/6wUJejkF
wEB6odxuasaqcv615R5CCbCoU+b+Q5U0WYBpWUl1HpSat3Y+s2Rxcs0bPsF1nKlx
AVRUTclERF/AO5hKL1Gm2H9k9YrsR6EBx37fWgUjduThcs8LeQs0Vkl3R91hrvx7
+Iow0bU06vcnqCnu3DU+C5HfQF6/vcHqnJ32Y6QANTIph44y/vX/d5gdRAELT31K
LmDzmkOsc0iEv9rwhG6K5glPsJjnk5HIPxqU4No+BWjxENLJfxvR+WtjYc/UwrA3
MgRSzObkFNkGxy3PUpuwZJPs9zf2bne6TnKntEuCZSJWkBMQi0f1TDT+/enl/wJl
+t+tdlPLyHDuJvBBuo6e32hhKc4+jxw4e6UxTtPFEHfhhsDCmOvb4/8B4YI0oYbA
BAqTSMoAj+LwIRH7slF9sUQ3OfAwmZp5am7T36VfyAdQfoGxohPHnJ4v7IVxe9pn
qp5H7yGlbfyt/jw2qFADXHy91E8eRJQaXNq4eOoo/i5Emtf7EdRhJ5o0b/UYgo2s
+4O2yWvoS6W+aYG2JNun+Lbdy/mKwUZQ08T67uRVSORD0ipOShXk1G2E3CCQl8xG
Gb4Uy+wJyp9YNAzZ0EEMVDmaphXKLuevfKHp50OOYIM4V/4Ch9M164qXd2MWc6sS
Te4mqz3XQuDYUlTIXnWSdGGjLsA+vpbPWO4eOIdO62x3hxEpkkGfrnoih4YLeP4N
0dD+ks9b3lbWWYZC+oKDtcssiF+9Ur0S3w0d8G424zbMmmwWWvXIb1xzxbVwutws
zUzjyrlf3RUKPVEo7NRFNfBhWXv7t9UmtoZoNQkzhUFjMr9pKwYtgumU3pXOvwpm
XGshpQp6J4wBwPHQkApK7qHaMlUsVVLhm1t++xePseVRjhDt6IMNdEqPGn1h+5JB
sjz7jB6eIKJUxeVXsfM8NYno+PDa60vqo7ioq2nFXjAhT7L6039+2WJ2gtUcbPd2
NWYRzU7USAkuDw1YWLGhLuws5tHjmHbmakj5xe9hqu4UAFFi+0Yu7tyguuFSDT8t
xJeF+Ki93kaknImJ22VcIllfeyWT78lFDntffxYI4FyyVueUWGfKDdIiyQXj2eqK
VGCrUCSghkc363KGMmTC9lFCTam4kUn62RjIs/OldQ4c3aEGF7+WxpJBTAhsr5n+
eoOPDsNApEM9cJUH/xnEucmxW+OgYyEYnD3h0rwcsWTwx/Ji10FOCFLY0jJ/OqnB
5kPHN0fk9jqKquulPptnpIlymB0Ovr5LzfCyqebjIeVaTsRUCTdbOUZBAbFhuCHl
XeXn/N3Oq10VA9RdLdM53Y05n9rnFF5Lvo/wKrtedD3QsKuFIVu9tW3QgYD2XMm7
5H2xPD8kqSbhMOxiulxkz12YWByUpKa6CaMX6vJABlGiyCzNuWuhA+jpXBO+FdGP
Nhk8pfMMk1SwNnTiKYsSy1snpWrUnH1rSAoeDirgDJDSzGsIsaY7kgDjB2BRkbzn
UAvUTbw5lgbt+0G0m8MLws6k3+inFwLOA1NsWrafzVw7gc/ae8hIRaOHrQsCE9yl
rjuj3Po2kGl6Jl/W6HN02Ywkg21rxbqkEV93rwopKA9AHd/4/uMYdhN30C1Fw9ST
H/q2VOW9bHSRxD4O4oSpFtA6jHADTbqQ8pM7qWkJgDT1bCV56gptZAxzAvP8ie99
sEFolV8bDynsbYzrVHtcKfsRCPh4T9X/39Z9mHzIIUd2Wzbv0Uug4sQVe0oERk/b
jc2OoXcd+ShZ1Pe5h7mZqu5i5N2H4C5ohawPJ/C/JcCirNfhNQJYYXAqurSM33Kx
+lk5wiOkT7jFfHVbQs48zLG56kh0mB8uykPuJnBssgKV6WZDgWsUdDzLQ08UZldT
SSpWZ8iDOwU/96ABqy51Ofsb93KLUtse+YbZYIfTWy1q9SyU6DBqasUC+oQo4rhZ
tjlmMNsV5VaVZwURvtVvurySAk5LRYtaTSPzIkkDy4RZqS3Q0CSFyJ/zB7lbmXUn
PzMmPGnCQVO6lT2cAkgggqbQtH0aXfujkh+yQwlrS9MV5w0ITO24SragFc3+ROp3
iwpw+mPMm4oKVE180Uk6Gzh2QDKZi/wvbS4T3M08cK4sBB2NS9jH3fB4eIe4XrgV
17cpPwR47TrVSKlulAKv7R3XS+s9QVegpFsEXII8KUOcTJIvl2M49m2x2P9PYCIJ
W/1zirWeFjUMOBQsPcI4JOax9xObj5Vq4l5eWk8VM8VZmWts5q0iaFDUm9uxML2p
cs/P2rJarDUPNxuOiLvkEv7UW4s5Yt3QRWGP3FvSof8QeZhiPrkLdtTo8+Ij4CwP
1xfuzAdJoA4Ee7O+putCxF5s5oxa/oLTqIpsHTmRAyml/ps0H1u4Vy8ViIYy7kFg
1yNpMjyT3j6OJC4zsXrTcTVmngn/xbvqyCGqA/JOLuz27b8OmEcw7+PXAJFfwcfd
CCNMU1kkDXZ4sSNfhDgK/oMU3xGfXyZecUsBo+jBu6dOyeg/Ae0iw1YwUgUEqefa
tKLK3enEcssN6YEeaIVWvvP8LuJnTxA0VkhSIwO5J5AJDjqsjdSmpvqJlSGMnm4j
8tqsaavk1gS1VNf6kYaQB+usnvQGEzig0amFucyNykWOltZdBNeEoki7mZYcI+Vz
8A0hY4tVXEbJIEIuYGNP3SLkBIcRBMGS2wF3FVhcJIHp3PiYFADSMfOWkMOAjvnf
rVdKI8FLLkYsY4ckH0ROPHJzlfgROIyMKAVJzJEm9BwJS4s8wSNHARj/gKqiOhkF
dt7qvz21K1BXbfdYfPfehEVaQ8rKhkeCch9rd1ZN6qWT9IMPxyxlH2bFUH+UXjHB
qzq3s+OSDWS5rYHkd153Doyja1qaVX9VM3r4ejp1uzUMvsXxG1rdCSvcz4FuJu87
RDJxAxWpmtQk3ZMh9uO2cnbZnVWPpi4XXQKuJQfw68BpVNazoGnN8r7rm6VGDOPV
Ns+kYsKdbph0LmGPo0UyuJmcoa0pi4xDN0As0iGWT6Ys8aeiDFbcekm8KlQVcWYh
wN8JZ4/LFC+CwJYGWMc2lxAciT8PiknncdjjueUdKuZmVsV7nP0lEKsQXhJap1MZ
n6Y21KO5xHgUZwofXvcBqXKOtm9Nh0G0ieVqjn5XdWs0KrNPRVYSVQ2rj9UEjJg0
YJ6MqUYfBiPE/7rv4W+PItd/nvIHMNZbcbFN1s0L24SRxgVqk2tC6LbST8fxQipR
onfsUtyALdgzeb5ow4IjaFVJg/D7SeN2MLEKpvuSh4tatLI/jYH/YiDMJT3x2DVM
O1i/z3+kFxF/M3S/KkFp5FCSP47l85Jr+HFdwG6n7do78a1+LtgwVgxykPARzU8Z
9DdgYfkBvO0UGFIv3XYdrojkjsKk6KfOWHrl7ckAcP00wb5Rmu6x0qbvEgBj8v88
2O5w1AInM3ctBtHii3n6o/FI5BP97l3iN/cnpOf+y1U0J9Sg/8hSvrahFxx7bz1K
wDZR0l6bkXaM8bpdfRxv6hcOZFvt6VBp+vndPjP9nCbHh3NhZc1duMwwqz/dMZCj
rucjgEN4UUxftTDtrGxVk39EAx6XD0/iTmhPv7sY043WFir1t1ehy/sKrWDBwObb
l0F+i+MCTx4xJAZzZRf6uIbtjr3ZMi2lmm32A4vWumuGGV/zyInfGxseWb+lhZcD
Wqjw3/t+OU/JWFTeadk96vS/7scxJZ7jUfThcod4Z5ih5AOUyNGdyIyzsPwyjclx
GnY9UwPslVyN4hqKRUhP84K0q33otApHPqWVJxPihMRaXec5TZu0SaaxZOWlAmBm
GJaSt9H/79UV9rpQGCrudqiNWAgG588Hvq9r/0DVfm1shz6oqTSxKClHHHBl6JBr
VhfdrMMOx44cUfnNAOYdaDN2Ll3awe0VGv59zxPQgxbyp9zyoKNg4VpEHisqv6qW
T4TwFqo+sywdVnBjt1PMiuziUQiFVPikdhtAJ4CF7KdcKSbcSKPTrbGz8UyzNP50
EPUVJTExPo8VwuvySJnuABgjShzstJAVjLCKAIyfB7d8oHUUQeJhiD6c1pbgon3d
xGUTivKbfNhaNe+By8F97v4cDPu5aUXAz896ahSInzFdfiuJl/m48RADmCEEYKvU
Ny2Pm96S7huCTJExrCRRVOTojCcrGscFg/qMfRxXbv/MvYcrk1waPIPnSnPeKDWK
PX9csh8qF44CqiixUviYINaqAL5eIYh+At/g+MFdGgWU4hNdzTzUo4s90FKWKCt7
SGqQ7ekVNdutDDWjMOt867SHcZX9jdy4M5ggERX2/XNttcSoYnxURFo5PPCoXgQF
Up4i24RlpcHUUOvq8L70gfyPVESbQIO0bqzaB5ffTkdG/9l7z/2JtGU+5GQc8+JH
30UfXAUo2xaDZc8Q0NhD50FLmyYVke8FdwwZmVwArsom6Mq7uOSf/iOGUdZXVQKe
huuc4qBROjSzOljNF00vXc3rM6EboVsFGkzFlOVZk8YOTSa9u8zQTOBKeQoJOQxi
PnOD4Wl4nzmM1JvhCRpjQAHBT4m6jjoWM2xi+u+S4rndrPWPreFtBHT2WXBN/pjn
IMrzL+j/IrYuZ4+DbQRCQAAGw7iFs7GooP0qkADgQea6komZR0xIhYwciRA4d0Ee
JwKyo0R9o+wVmB33zc2KJ0OZl2wo1lp6lob98Ng5J0YBjZ3nmaDJxopjd8ap6YbC
M4taX2X3W6zLDT/ht5yWVwnaYdOxjjM0VTMviwZ83/fpdZxbIbyIR2tIMHUllBtO
UP7taWMoE6NZSFQkZiVv8ICmzzNDopzmPmq/8La4NfL3K4qGMo19QCfs2XgEU3wR
4AJJYpNniyt/+NhdNpxi6p7jbugNDixeib/uqo3SRwg/F1L6U9qe7U5GZBEksG17
BAicz2MWWKbhFlEYWUXL4ffhwD5sZzcl6UCoklHtKFZSbmVz65RKkmAvPFR/0tbK
rd19QnAr7Q1VzAF8TuKfKCURuiO5fYOMJk7NSiUMszZYq0i2e5TTtHx+dw/oAQQM
OvpKNETtStQ4e8XTxUrkvYRUzipOHkwTI1Lv5UKq4B9SfpZfPq2+3+ubxXwrNTRB
NC4TC62QJrb9ashq8fxSwHX4RPBT3aj7gL1Zg9snVe0GLXedhZx15ov6YIzpH4/C
F3eli5eXQmd0D+ijMEhXBTPpQDRlybPj/mXAaKtV5tRrXuko8PKrQVwpIqcXO1ct
X9MHmjcPme7zrKcTFrHydVAZrcl0xBPHW2x+ioUWa4IRCuKJetPKjBzRNaqCm2pU
LJi8XSPiOhTD0/ZS0XY058ELsi/Z5z6PnV2vPD8VfqEJzLYU0IvLZDI8Hu0EV8cf
uOPbXrePoeV6yM2VoferzLgJ/G73DYf0vhibBNvdU5+u5oJacoh8QWuk+qbbQ5it
htw7/yXB7le+JSBu4px+H3MHU3nRHIjnRHtpyIXNxNWwni49Qk9M1N58NXrqn9V3
u7GxbyafQFgMyvyitSpW1J37xSyX8POi9uwYO7FSo958OnYuXiQwoPe9W/S80bfE
UWA9rKiUHNpIbnVH43N2YpnQodY/2p3LWFLwUlsEO6dwXSvIGenjvTUXzw99yXEo
FjdKDSuQ0zQlkSHN2euRean1YV+tQ0LyIRffqrXCQStTB5T995iPdlkTwMQtViw1
NlKj1kwxzUzJeHDdVa24jR88fegeIGTzR5qnYEf/4J7Jg2I12SN/hcr5P1o2955R
M51/09Tg/K5PtVuKpoQQxNyZP63MNCL2xr2l1wUD3THG0d36A/YVH/V5irkgfRJW
avrz6NKtFlJSiPDtHF/haf9k1V/K8nXipqIPVOuPswUDak4Q+uKe+62BTFEAbCWf
6BY8p+2C1KaESmTsI3MZelTUNA8OaFGBkMdQeJ1fNqwUmLFQVPmQwNNn1BAddkuD
2YRis4OzhiAi2iuE9SN+uZRneoj9y0U8n/gTV7btrNTrOa5AaV5TbxQP7pXLigTt
KZ5HsoWaKb744Y2G9H/aS7M8QmHayMrzV0fMET7VhThtl9+5Y7yPM+6yLsNHTMy5
rnuXWa03PR0djwLnPM5mf/I4XiWfRbsvodaaNdV8rzKO7aPSjm+dXmocMj07cpsi
h5R0Nh2s/bRbhRgDbdW29Yh0dfec6sxtl7RfkMaLqIures+FEgnxHFNvrjuJHdPE
J40Zl0beDExVTpSCFAjHvXyBCHPAe8A8lYiE5DZ1gPqw+70+QoRQPTjbELHWsVMO
I4mUEZqazx/XuinM/326oFtxdpRzsas/ENrxarUOTF2QQiGC+Pjq15k2DcsgYlmC
iWa0yXulEqw9dEbXM+PU9+qseTT1/cTHTYoxmfEL/Pz5wjMwJxCQgki7XZhDj8HV
kGbR7vgliGpq67S7wHD1zJwo19lbOrR3nzEa17aNCDY9cjrSqSfqJ/c+4pQVE7Um
YZtGqm/rH4FSkdrxK7tEhhGQQkHUc4uFOymqJwRV/vcJxIXXJ/ljnDn7qhzHS5+C
tH1lMMXgBgM7ZmqxEiwGJsISRMhD8zT0kq0jkA9FkiDYWRm6wb80LRaHbf8TzNZY
PFx6kAoe/9eYpHpCq05tOE6PCLS3GCpEAEfMpbe+3OCWCN+9rvNhhScTr8y+Awgo
UacbUnVzk3cj1jd5MTyQMvoiYHRiUjvC619VBIKeQAXwzPQk85eOwLfEIbQMr6B4
zgNTtTeXKLWsfEeIlil3FC889QF1lq4KxfxMVbRRmiTJSJ3IRFXp3uVmyZMdG/cg
FyrpTsJsKPTpfPxTIYWoCeNldtKQGzJHjYSgkd1rW8QTTvZbdypnag1G8mXomjF0
bT8cFehzIW0h5e4noTnzeGXIWivaUz92XszeIiCsJvJJlMIFLyvlZYZD3OZvz3Oj
qxzexUUdl+qrOFKMWaqfri63LXP+JDw0YSWXE9MUkel23k/qjwNRJIsVheIudyYg
n5S6rX94gry+EMwmmOuOy4p86czeFMaXESCPIpkchEzmhlHYyWcVEaBSpyEYYek6
XIQEZXPIP0xzPS9VccpjzTaDBqsvZDS3+oxCBijwoULDaNVChxF2R7eeqas5KqqE
SVIPnOy5oYcXZQ49hzCn9kGPyOk/z+WF79ZeihOvd/CkZhpnEPXwX2X961SSHxIE
0zErxyte0sbUIdK44ETuRQRyYRVAyTAThVOsvgL84Uk3a4z9rei/mR42p2Z4ihch
UVir2I5v9SGAGkJKpVQSn3+3s7aU3NGlWRs2DaIaMsRisiv5hF33AqD2+IgG77AO
k3TGMh2E28fZfB3G0iN4d5CVqeYgFsNyg3fvUfQIKnc2qQ3NFIV8oF5Ftg7E0UkT
BU+xy2/4tgE3hKlRAf+C3xTbdvVzbjCUQhiZS0hAfk1269fxTx2Vn62wKSmgkb5w
gw5L/B0Esm87C4/d0BVoJc4Pb8QyUMHPFXxOd9YTwBZE+/QTqY0K9WBVeh4E8f89
q3aY8fR0DYrX3pe+jF2QpCRhpuwzK9B3lCUiR3NkDUGsM4u5wWz1WIyh1C6KVH9B
YEUO9nXUIgN4iIN4awlEEnbH9pyz1t+Kiq0zOvwTgdmbcvQvci7TRDk4xWP9cKg0
nQPQDZhc68ZmwupFLc0jmsNkiFSXcWhJY8hhS7p4s0c/D0oVWLe3zgCm0QMBhtUp
TZ1iWiqWUgMHHTGedzz28gtTbLNVZ+LBFNo2r8LIhqm/fbWETQ4fQ1llhEu/9eAD
hu5HzIoVxISLFFEimnW3yRCWHaWdwhVQT97tkfSBktdySZIMyaFralUvLBKNiCKo
WBn32FxP607gmFRLxBA3kDWZB9gdkpXT4YsssqmslF/2zxK6nk+csX2RB0fv+/v7
KOc+XeeUVDPujX/8PbtZ/NvMO8Ag0r0UuzJ7p+F0ARq4Czq3DoMFGZqg2W9s554z
sbkkvcdGUjPgR7mIB5tpvRL8abTShMTRHoMWMTmtlnuNMv1zZXiX63z+mtv6uXBm
52+lvjANAG2hGD5I7jx0QC8x7Ppwfq+JUagf5VIG5v0b9OVhyOeiosQw6m5sTT1p
7R+DHV9qCkxZbt4lunHTbSRa6cY5SM0vRW2w97B4XF1Zvzcghp/0BgyCWmPNqXi1
fX7Ml51T1BjL7MKDlVV3zhX9USHyLQUhu8XwOufe+1HLWUV7rHoOor2tcgUuTn3m
f6Ey/+Y53qRZmNUzzIzRzcSyJVkY7K0fRGbUgLLNt8GRbtOBq30drpJnY4drfZIl
MXdxMSJB9iRfw9n51VqAlS+dDeHOm7F4jcjjBv0jtLdLOSTIug3e1YVQmghGuC4c
8prMhjsLb1y4PUzaxKDMJcDBUkIUo2PddiFRe1LQwTud4gr+NYfY5HUOUjEVowdy
F+tieDiRs3N8ujQhckfvpUusanNqlNE6ZiC+j1OYjz5iCPNDiH9HOUICGFX/igaA
6fjAC/HQ+peiHbnK1ZEbwhULxRiDVznxK44rxIYbdKN1qCrzeJ35+ibX7lGth2A/
G4k+kP+8FgH+1saeEuyWYHslyPKMtbvD5hr1LGoH5jNX2TKNIOznLL861tZkouWn
eJ0Y/CorjRNMpUlAbCY30Smii2tFmaoiulfI8bhkfH9gaJEBlkRbGkoiH8J4ZPWd
sO+UZF9TTN3BC94G+X6+6FBm4//DQwKggZzRYsXMcNcml1W3Z7zGVZRJZnQnKXp0
dI35Ha2mpAVK0SXF7mhmFGZZgH4iB5AYM4IVlKo6TB1A5WstOP1rOXFLeOZFA4S9
rfNRfHiVn8/Oen4hZi9r85dqUnkrBmxr8Heu3uY9hw7r21NACKWqOky4BjDiZ2k1
1RlgPd/qeeKBNncm1aYYBJ/syLa9ye0mADrrvLVLqswe5teRI4L8bPA185+bCc7f
usyqFgpvi1Tb8HLz4LPEMLUOL6jG4Xc7EY0T+Nug9+3sLb/rE1rHNcmo6njv3omR
zjVuKdMEBLP3kOT1MSyhu2IV3EWocrfEdw8W71c6NJsznpWkGhWp+nU5DCrWngcr
Q+TtDOpPuzr6JzfeHgXcY36/Xza4XZn8s4ZSi0NPDLBycGb+Dt0O8r0smHOhtOhj
Y3fuKD5ag8/zDuzIcAII9knX8UiTRNJn28valkozjRKv1dYd71AI4aPuZMVlojhF
wQZT4Th05KSpaXO8UOBQ/pwO1ZloAalUJPfmC+SJrkrKb9XM67/Wtu1dRDZqCZun
pST6GnjrroW0hIUCF0jFnt+E6vAp2m0xKQwi7BYZwnpM/BAorgmGkpgh3wAKwyWL
n/5NnuwlmcH/4E7MqtLWz4LYkXy+p6jc/5s7CGE/IxsgOK0Qt3GEGW2eH1Epg1Pz
fgohTSwIjMSGNgZ06BkgKhr8lq89r9CO2Jgz85GtUpdJc1kk+/bkd2UG9dXP4e/s
JNs+I990Y/StFAAab7WlEG7N2XDaZLhrQo7ArCgUMluskz+bcWN4n7+SsziReQHR
uC/k6uau8c25g18kcYVrCMecAAY2SXtxj7BgBjqDNsekWqsej5nUzyB1KWiJIIaK
h0333KW3xBZryIutUqc7laXH9JoLKOLU0yx0br6uZldBFBJxAvUce9WyhCPppnWA
QkD8+nrQvX/JTR9X29VntSfs7RIwAfKMUtBHJOWPDqFB8W+defSLPOH2BEeBzQoA
NJEBxOHx7vPChoFUVHoL0g044N7YX+vroC554Q02FAeH2epYjZZl4xICJ2jSfz3v
VwE9vAgClcKDCmiBvgFp3QQXp5jZtw8/UJzhw4zTnyMcDT4gX8qTU0TRvocejtkg
xY9H18sXVmn/3wTrdYYI2Euq+VUYEhgA3hJQVbPFY/rQx/1W8Iziv/orypeh+por
AOUKPDBaFOSpZoaQFEvvba+hiRXA/f6HFqhNhX0qantK/fdKUHEguLr2mwisVrz7
6+cpYVsv52jOZfsYSu9MizS4LKB/BJBcikt7XufOCXZuyGu2cwaDsd2qCLXwUbfx
ofN3Ehx5l83N4nxZmyid7GwmlLYUnUZOeg3C9sgX//L1XKUdfkNTW6b16kEss6hC
HTJH7BBevW1RnnMrZp95A4iFnMeKdTXuddOeHKNkSl830BYf8HIB7do6Kikn/x92
MUJePuBvOKOIIkRGPYUHhG6wGJwJdf/pSwOiftKkIzfk4tEz/1BGjxlkadKcABuB
5o/Y3v+N+FqvSkp94T9Gd3OADg+qw0C5BkiBPTwtc9qJvH+ciRwdHY4esJ/VX04J
YuXI8N4aG7pk0dy2KwivzYl0t1VPSuOgCHCPF60a1/8hkxnkOFlIpjV2cyFwKlLq
hjMccf3rv3rc4MWZlayygaT1g6fL7Hg0RZ8wqALlefLczVu3/Zk1/PB0yr3nOLwh
fUEssesmeISvdibC3Ak/p3n3qsnw5zwIxTu5QJpyna1zzxG/BotteqI5KHQWxpV4
ROVFKm6O0aHitUkMh1oG+8V4OpQJM7iPelNgOq1pXgeqvkGUTKlbb2wLp1XxGLrT
k4XtA9Nl7SXCDf0wfVKiBIB9gumwBNtcXus9AW4wQ65+4GHRWgSzly+lb391D7Rp
JezAIkKKBDKU2EBOWEw1vR13mYT5vKrUYMM9X54qFMzxmBb2Y/fzBojZvbcUb9/J
Bkf5vOr+QyqP95nuXZGdKyFX0Tf06Ylj4bwPvf82OIQZUZme44Oog/DuB5AhoufK
7rLgqXu/LwhLuMFsWgvueCf2DPPIBnvyFI2conHcDH9i907cq3JJKq72m2/dsTge
bmIhLw1AnmYTeafoUGtJ5aflHx0ZKGLXTOEV4YlW32QEjzQX2H7JCR071s3P7bAd
wqbaVBqy+S/RPHEyC13eEcmFveh25I1nxxY4aR1YULOxFIe7KcHq58uLs7fLjCYR
hoviZ89owJKoX4YPkcr3fC/q0mQOq3sqFBspqexLJKZlttVoEMqrBzJcGqGKlXSX
zZaZLl2kTa7nRLsMqhTmNd1JPO6VGS6i7LW5UZVpLb5aI8qp3Dy2L5GPiL/k3/AX
lkXzH/4wLD4xT38fEfjLSZwEC0a6DKMmpD5+EcGhNcJ/3mslJdoaRqxNDcN09N0F
b81/hNL0eNHbOUruXWv/L7CskDrdGsBCbeQ6WiG7mMeREGAVCZG+ulMP0you+y8i
oReWOM9s4WR4h/Au/KfQYRbbUmOLNe6JA4TS5+LcnX95cL1nwh56oVLVJfGvSpKI
l8nd33hGxqVIN+ZzXKBngQoO/P0XlkiznyPoC5v3dM9JlXO8GIsoUUpvMZ4reCPi
8GtPx+yZtgXK8b9vqA4BAWCh9O62cNW0AuvnjRL/RF/4wgks/S8mfvmidZTtedgE
i2yvYGeb3SG8yOUxfH6QuShnV+Esu6qP8kg26Kq07ieXZQCXEx9CUX+FKMenisil
UriuEpvcjxIk2zEQQfRNsv6SyKcpCUVvHkOY7ZpPhwgoDES5UT8ahiyNj0CIO/az
X6qtJIBHHWlXmGKM5q0T9EnoYjM+awAYU7J4WeZ5EtJJ7V0q6FA+e2ztLoCO6seV
YVhlgT1mxQe6tTbIWETfpGx4ozLV2a7gNglczoWRF8F0XbqjaAMF9r7UU5OCULYF
RComLD1pWVMlYz99lfiQyFCzZQAHwtlWBoDxQeh4+3h3t12vr9RoL+5MmG5qzqE/
895KeG+Nd0uDzpHWMNV0RY6Uj8jit5w6wkkBKzjkaAuDZsDXqF/rbxygqwJq1yl/
0Vj6h97OkX4F6ygzmhHnHmzuCUGu+EkBbM4SAaHgmtTqf6yUCRvHV/0RndVuxnLM
DNZ7tuuamtdDHtv7tJLzMZN3YWxyQ8mJOItIgoNMG7W0XqxjnY/0MrppEiNcgOCR
NNS5rPRiVcCQtp5koBIu/oY0hHX6MfaAjUWEt6Ahgi12estYIw7GlpWRtLvaoP8S
HQqi3E62OX1wlrB0umgEhc3HV0M6CbVEPOuDm6YVgLGJnZXtTAfMDyp222AI7S6m
9HB/buI7gtAuOfB01tKZW9RrBRDOSftKtaMbr1TA4IpufzAq+LLuFqEMQbOIy1u4
dGIo0lmxo4BhLO24PxlawMLrpbyBZIr8IsXfZAf1xHBLFToOdPVKcUgBhhKgXJr/
dtjBQa9OS8HErfRKIoQyuqDzX/K3CzGKwgcnATSR/OPYR6HFQVOQEj9SJwUX1qxO
Oe23bC+t+qMxBAckPlpJ/y0yFgJJUT32nHDaJAY6Q1gwWZqqZlY/7iD3IaTF6BFH
5Ab3ghwFhJPhiQ00oGcHyal/D3zW2uJxjxefkJ29aNzLG2XMS4xJUVdqy2NQT1YI
O+Ea1Crf0c/tq25kElmpWA7TlqMj3kMCDLcyla6gW9iE9Hr/oPbkFkqqdh6SCHwc
tCS2zwXjGqOW23TnjrWH7pHQ22h2pPluAGdzWd6OBY86EPMmdV9fZOc98L2jKby+
TIzxunyvMQ3MRquzUSbYilUSZCYoyjXFmS3t7qpVPnAm8tsoWZGLnAN4QoRrpQ0E
qcJBFEsJSiX3wHSv6oKY63eMNEkG+9p+Fe4NgpiA3Y70jLwQSp+9+MMgGBcu2WEw
bPlZfJXuWO132tm+H+1fQDLPVoFJYNTFxrgI4qtE7bqsaIFaIQZqKsGTaJI0QtxY
EPFFZOYcDIn7qAUNUDTdKykfNNRmwqTifJCSBVJo/owSH8P4HSrZBFSRHuJ6PUlo
n2SxKOh7B25uH5uwSM9GzOkkR1QQju5xK4kTNf9FysyDmC14YUh1G4duzxi5Hzpv
KomBA4yUq3L3sS2Kk8ok/Gfddxu6tkpIpYirfAUKM+nyDlX9gyZI2PXlH7wmfoyD
IaXRjXB3/eHMrV2ybZ04nCFNd/11chUiAekpq/AAkXcRJRN8K2fQBgg6nZEfwZzC
ok1O5GNZrOxOk26mLYt6Fw8a7TiyBd17NPqSDrUPkv1jcRF4F9abbhfOOJeONRFD
AddO4DPh/bSyZQ2Q9asuZVWSUCpdHUU2Xydob9kRnMxb1iC/qqWXp+6L3YyfiECC
kvJLM/pRu/iN+2Rz2j/siZyupLlPDWghF33nD86Lu5hTp4z3RxEYBq9thUuuIk/B
5PDL63nVtpuxd/udoGT7eKUfLZHxwHfkw8FHtU7qvJGG+d+FTE3ORp4kZc0riQzy
6x1bdz1PRk9KwqzjQOk4pLR5hGIdXQ4//kMnOsX1UCz1FuSLRnFQ3urMd+NnexHI
zfjYO7s0mRHoQtznVLAKE6WOhfVFTbZeC8Y9GggIZrlnYcOQVK9MZXC5qA0KFCrG
019O6zRcO7KuNgLU83P95hJlOcBmkUqKjaYhMaZW/2Uhb19uGUdBpSmHtES+xyPS
OVBaqPON503x7Wq5bgDBIyZmJb/I//q5aOJFvmpzFjzGx3NliKKiczuAcHTa79ui
YmRfRchNONT82QOlhJgNUdRr8CcAq5IDOgnUgfP6yb2dfZY6hAQORUqBszL8DBZm
CNaT9E8xn9KEXZkdw8LgpbBbaA8cY/Y0mqjwpybdCXJm8Fyj+5FVd4dKG78Q6f0y
GDjXqs0ZFptcBDIvxsqxU1Pfl2LZeaA7Yysmfm4p+6khBlOpajDVyNmMGYCFpWtC
VNw3ZqRvAaDTBE+LaxIrheTpyW07Qig+XdGcJ4HLHkCN+DX5DoKTGy7hDvEfIy/3
dqIiuZSvlwLIzV4sib3j2C4dCMBlX9tPFUE5m3qNpDH+GgzzQreu/8YB+8ijXfkz
rYJS4vLTTrhjHzJNJgZJ/Qg5Bp0qoR52QYEzXxfnTwCAg+fI2ms8soxWuOYKLVyk
k1avWqUTiID9lB8tDJaDzu36x3rqDO8XlnBhK+ziI5pLvz/AUbDmJOh7rSoXmMYz
a0PpmwKPhKIjzLps9AVK7inv/Z9555eWe7qmtr0TKM9tkkN/5lFIZRmMEd6kQPBM
T0FWKAV4LEwKUCGNemqM0rrB7Dh5lmvtWfptPxDmJ0xscEHaFmoaX0MEWtmhV37e
8luyDlw4Dmh1+oGWsWGiTcysLRF/t+IjyCrn/+18MxgaeFpLlhH2cVVyrtIbNCcn
FvOX2WlztjgKvZRvI9yGeV73mfwvl+6gCAyWESNQBMGphGYI0p9iMTNr1CYtrnMj
y3NdQ3/1PFUF+wDVQ+Ck0p1g9eMzaYwS4uJpnd0QRA9f9Y9TaIMfxVuiVldcM63E
c7V2qHIwzbUYN+9Tt5yjJhBdMSI2rxwVtSJAVIrZuP+9K37hwTXSAcxNKkOtZjoQ
WH7nFt5yRf1X+yT5steslCYo0hFkfsVRBs/EOKsmlli/V6XHX87FgHPrDkf+If2V
fdrgYqx5SAaLYnp0CFruGyVRBEYnNVOxMrrVOxH5DZbqY4dChUMIANIEyZRHJxsI
tbjXlWIXy3k+bW7ZlZJVNZ7ilzGkBcCWKJdCwCCWaWmWm07sBabp+7+x6Hj/eBq5
aob7mWE1wDA/GwQi5TR+dUsLZAwyr97QZ9fxMvcue8ngfjg/e2CNh1osKKyj+nOQ
2fhF6/E9tp35IdJf1N7OJPO0rWR91gtONs1xIk5EMfTYpIDXf1V6SDnt/qbjV/lR
dJ31wCq1xjjK58ZyefuI7Jty4ZS7iAbZinJqFGKo51UvDTrXmHJOmwwDSkKFRX4R
YA0TBsLxZFDx8t/HjYzjQnNLEmOjuaWrjNCeRk2z2kgidVMd8sftwj/Cv+onxPvX
2A4N3Uys2w30vb4Y33ia5jRCLOam5nkbZt/cyvNbwTwnWig/1ryNQ1L8SNDmFfNR
gTIQ2zSE/QTfUhDnw6SPqjYfTqMn6sz2KA1Ye0sr3fp07XjyZJFO1JtNvu2Bwprj
j8sk3i71eC2wMqx9ycR39UlxFK9FGq1v2pKqF+5v4clDVmYcyE5ig5Z+DFDbvHke
shje5SFGH9hK1bLUZOkw4uUO3MiNhAhm5I089uKKPRw7H+HuLEzG2R0azUPiBb45
YnCfwybXi0dgJzL3T1UxsbRnf0JGDI9KviKblauUdyaZZgQZ4QkcOosiKPEhCm8L
K03lHElr+/HiJ2sJXJkfO3igu4gwHEFu+rLxr+XNtzg5YFTvDBm52CwonCCmmHVn
2K+nx2PC8UUTBsamZxnrvfSxCLyPzZEg96i4eHykcSFN179onjMx3SNrdOQ8L4nA
+9UjZWJ5Y19HM4yZPYjCHuS1+lusJKAH09lte2fPbU3Om4CfNCoRLtnUHbWqXEbR
Gwl39tLTstQ5Tb2Z2stbFTSd2QPredTZFbW8Bs25gs7RKybwTcaiYe6djZ7K1EbJ
vU2ot8tqxqbt1YGm9cHGs0lJGq60Rp1KfJi+BM422nOkdXtXp6f5FqyGGRToGXm5
v41nANhT585nFDPZE2oWo8h5IjbGXFOeSKwJPAXFZPZ8cOQTII/rMzq9yPe00CUN
+VBPcxmq12G4KVlt7mo0LMPEOeuPZlpoitDXli4s3DT5gqu9QxDtfn8M/u6Yn5nx
t+Xeb0IlfPYPWgyOG38QlWWZ9jiOyfsLmru37YxGW72B8TSS9sDeSXGVpYZj8+E3
uvP2+yip5xWPTsCdB8B9WKLj5eNCmiOnCUqsf3wFdu9l5CSk6rrWfdwmUNUxzO31
BeMwrwtL8tw54tZR9RqH91+cpDKFwyNcy/a5EjBSrejwTw1cmLoSAWfXUchrWos2
pZ8Dz1hJRg7C7s3Y/0emZTeA+otm1YXGJot8ObOiDfyPuVrh82w79HaDb9nLi1Va
ulmwkZJCJmiL9isfnO3vKAlg5Q1v/PqBVulTxH91k7R7VCtfCDP1vfzSi/xFQaDI
CGkR9TkGrtfrvSpOlO7ZpHDyFoT1Jv8oWQPyQzclyfSK94b1obV8ZAplJLrO1wLO
dRGLE0Rm5QflaSjx0Fing84V4hNHk1j8CnE1Wi2INxR8SR1uI+HAB+6Gifj/e9I3
kOsMSNtroOjdlx/V3hlWCIHuLvXRtBbIwSLXvk2Mu6qxgQlIK+EGKEqdVWtaackT
MKruWQnQXbmvzh7v53Pj43EjW71JiWE6vvxvSpDs3YFJ+4hVuYrbXBFptlsjiyh0
jJaGqbOUNn1hWxXKKCSCMHmtb7NVTAaTaDh0tLDs/OQU+bV1NgJ7/M99wU/0vkYq
b4EqbGJ/miKXfM37LU6imIpGCjy3pypRjoX6eN70Y79AFoeqfDJklWFlCeaBvt5K
kFI1X1TmpqEC8veIkxoZazh3beuI8poyp5qg4vLV54xMlWdGPaLpo/HVULQi1aqP
SiVg8vRRJqMgiO/RWveyUEVEt28pdrLYnWfEueeTV+VvMgdwQRIIeO6c5VBUusGn
ziQmm6nsifzlOjt6hbNs3NA+DkW24H6UVL6zg0XBzpqVdNgezy2ySO4VfVzyL5Tr
a+a4+BFi/midJ0/Z3WS24DYRmADcBMusSxcb8MytvayDqzJ14dwWamS1VK1thtVP
WBswfZhKV+WnG4U7hQEsOd47ctdc/c0X6vRUpiV++p/s27Whlx4mXmh/o9qcXVuM
YmsF86foSlQenJoSYPLIrJ2h/zaRMy++y/yxanBKmY/GCEuzLAJVdoASy9PROnSM
ZzONBKel9dXGpI8euMvlLxnWPksefqgW1njb1XgjzO1Iw+XXtSVrIGehxAF6LdmZ
17V8HoRZrFJH5M15SOYwHLhE9Bscdz/hQKxVunPCzhz/q8HNUHF+U84RFMXbp/yd
erzOv4PpYvtd0NmQVp2h/kiO+aAQDLE9/S8TbUz8PjO+JDa2JDNV6QKvLlPrCxNb
vUJdsZWYomtw4Kbl58sUbJa+CfgSRJNsJn4qFax/9FOVU5NAqj0pS7UvhDofKJ71
rX9Y8iWGS1+JgM9gQaOXtM62dEIljhLr/l+7C3wkU+xqZlVI0n2tPqNafm7Hxtsa
WYqLIygsyFMjXOzqFXatU+MFCF0kkBNScD4VKzGqQ4iVJaKp6Ujxov8Sue55I72y
GyxUnn+duBTtCKz+dq2lL0hBdwJVXgh+AX9zXWtDx+aDN/jZ0/8pNlk8cdpBdJJ8
m22choRlmt/JXJXq2aYI8sf8xU6hMddhMmFEovLVPSDM5EN2ELBNtTuVE1j0/5af
II96rivslTvuuQ5C0/zAnHokktYAhGiW9QDj/BegcBqhIeLxjYplpQQRGuT72VKJ
cLVhHILz/N5iP5t1ijOt+YBJFc5HB+rbwgMlp6Q2M1yYUx/a/53Vr0PRHWnj+nxC
5DnjFAO6jFhPNU+itXPzGx/Gm6j6mSiOV8fqzm37Ji4lnhLfWH3nS5L6MxuZfqz4
J6CfphT4URYRrpNI7TuwEWxYkIWan5tmjpkD5qKrtjs1MRueO4wxrEwnELnO8Cmf
iPLjQQ8q5UZr2YYHUtvbGtzweApWncvFFsl+cJh7qN9lSKssnb73Feh0gbNZwmtK
i4BEnaRm4LahkbC1SHEHM71fcC2dRGc8Z4ItuZ4MDZc9SEAjamU4FCD75rSq/bdG
yXmjD9Aj8BDHT2Y+zYWz/uaPQ5ENr1hEZP9YBWAW+jU4XWXorODKHZATMAhdNVc1
Y9gk3253lTjCJHv+Wu0HO2EALulX9IICDR+BbOSukt7gzCRalQZ/BGDkWRGwZeVZ
+xYbNm0CiVzyMgYMmABu+B8G91E/v3Al9iZWturaaAgIrKItLVm07/Hdhe+9fBvV
KJCK6KLmQuVgv4pR/X3zlzQV8KEurOA7fGszPl9ZlBUUxOuNVzhSFqx9aSCNeJ0e
Zls9wCNF9sYWK4ZaNawfuUNjlwi++60gRQyay4AnJBjJIkn65qtnwRAg4h3XVWgq
B17ej++ZZJqPfPieY5Zjx7jv5R1UW6O+xQmnOuk6sTQOAtripEiHRZea2W9RrRMs
Lv2RVsOQJYCm/eNJal2jiGtv9zOKJ12Mv4pZingKoBRadFyEgdx2F87KF8PG30f0
MLoigOfLf3aTM9IKyTDlhUPyHaThYnJ6cjpcHiAE8SY4CYtctGsS0K2RXUb98FU+
sGPKO80J3V1NFUdBbNv7niUdPwS3Wsdm+oG0L0piVtlyMt9XniWiXz02nStwUDrq
AksvQx+6VsivsmXQ2BUBdaxWRX5qI/f3frF7zx5rDOBMu6idMn1aw6KJWNOtgj40
fjKhNxN21mpKEEWhTnhhHYj0ZnF1Xin13B9gxPZ+xhLpdwYhnj57H86BsSgEE4II
IxgbFV0dorrJAecZMyaSh6+Oh6AZKAY+WYv1OGMK2enjY98xHK4UlqgjIYdWZ5kC
wOCxCJtrW2GscYzP3xjn4+Ujnfd+bnPDmWZI+2C9PG1IHVnPzykf9XB5zOm+7gdB
md5oMYlOKJ0w+bIBIl132W4VKn7tjbru1EhA50j9QuK5auJKcshJGkZqz5THAOSo
J0oQD+/RLdQbfUxk/BNX/s2L+2YehhOIxkuO225/TafqZQSs8OHHPVmXDSLLdU3u
31VDgUXargo12kpTLW8mcVmxmMByrglGhiLtg1SnPR3Om3/RU0VQeFIvEgbD/m1L
o2hQZakUg2vMP6ehy0fJuU+EwiANNSqW4khoeRaSjA9QqzcV2IDHLLMVNDcbKmyy
T805eswKfCT+sOZYXwZjCv/Tm3k1FqnrgzMQ/HmxbDdI52rwDFfI/9DC4f5q9k6l
NMM29UFSeUQCianpfC/hr/C88VYsf11opG5bOQZulBBJt43Jm28wS3Eg3ae1BMNT
O9/2Y7tsElXTchP69/viYPc7HrffwadBySY4KG5htgXRJ6u9GduGysCT7aFj2ttY
MxtKlsfrmd9PZAGDoq2R/Nro/0SLFZh6L4f/mibn1WpTXWQtL4niCaiJpNye1T3A
nARDtBmJhorIt4ADAZWAR11G/aBymD6yEDfv0nfrsWb7vhHiGtQ4FOj8uvvRqLxI
Wk84Rx1xc3CtdrUjaIr3nGKD2PUbscPXuNEiYM3aCVdeiGc8SV5SpV4v5soa3/A3
sb6bozP9bAR24faVVF9rzZExy8Lw2aeIoWwWFm79ggIsBTS3jcZJAgBilRJtfJBF
hVnqjV6h3xqb3+Ba09ZmtGy0KVqvXOtVk0ssb2Dj5rtrLD3WS3YhxQbZIHS+URyY
PwpqtOTwW2emcjbiV3b7fBmNBX/GDyUHZDkyi6a2rTRY1Vw472iKMIeHXe1QJ2QQ
NqWnrmUlEla1HdfTy+OqAtIpg2guomhg2GyD8C23lRote11EmOnHcFodsywlaWMs
0KnsB/sXRArT32R5xp7HlssD+jIFsBn6rtTtFyd2D67DtfbCzLjgsmBiIdhE2zWT
QJ8W8NEejVDkipBYpxKf07HZZCigkJYoA0P73dWsEUupvhRRG5XeG9nopZL3ridz
kyIKAZWTgMi6Mh7t8NmKohCNPMWdbAop1LpqeAQKXcUPmMQg9bepyghFB3wWNgIt
5d3UEDnm4PEaJbBuOqOzJg1QwD58l5z4Py6ztsYCkhbbykQ4o+HCX3U/JgMwkdgx
4JQwbV10NdfyXzMl7jtMKQ6IT7yBs5nzTRtBf6KtJpFD9SpS//P6leBu6FuBctRr
dX50NWAWXXjVhvIUnOG+rJeXiPMDO5DU2lj2dsQjeKrTqDRvCy92VXHU940+fa6n
GPbIvozCMHeNV0SeKy+gpJBCKoQ0RtmycJ3FvZ3NoI4qoiqed73TPNTPdrlpY83I
dbIuF86vXhekQse+4H1de5rU9GiXHwV0Pp2MxE4leYMOmYIXy1sljqjbepmDi0Ly
uNaPRJXFV1Ydzap/MVpRARvVNX8LLFOlOcDF9gxUWkfc5ynEZQaNxz4qhHtZvLeB
zBQuqautUw54vkk10Uukly4d8TaRDr/aEouqKaM81VT8yYThsGUTRE3AQJpP8VWQ
IpJT9HQt+FlRJgP1KbgUwAGTLdWo/uVj4aGMQX5qcVJR5p8RVy2T/k7SDzoWxmqW
0xTUojneMfRadYJkD2iMTeieCpjC+FlESJQPHfgQIKJNe27hUUVQLW98kdSJCdlE
H3dCNZ45ZL9GVTx+Zqkh/fpkA9eQTa3s0Qt6+ZasjlKy5CflSaMfAyZM4ofZPj/w
hTW7KkMG1sueeFVLjkshOE6kiUTNeMm1cc3xqMEbIP0GfYA19rVAcTCMJItUf6La
s0/nOhFX8cBKqPzLMk4yqwUuv9/MVkPwpiI9ROrdwawPUN5Rb7x0BipA/xASnuc/
FaOD3/tR0fSU642ctK3l8PnI05e88YQKpgRPdDyvTXr5JtN9CHdbgZlLxrwhZcuY
zT0aEXAJ0O7c5OCQmC+TDil0TMUbDMAeb0kq08e6u+A1oN30toXfy3ewPlAc19R4
mAxiA6/CnDp3UsyiJ5Zgw/bokLfLHQYVa44MCb1QeST7895peyWdz5s1UkSYaXh8
oPbzq2r74SURynYDJKDSyIpP2unWMuCXWFhUQBC4L8TPlHhD7GZXjnAWBCYBwc0W
7DMKxgljrkECME/7J41A+BNoByTr6VUntMiV5lshjTR/9lMDX+Y/6PnggIeFNcNV
TmMptbgP4D9DWzQSBeSQbsWWM8v1hkagX4zLiw4MMn1UFPYXjLdHBfR834RjvU91
OQni0jXbT4wAYDBtxEFhI4JEDFJCRoY+NTgz2UPtvuSccjvWMAkueel5sSnbgv/x
RJQx3lZzrR5L/HKbW7HDUcVw+85vDU68wEcLB4oXbdVdN7wBXNENkTku+FIRSjvn
aOuU92/8elKKDea61Mxsz0kbWyhPRja13nEAsdyhrBYuVjKwGVpMTvFWBfQRVquh
pfBaOB9bcUhLSHapUjJ2yR0hzL2Nez/cr/SzXDpA4oacoHIIw/pS4RGoqGCK7dOu
N4/BpudnUxi4WNWhvP8cKuRMgWNImGV12EKvrPaQLANizAIdP568zpcZWj0CCdKG
6zP9IURa2BrVTpYSycnTC48A4ex/1UT3DFMqZWCiSXqh+VpbS88vCcdUsd6fW4YO
pVrWGmsc0N0uiTm9cvLsSTbQcrdabXp1hbNqvYdrkXnCyUzyLlRsekMB2O2CqXT3
NIElQXLzhpaqpLxE2KtSuURDf0dSlLs7OnFLmIaVp6I2NAOZoIf8bI5YsHcA/iwJ
Q1rjgZZozK4RucRm/XvPqeLdGQTQmSkS4TDOIpMPm4dC3vtlu/1KEgaezPcOq5Sw
sNoDovVdEj605ggg6aTHTNc7Rh0EcybZ61UxU5Z5LtFFvYkfsQCVnvbF4L9bhu09
fbbuR1j9ZNxDOp09SnyGbI1vtP5W3svIA14ZJSma0UTIaAo6cVfLBL7/8TdOkq/H
SRXSN7Iql27t927itQbU7S0a9q9DOeQLK6E/i/JRKiDC39m5cnIRIvHg6eVeyXHY
YicHE3/H+qQwKo45EbJ5oQqdDO0N+36eYmq8xPMOgx+p8ut8aBU62pd1FcxCIzW+
aH1WtG50NQC1YQkRegtsqH0l+fh8KqCSa14wX3ZZ2nR5cKo45+p2Q1+1xaHwttqH
WI+7VOuYr7TGHUz2yhhnHVu2hgzDooxNas8Q/pl14ZO406aLwrfL7QfwwJTw8STb
/rhWGlq/MZ1EgMImv11lpoFzPfL4Q/3Aj5WEGyLnvoTnhnKe61O6vs1Cd1skVpL4
uIh5y2U2lleJBcxWFDLj4hM3NmWEyLW0wUOvqTSu2ltGc4Za9gViKa8FRVjjUIrx
WWACsHHA7NauJZvy6HQ0x7Qw5LgbZoE7EvKZtzAX4RpV6G4To8oVDitLdCQNwBS4
64e4KSZKW5wOpFhMhSmi4G1NoLKESHoyn1aCc/AhZlewuvhsLT71cx+Ve4TVqs/s
4JoSvpDEumZT1ASUjA7OPCy2YQjTFIMol2WD0QqCcaKzObl9Uy2E4b1cby1vtHEZ
mMGKgxP8H40lt6tm3f4GvoXjqpX9uTva3tFiKYv4Jd7vgLtmRIIIySGFGbl91JA2
ZfOWw+LiXjmQlDLforoVvrdEth9mllyHrT6LEL3Qk2DL7qnMjj/NoQ2uAOhN/f5f
01+rGQG2i/xzXqPvX35SePXOvI/Op24SMRhLVNjiuO/alsmMBetrakXU4rerWQQ4
YZW9lQs4dnTHq+DeAIifJ7SihLmHb6hcxtiYWc3rdtdtBu/q1uXcANGpU4ZNCbAl
FMVl+jyexr7uggCoEzchPLYd0HWWC6XAUA51CYKHxbCcyvUgaOWv9wtB1yR7hqf1
d8oRb8vUyJOihflqDJHe8fXwiNXzeFYIGe4E3cCy9KC4Q01e8F3rPk418pBUc2i0
1vFmphiHJG7IL67qCZX6hfgUAA8F4tw7F3rnvVTcNmZWTzRGczrJJw15q1U1nLL4
p23WAndfsRn42wU2VR+bF85/QJucHOKLqaPipJ3ybDatezqbuPxvIknjUu13Bh3j
D2YyDQyFkof80PMZIjbn4SjnwZck/bkf/Oklt5wTM1uvcXmGvC5vTx4WRT0vfp7D
Wt7xoocd7ZV+QDLX180SN9QOZLWaucOcjh5c0pNNECAlYfuozhDrztUxrtbY5gIn
Bv0FkGroXfrhJR8XAo27AOOMx/tA/w2SDpG/VKN0Gwv1ew9TmO/5/zYKV6ITYvji
V1psOe4MfDrDA8tmDxyKAfvJxM3SPZquPAc9nrD0HAosYVIX5v/xq4jHW6ZXSiMm
9KodNdXzn0wEz0z3VKlgLfJQ2kPBE0ZwJ4hPe2NLdhy1/ZdLWDKF+a+35sY5t/ov
yxkASsQPpPiSAB9Z7VE5lEDYa6nCMv0Vuva+YVAngEgFxFiwDhNupwGVadTyEf2L
ldToUzfqi72b3C1JxvLGXKn+9reHywf+fGT2kczNxpnW6J24rbHRBa5hLjQRsMS6
UGJ8ED58b+oU0hXYdpvAHywDE/oqCQurlWt4rUKpsrpfZHQ7bXSjosxZDwBmDZuM
Z6fo8GBNGjeBcn4oPe5iMwD6QzhfC2f4E0nZX/nXOB7eFPneatbBE9iy3ZkHLox5
dGVCL0jcdjduCOyhroGZzd08BGdxUCR1USFAd6pndpMe+h/hI8I3oNrmhn617dWC
Ij1EWqjlfh8YFAeQj9DJ41HLJJQSplnmrn++O2hy2W30XQ+2c6djA5s4OoUbLpsJ
WB97M8ZJPo6S9AVU0VGRw7c+ocxm61N061KlQxaGyECKXy7Oc2mX50XVST4zukfV
4GD05+0Ukfd9FDCsRtugCvftYzy7P+rnnLlYChPYgZ2nUBaWCwnZBblF4hLweWQf
ZbWsfHqvUKJmsfyNSWKdsK02WbIOQkcvyrrUR1P6D0On5gKuEXh98H/8vwTsfBS4
fW/dK3ID0ii2rQOOmp3obfcJdxPIsqw6oyqvbryoAVxU0GSf8ODrOC+mn6KUlR5L
m8czvx7PfaXLWA4RMq7dO9IPke6AJxltZBYarrGSEKYPCFl+bgDbUQhQF8dsqQWK
3+w8GlOU7qSSMYYx1m41jdRUTH0yDLksagF43JU+Bq6zqwQV5pOip4Pw/fB0iO6B
qd2dUzwNHYBJrkfdTDUkLjfkEU59AMRVbonBS2Ra8vaZXAJ+X2oKeTVdw1csaTl9
NhPsPsrQ0ZSkqc94VqVkdWeUJvt0DoicHRvD+5g7d0WnkWqUZas7tzJhZQ6T4s0x
d6Yk+kL+544oj5cWwXXEBhq1f+6G1w/2l6nElzl0udaisHNJocICEaOnL7rgLHT7
GlI1QQJ58JbzodQrWNpIyjN5Jh2xeO336Ho4iusZ6QNSXgBL+gaMuuWf0FOoa594
VSOfKZt7SCw3txCYhXagQuPuQbuEFxIuicrq9gC9+jTCi+ZH+XFTcrCs+hcxcv+m
wuOseMhOEuuW/HySRGu2qhJ+XkbLKIlRHYNY8uXKIAu4kUPvu+Zd8lm7xnEV38y7
ENcrnTqwFhEEcUT7C6RaY6kLv+pd13FslwgJD+wm8prrjdC4hQ2mwum3wBzUi7j2
TUoAyd5GSX6D/9h/KkyU0Rz6xPndhvwQ1M+BIUv4e4A7822+9Ky+pzXPZu/gs8p8
M/a/3u7uQPyasplGJsDSzdv/ZMelkMGsfulFs5E0kBCnwWnqsKeD9FzS/6OBUT6w
tkINpuLISqU5sobFV3ypPCA39hFmYlCBQtjdWGHkop3THkdwU8LnVPJJgEiqwPHS
J7AJvoIByqHgRCtC4nwiAMg7hf64jgj8/RhgPhVklvuHWKeFqbgO7kLuFKGolFTA
XEQ7aJXJhwMAQIIG4JkxFdFY1zH7LNDsZajCCtUBtqhA6+WFsCBk7pXB4emr2gbs
SGvgqwYkw0lGY5s/7I5fERyPtDdn/TQjEnfx2n+OHpNbc6minM1yinmLbwqQHy35
kf5dyCRLCtX1zUDaCReMjKv/QuH0MlFGBujeeksS4s8CxBc7KuyYOmZWUb2nJnz+
jdL/9RSXJi6ZG/9QUOdQb6N9u4/Pql0hH3PFifeHIW8hkJoo7fRjkdK3BNlj39po
Az8K5v5doxhYKXM8OJoyK24/Xe4wtroze8tFEZ1YE+mMFpb4amcZBUaVy7HPSgoe
p2e7DLzvpv2uQlSGCjcwHIuQlwkx9M+IdLcwQD5omfWGvK1lKL1CasgxQCrYkAmK
W7XbccDAqZO+bkn0xuwJegE9S1/ZTzvucar4ovPbS15TdWgmCz/rnMNP/1OMxj1z
4z6cMR5gEr/NBsaPheY2YC6htMJKa2mklXDXg+rOmz9OcIBE8l9rYjMPRm71QD27
VNEqcUlLuwhk6yvzCH9q3Vg3b5mre9iaiUZ4hAAUkrLCv1tDiaJ1kMowLsUGTA2p
evsBJzdmccfP5xzBA/xakcezCS2TUwPFI/vPFn/OgUZPCuPUolv6BEO1v7LsHTCX
OQ1a42qLPryZFddtQAuAzt8VHD7Qr/ZgNB7y5bomw7uFwsLcSw4Vr/UfBve7u/df
oXkER1ap6nMkQ/BOPJIUxd+44RHMFKtj0ZYPABkGUEuqZqSl3aeKlHmeeeujP0EU
pMlpTAZWjFxXTY305U1MeVjWt0yy5Z7rUEBSxKONY5b0+ZmccK0fpTTxHytwtPWk
5XERMTMeBnOt3qdLkiUj4KH5k41K2sbOxmNJqLWbiDvIILiRXYsHO3N0eRRY0DnO
7LNfXH/MA6aeFOkqYW2IDKHvJLhEwiWxRU7EmrykDE5fHJVQ9C4a3JvQxDxa5HCz
9X3IL4gu8MRxtAVV2z1Pq5AFb7eccPttIqZqKvBbDoTtAtp6reOXygQyQoChabxY
k6iV1xtJ+hSkEam/ppb6ofCZJNseYN+ANh1rMMSXfRKPXu6dlDID/UFpIHeFTFR+
/f6w8nzVPM8b5OuVmPdbt3KIakv2bBPhYdlzjoBKZIXnkHYbJxzJNxqn5XeWfsVY
DHlwMiWacPr9rrLfOyDlbC0JY6495061EQjJjx20ulhfiLiUiyA2O79DFxuhmJ+M
JNw6JIYf+bFSnbNKNDgbCla/fZrHSGX79b/GZe5xO0rAD9Nh6PpVXcqOMFKx5y2l
iVmY32OYGZ/O/EPWKE9KgJp1j+dHawp6MCepV5JAws6Yyz0TiTkHiO9ZWVg80mGS
TVqO6vFStUTVZ0sbo+TDxkdfVmKDv0G24Bg1WG35Ncrw03SYmwEatCkildKidlbi
oKYtHkGF5TntpWOmz003C8xcVwx4/M6HdZdubzqKRroqIOY+0Zb9l50ayUhqfgFh
BybQdat8jsViOi7gyXU9Mcq3Iu09MuQrUuf2p+ENJHdXSA1a+unYQBh6iaHF9y7e
e+UgQewuHEFZ1J8SVfSMP+NykX+LRuN4hVZQiILCqw4OpB5kEZBk82rgqCEjSGhS
18+goH1Y/CCB1bFCyhNPD+bpYZqJVVfNYsL0CCEf4S0+u+goVPH2mNeKqzI8xWax
ozsdX/mN09N1DfWF/8f1f1QPX4Tbu2ydLVPsLjzbGq008llCOllfAXeGchQZ6Bbh
7pS9l5a7BH6mzx8zdKD402DjoffwvrT3KeBb6QLYEL+K+Mk8KL3b596Z6WC6ioc3
HYS/EtZ3B0uAfdYQDML6kzWHYQL1gvUpwy6lAfPQMeZybmVptZ4B5mzFxltNznw7
e/2WXwN6RdPWPAWa5F72X8ZJSFughWbE1IoKyVUip/r9wcCuc8OPPrugR2Rztqm1
TcyxSEPH0g5tmw4TydabnTSIrYAg3m6jz7cFK+WbVTWeBb8GOlzDdmJ31fszeVma
/GZ8D/Q4Ab9oi7b3e9ToFdRAR2LMTWDnMv8mKYT/9aHdUTpGL+ljmYCFl5VWPCe/
QedroVeuD71bNMKpWP2zvZq9zdTnlmI83nNZ1PYcK0jbsA+qmd1+2CQstn3RMUpu
M1tMrhua4nrxkWw7Kf11uDeWN05h8xQBqFvBW27TTC8ob8rqtbYUegTdQv0niV72
KtUAQaoPiT2pUdE3TdKFHtUpAJJ+MSSMoRRkuTggzdO7TH7zBjh6De/wBPl8wSQj
9C4s9OJI7DM4tAc4gIdFB9L7JaqtvMuPoiMG3KgniOxJDGPY+RwzyzXIcIPlNObq
EeqvfjWz8Kan7366tJQh3fBIRN0gbekAPVwuI6SvOdAJFOM5rphODfFOJWpakKow
SdL33GFcLpW2UDXtyjffyNBdHcMJQ0G6n5LMnPYzTsOIOvmG9F+ogRB6wxcq6EbS
8SVl+yLaQxoijjSTFiCznILWvyuVaYrxyqeQHbd6NJbIYuJ54yEixdhqLcqk52iv
T4B3lFZfVCpqpcPp2Ezvb3V7QZ/83bdY1k9YpaSL/sp8h4pCh9I0tM7nUEb3VbWv
Hx/T3KEQKY9Du8e6r388cBUnWxE7C/DhF9+mj2drX8ui1y4RdLZ2p/JOJ14S5nMd
uBNc+aC78sv1muwCoVf3Vbvhu/bYockEH7EG7kN/Eq4PAezH1VYuQT19jZydpSqc
gqPjg2Htd2PVkZC8zuAwJV5EhXZILW+rHrkGYpGDDyoWul5i8mDrd4Vchj7ybyXu
UsGexVq4u0pXsswXMU6WpXqUGI09ts8qe3HGH9eDIQckMDRjKc+Wubk236ADif8o
H2WOkljrZh1nZUTYdiHxs3LU9rNx3jtenpNDFU1fwGiGUuEzIxyi4l/JrLJVgvkq
w+7IByYkGraCTiPxQiitWEU/Oryl3OFrBdU4O4NTiJcx2gVPvbODo5LnOXavPho2
DcrWzpRMhZUMFiLQ+dldkifuBr9xXKAiN59FSGJ/KSMC4jg245iFjelzJ2A8S4+c
3n1bDNB99DEcAsAOfIcxEvpUZWYf4PIfm/fUfSAc9M6/8mRr/YAG5Depgh5y66Ow
kr3HSjGhRSt8BvfD19xnsNxl+ZXGEYIvb6os9zMIEJdUPiq4OCFPAVmmQKwUFawE
eOLd9KgB1nIzyBPFdzza8mvgvj9jrXlM24GSNJXoDU30lE3pp/eL2t9ZF4OyJaFp
i7A8c6URMCKK9wh8iLhl/WFb2vBhKwhwBI9VF0VZ/Xk2fO7yA5m4kDmXSvuzL1jm
jBYiF3T/TO2fvcY4UvLoJH6N1FTOqarjUxdG7i0X+ggTVZQne95TtDcRQ6uBuaET
QtZHEnRXkmnhR2HN52Vp5M3gB2EHoJRCId37NgkX3GZxss4401KTKgELDsueqqHo
VAofOrKSFCmjbbz7yVklfF7Pt7DVwIUHOIbBbRoEQDF5sDnYQ0tKz8pqMAdVJLB6
Sd/7KywboGVRfTag4RLabqsDD5k0c3kJBNL+Gl3Eil2g9mGF2iW7hElpcdpxYThi
wnDXl9+RiIL2ZTojHDxgoNhJKwBs6nQREp9MuxU3/ybghStAPtnx8wpSmPeku1pn
dD/+G+eSrvPJhSisSwYkC5smUCVes1DHfmUdcaiVwneCDbv7AqsIStRgQxUrO92I
XE26K7NcL5H4+phk5t2Dx5C75UOPJYL3qfkdM/SasTWeE8mIEDOXGtLtQN1EBoK2
zJPsjx223dqH1YWeVDK+B1G7HsI8FIDI4DEyI78QSosjfoxTLln2Rm9fXCL3QPqD
uci40TPTmweEnwUH0HKj1lWc9osOUBpFsUzKKp6RkOdyCUsVlj4EDNp2aL3fQIms
VsqLT7widPKwil/U6/slgzOCWQ6Zy5sdMFKys5j/6qrZx+IihNBQbfppBrPv+OIq
MW+MXdGBZUZvBUF13cbyoC+Ydc/NvO2ntJUERImEpvfdRpE2JVv5jIiT7UbLizLB
D2mTxSFHIa63e55GeiuEO5TGUxyzlXfz8pl5pVI2C9psHPwKS5irRtEJWdngbCB8
xf6AjaP29CplFSxnIFk5JHIA9uoU6WZXrY9UvDrEfddxH5oZ2KgkOpEyIoDlPL8I
LlsmGkAOqwEVdkti2n6gW4OVu3AIY8eYO8JNPPx8nAvqdH+uVhCvpjlH8xfbd8BX
ALMSCaVMVoTOhjUh7FTfRfTTMC0bDSBu8ziqyWAgTWEM/n+ADb1/Y8lVP6I1oDN6
/U7CMNdb2rAwcO9SMKvSFUms9xKnd/TS/9COsiYj9JsChAvQg9i8XOndAdHKk1SM
UA4l3/8iXOsjcJ/rSROWgDxt7mUzt6N3C3NW4bh28kZNuUXqi+lVu1VMO9+iSvHH
3k9eHy16q2R5RVi4TCgrnmTBjDqTVwjAKsgNSVQEs8PZuBezGWGlBnOZxFegXMHz
OgRmwpN2AZi3UtMKerDkBZdQwGV8+7lhxS/ZUbeTlQRE0+xh/pCH/xJzMnk0a0Um
HtDeQK7aqsFA4BmjbccRJXeqFLyk9LsC6p2aDlveTDzL5AZmbyVRiCIH2RNyU6Ti
nd/3/qHyjA8A7F47HxUz2csvaMaF/hiZpjzmoBD6vj+sryF1eXOhWlbYymiPJDww
ue3xRLAaeqH+kvcgg/AC2QgzsDTsVzMdfcXuLRP3DAUHzJZ8+JZlLmUdVOYxt9Rg
oyJxJOafFPry4YnGJa536Jvtu95LHAzis+PS78RToCDcbaCGvN9gbcGHKdCGyd6s
JQJrGv0eTnkK8yS0uHPt48fDFkzwW8wpqURxt6anKp4A1WqpNJ6Ir616XnAzq/65
gh6I2lwcIitudSnPgL61PTVZN+2E8e5m9cXNAjZPMCGurZFYmxNuUcWglzJow/U+
afnrX1ofL2T7oJ66kQp2BvnmtFkd0bnJXPlo+XvA2ms+xRkCw1Pli0KkRCIOjNHS
DVvXZJZpJk6pOLM4ppcZdbWjQFuLlaGBIkTHvCqD5/itgiKRwxbiCWP9Bpks0Uzz
jP7VmWO0vfvYlc6yTkW2ZRO10wYxdXYOnXZ6SOA3xVbLJkZtAZK62Zd+N6T4Ugrs
ACIyE7ov5AmMJpVH/jebB80ak0tEH+7R+YVKNGz11lXxV6ZifBW5Echb35noIS2g
4cFBoXzQ0KUo7ZgBiYLo1MC6yAbXUk3fFa0BR0Y5Z1IYHxJJhR+rGeSqtZ6oqvjb
GkGrTN7DdyjPCLqJl3Y4aRS+LdiKqbaxye4oFvZd7ctnVig8Lgs7LFF1rI0gwcE4
njpIHAttmaK2OQ1Ac1RfGQA98PJd9EacKdXoevgNAWMTiWRWW8zDfuggBwppQzaL
vbFjhozyRD5LPESk8d6hjORDqMiEOkbKnpOHATHFJmSqd4qFGCjEIb9C/KYmTdFC
lGs5D6dbx2TzB6vFGgEuqrONeF9IMwzsEQypJvz2TGScvKeES8q/WptZ3OUNwtZ8
F3mk3RekFKdnwkXhO+wAcSj88EpA5SZd0+2zvioPvYLqn7c/wWaaLCkpQAEbXI9C
tk3p2JrpjGfUMaCbVd5JS16F/w2YuJLI0QNPrg7X+QAM33P6PvsBCS/McuhKbfI+
duLgmh3194a+FxL4hRUJwAsojFj08XLG/bimYFm93JFyHp01rbW7+55aRLr4YmzQ
ClyzyaBYR3PK5v3CIe54QrMyr4dMOH120aqwnZ6RAV3S1wj2Qs6ZFRqBtbAhmxPK
Dya+0qH/SZKOr+dmqONE/hmyBEJNe9juS8yf4Yck8M9k3x6x5o79A5tyrM4T4rjU
GKAykU1cBZbGVFQs4lJzxzeV2cGfUr0bOKbnhZIzj7kPrCtCBXg4c1yjjfnYX0N8
rK6KvYy59rxuCyeEk6mrWDrqkPasafq9D7wKBJus/7TfMq3F9iJBnWf+VyOi8Bwv
8hj540ORJb215PJ22pAiaaUW8h6+2zgS+jZSTKEIQI4lo8ELbAd2sGmYxg8nekd9
WKBLn94bpK1TnlUn6zFskPuRRZ69ZJyd7S8LzR8z5WmL5iLtv/jUl6flX8N/H8p9
Ke+LhJWgwWBbXlsm7WS+dmYvQXCObt9OFgWTbtv15pKa1733kVF5YG3NSbpwS5VV
waqjERI7DRQcogS8DfeDCZsuBcLlAfqL1CP8egb4x52lOZwE7q4BBFgxICcfxkao
rGkOwHMsd0W+6EgssJ8jRm8DHn2S0AJvFCXbGO8yTKbDIZMWYhBRSzZ7q460CVDr
1jhNtQeKUslM3lE4Cuyd56ae+Mrk9mxZHkrpu25Ko9Qcp2fX2pN2QchRFPSLeht0
TYyqwONdt8pURU9eSzdivf7SaHCXAE2cV67bZXjZ0BUzDKEK64xkBe36bhgN7ng/
IkBYa1azaE58lmbHXQ6R7bu/GRNgv3nP1MJnn/oOBzs9mvwOBcizWHanrtz7pV6/
kCbk8JneXjmgdgcZ5qP/j8qYb+BXVk9IZhqxAcCmLKIhp6DOIqLlnCBx+RHnFxB/
pKwR9c6qA6t1cJZpqbTqSuopAcjGfFsev1aQvKUyjCDoLfFQuU4np1i7n61PHLob
dvHaq5IQ/xINUhBdB7jQiCFBtrkvwew0DCpwI0IW6WiysiJOD6HAJJSf12svqcVT
jryo6kqCz6/ghOFTWpiYc6y9JA05SBEn7hJSO3cFdANQDRhKNUdrRb5kjIMk9+iX
mi3wNX+11j1rJS2VC2ZA4ykpn7MTDXW75ar28/me6uNGytbg1Atg/lYXasl+pihD
vel5d+E/boU8wm2+ftxZH8JryFQ79F/uBACr1Rg9T9/Tu3+CnYQOUyfDg69PrJqf
SRpycMjS9weokjS3rL5kF5rBSFNllJEmLrdZ5l8vG6gJ+uGEAZO+vWnjMB+fcwYd
R9KAvomRmjP7ifnHc0Rv1K62IctZPxsXuG7tIJrpIiWpbAUlOKkh6UWcnEAG/3UW
nMnRPCLnmTy/nUsgs+lhOv7WDo37OoHKpVMM7nA1PXPVDSHwNCb5bIyIerS0jSz/
VpvtrZGpcNuz/zbQAGmim+aGOz2LupFnlrgVqSjkfwA5gqQUNiFJBzCmXmut9hJn
Gr2IWDw+sFVp4HJH1655+7jhrMzFt/fQyQaL1Q+gjR57O1kIhE59O4txLyaQXMI8
hAUBs1WszPA/mMZKeVfE5FTfz9xCA9M6Rk+nZ6tnt2eAYRONS0oiCtBPtYEel4x1
xncSxRO8XT0XyllAxuCtosA9EeVCSGMMkaFNoTnA0giWHeL9RURfF7bQ/93hA5su
wRQsSZjMQEOdZBLtt9Iy1YvNosbVAa5OGPUUSAL9cffs4LkzbVJ9wjn7tF54X7wM
7aWGIJZkIw7IX8MqqH8ItUokhGkZP5YYa4P2KHsBU0gcIcn1G5L0Jn9/HoL8ZvpX
bvk4dkypr6iy6x4sAwfdL2xge1Cv9DWfw7JI/8184fiCjbBTsewM6S7vL4CR1OlK
+o+h8LTwdYifEfzqbsznAENyKaTba9FN9fmOq3ACpgWJ5R2ut47FxjPfIP/MCmay
NmsxrQgE4jwbVI8QoTwmH7d45wBC0AB0IoFWiiydg0Wb3NDgfrO9RA3IbCxbn4KZ
MSHAUEr9fQ+BhOxAUshtCEMstNUim+Pu5OfhOwV4I6hCPH/MH3w8Ugp3fXRRU02i
6Dnwvu7ifWzrXo3/pSjDyu4J+Xpc64ipQmDxPuKb5GxmlKizrN7twj898U+231xY
E3TGlQVo3PfWWyNDs9ENlgmrHEPCgXW1xf0CPQoyj5oAWLdMwVw5REFVavNm59iL
71utnfYWSHxg115CF9PSsxe3qm2qngaynLtVkVkr9L3BDJGfYZc0SSYY//Ns7YdL
CtnGsBNEZTquI5n/KUrnsgVG6luWQAlAwJtrJuENpf+OYwDtv7jbsPWOJ19pBLZD
TWLhcP/uhebRryAROkjfjStsO0jjAhz953hGW2BVgnVvZpcYCYn5hihjuASk49Nd
wMOhMlM+cs8RzUV2wHxJM3bh54N9rE45CVN1Cs//9RYyDSTwrZWhOzkl+OotFqh2
UwkCv4ONwBbGc3xS5FCvwAFCryDE7tVNdbd9kANqK9dNPAdweXm1fDeKXb8A0Ile
kwBXCNd104mm+7FL9tGvr9UOFjZhuv5sgoF9x/YWk9NiunSOVC8YFcEDXgpjtmi3
aHG6cuwZeRnQX1bXZu34Sw4jr8MeCbOzvYWY7G200PcI4P2mHHemjA+BafJu18wk
KkW8WZhS5lf5PCa2/jSpR4AcfHu6zOvwD0bgj8LnPsQxhY0tCtGJHBx6WsBa5+NZ
5c9DJyryz0r3SB/kZxfwzmkJdcp7CCMaEP75u22r2aYezCT1FygSM4FXFwChxQ6E
ivGvlPPkY5SqAkfFhLhTUPG9yBiaT4gIOq0NVxe+4TN/M2pOjbiHtLz94YA3aZ4H
jU31ZyhwnfMMXAMoUJs/PvIFdRXsiDbeoNWpvdJoFikijplMy8yU3u1AFoiX6/GW
NCZorUF3M5hGQsophCmv91HD/fKau5FJnuQfDlX+Ex4RLcUyHmdA6X3ThSB+VR/6
AVt0d6lnn/cAz/zkazBUdRyMNXezZEa5w2+FzE9ogA7ExMjJ+OGcNU/qLhHMeV9c
a0wXAh2EyWoa9xs5WMvot3ZI96yA+20kq/f3h92Yuw4FWfJ1f8fU7/5ylrFw7sHr
m6bRJFx+nnr77NBvRS1dTzK7qyy/lCvj3HWo/fWWN+Zy7f9iSqjPuAiQZ4yYevFn
XvvVi6Yrzcn8Em/9HamycWETgWHQWVZrLNQJAGSBwDDs3JHiuwShbcdUdGwtP+AW
aUUZ8HeBfPtfulea6EQJsA499DmJ6gDQZLI3KMLvKTG32/yJu6q42tIkEnA9B9KY
d3PRwBkz3aheUEkYG3HjzN144mu9yshyFB6GrwLMErUKo3DeNRVlIKIxT585JVlU
n1qTEknvqD4Yw4blrb05sG20jW/nw0eFOLAZDECZ93yC99Q/lSOlvGuDO1xJ5PUp
q+zeDIUkiYIJhINut2tV37bT0DQCc0xXudMu6MwqdeHGBICquo/wyTN36NHa1LDA
6xJHEMsJ7kjYsRwm6ZukEcrAJMNjmLK4IPlrwvF6ftJ9rmBxWDDI8INMqqqKnd4A
Tn09pNo/PPNTlSIjqNVdN7l/t9s2E1SBWFRSNSqlFp8xom/sBwcd4JwCwHnYQmjN
kV1K/VBEupay2idPEH53O3kGoVkLyWH9Ig9Nz7nZ1i+KFRUADCHYKAbQD48qKEUK
RG8YDUcojJn8NvIKf+/v4KsMr1cJEFV1QM7ISQoBT44ZBDD1ltvbwCxviFdBck0n
HfWvATBAyBdkzEQzT9/igzUwiAY6QsG2N2kd7CwzrfaYYoIN+1t9EyNa2TRX0FP4
Aw1zCc5QYCER7LOUpE7tT0Xe0k3qR+gWeGPqLSho3NWTP7tJ1vu2OX7UjU1aDtNt
GwXCtOyctK8j6yHzZ/uyNm0lA9sBkO+fvTBP0/J/YPAEU6LuDh7v7fQvGElwtLRq
enO7snVjMbA67fkp8la5eAs1F68WbyS5Gzv3eLGdGOI+Vn8sTFcRqumOwyieUVHb
PxmkEEVuB0T6A4MB8yQ5+wwUMnkdPXyU0A5m+js17qyl7s0hDqBM3dhZ/fpnhHKL
NNtKATPubQsc8zedFLzJ2Kp+gOE+BqKfWL0yp3+EqQ0C9YfLJdkBL5FjkUIp3yrK
YCXMZmDSgSSq7S4mfM/EtlIzZ//NKoL/ExFpPXLbwb9x7t/ydal7ZhzYrGtDBhLg
nKtZ/Y42AZKYP7etfim1rXWb2xOTYCLRc1QOI0pY4k5yD4yHk8ne9fkfyGSlIJfA
hpNWPqWsXPUba3ScyT4qzAvggssHkpvVclKKFRfCG9G75jXZj++kWqZ9OYEKqyq8
lCkL5wYzS0BvgKIjPEMkHicbwhmU0WWIcrnPdYaJPq5ZF/m/kLQw3gZMfh7aU1qC
AfvFb3aMnWFkm8a+L0nI5EKt/hVaHW5bU2sF8p2G41Z5zH7TBco59t0jw6+Koks1
F4pHCeca+aan0SzsanvQOs+wYwEMcEsSv05ZWiNbTK4A1UjjhSQXsC/0ZkheuLag
j08YamBpJLTTtZz4fLeMfdUkJtuuDQ+KvTb7vmjUEcVx+zht4LQEP2o/xMtw+RVT
q7kTF/5PixUrB6KczSFP2g9xbqZ5If9leJXRG6eT4vR+qUEQ5gjj6nRuF/jTPhk1
C55CjIHJyxELRw4kzj/NEoCJGhrT4g8aAck+ul1nyOvQbszyR9yPLZevJM1g+4oo
zXoqGVhws+S1EvaIIa9Vs7ucJCIRj3xwIqwA54RwGnknWxjXc0xHo1SP9KDPBoQK
ll2EtXdpNuQ5+hkGFsjS8t/J0RU2wkN7TFLpJxvdE8qkzem0S4w0HpYtbnbPC2xS
YEhqnAaIhjHiOv/6ljaJrkNBGh+Hm/nudDnKt8/H+xDNpsr1qzSgPf/vHm8nymr1
OKS8Q8zegiboi09T1uVyd+2r/cIIlxOYNCIdSPL8OYC7tdu3GljlaaddOKz4ATRs
61gDbnZXQ4/GKxmN/L/IeBs6/BvQXyRZzpITQUq17njA0n7se2Zu5eoi0oTukjKe
int3Q+GlCfsQ1G+woDdS6/utOqPepoonfrtw3aAXc34V7mM4zhqjhaTqYXF1ePGr
N4fhDsIFb/Kev5jfPIzdNSQVTvl/5s+zbENGyhsC+sXR9PSn6bQBzhs2eeJz9zI7
ybmIKG7pHbOI1NWb41xZTzHbOC6HUi/0hXJHegk4M3TNWzZA999mAoPA6lFMVfqE
M7yBP13mOBq4jdkUW7oxaiNoHL9eaOhlu5vMe7vJTrSu/cogqG4aTjGEej7czi/F
10kyb7anpHCCf+rEgo5K87xVRGoqCaw02b5Cjfddp8XVMtIzyA4RAuOPNzj9MVmX
UCWGpc0+G0gOf3YuW9nY6Mo6OVTwMQrfekDSRJ7/Edwzw8jdg7OMRY9j6qxDCk4R
yAe/O0sa6VaGOm9AAK6hHtkV444+Fxp2anGv4yJc+U1e506P/77pUe2nGUMQmzLS
UaoLK8dNW3b4nZtjpEINRucnZenrwFwkmyuZHwhOZYGJrxcIiASGJTZiapbU+uVR
hrncJnKr1F8DFTDDVTLsThSgWcihaZc/0JM7nthLXycevBPYpNqJhYmnuH28AxIP
7/Y2Fcs0N44OZ9wW76OU3oEwvx/BdPihQhfc2+3FzAJhYeABT1kMwIIpVEgZZyO9
I166bMpWXdzbJKPxSksgp1WrPDpmCu+y1FAW1JJs7aZeW8WincA5JO3VPfWj0inT
Pd1SEbetPFPcwfJC0iQBujdpAmrHr+mysFiEi8J7D2BTmuzYkESsDH24pE9I9Pyq
wdw2sch5NQA5zNNAsGy6u6W2AQh955n7cFjKISteDsWm3+MCy83mlakQg+1q096b
EpdZHrN+dh0nhuIyOWzmjWGRWmpjH/tecV7pyQihOX7y7O1mkmZP79oRYDDVKtK4
67XVISaMKJZpCZKOs4w9JLlDWCEedSJLfQTT66YMQRCSjodsD02CR3bL86oaz6Gz
2iDmQmKtksDwNGZ5BUQyE9o/p0DCvP2Cax1+KklwX0pKh1Vi2/6VVnGeBp3hdaGO
EUdyOOlUe/lzBphue4xvNaCoewBh84DyaFUNT520sn2q0Y2otrq93TPlCSj14G57
qKKNrlAhG7w3ATwvWSfoGCENzGyAuW151vY53zgK58ZHpYoSu3kjLNvGiqxMyV/4
89YfAjNWkYVcWOTjX77cJpIZuEhXLOi0svkJrvUQ7uLZSDazPTVkTRgB3HoBaAJk
j8aQPcrYZx1m7Do2Hc+Dz3ApvqQtmqF5JWjGzw8n54npUZ0rOJeC28Kb5a6tZvrt
RwKnDkweoUoDhUduD5HtD1shVmfOwHuURKCKHGgLaQ0mRcDVBzToWn7MEC6VS5Ns
zwBolTyU454NiAE1g4Bn6uE5o7yk0L7RRgM1/QFEn6LhRtD9R9gn30101tFFXabi
7rLcgjV7p0KqONi1Ionmn+odVpRgL4M9tv9PpFaVe66Asl7TKT6RR+0Y6dScF0/6
vJqe5FQ8fFQMHmOqqYDsZgmG7Pz9Oiuv5aQgXroVvVLF3RQC83QffYftFJNALPFN
AruEECogppOJH6MbPi+HYNLJ0s2jeNHRk8ni2UdiadGfGRlh3bpGWkHOGyeRzY9t
qUAgs95Mxk0ejb04sAnKzdmboGI078glk4yz6o1fSXDwc7ZcsSWdXbPS7Ut0O9WO
i3pIR5k2XkUs7XHr/wwjG5niFZL3b06x+igDt0fd3Rlz0SZiqKzZFzPQLME1DEGI
WRzSoh7lATAt4blyFwbd7BZkWdXoEREMKb2f0TfbMPeKgzRlzzudOqsPoP5Gp+Ig
npjWyyhIp27141spN7xkFZCFSMg142p8YsD4i+OPnGJVhmSSFlonZU0bIEKhSs4e
/H/8G0TQmhKye1QPELeCUUnTNPcKIteIxfREgE8Ja4K/fcd6qStI+x2wR71sKmpe
9tSQ7ytCk5HVoEuBVQdHa1NajXB8YSVUjsV300z/BkzjfhW7liz4kqBuDYH9hZT7
5ofdKQgtSrRJuY78GjQ4uzioWToS+3hxS0vgWrc8RQggrZLO5X6n6+TZclG1xX0m
oiJhu4Uj7myiHqFqnxrvs/J90InyFU7NSHNTD3h5qUJIjNERPzB5SjyxLwCD3Wsy
fOK5UCdK1Nx4bFjZX3jgBbho0osWdGKrcObHWuQBximulV1iri2ODM9Q3X2zWP9j
Z2MExE1DrQ/CKOUi8/fiVrSiJ7NWYIIey2N6qPQf3DstInUMIJiMIZ58+WvIAqLq
Da6rXPEXKHeDKPs8fxmQw7BsjbH0+1cTZ5pUASnBkaudAJ1h/dnxc8DGuEp7ws4/
fJ3wm5o0+UjinYSfBafu+BJmaPX6kxrNHQnR2GJdM19ZlDzb29zihOg3sKN/g5gm
uhsS9pIfSNA9prrQWX/25v9zr0ikj5AuAyThokMbEH6rizaHO8d4MD/W27Q+JHmF
zL/OVKsQioGkBzDNnAnhyNi7ryG0aB0tMkmkNx2AXqfzxcQIEVNwhGfbG1cfm9xp
qB6oQ82robngQrnil/6vl+kgyXYf68XlFhRVGz4yllComJK7xgx4lRMl6EApYCoo
K0HwZn2OefY4mVHYG9QelKKnX3jk0niDOe+DRskiodpX9gSTIIeqSE0CXmyvFJew
o/bMuyXfGQ7178Jm/ippd3IvmsT2kp3yE92l5Y8kEJsWw3NS//9aWmSAGVQ8WiWP
Tq/2ec4yvnuUuJI42KRpm4n0YlO+koZPbIllk6H/lrA4AX+mi1pIof3DDFD6M0ev
aEqUwKCdnWx+vQsdE25CO36TKrSPtxRpjJ2PIUu1PMA/MucDbaJaAJGeQu2D1OgN
C8IXf1fJclTwEV9MRd9yD/hVHQkzzzmaXDQ6F+PM+q+Ny2ETUZsH0qzY6Omu129R
IRlshV+OMFhUUth+j03gBCMXO1fUd0fcQ6P2AR4OZyDDZRv23i+I75i0FxH5HvSy
NxVUHFoJZHzwbYYsmMqnXiUE5JHYKvWOVbi4P/OrpsenpYswlWzLdn5wtXejSPdK
4MocY8FveA8X/9oqAp9kq+pv5Kr+eYO06xmmnhg0loGixjHz0NaplyACJfh5lUA+
QpPRz938ET+D0XzgZI+uPCz/6tkihMYpfE3RortHc7tHO4+Gi3vh98FBS12XLzoE
OTL8NVwzQGypbYmnZYRdCnB7V/15jb5uTK6zoit+KqW8MXUN1EmUrsB5ZSRLHBbp
cvOgtNdwDWalWLidfgPHY2vmQ63z0Ft6dn+YIRISCiEgObRE8dCixbyOv38Ov5dF
eOK7KAOOVBxbsw6lf/SRnZMQO5pCXxnndx/E9AVdYYMBqd6HnVfVscP0mY8pNGPi
rz2VGRyrPCkWna3lXNeeNeSMYVs5rjAgnDhk6lutPQcSa0qR+APVylEfxxPQ9qok
yuLlTJjGZQmfC9NV5LcmyOibhymdQR8SoJ/GdriBzg2bTFAEMDA78kPV1l0Li5ej
yViAqUGsrZQg9h0oMPmcdl3gOhi6lqQRRs14PQ+1o0tX2A8RR5/SdJvvoTI8i0KZ
x8T1xaopdS9UYiQ/O5grhXq1/qt374fLc9Evcqj26gFkEisza/xcdSTLWHTa+jU2
9ffjC0lKx0GPXL98SdTUh/tjdMK9G/lENGJXDFZdJqXsQSyuW1VrAeEtD73HiZSt
r+rhl1hTVEnxLMgVFvBZxszrgXdO2F60pPSAFgbwaAfbJBMvl6GljRzkqX2BRZ5U
p/7vsEm/FSbm8XygzxahW8NbYIIOoRi8ijWtr01zf3cezVLZRwYArb04wcgEzCrf
JtBaZ1huSpZ8i5MSumr4RcJ3+zcIpjG7eF0p/FcSaLVJb021AliFIgLU1gcHZPqs
Ft9VLOVbO4QoWFKr1qdEO3czXnqoMU0zO6XmIgYJleVQ4XC30JAmLwyeoPt+b+U3
Yi2Itw1E/FklXM3aiUHcWDoJbTGypmsG/01WdhPHfRkX10r5aKzGJ+TogRLhGh86
GiHCbd2i4jaAdnnwIHcL9g5XXNFMhWk8I4svd/EgQjlaIT38MpIZeYfvCz5FkIZ0
4SEWAmF11NOilVFqF54jWoCT8HBbN/jgo+3q9gKe2tAGSj0cmR0Ax1w9OjocZ/Ra
b+wRRIhu/7xrYaQTI3uQT1tgdtjYLS+A/bErhoudz+b3qVXV4LukEGQ5y7F8SI89
NON87ti0Fpx8gOLEBbYNKKy/Kx+vnX0z7qNBYKAdEB0DIz0dg2HpbP+ggpiP5kdi
03iNoYZ3fAsxYEeC3RzYlUOnSdCjIeob3THueY8WoGWqK7RUu9F97p9ri0v7hhAt
WDUWzZZZmu7Iz6pGaB5ePWHePjDlHwlGWnRKTjAeGto8x+qe3A1hMNydl+lwsc12
6XgTLijCcvtaM4EgozGRHGTKSBxObBEvQDeR70bYPgKKscJFFlexnAUzeRIn+f+5
40SuvsRtHH07yoHYZczyetm1wXrNWgGxKlXKu5tVrDi0H/a3eL25AcRjxr7u1oII
oJpa6tY5P/H5E/Fpn0Eqz+jz6xkQ024u9oLdPuTZOIY+XUXFVFynWqFjEa+59asM
jxcHRNOKXtH9rX+UMN+SUOAh3eOK/zkYDCdzu0m6mxWcWeBfm3Dz9OhZruMtk5Ms
zyWbooc7R51bLCHf+OPjQif0XkzSl4QQq70vgARE4eqzLkgzV3OOuOHLg3NqQCr2
8ZjOiMiUXxIl5y9+R0TyVVbspQUucDPZdhulRDk1wyZovIjcTkKHL4Wpfnm1drFa
JfXKln0LJEv8ksrRcz4LJu9o8s4VIQzn69w+AB2n9hTKUEa4RRCNLyhuAtm/9NsN
icmOWJsQLpsMZJAW2S/UjmimNSsSAoqYY4u7SsUvg0BR2HmoKbtlFxja1p+gJWCc
zKXLuqJvpIGSd0zYUs9Fh96DFg/uhBoLoDdCYxn01Sz3tF1v2PZRuJjyK9bcKaRe
Sg8f+2OcU7crTarCxbyyyQbHRm6TzwTbKW9EtZFFNWqHt7TFBWH3yE0TVdE4bDTd
KfM8fKPxnGRESU8pDbjF5BGuE0dZXebiOKltCy9pFE6yw8WEdtIg9WD2AedQIYDb
DcpRHRPs7hwcOtMmFnODlUTys3oXAXIumFLalSynhJTg167+x06skK93OJXlDVJ1
TFhL+OqdEOU6OmQY+wA5hrKUajzjAkcL2kfMoxF6kPP8WkHTFu1HVWgH7RRAehQR
4QP3JL6Lkjdr7edyIHMfEjYqsAMauceL4yFTSRplFCGky2i2JQ3Maxov3G72baaV
9rj+uQdwicVowiW9eazzGcMF35Z5xzA+vltFYomyAAo1HXqRfVyGV6C22RPibX7b
1T0SUTbpPB8qWDgCLehoE739wnG4NB24QnjgfonW/RaTphPRrd1qR9IpoP4uky1D
ewTdhUoZZAN10zQkk7UTOIMhVf6SXsnEQ28gKtOmdkpKAVbUTm2BvfgF33psOQpa
KLStjDSp2alO+elFotGpt8TfyxFLtdeLdqgFfn3Fv6A5dQfDJmddGwmE6EnlRqH2
MuwlEeIlCMtku/FFXIGqRORn/nqU665l9PrXFM8qKlkXLksvkQKkEWztFqW3ZppQ
N4Qw8E8jR+y2nKwL64myEAKr0G37NDXppzZMXiP+k/f9iubcrE+oszogfkPrbfsC
z1fLCpxugv+9nOw0gXE2Oaq7VMsq13Ga+s4KgD5dX0zuj26WTBpSyqNp+6bzEXQ+
ptvtU+ZHFlzgOjaBvTv0UVmBCNSNA1liNIHtAtmvbUK+txaOHSNfz259lG9uNdIY
es757zdZqCSiJ0rFEKFs/oitJ3I49TaXbvIzvGTN11aB8H4mde4M8F2ghdEmpWfF
3j/ArXiujY34Pha0mrqnNmwRir8h48NfvRQatc7Iw2hnWn6LHo0atHRh7FQb4dvD
mycNEyyCtUrxYqReQ+V3bLt1tVqaeT8HHb60mc2EfEmbnFKSlWDrDK0Aw0l5HrqY
UIN+enT0YcQCXTvMqbKtV6NAETZxS8T3+kPZIbifKV+nkzWaJ96tYkfGqDG0OonJ
bsIYy5BUH8ulzfU0EIim+f5Z23FSpL8/6rXu+fMiYuQ8T7V51/NOg4T6ew8Riwg5
eILOyIXKcfH1iEENy/v50pvS1+CobNcduw2dp4Fbntlt5M9u3rm2HTYQQSFKv/BE
9IjQBlHprPMPGUgrtc6Um5WSSQGWjyzF8Sv15TW7OuXm9hMZXg4XBOAeD8zCWjVy
sqRIEHqpzflUznVIjNFtILnfZzF+3FgI8B2+tp3Kfvtx8rdQbR7B1D/UZOfwI0JV
fGn8L1WvpN7uesu598XxbjE5ufD/DgzcRCpW0EcrbF8PkVNtkeVkjNbz+9BWGr75
7CGxS44ihanAXcKAokCeKsM7cXG1WknFKCpQ1l/1MC6GBC3CNzeZD99Ta3mprEHI
NnF7js8skZtd5kRnXOOUKWHYBrrC7xR06DeKGM8eiTXjO3hnkF0WI8Y+NNVuLtJg
0swJDPg7SAXqeHVsZ2DwiHVKKVEom2WGdYYoXamGZOXeUfwwGDAymCO2Kj7LhMTE
lD5i8OUzirXyxTkXvhwMdUmFn/4dMUQ+K46khgzlGwbYzVe9KLVrRLhk4WzyfVYO
TEcA3hofTXHZ2JnMGvO720pa/YJEQmPvzMFRiqn+mv3HI0LNY41Z2bghHgGJeGCJ
TNbytTgaCRxvm6M+VNzPNCNbZgRVxuWjCOHMZL22VqYWZ8emqgK0dMmsppQmU/h9
uQCYUmmzSGk3bMJZg7vVamdDUDZMpPGvBLYyfGes9JXJlxNoPzI3+CvIOKDps4JL
ACuyP7Vp9F9vlhayMF2C0YeiCTdoIxk2Bc4Q276pspVqqcBubFDcRr0UnZXrX9zg
F6C9ZhLR1wQVGViMPzaLBbpSmd0HAgnRfRjsS2ucLUlGgDWBOaIzYWwg1VAkTed6
L5LR2l9hdQk10RiArNQssleSMJMytfws5aUHeJgIhaTw1v9rGabpgjmgvqluNfuK
r//hJbWz61nnWBi75a/oGYqo0GR3HDHAVwh+Pm1JpYThEtkOKj82nt8unQfVRTVV
ZwUDzeo5TULr03+el6Xgcgz8fTsxxKmGja9ObFT+K7JPwxCARwy4CZ0hiS8Ax4dC
fEVkaXC/tUR1rl6vahekNXMiJ7Y2F1oZEMLuFwQzY4UBgLCqlz0xfKjPDCInjk3E
+5YvBDGd45bHge0lOuEXLpIRRA10r286+BhHAv4YGc0rnMy/E71RgebrZRRU/Io1
T0M5bkwq89r3cbaO7Ann/HJs+0Ztw2fnPB3ZvN0xeJUgmjlKEskdWXuXioAU1s7s
98vgeE7yrNT2d641r+PD5K8foQkWpv7ky7rR/XlwmEnqgttFlarall0vxWezZu9D
ckoBs9roTx5fl/7VPUGXIWfBo1y2VpPBo/LIqQ2rCjXbEzycegCUmIzZUN3rPFPZ
ZSSAekUEX3xZ0IpmEWlz0R52SDgXMGFxeWoeSgTC4FuwvtGli8Om9vt9cpoMFPkz
hI4dN95vS503AqyTiVs7rlcwP7bq/QmpFtS0emZRdYHUQ9gu9aylP9voWzAg3VIF
G1321z+IPq27vONxvRq5cgQjbk1vOK9ie0BqzOLCdWczYbo92Ds5Xxil2jIFu9i5
g5rfNKRbdaIJ+6VC0D+4c/mzmWhFLRVV8gg7vYr1/xAXm3T9Rrm1pLA/h22a5JWR
d8LKdkSACgDlXavEiI4j9L5Ij3d2qAd8/v8Bd1VNtKQt0LMJC8rT8S7TiE6qHjWd
8K7YRm9IiBZV4tpvUaPvWsyO6PQfqpttrxddH7b8sZxZ+S0EJY/b8Pmu544sgVx+
9YnMJwyod5GSG1HNKP4fQIxQ5TIeZurafkT2Gloz59ES4IJGfB8GaROYJYOqLo7q
9KFv0msXfW46mWeIjdN2yJ2Niz3p6VDe1nDxj29YsQybUhdiHJc61lSs4Hphnw/h
gstPvYA6imdxJNjxy8o5ZFnuN7Iqfe7vuN+fAg/TBWTHYf3zX1tppTMBL/Hud2UZ
oLVCCapGijKdJpsSqybyPfc0HiofOS8ySjWpUdm0QrByNA1dH2iWoACEFmv4GTv5
lQ48ltXycL4lRm+7aXt3qx9ZUaBIp3QWD/zHkTAPq3W89RVFH9pBdkSzr6FufTim
HVHij9AvT2tRfMkSOUaWln2eNmNv69DrP6r34lTgfoYvsqoXKMW6VcRrwerGmOh0
xoOqdNKjtqm+4pgwadfm6cs27f/f5kVyfusF9PDlzXzdmplA4TAbc6aDL6pJ6jGK
2tjxlMcrlC+QIsZI1keo1JUZe8loXd1EFc3JkUa7G3TOUrT6jNMya1jfUJjEyMIK
V+3Mbei1FSI+sqS01T0dQLUlRpwXQWaNEHp+tJEN21gHA0TVJ6WiIMy0JyDCjXKS
G8UbFWiL7XK3NwTEZhonUWWxkIC8cBV16Ezuxp6uDpqnlihE2c6WPRzfB2nsAWRx
GINRLdBfxMf4e5ONo1A9+37EWrTtK2WBPX76AhcpDtOQ5ezQXtxR313RHPDsBFd+
fKGdej2UD9vSErn0r8zfIN72vVGd9bgRinSu/3z/lk16igt6M9x8QOSfz3q9ofYj
zxlXehRjWf57Cei/dBpvXvYoC2IT2+l2S6Pb5ZYcfghEHHqz4qoSy3UW9sG74b0c
Kgvqc7xeC/Yc5nPnXqBKiiaFNb/LHBpsFmEqp0e6HDhaTxkOq3UFDn2LRHX/5ipV
5lq5zh4KepaQGRec9iSEJxceYZXB4m5F6+N9R/sA95yFgB8CYCAZ/jUtbzDh6vX2
UWLwPvtfhndjTfxYtCHQy6Do7M8DXrVB0SUUqM3QNw10IL3+lsRq1JqqCsKUjGst
tRsqU0UChryjffIfOfcsfFNQLqjVBJjdALdMbjwQRqiYd7iPssAKj41sJ5bHnVlr
8lm+R0OblYTtkoQ8FDdWKOSkFUQXgHkkCSkeHm71VQCor4sXjf8eaSSFCGuVdh+S
voFi8MyC/XWRqh+RgNVsTtNtwlD5IHcI5yr8yCgtVeO3ffc0dH/wkB7C0ihlf64K
BRauM8VOcTaGQ0D8DdCidZAJxSS89xSg0aGuc/fhKu2WC8EQvVaM/28a5cdOMyV9
0rwKAZhTfAxoqLO7tE0+YeHnOiM/5pAj93YpZzj4TFwaylKiefb+e5r+tUD8Ozve
T0BQ8U7J/zMWksw1+KiXY6pbAy7FvZ96byaGtqcHWLP9uyPXg7fdYd7dnxi61F4M
RwDYc4DP7JkNUk+eTl2pFJyRiyYwP69UamZKxoEOyk7g08EzXtzYnhyYnfGvu39E
AOa7kIxVNUsNNSpJclhb2M9uCtpmlktzVSoNz2kuAwSGGVNUB5sbi/DCKcgnU9Bh
5qc6A1McNugfIOkKYo1oAvI5Byfno+a10oS2EShAaam8LtAri0kHPwbz0Ntj0YX7
K+1sMWilAH3IJ4SQorRM1DO97DAVOAMXso8aAi+0iDs3+IOFPxO32CgozInMx23/
RQv4IJFX7UOWlerE28n+PxIVuUZur1Odx9OpH/bJ+5FntZPc4gnABzlK/ovW8dot
TY4fjCNYV/0jH0tC3obEE/ICy9T+zAk0iJsflprXFon84k5OPOP51Te9M6KMHqL7
OhJtLd4nRId+ISoyXoJAcr5nf0JtKPdV4l4fAvy6VNh4X1iCWd2HFTz5mx8L4zPv
ihBN8D417QOm5781sG0iRyo47Tm2OyGdCzsE2G+glguHwLndJ0adOpvZ/0yyE63W
uLzc6N7Zl6LUNEgyocvCaCwjsrv0ZtuLO+ddgFIPVqrIStBsg8Vyp0O8gfyDtNZy
b0CZKV/n7ukG5iNVGEfr3s6c8X9/ghFmD68DqCwNh1xRXOcR/guFhr1EbWe+o5wJ
ZnNVmsxPeleDrH+BxvGyQBKHQboeBjySSbjb2663Qj/Nmry3YKqRgG7Cgbp56yvo
EMMz7xhrFy8waGbztcVIFt4u87bu7atTqI21OL34HqIf+i/xvZIP9qHcWif8v/Hm
l5ZSff66jEuckWOWGAw5c1+Wf/CF91wH0xcIyLCYqo7YBbPVxaEeqMSYYFKZJSNA
tht+1jVhfSKvhDEGMd7l9VfRO09SHw1JhKbEK1Nh7V/NRD586L6rjNdy0DhjMg2m
PgkkjdoTBWkMt8YKEhFZx8gnPOtMpNgryq1F4o1To7a+oS2X6xUEPk3APMzc1hD1
nNWrgPfy13Mg2Dc8UMCxznDleoamqtLQuEzjPKkrTrF0Jr8O8aKn0p5EZ0MyjbgG
fHoCvLgI9zZ0wg0AgmCjmmXiqnvYxgMC4zmB0evzX3mXcvrFEheDb55R9jluH/eY
O5y0ps1qfxYZ6KL/YmPou3X4wDAcD3aYoGho+WIIQ5n/cxB3SobEYZOwkjdZcOqL
/Ei+RR0sH+bP8PwoyJDpOQAij4rQ/IWnD//cUdtO/PkwIEfgXM54KAPuDipZKcpL
DXPTjWXwzp4umbmNkn1mLxAqgeCeq7UP85cT0JVnhn6d0e7FrbhNPT8bB1Rb7nBZ
uEen0tOmxs9bUL8nmeNPlI5Y5wCJApxqui2740sVFBG08CYxH59gtqtBHD7kPbJc
nHjiqDnqjiqgjGJ5SuiuOxllJhHvvgdaTdLpCk6o6NZTHuWQpFqYDcySgQs95yu8
DXqZQRUk+AwEesXI6bA9vso8GNqBafrKgEoJJuZu3jleQ1/0OS8/SGA9P72iZfAJ
n9ogCPpZqjFLFNLhMZQYegn7OwTMMRywV3xi8lyDUp53JZxNS1Fxi35jCJFy2RDc
g/Ir9d0Db4ly4ozqvfI10MRbHR8hDLflVII92WqIH6niE8XrtpwgA4Gd5eg48JZI
07XZhWC1nuBbYNMbJcRKGUtXO0ilCmjcsNN4yMAF33zztNs4AfHhAr6jXMa7Gx7W
AlvJEy81MhWbd6g4yO1W5dJMmV4ulHlDy/PxOKJwssJen3KvFuSuH0UcSADDdnIb
4FvhSL7HNPDGi4as9ixJ7BNHt6Z6u5aHrscEJrxUolasmiwWyYtXpkZL9EPEtXHb
HoPQ/ujAFW7VNqNmxpjdWYUwTIhSTa/vzIAf1gi5AKFfjzhDYs4dz4WxUbfoYrzx
OV+HRsI37m/H+sXSL/fDNKDfOIF7XL12QQuyoGi459gRsHjorLDzN1tDKFcStH/h
lNiFOcTFkeD6CTmrGFytjwwR6HJ7gBoW4pWIsys0jubNfcWkR39vZyJXPNMviRda
p1EOuPMGJpP68kL2vyASGu8qVaoUNllqEtj6/TQrrbKZ42wvirWXCrOTPdxkI4Rd
fD8Fb/Iawgm2OGK8UU3iF3TYOP7GKVZcnGFEbzuvCr2jjCrujlkqZwhwfrJvltEc
r6WuWXHlgBsWk/M4sB79MyY5oqFY6ITne5G/UwydDfiGMF9ZVqzJRghkm9LYxAop
ftjRtOVS5FIQsQWIpQ9r92VOhrpaR0PScI3HmVB6pSfym9sGNqR17tEHxlsHVUfL
WN3suTPVE58A1u4Ynpm0PQGdZERICvLs6FTYSWuK+eeu1q1/nEPb5jpFiJIfuYBO
sQUAXML6SLsfFSguM9niF5vyoBtaunUTadOAp5kU9ylRU42Uo9WlPOg5XKTup6r7
TXYT71nB3AI3ooLgFMoZ1vANs6rKTDUc24kFlobYA8/hdvVyf/vrp0CQOgwAOs3E
t2oevFXHTVCACyLeWBkPAymwaeHq7TYDPwBwpieGXTlUcQOQd3JvvemedvDhpC6U
kU53tI0BE9E3iaiw0SaLwlV3N42u8NBCg7qUmbMtHGGQtdOi564ziWlEmP6lTWoy
JsjtOYD48LKXW8jGxPvlVSe7LCpD9LFA1Astwl1gbHUlbNXYG7KpHJ1pTHtzgxk7
xPdf/5YTEizMtzI/fZlfinszuFpW0E8WUdpHXYGnvdpI/6n+SgJ+5gxNKIBe1lvk
+08pCN/rxNx+ZRRfSKXSY8BN/OWVuR80qfvjgGrhdWFaIYgwlFMFXW1HqxgGCNiP
Lw9rDMcYuA2nZGsImXwVSFNL9Yl1cLVWPwuiIpzeXGYqoN8LsKP4Gzmh3zGDbUMq
7vBo9wAm3LLZsWmxas/cUd8idkMOPvXhgMqgnZdbGhk3wrr5CzXlkALkIrFxt1Pk
LYtJdMnG6YUZ3nOVhYHm4NuWj+lXaUJVct0bnYRKhEbs+mru289le/pK//eqd8Qx
BAHXSq2gzJJEnQMwbWThuE0NhE3twVRPKQ9+umbzHj8RvXGQF0C3cJhwl12U5CTU
7tRtzBMszAgDPTfoAzT0fO6OhbgjTD4uEz+Ic/+k13zatsy673pu9JevXnvEecf2
S6V6peTpQ//MCk52B+ktMa6HxKfyr43nM2zW4Eb7Q0iGAU1r1LN33Hn8relLj2Ar
22yYXl3JfLaxjxdWkWh0RL4S9ux5ReqIn/1Y6NzlDs8ssUubfTwTdmyXHJZGVmue
RA/ZCtvKJ9aspv5M44mO3ok8epNv9hCxEB4C9kfUvM5MdqHA0bziQO/DtRffGJZJ
MMdFmpNFLq8Bq5QmSzxWZp/zqhm7J5BxXAGT5pFuNEElcXVNak+/+4z7WNealnf0
De38OU4KEyPITeBYOi41P2b5dnXur2rM5X+DRc3pjQ0QbiARLRNVG+Mt9ZjIWzMD
7eJaqVm6PbPf2Xv+/ttfys4aHD5XE/aV6skvzwOHuoHJVtu+Dkp/gZLASAz2yDix
lYkZaVNXcNptLiTBTgQaetkm+lCOt4AB4Cs9ab9F+Q8zEvW10y1sspXAhe8y7DOg
fTwF6kKXYLnQV/+PLcNH7/Kjzlv/2AeNbo7s7ST014vbVNmN5v57eXHTHB6xL6cL
4sKDwdZPt05eWiYJo638X1IuT+42RrX92byTRG82Z32BlVA5Xakgns1XURvHl7gl
scVSocMmBhgt6vclcyY2MHzwBbQiw1RziMQSo0Pt/GLfTtrgCR4FcGOdFiOrb+/S
+tSp4We2BnpAP5C6829SFsqCCxJUC6TeUMUHmexpYk46gjOqGnyM3raJhGP9Sy4h
TgkQ/tk7KZbcx+V1xAt1zeLFgL5LaBJJwRk4MSLnvuOs6J/9vP/E/PfyUeLd3LhA
ZbyAYotfAOTyKU7kFAJsRhIofiLwgO0Y/M09l8uDMbQCbQz5oalWzmfU0juNL9eL
IyAl/tmvb0/SOqcB7cdffsDz+XXX4QMqnlIxyRz58EpPwQaZtqbFo1abYyxOhLbE
cNKhrWFafOH3Rt7I8zGrBKalU66qtxmSd171aqCG/Ymx+ORqGgNc8h7of9vm0t8c
ktNXEotSlDWStKog/H47IZC9DjRq+BEg/C6+OyKrAJSm7x5dsGcsUDFIIJiTExiM
UnfXFAkw6+dBbNsn38J+15VYm7sXXWdZYeEpBtrTXNVWOXecvAv5ECDTo8dFS94s
yQrnjUxy7ckWbfKiJjqutDJOonwQwjGkcgZyRa8PIzJuF9/BGUO34kFbpuHRRLTt
9/jEm4MZz7xANy6gRg2jQGyLlYUF+77Bjk0EfFRqnxUONNazMB/lnRXeOdtO7k/Q
KatVVHMJL1CutnNT+eJ3lCldop/+Z86q7qvQFubeaC2UpnJDQqgR2Xpn9bmoOx7i
Of/F+jv6yfArOFeqVovTPnP/HiCzTneTe5i3Ilf8QrwnsZeHtfrpTtJlHTHZMno/
otmsPqt5qYHAWxGzyVQ4zCbRD3ws+flEKd9a5grJwwXmb8QG00I/52mMraZuJdnm
sXvBdWooQwAJY4Sn4xTPP6sjHrBrPPV/+5uJFA6zwxByzf3XXcBkuwHTVnghxzl6
qkar6AXMSkQY3rT6qvwGFDnMO78ZaPeIbGMBDiaZoTUQX95T01G+6pxI3AzbGnr0
7+GbB1y0XcBShCIRzqlzeHIhCWyjTJTIRKJ6tazZ71/O5Owc7B2mt+N28Y7LB3D8
bzUXWtbDjdKkIp8T2c+Uql60H2L6lOYLipm2JfyPkYg2Mes8aiF5Gm9hOv2ZWGmq
NYns5Uh9sKVD4VQGYKSXBJoiUvWmtZvX0F6aS0o3T6pDUy8BZHQpsw4T30BzTBDf
tsqsqO0MNzZvA04PSaEu2L8JzjmRf/i6FWHrMOuKOUzcnTqNxb6CG+PZo1Gkt/Nu
FLUqnGevHwLoom3sHWst+q8GcE9PX+QfG+z8d/QbEtnZsZTIGEaDX/c3+IDz1Nlj
DyQlPRMtoNbVnwIe+ATZURVsoSuSwoBmHdRQtAW/lV5Oeg1v603AvIkMXp+i0dFM
Df0nsVus23aTJLFlSjoZp96ruDN4bgRnzR+7MLPUxeAFunLYBW07SX2ktNtPF1ZJ
HZ4oT5i6i7lXGVWCWvR2m4xApqbcoe1Yaj5sa+ZwjJp40pHt0RQbvwW8Swoq8Kh5
BcdnUjK48zeP50SnOSUa4dptK6LEVYmx35FAvpcMWiSR7jUR2Z1hj9fiaBvMsYga
fuVLatmm69rqh8zyp0gN/IzjFkZqWROXYqUhUgVv1fhrNgDh+9d5JBJncUfzvn7I
51KQ+dLnD8OOtO5A0ebN57/aw4iXqy2y2iI58jI9fmemBs4884Ob6TXlnThW90zK
qPGbENx7tt4mTkOUUJGegdr36bUMM5cXa7bFTXT+jxeUGg/v+eGMxtGIi/OfHeDY
4DqCHiOlt7l5ueoPpQRN26HNrGjxVM9qZD416VAfdpDsjKps42f9vQtSl6UrJGbH
jW0rUUwY0cFV4yAjiGOezgTycGLcVPXNdV1Qx3RD5ORJlfQ6IZVHrApjC1GCDCwI
32sfbLZM00W6gsoMipqrcDndOWAg7hEAH3Ch1957iBXh9JKnbCr4pb2ur6DuoW3L
GCunPYdm4hobG9XtfF/jmOawhJnGK+G0tu8Dmh2YyabCfI1JBMVdwKbfcqg2S1Cw
iZ4pTO99U1DVi4aTq2vkMOZkSexm/+fX5NxEYonTBcVHyG4O5mwY9PbRIZfPYUhS
RPp7b5f5LC47Mi/pgcGiEDxad4etcImJbr5mmQbL48NTyasAjsq+uZ1kUi3lRJI9
OHhVexkBB7/QIrGSUbKlfBXkP0+5WZk3ucsRu9OFgNN3/+AtXAUdlBhbb9mQ+IjO
QgqME2QjAitv8BZY3g3JhpSHsZaBHtJ5l8pjaVQFuA/ilm1vR65GNGTOrtpCmxZK
Cfj+2vys/tlE/2vowFiX4XyZ1kD7alnqCk3cQVMZ+F2Ny3T2k9obkg54AlGxacbt
3q7vRX/WoSg3ILfHxE9lAGKuqINM6CBtrqXCwiRuyX3ZrjtOQUTreEqUKzEGbdsw
eULBl28ZA7IaKoOA17Xdm/O+ALWWn5xn6c/IPxKwMFZhqEiOafqu0wajAZfFL04V
jpli0ji1ld5l20qrLEY2jpmKh0LI1205VcdE5x6gTyuVZ5062OLSuc1mQcLh0mDO
dGCavrgGyfC7axbXztPq9aIW7nhr4MP2+exuBgVk4yXDaRmHK25OR8Z7pNRD8c/+
oxwoEGOhO+Ud+xE+q75EvAyBQFdz+Gv8RljAE3HbBUE4GHhTqU/2LLHPe+6WWZa5
ADIzU1eDuo3G6DKYjuFPuEVK40QjQ414+MgPN/i4jEBpa5x1NNBlT7feASJK5rY3
udEqUo8MDcviJt+lSf5lVaZGaoAOhaz3g6Tt3e95s1DmCPf+HCaoanG3FBKmDY4L
2rXCgJDNctUN9bFaPU1eEwgkicL9EczOHQ1g1v52rzuRNyL7CMGtc9lBarNVDuLE
CCosVSJyKn1vkM3Rmzo+5nYWqAZs5qORLqRv/yqmK3E2Fd6BpXprKqXerkBg1itt
Dwe2cE7MTIWLaQXx5MCveV9PVjgk5qluxAOQYNhzFoyadaehEReZGmjzyobchjRd
ZFfmU+8ZaZXayy04cTU8yo4G7KQUm38IoSA+nQUq3rx00gG3fUGVvUtueri08nX+
pBH5z6S3vBJvwT0GLzwh+2Upzr+saGEa11ARCHVB3iMHfQuHuph7NN9SJjvO8fyn
gaYg+aCQe80N+LcWM3U7Lw4acU5KW2rshC9PH8P8pb83DaqdEzrPODn24PtGRxFR
k9qE+qSLg4+lsarsrn6jx1qldhQ+bWbUn19ZfXLRQYtUpA1UIB4lZZ1xKpeaw1QQ
jxVdS/pmIecaE8XlV3VOAfMkOyj4y0X6exVgTAmHhDzhMOoLxcx49YtvJ8g2bLb/
4xfVO6UrkjmqkS3BQjo0A3TKbqYm6/H7RE1iUomKnIzIlrUhIye7PKGF8reBtDBg
y9Hnit1Hj0Gxk9a/NYZSYagbjXJDdrASUC/6SJvR2io1MrwoLjbci2ZOP+2V2TAH
9jv5NPhdCL2qBthBRg+za0s7Suw6s4KknNZjc+NBi96rirNava1gCWcyBwN2BY47
k02kRkOD1SbOh99zqCIYZ3KbpiZqCv1VrQgWXfn2OMUyjXMGi5TpkzctuaOEcuFQ
r6lWc+P2aS6rbGrXzDjz30AYwCNNI+vRgLrMaB16C1j6f6rOgtBtygsJzmTjQTHy
UULIsRN9pd6ZN+/7HZHWh8ZJ4claUyl5OwWo4ih5uV9Ur3+syMtzdEzk7HN+BLHX
CrUqHPCd2X1K5InLTLFHnhrooaoeY34Q9aws3bZnqaZ77GacSjQLBd/MmrQpOYSv
ZqCXvQcQ+cadWnL5m5i2lqfJYGdFtweCwgmk5PDkcWvKeDUgWUGL0mlslNaSaDLm
yNr9j2coTmtGFmXy/PPdActMzAw4INed53GK8G4OFe+HOELzi7dWNLLDRTQmIvlS
f+iFI4L1zmPoTYhc9yqEU35PnSJo4AfYKDg+/usKVVQ3Sbo1e1c+j7MEcna5k6/e
thy07ZrZdPlY563N5Zq3MEcDDUM6FbMXxpnZl3iwpNCzpnnBgi9h51Wj5uqLTd4T
Nb0Hws/KfOtCjMe5J19VdCe8V0GrsrcWtjhyLdgSAjGCwzROlH4LbQ8foMGBoDF1
uU4Mz9FjHcjPjH4SJw6uenPFOEOsi84k9XPQP0HtjuzhMpadTMGI2bj7mPLD7/4o
3296ZXUHXgeU5A1lKVV9lLREne4Ydrih+E2YpY1+xNoIgsp7aSAeZIaathTUd+Pe
+8ODZqw7AWfOsIZHR4RcQXX6iibCw9ojYWD9XL12P9O6Bgdz5iVjMfQHzs9X1FFi
pS9+p4s3LYmCgesGA3e26Z5yx/Wv/TL27C3JOiVPysKdbtLmLKeHEZb0Y85P0PHX
JhPmP/WK92HD0e+zSO5SJXPWLtQnJ3K+jufi/w3h1qI3loU8KeOgJVd5lRfsKW7D
pKZvHvGew+v3YNQoCACLihaKpktx6GSiEVg/VkOrKA0r0Rl4j51mAihDUrj7tiSM
Ov1Knhj7Eh6iFr+hFl+sQHvKZbRXKc5IuYsyxNh7lH0WRCn7SUSQLlGXsbQvZofG
Ja2z8VGZFAmX44PUMo0lK/bd322UZ98BDybPZu7vKwfCIQxf0GffGU7mlQbSRxeg
LcYFviFxtEoGxNvVtoqbaajaLxAPizSxWX6dSce/mtDUSnIkphH7okEz1Q0OUakr
tHUwcc7v/u5Trj0OuWfIvsNEDMEsK5RAajqRbwciXjFfR1QixgjSLB6fUuJpZQ3J
lpQlOPpvmAVh6UsHIrLrahG2HQSW5wIvfIj25yDRBUgAjD82GzOjZmUNPQwg4GIf
mMdG3DVJp0umUA3Mgif08L7D8NYeZiEf9Gh+FQX54hsp3r/MsW/+FyTOis+AL8oO
6Ds56EpQYNvgu3LAV7Z/4+s89qzF0JGWRXfEq9WxVHpgoPDp/KH3+LaO8uqxT8jV
YvcY9E78xGTHEiYHRgixvzRtkFUKAE7PuVHdOewDGwJeQO9csCjLZfAX1yKGTZNW
3GIZSA9wOBBW2ExjjxDwHibv8fB2xPU9ZyGJJlA/Hyzt+fuCaaVcY1morQ/nB12z
GPbjsgjsowcWQl3tClDQDz0iXz5solrU+bbnFlh+JkFYbJipA2JnhVE6+t9dLjxu
QaNq7ohxBftorF8OSrnA4juSkN61F1JfEBoaiu+brHSGD8wdWjUdSb3xNEM/Sdew
I0I5/D3HFNrwnOkPdh6fXPYvHrMlMiPH0N79OSq2oWkEVPAOH73IQhdGHlGtzQ1I
AtoASRvlFri8eP7zp5vhjtGmNabeY0Xgcfoday+UmsZ2Rp3Qi/1z7bjXOzs+VG40
aqaE4l9pvXEMaV+QTsU/GgTKPVlIHP1sroXRUk53klmbW9Dh0ow5FjJbh/W8hKVE
zBt8x2qzTfouvqy5VyhBl2OMXJGoHrnPpQQRCBsIx1iEwsiQf9ttD/hbUVs18LJG
gYO/jAzCpxNEa69zvloaedMGRmQZsooI27rmqZ5qeLKztHl3Sl31TCfIJlg+KoYe
oA2VZldIGd8KLQcQ8kbp/mqC1ywYEHm3WCF34I2t5msYkNX7/hrZhgwWGHu9TpgB
aTouu2A7FrgU8/U3HXXKi6daMeN5vm+WJQDsLjEdkBchbno3NwvSE+4yfREiveXU
KGOQHnlSNfJjHO/DAmSJIbdLS7P2o0q0e+hVz8U8l+dWuH0kWOp3Q0M04hLO9EkW
N9g1THIgLl4jh1/Pq70tdIgA1x91KXrLTAcCFh0h5wdBJY3QeGtSgZ9Ul2u+rR4C
aNujizNeKMHsDeHSpKEfwcEnLci87Q4TFHEseavHWE5oqUu+Bl6IJf0TkZ1qemei
ENuFq1PM/Mkyvl4wwh/bEOkFPX4NHRzS8KLPgYJ0TRLHK2zKSZgJL7Q+Aghg5vSX
u1Xs0ZgM3KoCw7MJq3lwvEBHAd85X+LLef+B6IA3FWd1IxPu192wU5k3s5UFOjCG
X2l3zcw9aslog8wecjzi6WhLs2zVYr8P0Yq2qNP1EGu7wpn5jfk5RnX3fl81wfXp
XNRjysB6GSFC1BrGNVbcXIc6zyaNk/Gv+ildbccFzwYr+KoDle0DoSxcys4PklzK
yYNtFrzP9Ts+k5D27cok4LFFZuQM3IpGYFFxPDiF1ZBB/IJ8NSGlINtmuu863g6R
/1pVZj74m1LhHlLY3qY+bwvkV3sHBCoosfdvUalh04KcJ9WKIC9MFlUKle1qmdRg
6KdyQxtHnPMgA8D4xB9JFmXMBAu2c0YvOT2z2ldJbh3S8noMmqTAAULnzUZV+6Hy
jC0YmaPJrimE46lXZK2AdVCpeUm3/Rzy47RlONpEu/Imv4tOAorb667t6xwHloC1
hzdaJEzAHpKhlenj1HUz21RT5tDntyFGbk6Noun+SWmEYH0GLsv+/kHi4OgdyA3f
TUY9S82pUEVY+rxVqLOfVMSUpyyn0cNbAeMn8a6DZkdpCieFZfCU8GJFFVDzd2VM
R4NYzJuvzMHqP9/p586yt6KtYjPEwl2YZtEX0uyo2XNOuWCBM4bXAd7X2vkeEnYj
Wpppwjf7NwDtfTzdOAf1pV/W8JiVSTOGS5y0Lmk3ttfVAT/v3vjoHBUd4BCvOkbW
zAgBQ+ArX1bOdgQDiAAyWLixr2N+iBxa6hUAc+7KVQAc0HxZMjx5sOO3qjyFaru1
ZXotUKIZmtwuLgt4FatgnfveBq9due4Mp/EuLIVEeSXVSlGj8ZSI+dKp18TG2Vs8
JNb/Hrjy7C2pnVX8Fc2OuAxvq52NTfC0ckvPQyNdz+52M1VSgByuF+kr1hxMLDjD
+Ote/hjyJ1j78FYSYH/Dbu16Jtz9GCBZuFD/k3szpfvwnQyzkqmwJu9UeivNY96y
I+d/pAzjJPGlHunJhfq4DUGGrDzse27XaRz070xZwrlEfnqkQh1fmdyBHwMZE3j2
qPLvrphCtCHk/TvkvYxLPFePLcrtWAzp6IFPLByVA7uC5S5H9CafinJRUI+kMQWF
au30oel/8zWLi6K82z/jH+muroBClX88swaFN5a9QCpYgXo1VMhuQDyQKRbDnaGy
303WunZw+biRbZjNnifpFf/3Q4GyLxJxqQ/1FQ4jLDbtM9CKTdD4bw7T1yL4BTWc
040jgH1Xmk8QpI++25kr1/Vfclp/USZebIcL+ZWvJJpB6dstuqcWrWVaq2zNG7RK
ax+5YUFzsFaOQIIcNaYxCG1AJIAxKtBCRNVudaMePil4qGrGVMs32IGh197NLdsv
oB28hsQCLKcQElyJi5g3HyAPLUW0hhPWoo2WyvydEXq+lyFOn3NHBjCdj7+fhGZh
NUI5hpPNPObUjOJskT/ujAS7IGs7wXvk4wQSxco6WoSS6nRQzMo1wEbuw37KGBdF
I3Hrhuzo4JYV+ub8mya7qOUZxjvoJy7PdLpAM21O3g5n4iMUfnfU7G5p/IIrTR78
Fe24teIyGVUKAdq2qHPudXCJIdqYgAmOJ0bt8fiE9BFsd2pAu9xGO7y5WHJbOpkb
kw4fztu78NdDZznUK3wQEsyR06boW5GE3u8uzSGfkU5yniWuOBJucE7stiePoBYY
Xed/eyjjt5du7IFmKh4Y1TUALBXEBid9/eUYtuY0uh//ToN1knzK6eqq/QecXzcG
wweAnq7DTJToir4rVO30VigNzeIsujTI7mQc9T8zLGp9BcCVG4cxLxB2L8Z5K4W2
EzLYV8pyDwrmVC5oReaWNqOwCKuknmjG58wCqU96dVSEmEXZQhiGFByIbLEI6Km2
x1dGjZL5zFDkZleUfVjganTuT5RamwoQBWXeJkV30HGdFbOa+yRgWIsCzHS0Sjqy
ae9fe5AIiQDqcGnHfaYtJwU6+L4gwPbLwkfrsXOVQ6TXleSRvUXsqc5EJDnTjCmu
x8oyzHoh3luSRKQYS8gcicVCSsmYan/RNOhDmlmqgds4BBqEDYFKyh0Z1qr1rhRb
ALqLr7lKiq72QHG6Z8eoZkVZgMB8smcwWQyZX/3S+BHk6DI2jM2XgPGw6kZ+NB9d
WodaVtaOA1qnVq3mKPTIVHuJG3KrZArmUon5aXEQprSdgEzoRt8IB+NCVNVHJtQZ
Da2fPXjrjRNGvfEkv/ME0NBy8O3x5Col4fMK49SCPa7L1x9tWgpxyqb5h2xq3eMF
fCUM9bDCipA86CZekOBl8u25ybh8iDQIF/R+uQQM/gAY5p0t7pGFl6TB7HhwUh6x
zVYwNukxpoc0E7a8eUfo4DODMogu5KV4llSBTfhnLMtYuaUXUGNdAOt1EMuCBjzo
c43u2p/07IbMlqohweFPjpiaba+vJYJAYWkXlGT5D8eFfmshPshVzJM3JwG8OoZf
sLKYmxI1uGqILlhNzPJWK2SLo+GzPBO2x134sYJ1R9LeOMSN9IZJDelpddt46jVt
PRYGbhnbEWF5tnpgdM2Yy47Mp1M6u0kKJnD694C6vub9H0dqB2JQzZkD6zDZYlPo
nuGuYtYiUrtIvnFe+ZYmfGUHylbNwFKFWFcm5jj/xk75mxbKhUZu+ScK5d8HF4Ae
qrGXSUkrjfSVmT36jbiyk2KehjKCqxjaqdlTM0Y2WpLkIBCZZrtv478qlMd5vbxs
lsPRycq0Flk8+2i9b9mokSpkXH0RUfe6Nt3qGgv/IGE5c1P8ELvJx27AfounOGS1
pM6Mb9JPEsWsnemt48e+Od8Np2CWnFBl/jHMm4QdP0h40KQXbMwXH3cobbp2cHfJ
5LhvzfOXOTCV2SxjpcMkkosbe0RZNrI6AoKH/m0YM5uNb8ut5eCKGzW79sKjI9m+
F/ZOsUlrJ2tLj8RCF2GP6UPNMwrxJs/EDqTe3L/ih1ePo+lxBPZNKG/SmN11UOm5
FrMYfZZO5Om2lflSeYb/PDV0ojamQ7w0L3crFgV/Qgr8YBPreEF4GmI6PaczgMXV
8oF0g5Mqwr6w+OaLASWYvZ7snJNPA1JbofeghITwzr1VPz8pJOBzGWDVTBxfA06r
3up0hvqypOKR2C7/rbv0JTMRqpR21yDweeZTXKe5KlraFYG2Cx2au2BBMx6uu4Hv
hS4QCDiB9w7r49/UWpu5FoXYiaJNkkopm7UTLxQTUmify7hbf/yDJrpwTwc85GrW
hlTzKrDugLy9W6JYLKsnb4DaxNL0Om0T/VmWOeg/zIcbnaL/CO4bq0IdPUw+Xw2Y
sdkt5fegL3/QdUE6VcEmfJ8hJHl4hlVM5YGuwU3ws6IdeQEr3heoDasuhz5mO8jG
dZjHvudS/6F5wcJ1TGnA44XpsY/m8sO6lBaIDAfjrlmieQXGjjujhO5KZeM60FjP
P6Z3glSXVaQEmbYPGZZnS9cY5At3bbSje7MsthwucxqDCaQ8IS5qN0KdU5ksMwIT
eppcG4hVil1RBxoh4T9GjPCP8i9ryEa7D5kgqqNkSayGaxs2pFRaopkEnDjt60IT
CaMcp6e1OUfyiUEKVfA6/2yg8ZefpMPtviNQbI9351T3da6VHsI+h1WWUSSpYmfq
koRm2OK9UAAq8hcpWslrLgbSi0CDtbCZCP2YiHS1pmLuJTI5i9AngQbNf0/gyxni
dShtN5MHVlgqp80pFzn9WTNk2YWzJ9L7+Xr03m1vpDDhNRuKbgiqYB7Qv+dHwiTU
Pjhylwmh9QAKQF9+WxAz8E121EuqGr03ssKSWoZWA2LXe1es97SenMQRM8J9IjvZ
qoDkjBl/VM6UaQPPVlgOs0kxkgH/2FeYOkmboixMPK+nnNsYe7Ej5QuEJniiK5FS
41N/w0gGYZmeFolmGlqse4puUmwmBzUFF0C8bWsNtGIpaAUYSBI46nnI0Khz482G
3riM2aLjMCYsWglIYxlftCtmjMGcP8XG591P0LgfKUNvnjrSg9V7+AHOca3o+nnW
U+D9OoZ1XUl8ZNLIv6UFktmpiQ+0M4lk8el6caBTZH2Ep0jSJyFI3fgquG2fHf0x
Gtgc2FXGgXmhaQ+SyNeskpShjBibF77ZZMeYgofSOR2qTirdp9IY1f+cqtEFbhrJ
QyPmq+sOBdILw1+YIYvbVbFC9Kkg6JwK8OvQL32v3pvqxG2t37cgj7pVWNwrwkdg
mxXlGT3K3xLWQgZLD2O8zVj8MrP4Nmsv4IPNx/xcT8UCHp7+xXvnl3VuFVKIlL2N
vKdmaf5UkeUjJbttm1dUNeD4kiDpYwJq4m/tXyMNoO5SaNJ5uWaq/i0/NUZ3tvG5
olQ9+8ntgVyhvLumdFEyicJvp8YCPkXUmkk24OluAgPwQTGjrrjz1cm+CsAuJiEl
QDpjAXv09kAf2p5xZ2TtvzGt9M4oX6L8gHV+QETKXe5s99/fiRWZOq/xB+wjM0/H
fQnEkFMxrCAhtUkp0b7hWTTSmIgaOERo9buydDeA37j1AUPQHkPB+VeIoH2tOKp+
KflQEm2Tychlh0uzSIEL47D8EEqWonOnbHXHtRTrEhC24QSTTljTCpbUnfaPyGPc
UgGLOrNwrGYkl8ayfffqYmIeQnYYI99IVYiBLpHnyIl1krG8ZyBaZoiHJrq3CQhz
eOLzFPJmbvKfKLrh+/TuFbIrJTwGC7/nI563gnELPW3We5euq5MEFbQEuKsiKkLZ
x9pOp91feD7QgMVRtL+vOFkDJhx5fx5sMnRXLZqtM7legsoBMNp6fpnz3g4wpTLJ
Lh1cJT65FnNPpkJxVqLbb8Hda6nPaG7tOGXcGx77t7UGO/6xyKrpvCfVVKHIgsrz
aKvECzsLrKpxWsBJbUfsWjmp8zLWUncnnZmS6BSh0Io6j+tDI0/Gr5aj8XX+URtZ
1Nkl5jyUMfmtNmYpoDTel+WiFc54J7KAy8kla/PiPRu9CKbobBBS1mj6MdXc3EOL
W+nby6H6lVf8y7DTrY6jTlF5Efmi0pIPh02yprESXWGKXeQu7jIKJKiDIc9ipqIX
/5Z3QAfWEehwbP6KpMVvdO4UsiVT9csv26e2qHtdGRy4lIbssR0CHmkfaXNE6sVR
9Uc8CdID8t4EI1hWkjQNh+4gpA2k5CP6UwIPY2VY2i2GvRO8ykyazSyXx5Wv7F45
mdCaKqoPkWmXi94mfVorLD0kORX80qshuLc42LsFlEOH/RliI0lLf7+kElWTZxxm
3DTBhP1GyiaEt7CYLMWXovxnSJT/hqunRGH1SC5CfaAtrZuCQaNWTVDE3aMiARTw
M7xaP2Oexe1IYWeaR7coB9HRsmGHoBWmqSsRONCGlIp5xVK/PznfkhmPBwh3/Y1o
GsQvnZvaw+w0M0TtoPfRVjfjk9ySGd3lLksue5gdqcu964COG7tvB5l+vJsnIl5y
WalmEqoPrZeFnyk4VGRHNtTH7n/+pWxuCtPNcubx1oPXnGzzoekkch5Tdkc37F7/
ACJQ3Poon/FoB8xstN1FUe1huSOfi9Rf044goQY4K31yEAHj8w3+gRI7BDAPVGiQ
6fVGuVLETSm2yXuiFunCxSnNypGZQQU+k/Sn4/8R9zkjSrHvJCc0cGXBurQjisM4
SrWb/UYaCIIKW9GDGUhIcjOrsQcftaj33Z3buPEJeJzH89L+Ha4ZjwBTbQvEcAql
38TDUnxU2NChIfvOICRsw/uiTqXeE+y5JkMUOLmccqpznJUQW4jyvzcVDyYsWHad
bymQzDBgo4uk/HRm1zpfGvc4b2ktQZqZrX888ZxRQ6QJ7zVjVjPJNMnxtf23k0Qe
+W5UAMFO3OtNsEzzE0HtFz4c0BeHHLxa5lYGhdx0ByuOkk5lsvorEG0eTVvzb1uH
5qR0GiDyk4J0GlkFL4kcBW59jcSpk3Zl/KQvi8lDVl1RxGzOSHIndASUaGpMgND2
m0a8rG1TMey4h5BGEiAxDBjqqTDI1/CEyu+JcnK85YmtnizCT3bIE+92uO36GGtY
pn35PfSkZcfKw51vkd6WnrmrYuKlixzeiLTos2UGt7LKICr5tlDZGEd/LO3ovCCX
KEH6+asQIWVWCWw0LZtGTgaV+Q0Jm63swUgW8Sste13ygOc/K+yXKtZbFugDc4cW
lEc1a0sbj+L5zHYu/vUNMb2iCVezFnrlwJn0ZIyM3ZXh+aHJZiBrD5niHvEvEtNO
TBjasyEKvSAACO18pbFPMpr9z5WZ3mGt2csVyB+svxdC3+dXsJD3TdAl/8ErbQtj
oHTZK+FnwE75yJJqpkxbRWsaVebktznWf2wC2NNNAp7C8I2NDv0wVEJXtFAYVgIa
yBUlIW1QomJSsjizxkzlrjVVsyg/Rvk84N9cBmPKDB4+Ge/rdywnsC+M4a6EWYmf
1t+isFHkRGDhwPPZNpdfkRB/KWIzmYXxjgwcbU9rXfz+EBuGIgbstT1k5sYrCZcY
/bPeej2pGsixUhtBkWsdJRH3TSuzTw0t16n1Ke3LYDkVqJdcjhF/SAgcZPNRvyT8
O3e8wyqRvZdLP7Fc5PJSOvR7IXh02QXuMcWUWefyGP2fVPKGMzepZnwj4dc55LRs
eHnE9hGvVleKw0ZlWXRRMelJiY6wrJwhr0OZiEO61PgGweZgMj/rmtdAFAGlmKuO
lvuKhWV5MS6LYu0fbbxkXCE94k/ASYY58/a80e8TtduAFSaAVxKfwYdPt/Tq/YOC
xXI3R9SNpXZQdMqHmDf3nWJdxLmfx8JiOr+8rW8EP7wIe2y7nT9dXY2O61vQ1Not
XBROyusSf4szQxUlXVbHFw7Q7M/5HS/v0CgWP6Ll2eFI7wdlRaFXPFDFi6NdOH8S
7x4gUzdCH0W2sRhuvVM7Nd7h7P+xoi5IjP2IXTBjwqreH05De+K6Dp0XcdjGrX3L
Bu0t4/TLA1J//opr+E6Lt8wZOn1oMbJZH9ZNz+k31lXdgLj+aY+o/tUsvaTKCrUc
KE1pe+BtQLA1uT0n7YvKQYy9xo3mwkiszUhC9TPjsc6udmv3tqZSZmWLVZsfjM8j
Hfoy98ovJTQWq4jtmpkXc9d6e2kKEjz7IgAojBz16dtOXSshPZ5HMTli5ltU/SL+
GTunoFKXjr3H4ZMe48q3H6aHg92qz0g2B+wJPBa9zRR9hLSujUtYFmZgBDhpG1dF
jPeSAU5OHBrt8phRLZvTAMU61WR6Ii1vfSsiCCXpVAEH67ETVENQo6Y6uG88hn/J
ynJ38rwxflvC3W+d9s+a8ihIc0cKSAumok0GUwRQtfZSRzhpS/1OJMpEWFMvOp26
L3nP559knjBcmRneZp4crQkzNKDGYzUzcSaTXExxSVa1NrMgwqg0K23eyh5gNvKm
8O+U+mch+yjxGY7xrvG+ey5EW3LUIW69BkEbNhrAIP58yRbwVIQNZf2Qdw3Wx37+
/J+Zpisb/U+pXQObWGq5Hc9mqq2ubtJBLPYrFm6mVpfIsdzpjL66hjNFJ4ZR/DHm
HSvuZCOzEQr0/GvZDtzw2iYVa1gSZF5Nvdzaqcy+A1TXavxDynHSdKzGEvcqV9Cf
1qBakKlpZqzLIdI5Hf9ZxIUnYc3j7ZKz9By3HtrxnETOnlAOJFF+I5E2vvv7H/h0
BR6NNLXe85XMk9Z6fyaQWM/slwAzNjUnHt1E428XuMgCaqEtrwifF9V04W3DbH25
Jxecw0LO9KsdQPshTIY9ouftARTk9s/6LQ/1UCz5LkQF3MnPbjdA7D8VgC/d1lYf
/WQRKeSe2iJmqGoAek/SLzVI/9Bw59GNf3iRKvi/CHN+AH6NmN5eigDocChoHKuH
u98JkkIYq3CFzbIlC0bfVJwYFGuAmBGWQqkHz7jL3Z1Rsq1pID5hLEFVV6ISuicn
XV9ghjwd2kmTD+Uq6Vo4XCcsYV7bnN4+94sEj5zZBbrnHxns/EbOT0Ho7/EPR4uD
hIZ5W+PzBz/KH+tqK/vVczG329sSiIETB5lB10RA4r+/Jtm3aNqFC7wLo60ZSS3e
Epx+pU0bNURb3qJBtLKS7C+rs81jsI9iFNFqfuI4BX/L03nxQ9d/PlYptWYO/R1W
KihLFF6oeo7F6Y+O881yw5O9CXGh2iV2qCX3OaHS27SRp08pRtuIYjujrwTo/Dqq
NKz/Zdqr9EJP952Za4zB+q85chwgApGbQkcbjZtXMYOOS2XhM8JbfEyqvIIT+vyQ
Su56HcGnUF4yR1XYz5uUM9wH01ci6pAMGQ+aVH21J8I5Nkbk1I0L6OYSTHpWqnI7
txp2EG73KkFuXXcCqifTSpB8lV+386dstaOpn8NjUNoGJpWKKYfz4CiL2xYxLJnX
qlv1KCYp2wJGlIpUIvsPn2uLw2pP2+81dx2cXgSsnm9aXtp3wJMxTIN2Kyr8R3oS
GLE4/Ng2e07OWB74uxPFWYlhC1JZAytdqDtjPMh+SKl5X8G8mPTtN+J9hTVJDJ3J
y8a0vX/QwCfETtf+B0B0VEw97mN9ZRRxlyo/ti2+nBfGOlG2XYN4BGgJHrc1OS1I
chgFeyuFYBh1X/X4AFYlcAzKEEReixvbXdP8fyQg4CreZ0ZBvJeaZQlmNbAXOsP2
KOJqJ/ThK+lorTUYpyLArFyj4iJLF3FB2oBG6RDuz2fF323SoEXwehaW4D5auS4N
VvjmLjLpu+LJ8bymJAx5LGZ4QjEVRkJRappNSdj/u+3BY2tt5ALoxim49Mo4Bw5Z
WNGFYpjnwEUU7qQsoCJ9n9gC9oR7m8dcr5p/YRCaDt9ykFyewO3HLpOe0b3+QyxZ
rF3iBn8pGMUjHj68xFRHw5evWBM0pXJMBBvFytlyzpsy4KYByRu9JZlnXxn9nclJ
KRRGGJChosnOkUC3XItluFLL8Pwq6hx/aeoOO8PryMP2wExAS7qIksvfrs7wNtIm
Gle/d5ID6Nfi9lDaOVvxvhMsPHUlPNTWZFY26Am+UKl30V9ikS2VUCYoYVRH1Sdu
nGagHPi1nu94F05Jzp7eAlp1xbRxqcit8GTLYbUsJ1HEXHFPsJX9QqQ/Vj0n79RT
iu1dOY1W2rnvDAt/TCGdkk57XgIgeVyomoCmKhc35sC6G8kGYobuhedNPdzj+H5l
NXFpM+MUDEDhjh+ctvi43EC9DNHeY+8+vzOl4TeR7bEV8/GiKNwVUNHteDKjA3Jt
WgYPWg7UqsVKfKXrzUrZnXVRo40oxR6bBHtVVG5nrg1qGs1O8JYEFP/khnowAjg2
rJmPtnGFACMSxjJZ/XAj39ha5S2YHBjTMbvWuQiHe//G6LN4FgsCu7+yZ7s1qdEd
Gz+45DEZZDJQEwc/tD4yYNHA10GrCeTNSOEvVcox+zqVGNHNVAWXaqt36sJve6Xr
hKwWyB1fhnd3hwXmVjsDRVSRjXPbj7zSD148YhkU0UItFtTsDi9R4rHSof6zez7c
pnOC2Ep9NnyiklLPdtyjniUWHc5PI2BgcAomnSEkNnkQ8tEuHyzC9MrC/J10Jyz5
H4TimBuFjju1RwFzrR+5bcB54AvVKb1RWCpPTsfLnHzR26/eD9GM+xb/VP4pk8Pb
B4CRlIvVoGKaTLJjTw5efZmf8gtYqs2G9aI1HT3iaw6uRYNfs46Xb3LP5ZAJT3Ag
JOI44I1iaBr31E4/F4iy2Q4Ad3bz9PbpnaWIL3beviSrmmX3BQWmv+WjyGWB8ih2
VDRcWnFnFixgcrhVcCQJAyLqLDvbTEJOTJVCZ1pKMsNU/A2PCSgWcBqsf10bUg85
2sAhZRYC/FpNd5tQEPzP5rvwn+7/8qkr5TL7NvMCwl8++5yNxTjGnFygxMAFeyK7
gxVLtff/rBEzgygj4U5lI8kzUXQ4LoVP0juivaU6bMSYxAZ1JP7q+7wBxYhjTa8w
7jg7QLbC5TEcYxztDdxT36L2yLhMNypa1EuIXMeD9ufYRMz0sFD/gZOxWLMuv1g5
W3pQV859d1UzeHHntVssfLFTkdT/zRuAz7w0bOXu1JNPWIYFYk/THJf6jvP2y1vN
sRu6OrZstOrO7DZ5ItNjFMZGNhriqy9xrNc8/J7alifukQ3Q+qSTT5YeUO/3hJgN
MSul+UFoc4EOB9cLssvVIl8co7K7qzu1FDVJKnOYQPPxE4o7H5fKNdaQJlaVW09C
AHlY5p3pi5UJ3VzN/vAwdUqJ/HBOP2TJ9KCOZvzxQsGZYBhO5zye//bjaCQKXSFx
yESbBtEbQ77MDvJ19TnZrY/unVyzOUFv21s7FPW3DeKGtJN9HSWaPKs/DTCc477o
AtH7Yi2yTW7HbQ85BcMyE7rU5BPjqjPAO3XRRTixCK1OUjkg7iKEPnNClN/ly/1c
78BeyPXValRHfAN9d10SStDKKKHPflrEfrYJZ+T5/vtS1wOX+ALUJ7oLoHYIxAJ2
ztF8e7dCBL0IX9FWH9A2WSBK+PT6vvDDD0lOi3CNiOzypANlKMhHtyiwKB2Ae68/
CPAJavZ2DTMn6H2JUTIhvMt1lhIjweD2NhNO2TVmaRd4vs/myuy3kjqcfy/GercQ
O/ZMRBdFKPbU8cn/HcdPggSwEww5MDWxAQK53Bxv6DknEMrHIqjoxqNNbU4AsBtN
TgxHTmBmMipALQcIu094RV26udb/JnL4boMarfsO+pG+A1+uXUi/dqy19/JooaQS
iSk+6btgmW2tOXm40wjenDu9vJQwWPAR++d2EqiFyWbDVWjtuHIM0FmzN0Co6c0E
8LLdAhyZVqMV3oKtePwh3T1c8SSSRDWCzwKDvQzYcQG49HviRomyRnc63reUvuYc
Mu+WK0bQu9ISp58ajvwOknXk3izXop0RVK+FqV1iItk4XcAFkAJ1dEFX3aarhtxl
w+1AZ0+zhPk2OO1nsg5fsmKpg/JxynaMK31YCXDXulP8pT0fj9KibUe4X/ykuuU1
JHLCSV/9cPdkj9w9/VMt8yXBB7R6qCntScrpuFlhfO0BFX0zOmTBMVq4Z22qBfZ6
nLsGg0fx0rOR7nkBxdlpDDy+WZId/5OCW8rHYXs1IQmUfMXNlL817UotIkV1gNsd
ZU50Y/bv9GAr2AR/bqIvKS1poPifSS9nz/PbwwgOEioejswFvHh4Rh6cKYpBmT2d
ekEX2zAjXowgIvyGg7fWKpF/N0C9u5ykTy7Y7i+I6migO9h5g3b72LKN3oxSLlLC
O+WuDRTyB9ty9G09sZ0aKxph3PwzV6aCbPlFibOI52UbyoVE0g8Tz4jiReULk/qO
3yc9mLm/wxO7LcWHl0E1gTkHPaegqkNthVnVb+HShvnkFjJq98nhZZjkwhUVB47s
xqNSSC3kB6+lsB+uVs2UuJczqHdkcCLnRHTJoVXg1c/wttsY8etVtwycyLSqyJE+
hjK0iHd3j8JbZBiIL/UGVwhISbK0SjufiY23mBaNWIpA6g4JwevhFxmp2XDwvhXr
WxTMROQBAwXDfmENO5oDkiMe6qMa0dpcHbG6HTz82veUIvaPWUXMsGK9yL000Hs8
br9p0km1RpdswD/Qy4nb7xpNOKvIATTS4wIZIbFHZnnVYqQcTthDNIt0orj4f24d
SR18kJBSfMZv4FO8sCzJoQoiqhpNLuYUA7sNB+kt0OYS6FRjyVIUkxXeAJ/wKM87
X9x7pU41ZBqm+1MoqLW8+KqW8/3zvUXa5Ec98EZKXnEvZAO6gLDfZuDNNhGSSYgT
B9qx84rM9F9R0dEigY4bsKywrNjJCvzYWj0lrU8FYbCZQqvLFyaiUU8MOFrPkXKH
RzGEhiLYUWMBrkZX0R6nHdX+ooAXs09BIxT4f5ZPVjMmdxTea//Sn+8lQ5unEo+6
w5L+Q8YOixOLFua8u8nkvqfp+ZwJv9WpU5w0wrGlHQLojKTng9gZpIanV0cfQOoZ
c+ktB1ZB7SEH/YMPh1V73BQ0uz8AiBxNsFrC+wBpy/fDfHeyeq2pnlVRWaBPBOIw
6mQeVE2v6M05USgPZll8Nd5E6jgDJZitFpPgM453Ia28x8d5ATCWHEfZsPLlNPeA
XK3CbS8UJI1DYJcGpwqJ0nW6mEytVDvxIkTa1VFqO7mNA22dvyqdQItmoCIq4pXn
lRpFMn1rK/uMJqiqI3YkZQwc9X3D+MP8h44N6ElNffWqsodnZj56FTvd9nu4Oz6G
I1llSmaipyXtGGUtReeXwABNpCl4ZNmJQByJG/PIqd+g5rl9BuMo29FVJeDx6tSk
7WTBYjAoE1A1NVpXZTD8eHkRqHmKO+P0ay9f70HWF8wv+gQIWmJ0Zn/cbXLfb7Kc
7sGFMf/c6k6C4U4i/g8AQYv2uDGB4RPHP4azwWXWgeHKqhcCyIuQZR2vcwzBeDgz
eRE4D6Y+yOQHXi9ujjz+Ku7wb1SSKZwtHN1oIDlysbP2Dhq/JsjtWSajU/fDho4g
BZu0UIx+o/Znokx/VL6PwsDZSkrW9penwyMuia3tT4ABJdJS/kuhnOPZXzKc6Ean
iHU0PfRlqYFbPx6CYpFjYij4QLI7cc7mTuGb3FoBG5EPvEV0kf4W+y2h+cDoItpm
79dDoYJt9gmAuDP7wSGz7N1fiE6s/vgEcqTG/AYUxU5TdLXNY3wUwnktU87u7ly6
yt332w/4iGnJaeaQVuHJNdrQxoo3B6XZAyWNKPeA8953UOCyLPrUFMATPSwFlA77
d8zl/d6XUKWIlOiW1ZMaxB/5bXK8/u2lvbvMeZdBwKlo4REhOdB63bD7b294Lf3V
aLUEAAPiMeLltlaumvtusxAdASKdyuF5hRerQV1IkVpGh9he5gKvJi2rLNNfYTWD
VqWVImP87C/DUlnHDpzbQA8QokjGEXjVe4TGA0uCre1pYz9WNe6ydyh0stU7vf+r
h1rSs8Q9HCso6OZ1myTOtT3bic8y+jt/dQhyH0TH/rw6L5DqZHaovyr4pDMk5ad+
i9u5zg4vFADYi+/cAgqjHkHzzaUQp4J+K6zUk5QqKO/ygN8vJoU1D85EH9FUdTRL
n4ifatXkuu8FfToBFLfwD5MUJn1m5sDzdMXGNvjzHyUsjBxv8kIE8eMoN4Sjk6XU
x0i/CEvp5D5WUAMff6YVc5PK0WJ+XyEaXfJmwGWqIjMKhf3b1AWG7DQvH30Y244P
dKgRY4cOTTw3TnLSx/clwiznwvlfzR7r+4jIMVA0MlGWNltO+aRxAQ4UpZ7CL5EQ
SdrHIOmBun/wGS7SJ+xNWJbHbVRx9m9Hjh13Kxb1V1rnTtGptXaavsLuevb3tSpz
kZthGaS7PKDi3LlCp9nZfkPe07QBLmwYQrIEO+iQ6EzzwayXSbVErX3Sq4maU6fy
X5OjivdPRYVwzb9lt7BRWukIlnLwfAG6xFVMXzq55sitSfsHCn6t9vhXkb4o83+R
L9s9WHE+DGvvYS/Glw52z4rxiQqCB7bVnnCpSUs7wsTzhFrCu63Jq2I5UZhHHsSz
6NHtDOt8y/fkqco5e46ECfLR6lVqB10roZV8GzOKUfgMb68sYbQbB9Wb+Ifl96jk
N9LaU7VVOAYrIWSwoV81X7oeyv7rXHbhmcMLhPMp3jCRWlVkkyzGz3DNtVWX2TPm
8E0zdQdGreGpo7OiuEMEy5ordJSNUTNvirlrqW+OnX2SPkOR41rbrn4dft+17JOW
YeNCab08ccYq3p8aRKJ+LsWv4B8YXZf07B6X113G21Jtn3dku80gqmWm8TClhJ1i
J17EvKQNgxBoJnn7w8eELQ9wnWFuL2dGcdeS1UmL0ud52BBf2ZsxUPPrrXSH+wis
X9N3h3nNgT/96jthBvSBfunDUOhJvEcByrs0LxWhlwX8WLjc+3GhbkvRqCe1QGkt
96BxX56panah2CgzNQdDyAiC6HO65i4cNeXd4dm+MSLEnjGtEBLcYN5TqyfCVuxB
0+9WNKc5yclh6ZcyD8nZGqQMUJfm/6qPM6y+JFZ6hMQ8y5ptr3wNpvL9XDuai5t5
+4gDWBfT97Ek01tfNx/Td2nxjCvm+RMGL9qFoctJHXT65Oj58qiYF3MNJpbdPnyP
l+qwjqo1LdS09EAv/ng8Sey6hp2LSExpUECd81gpAnpu6jzf+Dt6QKk/iDTsAFOw
ZRVA3++WiDxk3jGdHxP/5FIHiBiVa0bWXycBHgq9Lz97cxvfHNGp9pyDmoFfycf5
oK/HH5EtA3JOV1/afAPcCDGqCYa+fgvPM4pr9rCDBLKuUx8CK2b5FJ823RIuO7DV
Ym8GjjBNR9vsxoStQW02RVuAM/pshY8jJsFFowohDmZ5wEqzm+WCs4kagvv3MVBJ
kuFHkoQjmAcZj28eiWXJRZxnUJYqxa6xCpiSE1CtBLBG3TsGUD0gmCCYGOx+KaW1
Lg/316IdT2peYehBRFfm1q5X49/cM0GxoodDLTCBD3SUA1xqADQ52yxkFYsFx5xh
8vNZooba0zrXREV2R15CB0sADOFXZJP3+VGhTtZYX2PrbASOk7T7tgEG66+K5psC
J8v3qRCDrm8walS3950VZ2hmyz0Mv5tbswHCuhULIzXrGUCaY7XQlDtbLvUuvzd2
KRnUNMhdhxrZbvXHR7wdX5jrnFscW8+XGOhjGasLHXIapt1rFIBzaccPxd0RYPxD
bbdMDfkV8Nl7CAgOCVL5IdsJxXDCcDdQ5f+sFrc053f8zzMTE3fiDaM8Gp8uaZfh
vmDabEYq69k5zWdA2aSj4jendVCQfB8hfVgMWijbb5vuGK+czdzjDTCyrfLi+dmJ
KYyF9ehcwn8Inz81oBs7aX9IBtTBnTMql3QDVj/zy1IlPurQTiMLUTuJ58HhUD0A
3aSbOirT1zq7+x4CshCd8+ixCsT61dMmvjDRAZFDfzwvnHaiX1sk15o6katCsgtX
46ppIr3aPBH2ElDQLOtH2SqxYHcdtRsZ+7CvJX1CjKN2CvPZiykhcRVfJsV2D0dm
NcZ82A89V/akG+bH8p581tvOB5QPNV7i7YD0bbaQDkYYkBUBGavemeChaVHJMguX
udKb/l3mDSHi/U3xlpLENZ2JIhOo5zVaZFVC0kO2oDKfC8/8q6CoTf2mCSo1+0TR
IdgGoYf4iMAU6ekr88BT4tQiJMvjZ8DOWRlU5/hDpTCpZ+9S0dJIgFtNIAsLkfE4
8OfbZKtVoZLDf6F6yqehlHPAsz1DpbtzmNBH1lklq3XtJRQ2/RMelxTmLv9rrd0H
KKGQ/pvqXPrZkAgzYr+adiHQzg2CYv1O5cg3EzYjJGxaZfyTHAQ9g2ufRI1Qijr3
E2ilERf/Ajr7VsPUkV4oDAKbpAxFPQE0Tgs6LJqEnWDbiGZdqnjUn20d1j3/Vnas
tzoLdQsNQ9TRzlxKbCeL+fxkTdhpYOmy+kIouD+FVR9Bsp4M92w0yzSM6UAvToD5
2VjSd2LtvN1bAF9kVUvLh8Hk79HM+WaXP87QFA0XPQP/2+1CTBhAi4sjSFkfmw2Z
bDw2pdlUMk/NHxDqiQHufHRetotrQxJXftqfMoslUmR4uf7JWL/v4jJyzc5LP/o6
FJcIH+CZCGLxU76eJKvVhOlcfBIDci2NnSiGAoOIvpqQfrTTl2GugeR2p1JXoCI7
5zwDH4cXgZnJrddYL1jKuE+wFsmYi3RXXvfSATCGr1UUbgAyQ+Ny0bdQ5AfcbE6Q
4vObfGFG5XQ80x5BvNKQMPeP70JIeMAYIBoCQuY/ECwLP/ONkVvT7jyeUMNqSZKc
QiY4Y528IZ7WIwvpKEA44B38f0/ge+as05rugy1lSO9AvVa8LOVf8U2oI7h2Hhth
T4inAPSAGoqpqoV5GEi8Uctcal4GVca0SRMMrlKsZ0aubU7HVbme0EnZMCyYljTV
Rc+jwxERdZsMGHfrCf+TLE1SVR24tZ/uJuHB8porGYcPC1oJWmPYaPOo8qC4SLZu
sgr4f6znf/w80jdE7hK0b/1NgwOX5N6LuVY9W/eQWRHYlXmYL1aCROsKFYzQ9sxN
WtgwaefvXPkHgXWDb5A2EWobygX/Gd/l5EZqrNCe78sRIIr3PBZqoGjLtjcug2/a
8Zk3vG/R8732w7xAImWtvnyKdxKgvXJeuc/xQUgjlK8P3ajpfNAbZSghprnfdXt3
AMWWYy/tsrAhKO6IwYlv1pHIFQ0WVIILhYLYLJ/fkpP4Q+akZh2Pkb/rGb1+Mh5V
wPUlcbxnrwWLkJJ6T3NAAIRWRczTm2/qQiEvKNgoUj80qxBHvOI/OTw/e+4oy/ac
2TLEZCyPfcV4XyTeYXa2buK8U5amcPcYEsJ+HHop8pie2n3FFH7l6E9obhAs2Ct9
M+cw6EniZIq6hE2rSzVL1jYN0F6HrUeO+NhBNtt9P0Lz1rDV6S7+KkZp9InSFkds
QzFZ7tLdTpHvP5b9iqC5xDw4BqOsqgawYaySNwYsN/pfw45o+KYSDnBgeaxgb3ua
Mo6d1ZxQcvKNnrsJaBbSFFIJ5eL+p96mwOsNw7xwhYOrxW7Yxm5KA1sRcEgmNYpN
OM436VOZSYuCFUlOD/9qRiCrrNG7rm/5uLXwTkMT4tEWmN/p+aKZFzHLyxwW1ttD
cYew1WjzVbFesuF/i+JC7VXgciV7mTDYmtruKO3etatMTBBVIpCykBPhOmndrdIK
tIHVGZ2SxZSmkkU/stpVEy6JoGHU8X1a97bQ75z6aVNg3c5E2ZnVFbH4/uAVuA0v
3R0oyOX07nf8oZ9IxbBSLP66mTcz7V9xf55uY3Wb306mFsjQarxEo2mxX4697n6a
Or+7/WgQU+N00JIc2JTkU7ic5dsO9RcrohjBHQow3PrfeVdF03f2zVyN3mGQVggV
DS6EOkwHVb1dQXMtjj+rcr1De/G/6vLPCrsoil+tHrwEKKhIDSBwgkzgAvzfV441
pRA4xMr46h26bGqZc2HZKYDk78qBfYDUYxDnr61HbX8OrD/PQdny+VQXtBxPuCrL
+0DkAmFdX173Qj4bHtTIUy4l5P4TD27MztGSGka9MlGd9up2QYC0mJ4hD+/2mobG
wDGr6vit2O5qt8mdBfK3E13sTbcVSgwkeCkl+fRQXP+lBjXOHZ0G52kO2V15jL1/
UEmfXGHCOqcSCjWJpdyTRSSacWH0Cf6Bh2z5ursjDcSYoHwpnzkCuoEWrMhr67qr
vTLKwQabyzvv+G7DG/JvG2XLdVopxziqCdJRdc/NYfO0y5TMW0VfG72LdW85QdkR
Jds60NY81J0RlI6MxuYCbXFa+3oU2/SWDPeDnUbgG31UXwL/DslaMN997fOd/or4
IUA6KzKxY/7rjxSCw6FcG71z6hQ1uSzaGXDYjd3yktEuufOUyMPmuBLX9DGeSu5Y
SQuuP4Pmoj89CcNlmqqKIpaezQVPLaviLZk6tQDtrEezfStuxUDdTZdtCssLyF/J
DhGc2Qp7aRflOlVlCfv7cfcK+NTGzQN5Mo+jSrmuWszx4qLF7ajqXar4jxjYwxRs
c0qpJJaaPEr3XklNkmFVTuxMmwqUQ1YKGqVsLVUnpgo2MvMBJRelS1tDkGylL+YO
i+iDiWD9wjSQfFbJ0fUcH31/65cLpUUh4g3c36BQnMT1YB7zgjYeneZoY8lIbFyA
IvdtbaRYF4+wZJn142Fy96b5CZDs4+4/mTvA5F7qe0U/ZT+TRMxT5VEFqeZp7gbI
1zuuyWWLqFLH8LPFjbW3vD7QOz6SE/nBGrTcM5xMeVlmDwHk+aYE/6aLs+7eFtNz
f1P1q0nqGliEvLI1MNg4U4H2cULml3OuY2vDc3bQDZ/JQNGBtVsTKI8DGO/mIjUF
+Hw0Uof88zOfqvk6ffaBc7jOFx6t/iisQ++25J7vJ7d83uqo/dcp2tw3iCAcI5rt
vwvgD+pgoNVQsa8lsqXMpYJS0OubeOpCVVY+zMjoTxcwV1xs6vx3xLx3u5sfjdpg
xzVKTa/5BMjZACPFu6mz3Dviwxjcdn1ywhMLUdQCP8mFutrQllN7CByJMkeGpO9/
kK45+DuNiB3RYpf5BlzgonLIMVLn2Uq6Y7d0XNrXMzvIeis5YjlAs00tbEnv5XsD
D/UAcM+gWOO/uMUw7arNuXIPwMd5+SnYTbLjg4sWwJAwVMi3DpQ4OQzc2hoso8Ry
tDN1qAEgjAcVRJVgKd1uDgzM17N8CFvoQYY186okFBXgMM5G/YtNKCt1eOvz/7f0
Qquv+Qo0ne6pzR3IDU8+4EKG5He1pvM4YFU1cNgorWTG7geJNCMyFqng6XjI1PkY
SEHcjW7x6M9CJvff6CRqQy8gCo1sGZ6/MsvQ7uRYUU5/UAbfV5YKgwThpY0+UVzE
Irty4g4VcM9gNSE6fvLnTW79CtGukRgGFkYj7hK9nn1sHZ2LtEFKLpnfylC0rOMa
xIY/3cXkacCTtyCgD/krbumFmCEY00YR+WU4ax2KgqEtz4Tgk+Tg7hIudKOby9TB
eL8O3B83rrshBBTDQpzGFeAPCLEqIlaqtRxUq9xJ2906eoLHTnBqlDWMrXqBpQGV
M3BiF4yTZmm4z+CezWShzZwIdtHLfiCg6lVFVTll1HsBlih+HLFwcZyXb+Sfh6FT
DL0zuueD0PN5AojdWIeJ7Ke4CvlSNIQwUKEP1rlsP9WJg2ZWcJtNWE7w/VaFqP5r
NUmZj6JdIIuaPXi9vK8DaXJdCF+if3/N3tCkZ5fmvDCXrZqFNevG6S4kDM477KQH
98Y8f6s7zihdjWPA5cU6l6dlvZFPpfCmdmHNSmn8Hfok6czQiV3J0IgERPPDC8Ol
4V69m9n/EHPVoI3mx2XeuBbLhvY2l9BXJBGU4DKnem//sxBydhtk+L7kJPlPCpES
OhSSxK3aaZkf8/2jMTEdJG7PebItqOgAWlM4Eo60NEg7vsiWTWrqq0sMIOQuwax8
gp7ZupwkF4KoHYH50DjSht8RYx3KKXZxqRaidwJ0uFGsa+3WXx2gjzNzKzkGDI/G
Pr/LH2ZddkDkiGnmKmdOCqAzD6aH0X77qUANOL9IaMKU939w9PI0lfbstHqtGpUW
hUX2Mv+PwJ2nnLuZ0vkKDcfIxFYW/fwcT761chU9W3ZYKDELBjhzszHjLmdVT6X/
4VKX45Ouy+G6Fc5mU9SlNhzwMtinbhoap4W+Hr0N1nsoegAklfKslUbTgj6lYGRY
43qfd/4tyuRU66buql2EHncucUEbyWomIYUhUJVIM1fsgCSMTf2A3mo4skSAwITH
jHTsJ6SBRZoGWBi85rS5cArq8EPUCt5PzuFVDyrvgWQU9gS4PsmKATYTJjBERm6O
v78YOlsn+ixl1cVfxKD6q9dCHSvoOknqq3/LrU3mfZ6yaUH52e9fYCXXXxdt6bP5
1CpRg0OgrCiEwxfPhcu6GCPjtFOvW07NesSzp1XzO2GRBU/ty9RJAfua1PbrDRC1
JJxQgoKKv6o5NoHkxek/a4LldXmbAFkXFi6JgqTllqt3unKMs+m3wexkUeZEQcHo
b6KEKCnzBULWzZ/D2BJrQHWp5DGwkMJ5cFXUxSAyFZQ/IA3NW8KCJLPLc2uz0KCT
w+/xyWWbAc0RGY1lioaWHC2AuD1bFkZHOGKsZNv9ySrDdJveyYyzua3kq9KVaffD
tYsWhkfcP591h1cSXzfV3F76CP71PQIifpjdgvPdBXZQzoolP+35lbbcUsr7fVXJ
sYyrNb0IE370L/WQLH1GuZhtkigHTuLZPB1eNL6QJYxbdsWKPP1U++C/+5dFIjBM
Lwv+PiH1s56qMvwJvYMvVmrwGHV9h4dlQw94ZezZ0kVU2MxkXAW4+xfDGMWfJv5T
RRmKSnksO4NEm81o1JaljxsAqfOu+Nzcadhs/QR4k/9aV/a+zxxHlBCuy/9NI5nD
Lc3rtYbI4k8VSXv7k72YhNuOOovXzlvhicNseAnZVM0Id376pviQJgOFqp2eI4/r
4Jg+Zer0N+5AVQTgu5pdfpszgcbnnR+cv0VIm1GVj0TGW+PG1MA61E37+uzowukn
MH7VP50lRHP0rGAmKGpr04kFq8GM9guxsaemes60M/4GtY+b0I9eUB0pKLt+Q7JU
fdYBYFs/rUu+MEExJWQMiNssT4MPcXDhMw7Ry9XQQgrxRnefcv1R9QPbER4bk2YB
BeUcXsaiFRKQNp0UGcVQop3/+prFt1o6K/ikQ7dKzfYPeJLEMENOCT0grvIAsaN+
38udyDUxT/ggPu65LmfA/DnY26tikDPXStCvwiBZOTtzHUzSVy9+CUkW0oSdMa9C
3xmFk70WuGDlGYlxAgRumwlv64p+yo8VSvUyOPiTiklWxVslwZSkXcxbS1tyhdbd
zgF2SK/Kg3F3vu6tZz2q8Dwulu1Xwf/SYMMbJqPHBQKy9VwozdD3nyDPJ5usrNwo
siVs8Iibl09eiPOcA9CDSEpi+R54BV7dkCJfy/T/HTZ7NnqNerOidO5szbxSrMlE
bd+bHkxp1P+4k/gt12Bu9DOSLyoDLb8As1UvB4zxqK9HWriRzd/IGAGHmUV1DRvZ
iLd8b4fngY+HafdJSXtMi+XOa5+q1hL2mvvtSEdaVrAVE8uVLyQQKPTfj2pvZwiI
yXpgXAlbiccGyKDnTYzxSuVzcSienVP0GL/SYyEokNP2kpDUO9NwurWB8ObYgM8d
0QnwuLaD6EcHK5Atw+eAvt8SGcODxfTzYuqqosm/HaUJ+ggw0gN8YABvtlJJ1x+N
68CpTOAwTIK/5nj3UNTqtIxDT53K8OlMbpeR55K/q/Wq4QUrs3PEsDkSDTdq4JOb
AH4avxrL/7BowGlVHb92iwhTduHUExBcBmd9uL0whyDGIjvVdZEIvczGkDE4oJ8V
nIhZ32mtLRQ3xFnX5ZHRP8i1MmPzkKWeRsMcvwzAnS4Y36nzPsGdQqe55qZqOo/k
ID1adZHq2NmAVIDMs36UZWJyTx8T/nUW8rVWqmn4fsWh9dwLXfNZsCR9p3mQKFr5
406Ia6ZjwsISrJgiDvaihh6AYKb/wW+xp4dI/J0fzfs8fKdTzMonUNq+0A54J4tE
iOyaTxIhwo/qtrI6lKpAMk08s9Jkfgt0X1NZ0j6edGoQeBKWl0WsR6PLo6bcC0Cc
S72giaRlKGDr49YYbEGCb1qQoR/kwH2LMSzjk0h7wMw0LFCfBSbGVQWhdCELrx8n
OUQpuvsqoedAo/xJi9IVWe8o0XjAHVIWisdh/RBP8k5hf+bTupfM8V60a/cYmccu
MYVnCuQWgvT7Qp1kgu7lGb41LLWqYuWWFeosvvq+RlRL8jmf2uSTbQD1GvatUbVP
pZoPw+n57e1qbo2xsR3ze5lEZuNMOLMg66nQLmsG6FYGB8mMo/rm8WZZoDDDJgHT
fZoJo6agkH0Os7+4/2nRbEGWxBlZmIFdBge1rFzzIaWNdmMwA9QNUBljCLBObx+3
MUwJcw78hEqzOIDTq/Aq2WL3sAwXNcehFzkLZUj7WqTEBhGEYwU19sy0wVbqzLe/
QRffYAQnyRswA0sfWzEsJLHKMJpFZA86jpnRZJXaqglXZTFwlMiTuybGxBGjN6sS
OsrMbpOslG2aI9q+2u3LEDNJjP9zm2dkwEFMgfauVZJPosZjreldIKcD2KTz/oFQ
P4Hm08ixwMfkdAt3WC/PO6uoQBR2lrYgkNIMPseG3bu2z52JT22TQ6AeA8dMmT/a
Ld4ao74aat6FTujiS/l4hjNTINPrG+oBlS1XddGBtHqhjdSsNc32IwQF6pEC3sRI
J5KCyvoQiVIK/CTSkNqmNNB0Yowm3jCSmE6EEiZNZ55euR2InZbM2k/n9Iy0Qq7N
VsofLgu1GqJ9Rlo/77Sh5qSICV3pR05vLju7NO//ulUbYumg1uiQdXZwgKHZntYN
BGX1CH9k2m5uIVdygNtJlaU8ZlZiIe0acLvrt9n9wmqi3VA3a/D4W0okUsUiQgxR
qVmxi5F3SJViNM33DyOI8JaE7bbBd62qQS4z5ba/A5nv307unJGqCTkFFIDzF1ht
QqEqMdSALPfWPANZPwx3cUiEJuS2MpvPqy1oAjUXDmymwtsiO8uXttmu2XfomDmb
Qiq/ATzM5e7JFeOrv5eTmf+D80UwUCKuM3xXXJLOn2aUbW43mLzZSQzfi4v8Kzmp
PaAQOZn3c2lq38cr7MHvrr9jW0NzPBVi9fXyLqvMmMdemSfvuRCAdD4xZdOLXxv+
jtpd/8I38skmTfAiyE02iS7EiyODO5gvzoH0xz+T1BaFPsVDLKJ3bGC8sS5XxEj+
TRcu9QegSbasl+c+5W/Vksx0P5WLgHVn6w6PBHvW1zlP6gPHmCqT/PulziG/wqXk
ovqUFbdVq+SQa9FET+nQBoEPU4wHrgoNejvthF+i9fxlWDAjosKyUdsDkSuodEog
kyJgyrnHFkcC5idYjlUQejW53eaK+HRl2dY8Wo49djFJSbfyH4SvOFZcdn7Gl+/I
DIGB5uu21qqXQjJ6WTE0OMQNm9gypZqYBV5FhLDsDDhvId2tXFoZV2roNjWSpqir
eEiDMK3YQ3+xoZ8he9D6rTpsjovzq/J41Bre7kimBEMYgYOTklQlWTK6J0gLGPjh
5or7iTiYSYt2q2EfEKQjgQdByaDtQxl1Esxx/lZq7nLECaB6gV3R8DopuHo3y0/L
27mSAjAqlRXbGK9gjrw+h0dMqWR5QZ1MYqpqMzH3d8NB9cWw6hODdz/XaiWZ+mCZ
Vv5gJ0lNrgYYXxpZ9Hb3xTgg4kbfpXoigrWsUivt6YWqvwZWCKoQWCF1MChWlt6/
h7wLU8QD4CSUGw41PLi8QDeq38ryZsrykotGSWgp/uBDN1YhuWG0SVDc4M9abnWO
p5RRAz1yWQ4+dQ9QnCMzocblFsfi8ryZgcEpa57IJ38XZ0+VCm8wwz7vHvH5VTV/
PdgEkA5CSmW9zi00rDg3Hb2SaMBf0Ui6nclhNO4rBy8MhvIKX0E9q3SFEBbpdAD/
dJOip3tHrQkTjjuYAAZ3hNoVd5VqsPtfNRP29VpFh8lCQjhD5AaoyrroV0YhNZFu
slHxET6jashoLKL9/EDQCNAArlsWk5v9hJWT1fyCfV9XsCj1MFkiI28WNJsXr3OQ
NvcEwJnF5qV4CmTdeieJxBvzQ+2kn+0fAnMXvcDLiG7ZT/NjTMUkoBJB5a/v5f6v
nMtNsxfQjz8asbygmjeoADZt2PyRl2SosLGn0aonmXtoEcCs8W9TeKwvceZ2+g+o
mv4St/ZKIcuc97NDZWZ+a4woOxjTqXL3IQXnONZ8Pu24Gonqb5dl4TmqVgvnTlCu
RKSFWGvVJ6tgd9y1cqaI8uiaWpaSOu1IzKnEcs0jd0uMwyajG5OwXzUhWEScXyMI
bTB7eDBIkaRuPJEmn01xTadk86yfTNlzqLnY96nEVNjfouLhalLBXgo1rlx5Z0/k
3YfKnzexgmDLa5uVfkwYUxjmNE6jlSgT6gp/+2UdvfRkAFgXI5kAsl4Z5KyXSQxP
+kLfZmmnt0EkMZ3M1B10RqCXg5k6Xod5GQze+ZqPuqF+4tX2xQReznuoXD9q0L4C
vi0oTLdBxeKr3szP7dOhFbKEzoO6rSJhU9s762Tlq+1DDUnQtix0G4WPE1AMDD/p
t0TU0QtsdPJLxaNihOxWagQceMrUCkl9WvoqMNr48wALnVoVi8SJdg4w1/hHhN15
XImRsf1FucQsnktng94hEPFWoZ+23enA1lMaZHRwN4+wKCkcfHTRE9uxM3iuvZgT
F+VYvcxSpa5V4qxSz3UnVdDe6fnfDgI6En/oucyu7lTipbIyr7XuCXZF6RzX/gh+
Fbc13GGoAlMg+7Ch5rTbYOyF7TAKtWR4ul2SUtI3Z7+s6HeB1XDbSM/iXsbwmJBj
/t/i5pTRB6A/RevOPUMJtx6yLIsAHg90CBDLThTHPm2qXOd1FZR09/PpAbCCnaU6
lGirpnSZw4jYfp9yre+BsPtiKjjuEZzY38UA1zoNzn53IAqWv+nIdHGE5CQDHrOr
QJb9tR/LwCHQfyfTYq3LHA32HZF3Sf/odgxFyF9qxHq841AgGRkunM7N6h9PRLaz
MfGzpCN0d4AILJ4yQx20uh1MtrVkRS8us/PmwsMFnpNugxzYQZUojMn+zuIWP9BS
MdbnwTxL0rqCTQoRJLcwPqd5Bb3lMaDjRxz+meu0WvYk2sGpIqHH4hZwcoXXV8ZI
NozAkzR5U0QNckrmL+WZkBuwofP+HNEURbxsTSubEPHfjuDqsEuOclRqBXmM6iNd
ZK9F+VXTWEbdOclWIIYyHjQhK2ex6NCsS87aYeoNE2V2fj3mHa0PojWdojNx50qN
N1BuO6eoGNf3GK442+Wj+8wt5SEiaTDqpQwz+BiXSgCZ5sX/kjSqDwpon8IeFBoK
Ozf68uxdalif8sgtLqLcMNMnj+jhGxYLVp6nIrLyN6cNcxaUpPky+BPSas2eeGey
Y+RtC6G6O5X1bdkBjAvzRkME+MKrOAmBhLnyFG9l8EjkC7vYCFnIcKuAigeIwoqR
X2ES8j0sPJhhvSWkaFU6aqyVG03eXyJVcKA2ztBIpGDDlCcdyVZQbNC0sebQv7QP
If0Fwhs/NrTNp9y9XxyZDD/O6+uhU7oqy+suRwKddAhbzC9TDCXLKgsRqU3JG9l0
2wvRj1ySl47vBayJjkE+h12dK86uG5OPvj6FG/cu3R0QQOoesSm7/ndujFHWRCjh
Oxk3RVvtZC2tV9AViRUpsz4vgdGJbe/dVUmG2j+WQdONR6up13lQ/Rozpa5/HcUI
FmZjAlji6u2nZpvuX11NJussPE7OxfBlsqg/ImneOG7YxN71IGRjMyw1nix7iBc7
DzA2Gxce3QyqXlmtD5PJ/vLXv+aReMgb2jzu83605UG3el8bNWYc58Vi8PrJerWn
FMuvaEb7d0ClkpiNstGgyZMsmVvQoajuf365A4BBdVXXOEdakamk0QaSTabp+dL6
4wYQHHFn3zqGf9NElWfQEwG1B7GM6frdIKZlaVbuwkilJgfxRep2aBVoheFB+w95
eDS3KUM01Prqx0ldlajT0w2J8YysacWjiq9CeauCQnfu+Oj+9LyEODnkpboijxyI
SwY5EGKg+KE2bLAX9PVa2tQVdJlRZi0ytNejcgeJb2wWNZA/ea/br8QXd78hmJ7Y
1VZo292oWocHLhrrDJHClpwxrBjefkFlFXjcdkk+wCxG5pzHj/9UzlqNYFmr1jR/
7q7RyVkIImoBNEfWdZ9uBr8i4ua1JGI0bxEXqHpPhTdbHzEqNqlhQjugE6rZ2pCV
NyfP9dUYkxt37eTX15VnGkNpL/3OvegrugxP5E60DWaYd0y7Z6scbBm2/bPA/VN/
aBDbeK4+4Jc7LWgP/EpZMyd3Cnkzwdjc189yXHXVlWnhRgEWdPcBya1BxrWX4y39
RtbPeGe8gre+/2k6IfqG/6SKjVJci0v5DemSXpht9mHLqOsa5X6jU3TYye4SrNOm
78JR3FcgomYrsa6qQ2GChvZJ1OanNhXro7q0YP7lBkMtseLjUj/YLUh3wSITfQAE
0Rtl2aGJOVdp7AO6tH3hBPW9BDfvLCzy3l0J/e88nzrRCrOC7JNZdUbyiZZ5TMbB
ce/Ot7X4Ka/dYN1019BFpWnBJUsNTaT0ztQXgDz9gNVSq1PtzctmYx0LOl2eNl1N
hBE5keXBuWTf03RUfiycpIS5fZw/Ga8Vtv5YTluPdEG9X35RPOdDz2arfFuUVDGA
YCntPZPrAZhfEGZnj4MghYE9wu5C20pC7UNRkAqY/ZLy32UHOxwzVJGxdG0LxuI3
wmt+5dyfnGThMnL0zUwHMB7oxfg7XygQfqF4aO+iunDeb9yVXuyzL/LBVv8nVJZG
FyvfPfUig9FCHtAWiIfQ/t2gc4dHZoFhZq8V9dQqsKJgRl60Y5rXOGfBnjdzyfvP
4nwfhXcxO1ViO66mTQwKG4yRnhKqY7SGdvLZEhjDYy0X69lD4MD6/U6XyB1fOa4d
LiYKQ/TRhebPaQOPNDFrXIHtsp/KCBtg4Mo+keUjy/pNOhx//pTc1r/JHnma60Or
Vyd8I6Eq4ujnhKNEg9z1DMsgHXhQWMILJPA7N4o/hXnmyb9U1oFSmZH0iH3SO8vU
YdVAs0qjRKEeymt9EhZmU6YuV9shz1Qwr9QoBfi9XD5M0hp1+tEFymOWybAFt7hG
1jIr9B4/IlPKgCxP4mVKMWPOwN7MTY691woqrl39ATMz1dWb+MjRyYwHj6rWiw/q
6Eo86IUDSpLbcXZYej6EzJOoG83o7r3AFxessceORFAS7ggbvnW+SfG9TAEDe6ng
tVpLkp+9eRrZmBoqpPGNHgp9ryk1pMS0zG+vaDezRPBWByMupkSoVz0S0GU29++F
f6xazan//z8WT7TQ9M0BkBwQyesV5hk7ldgTN4JCgTqTGa6Gr1zyBE0ImNYQru6R
sZ7B8Y6HFb+qESyPUfDpQqw4oQV9Zv58L7jz8JjcNSOzoDAZkQceqUMo1Cb3n8mO
4gKrQsuJgAuYsONfRopgWlloW13tFcAH7DG1NqMkqMIWrUiFxryqdRWCWv2mylpX
qP4jV4MAnfAcwniw7f9mdS/IHq8l3D3upe8IqXX0FwmOPrkl0TK9aA3tqoHwAr9S
C8Y6CuptwxPClMTUSWkQyTQxdTgupFljpU/RzfI7+XXLXrZPDU/lZka7illGtASi
tPopy0hNDP0T8vZ+SWNd9DdZ1V5DvDw+THWCuEU91RycR7CXOf5AzAILN5Q0DZGv
sDvTBjyxURv0N+FTns17OhKKRmWrLqNEQNqZtBKxJAOiY6+cksD1N3/aqqenFYJ+
u4EK3o7wUwONUW89cohLCyUwdEUb21k/+TqsgWnYofHZKdMj2miN/3iOnvVnuq4r
utICN309L8KxqBGGUwbmBQ+Nqso+gOKi1i7apQeFSlmNBqmHdy826b1uM0zRskU1
EdNoNmoJFkYhcBM2HGaehDyp7j9WALVvbCu00aJ9eLqj5G9cEBA2KeEa/tMNRI3i
4chef4pin/hRYhurVzRN0pk5We+a6MvuY5o4PZJp7BVuEf30wMeMFVvbGO86RSHR
vtI43lhY3uPLW8F6K9tUmwEKb3Y3OI7OaE+G5q99MB6bliJIORDEAa3XjV/BqDpj
3NmVIMzYGUU/gUPW1FMQMauYMs2LBtsTQC/Im5ip5OwH+IbTk9YlnHQobuutyYUi
ofIpcABCmpGPTfcBb4f/XxXcwYdETD8+0rervbMBKo4yi7xbRb4ENp2+XPC8cBP8
sP2Vbz0E/o5ZrhjYY2U4SPSWTSphXNqQ8AtPlxJdrIGVmsA00fM3ivImbgNeXs8C
EDWNbVb8oxKMJ0T0CBI+dP6cO6/5AvT91UYofPE9H8ML05eZS5cFWXgcBOplK8ix
oOhbFk7ZqjPrAsES3LgJYqoPWhJYQM6f5+srdJZhVMqXqxlsJHAAUS50kJl2o1VE
f5Kf2bka03ouk+rRotgPq5bbyfAfBab2c1uUcXj7lsL57sSvNLKyx7qiirFC9Udw
Og/FAcOjKJgknHKSScvI38f5RqePtBipYQaoZReIuqEp+p7UZ106xnE4+q20UIug
hspHIHqmzSmsWwFrba8ZqgM7vcmrUuEZI42kPUkMNZvzKn54142RV40OZ9+GXx5p
AI7VZ6YfMLdAPRxumrG348hZQW+E8eqnFMuuRVVp8dNfVN/NTKQFxSe2AsExggIJ
JfRKjZUJXrwDK4ig4G1/1fXmnorafsNhiMRlTTluDle3qrinuLElxgpE9/joKh+R
GjtqkDpZpTQHVsPS42VaRyv51NTZzOSjQEOO+BWNz5MuahC51iHxUhzF8h4t9oMf
ucA+nONgWTBTbZ9BnBx/shdJhix55X3aVHoIhtqSzqCk4Zt65ueOEImDFMW2y6nz
MBI36Pw7OFELw8a0FUJ9gyYPnKsWQjXPEt6cUp1OcD1y8onNLG1XdV+Sp+nC27up
G4csDZI6taKy22WZ4Vcxnnq+UJhVtSv127166bO+U7Dh2CgUoT/GuZNw0o8ngKxB
gJ9haBxJSnFeNPRz1V5i/NZbreEg2bbKgoAH7XefTqv1ZIoq+ykCnJ1HO5Cj0Lh5
dcrfG4V/1qlsmP8QZgknDl5yanB0T45dpWOM5wvhI8XF0EcHmXNtgNf/eo8ovvPp
rnDdrO/cZuOieUkEHWk9B6BF/kuI5NjVHueMa4X8WuFz+1jYadvUSvlDt4b9hEJe
PSTXiEuMqidunVwKKzDGUNCEa8Q0RTRjZYQiuzv1Wu+GdC03wGfFFCzsDBAdmrWV
/HBbui84PRFdthhriUoLbF1j1EGeIN6cJrX9/O0h4E+7et1Vs3k6BDsuzcBcYOXs
gAl0uaYoFBeQyMngsy5GS0EdCchyEFk4oduCaUkkN7U3pAWep0WTLqUPaw3lk86y
OnPPqPkiMVTazqccmnknO8z4gCg8312SO1IgpouegYsMqXSMwUL3XoIiC7sBIxQV
S+iTTXYAn7v+PyF/qJ6iDtIWiCg9z0egGpT5RrwqbexjSq96dy4IMLCjLCajScce
510LE7fJagGvWUNVmf04GAFvHtkw7O2mhD8As6LWR3pHcssdfVtIdH/UVyrW5FkL
esLHRs8njReqKIJ4VmTqMGOeKSqRfQqKPFOouY5TwYtl5ce0f9T7eVqZ/V57VXD+
e4yXXc0KMZObUSWwms8/wR8XIPB6QXTZs4Lmo4FmpMPuH/MQrPf1it4G079rVmzr
6Gt11eE7vdoeavHMyO8CrTwe1BMcG5OBpPEbTBpYLt+2lztirgN7tTrZvG6M4xAM
nqp/Rvy5+znAk6RBiY609O+wrmyRp8GkTr4VCsNzzYAphW25DdJpzfjkxNJKyYOd
iPm16KkWdqMkZ8Jei68PLPN+Q8mPDW0TrEM0oRGZEWW4mgoPbhlmdljJDMUdkBKS
cs0V3bL1+khVYpt54B1KYY62BX1DZs4AT94S2zSp6sM5oQ9qeO7lhmDYKNmnHW7m
YWzR4x7YKyVThYtgiYJV9aNbrOCRxmrVJZlC9hFF4bwANFDM//XEqzm/YHeRI/sK
KRNPZnLKzXAZahzh/jaCe0uuZfiHcI+2X+Cm9SrWYMLXqAQr0dqZEEL+pZf7eONh
LwmBM6Z3sbqfY2OQ3+7xMC+I+O7Rgt+83FFx8wiaFtKGh+BlyL8QKR1yzm1Em9tO
cNlV1y27q9sNZCVZ3grXRNtyXhkmww/GUBiglLqeu4917+uLTuQkmsb1gRP+5rE2
Oegj9xd4czb0/P1ZWEa+tO8t0fqE9epC7uIM23gRbE802AJsCBq3LCXaewTQtKwt
tvH8Juza/AjJHRjbyzxsTZ26rYqy70VEgmhvWPqmkJwf5rnZXnakxy7sqXCxckme
MOZfiiotaBefI7uhVbLsj7b6SfjGjLP9hMtDTdNwl1uyYyR9TldxICw+lmtnvIoy
V2kpaaZkuV8KkJv3D1BHGKwsMkEjVgjaM+t6xTVCAwB07HaSKCZNkj4pA7WXTQ8n
HCAi4jIVFMO0NrlITVrQRvzqLhm/0lTTrvIG5WCT+9FjCXnyN1wYbsiv5F/bcm6b
/WdYBVrSsPS5sk5hVnrfnGSV9Tymf5wIXPaYFXISsS5qIDknGX+zQ/RO84ZKOJ+G
WgdzpycpZtXKODPCU0t9Dk0R7UI+tyeHl7a1OjxgGxzYpXfUJsbCjfm++HecXD+6
qCl2Y6P7b4bvCSYEgdz64m3lSXD/vWfSpTTpsA7e3vhPij0camXWDR2fhQ4rrOAA
1knY4o9an0yZZhdaxz40AxrnqGUM4x8WtfmMWZeYdemfg0gcSRmmHp0dqbsCDyrT
IjsHND9defkRzVFl4A6TkODNE29xAVp1TyuV6lWamnMMWooZwaNzRPQru69xtNZ3
waI2Ya55NeoIK/zaBF7wrQZpE0mIBAnYx+8Kfx32qqoKMwOeRZIq1ImOEn3HTw3W
4Bu+wytTx6tR0f+nR3CdIOZmZ76VEJOt6rg98C7wjnGr2t9O11+q+4axMzgofQNZ
rsOrLIqbl2JgHPW9nq2jskqlyZbNrBsdFKAKVAwMzw68DSZowpr41nzSbuk/jPq1
oXwbIakRxxWN1/lG/i5M7FRoXsfH5IgOiXWp2RKyJ0KhuAsfFZrJECkZBr7U23A7
J5Qttagi9X01JIhrrRbTd0CH7KumuiNpwsgdy98ZjmgF0wmtKtuCgtQlktdsCcnI
M1TxkCnaSZ3kckkiBdkQdU6w8wZMvZhOrgBRgA62MVlsThFEoCy74GbtncPFkIOy
pKCB1HiURywPaXkiA6kWXKDKD6AVmwiGV2cW1KzWyHKeIxvWsUPd0hPm2vs/e4fu
mALDocGoU2Qvdg3N6YWW7xxMiO/MvAIBAl7Sr91LChAMMeTthSLx0fd7y2TTO8Os
rWYUM6DYz1ypD6b4Siq9fMZmCN/KbygaXS5ljSA0ssldOfqAZGw7xmIsiAD6yQ8R
Tj8/gRjWPQcdpMrI4yiT13KOaoiNChyZP04mcP/OqQ1MPTjykkk4EAQxFX6SOy/l
mIRI38llYCCKA9AWDEfFkm5LFk8dWr+2X6K1YaZc3Zwwn9gJboH2P5gb+EmSwznr
sjMmiMxPkjJQ9jF/imkiPYtvt7oUCCWoqkDU4gaeHGxUvaFyGr5ALg1ZCOrSXXki
kMdw3ChZYM6+6/iUwyRHT3rHcaRpEdqkNtiAGocDbgR2NLY8Y1lJU1BQh1MV4S/W
t3uNiiwNGDJtmuJ2twP2d3wW+i2Z/TAdH7rDPj3UYdxgEislBI91cUoup17aMhw6
7pRscikPHa14jC7cRy0BhLEnlsEA8J8Zn8YtMyLx4FdF9LztSfsl1zjvcdMrZNRR
XB2LB3xUWKtgeqZnL95I7eSFIO0OEWGm9gA1v/5N0E/m72FigUR3JNCBzxtL/VIw
ax7hxYF04peH3FklvG+nUDGiOhwfv6/gbojnlkJHkuh+53xh7fcW5EuAklc0Lhqa
d5JMbGJvFjF9A83jDlLxcQqWtn/hq+2wK2HOoVyeLNmJBJWSZb3OYvonyvZL3UqQ
jamGOWtiWXrK/XCU7pmaLhBlMFNwNKX3RILhMX6S5WdyHHcEf2Zjbu63Mc2T+You
nUtLiAQ9iphiOjyRLkJ2q6d2e1OF/3JevJX6J81TtPSIwJ74BS3I/JTaISsxTlha
VmCI4KCWkxPn+DCKD40q4v1K491tSw8PLZJiNvRa97Co4zeNNPNA0shw+RqLS/TB
Y8snuwKYdUK6QPTsD2hJjkMMuriMLsMr+j6exqd7qP1pGTnsWdD7/w6ZYXt/miFu
qel3VDLYM4Rp9I/wT7W4nHPWuUtUN2Naal133fehmoEh43FygRBKtjcCzpOL+9K/
3AvPv6/a6yy5ArBDc1f4IZhEqRumZ8VuF+2C3XbKeGH9eh/NeGt0/nKmDD/UG/aK
4NrxlCMHe1liHG4yZ+gzvD1vOiORZoad67/cncKUwjKd8+4ZSjgs9i8zUn+Yd1b8
pGSZYB8orXfTD+FFfUORXwE8vLCNas8yo6YN4N8Px/WTY+4aaMQs+UqQrKC8Erh0
WH3RWEmzr2jV4ntqZHveiLKQ4d6NFY2XD+sLaggu5YSB+mczJSDMQ+ParX9/BrBU
8TBq9APJGJ9Als5HA1QQ+x/jgeiJMkHpC918nPTUKTrkalH2VKQEUWCX8ACAM2Lv
q+6FY12ddjqjDeh8UvfnzKSST9lxG+FmDStH4FaEYYZH8shb9zsrgK23kBVcYOCt
KJVN6EaptMviJ8vr7xRDR7JxHS5pvOQePPUb9h2EJ4tWI7Nsdzn7cU+JH+2bRBZf
tshH2e9UswTxvBoooS15HWKs00d0qxww0/trQKPgg6TCRkJO6B0Prj3WrFn2lRMx
mMBhQIbbFc1xZyegRm8JxvUgz0rI3wsJSdji0PqEx3Ol22DojvGwsRJ3DzQLk8YV
NSN+daHYzFz5w/eVFgC+mSsCQ943f0SFRxZ0qfQUHyIM3ehPt8DHkrGTEXwqJ90A
lopY0LOt6/Q8zOvG/jw7ukVbDYDRiEVTS19Gt3vhcStoXMq6webJfHwt86ZgrnW4
xE0M4ZCT1ll8pmG2RtbLYl7iCooveJv8Q1LhYedrSYawJFlvZKM1LjN6AVagDIFA
+ul7J0Q32+ifYlzUViB1wzn/eJiKvA6uizz9JiKtN5nr+UHyRHpPEV3C7HaVyn78
4YZDdWZgnAIUW1sfdjxfQ0PFX6F2m7stIknx9VH6gn7PZMiSYJ/dlIZqBRzZCs8r
6Gl29t5IJkYMk1ZUrYPankk556fLtSI0JniIiSpEHyoQZWnjv2LappMlJ+KwfHWD
8kZmyZ1/cewdyfHYNbOP9ZBOv6BHfc8dQ64ZftuX3riWlFh9ZXF68erhNnpfjFZl
d8vrku4uCCuvr01mWclD95ejc9nUDrZgGRPyy4oaLvK2WfnXjbc7lOGD0OYUlW0q
ghepU8pEEM36wwKw68/hkCdoG8Dd16l5FmzoLwZZ9twU9zIyPJNts9CL4SFJdhEQ
umtPdL30rKIJs1bsfgnRQfKy4De8zzX6An1heuSQzkQylP1gKV++OqCuQGRiNAPX
u0uBE2c6kJgYwF4VBM2Km5Vf+xVoU87wd58EiiaLcsRrd+BrvEBOHezxrcLWUNDi
SH8WiZKz9f99IQSd+cmwVPYqyaSgb3gLJAFSOMDJTFnQvgMqlalldiAuI/OxkeXL
14m2POXIgpoY3X4DfAHElaoZITuYj78Q7oyA/72kpYbmhgvPqsRO48DXob42ym5J
M7t1T8LrXF9Hg4nvKdKYkMpAckqlQwZ61Q0qjPKLKnGAHuHzKNCQR3kmFlMcjqcl
j3zsDk9NRGFUV/1iGOhn2vIKtXhFphj1pjDqcO7bQxFFa0AEmGrZPJobFSJgWhZ2
g/X5XtsO0oe/CjUiwvLA6E7kNHk/hPamsWG4D5zGPGZMohEVZR7t9UhWkRm0d0nB
Xyn4ftPFmF8crP+9Ktry2+K1Kfw+9PaiWtcuPEeXzgt2Dyo0v1uSPoHBQzgMh3Hu
y+xUrO2sQ50d6kVPQ9bo1uq/F1fEWljKqFHZYXS6lQVj2Ea60gzfl3F7jSFWoaFY
R/9VqGSSjv0T9ml0jWcBppXoYTy5V19NhKU2T5VfXJ1wUvGBXOwY6O54JcfWeZua
2oQqp7JyptDTzlOkjR0tefH1oRW/8PAdJE578C5PvkEHkbT9goteSl4FQdyN8ruL
IWpDBgy++RkQjJwzIftZVAlbJW+xYJHFMmeFZF1uaGFq9exo8fFQHWmBpAI4MtD3
gZaQjuFwuW7EqF9sK70LSL1+qqW3sY6dLh0+PXiIondX7rY0y2irO/4konqud25c
y5ui8n79IKVdLw1e93BmFOI/gNOs137Cyc7Cn5hCW4O9SLi2HnSjoaYuF3yi79LR
Z37NBabOAdSh0K5T8HhIwYxxOiK38bX0gqYISldulGwcK3Cq6AyCwAOm8nivzxWB
r6wKGeA5NfQt7XjUxIA61bMU433ycQjcnl0K/HaxvhZBq8nx+NePqPwHplfjyweY
moGBe3UxN1uALu/8QawONV1PveltYg/xmoksBprOct6Hc+OV6jOfxE10sXE7Vxlp
cH816cAvI2En72VgWW3x2LCldHrYsjaFBct/6/wxXNDbOFqJx1poLZnxe/pgZcaX
Crgwz/uRFMWkjgtJQS2kiFnop7V/7MNXR7Z/CnoZWaVB9nd1J2tiCm5+lUy824rP
`protect END_PROTECTED
