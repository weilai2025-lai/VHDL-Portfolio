`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1u70mSAXhK963b+UFTRLztDEQa83Bz6SR6abWEJqANsb3G85/vBzCbp0kJ4ajjj1
M2HTySqWShPM9Wfdt6iAMZwtZ6BGPHrqRzJuO+Vc39VhfSGA9qYNZPpz31DoIlj0
hukJx4vweNPj8r5+FSjHJbFNdsYM3wwgA7fNnSxL36CP2SR71IXYFbNCxM388EgF
pMcpFcEISJAn1Wz20ovq60Ws/cN8vGwyanaIwrCYb2tJ/lvvLK8/7bjuhBxI3RZo
+8FpPk5USIJmfDrVF1UbASlWuTwpoFYzvGdIm0vL2gDSVf31mEWoQJU6r5j39FhH
vf8IaQDOiZTsiATLsgLg/Jdf666/Nf/XiYjpTRc3pMLRKgF2sNByct1YGdJMtpn7
go8Vf/NOVb75Adpqrq/eRXpBuBRrjXjRG8Bq0gs+hj95UD2xwFiRsese8Bp1CJBU
c2Zx+ll+nwi1iHMp7lzWpwBg/6Q/U4Haof3V5b8lKbpNOUEPCG+wbntzIZpj0qgy
3zspCUxDwgEAlv7knSdCxPgLQ/yfncpgX4swltLV0bR2/CFgayZEG6cXLfARHcaZ
cOIoKEtR9Pnx8PMB03Bk76c3K+PROiqNR7byILNxeQ4Lae0OnEJwROvOrLcSpimd
21O19Nt+TzDGhGgFLNa4JxTBHBwDXwIRMPbsj83l9jenkD20Vse5tMOSlJS09Lc1
tXUYL0f2yz90z7zEx0XlkFL3+Vthq95eiyv3H9aYLl/0ZYOVqpY5lKF+Clf7njxz
KoTqUJ4gtVu3+DRMEdjayhxkFrUF9jAf5dn7o8NPQjMJTtDlZa0JxBb8si5LzJ+K
Nvxly9UvNjBLPtxd2hQvjfbKacT/NTqALYllAoathof+KcGHBCQdGuXcmq3gthZW
SBW3H6ArpOPZksWkG6NTbpZZbcxG4Z+E3QZiKPEqf+RyG9xAJOpuywJFKOM0hB24
n5VkBxV0MUSEh83/AHofhrLVXTuV6/jt/1Rcn2JZZmEyfFsjPCTEIoIQWdUAoEIn
Wb1S8Nqsjg/upVM3L99YusddwvK8NRxelfP2fvpbk1Gh205ZeKJu7xUqdnfaGa5X
OOyk8LvSadMtLPY4u2U0BIGqRcmRMwX6enECQMDWk2PhPNOsMwCsBxBsoRRi/QA1
p3kQLI4jXsnVGH5+JzAGOo4IwkcVDH9tVghufsNOVlPLhru/6ZXQRX6ivxcHp/pL
eW8rlCiBRcMY9Rx8WrYYSMX/EAfJxdW3mQn0mJKqDx/Ajl1P7PBd0YgPI1LcEeaz
yBslsu3Ouwjb5KkCAcawHRz79JCSnKW+msTSQpTgLihNQ5keU1AnI87zN/glQRo1
1fNz+vNEM59Pxug0LR8TGhxpUxCbWe66miU+8DSQihxT/tFZd3ICqjd8umgJQZGh
YJ13v25r/MjfrFRaKbf7HHMcoulqWgPMdxNMZwn7b9QJeEbC/WG+LdqCQ+gMYc9u
`protect END_PROTECTED
