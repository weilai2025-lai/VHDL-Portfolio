`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGdFl9K7x7uJ1q5o1pV7NItQ3ktu6eLVxbfrfjOE1eDuocsSN1n71kKq3obFXtTL
7mN4AbLA9CAD8hB+bFUxcrbu1SotCJZxDFZgY/r2561TgdPtdMznS2vAW3JiJ9dj
wW3dwbGTqY1UvHNpKMjwEZFJKXZDypQf/1YVYDRwW80EtdvxoYb4P4LA+OSTQzYj
iqZZDR3IDIUB0IaDl9NXgo/3Izb+xkJ6ggYlmyYBh3iDJLFoZXlT87BmfLNkQwFH
OC+qyczFtgXiPiJcFLMUDe1LI/LBCpX88OOmjYng315bl9TDby45M0Oe0+bBSBwe
zHssIuqlSYpc2MaNzOaT+grTFh9AEXNlPAXE/F8448y1raY37oyt+XDIwKvK0w3K
nREgBvn5XSjzT2Xv9jq5tPz/axSktrIylrf2r5G4QHbTrHCdqZKlM78E+3jdLuPs
Cf4wacgYmxGjqsXb+zN2qCDmQvJqDcCOnz/wVakk43Aw7jfooLsHF63oCwJfFzZz
eluXKlcxgAPEZWVTGp1UYwBnBa/ZN/x8DBdnvwO7T8sjKUF7FSSdsC2tn0CHhsNV
b1NrdycLtxNbHkUI7AqnnZmQj8dou0mlRW5cEsH/JRVXuX7ffgJ5vfnK1jwFAtRk
c8eTabxaXqS91ikdXohrEUnq1m3PY1FDJ0Qr/xAHggz43LElzdZEh90KDO63zO2L
GU64BPA162czQh2ZQIJFRBlEBkWsD59ycVtzt+AD1DRO6txN3vmDHy+charX4d6r
9/6TyK8nDm1KlPFqngwdUSDYwr4HW8DjEEUsCsVIzv5nM3xkfr8ggjchtcVa2pYQ
Z7Bbbi8Ww09FcTe2Dnr3Lg==
`protect END_PROTECTED
