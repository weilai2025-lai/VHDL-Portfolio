`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Z5UAbs8lPyO+ph00qcsZOhM8Hzx2gYyT/GUSujxrzEYmrC1LR4pCZQM0B39oKp4
r7dMlLbFWTp/8yYR1dVNM6aBq9x+RqL1WtWDvIXoIXXih8Bc5LWGVyDBJRLjMhA8
3IaJAKS+Hcj/VOmnlnsDRlcvxpKh0PnPP6bR6tJqUSQ7hBjroJ7qG3QKO/265OPm
xrAO9GS4KYnvXM1Igz2o+nkjrOLy9gqbYTMZJJAbZJx4wtiLG2yvxbBlxZv81RUJ
gxlBiPVmQkIWhI4N0DbifnfzqRjIBsNWG5PffyB+fOIazmlOE6QkdKPcSEYQUpkZ
iP7I1qYyzMDasuYtkFfzTkatHqUAp0ydAVxd6Gf/lScodXh+irgVH1nLrDUYnLyu
N3zLkoM68zcGPsJU7P5BFjrhbTo1ZvfFaU6JhSxIcDgGBcUULb8Rqh2//ucZ8Pfl
6cFwbd5BLhsN/FzQZlEAMnuWqX75YkHzUxuKbatgj1kS8BBmsp+WvCjSdnhbSLmt
/j8l0F4xRnKeHkhP2GJMJkKRGD3Pk2dpdRRieZHD+dTzqUMrn8gKj2qtoBdbBfSF
CHMQ/MGAAV2eb9dD6tk5v1dHvEZ1DmEK2PzEzqWy3p7Fh4QqHe+ES6+84sOuu6RH
NMKv+wqug5C+6rjT9gfNQKJihZfYbGqgfjIUAf2WbuJ1aMPCM/NUhZYQJ9roQ1jA
kHcLFo23kPRv45NyWpl/IX76zlD9OjhxdgMXXPD+Nu+A6uoBPp+AtuWEICs8LVEg
`protect END_PROTECTED
