`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjZh96mGQfnaMvT75fr+r9bxqtt4dJndj2xJvNzSk6QhG85PsTonp/BGJooWr482
qPb15pqqIEwItIWtlWyTFHTokzWVI/Qj0K4LQSMlJNB1aCEbxDDa9mn1GusnZfTg
f/Ys3fuMCjZwVPqjxhnGAzh3EDNPBILh8WgKDUBXPoq27649bZLGGt0jDrqhDprj
9e8dDT4Oudiyo/n96zYAGneITP6lufGUmCham1ratp0PCTHQd1y7EwrvMwJnMXzv
fAwSJs01r47TgR1Cz08/TlEUBvVvEgr2vSSpkLgeK5Keebb2mNQuLiYjFxJY1uaq
wi/t8OkZFYhkvRRWFUaafgpECYzftdCJNbUMAWSDTFkFRLwPgoftr7FwTvY/bhzK
vdScDaTtnIoNIkOVZUqzeOtUEGI8SouHfC3f7SExWQfOg/3SuYmkmVkJGRk1okYh
nAaZ7gbc01f2MhObyMvn8KMstK/HuYsf81aJR0RPJ3P6zgxoueh0FY0s97SCKbNS
2554c97Idjf39sX+8FiZ1olzZHmWeEkDcD1ibHsd/tYS6Zqqq9tCTmdCU7WQ7VeG
tl2PrlCSI0D7Q5579wySf56dRJ31BrTL7y/6ftZSm5CH5zRgRpk7jTkXTYSSyj3M
OmCAl0VeK/x9ojS/sJrS7GsFCnfZPmu602ygYIcyo1HjJtl4zuZp1E8S+ONXBZvi
7BnwCtwc450+OTmH91WppdbnlCbXHbH3qg96AnNR0cGYyS7CfEr7jO9XZI+1UZfr
Qk7B/wIIghU3INQeVE/xaCx7n/SOKNiTi61ZTr17ku6PLirRVYjMlGz4RZqwHKiA
xbDI5lFVUFYw8igk/xGstaVePV7S8eDf8XzX6Zdh2OCNkVb46GfCFNHwMWpz9Tha
TBHj+eYY+eFtwI+mPS/2TJ5IV41k8l0Cu/2+Vzsg+Eu5BJ9Z0btMpm4uZjkc919d
5X09hD6HV4MffGt+PDv0PxPXNq+cj45tLF3WcrudPTLHeAmZFvY8ROCACqelhQzG
qvFtpPRpfsPQkq8br3r63ynpX74D1T1CSGzhXUwCFJGZD3tU1NW8YvanLsm3th6b
yLXAMWoTHiH0plAAMBmZTeFxj/N8AUx+2PzgBTc2npibMI4x6aa/po1DlZn2NVSh
mK1Bf3HPGtP7/4kHNpkWrGhGq8NSDYYLHvbswtEY6J0ltYg8TMlP+0djZHNBlfoW
BxGl6cDx/eIQhxH4GaqaiYBshNFmQK+JbU79ZX7cIt7hMv6/oElsGxdCCsrMQv+E
QDgf3T7A9cVJLifRkjHkht15Whkubm76lcPhzA1DC2MUXAaU7V5OGHosf2O1GR1t
ePOQ3rt+wDjEhHYNlx0TQawKsJ6nZ2TPAms0yVJyP1/swFJfxu3t+bq/Wqyfg6Sc
PfVbDVayJvHPHd9mUeVfZlXIsRhhTzlcwq1uYYh0Vgu3ze+xCYSU3nr4e68Ax16p
tVyxRdmPu1CtAYYmeuOu/NsNWWIkq1LsDa8KebslOiBOiat39vT/r/75TkxPPm4g
aGUTBniWsJn7HxUIGRDnKQd8ZgZQyPMUdi69dOLzJ5fz6/3bAjcH1JOuM1/3vlvZ
HO+ayRFEdZjMhP21uc0IGFfV6Ht9yx4nJuzHO0sz67YV6tIdfkhMqmXh7eEp6JQZ
lhxnkO3mUiZBARjC5u02PuFkhWjzq57VrQ66bnN6wlM+el4F6uoto+lzSlkP+yYH
WaVIHSDW7FMWgK8u2ZS6GGGVgfGkOYjwwGaOaHKlXRzqU//56G4/FYxSoaTeSmQe
+LEtZZ/VT3pCRegKkktEeHLSonUdBptSIb0lIkARuOB03vE3H5vUAeaB5VSLYSvS
6DGWR682oNjZ0JlEm5v7X0k+SQYJ76W59t/jKnINVxd0aAGG61yMO2UP+f06T4wa
m7d98+OQ4XssWvLXFD6B5eRTu3Mizb1SCi+EqV219d8b0DcIUIORVk7pG8SIzFa0
8wNgtTStOoew9A+0FzZedJ2pz216zSS6lLzb+TKp2GxtjgLYcafU+N9tmOM48m44
zRJKxU/XEDuFZbEoqay/gN080n2SOU+whjwfqnjN9M18FCQiDAGYZ1COd+pFvDQA
yhKDL6B87NhPrrM0I9+Ehubu1kYx2b93DDAzrH++5dgIumq/A/PAfUm+ya8A+prQ
S9z89DstefYZExzufC7+NqI2lwkq00rvt90eOQaBaHF1dGYSLtJxgaEHdXKsuQsY
qzM5a/ukZcv/WE7z3uXv+wPeuLDd8pv+p0lKwareFBAqnmI/kQZ0Nzc3nqNjB5dN
ugBcwHx+BI4QYuHYzy6laSucVES8oeCgfkrg/KuPh8amjsp0hwfSTFexpsv2g254
kSrnImb/hjm3EGxvBAiPmB3x3lQdBxNY1V8eHW9VfGMM2rx3rjvBYEP08CgA8umP
ynjkCTymjncYClvICAt8GV4erA+KQclPWGRJHzNgbBvJ/icLyzk3bulMsI7dek6z
72nXxcHwIasIf8PrfGQzodBE5JROmp/MRDvl299mMi3ReGxGAAcQHlCpAtsl7hJC
wFgIxxpKapKsLbmDlWrJ7svZ+RMl6+KoJuNT3jHypOuuhfAIgtNbhYuZvjjdd7tb
aNf3V1ThSfrZCTsoovjrbpaWfqBRz2xg0oWEk3BpiRhSWk71+9tSM4/gUyK5WYao
/lalU+tHCuu806n4z/ArK75QGJhPPuKBFdW/3gL4bIjfIjsfIcR3YWn9oA9Zjpkc
958CBZoN8fEgIh0Kp9yBXuXi8gdtbPxRW5+JXNkB1JKbppDqeiuTVMBgDmAN6j5A
2DCel0HMinD1ZpDQzu54pi30EVHuUHD1Kc0axAEIQbcY7exQyOirmqnypimikyXE
YhIhBBK/+phaZ8QplxIp8YHWKPDX7nuDkXcCu0iv3pywQCDi/lRz+xTSwgisunbD
afOEXZIw1O8e4y8DTrGsxDTGsCiF6xDIhPIWglZvSQssB+XpB/NunfGdDWfXCdkE
t49p9IFcnQM51w7KQrC332QgpMhKrYG6a0s1tdXzTNy9qzbm4NJvRd39Lz+g8JmY
HPoiq6sjStt0nIu44G6PZjnYouGKCY7ybkEo30T960CmJjcjM7nXZzHkuiCM6Pji
9BXzKht/vJtLtIRSumlZKfy4YoWCqnRM80K4s3dXIf4p9sIB9xhso7Zkyzxv79FV
Uz7LF20Yg13Ebx9JKEAlCOzaHnkcN1t6ndiTkdEtulLoA8SNAJ3XvljPONvbHRMB
PzRWPkktZC6+OBPyr0a85Evzsjyaf9LMOy9NTsVcdaiIMiLMDw6M9l0Rkpgcrh9q
Fi/ETC78t0/TexDsf7CxBG5THV20fcr5m+AZgpDBQ0Xsr25vaK4abgBaYuU6yTKX
ek60H5I09FuoyIlW3u1CqD20bcPNii9UTAQzBY3Q/XJyubQjDwPf56Vr6iva+hzj
3BbYzIy4r3vlp9fbuntskAS9d7U2iTpcLXV/K4dma8pOREXH0KqUi/UJQgP8IFkE
KATX1KDpoosGVSkxauLIJxO5nL//h8W0NbEF6dA3xjwFc8EfXPouLQ1YipbajQsp
OjgmSVkxSEzfCOmdzRKUlSjxED9tWHJzeUNA5/JijCMeRUWqMvUPAUwfqhb1lSnM
R02rd/PLjibJTcWuize3gN4zG3iKlfDHDyQWMIvTuM8PCDvYzfGsBelDinTdPL42
6YwtzFerOHGNQHPBVdlbfA==
`protect END_PROTECTED
