`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sk1zcjnZqYBJPuwjNsu9Dns7IYvD+UYPJ/DYLsTbyPZOyoeGEStVQOQa8iIs07aF
Gi7tci1dWfVtkIZpKLBKWoCr4uo7+/FnpeAn1WjRRfqFrVCAejux3nVWkNRJpqQi
T8tJqzAB/aDTmxmL+f+XJffH2Z5Oi8e5jcR+K4MpgbyqIKriaQIvJ5c2McD0lnMP
80A3gErYhii7HewNnQFmqFaDQo+RJDFB8OH20v4bBpeaqvbqkndVKwnZz7OQ6u5d
uKFJEk4M5sA7g8JnfN7ldXaAKkd3i60L/XAXz2yNZrJMETsPFipHEE5X40k2ZYep
bi4uxdZcyxh0nj5jDFZzSDTohDCOPLXPmgAoU6+qsaFX9MDd7PhWuvdR1DmUOl6W
MYMdXCPVyp7j5QNC/aJGS/8UiNdNOrhFi+WWKTiP1st79LalFaLpwoqZT1Qo5JnT
n4SwD19F2abRd2xyIPADB+hwGVFdScnU5+H7Riw59YZyCyh+NuFU4870gUS/FvVR
KLk9eX6CJjyGfPKxjTNRRXI+ZgGCrrToMV9+55BUkd1uixnHj28bcyw9fGutNgnz
KxJcTyGjGQnuXfMvtyVYODmtFketCd460Gk6CBn7ZbV+8gZw9eogjWJwtxD+ijYz
ybtA3WswPKh3y1rDAAi/i2V64cleUkrXz5m8YHls0S1MRyLbrq5quurfQ852QXt+
WIw7FJvxZr1thn6rMDKMZtb3/3XNuAfAlwsOP8Hko5+ynnxk6QZLwCpZ3HWbsKkq
cfJuGolo+9xGtUIittjOoO9no5KM1jqL+6TECPpEH3YsL2CIDbnLbOiTZBGxgJ+Y
wUSvojVmn+ZpFJc4VB4E9yA22SMnK+GnnEz9AaDsYnaM4eSA8z/dY+9+yutjDlwy
bTXz2EQlrdmug2NfKZhe3GBarTV0WLT+TyJih8dWMnebiE777UBr7b7BXRqwVBQG
aD/NapUMjR5pIS2b80gP0PJvhANVeYQiVmGYVwoVvhR+5ARQgWk6As3zh/HeT5pz
S+X9pesUD2VsSRaOef/weVKojYwzviVVV2FVDBSHSH7pwaikqkeWhBBdiaDBqkV5
Nm3QLGztFvaNlwqtHKdA+s0VqpVin1RSMgmqHPBsEcyNOKsZhSBnu3Sc0yAaLa4I
lofTip1ns5M/AwK+B0Ajf0zF7o0opq4tCUIUBFugxScIzhSkWMxX1wxkw6dQ2Egw
`protect END_PROTECTED
