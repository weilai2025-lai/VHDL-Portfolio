`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kE8CCnTF3jcmFZUfMaLwNJvTK9TEdkusQ3Crq5bbp0bjcBf4yCuZSjkDqohcxenM
LJ53ycp3j9xKnvaUpUQQjHmtIXhNNdy5DLU1i528xxJJ5RlvYBv+2MFlZ2SywGaE
LdUTPfsak2V6/XFDTey3IvnpMOGv2cxwGFOrC4Pn0GEoUpqQfK/FlhxLpl9FVyAs
+FPhUPIJAjfLH9gAcdWEw8QPnRPe/Mbl2Bi6N0OA7DqeofFrU5MpmoOY1gA46FBg
gksTvHz+gx/9hDn7FsRzMxkBKvsmJ8B5J6PH0K8lQq8g3WSJepmdT3O+tQY1/J3V
BWzddVMnCFcOWBNbSk7c07Qm4biqKb43Maeq9ntXC8cFXAtXZX/f9idNaK5X3ApA
k2yqhzHoJzSqi98Pb3v9qYoLoXTBgy4+DrBSxF1cRZhs33Ea/0mdobxkE2FcRdN6
QydGMrVSwJcz0yW1Hor4hyKre9Tw+Om8jhYb9LpR9+RKx43XS4zmSRdY1pDCfFVI
3J2St/F6EPJHbnQxi1C7Xp6MPMxmMCE3PeDCFxus1C9zpyOvwqRp+6M5GDqqhQbe
flF5wD1cuRm79BLhFHqyUYWmUusBzp1cAlJ138WGoulpGU/JPtA+FkqWkeg50TOR
q4FAYKFbbfKG+Loebmc2eyj76I2623LNq8aiCdUU81iqDcm7h+++QeiVUoAYPEu2
tiHE9kZ6XFcyjD9wVoyRKxtssEpPbMslJMU5a7P98Vk0cd3hbmsSt4J9RQ/HYhtB
3/hdrVIdErH3tVahaj62RQEnYcZ+HXzOVY9ljHhr5bHr/3AHtGahAbGm6x+RzTVY
xzA+3cZb821DTRt/H7kKQXyqC60GebUSy485EgvxXqUXAN4KynSgZzsXmSMbmhlM
+8+ElfdmE6cWjMAMNVBQFygWbnbdgExVHUyuujT6Txr7JP7VYFM6cCYS5gpd/zy2
R1RCfN/rGSJPRmAtCu+2I6G1tPBzQbCtkV2COQfV7RpLhAozSdcZE5SFs7g6WN/6
RlRkWyYO4cAyvfgcfm2v9OdlubqrPLD60r3xL96ojIAGZ1/3+IqBQExno6eCSN5h
pT+MdDS6L5nVm18LZ8HUESenocLNVGEOJOMzuZxL/Wk0gZYtY54hUnAycRgMCYYM
y0TmAWTpRAuymHpxGvEQGF2wrj9vbinc1J3SU24txVNzLNXWyZs3QzNoUv2dInSF
EY6zAEpZsIAeirNcmg82aNNBuWzsyxZ0fqXmFwUFnKtGlibJiN2jadBqYasDFw/s
0HswBpBEM12tw0LsdEqePZloQc5Sa/Hti6xT7IZBc9FwBy2ZcG13fui+E2HzNnUB
qQ4vjut+ENQug5SzhPNvWuveaP4KBrdYWDYagHPbHj5HBmxrHoSmXciXgMGgUBxz
bBdBjge/bLASp0j6jdcZQK+G4HR0OfpIsbtVtFWqmfDQo37HjdU/x0X7amgJXs9Z
n0clC5tXa/wyN18Ty6ABT1qVhkZiwUkNrIRi8IWZQxyjA5ATqzilnCilLnUjxO2r
+pJNp2tzWtkjhOfhR6Ax1gNPPO9G/RPVNNCWt2lTtg7ptZUKq+m/H0hF7bgrdYJY
5Mc2b1PU8u5A3ZKem4GB6B6jBNNuQe8T2IEzSrZK8kEPqDw/ObNpz9NvnJxSPtQV
9nJpt1VKT/2C20hyF37dU1hN8+d7Xjl/JnVzDkmDNRyV11SGVDbcvLZNVkxutd8c
c9pCSnnjSrCeH42njrgXOYhPTTj8si9CsnnPiOcFnPGhe1Klu1vBN7H5CDVPueeS
RfWHdDv4p8rZhXvysXMHAjH4g0Oz1Nm+jaZtySpi5ZKqyJclnGUj4ePaYjr0ORPT
85rW7XGx5veI11fx7v237nhQl10y8RjSU5Hq8Azf/8Q0/7KbOAHPtT/OBSHbxRXW
EePA697IpNn+uw27RRz1Ag==
`protect END_PROTECTED
