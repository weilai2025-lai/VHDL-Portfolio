`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LVH7MHlbOzXUqpe0vWfqgXifRhG1BCPCacJADpdqIV5ySOGpQbATlwM22Aimu+ps
n28ERomOlUuPS00NuL/sPM7SRYl1sMuS1dCl5qPB34KZHh4hPeedq+gFaXFqPZWU
8QTCbw6+EG9Tmm/FzJhUs/t4KrqiJthH+3sljbW/AR3yIHAZa16FsuFoyGPqAXlp
DoCknFEK1ydxygnf3h1K407/ZH90f3KGw31lp7RhUf0HCo3CfL2iKGI6r5bn71AD
f2X3uhpy1disOCthMacSQSahjxTD+ULxezEGov/nJEIebLDdA4k09WO29rlYMqJN
guVx2fFoe6vepsheSsStzfU4kkYq9Z8rWK55kTXAFWjxhojpQumtydl75Qe2ym62
An7qQLSEx/CfzFDOBtwH5Hl2xLYu0qBPQ6/O1mEDEgiDxigZSymWyURkqXzjUafs
0e1DSgSBSkgmFIlFR8YCfq+BV+m7JpZ5O/R5Fb5bRe5Mn9h7so4qHyH6ey9fFdzu
yyl2estAUWmDfC+3rPBIgfXMkD8b5MBgFtbTeamG8BGPYG8awwbYDzJmkQ7X9Bpf
YUSUc31VQX//x7n/nTPO+mBDZOSb9ZwB3ZwJXI5p/EzccXP6cxD5IUN0cAqtuvZ3
yr2M2EDegtBhswsoayKo9/MLW/sf3tsDNcV3fupqu47oUJX/3R2f4iwcFqAMfHTK
QzFYl+VlfG7ihMf4ePxGSivHlChW3SFUHE97LvBTsh46EJrBufbYNM9BcMfrjP2g
b0VBj+6QzdIgHt+iWbiaRtetuMybijmY21BadI4YgsveyiwHMchu69ceOJOdk7Xm
fFXVBRFz9MKFwH9rU2YhPcTesWq2/9KIC1hSUk9XiPc=
`protect END_PROTECTED
