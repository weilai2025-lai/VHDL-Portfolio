`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7KSyh7D1SOrQiMvhJZJJY44hSAcxF3PvjUKIiebBglwSI83rIOEJUz12smDDwlar
Km/R5HVsL0ANppXSnf7wjEqsCkS7y7yDOTX5+XpuQqzGkI5NrZfJ66nnOM7NHCsV
34XkT0Si/nGtRLj1YW5b5GHZuK/qy39oCxbJQQCTc4pDz5+MzYArz24FsimZht3E
boYuJsYyU+S1sYGeyWABhuzXSLThIrgseFNuzQJ+FC8FRX4KXhIBTf2qYhDil5QC
L+0EG+OQXs6lAUYYPgC9XtBVzSGFbGbFpuB16+a6ddFUrLyMkTs5237J4ep4Hqr9
CfD/MQCujROMD3WGPPbZBCC2NJGU+feUPKuNzseZ9HH6ZaGbH+OajMpqo/UU79AF
6/APVsFz/aEKniUyLr4m/b/GF/2MY9m+s1kBVhcySnxzfrpabuCrPxRNBIPQPj+W
wTUPSkdrSm6VpbU4HC34gRMpiTVstXxFEGxXQjHra7RA4R9NHNROABxmUgIYScGT
jixePqkTTPe6TmZmyKx/rtnNC9lzJOvYQiTfmheMowuFEP8nVn/nalrNPwdGRxb/
bpcN39IRyiTDtlXSVZz6EH0rY+VaE4pS3oXerz6x+fxG9r8i1eqIPLCu+GksHuK4
yWZHSCVwl/WCAhP/sxNCOq1ucjS3UMCiTrkrMXmlyqRfXQp7hsM6Klb+H35Qvg/C
HjE9tt42jorXflOrXxQxUChRnZ559YpP/nZtOD95xWyv68QeVnmK7g7UiyypXtiJ
9GQmAHCCMZGMwTF3VXGEN1zRDyHKQWcC+4rZL0iDmGSnzYr3B5xtJeIKdHx3e9p1
4z8t9gsLCJCtyq04aR0s9ajRRMMTclmgDHd3uZsXt2bqN5Hbhmu5zj3lHxz4WM7T
1ljRT9DIAhAKwBlJ5/feSY4jnpTUsK2ygeGGh9kC27oEWUm6f/+TAXLFDNN6L5GO
AWMawTHHfno32UC+4BVoy9wa4VzwREYeV0a7j5NM3V5tAedAdOpLu/ZY0WcawMZL
9dyghpsJdsZHHjiJHsSjihDX/Ckz12QX4MaTKonxjkwXI5myuz2r2aDbFNIYOe3K
LvELX1we3ISZ4HvOvHqxLv1xecz7I6OtY/3aiS45XJniJivUtH9CjHhZM+U1NWfW
zZHXMrPthLZzMLzXuZKdwApQVA7si4zbOZZxGuaj8DMr0lhcYqHGgRGwWpTLztij
PHWai/MTe40XCWCLMK63myfu829DNZhoQz/I7lt2j0VfDxfTV01O/G8w+S8dJqBr
cAz2/WCq45vQUWh59tD1D8yAbkL8En+MI6p02e7slhqrUro1lnX4nJMO7bGTMfMp
HD5c3VAndBCIRkifzWbBTLTb9sv0GqIUY8ctv5qOs1t+NrG672pe1OiSK3D+Y5EL
5jiwDekFOYSkoIVDPi4a0M2+3Joel4i+nQTzYd7nEZALscsekkgJzGuRUMXxIo5c
Dj+CVy9tszS41mwoNovbmQNQ9yD1u2jPw8dByv0SmmRaTkonfA2ueCkg6XFv0Yck
GiV5uSy33S0sHgYH+jJlJwzCiPznJJ5lSY3TBLQkPu1O6g6NJI6SalZdj3CizBWz
kp9/Y3YL8ZoMJHywTMsP8IZDk/JtZGGG79AZUjm4U6JI0hdnM66tBDC9Iah/2alR
4mYSWY5Z1OBZQlGXph8PjtAiZzxrODmWBuc0lIC/Y3xMZQojgm4YEFXEMi7vvoGX
bPRZcSafGqggpq2MfH1h6Kn6P6MwTmg2YBoeYux/RgkAt4A+QaPR94L6b4m9hMnn
scol7jHeMIPWsNdkLrdEvSP8Ta6f463iwobwXt+Kqeb8Ix8hqtM1AH1PAhmUDf1T
cBT+HLJLOZ2US5xl/JJ/BPQPey/TFfjLM/2Kz4Kn/hWGGByO2EG2ORnMm6C7jwLU
LaOtJEJsMIaeU0uc392KTVtioL5o/9US7+qbEGZXKbafs6+4KTZtpR4L5nfooOwA
IrMIJN7P+5OEDqMOlwxWoeiJ4pjc1JBEcI3jA6JAtrkqyzl6gXT6wVXQH9H0pLV8
qhsLhj6xde+++GZshi/ZfK5Dv1WdPJjWR2KSmswfYQSJHA3Jt5/L3JN4RPe+98LO
A6LRidTRH6IWm9j8wuSiHr0mm01x9pUpGBLZGRcaeoAeG5kR2Glk+R6lEZPhzaIB
eXS0k/qp7pA+t1jZs+uML3P3wJyft5WCV6VOeRWSbtXphw0EOqxr2FwOIVsDslUP
1HQD/u0MMVIerpQmaixW8nx31FHoJQdTiaitIvWss9hoLVQMTtK/cgHDB87r/AZa
/91XzSXT9jc6deedQbxJO6vQX/+LlOMn2ppIdkuq3BQgKVjEYIlkTZhLxBxZcgDl
oeq95YGfl9gRaNF3Th8IeZZDQFUdKm89AsyaEZTd+vDQ84jgMcPUdaOhx3+VjWvV
0ZvkGGCT5GyaRCU5UfQgnCfA3+8mV/U6+XZEM22dzEOLjLS/MJohvwvrcwvLiN6F
GujUPvbTjJcc+6Scox3ZR9ixLP0OJEPoUzhLf6yf3MAmxGXuEDeA7n2D4bUYccVk
u+2m46OFMS0Z2u++ML5Xe3D0NKp8wean42v95XsJBM19GpOTpY8PlFb2J47orhGk
LcXoYgsQbCrLJHlcFaU/FoRWOnQYeHy0rZAmazCDOsqzscbpH/DyVVeImZmNTbSM
i/aU4mzYQwrFt+ghgWfpx/EkEuEKlq45ok6yoCGK7VYvHlKI7lo/o9QBfSb+13A1
lDiHE2REq9hwBDVzkPr9Xm3VtfQ/tj6r/as5+0t9fNeI+u6OLk7Nxc/SsBnVhpig
M47nXeta+BXIbYrHLcQhlxQjzxdHOpM1G3cgBbWyVGDMTNkBYZ7X2JH2rHCG+1AB
Aj+Iu8MScIkBckI3OQt3exShtmaX5SAQ2corMmgE/z3BYBkmzj5zOHXJWguh/Wj8
W9oPGDzPilnMYpplOJ5hTxci3qMnXjWaHO2ip/kx1AEHUAkWACV70cL6LZ51CkPC
a+dn6A2AXt9ul+iV3cFw5OeLZJosXKAHx87LV7zOx0RwZNJCj8otn6j0ns7py4Qi
Perf1P61gkNRm5jR3Un6v2s468mY603JDWlh5wWiHOJNoSm69OhRO4lXlA/H1R97
+HkrMSTPnnA04rQm6VH25sCIi7bAdZUzZqAItDvJ3TE9H9rk73oNbfThmelqjdBB
v2pm5T/o/iWaCIC7DOgzu1VAtg1fyzQAxC9OlSys/fDSdkn1gWO6VW9JrOApxqu2
2KPFvjRhPW9e2tF1avltZ5l19r3b0SbM02SDLaH25n+/pJ70UOxY74CUAlLHl42V
pi5kZLnWNxCpRv9fOAi/TS/o4eHvPBl6ZTnRyJp8+A9Jf/zU2NlfZdcrbbxBhTiK
OchrPeLwwP883JQdajm9cZm780/+AVd++NiHEUXoUmKa2Xf/J/quRMTgNZaFknIN
lQ1az1KPAJEUVovW1dHryN7bMWUC/OuxPRZBxa3y4+Gw48idVyPAgWoNKy6qlefp
4GKMJF2Mm7z+01btWUHkHysHOjJ9+vbaomHF+E0f0aLuO7jw1fhwUEiPZPTKbwca
/bSWy0xJje/mhlJnQjI+zYt4oPdZPhTEwu874yfIL2riUoGjbc07bO37FHVb6Fpc
ZZPNR2UVeKVsfHAyV22Pvkma9t84u5tHiO+a2m+0GuaSrcAiERJBZOC0RDegPDMV
zztehtovWIZBvTxbG77DN1H2H6Ma2d/F9OTQ7kU/14TgE9zitn0OsdiYFXUh5mBl
x6CxtOKHa2Z9D6InGYrkT5ILXw9jEFYP4IBrf0S7Kb8vUAxZf9jxX1nd++AKUH3g
aHuG4etb3tYD+TRybP0880s8/uhsx/CJkN60UXY1gFyUaZwAaqxZoU45tkHr/GTB
LpUeeymtaTLhnLQ8PSESq0z8WmV3XgbzAmR657ZqEk4BvWcor9GKI+8WqLsuZufw
e/JAUlMrmftd7p/XstB87ojAinT61Qym8NqpYNteDPzwbQOdkhlwSx/xH+remfil
5EgyoFF/DCnQIkQiwD+4LzOHzUWsVzhIWCPDcN53DmK3UHCcwFurI1NBykjW0pJk
g1nDvzDb1smjidvDLQh3/b6FQjc/9nXBtukd4PEH8g+pigEH4Ce6/8jKe6HsI1qW
fdnw2oaUYDtp3xT496XeFIQmozXy6090NwjpGRhu1S5mA0/ySW4s41divi/g7NCF
0JUj89g1VlawNlUxrr1HCxAMcg2Q7Vwprhzrb4VdQb/csT3jxaBDKjtN920uNasR
y6tRwevm1Puhl19fiT1EH9U9yq03vSSDmVGnY47oeAnpEERx9ReAfJhvVahDqZbl
nDEE8KUWhyamCwFUVnynVafyYZzYKCHDfzWM6dWN0qFSB8LsBeyk1uqcW8aocpPB
MQVvH5j/o4yRp11oqZfLqwaWi00KDfvnWSFUJ+DlqbiuaVhPNz7bfcQoguMuUJKI
YPXvVYxsMFhXdejChH2eYP5D2yhWDrgWTPVK8lTO8o1HyLWTe/dh7zb7sQ7C08uc
Fbr3/aGk+yw/xqKcIl6jrjS5pDINAtt8NXZpO3a5pR0fxkHdjtlgh/0amJcJ/PDp
`protect END_PROTECTED
