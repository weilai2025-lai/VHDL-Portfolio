`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ftcdSSmhuko8Q3TWRm00va3n5QVD/bLNmQKofy7n25BqBVVeGuNPeLE+5K1auj7
QtYXkRQI4WQamZ8NOHkFwIA5s3LdKMN8YNLVcwyf2TdloBOc04gOfrbhQcpMVEYg
5aFPPm/XxZpI7e1hdwAK8gf9IWHWXKEyLcG0/QBIbb8Zb2Dx5v4wWlzTxN7Pfgl1
aWob4WiFhGU5yuoEnfVvv1RreqU1MZ760kBUgAQyzSxbDhO2sJdKhtauki79RBd8
yEd0wqSG29ZjTW0Jzx1UUylltTB+48V653WCP96UsYeBPvpJBv+B1E6wYCxyEwCQ
UXA6+S1enDXeCUu8zvj8OTxwmu1n9hmTuR7GbEVZMNZ9L7+dfhdOoYmazJZuQXq9
c6Ls3zmL4zH3W+v4InS+EEAw+UYotC3cvPWMTYgmFE8x26yUvvcy2JCq2CKfdR6f
3b62vCA/MYj+iPQQvU/tvRSP8RyXWAFjhc4MzaWLaqs=
`protect END_PROTECTED
