`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EyybSCBs8Qr5qRg+ue4IjaMYYgHK4P/b2sVupUyTpT5xr0RmdaIjnwVDH7Z5XGTE
sMsKVhUd1ktsAqjvRV6QIMwG1VTGUo9JvSqhQjUGU5tdO/mADw9C99ucAsTFJ14D
7KY27MAjXyoXymONUAksvxsRdLAi7FJey37puts2pv9mMFC9ESWu+pWt1PXalQVs
2nDgLMfu0xy8dsR/XRk0yhWs9uAtYLmx4SLyvstmr6RdBHX+h4SDOPzCHJurcq0n
3th18fFEOT//8oDNxHs/plIP37aWyP//27BCpX9LxoWag5yg2freGa396DfJp6QI
Ysc/IZHViJMkLYqLBwdHkhMsFJ3VThiErdGUbZweFb8VwrLO6hA+cbLiuXXLnG4M
`protect END_PROTECTED
