`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lx5cQ+xvGVxmJ2aJ6ubRPj8xsO6PGjfGtnsmPOKBOWRV1cxukHJhSbJVo2+T5aA
SSw/8RfZHTqWq9rMLnb1luG9JYGFzVoITnPaWgesFOVm7nheICYary9yWyuA/R9s
OSrRYHaocWxDOrDR/q0+uhzzYcv9gvo34NfSVZo2xMQTwYSHS18/4gPj0afuU5oZ
zXGT5eyfFEAvQBmNNIQ37NczX/DyJ1550HNUBgTGBuqmSNzumaG8uWGF3Kz+cy7Y
NAbNez1BfJSb2v0xfkDVCtRRRw36NdTF3wiTUPR0X6einQ5OmQH+jicwr8/xxx36
ptnNXUwp1LeEHytH+v+ANFzKsalDD2rYTKtY3LUdie4tz0D9QEIHFBnMLili1fRk
5n5mUxWcBwdWutdeWXHWGoLhoKyAMN6bcne+e1nmGBhZDzT/61chiH8OHrR+1BCB
3Q5/EBAYHch9cJ1i9IAAL+yNvyYIKAGVih1Nxp3vYqJiqutMAtA4j1Tdakbwy7wP
tBLEa5TKaqwAhBMt+3WpAyA9/eFynToV+4Lz2VPsARy41p5uOZVUCdpsvfwjt4aT
s+jh3NCnZc9Voo53ZHqafYnG8WUcREKl+bK7ecGyPojiJ/NBSwqOdBEQG0czfKy1
o77qb9olIvIDa7fuafj2j7clz9kJpvaGF5R5/khH2GsH6DSchbEQsNtszGgJCOBd
tScLV93G6M35h6AV0HINiFW7VNe6hfqEqhX6Z4X8e4UpZxpyG3aktnjW9IiMSswC
3rOi6Nnr9yxRPgHNjIHTPMrECODFkHfrMwHkxJuOYdGrbwvQUNYV8XEHERPoRb6Y
7dl9V4ab6Fnm6QuLBTBU70ZaLWwLXiVxfLdQe/hciUhtjRns5AJeAQ/V6MBdm1Ac
2beIPGTTpRltIOLnt1DKqv37fAqm1FPb7aCDgZpAtJiq8G7y/hgj2uSftlNFzQZL
aer6YMfriVvETA3DkPU3/+VwuECFWzR4do+NFkba3u86RlzMtKFLJa18nKSPwGly
/z4wayLw73zHIDWYsfLjSWaNAWq1P9Un5iH1QU9rmM/wKJo5Yo35nU4d+PdE6bbH
HKTGu8rKWTY4biPYSafaXhf6W+fJ2XGrVtBuULPRe+8tzxhbiXtEC5cD6AKWgE7O
lqqIntrSfBe/cPKIcbfrkenTBzgUkdYA3guCp1xBgtjaO8SfAOyU1sLBKCT/isZR
tk24b+HgfBlMrz+e4HXLvdp7m3xs8cZ6KuEXwXbnoD9NFoyN7rOPyS6UO0wGUExB
Hq55MOi+diRLwWGDgduXR2rpxcTx3xEh3GmnL73iIiZkYdUZNg8cJguMHgeVfcLM
SIfbW7S+9grrx2xiOX0l+FBuZcnvN1Y4bwAPJSRGsUGGU/DxmxP+JuaOs9qH5RiK
IypiE+t+95h/13WUiTfKnIZ3VtsEpMbdQDxKExrUJzVEApWSY86/eONl0d2zd16A
AfzeQj3WWPyy6P3W83sJjFio7CfsiFvhpQtUcgxuV/HnhHv9aTEdV6wEBNfJy23r
hHjqMbrKeZ9lNba0y6l0WBm0ZUWUjrCoENeqAjtCSHd/mtoLoPSaPAunC5gMMFa/
H52PKISSwsCT4bD11RhVBDtCTpSlG51TnRIFAVDtSCLVPtw/Wl/ar3BwKCaydMjy
JrRMZxyxEHOVIldDB7Lg8kDtOFuCxOqM/dHobiVjT6hT3eS4JuBrt7f4R0ysJVmC
9jIYgs2xEW7GampYCNUspE1hgZ+Q7mCCV7EbBilAu9MlY52ElaDs67zjvJZyyxU3
4Uy6Xax/CgN+TeDqIKuhL/4jNDdHX4CiPl+YXzE3Lv0iBWVHFY26fZSdJ2W8bmSF
2tK398qZSJ4O4PnFdPFOXOb3vSHOnP+KgvNwUUtnt8UW8okjtz1BkhApkriMc7Ga
BGn6PPznxENVJDzxPypx9Q==
`protect END_PROTECTED
