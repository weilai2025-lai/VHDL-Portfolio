`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2NMRgf+lVXsHN7NXB1UCCDvtM1Od1Qo5eFtLBdXi7MNQO4c6V2YijiJvdHUsl8kB
7PRCe6ab8EJWc03v7FYyOwtPeZzKxUrhXS641PErqd4uKklZ/0nJlYbB25VyyKqO
sJc4Pd2ValwuYlZsfBMdAqUmX66KINlLN9/n6QVvOOjXMDggnP3phpMr/zogbSuf
hv/Y93H874CWIFg80iW1YS5O1bGlcMqnQXFuh0VCM3zpXpqWUuTCKEuzHXieSeUK
GCKXgCjPxSJROgA3gSWxOARXA98zxq6LPTRzeGk7uVSUn12jKVj6VKdc1IjGlsDX
xTBpDHeVtmR6hi2d/RIz3kJTJYIR/tYYB+ugJu/OMaSt3BaII5LVIPYVZ1Ss9QmV
m8Y7miDoIbou1ofd2Z0tCBzfYJOvG5bDqKGJ5N4R/U5VYEQKAXCMzOKJdVei/L+L
SQc3neXI+X5tW4fJUiX6FHmsxmoJOmr0MPyadqU5Umm+0SjppvcYzFtgsSsiAV3B
OmoIdX+2xx47G/NdhTcOituFNhCppV+QmVLYjFkAEaOjJNbbOvoZjxWZaIqKmnQL
tMKCWZX7//Fpr4tYMqzyLUR8srFQ4aFfK/0I3YiNTQ7u8Z/JTJyaqxsxVHAu6z5V
VCnyzuRRPqxR3kdT4FgUnMdlNP7bWzPUEZqVLFJmKml3ZfCWD/q9/vekHat5Mmtg
kX9H0MNw4KCRhlVFXMkDXKeKySMus+bInOVvIdpJtBOHksZEbfUwJEDelrqol5Rz
KYWsyhMo7xWHnHoueMb4+ZsPuwV3MVxPk1GwsbXUd2SmxwWeuElfdEQElwM43JSj
e/i6kKjHCFEyz+tsheJ2Z3ltdR1WWGaxvyXHmOmSmRI001YbBZ0hleFushwBvN33
G2/5MPZLAzSs0MK0nrHIY7UXnmDR+jBZAjV3jwqMz9SqKwFDuJWNslOaVUuVrLCT
zNo4f4AP+ddZH8AXZraMbcdb1AQbwh5X9lDyFi111lD386+9PoBH18lNJ7xpttLl
joDrIWXu/piKUSkY5OceB56tbjyzg7EDICJGOiUDsuusbsgLBvi5UVOPBn3Ul3/9
DOmQ+wSicrsx2xhXR9xbpzOr9POY3sfqT0dh58IT3eWSEKrhlpVVszNnrAD7Iudn
tCWMrMQImxEhCu9KC4y/rYcYA4ZPZgHZaNv0ZFHRFidGe5FlPYe9hQLdix5BqY6U
15YuvkTAcbSNS+MiLRiDg+K2tvayBZF/gK2Md06y1myTEm+/WRohchL5x4zmA9/s
gsJPHkrHVEhLG7/oDrZdyHcEjmruiVA+6jpyEsRn7347s5A6klbgnTpZxJZ5M7IP
9Pjo+Fmw8JAi0wV8YKn+/w7gBYvSvPY9RWPzrAzPSULszyVkwkf1uKcns1NJ7n+W
i+oXTweaH04oer+9szOeqB8bMvakaSWpRSQJm3b56NfB1UMKMoKAQkvy0KCKrxh8
kdmKt5MwEt0GSUQ2JbRuuaV1Pn3F/FWigFY41htGMU2D/d/n53w59raE0bAzkxX7
ThEyQtMh7JoNIIToe+0P+WkiaTVogt1LbNb53wHDbOSOWZf0IEJ/leYuTmJlfDZX
jaH+WLPEigNXq/K+od4wR5jxb9b8ktCQpEi+Bzyg6rhferug5mSOp0U+5fdhGX6H
NiBYSGFnEy2TcW3Qv6C8S7Y1qMhELwZARVTnLIzOwGcXAEzvnwrT++zOA0yFHlBv
9PWA21TMStwCO6XIvKtPi5ORhyQO/hA/OsbYmOVh5rAOp8GFUJ8Kd2BDOo2P750n
7YBFG/WRkUN2m4H8nX58H/2Ju3GOMEmzVHdmxSH1CNKBybv9Jl/3v072UopopU3v
VYGnCJjbeqmk2hQz4c/F8gt9sEQa3I/05pJnDZs7YBzZ1NAAMdNSbjKGVhJqlyEk
KC+66oOioL1/tleAvUHEOEeVgvMYDihBqeTJW/Xms8CDp5brmenev2JBUMV2x4Ki
CBQg7kOEYmMhyZOBXwZKoM/M5QAav4uoH+VwiJ/3f2P6q7t8SuKSnzQBCVyrN2aS
ceNxJfbvgYGGS0AV2of0HRsvHrvFePwecQwJiF8Ep2sYcSozDLDwF0R0T+ouPgur
mWRSSFS3MdWRO+nMcKxoO5Hb+Vd4JwbAD2U5Mgjyh0GP8R54ilApdQiwqw37AH4z
9SwtsZnfZMVaPOkNQyhYizCb1Eh1piy1CtQGvcPZutEX+UH6kGROyk5nL2FiNk8F
hDtQD+1N4salUw7nnuRlhmJ5zAu5teP6j6qkvNUwmWi0fiqIdFJ2YfvM9DZjf9hK
hDa7SbWxsi6d77OaI+ikFgMpR35xkvELpWKkswM3gKRBdVTOYqa+4BwGLVMQ7pFy
kV6/FVpSzUlO2otKwTzdWazyY0pLH1XAMiqipe9zdAgoOto3wsVz14lN5Xt0GkGO
QFJTKu7X4Yxws5mgcJqWSWc59wJwSiFgcTu5GrevUSRM4Lw6fM/LLxsTt9AgtaTg
oVSnZxLc1f3SD8IaVMLFFes9pzLR4RECYrfEf9aeiNqsneqTG9IajY9WdzxwNwsH
2xEWZ6RVZGGnLxexhLjKVPVuKzbzlXYFj8uc2Divk8W9ugBBRGaK8K0MEl327XQ0
sc2AFEaoqIviQiabisC6PW6mKibwsp54j7V8JzlOyUGxG4eqD1bCq+NyP04GSZY/
raD05trcbw76x5mSAru0Cr6t7RD69E39FbVL3lTKJ66F2T6wVhhnNCV0+y2WsS1M
0cjIjF3a1vcM6I+SK4pRsk80nRy25IYwqofPaPpw2bSERoGrwUw8tavRU4vQV3wf
MjwCK2ZxRiWXBKLaFVt9fBEzSjwQdSzukH6geqNew8gVma2JLmf9zVHFG28ATouT
eFLeyNPS73Fm6wGFjwFdosflw7voPN0U6qM3vITtVBeLQc76mMs/lEdql7BsbRri
8APwXD5zeTAPVTuPj8yssjzzMijJkidi3p9qKocPA+y6GJC3+VuZX4m8JRqiDUak
Kf7pmzlfyCNLSkcZQTQFlFgiD4EESW9VrbqEEapXNIa7gVzHcSvkwVoIpZpFqdZZ
y1YALvTTcER+AYhNnlFM/W/Z4Y+dDyZtRbJDwHJ7FGJvvfXG2QdNs2546xuFmAmj
tY+U3sVJAevQrbbfaAHJLNXa8OdY86/lL7ug9ya2srgJ3shlZEcDKXQWAY9n1vvj
s6dR1cNQjV8GeeLl7mWRF9mbqSN/HaRfdlXGYcp3p8Q/9E0TlOiX4r9S0zlpcQ1l
GzAnvCLqVTZDfhIKUvlGXliBdoFfYggXtF7AjGaUw+b2uwuswi9SSRLTDfI9iQ2D
eOjGLo8mkTzglCAOjpz4vSWK5OEoqwvs6TPzAWxS154VDzzRBPsrOakurfmxnnsL
FP6LjM6Db3o172EpJGw1WqAgpTo/VE80KRLjIEoQqCNt0IcHDDUFHikhtUGi1lFw
u+B0pzyKhLMf6w18l0OF9HTXJgZ0GhErLfOtcqds7Op6cmcwxybWP1T9h8SdCq5i
17J704mzxrE/nK1LKK/kDb2yR9wNf5Vq0Tn2HaMAKUEHgcnhdeR0xWMNz6iaErW4
XQqQ2yZkh3sTJyfSAUhF/XSGhBk2MWGdTa/ZjYsfja0ciXpyZr3wMySFBZNEEbMy
s1PQOZ1CiPMwJ3TIyi78/P1ctxrtJa7B7dDdmzJxh5wOOUEjDa3sUYxFNuARjzWO
T1nvI8t2fH5DplM8LzaiKmrZX0tv5k/z2rqjBiuL7v4Jjdl190oeWuSBUgEsqTYo
yMl4z0q5PadWEOBUWJ2YxjWMYG6SNWvu5Zd2BBg31eEN3jEvLaqjb2td4Ipjpmfg
vcYyApsVf9xoyyzS1FHSnif7gFjAjWbVV6myk46ANaMQwx4BUH8MMt1GIHQgBUDY
oWH1AE/5P5QBGHby4Q78gJ1HgyqoKBZffAcN3Z4U9CxqcAVrocnfWlbpNKaaKCFb
hPGuQQ6tlLTOgWmYnF4gyb/HLe0OCVAMxUsiY1hZzOZgT6dmtbZk+bdQl13H45bf
M3XDfdXI4TiF8dafDl5uK5ccL2zQfCV5dhsfkjmYj+Y4BJPz2J9pE5FOS+Zgecm/
EoWf7ErLU15ODDdkMGWpPdlrEPGeFcWtKp9+/MXUbKCFighjw/hhiGc1rIvsEu9H
UoJW7t+h0XczyyCeNt2YHXBzwk+u0ukWy1csonw2w6V27wQxAV6DGIA5TsMtqQMf
0ESaJ2wBTHGeBW90XTPJsN+aPmddLVPUb/MPifIyYZHI7XzUNHLc3GMgoc2RngER
9iXSIXDKeET1ciXmt9ZeKVjTkviw44nTNZVO52bXCNL4i5vRhLeMzz6uCILhXhCf
gA+uraeRyD+A9oKvWM1dI+jQse71mLgtsHDewblUmIP7mF/jNEtYiaz2oiiCwy7i
GYJxFbanWg4zaaqjZxz3+c2ZpB1naGrOksxXQUQLXMSjiKCAnxaRRqL9orIPJqx/
S5ncm3/GYwPmpYAAAl45KfqhrjbHZlGeK6Mwtg5nBmpQ/o1GaQcNiqfSxrIEwviL
uWhkO3lsXqj9UTnbtz7WeLh41yx3AEtzLq3NVm9MvIetCHlvjGMUlpAlTIxfC7cg
Zf58nzmX3BuPwRyjFJiPcbmMlDnpIpgNrw+gcFLJGahGdnUQR8JX3hABBNkIedve
I1IqGFT6Y1UjYWSyRyF5wO6D29PwOxh0dBb1urxdKm3iySLkX8QJjXGmA3SVCese
LVNvoZ+6zhOkxJTsoLqegq0qFKVX1l1WrncBmjTZq5ElghOcB8EUefymoLwyaqAp
ITFdAwD9SbRM1GDk4zrereZtLQbusLmhYU9T11NeMrSOl0joG9Mr9fy0psuuSROI
sdTgHXyiqxmkxnqHINOScMt6ZOsmP3CjbzncbEE80UgQ2eQQhPR7QeHH+1zRvIcq
GHfnZ7nVDo7y+tooVcFxz4KHwYbWZuoQePQpaTZxDLN4ToQ/KjlcfChUjiD2veJj
A88XWpA8StWqZZ0PjJiIo7YSE7WbzS80lOUScqkvOmdarEBzWR0rkwvKMBtK1GdR
URrkW0supaL8Uq2wxgf2157woeuYMTcDU/x4AWWzg70pUlGk6opstSK5GRZpIb4O
JEZGmzQ8l+MCrvzkmioZKs9Uo8130H5OfIcNFk0DSVv2JyrDYJNYkuSnyxvyosQ/
F28dGOdffUj8D9Ye6TDEkh4akI1FaLG1RxZG6MpPzGU5L7ymop5gUHE8ltgQ0R+V
BYUEfN97r+jNUl3SIkxgP/Cn1+oi9c0U0KwnSaR+BrlQKJMY0I4oTCrBp28u9C38
nnDuQdtoYzURezugocQ09npwlaWhJFaJp3lSTJVvFWGCoH2sc80OQqiTmldZ9GJ3
IH9sfRWcEyHANnIo9Gx9M8/m3fqFY0KQxjGg6cR4Xoiz+fXJhkvly2K9JZnVbJmW
XVHZOSMArXomAec89BwQUYiX6EjEpuFtwTOp6AUISl+q9ueRejQiWC2QU3pVH7AF
z57HAtt93+EIAXKxY1k0L45BzAEsKaEBWJRoROp8ur+HVFNsabMC5h2ACFiMugrG
LQ9NFzkGJci+rR/WNnYAwgUIyFQrinhWUYxZkW0/If3Uwscipmtk18dV30LOwT2q
mfzJQluGtsKxQoXJJMP32AHt5dCsR0nd63PBel8vz7lfjN06w4MRzG1w4OOIWkwn
xP7kMIAzg0h8ETtNI12btmtxHl9ttvXg8oSHa2oZXwdF9Tl9EgSR5j85uHcFIz+y
1qjEcVUH+aLchpascbTWZrgtqxMXGbPQ7omiVtsbzB6IVMXnk1uC1Lj40M1TkyqO
yS3QzuFF8sr/mEQlNzptcQhenU//gJ4NEiyyVbhbGffIsfSNwGQp8l9PJtZY6JoN
7/LouT7MLrMWIOSxNKlD3n3bY7f9KG+Il7QIs/BmEXwCAX4l2vPjwso1W8yZdDGZ
81CauY2xNhTFeP7lcO6dfCofzz9yQgOZYMufwBgxpClXkMrXXjsv2nuXXvz2GH4p
oZwr+wOYIg3lQXa4pGpeIPtrL3JTAwUF7MKQ/bdn0tZ4SUQ4RrNYKf5NaZvkKS7M
VWloiGqpaZQTV/nen+8exkAZTeMDdpJ6WfQ6eQqxjxEPAFQtJnyFTwBwdUHdcmtw
tGtK+RLry6T01w6KxE9FghLBbqkNaaMH0NMnoTPdOcWwz97qZbqxRRQ6+6MALIEt
Eb40IoYgTYB4Ghd3IW8bh99UiV7yNE/sTtb81xLa/N1Alt3YUS/n+dfcCOsw6f9U
dBdw8tgL1kb2hEDnX/z+vmdWAHO8yHtI1rP9wmnCRCvgTO9fDnYIBfs4pwmYbDOA
dc/n9NsWDID0KsOUwvYXmnprzkbFKJkMw+2J0b2oO2GLXj0aZ7GwdkxnFL3x5F2p
wh9MFOo5G2ROgohG288ESAqpu7QS5QILcPNRbABRk7AiuoUkefZpIh6B3At1TP67
5ecOuMD2a0x3Pz0fUGKoMUGCJDefBkGOwjsrtYyueMSiBoAuBJu9zSNIsJyo3V5P
ISxIgX/Mizx56mjzrvyuh1rl2VKRvNxECQoRvTjht2EaRIgXYSC0SGcG7cmauxmf
7rpGjFKaGrZQiN83SoBtnjux4WSPdbp4fdxrXb7VJpBMNp2vWHgQffst7UuNug1Z
0b0yJ60eSug3P33LOUgBZ9qw2YCCQOeW9ES6jY75Qn85a3BugXnXLS/nNyBRk1l7
fnB0YMr+pOe+DBnLMCZvlOp1iFSEblpBHWO1PisUqu86n/CvJVz0uRlJkrNsY8KV
N3kOeJ1yHSkUXZMhW7Tb6JQ1rW+SjQVefX1Bsyd63ID/PsD6xYKHEU9GNTivAmK9
`protect END_PROTECTED
