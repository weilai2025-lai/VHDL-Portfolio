`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAjwIKIXiz1ruEk1nIPTDnyv+Jf0Mx0LbmyManQb12hOgzIqJHCW8GaZLiFBC5fN
9hOxP+qfTKnSbPQoUvRq1bwO8thIjwbkztZI0fGiGtRyFh5q1uxJlH0d7em+mIFm
HODhJh6iSLVCCHBiXkuxWYuUV+sTJaE0CnnYTCWKz44aLXH9ZVF150DWAWOEtCnq
6WvDdhLSG0+wwzeafohMK7xXgVOpZJX6IeFEH1879WUR4NV/54v01gniptYUfGxB
jNfL3pqvtx3FyVFHUJq6VBGCzBwV6sVhwCdJZlG5aDm1yK2yY24FiWD9hKq6WQfy
wmfEZxbC8EkWYZp3huD18lm/qernxnUFqgOeyKqudpmnRJumd9Cz1eQjquUFJHa9
Nq/hUUjtF+wQPJHFU4k+a6RIHTDcohKEoglCpPS3wYDD4Y1xKhQrMmPKQhCVRKxq
oKBbUllRCxXRSrVM4DqLuWrGZ5CFT0N4/cBe19ECApKJF1IrkpHRtgfOINvqQLff
FKBVuU1Ek0qbvmPy6DNgVYZbVCNK4huD/kpfUcRSm73/TCBvyoEUUqEhUqy5LgL3
kN8IoOVuzlaZYaT7spaBVllk0DVbBD3lYHId+RcvSzipTs47k7M83LXd5CfBMWeO
2RBibyKspSI2QlAoK0xXhiDTi7EBJzdj90LwBgqNb9q18g3qs4ZNARtoiXjKeCLW
LU1GtaWPfsvBxD1FcCBqO2jjJjOv7vJlqTgcr+NSOpe/gF0FMN7V+cZQzbR7YQmB
YCrqcA+bporJ+M6dw+nSn8cAkU+myBB5hKMu6I3Ej1Kr+qFNNvozDVx/x0f1UPUA
4Xm+UyZ/7xczRplWb6gZcUKCZoq5gWJ4o99SVuQBBbPmJMHvK9AQrG5/c5Exmles
CnrZ3mB3OeegwuKAbGReyzOustt0GhdbxI1NlJK0fEuj4mCygDebNuCID478pSTe
qbxJw/Qu7nbaRP37SfQCa4TL2zEKW8fBf4qvDXmP1z9uR7snTs92E6pikz4ZOZ9u
w8Km0mONRHasIdnsgnzOMJz7oHdixM754MZsrJ0evQHGQrPWl1ux5xaogvKtfUO9
0K04xYS/a7BnLp62rLijCBJIcmZgPcmbm0Up9QJFGjpjk3UvRprP3gdXxbkvsaFm
aGpNHc7kuh9K4X7q/FSmPZaBiM8EelDG5MdvURvAj7IljZ0aGdPR/AwmwWW8beF5
tXimmVdWA4x0DckU1bG5y9VUrxjfFJOjuCSWja/kShlfOJSuSCnnbe9HihvfrbvN
1hQYQVBmO3l1yWLIaG5sgHU3bLB2kWFBsFLwqBt3lWTcrs+pFcO+OHsKRaHofMKD
YLB7LTLjYV27+7hMIvJYUo3mwkrZSjbzAJ9xeW+VR1fr3gEVadCpJ+JbKvTLFOH4
KvRsJc6RBTZ1JF9d6ydUfqm9VUryVr3akkAQVrHc4Hk2gafzY/GLH8JfvQ7JwWhc
+eMUEiWUC1Mb1QJBeNRzvjnE1CBS92VQvzqDIhOEOk0v5UuTgMAXdCenPSV3gp4I
UGJW9UfY1FNKjkO0zzRMHVafA8aSSoQ78tyAxioBEJtYDstCbmbb9iWVvqI77tai
95nD88UF6FAvt7dE+l6V8lY/zKWUB3Dj9EVcsdxYWhp40s+/jkFJsTr11e3k199a
v9b6FF3h7qncHaTgprEkTk84F2qXDbMLpLrXv/LEK7idXY0mOipGxS0pvrg386sV
KpgBimSB21ZGRYfglKdGGutvGYZWe44tI25Zupvlbsbs1qmakBA31290IqGER2Ym
bli+HlUaThL1Kffc3izPj9losXTGUL8J1iram8LuGgT5D6OpC1SdcJCCz7dgXPqD
w7VM5MxV05/57XCBUy2uCrQJ1kpp0RLZYGYyqb9Q+avNrPlbhmtB8/PXTEEmfDZ8
SAGOTFEMyU5/bh5Ko2vHMB6el50t7K80w/3ui2P99u3FBbi8RW16nLffwKrtc1SP
EvK0z+KHWHvfWz6l5KiceHUfxGyA77BRyFCxNuQL5udv28pXU9WUtOmtXRchO15L
dDcisv+xfwm46TJyc1rRj+2hgT/uMFhV8h1XDOHmQptpw3DluT7dnU9m9O4mgbv1
+7M/uGi8tuIh8iqXoukjTRcerWpGs3Q6wAmd2L3TktjAueJgqs02gTN0hQOkPk2y
HuK92QLWT1++Oib27vDGsyMUv/PnlNn8Y1vHTl0qssVQzu6DchdwPoJUWIUcBZ/q
z8iVaoNdqdioEq+jKfcCBDFsGc7uW5l6KqOlA22Gzx8E86Ig/3eCFSTqPLY6LGw8
QmSc6mhVX7vdPlMgiEI7e8Kf4X4wGSd8uGvqnKRXQ25CkqRJRnd/bhUg/BZwYGo7
nrXJuPC60aqiLecCCZyUemoE4Xs1gLb1GBwmxm2PJmZy53L+UabpWTLawe0DcuaI
RI5BHSgRuBnmUYWpfT2qT3pcw6q87kJVnlcga2iJyvn1IwdyvrGU5XVzIysa+/sv
6M8B8or3DdA8U03+ydKu2Sk1ojCKsGPKUqZPVqSXomnt6QO9C5Cr2kECKOmCW8Jf
Vru7DfgXOWkf0P5zrOc5ERqH16zR5eMF3ktWufU0p8jOmp9tcgs0dPK21XzBnN7C
Fc6EayLU+XjcylilOk2XEPcYuR6CTcDlM1uq0pbeL4FNO6vsK5bNAvJkq2WnbvmP
YSZGjdgns2Alk630VAtXJ9oI3Of2G2tvTI9PgO1W+2DoQHdfFn8XezttXkUow+P2
yb6WObDnwU0QCJuEh+safEHMzKZZ7BfSP+AaG8b4dM4NV47feP39tjD51hHFWCvd
ieuB6zzLvEnIukvOXrund1yiip+W+hOt9Rrgz1UmAijK99wz/Ax17371VavBcPpv
GbCcyQjfVXNNIIG1ph4oYEeRHdH85ZDTkQzOx+xsmaHZC9lQ1LAiFu/Hmlfx8IRH
tViAeRJwDow9o3SRcN6+YAFzc9oew95cf5S4s383jiXjYc3dA/c7BUuWLsCO/Uip
aQX1/k0c7FJY0ue+F7wTYIJrz/NRT624hPAuH+O5csE1gUpWdfwK/AMAOW0NfQU8
zVQxYFKEO4l+In9qVYffk8w18ER3FAywZT7y+oECxWlDGCzb7FvounahlG1Oy9ZI
vZSXVzH2XaBYCLLpcUbktOgWgyGPRZH2i5N6uo5I0hkGEdEMDhMb9AgbJARxQsng
jei1BN5eS5k013CbaTF/t7MVyyLhT68S0vIG9tvdn+trKOpxHBDBGe6EUrUJD5Ga
Ve+/6NUqOOuWMXR9/mn4MTRQ800Oc2BBO5VISxRJjD5KtEZByB+9LeEx1tT/qMUy
FKQ75vKVzHZSR7Lau8MK1xbjcxEyhc4zPacd/1HuZnXWdUTRJgWo/ylgPIOA+F2M
9V+XLfFMH7gXUbI33QHynUTML99Fbv9tgyVoLnJitEN+wRAg8h+xph4FoeMLo8eK
hOqnfgCw8ZqAZip0Pj/QBNEXRRXrVwZXOuEQZwLGuNIeGrglQ37ynRk+wrkj4jHl
Bx6clyUj3N+GP9s8CsVt9CH9F+RpTRbqpZFr3D6pybIyvtwi7qbCwexzXulV9b01
UdBYJvvPIMovn0AjR82pAoUJXsGfn21261Dq/WNOw0DJGrCb/WXH4TrK3h2N2w2B
AEb/jWacBKKrjLP3sRonGBJDntkkX6oi0fLpntm5jA492Hq1v9zbTYKquaFMifxc
eaomJjHZF03SG3kT3MHHCVEujSo0nZp9zktgOmBVZo1giaqHKo/nUzNX6MFKTpAk
LeZNadk3Aejg5KLS4R600kqsPD4CcCItRyNOA1oH2QXTOcGgXa3iXMsIJcHe2JqF
x6O0/IN7erPrziJlbJOBXiYggDNptY/jiyasQSgiqPAu27Me6Pls2kAMTh3LxHkH
OW80R6tAttAEqtwpw0RkXxPNAwcnM3I0a8eQ+2sYtJUr5kf6FPsQNZ+hSpCzmFvK
LkOaNwMv8FAKxAsj/TwV6N9yrUo+O6wMR4WyjnIhcae7iRW4egS72razxWIhyxEv
C8ujJ4OUVUwIJfTFRFXmcXvZfcPWC0jSpiJxtcEr0jkOI4QHz2r1I/9J4Y+213ro
kcNT2bhEggGo26dTwPXb/Yg4oPQxdbqAqfGpEtEDIL3JDnOhmsX6IcWOPJOTy7Uk
JLKw1hz7qntZO+tr+2QysIRjfHloYo8ShzTXZVwcJvRsCsGgVQJi03XLfo6B/Xms
fWTex5y6x/XswzBVJxTvsc88gGYyA9oXQksJzObiTaE+3JwKA/VfEGd2z2rOptNH
6a4nb8TNWfg2Ad3Nn8XV+60g2N7tXrWaZyy2mhsqgGPAu8vIChpyhjgYeX9ExBNW
N/Ge5upAm2jm/A34AyiLJgUr/onhdFea8X0DyZqCP6deupLK/eDdg08RMU2KVXZ6
7+9hXiZGfj1DI5VcL6FJ1B1PjptQTZDzNmf4L1/qSwHmkAfFVXUZos1xLZ6MbTL4
ldgRYwunBfLJBm6hj9qNSOgEKAbBzUb04BguLd5QagSwOxs6mINTtVyYbP9hgRgm
43L8WZONKglb1MmG5a3TFqa0P4adgrE/M7SitA+hxy0X4V325CjI50oO2ZVbPBUR
mebQaic48uU9G5pPiiD+f9bIPf4uP4xMzJ+nA2fs5J9CQ/ZxcK/lA9NgRLKsvrXJ
CeBHSiVv8GAIg1qOvA8lupeER9yQHUoYOKiRBvDaRm9SpIRtdO+VnhdQhrMhcVJ1
dljqThopnOorUOzeRZE7/a6L6zc0WDzGg0qqd22ByRhYXrmIy8bIZPn0pAMD6Wjs
HNypsPKT9+LhtAdgVDdoTR5udZBrexKzsPrqlvaNM7DW915GI9c2ZfPc3NfjasiS
yeHv1jbASne2OMyy/oNHxqc8Fn67pouV7oRDdcZMQjwFCqiGZsJyjoeVdu20+i5w
cRMJx/CVpPrjbFya2gg6aG5czA4R/2jeLTRT+dhTPcsoWb1LrfMGllhyUomAkHQ9
kZbvbkw7XvodrQoXdUskQsU02vNsHpH0IHGimeb+3i4DOr/Wuii9TgWf4fVQ4E5P
fbAPKs7Imrf2gzfObP4nZ1bZ7QxJc4Isq/1aWhzRDNY1M7Gy8rNsNY0/xnv7LRAr
NDuTEr8bq38dF/dF2KTT8kzhu75oF5Kv8eiOWOhyZS5+aomBB0SkPGDQClPfheEm
69ss2f3MACoa6PeLAfpO4RWNDZYsB5pr/lA8+754oOTD2F6o7UKIZsSsppq5mK91
NEMUPjpIqR4MDwN6lliBsycmkE8jjWJZ18DQNIFxxzMtcxrne4Qz+vgydczH/T0C
ql3E2zV35U7jIzoJIzxWdrpQ8t9GHe/B2hDE/M3oPKtms4I2XxKt+cj842ONqtGq
3xL+hMJiZry+dXGwaaPFmAWv9abkHRGQvHGzrKrO8DYlLOVQHlHtgDOOYGCLimcf
eu2mNvXaR0Mz/AyKOS745SfU0HtByOTQT5xdanp5RQ++fD5BuLkHZ3ESazDrAUDW
3wqnvaBhkHPIAfaakVvjF/1vZxxZZXgUzcPe9SNAZE8d8Vn1Dr0/GF5SsOpyU7DN
oq/9MedicJWTn79juowmSM3sIoo6+oCIz1t9hbMT8gvRWvxUTT905LEINMaHR3og
C/EpKfPmPJ+F+te8fq9Da4eEG7/3s2QqUmJbMDaQzE5U7nUuopzKJUfYF9B5gyLQ
i1IL9fey4B+jxiXGEhjZ5N1p+7miplrRGNN1kVUBc2by03o78gYs+CTU288qoHJF
sAyaDPIyIhfnvMhE1IBzmwFEdgMYqKYGBwEpnsR4HkJVyEysoBdv8uLQ0hALVXX8
kUzRzZNNODu0ocfAvAw0AzqPEFz4jYco5a8bnpkcTB6ttOKRiPTB6JxQf+rDQhUp
AjaG82TV+eKE34X145RX5cTaLpDHOmThLQ4tUDvdjX38Uwk3I5uCp40nyqac6quT
JOFvDbt6PTBkpHjcUk/UPUklD1dzcJn2mlajSJtAAoT4SKZI501xRQQlpa6nVhwC
eX4nKhKGmi/3t2jcV/M1rkOMD2F57nmbTPlYw6GtmcVvv5F/6C/rX9r95DVvg4TV
MNIQMpvBX0EP6ixl0y7ZOvHaCQiesi5i9XwwGWEtYvdnaRG6YAnQmpelekLzq90Y
oACFN3KWA0WJFKWFblrp6msf6/EGNW7vPg8ctOqxvhjCHbiSrRgXBAof+Ynnf7cR
Nn2op99g9/8OP1b1ZOhQKdeeOq8IoRxKaDhmjHa4in5lc1k9M4+2robVMYTiVXtX
VJosBIDIlJgkrSeqJvferIyxuLNj1yclCy+rxJRgpehPlbbrAPwBqkaaX4WLqad3
H6guK00eEuXL2oFxXcSghQ==
`protect END_PROTECTED
