`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7ePAFNXUeudwZRA0Vq/eSyFdd0n4+HxvXtmNI2xqQfPgj3WxC+P/8pxThOE0r96
qcOq1HvyXUoVc0F4FuoqM5rEs7Aej9xM/7F+1RGn8lS5RQd3TeMB2Av70H1gxdGv
M7PlADvBYa+Ua0cudurl1IzpyyFunF3GIQPq/iS5RuMoj3xTTHjy+C4H9zwIAttn
NY7alpuz4+EypW+fyggzpryBMKhEn1X+JMNM46XgGVAjVOXZ0evGG5dBcRq1UBkx
IUL6sL1A/kR7tDlUZM9C2zSjBdSYz7ENBenRP3lS1utb0XKBO3WzpDibubvr2aXr
Tb+1jUYYgk3Ib/JuG/VgNjrobPDkbt51LUVG+bTivUSmk3aeQdcqL2OpLnIizFKq
m7fZsCxbxjfuWeMIEZC6T1LwC+5Zp2D+ldfzIKNx6xm/wpFGbOFxOaFqWs6PTakD
jPxetodgCoDsi7LHcfNPtxwsHHAIpnIPFCUY6k7tTPBFlWQR5/x6lAd806j9Os90
UPCDZ6QkrDLTSz+jIpW4f0o2MOGUHiVgYWkcFdYZvRVnprpArDLhu1Dvax0D0rq8
at+MKIbB0OQEQSI3OFGl2XNA3w1S8KCLwh7zuMJltQm6ZtzmgTU3/Z3EVIagEGGd
DwyolOrWvht3OH8eZn6cc04phd5lLWsFx5vUSu2U4a7BpCN9mUI3ZjtsTlegrld1
VCC4J0XzVt/P/bw8hdgjgLDnTUZ/ngF2TOWbAYk9MIX1gnSpHnPsB/kdlMS7mbB+
d4Tu2NgisZwcRwfLNgBNHEWgze4PQlGWyJsI/8wNYXMXucUYRXlcUAZIFQjqnSQT
dYJVNT7tIN2jjJH1+W/dvUGuM8ehA4uRqy/PYbMo2qjHYN2kcA3oopkjOxXjjVmT
`protect END_PROTECTED
