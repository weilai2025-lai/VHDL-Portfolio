`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y27mPiHbwRo2WuMLq1cHroSQUbi4B8cpZZC1jHzOGBDO3fdFXoav3tSKEzf8OCiD
TcXsEhQQHgxbE6ORCBo459P8ebGxSK40KPEqyyNki9QHGT9PSONIw/K+QkBd5ENZ
yN6PKKzMWCr3C/I30CclYv/Dpj9b4kjKorSZCK6AtviRjnwVGNPgLUYeAYSwrTsj
`protect END_PROTECTED
