`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBoghDk3xnH9uy43T6RZ2vd3x9HnLVtXCb8I/5o8+9BQsY2EiAil4RjcnNKjrkH0
H/oNhV+Jo0RTuYMBy2L3+TijlJ50qLbgRS+JvpBHjt28BwO9KZpWK5lMdCCwTKsg
BLUn/dYnUkamycvxYKeDTgcheQqZhmvzTIyZ8QdWuA7/zetGBFQ7+i4xARK2vj9l
HFVSpMfQW9alpL9PXoKmNuz6AM5VgFk9w836B+SdaFTm5Jsuo7ZTm+0mDqNxecuE
0BOF4Nn7XI8wUq4Ub20rq3sORbB62FqNoYTgrNvoWj7f35NlA/xUuC0tNGqlgW2M
HgclfiIG3sPmMSjFbpTxkeOqFYVjiCxTtPsB+EOrzO+tpJ2iHi9A8Weitu+Qa+5b
Rrx5yzXvv/dwWQwKsTuvwC5rzU4ZnuiscipPt1fZFqtqJ3xyGWFDZ5qoEtFNQmvH
SA3TMak5pEEnevMQpWldXnn55dE/oFXNH4PwPDZeBcOJSsAaicfy72G7LXr8RTYZ
wNY1uJtazHNGXvxjET9lGdmk7wAeL045XIYIi+PcT89dcvIxZCzQa1BUE3NMsHtS
B6Ygry5j8HmmaPx7AUF+b04IiDYF1eIxZ/z6Rz+2AW/0ysSczXPq0eB9EhyX0nY1
FHqLTIFt+2+PFXKCemQzZDRCQVY0WWmyPHlrW+X2f3Tw8yPeY4NquXcUaBYKHC15
xW/dsmYj3NFbjIBOkZ9bpuFZMgJaqjE+ZLPuCWHO4r8IULntFBzj2YKmAL1qv4Gi
O1iC3LM3faaweIA8KWCS7N4m8iuwgzbDJ7xi+MC0TvsaL8+V0OdJPB/u+hfIzMJ0
65LMIktzbhPNa4DCsws0ue8QRAYgWRZRdm4+MigYtKVe1AfoWn3qqxBJpYfvXmJq
B7xE9kRt9wRcZRMTSP1LcVFNktnrsyh+pD0xWjlZo0XH2OGWXb2/bqYKwZVlkC4z
H72edUqV4a/GkXWgQsCrGEGmVPtwPaRNDeUe9GKzsq18cgeO+8wUDnTh18ST7IQi
tPEYngXvAbYhr3gon9MTmuqiCFtX5kqga4q2sqLpmoi77MZ+TAOhrN/CyB/FbZCL
GMhko7FkQUX2cxmFzqo/p2d4ZAcCkbNrUI+Mv3ve1mGWlXjy///nC9qeIXv5G120
Ln0RWwsnrZVjopEe/Ef+7Qwf7za0Bs8S1yAZ8qTEVBw7mG5MblVk+7tDijTpFr0k
fjSB2awJvKqj5Fr6QxnPCg3X69LBD2ZckvGBrVCyEZLLhbzGwzVOca2DEJIQqq/v
k/Tb9x0AUZmTbh1njh3Z2OjOjI3Hs96whez5lOlBAby4gyq/KpV63Bh/gn8FJSDp
nEmd7xzl8n2r2k73tdpRE7jJ4c7y6WXvEQKVLmXnUnwMH7t89qzBXUXXH+CkUvo9
Nuf67iw+SzM8AmjfinJBeCZMgou94jCrm6P7a2fi4t7ykqsAX8/Lmn88T1e58E9z
Vx61UOloIxQ9gR3eri95ioPvssFyd69KeSLvzd0PfkJURbf/04C4a5XDDqetFAxx
YvluICtXmKOh3DLFVqJ6Tzx1zsTVlGgF1cBCQyMEGOb47w0mYlize+UOBNvRt4hM
KyeAXPyFuyVHGMtpxuDQDvWwzCSs7AZc5cXV4S4hC6WWhhs7s0T3pEfJvIhGgKfW
GoVf13I2n5zRgk3sIeUqxYRUIRS6StCI/olFEwWL7iephh2hehxQGzHLF/M0VZq2
1TMEi0j0QNhgWAB2BdMDfxSi+FnYXJ1htv/HLZ+oUsFHjbypm+1iPzK7845B25Ci
V5wc6qjJnmTUwUAX0qIJ+ws2lyl+YB+jSqfpyfmFzaLUWp04y8Hay+H4uT4ls1Sf
Sfh7B5iXghYU4U0UBZTkwtCyJdzevLedTpVTGJRIzH6P2jagZcExTkFTXRrImJGl
zlfLvVLY/dlFlEgJBzzLW80FpQpml352EnGasUg2jRa7pJH0MDO6UG8N7+7gz+Xk
BlubLgosPSfiJcrv4R94TuNxlN7GfLvyrRLb+S0nsZhhEzQoZpmXo4Gw625t+zmi
ghmAmBrG8DcvuSrPfd9REWkD+XT9zX71okm5YNDlPBSc4TYLa0Q6c0wmr7EndOGB
EsKgjPpW2KEo3mOjBXXstv64G7ITCOMnnQ/bwKc1cj+Ui4jk946H2mTjDr9m26xh
RGMDnDn+BsijMC6B43VviaY9dk/sK3su8OYzqCD9stj3TloM4QVYHjfoVS6TQcMD
7FVv4Tr97+6m/MbPj2mwWDyR4oG/OKa+cQivnLXjr3uvQ6GezaQQjtoW+DwGWqLL
AdYqrp6LXRsijQ1rbTl1V532OCE9kutsmNAbTTJMHymlipWDQwGwI2ahbQ87q86Z
C0jcB99bofk3OTVaCGx0SCxHIrL5RAsuDfalUUPoS2YfVbbxCYj5nGjhEne0h/qI
4eDjlqgJ8U0ucuOu8OcjZ3Q+dvvIJ1y6E4AhHQ9Th0KgQTYlocIvFbsIDjDar+MJ
YwIIzcuvLSjf946PZU1V9SH+yFZ5+H3uhVtWbo+H3IqOdtcSi67yKnNeafuLRoD4
+fg0OQl+dLyVXVjrjrfORf+vMRgea711o4uQOItzMvqmRnDJePMw+cuw3GwNbCF7
vZwG5iHBRp2AkWniK5mvU4ReGf+SV8j73n6nmn0ww9fvoj68fE+skxtNKZ7Wlxnl
vaSlM053XigpIiiIlJbhLnnaKdp3XuOT59/PuESPExc9IYqY1Mocw8NU5WbqwNbn
F1f36rb6bQW7n8J0H2/bs/59IKO2YSPq4u9XSYSR9DZreMZ3toTDcshnaXlrVOz4
lM9QaIVa54l+QO9U7bfNW4QasEiOHrEI+YbWhKaEdZnGjF6XgG4xQAfIXPp6sCm4
LkVSxBxuGEikpICaiVtotBR7IT4gzEEEgfJkBEbtgf72EzVfJrNiL1CJI6XyP8c0
XI8av1jR23gZbyrr+Av6y2T3yCnBsSVBbiY6X+6HsjvWVuGk1rQkY6xaNNWE9eLM
eZphqwXxS1EsaIsdpfMJRY9625JG7NL1+6afavn17Di+6fLxx5zXGSa/qo/BYsFv
QbgV9kd5yLRHS4uwgpf+BQWXD3T9BmebfD4CfXsHCG5ENtQbKmyvky0vqHeyjHQg
J3M3dOxpeGvqv6jYONTRBMTV2goLEFYPPmhTB1J9G/6Kai0tnp9P6chfSY4zx0zG
kFiWiOPETWtmsmuFZYE0JVrKMRNiWNFoYLlqoewDA5sIC4YwNh0Z4g4muihl3wR1
bCamGOcIeIJysDR/RUNCIqDPzFRzeCLWqwismNfTUvPHtMM6vatufd+SjV8zqx5o
l3bOSrK46ZYsgF/ujYxn8DV81AGdVhxakoy8a473TKO1UaqnfDK2RlrF+gVxHTXn
I6LRuv5O4QuXzifbdwfo6jZMiRWSnBunTyIGDKTHHVMG6i6cdeViqtwVMRZ1bMpA
bOeubnPfeB68B/8IZLWwtSosaUbSVDjFYdswl6NsVsue8bRx/2RGhvrFHKDjFV7f
DUx0tVwIJ9dsvL8qOYpvaJGF+uAcm9LylmpoSgRFtxH6RwY2F+bme/Uj2ueG7qWa
pKyy9J19+1FibUi5E6MxsBILwwVS/d2rGU1NS9D2d+/GnBwSw9w+tyIDy0DOBTFX
3P8bed7Msxj3kLS42MQJHFoStMOf6iTzcVGKx45HqjLjgnTYuhaEk3HwTWrUiKW9
1a18lh+SQFayoi2kbg752H05caKE69a46907snkhzaJbWiW60ibmCPSMv5XxYayH
9g7PkTl3CM4clNszeYgt2i9/P8msd1ei23w6ynxe27JfhLmXBgJIbcf4TmXp/Ath
2fGlGwjWexcXkE0RYKlDoK0muuHWiXH/FHRnicgFTMwudIfOxjPr+Nyn/M0XNAVQ
9T+sY4aBfS91WyRlnNVgsLvaaMaW1sPs23UkqdFYOD8+vr2cmKTI5/z+2FS2IBj+
GqIdGblYvyzcIDDtIeCsztr+M5V0ZNfewsyQfEGTsGNk7IQDL8lwE+GJv9Q5OXYc
d21DvBFXD+yQdWtikuedjOTtUPo2o/ewnjuFMW7tpMogwX8/hiuDnxNCQLRkB8z9
uAzUccZYmRph72DWO4Dpcm8PXUYwgQitPcnjbQfb7ickc9P8l0AB11GZ3+675I4e
/q7eEj1GVxhKkVL4JbvPS5T8BSCpGwOGVFNneYzKGXyQI1a/OIomGHdvhl3q200M
MYKOZNWrxwbI1cCNt1w3lpervPqOnHZYAy/pPIRBhNI7NA2k61RtdEhgPiTZp+4b
KCwHfzmoSVWutasb6vO84g80sVB8vPO/YbrRq96jq6krWZ1kTyaAnKq12EWBc+8l
0VETly5G5/JgLj9PdmYtpL+fGiavaLC+4jjJudVe327+QMKDnGWw7Qpiu1yOjR87
XxQ49NvlEWpVl+GBSQOJ/uip+JPGg/SoR3yCMvVKx1s98ejjGrZfNWvkFGjc5m3y
OBGHJc7NkkEmO6fOnTbNrIBLIifV6/aQkQomwVdJQFg6G2IlW7QIg9fVREYueoCz
cqPC+51jbzyg5HdBAoyWOr30nVMLfV3B2hrm3ongKSFOfW2R7KUhR6bfDteniGZp
ab9IzrJCXp8PdPzyVxOCAg2NYboONghgEaLxoyRidm9PUB38ETI6PIIE8XBJMjLv
sKDQctXHDE8ZMZRAFxWklWMcY0T0Z/QK+RTbUgLisO8YWU+ZQKQlm5iE64ce87ho
UjPDxvtMJEwzL8Wbe4mnkvabMu47EqCi9ljfPkFgUoAyW8QGrf6NNlcOmxFuXH5o
UBe7s33bcKCKSOLh6Z0kOPWhkVg0d+rsC6IbNke3HxIJzkFHTv2jiog3e2hy4r9d
FlEVBF2RHS127LxLcf01TLBuLh7TnMnet6D9OsKajxfru+VVYHPxsZNIUkoYnDJ4
QMLEWjQ49To0ZsvubHjMsnAMMx7ixZ8co1VtIwjj3rtdFzDjhP4K+foKL8eSgeMl
GoJxTpwQ+mfTF6t+ugN3bAGsiuvXGYm761uY90y9ke5/nxMHfngmLkNIN2zRGTlI
8u1AGwrT/bZBSF0CJMD0+XSwsKoXrOJLmKQE3wTuki0/fnfcyh3Rms7lfR3/VQ+t
CWdgMAKQY2l1LdMKeLV5NDzpr/3B/1CO2XiYfuM/vig27iOJwzQrNHSJYMG/MZHC
hONU8mDN+aTNHLGuL+G/WqdRNJPWEWerdRbdfUWA/5lxIHbHWeqjsQQe1p7LmRoL
PdlzQ7iKFdeU5hzY0Ub6nRICyBPOk9k+Z5pGmHKBp6VhwZQPpfrEumuq7ejpMznT
UVWAJlsyF4iof7ys+1ev7Aer82j+AFaZSu5nzE+4PByNMQHt5wr9e8fxc81D/LkH
IiagQNQRXCWG7P5ggOU1E0ZGxf4bHzu230hJQ3aurGpU1x7bN21HQAjnMYxDTx1o
F07yEI9A4xcXNO1LbM/DiYVkecjI6/jWMVF8ta/OsiDxDvi+akfTdwcrba1MtT9A
2cilfiXL+e2wVs9+elg84hw2YgxtDwMCbSQOWng7tJItkqYP4dT/D7OGCEFDdYH1
89+/CMko9sqcJKeuP7Cfvbev6HhBJnbbpyDQ39XdKjYYrjmZbUGG17PhY9hKijnR
cJWtpADB1gB8aDSUSuunMbeGnFlRlfWka8rj7z4/tYMVdq/26D2gvz5bt1dPFWjg
YNsOTpRrFrXMp22L/GQiof+lXXzktCpfCVzIb6dZtauXW1caxe0tDY5p5AT4mqXY
KMD3O86DRpUIvOtaCVbDW78bf1NeU7uxRlTP7cHyE4QwDhotOEgIFzheTticO/Cy
DhnDvC1n5P4ZJeramQHSn7uwYJqpc0GIRVet8OFNiDe+nLrnGHJnZHZ7hHQpFtVk
H/mKpUdQPzyopAjj6CtXel4kXKek76KAOiTB41MBAbLk00FFk7aH5pcfGGKUhj9M
4K2i6vRZo1rXmA5LqG3E9sUhL0mCTEKoo/MMDl37HvIuOZHiSORd6h8X1KlMFaU2
f7BVCBVBn4s3EcMa2GoUFjI6cEpjO5TVumfjgMJf/7CSLdZekPB4xBDBnUhTxINo
ub4y6nE9esgaF0E7tSXIJ7eDs2pWGcjXGysUuk8cdp7zqbUdwZOjYz15vOmSM5k8
3BEXBBP4l5zPhaHv8L8xLZX3g6LPOf+i5JPB99Kdy362jxFjXcghBVzooVieWUdl
BKajljHnEglWGeXXM1A7oAMjp0bDxhNPDomoD3/WE1GitRrixb9wotabmt91JtLQ
9Vr1OOHt1q3b5eWv4OnDrGYZkOF6BzwJ8khJlNlNeaS+1ssczK+u4MBhhKkPCtRO
CP+qaZ61/ESCILjIhvIJEg==
`protect END_PROTECTED
