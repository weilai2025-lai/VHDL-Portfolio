`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLCKX+KPNJ5cvDlzeB69LkpRNpoS7d+UdIVs8Ks2hig2xQOGObMWcs2x8cyMDW1h
L0Z5KeXliLMHy5lyrwc51ftcV14Ee+Zo3e1NfcWfosmlyaxGAjm2Sk4qc7ENILpW
ZL0HOlvetPnKk7cPFsjKipl8gtHNWYD4Rj7M64HZTsyIXxMppyxptrHNumdb4lkD
mOySMshr38MQ5RiDSgA+8Li3GdDTmQTuNuY9TiKcnhiH+6v1hJfysmGYTTT7GH2b
5sbHcIKgWf0NFnUNU1kb/cXO94bYTgAh6+7N1Z38R0NazwE+IxtiPb4RGeyDREnB
s2s+hb2uRQ4sS+Y352Rvnf1H+FfXvrwCUEI1qxoLb8awKI0v8b8D+Pa8OKsjKDDp
0V87HtA1oOiL0EI/QbG9F/5ScX38YYbJ7U/SZH+Bxh1vQEnIgv/JtC64HKlROz/e
l+NMoSqNE6/pjblePUiMHjuzqMI0Lpbtu1edIWnk4EOEzHhZQrZisPh8/yYlskDf
wd11FrIPM4WoFGY+5BRVCtVvKATlZZ2paTEgtJ9FzLi0kxWUKa4NXEbvpIXKYqBP
zEYjJQ1V7Ui2WPKLnnNz/49fNb6ZvbhpyQA5MrSgP378ajwyzdUZ3aslC8JmOvQ7
DdlRhGaQ/vB1tCT59E7Tb4OQFMy3Aepn1jD6UXly+fgr31KSnDLxaXpK/d+fDgMY
7OArNzwTCMC+c6gWuvzFRdB0UX/w2yVpSB/ZYINrqe5OF9XL7Of/4pXh8y/eowFj
htTKE5b3vZ2AnRe6fbCB3QHKC80ALmV+yhWL7o7Py/Hed39rKdJE6fD8BTXFIFC/
Bypmc0glIE6EV1nBndJ3eR4RaU4ws857OhSD+kyFKNajEIlVj5qRdNIkPSfPiJGl
fipjL45iEjDevnRg92xDsKPzDj+Dysq3yjV50jIXEclC5Cme4BOXH5EY9yOWMCLz
piAyc1Hm686MF7EnBl28QVDg5woAiMcxjBB9Rmxs9zJKMi2B2JQIoLDViOdD02Ji
fjn7yc7ONzBB6G4huXIpeVNjF6Wd5+/RNn+cHefOrkprd5znPFqcCNa0uO+XcW8T
RhZhb5ul3KnP+2N8hs0gCJvhReo7/lKkqRxibEw7N1ggnBlB/7K1SrUlp5C22ZWu
BAeDQsj4F0RvfGkABty5k5TF0I/UEqZYZeTlRYKlSyfS3L0ZSly6P8aroRvWgGW2
kinc9hd8TXutSgViZMa+E+h1dQo36NGWAbpGJHhd15FPHjO0fAiKAOdLn9LQuqsD
6uIGTltRLQFShSonMWXMLTKc62K2JDealv+yKN2sVo9w872NyODOqTNuCM7BDZVU
xBsv0vQSa1q1vNIbLwuIC7QIuCJ+p08Yi1gqXaaYHCPiDhkDBZHcBGwoRJDEeFV7
XZCatIW2pq/gYwriWt16j9g2ZwImQDAXzXVp+2Xy3RrpMOQ/qpaN+A8h7JWNlKjH
JXlHFIvRSAX8oMowosFP9aJkbvFx+xe7hVJcfLRQsHAwCcJwymomeaJYmypPl241
yPBsDxtWpMBtkGEz8JspaffyQa4aodCyWPzolr9sOe9DBXE2uxtkGSjCLtgwk0/m
9gPA2CXFqR4wsCRYrI93riDejaNN+WX7i/txLUQ5L73P3+tKvgd6Bp/4VCBzk17H
95p+nIvvbJJvLoXiCkgrq3NcXPMHeboqm03uRR7fZdf87S3M3JXUkgZK512LZfzp
S6TkY45vKj5Q4P+cjbIWgJyYQbNOBEd0Vc+RIPObr5BNMRuaZ1mkJTg6Gw9NKuIu
gGByGsUpOj8wesryE92JIXBmCnSc3puEN4awfjfQIGOlcacnPeGLu5XTjgGHKUdq
Yaj8qHXFz2eYGQkW8dbUaDPkS3h/h42PkHdCyBC3+EvDd2xve787OE0uBnrCidAT
dCh51cSTo4TBD5Gk82b4DgatusLQGl7j3YNT35d7RE/ZJW1c5XmYKFghk/E5YrRT
0Bu+RIlydCKrg2W/T0xovHvGncrp1HdDWUwLG0kTGhDK0EqL09peVYf8EEx9tOU9
OAy2/McUS8lvTXmrbHXgiBhAAaK6MGomEA3kcl6dGlvblDokVE4740bsLcWc6SZt
v02EIwSwQlEnHIqV/aSlL/mRhqaS5OKwpBmLEYzZ7kSMUnZCdWnStRH13sO5qYu1
hPO/WTcgX+ntHbhBCpgH/Aboj/SOFSdwpAwq7QYznksb/2DTSJ6zN2nkV/4rqy8I
S81McRmmEDkF3zLVKCXyjLxSochaXRMZdi5RRk15QHyeX10AEKzvfeXBKik1dxKu
XuMJNz+MSoAILhRnGsI4meUB6NqID5c6bUGlbzzUG3kfbCB1FPfxQ+0/8+C8zMXQ
TQc+8psC7P9OoiajlOmWFmqvgqT0rYHuseaAaf0lNC4GURjwi5tCDDjYCst3a6sP
ixw0beCm63e3eqG00uJH9ieKBcovt1qSaiED48w7CAbePEr7y40TNrBuNKwwKqFQ
FhHwFmAeYPqOJ1pPt8JtrnphvZRjp+q+7OPDeBCD3yPsbausAT8iUUvCYsHWc3G4
I1xXmPvcoy//K0WR19GW4H6Y4aBIatzX1q98vVH3auo2tXxXNOIMzN03xR69g/xv
UBK7uKXz4cJ+F1R/VhQdM3xjqeTWuogGI7WoZsWxppf6NrAIXZbYx1YunY9y7jnC
ojrUby2N+CCnd9+TVKEgT3Mce2iqt04bhqwAz2WxyIHlBTCnuAP/ELv2ZW0UnG2j
HA0bNglQVHPZgvSk/MnOHJnRuUl+LGyyr1oaYBRIF+u0NOcV9H+tdxHVkcrW+ScQ
yKeJ+KXiNefsPMjg3Af1gues9WlVlH9IcvkSmFH9nIygfQjaS3kRC/G0RGqKt+Sq
c2pmnRQOxbAIWDKKfqDbDQjmAujfB7hliuijFggn/6Q=
`protect END_PROTECTED
