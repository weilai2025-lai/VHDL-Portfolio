`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMbgX/mISemFvmE8IRNPs1uebd1jSf1SWhSi/teigOtFKveuwwxfRWjV24TsO35p
nKDRIJpJQcRJsTA3LKwbmY0BuegdL6tFwALOYMwQ923xyFTM9DqhaNDqxgWGCS6h
eis70WMoVYxF8yrRrssedTX+wF1Rzay9fWbBKm9TKjatjYKCUlLI+NUBopqcaiW+
fX1DMGL9sPNSTngRGixj0Vvq1P5sMjrCXABFKd3RCTfRHTODGzi+xprDQyhvLqyO
AbdhXxlijl/IXnMS3a2+8OspLSLyFi0zBJoOK/+DvNiJwB02fggZwTvtZhpZoqPY
7B8+jC1HOn9vhAVAZPiwrHWdYYsh1V8oRTwG2u/9KdU8Yj6uQWitYBX/6wz3XvGA
UGZR1Labfn5EI/DnxqXA6v1WaPnHWlInmju44iy1Og1k2q2FKnux1Hdr4BdXinsO
htazKOmLaUr6djKLZVKtj866pbTeq71wRwPD7KAbk7A/5GfQ8zCQh3cmtVsOidLF
eY+By7qlVnkM4IU+wU5P8w9eII96IIdHh/0/ZfHvVYdn698I7hfqt+NKwLGQKZC+
TyYQ2KtDZH1Vg+pD5OVqQr2GvE3CavRhTvFKi+OWsb+h/E+wUp2TtRrTEtTb5H60
6VHABcg1yiFr1Z8fh+YA5ar3CU4DbMc+Xau9tuUOCtpKeyHJWC/fhXJRUnsEasrw
ruT042PfisrNnJM/Hh29noLXnr+AzmLOEPNtJN76I6weMDCYZe+Af/zsIe07Mr8A
8T0rkN6tdoNTr2uCbyiVSlQPtJRPUoItHJyt3BR3TtqjN8aPDM/rhWkGgcoMR38/
PEeVCDeK1huW+fe7HJq+e+Cb0OG00iAC2h1rRC6nlnO4FJrRuQJqCn8bNbhtYRFN
y1Tu3rnLR0d7WxrZhnSkocHvBvHe4Pg9QxilDT94DiQca/0TEYlFLZLGd+xDsnx2
G/VUtxsGyIIZ1zlY4IvLt7C1+jnAdb67dycnEpqRgBaO9YdQUTST6aKIqyRo7zzq
aZb377nqo4rDcVFjY55nCyqpVz2oqHKBMSp+ourgV24y19yWe0Jh0903k54UPzhd
DXTw18nwHltoTxKdbd0G0zHWCa/U/YoDsm/aDJbcdZUzjq1v6DO0v1qj1ha0wBk6
2U1tOY6x19+DA4XS1iDW/TzOfTbgAckNNRBKch4OqtM1rlzG6vDkj0a5E6ptPawm
Wq8oN9Kq7pzFOxbI6uEDFjsyFFCAx4QEYgkDefnPbVoO535kWDbh9ZaWlVPr8X19
PuiY1mNZbUsWNF1KjjgGJBiVkcpVOQ+S3DCIntMvltgoN4gX2JXq8dhkH5/KQFDT
6dh6v8KDF/mjVErADhv4UozQFjw0WuwPAGCM6gwzI6caZzxwZj7ZLsV5VA9fW4Ga
ScsEF/b3HgwZPSj7mKeHsbF7qTD9S5uB+8twi5QiFBgwSwbLyXsdGL1fqlHNMg1W
5/Hd3xUfgqZvXGC7XLFfIJQwxhneg/g0geLfu8rLK9M2vX0CYLTJFsx4Xfi2HOYo
Ty4b5Mbd7QhLVbNP1yDnmUKe5QcJPUZZrvxQKjcSz2bVl9WtfGfp0V2flnpo+6WV
+NHprvQAeYi6xI1PXItGPD9d9id6Y4ndwSaU7JgIZot+bVl38Zs4eDlDKcwGbTbj
dzKwabeNyH9YJJUR2XCYLCQd42Mu8OyXUEwETcLE6D0AqStYboAUzp2ef+Gfz+w6
xmqhQipvkFO9ib2mqjD5HJLzy6UO6EQnF9tnuniie2K7C/q5R783UqIGdy//Pm6j
lq8eTzo9h4PztrJE9EgzUAGGby9BeoOQoIkNWr7MDFok9zAMPqGNLKpPEONS9m+0
d4HR1dDzJmP0JArGLq2tF5XPaiIE2ziCCaulyiMn8HhWwNt+fOnoUjlAbI0WF31s
t+pch9hTvKWWrelm9x54nOekipwZ7x81mB/FVNvUEsI6Zn8JTT1xUX3YY/jAN8w6
epCoiqbtjH19/DYQGpzuMq0u75VFi2McqTXu6wqfEHhdJP6A+fblVbtr2/aNdwvz
i3mAz9FlphjmCa06Bg/4Grq46C1uwuZv3bNoNf+QuKZ9ZVv31OtC2xQRf1BvEq76
j1pl4P/Pz3Ka6j3VVtAXoO/PLSx1PHReRS8nTCDh0+oKXZrW6bmi5kd685xSTKiD
k681CCKEm1k8mLJ+nahJMPVPQ5XgtXyUrt1C5JTQqJZkkYbpqMmMSOyhmUlbUaLK
u/xqcUgUUTw445ifvyfpWISjRi2XCwb2oMzkmTojr3vK/wi5KNiNtHPSENUIYdgN
ZP3QDmFHbmOLwr39fOA4aJoGCMl8QUMnqNa80N1ChqG2Iwui7hjvq+Ied4SvAmjp
ififauPAfF1leB3Q+LLfAvBSBDOKXJo9SXXWPM6bnrZsJ97UzMl0SJaA20Awo3Xs
rGfxfHThn4Alm3YRSr6VE5YpzKq15lmTEEjGuS+tcgvoEzzZLZjS+uC0QHOq5jWN
6z+BfFTOF0WTAO+DEua2k4fq06Zt/n5LokBK8sU02TcwasaLpcbhqxiREHWRWOlF
JDkFV9ljiw1ZbCcSTN/BQ72MGlSSfQc89fFrYa51oaKjNzBna+SEBxAAW1G8Uf+/
/LCjQcZAmpKbeQE1TD6oMkgNWSKDP083ZJLHfG5lZ6eU6moNVmlAnPgxEuL8jjMN
PJWqTN0WBlAMuVMWUFjdHuRwHlmtP7yNGzij2s/RDncn/5f8pipOgAMP04+wX1RW
EURbKTEFrIX0kTHC7+dzmgwwsFF5+/49/DdWQt1L80w1Sy42wii+HwizNZnEYklS
zTbPhZ1SzL5UVdENZSocOKqNK6pYngu9DEYGmDdo0MXFjoz8/pKooUjIa+zme3mP
emOURgZEQzwWeqkl6xWrVV46sW098huc0WCsJL50DBbzMQVnEz+/qIyd2GuyvHlS
WjHe8tfGH1IQcFsbuHn8UD3r7gtaQREQuCwTj5v0nzIx69vMyv5gMzMTF4nklvqJ
VHZFOAsKdjblJ6BveXJluPXFac9R+k9xQVQeUkQeW3r7mMZCIZQG0adYN2sIBFHD
BjEc4+zf6SESISweXnnRly+a5voxdccWeu626m0q6lfwSjah6MkFM3zRBNFWK+xD
OnBNgatUgsg9YGSJ5p9IwPWNQY17VDyzLsYjDU7gKNpaHFt9ZbKagRNxyp0nkm1m
KhDoY8HdH/mgjL+J23k72hhL8fX+GVqVHMmwl2vYXlz4cw986qBX9uop4LL69pes
OQjYtC0vldufWElLPKF9mOUZZpqn4ZO/hDf10deb2fwd7HgxowNhzoM095gvXgji
mBQbuzCyrL5c2H0prCs3WsGEvVRs032SpBenmamOVhyHuLvvHmZeQbsNhvF0M/o5
DlUYIK0WZNfhP4Hjs8RSOry6uRFVLP9rIx0ekYsoGXrfFBevo25fXeQast5k4se9
zNXUS/NSWVH4xsSk9moz6NG2xzlyqjc130LeYQCXyvAykkdpVh8iZxpX2yNefkR0
EKITKJKImAOo3Pw/sC6SC+M7F3r5AFQYFBFYQWYNhMuw7DpTy7EIFWL5SNNKibxK
2OjYwkE0eGb+xsNx0P0jbddOcKnATXpVT4frJdhaaotw4yXG+5AFUs9lbL6V+U1y
BMXMczdbz5oNkAUb8WGrYjUg7yWxvSjEYPtDgxpIuW0Q9iBcKDIOu90PCG3Ij/i1
53pg41Z/M50RYrNCblHBbRl8idABrxmUoUtwSaXQ7Uj/xu2x7eCeOVyIv9A5OrW6
ycghh3UuNSlt2DbcahPa6bHgpnnSWXXO3t0lKWqzcw6wLS8YZgeJvYkfKvHQHLW1
UaIyDbAVeMO1cp6eb3PBlsLI7MFJ4+56726n4Sb/zE4T1E9A4rTwP2MhB2ZYsYsF
a+GGnc7p6JDNgb846jQGRv9Q5XIhpf6EO9cIDwEipwUBcsZxZZvDt/82Z6OYH8BG
LLvM1HsO7MXm6W9Gk2McBiLKp1OWWQDVzKKGHMFDV97AXS+TGGzqZfx/TJ/uPoty
BPB9s6JbA/tTqKbHLIz61WHkjdWMM4h/P7bwzw8aL3/iQS1LCtXrHCjPteYgCNJH
vLEKSmpFR9wb/54fnVfg6PJuMPzgFzMoSBEDDvuvQtVK/ulei/oxjWdCoZ1V8kbb
E9l+qFHr5l5V55rYueGWTZfy2ou43UFWEMem4EIoqYPWjkbXhk22/SLG5v0WxCwX
Km8MCMOlzZyYmqpdEUKdgmQiVERnY90FNAIMLs0kmTrUQolepW+NPz+toLZcMVI5
rg9mbH8BnuTBTFDZ3ywfhM7HO7OBuzjLrZ7n5MmMXQ5tuLCXKHYoT0VE8CpV0YHr
4q0Et0uXHXJ+NetkBhG57J00Q0ZsCzIXY1jUc65UME9LU+ku3MyzMOT7HrjjRm5G
gIB2Umgyat+EqvKffL0AbC8yerT0OlnlmbqhsnVCX2YLpM1+aJgCSykTwIjMBBIb
GLQ1DfBszIYY+xw3SBPRYdnJ8JBuXFEe+kNQwBL+3DVIRSrVWi8I6RM5yTu8Z5Me
bJvGHOK/zAgmas0oxI+SW9gLNglDba9FKBM9kTbYBA1HMtwhzmOev1XP4JFsEzmO
CdmxqrJaibVOKwqA5Ih5nduGetQHQfjgWde577xrL9RP9vlsw7iyLeZegEXABzfD
mKQHNQcCkXR5Xn3mWBJmyU7JsLcuHvxIIj/MyX5gxthgzosq/PhkaZq6SHjhOFSQ
n9chnx5jlM/SQVg4v9Ercqv6GiILjFAng4pR2iAQ9srK0qBokOSARr0JngW54UFL
qG7Nh0paUNVQKgeBlqhCUj15pnVXBYXf3VPnQn0gqjKWYZreqdOj6UriffLvD4fA
ywF36zjIPVRn0sROyNXv5TvxOtQOTCCrIy++z/h4tmbABQZ9un+jME0pMxQF3XY/
0rz7jCj/X/7qyeydvnxp4RZAMjE6rBCirtnbYvXqojmWzovTDkDspG6mfKXBcs7B
6Yk4DT26CQRBICCQyVofPV6H0HDqIul/Szvf9sWBI6DHiNmLR4/HWnxeNqQBMohY
By/qaSGgm3EPgvaPIZX095DoqbXZ777ffU5cN3SbwLH2EzR7v7IN6nxIxjEU8UQZ
MPD8ujZo3RZWpjmP9WlXHHIkmLMrn9AhL1j15EQHXZr6opEhIjnbwPEAZqYDgeiZ
S4edANeCcsgHOx0w45jw/n0oGvkUIZTIoNaaRcL4nHeTF3d3+l0Cm0Q6JDnih+sZ
LG+6c/MqH3yBC31fEtR9eg==
`protect END_PROTECTED
