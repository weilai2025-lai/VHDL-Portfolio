`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sn4eWf+T2nJm3YMOUg1q1ICE1juZ3UjvNSfSnRhdmjeQu3WCo/0hjRhGcgG2Nxu+
6yQwFlMSWxQkJITK7K+gq1BYolYSuhJBhaHxx+a3YI3zZagW6/46Nhxbksecfz4j
zKLVWQ/MWvR2Bo/1jozEa5+3/QjB0zw7/bw+a6oGgvVCN3PajNSSqpXtRsRj7EVN
zQwK1CdIK97UM25O6FEJxdQCsyKMqqu8pXIfHzc+JdVj10F9pq3NgE4gBIKLQK2w
hpFco4JsJjKqu3z02Ctfd0THOvth4XgqfQOq1MKAosNm75M68jI8+6+S6egiENTg
kJo7LdPIuIT0BFX6ZRA4RIPl7o8lOe/E4wuJ+TIGafiEnS3xxmk/5iQa7+WFKFXT
wHIpJVi3e2UhjE9ABNH4xNl43VimzZSPyc+9qOmFRtLvYyX/S+pQx/8hUZJm1yDu
WxPSSJDtQqrhkqp07s6ST/WiGhoVIyvPqUB/ye+8JsOOedlTV0vb6HzTnyVhCRRR
RxIuQFLBrWBkiMy4rct/AcfE6TGYQaXfD3fFt5Un3yDhf8n4lFkVj3jPcpDd2Fpm
YgbqFgJW9FebkeZmLaN+kMOfe1xJza8/UV6byCYNV1YeaRUtYJPUrGbb2Y8d1L2E
Yl+f9gBAVa7PlPzkOM2fiwZJDCx+sog28KJprfMeJPK2OTzJLD09YavJrKb+90Ww
rT1+DB91kd/Qx6fiJ7RQaLS0xUNhaeIEGdqY7mIiodxzpT8QH/+WSu1YXSrj4S3O
WVyle81qAfK7+whadEPZMAi6Idr2fxUL2kKD41YXRgPqm3xDUe49dNlV4lhXUu+2
k+pO/FlXoyskcAbmH4VGuVcoteATwcWhaFz/QwqucmdlntCV19CUNSrttY8xfxLq
KngZMMcbIliANS8wAJoXLQXbBgsoQXUR9MVuAoYNEVoBOfb6bDk40EuFAUcl5ug+
sQGEthHRl8l1BifxLynXVVleBdnPAXoo5QRuufl5kV5z7zux5tjFdHGu6hqEzArL
Lu6VH6sg9WsWuPPvytsMcLJfa/iflCCfNf51HgYk1wn6/sIH8b6BjbRKLUpgIHMa
HmZNSBuduPfkN3wPrA5TnmqH0Wh4np6fPfaafA3G8mbvCt072nd9ik/W+qiunfd7
D9QaXPmRABsKYezSfeOVgQJDAqH4gGEHLnRRXVHPJGPc9tFaoVzMiF0ymE11y9Cp
LrWvUtryABPq7NC6xL6PM2mZ/iq3AvA9gMpho0WY164gvaP8VWmWed9Xd5wRjCss
QE6595YSvagLVchbuQxFe4mBuc9dQuhegoaPCwV0t70MeYD9bAQt3E5qp2VGPeZn
3wJUD2dk91/X9MaoKkVkeDkZ6VEoMYFlQ8qWwHdUmJ/bc7UlFPJWN/t18/N9o/no
1+GHGiNrkSkP/Fj8igV0fJ8EHxzx69l2Tf9LvEXLsd/fnHvO+oZuvKl7UpeCPVhJ
M25WprmCvcxteaLUBnZ5gVy7QlEQtSFFL4yKUxhVp+33kawtcpXMOXucTORMQhXx
LL3RpE4z41XZwSCFbfUFsu+Cwu1Yutip4JkzHqNZWknrP0L601jTAMIz3o2Sg8aJ
mPohvlpgEyrgyXsbQVmWhu+L/ho44KzzKsafseFPQvAzDEomn2YRPjaMS8XxXsot
Lk/DxJxoTmao0vKtezk686dso7aNwhDTSmtHcqmAdZT1jQZpo4bG1IhzvMATyhza
QDZVVYTvn8VZi431Y77UHgZa0+pcpuKPIkaHemqf48VTuDHvvgfX8YOT0xz9KDgB
BBOPzrDBNbseNv+JHYFVkuURuM5SzsFMstmGYsnP9Wjko1TdQnpV09cBZjvlb4un
VnBcADi8ce58goAmoax5xPm1SxdFZezXTCRltjPsUTqPhwFNPjzRLu66yGI1sMau
syu+sg3zvsmngm/+1HANQpBgk5WKaAhbtiQvDISTLmk/gqUPu8aWUobuT6Hlt8qR
5tfnHY4WsjrUo6uJ2bjCNNNp3XZVZgoZ6EBbWO9ybBz/hPJpDGOzjtI60ywoPdfW
8LMM+H0sxkTnDbMwkQTqYeUfztoh2VEZYD9yEHJXyiCn610WpaPdWASQ7EJnxYpz
SqfYkIoHANM8VGUYnGKrNjRca7nmGK0f5p8Wwfi2OMMAUvrAkrFxP6GufQ92mfEN
+vcpMVce67JBLlgdKmOJst0e185+ONDhNR62tDHU91VFiuEL7zUQlATKajRgeXtf
NqJ9yI7lgFR9sufooByZdegIPaS76kcAR5X8406VyX5IDuaYjwnNceqX6L+Rxg+2
AkZkBCKLHQxTCMERhDnN1bHB4FQXUwFU/2FwAk7UPDtVV0PHbloSIIJhdljJSfRi
+cmVN3w1AesYdH+NqMF3ojIRZwiMJ9+HFIBC0rCgL7t/Vh64N/kW9WC9B1M94WB8
/oeBX7nec1eEjvi4cerl4U1OE9Sn9Mogd8RdAdyuAUNxv7P5W56vG6L/PQag5IVa
1U5cVueK0rfldjwOxn9Y2ImPclB5QEjiR6XzzYy4W8t8ZvdIvZff+KGaC0hhZD+n
6LHFJP34k+6zgZKN/LfJgFvtl+S5UEeH1fBgrs5hBMzWVKiXbb/J8OkW+Mh2WpjI
+LmRtNfMQM1nBUSGUJqNh+iWgbrrzZyXitmO+KwZkKxUsQdYtmm7Ag7rnv9E6TgC
i9UyRD/S/ZTDanb0Y+EfgKXlZgBhHPlS2xRIB+eUSejTVcoO+J3np4zbMi4aacL3
v9yaMCWmZrpyf+forPN/DPpfINg4M6NTFwf+EAppCRXxRo+nrGtTA/43KQkWd87B
VY0OVjO6DBMSyE8PzRve9tLtiXkCnnOfNKXZ6614fBrrAqhKrE3XWYa6IkogNb/Z
CDbkCgbE8L8jdIC9yijZGOSF/gKw+WTgzE14y0gWcvn+mFPF/JxsckYLBr2eAFWr
qxVBgW1bt5rRE5eVy5a8BtqUZpfinSooPt0DOLnUuQ+v65PDQ4yYLutOV4vNKKyu
BNQRy+2NIJaq1pe3qy7USCMW/o0NxOdOVbwgg4dYbGXjGunimrDpVuLa7FaGbMny
psxjmF80bUtrzoLOQT1FUtDOwl8rRO6FkQP+YKo8GaVqRcBkrvS3YEujMTSe8HGV
yLrCaJ3MelVoU1MPNJyFXEkL1Ngzv7em68oC/+37uCOzUc+cAI6guDxv1v/7lrUG
5X+BDfVYDmUBmyAjIhekxPm9h9hlvISqO9SYxPlOpys2jZw9fAyEPRm20kSo//kn
WzaKxrCN8lCXehAfvDYe4NMla/arGejfWOwxA6iLbbQOqWm8kSoEhbEkNjYxprua
QSTY6oY3dYVr5aXrT1KaxMygTm6jmyYmdTjQh+LYjzEDYdtS3fHypAYbHYueRLbp
oXosiJLAxniQJusYtj1hCMdQZBTxkKChlmWEsMLi6oG5GAYOf2Xw5pn7R3xTOe44
REaZ3GsXsTrYa/ykXmCayLUQUYtu4PZ4//5V/45Li1QNLzEFxwEUmL9n8xhDD64D
0bTBu788kqDVkYt/qKNpvDFAjN6i71HvJ4vaEfAnfgwxJmfwxh36Ol9OAxhStNx5
0wCP+m6hAPRlEPzgkBV8ZvBp9I7AimW2SRM7hKX5EAlIcFKTrk2hkTTm+crurwCL
pu+GkkCu1am5Lrswuej3cw==
`protect END_PROTECTED
