`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
plIcXlYM5Vbtcflx+H71zFEsEum5xL9LUtIew64WHNsHgc7wsjcSpD8WECF4PB1b
aa7d4xIGO5cja7IipcMCoZwR3ELf1iuV6QAGN69u3J7hSzpZtWSFt0o4HNYBHtuL
mGRmpF4cWwQr8BbTg/l7qlfkSEovavl1MMqsF5gawoVvTyiEHKSIzMQ9aFPvWl4D
Is5sWREUhEv/hfd+zIamMDTcug2nHcitQ+mGCQXqCgq9ygj0vy74n5q1j6ZYJF9F
dl58/0GdXjDtgOXIQx0dWAF270BHZJFG/BKF8IErNKjsGDEI4D4jSHG1wfu2HoCi
UVDf6LsgcQSLS2sMwnKl2jze9yoGiJxZxeSGtXgdTzfrWJK9S6oLBmEUMeEyjHdf
9JL27e8Le3opCyGz0GzyZhYf/MXjv8Qm3nLMMjGqRHpmz8mJ5yxCiGcB3qN3bf8n
6lgjCE1t4j2wMrmtFiTqmJqt529mleRp1y6MGRqulCQ9PzcM8lPHo4XlCxCMMgA0
FwiPYM8lDAeEw8kyeJovFznyopaGW3PUBHIXUo1/ELt2jU1xMkquml+s0MGrY20+
HD479tfhr2mTZsAzzkJ2ZlfmJJKAVxmZYF2+RBYpOsDX+KWMxv/ee63fhrSehCL1
SnEHG4lukfslQQbegg2hk9nuIYzgJs6nEvBofQBXect6asSFg2RwZ66XkVONRHvl
9uz28u2Wm1z7kt5G+3ZlFCDS7oc6Nw11udirsZ4kGUVizktzeF55tADdT5EDex//
SNfJKmS3jBDCqdcp2JjCinIXwt7INn3azCFA2tbNqlV3R5/88vgiPo/GOi4+FvRa
wycKQXh8U/1RiGQnNG7f4hoZAYM+Jk3nIfHN7cQiZaHluc/xbuWp++LEbZ05l7Hy
lnu0DvBZ4SM88mNYHbdpLORlPHYX5ljl4leEOeM2QS4wjnhrrxZSZQfePN176cy8
mqsJjaKCSKEHvsgtyR4b6ZEoTXquj8AuRaL87kiENe+YoHS+gSwLEThe3mBs5yWF
NjGJ++KjovFHj8RLogX2s1Oi2UxxqqNA2EUfPZZFxz1YuFZJJ2N5E06okgJK3CBG
aIUxoEDvaR1FsMFve1+Gi+ZHsJYH0JnNK5t8Df6fAMkQFPcDn0cSKvytnSWiadXA
f5hMm2L9Qz1/RohwUbPv1jc1H+38mX8zZ1R+uhaN5d5YU14w+90wfFgth7LweCLE
AjHA8/07bhbTHjjoZDxVS/zs/DdTPri18LFGawfKdGgkLBE0blaDKpfzyELA1/F8
2CaT936nyGEHl8LInymY+tVEU/BOJqmlcUyMgth8SW2YCy60Q8HS9zVbSJ/vsLQM
teZkpQLW40OcJ9N4TlihcJrywf3zVTZ1g6ohL6dQbbiguDZQ2t3Or1mew0qlwLif
mjWcLFLcBV3fZ623DXwbXjWKfHjFep/aSyDblZ94rSw=
`protect END_PROTECTED
