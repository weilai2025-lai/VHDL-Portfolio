`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dchLyhzmHE2wfjSQbGGFKLEKsObJFiczYHlTOQd08ywU1VZXg5ySEfUBzyRGir2/
PX4vZKQKWD7NBKCDFGYIc146tz3hSljUJnlDb5qm86k/Chn48JwJf6BNxtwIAZRc
onYuGTsfcgw6XApQmow1qjiTtJQJVptvVhnXhERb8SPd1gtlpLm5HD23D7dLuvxx
ie3W+o0MuoxP9ihJ5easyx9/MDUc7ujTNR2841PY/IQZhguhwpv7EDDoEbjPmiMY
2dCxbv4OfCKJG0uf40DSFZts6f+RH3dk6JYOFhrU7+yRahHiL6tFjmL1yocKApR3
ydSIwktIltHpNxeXa2zVheUIOPuOgML1vGo91GPhAqvBoSFjUAs7Ofk4QxNBx6Fv
jRfz7PkP9UJnnjlX7SnLwK1NvF7KjRgk9vS9dmK+M2yiYch6CnItLbwKMfZDBD/+
Yg+MAD+lmbxJiy6yfUXNub/Pvc7gnE1ESXBnQO7XMWlBv+wZeBkoI2iIqyFc6BuX
XBWzAA3nDjVGMYPEu5j0gtpa9BCYt6tsR4FcgeKJiRgHzoBHpP2pcC8MvybdHdN1
fgXYJ6aOE0KTlXs/XGWJ5urHeN09lyWkTfD0u7FVT0cMebiMTPYg9kzveUxDCXhr
2FUwlI/375LxjOBPYOhTb7WLPA4jUYHRV//BH8Jka4PrUA9JPbOZnUMdfk+h/c9R
0xS2EN7DRwPKOlSsBBthmeTOB2VJ68aU5IqRswut1hY8IBRK/bhpg1OyOXd/Pmat
Z6VWrerI1QwYALthzd+t6EbchydO+QcXIXIsjznmINLaAioqppIetHCB710CnPRZ
M3+i2S3o5r3IaMymGkRg48DD2dPJudqJ0sViHId0GhWwjT6/ZwgnHmh57I3jNFj+
Mg7mrcmgQxRyRFA6lJLbNtY5POrpiC0jcBJxNdF3B/GYp7mFxNQD025BKuLq4fHb
xwpg2/v1hGNqmk31bcG2HNO+AtYfWXog2q072PzXJZOSfzDb9x0t1kU9pzpzuEJD
P/Ol+5P2RrCiPi3qMK6ualVqa6dp3Brnhbt+n29stfcfnLZ8INQczMXS/slK9GLD
B5loB2W/zNo0f+uKg46jmuWM/aqi4nyVhAKFuWrGnpWFszGYj8HkImfqQuamF+Tp
zl/cBOnzJBOE7pfweMGML810O8l+BnV74U+3Z36RKgM1msigMbhoGrowkPW+zZMX
LtZruPLqCVbvRXIFjGieAzMcXgnOON8EHVRludbzSZaTYhTZ1T7WtakR6GLEchWX
PAbWdnb5M+zoDHaGXzJG89Mm0Z6B+Q3oVHIg5eeuhSeeCUAuLp0oRrJA20OVafIe
EuWa+bKk4YIX6IM1Nc6gJEy9GdEtbriDq6CqCFJKzxLVkGEanBeoJuzbYDGQNHIf
jR0uE5VwROumTH0bq5GcSoyjy/92soqohXAAGeWJyAPEao88BwRwtV7LuTBiuUiI
vQKp74Ezs9VD9QW5n3MNaG8EGvrbFUD0CCkKuknfYQlC0XCePeHLhaG5dPBpOWku
bwaUTnEPgA/zEu4ENok0CvtRAsW+3CxtLiTKqZGu/zTtbcxq1BYgns36S0YpmeKn
89TauV6XUn63M95zW8ELOX+X9r5I1lCkutIgZDcxESsAjtvLJ7YriLdVTsudiPkA
welk8wNlU88qX8L5IFe0z4k92Ryf0rcBMds+RYRFWvPcLkLG576hAsICb/Qz4UMg
WgHwz2Zn0wPFzCZI1e7Q3Ra1bB3YufHg3MrxDDOKFBjBzpbmhJm7aGR3N3VJoWr1
n9FlbYC/nNxsAtf0edUKjz7LD3vWkKVDtWfVU5Wqo9DQw+sr4ARXwL+HsPxLE5Bu
spCDfoXKvSJD9hw/UW+nadniHdf8DledQcst+Z6BKVuzvnudSjtx5f/i/de7V9Ei
EbyFQKbXHiG4j0LTRww4vUmI2PX1jTYYpzY5DzgW4besECXS3Vtpx+p6eLmIACwM
mwNI4mviV0mjMkhPaieam8zhOK97wdpEIH0jKkSq3lxYTccmavPDeaK96LokTgEq
Zj5GjDH14TojwjutS+mz0ytYPNddeYg77ZaKWIHYJ90hUjjhQayPgozLBH1B0Edh
Pcs5NMTI2jkJ9gYgk4eyi9SBJyw4UkG78XmYWmW65drHpa0XHDPTYc2MJB2c+P6Y
ixLESHWY96k5tLyg24UtRh/pPeiN684XbUmgmS8WYXI97Md18GSWG2IdixShtcyd
sPGfi88SG3Tkzb+Mmli1mmu/8rvEDMfvO+hrlrA3DXp6c5o6YFlGCCqJlctLHGoL
oxMCXSRITf1mET/1Q4NwlOnqAEIfXfMzRiO1nLD9ydyAuPEc+oZwb5YQ1gzu7Ioq
zds8RwMXXpONhCc3VPucibG1YHN4Dr3U9116Kd+LDEocQH2RvNcacMtxFmFgxvEU
BZtZGAK/Orx73E/E9MQYmsYUkH9u+QzHS3cum646L/kXmzXbwu4SHiMABM3eAyhd
gWt/asQXX0rN+0IMkhXdCop1WP/f/vsJS3EAVv1c0h4UT7A5i7ygotb+gV5SEeiu
Z2c0R7GeGeYfgAwcQwo6iFQOzvFeEfY3JDMU/byV91xsmPcOeRWyFeqbeimdHlM1
Oi45tn80Qj+04qkV9T4Hh7qMQv5E4N83pH0W8DG6gh9i1MgnlzsY4zRbeo48kZOi
cxDVsw6gdq3rK66HFR4O4cJd+jQ/71Rpwo/Mjjr67NuKP4qYTMJXE3jbzp/xMDn6
wg+cKSKbZqdGNVmKHu0za6T/wz2vVe9AQbc/SJoKRnTZczd8kHFTwfZSEm7FJlv5
GhpYGheX7CWStbErxaITMKLyXO1N8wZ0TxbtzZwE+0XhAvWW1wwl2HR/Qn5vPA+X
VJuwYR2JyXg1EC1auDese5L/q+NjDB4ovOq8dPxtoJxSMqoFWq+TDjfO3kg5+XbD
oV9igdyRl+Xb/zcJ8qS9KzVpdu4Vj/L6V9PCbZa3UcnzGHCBC0QAZKiwTKEn4Np/
+f79mN+qApWIAKFKWRlwSu5Zu2WRJHkA7xQbBYLL115EJPmpHMm9Z8Ky53Rlo1uq
UmI1oIwnWOKEvwt9IuG9JsknI3Ik6Ec0kWLTsyMqnCK6xpeKECie/HkdO56FPyDU
c8hBo2T6oE2uHmwq+q0ezI0xw120tpYyXUJD8OatX/FvwS5rBb9RMO6rZy3QJq3h
n8CIzx+ICEKkgXVT2Vr/lTy1JGWmGi+hvPsyhRXtoiYXzjOPDld5Twuo4LvhttsN
N5MvKTJ+0yNL3zhqND/Ib2tZo3qrBaN4aNEp+iSzG7MwRGFjGZwqHJiNN7hBV8dy
e7JUt/w9EyocnhL63CU/PjCh0Gua+BA0+37HaCSDFsd9FUmYIH5J/YU613Exw76J
mNygt/LvhncSnRw9lMqVd0MworJ7JADwedyH25fqWSiRcjJ3wfhmOL3Qr8F3kWaB
wsqdHhNRf2XP7zRLK9LfDfkXTK1WozsUTxvfO3IaCzKgKm+DVHBXppx5grm1DLMM
r40mEe+9/J4t7vDK8CGw9xOkL60dNO1Jd7gX3w+p98IZKDmgK7LkNgoL5IQkCKqv
pMX+llbnzJ1gvAIY0uY9l1kuZVqr9Kl/pyi5MH9wwDwQQLuHtCtQSqkUzGGJ3ntY
hO8XPh4+m7srgDdzxsnjW/MXI8wTgg+heZuGJOD0FR2dpXST1UKdQ1AQAZpUCLNS
j3ezACa+G+j2gGCoB/+aqeHe5ZHXnJ/fGrasB/IeNfMsjOJ3uZskgm0MkbpSdb3s
SuKjMgJtUSx+estglfdAj6Oi70NgvyU00jwOCpfA98wIfZV0V4QY9P5/+3EX8ABI
3yvUOSnhquOSXaQFzQT+30sf8yP44K4ejgLhJfB+91IE/coC3ZoDEeEERJLIv8D6
NrClLFKNMbYFKcFpa5YPu+kAvv2N/ISYuZFJMieYzXksuNCSHXaqK0yUcrHs/Gmt
UARxI6xAUcGFqr5J6aaJ1XznAaf+6n8z1K+hhD2hF2Blevve+wMB2wU17zbuxLV4
eI+m8LV+CGYm/UFfk00Ar5kqhzwIUlT4yKFgnspfGo4J39SQvpEni+FeEzPqqHkv
6dP2BlLkWYjPb6awOFJnvx+6B99AKbflAcBEKshDuWN5/74RORTosvDDQtRf1eNw
fdcn1dI3GVkgBL6UtHBhCjH0D79towaFevk1trbRzwDVfLLqXdb7EPFlYip+rwui
SoPOUyVxW8imzf+K6ptJ7ueokHLcFSPk6zMAH32ZzblCyzS5eZ2iJpw23SmEwffu
EuwbYEvgRg6sQtDSUjSW64InO5zNPrQfrqBsC/eSBsbXaTktybGmFtHVs7vj0D8g
t0imgvTO+DfXmQ0xkOPWhT3MNAIZIzK6/guPvAyTq357VY9pTPZuihqasLBBx0bB
NVyphJjxDW1wPxP8zBa077IE7mqy1KJHZQKtCq2sLG2tvIM8BmEpvxLJaTyX5BA+
Sbm2bHBuJlntRQXVTy3TUrpSDVN+yNunwTx/6DYg185B06gq+UtYHKGipup3qnqj
j3coO2OUaq7AgQ8uj466o7FLSlyIbgnlw9pTSBULGn0uvsgS9T4MedewdbpNqkf4
6ngv0vOKxvvbw0QC5xkGtONfK0r8pdZAS7/q3jGbxesgq/LKpGo5ybzy2wU6G7ez
9DFuHST3a0Ta4o99Ig4xVaYPsIRrlKXqArYuNadKJ7q5WGn2tjGbpn+2XdGK9rv5
CleQVUojKRZ32QmhT+rFM6Ep8CCkymVU9R8DFokFPkZOpa26vVF2EYCqtGRk1evz
Ril1XgoP03FAdbhwdbK9zL2C1Y3w0ZI68z8GbsQwG7n4/OeA9GUDjZoFT8Sk2JQg
fkYaQP5ACzxNDfh4QhTU9TeGS/8yhvniQ7x0ahDyfbo2y1IQ4nuFyq5VtNlqzzWW
l3X/xObj/oc0g4yRJCiHPszXCF/y0oRHSp8mMwjD9QJM9fTJi2EW6jkDIy0GWaEq
1U9iDJzDiCs4KRXLmroLkIeCxtZ0yQ+NsFG7VRuVNXYeY8ZuhK+saIdUMpVOQ2Y7
E+PN1jXmDEtXHAAfLhU04bCmMF/RXcGJCs/749l0nXDW5ePL/334cNV9zUlTqrzM
8rdyrrR3PLMh2GaW1YZ6ZPfiUN2m9y7nIsF0PetJWmD1Dz+8cVezl4E60AmvGkUf
EGDk+C7nogwPEQqCWzscq/TSRVf6TwAmfawha62/gzReCJzIB8EWqjnZgmY8RxOy
usXzSv5xfQwDpRK14hI0WBP0B+DJhbipRB9UrB1oWFKseJs2hc7tQ2CMuwbXbT3g
`protect END_PROTECTED
