`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jam3UalKhOrL9/m4yy9qpEgqegH/lvechkpU0zOLdnptXeoOUmfN/P3W1TquApx
Mg6l6mqSmDcXItm5gpPPLmlsWLdYblkTiYj0hU3mOyfXnDOO9vKy93a2SlXny6bX
eKqrB9E3MgTpXMj6gatLSru6rszlrGZgBXJ3NbgUbYu9zoQwlnRBa7QjFaFPhq3g
2uRWYgLOVleXyeszWll+Zeb8tpyaoOnoSjX0peIiQirbkP4fvklH/x1n1Muo4Hjm
vgLRqzqCnm3e5YN1HihpWBHCx0iwRxVwhUdXh2iEuFsYYk1X91q+7IcjRGcp06uA
3b1zTxJcLUw/ji/tNMrnw5lS9m/NRyP+OOi8gPEInJiie3dGogVaQH2GAY6uxhkL
dUHVa2KU28OXHP++s+NNvwJ2cspUgwLdx2jgv2bgYNZP3BD/nL78+qGcykj3ODGi
2UmR8A0+uL8C6+37tsvkXAz0iOEndVzEwuyZ09RpginyGVbCElkRgfAZGNokYrPi
cHARnut2f0B5y7kQsvlho1W8PHdBCYZR8hoi501a7m+glrURuAm3UIr2taSM3sRB
sDibMZ+3Of2TxTo+WPQprLyzKv0EKmeAPo+SLhE9SuPNX9oP1hPuTS4z4Uy6X6wr
MKCmaHF/3VwsNxxmlV0pRr1OA8frD0F1CB0qUn3Ef74mgA1DuRM01EtBWqyloU0D
dxJxnuFfM0hadQvmfm73c/YZuH5d7XCWrmU3IfrwEq9KugWU0T9GZtkdy+5N+603
P2k0u4M3Z5oBsp9okIc7sQ0Caxqz5YXTSpLtsnnPYvnh+mG/r2aLCCEykI2Nr2TQ
fwYprKRvY8OJasAzqsInx/5EF5v/TuPcRtaXhKBIz/FFIvV5S70MZw/1WMIypoVC
m0MxfJ3O7OmgeYcdci3SUiJPKlRu0BysJtJ4n8rHAmR0oxEYnNnBb4fQeDXrpwbP
mugdnVo5xdnzeaQ5iius1JoustQKDNSQ+Qan5NuBLTjhEsKblxO795u7N9J0llWg
BLFkE2BnyPA28zFHGzNQItWkJNqmqBVcJJYYzYquc4TfJtcXweeV6ajVge6q8zfV
Dl32DW5IN1I5OlL2DOFqd5skWv8BBvJOf31Iv29EKMDaXG3GihsK2mqzF642hv1j
kbRkkca8yhnIOfs0U0KQs3qWzipIvv2Afj8n6lGrl7Y10C8rDcS/MCt8okouxJA1
D6hTMS4N2UQyhKeLTqjgVRCQACjG9kq4Ye1xKjA5uXI7zcIB5svDJLdIRPSXD8Tt
EmBrloTa5SxW8s9DvkooW3Xz9aY4ZJ2mGZI7r3KlW9N4HmIx5BbBdtDAe8fGVCX4
RArUAijk8fk69mcNFjE8GKzu23TLTyYQeZ5L0hr1eANweRJcHUS8gwpZhyckCHmA
IjoRud7xzNcnobxsRqzcb4CZpzN/vid0W6fRXok5FDw0ICsUXxNdnpYNZdjWxUG1
xf7IrDRjTWS3VqnDJqi7m16THUYXP9dhdWqlC9rdvfEgcS6jMfQyJHn5KLCTT5z9
+/xRfOPlJ/clYWzvql8xQCawFwleCf03rEjNKILSct37VT8xZQGt41GOCP2oDO1I
pwRHSoWhviWWNJo9A9vUEjN60Y/Ev+KJxp6try0c6jvZLN/qMU4RYsss0Ukjzf3U
EvWmLmx76HVH4gCnrg1QN61ZIZN1q+MM8DmU04hE0824jxqKf/BN+EOqRZpEFct3
y14FuosZbF1hrwfLF8LevgReOsjm778DSZPsjZ42CWgjuw3YIvivaeHZZA8PYYHt
+MCB5Mm+7tRvzso4tL8uYbvtCfqVyQBUS7ZlT27DExo22adRvRLE55wyQ4vx2zYT
Q9vGLn6YX/FaQhXJN3RpKIt5SB6MLEf2bkfi0D86VO1ZwCWYLGvuRTTzrIbNyukH
8X4DoIqZgWoPMhoKZAmnC/gwMZmlcPEtasWks3ryur2VtnQgfxTzzpmnpQN9WWz8
HgBlXI0fT/GqxukNRNkO/9o6sK850muhn13vSfd4CNJcm+s3viVfY63em7TXUTP6
wLnkhCZDBkigV29UucqdW0IKp+6to/LJC/QhwtUk25CquvZKuesRvZ8DqTQHt54B
oKHVJ4UsaemeXQJWkkPBVecp5IzyfANWVwx8jMOHLk8N0416zcCfcAMFL8hSdn4j
m1X0XhZSSHC/+3dh6h56KGgc6afHJ4vLKhZU/JCadX/1QDI/nccmYu/oEeOUjq8T
LvpltoGUjYCXDpR5lLBPPKgMvi5iyZ27dz8vXWx98OhdBC999tsI09e2KcZgJTfa
5io3krkK9QBSAt0kElx2CI+UOBa9Ao27AmfuMszhP6mUSnSBbRmj+q3qNw+trUPZ
TMC/Au39205XnvlWbnPqtBTvepLd7lOaxXJ9ydCPG7FTyQHtOJRY7NMp9f+7nb6C
qxFg+u6TALPoz85yZulOFvJ31wDNzWTuGdKGJw1ASEC5lsVFZH0Gzf7sxh56I5xv
Cg6lM8Sg08ofKQiIqaMCw5yP2//hC5kvFDfwiiIaS01UVxRde2TotIVfWS3zr/n/
XS4MgDhJgMvdAsOGy5A38C6bQabSsg5NTDeWYJBgpCgtu4BItGbyY+droH5sh5RV
wrdUjLiJJcppnrE8cgt/x79ik8kulDzkxOqMjrfA4l1SMAjyMRqTQdbA7Em5F9MI
OTJMTNvhrsONhyidcrvPQT11mtxNunClqYK/ZTx3GnZ4etrtSoc+fDKtLijXx/95
hVdpgVR1toOKptrZB/zylV6yX7FWJ3KF4+gFddF3nDjl22gSPoJEBIw95E0NOHTn
FpUup00HeuiHvP1YiElA5v4gCyMF7xijOq2PnlL6Plsb0HnRUUrNDUdX6sZzSeNd
9qyMkMuxStYvpa6DpTmotUdBpldQhW4C7WifkoG0yuYgrdNfXlIMhrc4sa8cE7QZ
xu4q3KxGc3KoLnyqJ6zG6iqTv/A+kNFQK/SmwrkcJNuKKdsqGmcQUypIhktObtFM
C48WstgtVIhFworThV5Ms4PAbKAIehf73GC/dIIPY2nybgKM1KkQq6m4VwQBeL2c
9wuMHlbxALR203BySbyC9bCpmxvGNOXn98iZlot+reOuiFmW6VmOzkAk/eTSlC53
ly0qIF9lQliIrxdX2Hdd6Q96yve7HTyYU120BQ+qsR8GBXMACU9pzvZewipV2f2+
9+xIcgkBRqVFI+okNvUQRMvxXlc6hdktwjtSJQzQ5RPKeO/UeCP5FwilyV7mkTFW
zb3ywQzTddcFVNo+kSD9ZOt8KWL5fn3NFyqnWHg+SzQ94aVE0045rEtSXLvmBq/5
Jjm2W9kQHJKcHdiBCTKVZ/o69qQU+Lh0CX1mcOaWHgfRkstbFnUyN2ok7F6LO4C7
YS4AwLDC9JZrCQYpdtmY4vSqjKb2/YiaCNBRoWJsG+yBBg5AtbGp+5hvw527wisT
clo2hMD1fKWQ5Aj/gqRWJAqykkzQ3odY5hLtkQaJkOB2kQVzVI47Za5LkevBcb4Z
S30VOWtqKMBgyfuEDcmK2XEufeWL+mlZYKa7aWutRXPShMmV1ay1/RLC6zTN+Ypp
pom5NTP0SsCQVQTYOW4EL/LDvEk55I8KjRS6XpveXH+9mkmRQGd8wu74aLDMZS4N
2rpHFexa90ppwcoo9QBqkWy2DELDuZm56ytdx0xJqzioLfgM7zJPQLK3AaVRm9qZ
/6ck5NbX2mCP3LejWdbl/Q==
`protect END_PROTECTED
