`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6yZN+mEqFWNLoYaHZWe0/gFeyzaDc/SVDxlpIvT6STUDDDBsTnWRGGw9QUkz+dWw
audnksiMTjgSBabZzqZUME+eUgKG85yw8nQNpWuNNXv7YH+jXcGOlMZtZ6m+SMmU
zzBgk8857fyEMWVcOKRoF1aqQvZZ10M7KNKirqsc1KPRRR+vBBZKE9IKxkwoLjyy
c25Ya64w6oDmM6WBISrxFGxKcOVaUThWRltVzSMvuOEGrAGfDc98mhyFLirdy7rM
W3FJAN7PAluskndAcvEQE5ZHL0fcoRLnxo1Rxsvsf2aOTvbynb5IO/ZOYai5IZom
VALhLfDwBAZAEu8q7YKETxoXz5q4W+DHLp99Zssvp9sIgIZjo283EJ7crc06/jAr
nw1FdtfAXyg3kFVxtAcqrWG7szYq3FI2hqWkghjjt+mXi9Spn/vXPoLaWKeabL36
BJ4DlInh5OXsKjGclAg7hVT6oGFkf6I2uv0WXckWLgzcM6bXqOgWIJiI3Vf0gQKs
Oa6EhuSKVr4cx5xG2pT34Kk8YoPq2k8BR9J6hzdHwuk3yzbxuoCfRIIfHl5iaxWn
tcSgbslR8fy4GvC7hLsG9eoM2BgVSZGlgVgHL8KyTMQVG3LGGInQET0zfT49rVI4
j/MWHv2eBZyTqEcacykGI20xTsm1Q9sKQ1Jgoiyx7hsRZgf4mIj4mlSLll3YjyTR
URw1dV6qzsCSBHVka9uG2f5prv4x0F8UpomgURx7jwrbHzguvgzaxFlKu0Jc41bY
RMwS3g2uxms6Ei74im55SQ==
`protect END_PROTECTED
