`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
deiMu27BZt4M/Yb8QGTTA/o3q3Qc/jbXUVQ5IFbuqfLqXxvq0HDdlQ4x80ZLBJp1
JOcP+M/wP9mLGhaIX5hLziG5U3xOjT66rwrOxzYmKtvuJdIWnTf7Tzq2e9Bx3LFy
u1ghNhQMK0m3RU0/9oZio8L9TEOd0Zh8SeKbSJuGxsDRPXplTb2S3y8ig1Y5ybVl
lThdkIkYyWIEErlwQsYNSyjGR5HExG2weS/NWLUEeCntX2i3rB16OA+tCmT+flEy
NFYcgeHESRhl0d7hdNfpxbgrcWOEJvkwJy85fUV3HoLnQdn1UZdP0D8/rBXqTTqF
uzxlJvF5MP6RTGmchHBBi/KA3mmveUYKxzke7bphpD12o9H/zzJU01NoLwq5tEoG
k3Xm7lV0HJWEUtIUYzIMHPOzXxxpbor9xWBtHdW2UONTYnuUQf+YCSgFc8oARH3H
pg+vGpSEAmRrbaknhM6wSa/+aoBSWQ+BW7rKzmA2zc9WJnM8w3URNXCmtufeS7T1
UNUOngAVoIpCrO+2SXwj/r25OWc508WQpeww3Za4q3stsHyvmAiJbj83rFURnXxL
hfGrznGpqLnXbtzuGE2Y2jKunpV330wxmxVqj+pdw13ZLZeZq/NSZjS9FWara2KO
l5zx/ZQOgFRQdGeymsoh1nCJMmjoB9wArg/BNVzJ7hWYDAE6auGOE7hrRRo7Dgb+
iyYES5qiWHjFMslOfybFTmDIFc1iYGc7w3H854jzZHJmsuYcYznR4Hh0AqNciDDp
JDNFE/YRHDSDSpbnefiptsoOSiT2H4FWGx4bvznEqYQfBoSOctcb8tJoB3Ol/zhZ
mJGG4wqTBA71KLLs+H4YvtifPaeiiVDBp8gNvMafzx9XNpxZAS5jvyiqDNgIBLKz
oKo5Jl4eQgPDXX3Y5lKMMjjmkDguiX4ldkj+qRdwjDmzOSeEnCHn35hgHAuCweXy
RKSPBXTdHTR57OXGvL3eqBxm6jajwdhDDj2TNIrPSqZv/CP639K3U1enp4Gr9ZYj
PkM5uyswW1N/6pGAjO7ZCtc4BhvLR5VzrNfL3H6WHFO8sE+lT5LPofKrrGcOZeFh
crYlsuRlPMS/7To3ka1PBHwzW/EejxwORsKSgFYyVaVfE3Y9yQsRfUiREh0Iz3ql
DNQAIP1Li/QgHHTq1fBm3Ejh48efsBqf/ETzgn+IjtM5LQscznskAz0R9wD5lBXY
qOmEwDKCvFsGLgI94Ed2np2+VjD8Lu0UcfXZKgOKvwnT+KNNis8dYuf9umO9Gx5s
gJ68bp2u3sauf/YU7UtoJNAGFixzbP1VXBjZUJ422OZoN+0MZ3jyb5pQ3EgUGaL9
p3i9dV+E9mO6QcTtKdFxQ3FfOK2ig2gvuQchfKi46AMBDO07OCmnrTxdDJU+m8aw
7CV4ovHtUdWKzppGkT9KH3sROyBBGNEfPQU1VtP12npzAEt+54DtfiYALexkD2Ln
AP97pCFDgfLFFwS/lDZDML/IL/4wLhctYDodtKNM0yq1tYL/dY2EvIpiWTGqJN9z
vu/MlkC7YJ6Cx2TCBZINRKPg92at9jv+36+twiLM5w8Xh7NVj8nkt1cUPraU0wlz
+HmfCHRlhb2pKZwhA4JxSvzJs/zpPOmaWyX0mef9wiXkZpWoVmk7eCM3wXp8mVMm
h/0RL+MmDme24SB6PfYmATDvNbwNyaH5Hr0vxan9sGyZ+Yj3Fq88+jsZcluFnseN
EK1loFWNOEvD1izzG0pNS0mbUtWz+Em8JEVsAA5sqJZ8EFp+AoVT8wSzzFkh6nG2
sSShqCMwHCl7EvNWpeEloRlKOgJ9y3tBzDYyfHFvFGdfBoF8B/bmm4RuYS64V4rQ
1/3NphrF8I8cMkpJsILJIO47xQfm7r3tcFaWMS2wG0SzB+Vm+rkO7VbqnPzcyfxA
Pk1Mh6Becw7xVWIBPCbte06nPONQNY41pDJk4Mm9bQcVDvsQ/P7HBKjgXfSp86EN
60RS0TxsplyA6+9LqNP3cK+2f2zJoXzLF7ApqAFoJUZFDfYolKOMBrh7ctLKhGue
M1DglizovUoolIZodV/ECDBOcbwWXAdlyytSb6OyGNGoGsiTbIymt5f4e5P/lMbY
QrLtwfolSPL5zOaP73Yn8fqMasbRVONIzl47mKGNnWIl3/WFwO3kenXTbxoecWW7
94itlwxjU+PotDdd7i7LHicye6iTqPNsjnibGnrzMZsp/W8T2Z8rYZ2taGRShNzO
s1TTWr37s2wrBV/8JX4bJR1Jz9pFM9QEs9XQ9wKfmj/jYUe0kEAGrlnjRaSnh8x9
5ZtTJr1CFyFYOT30417C9XKyObxmIv+6AFIa9UJAEjT9wUuQZYqJM8W7YJOhEUi7
q/Jke0Q5ahK089eRbZF6+06LrDsG9XmenvjvDc3mK8ImLp1UwMUbxbySo+zIb0Y+
pjBv8Hf0WAbRs8/n+vLORSoHIfy9rdThyrgUZesV8zINqt3e353I6jyxpfUASbnc
dmBO6P/MvrvFSOwapqzKu/4APmYeBuPbZawM6h3H9rFJTaQ4qmNKRp+6msyNoSTG
AHD9CRE3Lk4R47xSXJ+ThKFslFjGASLWd0sOT3eL66eSP6bJ28v957I0ELAp+Dlj
XNuHlDCJRX890UPt/FlCkUaOxsieeL1gMMdJMLwT8eM167fcvTm9mEvSxVuTvPhF
4lH8qPJKj6wj+RjRgTf+56sgn8n+wFNXhdgdznNBct9KCNCjBRHIlAflqy2XaCAx
g5CoEOla0JNsgzHYKlga3kRfiA7EDqmscz2I6pfmbUVmYKvqJU/8o86zIaXmJ5MS
nfr/wmbHozyeLih2FU/83/zhkf8J8kChx8TWsAWr7ODd7BCnnrEhtYpMc5szxpq7
xeMTLZWgdTQoVJ1KRIncF0h7T9rClDt6z74RvqxKRQ785aFFW3lGo1W766VzYPxw
VNYeXfm0LpDhhU4QJEW3MfgBQY243OPGeHbMbsOFzRsMJJrK2zFfO+xwjqY2juio
rT5PY3G4w251sma8zdlS8LCGAY4qrSKPQDCWjnMmRPhhw7Sxzq51iclDysnrBtjp
1O1R4ZKhqoOtegViM1Hsu2XmDL8yVCS5RGB1rgqoB6EdZShXGeqEQgXWZiSVZxEM
Si3G+uN4lQmJRpbydSAjibMfb5TB1lsYqhX9xqsTqRNMDCtRHRCRH+jNb6XGLb51
TTskwn9lcNzquiFSvSSACLlQg5grcnYglVChk/jeUc37sF+htnqpRWmnYqXB9CU6
bMZbGGDE5RAiO3Te1ry8JqjGi1WZv9k86CS7BVPfVSB5IHoJciQZeHYxmufdx5lq
P1wQEhFKSYO/+4gjGvKIvVdebsVAa95FdSMFaB/SUxpNIqg8twA6IqeTTvkNdzEG
gyte4AXMQjxt6l4IbjODl34eywC5hb2onh/+arZkj0GPDWeo6/uEcSmIguxyc+3Q
81Zox0L0AZYYeNHaU487ks8VMVzAwwHeLpOIJl8xIOAe5fe652PEq/suIPDOOA8/
fu16smT2HtGhhtxJHQT9TUi08aRN/lJ2k7/hhK2lnh/ZBjX1UyuWyFiiEpgZh118
tBd2i00aoEU3GZ0BUiCzyFm9GRjKfT3g/xe60zVe24t2bNZ+QE3QFc7kQyx8xNnV
oC7hQSldN/3PPvwQ59uZd1lRfM26et3gvC+HeMR+V4vfYu3jc3CPID3xL0ccCv+8
NJ4qzR01awGCjXW9bdsoqJ7lc0vMbPU/Fabqtz0xz6gapAt94Zsx0zXU7Ct2ihOh
axOYismdk1mkc0MCdCjkHt9/000J7NM/DKoQzoeKi1CBBrVFUJAJU/L1PCdZk17t
jYCopFyv5cR9LIpCGPGltAL/C2bPn4Pp9L9cIT6mIFSWo+ALE8Y1A04tldd8+DXk
cCmqlXFxfPVzHlO9Ense0BBn7E2vtd/w3vdkrk0ORyXQ9uJeUKlPP9i9CzLNuSW2
VtfAc6H7Tlj97rRSb9Ou5HNoSp3g05w02EGkEAMjA1gVVOKBEZrs/3pMNCosl4bw
OW4iCu+0w6uzH2qnywBoFvK+B5IzRdZquPsCC2g3BAbOjrAzjvN7s3O+ofpVzFmc
s9iADvEOFAnZPa5uFSytSHTyMbCFSfa1tKzbBCZHh1HP0Qk2gI2ij+XQW7UEhs0o
2EuINdbytwIy4rx9u4g0DDwgF68WNJpa8tt7liijGbewkFpsWqRZgy56qR+9H6wT
/2eHW1dziUsd8cQFh7YjlbjMgzeG9Biw8R+dljpJqj0yEaZAtVEBf9LY+24ouU5J
85DSeXgTbx44U4lm77SSK48vE10t1Ly9YCwtdEahcLFKHJ9qcNEHRQsLcMAlqbUl
r+UJGMRG3G6opk2ZPdDlbp0wps1AK6zPKS1Y1tnbI9qk6uJCYdzAdY0nMOkyRYSS
fvpocGwC13ekQq1QN0luRttCUisGv8rABPoSNrjkKLBXKujetY+nMu8i9j2Ge32T
V/j9YKYI0XSs3nzGI36Mlfa3VxyE+UWL4A7t6/32s1d3CEDYO0bxcyDYFW73CzuQ
GKrAumn0CLsA6lzeVGEq/aE1pQrStcULmKBreNcW+p35Jy9XMmYg3cn+mW8GoNTV
Mz2OMxkbzT3b8+8qE9CIBJ1ZCannbeeyyjVv8w2MqiUjSgYxY/2JMnZzxxToBYsI
FpEFvfhS02xI6nrUcVo2wRDT3ODNKvP0ZV2C5TF/VOJ2X2ne+yl2TwNGpa703uFk
EvapFxP+5TLHWDil0UFnf/C8c0FDhqcOI/n/5qgARVMLpy89c2pllAnimdD2pnmM
sYdjG1OM9rRYvBnHLcC5UxB7eAlVuICz6QrzwoO4YeQCzIR4Vodm6EzThXoQCVnM
5G9Y7mQsjL+h/b8YezeKowOTbqwp/IT32KHP7tqaMpuljzdNbz3ApVk+9DOHSBSz
4jAKpKrJTcqp4bo8nXbZrQNWA8d5L7yR3amuH3Pv0dQhvGebbeV2Yh5B9iiIcKDx
EtnQhcGiOiGGoX+ViBfZ/l1wwHv+pZl4jqrecOw0TdcBlFP1qtfbkulhAuaGwRd/
iLMv7vbnIgP65hE2N5ZoPzlNHHIhdI55ZPRtL/Zppo7IwYUu9OTMSX0OSIurCTbs
SEkAAVBz+NPA0c53R8nCSSfnWB+ZXpzQgy5A3hviBT1ZsVPLViPXbI0vH/47h3e/
xIB+FGiwN2JHA6dzimhU2uYXHvLmVjYjHrJLfbkNqYtQeLYCN0KFYJA8sI7PIPwr
q3P9d5RoIhAkg8F1vP0xBhGO98GMn6lyMl6RLvvZBYOiCKtAMb6vHN5FpEUwJH8V
Acc3x6dWt2XR4Y2zOPUeQhYf91++bq5Or0M/5vZ+yegIYdhLXKOw/2N4Ti0gIiQt
jrqDcfgw+pDAqoGUlFxRS3avfE4z2+TiqdTotOLUSxk/AOdruePu5WzdbQuMKCet
CCT9DKnGTYtZ/ZFGiyZtNn8/crlx3ArWRoXhvkcf8+FK90AdfO7T3MeEq4IC/Ak2
izuvo2b316ltB+vBuLkZea/Jku69bBn+6q2uIfvIaCHelIy0X6CfZ7qLbl1G8kZR
B8+sXa0w/viPF1+FtJ5Wf6vllB5rZwZAX0hRJdubSU/lIOF5qRywN2F08nd3m0WY
eZaVMh5palm54RtVaeZI4A5ccD9PmRLSGhYm0gOAkW7mh3mxEDQGwzy/XqmOslBs
WtRr5moFNEJ1muBaItYCJoDs4EefIz7kwfpakZSsjf/j243UKHXUt2rrXGhGTGHv
Z563pHoEuuoGthuv9F0xgWnj+WBLITU0hKtpREJuuV9Q8qKp/uq6OrKwbF1LfZWD
FCibx3t+QtrWHsh6nvpoMj8wlv4gKP3pkqatTFOsgBgvz1EbiX7kMNb8rTatWvVA
MYKd6sv+XYXREe2qHglFRJq6l7Cm6pI36ACG+uJpe8+OkKiYUrJK9VRqUheO9BXp
pmJDAagelkWwOU4ubDsEtU8gXvCVw/rhAADpi4EiMdVGg2tYrnczY3P+AXlgmUV+
jwN4B9ZenLZUpnnGrRTv0HavEGVcqaaiQZAUvKjQRJ1l0g006vVUQzHL+rH/WBKY
4GN6+p4Zzr9ZuYUnZ75TUteeL4+TCL+o/QdOVe8oHehHiY1gli17b4U8GtUjmCgu
lgSz93bIPpEOghoVhG1Rz613ydKern9r8sPUjWTlGkEnr1CTWdv9TA1cg1JRLVXw
Lx9JXOpxUEqLYRq8coUfYRNAvnZtDDf1f7wB0HF9Dnm6Od9nq3wTZG3SrbzIDtDQ
DA8Db+xw+24H1I+DuHOBZIM9MKtEMX8OqpiUphtlg74HAReQQwDWLwkJj8WMQ451
PDfOCMuZ7HcnY7ZsMA/XlylNPYQeJEL6Z/7eot4TA2zqL+NFabVSFNx/7TPIywIG
Rr3OaieFf+u3zl1maBLOzxP7G3KXInu+kmA21snLwROz4gnZkHFE3q/sVKS49+ht
eVLzXfzRirYMq1qINqKhknQYtD53Ht4rHfpnjDVEGwz7yvgei0nogojU/TSSOO05
+eiGs31uRiCwaUtgxK4K2gxeRTZHa0btpfQiqvL906YX7UqstdTtCkQ6992azOAt
uakS1gOE5UECCJ5mKE6LWWWXX63QOPyu7X8U1cM+lkU/dHArr/d3ELxrvST4PdnP
jjiNSPnxjO9qE2F2g7iOftn7Q0jdyPAz2IcYmxINPlvRwMuZIbIFw9C3bxQ07Oqi
D5Dfbr8c9+V7AD9BY2qsLnry/+NkqVeXDXbLnbYcUq8vLhvk6zjuhgrO3Cjg7G1J
Yl1sgddg7J4YN8UhlOmG6brrj1VNmtLo7aOAEKONvnCcT0CE0c4x9//uer4DKKKQ
tjbkl4PrlAHI75mcY4FwEJoe7s57LWu1yCPcCte4V8Utb3vzaKD9NGBDHjK6y/AP
XIxQuIkHH5cLz25PCNH3xnpmjXPfjXNwu09npFNE/Ka1VI7vZMjsWQZRNuEqA4KQ
sOZhj6H4wVpI/NwAilNlkXBEIB2q9a1wtAsl+H/+sw/euvksBYaGwAQZx9fFcGKB
GRSQfNPnnPSLCtbHg6bawzSE8bXkPjxGPhMGksfx1M/hT6/aRccfWPt8H3fwz5TW
ciLY2PyeCmPSLTpLo9RJZWAuknmdmeefLaANt6e/5oqrrshu6/IoxM2eOutf7NQf
TkH9vxAAgHlXiGgzeREAACwI6rz8KQL1M+BmWxA5gnWQT7Wn2UqOWwRtgntKGQDH
k0IPZVG6AqlHc/P+rJ2O4+4WEJS5bF7PaIoAb0kc3obrL7uhzBKelzjnZnbmFg4n
/vsXwgf3nr/k/HTfEUcheaavHJPr/EIffiXtgsCFH/5OUKEmvkNRoRnmexpqyoWY
Sipgj72RlnPisMAmOsPzaCmjPn4pTphEkxVzY3DUA4t02tHfBe5ThSKGxUsXs+Qm
Akc94nYZFeqXMKHJ9ytpRTl90DiUveKhCWLmnIkSoL8sKxIVTdchgipynskPCCDz
jjaA0HLTbfUS7Ygm1v96KP0XhNPBqZ9EeT3tSkHq8VJo8KQIhqQll8ekmktmFpFN
Ebkcv+thpZMct4R4kf13YSLtgp9lao7Ob8Qfx4BFFuGHBbG5Z2RRuz5zTNXSrmCL
7Tgda6/xpaWSUktPi0a1BhruHc1BN5hnpY5c1HLETuZvs8yXAvCz8xxBvxaBZNWf
fN+b8sHeQAo3SQgkfBQkussD1lrTzZa3zv9dMmP8vdp6PAv8ZcwTBTKkwTr1s7mT
cPXR51ZpIn0mcAmjDUxl2FHngV1/i9gmXw2BlRpAifQ6X3eTPtqdSo0L/6lJeVv/
ITtjPGfVF/azbAFZyDFsYh8VDi0iFDXFAHAjYyizWVpPoPImuU5Cc7lB3cEhpwIJ
Y6rXm0+kthlHRO8QOcsCO4IToWuA3250V5+NihxsXu2rgrTcer9DxtRYAhtcDqlX
mk8MF1KY7GNH/Q8cHEfuEcLIa5td92M6IxLsPOGJ+zyMNCI6tHy/kQ27B0h11Je0
gCZiw3YZkf0SBFRbHAVQ9qverHabZFjzZ1NgHH4EzdACSaEx0ub0cRgH2g8bbiXT
lM/aCAE254x3yiKnM60H7e3bJWiztoLEgYriQWav1z2mZGD0efrEPapUZYmL7bV/
h+ShK0UQoDHg/W4Tvv6uGDk9+T+HpA9e9p9Ar/ylKg9EkZI/X19/7KraIghc6eJ5
WhWDeqCYRBtFCexkmeTixE0byd4YTcTpkFmG+1m82I1pIbJk/BzBEOzpiF18gWpI
/m0SVMoxd11uFEmvpGUTCqDRjV5NYAJDybeqw1C0h0JPMWRLM9JZe3rKkJXA5sh7
1t1QWTnwgrp0KW/Sp1AysxLXRnRqb5V/pZ/4+dO75G1zaYo2a9Z0xkLamajqPni9
/nccCYvx+igS9VZsiY//a9w8qDmvvMz2XCx8vKJ8YUJhXapd3v4XOrbnjDwsrJDO
nWE0cPe5KPox6ZbFlstrnhtM3LPLHI3sQZnTHARXCdykKDduCaIyKxxjgRms/HBp
yLCUv0jvc4w/iDv82C5/JF8c2dNA1y4PxyvTOYSEvIozbfSiW87frRh8LoALTqVt
DdlVt/vNhR4m4/6lRzG8xp+sspTmCYcRNCacNfOToxdF7LKRqxbJ1DM0+vtAbifU
fL65DsiEayl48Ed6+gSnQRr6CqFogGYrw/AfI2lTymxNqkcNwl3KaISIhWzNcUfT
QU9o1SgY3EVhOszsYUpH1gIYEVqF+w4xvg+eVuJAYm+d+hhcVuMudhavi2Hkc3u+
eEYC30Qf4yHqa1n1ThIxZbHVqv3ct8YCYXvt5K/Av3cMwE3y9CYWjJFdSohuXgL/
RaMYakqAswkWugj7ryaMaYkburhFY72UHA6mfkwgYIyX2oosb2K3dzhuTXjFE/dF
0I5siBEfmxT9JbujrMBr5tIq8os9cXgdxaCovBGpcpj49VGRSxcgNLHpNmUHBLrf
Vmb5S+kYOem/FqXzLsdaEmufOX96B7Zr6dxZQPq8dwj2hKQEgxwiT6qZSOI4OW49
swH3IIeI81xejM7tlRdrGvK+4iqrfcLpOJJtrBXwhUjYeB34f4O6gleXoo61W9/E
3mJDtNDaOSRubmK+CW6MXvCLqN+DIWIB7ZA1j/Hrra7APDPLPKU/E6cERy43k5tY
hbcXdlBAtuwLhs9xTV5bu6uNDOTEvwfspRau1l/qixaxPgx/Aag6FrtYZaqU11ys
6zQ827/rYyQlmcqBTiRDrIPa0RBbztWOEu5RFbbF32RVw57/fJmSTUhAXo+FLjF8
5tYJ+wY1fYZdmW1995oin7qyefBPJhoMidz7tno222CrwTX2KM72xhkdLW3BTOef
wh5lEjZGDgJYHkA38Vv4YTJtnkS9ityqsmC++Nn3fbcY4P0eOlXVpQ8ycvPPRgrA
2xcX0ZD735Df4vc9Wgg8zKKWB35f3y76cuHlAGswEuSQ6IkvmoboLJd5xT0SIp+K
xvp23SEB6pU21txn3pImq0wI3EeDqdYU3IykvMvIb+FSRWFLWijxs9jOXwMGpbSb
BfZyOfi75208hA+1hqv+cKqVjl4ksXaiMSH4BHilMiyHCMd201YLN9NZfp/n9+jk
2cZgeN78785aNi9Pe0m3BlV/fVZywbz8NG0sZ21VZ7DjtLsfjkm1VGweOSrla9Aw
cM0cpFUBio4In92xz0s8ayv2+nGYlqzn3TMPMGyjD+HKq0v833tD66CKLYbzyBne
cZmeOLYAF+GyV5UepSowSCzeQh1ncT9/PPEfEUliZKTnG+cDdwuq0bdcGLd4Ej1o
zDBJwKkLnO2gRJUGHRmvr9/tB2+6xv+o/hXiPug3m64Cjg72DrXUhohFopcI3OHr
6bONbWmFHXU8huUZLIOsNikWOt3CDmKt+P3X7O+9SN5V+s10/vW+6GFeF46skTTm
fIfrOMBGLi9FW8x/1wAMfzESjz1T8dmrHDQstpj3MvLkHahZjPKSZ3a3dqjGnMRb
yl7kdU6iWRiLB0N9SxTi/EgH+Oo/BVgjmblJn+WzVm6MaAJ1uVoJQSZONFo/ydLP
Nl3xJpDB22IyGOMxk9JGc0g4h4a3yy1slTXEZpU7gUB/W8e8fncDVksL9r4JDZ/k
NwJyBYywngiCFe6UilC57RFqXPoagEx0y0iAg7WS3ta467CoboZAdu44N/dRAaja
9fWPq+N0NciY7gBNjtEoaklX60uwkP+4SNOaiyIHjjlAjh0hqpZKdstiR2FvmVQa
XOtglqSPOWjERIxfAlWJGkB0E0EwNN0jE2LtrjddZ3lmquGI3ouUzSo5EPnv+JWc
J6Ney/Pvx6rp5m9lQqOVeOdxMucFlqn9Bia7mUASBXmbeC0NlvLiPhEGktMDs3JM
EbcQdVUYgyP+o/p5Y45A9+FUbkLTgRiSkLtaMBqBjgYaOS0PybAM/uk4JeJ6pOAk
wNGTexcwDK39yw+KBrRfleV4zS9XSNVKtD3cnYqVzx8nXfxko0QNuK2NMt/RFz8U
SDTsdVEV/57NuwmCMVmj1zJ+7ozXMOZE0K8atejafMioftWp6SfGp8wBriUKEyzg
G16K/V0umemaB1VjHNhFUrONwBZGuupeO8IBW84GN4FoZ8d1sQDu1z6wRtEMNfka
fz3vq6fQAFzHgaoXfUJDfuO+izuwh5Q8oyeOhc8FBHYLejHTJOM7eyYW8WiMiaUU
pON8acXKt7/sxpgDl0BSmxlr6QvZQ0LEJRj/OlGiUssa5leDOHpgkVmAvcEY63tr
Vt+tCyAC/dl8rTwyWL7YaH4jA8cwkxbGCW4Edwp8k0f4GadMWkM40qF0mv535oSY
a2Bc1XmqnP2aT5apb/bEgjneog8I13wi8Hzx+Bm2CtVHOWGpw1E6BcOUPWIoO0J8
oF4TUw+2guK7FA9bA4y++VTkkI6PZhd7jSfH+QiRs9dN+caEU4BLKKFCqjYKsKh9
e6CXOH86WvG7Tz8PoxdDOFEg3T5VIb0mdypKVCXU0KQH4XdWxAnD6v39EzAcB/St
URn16p/mEIPzStMe4WlVNIgshobJQL3LPjDsw8bPsZpByt254o4V4pdQyGx8v9E0
9P/kBPV5J8kz41pRdMtCLOfP+1VdQhqIzVzsu1tGR37hjr2Lrz9li4JjnPTRvW89
3ejlrF50QelRS3DOSOjGWvAwvXGk38bGv76igMtbCEZGB802e94q7041Vnj32nEB
U3SgPhr7+XPGAZ9c8BhwO+QUFTQtwgM145jjBViO0SDb4eVkhWI2LTVPfOUV79Fa
nN8SsgnnJlpuwA9BhoaxZDLd1vAeeA61pbvXxzg3GJbLshCLXz9fMpwANr+QAJZo
x0sJBNya1/doxKrM45ki4uinFKkhpS0X9DYef+R09xev162DY90pxArWWjsmrZu+
iZbnDk6t3eb9qiB8kzXa3Bd/dCDNZS8IusNufNQM5esI7SHgR6YVg/rm/LHusQcu
fzd4yjwE8tpby2f26KPTBBjWUeTxx5Qd62Akeyn/6CXEAuojdxraqDtM6O0T39YG
gwomnTOZTHC8d3k0bM3sZCeMxNp7oFKum2v5O+Ln6Fa/EfKGvlAGJhOLHfDiIHCT
CvhcsHaCC+jOjIq3shu3Y5k4wKfufO+mMVXVYKHYbYmZVwbNEoVztvsHWnzwLtCf
oK8QHZ7S00pjwgsvPpH3Kx4C62RX/I3ABQyen5fyiwaZdWdicvZLgbNR1zNkZ9YN
dwIOzVMJcoUz3+kOEwEIWYV6IcpggcI0y9J+CQmfeOB2KEfXgUMDKVNeTUANaH1F
MYl7GPGKH5XE4U7tglCt0VfuKE2SWc50ueVZ5Cr07Q+1FxWb0bvRR0jEX/WJH5jd
sGbLQkCgTg3Iw8ajSBFX8PTqXc/j15qeYc4I5L53PoHk1BuZ3/LbdH6m/mgV/GB3
IUxoDlkTvARMJThBTShRyRk1IOyrdzdQX4p1wB4xHmlC2Ct0vn4JeyVRecuvTN2b
cbMmFRM60qFbqkfWD6TTKA91E5pjNooI7FDx/JsWNiAn75p1K5KYW+4mXcR1+7As
zThZq30ycmYCUdQxLkOEnxo/Tw9aw0AKopmp+Is5O6t3knmSogJlmOPgLBNGDX/G
m3RsHY24yoHvvlLbUg7FydNbK2/16pNM34mUobxk6jk/ZvAu9p1V/SSHUm3YTpZT
A7KMPzE0gjTh9KN9xswjmpJOd2VZA+Zra/xd0FaHmnFHlTD7MClEBKs63rjRw0zC
R25xCtd/S2imyi20EueE+lNiaAg+X+smMR+anamm8mJ4vf0xlP21FnZ8oAniiKoD
NrazgxbWhBs0GWf9sRdU2AedpTjwTKXpm39/RNmIn81fvJE99rcioDEKQdTM/POO
wym/J5ufS3VBhDC2YULvpxRPkJaC3lab8eMnW2nbfTo64rwOLLUIZj57hXgE+nRq
TSbH4l1zKYzcfCOu/Q0Q1YS7p1uOS81z7hBFzrGtEFZQ4Mn4wMq8WuLfnj/5e5bR
hHNpA4OWibf3zv9C52XQHIqcl0Nkjz5PWq2pL4OJbU4RqYSPBP2mpZVeDQBk9CKA
RWISfqpKNtXHZEcGedjGGQ2A+S87QL92HSDyCwNTJM52bffRozjO1QGL27FEob1V
YkFncPeoTOWVIHXMkwprRZgPPEZqeVqe3ANDepDytVRBYi6c59gNfgGugmU4Vdvq
DmRy4LgwJblDqzjZgp8HmS4maVZkrJCtB+r5cReYDWEys5GtkCG8TQS0xciw2ADN
UrWpGBZkREibf7SesIOFNDpgJQkaL9TsDyPIdz7+pL6iLVERvFBdpdLRgisFgROb
Oi5Y3yCIFQOZ/3fEtnfBCU1wyWW4PyJ/QrW5cOKk+N9eSKqydqpdHVPdUfpVDktt
Xj1Qvb69fpkGknVuYfGfgmPbRq1RnHIFxHZyN4CXu9yhubmkfYFlCux+ESDcMUxt
EUd8THiUEmbyqJ8pT65G8rvRG1IIJvRDZsiq9ykPpg5Tfym4MbNR2bsqIe1NcAln
NfjEBnpVlF2tYNaunb4qK25ysmcn1IKOn8FvcVgSsTijhExDqdJDFiz3BLef2rZT
dDFJWE4JAPifjq49WQiKYE3ouPLyKq0bOyKuc0/HKnj149wq5vUCZMO84YanPJHs
ykIdO1zPKYVHhiYEhvFKiSPjUo3UODo2sEjwOiO4ZEU1SDetlGKUKEmS9lIBcCIl
67aWSZIkNljEkx+69gIMqP4Blp7v1ryH0KW0xgboaW5a0T1PcItlXJH6RAA7bUaH
PEIDs7JcdtdTdiIRef1ZOG3knhfLzIBvyFKSh56HF0ungS9p4jv1FwCxwsdtrxLg
71ojouDlNs2iW+B74vHF0i+ORZFhPeLrqqwerlgMRyvrmkMNGeRu5UDFFZfOM07I
/0hPTE+B7H9jYIJxFBNiHnxzaACVbufl6uU+AK5XchTlRgMFjEYJavgXjpyKR+Qk
3z1Z1IwWAWGY0etg6II4h7DBVhY6LfwidMH+CaHZ3UiuNWGHiFFNWcHILBVtT3z2
9YOnJ9kOgGRtSw7A9JkZHYAXMgaXtafFfN3HXO1qsA1DQll1YQw/F0YcBGzDhYtO
jCn89c2b24XtMJFA4PHAL1Ztk0GokDb5BKQIJHCbcFBAI2XvDxS4JOc77X0euMIs
n7Y28cbjxjC1TY9XR72uJTirzmeBQbtZJFrMZM35UcNm2/yqmOnOAQLajE2pY+pT
W5r5fYFyf1/60TYfCDX9uv5qnNieslrEYBzs2WqWGCy0qeSvFYyYNmfqMO6KIk7J
PYSg3G6R2W5UZg4nQPD1h9na3MhJOxn2b8PLaMPx25NdKsoIPymqT1ObCjTi0uE4
C+yAETbsa02L8lw9YP9O2vYVlBDRAq6Jtbqy8KwQVWRKzmYalqjH+uaHP/7UpUHN
43CxEhGFVX0wzKBzwHFJrtyDpNzZH55f1O4AZfPEOj6c+Tbmg8JAu1Cu847/k6fJ
8n4236nwXL0357TEyazJHATC7SV6iubKCcnBbjX1W2Kd/OFADFSrxwbsxedve7Sw
FKQKZAxSy4dN+gWn3yaiNtmdOQaV2I1port6o2tSM/TkH72qH4y+2rg3zjwSy7VF
HjoCkBRYvGaVruP34WopcB/cvYIRUbrVpOnSLMUokKT+b4rhEcw8iNmHcNaj8glS
R8+W41arJKzwkkE2SbYKErE5YRmZhsltAIW3bvO5Visnvy7/CUhc8uwkHn0leLEx
9XobPFLKCvCQgyIURxSwynKDX9oYRK6mkQy+oZYlISNB2pK4lKkOOuVVGdMakRDO
2euhcfEcaZLJG1tZz/vp6msrHWbqy2fivPkbvcXtzti/QyLtjgWsn20OzQAUR/1N
uxIzvCWxCHkhHJvxsyCw7t2QJKswXnu7eJfcRZyrjPR+XlAX4jHCld0HNnVM5wrP
jmHAha1LFXduskUUtTOvrBoDSmM7KmgAanVrseujswCBtDigVWGPuS/IP6DL3/fd
I6JkPmEzSMnb8gHz5MMtZ5AOfkoOVW2oss58HEoN9BXSvpNo6VFUYXRyLruNwk33
ZwWKS9u7P8FVdQ7gMXfpGcD8wPFiwloJFSjo6pjqHpNBiEmTGh6RRQTp0pyX5IUk
x76j1IBcPtz636SzUXbseaUdOEbrRG/GTuhW+fq5bNGoc+QH37NCnoPiv6TIvOTg
fCQ0ST44u0xMvqZnFlPvr6ZrnkVWa/tDRTZXFUS7J4FPHC8IaH5LMxqHC3s0eTzI
eSlHmrt4xtvHoQX7d+FWn6C/AK170eC2O2zpcXLT0jUa23384wQE2Rpmcz7wV09T
O3B6g0KoOeGlDxfNJX78zjq2zFqa05Un3dLThDG8zyu9Grc80kn/HfCdyr1tumpw
HBPVvfWBBLmUrF7AYm2414w4ds1V1jPjpZWUL09M3Om9dbqvD3EvRrsAEG7486cw
eb8D/Iq6zQFPHsQDjBN2UX2PWlI+j83R9jrNPJaPYmIR2Z+HzT8qXgD6kpmJFpP4
2lYtWfdraQa4+2YovtAVfBtZ87qhqjM/YUsb7WZqA/LSdVZrE4LkuejOuLR7r0D1
N3LJ3g9kLN91v/zPiRxBQRhqpVGgNLAy52clmLxsKiEvdqZuXgXXgvpOsDVRtSAT
yOMk4pTIzf3neBlpuTl8P6b/Vs7VNfZ4XLKWfxGpi6tvSDqZJZJTVNzByT2YIASR
kd1kLdqAj0K6HwJskIqdE3kcMhQ4uxEzH9Z2VIosgWA/pWLvPhaRKrrlbeFm1O/X
HfEFNpDFGCaFnwD+zxmMLJKA1DTBKrpX3ejY8RJUqd0CPgN1OKDYLCYGKr27iEhH
ejx9SZuq0aTsKeWVBw6pinN3OJfugC1YTeSADpQjI6kxvcrFPCr+OniXK/CF5aJm
4X+9WySfWWH1Ys5qI/wsUCcaR+L6LZlfyQHF475F6RkCBuspcWYgHMWGH9AvPoNv
BJTlmMrM7BOqyxdg9RalEgnd7GgllCWst3hSMrRsu172NL0TdFDyIjdlunbrx5qG
0fy3L+dnCEyp6Zqmle9DEAV2hR2sw1p0prLba8+JoMh1Hi8OO8rwEIpM5hhGl05T
s97kTBtkdV7lqkt/opNLi4EZgO80MySk0BWjzCLDbV13yj4FOJvm+1djx66rtmJ5
zgDTXnuTMgd2yiPAs3gz2p2d4FwewhoR5meVKj6wv35VcN/vvDjiw0sTflaWw/QS
pRpb3vlq6YUq5xyOdyetiOkGemRHOsgqX5gTmJGncN1YjSQnFsQnPE6WhUhg9ba1
XtxrRjV/WQ9ZFsCiz4OZxAdLRuAOetiBgbY0j1PhFKU7nWTwNDKMj6Wyd4CvPGLn
s7Icg1DHXo4ZRqi4whde1PnjMg/ZTjnFCoQqfqjlhE+zv6/2jR59jN+sy4eVOsh/
SHdMExH9pCGv3BXAyffOJ3NqwfMEaETc8PgxJKpoyQXuMmka6lcH63tQjgrnlYYG
OvXDXe5dTijpwPh0g47DikitYtFgdhWRW9pIN1Ej2qlqS/vw5nIMq97YYSypmKec
M8YKsMnjbRUf1ak+Abb40nV5fDhDeccCJvvyeiyvnwiHypkAJmZTKqgBo9srReAc
C65SYoBPSqV0JLQeqMZyhhb+Gf2tB2+JtxsL/hTMP/kl5l97IL0n0F3dCzaFZ3wF
NtnGZIXiIXQb/SI/WR960JaV7fgMTi6F4m1rJAI7t64fMxTc4czVcB7alulUgO1V
CpCaWDUq+VzC+Gdz144AvwPLzH0BHZsJ7YMAcpkkb1Wev7SODKAOWbYEn2WNfyMC
Wiq/puQmwkYFrjrTpJt5iVl7cC4VHhqOnrourXcBsa2VDuKXjUi5RS+6F/9pRLMF
1BEJ4qrPr7+RjaaMy8HpRsg2A9i/D8clWLrU8iIbRJCG/ApUtsxwLUz4/FmvmK4+
r7JrY9G1huItxtboR6fCLucMnG1h01vtia157zbLILzQKRXf256ePnr+RlZjkAR9
Y89iG6BC6QoeCMXFt1LIK1upOGruhygFntIQczM4bLuT8AQDkSd6D71+4WnUTCg0
vrcrOYs5Qql8EfpUbK7P+IZ3OoEN8u+EZqzQFVdEpEChd0Mdbr9jHFK1TmS4EC5q
N8guJ4LjEk6sgfK+d82InWuLTlHU3PFAteR5Ew0RsM/2ve67A6rkaCL8snWDjRfb
/beT1BDiQoWsAcI8DBNHO6+/jEiLcNOOjUNDiGyyYQ21kVcVOVCtP8IG//E9Ew8r
4Gtc3BjfEqgyish4mnmtqXjTn7KT61DHac0M/UiuKyanmd2bllsKjhh3JC1zuHAr
/F4FGo/bFeu7GWStMLVPaGwZlVXM9OZ71mDFFScrA1a/88N6Tz3Pkf5pZLlx02RS
IDTpQOZj1bOBxJHPgIZ/5OqKufocZ91QXw4OIQiStnIK8rPZ4LXd4e36Nny1vSQp
vfm06q9rBL79J4XMgMnSa1p93p0y8BqkFOgdju+AZBydDjY63jZTwqw8iaJ7K4Xj
IYP0giWziezUvGBNNwQx5X+nTey6DB6skISX48CLJ0Uali1E4R2fVElRXj9IIpKy
T3kE/4OBNSBp1PBnhP9dKQU3Yz0Snyg20H8zukEdaf2qh3FK/EXqQA8B/CBn3fCa
r7/wnBwKfw2SG8Br2lt+QQq6sQozsWkYY/NvIP3MU1/TRJhNYVEe+qBHAfUdsu4v
WNFM8hOAFQD/tA3XEykNhPBhCJfTaEDb/UR5842/TGr0eEBqWtH1H9lR17BO6Ssa
9vmZ+HMEUvZH1iVR4KX5BnoecjvrxD7dI4orxkU+vkLGz57vQfPhRPOywq97A4K5
jpJ2Hoh0Loo1FfIb74ITJJyqB1NbE9U+3p69brMMHCnWyuIwEY4fkAdqLzjP5ABq
ggpnsHi1MaSZNqj71iw/ni2irxVfieb/YHqzG+dS94yorQxUbbxDFAkgzi3eKjXQ
AdPZW0JcXBMRoss96XWyY00U9J599FPIOteAh+d9xS52/eo3Kfan08hMziBIPazh
QNgTmFHISKlwRYmK6//sZMA7RLEVcO/XMc1zi1HmySaMD7vkPHIipRTQ+LibOLRg
K1tf6gyjY6kYZhWh4ZpHiiFG4qDZLdLH9KSls8S/BG75p18SM6b2w3xmb1IouGXe
Cu0mH+TXxeksrgHzlkyqgRRa0zePzE8nTc0nIl6mZS+S9ULDJHEVK5dMj4kUwfG1
13NF12LHzP8FW40uoUKODolQkLi55OiGSdVvhl8brhnbbcEZOIhgI+e9ce6+E1jM
EmD2o1oSzXiD9xAEsrbEHli7M1zSI4igAx2FHIqCliUAk27cl8BRYvEYkvqceuLq
kSkWtb9f3ddsIP7m87UE/pckqkw9OWE6y8H3Yn5MbZfITKJE9WL4JHWE2X12LOWr
dqIm0MTXCZRjIrsE6YaHVZHUr8S40D4UXSRRDpH0dDYJAYfx8d9IbhegWU9JL32+
1lyZQrJVarOQJv0AcaMxqwcSZ/FAAtYx9Pdp/4CVw9peFdyOdTckyNARREhxb/NV
tzRh4szxfVwUAyySi0VJ7oBdXawmIvgYPPJZ/yyTXnFdgFC4jox7nAYxLc4rNUJv
ISuB6ZQfZF26mQuOxKIOpIPWx3yA71XAAJ4c/XigZK/wZs9RrFZc5Y7IQMzbZJ2V
wEsMQS9Q7W0zo7NoPAQqplkOUmn6cV12tVJRbg283w8oQll5ArCVn4J/Qr5kricu
rBE5O+OHWDOBYGqnjeHAGG26v4plnOGS/jyJGnS09Xo4N5ZypaH/x/1wFpMyV3B/
tyL3xf5DatGua4GIh2eC1DAg5hVKLkRErrNTvX/w/JMjlUNkOaufjK1qBAVSIOQe
56BcqBIex6wnUCfPpwXjdJI3Q2Hp8yCwjMLEJZMSMycJzp5bc88HJxO4sgTLE4qD
XxEkoZGDSCxqB3f10DDRilqFWHyyA4VVFDUX6+jxMph7HMgxQ2pqMRrWP5ykn5+X
Vio9fmQGgZuXwgz6ix1XkNut5BaLNpaTuSjtvFLVjWvbq8medxMEpOFwu7c1l5HU
8W0JI0sazLH95kZgH3x1H17BzlqfZiggLKvcG0THnIrzij4sy/W06/kNjtqJBqlW
nXbeJsDO90B/YXXKc6sj0tyTZpjlyvD5oKMZDHTIglQ549hNnc5FonB5kG8uCONV
mtiECULpqapffU3L8yWKn5+5cCFXkiv1Xg/67Hbrq+2yUvTLqPZ/SBcly/db+Xlz
1CQUCpO6beT8/rv9NAGtwgdpyMSdI6ZjOj+w6ADBZ9IwFr/vpSbUT8TRHnayioqD
P2usGqHnKt2v+ETbyqEl9zSy744Rgwr277Du5Ribjy7AyqBtAcRWpqeV4oqa2G6e
w8OfKfMnNhO+qb+y1MPLIxq5f4PuAMzj1gofOsZV5s3zYLcbp+hU5FC1DgTYobHi
p1CE3BZq4CyBlYTiIEhE9A2A6gbjGqbGh3YL0HxlQHN3+yxTAvdqq+WJLpARatRC
K4XQGwJsPwiR1np0WkyP53Pw6MIkHuCwkrgM17loDG1QTtT62Ep7wzOZfyeHgIO7
imF5BlOWRJLySnX2KwwrzdMM+QLqNNWJQjJkpQQb9Rv5WjgZDhpPkR1/7PuxBTm8
VIig3un0sDtXZ6f8mqxM8pKvWI0sNAfHHqQHbVHZCnGQM1VTbnU0XdIT3szBsPhb
gVwHALQLx68Tscrc9/13jrWo4apXBTIWcJeMG9dBZTtd2Cc18sUnNEENY9LGRfck
O+ot3BK9cyiZaouNQw3FPBY+VUDANwSIpxYh6FMSX1yiEAI9GtljsAFvGZWFcRmx
t2eyoL7ja8SB0v1j4AmbFZ1YIOXyggLaXQbasWKuG46Tx3ejdLV/dFEGs+BRmmcs
H3YO492SvWfs6kgEEQNIUaGXYqtxodKG8BNULKtNHgB9DnyOYH3FQP1MLknlSmZ7
IQPHV5+zLdG73OBLz0uk8J7WGiC3m5IzcIR28KMWboW1pqJBE2IuF1T3i/N3Oum6
4C/oZKfwS+P6Z2G+lhF3v70wZbbl1VNEikTgg9AfIz5LeOLcPGT0il/cA7+GiFu+
PMGF6DJLMH7JEA6crDrCda4GVonVsiZDUsXc0peCypiI+nb4nq6kogzBVKZFZsPo
jOA1b8ObsdnLgtGtDpVnxWPquLPA+6E/aowstEGVNZmN4RZR9wkI4YSNueDUReJe
ephIjoUecuxUBoFsm2lQ8Iln3qsGP9Xg6HfSd5NE/dziedGv9nto0zigkyHrfGVI
ujSglJQDZllkjQV3S6tIn3QK0z6esTY1mtjoDA9G30D4HV4oBHsgPT+U8Rou3QzG
DdIvhUPGlAcPU9vQfy5jnh8D78NZJrSxblbRyB9Vf/rmE+8V5DOLP4XJX8fCQUpq
MlzTqXyQC5hG5FO17t6qVA==
`protect END_PROTECTED
