`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zs3EeBitLt/+F31xVfpeDI4G9yrAFXqDRQaRRoeDhgevO2J6L39fjoH2dcDrSwoq
5h5Qr/ThbWyoqXzsA4SMo1hUDelUUeBE7eS+YX+6r+WYRuWzF9H/FygbwPU3TEes
arEgLRbMTZOT12+bU8v9U4INtR/tYVFvkMsOIZRX5nEXt0dCPSOWasm8NjBHv1BQ
wClbFiIxC7PnZNRXNDSTrHXlwYMCWmfHbq28D3IprRPtHTdrb++eQvXZ4F1o6ENz
xPiUwunho4kibcTtgIJXQe6k1iqlcUWo3YJU1w9ucYIr12Zt4qt39PmxyQn8jOBd
+cAxHNgKfvgU6x3ZBeFj2Hm2W74gmSVfSy78ajj3YDAzCR2Nlp8FKWCWWWgB//31
EbSvjBDh19Ex/zb6K87wJgTORa7WaVBeSF5tS7ZKzOteNJ6iw7IfTX8a1BpKXR1O
catw6fJGiOR28U4Fom/vZzatpuoIwwgoBIaH14wNCxO53VG5HYaeqb4pJ5dxjS+0
q84OZO9U+St3tcKd0jt8e3OhFLppFfX61jS4BEEO+L+x5ceoCtz54AI3V+N7s/Yy
+QT3VSLmVWeZCCjxsu6YO3zz2W9MNtt0G04ugvmCEIjhFpIGLLiIT1ta53v1oxK+
YARNo0ky2KCFb+guUYoJBTyNbn4dVeIwxnTeynRgqotAIw6/JRTjplvzFisMkp/k
jHrwjo+0fmyxQwTVbOUhFnGiTCKi1mqk4qznpN6HriArUM6r3A+HMZvuDcbd+M25
oX67MuIDYl8CWLtgr6rGQrEpKec96hsV6yr1lDWMSqm7EBk4YnrR3joaXOpguWZ5
FZwcwIF/H/M1mM6HQx81+7X9GbdDpW/icTodXv2DeWHmLA7r8IopZE/KNS4sMfqG
EbeMW/6iwDBnYoWVKTN0K3xzCpQM93Iz4dA+3XiAs/sWEbpaAVSsQ6Gj64eU85Wi
Ti2+ieM8txc5BSPYet6g8lm7qwFTIiBcKcJzbBlx7L37DEnfiiVFNsg0szJkuahR
RByPoXHplWPR6gUQGAxCcd3aUBsmfptRBiMb8fA//T7VsdTX7ObMW3V+uUfG7+12
sZ5JcmL+IOTggoNsQZCvyQUGpsBNUFCe/lpQvtJLOsQvh/usTeMVQyQ6rfNGvH6P
T6B/NdQuXbk/zEk/h5Wh2qWAmKotC+Qvaok58nwzzPk4xfLR2KeoCTAHiD64bTpg
4OPUpqTOcOh7JhFm2f/nmjIVmqFQOWUJy28CHrKhBaAEqxWao4jhq8V++Mk2OOmq
OuK9DyONRROgxnDXnJxcD4Cxg3HH3gYuRctgHK5HhiuFp4/jJtQLW7V6zR7JkQZc
/Qb+C3B3MgvwHzGLzOF4WLcvWWZynZhH7TOWx5P9kqS17dNxkFafvb2DbEYJOncp
OHN+wzj+alJVWs8wvZfaZlMCXfo61rb9hvfE54RH6oiHKtbrrExG4ST05btZB132
KYhHei3Tgp4DB9oRG0Ju9nYn3TzhJpKQkmut7L8Su0+GWSWCA85w6Uy4kNq3R6RA
fJxaKAm/EzgBM4fcDeuys3Yuu6VB3xw08PLW/IGwUs6+pynK3vizT1e4lbmfWSWQ
AIU5XNEIfmVc9/d+rDjR99e3V0+cSTaIj3UkxtG/nEFSqzKowYRT0dvm13C0L8H2
0bknts0hReZYidzRVflz1HXE3Z52tP4NrNcwcPRz0AMIIx55X8uhMTfKLwawPX7f
pDJZ9swZZwXdGedu3F7Z0aYcvbD8Y9fDEjwy0ms5g1XHXj+0fXXsYwcxg+cZEJ5A
WOyP71KWylXozDHWXZXLQsXQcyStHV6y2OcsTVJ+rLMXxxPBnqbEsbIUfR6abLJm
LWqhZCvX6BRDEj5uPBOjcphaD+9uB8C+cprkrlYwmKV7oDcWqWn0mW/KBGXRJuSI
l0AALHZytyMb54/U5h6S4Xb+aWeo+VteS9gtWcl+ElEc12VAmu4y700F3VYUrcAu
asBXgzQzd3gAtlXfcNLEx2NAaTnSLoSjR7SZIEyHaaMBrex9mbWoghGWNjIpS1tr
Olyn4J/V0RlUTGaJIjxGY11hcfH2zCTtki2o3JQ8Ka2y9Qc5R+yWg6eLsdn96VqH
wfovuNXO4BpDgCSE4tPZC81AY3+9odY52Za3PXfEuYgAvgXkae3z1KsMEnVdTDIm
YKM5wvI8bp/D6EcFca5FQmyJqWb2r6DUzl8g9zENJRKea1T/qgXrv+kEIXsbHtKq
ZRI5hTQ+HDQUHlodHu47zHpBjelCyn3lpQnzmdjGaAeWl4aqVySBuP2J6fBRuna5
IIf3GjN8aRTGcIyXSBiyxtxLc2o/QvVIGk453ssPB4S/IQ6YLPfGjS3u8loafbjw
lx++/TnX5U2OV4VAGUbwcvL6LL0I1ZgsXB/rDB71OXSQfx+NVFf9VfjupV8RPhqi
IHz0Am8zFE5QzWUjIs+BkJMDDZNZvXeguf+JhkxEe6QVO1WIgMensPtcw3oY4zuq
QOWxYfjiwnT4iBP3EQvl2VIyyFNqPnSrRZTpgO2LXiNWJ6M9MddMXhTmFPYZiC1z
WvSyRRKUeXmw1txOw6HVr+fAo0nSEcrviQr3Cmx2M2TA5NRtzA2u96shwhQN/VLj
9+mS3QutcFa+gGxNPD3fPs51M7F4bxT0ycyrEeTSHlr9vXmwUz0LYt/T1o8NVnMT
jMNky2Ped/SGDKPQwc3q6mT98PtsoWRu2oerZt446G1EBNm2oTEu89Om0xHPkDDS
wshtw8RXi/JyB7wz7JfiF7R0c+G+iHUGT1w5Qo+gCc4U8SvHSG88N47h/faCHVfY
AwZQdbbbSX+yiQSRCo9HSyztfIFVac/z1BdTfHQDKuUYGupeDgHLIJY5ctOL50x+
wC4wQI/9KSuddvUE2+CLCu1ubMu04Jtp84x6cCVzPAx+EK1TyTAyR3E2Alq/c84M
tOWO9V3DXKnmu3tgXVxnQF1sNpJCt/8D1xlsLvPoT5zLzaWdefiP0vBq8hc62Yf1
UxHOyZ+/KksDE8EOgEA/FmwH+VN+T2gILzTuVCLE3hcHEVvp2v2T2OSZZHTe6CF7
amw+2FyQ/sKmZbu1N5MAguEjaYNZsFiG38ZhqKi/jBS40owuxoAvKUCFMynkkq3J
QY41nHYWmDKbCOs5Rtgv/ZGEM/WqJtHPSxeDVD53InoUqSAW6t3vU8KpXic7SBl+
6/z2m1n4QdnjRGQdu5fKS7wHXj6Tp7wlk9eFgU56OV3k1xFQ2tyBFegesYWfGXgu
6dTt+iT9G6SnsealFOKjyUB8qvl+305M0jEFzzJUxQuhON520bCz4D/rpkbSn9zw
+BThdeHITpwgpJKv18cDEXTZlhwKw3ieQc/RLZlqPGRTfN7YOvMTF4DJKc2b1bi2
eJVE1LJCx38/Tkm9iizzKNt5VSzZGUc8euSNsLMViEtFw5Gr4/EX0L4X26gUX1Lj
5a4DOTnrcOz9bDAgLz4C9IAHrScSty48+++AVWzh5GsCZfYyLvNWaTHdV3OPABW2
K0mTen9QWg6pzGcw6op/JpgYGfiC4aCDHbCHw/kwZaSAD2kQPoxI+Ag/ZbHzjlhb
cbRalEBuY/LQXyrfc+eSV0ypBEHxnvRzy2BwfJWpPbct82ouQVr3JDes2r7s4B7P
kzWsLZ46SojueMFrhK00loDxj02L/Rj/kL5qj4nzXXXrEM7ldGYTbfXqBZoYdDwl
OizYEIVdNtP0+m9xrHDItr/9FfIlD+KlFFZKEzmcsBLMLQ3aVRgUw3SelZiIh2F8
lOdbNBXdp3fsC3nTKcMPmBKX4DefXlBCFWQLuo2KzfnRoLsFbKdLldWgbDsJqjXf
qDes1m+/gX9j13DWRuFNnw==
`protect END_PROTECTED
