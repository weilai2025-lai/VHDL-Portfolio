`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
td0Vd0yVqb89NU5NdVe07wRCZT3nZf7fngiJiVKuNKNlL8p7g9m4lEhudGHTKmz4
wC2PPGTe5eeis8w3LrBW8T+VugY4w8TiFzvjfF4qRRAdjixvtiaQdzGsnFc9MK07
ppNak+ollo2A/JUDuZ5K0vA1Mf9QrF+umKtSbgEH0gigvhP35OKWqldYv6IA3sqt
GuCrMYh7VujmxqL6VnlOwkPbHQ8uHz4K62bteFE/n4tVVQtr6wSyzoIPhsPwWj9K
orjv+qVrJoDNjHwyCT1YjLa2cyTRTW3TgVZH+GEvJNHn6+b5iRy0fW8aNlUD4m4k
nSa7jxc1fz0ZluB5N/V+3Ni3WKbsJs3X9QaWHJ2zUZgN6ECreMS6k6IpPMRAq+c9
Zo4gOiaw3q+2TS92/LXUMe+dJ0y+JGJ40KI25BRTN9sUfsDWBP4ecWwZFJULZE2E
lk5PQlD5+nGJ7vd03l/n7fpBVN3y7/sSbCCMom/zcHAbz00F6hj9wN0igbsXt4B4
15CvKlugOG+ub3FSHUG4JD6mhCwg+vqU+i1mGVK6irfCZc4rn74tbGQOnpUDLmUs
lB9qCc3ERgqZrl+KTRTK4oEfQP5yyB7MI33QbmkzYrqspnW4rJIo2e4f9hoyj83C
G1ZTKX1NCuVRILl9h36Q2efOfVp8m3BV/pgysZBxAcoxjcFZiwgrhG3N6R+Qjd0j
YhNRYmDaLD9+p+tlkkoPyzjDUOdZfkvhDabfh7awzN4BUY1rniTjdebBguATZDmV
Wi4pKL62oK2x20sJzDu61S7hkc1Xvrw9WLK1yTioBYnPK4nZEAhKcF+Vbimrq/ih
omuSyzYCZkd74A23BOWESH+xR4CpWkwD2x7FPMEBIPv7V9fb/nv/Se9yWsKNlcqn
`protect END_PROTECTED
