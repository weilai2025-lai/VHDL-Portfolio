`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Rkouuf4lHO7Q/RzLt5607eBxiJOyleDRtYcgN9sqBSbPJxxq/+AHtYQ6lNuuaWD
Ec96ZfuVqr0NkuTze9VBqsmfVtmS1LdlJman8IZF1NdNaEHMwZcODdLkq9j6bgFw
sESNWNdE+/W0195d+iUQnN9piQc1Pn5cMP463Dr4DdItaXy+hULJR1IO0rH8X0bq
jSY0h2+SAbTdjltlMZBKqM5hNx7vUfgzGBbOZNVuOVlZ9CbyduvMqYkP/NP/YCel
L9heFr+zG4/DglboHGM4qyHT63v5rHJMatp7HZ92V62wAjJdQtfub7vaSPgSO6TJ
1rNPA5ily1pchQ1DKwNV6IF91ymy2M99o8t9G3yG2UMFBRTsgviSbGe7B2Wuz18c
rZOYyOp+Sc8HKNKrzudbz6JKnNFDmf2B9OBPIiqDS3Wyl50Gido19KyxWl6hkvp1
YGZ4H9lwuiygIC8vQGlylojuzv/gueSzGbb+wr7GN8jzwiGkP2NxRVGcQrItuKVr
Af5AHq2qwrLql0iJbVeukRVkLA+um3UiYmmFdaMg5/tHtCx/EIio/QNKq+6Jnh87
LDruD+h3mJyIhDwboR/6EG7MOFNJytLXH+UuIS5Jf0i6R6x4JcLUt6404KA2wpYb
Jlm6SIgKhvCYLVFACt+93UNJ9O32xSS3D5c0vgWWQvfOp/JCZ5Gp9qQd3yCTAmm3
C1zn/fpwXv9229vTD2Op8ZhTnvF2RTFZSYtj+olAOelIVNm1nSMH8w0UC8Ii8XAt
x9hnG8LR58PTsCkWeXVUDK2nuwO9d7CAClL0VLu6XleX167rr3qDOo2/6WQn/wn9
08BcdeQe1zX/9pa/MBX1JcX4KIg1/6doVErBhBkqO/RWHDhPqaKEA/xxKTRvRQdV
y8LKvoC3NrB0HTA30Wj0mVahZl55qQCTBofAi4ZC/xNRkhRRmimVnGBd1tI8HMSd
HF4n/ZnXq80zfIIV+XIgLEQvIyukO2LhN63kuZ2SycG9YlajG9xwR6T2egjZpBL1
MY8pqGOilRwPbR2FtzS8dsdRL4ZdIlKmwKdC8COh2TsjB8tvGRx4yEFH7mVLnSXg
EIwoiFTfheRVpC0KVxZrksGaxipKEGCujXr4rvLwX9/YbVZtNGTDeoC1TXxeTFSo
h8jo3JoCL4/vi3hsHvJATlpKQR9DGHu+UN4h1mhEGaZ/ngTwhM8mmEzNr+eiJHiI
sANYQ6V/9fp1nha0WKNhG4M4wHfPfh57ZNtqyNtJUCv+ldziiksZ+lOx5gK6KCTd
VorHnltKpAXEhn1mSdrFSoWx0xwsAzt4shL3e6zuYfQ0idigbQRdBLtD3ISSceHW
eQapWAFNppkiISIgMzoAnv5QjcGwv53oJeLe6fI7ymSUUYsqXYOFRrchNJp9jRJ5
YSX3nn77TbkMvurI808rd/NNsYWLe6xpXJyLhJKC1Ld2tGJuX1jUP6GUXaUmwGGT
myHEPI+FLxMygixxejL8InaDN8weLlfFEOtzoZFI6/B2iU/TkhFJRRd0W7tgL5Fu
4+QQVbtU6BFRGtLDHgKpk9T5E2d4z41Vx/Kq273dehVVu4yz46hdJ6NmDwgmhBid
vDsaTPwUXLZYAhwhz7tHQRwZp0zauHrkry6mNYsgWLnTsMLz/h1Ni28XeTtIiR/a
cpSqPiUcDLX1bwztehP6NILQL2rxvCB9/+nhTzKRf7wcRFWMcVVkIsu5rp1HpJTQ
CUsyvJKVfgS0X4ZH3BsOkjCN6/O2Nhs7tS+ur6n1a2eZn09d4d0Ks52v8F9pTRws
UROx6f6brq0YsrNXHNdTMNEBrszNBR15+tXhLZnfFTHFVA16R2OlLNbQUUUX0qK8
BfJN7+4y13KrekUXI0hPwaJZkIvsYsRXDwXWGQJqEE2mJQZxHxNWP+u/9CHfycGI
wJJZu7EYnjl3ov5Hc1oB6OjsT8yRwzOv/pDJWMsiGqdrXZGmDew4r6l+usUMtH6w
qd3t5qA8AaU5MS8l1ptlCv0LIwjpcLcESLCJWViVcQ2mXv6qu2JB2Q4U/qyq/iGf
4jMujMVZVlL/oPIM4LfFfPWrfZjCe3rtq6zx6nd7uGXliMHgdRHoNmWW43YbWZRM
dqMEz4fZBoj/PZ2djQ6hKmkfj69x+LQjvgnsz1S1aV0H8gcFaaNw9dmluNkqa/xg
eVyMPsKrjB9bq2jYP1eMa8rh67Pz2gOxENx93NV1JCogvek75AgwHCPkclVvN+rw
CE3hUyvnWHPuolf94zvf8nn29q50Ex/uzjkYPj6jLJyf2MXGFz2szSzHdT3hzjuE
tN7JCj9igTAD3tTfrneKLRK4QVF0ue1mrEe9FLxiCIRIklhBtXmnZhsLwFH9gi0k
3LVJNNJCuHPjdglyDZZuVymdqUW2m6PqMPVvbKShDb2mEln4B7m2xHEBUdj6Z2sT
c4c50LfbsBdxuusNIGM1Q9TTEwJV48btXGe0VMm937JHZxw3Mhv936Nbj/hVH6wE
mTQkznyUIMUCjg7iu/jEqPheF1qWtXvlt9L+TIIs75QvXvaMiGRSG0dEu5AUMk74
X9d/L3yp7ACD012w7kVIzV7h9Sv8xTsu1kcRStFsVtIDusGCMLRydYdzTLasa4cI
ORmsYT+uSV3M6ft4SD4BPj9KEpcGOfB/tOCXjhLrmI1Cuin5W9V668rhDMmCBTKF
`protect END_PROTECTED
