`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mH4CvsLwKtXmz0M84owUZQd9FpqwUM8y0BFwEm/kT4y8EiPEX9fdvLBqgCmlGz2+
lbOGAFOQKOUhdpVkv6AL2ErfHl2kjUNjM9VrsTof2PhuBZ79umsvqax3LZjh3RMC
L8vNJ55Ea7xxhNDORUfR2MEV1+benTxzpB9bNtIEikqGG3NHQXuwD/5AEVNaZQgW
oxLVh9V3EYxT+4lUoClCNufVcA1C54iDIFRttvB3DmHnzafGG+7qj6bJKQerugqx
lj7bQ8YEpU99dYSdg5wsShOtPbkFkw5Y254tt1ntrT1XVPFjLQeXnEKrCqvhKpyE
Fn4zhqqiMtxsAx5f0hq+dAxKX7k8M1tWdc2l/fibAw/8dJ26R5WrhWhp+5xwpmPd
GL/TnE3Xenexljpe+v+jgOFtwaDKvuN4ie5VH+9TbtU9vGGw9UXLzRwghlfkampa
TbEOjB/vUfCSTVl+4UI6CxB4KS+8GFXG8EMx3gxC9+VPbwZut/2HEPX8MMfDmBqG
qPjr9Jt1jJF3rJnQcjCp6anRhFdmXRVw2AV6EHHR2YD8xWualtN+UTDhMWwNXSc2
dFFV32FNfwh/ndPXvel4fbjrDOfBi3rXf5hwD3am7XpDhFegCU9EvnzPZ81BLmL2
UvGTdPnZH59bTLa6PHFOUURa9wMoGPeGrDyc4DH5/8RVB9wqtzELWvhr2Qj8ZBLt
pHNpztxLcFchVTUDUTMDoQDI2lwSYV0VOEMoSlXMMCiWWyUgTf/nPhzDu9jK3wU7
+Kc5Ux4iL83Wk4oF6xb41VqfxQMrft/L1lbkrHxhFNmcCEQIIYiGB3EGrvS35x+V
Guima85YOaSrsOZDGoNPBQ==
`protect END_PROTECTED
