`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RftWcSOyDa0zglV1dcifxrzmRUs3nBybNPA2nsuyZWtgUnUqm7fjizlYoZJMgGRs
s9DGIEW6j8KD0C5XLq4ynKznbXStc6SVa3FKJQ2FcCz0gChrHQ6UHYcJGzw+wGaV
eNlT7EM1AbVEC2+DnTRIq1gy8ipV49MFOw7y+h5YObmy9p0zDyEFz9BWAQV6S/YW
9eJChyRcrHvgaU6kYrNgiPCrrLFTeimx1LkGk0+0hrFvXl71S3n7M9My/gmaiOej
rjxRZpQfJ1a3T0rzQM5xBA3C2gxgwJa/yCUCexe8n68fmZJx5QCy7NthhEJEeGEI
0W90Re3ZjiHn4JS6UlpP6Sn+pbu+uAsqG5kyrTCVSi6If4ZPhzuRaM4MrWtaf+ir
wHqKqk1GcTgXHFkSECpJhH8E7IvE3gFTxdKkJBgCBi8J+YvETU0yJtyt7eC++pNS
`protect END_PROTECTED
