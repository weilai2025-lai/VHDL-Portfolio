`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
heGXY/KWndpx8YGvzFMObKsxKdxFvRhWs4Bplw0L67bY6PxO+Fvdhi5ew2taGBbU
CyHxLyMnSg7QzkvvshgRWltW1IpUOcLeY3yM+UnQ0jmzlZ3+UxmaA9+AL644xzSh
UDjfRf0JybwkXn/fUqb2HoIiG6NV384xzVQrOrm59q+Zn+lW2kYRqdmwoRv71C6X
9uqAPDVRsBFouymoIzW8JV+BGvZ3StC/YChadqYFuhh7ZnEPu+sjmS/6dkvjet7Z
HZyp8/f+OLR3+RB/Hif1lqz+RiNvIWNuHDsRGyYXqDuL1MlKxVsaSoS3KjIcoITd
HWEW2CyjzZJmyPrd4Kiti774WG/vCCkkBDL0f1eyIvqYeJZIlwt5LdnTwnT7Bk0v
ijdLxRNTtrsDiwCSa2bW+bb9iWo/7ixnzjP8TdnK68mDYE8+FmwZEI3CYjt4XbA5
5FWwHRcWFdS42y9LkK007N+k0ASyHuL8pzh022BtiouK82UW+A7Px5iJ1pphTa/J
ws5b2FTjq4ZmRBbDnthVa79Uy5turD9EMdwmTAkbWAY=
`protect END_PROTECTED
