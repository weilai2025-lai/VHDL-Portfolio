`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8X1NMjQVtflKRf2E2KGDb5DE6gff6gpPjXEHkwoEK5ak+Pijw/ryQpP0IBKYVd1m
JIGZjSCEaHJT28tw/RW5KEdPTVgMcx1tRjysdFM/sirL1/ibGBQ8j8NY6V9bn0J1
FOYBdIYAPDGHaqI8MQMt50JwBzExeGB92lTfTRIjWMv5zYoELc680WvE2lMv+432
Vhyxvx0J8ldMy7tOGyZ85q5Xjc21A+BBOm4MUS+QiIUmpkuXN/bXurHXs96jtCIE
MMQiBArj3S+oUssbSbbyMel+wx6CCtCFHqjJsMlip64d6QM58IYEAgSkkoYhyZmW
gsQLess8rKAJ1OHS4HduHwl221BA1CvSPV2xWrJiqr/C8vhN/ACanCvfITIm6hsU
zA1kHgFyQxGedB4FpYN9Q7UE6PTg/b60tcJ2mdHWrwJ8g6A7UxkgVkGwSo4/Sa5o
1WtzHqXyfgPqyv6be0IQKDvNqD37DswDGU+N8+aBub0xe8+0LtjcIaPp2Zzrhhru
1D5/GF4S9SIjg39q3asJV6I3zAOKvGQu/hqn9eX+f8IaJDKuppz6vL3oBsmWeKxu
O4kQheuvZTIhpjlGET+Z0Bd0WSwgy/hgIRzjowOHYtwjtfk+hfjVDbPkj9UNrFbY
rhOuzzS1Bv4JiKAnqKt9G7A7dE7WMF3th9/jcHMGO/E0Hg4auEueHO7vcUwuvIxU
IxA6/8fgVtpsHHaNVCENLlYZG5Dd64VHNNALuGy7zzQUU9pw9wxBOKngtuX8xyvK
zUNCQlOpJA+gFJim7JEETxAjUnGJSDESaXkL2nanWo+ZmqdLzIabHAqkPg24zxwZ
17EYaXvDFBOvA1heA9cst3n9a1vDi0a/qIcwk0aisled7/V82BxRy/ykyFKhiP2F
GXDHIO6PAKK4eU/0haz5SQtO+8EmbMaxmYjtM62eqRsrafYPQ4J7FCx+qqOgf2gg
GdICJywGVy43lwWWUTkW+P9K9GIfSh2/JfUwDxbsH0O16vKs5hzEu2/n07u0IKEw
1c8ISOCSdIstE9LBMcHsMh3L9nBAlNROSpbU7PlCE/X/1yW/aorz7fiA81G9Q5lZ
slE/IBmxIl0Pno6AgMUefqzHYYAVUXhfX81+hi6iOq4RN3N8aDlZuynPW6tIJvuG
OzzE/3vJB9FMn1wo3eaqNdtObNFRs8ZRczkM+jkvgoAoHIi9Y2Z58pwTMKPgGNLi
SjZobX6nb4H4IaRBvf4tFHmeBaVkI45lLi6STyPt7+qg+qzTvteQ75e8lAx3siLI
t9I/pO5EbUBHGC7tpdNgv5cDCnfRxvO1dZClBmxwwldDMgMwge1vcCyULl/+GOZP
EOU9GanT1/0r/pYlN967l8OxoVllxqEoFAJovSOmmxzEVVSrn/Tyqt5PU+lKPQoU
HrpO0AtZS9lkesljSsfkzlkK6eUyrbppX+Msqx5hyAGxH9NUIJ4gfJo+cow5GaCm
WThLpAUYxod/eFD7rbo7c/ISU1K+aAOGAOI/hPYMse+Evz0CYntmdjjcz07ut1tT
dAVX05iYxaJCKhqFkg0fCkX0nGsaAMrmU1eYx8PBn1L9NHJicXjxdGeeIXWcQ8tH
3sLMPtmBOsGne7aOatDdJ5VpPe7K4XOLFd6Otgvy5BlYl0nuu2wGRw33nS2TGuUl
i8aCwj5Aj50z9kunjf8n1P8tJkbIeZxK8MAaxJYIkdXLcgtMOsRbHANqPCN3foqZ
0P+CR4aVib8wm5eN8Y0pjwhKii5mLxrk8lAPHjrPZ0NlThkjrB8KNrpWtbco1XgF
oJgQ0sqlJTS6mACkzxA/zTGs2ulnk1FcCOan0SUxfRX3gh/LduhPuPMhgK3IhyhI
QJuldQ3qHtNvF7tc4NPAz1Lf20W74S2Oi+3NlrnC9ZTPE6vP3Jf3cwkPLKuwIf9u
74aynBLR/vAxZ5dYzJWPZUjBEQ4St3vwDvElUlfamPhpoWga5+cXBExWNNvzIpex
ShbcazEd1N/Z66p2KmyWfA8JDGBEUe+HfPy6ACp6mcZBBkfZ5tdEKxoifoipXq1K
bqmFseWNfTeCHLdEukbJK8hkO3JYsiwCdDSuAsNFNNeYei/ZCOZtMMBrLBK/j3bU
fGnptOX1dfiqM5IginBwtW1Crp/1Q2Pygu1K0kFApekGKwhmcq9O8+G0jy4sHutl
exns+NjGGrBKKIZcrQAzT1R80DwQm029WWs24TDuYva2yXfm4m5dZxRC3ryLNWHR
icjp42fVWSV0QodbAp6f7c47nm+hOh+Jza4Eg/pio0TUQ/7kWhOc8JDLhLMr2T9M
0Z7ojnCuf+T7TT/LJrzfK9O8fC7TiNk81hfRocwXYYp3yhHqG3x/hdJJ/7vJBbaa
umDGpb/gS4XPkoj/xKUaSMqtOQkypv29Hc24O5xCXYCINDp7nN6uTMRvWYkunnXC
4ZrvwlFz7ZltVE9Dzda7TK576jzV9Zkrgmf46tzqVRHpLhDJaTal5L5tblPYGRRJ
oJ07racUQRq8El8Rr6pZg9ypSNsfHU0e2c1/ixKA6AhAKVoJgWgijIAcsnAwdbDP
4ihW47GOFvglRHP7RodmKujHClaXZyCZ70NVvaI87JJAhHykQBEpOgaW0Jyw+pJx
siLDzPjdSwroJva7pfwqgDVc8r+qUcDOVE+mI9sWL9LPSf4kCQySFnAJKR4BAjmI
++Htti1BHc4cn74KT9SfPUvBvtcZUHaYLFa/CdiwyMuh8ZJ4KQGxUilRUGnmmxU1
360P6/Dmy3W9ty8mn95zcik6g06Dt9lCloksb+op/1Z3gtuNILr0ufpDUloMzpmW
JsEF/Alf/hn6Jq0H/EcblL58uFmGjCEVZLHnaMo4wk1mPajqVjwxQGNvFQiXQVM8
JDOeELQTy+e9l6OW/9ZfKGg4uOWuYhlip68rVmRYueE+IGOu27wA0TvBm9nOwk9J
LDfewrFz6O9TKD1EY6IapCiDFChhwRORT01GFX/CC++WB0DTjnG4R0dKYFi2nBFT
uf2ANxzHU6NeD6exay1dTmlKnL9GPMLyD/77Wx4m7JrPXRIdTbcGRlQWqF44iVbk
9Njx5P+QAMCykNwga2iKLuzXAprxuaPF5odVnn3iEwXnNsdKFwkFFlRdL9kWaf1/
Dxpohk9Q5F7haC4c8lPCpdIWS803KDAaVEFrbmRq7F5GxBxSqJP//q8+Z7ttXfLQ
8pctaNHy2TfB/c3whjTHEWJpDqRaI64xKar5k1HvM+TiWtY8HBuQQXffOS23064z
5bFVFF8h3VFd/0PpHaYo+dG2/0J/juWi+cr52qZSWTmQDhJiP4sc8CksH4CeusGH
ot3osMQcu/cy9eMw6p1rMaAZZavtNKkfZDNppsMiG+z7hWZx8iTe71pFvw+P0oDm
ngLxEMLYpZN2jiUpUfB3UP0GKkVZYGppNYpzGDbGUqhpYIM+Q8aWvunTc2RPJymc
Y1D99bJNFUVSBk5LE+h7qnY3jS7EfktSnwHSNkvvjTpgWTdsGEQTz/w4K4gJcnnr
ig4Hze4VVNGjJ1DT04l2hRR5S7+TY2rkptyRFmDRpFTq5OaZcVLtNN0yYrFE76Np
rG22U0oMw2aTvE/xqSx4eCpqSOYbFjIPRnOEizbw2hzf+hVpA1A4ZgPoa9n7VfLo
DdO/9fUiWqKeRstCqp8m9BCeq2JBmTtuw/Rf+UdZM2MOQwySpRfh2kBB1+6eWYVu
Z5YSc1iQT1uE4DHsklCMEitRmzpwgFGvWuWXwRcANOavbYJ8YwHG346lbSbGaVcl
REprEYonA6WP4UUTN1h0+RUFfx25HfbpjnsceAOwFCg8PJGhFr7vafSFrwxJzmr3
SNaqLsZTJ1g310NAdJw1wAX9pwPpMFtLDGgqIRDdqlCwESWKrgH5MK+DNDM3Mwr7
qgkkWls5r8w11ItmjYXVjRmhD0V14Wlq3kckmZMXcYxC7cGUxuTv12aHwqwhRIOI
SHtj7nldfRfllmij8QYvm+JENFANJdcHdRyM1HE4jIYXQvFWC32Dp7T9jNaTxuXf
8H4XQDMoALj4LXSiVCpiFQVB7803PUWyGNnVkJAQNs8lzCKyOMN/7PT1C72L/QI+
l+PRlqRE0yEwUsKzlbGPSNi6IXzPJPgDlt9FBhthz86iu63tAKYycygudyzfWugj
F5bZmXb2gxxBudFE3+/YbHLj9YMKRkmygFih9Nx9DdXzKDTMby3RMh3aMiwa4kBh
eH4t87esH1gKNHownP2EzkrVb6bFBpgzHra/DsAgcAjuWZT7JRiQZd/P0hvO9Oid
J7c7n2CkR+kEbQDIDTn7jwpuRuhqHWPIEXa2Yp2oqs/kxGBeHEqf2oqXEBHG2Tf1
dPOX73lt146p5M86A81yY307r8yEPbAWJ2ABZjZAo9v3IX1unmScgtIxo49U2D48
0C45tGS9rivngJ0Xrw5xeX4bLK+eHy/2/kHUYSvnAxwaGJ636fGGCwyrjgEhqXvb
abwlZSmJRHCQyC/woavQzO6CA0MgjFqWDZucVFEHK5vWA19d0k3VB6M7KN8LKHMn
cUdmA610J/hih5Y33FNNwcjt94mE+3kqeHagSeC7QoI0d7rT4YVDSJ3kpao5PJR9
/o4WbkqwkyOnW1Mel7MzqvsMmicTRtXzQ51iWpW9Rnx0v2MFbLu/UcL2+rxVO4pg
gst2xiMjEG5bDpH2HsyZAh0Z3h2ixj8NCCGXddYkhTjZUl2/EuF7pc4tX3Gy4eAb
Upv7a/tyJVVnuY/ws/ocRQTaMU8HkSl7+ULUJTBGKGKbi+RZVKvUF1yyB3GE5Z31
uXyigttcyn4JMKWrlSdcxJAmGsfllJLI6nWIfSU1UXVhp7F/BNu7GOm1mVSeAepN
CCUTTcOUsGqP7DtIQu4/3OwMYUfwCvD6Fwtbx2VnJIEBFEOl57EXLGgPEzmkSHPl
aV4KyuaBJeDyufj9yyXhLDwA/gNEZ7yq8JtMwNgYhUjdMTKqIXWjBFrtfMdV8iXV
k8yLD7nbm52UwxVZlSFHNLFxALurA4sSjlkDpb1ezyoWnHGYUzSbqUy8O1ptjO61
cfH6UwDHLB1LMEOwjpliDL0lWM0jN+eANdojntg1XQnZmzw3FIpgXY7SDKS7hVab
vlGx1Vp2ueMluslskoijRocd+0s54jz83giMeh7PIAM9K6taR53ScEsAFv++gLyr
NsC53YyoZR42JIwaCSR53ZPiem+p/SprA1GmhG1nWMTQ7SMHp/aPEwLFGvNM0BAk
nb7Ntp9dtOVIuFZca8HATmXvMQVzUGcL/x66fFHokk1w3SH+kAZE4w1CqN5WjuXG
McbigmHbboGFJfnUI2D6CEdXy/93o0w4Axfw+2p+LyBwQh7Pqi2R1cuZWg9M2PjY
KJQzOWULmLtRY3qmfO6HmRGU07xs2ekU7fIDKbJLmZIqbx41p/aTNnlsnqc5gkof
BtoTCJvy7P+HU8NC74qi/ocqOpq+OwpX+9vIwaJj6ndKNOeJa3/iC499FVThRdqB
oY3WDSUlYnryNVDtFs3Ubk1U+GZ1dG2jZ2usowiY/OXiRFEIPz2A5S4rAbLy5+df
bJoyZukrm6M0BjRWwqR21+SUgDUBRx/OPr4XnuQgbr8DVL9F3Hry/OZcBKhaA6N/
0tyW9NYDMBzIOjGBV2lgaLnr0qUlhxWe36GSpWUAgzsWEIrV6TiUO8tvYT6KHyAe
xwZ5tH3oMyvzlDgHBRZ7I4jcRgF1JGpA2eDMt7Kr4fVfB8SlOpeeufM4U1CZbMlZ
LDP9KtnGkwlOyvTAI1380kSKEx2zyZ6yBSLzh+O9hXcq+00JEHNwil55dGqDi0yz
2l7bSmm8T6ec+u/zI0ky/yIK3N/kVkJMHY0c/6SmMXCzX0yHXhmoI7rO6NDcIoxE
gvIZS6Iqq4sJvvg8uugxawkRlvyTbSnlyG9ZKn6W1LPjW7PpTMW0ntBonyI19t1Q
lPFSV0pbjv+UgfjA6vhYUrOzuXL+XHrIJ8ZLZ8h33b1P76WDdCHkNR0iwOU+d7Jn
QFS6ftysAQaVbXpJGDfi4zXSXT0+sBH/hKzzyYNQNTQ2QGCs61t5vSgJ8ZVacZ9j
ED+Kg0Mx4NDeJvu7jwZ30PZzOv53eBQJYT4MvKgwhjKUMHFzDisjv5bvi3iYG57L
gPw555cVj5xYWlmohLUNoL5UT0/JSdFDGUmuy9LqDHujVQjcsAZh59VbHxwyjYNn
rEV5hlqCKIiKfL3ZjDigXPfMkw3fXveXpOq4sCRhmV1qLRFDb4s1oXb7lCyvk+AB
uVUSk/t8E8iEoPMWgWmXli0E/FdEEqu6NBXECDeDK50oP4Z+iy3EH1Shrhng6w3I
PN1CRz7n9/E3QuYjCAYdsBBQpnZeEgVKSqwnjq/aP8bRiHrBxo0R6VcZgTAseGCF
OgZPSB3ZfTepswpcSBUzdd5zuZVFqdjrdp+9CysodhABPdC9r+x2C89XnuXEUD7M
Y/w7DCXYLoYPZFOtYlHhXhvQBzCPLMJZvQK4OSlrO694+RGz5pssdP/KC7ibdqhD
NejuDacN4ODWB/6blnyGGs3h+deQVZKxWzHIWam9nLgyE5BReolVBrT+HVxKrMOm
Xiw/oqgxFBrcwyPfmKt/K57r+vxYMBv3FAz/4FFBLGTrTYCVVxTHyrdbNOjNgNZc
7HelEEkIUKz4W6O+BYZE9j31DiQnVN8Eca/p61v1+J8I511j+TZa/9gdoyXAu615
kLvCsPx0Dck36/IQ6TvmUkBKAWmFj/IzMUo5jEyTjDnkpGcPSt6vJRDYfyrAHsGo
xuVJNuP99jpPpYO2PoPSVYYV2t+cn/6/xhtcOkX/2R156pjB9T1HEEmbcuUpatQW
hkxjEROCxZ+4V2YLfynTjDlPk6Ouwr6VYausmt+M3MJq9vktq/WmHnHS42SOQCkH
TodnSHoCrrVYw+SprXcOnKdcrxGy3vuinV0byQqbu5U7FlJJ5nJnIcqi3Kgnw6Id
WfVAxDXer1z5FbIlB/7mC2gdpb2uRNrkFXpy9hbF6b2eBDhGozkqfFvXGVCqvIVR
sW0dG08A+w6S1tEM4SPqiiH/4YZedzv3gOnW2+CWN/fqEwMO5qYXxq+5cUKBnDvo
8XgWxHKI7LEA2yfSOPTVSWsp4HKulEeDWGYiYaG4gSd42O4KsnCqUTCToVUWKErU
WFi4G1EfpGvfdCPNogk+Qif7hT3lWKonL4nMd2UDs32v7XDcUD8hLhChah44nUZi
9wmt/Aop1K9WHPPyEa07vmhx28dZLUiJ8pC0WSWsJx/M+k39WwIdO8QZKHDTG9JX
VofI4BCk1lideNNTDMNwxP5HcGQIzOY4+77o/TCydd5c+Y9KSruN6qyFA2j6BtAD
Ke1kiySvt84gc/OsZaGY3Iyiyp7lfyHlT1QY/QBDs3n9/ZRElTQMdZFDDwb1CxF5
tq2MSI61I9Ugnug2tk/dmQ1oJrkklJuF/ZwEwNCFYYybwZLFozcxe3Wjeil9dNj9
YAKMaToX3wQHBpHTwslDl++4CGEqz11HJbD8kGoXl5qZApK0Ff/gNBUv9Kl5Q0dC
r+fbUw/7gsH01K1wuwOyWmP0FgElre4SiQH+mBWU/zcGPc6qgVjKhNbREvy+tBhm
bXfkB1/Mt4m8iCxpMkL02sdfzaYF51YS0RAHBnzuWCI9bzOGSfbeoLFuRh9lLL0O
1NQG5YiTV1/O84FO+fhFSR564Wnp18fHkvEFGLe2b1/J3xmQYWJ7w62ddRJPbK4w
i95zyhtUARm7A0s7mB19r7jS3WFkw1iOwaxAiAaqjax4BidYUjyJWi9TMsS6g59K
V/f22WkHB22f8awwhW5xwS8RL4dmJ5OwCYnPP+h+21Dqfst0mw+2g2P7oHcpK5Pq
vjLjJFVSCaL9Ij5Nhb5E9zcDuGFbVP0Ygc7mSx6/0GKaWqaU09or2LDRpTeusmJV
GRLjQny6XkkDMZBMEdNXG20xhVG6KLRyR7FUIuL62rOu5VKyqlJgU8fD1NeXmR53
yYb+yEHU8/SCEdsn2JkR4Sge30/x6GV2AfvWLMCWpGgDAWX8Xbf4JdbUkGjZrF/6
VQRoUuhy7jJRUaVPEiyqX5C4WU1z9hwjEsTDEzuOHOoOhSdSPwn3Igl7BAwwecAm
b/WgZBsN1ub5eq5x7ezIifpFxN5GHMvAyTYtBvzOtU2dsiVLrYhHXfAAqaoSCYZ/
eefLX3ndhdNXXj+m4iEKSIw9l45p0ewRZfXDsayXMIxs/SU+L7sKo3dTR0/xXOnH
/GLY+s0JthWmdJs7G7e5bQb12GAwiFCqFsy00v3+7JfXvZzAg9IF+MoMFycihIGt
jbRgfjtKV1OpxdRny1/UPOruxNOq66quMDIK7mXDBd+mmFv1hcd2DGtPfF68oZNU
bAK4RPENY8JGr/bsgb7qzo2axQ5MWLc2zq19X7YWR17mGlPvZr8uL+9Kqenk+pkA
Coy9iPmOtKz6/YM6cG+kb/kvrs7DIUr9GJSY5McC0Tk5gvpVTPZ8PFBgUBmkT68x
G5WP3lTay2kzecahzIHnIfV954gldI3jvcz758dwF7LfjndsnDKmLCPQtxOwiXB+
LkSeubmiYHYQEk4rc0XfPKKddkCLehSvArdvzhpHucaT32K3OlNdmu71QUT0kExm
pjwYWOui/6NJVOi6TYOfUq7HN5lmMNGbBo8oujOY57GgQIXH65NINu5ivZ7IhlQf
pw5md3fkRbQKC794ufucFmSJHuF29HAE7evMXQ7QBrNUU6A5ZSfClKSoNpFfuGza
A9EbACZOEC2M9ZaDfeSXCadJug5rMdADHHMzyODFLA1AZ6s1W4ygFFbvpNQDN0az
2uDpPQvOLADSxmap8+er9XlyXdQ3SkC5FoC2R9c5hRKMlmDgMADXy+MM7/dTcqt5
zrDvjz+5c6E6K3IZQLVH2caTgCerrEM1SQ98fM9/KJirjyFUOgbAneSM9B8NsYAt
PvtPMxfjQn5AvAcfkLBYtHB96+DZOgPk+dHg6Y3MgaUj6J+0xuwRHORFT4x1O+b7
ogEc3DrVWeJrsrOaLvQcYKU59teTBGlqEdleO3YqoUklOHrn0cUeG7UYSSvuEbV/
XLKfm1ROizb43HL2kyFVDibYWQQA9U4lD7zFxUNMdUp2jeDkWDjYYthQSPxqgjdw
bg3bauwoWBOHa9e7K+yAClZMDS2HAzxAsxdqGWEMUkb9GjIF8jC96BDgqgzWpibL
TsirdgOcnAX0Zkt3bE3mMr5xB0nV89/OF5R+DtYMtmB7GtIGDuorKD+aA2vgnY+X
BwXFqNu7TNgwezMJNIUdSbIuFPO1tuyGOSVnPdIHLj3rYZRd2tiA82yCpv2yiDKx
7vZLUNGEgLiYoGbgdBToAfbT3ByakOJ0M1qCacMou2RQiI1y4GzlSYAYZVrlccyh
t8x2oCb4EfTqkUzoDWg0HLn0ib90LA+bQXYiTQ+QWd1kLhuA6rkNwj46uGJvUJVM
fyU8P0fAZbmArjhwyOgpg4oiOdJIRu8i5r9X6J7DoWAQ26mVXB6cp73OzdYTyqqQ
fqmiBGVQotMstwgOPZAJBxtj9qDiaNASu6xXdfTT/8fERGDX51iantPdFGX/kIef
EQtr3GlwACil1v68WV+VxCRwMJkQZgmDlTNUaLbaHseJKJZmCZ0NYS0J5ERdrPQu
On7bZ9SEMMjMOldV82rsuMcBlkAbYed1/DP5YAWMFaBMw3yDcmXj2jk0MxI7uMmS
zX2hTZ/99VDw1RG7OKGkTrzwYpFafaNmu0lv/sS/nB0ZNNbd/d6SNP/BFXfSbEps
5NQxLTTeT7Ie0HUApAQIAKNSrD75RCY2FbfrDWppZNFUO4dheTd9C2d8KP1eibD6
//7OznhTQiag92lHrkoajN0vgNQGoHtdkWThQQsVPaUWzcNO8LVsY5ORhVBBZwGu
Nyc7xCcKUkC/bwG3DxaJ2rHaMRq+8xq5UGJznicHyD74xjwMXMjjK9GetxsWewKa
Jxk4ELeXogO9FsaWnnH1q6N5RndU1xZFkCSiaQyJsNo5s/MQxFq4NgknVtgstZkd
/8wEdDGbbdq3UlXln+o+0xF681w1YP/3pny2O//t0ivFfSekpUGZd2tARXxla5WT
p2OGFTN03zdy2YGpFcOWj8UJ6EzOj27xOSntramg0xMFbq8MGA1zIUYUFABHuG+M
rHBwjJuMoyGidiWKDAS06jDcMouQDs3CdMEl9jS6W3GXvRyHBgYutktClEUMGRDa
XT7iGpVFwkSij9loKW/hc22cLOtrY7cRzSnx2Y+7H1fbcRHaZ9uLWaTdkI91LXbd
xUUBeufHGxG+IQqodcfO+i0jj5qyxDvFETDzMDz+MEZts9KjjLsCG7pjH+U4Qw1+
93yIz65IMADkJmrXs9uDvPJUITCaOf8V/J3BMEY4P4xed6bOuWCQZ/0sleGp4X0v
GAi8+UmwF19rFbNDJJ4nEMpFp0W58ljclC/X/G9lDI014eh1Jzjrb6TRCVXwQPPW
0xW/HzyjEs5B8CsNzcRsYLdpcja1HmtUhujnhAXQ1KJzq8cUroYUoazKsWfH+eqf
sul7r60DHo6Cx1J8AckbRqFF3jwFfV9LvW0UwgucONmwEn0qyCUi7aonsyrJ490G
nwxxXMSjsqQ4MgnNkXr301mU3fIEVGSzcbxXoPh3mrXCJRJj2iHBhVZ7imz+/1cP
9SqvvQTMP9v/5YU0WQK3+gHwkVTpAxzR1I5kpQKw0AI/vrKvPN/sfJPbeXht6zoA
X20rN4yqJh7HnP4b+HXjUbWYYrPCpNp49yVtzpCkw4fMvDN+QDZwhQToy9XRA0RL
ohCRBvYNCzF0u6d1gkzWGNqIOO4F7Ch0Od4jGhQtW+SokdFM4MyOfdSIz9ht4jr2
iiSJAMqB86uVIHmWr0+8/A0hkK9IosWSkRIDl1RdAVEvKAizZCj6LKLR/OqW9qi7
JrDg3KzDENQE93VoEZ3H0RZPIHMQIan2RbM0vwWQHQVTMPfdA/7B1h0NeoqH4r8P
KlwNdYu0SRTupON0kMeYsQEneftaEaH69zSe7pI2JnwclL7FK1WUnG+0sBEf6Ka9
8b/P6kxF1mX4L7bm7xneA6YANmlpwq2IXBuccMXO2R42Hu3Y0/Wqy2CXmkMooCRw
h9xPFWmLcubfKSGbUho3Mnk/puSckn/r9eNOiLV1GoJOEP8lolECrz3ALpPjJSP7
ozHSrSR57drnTF+mnq6Hh2LcBG3czcWSB+fZC3IdMJ0dqNJAIFCkXiIpU6dwUSKE
LxieHcm+ZoVfyyUhQk9ubRVtIHjB91r97McVbmetFc8ERB+yG7zH8ucBmnuBoJai
p5WygwX1yxCxA3Pzd1ruVNhhvxUaoaTzaDluGr/xKQmvc+un4d5CXGLp/0budjkb
CkbeOFl9t6s/ZWa2heCKzqW0qsFMlz3Yybf953rwCSmwyEGZ/RiizqzBavjB89BL
vK7h3F3HEBOFf6MNnO6gAwVJa9rO+DnWhYNP8iFSlCmRhq2783o8xrEEiJYdseb5
aUEhNnPYPFRZCQoXI2pm6lmBNS34Gq0DrLKBtet87GEghQX8VZm5D0CmOP2C4PGZ
k8/c+Zy9LQ3X3xuZj1XhnwgzlDVsVxst4/Lt0DxICm1iDu+3nbVtl7xw5vczxNK9
3XI028aAuL+7zX+sZ34OAEtTXDhU4EApuMmHCLJ+c8sJ4X5g0RXPfjnMjdjr/8y0
/ZADpqIhmb5PMmSFTgIvThH1uAPRjW/ZRYae/EXdBK8ytIQ+WAz39ddBPq9Dd78g
LFTd16DyDn5iW6bSHoHF2Gm6ESW5FSuexRjEnrj6eAQbhptLFaEoKQisi0yinjA1
OX+E8ymZl2FYw/4ln1Yy8GXUT4UUlAYR4rAswL7VSASA6DcBdlXBkTRM5F5e1/Vr
gQxJ5MrqKEbk+7Z261DQyxjMzhNMqfP8uwsXNoAQWXJZ4Kg8oMzxwJ4zHmtmVeNt
fJlcRWD21rmHzmehRc/W/UMPcxpKMtMeWciF+3q9N9WPCnYEW9eUYXfSkESiGHaf
5hibYB1LWXQe+rIrwk3gPrBbBNH1twFoURW0TVxkmkzTS2zwSj6da4mn4RQ9CAKI
fEReseNaTMLHq6QmLcN8cMAamWZnS8Y+jtwHw+4uo1KZVNjhg0v9XUE5FtZdW025
YhH7ZobkaBOCKFC37vd7GjjiqWOBN0UGwaFVp3Ht9dtj1DHQWycRPrnIjko+lsFx
TcAEBxRbti7h6Ew5liIf588lMt35mDpdM4BQCrjxlFGiuNKsW8pymj1o7YtBZQuv
RHkL5YTVhDUZrExREuQ1023TLBzZTOtP4qFiLfI341p5U0gMbTPo472dUM6kwhXF
JjpqIAGTZ7YNUOTwXVQngIeqGkoCHKd/rkS3WYielGZ8AgkLu4PBQisoiyRDURV7
oIwmw1ZCpHlNalmHnRtux5A0UJc44F6f6g+h9fp7rvZOUoZYSBQWuYbWrleLELt6
chN+MuhXK95s87HzPTkfv1egIJtCveemblnKTns8mZuiH7XrSyETqJ/GK7CEsE6z
0/bivLPkHeiPRu6Ae1IOolfK9LmzudxPl+WwFWaRm02CRBQQ3hG7NF3K1TaxRZ+T
Twij1tkildlWGjKietI3S+0FjS7glrlVpEGb7SwHBWHT1S+vCh0+FxhAgNSYe6kI
XcYiVrWZg1hBr+quJeIgpw==
`protect END_PROTECTED
