`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQXwfIEDOOB/6DN+a7obUl3CzTaSS2BuvMOOugVMvJ8h1XWbVWUpccc1Z76qBg2m
ues+AMyg0IFCtjwZvvo+N6KsKN477RDPUtbCfFpuWhFpWwpjtFI6QnwYcaWka4Eb
mqV8pvnTu5AwrccTSpA24dOevgZnGu36WyLEIRypfNz4+b9ucdal5OztG+z9VVMx
M6QPVlJzyInE9FEo3yaFX3udjM+5pQgjOi5YlLdkMg2+wTdG42iyU+7f+KUloNSd
Gq3tck7E9e3F3ja2BVfJF/tpvsQzuZ5ORNnhOQieCZlpXiczrbh/ccI1sVrLJps5
X3AfSCaqamYjNxTg3nOGApHjDhBIzDIg0LlpvEyRHb4sLGINRbh7Iz0/CCo7BH6c
gWiPvczDotRDdGlWcbYNYGbiCcut47fi6YexMYzEb2ifGwxsUw2cU9SntC3dE1mi
q9xsXNSEliuMTqsEZfZXSVpe5ymZRDtZsNQIkYdUvBzCoo/DNjXpwaJt9r2pixvw
MRdD0ikGMmtQ3Qa7bP5ZUQP4Dv7Cm9TmMWqhNIHXSgK9WxljFTudVplVzCKm74Ed
wfGxgU4kaY6t6WWD6qsmSw8AZM+LjVoCowkDYYApjSz89+3AYOeJ9FoIuttBx3cT
NB/L1rkSfWSDoJTdB72m/gmoK2aTk+9EVPBBjFbF2JHylP0KhXfxZpKyS5s8Se/O
bwC+j7rXoGWEqhna0jmxifr4f0RX2htzNjbFFfyccMyTFFbvav9crHAN4eFPemzJ
bFgQnX+muC1Cq0DE9golwsVqqvOYrfnFPkDcB9W0SJk4zw00hF+bN/ivFl+qe29o
dK0BqxFbRRCAQLad8SASyFBsS1NJIX2rpcWF2TQE/9Ae6jWp4gQODExZGlG1PHjB
jb+Bhp8egkDPAXErBbAxXcBlHct5AQ/27pjulaJmhR80SlBn0Bc6ZbVSSpu15Kkw
/2W09fETJDYqGhyFpkAaxITDQ7nPqG9YBnRXt8U50Hs4nEEC2q5dqcRkIN2HswgI
4y1JEPqDCZwZQjhe5+iRrCTmkn/Cz8XzbECkeqwb6226fLMDf1qSwjHziMmsD1dA
FNCDVq5uDbcq4wPCfaxp9BLzCBsX/UvQljlJvply9TNGRHOIDP2rSppdnCHfczI5
O0f9MLVOA8q3nFNGwNesdPjE929EETUp3znc2bAK0LEdRHCRutF8v3lXq0C2CaGe
gjd5vi+Pg05c0pXxdXdXur7e6OTodhHflDYVT+6aXSincgKQhnH+QqVI3S3jfj+5
UgJHJtccnm/KGuUwFhzlriQpNWWQWpOXyCDlNZjb+HCWQbXNNu8+MuIw9pdR4r0B
LwybBDxhpiMs9BALwYYbBnFa6PQvYBWDro6kjpuUn3o=
`protect END_PROTECTED
