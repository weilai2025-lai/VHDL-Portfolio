`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mcxL9vMiswZl8lz+sIeptCo8bZpRjWz3ugm9t1IhuUXbPhQAghnUgWatHcrhG/4k
CVWB49IphMbXgigXgqOTRf7qiHMbZkOtX0p0KHTKY6L1e/AEob49lS8IMlli91rV
ZQo9H8M5o5E+Fk8nPdVteHbZBrOwcG5WIKIJZdsnnn60kmS9MWpk4LPX8NgnLfgl
Yyj0nQRU2k9QBSROEwvOGx2t1h8Oe2hMPDT3riSSqRHzSXbzrhuD5cSyfMOpoiWw
75h+jtt/QPPUsaU5T2VDO220OUvRGiTNAyIUYxrdD0zFD1s9T8xiN2014rWJ2HPl
ZrRzchSpuTUZBay797txZMaWxWMhd14TeB/Q51efRoldRs6gHvqT+PF9SPXcejaz
B0WVT8kEPTVAmmLZFLNjEgdIwi7un29aX9fOMn5l2EW+77+Yk1OclzW/msEWbfhc
zhWuPWqYwfS/jn2ORaZst4KRFOSyd32kMXfBH13Mrm8qbL9Tz9AYA3pvFXPh6+hq
v+JCTCd/AMGBM5iSAfwmETmECd6HvaK1eWlo5emzSzGzN7GA4wWksUiU2gATPZRM
0TYpbLR1Uf4PVWzBcjuv+ewgfTgrznXgorZ29pR4fIApV58HC/M7UwfxKcuZxYYD
SZEiuuh8GzFFby9zilGa4Hit3uQ4SpMcL0ViIv2NCy3x3Q92iwfJpiwuzRXa23ts
u3n6y4fbdFfHLwEqr7ihu0XL1LM7IHkZyvdWQmZnAykV3DD71ClU2Je3HYCo6USj
pDAo/LLC0bgDPc+PtODln5xSfFuS8mF7S2hKaNuNDFxiSIMpCUf8W2ydubifaevN
lnVLsCi/e2PNfmgec1p/cN42rVGbEIRJwTQf4GzcVS/DnX8YNb6bJWo8ufhpK6je
AKyGIwakMawSW0VZHhimJ5on2eQ1bNFxdZo9LIe4/LCsM/iC753d/mzCG8i+grRr
zB/ZBsLrkj5Ydan1PVGN7WkglAydbR2NVvEObWs1ASlqE5qVl1N4jW+oEkEzwPgO
c+V8Ywav4sHBcgqACGkf41riRYMHIGbV8/S9iuS81zmAP75YfwJ2KHooP3ippL8K
MN2m673KlTaEYlxm9EWJay7aqzFtp+BwPDU5ADqZMhGjONFr+82K9TRIFmyHMDx0
6d7H7PujaeE3zMDs9DahM738fpgSfd2UbG8R7B9THi8l+ph5mR5rT1DTOpsDrARC
edljvil4ZmSQXRAnUpVT5uqL0bhmTQLUEN9ikpanasT6DSicOm2BRFUkuevTcTuy
06pPpXktrhR4x+9wTmztRv9Fpqct0WLCZhx3Qxzeg/BJPPeIlwRxkwoLXcltXCRw
w2ZcdoOvP891tTvUfW+XyFoPYnsLtzHnS9WxRwZFb8YqvdEpM+sy/IdVMknsSv+b
mO511jsSfzoRa+Gsf1+Yrjd/uvpq9hM0yrtmHIOYCgRUATvZtwAwNIBt1JCGCs06
3Wu47+kH2cn1vKdNTxyJR90NLh/FuQBtApahORJwCmvCNQBD0fMaC2y7apw0ry5/
hyJ6sAtftJFls9DpylEKfT2qj+JvtMwIxqNPTLh2a1xOYRf5m6IGJsYzkPRrkFSE
P57SMiSknr+M9xgvsnry6qFSs43lDqQ52To5aqOxNsNohotufT8qt8+iEKYPBz4i
F9ieAtn1FuxAJEyrtiOzYXEKoW4vvLWPJDZQ105YVc+C2gzuPuCpXF34YO8SmZha
0ZcjBmFTFzYOLvWV/gbkZhG8DUrw26VNf1hwxcBWN2cMqLG6ldPy6cNxI9uF2egZ
PoHCEnen8YASP0xcjaZyiebabsN1f0IloKB/xfAGGxyr+Z3iU18kcLfQfSpMOB1a
ggwA4YLI5hCh6+W0BvG4ibRYXijSQ7UGaE6Jy+fvzeQ0eVJUwvzsxkex3mBmnVsc
mIeTJx9I8jV+A8NwiGJAVLxFXTkPDEmAHhaUYRvH2vHDxhOuo+v/CxavoSZY/rkd
kdHW+DVvra02jg/RGGJo+jIq7Wlg7Uss/pmGcuS8okHv1ZqoWgCVCogxuDvMo7zB
jgE9keiaQfqYs5XAfQoxvB1Wz7FPLcHEzLeiXIZ3ReXy+glj846j9YQ+IikJTUn6
kApUJAZVV/gJzZtyGfbB5ZWuCF4RkAnn4ufsyCgIleZeiyy163ENJnOibsreDsQc
JffME1perusErQjGS+IFQ6/KjqAMqSOHM7RzLjJaEsSTM6cnCj/BWSS6Yq4Jox7Y
r9a918I2ZPO6+JkLgzL1ZplLZpS/f7gt+e3F6tsYccpYrOHmwcxZVFhrqTF33kgy
qcSHf6gy+qASRfllwDoGojLvXBidqJZTEKcqzrd3zUKVbeKkBZk82n6TvmIKUw2z
MmLqzvKuP07hqx8i1PSMClgSx3iBnL5Tu6osu6/N4GZFsL3hYpM12CzHZhJXoa1j
JBz2yAKNQw7oP0ZDauh2pY7jOXCz4ub3Gv7qjOksIagehk3kvs0NrO0/A7WMJxHU
rokIMgqbwzBQdQXkx9az6HyJvyOD35Caz3w4+/1x1L95G4B2VfxwoycjKedKK9mL
RzzZK30kGMwqpHaSI+OmVYHJ+SONfV2vX3nY117bP5f5cZzve5dZP4RfMbkYzsuh
hcORNNeGI7RIf0F7z4p9cnsiS26daEhwhaxAuXcysGLJxAqFSHnUCRbcvHcQj2Vm
92PSME2PEoR3KzvDt7Q/E4dmeBbrq2Whd2oeoxcaVMtgCPIncl3RnQVmK5NPFCSV
cfMmREG6o+fdP5cXvW8yp+NChLoHuCzo6b2FKRByGTbIt3YxfvoKuSlQFG0BUDNN
RalFE5o4HWucH1WEsE+3Te77wZdQbIhJ+lwbprdLNj+/zCzl24PoZdwuBVg4NoC+
ph3br6fHsXxq3WsFvqFLbtcA3ew7qpEErZbvrPkrE+BVunMdR2SDZDg92xme/R58
e/5l7ZqrjGapW7t1TueoABavKTnl9Z2pLwkpcIOMLG/aPT/OaXjMB4LPDoucd+o9
2C+MWOx/bbENZA/8kZDte3Fw1IbajQmbeekVdSA9g7BngYWAZlv1zIiGIGFVVyh6
c9TyiYwpWJBkBB4tu2j76tx+NWDp3utklzYbMn+j+/kCwRwS/mmaJtABqF+vbMai
UArKlrNOwm8ob4eUvWapNiSWiNACBq7mUbR+eL7qCEiJCYChYfqTZfqL9lAds2C6
pl8yEjpV4Ve6tiGGa/fvDvJiexQRKk88439mR1LPVOYsUgBqFJNrcZH5hS0hTo4B
50c7aWwL6fTvdPY/mKGx95KLpXB+BskYnRyGUtii/i60do/mEeJfojjXNvhBHKBU
wfCDuQjMZ7zNSjFnwnpA2c2te2e9Tsdydx4Ftj15MfIuae285xnPapebNs53QUEh
EnCs9D6DfTII5Qfxee44d0teEi4RPxEFbneg6Cf8CHtvzVCefcNvGzvJOrsNAV6v
vpgQXrM931Ra/S65VVcMjN+NxD3bEzS4bbe6ygBUuSkquYR0UdOaPqAj/yVJT4uf
FPak8HsCDyTkTQl8LICLccoxOv4hBKtwqUsgVEJGxQPF2D6Zy6LWmwx7cVLRNVwu
WUjW4ALRrWcf3opRtPRmKqsYKTF9vUmF0ZR8M2yzBYfwDPwCcwAngigpJUdmw00Z
3ioBKPOEJJqYSLV2Qz6AknXDr8eAYFzNgs/Jbtx+U5pPelK/CQMugFhRFXrNNRZA
lG/v664M6+QFane2W/Vy/LlQsSMS8MEbLhdGNAQLsvXP6aQ1NvaoPtDwCKGnF0kq
bpnMvAckzZOgc5EZmFDIMWbwLNbQ0ATx2JvwlLqnlrmG0igEyFH1MvKsj0JP/BtK
4C620H5M19RimwStNeZtsQycUA8CFC7tzOQXVJCGSzz3wAg+nPPCARHCKBU4zppw
fJxbnn2kfPEkF0hYUHJFBZrRi6K6+ExZKuiBP5uqAS5B1t85ZK7BFSXv5JkcAsbS
btaJ1g97SxQLwXKIOSxEGhXXMd5sm2ZekallL3nxlBLXCbVJyviWLpUCcUTY/CVN
8pIXaCv2NaGUHvwBNDJ14iVOrZ6M521/1PTPA6K5bYnd+O4nyFT24w+cgagm+pEA
slClNBjX07gn0L5/zeR+sef+sdGsx5/HbRu0X/yYbTnTFP7dZqL1fCwS53rhVPLl
JuIYuwv17JqmUBTAAftYr1O/4HOyE3FTK4wDotgmPlSIV5K2ttLQKzLlvf+pZYNa
kZxSCWRrp0TpaN1t9vUEkdnQbDb8UjHsGWJiY7MV/LRRKP/nybapKhYnkoMG4T8S
dNVTD9xRkrNYsz8XJRmiquUj0RvzKYdGP3xDXdUulswCGe/ubKb+7ZE38scSJfMf
++xP94MT7dcQhrg9qsRMidoyFlaURnbZUmQYMh/R0k34EKLFc/pqC3SwqGdnLwYj
uotBbhgambTvh+D3CtGJzumRj5kKV1QUlc3W/Gxi64RUQ5Lgrgc7PO32QGx1l2KD
O/qVQPbYhENbzXcUWKFd4K8eoCWQblEUbE3PbHZ82OxVf2lGQ9oPFvN2epV5JLI4
vvx2cxRzddxbJ3jXzIOXpGi7Q+AUwYGxxrPXn+VWXEjilH48L3yHxscoQrzF4kj6
PItcQJYj76QPP28Rd84fA2+T7s9g0FHlRStxlBNcG4DUOVtlpDBFtV0yQN66pxpQ
3+w6Oc9P1nvgr2YGn5klxsQfF28vQdod8XpkN9lVpE4hh5RbqkOfkWJYCXMipvZq
LpUYXuD9+6jn7qwfc4/0aSWYUGl2O1L4LqGnW0W314ZkUANLMiOpVmwcBRY3649E
JLQgw4ZWR+fxVz7GE9ah6MVqQphHmgQ2Y0+ayTUQn0zUFnCsMSGDdrN9vTSDY6QU
QoROyX2bZ7oEQ9Rj5uWKNxVznzL64HppYb7LrY49lMab1Kpx7LW2UmjPuvrJeU0E
p1AUtuUahus91hyUKlfGNxOXNr5iTWiFc6i/0O32Qr9G8Z+va+512UcQkeXJ3CxT
FpepriPmnR3+kGOZXClXpOA33HZzb56moHLoCoQgcYGElDce5klnpfzhIcczSXJx
vKKSvPKhDGMxqU/JRdjEs0WvwE3upCHMDOGvQLuHh3pkY7EdEErWGN3SVG3+D3bN
TJkQNNsB+tOo2uQRYpm994/RKKuu8jzPOU6wa4ps9DxpxwfwNHCysMctrXwwCy4B
PoPviBPTXWda5gNYBxMAKUQXE4+D7ZLtMy8AgUIo8H7NfFVb3xK65mcqVe4Wwjl5
DQYIMgi82AypjcBO+OmmFrZeVnTTR2tyNu/sbOrwpFMZuTcFjVc3sHfiLgN+D5xJ
lhzYmF69t8EoWSLF+2uhVlNLBH6Y/zXycVHUmrIFUL3uDKB/hG9rTZLrOqKJB5Dz
wLuT2sskLXwKCiK1yeARhEzuyNqvl9XFC0I6uFS5cA9rPVr5k9iWm0r/sluvDTJo
bcEUhczoAOsQ2eBeBsFKrovq/afvZNyhT6MnRP3ErXQ/Q0w83+g0zRcNfoYnuzSF
7x1ZI6SqAoz4WYBHaOXB//URBAMwPydlI16/AB47anlc7YYOH5xQkkmIHQ+wMwoN
qukPfDJtx78pr7hlbySRl+RFy0Pdh6K4pnTmVVdyM1/DCUHwpAxysrDpY3pYXHYQ
YLyfkGfx4BuC0qHDg1vimL9o4Gpi3g0jPLbn1tLRDRsUYmL5ltpA2zs2/AIfogKd
by9WM/elrBKv4EU1n2I1glM9Ao5omfYS/BPq9ywtu9SfHuwFW/VYaFd/5zFjDIiX
GWnZ0vyBLvFsDDrnqbvb1RMguOY2tiCBc2syfX984NerldaGwF6CgdxOg4WaH98T
3hHG3VuThOwPhlsMdXOF6R0lzHfTuryFoKch4ciOi6sCXitMrZ5ezP3x6ULdG973
8t9dkaJHCNgkv9OHBMpGEv2QwDtW1chq1KHT5pl8KHHBZr9HKOkTsm8IrBoJIF8U
QjsJNskq6kjuFaahVR6QPvRb3CN4v9PYA3viZJ5SgBjAwWYWe/669W5tPKF74Q7n
Pp0LMxrk05LAQR39NeEo5FetM/d3l27t4pheScqNiiLLTMvyM3NxJqaSlOhk7U8m
1/MfRA1jv4om4kLoMVu493agb5cST/BZfD1WeCSMeZ7G9CYQtmGVkDORr8xRaVPc
Hw+Ld6vIZ8imfkCaPJQfSiSEWpAG6oO8IKJujqoc63hzwSUGHWiPWgPkXy0D5kVg
5elCdqb738S6nuSHU/vWHDIPRzUAqiTlNINxMZQvsEmZY+H5OvKwm1PqZBiIxqFc
klCrRFiRV4I+iUatUuauLnWl2Z0dqqK1dp+bAefeGJMwDghsOUy8lX09X76B4iqP
4Lo7+7IBBYL+VVbopN+aFg6irjlTg6MhB8akGc1WEM3F+LNP3NrKr8xzC7dfznGj
iL2pISyaw2pdCscsoTKDOV6/aHKk8eW9C75m6SX7AdmGIOdSR+jineu8CdHOeuc4
J3RaqtoUcz3hi1wh7qQbOQy1LIHxMepdzA0SXb456YOv/UvvhfxZ/56o9s+6TKuk
ptvrAArH4XqvCCTOwJV/yMvv08KqFDVpDQI4tbV81azsdoqnzNjZO682Y11T9nx2
egKWR1PNYUjrefFfi6tXvBvFdpYx+15512wmL4RXUXZGz7DIyxuhx8QiBfJp6PCL
j8kGvnhMwYz1F7q+upVYk3LQEKFtleFo6epcZ+Gyt+jrtWHSfZdyZBa9Ama3VOK/
HvyoXA36IFMS7uQUc9u5yEJhmQs6ii6UnLqXzRIa5/z8T5gubaPZEJFiupkkk3nZ
/nao9n+hcX7SU3RIkVbdqm4KUnYxhttKFv+6qd0S4YVmaktMbcFVuxg8BPSEwOy5
w09Fp4SPe/Hq97hGO7yMFUUqw7WP69ZgZ4/0MJ7kMxRAyxFuuvslMByKAuSSnwjb
ln9vBeT1VpmcLpgA8nCAkhs/MPd28lFxlb2RiGwf2YzPQSGJ4EsFnHt8nLts3v9y
2JltqASuyM7yutU8CuyWCdx297OzK3Kw5jMGw0uuHqg85W3/WtjrlrOvF+HN72XD
RQf4gahlcRq2yCd+teTRVlzIk3ChlF9n5XZBCSl8JqrvAE8Nz19TpxUHaeQSi2J4
yUj8CVxWIvt2vHrlFfkFfrz30+QibSl2GheeHSn4ryrlgEnr2ULAHsQW3bhOZfG5
2nLm2TPe7ENWpNFGewtAL9d5rdkllYa49XmPYguQEcB8oYAbxrmX3rglyMLOUJN3
43KN4+Hs6pqj2lhh2uh0fx56LHjaFfccE45wfqzhNTO5lzR3KbynMJsgi5WAJvBO
hfX24bawaB/6F5k8gwLvhGJtJEGzbq9XgpEFrax3CJEK7H500XNF3R9Y3TUGApqO
U2+2cXRaOiGqRYWrPJhfuHnYmiofbc1Cz93uo71P7FWHPMnBYGF+Gi6i2MVy6G6L
MQ/p+yVx/D86vlzx23dHNSYix0ge/SmoSzfnwf6G49SdAlfx9FwYabYJMiVn+KK8
2R/pmQED81HcKhykXwlyQvdvzcda9x6CNZoOY0D8avTREEubQh9ro9Sjktm5xdXe
B0sYACuLeeDyNaxbqXay2ZwdeX4176HqekWnvlBEAKvSfGYUMt0A9J8ED1Hq/0/U
NmTM1DyA1lf9vIqvmgWzcW+K+wobhrAx/HXYnzXkI5y1lI2h/rzS4xkzkUoz32WX
szlMC88IbptHuQmiT46mKYpWzvZYhX0j8j8L61USpD1NXI+9sCG9n/lFfU5/Ymbt
rAlz1nCjLrKMnMGgfY/2xsv6VeEMPhJmdmMUjoVX3fUb2OFLA8tAvpmrgxfhStay
Dm+xKAujqKgJYbl6KHV4cVGmoDqkkLCd9Ibu+ARfR517e8fsfZ6vzYZ5IR/d+ILj
ht4GBAOZIWPLpyumJXkRe/W+aDAmRFC79zynUaoDT2ZCMOz02z66u7dl8lKYvkYR
wg7GxfLeoJ6wM0Misc8DKN6hOJAc9JBHl0r64rIVUbMuhdSP8mQRHizjoi7WExVx
TkrOBTqKstzXzVl32llP1Ndj4B9jbKJOBBfZZSEQ6IUfHqE5HIaLRms3Hkt4tqOr
sBLPJ14D8mpitR3sy5JL+Liqta908SdgOGnaDgfLDFxS7ULSRwR5BSRYxPrijoiJ
U8uv+cFzV0BzxOxlmA8dJriiIz0TOJo/75+hURV+b79dyvmeOZsvXpje8SAUDNny
Bi2LJlegocUCR+j42CA9diXI2WcuQgIrQiCei9qkbm4RhvoqcawJRmjHq4FqXpKi
7RCM5OIEHyOyLmmHSdgw/i/hqlbBKaJ19dHKOufhY9Mck0RPjfmnQ86YZ71u0q0c
GQqgsiy0vQWP+w5P+szP5v8q+Zt4Y4z/bo7nFLXr6MHW6F5u93/z7HIxdwS3T6cU
kuDTi9nKjf/ZQ1W7SuNGw65l4hvkJYYuq3PaNDn2fR2SMBi/jO39Vd+3wKKYPRzg
igbZQ9pxNoHlVaaiiPxYFQs0UZy08W6GktKBRqnCtk2QA0GCk1mT0XFA9khs372z
I7flCgbVDdXU0fchB03MHGCzli3IBD9KoR1GWsJbe11/MeBdkVk6o0nuNeW/MM2S
ZhJTUtFVAyW3uovtRINbeWkcd9sS3n+6bG5E/IpDbOT7O8ELIhjf88NvHFAt3B3Z
ePLYObBp6f/YDEZJvywkhxQckODccHqcxcnY8lIZvt3D3fqs0WLL1eCinvPBO7W8
fv1U3OX3CULM1L954oDqDqNXCsxaR6vLm6Cr2Nw5sGADAbY9JduURRUvsiKKHRog
Xc+sQJMgcB9zeqZy2yRrRuzv2aKMTJ6WBiYTakOq8SK/TBUmmL2mENbX093dArZq
4xDaCLh8aOEKYISMX83hTPm5IeCRWUuyI2ofwjBH1HWhfM4X1CN2oMVe2yCGX8xx
dYgXdAD+3XynoC6hxRzZulWKzyQXaXXhesgliRhftyGG03AJL1NxjlJupqyQVLt5
BIhX1AwBlB7rQgClINwWPatmhT5czaj4szv9FdZfRajpopr+rVvkuoxEwysWWcIQ
OvgOL3A7A4t6AoMUWuan92qww5LrdcgxZ6CxbnrFj+1GQ7cDtP/LThgzu42pJDIW
WtQ1mx//pOU9IkHK4QPRntmxnHwvtImVdQz8IWagCd+XtVigmMCqtAU0CbkSJoAR
QdASRKck5u1YdM+u+1gxbohwy/xfIDTlazGl6t0VfwkUH9qlaxmimlucN17DqH2y
ilDjjHzOqBf2cacLJJGCksgnKbVxEAdH0WRabT0FKw4/oMYDw6D8nZgePyIhBgNf
2nSgZuXW6+nbQ6gLJG8+L1qMFWmQmhTcvGitOTcy1/26ghpA8guXXVX/fgrhIW82
kkOFbtH/UYOMNsFPJ69Z86aQRy54bcnAMTzLF3XowzRbdRBe9eLh0f0L7Jnk3X5q
pXEYK7PvUhJE17Y6vB16TSGAK8HU9edbOEJBh9arN22jwpRhdEjzBb1MhiN2QnJs
Rodrd0MHYiWZznQI/lV7/J2gEiB5E9jZUiJ4/kigs5M+sE22Vb2nhEmyp31K1Mjr
rJT2S2MkxvqUlOepz/0rps8zOoUXdys9Rfr6eNKs7w3TaQrXyzbLod3qQxsCpp+U
tuqIsDbEgUTp/lDDvN+EGrtgJd+v6iuIakpkNOxM7RNy8o5tmKcrnq1tHAheCWOn
hGCwfl+7r6g9Y+iaSU8Qhe4kr7NwMU2N8xecGQMacbasK9tTIV4ovqoYjDzYHIPX
RZI9vqOJxuEHnf41MkTy9e8210DWFUDwlPfYs+qINGY45EPRCf1F6T3Yuf+CJ74O
dWzQ/JDfjbbsrFgxyTSc8+don7vcR7qFrFrEZe0ocCI4mByHAvQaCifyNdVMQIyc
g0rcyGPEL1EFe6zMHzsrvxE1mckgQQJJqrixTjumzi7d5WriKKkJXqJOVhXiGddA
+l6FFJyyy0evPm7v4XIFhKvrho3ruligqUtCCNK8zMlMaxlMvZj7DKso889VdJ0L
yBxt/Ad78AmcD8kkA98Rt7u1JfXeC2nthln4jX4XQ/JrxhyaQOPqb48wJsv2d9Aj
G44iEbRLM3FhPpP7tbYkhdPiXlG7DvQL++6p0KnOrZLQ2tDS88L69Ozc8vf9vtMN
MLMDKa0f0NMAJoROVDe9dq5v1ZXFJJQtntwm/gUARC6cS7pz117AVuVi0s7H1jgN
b7zzFW6uu4r11D7YHzp0CizMvEE2Tifabj4Ed3pMkZrLtA4y610+6mf1SO/VzdvK
/5zFvQ5er8zKQzNF/hNJ0eSaGtvJlfVNq/7gX5ypUJS5q9RI0p4CPmXqshlvIu35
AQHJUjGq+fM/19dfq7JhpJdsVu1nJIdbr937e7qIzccWXYJcpqd3HsBcK9F2/c8X
DoZkBiSxzFrdcFwoAm1zlszG2dlhk8cvaSIWFd9ont2HkXlpjEJ9wyM5e+nag4qZ
d34mMOi2e56BxCrw/wHl7DV5pCZt/Ie6ZBt64xFQ3BPaQNdPBxgZxfnmsffQqdWS
OfrM1LLTm11l27vdI184p1iVHF4Lauow8XOt7F2NZ6WTPkpPrcCj1ld8WK71MUzq
IAzGD0RaXl6r1fc4SNTgFQsUY2mKDcSsA1x601V5C+/lHQce7+mmPbqQBqeuriRl
Pumtz63qWAX9H9BTA1m4AeagakiIJsx4Z9d54wNofQCadqoQKKCl4TMqzfvTWbYL
R4mzwAHoZmwHIihUXfOz3C8K0rGcoSm+k/rUP9gBSzF8ZNS+nwVnkf/asowH68tQ
Bh3IBUZXYMSeopcH+9iGO53cA9hd0sg1mgiCg2o0lVvosNa7Fzx7f6LCuOKAt0Qc
D+Oh4/zo83TkCXIMyvs/pO23xaJHjUCn9rKMNyXdGd0=
`protect END_PROTECTED
