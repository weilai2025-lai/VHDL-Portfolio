`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zNoGrf9dIB2hJ/BjT1ZaADpyBSEC64QbSAsg/bjOugaz/etCBVqIW2FehnO6hjA
1uGLivZiwMIhIxoUksyLGuGl3selZL1fjKXoOxoEidvAPdPpGiWvwk5qiZXQVtmN
U4KU7xF0T9pp1Ml/0Gb+ZFQvrnO7atOnISBmS+g3EYteHzNeWoBThvii9ONRSwI8
QlRsFdCOlzQx1AYcnyMB7ZEwvWuwhqUHbmQo2QIdFrzHCir6ejNmRAcPMdzDPFlA
py7O78XAof70BAvp2iYXyfS+UezNeI1Bosf/3vdHW3P4etG/cFr/ylBMFxtG4wB7
m3EaWFTCJdiIOOWsx5JQJYAK1ZtehBYG383lVx5mGM5KYZkGvQEzIAmawXk7BANe
4/dam3PJJtUUSL9q39zcBe5fXMil9YzFj8I8DjwPEDuxlejzWpmNgBRhOeTyF2BL
IMC+ESFxaVM4IVMUVtTLbgGb29xZ8C1PDqo0xoFwJq9DqhzHE8LkSC5FU9YZFkyq
`protect END_PROTECTED
