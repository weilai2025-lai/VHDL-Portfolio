`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SDHrrZuFo8DAi855P+p4Y7H0bZMQJsFN8uK+gDRTEWxezdmXaF/QfX1P3E+Uk7v
MW3c338IGaDPJ0bAZe4t7Q/4yat8HL1IXf5OtbEJj91iBhK88WnMPqX7GasQ3MJ/
vhPOzVzfWx9dS0YywHIou8qFqXcp7R4fZ/qSm0HULNAFCD1INTAMWugUWtZPJhor
5vEjfVmFtx9cDClxTKMoVYD5b+IAohF+FDYmMOhl51rd4nJu3K2N7uccN0JsIoQt
x40QRpJqEiL8e4OiSrwnTumvcXZlVnnR5h8xX3gWmbGaZt4gxqYsCw4C6P+ByUU5
Y6ssGmmBZKpeRn40ppBK8h8IEylDK3KQ/1XXUMIr7dCtSOtssEvdDWgj73mgMisW
7V8JOltR+Tk/SPPivt1clWkR//8Bk+vXJmIDjpQnuFut3FsuJWBTDYjiRNWZN6N4
c2E4jPfhc+Mq/xWI1LJ7fkRWiZmH7FGUaiPQVKc/9B08mgLmV3FdqyZgGVsMwXwi
em9zixcCqx4W2H1uirRq4qqFpmajeyVzAPG3YwFLVjq4uQ9bBESqHKVPRJNmdymm
E6Kb6I2WIsQmgcSKrNW1LUNr26Dav1gBOsThCeo3W+Kyiy1tRiiD8/K1MyjDuG5o
Dkwu+dZTVxM6wRFSF3AzBYueWdmAxuJURBl5Huk4SdPB38av8GDZhVGftdQatUSz
oHYQoPcQ8IVT1dEsJZDxfsMU2YcMiQ+UkG2vbJ4SKMJzHGOyyehUmP+fJFfWK02G
7mg26dveZBRk2jqdke/XVa+v6UFE/ooRkaZ0nfVseSFMZoqGKfk9A0luQWz4J2Kr
RvND6Nt3hU4W+YHho0iG5+F7qtnOcWQM3E93rnkur0VqPeQF2aXZzTMW7snxCw2V
cnyjRqOxx8JLGWe1kQbvfMYeFGR0Oz68BYZE6JLSRmYGQ09WzFSNIEEkm7oB55Uw
wwET/CiG2phCf++ObWiaRK+os5RN06YI+AdpZpMZ77ZE/CpNYCl6nYgFufL3DDhd
H2NwHkvWBX75h0ncTKO+fm1dqvKBOcbDg6HtbD5bnqnaOOPlNJxdgVWaqQeTLHmj
3lcDmjY2u0phZ8UR9duYVe7GGRUfn1KV2T48qKRxFahOdJSGTmwlXoi913wPJgQK
p69mKAzhgDkFAqdIuQY96m0kk78qIZEMHPRKnkVCXcD0PHQxPSbKRqNAJA8rOPTL
YUxyytqOduzDyGqPWBPsYyhwWp6WIpDfdE28vOsAxitndyw0z7yaJV0SSefgigRL
3gSrwKTfxjHRYKeodHjFvJQ+iyldKCwyaIOUQ0J6qL2LtNVRfCkxseUd22Yjf+q3
kIJWK6b98CwQZDiM0ap7EJNupmyqFoVn8rdKicPPqykvlrQ/hMfrcfgZsphI56RT
qb7adbHeUgOrzKU3tu+NXgUno0GnSob7YDPWelZe2ofEuvm2iPK81EADo/O6x7R+
eJtiVJhXC9imerfmTBbcqKjjJODHOlMPzhoXRZCQsoIKBuGrDUN4b/h5BgD/aRdW
PaIGbbhRW+SrmjppEs0VajnXvLbqZ+0AkTDXz15xN25uLKEkSeEzt/e7mJUWED/x
18/30Lsl+10mqJ5fqkw7ySFWGDzZQ+RIx1HRZC1qUlAmbSB9igZjcycnSNX2FClb
a+vaJpCT9oyO9Nqhd9E4uWEPItTuzkpStjJJisDr173Ff0/iEm9AjVFvOQbfEuQj
2fx1GiXA3A8iNI7wtEkZ9H07V0jWkHoDaOq8+JZdhxZVzkToSUPw+/CRm9X3Urdz
1ZpwIMUy5eyTXJi2Oab0E7JspkShRSr6EqQdeVHcxeYeV8p572t2DE2HJ+epemjf
yZrdsBlwSvtiscRHeNsYL+ZBY/lBeyo14jdF2Lrh2mhqKgFyn14mmTZEABCvibAX
67yo4oCU4h/XAqRURjbtdRG9g1osmOXBHiRpWW12s2TR3agAbTXn2wDeYTmN0o2J
0mPTAt2Xgn2H8piqd1C6TJAKXhdNOOlulxgaVJULfxzHgJemHcoZyAWVHqDOtulJ
7SVpVDIjfttPAtMYDjSYOzYeOgeiakmPaHjoY0ZvddiqC+mKv8Mt4W4F7Ww5haKn
AjD3rkK2OAV56eTos8sb2lp8NbcFMvSiKi6rsmqNhJwePsghC4MXr/3TxrTuzynT
fhlg8HjfAJjTASOcNVo4AYYYOJnoK88uvLldiqBLPe8aKoU3tLvnBx+OO1oStV3Z
405X7KRiMZ4/mkW1pzLVKxVuKwee61IvPab7ixQMBqq4YVaRcV4vb+z/DMLbScqJ
QXhtq7y7a9rksuHdO4AwbS85AmkDLn57tC4S0Jf0NKgy+NZJmdKyMPnHQh2nJ85c
aX5KTu2cndzeMLH0+FBv8IH6W10UPjGI1FhTIwh3sjRMSqSvNS+5BsjPgffgFD4z
WK4Llq46aq2nXFVp1OqexxuxbgF+qemC2xZN2oPfDs99itIc5uP5ODz54P21fz3J
pXV+y/wzPTdC7YcCtMORCc6oMWC5yVXtr6yb0gPnOHJRHUPbTlDd90qRGberivQQ
2VQU2FPyOUPzmxwrp4Pr6CEwui4YcL4YZtFB5+mD1wpACJtuCEhLeStzRxzW92oo
5earAi1ee2PAhE5zncPxknRRqL5+WUHZN30qFIi/A76btUrVk4s7+ljplEAQQdNG
1CzxlMa6Bt5R8isIZgoBZilzr7ZN1s/Q9Qw8z9VHTFB0RJwzKHroDrL3xPKqjFUt
ePlgz+ONNH0W3DrtVsR9hweR3w+Ztuf0odxcwtM1utmaAb64hzaNHFMscsFLaKak
vN9sqkNlT1EnqsEajw8ckPz8iHx/7StynKGMPao8pGr1FgGcYBkV5LFdXrWuRWrw
yTL71vIxVsivlCcjLMYF7IEfVIw0GtbwnQcFeIsFT91bNwlUGPpdZ47173zQN42N
jrqs7XSCXIz73foqcfLWuaZqsygPLjDDY7+BTS8jI7XzerkY8M2SyObeB9SsssHJ
tZnhaLAJwkwccQPUh371Fj/Kt1vos4rSFD0Pdbst/Z4UzvV/92JmZvgJAZCPRzRh
A0EIGyHyCXNy685I6FwIJXv4IRoHbGeTJAg7EmJ0H2o2opDbP1iQsovl0sycjDCX
qWVYR7u9JO6bqiqlD4kXepINRZr3AaJM1u47uvhbgieHUI5kFFW0dZFDEx7T/E7Y
D3CjitnM2h2u7CmvhbxZ9/yscgFj/eTPANCWdquzN+rNptrdkSJYWmFFoAN4aH/v
M+w8OYPZeplT20m9Ne87gjVnsngAGOhnhokFH7XTL1UtU1hJLCCYf1Ncqj/B698K
cAmD2dIEQmivvYurUMkrgtyjem5VxQ9ODgC3ZwRIxJZWHUgI+V6llgNC6l6wuaHo
vpKNe1TYx8UiA/noyuHCqpQ5AVUOhJS5QHTjr+/bK9xHtflgFxdELP6rkRl7vg6+
bxT4Bu+9nIIA2NTJDJ9yMK3lbfk5S/Pl3lN/p69/+O8yleODGdKddSBCtnA/8LAJ
O1LATYWuLzznuKm0+/1kmqOCCH28AD33LDtyJtqHl5/AZio94VpsMddDljCuxMf6
+aRefTpuhIyvRHsg2BhFIsZusaWC833VMW37TwRjNB1oMv6CjluTDw7eQeJ/PxRv
Z4LBIDV6AAZnZRp1WQUlGfrA6KvcLa8vt+9N/3fdDDf+j42920ljYOBmDDm5nH8R
nuMwfFs5jIGJ6j9fZVfQf8Qe+nD8KjXALmSmpYN4gH44TrBqpfdxsmuTzNHnqe6I
9fyWtWRynz6yRR2mtCScMLyCP1gdD5irgpP0WU+8pafnjkk1r/Bgf4PKte4XrGgh
Wqgz3RHJG5d6A03B9qBpAiOF/CSEZLCbdqfz2d+UzxoI1LSA76S0UMxKv6NC14Gc
CRJlz2LQW9TCc8ijlElV5783awWT9wvcdfYZ7cngWulz0qJEoKXTNCh6F0U0wxK7
P1PbCpcER1GJ3yGmMCR2EZcZK59BHVVj6hTxLCB2ngqxqughaOBzrcgtButsS8vJ
6nHrJnNlurt0TGKl3QlmWoEogjznUZnlr5UFUv3SiGyrOsYuYV7wgraKjo+0+3x8
5Orf3T5NPAioD3X61IXA+IMmJgtJ9K+xKYp2iEd6xB32/uq/h8ABetHuGw97RHUL
nqgkAoL+Hdp/qZf+XjJ4uIzcPCoaM7gFbYBiTLDOQQ8TCZEieAN97y5hdi18mrC2
YIZjkAsdBVnFVz89plf9BUI2Qss21LYE1f9VN/uR7YRDtp68Mb8iio8i1e3MZi60
iNX7pvqxLnV0nCMtELy6SzdLdW7Ep1s9/SU51prAfXzKFeTRSWrx7B29iXCPsqIW
SthUyESGdjppH8Kk5Qt+QTlQGzDbdRic1HHhDnEn6I/gdgQHrWmbgXx/qLaigj9a
j1lTeLQwWpZhZWjCBhMhD4c/PKynCKniE6Br027VG5/LnRBovhFTwmHQ16wMuVd6
WrFEV0Xgzk1qvAihMnRZsAHKdwy/6MoqfSxG8bdg510t/2MfT4OqAhK5TpTktLVN
4ZUkzqeF9gP4zk4uwgP/WBpo2A0fdVRIUSD/xJThLPYj9M7BryDldarC/p0fBF9K
/9TZn7VYhaGn7PJdEKqf1xOvP37X6FH97FZIwyW93A4bQ5BdNDtXuS09PpQOTpNt
QniGx6X4aAop1TpKY7QsGTXWz0Ls0LV9ZGKdQFufGLGqe5+5hj/WUJFOFZ+3SWZf
H1vnEYtWah6GewWCNdV7QaYvMOXeAPSgSljXzsnnNVUDLVb/7TQGm9jLXcydjWIc
ctPVPHe0ZTWcXQz3LOespWe1wTYwm9OyH7/QiF9O80wE11QdUS3vCSHG+SMQPogw
XHIOnqLi9Sy61SrweLgdzb77XkPCuhepR3+z0IcN5HuVSmKbG6e1AvR6B/SyP2FZ
xjzjQR3YKX7KIt3OloHk4YI28LHFe/fSu91KeVYiOv0srU8iNcZZrT/mGv9msycu
0TklEKLvru3V6Xm9jtCHbZgmQ2OgkN5CFGe1WjnjnTUFCMKjQq9bdrRTN8OF6/BU
xTQ0UgbaO65B0ffHBhHOmnrS1Izga1WdM+fuXn2IlVCcyo2G5QyuKRVrWRvY1qMd
zYfZpevetI8coPObPIDex2yG/H26O2lX+Wf6WejGB0K9qbA06cIz+zRBl+ilFTqK
xLThrU+pCnzhBJPd2lJVUaLbQGzYofLd06v9eEOkBxysHwQKORckqtfO9OD5dfus
ZY5FD0XC+yDh8zt2upWx0v9uZkXvdH2kGuAJj1ca4ekg++hLcE7Ae8529Y7KdXwf
W39rN8UqgaKWfzvbbX6GP/kVzHZE14Syhrdpqn7mAAnJTY92TGcO7vA30to2R7yX
F3v5ZJdfrGJel8fr6XrxHesEhboZ1x3/B8iPnXFo1P5e9VxYFWaa0qkAybj6psyR
bjOxAzcwgy3ajbbC75w1q63tUtjE5BY98NLykonB5iEZqhK0KjkiyzdujIbO+E3/
b9ylEu48t8DIclj0BznnqY9unP4H2ldTMslWfdIX81cmxRM9ApetVxX00JU7fERn
6oo9FoCEdM9LH0jGf9SYKv0vr9jVZXoLCxX7c7AGeKcB0CQFAOXKy1eApA5kzZIO
2Y/i8+6fJzXtDSIsvOhlwjlIbWsp63UaqQmLTEE2c55gPY/38HLkufhmsCXpwKvZ
VWZfqjBlpSnUllK4QY5Lo8Xd5u3cVtYmjO2ocGneR8mjELmJBGveyqaFrSNermPa
LyDQHwy5yOEZ7NtTTOz4A9do9n3iQ3If6ndH2RqZT+T0rXQYS6oDn1flC0ZAu023
YkjZqbDxc3XXPNayrQOCvrusgHr1WBImCA4iRw4zT2jp2Cmk1vLuIaLPXOfk46nf
JI9vVQOjjcwMe6BCj2FgAPwREskn23oebC6YLqXSjDSBN5v5/JkkRbIE4Z2oXwsg
imloVJAcNDEgLaC69LZPUuRuOIYuvxxhg3/J9toKero7hxUGtJVXQWORGitSvIb3
`protect END_PROTECTED
