`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Frk5zVt89lM20bw2aLiz3dABE/5mW2qCfgjPxsYQE1R94FDViMl5PWiWIRKsxG0y
YWhFQLAeC4eEg/85LUSAftQN/gmIEkz4yOY+S7pUKSuimE7qni5Lu6FeIaGjn3+R
fZUf9fN6nk2jb2a0fzzMz/hhsZIa38MIV1NOy0KctkBcskufhD5zFrXwLBfq7x/t
Pj1bZUdRo6v1owE3olaNvzYkvO2voudWxpg+qI0Fj3UIQbvinWiTpgoQDfEuwY80
N6c2FilNNCygVGiBfUubMfH+RTAmXsMwpl+X/+pP9la8OXGsVACLzgFq7t1pOmNO
NeaX6LU0uiNuJfmgY2ZGq/Qe9xij5FDB1neaHHje8yJHQawn1BtEFKTNrHacHfjQ
30ZtqGcZs/DiD7ZGZV1scvT83ch3fSzhgMmWrfwt0fKHASBne1s88T9dN6HlB7HY
89O8wM/e50os2gOix75QcvjwaAbet5y7FgbriZZronUofO89rqUOSmp4rLnlrBWQ
iw+On88Njk7yYBVAld5gUU/QQ2HIDkCPziZLMswHAbbPXBwOj16d7FSrIsSMTL/z
qaQnD7rar+hBha/BRUW7jDhA81fFmYb5FumhzWNPlDHgcu2Q4l4s1eRt1qhrSvEt
FJhHC8EJLEwX0sfU6J2troTj0gQlByGlOM+rAVHeV5ZgDPxqIWP5mD7bvWbuM4/i
F1kXja5o47qZyTifWbm/l02g4cEuFJCZyqSaKfNEI3qvxuxleuix077Vl8WWEPgc
M068gBkgN5SjG+6+3gPy/VnQWXH0yawpXXgDVzR4HBu9DLlxwIlA6otHJooaLLKe
ZYOS2ez81u7A/q/M9KqdpfNZyiGmfVl6wa7U4syT4IgEOZC9UnLexxQSZYpk257n
JZM4oGAGBHGRYms8Fquh/MD4HmDp2XnudLXQLevclVLzfVmiuq+Q2sXBp8X/cSHg
dE6A9TfbWLX4bvHrVH/5Z3IEgilqHY5o27tGO7rp6vBqH7rYkg5eCUcX7ejs8Skh
88O+OBbiVWNWhLyWS5oOUUpz19Aofc8JD+qkKHybUMNFp2DxOfi5hCChpitMDWtH
3RExeTVkMogJk1gsOv74yGxckACsdrmTXQiKUTi+AXEpTF4x3IPrBOWvQWFWEH0B
aneNYyN3KlNR/ZHc1QBkr0ohANz+B33w3Oc9rkdWTLmS+hyXZJB+ugg18WAtkTCy
7WOOxkpi+K3h9e6iHVoBTIlfW3OVQqczuprrzN4n0rn/pOKXpUg5LN+ZkkIz0Oux
1I/mGtTZON8XaF/xLP6Yg8EZJntuQFzhRQvWhN4j3PlhAO4XSW8Fj0Zt5eDiibUi
IXh3oly3ZAnAeXSOVc6wmDoZjhzDSA02dePijQgNIvmjJXImUnsEeEq/8ZP72je+
4ejgD5fXmHCRzJ6YPH/T57Hj9kH8cD7unZAFNOdVJFFAu+v69uVSuh+k1en+jcG6
XBkM/fjDvRL15070PmMVTETIj77L+ckHl7vew3j/WCKJWQqt1brtyldb2C2x0s6S
P9WXTDzsbKehjaMB4Oa5TUZ3r21TmOjrRbcH29sYzlszbCWcK8Trr3wKSxJ/0+tl
RYOmQrWyYan1d2kIFhBa4jTTMbtKO7CNvUp2v/V4MbcaS7xrOobuuSUNucOe8Q8P
7MvjQ4l/Wx9X6HC1hnQGAVYAngq7fGwJmdfjU04GmJdxT76Zyw7ZNQZp9sHlkdCS
WoqByq9HzzmrGVHxf+aXIil0LoX4jlWiHpCy0/szqVuojETo6t+1w0MA18ztpkc+
vdT+2F2fyVHWL0zyQC9M29Q9Ok1eD4AtnwkIQPrKDscvMj4Z+AEw3RWaicSMnox2
c9lRfsYf81T9/aQNTssrWbP5WJQjOoErc8u1Rg/xSeJyGBsPgDmAJHRxESO4APPh
3hDBB+b8a077YNmRBk4bsNy6+APYdQM5xjMl59OBRqYvGav8t7sw2NcHrjpTWkhq
vqYBrQNRCGhIaRLjchWtyjjbDlwx3rDhFYuBHSGcr58qTGxOmAtTn8lZQJkH5HUF
eMFrXTpIWnvGsp5zuSKXuXjgG2BcRQYDRPiZmcRVtuEpk6pVdl/fZLy/wUe/+3r+
G55tTTaalEDyf5vddvbdjh0a0JYLHTaf6I5lp01/z7qKjjb/r9CisdcxQhr8rSHc
d7yQrlHX3+K2izRjHkZKzA2E6eqKQK10ztE8vKVbVWtT0mAPY6C0jGUznIPfYVkB
9eYBRt9UY9l8MvmELR+KMRiNErzEKiPBldxDAHANaa2sx4s37xVwLjcLt0p16jI/
NE2gpi84QCp/1u/J3ro53zOTYmN2QaO9M4F+Wm0pypL2Z8OVjhgdieFTPmhY7al3
DEYI5fct1nEChkHxx4ASWNCgNWNAjKyUTzaaxwMpNPpp8yN/a0M3TvWeNd+m7zmi
t28cmWavL6C4dYpWJSeCSWbgayUaasSBuXo5RWUblFL1kbCAm/7nr+aLwMy4hNRE
BmO/qCBVXoCczQs1QdslNA==
`protect END_PROTECTED
