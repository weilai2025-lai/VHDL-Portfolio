`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFDSZ48jzUU9hYfOqYORw+fgN07k9Gx3y9Zj+iOFPK80uD/FjdSN14iwzq/e44By
0cB86XZT8QV+a7SMmMRZtMHzBuw0xnTEZ3dQdiEU6KGVjRnmn1BLJ8ibW9i1xqC7
PbcUhPt0Th3fq/R1vWyGR0WBKfjUOIPm8CL5+PKRkjYqB1v/uz+3G/+7eXQm6Yb8
CWVdK+CrzV0BSeVLXqj4hYu7OHJKfE7+kXZJhaC5irz9RC+lqzwIqjX4EP8cI2N0
qUPsubGzRLQq5kWmjf0nuM+6e/H9YA/7rVCFuWdvoauf9CimgECvzzZRCiQ7uTQz
EMf81ihqgtHzMVb+Umoe620/YB2WWQIzC5tcGIDLN5IdzGz2fJymAa8VxlhbeWsV
ke230/9Z5I3MtN2gupQSAiCY+6FMC6TAUZ0zfsuGpIs=
`protect END_PROTECTED
