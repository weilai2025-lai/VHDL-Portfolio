`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uB46tTVTyGvwqEpT8JW9crteq0H8GTrZCrA9LE5IqmEg33zK59ukkJ/EorSLy+fI
uwHDp054lvIYnoW81rYCPTfqg6MUd6L5o1n5iQVlRELV65LbbHj9VdJhijtCxspj
dLouYKj8+8VMFllKS72jf7CnQorvYiCJFvPUMXaQdHLBPKjv9a+uIIjXAvkB6KO+
dqOgcFCBuzSDstuYEOwSmrjQawFsrRIVFrGM8gq+rfbi10aQ8m4yXLJ696Szlvfn
1Y0mz+/FES0Pz12uUwADgeGwm2WZNNm+aXZXbh6wIpnjAEPk2NC3hn5QG/hpBd39
TOAw5hSEwLX51KehboXvEV11Hry4Hhe2bg0HgQO98ZlfhEwq5OdQfMlLs8aXGzXa
lybqhHkwJmdnY2sWP5WM8HU8jrggLhc93fCNap50r8zteQcznNHx5Nrbo/enUO4A
DQa3ptC2Pk2Dzkze+hhg7ufC38Ud8tKynEygqIA/7+b+JBitcI8YTK0QG2fcoW1r
NKLFEIkjQ6HpIsA8hKoxnCM9UPbAjwU4HMqgbt5r2uQYb2a4w5hLAyc1SiaP5M1n
55qM1TIfWpAtMoF/YKrEO9F1QbGfessMoS2rX8w8JLYvisOBnPBqEBVTZk2Cv55Z
tenkkQodpB3qfH8q72DOk5A4LjrJk56+H5uLQ33D/dI7zUOBL9CJVN1Ed3xEjIAW
fiXCgokj8xS+j3Nw6U17lgzDWnRt+jvjiZaAU85UxKbxXV43L6bwy70diUBjJSiT
g5qjLwuJeWUOqwoK/2An7y3ygqjFpVEV7pwu6h8wPZO8OXKE5wwOH1T+DKPUx+qf
aN1q5lWLgem7U7JAaK4+t/xNW/DTIQAEkWww1vuPS57Y02zp/JA9a69pok1XavLf
LwfzkrkLwlBhzGTSdTDQUgm+/zAZ2uIQ18pVEXFTW9elpnx8lPA8DDcDcDdBhFOS
SJlRPUdH77kBFPwiUqMvDEJ9JW3Wfs2ereI/dcfMDqSa5QIBs6cmzHB1nxjpleul
s848b7eG+R9NkvlKm3uAuV8l1h3W4HYTnaehpUqXOdVy7fPJil50FBXQZJgQYHTo
RP5OApTl04KkYu64TY9EuYvAH8JZj/L8cg1NQJJO7TfcVrno9p/yvjxVYTeGm+2M
lTBJORg78ZKy1/AhErhV5W6D4jFjHWcTKDvItSQqYMA1OmG0/bRDJJUXwVBBBuYl
8WuVjOYG0izBCUTNV1gf/jbJu4lnsLY7Lf1AxkgaQU01rTmKPdnRgGIeiNQeSI5n
YoQT3D65m5a9/mgHoBkaXWbs3zCwue1L6sFCnnC5ydlA8Ku19b7aZ5uZY+4ONrn6
dvV8qit093oXkPw8aBaEFsgtsAsVO3u2YvzrWPgXPbGWNmBITS4o2zXq40N2OJcW
glUtIHhTSOYvxuTdNxyYnDvEQ/W9DmOFNgcyj7QUd2AQoNig52ExdRHB6BCZO9Rp
5GL+1GR8lGFFWmISdQy1TneIiT8Hm+45fbGn63nvxquFc9h2zjtt9TaBG3ALA2/Z
xanXXpGrTZLnThvt/atTdU+w1xBN3oThCg07X9ll5skrMSCXpztpjlJaQ7CBtDmI
5X2cSWHan8fxFzH0J8ZbHK1DAD967Z0cQuHqakR6a0Bv4zKdIUwYgiviPjUM+d5x
`protect END_PROTECTED
