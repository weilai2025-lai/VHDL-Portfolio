`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdxdOKsfLaxAyC7Sq9ahU4Egl6/ASb1n36ZKEzIRGb7KE+//s4dSgzq2Zp5QdTGv
8oFp0N+MHUrn4BH3y0N6cVQSD19o71HVuTygSqHD5xVpXUEboYxaHTxGEwdASH78
dA2xyGf1RiaWEqsH1avwbKz2Vh/DvBpWQ85JrSZFmt6/gGGNMJwKhXKlw5zaFbb0
SQJaHar1FmzT0bJxn7Ci18TsaVxxIWqSWLcRr9lLm4YR6MywTvYQ8on3ERLwFrtm
okMZKjwEz2GE44yJdHPDqEoibmAyxqjUOGQfq3Arp+i+FWpNDepd6R3+JgGORSU/
cDIoxKGNxS3Ih848ou0Rq6Rz762uOch++0nPe3VjgUkjtKBhUMcwbYNIGhpdjChT
KNxrdrIHyoHe23obxZ9V5TtyMfl2sXKWtFdsb5umPutJLlWbQjwQc7ZZlWiVxKm+
6v3N2DyW3u98oKNtASMQf38qKq4GxADidN0QV8MiCfDcZlLngtfaqkNjIwWsqxgA
IlUOf+4tfaPN1B6uMPq8uxS434LYeSQpMbWuZve/xSgQ2L2YPyBat+HRyjHw510i
mQ7B5uUi2yH2EY0Q6i16HtEHOnXRmiL//MrzL1EAfO+pFB5DDyJC7xsRX0vsliz+
J5vUZpPxJb1cp5Kkh1sgsVI7LLWIBPtFwffLJcrHb6oq4De23OGQAvUqMaPud7Bo
ePqzoOnj4bnpC431mc1EOkhpnZtjDUoX2HlJcDbIXUmsJuHQcVMnUD6u1hQupqeS
LYOpPrCkquo+itLR4XdlnXIIlGu6npQDgDQ+LH6bjQfW35iYM+qtutGpFNiE2fn1
TvDHWYj97JGE5H1vzIPdwHgJwtPEE63Ay7Zz/navwqXpEyGaS4RMPYrmdTJJ74cW
+OKBMXlQ5v3R6V1W8R4c6Aoz2hdnvJKRF49jbD74L3c1NlOIx5PfeGNoajNHMha0
fdSG7siMkaLo3PxK51GZ0OVnYPLm1rB3LilNeQFbCKVWEB7ia/9bSAPrBDzPUdK3
E6lOYJUAQhjMD6jo3j1rTWSJ4XPdj4VLxia3kNEIJ5DgMzWN8RrONBNROYFBnFG4
w/D9fk9VeDNhh31jO5GaHzG5eclxL0fpL0kGwgVeeR0PHnmJx1es/kVvy2bU82xV
NNJTMPdgySFXnON/IGeZMhQ6WfxHLFVGpNCY4EMFx78CwPX6bQk9o0Kv8d5/GSRJ
YM5tzgRTzCVggrvpAZGQl9zU0SjEtQ7rMLNU0I3TAOrdxqnpG/uB/plgcvdO18ZX
JGRTvyxI9qHQxGHkSqfnFja755aJyVInoj8Jp5NuVwp4uKmyHjg1gGrLIqk0u1Ed
BlCN9VlxVcox/RY9Od/q6szeIhJxX/57GJ6TRrtpUAdqIBGe0G0XhwtcQXCuQ+TG
8YhELDDrGzeeYvoAA72hQxiLoVv26oX+x0Ap/BBMO+1gfQPSKBV1l/JjE0RP4AYT
ySaMi4SS4slLCtljhsm8jHBrELeuFSDJC1bw1z+Gay8B+sOeskzVmFlSC3jBSbLr
3PhdtamNrIaYsvhQ/Bq4/EvryB+kh+pr+6q+PyQ3lEd8BjcZoQxbEhKoGuyUu9b/
`protect END_PROTECTED
