`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFASrbn7nYSsau2l8b7G4eznSaKIIPYnL1J5RnenUiLc167SqJykO2QHysl0XnZP
Sb+ik6JqxOhSXGGlpZK74QJc/XLlui9UVd3V1lGVjhctDgo+Gn4PAVwQCf/LNr5s
zaxJeWeeUuCrUDooOTO6gQ4MKaOPJ16o18iznuAiW2uC865imu8SepOzrVyeMHjP
Ad0nRXgpmOhVA45lMKwW1R/5qfj2nllrM3TPnXEH5PXtjIbfH82lotskyumSErWU
MaVDuBTUfoWh1begv+5z6tPaxSCXFZXG+zdBMdT9/bVTCuO9uwotpJLCVJVoI5cV
Wpm+sOP6FwQ8utlfF3mtqlSq9+WWMHGC/USN9p2he7QnJoDzuzfUt8YYekRZRYdD
YZ5FXdEqabZ3qSF6jEVPC6J0dxobz1PCKETlBjfmMib7iir5RCBYaekX//fNRhf2
EocmNT2Cfcd/rnjcte4OICIhqjRE/4ZI1rHHlMNFFHHQ2N5kWzFSo4PLuYXcbnkF
SyyW5FI668udkIYAh4jHzgGBL+AlIDsJ8gw30cLPoYhvVCKoMIj0nhTSokeSuCvz
72BcVaZQbQpO/JQ5QHhIhVvB7h2Vo7yE7E4Gva5imTWzcqZvYSqpJEVsXbc1NQj9
8PGNuZjxy9gtXZgXtzZAi9jsgd+QoX3awaazfCIuHiTz8GiPrcWpWLRTCDHJWM72
Yt7gK8aLJfUoEScgU3AUhyrK8P1Gks6i6MrB9LDrtsWTCZWeopnrbNTfqtIXn/pK
3dYolJFkKTg1ioZpeldaX7VfoOYXD664TEN6hiTnsYi/c8SyMWtjP0dUuiaJ1GGa
BPdN013YdeQZVBBZv+8WyDd9mg42L6+fGcTZySoHpAkwrPY5Q+Y9jVBTEJjVFxCL
2NTHzxSZ14SQcEP7NUcBCdQzU8kQVFlLAuHWinfHq8s9ZZG1E8un2HeNVBqW6rm8
aq4yASVEKKGhYEcgopMpPauUusPGQoHW8/IDyxF7Eg25ci03tAm0Ehe+JDg2Tmyg
VkZLJIwFCVqaPo+BgQoKwMbNWsEdv+scajadCLT9riDOw88wCmAGUPFSBWiAjU7B
GGIjMbv+BKkvceC6oRfwzNDPZUnakTbi+vLEnaTQc3sG5C5qKYxQ51o0x4YIG5iS
X6tXlrB3fc6Pp7XFposHTrZLlvACIfS5C2M+eYrQet4uWKaO22m/TdQtQNB2IJ/U
pozuDRNd/we46JHSTl7UfA0PMEhv1z1I+rWZbeAljXM3bpVKlyPLeklcmlWuftZJ
u3SKQEm/knfLqBMAngiifSp0dB7GKnus833PeVq0Qkd61oTSnRVXq0xWMwere4Ag
43Qrr0Aq+OTfnpFPiM1EeXu0LWIvHWi0y3kZNCvlZinaSbTUWrinmJZXPBZ+Yad2
vx+B5onh50K4aqNB1YHHtokXWqD9aD2543+G/yXbnDO4Q/PKrBKinfUOrjogkxZ1
XiP8L3In3dTLDorMMF5WLy5gpgGjEHXOm48bY7w34Bsb1KQgiREsI8pSMX8IVrKU
m/HsANTkpZLLo/iTIX+DfrT8LA+CO3kJYHlru+1d6/X5VPi3+6qxQKWmFc+rtVbx
e9n4eIDfVcBhxAKZcYgbZD/t8WNpzgwEPvltHGFXAo2lV6SLvQTEw/OZfrnPbKKg
BBchj+si7QqJmdgbqpJjp0M9La1ePblqd3LpbSyTyEbSNbq6DWwiF1NFx8507hOr
seX4QaygiLlJE1Xt06c2YDSt3Nt/dTTBwCjd+S95YBMO1iF8blRMSyLNl+qSTWvF
f3aF5i7aM0C2h7cUYpsENZ9zLuAg+XF/urS6QHcvbp2VKbDmMTUUmGyPcjf69Bhv
brneRBPJLbnkKDH8T0I6/zUk8WyYO9z5zywlY0pgvDKqgAjznbK4dAPKVqzORno5
1Fba++qNQxJCJm+S/2s9pqa9HOW/Hye/Lp7EuEuJSOLdh92CMlOjAwjDr4d7kUy8
Lx3BMsdnU/wiAFVX472MlJHLw/6FgoRHJqaPdmolduOyBWZZvcVl30zVAAPbssN0
OOTzqSAjlOtILGT6Qs+wUZ51/4nwSjZuqOUCzK59lDWZPoSRIU3Yeazfb6dHR8Ec
x00VVn1ATabBMeej4txzWWuaCG3H4kITgyQIKnmpVSdAnxBPB4dOqV2c33Imjof1
K+5EI3qDpRvmeKskn+o2xGsGh5LSftOIgqGf14YWDzqXI/HGn0xdUvF2I46sBhVe
+e83DcmBWAODQjKtjM3ujEctRZktMS7Zr7ldh7xy+9UFV6hF6tpsaDlsIM3ckaMV
/1YVNQr+JTWfe1wvmNbn1D2ivzT5lOD3fP+Mlsfn+DdsAYjUSCuiLpgysaYYCXnp
WxdlYq7BJ9M9JX4iWaeYH+FnjCvTr4RM8KdAyDSVvV+L74u2dj1MQwqDb7ehD/Sq
`protect END_PROTECTED
