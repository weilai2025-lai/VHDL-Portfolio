`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBY0njM68p3nTHCGrNlC71RRbeHUyWVTf4qUX9x/EIwC7B2UcNmpBeVqixD5ammk
wxm4Rbf6INI1XGzB73CsIoCcQCrH4vw2OhYp+1eLgHAU0/fTuhO63kchI4LiW9iD
nroJisgZmjXWbdwNewcyb66YBGtjhE+/mDDu88AAYWOPnNPGJJT9BurJXqCh839T
eIn55nHj3oDtGta0x0fJ4EuUF5CcnqM6EvZZj9CXg/6e+5cTPJvj5qbhhAdUud2s
FsAViJaO74n6J9tP+w9RZCTMgtoJWxulPCaP7TjkYpCu7Pe81qlMpAWg98hVyAQl
urMDwOzBLPdt5ew1cNCZ7PvLBfqFibxZUpCMwzOfR0+6MQzkvm06omu4morJDSPe
RvYuTlT3zhiBmzhmaMx7eGh5AXHLnwRBAx16PJPXJHxhWsgT7Now+sjUFbneRV1G
FTV7nZh5EwQKn6Zv7rkxfA==
`protect END_PROTECTED
