`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLVN1oajnDKN4nX6BKjD6iS8mZ2s6jVnxEh9tNEtIuKNuBRXxbMkViqHC7/2/V9q
l4EdpB5YjEC5cEtqZgAS+0oMjPSbr4dRbtI0kRRFc5EkBokd54d7yKWDdaLrNl8K
7Dw3u4PrENQ8aKiyWNzVflC0a+2nnQ3AZjeT0enJZSbdRYQdiSxxiiF75PJe19f/
le2NBNZa5djJI9+vvmtLRHFEKuuK7ocb0v/JWj9lGp3wE7X4EL8nO4omMSy+ZXF3
616OpRiPBcZLo2CjvXKsPFJmoTrUrOAsOQXA/UtMRryA7bbApYmNb4zczIpXhPJx
aRt/9hDWyN8JdAy2gapGsRef847L46evdrfKXuQ3DQpR14zGnc4Ub4wUWLSKxT/v
spEf+R3G1980FsgIqGoHl/oqbKTHRZPEiZ9hXAgVEcHP9VLe5dkkips1AdOGbn0Q
OrvlpK6fJOC/SQmd9efzmzztMj6HfHj+9fud9mwc4BQwx3Snv/pYsh+iu5A2/fnM
cY7j+J/tpBcX4AMxaMjPrjgmU24ERnabw+qZu71qImrxJryqEADz2/sW+OhlC4aM
U31HJ4Xt6hULsPs4PJAy7Snr9Lbm/QAyKYkGDfBifUmpsMXwgAJ7UgOXUxwZcA18
nT+ITZdO6z+7MRTsPiHq8Ee46ImQEA9oAVhz9M9s5kIzw/SbIKC28EG/UhCgyrmc
8zOS2aPaGSqDOtDjss/szi8XGFgYx+BYQ0TOT36ZBNhS65RGp/7vSFqknMrj+LDa
OGm3/WdmUHMUv88alpPXRtLTPZXsUOEh+0uSGNwfWmNi0//8KRTObsJe6sl4RdtB
zYk5GXJFQiI3vIup9mWKwcVFZ2nXL1a69z0I3rOzr5iPc/K7kvejfeo6EszKTr2/
FguCocVpOaO6q011ldRlh2H2mHiLEuSchsfGprjxhO9VfFHmVmocZ3GoYrpuBNtm
Wb6c7TLYE4Tj71qQVGQsBIacwcasDYRyhn2tfmV9LBafTwZz0kTVZLaLaCcc1Lyz
RIPk39AdoIt6QG9IxIiVHe1dgBnUWQ/g+QJoNiZyD+XUqWHf/oIYRMeSAyW8IhDs
tpGsIeDs1kFtM8xw3VuXggXjGHQDsmyIOtym2ypHRdTZPWhx/z332t/oKzEokfVZ
OGbOqwkG5p4O5k+lrdP0vKsdeR67/xfqnUxz0yriylecNQS7G4Nzq+IrGsLf4Rii
AP0FFqtTlCWi1pr9WybixWLYdLfUlpPvhlwIs0xEfZgQg8zNEeMX1Tw0iT6FVaaZ
RZpB67MU71J0+JwZ1SDVyQ4pajfhsFs/BFbzhMgQGx8G2O9dwhL+DlpUyr19hQqr
XXJi0KhqZBOFD5JlPPyKYoVUK5zo7Z2MgsNOO/WhMSGs0Cc7ZrfJ/Ecj+eUgy4fi
ujGBijpt++DP1DEM23TjG5MFjGtqUwMIUaMD7+kPeKps0qu7G7RAUd+fkFT5nui/
nJVRZDSdSEv2g7GgLaDx3kOWWiGvItt8h6FRoW1uEUc1xd/yWQb5iYduanjohdK9
6vvLW3HM1c9DcQhrAucA3SUZVNzk1YY+jq6yFdxKyCYnll0jUihv5kQBpjb4vKAe
VKLObQIvDerC5VCvOTBqKIGAhQ6M4IHkhEH3EYpdb7f5fYr0u7S4h+ScWqI2Ie9+
m4s1YLJBzfdd06ufwxsHAhGscYiQ6wgtj3OM+MUSOYUxtNjGzv9Sp+bJwZe0OrXQ
r2RGI1c86nLL1JvQU92iMbg0rXB9eS0u4TKDP3XMURgt1fO21bhS2nXcYLhxz3hi
n4JQNjSep4N1T+xuYhSGR+yC4SaFP6SJng23I2Q7d4iwZhc0JqYHehYPkIpoK7mu
CAkGFhgNGNUX8UIF2H8L1ajCrdFuhPeS5NHNN0WQ7RU1yUlK61rQVsCXahojzXJh
2jj2v7zO6Q9htPDvRyx2pjY1YcO0WMZUAPl9KwubAHcEux2kz+V3UYzjUHchCvtA
wSvxo24VrbFTyDa1QJE6ruYmICrIfdwke9ueQkoZNHfYceThE8WVw+yxBh9pp9vt
Dqt8bjfl47UAdz8S+q3qkSZ+otZHW+NvI7iHj8bkJLtNESD1Up+mvUHKrG1AMe8n
SqnJU9jDMn9OUKLRXNyFqGqXY1D/rOoV1l2FIJCCBz8oP61hzq1S66BNKqyokuuf
z6ScxwL3Xb1Dk793NylUqii13fjdX3KHf95u+xwrIC7Q8qmQ3vOFONqnTocGvd6I
LgONb1PnTG9uR9ZH41HQ9Zb1pAfcDERfKQd+ZcQhyWbpPcATcFIbq7oA4G3G6g4t
6e1BEfwsUxj1azMidx8RERVFTb2IF9CBMYbDDWdmDXJX3Y2ZmtN3WSQZPupCkca1
280rpQVvA7yii9rYwZr6snrulkLbMm4Go76INHdDZK2PWvQhOWZEJXhLr0RT0D9F
XzLCBNU5jOdqjsNzjhytTd/bNDgiIVhOgu7bcuH4I5Ex1TmNUv2uq+rJW2mpA+Ez
RgiUlS/moER8aYupWsJizis3/+wVesJWA3J3BOBdVIKyJtKFKbz+ga5/EyzpROaj
E581to+j8kzncpKgkWaRP6PAUjhALXmxLRQp7A0jrd371vH6U7ItnP2SIrwN7GTX
zCBFl7i5DnV94J3XCxNmn6nfdjEsiFk27avlXZCcgd6bforQM6iFn+4s/cTXuqI5
QL0XO6NKCDEy9h9TByx3+tgEa+OqlLJCooq4bEUkAa/nvZAHwtBM4xaGdicwGgy6
NZhobCdCj7os40ujxDt3mFC3dWjX2WD8CPF/yKZ0YTjovxgfK2IpkRe2LoMaFNIq
nvXoyMw8H1vf3/JelGA7jWuFbfEXnN/VI3cfVVbLznmFVIeELCA7UdpMbqqfEOew
AOMx7NQHDURja/uczoXdHWicgRPnfer47UO8SXJ/43KtHE6k2/1Jq+9ApM8z/wiX
LgniWRjm51sVu/teS/k8jPD00UiEv+ruyTHByqynSZTJY3iCgiQdkAmhvGCwjhsK
+H6MFo3r7+z15/bO3Nb1YyVq+wOFMVilsEuxZNL2jUypWUAQtJmKy5rH85YoKusT
C0QHw4IeBHpsRu2nD+OLyCv8uqBKeOQ/ONm2Oz/5+VuuzYYap2iQmZ571t2nJY8V
14c6K7e9RR05ohtnzA8hfx2NEfoBl9cmbeaqQWr4NNEg23caFPhLZiSeQmt0Va4i
5MJufycBTbojysWePs1pGe3MIDldblzYV79r1Rt558bEd0NQGUUdq7aZhFgDni70
6G7DKVWY9gRUjBktBtItstg3mEKTRe5Bks7KuhXOWQQbBPSQk8kYjpaKSWvsqybW
zX3cdkmd1/YDYmPEdG5vYtY8mCzdei5RrUk4ASrAGRK+9fJC48L6LlXFjrPaJQOm
paYSxZ8soROLIi2c5RJM1mJ35pXtZ/suDXayqo4eVt3gooU8pFOG1d70zY+f8RcB
jKHVBT1H6GpdVCCnG8XwUEj+C6g4zN4tN++Ew8k7KjMieYn0jhV472MRQRYC3cyV
kAXuiR1CzR0ovcsovho3mXL/vCTuRh7W9v8dSPoJbb9MqQnvzPmB+9AaXCp886F/
NY4RmgGe5GyxVK8Z086+rMMBnmqZsfkpuMx1Sx+Ap/Ji3dSJuoHdqe7m8sOQiar+
9K9hWRZeaZCbl8uAwdEJ7yK5KXSAbJ8XmY2EDp/9499P/SlRd9KC4iG+O96i8SNC
tLKOqesJioQqtWWZa1wc4WTvTbuY+Q7l296h5Xz38iv782HmNcZc60XoDueryrVl
zEOLEN0sCevzJhXFnUQINev0uxTVp/DmK5V1K4F6Fk+T72vCfCnr3873O2LLPx1B
VZvevjkGFZ8B69va5QmWGTKmEbGHjoRIHCiBB+lQIHDRti8k7zczXn7geLkxpeyJ
ekQdugRPVIRXyObRXzLReZdYyKbqYsdEQNdz5TxkB8cvO4GEl3oeUodc80JwZaWu
P6HW2vl3YKIeMIRgiJoSR8AXvsMlol8epHhjrSSJ/hUKeMSzS50p1cG/uJdyP5hn
ZWartOxZdMwBt2HvvDIZaB3iS7ZHueA4WIExnFXb69+gaOtOwT9W+qM5WX8z4e0U
smal+x3DWtASr3OGsM5I+qg3VAbfXr8GsT3bHSFzMfLMlt7zdfkHN3DFxKYuCNei
9je/2QHhnWmxHKKWWgfn1Vh2BidLttgLb40b4hYk9LJqu++jDz6Xt3+26SJCmp6o
jAbhShGrmj1m5TA7dpcY3DEGPaiYiUOfhfcBT875G86EKSE6co4ZcIKkvGV6tz58
bSxCyab4Y/bEr9zq66V1bYAKopWk2TAc/YF/RI8C/BqJphbRUJF+LI4S87G+/XHL
BS5dyOWFVaZ2NAbjz/r7/eBtgBdOOCgRBbBjgk+9etXakKph1I4irpEC2nCJXoNe
tLGfEUgu7zYs6Yd7PjtgvtxMhefNeWl6YBwLECojrVzvh8IayB4bLSl199iafBYR
DsekVebULF2Zxv07GRHRMgonxMokYg20cVCYcMCleLhJ5aYqxwQMUflH+b+BFMXl
mG1ub5SShP8Z+fzrZWXsPwLTuSUNFiB6jbALJv2ecRTyNcyHCC7gsg4MShJkT87z
bo8rDXfXRsT2UW3+g6B0zb4yags7fQ4OAXfA/Xr6wwJXd0qO5gKnusAIogRXp80B
/3urP1tlgo0FLzuS9xPSZY7bLfi8E+TUo53O2H0zMMdgRB0S3OardAL62YCqAHWP
24z/gMsU6dhZwhBE3nH77o3Hpbu/PL1b72pnrstRwnJ4k118A+rwcrlX058cierf
HolkuNUPChTgAVeLT9sZPT34uCpGTZFg5ACOLYgru/6QiSbyF18aQ4IczTbo0knB
Kohl1SwwxAkpUVu/qx82wWVCphQeEI48YFpKwJsoMQcsGgoLltWENZJ+YdHF4jkP
8ablmjJAkw7xXJdeNDNm0nS1yV7YSvAn57cCUAkPVhs7RVZPbGrwR+iTLsb1k7t2
r3eL0Py/kcqJprK9NRE79gd6yRKxPdRushKwqW+AuOkUlQgtyt6oUX78cL07xhl1
anEhfiv+FnaSos127saMlKJMTLK7pNN/HFRR0aHwjxOmQL9UxtchYUw1pfKT5qyn
HTg9lBTXjiHNgFUlL32YDLDAE8XQP51fGBPwUPSQmART2onZBHc+8m9EtGj3HMxR
dgkKD2rokERgknJUeIJAIvXFuJ3pevp2kx5FqHd1pDoIMPqkqOBmXEiQv92uubsf
ZmIhRIeQsc8Mphf3jFEyRxlTV1gwd7enK78q5wqV1lWKodcT9E/8SR8oPMGEwqTE
jwJJqCFTc1Hs2V3yKgU2ZYVqpK8TS5Ps2c2xYItjFwMX45cqM/HCAIU1qxBZxHTP
LE1lKNNw43bPP4Th8JMrToNVsffk0gykpoA54xMdrTo5t/ZsAfKwx2jpO8VDFLVZ
MowkBo8yTcDs5HOYLJYCFU2A6SHE0e2vWQDIgHzflTgL/+ZQ/6/eurXByEHRGYZg
HcD40GGN/5pnM3QpRtDlfJuN2cA8TpWAZmmLQGoeA507O+5+362PXWUBd2lpQA0r
L+/bXdJ6tvvSnEBFzv69i28nqN7UfWHGZEGUXApFDveIipH4vvn82XdxrEhRJCxd
393M/Pv/M69E/c6D8hWXxuEMY81+L/yiAD+BpbNKwnO6PHcBqwruEYkbz7uAr4dk
1db9bb+FvY3XxnVeOoIokNoQd5cT3E2G/feqzDI4cyjLFUzTMrsuZyfRsMYEhGVK
VimJ6dwAaQl6jpZbSy1vGetdFpo6nM5xw9o4KIOc0Cn7VcydA//qJnmjiimJc5WT
4OcaKCC/B+O6VXtL9oTKoz//6i95Lzsdp8satB4JVNreJZA2zudcQrw45l0OmueB
DgFiRhPE6nmMMbEeyWetU91IjhejfG+2runy9SjjAkgpqTYlrQoY5Qtqmbv9NXWQ
IBqNL8i5CJ+MgaBPEeGwYVXWS3cxnXHzQLleRFTG8JCx0Ho0k4n8SK+1OT9KcLLN
92rkf8bjzgpur/xtvOhoR45s2T+dZ9Nu3Gpcan42h3u6q/lDEPh2LP2R0BCQF+zl
uf9aAXrswFYkx1QKjEd6iTDg9FinieipoBhICM4O4iWOcWaa47JCHeIMN49V2EiK
+BTq9RMuoGdV2LZFm+yYyyJhWfgo8PL8nz5oRY54QqEJlSkuT61drKSpxAKhNby9
tVyhSpbXXNW4oDCMqE8fXSOlEmUuZggB2xYlQBLMKaaALBnuSiU/NeVJIb9q6dMX
ZMyFMq0NBaW/75hNPHlZg/ogutn0+nVh40VIePJea8AeqsQxYtZwfA80tNXGmGuu
11ozme/BiPFTf0/TCE0LNMEKjKR76uyrzZECuWCHa0abYAqlStzSRkoat2w5RVZG
+bPgcrM/VuDPE42zvK9nfNNwEPond6eym0aKlZJBBLFpcSCtoofJbqOZLy198xj5
a6rC1zjiHk6ForYPBRJWHW8t6gKVbAvpbG53c/SRFG4pWV0WQ6tHnEtIsaDhdgmK
nsQRJsGYR+RTzum1yMgAKspp/FesOvEvIuNLAoHPxxjfdSpyjPK0IlSsNFa2xqgO
CGNV0VY5844i0IYTFYnOZvpHjxV8wS1WhGcWll0nzhjqdXkqimDMtyBkIBc5QdcV
9ncqH8sFOWYKQ6yyXtigqZ9Nrf8Hj7eKFacCdpcmEgR/uBO/NzfFeP3ZafgE+EXi
mM6WYUt4xC5zWRz2sXDEEeLbrhDu8pDQ/JkilCBLqDcpGrsexmXJ1dANUAZCKr9c
s2O4pv59vNFoGWM2zuCYypVpjHAK4TOcvhfPa83BkSJSgsWQRu26Hnh4uRxiJE5h
Gb4czioo5FckUWn4sfwTe9yZIzo66X1kPlkcZ+L4UTDY86J6fgVjQTkhynOKPpRx
vBl2cnOXXMmMj+tfzpsyPnEM2iE45yCQmblRFfusz1FMHss/QV+DUS0vBZ6uhg8Q
JuWhTCQ0Wt66JgvSMTukUMKabZQ3BLUuYZg7Ih/drgrpVnkH78cprBaO+AmNZhxI
qw/tikwNX2OaIzPFHFFQij6ngPoAMj5K8d9Uo62UcudO/MK+GjfYXIqGqvJ/OZny
NneYPIdvHrP0hJoqtBjObbGRIEz4SOfau5Jb7FdCRlMJrWLitSh2aepmAEuSBbgr
/Q3MWyNDt3FoHuiczq/EwHAgMmt+HMZWQWTvtmKk14MpVjZHmdZl2LomUsXJdLcC
dr67puzZoIzZmgEE/4K4TPIgpKjzRwm9a6TpRj9Hm0ETJx1yUnN9HyFIi7lfpPKn
2LLDVg3ylf4+PM6bsk17EIA3C/BIeujLJk+MWB2C5xAG0AYbHMiIqmF36/I/vPWt
DLAApsvxcmsiXQZQSqp+qLeq/ttddqq1/hvyNTYIrT0b9TQpGYocRpUFm83A3G+h
dFxceXf/Jyya/bbqD9fEHAKkIbJydm7xzzIam8boVXTtguuD3yeZyrtLjiYG+dLu
ywM9180XSfKr/Z7YjkXSvhZmkLSDQBuvzqNFqVUMPnHGGGfDkIG9FSR8dmbnM53/
KYX9TTcjMX38WgP3OANJ5Na6/Y0lMHmlaGcEhUbXrWoydjT3w4PiEoAoZUTb5ePX
uhrSXj/jm62YxSyoMTai2Ln5ERr4Ij6+fqfnLz2Z6bcoQRr0UeHM/BOUux88D7lS
hqVF2HaAn41m22a3Wu+XhXvVZzf/ZRppYFnVkQG3Xh6ZH3B5tipO5R8ybjYHxVSp
T6YRR2PhN+g663zoO0y7DRwKYQt4M1g6QAWfUJJ/Jz4Ocx6NeZipWS0nx9ZX2ile
wTjN9exjMiryxASjjqHzi4fXN2GWCjIKh8USIVb0fI2FGrZoZkhbZqHq5WlEtfkS
+ADdL/HoYSjJzZndrShW6J87gGMDiw367SB9zsRFTkwAzqLW8qqkZjXwGkV0riDH
72VmrmEc6nYoZWkPz+9BPqFkitHf2umwFQQOxXlBZs2ZkAvLK9FylYEbv79iss1x
avHUjQMzidWOIlzRQqGqF35XrrzW/hafH6rkyIy4aKeX4xvuUFUsUbrUUIXXH+ZO
dDNb7bdg0/ae7ItMeqDmd6zSv4NUWs1cagWDfkGPJlcKA63R+R8DAXG0dgotI5Fx
o+Qbqo1/AhkpwtbMXQVz1nrzKZcRHrdemwukPGIyhuIB3i+eU3jgUFHNN+UQoXh0
wCrSMVnAlcOWMvi78XYUQIDBV0XHRmEMrH4/pNTzWKFbeQdCpf+WuZygDkr/PyEG
kBQVJqAaKyaVv/Wx37T3tQAeqI6G/h8i4ItM8Ef9+OGyPfixsCQr5cTBI51EUssC
pYJfTe6q8+i/eIkdydHWtJf0ni/gfkuc78eT4VLL9nVNapEt7FSIKP8FjZGjJLwj
H3YktYprCL2ZiQ63rpCXZJvEj2nVJmLOyhX/nQaQejPvj1FA0c2iNCH0yVoMuhnQ
Gc4J7jSbI+Agua987zv0sWt/jv6F6dDRTtsylYKGo3F4qZnKBcOUCOa/fOFDBQMP
o9EhxEq42oJfaU2AhX7jG7LHxFfiJBQePIy7q0yOLpxDUGK2q7adcQEkooiMPutH
4CnkhsjK46F34NlvNpUrz0pXa8yda0a3k4Cma4jMaljwh8bK6k1eGnbJT3DLSkoQ
MppLfj70jfm2OCujH643Pc4DJh6sI3mnTSy5sx0Msz7quZFM5mQml7dB2pbUrMtI
pBC2jyFY0XQAsA88iWJ/bUSCst0IXe9xiN6cg4RL+fLaSHPq1siwWI8f17UMZc9h
wjy6g546wohVNc9XYFoUcYCunTsM9mferUYUe6OX7Un+6kStP/eE/0aN2kUjm8V7
Tqnsa2hm3aZHJW0LEghYLsHTcAuGpEvpe045wbZWNl+XBIxvX2qqZECeDaDfx4jj
qtlCAuI8IZ/Nwh8skSs8nA9CNzjLC24LLH7bnlHWEoQNYCUGB7BwPA3BbczUKPCY
t9PtBSxVxDouEOrxNgZoann5IVppF22L0VdGvvRLi0as82fOPyNiPsg1IzA/jgCL
4rpB+EJ1EXznbqznT4ZGl5Udca/48WFn5n60r2Z/SzdJhLc5b58WKhw47srOQBVc
jgEjHgBK/d7Pxk663uPdNtcSMEPTv8HHup3Vm97rF/GMDADfl7Ral0Sbg5bsDBC0
XdFPi5oH0Q2YBSz8UAj2sTrx68gLstcOeFtF853/GHxZomVVFYEcRZKPTo7Cf++u
46FTC4t9jG020LRXyZTVvr8I6JrBugy0K1mv3tj1Oy0893gfdn9/HuNOgmXXJoH1
P+aLoLQrAj037jyvGpYcsxqUXcXFdotNPBJ05a5x/1Ptj/x5VfKfHNdPt9qifFet
TLq6V4XT1hT5zk77ab1LpjWzuPmQkMo5tsRdkh/IhROUNgXn4ziBSwZpBMuDYo3X
uaC2+QASKAdajEdNo3Re16yxp0RbzMPUW6C9ZN9mzdtDWgZZhxOyalWo/SiZSHdk
oS7GoExa+YAGaP2/iEvnbOMMFOhcrB6keWE9WgjbumKEWtjgkSPIKhpA3AglWqJ2
dpvkNMufHTWYVyHZ3woI8OoRjxs2oU1fpzzYAPDINvzmVTqJBY2v1xjOsTx5CGwe
vKF8/EBipM/+aP2Y8K/yIzJtHqBbI7t9iq7OKEUZV7dULIlXxHav9PEIJwBCZSWa
LhA9x8IiGwuqGhNd6863piuhAK1U+MgR/v6Ghr1zQ/FgfitxEWXU1JbwvVmQDPRo
5qui00gqpTudxU0CYCGHA/ULiK40JP/CAQbOQQcu/mQvhcoO7FZEamgrCHT+eCb1
vJPpVfQ4XPqk3bXhC5wnKzsu4ECousVRL+LIZVdWWmwXMcg386qAWh1He4u67lmU
Bi+OzZzTV/qQyHXaQG7L9Wn/pxR6rcN4o2O/cLbRlrpwXDMTJ9HRYpzj+ARJTkxO
F6QEd6PPS9plQLT7mc2TEkcRpOFJrC1nOA17fkSU6Gjwg9oA33anVs+9PSeZZhBP
IO18aZl6E74Pys8stTN/wMk6i4qeHSJ5PXvB0hWYenKb3aGeuDr41Xy6onbtviQe
xe9HXfEonHw8ze4HFRVRAAP6/fTQhVQ1SNZyjDV9101PpNviF0maza4F5iQRjuiK
xXPVoiupbxh1VIwbz92p7YYDiyhhyudfDfpcEWzyBN0I+C5eTgn3xncHnSC+f4gG
xT3NU1jpnAJCfty5KjYHuwUV84p9Drh+Ja5V94QCc0HOOMe7YxIfJYIOF/YHxLkf
OvcD5H5nxELT7wUPT8kWInItcnGyWfey/jskbqEqeu0T28jX2K2BS9kDb7e7Wr/R
B5R7lrvLNGvwdAiRmhhOX1TW2YWC63U4Oqyrb5D8YiGyKkmtnNQ99HvCONetTI9w
LuWknOigW2OjYkHztVmK4aJ40tEPoo0FkluX+ZjahQY6Fq/XX0DSsX6tXZSgDQpd
+SNW8xROxw7xYDyhkHK1OGRG8a2V/e6aBPuAFysXuQSkQx2atLwCowxhFnNVg+nP
xSsEnc+b+fmlwJQ6NJDjkWDbt6xRQlAvAm18QgF1yaBWKwgFKNd3S3oznXs9+hcx
yWfd1qjeWJl9ct9jrvxCZ/ImnBFtS2OM85rLcut8is5RYZ0pbgWMh+NJywH0gOLT
euJ7qStbel6oVuCu2OxdxpcwJvrYhzt0gtmQwzOi4xQSc2EQtPHr92WFr8X6StrE
vgjmi6LrpwQcP5JRSxJJHJdMro/ZE1mVaSLCjp+rHS/CRg44w52iDC1xNTzjSrry
XyZ6F/FlUdxYgagncH25iBedeD7P79Ba3SOdYng1HQDUru1DyrPqnBwweFltoN52
t3RC+d6jBb+u4WO4vL8PEXyhNp6EwNeVqRoYQkmDFMQXOTNqMUHOC6QiRVutn1EL
b9lIDHEnIRBBWWH2CM96J5JVUtmxTwjfPfW7Dvd1Kfc=
`protect END_PROTECTED
