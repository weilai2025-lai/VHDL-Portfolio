`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/XNULlj6dT82RkhKpYpJAc4AzBziJpSlQXD/U/rQ009NwwK3GArXVmjKX708AVs
EKi/PatO36HqdVfeIm8xd2xzbqPOhu2y/sHdeg9CkYopeQD5DXMRIJzFYxGDb/Ix
CfA4y5+8bzpYDngtEH0WLzjnpi/1SLaR0vkZzf9Yy1H29z309A64QB/3T2EIt1vs
CzLhXmsNNG6lF5GL08flmUkQs6eU+ZJNQ5RvosD12MZzR0+Q/+xJT+UiyMptqQk+
hOJoKPM0Rmr6P5sEowwIeX5QLQyrgu1mSAaLJen9Iy8VDy0HnIAG99G8vxYqVxN8
IA7qWRPweH0tpTa5JLMHNaFVZ3sUJLJNOMdhi6Sz8vlkxd+VXb26ofCRLxtQMjsc
IooSWT1/NR+7MEMkDxS/mLwxfTq0ziTHAQtAUCzI8zfH900L4qh7OiWe4nd9fI7t
z3WsuzgT3kTCfHvr+gvuGgzWykIUi5gElXJY9A8S5nOi0fze6YSdxFIl7hxYyK3/
dr5eKF8pK2VB0mlYmLeVlbfaoq0G9CShP04kkGe6Y+Ye7lpYp0JJS67dvz1xMBeO
O7xslT0coTDRFQPO7r48NI8VZXJ3ewdMZUK9w3yCaHVRQosHz62XKeC5lWD7HNET
lXZuQ4D+bbD+cwlKcAogQeJKYID8HABzoJUv9s5j4BsgT4xTTaFgIt66stSwmZiG
8J6Pw+n20X1EHdevZ5u0nB56CeKoNRtsEwqzwu0WStxnYapa0uE0B7Ce5Ca9Cr8L
v2Txl7G5dso1n4F6GgfHdmt2Qe/Ve68xB9mPTNJ6ako1vGdRUZPo+jJD3UHHryw0
SqyOI2rXgvRhiqCQBZsqGLy4g5oHr+AZ6iyb4GKpb8Xed3DvRZGt2RO9vejGELhH
aR4FL3fw4Tle3GwatTXllPKFDD6YX65dy7W9QYQJJP0idsl/H4bgND3cm03jLgRp
+urGPw3CuRyV/23aN7aC65q9iMABoy2xZL1XzTmTHTSKQmvXYFKYIiGmBFm88BPJ
V8V4vSTy3MA4D9i1HMoO6+RQ2ZNNG7fg0KTaiCd1Zm0Fmw3C7WLOCWpKpmWQsEK7
hQEoj/iJf0SnU4l2gmRL9SmrzbVYuFM/GO+dENVYqGZjTrAEwET0kh0p29jagP8a
hykI1nWmkOxqRoA44MDCzpGmK/cIXuq3OpspcXUEZmNdS/1bxBJ+HraY1zfdoB9d
aVY3g4v7VeGZ3qIQPC32t7H1nE6GyLn/zPUD6cTYb56TlDQF/rNycZDAEip5Ws+Z
27vIkTdCTJFvPlSnhteqVQjxlIkKZCyD4XrYJC5+laY0I5FYoVpysxqtJykJy/EQ
AiALjWwx8+dYUiyAOHBrlO0lrjhpXUwmNw4i87K34XCQoB5vpMoO2KkXgJWu/JOF
/noEERFopSOIJe2yIDlNuTV4Y+OaJnQlW/2jlwMHbwLoygkksPxSBkZ2zx0KOrnj
yYVZA9dbAaR92aQHAp9Dcv5y5E9h9WbK1ndKSO5pSsqiT7OzconcTTv7Oto6PGxt
c7DLtJ1sKuBv+nurOvQGdBQnn2cuvsOMPLcjrLZRJ7Ud5R3xg1kkGKa0PidgQ+JJ
iWmXXdn+kpNnq92JI5ECAIUN5VGIQdtW/kzsg+DWp1dPmAUtVZgKznwbakUBjHHW
t5X45cKO7PJBv4I09BDP8CUhQh+ugp5iKEvKNvanLkahyQq9uXcA2P5kusYATaGw
CiNYNEu8ZEoidv8IBx9UBzHNqyLTFeRqDYiSy1mU5DPbXubRUD0Fw/h1T1LEQYEG
OslrvL8zoo32RcaOe+VL/bxmphgzLaV/pgJ/TzAqir+o+XJ6IrbJC0YI82J/TUfC
0LCSnMJ9+dRZflxxWWEgSZ1W7C5iV88L9YBgYjeyfcQ1MeAYCrlzDto2gE7Bxzk8
r+ScMJ+HDT9gGMgqrXBxViQNCvEHibItnv7mznvbyzTVS9sdY7Kbl67E24QyH84M
6n7+Doj5JtAcFopeSeqe273BMCe+mKj+edRCr0zJeGwM6+RCF/yK3PwjnBdJWV0w
6K6EZPdm5/mK8MFo41re6HsUnSHb8r4bXiPd9BrZcLxKCzjtWNBeiJf5oMtzIrjO
CRg2YMj9/t7M4VoIyXSF28gQ2aNvLrlkjFf5kkLWaQ2E+Iqh22TSj3EvlPZyor5C
qKGBtk/kSBKcp5dgycdlx6o/+I2owrdHKcIVRUYrUCo4a5bvDQXAz4GKph9sAn1e
PvguqtWojV+GKSAjOSmT4VtFJQ1AGZCcjyBGnq4CRvllcoqisKIRtgnkA4THE14J
YoKjhGY9wQrSF1uFONpBbGN+FD0wBU1LN5qHcE4fQ3TslTgPS9DS0ByurNaq0OeP
K5sWmzPUPgu2VCZjLkep9T2q2cWeS9zpXSmjlOPN/U5G63l5EmZG2PDIR4vi2QHz
W3o+mFJ5PGtVW+Y6atBSKFaV78E4BS2oBhKOkDcfVmhpMlx5/MrkBuRBkOxtw/Pi
kj1o9P/y4D3f9gxSvx2Ap7qQX6Sqqo7VMhnueh+EyvrHK5+HopY8dg25KFgBvyLo
tKkKujj77qsbjDvW2h3bjARwlhOrt3Qms8wHy5zIhfEthildik26ibDfSypn+CVp
F/eu9huK2IBHxyew69lboU7zIf2aMTwj3To7Ybbeot7dqABqcqMcERj+iB0kGjZo
PM6CQitU9Ax/rZQ9f38xLTg4c5k6KMN92vagfqY8N2R7ZNMcDDNJ4PV6h3vdZizV
tsHtG+JmLHnuIuY8zrsTBdYK9vJ4pYRQgZ0Rr2M7Vk7//k4l5QwAIANkIlafMq8N
TwdLvCTE5nYQXEb8R+0X/lnOlUH76ifQVmsqLUWUkp+NzqvRk5qfvTNBPEhzyC4R
n84fEUHiylnjb0JJcoIPwblEruQ4ipd4sJ1u0WDBABmfFELcI2rfUe7y5uQL0qVZ
2tpOm2iWVsje6iPSYHtFjgti/88dPMla17P9vdREFF60ZgxEhKOGclgzWiC7ihp2
HwqPnnGMUvaxeHBZ4/tYWL8y1UCEVIgtB4FrpIdpbQLWgFffQSuLiBCvbsIUpC8O
WFu2+aLWhQFxx7EhmHbG0NgcuUL4XLK6XXA8D1p5o3igNqwqA/gPvPbgj16V57+m
hdZLfVJwVO6mTA/T7T/2EAEbVV/DD+wRdGbIe4HPWIWsFo8gd/ch44LczCCCmsP+
Y/aFVU+TzqLzoQrNdtgl8ubAPyc3NSJM5hM8GvW/XlYN4bTpERxyDmH7y2ZfAE4k
TlA8c7+1P90AHc7ES0ZXP/zRQEXOBcAdkikpkvAZW+yCeQGMX+qcOUDxTodzEfT+
HUgcuMYXvEhNz50F/k/34QdEWaH1f1OQSOZko72KLfVik7C/W6hec8Njw3q32ZHV
1HcqhHpSBPSzFNI00c2ajnuaOuJrDfz7tAG8IuzGY+AEWJ8z17wcEUOt3g+tJnUo
jLsAF1DfQmz//pAQ2B+4U5h5a1S4kUPpMTbRNW87cupmQIoXcZHMpHUuK3AmueVA
vDEMgLQqXQ7m1AqAybW4yCZjydnJNkR1D71RKAxJgwmA5AD6Uvu4ObgKSaqyr09X
fuTsoyV8RKPRBfxTm80/zzRlqG3vdcik8EoF3rsJfoIiyloF2Kaejg/Gb7Rr+qiw
VXye30rxLYiG/F8IFCtC8RNFWoPSVzQ8udUCAmGDfui0kDtPDHh+TzxecF43pK83
u94WoxksALyLbSnOFXmjWdfBnJrCkTM0VVvDT+d62wzXvG/e7WEtX48DtRspW5Ug
Y5mnTqboM9QO5l3He/YE//W8ugMFvJGm/T1hb8cwjh3fkvPh32y6b1KZJvAiZ+7I
ZfB7zVDHl50aCUdySTWGjEqm9gZ6T+QVO7FrPhtghDnNc/3k9r2WV1iIFUzGoM6w
+ZCubFKsM+aZdsq1eTUA4lg8jcaU4zOMbfqCSu/J8uCntobBCdo3SAT7ZX6A+bH5
v2owBLXHT7BUfq0plnjAgXVXM1MOljDU0z3dron3992gsGH6T6UcvPlz6qjZPk5H
RE5oIZm0ii6mmszATQ3a6qw+NBrJqG9xxvTuUQmvEmwkQzoCtEbM2anCxZMI3NxM
TC1x4eD8/K9OJTuiY8GURzLbQTKTMsZqEtJ4W5v/WOb4FUYCZ7sdDYLD6b9+ywse
dD9Z7wO4+kFLbXEdLSFxcYYmvJu/hz9P5/ZRvqNMdH6px574inkIzCPfDEKUcDTW
XREgPaS7TCIUd97T/tNXZZV9VNbogk9Z2J/aUgqKWAv/RuO9xGGdtFb1ntKHWwZi
0LxgTwwmrJn7jAsrBbY0uVwXMpK1N7EE2Z1HfwiBfmK7dq3zT086YwOkuOYOG4C/
iBNWI5jcVS4G52HzuA7UvSAXIgbZGoc1JFjhZco1Z4Cp1sLWTROMqlZWuir37+YB
GN+9OZSE7wmKcOlfGjxOqcNIUSidykhqIvg0rUP2diRpVx9AtvqhOTp0fI4KPlmv
h6W7seFLOsA4Q8Hy9EX8UTia/QkL+NXxgEwD/0uCZkhBMb/rkUTisTMyoAZAm1QZ
DB05cp2F+ESE8x7y4W2H8cS+aPfvlQnO32BpMR7aMIQnu1zgRAj/GFalSC2w9Dcw
FRaOlHd+0avFTybNCPmOwY/DVq4NKyTuZe6OQpLyCzu3qM0lcEB4y/MqhZ5E71Vn
7AdIBDDbO3AmidoofVTRoSC6WZIMmOwM/NpASvZ35ShZPVQdv5gfyZPxdUz3og/K
X0QTXdOv+bYGfi1ErjNlQbO0ooscmzQrwh7ykCqbAz3EhpPD5+ZwVrvwE3SbLpTg
rHABniJ/Cyj2BKRRFy+jf5kjcXxbYBm5iFK5N52+VTlvTGuSdEmQ2l4xuw8p0CCz
1lKORlc2X9U9rzqnfy/A+wubZQtOhIrln5DuK2yVJhCIdUQJE5eKl5NdsIuRPzmL
vnisRTeknVFbTn/d8kpcTnqmrqNggJ8lzH93nM1RdZydZ05T5N4VivN6BVFtrI8V
XiAFF3Rxoa9tr8eWob3cFC1StTNAr9dIJa3WjVZWlllcqwTpCgnrM6O9mqw13xke
bKn1kKfhD6Lw9t0pYbd6u1oXhRwiZkDBFAK6FWXNhJQei7atVLt1utkuNEmmzYc4
/32FVnAOos8pqkAncT0X+XBtqy92oWEzADJU+OOWwbKrJjNoj/Vx6FO+zy3sWiD6
9yo7/f46sSd2GisUKfMmxs7xeCeF4qy4Q7Gn9t3+U4jYf9qVokIBdsZs1xX2n6sc
IWM7g9L7v9p+3NpHf3GMinY1Vk6dxPA0BH7aQ7t39o7MHJzTDRuHGXfJoWPln+Gm
jljyARylYoGbYDVsOrlcpwzbbo2agzOPvY+TatkkFL4ZD/CUAV0BNRZJ7aC4sF1j
ZPrDl9X6MoclulL9prpFc7BvArNYMS0i6JP3MAfcW31pwndpAX8yltaPHdxTQQDA
OeOsEjSoacbq35HTjg6Hp+CXHe2cHHO5QlG/jUSVByACBIKSH+1KeHyeMxr/nQSJ
kXRaOicflSsGNDDPsFCq7ceS3bUKI0d8tFK6vO8zaSXb+aapEU9L+j9IU1msvWwp
sKBu7XtBlCqzvQ8m7sxXJ9AjS0TXONujyqnP+xn2onyWYx8GlHzVmXnzwW3Cw+nk
Y637AyMkOMm7GZQJ6zzZP2i7Z67XOWaTgmdAVybclWFfcGhnEJrsouxmCpmkVT3W
Nh1aDW79awrRXmMsoAvJHiBe2p0vgqO8bO/Y6Y6U6gQIbibYscgEE77w9E9zNu+4
mmVG1otjGGjpPihxGhAGi9+uNklQa+zfoP7tZykRS+BKN945Laur11SWpV9bKBBx
JImYIdb793PxtMJO4K7WF4GoqB+tGosl9yg6uUn7h6XvfMn3iQZsjVEjZZBD4tEQ
8p8s6W5N4QgQcO0u3DQzE5yeVGWrPeU5lhHq5UlBRD6M32sb6a2WAebU02K5+yFT
3eK6VHfPNgdWTXTUub/V/+r/jJ+BqnQMmfeVyu+KRhoJGNEYq8CTQhbeKQMQvnct
u2MF9tGkjKGbqMqan7Fm5Hb/uYy98h6psDHxzJM0swSndGZ6DQhcQWxYzovTydYI
3ljsB4B+KZiGWnOEiC21d9hr1/5ZC5XtvCMAIKCkivq2R6cJGpRMn5g5HpF2PNbt
MRogl0NnSBhboiyWT+8UlyiZSeDxM5HBWJpMBJJj7SsrUNjfg0LNHwgrmHkSibJW
8lvWPQBuA7vyJisfW3qB9x5CaDJv6LEejLK/ujFdSBJywDugeL4qn1fpYvdlI3/b
Al6r/UbdQZdb/6O76NRPKLJ40sVWhbC9jTKbZ+E3BU8MYZhrsNif0JeW7eOXFguo
82mxwUBVGQjcHwl9FbVuPp2I3gh4KfUlzS9fZh+ubNU+ANss8ROCi3lOypTgth2b
G8Lof7B4Y+fEhXzFhQKvc2ztGLp7OB5mFwjn6pw8YfpAv6zLwawA2nUcTx+WCJo8
YU7rjKd45ZvaBMEa92gd10MTCoilX9+vWAKKuqkucTfRzwtYk83ZuAvWd1XgxE0H
am1Hyb+fafGXlrSQdL+1uM1im8IrDOzIpwi+CAkF9l1UeN5nrJOMtY22BSCMgjKP
9U/+KL/JCoXMgR7vGstcAPj/wigKuFHSqio5ylI8xgf7tjTSSuBHYNQTqDnAW8KN
93NGJHO8yYE47aZVL2+WkPMqpOERgUpJBKA2hN1LsHpJguulmG6gbXPrc5OtqBh0
L0clq4M8jZzMm1ElEwe867qeDIv1zPWSNQ7Nvt6FgRpK11AfiKu18sK8K+IQhVcc
LOHCElov/zYYp9A7/1+S2upgune3jFiHU/0HyYM75mgrUp2WXzK2R+IXiuqIMstt
3LihNSWj4Xx1CzjFMiu5xohnJi7fzpJLUWV5VMswgmlM+vH9jYM0gGaPLSXOk6po
ssq1rISMaZXw7Kk/+vXnxVg6GLY/CVkQnRSYRLu2CWptqj8fFe8qVebPmyQm2fLU
rK4UwIfH1m/CyAfQtr5VoJSxakkTYSHNJMCulBBgYB4IwbEpZ/Lju5Kr0rF7QjeI
GbLCvQOEc1U82KEd0bfS2gu3ET+aP+6rHyhQCfALsRXeUTQcmod+Qi/+WdRDjEHH
BrkiVcZeiYPp1wjs/w6jsDJ48IJ724T1nnJDR6KCC3hJpPnjhw5Wk0mdDq4LGXcS
XMLJkoTmnIges1Co4somMzsHQ8/Oa4OT/LaZ49WR2wTyO8eHn9KbGWl9wIZP/pck
hDnnpROggiDZbDjUFyCSl9rc1EMjczPxnEn83dGAfj8=
`protect END_PROTECTED
