`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XsjzoO4lQ7LyPFejZRexwbf8udTE7zrn0KhaiuyRGkaIYRAPTxeZMmRMABYMzHsK
FKNMI575zE7ytJjzvZoaqITCAQmj7HYSsBzI4L8Yugv7qd8D0peSz3HxOfCF4lCW
Yn73JXWTszlJ1zUi8j+ADRjBimYBWfKPPBq1+JECvaNwxMwveXHOR5JV/5ek6Sut
EUahyGIG936ljpsWWWh1WU2hRNIf6YB2H/gXcbMAMfKRisSwYqFwfk3l7ici4UTQ
IA52cN6l1WumsT00wBehak2IT17uYK9kjSISu294D8BojU5oIqgFu7Ux5hwdybz6
WlaAwjw18vDtquIRaJb4E8/93Ptlm+lQr2eBx8TGfI3qEYmTj2TwIIwuC+vRuOG5
95xqbqzbuAja6jBOYlK3HxOfTgMMb9eQwaFoYsdUNmuGecczE/qs8/iNITcD4I0p
nRQOXr0HSGNH/RVzS0MFWY2Cpi1Ka2bxQQsJU9Zih0XlgIJCJ26K5xzCRKUb5KhC
bvH34Bddwcg8wzyz2RvEN5N7M60rnLJ3KD65G1xwOdQ/GzQ2UBAj9wI3uGLjpLaC
5m8UI3lZxgEjZo6VZvIQt1KsT3ibSi8SYkjuDv85aezAQTwLqp+OvX7nI8ZyneiR
jR9nvwoqepfIP2ssVpuxHGFLKa/tDCRbdDNOmxoLJXkQnEvzrwCWZaQWF1a19eCD
+VyiV0Vd/wxvo/ybKnRizECNR8Z59Yy23VRaZs0hQKvxbyKqGE0e8ncVEbkfWu2G
15Nu8J0y7RxK+CbJbm6FeWPSaRWKOFnz575jrVggPlS8nAjpQclkgD8adtPu/pXS
a/nr2qgRY+ZkIlB8Ze3RfHU4SPujakPJM/ueQ5LJWuD9FaK+6mgMrWnbb3Ml/7Mp
111mCLbvHnKqiYiuyqeHW/jSBFkelDECdxrOB15U4XCOJEmRgHSpjv2ghDb6edZr
p3CYh1ZwItZpnqm6Ok01tO+XlSgFj8LaaY7tPT0L/xG8CYDdwqZRhp1OJqw6MLcL
G3a0caThK8hSCgv+FE2p+NPVpXMmwlAnPCudObEwyBVOriUWHgD0CD7kOxwFolA2
SqpL4kHt7DiSP9ab9hww8xfMJTklGDcJQzCZjTEyHRZvXfpMDqqRwu260FnLjKin
7MxUOZdY75X5jyQWS1Ph8pGhqPb2J8WzXMuug8lrH0Pgbof83NfckhbrUvEnaVhW
MnjQ6wkrE0pqOSppwp0gZjvMaSgmvV67PakyoSdqO//2siHs/ON6u+BZ+XzPPN6R
H55/dhEhMY4Z21XK1Dvk+5jQyJVWNWClGy/JiRTjVxvJ7XvRzZlOjU9EdsC5eb6S
vEYNgA/fWzXUDEFIvgqMxMARESwJSzgDQw4BId4v0aMQkWTfnzBrIWtRwig6PZLn
vOgpSlY38a8MymLuhFMZ+iYocTpNYKP4m5syw83cpxKKPpFqGfNJXeNIYtj0Vo5A
crfiEtYEblCtXyD/QUNLl1D23GkGeOMTN64DhqZiYZvYFCrh9ew8FJOvBLuT7edn
2ludf31qt2yErOc4Bcn8ZVqpow4ofO97z1w9vfP0CbtHvL2v1JD+u1yGE3o4vd1g
Ub2pdDOaI2aWC2caztllkGTuzb17ATp9vEB8IL6pSMPqIfmVwE/2g8wGhpkoPh2i
oBrcUkFvURS/7w/zDYsu4ujpUFtG9xboDsC8S6aSrwpxWwa+lXaJFAlumACgnGz/
u8kEh07n/0t8yaTfICMgkmIGpYTZsLgS981GstksOhQR3qSm2YYeVfy183sdoi+a
B9iC4zBHo+rrqZCyvMoZW7VlUsW9TEgiKRGRAOO7dF6ykTemhzU4v/xupXFsC4wX
TBjosxI8rcB3HnGOmiUHwf/oMkqI/UJoW8WPAprfUw8sy/SxxoJckOB1c934Sgp5
F++tLgyCC5oYJa4Rg09YVyT3AKLJerpsIDmhJ/LGR4e5+wHMOPDcMP+1ICixbNUR
oR6m9w86DIbLqyK6rq7cVe7zZV6u8+e2trcRTDZD4DhxcQ/Ak6VXOz7mXuPuMCYt
CoNpaDrWHDuSUKyszUlzWTfRj/7zNdmyGE1zA+IF4iqwYNPbAp9E3/RkVP8DyR2Z
U/BLy/XAS55QjvFrf3bStjxIhCov9zqAfT9iD9Ac8lC86h0YH6O1Z2YJ79d5TR+7
ufptGhNnKV1h7S+LHImC1Nng9YXRq78HIZ0GqfN6yG70u+5wzZBsdO0GiyyYCNws
kYKAnlpO2e0wfnhc+Gm6s45gEqTbX5XeNfM58Wvc0CPU2kE0PLsXhvLrSmgw6BX1
cGNr1kEES3BnRRkrBKKZC2bFwT9ucxMh2/8BG3K9oNTlJ4Icjg7JIflQEKMcekHO
C4Y40/l2TVibe5T6XZT2AGw0kz+13bqKHlkNcpZfFCmaDVjdJAQXOeN0aeLs0lOs
DbwcZrTse0cdD0J2MILYNj74QgdOw5g8au//UlBU1Chhvz9jQ8bC3qAiNCwZjdeS
rosz5GGYf3X+ekTimKa6H/JqpP68vA/UL37aZHN092AaRqqs0hzFE+Eoyqg2kUji
f3yodnlstd7f+icY8RuT/CObunHzWHsvoG9Ivikivon+rl92x4qEK3NYgZndTKeK
qhIq3NG+149jm+NfrL1xrSx61xQofOI9TBvGziRHpCZUY2UndxABrIC3WhOf6GGg
X2QxqmuoP6mdXYc9zRP4yk6Oywf5SmAXVBO9KamaZmgri0iXIWMg5H2z5VbYk+pZ
CXvtPNqN2T5QdhOJiHbJ4VMcu7RcArYBeXjOdobMenYq/svJzMMPXwKHhJRX4eGm
J7O6wI2XBb36gtKELuehF7czoi6HHK5iTZkJ181yF7+2b+PNqEall26VPZFg3hdp
+hzjBybhG+tgW/KtHPd6E2Qzg45F5aPhweGgqe4BpPPTIN/tfzI0zq2CADVrtaLS
aNpdtNU6ivOxZzNLLzG3UbhgbJUHfJNR5yy8X1LoPwI7K7FzFC5a8WYl/vkv0L1/
r+50Q5TYelMy8OjsgT1KUjCe0jXClTp4DATP+TbdoVRikmf/yRhIiX/Sb+VaCaUB
EaCv/DV1+X3fSGM8Duvt2rd2LVWcv6KQoMldEm/hLG/hheeDUNMHCdL8sEtNCezQ
E4uKmmTpvGdioDtxeg4eaVlIVu7/2ZHWxbDDTRzKE83/VBFBVbsQtct5h3W7anlI
erFMUQ1CTg/cQK/Tal9AgiDHSm7L+R6o58apWvQ3/pV2akk/zCG0lw9C6O2jt7SB
Px8/g6gaVBJbbpNMzH94F6/9OxuCP+mSD6gZJAqZWNmbFDeNvYnTP3OFqSzUKl2i
Q6gjhsuVPKWFOx/EuJWQ48J4lipCCDkqwdVfR9rgy2bgOcDQpkcWf41MeIlhHkaE
8FvNEOn28TNBf/PbCRVKNQfjup6VfHJOAROTK0X6j2Px8M2FiSTc3PxLoyIx7MPq
fmqM4t3WzG/MKX0HJxcsz9wujNYOPDWFHrQTyCnL7YoOgacVV5hU+ZcsZApGjrAR
j+JrwIb5Gw4rqWLzMx3jw1aXpiuwAspaTqvgMKKehXpSWFzEpyXUqG53360/CMF8
hCINnIDDr+wqoQYhZMjAahlQiQxHveV3L+uvbCHHs345AtYShOQJWo3o06varJg4
D+5PRVCZgs9V0f2Zwr2ebobIOdTQKZZMbIBFyYSGNSVo+upZJnLNQoEGIpEw8m9F
x+u2QLUUUe/1/8KUR33ZkUSzEd1cFbkPhIr7RsuJsgJ3gTXBe6sGZcnPhqA2u/Yu
6Dxha6GBM9F9ACwCppXBPbGf5l93B+tyrj2DMAyYU1Bh9FLtJbUdG5ghmyg0f5Kw
LP8cJQWesPf+AXoxFCRrr+Kts4lBsEeXl60s/aKGglPdsAlbkpmfIIgEnJHWoa7e
gHCrHhd8W+JMbDhxTxwINsxK0HN1u2e+Tk1W95V7xm7vHPD9zFMZhqJM2mxl6/Jh
CQ70THkSenbBMok9j0CD0dpBp8YeXc1Bli29LSEVziBiur0Xy2s33hVGh3YfYQ8V
a4xuXKnz8CszoazRhBkMJWyK0qY/iTzhiTZJv5lE9tdMixUvE97KDBWk7k0pvv20
Z24OrKQ/R8txZIFUgGgG0rAsyLN1JoaVjfG+jdhcd72EQxBODE029TFqv5/Pv/B7
l/dHHUDJqyo+4qoJDWfmFz0CN/+vYi6woDI/J7PLsNoVtwSC0MWsfeZ4QfiN29Gi
vB9rTyMdMSd9/ZCiGWvvx1ULiwVpxjFklDiwpyrOznAWnyekDHoeDpRHlLr8JkO9
`protect END_PROTECTED
