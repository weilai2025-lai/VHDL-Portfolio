`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUw2qriqrF+aiHUKTpgTq+IUMyh87sTjKWgugFsaVoRI09evCTFWSnx3P/SwRYCw
KqG58bQvws/XgelhHmztA2Jv599d15Afy/zUPysK6CRun1VabnnRKy+EENFWhOy6
Uc1W8El7hltD2HuD/M108iB/jQIX9/OIpq3HUv0IABXlJ5qMXeqh8PD5GHNDz1NT
NSLAnnUHV0eZFqgHxnKMS4Bn+G68HjwOW5nHwkPXy4id16SFfs1eK7h8Y3eWmuEz
9+uZxhsh2f2MASsL3/Wo4miZ4kQy5lsIAM47lAKBra8zFi7Y2GjrycFtCYm4cttR
rk4124Ad5EBA50PBArsv1ySWI6mp6JowwIwe5UyU0FSMbZ7SG82ICM1XFMv0MX6g
pmmDor4YKv9HKC+Av/+qn8Cw57YeHEK2MEd7R50U/8wn6WNNun+pqcWO1uJcOCQT
XKMYo6IKKcL221rXxpA5xoryHVttwCr7MV4oLESNaAVkZKZlzSjhEpDXFYN04RLT
pjXhUvwRNmj3DGxJmXhBuBnxtHWwh6545nl7bVXJgMfdL3ui6y0vhzTLJrwUu5GM
i8w2WYGIb3qlpf5+5js9DdFozuy5B1/j0nEK137v54Cy3A4yHBoc6oJvyHkdnMTc
et6zyOAOw3q2dZ7k9+vrqLDRz5zMRbAvLFNG0xdC4URKH+m5/rwa+wMPZfo17DrE
uBX3haYv0BfVXOoqe/qlQILgJkiI6iPhq4gefIXzOYSpleyE79rF5WKr0QOQfd18
frdUyQQ2RYM+tEQudsA6U3ZrW4UbQWUdez2xeVXjPLoZrx6oFJexI130NGaU/rTW
ht7KhBHxzk/ULymPWzwTyZrUxmAxQUPah5JXGqNXKSb6xL7i+IANr8GC6ccCzcWe
v5zXpRCeE/4QHntJ4A7ke3E26Y8GjJYWDt5TwMpWmiSrR3ncIbvMgv8cUTABdcvT
+f3p4QxCjialuqMJEp3jgrqOZ1mu1rCK7qHGSYexZV9Zj1iR0GSsJVnY+2F6efYj
lIBXB5zoLiNp8oNm9F94TYjf/n9kQntmMQEMNR9zlUGU4scFGn/EKtdzGX36QH99
200JUxwJd9svvZPFv9zlwNzfK0wc7bU/UYFIvbzmJR+m7BfKb/LEaMw9nAvftmG7
evknivyak9thzKnLe8UGAw==
`protect END_PROTECTED
