`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F63+wJD3JaUmHLp2tc0nxSqFxbvK883VdEhSgzVnGFoHVFlhPwyPGjkgHXv9V7Wb
H2uUfhOE7QPEtZrZVHMf3H5kPmiRTAS3XsfIxctfcjV40Tp05RWmwx2SUanZUFUi
QlhRYgAm1t+RLNSKfDJMBZQqoBODXdVY18ExUbRRglXlVFl0VYcbqt0kW197NtkE
YyLltB3M1ZybQap2jfpqWPjBNf1vAnMD3ozn+Fl31VNmuBFLj1eBu7IRTgSqxiVo
vc9wQ4w2Ycj5mABRZkibaxCIuEkNqofUVvAd0GGop60OyHFEu2FuwRmDp/pCFktg
CJuxyLVlXGP6BzTkuX6plIVEtFJ5cU+dGdNcjcsbtGjpkJsiqBv5Es1UavrMdTam
cJOApYulHstm4LP1jpXdGBpWs7AjP6cBueQ2mCzP1rQhkLQ8ZGjl10cJS8H21R+N
9LqLZ7/cEZU/eK7ngB4g0BdciK13hkh/98YABMGNNEhnWwyCNaQ0SRtaqsZFXAjR
s0Gbyzo8lmThtwO7wQjzQ5UMuZfsG3gJGj93pL552q1D6rINMtU7HodC1PO1ZMdI
JK7fKzpuNooTL+BapDLCO306k1XaAY+HyR3GDr2WZdCNos/H0dBpQc7/rZ49Qxvm
UNOS6E/NSXs0t6BqdnVHpQL6vwwn4xYhCaZU1t7AK/tcUeNY8jYf/9nlxnQoxiOG
bxIgB3UEZzPlZKLvJ3bpbVzyAnx/NAtmmgmnyE+WcodRoUMqvSnYn2bJIBVBbP5I
Qj0UhUx7DOAEE12yXxzeskLxjtIN8H44SLzx2t2EgOIMFRu54vsIgBjGlMuAJYmH
3ykbpEvwYQYmxImNc5QQx/WNiPhONm29shhg0E5Pk3I9PjY9SovH8w3/Z9oOPCdT
UUPdMxugvqq6cHlTXpBKH+x/fR1TYcmgZYe9EHpYU+klA1Dy2V2nMxDaw2scE+XN
4U9GuP2LCr1U4NdrFU0oY5l9e8laM3W7Z8dUVPAw3gCg54Kk7aSGO7rduYCFaGiH
99F8Mzu106MQp50cctbX2L8kkpCA/phsOPvT99OoMBKFJtKIZ5pd+85Dw3dwUeTy
HOGLnnGREkkGTvjQSvXVCm/OenNKA5IN0fUdWXRS5lUoS0WJsNoX1Ah1udedBASX
CO4E9SgQQl0J2Gkh5FjV8vfHJveR00H05FZ3EdbvW6rHHMZQzKUX1FjLBfR9iuwU
iI/kFSB/VU60Vhd2EvxQwYHj1SLMqydVGr0kE9ooyQP+uMup2BFs7HXF9EgiAmTA
Wtki7j0tui5TyU7oKCp0Y+koHXLqLzYf3Rnq0AaAj5TJpPJCjN6V5//AGK2JmnJt
o77haaY/ME2+bUhEp7Pjz6FbjRzllbH5ciKYlzHS1LhlY0QtSWQxzCzGrs3lGl/o
`protect END_PROTECTED
