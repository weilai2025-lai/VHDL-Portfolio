`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKwu8JL6hVPZLpUjJDCxLGajBxU7xwn35MpxlEmpH9S1nANQV+Djm3nB91A03R5L
v1EpaivFfi5xVyixE1EkIisWAJf3VuZAbHyX34tFH/pwhuu01bGlwCZvAGi44DPW
EsC+wZaGW9niR58E9G4z9T6NUTWyFVCY3N8KHBAVqLuokwmwYBK0sk4JxDFyEN6u
qcOpTb4hlILYgUBC3/7nuKgkozW1WTuVyAgASPvU8Rt2uxJMhqzgcJDosarfi7zU
9hoyq1ZufDM3Vo7oI53lzHftU4y5wy2xUU0y4AhzPqj2hen4ZXjDstXDuJDkrxbc
KZqZ0RAJARiLbmTYQ5OkQLi6dpXsX3wBA0lEUM4SWbKI34ddSvgDvDIBrf3WbBld
vXohiNKsBNOogfM+hTBdDK++sAs4+3O0tfAuUbZ4N0OO4QdjWcIZSwLSAYVjq82c
IIb4Ovfn7f6o07/cPRj1XV6cG0Vp5A0r+yvfo4rxL1LfKfnJwyY70zRU974zOjcb
tFE3yskrnlZDORy5YXPlpAP8YO6OxtzXWI3ZeE1rwlqEhf+aMgwz/gHJCgzw4OBK
0QKdm37ro5vBMPXTLPy6TDpPrNj5ftcGLEM6BCfPpfyY4GpbnTDE61YZIrTaqrNS
JZGpg0TzwLKRCWleVozK/20TUiRaIKC+V4EwjFK9kdfBxIPA6WOsQEeWP7w0q51k
YoND/FXNerI0grYr/LPtHFJ90iW6t9N37jN5q6pOfJI=
`protect END_PROTECTED
