`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esl0nNhQU5etFeD636a6PpOd8uP5p1pAd9jYQjE/p7fk9Zr7YydDHo5/b13BD7Qb
ltMgfzd5rUzP85VUMZqDeO/8kBaviN6nuuS0F8psl2Z96J/8qiaONdS0LqM3zFOp
diYtxc2/wdnOxYgwqsFGv+BgDHojTssLcL1v0iMiSf3bUlobJ+/SsMVYLdm+NSb9
FK6rHpnaTJerqLX+LRzfbiOgKTQAmdOUxyNRLoS80b9q0ut3zqzO/cWYOfkAhH2K
T2hu/AinjdEmlpIQ3vHGtDUJsEVeh9dGIKqJSvcEepU39IHN0HZaPAnvfffk2RBk
K4Ki5F7RxC97LnP2szWMs8gtDsm5Tlj1Ua9UfaEKlKALY0kwKzHUlrho/K3Ba8oI
RDPNk5l8Mq1XCwStbpqG/kRRSE7APxVUEy0Sc4vQEgfolizmo7U4JRn2UCBkckkM
XdFkaHwEYqK1TkjyAoQsTn/UUd8mjFrdVefq+guwPp7FKHF/UZjiWCJgIBPyOgDD
pGTZR37GyEvYMtEOurskk2kvADpWB9W4BwQ0qAVGGmruz41s66wt2tMWBlW0MKPn
6pFTq9WlCbCqV9dW8aZeG6aTr9ruFtEHM/1LaF2P75IPBF4AVqZTpiiWUQhKT1yr
1TYM/dvbgMAC2DMtqlMXGM4sjqWjNkZBgY35LOc5BqcOCNMTMbDUKcKT6HQjSJQP
UjrEZ0H2ujF/+Y+D8Ez+HjjOBD4ZprfwPW+M75QWL60=
`protect END_PROTECTED
