`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6wVAs2Wa8HhCwRiTZzbAYa6Ysqk61Fi0z1JVEnfS9mc/fopkKvwMPxamG7rx2OD
oQKpBuOpc9Eoyp01ohxukyE32cxteHGiYupdRdU6CWOa4o2QbambA1/SJXC9j0Ff
8XmJ8KtiMISQKa7bOdo+xmcBPiZqM5FARET/jVkW4J6LgFhJFS2HpAJnGErgsQZ8
v89GQXh//VsG68Cj/s5Bocs73tm6/r0YIM0fn5k27VwWsbxbzUF2wBli7chJ5pCD
1ANBALQZ4NHp8Vji/pmw9kpz9yNeazovXo8wFaLRDE10l63Q8/NHdQ4tehR5gZiY
cj4diQSTbZkIw12ALYlGg9/DQTXnrQ/M1AXgDRs/QWZJvB28P9Yef0VDzqwj8EnF
Nl/AJbDVjl9SrVuWciUm1BRxLOg3grR4tWyxzpeBgTSPxLUYbG3BUR/Lk84xpnmu
ZCQTW7Mh7FP4+S52rLe0j/27AFcSy6V/DxdUSj+qwt9PIYhQ6w+bnGQazX2zrHCv
KfoUSoYIDmfyiPGAX0X1XH0uJnKCJg6N347JkiXwtAMXXHa0rAvA+rk4Qblb7bRb
eC6TMU8sA31/1UsQUPAezn/meq/2l+ZQ/ytqJUL1XBlKooS6Kr56Kfn0C/vCFDYE
lZ9wyWle8B6o5Ff7XKR7H7thQuDuqcnp1GXwGmhrzbR2B1iT6MHumFin/04qReyc
`protect END_PROTECTED
