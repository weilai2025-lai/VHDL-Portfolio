`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EnCl+4tRcyMxQSu672ttowH+vIein7dXQad8VKy4nc0Tw4zViBoDqm4aQPEYBe9U
9WkXrjS9H7LI+d+f9rohWv9LYwo0D11DhU6NJ1yjru4Oqu/QSCVAaIYL5irXnPgB
3Ffxwzmnp5J/6mKpbDbtX4xfOTeKI7yhpGsMqIDixniuM4bgufi08R4Yu8Tx5BYv
mhh4TItIugW1X8aKb2Z2GKaxXjFnZDHqSeJjgQmeul4we+ZvuTS1kkp8NBkM/k/+
k6SNchO1QSvae32Pj5Zap98cWzDBlCmHXkNuxxND6kvtk0kdHmR1wMnFVKTUhISA
AQ20W7pQrTqCZv4SRn/e6CUftj4Uxi67fzfLQTr0kSSM6RR27qN17q8lB969YIB6
nM8MmwNCY/L4M5QOKMp9MGkxr9BXh7dD5k33qykrzaC63oK9HRa4YFOObWvTKeCG
7YmXTfk03GyGKuDoun7v/w6c8oEyWF8yW4xsaVnheBEP6nrxoU+U9f1RjysMdeFl
tmPGFXAN9Dj0gisj3fF8iZhH8+dHHHkuwuWGxzS/6S8tQXmMS9mfWV/mJgUb+lQs
1QCYCvm/2I0X4Wrduk6NV7Vdb7c0rozGK/G58W8IRyJLicNpl8whNNpcpOmPis3y
2NcNCXay8sf/4ZpDk8j4l5c59cYsak5S3GhIToaZEA0HUyNqm/k+sQqkQ1ZanebC
la6GE6UMzsuHmRxVt8vcDX4DERGKZVoiaXGsctMtHG1uuG2rpUNq4/9p9IocKPKK
cjWwUeM9IwEzjEsV46OJBOC1fpixsIbxAoLSkH7a6EFT5NzNMZTDQEloyB0Gq2Sj
yljP+8MUgBhBjirfUB3hvJ2WsiWiCru4I8BkO9zWn0u13lOlYJczB5HosQ/3B5SB
`protect END_PROTECTED
