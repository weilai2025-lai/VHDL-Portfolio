`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gair51HWDM0WG32VeCQ4GESahEgbqdnL8Jmyo7dJIMtYtoYbTaz3pV9KCG7WBVe
vJoUgxoeFIbyyeIX+IQW4TmwmVoVz/OmXJXsKjkWgoG080HZBaWohs5GnqoKedJT
UDKLeCrEw+jbf9nKiT5VskjOW8sz1cZgXrJAc/Tb3D5CkOu1FgQrG+gx8/M/JNE8
`protect END_PROTECTED
