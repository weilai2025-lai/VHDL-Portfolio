`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ynbbbE7BAghV1Cv0gaKaBTWBTPkQZjnDvWD7otFBlRI9e2OvoMwe7b6gWBZY7vmL
55lcOgpXa5h4pIvTe1qo+9JOEUjbbQ0RkISGuCwCqCbktiUs6hZhPxIoSHhaYpY2
2hAWeTYdaYVTjxAoXv8oOWGK+PKUhSGjxWn4sAZcapIDgTD/MqIdPVHiR0Hz+yga
QCBCZ+iqxswFm8s/CTKW6rBVdQplIcZfD5pnQsKXtkcPspVCuMEkg9jrSmHVldyN
IdjpjZhtmLzNqNc3bvzbVYTZKYCQAruDCeOEDlT0xgh4rk0dvzn74n5gIA3bKf4I
QfTSGl3d//Kdx6HWgjdFypzpA4hKSKXFkr0TCblwGcqa3IpKc42lYrprSRZwVCoR
jw/+C8lujAAFDT9yM2Fio2AOc9h1Frx7aPVqagS/kuxFgeDwCWFZtRbHdh9KX2kN
LDE0+wqYP2wC83ug+N7nrfWkhE11nGeGaCVk4OL9rmHBSmsyBJWeBCnktVDMcS0l
d9xcpCai5bg7b3j35VR2mrl/kduthcdcXCu87YKJPSle8ciDyQh7L296YbZ+RCGy
uHDKjhNwrlV92rHNHfYKUV6QP+XloZAx2VeSmoxWDHaa0jo5q7J9dbQ4xbaLrnVa
gfCgddixkfxsH4aAq8LPpmMr0P9gFIwYEbZQKP7IqYeaGIFaPTpAEc61EY2i3NXr
PG5YWG3dqD4Qhw7+CNHjy2WZK/BxQCcVIS98kN30dl7BxljmxOmyIVKcd6P2xkwK
g0B2UDtPSMeZXIMnafVSrTqm6g6nJAQL8DpNArqI2YnaTPPgseAHhrR+QwuQxiCC
oyJ7EPBqWKx1+NF8eUruDw==
`protect END_PROTECTED
