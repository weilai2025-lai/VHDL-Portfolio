`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3aGdp5BL3DUO8D5WP8A96LENlvJonziT4UuJAuJs0s6bduuxgkoYoGShlxNr6E3
03+PnGhBHjgHdy8hgc9Qwmqynu9OBzMun0wL1CcEZwmw1zqCcZ9lbgJBKRg2UtJC
t6lWBLomFWWLJXWVgqCnHGEZMr+jFqeeY+fzaUL+p2ATHXK7UEd2bwrZ3gY+oNAi
P9GNeKaRNULCwry4Oe1AukF/p7RdcTtbuz2RX996a+E+0Gyxa86a3IMtcqXIhLiy
fLk9nImzXpVGfVuPd83RCUyfwE5gVasexglTDdLtQyUHIJqpP17KPnBXf3J+b0Wx
co2MUOJM8yrg8jDUh+hWPUmbJO1udt+m5KuZQE+HU3oJ9i9/vyczRbYYFsvgBoOF
93TdelFXOc33JSLJmZoo9Q==
`protect END_PROTECTED
