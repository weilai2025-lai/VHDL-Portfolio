`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAc66IU6aIoMx55diE6Ik+1l90TlAi2aEwcQCDjUX90NZT7fK5oizLN9vsdOIgdm
qajK7L7N8/elv09jUzrATYIT13RtH/RuPH8EDyHpZC8kxKZBsi1wuek2yAfpVaty
bEPWOvFzXGKhPXGndPtY9wDRljk9Q6Xrvn3nz0nnP70rUR8WmXX7DeOtLinpgKzo
9UzKMFt7fJ/n7IswQXRghO8yCfmW5b0GFsZpM97qnxqYIxqhKlV+jElz+Y3Gs7TI
qxN+s/pDni6ZZVVvTDf7b5RtF9PowYt/5HN3Qp1ugQ/UU3tUknrL/7qTdjdyt9Ax
c1Lks31E6C/4th2r56d0akTJnMtLLv/hoQg+khORMpHoTWCdjfqJTclbWM9K7bWM
Zn2v05o2Um1qVAsWvdhhUEI73sD7Sz5w8FPkGFNPHVOLf4MBRYx6R4V1wjHepfq9
rfI/ztxLmoGdncWOMo+3pGgXJT1yv38X3GzqkKMTu7nCs0Q6tP2W1yL0XBDS4u02
S0DkL+HGgE+MvKUiXj+nOvq0UtZebSy1s99mjOt9aNnjeMD/1OvZ1z47iJzywoxn
BSquBgg+C92ARIUP0ym+hVqWuVVWX7Fmg2CtBZ0Pu4iln/ytfbnmB31eq6X2sLo1
tUN9JKD3KtYW8PofNh6xt4qo8AND1I5Ng8WKW+odu9SFIbKaezBpRMjE2QUbEWXe
IcpRnvx0HsmpmaaEEZOpWgdllutxCfLiy9H/Tn5HUPz+3Q7O++wPkXIZqKgjkBij
QLX3+Yp+bsElMGsvenl4Mz970XH/rgimmdemECzb8+EmccVCycvE9FNaFGqSHbGb
+bXsv3TF/V/TPvoxeWzuaw==
`protect END_PROTECTED
