`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rojuiXGQNn1PPwIAiQBO1pW72jqHijMPtq9L8nKIFbo1ziDTcZ1ycJcyQahgM/lg
xnK9JuhUkZPa8bA+Lv83rbGRDrDAKe41So3vIzGKupVNPhCoAzAnMgXDRfCF0r2c
ZLYjCSegpk0OlGHggAttFkBj2Gd7nwbKPUR5YxY4g1h6jYFh5dqxqZWggoO/pYNh
C+L5qHMpAh1PLIxcYZtEwVG0simqqtp470F+Yu9IWHS8tn79g5pBdNnJo44ngfTH
63exHrc+RmsgIZnxDg5O5JBLQarFewWdQStS6rUdqtKU0TyiP4xTuiamvRPJnSdb
nCLbEjLJOWo4frbH5IgC04owDGqZWmvL2yNRC5jf5/VJrg9KRhbtN6Pv4u2V7sLR
CM8FdMWJfMJ8BLPpAXk+PYTz+RuICvwYj+4PXmDfc6QVeW3bey/jYJaAQJUQgzui
BHz4Ybt+naQtLJyXWirnWy0ZbUWwT+JBDxN/vUlgoqIRwG2kOCli5EGzxUQBmGr7
DDHi1vEmAVd9UDMo0m8SWPyr3x2s/RVf2qD77XWszzbKfNJaXLo2bdTlmIMV6spb
z0qFtFfU3TSLkA93dIgUPAQVG5uWq/JCOCiP+rGJFWZg5pf/IBBbnpOULiozyVYF
zelxz+b3DlVtsK58myMs15pHP3hz1QedY5MRLOVldm4j7wenBYcLCj2WoF6pcHmd
D90ou52H+3kBMYjxdLFoNjvp/BHMDpVhzyRWKW3jO59TBHc1ruw9S5taH1ZEfJ0K
etphpsCOY+YocC4suoWtJIdY8Wys6m1MtILGFYYK3Vx4nL2+wKWGeOPBFX7pAQVT
QQ+5OMJxPTFc2W+lrqV2TvdQixZ74EQpIuv0mhpy1JQ2Dr+SLurcIE28a4G3MQ9h
JxEgL0ryNr8ZfWn/+JEXWVH/ywYyb3qrqp1PUGtehmE2UeFMpaL5cbdNhqoJrmJd
0KxKUoaVW8Hh7fMJwB0u6wPHlP8xKZQbI7yTfpPgsqEXjNgwWV3Z5m2HAb9d9ljD
XdMYhuS0yxOeGCM+UFzDc89pxISUeXjEnCPP+veAbBV0pSw6EKQQgiDk/4T3L0s2
p+tvyijN0rvGSBB9Apq/+w==
`protect END_PROTECTED
