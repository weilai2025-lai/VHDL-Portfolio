`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ECoBlnLmb7IZtHw1/lwCgQnoieaMyG7oIxVRasQZC/Qt/06IvnlofUdFssgPCWEw
4LJ7SH/yyt+zCNN3tXHABSfl5jhmX4m0uH/itgk4LdXDrO0BMr2cjDvPIr+ZT+sE
Jo8trW7lAWBb0ZN95ISYEo8IIXKEsl2/af98QtnOQ1L0F+PtJCfcx7ejLKdEHAnM
WsWeFIiUyvI8dYc4qkS6Xb9PUe0w62I5iMM+Mcl632n16tRpbZ7hMcxL9FzTEfz5
MpE96vcsGq+GneW2ocS8umhmx/XLNjpTdNesJvDfiPGJ5kM3dJfhYQWG7UdtiGl8
uccYNaTxKy7DU1sw+iqd1YM1oQORsruQGyBGkMTj1H3QJcDXWpORiS+xHIb+c/X6
b0cHU7cj04lj0f6V/b289o5tlyBOfTg2YRiruPeLa6BiPzzxpEh0orS4C6F8s/G8
s3EOU5tOCAm5BbxHRUCQywzkSNKHJoV+G900OcvWmeKFFo8KuOKB1J0P9EjDRFOQ
74406wznk64HxLQKAGWzrx2lzJYoiaa6jpFCMGy8JoAEg8Mj2qL0OkYjaC/Mna1G
KPbfJH3z96VE+xNAwE6pZUJwVr1l89mpOuoOM1g5ZVkfKLe0d921ZQlmWURhT1Cd
bGrqBXg0bMbxe5685b0Uf5E2vhR2nfsnFuCd5kAhHNweoDiH3n8c5JedJFnW7sDl
z8efjYMRt5TmU0/uhPkCPGqMB/4M2qJZnzQg8JDLyJ1ihVLSkJ27RF22yQJhgCUC
Zq+7vhDkxh+bM7CF8TpemlVHYUCLGHvTxWN990mua34J1ihKZL3+Rmlb5zqN4VxH
fekFuBlc5EypGOEsobGLCU8rmSAmsPHTfCnfrbF7Zecm8orKbjiZv+ifR8udCPGe
hSv2IYdinArsqdvVRlXIgDsBmvcb8oAsShud18A8nE6nPePE44fq7MmOHRG4bMx0
6bGe8PKhsSEi2gyWs1noZiKrYEHNNxfdHPUTvwzcr3rgQn/M+YoMT1q+78C6hKUg
BL5gXMK8krplwDfkWZXwAeUBiZ53TLv4OSDLfRei61Yog4VKmSZJNzi5txScVJ3S
lPq15FMGsJfT29ZIaTp4zVzNOeHzgodydI5ek4uvqmifi907kLro+YIYrOWz4EQx
+llpk1isKeYlZrP56K3jAkosB95WUetKZD1uiZc88SuZ5ua2fz3M6oQBLiJVSnF/
M++IHPLVGoPYyQFexT/ZCg==
`protect END_PROTECTED
