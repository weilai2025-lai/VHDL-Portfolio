`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1uNkYuvvl/oiCSISyg2ZSCAodEX/8NieP/ITf17LSQ+tLpLje4KKTuSiiDjHmeU
SMRjchN1dct9W6YiX3YkRUPePpiLJik5SiQf/3QddS54qNV7TZtwui81qypf6ovS
YPo9gDua28EObEn2bKkVI/oyh799DTwtvpjQRYxU2jqCyh1gkmiK9NXPhVtxTHux
t1gqHoZkLjptnuA7GjQ6Kppqq5jmolJaBA321byBCvZnR/EcZVheW7o8jEjxmXqZ
ImX4Fy2QKvUNY9iNOX7I3BZgy6WRwdFegGTMlQB15RkjDtOIQEJSrV6+y8gfF98a
FmnFleDLycLOm+YT2TAoSTLrZX61u4yLCjeOX8Dzi+0LFWEnxDunuCuBLnf8/Eaa
KRUBd8xJQaN30WTFSw2KEu2zr4yJhS9a9SUM62giQHoXd++KqHgQ3AQY/t4JdAX1
Rm5fQRQfSsGqyvexcyNPpghmGGOAotKa9etR83D5OgZ0g2aBAUblTRjQPfVToM6a
QCdGRWWfy53lPRH2HiOvwoeIi/eMoJi+9ZB+xq1CsPwGq5N59qfl5VQZPLyEKwUU
WdgwAvJzBEDpicmE6QSANAmgUOTvwyFG+e9wi/pr+z29GqmsBIJCkQ6bixfb+f8m
Tski8yOGPyZWPCgYJkZQgSWBjgFysIt0GUaMnMjF2Hic/fzyhUWiBcDR8iD5cyMl
5FXvX748o9tOMMIQywSGCoHn76omTefavd1azYip4t4FI0rD5fgeEvkXGtjl91nR
Q635DvCYCJOdWT5I5rHrTITPQbo62V9eyOnmRlf7lCmQzOzBSRQyEDZMZNZXrPWW
WaGzs7RZsIPIkHVjRN4+7W8CG3XSVB+jLJsY2OefzXb1XzhieXT9vZjZfn7sZ5cc
H/3OMapjs826ZlftmlmXcv8BKn+YXNDaFGtUQtyq4CLUSxlaMOclF9Rn0xYcqS8r
3lhTeYxvkTuTeJxvlpGOhJ1erZnlXKTZ4+Ham94LgT9fp9O0YBDXpRi14iTbhBpG
EOhaVNdBy9OFqj5YtiRZV/WWq/xFyqa3dQwbH+XbAX4iZzj5k8HaaPRiAWR9SVDg
HVcugixMpi98RJTRoyqP8yb81TuhQXMQkCXVeY8dOGhtE+jftZ3eOt7zrxcYBDrI
7fTIrNN5cuWD3jiSnHALiC6/GFgCzMS4yKgx1XTkpkzpZiV7tQkW0plbg7BM7gNz
ES2uJuiYXZw3hj4waZRCRpf4k6CVIzc9PhAWsi9OrF6ZIaAdSRqp7IaMSYDzo0O0
rHCw9jLZECXRc4X+DRbZA257/xgi4RihgsdUV0mwhbwDvVppFs+fw6hj1xlGYZ2h
nGrDP35v6mzUuf6RkTb7liFYNjDEonmGgakcXc50H+UZoLlwdZDL/+Y4hBHHaqZN
OBhuxIG2pbGPlpDNURBo1D0BjngRx5zeX6ETTZWaU/ZagJMPx6nU/2MPMVLrFrqu
tX5VT7ZtfjSmcFt577yK7FWqdnX4/TybSKsnGe/prvvLe6O5yqPGdogck5mhLiNM
xyutKr8SK2pQcneKz2pio5DNhsFJiklJH9c7n9tAjgDrVklAJl9B7283zoQ1bgop
2KLLQDuk9Eo0qTdewBV6RLObsVMfjz2tWxvGWrB9kIVMUzIzUPSEpALvAs8WPNu1
pYKfwQMrUsb8IKcFtXAcd17Tq81nvpaeWDQ4bk7cxxLaH5ZA8Iq0RNI1hIU3zm8s
v4VJ/tJcpTdtOEM0nB1rO/SeSXmVUG5j7zCVa1KbCVI8gt1XgPYVpnR+6wcdoGtF
rYlPY9c65s/RJr8U2Okaxw+Ozk0YxCYxUKnkqnts+CMAlAcp7TfuPQQoTpDiUPMr
TN1vULABnG0FBNuyQbCgTupzAXmxLTi0ctt70datCeOLLYafOWaYoGPzr2VSjDwS
VtWisTPhg6W76K2LlpLWeZdiGmf0pDuUr5ErEnbS6+By0dGqGa8oQUlaJY+sPQFX
K9lpvL40Dahxyj5pduLauaFNSszUfyakTyyYLqWUKS9WCs2XNP5TOU4TQW6zJVVA
cHAOlwWubn52SoK9eYeBrsO2MEtmZJyLpGFeGlBwPbeDjfGl6+//1ILsEtbXzOK+
simNamJAaidk9lOvLigHRLYPEYiRLCrw0Of1q3PooYVu7rlIb5CVRSVs3XnJvvYE
/wCwYPndFzLE93ICPMyhDLU7XdMWHaqijQgrgwnOFxJl2LlOqwbM6JSiaM/Ixy77
eLeGn5iF2rQoU1gk+x8UZgkbX8I2QHweoUxGXHLwj89uy55co9WO8iOZG1fs7gJ1
W3YD6w4/O8826QlblSCxryMxree91xS4OvSwLt5A6Hzt3PImK6CjuVi1qa10mWI3
hosHvdAcWYqIyRJ8ANp2tmWtOE7KVqYCXxpNLw4rjGHXD0JM6Xmj4+MAnqaPbZ8t
unWIfym3BPx/Y8EdagYcMefTHXp8URui/hOmHOaqMJs8nrrVxS89cxVpET+eD9xC
1jm67K3wXFziyTqkiEwyhjHGcsFzjFUPmtMvGPV5uqz/va8AMWPpMOkjLm+GQlpN
B2GISJLunGnUpw3NGf1+E0+9czbBTV04VpobCSqe4LWoq2qAbLmfO5G2RV5+n5Xs
zJg2QlK9aYeuT2veOIs+WV7V1EVvyJcRUUBDzz35yxSivu8ll7YzxPtMzSAXm+K6
d2aD1+PxdDEleitoaeZkj9nFwbrZs39f2VqLzITahKQHAjUknoiZPEJrWP4TzrtB
IPo1MdAy0smeHTz+HPa4D8XlT/ieBsfX8bJHjJ8C9qbB1ZPXjfpmXe16jr7F4cF6
q5WM2fj/m3PW75BqdxUJ6VbHa0zQmtNgk/U910iREzOFE4SRhgQbpnI/eSejW7JK
opO1zyR6a4ZeRl4zhda+O7wglkdDiK6zSKjZGVFk0Wy1GTDKMWBiSqDWN3dWA7L2
pVJkei0ENDAJ7uPCetOupjfIcrQ5RD7M3EqgdIt1f+ixB2ei8PDse0OTQLhilv/m
ZB0Yj3SEJA8Mn8CNouh5T3Vx5Vj6H2k/UkjtXY3XSoU740fkDdBW+0c5hXKCl8ls
WyQX6pT1uwGC2y6etNoc89E/GC1Ojskssabmp/iHi80h+GNT6jxq6UaloPDz/01E
4uQtnmTgk9U5UKko9tsi41YsGJkK2cwOdTQa3axfY+0+xYaf6nV6HQT7FHiMoIDo
a+efZd8e9/xOfaGxIJOWi6ozw2bJ5d9fGX1jus/a1AsRsj0I0FgBNOEHweVvWgVG
UySBImBDG0gas398sJG4LLWIBmKH47obUIqq4ybWS0JV3tLBP+ax3SNAvdQh6r+x
HlAiqhgZdxmgZUe+Q7HAZpDLRiRIzJqYcXaR384g+ajZ0HJaLweWvn3Of+L42YwU
PCEvJqVRdE3/yHyzNKGt67PHKGQqTUWflYJMBMDwcjEeUo9dj+cT26h60PDi/Ql6
Km24WVRwegLM55OeCBtOdUZoIqudLpJYzaklpeBktGSVoMg+Y96kOIIfLEW1tnm9
2xBQxFRa+NMH/YqHX5KsvRRHaNM+03MAm2xigOZ5ks76qraJmGhunIY/VT5/0pL9
86t7zdUn7bRS5T2PWkpDRVSpqgebxs20MnU5ud8/PqYweN5z4uZz4lcdFFCwsADK
iB1PYnXjbIvJo38g1qexIOICGpLJyiFTsB6CDuD98JbTDL55EaHMnBjtiu3W/XTe
0bdENj7YpX2AhSVLHo/zU+btpnGbSOtg3Fk1DIP4+EqaaX8bS3lyXHVxdnozJ+z+
l8nDBfZxE215CuzMqEtC6/UA3ExCZgttQtButqwn0KgYEGuKmHDoz5mVRiQnmZGQ
7jO5+SH513wuL7oGLqaK3pl4CjmeCEOidXPy061miwWPbXT9Eou0vF2RuFuz3gDY
6W+WeaS2cCnXfejXJE/AntbV0khNcqSsCUTEUnbMQ9wI7G5J3HA7yvWYTAgDBATX
0wf7OiooHbnCOqL/2bS5NRHWdn5daefNOb4PSJCy9EWMdCLSdy3GwwIZYod8IjGw
VkgohkdJt4fu9Uw6kLAHhFvLCeg64FAasKlVo8UcPtltLUZxAiTEdu5S2DcQlFgH
PwHqKlvftGSgkcYs0IiUMw4qffEYFxniz4KD7GMd7zjFuV/5CSP7P/Gzw2butmAP
COg2fLddu/XtS670NBcZ2ANBnzf5t7LWXPybSnC/ZjcW5/dgFx1EB4t71AoVglxK
Ti/0Z42TTGLEWGyhm5DMTmhtT6RSRcyIMwjmlfzu04P29YAsP0g8ei7yJjmHBiu1
LU3cnGFyLM5rr9EBMBK8WWNc7qA6mwpPtK/+hEsMjNfrybZhem/5kxyqwwycQHqI
Mku/3ZiKXSVtc1MrpATbtAnKwpDuqFyo3vSzFtYyZAWSTaN9UQ8NoPP3slbV3yKv
ZqGjMGTdIfRF5fZitI6buUjxbqx6ADjkNkv/yamBDddzME9jrRBQF1n6BNqzoarF
gl8N50NCtDVnQkno3JZODNhoAn7M7xmKDuvLN3mqBet87dh4cuj49OE12t+3uU07
K4SwtIL4vB8N9tk1NftqmjdwroGNzOX/Phml2g9xxXg6t3b8T3HhqhiB+Q/x5aL4
XjCAN83UpVmKk3xk+pka91yjo22IdzT8gkYd2c6ZsmuXaIJVG/nL+2mAd/eIpLZV
DLGwq+LT4r/wse+4qnj76Ir4J2XYqZQlHRyQl03sP81L3sfxT34TVppYPsU1IdYW
5+YV6z/M9WAXbTPGlXfYCcUygJPgT2SOJR1ggs3e9DpWSlWi5EjwPvsuW895IVni
KvQRxKgeDd2kB3HIoRtQdBwY9ly2zmejOsCdSaLbvJt0VxMSihrY3FHJESiJTVh1
co/09ZKMUl0Dr5CMQJScUIgf0eY8BaqB6KNrPfMzxtaZ1vW8I7xwiY1WHdPtQRrc
h5fb5GYIXA297rzSnlF2LXi2bWMCN+XYc0Y4qg+V4iXr84MJoc2XFYWpUw7xT7m3
gT7o/xKC4JO/WbibnPauzn2mG9c2sTEdCTQhebsUxWHF93dObRjg8uDVSqtcumOW
NRS4lwYA+RJnr2c2mTF8MRZs7IosscpEFsEbTAZ6bZEYGPfrdZjZsewMvZcEGhOI
UG5EKtCUYvyYOYe5RxFyezMK5BsmNltjb3rO/7R5WDfIvpLeuhUCHWkZNWNN/vTZ
FvZHYqhkww0a0MfNwlfICyY05DBGf+xfvvcZIixvHRiPW7toq3dJJVmCjAliyFaU
99pOsI2Phoi27mffDnfW65Y6XhfM5dRRCcutOLQYHx4v7FSKbD7vOrQRSgkL32yZ
3u3tGelftRXyLWxkgmuNYmKVlZ86TdY5mNoOCR86XjJiV6mRrm3zhR1oYMkgShoa
TTr4pPdtChlAfhbn4nB9W3218VP7piJxZyOI9CCYHIT7wMW3+0qwQSBQn4srytwx
jq8O6TcTVOyscPmDxnAXGW/h4TpxIyfocOhY/x4m2TRqvTeb72pmLCwUCyQd5LKt
utZafOAM4C0dpUVo8vwqcgMKibQpKLJSg5Ktmvm2w1cHG0MI64slm9vrbKx3xIeP
UMQhzboWHhsC5cOf5RpM5xSQv1zwJwvbqFdsoyj6v2SZ2oPaBNRo73zlOjuTz9Yj
j3VJxJhPZmh9muEtvQkLCfrC3LdXSeeMjG4Kx2oIa6CuYGuXrwuXddvAddeOaKHe
fSClgBLdythGGj/yPbGECtHTsWk6xCkGp2bAdMlb0YWh6Qcfem4Sg1d4aQ77voRl
5WmbcudG1NdF5fQduCixbFsQx4nlIqrDjl/NluLBxzkGS1eoUsc0HwI+VOB7j7Ze
ZC59pCCB2OdHJHGAJqei8Ah//iOCSiNzKyhyqkQqBrTbnUEl+yQYizO/S0PTm86X
YAMA9ygg6hqnZFrJev3bIQus/XY+/v0kTEg84fg/oWX0enbU1yc3mr0rqdkC6VcA
/7kESR0z/dk4N/JpduKy37kPMcCq8thUJsH8bQM1QUWYetIffjnQctfPQxHI051g
WiCQjMrY79pnNCvlFuB7B5OZVlge4VLTge8/4ZIRK7caJOstN6Sag8iO25f5pf7/
s1I7sNPxAQ4XkVMw+JVBN/cGLnroz4A8nwDGeUtMedym86XHQi6g729bVzIWgwQZ
EYjgw948wHjVRJf1p4lm/PeDJxvgYCxCCLmw+6d1NREfzBZ2clAnicuewWpVsAPj
TzwOiiLabc7H70FCmzbmPAUNMBVAkU7QAMPah3J+ASlzLzND16vJ3rD/EV4Gdeuh
RzmAWWSTK43Hpvrg17f7BfkuuXK9xzKPNBVVyfnjlnx8aQ+YoGvmTCfCJiiUz3aH
iptfCmSTnUVllRZm2JGsxfRvl171vfwuKApfsPLcqXuEg78JItIZJMcEFdOj6pXZ
I+7WaRT2Qb5RV8rnnlpuBKSk12RPfoil2pHXknu25S7968s9x08ZAhN0bi7Bq+9J
LSygJDIj6EIpENsyMstKGtZhEKIXcJU/KEFKkcxk8YKRRgkMNr+KaB+ssKbr5zkW
dK0EAAho7oh9s78Yi6S0hYmz1JxW9fWIIGGIUQe+aRetc6rfj4C1zhJJyoB/YZwa
9n1HjRuIhuLfxATWTekynzgKgefFLMGxqwaiYPaYj5XedUE/cAt5lJrOzGSsgtsR
p2y8gjn1ZpmTvBT4Ncdl+pPt9OlN1I9JNW30+0l8gK2YhyDybjPaZpUg8+1G4TE1
fDkIYQ8IJ1HUFeroORWqHHkInvmy0lmbj8Ym7T7fZ5K6MN2Ahm8/+IU92H0pGstF
njYZP1av+JXR9FSAWraQXfOJEFlYQmbj9KSDWgJ4VexMyxwueKYSxpdF7AHqyvR7
ZUfyD0yBhor0utNKAUs255/FQtxK5CaMaFRz/xG73bnyAJgkMLrP28B98brjl4Pj
ZBaqBViRvCW6RfwFPTLjRNAurIbFln6iUJ0X4W+OympGS2RyJ16CaKcTeMsbaXbN
YuS+bP634fdW0oefm6c9cHSYd5dmPtFDUMf8rKh6JBTJEU5z9dDselvkjjPUrpTL
V6RJut/VIf1A7AKAUnK1rH5QLOeQS3r4CCZ3mHgVvZdEy+1yZ2jm0jVe0ZaMNXce
MmkahBeii+kPfGipCXhTR6mVc3w/K2UFBCY87zeHD0RmhohbMVVvY0/goDlziOSj
kF66oUSL6pQaPSkJAmBqUBr46CuT9RgBtoN8qistFw0V7/pVViSDbzI5ZTihPaCx
Lfsaw1mKd4IQ0ffBF9scIyQv9R9G/qJCCKUJH8H8bdMSAKBN050V5+b3RKemOo0g
HODXtPtdytyW07R+8jPpEAUYb9MnnBtKYbISw0T8MG+7162zeLCaisxG71CxlAHH
IudlM/6hBpYbP5a14f79k9Jn6svE1jJ77kLC/qFBoW4irSGBd5XO408OVtiHJdx6
IRyjeDYYtg5AmnJPtjEjltADDveRd6M5syDkqPGprCwtumQ0ZZf4FgHy9XZDEVKZ
C0tDphDwhPBWh0mi4bHf8RFKu3+kBk2+pfPgIWJaOYEyX/yT0y+m7U1Bp6Lzppq/
UZP7XgFmmYXqhNOmuSMV5rD/k2bi1tFOZVR/ShQRtTt9WPfNU4nTgnVRxCkhpoO/
5/+uYdLJl32K24nqjCguBY4qyPeS+ZTtLM13D7iNzOuBcO1OzX58eKvepjZKl98x
GKyHoNdzTGbG4Det4HBXemVTufmUz1+9yQrY57ArcZfbZn3rvHb/S5+Mi/vje8in
DUOjF3uame1O3TlNl4OJrEhcM0lg8LVhas3Qa6XABuhs1D1jVf0m6v0dXpPtQe9D
FVAXuFIzTSjFkomTFo9/6m1ClHyjcb2OxLbCLupMQ4p65kXKEXgJjhBqPyP9h7rc
4eve8sYJuik7vUDmUcnIGVXgXKBE2nBj08L+qFvp7wtybbjrmZMNrmw9AT7Xc+pw
rl+W5XWEzA4dCSbnALJYJbuGEOtVQYjqV3M98fR9+8B3xCr5O3F8ZQBbCbgufao3
WlPtER45wq2hsR2JSyd+cU03V1nnQ55E4+B+MzVn7+gJBH42R4WTTteKQFRaPFkc
3ByymP3unaM6u8zMW+xtxbVeeDfgosnq6FO6995ZKa6jDpy3oTglIQzwh2xDtFBs
Wc/Csg7MvElLSBvQRU26RfQK6V8Da+h+gDKn/mpkeKuq2nb6JfiK0bFKDxO+P6LO
/INz0O8AiT9ph3Sd2NXI+q6yiWLYKx69zcjwW0X84r2VwebtKJNVquF/aOhttshD
hFWzKLYqdo5F/ktWXb7dYqbM6lqyuXsU3PPhdtVgILQpthkimucK4kOWQbG+F/SX
4i46ce5prcyxBa7k9VCCU4dB6D8IBuH5ce4FEbr8efC8D3quBHgRiG9t1CkdaZa0
GQ2UEsMbQSZtU79u2AqzhtXR77EgWcyef1T+gIZ84MAb/+G0qinKIBCyZGlqIn4a
I9HsP6mee29o+IGYRkPrkMYALf5ZJ+mlvZV6MYczSdYsdeN5BHIVUrUCrgfifgV2
9m43BRFEVmG6UJAAnCtd4jdax367sjU4PdKxH8ozTIjlI5BLw/wVV7AUgY4yus1m
05B+VzSY90oAElP0TRxkEyrtiF5x4vdcVcsZp03R7Q7YU1Qog9QQvDtcZJCrvjmy
34cyPDwgUmUSONvZeu5iBuaoVFt/wRFPQZVNQqyaFymCS/RTdta/S36nr27rVwC1
W1sdGA19Yfi1HqcW7wgXygQHagUH/oQt1tAaSbA8nLdhqrrJ3GePPIbZwrzoKvHu
v2AR4ho0wBVYF1TbGp2Ey9k5cKHnrnF+jVwJ0bOgDN1kafs79vqY8cU+KPgWvWPk
fao9S1TTAIilj/MNTFmigBGHH6nb9RTnfNraGWAMYe5dTJOx9W6Cd9JWK0YTGXp7
mgKKpyrOWotYIWqw2J9cexcf2vXB4e90PquJreIR5HYXI3F/iVRNcdZFmj7UpVQl
A2d0pOBtKTRwZGLRFC48CLJ1MX9e7UpzvfavSEZw5UpFXKnG3Ks+fE31f/K9rWYX
3WA6uYAF1ADBZXh2A3CIrfx68aThP2sPoXdY3BMkv7UCtkkp/j4fN5/Kxf/6c0a9
NNQFM1NwDOeCTCxO/3hFv1QAMiodjhGO71spnWOFuxYE8AuGfFyeFMebdDAvj+9m
9/BIwG0KAeq8yn4Xj/Lcuru6aqi7iIgZ/hjX38eoSDDlbl52Z3to6yYscVGtfKwD
YUvwNusHnOv79nH7J59oQMQaQg9jAXPsRbLghAtL8kvVmAAz50P4b3wAdGbtOMhA
sIio7e+OH6MhM+ekl3Tra2DiWBnrV9MfuQsBj5qpC5361CUrlCCrgZAf8vTtiqD8
t0nNm494YujV563rQQvESMpOhbTlvLh8O+8RhGIX69xd1lkLzvNC15gX9qa85U7w
HHZc47+tL+rFiGFWWF+lbtp86hIyi+ID+tErwJBGA0f7SmrutG3jgrp/jmlfuvBe
vUYnK2jxFR6eFitQiAB5QGebmiC4hr2uTk2egaVDAo8Yt8Yl8qOYvTBLwB1LcWjw
TcODlukWfuCZDkT8xz7Q4KVCuQ6lACuI3IMJv3LO24xbztkpq4pvfriXpa8Dfkj4
MeeAMkTYhNtc5Fn/8ya8RThgt6/U5uSUC6TmEfMhf5awZy5MEZOpe85BZhJkSFqF
mHibq1jSgekojSrNO70RaLCq/fd+ssh3SWY5VDre5eQBtZ5dtN1ZDpZIUFFYWJ3V
vl4cg415Rgc+90lKjHy7e4/Ysa/kh8iJbzxF6MaaH4Y4LUGI0+0XplfvgtGRikMG
KPCNHA4O50mggZncFMopu15ctvnuSGVg8wbef7dTG+qc5WYsY9DSf60+yFg/u1zW
SE6XwjK8S35HDgWUwLtlqSOe7uq2uaMyfB8BlIZ2r0uqe0PrKgyX3klAcpiGCxSr
l2rSPUeLlo8r2FPicwi0uwzne7+/yiY0S4+lx1RIMNzNclgaznVeFizyLvqr9ezp
lVoq5y52BE3bK0BgcMD71dw/fGM2sE5MiVSzNkdQBGSmfiG4ujTm1hBZh0B3lwC4
8v2MtpJeRTK+d34mbFtkOM2bo/ZZx5idj+lfzJfyXKwWoumgp5YiKKUkHvJRwseH
+c4qtSAXWEw09bGLwOErLlP1vgWSnbIKcGl+uoZJtH8lLC0+G3Eouydr+Fe7ZVqY
+nE2J0whqXq8HPVDbu678R4PKriFWqRd1QywC/FdUUJefE9QCYX3kLNuWe0AqVDh
7Jpcj1xXTh+5nw2G0C25v5r47bYyCiGaFGkM2xNtY+ZD3zrPYdMR1qu71WSbvXkE
lOkn9/hHgWJPx9tuIPPw3MRXucTB5xyPdWyvaS8ZEvRzgRiSTaOSKG/O97pqt/64
S++2DP2Rxfs/CNGhMN/l+uVSfALC/JT2jGGULY7HD8ddzbsLTDFDSnZjLrbdbXRW
0nYMNIzIblpE2lkLF1zpW9VVH3nQfDJFdZXg6/ER4ka6gmL+EKod0cK/8nXjYhh7
aKoVY3N45o7uvYkKpdBU+XKRD4lG9PjpCcCN9Hjw2QQk7Q7qf/oK5prp3NEH6uVc
WyATfYxKn3De3YKvGTVAAM9y67+BWBf+j7mSfTiLdoiuqeBPF07ZE2hcqvXiE/qu
mJdThlMFkRP8ZKbmvzqljToum4yfKtEiV44qChuGLs8vYEMxYUpxD3RyHd2qxBqe
GyGCH1H913+e6ErQ226cNbIG873XxAq0WDJRNqgnpUANcCYDvAN8SkWJC9R3JMlJ
04+BRaRzEZb/PvUrqaBvHrk45dbuRAcwRAP7t9b178tuc9pGyyKhC5GTHzpHRhdl
K9TfXgyd70K+e4dijKg0gVNbF9iP17Hc+rC80/Ap0dEd3i+a7sU2/bTJUk2iJkIG
TFPzTfqFrj2vQhOZcn8IqssKCOEk7S0rQL10IoTYmllr8Oyo/ZJtl7WRWCkhH8Vt
XfnPnAgqdzhLdaQoVj8Qr6C0mzgmseG0MumqrUF0ipTT/xqPoYA8skDVzW6jFWir
gUDRoeLwSclnAj25FbjFl5B6tcv5ayVEOntQLtveIlOZZcsDiwnpv6vRYrlchGQW
aIymBGV1I7RYRiYPbKB8xPwVi8Nm+2Ct1M54KLmjwBiIw8eKqOr69kBWokFG+rBF
mnE8ZsHCipDtlPwaZ6HMBx8qMO1vYB0EMguDy86Ag1kPByGC2J1jRg+CSWbxOfFH
EL90oJKusXezLGd2VBfDyKFHsJT3LLVkxKd211+VE6gpE//pFxZST3KD0pEsZgIk
pSEX9lCy4+LAX6szrJZSMMjYC83/tnJnm/wwe9cuKybnVlEwOnN41WZQ1UB7hOLn
1kDlkxrsPK5uZXfELQ8nRIEGXaikRiILUyoMlMZrLB7gzzlufYhND74M9FHWa9d1
kKHSXv9L7joVsYlre37ZEV8qcVQ0Fo4Yyho0LgpCwnOAWGbG7y1lxTdGlvU9J1h8
pDfvJbOFir0tTPGcR0Zhqm9o0R6iYnYHpE8ShYERcYhQj1G0l6QoF7iIjA0mFowL
dLJkbk+xowLs/l8LGA8OWH0/c/mOfAKJOBWEWnGFrZUJqR9Wk/1E6AR3EAcq6Dhi
GgaBJg7RzJCPqEcKFQ74Q4f6qR+0YiaZeNGxMkVkb6ADi5xVzksix/ld/3Xqzsh7
eCRnXoFfCHcsUhT8QapFgblYI6xBOtuVEucj912tc1ukgjZ17YtP1XN/Q082g2z4
YP8IqKqHbANcYd34zJn+U+/eq8qn6IhUxIZlJsJ8rG9yMXrUGyNDzbYl/aG57elF
FEWKUoujbITshkYZK/5SApbDKoo1KMtzbxmae3FjvLSVa8cjYIVo06+It+sux6F5
d9FOqE2akLHAutwd5abSYU9ixyOHUSllhkh5Hw1YJXpHd2HeWsyUd3XHm/SL0hgi
biW+jbBx9Oe19uv2wjqh0Q5kL9HOmux3taAr3G7T/EVJ+kne5QE5vF8KQ7QGUpqL
RlBDEyBsS8glEOtWHrRKeTzD9Muw1Ym5gf4bVfuFcAEkqvD99UAp+X+ec58t5U7h
eKIKHzZDQVDq8REmMG8PCWP+DnG/M6nlBzfy4sgyKLnb9YGvRza+n+v0Ylt3ijLb
mVl3Q21pQ4qTspc9huTmvGb1i7zot4zjYeYMdNokXbtNKq4qBxVCh0q+98QNcJjk
YR7YeQxRxOCv/+jiSiFVMOlwMAzZ49OwqN4At0H/UJLOvyWCHooaO6qQhA1a0KGF
1X+RRW2W66+ykoSzdLIwqBeCB3ZNgmKMGhKrsZF3tDm3G9Vhy07i27x+BUqM9/zN
6RSQ1ZhVgDjNsDP6BzU8Vux3q5kdPU+Hapgiy30MQYE696YsAIjbotPHSVQ1uMX9
UqudwHraUam5CeKPahVZM6zFzrPtm+bSFj5w8ERxokHAXrHj4irHL7v6bL164Kss
dxqrYy2l+XDpeUi+GKdtVKGre4fljg5aXK7PH+iq3qWW/X0I42L3RRUNICfvkvOT
nZLvJiypLIcP2lwblXPRxIC1YtxGcMdPxQKkfZbOZndzZrMWRtcCjwbRECxltSYq
nhRrir347mhtgoKLvVYTsSL9S2dxkRxgkPDt2xZK5VkOnYfV1rRsBtIE/5/xndMa
eaxuP7g5f0rVcqnLog9oUxtzL0CNIJAClYwpdamECpAtwSN75VU9hw3m8iy7LRwE
SpJwiP6kMLz/hX5tQsmwkSqVik7jj+weI6ebqm1HN6PfaHXB26O/po1wkjmTCh2g
ibiCoSCYHZWEUAmWoooLOAYv9wsGpjQ2eEreZmOHdjaTzIrQEK3grGDuiJ8VzNmJ
/QJAdpU3qCKn2I3ER1yBGSfEKpFEx8Of+0L9hY9mRYyArfz9JZ3D9/6UO2b7l95T
aQRQI2l29TzkF0DzOTs0hx2W+n/i5EHf0Jv++/T0pTo1KqeGDhImOxJY61BYnku4
LxM/zXpIQxyIyxa5O6EG/SZ9K3eoImsIRVL+s3OVbEhC3+i0MUZ3k234cMGOpPZm
t+6uEgfIvCRd2AhXB/YXiOJh5fmiDd0/7gUKLoHXtdH2tXdr92vLodm7J1Bw4jfm
HcSog3ZJnBuYBxH7LFrc5Ih3YtPNeX0DeZLRCcmv4iZyZ16DI83OX0KOkJd6EZhG
8IRcrZJctNAErAsG9xJ/1YKPbbllPbUlsLIaTPdOf7iEUPA180TPdYVoCtnP2ucp
HvcOXbCzWKlLQjCMKLSTs52uLnUjRKwQVXUYCEBc88rmpnIFr4pIIyLBiIzPXxMi
qq26uV87HjgO5utKPJd7Rqrr6FTtjPUYXVl2Hh1BtwjQ5pG8NFwb0nYRY5M+oudb
tPN+TCJI4+TRmb0eavpRBZJg01eZsDrJ4NrMMalFpJbyE7/M9I9vf00epDPou9p0
ciRL4Hb0by76mEC3om7o0++zuaZ2Rx0V6fIq78o+SBSVYSQx7EKR8AOP4pNL3WJp
p5b2tYspVNS4AvNOHofrdCLRjkSKlnJZc6HY5fwWbxtENUl/IKmB86BxkEplaRM/
SVz2qVimkPgm+G6NgLuXapOxAyfuReTahXtaJF99xuImHdS6XqwH6xWHasy6zNti
/O5vOKjLioad5vEXq2GKNdBuNu8DMPXL9CWJMBvRv+twkqR5tRU37OlsVw+WU48L
X5gQC3XsDMIDEjUrPnrxBeCLj+8ivDgeGuSgDeSni/eL9imeNiIEYUjo7KUMGXAn
aslRnQjxO8M0sVlOwng1yf4oQMSP9ykYFeOuvUPIKhrWuIjYCueCQBSh7tt1GcmW
NaiUi5Ej4glgp6dqbhiDFGcv9XPTZl2QHdwxKpHpoT9J/0GfQZ4BxWRxXXxcFDeK
byiEZLvIpOWLknbA4fCT9wN5dN6uj+NuvBbQ3Qc2C80s+jpkk/3xPY4fSJo+o3DJ
EMLKSeLajJTeYuDPAg5eL7eLDzXa762mSWAqZCwWwsdT8QI6hwiP0926g5o/UDDC
rCUbNXlHmgIWtYPZwKNEfUhjOKsBB2X/DSkU7bTqAA+kZ2/fzJA3IBkvgrRb6O4K
mA6kWCVTIexYHUsyLFS2UlJer2gmONKeZ+CrEGnVhyZKh1vS+Wi0mnOAAqvYYBX7
2fypnjbazPkW9nIGgWqCitmuOFIFZKooWoiqwrh6fbaFq7pqjNFjeqagFyRbZH+a
T/2JUx6kpQCfgUgo6oiI/3y45KS0/4Cxn1EMUAicXK/965Bjy4RVP5s2E1qztbg4
PSE4Jl8y2LloulNQ02ZHy18pB/LRNpoh8mwoQT5Ifvc5kz/fo7rq8m9gsZoJpQ9D
3OAv3F7y2voLn99Awz06XzTDFTX41reu+fYS8m8CYCoxyrFo1oQPeMxySOzKGJsr
TQYs+aSZCLuiOmw/BB9S/mqs3HJ/MWeys1kBRZaEi1rvL4WzaNFdPRvKz1oFluTu
OC8FEZ2oNvpYsbxdsKjk1lvPt7MstwIWC+4hDZNbPYmjcyqIP+Emq71tjkuUF/d6
jXxUSDWszgRjIWp92yoz9IhRGvlveHJd/2n4RLT8XokjdjlaeF0oiFOdmTAF0ppe
08+TsPInoy1FAJbhdajSF2FcLdqEbjvi8+BgMUaR272K+zqJKLATfexzyqsXca33
aBcq+ZEOf5DoEsj5lKec25Dk+Czj4+bd1nwR6Ey6tlvfcMXTAQq8mLBVO1BG/1sX
l0c0slGrgQ1RQ3787DDt7LB5rNXN8gnfxdZyHvixE4vBZAVvRoYdsMeIhST8UTod
tlgAttpEfxGeX/WDcFaKJGJDS4uy48X/ZFswh3lOgEpvw74pDr3tcI99uzVYO9Vq
pbH/ZTi9DEB7IolBgoxpv91aFOLN+yJiu+ceDczZ2VqulLTjbvyJQN/gdh+hC+Kr
wa6jEwjudO7mhgofdhzihf0LwXtVlHxQIZNh2KvLVuYnnKIjWTqNKvHdwNIq57nz
/hLEAIJUrSsKyUlXRZwEmsjklIoYg7RNk3y/Yr6kbB4eJkWlXREXW166HaZllhCz
3j0+nT6whzyKmTHPSbTZKvlGY4t4DoKlcSj0xQVA4jkhnd0Xx6WDmRgz5kJASAgW
guip2cU4Cd1QA3VjIFBZ+8R3nIiY+Yboovf0beVreZvUHtCRS2nLwc9cMutshO5v
s+nCVIrHFeAJZ1pMyH+Ye7jvyIca9kg3Gj8LYrOFjLVaHcvzNlYQOocjpa32l1GU
yxJxtSv+Ag9nf4oKLKZSdJAgYClSDqfWmFoiTIg1zmdwJ+629yxFyvT+rTG1EQoS
sUcIeBeJT57SJtindmYlkesDVyYi1Ma/VgntETaRvPBlh7KSi/FuYrRUXF/jiPME
lac1JfTh5Qttd1ePwSPfd6kkvCSoxVmEb5krZtQw7Em9D24al06sBNI9Cx74hNmz
OglKssHxL2v81ARNrTu3VpmRFetZ5urMp7Jtk1SrLOaam/hnaVurygtp2+igAAkc
Y5OIL6HqsOYzMAt1+zDRwPdMcU1Ux39DvzzUetOqqF+T8T1KYLieayu7QKvL3fB6
J6was8Nxrmhepej2cvWQNnvaXOGNnMOu+mqlZjAdqe58YAg4rjQoCKmL5vJ6TXCR
K7qp9MQO04pVn2/juPu4j2x/pMw8Yqma6Qcs08mmph9dOi5bGQy4xPrOxBWz+Bxg
Vfz3MWYwhqru+5UGCKzn4KeRessE2p0EfSmk+EMzSQb1n4zgFrI0KjokVSG+pAWE
xb4tP4C1QPh1TirY3myA4eszDklZ9l0oMs0tL2WSx2ae3RoiUjrGv/Le7PiexaoL
njqif83IURHVYTRAr/abuagMN8PXwlEjkiuLBs3fdGG37SXmBTsu7YedpskJmlGa
yJpIbcBPUjVCRx/9n4XWDFJxManZy0haatsr0YL1u2jaDRC32COT5QW2EIdi4R8p
bnCZy6dI1mj4lyLydxIJoHRRqXNTZdPirboqjAcDvASs8gK6AP1ZEzikqyCUEy3w
q/NouI805IEofKYBmvk5oq5pSYKllZEniQNE8Dq8ZzXN5iaj06ygi1BQvKBFP9Zk
e8VmOstgRrgRA6afzNIgV+aMXyzAxKvot0jaMckp9Y6DNFfNqM5Z9c62O9rbmAh5
x8GmQGE7ivr87hPZ5t53SHzD2YxLuVgMjgvyqwvEPt4Dwn3cFfshAq7MbCM0f3EO
WVLNST16ryGQXb1ZCm23ULnbF4nQIIfpu38erAzIjdUjaoXdgd7oIK7YBmigR0Tf
OcD3X1eIt/2vBpS0Xn0gPkJpBrhKW5T9u4SKJijWL62A/1FHXCyJXH8gcXTrB2CY
3s9f1JznDOoU19rr3FRazSbfugHSEUQP8ghTKgAvnLf4Nu8Rw2WO2XVgy31lIJ0+
Oaqz05VLZHtpGZumbGOhonbWpaxCcPVSMQARlksLyYj8ZQXhqcWm9/ggQm6kmS6h
nI7+Vy7qYmk1kmxVOLipmx7WpkKfUi8JsrShDfbgzU1jjcB4rbmCd+MQG1VkSMUK
ok5+3emiJV3glredPmYxlw/0UXctUgfHQDgIAgUsxo9AJYpFLoY2BJQDFQqWfOA4
fVWebiKKxx67uno7cq9Uc/iiXJ2yLNGh+0HGpQ8ixG/g6rVAuvWKra7oCC2JJQQ3
4znjkFc1fyYPK8DleQfHJx/i65zXbErwSZy42e0Ukf/eS1Vb3shvh8LKysJU9yKx
1nqLGaSmMdGgKmFgnP4ubvN1RS9h9P+BB5n+EPb8sGjpO17PGifl93g80bKQMl1D
kbc6a8/rMQkY7IYiT5ip3SRwne2jsV6Tl83TqUCGQIKkt1rc6wDcUTfwjq+/vIP4
7tHEbgbO+A5Rhso9utRCfBni16ZDRRVeFsywR2jhc4E1RDb8+82PF2V+aarpJ5t2
l9k7SDfMVCp1aBOXkDm1GFOnzcvgoRk4lNjLrhg2hhbjyhD9AgYAp16vOj0seeX0
p/aLHSYzCxWIhmWIbrW1NDGdgGzJPpaVhJQHfTBA8GWA9geZnFF9xpyZu8zef1AE
1FXYgvtuoGg5v/td560jXVwBc4w96coQ6lWef5jm5EKi+DDu0Hnj6AXppJWmIEPZ
BCeyFRrdowrDLOD6iUuQTHmoNKXBW1YZKmfswTE5R7ccjiY5tGZS4QJstzNI8Doh
Q0kHnEmSnYJF1kNldwFvtdyy6DSBbRPUb5I8ugyT16QmfscnxR9kqFuV/gGYs/zG
5RoOgGDcuIu4R5cVft3Qfm1ypL17RHjSJu4b6O9/Nn8KIg2CH6lfm2B2ZllSxqv3
5KaH2SVyPRJhpPV49nPlXVEv1xN3r+hqgIsvrgCikFlJtPfNmSo/pEdQ08dSyI5o
/aDOyHHuwyqv38OsRz/IKFU8vbCWwoc8P9SNRhR6w4Su6Iv85DqsrhN5DZ7h5eXP
ey7JfRZNWrNfMrhOS+OC861rExFO5qrqxvkuO3t7ZpxyZ5+aCedsfmRpSKYjbzcg
FWWpQl/tdYM1HouuzHDffpYwXcJvzPNZUAMuGEigShsu6l1pfIkJFrAWKkx3/CxQ
5rXpCs2HGhAuA3LPAGWSI+1DYZQXY0y/ucD8Yo7O0E9s5OcuDwyyNizAs+9+CRWe
hwcLhC6bXRzWK7Yy8ADnFS75x84tNHH5hQERdhmt+7WsR0HjrJJd4TXoVUTMkp9t
1vdOEcy/idHiB1FFXachPmR2+c25BL9amukBQnGMefMLWoyyod9WQclB4vjo1Rsj
XX2MkJgUMFdU1NlW0+j+kLk5Vvnev7vO47hRGUkvVoJzqBxKLcVWQ+G7YExTZv80
wyVIhT1NlOVpEhE036xP+/XGJoK95r3kxI+m29G1GLzxSxojfrjSbjK7/BrxPiCN
NvQ4Q4IgcPUwCIEi/VN2o+rVA2YENhIq2OSG1kP2K9yQuEnextL/ho8L8udDIFWr
52FmZswCg1TF33DcdpUXjVo+Aj9JyY9FzaKGF5YCCUm+x4GPMhiHdg2wRMqzTxJc
QmMn/S36/frmh1fwRM6DCfrg4cy1jaXBZXQrueGZzjx+37vk9r/DqyLOL71hmEZW
LvZ+uT5wqID6qgcn7Fid8ghj3cEsuSHYcq888W5GpsrxIoNv4c5Yb4K6h+TOnudR
6ol3aJ8kIJuSGy8JjJRBviOtuSPzLawQD+fdUYrAKXF0S/d0BCzKULxSO1AjZlUs
riFb5DVaXShc7LK5SJshlGlTcxIXLtrF3JVB/H6MzdukQkw8Q0SrM+NbrAQns7fm
nHLBHyaUxNhkBeNNHJq2yz/Cx7lW85XobDxhj1NAa9b5RuypplUnQ3IXf7ENym3O
mPAiHVr0HDAI6OO+qvXsnyfrTOvy5/qj3bSfuIf5/X9lvREzDxn55utaHTqHixlz
6jp6qhBpuimqk07Hh//U9kjLeLfMrKp1E+dhn25WAYBx2sbistxLu1a4TYiEhS+f
F1zkl7PQ0jhZEIKOHXFl9+jcWdlv6c813PDWvGUlZMpV3JuLyNU91Jl3nyq/oKLv
rDuUhxN4IkWvOP71XWx17OC5oEajuztRus6rLdYSEtP0pQQ+TQNTmpac3uk8N+Jd
uAasuj9J99CLCbxCDP3LXY2kbBB3CBDWB369OVbYdgfdC3uWUcbTMp1megUm6T/7
h+xBp8odOt8PwIa+Q9UHnIYIZnbGvIYXipT89RaeCCklejrp0M6GaZMuEAngC1Fj
IrHwJn4y8C+dtzSh7zP8U1t/BfUMI6ybPonKl9d3lfUbZ2suU3hTvjZ8PTw7N3bG
BP1Qri2yChpPTYaj39RO6wxgBr1TI+gT2O+G48wgz0HQLYO7Hy/X7YnSN8dJ6t6Z
UNMVqosFs3088gaeYBXByZfiNPUeP3W4vgVlpTGUs6Jt/0MRc04rBFNN0eg6X47c
mrQBcdAXfKKbcNwMJ3MoUsDdQD6g2skomH19j5tt3h+K7Rsce7000i+h53FcI7u/
za+/SFSI0/29sex8VgmPX7cNT807B99qwONvJLYsjdgE1Np30EejxL4sx9IBlw9E
CdnlLrZQlBDKJEylPqPB2GVyXvQI1AmAD8bGMkCaCsNcX/mtA0mwVtXMvONhSeUu
f6TNpQEK2aNOyqegiaVo7qCtmXLg4tM8AdGdhr7f6g0sKyixAyKPTOEVE8KXcb/n
jIBP/3c9RNesgTckEF+pR4cS2uIpjQzUEtkTOWA9+/pQPJsnzJHUtHK0Ut2pWxg6
ZocB4RIUKkAZ8I+U/+ttwmYIhJkLhHbMzUZfHXuBH8rldoMOqniWSKyGla8Fatbt
HHGi6yA42+5L7kGk+9zKt43ZPLyiNF+46ZIhkMkw2Xb6wNvWr0DXbhVP0qPffLqF
AehJGhJkTQfgagmWzi/hxtSmlzNoS4j8FKhI2SOOd3+NkjTXu1p1pcsYVhK2zgd8
qybo/cYikeIvTg8em0xUC9FZi3vElSevbvop8rMm3bm3Xx6C+vMEouTJ2nejNlCX
sEvJwxEu9H6QjCZtl8JJjyGnx0VksGxh92rsa/XUASy4B4H78lJ9q8M9/HRlpjvH
CbmTdEYKfArjI4OShsevv1ueBDTXV/F4rQ1ukasy7kvU0N5N0OI3FelH/TCgR8+s
rMqIJVM/ay2DuYyZjQnBWjReB2qYJWbmRijm2b4ziKgWTOeAJuqTpq7OcnNYeZUu
SFFh0Y86e54hA0pmlwmUmSCorTWVVgoxR3h5gltMaY6Ad5GNdd/nc2CSyJaO8jvO
iwUT1+vQdvd98q5u8AQMMqFLfa4Vq20eyRhRnNMyyv2Y9X2F+FjT3MMI9IiSRv3E
8zY+Tp1u6yxK1EppYeFnFaSfMHXSu5kH9udMLxnqJif8bMLNe4aOxM/mpW8fHuA6
MAa1IjoACxLuyLhVBPg+f8aBnfVVXK/VO6sPPfZZ8ktxj4XODbtuv3QH6Y3/NJxq
vC4+9rzPKR7moDqxC3Dn1H+H9odqb/aVsT+ZXgCZM4m/xGVpBe1Zm0n1SXOfW43W
LStVhqVBe5tYuQmLs2ba3twvEzTPsiyalD2yHGPBc4OHz6Gwf/XFK9YlJ3AQj0gR
5dsL8jhmjgePkw5H9OUoJiVvJ98Gx/yxKFDgJnCCSlk0xh9Xtdp2OneiNNXgwnJ6
rEEIdyN0KsLy/OvDRptaapWleVW0vSFTw6qayHL2hzyBBI84J4vJsljfpRZCCmNo
nLTBKN+4ovgAV12zcOPa26LwXFH/rkjlQn2l0xSvc/JQTfO/lDERLhvRkwKQSUeT
DEScfJiu/KtOoudjwtD5mx7HE+Jud977WAAd5j5z7BE9Xmv1bQ8MedIJHb5wYjUu
e1NJJu5REJuZ1ms0Fbk9O3+MShmp9Rp5bHMtMlcpJDfHG/VP7leLtBLjizwPPzP0
5/OfHorz/PRhkiNng8GtF6vZ2fqHu98TTZsn73tIz06lXB8jXOuQFuJVoBtVRcGo
ilkIV1WDUx8ajuqg/kHe9c9UsG6NQ0f+DdC52vtJi0ERvoXDyrASfzz/S0oKHf5Z
NGQBSPAWmDVIBuBczLGATNpI8VgbGyGCS90MVsh0DmVUt90ct4I82fPo+OyeFufm
UqyXbrBwvJge7I5CFAAKbCAMunxhy2yogUz6f2+42lO2Ud0vepYcucsmfOQfcXfq
ylXhdJW/QXfni59FgDWnXd7TijUE/kMSMHcCVXvcFC56A8gmd2nhr72hnpRn6/8o
M7QetuaePjOHs+tfibw/EYVdD1/USO9/4FAIo7odSJP1WhRgQb7OU+sxyKxx0AmB
7m2z3Gjm8w28HCxzpZChm5HQh3mFtW4/g+3AgpxVYMEEOKie75YVVE8mvN04keIB
IiANvZG1NA+btSca7QmKjmAYuu1da/kz+xbX+AVB9ToQAIUXirW5ZFpEeFFFClIz
ZYOb9me7s5IFO7LXSoFZ4T8uJaG5FjJlwicCuA0mo7+XX5LfdZl2hxUWq4M5YQuc
EUI5uuEKf3qcYcI0SpX+ptW2opp1JbteCutIUHn/AYZmDsihhaZJ6+gsZAm4qygH
jfsEsZW2FK+iR7aMbt7DzJl7XT9sfBDkGGJt/LTgQXHIz7NvLjbNQit4bEGx603e
b8G2gaB/fP4e3kHalRedDiqhAPuZ7K6QfS0y5YIYEgzzgJ1L2kM2EojazedSCx9E
J1sFWiRYYcPjRCsXTuznc+U+ig3nI1z6enH7CjZVfyaevdlO4JUXa22uj7j3EeOk
6HdX7EPVYBeYUJgfSVCfRGsS0f0DaMXS0sqg5gl/55Dr1Pwv4CVw8bdCoGuxPP4T
RNmWVd0KcD+fOALmToWygQxoUi/LkBr+EfXM2TMIBa59Ua+6+qOx2h1EqwgnMxAA
59FZzVIKMZ7XeRGuAlYUdofh0u77Lad/x33hHBujeX7Izf00v8IgK6rrzlNtCyhw
VEpm8P/ReXmdqsOqprWD12gXkPbY4SBqv5PdM2WOrfPZ/mDK52Qmx3SdO7ZcVgup
H2hKclG6Mpeq9RRsviS+8rlng4CmfcSMHHzfnUW4ovQWGiiuhGnxRmpx+QkhKH46
BE1dv6kRLP9K2VpTa7Lut+jIqtCtZXSRIHjfMhrb/wy0pCjGOwt9VFCG1TzpzgQy
i/XKdMNF0iQXrw0lDp3nT+q19yxeuW67sti8kxsO0QFZcKJTZ71Q1cJ1ITurE7aG
Vwaa2g/6zwPf2GLli4E0ZhjWalf34XAYlDKzaAnsGeso8A2ccPqlPhfyrcBX4dGu
XsTSG66WvTg79tMze5GNM1j/pjFoFhyDrBUz4zUfDNqbgqrXBlFVKG57eKsUsb8O
cvjw/t+9m7l0+TRe21gzG8KXPeoqPOtp8sg0PKZI/tkalKBIqbbt1zDSciEFA8VQ
2tjuD67yiDztLTeL5Hs3PvhAlRQHyUpqpKEd3tXtRqJs+tUOQjOl1xbBOK+5nGwp
1aO3HyB3IuTK2mYWcnh3AB5UAtpayRr2fCJJHac3qZmaSEpxep6ZIq3t7RIKfKwt
MK8wDoy7B3DzvlXSplSKm4z9ZAIYEa2bi5JYKrcEt7U/x4n4/LHZ+CFKookYrA0p
VTa/YjbsT12fndUhsF/RW5zWgW3mILSAUWARhnl9cJbPnQxmM5nwCeplqbzndlTH
l906IXvYp1+sm7ZXGXxk+GumN6/SGLqiVGDExNoNBkgPaR5mS76Aa5CaS3tPQrxR
aAbxuKINbN+sdo1wQRNUsLRq0wXoj/IYPibXic4hct4bZNKHu8t4YBJ4dCfxocaf
5cNSuCcKSkLwqdjMaG/N8VZvJ48QWI0+Je655NsmiFiu7fo4Pc3sbEe2Q0FDyYRq
MabXx8Oh3De3mfATLyJ91C9ZCjf5/uL2L+nKQVw5mHLXIHR/0ywvewNDdDv8AI3O
IubfoWn7qLCqTLYqcCAqvA==
`protect END_PROTECTED
