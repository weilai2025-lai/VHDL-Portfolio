`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GXIjYSisMem2uvt9sRl5UhD33ga4JIqxlQ8F1+LK/loEy3uaFTYgKrHQfNSFlJNj
fTiy7qgPYy8OAItxUEHN0Zlw6sA/VCXO2X2W/p9afCB5Jy+p0FPEzV+C18Y1dTJ4
oagESfV80sX7fd9FWTbrMqPVkP2yuVQJFYqokt1vVqWXgji41HE1UjlGRcB8A6KW
4eby5foAzzLRNX7yDyJBxyQ1faWlSBuX19mkX+DyUvi4YHqzrZZ5PKJh7RyiG6Q5
8E9qWP2FcscnPDmEnEif5bJ8HZtCstDGVOVRPOt8bcEIP1kbZ2dBsO2g6kJ2kRlr
4JGyq5A7h/lXsR71Hs/EcLvLr2pYEsO314XrAKANEYUGLStayElkkFSfylOmI5rm
4yMFZGxYa/Aq3h1wlXIlWVT1e7mM8WNfozJjpTELaL7txHmm0ewMStEBXti3vdV0
QOKB/LdUS2sQxt5Giwo9jc9xUOovyUttY92RODpLjfF5692TZfk8HbOkywX1owRZ
7y+4MvNk116bmvK8bXuGe8JMlonFaUX7oZDUumhHy/CYsF2CWPMYK5FHsmeGX2Ji
LQiwVsFaJVOTvOXe+gniFC/rqKsPsPTUxu9mSFoH9oXAlqzKheBacp5+D8rS2HAr
7BXBOa11tAtQq1od+YXYa51OBmy/eiM/SNgOMChi5T1QF9s1ZKysgACDT1mMJQ4c
4qERA8EY5A8MXWtjvXM137i4yNKd6USSouhMsh2NSbf9c9a+CsaCqtvFoyPB/jI2
YmN7fDVO20e59mCoBk2TBMFNkEO2fZn7Dcr/OWDfEdZD5e8118gD0hviqEoEvCSd
VEVKkMI0qiU1LedNBEO7giO6C8GFLK9ccHWMAuUB5dJ6lTtWJqAnXiq9SIkSDuRn
6JaTJCQ7chmobyKQllfqLOg7X1sNMoQzWEou+wisYobGNkJ1WF028pCD9YE244t5
WcKItYn3epNYAzBl+8WvSbA5qMr5rYk63Yg3z7UqscNPpr5maZkKttHQUJfZJRga
kBhaZW2hu7SsT3xq2SOkDLzu2Xliof21vVE0r0mctqFD7o4HbK2U5Uu1DJg8Eb1D
jbA6PVOu/C3FHg/K/PxQwwybEEroVgp83J9wfoey4CO03uPZkM5rDRPC39uLPCMW
EhCsqhYeQjIwfweog480YgRoiB4Ya4NJzQ9o3cd+cSc2ZzsqkEcNw0RtK5jRZqf0
F6L/sfv3cv8dCXZjYtl4hAmiBJMeQ+dy5+gyv2dwZOyhc9xFxudqijGV9clPJZW9
oTTCTEVKqcI0h1QjMojnSPWw+5vumssCtOuOp1JLFZmpbkSjshzDDUfN731NTX6O
CdBTKAl+QhjeQVO1baf96V7XbNA8r19XhSrMgKezNn7OwOqCdLP0DnP++dGQGQbI
DPuo8+RJxBvgtAPgA/LVyWQFyj3jw3IPc0spTVvnUdYdp4RQzvGVVXtisHeQxbga
nuxIpBJ68RQJreKQ5Kazj5gbtBYM6PKe52s7HgoYVPvFV/QcD4wkTD5nd+YAzitl
Vm6mvyIuZOCosNbWc4JimaWts8h9n124Husms1itAZ0LgIW6QMOybzW5syQ9ugui
1PC+8lPBisEIYgBpjH5ti663yUjDGyY6QfY4Ilv0mOdvGd4wGMCs4pxQE4ncgdx8
AptFDe2vjsdBbEWku0pMJUY3ATk4w+iGvgBkNv96vwW0pYaS76x3kXaKihaV4Tqp
v0Ayqx3NRYtKxbTStFKKcuoGg0/F4wnD/NUpf+Ub53Azw+4J9Jp4eeYlBIxLkY5V
CByHzbyU+b5lMSxnxdto+nyR/jhUuwGJSKvHttG+8eJT1CMVwSG5nKQtz98ToMLo
k5qYvrUrtgbyXkV/Kd5eYhecU7NRKDBZN1jJCvfJZ7fSVI7Oicc2W6t2HgVDTNxH
LGPzSEATWuRA3EXc6iq2LqwR41n0EBSTmcLChPY5x2hv6m+km//wPQgoiToa0oD8
aQeieMjWTS0oV3CePO/c3g2Ou3IqL+sqGr4sEoltGubSj1bhc/H+/rFjY9f4uNHn
GuFkwDXAkyVVOYUyDjfokjR5TExP04FFGZFNWi5O0szCoPNnjocPOGGvhB3VuqJS
tSHVw0nqN64GTkQz3jc5/XAWUO8dTaddy52aU6LIZfxnQxYxiGkDwpqZKFq02mWA
MxCCO0WBXEY55MHmf20Il4QX9p094G8dugB8ngn729LtUBXWAJNX/QXKsHaBudJr
c3MbRyqwr4Y0crR68ZLJ7oO65ojq/obgxavR07cSdCsug9HiRY0Hd3uZIPbYlW8j
ZOFfgR88vsuD717XSMW/7F0SJIpSZfLgUrd7+mWpdBtaQY5x7iRJXWcNxHgAQPje
eLEVcgkJFq3GDtlcZPq/HMoCGFr1XW1bXBGa5duSHbHqEhY48wj0TBwMY1B0zSW7
+55mmsYKPgYBHrzJ/gR+hfT0ewiwQpxjBNBT/FXiYTc8vo572B7iXXhZN3LGgZAn
GH6/VVfz8ov2ZmrYSmd3TA==
`protect END_PROTECTED
