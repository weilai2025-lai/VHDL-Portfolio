`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
89NM2PJwclDcX3W00aJQQNnrvnW8CThU/WRJdiz8XdZ6ltwcpo38/zIDO6AM911k
uGne5Zr3+XxBtzjW+4HWfTiWqYHgjuXzobN1T+e0qZ+ROJOyb/6eiargCt5qa6vK
/+1x/ymCjFIeUMlZtbvuoVyv4rvWZWClXNLGXZTul0JXV8Ilfau48Kygvq7vOQip
IaFUexrY+IlXEkLoM5qnEjWK2DAM4ewmRmMgmBMZy2yJzsfC0RsyfGyE03g1lqz3
SAy6NiGJtEPOtLOSiSTfHA6nh2s7WpWOfw2Mxf5gG+DqiI9vbqhwQX5UOixID/sX
8gevlvSH141RYJw/25rKz8wMt/giS0IxIOv0WhjErKbvkpWH44Eiwn9X/kQ9atSO
1t8NLT9GnIlINB9YQomxI4S9Cl4X0/tn5rb5pIEtpDb8dsyij33j00J9g3xLAWHW
FCgIbMaNjdGazGk5EJh2c9wypnHHIBvbT/3s3ImD/u7tpL1v+qro9GIa4kw8V3bC
8yWFVGlMlLo/xvdncpwy2yywDGYGItoJrdi1vXG4JrokjBz1wNa09a0Bl32EQErU
mzJGdD3LiGwvkj/MsjTNYmHnsMMwiJSnw5zeh/1o2M0MRAp6baUydBZb+slPGosR
rZrqtN//teNvFeBuLrh/RbFfdgBgNhSw3P+W61pZo5PRL9g9/L+xGd4RbAX7cfF7
gvcu+4qEyUUYMDJMskP/NycZ9ED6TCB6wY29c8lmkuqHWf5iydt4GvzootkMs8aa
4km3T5Qy4G+bcSb0n1Vcq4ReiCsPfk9e0jqwa/2lIxfKrBpEBLSAErXtrgT4hxh/
Hx4/fD9Hx0c+bah8C+at0j69m+ow6IwcK6pTmTnZQPA=
`protect END_PROTECTED
