`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
af28cq22rpTutV48btPJ9+lWyPLgGW8gPw5njMQmd8HGYKHM0XHY8DyFN+FQ7v54
ZNNWFGmBzjEFazUwczJtb//7e+I+CCFOpl4SE+LiVdIaHfLEHpToVNJYSss8p3Mw
o53o3pD5QSbmuo47cagIrJN/zgWaey1CRPo2bfPSVS0oSJcVd7FA5CgvdfDMZ7mf
MO5Q3qApYYMIHKdMtnWV0n7qHCP5dJWNVJ8L2ZeCL635dEWT3AHXAt8tSyqgy+13
f4dQSMvYc6rKhbrM8nTEIBY6iHqRGawRvvvOP7CcKnOxqdTtN3SlbkBAyIijjMBC
aMac0EeeaEbUSfsD3HVgdvIfHQ6kckkj+hNMzS2iLhvyrBUrODGQ3qGo+1uKZ3FC
kH9leho73ADgHspSnWANoeOxY7YTpCo/nI6HtcgJDxoZ/IHijKHP1BjLtF9TjJuZ
2+Q/AVhxSbrzKQbCs9r4+3l1Fv1JTGLYjfBD50QDDCs=
`protect END_PROTECTED
