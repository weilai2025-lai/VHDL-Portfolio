`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VaEI0iAO5+D+HDZqzM6jsldLs76qYQOiRXtjKfdjXH5SLbyz3cRJaQGzFehN54xM
r1jJtVlL7Y+hJEFQ6J8Oks8k+8eMHXbZ8phW516JXJn2/AbAyOksypv65HeKgS99
HVCtB7khQb6xR0wr9Ze2UiDGDrEDADMioB2RUgJWjFnXiLe4uHLvTP1lYUpsYWl3
zMmldlU+6mseY90mVCYegkk8pCjX1C4/bRgyWv8IQcoPqRNhQ9jYipmv0nyhzflI
78LNGXggo+RaIlBshNPqFxbapllYJ3M0U72U5wa19LmpgVmAVl6DcbgUSszfq7ae
//bAudPgPUcIN4M9zbjulSytXEa6cntrgKi6Br4Dl1Ne7M6YgrMcEnbYVjcHLFGd
DTrYwvSUSdTthxfM53ZYWkOD189Q3SXQ9RfbM5X4tcqXl20d5eooBJtEfgOCib1p
Q2e1DkVhQcXfuIXQs4AxT9FPTlp/k3Cnn+WK+Ib4fRCOT7eYDoneS5r7s7kZD/QL
MzXjdZ9YN44JU7yd3gDyrf56BE8MPWYto+QaEuOWRIMCgYtzOhUty3vf9Tpj1F5E
FqKvkTprYx5KVUr6nR4SQiX816J5lWnd4RTf1/kVYnxbQuvLerOGWFth5cjgdMah
3wu065x9l2YEGCZ/WTze5INPp1TKjj57GRB/hWJGXT2H7F2c/LAsqynCaqcmzVZZ
z5/fQ41tcZzG1BWAMmU6avMiMqzTo9OuS9tuv8IHIIjP4TppKVhieF3taMgebArA
DgWFL1ZFMFqmUFbx0rB5JDSPwNLrEKMa4RXB13a//a1BxhAo8smt/7iJcbDu5LdN
MNKHLZitUTDz7IyPGMEkrMAkEXFTvLzHfuHrMfC1HEgeLwjzoqM77IBGi3Q1BEZh
OWD1hmI/90zSOcvW6ZcMMC45CmjFMRjBOo18A+pSBlX7snJwsgcpLFPpaVOj8Dvb
JzVPJe5IcuXzP8xcdSm8SZrKcha8XyrqdkR61/MzzFOvegdzoAbM4+ntZKuTCyz2
ovlwCBJIY1+XqV+HutM/6UYl2KLiCxbGr7gNkLRxZyCSM2wmmcQOcbzpZArovr/t
`protect END_PROTECTED
