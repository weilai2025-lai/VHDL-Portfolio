`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DF3UmUERN2tIergWZBl8KfTwyaUBURwo216t+wjCvCdFPYU6LcUGhOPGq84YKOiZ
QGuBLbk474bLIOa34OEMpoUo9XR8h59Rh47gxN5Jnr6AT5+BeXTmZkxnfg0cbn9n
9UB+K//z+jXYE1ANGUr7m6FiK1Czo3iNiIbUDOkx8zzTH70uWnmoJ1lSLpSUeXBp
Iizy+SxomMxPFt90KhfxBon/Ck7sTT6du/sakr0M7aJ2c6HcVYA1PngO7ZpP63C0
nFB/KUiFeSMmW5koZWIejc/D76Kd1IG6yKGOiaB9esNsLBJV1Mey7KkBgqGY2x+O
w7LHSHFpsb8bItoMM4eag+eZBrNtmSXwkK5fUg47kQqiKhtNqCUHmkh6oF73RVRJ
pU8dT8htm2RpNkw8iuiyTGFHn4iY5JZoaE0xLjrL+USi/ia9dE+USS3OyqzrWvuT
2SJxkYR7hWa5P0rsGdEhsMQKOK8pXMfucb8dxra4MWg7n0k0tP1FNMZejkez0gfI
zFhfFJI+hqYjTnjQiyDtvWhv0NGU84YclbIkJOigK3W7SXwtj4b0rZfWgew8zMs2
JdPWh6WJ/UZDbD7o352OH4c6Ilu5uO6QsMUJalZybs/qM+uuO8oiAlcPtfZ8RSEB
Ixzqz4lff3bVYuX6pA9pZj/uEy1YTKoBVKF15ix0GWbozBGsBzvqg7qJ8G9o+zJX
fDWwLNxmFdvtFWDbCa+LUUyzqBuW4OK8pAgrPaesPQbZRHpHfN97VAbpLyGuBneL
nNuC0tghNvYy40amrSNW1v4IK3QrX5xFsWnAlGi0drioRijsTqLz352xDb2vEcAH
The93ZHr9dEUMcO2DYAvHRDr8FPZJsYduuvzbVdy2cIpVejPnglJSu9yvu6M7yHH
DPyaNw4n6ojkckf5Mewn9/ADRcG6LCb7EdwL49TscEVsD6M7VzbTIlkRn5nguQaQ
nzqlapDAGjk14JIuIppxe39uxtx5S3xXYueSy8M/muqM5K6ZEdccKfoQ6byd7WDF
rS02pEBAkYdmOxDHiSPzogLXq7BZUjIkwoKfJqwxkQkecMXdkfYS1tTRorrvtaFT
HqKz9fLSV66TUVyWebwVZXL017+rw69gQvY24nR1JKdY6I8n40bPGj97WaPkZX2k
rto9VAUHavUAk4gwRCXU6Te8Z6lEeK3k3v7H2vZfRRJEhPy+52Y4OE7YHjSof+p0
e82yZvsHUCarYhVRj0Ygw6//SyLI2ZhLGoP9kWvcxW2h6mbzuYJvohwhOdBKquB1
XtNTzMzB4Uw+I7Z4s9Sdg1s+gGFFGCpwUGTAM9gll+WKoe69s6bkWEAv3FA9ovjK
l6G7yQ2289uJ2/XfDs7Hz+BSTCkevAESiGtD5wBByK+Rp4dclTccUg6vKagflWvh
9jmXgoGFUbIyFwCeYlw2jzxpuwrsLJlOmkPvlvTCV+K1uDvCCTAD0wSDHTI6hzYY
9V6Qbv0Uo0USijjL+4/pAfF9wFBhBB0nqro0Ik1EYiiwb43uEnKa5I9NlsaFlgDN
x7Fd2VBkiTd/eRN10HhEIPPrOpHH/UJj7pcg7M+ylujoaeFXQCPTIy2sO/FaYLxh
lUuDFAW58v6pku4PmrBYbY5t2UyRkfN+XohEQgOa3WZeCgY4g02CJLqeJMoqCgKn
AM7EglzddLrM3ZNIgRK0k4TyI1r74bSoVpHe7XP6LeUSQID58tlJX4X3LpEw32vl
XZ/dxEzuMXyWT7wKYh3YpHao6B77IDMdsMZqgpZ21iryCuWDmG/0l2rwu6IHD3Jq
Upvd3Psd3ZU76rxvSz30W5r9NyiNkeXAL7RvKzzPVsvjInvc9JOMYF6U8RoO3EUk
8M6k5JebDajFiN94IgHOywsKvgN/S/iTI8JQGHu7erkUnj6Ym/MbOcHQCngK1tkc
UhrSgJOS6e4M0rRVWfYgLoN8N2ARys2cwQNsU1XGH1l+TIgrfXIjR6OyZVi5I4qp
ZeeiBQQSIt9psEIUydQhxgTKrn4UpYAvNJJsOOvfjqC4wY1bJXgGOi4d684bKBYg
I5Idtl/sVFpumzXaguNhVJ+7RNdYwzUvNNiDzVJTMHVhpUMrZqqxXv2oHQH1h0OX
ZFOid7+h+/ZXPA8h5FtAae1zxm1vJnj+OyhpM8K7oixeARseJZXVgugDFrYhcEmM
TwjieNPOOOeTHq9Ej79xQygd+Hk3drJyZPFNwoPKf0EsmWeTO8CZlQxs8rOtuqzn
VKP/9Z2f2Lw2S25GsmbQFJF+CGTYgFbsu4qKQEqEJsuIJuBIYNevZD7YYfzPfA4n
viuB8mDhrJFPzIbSOFcqCwzoMwMr+3072X8tSaYvVG+RrVtlDyuO3Vywl0nYES+8
TUl6H2Qk5nss9OT8dJjtYbZaJZEEEXaELYlEbjUM/gfyDFJWN8BvW+JGVaKwUwdy
XoHLL2obhCDcOjsAqujfDgLX1rKitW0vzPidVDQf3A0BitJ+6q31qF6J6CXwiEXn
KzkAdN+6Bkj7Ilxe47aRRoAkQ0Xf3AAFCCYiPOdsCQxqaWIAtOm0y4aShN1cwqyr
hHxB7aF1DpGdV1LdliqeJQGrmlTAcYqsb+Aq8EWzaauv1dFctkaH6EFqP1XON9Zk
yRWJdpLjU0cmB+lyCSL37UemYbwTjLuWmNjMw1ILn1FPBTWPVRYsNSGRA+XTucnX
YtdnuIupihNIL8LUcH50SMCBDpJ40fIsdpZKJ/M926tbKXOESAOQqXsYPOJdehYt
rTGiitjJVqKkJJK77JoJfX6a62vG0AOYEuGxYS79bjHz8u6UNqE4oDXKfvUIEdzp
g5NWnXg51OX2A56KB5C0taco4i2Zh0GuvlqTA+sHPkZkGsW91pAQuQBMGB69SP95
+FTy2BdG1gV3CFRIwZhF9scwnuDcwDOIiz16gqAQGVxqhA4fhylJvR+opLLQeTQZ
UZOChJ2oZGPbiECzHnyyhxCmNt7dha0a4qP+HJ19ncRbX8Lul5eO8ljnK5u70bIb
Gbr2E2x195zq786tklmOqqS+28O/o5YjQxT0ScTO92YtD2wNahoEHkIF6ahdBkR3
oRuscQYci0k4Xt3aXTUSapEu3Q9eZpNP36kywxB4q4SmtsSHOwqEV7jjg+/tyXuT
lOFrTJsIBidLb8mFlYJAQ66iUWMyiSt2aolCZBWoTJg3nP+7LaYiMW9odpnHy/7p
lnPjVTiUKPAVpcE5Xuxcplf9Gi+npxddbDE1qNx8+RzFxWIiWplpNt08+64ojPop
7LsMnp7zg+GKzs56evU+ZDya0l2wg2P4D2hO0JedQUtIvfFOZZSe20z8zaTk1QNj
71tiKJEifuWGSiAVNoAIZTIaUSio1a9/M87fkf37aVsDrg99QR2YSSXtJiUqF2mg
IVg5zrvdP5nfCf1PDv0NLa5flhSWJEJwfKKtdYTXkio0yXWVOuR5i0mcIizvvK1f
4kPd89VZgOgny2ItdVmaF+WN1KRb5/zxqG3O6PV+MKkdTiNEfCjKaMN6Dzr9kAqh
LCKsQoGh/ry3dJCYvcLuB/2ImRQcLhXb6QQDbnwCkPmyq6ZepOd3ylmPhwmMSRJ3
OjVMSg13uhyCkMg/JR7SysyxXIKsWL8be7QU7Y3Lgw2kmYEpsEUgWkq7btPhQEu4
AoKZXEdlMJbEJfzzMirlpRDu+Tr7Vjgd9EaaTneCsRMOCELm8xPo9J6T7Qq066Yw
KQQhI5ruK0NDw1xKt0EzvFBWVz3cXHYSdiidskdzPx42IJHh+GZEh6xyE8PxKFuG
FqaZaJk8ICP9HOIUVRD/XsSTXZ6Ta3haTCEwhiA2ci6gNIkotqqhdr4eLjTKnGBL
pCWNNlY0maFN2bTCf/cI8uEbl1lDtPw/EnOLH38zKlIVyG/9ZzET7iz4MwkedlFC
wp1BsqlcT/jC/yACb4r8ds4wpzxTQwQdqGUv/xVnH3nz2Tnv1jbqUq1Z/RnqpbE8
3534luVTjOprrH+ZwhaEvLAsJFr9E5xQFOmDVRYDgWSZUNBF3Y+tRRGPsPSgFQff
L+JXXyygjfLOqHHM7PJ+K2KKk8uB3CmyILDSQDWF/2PLo+Fqpf8IohksI6wXqjan
gDAMlSxk9H/l4XHmeze1pOT7NeqqY/EKMLdzxZsZYgg0BrxV0MdYIwiM0g0gcwTK
dRx5oFdSq1usQFMunLB2c21vVyzznTSqxtPYvLKJ+OKvnIEh/Crl/+pl5iAu0bBB
7vOc3XIko1MfoNpxEPC3ovKuHuqEEV3opmOjfi6gQBNRfTv594WZUeOWdcXA5GeB
frg4uZC5Mlx72tQmf47WWkDXCUK+TofIMB3iTOcCCKEIGZj3MUxt70e+XkfYRKZY
UZNArI7jbX1Xub3RjsWW3wTAePekNBhf+7eYnUGUSHzFozjHRLcdfk445je2+2sX
oEDtRqYwIl9Rtfh+qEmh1BIki9bgV3GH7w0Exnss7FY1qpj4/nq2451PC2AanQcX
F36LobSYcu4D2HrxHNN7GDtkGEjl6b4KuKcvh+j8rpuoUdDs7BKyyKX/NjRVzAFT
bhNkR+sPP58XRGxQwOWAtPNNblxY0nkyOW/Lc7PDE6tB24wztewjlwweXlm8gggt
tAIRR7vhYTvGUGH085URidb2t5RSBO2z455BbFMq1cwQIRC6OzNbkODClMyM+b4p
dHCKEY0OGgRMIja3RehVCQ/40BWjxM730W49VLr3eKq4bD42iz4dzJ5lWJJ+UOU/
hQDviMASh3TUpbrwCdwetC8ibS4pvyZeyJqw/Nmfol2vxcMvJ3jJWg4SiPFAbClc
Ammr0DPAkP/V2qqUPMuj8pIyl/o3Rzy7O4bKf4HFbSRbfWZX4Ft2xDI1OwLym4lJ
5hPIj/zF7hiIY+zwOz6fZHV40UU3FJXs0Ch4WlGVY8+a/RY44r1C9ffuve534g4r
ID258sDvpF5Io51nvXbrxQImCNO0UUBovKrXczWGfbyit0MRiEaFfwnkokEMpeEO
NSXdXxPRt/LIXVqlu1YHpPO5hVbuagRcAgScKremoHACx4oKzoJvx5QzMiLUS1bB
UxL6NNZrVUrCWU1/pfoxTquQLVmy+zLIXYZ3XrGFa3mxF/2sDYjbY4lEoK8BzJL7
s0wsqNonvf+C0puaaR9A0tL18sIlxZ81UneSy/KZvqlWNH9LBUhsGzmLVOqIREMa
HfF1ijhzJxk78N+Ts55+8j/ZXImgRL9DaPV6VCZGAXY8RgaV9uyT4Y2LlC2w0A6o
VV29fLmwPAOG/EqJm1EEgQl3qVQouJl6mS2hxXqNCSFVyE/GmitFHRtF6FsSijKi
9YCk5kEkq2mWTJc8XKmhlmMhQFsUVfvXX8Gi7WC3iQbN5ofG3tjH24Zr3PcB2Y2Z
dTPLRK6q+mo7uJykGMGuNKkVtJq9G9ezhBh4AIgRXq4Y3ROktkNjAEf/GV/zIT8Q
WNhYYnXiHx2JnoKuEVlnjIyR08PMu2IEnt5H62RPAOlRs+g+q5dKk0kM+Og6JBdB
E8Y3YnowBQKrNUOj8eOF+NASN8QHYrsvnY1CNo2nSn+b4dwKWN7uI7qb+D9veLca
vGK5/AX9Tag3tsvssZSGEVmraW4c0mnra/fCWEAYn+0rrq8vqeT61fHx+2BrKX+U
hPNFRcRur2cRVYhv4I5COivUlTZNHSEBDZ/Qx7A+Gzkx4TP5Asp6LZ21sAO46Isx
Ac+HgL6BRzb7VShap0ohqtYA7Bag4JKkBcWWmYepJjVjVXTSlFpJUa4YEq5sX6wQ
ZLjIkelZkkJA3Dup6LBudz/hxUL6vNoR2ZKAnHN9HoOqGcXia1+klG0G9ZCqHl4j
faOCLvtUnWWZi2b3Vap5PI8AKW5Pq+XlHmcfa/6dDxedlzPR9ILtXxT0Tvif691Q
80I/UxJR4UVfDbq0mf3jpnKkelsGNCto84jvBtV6FkE+S8pnM8xxrHOZ2qqajAmd
mVM95AR/O8sxXoZ97Vtg/gX90sXllz2OOUaUwaUT5dNq+BujNj5Zm2soxjGvylzs
/wte0O56qGqEqSLRsoVWBXglci6b/uMOrnoXwU+MrF/EnJntNSsXdymCIeF7uFro
HnMbMObWIT3P+wDW87wTjYPnwIeAZWCrAY7gUi/RWce0D9YUa0lyTCwNbyTRkAE3
X4FotbMp574DNmJ8JZeV3k+0f+8rmTEFfHg7lLjMf9rh8qnt25PM50bSq67/axDy
bg836HRQTsGlTWa6Ghj2q3/+VCqchwYRmCiwAyrGVZsZwFuiow6LydsQaHEABi4a
F0PYJQdf7bobQobBoo8lltSFm7GCZYCziH2d0V83qGdHYvOdzNXsg3PX9eekAdzr
5NPqdxjYpzzeWUqUntyDzzF5/EXBX+DaBwqGsLBqk8aJLdPoG7H+PZ6oayxC6DHm
WIs78EHl1tuHEHfb2XXBjcQUq0qATf8o18xfDhGznJnj8KGvjRv1r7UFXbL+vfBJ
aQQuxqTVCxrNm8W28OtT9V9W8qLtPkbfcHe7i9mEJjqUG9+/YFwuqkE0DwdY5rlB
ka0JmQl0U8UfErsl5DhwDopc8q1PizGApO4LhV+5UwmaJXXL0HlMKgdiKUj4gg3O
HOCfl10BfB34sN2xGK895lenBFTpovQMbDRFWFpWu7gQnV+9pCf7N63b/lokdTJ4
fuFaWmV8fVFe0O8mqr80aTvf21PEErBf0cRMfIz/xlpVbjlz3mYywPuJN1txPr/S
hbjJyT0BHI2CkbU0yKoctOMG+63cC3NNkW8JB/Vnzqg5rPMnCtJEV/wvEMP7GbPy
PSy9FsGpEiydRUnpWNliyxcxxVOm4rCKFfIABNT3Q2eFPes/7+DP9lShXcG1HYaE
WX49rPwNcXQDNeK1Icwb+yhQZBj6GwtAEhdB3j1cBmCr6rCmDodfbamPHtCHNo1Q
ikV78arvhRTwD3SsQRhOkpuy/Fj8XNfaEfsSuTD2mvk2FJYG3BGlVICOKRol78u2
v8eRu4n7cZBb5cjhxbM/C/WANw9tq3dtc/LsKdl+Bb3yzPyBmUVTWHkdXp+HWap4
uvWnepKGMmv6EFkluL+wEIe/ThJZJKhdQCEQlmrICvUH+gmi20VIAGLkkZsJ7d9k
qXcbOGNRdyi4LcmyDn6FH0rmjqFauvKU9v28FJdhCXhu0U6ZG+u1IHB+MF4vWEn9
D3gdGljDnFoiIcAuMa8qTWCFcDAiF5PR8SQBN4z62NajjPsTS4la7I5gUExbaCPm
bKexMOK9JZDqFuWLzmYKBwRuDjNtvzykMjeJUh3mKBJE90C8jI9Arj+LnfucttOI
sPb8k2oFdbadJVby/wzltpjQAwI6pO85KxHaOsQJrRQRt+P9NZbiQQNmVRMJkGwi
LI/Smgvm+/uTUxVm6Z1mk/didy898K5jW51+FdgYMZcsaP9aQLqSpvK/r6aac+p5
J8ZaTxHmrzhPzKGwi6d07SUVu4a6A7Ux5JvMT5vYe150lYh7v8CXTvdJeEh1ZQJP
NDqTMenVwcpEOA+M9zOzINCR3DNHsYpQ23e+PhOOWwI2Mxk5ww12ba2LDWZCFw0s
xODLZtLPjclbVjbeG3/EW2qH2W7wXFgzZ0t4H5SEkSeD4ztKUj63QFAL9Zw4qYUl
im309rDMbXhkFp6p7XgASm/ZRUAZG5Bl0XMHH5rzBcsFvXgXeVG507w5RQ5ouB5r
Fj6S87EpNdYjYPXEQwt87NyJMmA/g3LxTgJ7SIVg+ZESh6BJgP6sUTuoqFPfhRGc
BE+JWpimhxCG30RWCrT+DR3hnojNRvlBis6j9vZDXVQFHgxKn4dqV3eyPL9JjskR
fb9hRgyRAnT0DOO3Sy/GoSsUD3KUVPTWf9GDFDp3rKLetPJcs+9grsFX0DSvjYje
DM+BdkrbdZRuoybW//hUTBz6XIMiLkcAwMBeKkOjfuJLTeI9i51R1K4gpe2JcXwj
nOFhjl/fPYVrc1F1/b97nndTXwv6aoRsu8qJAmJYN9izz8H8R3zIfmSdGN7pFMVZ
JBRpJaqVz1zOzFF27f1zEzMKRlpIt/Ko6EzqCTB4C5QjVim3GXCqJL2yEGmE2PtI
gy3bkpwLsou/20IH7Cmng341oDVjc+74UI59C6yjMp7LFo6Ha67MBPrrpyDUbypq
6HrT09dzv/27s9J/esZgK7QtENua4WdCA/o57cRnr8eatSfSdo/ChCV9ZiYXph3x
4kCUPZigSdIHp3Ulda7AcTIqI/eNlgbhio2ERFYn11tCO1ykwWmbp2XZdkn9fqhj
nS1C+zd2sC/439ikm6xNoPqu8yTgpvN3s8VLZComzmrVm2GKbSq2zrWcMcuEg0sj
caAJp851KgdYG5ug5DYwWQVn8AyZb31JPnZihbmjDJQYwIOwXMTlnrr0m5pYZ464
rJAkCPOTKOGDlTULBQ18kqGFCVuUyjHPDyVcYP1kglvzAKuf2xy52SOBfamcaJ8U
hLb7d3xzEO68PkuPJtmH5LlL9208ak8jqJxKbPz861eC03cEtVBCc+KuQjhjWyyc
WFSnVzHIiyHGTel7w7HJKpbIQcgKOX6KM3p0xoQAuG/wjwzUVpU7zfmQVukIKM/i
P5brAx2T63t0Jk+W9nI6EXmi2HGZJph/4GpAPK3sVnsj2FAthDShr/GfgAwi5mGw
h9wk+qf0YxWfR1yJa6YAe0uufqkI6vQElgVoukR0nZK+XHijcoLXgYeyn7mFu8sc
k1RfG4ga2YKElg8X+WkIMhx1tENpGEV6mMsa87bps9UwnJKL5BWbbj+JVV8pBe+R
gpcI8Kj/4F1Zj3AMksesON4FRSpcghBztv3Iy1EnyB5SdSkGWl3X7/Pbmxek7wSm
9/utP4fCo/9XFDjgJU8Sfn+WpjoEzovjBhUQH8qAQ/Y9NtzrgnkEcdUpELl1xODA
orbuL0ZwGO4+2saSYpJt9fK17Gg3hiGvv94uRXzoZekUdK5A171LtgdWLy8bcTB3
Yn8td3sZ5fLGYnMi/Y92mXSk3wNwAPYmD84LLErjTwmbVE33iXqp0Cu6lDDuu6+m
cIn97Ssxlb/S5LMGOMLmG2F9upqtpKWio0oSusD/Q7z6jipAiDf4DInMixbSGdVD
MNYoGB4O7hoNrDbkDzkEfOREKFAWIgSDWeYIfi4d2OTKy1SlrlPRL9ggYhL5o1oN
zdf/HyzBrmwG4ZWd46VsQbJTQI8v2Dy+LIinKfCRf5TwKdVKRHKILurOtnuUunGk
h5owbkir0VbO18zbI2Zc3bFSFm04RLdkNCpsTYNltEs1uSjJGSOqiNM6Nt/WNjhA
9CibDd22zacnq8X0erL7o+WKpTvTHw7HKYnEqtKeo1YNQP0+BFhPpNCkUbkoQL9e
dcgo+cM7Qv5K6EhMvaYUj5ZpxK0d1YLvRM2IY/tPxRhoJOew5s0JnDOqq6wEazWQ
57UPZR92MXyJPdzrUD53Mb5uTZFD+7eEubdAOWkc1w2DX8t7SuZuhqBQpO/EIwSP
eOAQFMn64oLkrcy2sakOW0kjB5Q/SWVtXVnfXcbO1JALctfRl7Fz0X7UQ4AaFzw9
fDXSWLBg7WUI1sFIRBYq24zvv91P8aGnoiFgamuP9RBCu++E1eqWQzlueEtqPWw3
2XKMkl1BuAToQTKhRhuRvUTv2o6QMQ+4zkU0EkUXQAFseZpjkCRJm4J0KPOUFtBr
fPan8LKvoOoS8kbwZpp9mWsZVtbr3tHVbkkQyHav75VmA9Kc97lZX1dzyvKePV8Y
UtzoZXRWLSenstS26rhvVT7JluPDAmkJ5UAEra2ai4wzTqfaX39ml9lNFi6Ph3FZ
X7DtwCNWipjC6E1xO1wMC1xp3S2jr2Dao2v7Li8z7/+q8nNwiiA1a5OxnO3z2+2P
I/+pvU5eAj6kIukt4G0jLY6fMwyY5f5p2Unfm9ZOCGT2jP49d86vpQRpxeYxrFht
QvVOZ+r4laWwEt8nLFFbEae1vLYG7TY8z8jJm2H+VyFJwvkte7icFtIiHhDCO429
Rg7BRGKxfdQeJ7H2N2tI1/ph5bouWROMgubHbycxDBI1lLZEcb8xktitZbufgw3Z
zh50st6KG27zakzhhKnqyr8hLZLAa/h4HEXCr4rbb/BaCZ7XLmB2ejE1XJqH0rqE
++LuCgjyGRPB9ktFQlyY6jlBC9uVZknQP/MjeJvj9aXpIhnwg2BE/JIzdXYF1/Rm
PAMFZwUszhqK5ZXuz3c/wyEzrILrv1qbx6lIhmOKn9VVo8wq7CF79Xp4H/BmBKp0
0AicLbxNSLuNintatBy94hUbSSNF10QZXybcw6iqqENVpet/OFC6rSBKAwu33r0G
Rwx7Lo5BN9ajZUALiP7K4H43cLuHlZPZfXSOMPD33gIR7JqoEFt/VJmqgoVw2XB2
/hYYOlt3Fxk/K+SpBv18+xRXxMFRJmHVPnJbaglUlX+N/PXHlZVZQnu8WAmhMB/w
7beVBe1OkI0bIwkOFb5KyDJLwto6s+DNsXSqfGw46BJguXoQcZgeLMWLx+cLEeqH
s8hyIIgHZFmHQt0oWltC48ro7vQ4KwfAjZ24KjGTma7Htxab+z5yG6qcvlZ1xKZg
C7RFUF0Es7wKzGp8mKyzud1PP/HAQIWjUozMEWwlrl7PmsAsZDhvF6iz/oUSD4d0
sCW7Bx8697EF/WpOzeJ69ugD3P/NNhT/gG0yehmt1uo61yhQv+RjwT7dAZM/MaEQ
7ExY5mtvZQ5bWKI3T/yaVMiwerV/NCNfebNRV+QoYi8sxKkFm4u/KuaXYZ8xY4eM
r9Jyc+bO6PbB809Ac8i6fr8Zx/E4VZgxk4y/9M6zSat433CzdnioH2oj1vuagXre
kHny/vCVbs6UihnnBE5nbY2+09yAyU4v3ieE48PU2Lwe/pTEejxJzwczY4Rjk3iu
Wg+f2IokSZW8tlf5rkzmjhjfJBDQyGJ/JbU+jaffQlwLEzP1KnLTp6VuEeb8OAtU
iIGEwew5390ZFwpLdmEB41VO0Y0ANxPLPcsnFzFWT+TFK95pjWWVaxlRSnERiskW
qW580qNoO6Ct5UOeJQ/lT/O+dMn31ykjuH0zFukmgy7lqaFC/6TsGELO8ZyT6vLy
Ylh9wAeIXcQhOneqOJGlS8BQEDVho8oi96sEFtAxGNSjB9Z0TVTbNWte+Gw/2imP
VRVUCNZBUma+6eNt3zAQVBGj4/qaJIfBHn9dLMP/HBbvbX10qWHJXd7ZNPsVlW/2
fSJPwdUTRgUw78qhHPSCRBLxBq+cYh92fvWWjUw9i01Vd7IA/giwgTJLc8J3Wj2y
Wnl6YpnTXUuoO1U1LL4Ov5RFK76btxkbAzS8dK/SNA0fww80vfmWK5KVnUOytGCf
RnDQYpUT6uhHHYzpjNviP81VfyYnPWqUnpnGy8iVDIitbUpl99tRlD3Bqr+jjXYc
MGPG+3lzl66zPK6CcwWpvPEo5+aSDWcvqaXWif6uko37jUnwJr236FtOFUOQFDkT
zCoDG3NbuBZudSa8Bz3wjc3MxyHLpVyO6L3M6CjnS+3Pf5HgUxgFWVmZQctHpNA9
nCEBxCUg188AF2VLOg1ekQq9LXiCgMjsfF15EMVSlBJqVp+55kHrgMMI5+bvAJb8
6y74z+52jYGAbQnfB1hmvh1Zn8cANcRhESdrHAC7qO9xcnnGyprMwEDPcpnDkN/M
husp6CMSw+4Ov5hAS/rVJWpczVZNwc+tmcfVHuQzAXyCK/pcDxA//4R51R2mchFk
4yF+wsZs+pddKvWKKsUfWNIqrIDZSXdXT/3WsRXldlnZxHV2jTsRZvzydzuLlT+T
dEfUL2iBiwO+3Epr/MGMv8JM8eA/itWHbpvDW6WYVxd7MiOXCEBMoel8f3qft40p
Jlp8KbU0p/5qTUuubqcoLtt/pbT2A4nnW8Brdk9+0BkY/hOfe5j1SNjDFkXxn9rw
mMSbkHHhUEJyj+lWLqNH69DcaZdKcmfFG2JUSE1CzVy/4bKBLb1EH6nVp/g1eLMC
XfLHixBKJMndkSvlRw7pONpd5X4Dyk/ksxNq1BDfbKhh3FfBhvnbgfJ+qy0oa6zr
yKEB2pyhDIAmMD6ey1D5x8UaA63Jy+j0JWmHbjezUFINJOGty+wro9yQAM3UmXB9
oBtnocHE1FSMRy6YD0Sicfpqmt9EzRzp2aW+oYbXulRc3eZt6V5eQllrMe9jDRpx
bjQEZBdiO5yjU7KOhEaHdHE94pvnqEwdt2A0LcpA4j7jbpSWWaK4M6LkCwDXspjg
4T0ZmmrW0o1hadMmWpWjbJAs70qoInj97w7GIncGQTCOXY7lrWB0Me4egkb+Li0g
p2huJotrQyN9nH5xvJYCXZ8J/vUcIPewFZqk8DP49aCuOQ/4O8zBWkfikD7cuhwK
x/QZabCFrTB3KTmZBYKpPzWwxd2Q+DnX12trrUGBpyqls9StO2caYiDqz+tJzjqA
ypQIslpPQ7OR+Bj9/7Puee3yXneQlskVHQAzol7N0y4FtaJ4Ml+S2Vhp3P9SSy84
cubNkhweZPaBm2cDpVsynYxezAgJvt0VSlLpdOFR2QGzFOIXX8NjcgixGhigS3Uy
ItWAXlXxGSgUWsWBQjLsJBN55FFSr3JzEJ0Jk+/4UPsLLw0Xo5lpzkmsAd0FRh6s
DaiA8ouF9f3QjUImjloth0bn9loY9O5615h9dKCZTqron4dZ4dT9mAtB06DGWJDa
dH0zsEu4iI1V8VsXSQ1WZFGeacBsjLOqq12Y0FgU6/qRqlAvxQaz/P18mP83lSUY
tV4Z5YFH3Qnp4Er25saxW0LWW8pBxOpnCPR8ghm8FUsnsn+HGwl+fQVYv458yUHu
QwG7zffr4pgir0M2lWYe2hSbhYFGgCIukc5d/Z00zn22IFz02wiAH47pJSh01U/P
M/Ns3T0OGTtQ06iDYHPio3xOl5nFuMIQfpT/GkPpWsjDS7fTFR9UczMCM30ffH2y
gIkXQWRjmBFWfW5Woo+lfv3/9KefeOEB20XSMHw6dXBaaKZ3alCmTlu+srg5VaPQ
tqvKFRTe1jD8lDuKAWq+v+8jIXFVV5DPA3qHET4gxiiYMozHcxk8lIwT4Q9ORatY
dIho+3RBrbQd0TM0tUEFn0fD0wgj8VrU/wXzj1xMonifRXUFj+/anVubosZu3wZ9
ntmvXpraAO/ltc8ewOfIQj/FKUpFa3/GagNlf/3zUl/QmTHFGxbo3xoO517MW+he
Y53PaVDydAkTlYKK73wX1bHPHxh06fRT+cRPd1UXMBeU+PGSrqL0INoA9ScWbV/5
yNHba+ReCFWsZJ5gcu7Ad0dSQBZK9rsf36tsLsazG3qByzj9nQbdkBHuPONkiSa/
YHEcP9vRIlJoXB5wItUO7uB5H9CrSp7OY5QUSQ7R/OWlKigxgFrJdL0jGUjpLwOA
t84mpSulOoFC1BK1xCHKGkz6lfIuKYI6jUHmss4VuTp7ZuS7L1q9yQXedYvcAwb9
EYSpX7to9enNY7z/ubLfB3t60YHjjByWxelJQ+2oawEsrh+tjSAG+yLs1LthGExF
4oYIpkVfuHKBhBAdzbUVfijbrp2kYOcWU/yKRVqBIUV+BkxqT81x5wV0nEb9fbKd
AIl1UjkKmDOc3gTVhCUQ8aeexVVf6+iedCh3f9czJeKImfolDyi71mpv93um3Dhs
rUJ0srEwFtnqvYFTJpf45r66Jh60c/nK4MVO7is8K1ONj+cB2K2ITYJoa5ATCvFc
j5TsQ6OcWtY3cfClXSzabbmyOwIfqQ8fE8dZCqTPxg9/l8JH3GLK3qg7Jj5z0i0X
DBY7H2VdaIAx0/R9OVTThzTS5jQ0KCIcAR9L7TQkfyjgCvFqEp/T1rn1FQZGQXD8
+F7IQQnFPLY4TbaY6knSgxNxKlweKR9T7jEm1+g0F7saKdvf6rPCTuTGjwIajj0l
dsO5utYWYQJ9AVyk+/SW8ASNyOvK9wMv93JV7GspGEGJD6qrYgPtiojebM+avqzW
jnO2rdQQBZF8IEQ4gZqhd31sMOLNTdYYDmM9zO44AGvfI5iaQdRQ2ydsd+bpUqtJ
yZfeV5SMrmhhnFA2kiBvwM3aFZyvNCeED+ziWUjm7K9qnbBCDBsCye6iDGh9OuN0
UuBLSf+B1OCrB0wu65uQO/Wmxh3sTacnh3VXD3QeqbpxM0RYfIT3WNxvTAkfYfmX
btMKMUkg6bgLMrjU1hnj488ghpHYRqlI1bO9nHhB5PV6G4G7BslFgwl8WnxU8yIw
GN2d7pP6WDwS7958q/qk37bItpp1jgIjTaLhibyUFlDlwuldyBVgYm258lUHaxyF
9zGjPZgz+jnIKoO+XShh/LW2k0Yo9mPm+MsmYNxawNzRqQ6/xDthzjsywBesLzfl
qWSiRMt0MOnoSZgwGquRRFCfkCRFaFaHiAruQLzSvwkkdqX9vDbf9XaPSUcDBCIV
oWJeL/0ynYeX2mgEGLwBN52osZosYDr3VuT6KeVHjzuzoOns6rFizins/eG3gPhY
fBgGgBh+d7/7SiqR6RyC+ROUAEEsHnRx07UEdWSdrZaQSqm2se5/dIKnfDZ264+T
0cfPdUVi7A3y6RvM4XJiRdBtcAsN98S/sVUaodWaXNh96HFPlZLrT+09OQC5EIAU
AF1L1ufFc97Rn4zngcVCEMpGLRGE5+1ZhdAKeUZdhZx8fOEFSEAougqDHAh3nhYr
Nd3PeUJ/ToFnJFo6SOZtbr1ewe3Fqsmn1d3PaWmo7WPyy15NueRy8ZkqJI21X31s
5eJ+AFVxqH/13aNhLj0Ai87h/S7iXELHycS8grNu9QMMN14NUiRwCJaiaTm8lIeh
CQY/ZjwJV0M4LLQG9a4+OC2/Z7wYGt+LX9ihru5flHfN12zmz5j0MchMrLBCh4sx
SefBwcPD8WmWhwJXfM6/B9XK5xmCl9dBTThuAljdFWSPYhsCRhjBPXPDX/OMbgWq
m4/Thuaz/S6lxA1AX7+1FwAKrpjwCpe+nF4KAj7nG6/nYWX1n60NaelIBp5dE2FE
Zj7KDrj+QCY8co0klhubjwhvrA0tvlMsUmQDRmVJMkT9P7xgV+8JvLkC4tYYMYib
WuH+gc85HvMBulc8A2SAiQuw2oRf/QssdApq9qjzeLqbG1SSSCRMkCpfgLzkd9IR
ylfjDgwZe32ar1dmGfkxhquku6EBcLkExupmmmiOZe4nu+GorPEv4gkm69rayqnI
PI4AuKNQ0r6w+S8xI1pJew7QwXpzWEY8ueivn9eR5Hf6bg9wG0qg3z8acqvnT/r6
UuUG+/J0wiimmPV0WmJ3e1V8YUFe4sFbSVtGH6nazXjzdh1VOv202jxiunxS/EGl
N84BGHY9viRwpugvLvMPpxN9lfnwbyC9so4ZOn1eLvCk8r7y4mROWL0DR1f1UdVW
ZHFgMMnL0XDpqxj0du9fQAf+ZmlKZUOyvT6BksGzjguZqrcMp+ryZRVaUHiNDsOg
AaWG2POpFGSEcElypRoAO9qyoad523i55IMsDkyWHUJZ9xWEZJFI1X51wHH75jJt
CAVEFMaUTkaSgAMP3KSreSjbhot8IY7mVh6crsQuttDzkjXVNPlAiNarjzRRS6Xq
1kNFB1HAMQt/QArG2uSkgwMya2mfpi3LltL4RSLtqy38xgQWSgLdh4w/rW5IsAFV
3oqY8+Z09cdFMLEuXYWwwLjSubAVBMcL1mLAOMm/Z7Y4PiwEU885NrUphJeamJFI
ymNOfI0L/5cF8rx3f+fzW8zuU87bcqccQ1sv6ZhJmsFfQ9qoOTYmDpxoCtDwi/sr
cZ29fvMfhB0ZrwwFuDJCs34Ekj5wbJQTY1QeyrClhUk+2LWV35SMOqVwM+eDdjMU
vcGObym3AOFwyXdE+HbUzdhEQ/5Td3MR3yKnnelYDoeJFks5YkQ2JYjFrWXCLFGb
nY8HgtuJpqX0h0tBTbL8HlzZ7dQo7qjLoGBy1P5u7NRujV4UzEmXbz39Id0Srn7Q
Cn1HTEijcznDZv13jjijL2Yw0WQHBeFQ7wEL2ZiYqE3+Gdq649N4mFrzT7ZXzpBW
h5JndARsYgfx068dTawn+znaQ6kEtaIR+YbeCARS7zZx9REbhhhVbbIlHmEWRMbV
isyeJmMzYnEpYdekPbwH5tOwl0R2NDa5SLMGtbPjPuCQ6bvZ1+3a+kx7ed6RoI67
/Dah2z3woC/QH22KTdTplsQXyD6UOeDnZTrTSw3JEzeC5ZA1RcnCDZA0IMe105Kz
RuN9UlWybeWVrH2e6ok/UX6BDV0f01p3WRoXLaZxLd+A+6jVh1j2DLsDNCl2ngEO
4kOj0wn5sS0F5Dwt9RPWNIwUPVKWJ3tNGqj/tRMfCp8XqHBtJav/lU0p3WizJZbc
GiDvv2hItne5Fd/9D0Cfuz3iHNbt1HA3iHYWOoQhVbtSEofFlo3Lnre8VA8QCH6E
xSCjO/zdJP8u+HtGLB+uqIWE+caf1B2jtrBQChH61i0SFpavyGUqiDxirTOli2Tt
HPjaIRUFcT/Z2me2gswBv6qpIbEMvxKlk1OhTR/avF4ZYAyVxooL5ceNKqtyUtdH
YAT11+bEsns5Z1mSRvsdmrbozeDRoM6lKeWVGAU9j95gwGs1lsRMYxozc6GbvYjr
B8iPv0tmC5jMeR9R/jqupTNnKfYWATiYXeQvgNwWmOYKRGRyRSJR9vLdPyb8fhpd
uOzkp/RDXOXAgG9m/+UHDN28gpRp1rdVQtQci3yjF4LyPQGrQbEf2MxLtbHDTqKR
W9E60061If6n08n5u6iXR8u7WMyybyZorl8z03joX3dBT9k0S2gsgR22Di9DXEmr
728mqJw0jHnCMXNXA5uoFxFD1nLsXsnao7cd3yHukfQ7tYkixh4tbBJiQCqY3kwy
M7foOJU1kOVYCo40zPB4VGlZlNZRDMQa937DClrH+iIO41xOwo5cuktCvegagAq1
kTtzXeuMfrEtrWVshJDzbiCqstK8roPEEso0YVAYwVgPzpdR1fM36K/eq6ltU5s7
P0Bd//Qgq7Do/f2meaejyOg+ht6uQKxbd5pcZpRqd+34Pi8e57buz+vrpU0IueIK
CTzLKgaM/QFTOvuJ8LjIQIuzwuU/x5ajiUKuvqHmGYS57P2STQNswumod5W+soyk
FKKUf0fW6z8OFsZtH1urr9k/Y9mlZ276ygNA3IkjjM9PVRiDhI4D3WvFoyd3GFrh
IPLCDBmZb6de9MQCLRl30e21KXr4CaQ5eDIphK3UTWEQW4rB5P+ZzecItm7KfE8a
xfPma2MG97eXuVXhY/lIECMd6u6KCDKsMYYEz7jPTBAGiz3VXYuY1hSJNMnhsNxW
Fs3LxJhj4gPxflaG5qtRw4tIsv2u3hSm9VjKHb0v4DYUDJsYNuFSQNR4MINZvNQB
r6+zC/KgY9DAXqHq5hCBZNyCfCpCe4piBlELnvmrOI2BIdPWnwPg7/7BQDwjjXGk
t42k/UUZu7VkUy6efzkQifDzCiuJkecGzsBrnIvrSv+YiOBNg3j5xWal0bmAxmKK
TS6t9VwOA9rhFjnWmaQqo1bN+h18/6ZNuyY/pFVAWgrGbmR4IXd6M0JSX96cCNk4
FO27Te1a47vslHrC99mSt4GVDKM1zKYYrQP4Gkjle8KIL+v2TRV8gno7n+XFbOsb
fV/JWfGlNxFm+7ObdrWXP0RJx1I7jUEShaztyBrQt/OLJV/ZeeSWKZiq8sCw5tx2
K4Fxpdm/709SdyWCbbJPjkXenLn2KvP6M8ZGFWeoIupWJUSUqujnSWGOhvNELGqR
Ozb3e0e7YAtritMVO+VjWBI4vBVFiPwf4K4G2mcR2fZXPgaPBBrW+Oa0KywKpahr
XxjQKm9er/i0K1HUI6sU5BzVIRHxfFH8avgm/tzCw9b6m17EHYiAi+cqQptyb0Sw
ILS0IBBA9KXiJXX+58yFO4c1hbk1L4mmd02ihxEVozYReBafrQQL3nHRchcnv2Yb
DANtBdf0iDst+vmW81qBR22vjpMDCMpAS/oxwxq1wsCnk6oGHfa4uMsNxn+ydu2y
oT9QoO90Pwwbk9jqD5FzhlRdt3ySAhBYfhr6ulx/ZhFUkJr3F1MGR6nA+aEugU2c
N30PqJqii7YdBJmySIpo+e3Ais3ZX9/i1XMSYVN19rEpneWN4pLAnNOORmtzpoQX
cmlvgZL3DUx95UboyH8D4ZjLdhj7/eyZtkdnxEw48O3ls6oI6MEAlHDgjNpPxslP
RaexhuVlxx88mIfRuG/DjD4O6EwBYy3T0vR+RObVGa803nnLD9+kRFFXVg1Sm5rR
aY4b/A/qk5mA4vvg9AeSl1L6QpQxxktQIN8WYvBsUNV8S46xDkWdP0MAPrUvE3GQ
M6ea5dx79Dpd0c1PjzS6g1fq5qqCf5AiWohDIRE9BgNlg+2Sc9pwmZLenAHwP+qH
2nRAx9lJYTmNjnDFtoG8B2kKjbYtE1aboIG47I8H/EYbTxrgnPfo/Zt4yX5kcR4Z
xUM/Lhqpz1Wflp7uDfsY8FA6U0KTH/Fl3ofcikWoD0Gr6YRTg5hl6IBxLmkalqKu
u2NcBx0hk9P8YucDLKDXQLoIEA7WAILZluIumV9jsE75dy/XKC9v4XlYp1+1IOIt
g8RJuwW0HvA6vUrwrBIjI4pXe+vmD0K9BhvpP21AZt+p+en/OvYLirNP4RtEocJS
KiYWpHiqYjJpAG69x1JHu4w2L/36eXBj6IItxLCDIrZFrtsHf9ezSR0V0fh3cqy0
at7SNfQKxOSusy/t23tv2Wn5ugzHFDDO8TMQev0TyXq/vpxsDjDSmqhj+KN/rhQC
JUINOSsi1fkXHfgGYD6rInS1Mll/Jgf4xOBQHrUwCXH5t8ID+sBEEAr4ujLLXUfJ
+fuRqDzF9BsUMAOQMx6NONMDYsWO1NwSRITf+dVSpjRIoAtaGvq3g6SPKOshoVq2
560roYJQLsqrAhdsHXejwENhOjXOuIPBo/IiL+Tqc08tiGQjPr+/yAh1Payk02L9
G74cnVP2EBbbUSWYp3TaFa+8VDrLb5a6rgkhE+mms6/g1mCXdz9XxrrUwDzT/cE6
/Yerd7kyh/THsAvO2bXT0z0Qcykeib+wph3hFzgRJ3D1pTeIuERkbBV+PShYAkvH
2Hq3OdxhhOzhh+yl4tCbTxyVEKP7yg7pYKtld8Ko/LGrcNXoB+7908rus1jWFc7L
K09Kk4nxvmBR5UzUmkYIXZ+tLoObhM4rdrJv8nezgV4by9AJxmQt/BEN1N1cq5Ng
IUkpHWo8JuQQaSan8UE2HRQIcc6aWNx2nwIH+K6Ct3XyCpfYfgr+pgjnn1nOsDmD
bx3SYCjc4q+TQunrTAm2+Nx//yITzfQpT0ghcYebeS0gLge/R5NeU+OiRk1is+s6
01GPaSSIcZa/3GJTIGSNIwl9/WBB3+Tt5O19nkpK49g7n7rgORcjNNibVrhQ30TF
dkcPVu1U/Dx3MMwEmvH2FZkAhaUckRyCWLMys4cT7pztJpvYLCjs7KBYqXXW8KaV
smvAjbHlXTu3dEXQA1zjrYTmRR29HarJBIqs7ZKn1XjK+ipQLd7VVvIFzI1dZXaV
DV36NzMgAi0OG9xkAGTXugyiGc/wpX492M3xM6tn8SiiK36TV4JiqJs6BrBM+gVC
hznvYklFSk7tGUuQdhdmIp9BbzK9HGKGAa0xLhRalNK6tNP8oNWr54UbMfZe/CP+
Q/Okr/I+VJ+n8BaAilwtydieCumWncv0WmV9/CYjfJ+7owRF13pnO5xXYXn+YoC4
BK0VxNxmxfiC7Z4Hk4dCEyfRD9Dy8EC4YO6EcsztI7AiYdRlAWpy/eK5Z46qxpmF
qXkF2OpRY6WS1Y0cHFmyWqvWZBQ7Mcj7C1NA7uIV7BGjj1xokT1LIf/AKe/M8YMl
CzyJRymNBRRtBnZXVfHAxjYy8hlR1+wwTJmLFocQ2AaLJzCV4/LnkihuYwL4yFhw
kiRF4dpOYfTWKMf+qr5Ws3iKbrmOJtUou71fV2y9Hlm21oXR8Fvw4y1/R17tIhnz
Drts98OxpGGSfGJ0OmvvPbXxEwSmh73KwT9PSrur9aWUdC1bHsQ0H0g9Um1AKcF2
v6l7gsSb1xENRQ1e4FKfOGKWauz70RD8uDByxXIcjDH4DeUUzCOXOEDsP9hFjkSt
o5ym1t16tUmKobH0NjpmIV2jUFKnrjAVLfk8HvsPEiYIqMAZpY1dqutCuk5yXthE
Q+lkXnodua4KKSVHGXJetBoCL6XtIniDP3DSSoTGqQGv5ZLue+U4Id3LGR0m4/gJ
uapxdP7eTx3M+8byvWfI/L+WMkfXozTS24hjB1biJ+pgjoufftkqdIcPQhw/tukL
yKFFFyQgsRfUZp/eFA8Dlnx51l9Rad3nFu5N5oCXbP9WHHIhTssvcworBJ/4bv5x
oY0vnuaHM/DX9gE77TxgderWXjJbc6a3IyZX5hB6snvck0CC6CIpTb67QezPeH0O
QAT3YHWHEwcWvPsLSNPI65FWQIZqVrhYCE33KZH5k+ERaK/I2cljezqd3ym41J29
ELiJDfympwXrdeyDCvjt+DWEX6QtW2E/1yQ0WdmU9W545qk7PxHidErgLv17hAjU
T71KHUi9xFiqLMtH9YnpNVF1WoP4/whGKMn1inZ0W1hd08dzEoCUcJ7ezsKY/dks
BUTOxnSH6siyuRlwl2wHWYd04pcfQcwmhjCajBZpL70rTbjyptqKQf0rEJl4ay1l
bqCWeD9XstkLYNfolvjJHIA6MvQ6bLBuli+gMYc6SPZ2gm8C10tgTDTUE5sEEbzR
vm2UtsDdOBZ4HlwGqEUcVxoiELsIAoSnsROjSpSNQxJQYQNAaArWvRXJx+ENld/y
SS76hkVviytCY7TxPyWPBYHf7C3a+xttvnQlor6gtljgk1ZSzawGYTtzXb+yjKg5
jDpG7gsLJaFD5mf7jbrtl7UDgbpLsBAUq/FzP2zJoaurkzs08OCqdObAzfquGwKt
pyN5mEOHr8ZqVjBmFWZ2pyGUphNLLlnbeT3rFOzupiYQWXyM16/MdEM1HgdW09z0
sTRnsU/dFvDBxPKqtLcilfsAPB2w5OEUJmPvIOVWAbMrEHkyxz1DLstxUnfpwtMP
wvWvQWaeTA1av+f9hjTuvSpu8yXvoZN3l9eC6ShaWcUWztixho7A0g5xnxFdqChv
U1uXdhRx+GNOz5NsIWBtE8KXhCl9hN8U+VZ/ea9rI6RIkIXLrWZiGXWArqfiYQsp
gN8qBawwCX3ZMmZCSWcvMWUUO0aqGc2I64aSv5uFxy9fczfppDxx3n0OyNXlrolN
aK2UOJowOEYDBOFkE1wz8t+2er4PW4y0lvBMlUcqzlAjzUd31cPimtdfqfpaDdYB
g8mpiFNwjnYew8e309xhg4+N/hSt/1btN6tAsOG4GiqgVMgn/bFI9Kc17/z+bX6E
WwC+yX6a4jjttNEXIQ6aKmJpaa7V/nhBAqfP+vyMhpfDoI7QaygXLPTQYf9NWAjW
v1rD5YBdkbiXAGwsWvnTSbmL2LRlQPswWbE2C5OJ9eZFKmp+gCrxIjsbkfZrXEt1
7LOgAZhX8ZixmTYpyjQn2AkUX5necZNR+G/3ueGImCE2Yd0qcI7XTuCObUiCzfyH
TYNSWww7Q6qIIZaZGZpAiGu5/HwQNbys7/UYOrCdaoPSudUqu+jL+UlUX0MAaD8j
LJEHeFLRjFQhNVJYdfycBMnCMJiYXxFCtzKYjDOmS1rjYUQuIUia6qnH3rRR5vfN
w9rXODRP27HERQtXmcuNifsqaQ+JlkBlhUjk2/5cSVtMoey+lgT8+tZuON/JDC1Y
qO0QXvpmajV67r428lhMVn6Zl1lKtl7MvgmcL8CiEldOz/S8qBePWVdIoXsLMo81
CjgnotfuM/ktswmzLAnmK6sHaH4dwRvknBxO1hJHnu6ZdfH+sPSGClGkWV4v1YmK
zYzCqB69+YJzjiZ1P4XYVspJ2vPg+wkhf5F9A3Ko67E+6+3eoGPNn7Z4uHxdW43g
c8fRxCjMpEWZovy2WXb6DUTTPjEX9KOL/kGlZYkZzJvpQzhTL5yJ3+SJfUicT6MO
ha8jOrClV8yfgRA9Z89G8aQ2gLzIpbr2xcF4hiX+j2h+abiQ/OmKVfsTR3jCUc66
FDecy/vaqsSGTzdHeioD3FRMsXHTvluUUE0cFcqrUYz3wYEwGIuTiaGbf3HhJj+z
Z7HgOLAW9ZBwnEXyH8Q6FmqyTybZvWFoBnR3GfVM17U7pKZ0c3IARdcQwBprJXaD
Z15qQp0Jjy2GODDzdJ440Y09F3X+g7WyFpar6d4JVw9AA+vpg4rdbiwAK7Czkbra
rC2OWIGctk71PcOe1V7USwMkm4GBoum48HsURpBAh5N2nOBZQM4ern6mbGJQG00a
Lyf4ULYu5UA7KOzpfzK1oVDiVTioJ44FCzOkr/t78uESHxfe4zhosRiYNQJ/1LbY
TgvGNgONPHscOsk0ghLZgDR7ei2ULlZGjS8Z1zmvvkirILHZMfJivHwLIfJSCwE2
BWQzNYcvcdhlcTAgntrZLmRhI7qqEx6IQjvb0BMj4Ck3zny6VuUiG1HQbuPTaImZ
FcGDWihcQoJQbqPIlxWCsNuHZ+gudtXMgjatq8p7cDZu3no2LPiZ6Dq/fhhgSYcL
eNp48HdV04czb5U4bwWnhluWsTg4AjOccUvhsO730XEpoelsnwSghGBudL5rhPRr
2+cRudnvFaNX0b7YBJwmyT22i4MXxR4fkJN0foCNP0g3i0n/la5THAbCczkwBvn1
ZvHWq/z+VEgQ1KfD+1UqVn6Viv2r+Hqec/7g27gXdWLh6lvO/bhFQmW8KxaHNJcm
e6PEqu7lRgVVapdkzUaM0VB95tHtfgGk1gnvTw3sBGuigkZ+ie273ZjwXlVGhxZo
3wX6QV+c2iYrsKZjwCb9WvqNWqEQJTutxYvZGVDQKcx1CfRTFSGFW1s8Ev8l80An
Q6pn2GddUL4jdCoZS+cBx7UQy9dn6v14NipanXQg9nq9s0qM19qKvdNWZhVemUoO
Bmcmx8ISddtVGGhqv0FPbsOKSebbiA0feDvVk4rV2VXiJzeSltVMFA3CQEhikZyh
xEPgRwployTeOWA15pwpN4ygV+DSBm0vMYdFSBo2V7aKSOduXdWOeB4BSTWrP371
ZXt9RkOuElf2VSYWSqhaQCn/ATgkbao0HzA4KX6c5qHudbKJuBcPV9FObmjvoML4
hhixLo4bBUyYOYcoIOLOWwingcM/ve/puIK+yMYqItWNzzUfL+k2O5QOmmhWGxwP
qtxmzYRsZrYPd7NMjtnklzTbRunh/F2t+gNPAGxq3jnnPWIAvpXtA+nn4MJNb+Q3
SrWUg1L+vEEpqNKPMZU8oWrGPsNocLNagfGDwupHEDETN2Mop3rJ4uzyJa9YfoB8
pH1B7Gg4bP9zKFkfIZW4AIgbQ+t2SDQnXt1R6Ew5qUYHIPdPjPJEUSJBHYjM51OP
0hOFKbziFeak4cDrSeNzSYYQZsB+dyM9HuY66ZvvsvuwJXa6KRd8DNPw5nhZIT+d
x7Oe29J2gSc5Ssqwq1X+wINxVviJIgs1LREVWwCyx4v/4wDiNoZk9AqXdxSWk9mz
9ZkIwsuPZT7DWuxFYXOjj4Cquv0uZ9PN5IumIkVWt7UzuPcYhc12T6uEucB5H9vx
ZhWLg6p+TMLZ4j0z+S4zkmDyhoFfStMPw4SVgKzdngdNP1lgWSaDNKLgg84WsEUk
bx0OOMITyQfl/1dJsgK1yz8DWDzcT1HrDo2Ke6UamSzxu4z9jsZ/M9wa2qVhZLTu
5dwnmjMFKvQSl/gzzphbGWCpfMblwOktrC4qikCQbkGY2Ho2VtXl6MR1ODmtjsmN
65+s2vFYcak0TyPZqIr1yfkQDEcTbscFdSwwTPU1LXNndiho7U90IC15eSmSEHq3
skXwDuAnWvu9flhjT4k7I5F/R7fSI1eCaO1eVhnw8aWfS0ScipBaCGSqZYEXE06i
YqZp3C52F0ZK0t3uZF3ZktRdv+ZXuLwZhKqQkSidMxb579dfBJO/z3vukaGW2Gqt
leoIe15hCPAK0DKRwjBF1/PJGSefiPKntubAgNjrZ2s3B/7P6NzSNbD8VacRKEj9
K+0bAaCjZYhmKH624Bg1+lG0UNwWWbLpZSQk5ilDGNwJpSQjEj20Nq3s6VEkLEw0
SFQuz4QOqUzp+brrT/5ZuIq8ng+MHabdl6bwLu3TaIOxnO414oKKS946d+kFE7ze
o0qxWr4YUeMw00V03pofMQtyt+VZ4mQjiQBvtGPP1ERCDbFdqrST9EHagXY0nwGF
E5eYfPp9mhTrAAYjgAzNDB/ns2I0CXgGMTNZaMVZ9rWSSMHihAfI5KF6Wd4nPYvz
T8amDsnRotGlRkTXNuVPvLLxY1Ey8F1AGFWtM5Z+W39Wo2OziD6oTCAj47joJqI2
R1m0exI8pAkfN4F/QxxQjPmX2gDSSqsoIeZHXPoqimtRn6U+AsPmISbZMbsE8uGc
eeQHmniXPY0wyL0I9VHDbugLlSN95+K+TUrFIoGvBW8NJiSRS/zdDx5mj+2sJp8W
W/GVI2fyki3G0ko3TA6TULdWGw5qA4a3zKAAk3hbirr6fCYmm5f6/Ld2HpdiEg3d
POquLsv7FohdgiqWCG0oXQNYSNTwudEq/uxfEedT+nrY5ByUJi32PYMxd5p3fc1Q
J9aGuySI0/KB7mcbzHnPqZdRAkkiNzN3c0n0f1Lcvv7mJXwKpu4CU3i8bRuc/dI8
awDN428MgexgZuul9NUD+HhGoPNMKc5thJO6ObO6MDZVpj2W4kGEh/zR08qtYeXn
K5fh6edcHpv4TMD8CV1JHUxdod1ZKepLc8vEwbEm3D7ZlCBvf5Qr7Cpbq9ND458V
UgjQNL3cBkvkge3ZOaw5V2hFDPgpynycoYW9Uswz+qAqbcpbTMM0WvfORWFz66YN
LtMASrxW0XF2OtFGETgmssD2WaFhNFX2FXb8yR9W1uJqSBOtVui3YzN1pSFpkkMI
eYXYxI/YOt94pMrKSp0F7D5BSsZkzH8F7GOtJgSZRgjaIGeR2rTDcyoXwPWj3Qvy
FFlMD0HZvN426MUiARLcFxXSRe3oHah4z4fm2AaM+36rmqneZQz8ZFRuPmOKA/bv
eGdEIR5ZdgV7CXoOc8SBJOugtLXVEd+EjLGGTdz9jY/igrcfsrnNTFWKErHQ3UoL
EfvIJiwCM/eWfTRLKnPBr9+XZhlHyDKLtf0dd+WLuiE33gliicP3dms1pb9gSSfe
BbC9z5dJ+c8yZdlrg8HectOnnisnaoTnvOgBFekhDqFGzE4MyLdTdumao73BsVXk
xeMOOgvQDotmoJ6okpgrkb9ChIXK51WZy2TtxmYGwVjzWtKq4FAgLtbeqAGie2a7
ySHOYcYV0Mvr7dSIsVIN3U1mr0oGWR1eS2SswR+E/Rtr9AY3O20MWrvab+d111z2
jNQr3Z6NT8bweQhhmPGXge1C6iDeby36iJ0oO6uoQeLkcbeimhMt7CeQ+/SPNyae
rQ7BADqwvVkP8iekq1jqgm/3SC4qlVKBa+0HDXq5ztIsB8jpN0igo1vLcTaq9OQM
whpaMJo32+BeOUgoHsVVKgouhdPNX9e5NMCCRLvVbs1zfV1iQM8MPfchAohLvxzO
HVhlaMgnPdQPeoJmhRR5Lo98k+2S1VKKQCruRP5RHfd45eqt5uwizkINyOmXnnLB
A/DBivAobptKi6qlDd2u8qZsKIb1sDW/+c6irw6cnYaplcxgjS8stqoIBORHJyqP
kln4MX+UlaFG9uXR/rBXDq+YNMCYlXndh0/NHJQZoE2Tq1z2f1oxyCPeW5RgDglr
DoHLOi5vUQ0r8dxp+A7VXIGxQb3Lqp65RHjdUoaHAX1QZbaB3/azZ183L8gKT5qs
bEG0QU0xV9IbyiZgSKhi/KaXF73axrLOnibkf7WSlGMEtfBKMU3Cm5lvZxTDKSUW
TpmlhsFSS/OakP/dA6S2i5PCUyadKBunw5Am3FipS8Mybo6XlC4xQ7H2qhE/sgWt
wXq/6GoTVpRP9TXK8KztfVRKeO5wKw3nB/Qd3s9VUCwZUc0nz9OqFozsMppL8ecV
dPGTQCg5laEPOy+8WXbJtDsqoN/4XWywzD+BqAk09u0neS0Akdp/AU7rxfLHITAl
jBp6CSgAiWOMb8II72Q+DJyOace7vhvDu+Bitns+QXKBL3FQkjpLuR4vjUOjou6S
uZEAx3FIe8gKzAx7M64xQ9j3GbBImIPD24XnQTMSKbVnUcRglAdN2nOitdnpGKuv
fFSD1hbwcoQfHz+tF9Qvm3jbez968uvJsnuGByfvRa5t0AAKEee7jbqbqx9j6B9S
rxYbiljpN17JJX9dE0HZ8XMVnG+xi9NED1cRz8Tg5fkr/4Gr77Jl8SvvLzow2UKd
WQ93jvGWk/xNMm3CD6aRgZ03ILr/N06PZwXfhahp9fnBqoq5xH4e4KyXhOWG+yWb
vq0WnCSjf8DqU+6YHkCDrBccWLVz2OOxVh0X0JzBnn3ZJHSistDiaBy+l0fisU7k
8VSh+npRE9MQwCRJfa5b8N/shtKUZz+jWUttAhRX9CKyabgzOChLCAhBLDiWy61+
UlbuRbZmoYDJ2vIrpQrOxqXflsCUlRS4Uk5qnjttpfJYF3QDSkc8Q9r+IH+fGgCt
YjjkXBZTpjw+3h88mbcTGnyJBDb6ACD+JUh5AOjW4pS2JUsXdH7vkkg26BQ+uEDu
qAjS1mTJFq7pzwHehEq3n5CYmhuwKg/N3ERk+4j7CxNtHlvU9w5AwZsfSVk2YU3W
EeveKd5TyJwPmbphKwLcHwhNkCNR5jTKEkQbJscaepyCKijzvZVPpzpitnBoVhNN
rd14mt8a+sb1VtA+4KTUVlUcQfHvBo5JlKnIqvOb7x6gwBt3CM8HYeUyoAXaMhFY
TY1OyVZs2iAjSBzZXZzjAP3/qUuAWKVAjThl+MSJ+e/52ku4lpuGQsqpoZX1GbHW
k+J468ujScPNex6ggtueU3+vWnb3VcnJf1pdfYqY8eG4RjfQuLzng/4atgbXA4UL
BNaXXbG/Bm1EqNKuMuWGwqiyfGjL0Gqo5iHXcd/yfwz5dZlV1IRmH9xcG6xWeaV3
4M6asD+bDyuAMafqNJy+kqcUAdLxYCxHwQM/3V+XKUl2c58msbgerl/NEY96Zgt+
LFWHibb9URRYBjXsZWW5fZRAnud73Gqf8y//G1dQ6Qa4eqrxnkTkmxwMa3PdCXQU
BL2Via9iTcTlJSOFRyFOCkc2dMxUGaZXbWqGxSUexOTWAQhMed51wxFeC0lXysaE
FZx5qOBfrARAJ/jeto+B1ul6T1JsZQgnkwTUkuYDEY6njj22XRYT27yvYTY6AfGG
d5q+wKq3q2AMdBDrgn7S52X2H0oX58ngmK+8rDiNMkftYnhZKxzzVL1GsQ0IcoLz
PjRuYRS+f6ztouPQHliTSlH8j1aQSojD1ngwjTMQtPcv3NWWKuqtj4SnWA8WMcaJ
Kl7O6cQLINWjPmMiWMfrYr7Oq4ouZYE8fo9BsLOoLHCaNhOwk3JDFbpye9l4Mu1W
gvhaUcTY4ChExyXTN3cIAz1fBehJ8BAOzYhN7AEQm4HKniHZsOSH4Mb8VH5B3itH
XYH5XgWAhAxVsRibSQWgnUyk8YlrIl8+nMkFC51OqkzpteUBpFO++2P8fsWQy/ME
8ii6DXR37ctacg1S+ErO98i7QVBylkJGWrVogu+t8tJ79iExtXy28nIxzu7MAC0q
/KXPadUjbK/UOcnqBxQ11UIm/PtUbQie1NPDfhuKWJyN6X/zOzzkvEsmqbh5g4zG
H274XLdsmS26EJQLsLkMvAdmgextaTtB9yiCHr7+6oBQdy66ihea7Pdw968/Lzz9
fHXk2gLdiXZPLilozw7OglMMp78Mf5+CD/HQJ3H/88Nb3hqcbRZK8ygRdhWCETKy
24PMtvOLlgJN+HT7OxJ12Ltjbfc7JraAcVL6lbTqzYvW5ibWRRiSXtBF7IOW//7b
dKNJQ8+Vn5Z83DOAHRb/LS+TI36K1JKZGBHQ6qrcesyV7E/hfW2Q9l9HR72Rol40
A8y7OtthWxe4FE/vZKUjMu7uuNSviqB072NaWqhjZx3aFd/2a/act/h3lCQq5E+1
fLa+AR5iaBWhIdkbSOJKohgqkKTpbiaPuLiRB2Re8YI2YCC4V+9mBpjTIf19EN5W
5o/K31hp5FHVUtr8oz82jTJZfjXws+lKo+NtO73458Puv1k4TlY/C92dSRcjyCqT
DbFgVaBMIRwtYnUZYs0jyAU8qXH5SEENsZhhJnPMgsTZm4ha9c3lEZSTyiIAqHJV
hiF9eK2nt5GuohayX230YfF6RgkGADFScRCFoxiw9zvCR1u0bV1ZVn9ImU4vcXFd
qZOOkC664Rc1CUQ0N0JEAw8ZX00h/5kyf1SW/XJdbtetmNMULk/1Z2wEjidwfmfU
WNV0SrvRokqHH+KLpsmqfISCYKLphGuVQziz94Qp0TjTJuY1klyV18UvFfuRi8Qu
oAHTUBHijI2qgZoJNjXPUUUyUA6VAyXxjfajSqK3AQGF5pizA+kz1IO6780UEbs4
Fey1nVmBzWEo0/cbIPJVWitkzk3NMLqCFYMemyjO47BYGWrb2FW4RGVyYo1pAEbq
L+9lgXD4Ty9P0o8CpHzRdyfMk6P3EjIXH56QT+pwvZUSbjOGcxXyqxjL2MJ8GyTU
6vV2h7t/tH+LEGI23lARify6ocryGtuMJROqKI8YIQzGgIWvFx7ffvsOcKl0cSKT
Ji3kvuqRSmEFcq8QVc2972azJnDSXjtHbemxbrh0GZL9Mdt0JY6CurIwCh8zWZuO
Nyw12s6wo/YIqFnqDeMzcSxBPBFmq6jp4VjLRCNofFK+DqIWywB0j3/U/voJX5Sd
U7/e6Mp2F1cicRKEIBwuBVYvKmwEepEnReuEaNBMHj5s+WjpTQOfCGOsSFUJP22T
DgeTMsBPoagFz1tYMpFREGdrf5fZ35ibfObxrwv4TY1yK6c52wki9sfDOXI1m+q0
wPiqpxyl5R1cUErgVbQar0hBiY8YeBSECkR7YzL+NFxPwGyghj4eVpQaC0zvp1PX
x/zlnqhPYHsj53Vq+4/C4WNAUXN5yGxEBcLPrUddcMYTGzdAvXtlEbeM+O3Y8tMF
KuMTU2RXGJe/j7gzBft3c76ULs3P99JGfcS1a1ddtHW8ApdSNri8gBt5ZylxREKn
PrdDnJDZnc70Huk/DKq/6RvrbDy8/pQA7C5uickA+3+Zi3mrin3UY0bg+ybLGsOl
LtRbp/7pCnI040ky48jBDYcTUsj3yZGsdr3bbYY6efosaBc3IpHyDPat6r+3e3KV
3IB1ghmOSh2lEH2MRszu9ABy5ZzOVxTiu854ekowWYwqiW0S3aELIC1ggC7dEmGM
7IaoqYZy9GML7CBqFnwB2LML7wfG6Pxe8gOtM4QjEqXFlIkKKmFWlwRhj9XeoYqC
NRleobClOlY/TCIXgo+fE/BND/Sp8jQNTs6hVebSLriSlwwOKncXETMRitMHAb4T
wSPJdhlBl5dkqvF7WM+a3oqnKFTpUft+C5H9TC92Q5btI+xfK/MU6F0rRDOjCN2W
/yAZmYkJh8ZzYGGqD/zuXDabt4U+sCv9bbvI7J28tWJiA9v4OZbIvT0uCc6NRQAt
X0EssCZ+ztd+yDPM19q4sV8FU6bkEj139Q+Xpe0Tr0axyHv6+yRErTd0r1j2KMlu
NWVqIMglg7sBbwzlLcAGpBQUz/GUFxZjs4bCmVIkglojvDb5IAWcsKxVmCfsV9vI
MPDfE20FtZ41UqHg+kaTRIJg2oOIOvxza2konZd/L4NuPDGJanMNOnhasuHlh7SM
IHampJdCGHDcsaGJEIKHdPo8328JPAUg2RPzFu4PEFnvASOjpwktDPMbdCQZKYjO
WViY/E13HwDjAc7hGRCq8RiT3jmo1PKFbnqMkDnX75AJzzTumfde/aQYwvigehku
esvkVlxMStl3krbzUtN85KrxnusMKIVd0JZdgt8/Au+rpke+62KOE18lDtG9zhDj
3I54X1+k5m41lr3P0QBZrdEyXLP2as1KqUy9ttMEaasFR9wNHANtTdYc8zVKOAmT
rHOZtOf2akU+LhjNmcGcX42j3cIkQMkW2yDj7/ojR69l9kAphkSp55cEgTrm0pn7
RqImUKFO1kXLuaCvUKAemalH0OtkS4kFhwXAIG7P84mWVFq+O47zpY8bnX4pJUMn
DRsz+khRWrydo9LQbHX+yO/GpSOh102YolNtrBEAbJqpnxKnuPYVQb2Cv7sUAeNj
eedUsmTfnAuUdFuEcyg2rinykybEgZe9gSxDFv8wpg5Oi+tEVxG/1rwdtmF7NKZ/
DbK7jbytWa4OASNbnvqZX2YGwTZIZgrfMcguqvn8MYgtqgj2aTtY5KWBF7tQRdIg
di1Fb0F0hiQ/QLZ0nhFo/cfiiD2U3XsoNyodRfVH5AuejVmpL2r6xWNiBCuKwYdl
iYVmx585R/V1CbXNcYYiyvLqlTfYuG6gQOxYI0gSKrQBPtCOmLbh5Cj7caEMOl2y
mv8WD+4Rvo2tAji0n8lTzLbXzKMagfb7Eyi9ZrhCtlOFBlPwq372D5ou1izMNhIS
6Wmt/4a4cY+dTVXKqVsi1LWPVPfGxgYesllSaH+kK5VEcDOv4NdVpamUuLD4UvE5
A1gIvgi/274BbjfkDAJFwfAspwV/ZNbRmYxizQZPrCa4s1GiUpj67M8nf5lVL4f1
DibewJ3qIBMHPu2BL+2FYkNe1W/JJnwDt/iSC4CYEe27GEwGSSxOCh8ncXqxWDMt
byLO8EgtyES8WYkUaBT03dmpoCZREfaY44RwL7we41jdjqblNxt/kKA5jXH1P9fx
1RkETaq2SHVPn01g1ZoyrzhIK9vKtBGXhYTawEhcVzeqwMwWWKal3xROt1bcGSoY
kZdA0rqy7r9r4SEqDIO15UffQyuP2KDXwMT4mURBjhAUDehgw7C4BQqf8Y93TTkw
/eGq+nrY5BQ2OojYkZmywzbCghLfFD1IQt+v5t9nwYUC0XS9fjrmBIUjf3A25uj7
7887YU/0Xy3jExtCUDdM4CqSLpamldzrrOkgL36xREJOOyFWTyd38qtxRo9J5mNw
X5KKePSkK7Ib8bJjofX+gZv88kyOmQOhqG57CFz2DTeLkuMOSVU/NukakNWM/58N
n5Bi0GmdQtQrt3omfTTf6ez0nJzxONR9dyWIBm8D6W1xF/xbQ8g3XXdcDQDHALAI
KsdTds2TLO7L93hJB08RIqV4LtgdT5dk7TTtfJpNX8Z41Qom8u4QF7EWaJZS13bL
DfNe/dUqwqWcU9P7PkcdKp+/gIASh9ghJUERLGtTdaufDFs+7q6mIr5fJ6wC9dNQ
9dsEmIO9v8eVOlfRo22st3UkvTKhHyqAlOTtGO1rIo7kY4NGuNIA0JjR0/0am+5G
FLYGYRrlSwalvZOd3D3c5wkzpPsnxvVLK5nro/udqpLyKBTKyDNgF9CgzECpFbNN
wY9RLTSJxgG+ZPj3dvw/CyeMAhjoNcMYQrbHEyY42I14A3x/990mKxg/k1oUioSV
8FTBCh6Ucuvkmvv2mUTcZzKiVXBHDjtoJko9nN1pwliy9BUIV/7LuHznjkyQilmU
fumfadTVNf6UbxAgj2WvsVEXrEYT7kZOvzrKsL9r88OgH7XnErj+URQLzN2J/YCQ
0TzvuUN8YyKa5/TamrHgp0515wNlZLxuSYy0fOrHLZFszguNXSNYSNTB1pT7cwWS
QdogQeFsKtehlwRyArxfZCWZwX6WhjFA4pUB7f8qe/iVHF0rNNCAtECSj06JisQx
jzUDN77O3NPhL5o7y1a3mjvl3jZxNA6J/SPlsyIT2fg4BfZH87ol7rzxXHVxxSpm
LL3uc1X9oIL5QMRCF2Yc51330jloSit0BEumebkXHY5UFbKOvO7wJOwz3RCjKq5X
oKbQ+tuG1lG7hkKbGhHymikHuttPo54a4qyfX1TzSSFO0czSgmWA3Joua/zcrxiC
anFZh7Y+zRh43nY+JXjV8SOxXxB2GEzzZC2jg4SLcnZjLj6NeNUPDYaKbRaMxRnl
pU7YnFTwtVE9g6D3pjaIgsjwv98lfef91PCerdROUQiIfAmwAH7VTSHu0jOGXjjf
yohJWAR3w1OZPzuku3ToyY3KGnefp27JNACwJ4QD8YRyBLe5+iYZHgqGXjiX7EFB
u18dZ81GZhutYqXhbwrqYLiWuUOJu1wOmZWfxQhS8FoMgdnCb70/54M2UsxUHYEE
vw4cc7s/X/pOpcsIUIT9MdxD7k+Vf2DLRXYvc8Hgjn2tUSglC+d10QkTOwtMcS3b
Fd5uHeOdOvT4gBDpnKytrRwv4Ji8EJ8R2iVjRjCyiIHM3qpHNZfUHVRBJrWpuufs
yQ0KTIpwtMzBgKL5F71ZlAv3qV/5mnZkLpNkjwd+G5iEjb0smQCSoBxQDYoWgXO3
cWmnvEYUxE99El3F3qismHM6fHEiAErkchSGSrM4V/0Pd9yKzbqLiUCo8DbqPxVM
NeyAuFKX3TtGdq4aS2w9+NaqTei8f+k8LcWnIYHhOfTxcjmh89/HLMfcv1Gs5Pw1
dXFU59uZzJUuVhEmHr438XQ3mBLBQWvlxkKmzPcIqbnoKD5BT8juQgkUFdjKPJsO
xMS1G+OnWj53ddMob51iKp9vq0DWqOxBvto/ifr3a74Q7XFVCDz2tx76GPantIiZ
U+GusvUPDSZntzFomkzOh53vYFNqHPq2xMfXsDm1cDyAeAk21AlWA/un1K6PdOMW
uT80ZU7MqzINRmM0jaM6eHYeSRcD6KwtOtZ2XTji5Ml8fH5W6O/CwqU7op//6Kmw
lhv4jBwvPrXz5u3EUSP8uYNtWVAS7hFcGoInZwcD93ExFeUEPW2JaH3mrki/faDq
aBR1OIcv+9im1gqps7AH3JellJ6QHT/y71FTJJp0AFfe7d4AubSA8tYHpoEykgSP
bo+8/Xip6v/aPn9SLSRtAHD30mJIgH4En4WRySzldOlVyedOUifQkuyitsY/leJs
kbnPIl8UuImCfQnmihPVVUOYGvbynTl7o0pP3RJacEVeaBVTvmGfXqQ5upDfZILY
6Aj3Tj7wdjAFN8HAPLXRNFVczmngfuCUOaVZhxPwB17J/pkJYuxLEmyHZagVODmL
m5VTBa2Deyi6uFJRFriUyzxL1xMNK+Zs15/lbqd/1FNfGE5toopCKQwkvOsp/yaT
oebyw2ghhAHJ+AZUJ49AQGLXgLZq1OZVyIq4gW6uInQlDATk74J4otHZK5oxCftg
Opy07IWSZ+zUMeZPRKyCd5hfuZVt29DXcEH7/PtURPSWjEIxaY/y2d6uCIVAHxFZ
tWk4kOzpIxujpYRlDNdDt9lZNbnX2Nm5vtz6B/c5lR5Px6br9CwN2qOXFsI0BhuO
ZyNPBEeP+bqDTtgihCYEmkLFr75cfRMTioRWvLQBt3y3gk0RliJRh7YNHXUgdOAi
1mdLnzJYQ94D0s9E4qlOiWpQmbc+WdLo1YFjtUJHWp6A1K1mAWAI6Afivt1yrAj9
V7m7xtxRQR1BIjkISfwKSAc+y3rWuz16cGRpRRK5Fgk/y4spnyOLNLDLYZuJi/0g
MDUdzNVgoS7E90ugMr/nQ+yL/ZiLuLnGzYRpPhPSA7JaDBJ1Z435BaCC9CuR7+k+
EO/KUQDGMdvrrEFzQkIp2LSXMK6OCunrCsYY8flCqX/WnlBaXcCPmDX+o7Y9naXW
byAGXYn+tuA5AWM0LXjt5SbleTMzJ8KbGg6B7q1QyGhe48WVY23RxC8S1a3hDkNN
utfZSpTrcN8yvPv3OVM/PQWTth4uaPDdOYdhy1YO+POUcrGwaeqdKmNtUd9S6qI4
qXY0zmaxD4OyEreNjwvwAXg+VfzR3uyD72SUSUfRS2RQE6b+hos3BPA2+YX1QYtw
/gVkKAipkz2nKhruMR/grquYN+v8tzCNIF5jifp1CVQavCHGMTMeC7kqD6HNNYNF
YFAO3+oooeIIe47pmnjiI2aDs96XPbFD6Ntglxf8UYtwMArhz089rV+szjrs/zOc
dDfGgaiIPTdbaInQpKCq1Vtlur5yvAG1InqR8QaHhqTS+PfO1vv6uXYEdHL5pUrY
jsQcIDeyfT9E2H9iFpL5HGCTmyoetM1FufFfCqJwTthIXOHJuoO7S0XL3e02WP5J
tWTRq0i38htbbzLUZKXGPj8NWYc0C7xwPMbHNeNm/pypHbjAAN24j5n9mXitlRj5
JbXWkuas2Z+el/wp5tUwXJKqf+1hu0yyWsOld74OVwKTEg1NJYeU8Oh7Zl1c7Egl
tyk8hnjC2mDApGVz7wJKKIBxsPz5W5kQG/sUs0wYJ8op3mEr1LYWhsoL+IX+KCAV
d305tg89YBEik0TwpG4ppTYjE9/rwkG5CagRqREwmcNm9uRObtOeiEZ5oWx2Sa7N
sM+AO0uj2JnnXTuiZwMbBMWXQktcHbXzD4VyeXrBwYRoinEPJ2lIPF/o7yiO8vOZ
pkVlYR9Psn8uNEtq3KrzvvNjfZUFCCG1cWb51uoI0YUUNznubqQPENerco14mCV3
hWGXaSiEKiqKgL9uw+uejWC7Dr7xWAN031r1lgruzuMgfnECXyCp1POzkdMlvqTN
JLEsPtONzH2i2eoj0xbCahayVQ9SZVcTua3788R/UUXn3nXAH9nwp77WrclmbKR/
WkKXl1VY8v3ivjDhEpQJNJvuCkDXC42DWuUSb62cXRQQgdOPSOQcwLKojCyI7EW7
AFXDHJS1NEui3BFXVtP3WMxq/a0T/Oc3dL/oY4NK02iAsizQf/dtQ121bX53N4As
DTyatx3mQY4HfUpjnQ0vnfkR10UnGZTvXDAEetf6HExblRATt1m+/uqfDOPaguPI
/vTiuGqFCxwWOpbOFEsfTzx6auUhuXmrGBJwUwyn8PpjuiFRaMsozpREGbYSveJY
rtH3Vd7IBqSLMzYw5ftTalX9wDJl3qW8iTeJ5CO59Q3UWCv304hldaFtTjVJKESY
di19qvVlRzSZwxdK9d0r9dPWpiiRsUFUmKmt4PE6Na12M5tQ1RCuVQ4rduDKe+Xi
6ZembxI0clIiHGAPLRS1zBYlAJuysRyHHzLqS5z0f9k2bWk9gzVP+0ZnXUMuV8P2
52qeY78+exaA21rxNzc1uI9XFngLQdc6wrVKCO22j4W4VidU/XTDhBRiTAYozB7S
HZCqkrrPPs/tskRWqmpxdpkBz2gA7jSuUQ1wkVAjvGdYPcb2JDpGj4A5zpbdzn2C
C6KtgC88B/Inu3/KHi/y4mZ1N8mLnQ4WvCd8HRP7ajK+MTyc0H9lmfJmD1X52Vlv
z4raLQbOWUETC+TgSn/hpt92VLZlnZvtRjPdwyoe6uh6Kp1hRYYQlmUOL9Um6T1R
FfqQiYokipy3YeQPQqdqXIsN5CAbmZZXcHwV/Sgo7/DntmAlTqucz5hpop3Jsr0/
7D+WA2S9KIfuLclr02R/YonVrPyOy0Y0Ih5MaFlBLcsi/HO9LkRCWH+K2SscaSUS
BwHulAHsHanCQZxZFeZbP888RXcdg4IOmdvN/hm5A8n/ftU9pea2FwEOpW5YnRj2
te8MOZKhTMhDN2e3EbeucvX1pD3vQ/J7XMQK+HlmGXlaOH+w5sMWH53EVblSpmoV
fiQUZSRfanr5b2wANBGiImGfw5g+D3aLkb1OOvhg/pYdYcEANga7SeesRVW4lFAU
TzZwRCY8LLo2WgmOna80jJ5ZzDAPjv1W/hiUgZDZOc3aKCrsjh2PrvZbw5jzrQKf
48nRfJWgPUqkCIUPD1HfwmN4tMncr3OSFpBNt3EQH6midehQDPb5J8mtaIkM+k0A
R0q6x9b0ucrCDcs9RV75PnjpZHSn35ObWif3Si/7ege8Xx32/I29typUQAwn/dPV
pDPH0k5KkDQcILuNz4lHYa9lS7MJufgJ1VheqqUoqHOYQwJBHTJhnYPMnMDEbjyP
UZN2hSrr9hPCeXTbxLhExBrNc7WLn9kNozdwwNdkgdRCRyAPupjicAAGt49jgYQS
XTKIGddJEG3wa+b6kLnmJU0D9Db+bhkzjjQgxMnfoYAgbRYIEyc78RLEl0qItBoQ
Rx0geC8kqwGm+UZQLSizBxyEYwnCTz21EXsHC7OhOqyS/J64cxpHkr+IWABrbAFw
r/Fb0vhpUdPVqQia++aV9Jo2kwL4Ew3ApwE6cUzpsSD9KZ+hJ959qH9bQSXZHhSN
kXR8r75S27v0nTn1/ccpcYQpcu/SuyD7jJEVAQraHZcGe2O4/s5r07BNM5DAdxoT
uaUwKwIANWa+91MK8KSRDMybf3/kMSR07hKxCuOM725eZ9jliXT1cilAwa/h9CuB
oddIGcXI3oXK399AGUgGK08B7aliewmCJoarYlNJVhoD3uXJgHBX2ERDozTZPyMx
eO/Q6Ix2e3d6LP9H3RGV6kEPzXLBtNooZauTb2r0qtrXcIusdIQeu62KugqNarcg
+9Be2MBbp+KNCftXC3FBgMVEX+z4njP3F9v+PySEEZVfTtY6GpYOZADX0ZZSp+i3
2rjzFRGtGUCNqpoh3okGK+E2USN1LQfFCc4g7FN6bvXpiQ+MVROFTghiluGuXRk8
DoJR8L4acg8ZXVu2C+dMk8AiN98HGfmIrpsuxyGq1nqOp9kl8kAdMaIyUytIHcA7
tqkGXWcbY/lsaS06nhMk10b9Y5nQbtT3RHEAdeXdGPL+H+MqSRaR4WSRcrbyZolU
/CNQDp2h4TDJkYtNCqVh7MEFD1bIMZi6TcobEEBSK9M37hvx3er1D4oYY//Vn5ck
/D6VsfVeTqNBIUgPi1ppveTBC44Gr9DSVTAeAVn3uUFW3nuYYxboIuo3sBZKchGW
0ewWnFiGlsCwlAOaEXCII5Lq13/MCW8lw2Gan6QgNPxHVLiO5LnXTMHlVWzqAb+R
bSEL6ccS9gPemWShCAo/s312POEvwAr0OHDA0xdLA6AtXznXfRWpnGJX5L7TIehg
rcDkLKxw61tJ6LgD4H3iFnOK/S5GwbKeyz20GrCU+gXtfevs3u/piZpXq+Xn9vY1
ynQsiip+mb/XB4Rvl6Mtu9u+EM4GH7cDM9rO942a3wU9uOlGMHTSgHp9DhGggjfH
N8fxpNK9QsxM7IGEH9VQCga1s497y2rrEvl0DHtM2f6i5CVy49aJ9UirlPbI0vMm
UzvtTY9ZOMxKlj11ENtp80DM9XgS1bNynqKTAZcbKiuReL9EPvh0LH2RGy4Na0AV
qSY6+nRSrK3CEQ3/8+x6gYmOQxvZ9OwSdfSyEkoCltRoTaZPOMLFrEDMMXbD4Xon
tiADKcut0muf9HwuiDgiRCqOcLJwtir3SygJbWgbNDQCG2myXitM36Cx0nS9KIYv
u+5cpkiTLFn8wCGulXWA3BdjrQFKkq2w+jKpnSI7Rz3kR31KSjATiIiNqW6ub0EI
alRffD4CYHmFBN2f9hURuxQnkfGBKax2wWcCpUGFAuJngD6101Vq2KZuJKHZPdUW
nibKS4zCTZQ0xCbG8d85CR/2oh2gtEQ/E1GTNOUL/k/KrE1WzQYN66HF9iix+PKi
7lJHj5oFnHRaY5jOBGZjpU9WUhoXWEe+hBoZE2eGlsIZX5zS0PjxTUmVNz0qprcH
X80R/YXfCuDrnJYw6xWwgszuoNiED3z8SWpsth9/KsFLL+HE4fLIdb62RNoSWhsv
KfPR2SlKvL2RbcMPYmK0WuEJOuwK3SqwI+6acE0VPdVE3Txua4MfCjDGyYQpCbOa
5XQJlEkvv87aLyyKq7exfDBoLl+z/kZvG5amoERZ8G0WmBXzAEufA0Vnp4JsdzSu
uWjpJyth4AS5mW4hqhS1i/P20c2ITvf4t8SeWGsUOcg9Q+7V9/q/DEyn+mU+o/KE
Eq+JFZm8r0SyEkL/rn39Do125Tb5plYUa/SkF16w2JVLjcyCugYn6FX3TnoHW7gX
LZ027yrI0siKNkdJ0HpuwglIRl5wr884zBROGRKiTo1bs7Wps4T+K8avqfNRaal5
Tgp1s5+FVsE7YhRnA1eMuL29/FZ9aFHFZv1Y3CO9SvRbAFxL7xxxECgJPyCi86wd
ZkFQ+zhdu+zkncr5i7A14q39ylleRUa5mQbnUHwuJO4c5IWYiYa29ZgQh21IpiYw
LAr8B7M0IfVoo/nJa0qhJJ7hLABdTALp4aKtRzTyq96vTMqV5O3RhuyocDw/+woX
22fyG4vqVL6TRlNXogQ1buzCEB7hW88ZO0NQY6wQBwTukj6zp/F2/MpvgoMQ481j
EeLlfv+VRzI4doYNcIMfCcIUItRBYFpo+c3ijy9ixCJS8Oh7xXyaO4FLlH8utoKr
Eh2chTQ1dhkiy1u8koA4sCGAC+JOCFeunQQdvW+aRDzVnuKAxRkF9oGXKOT1AUrE
iLN/pANMzNviPw2ziDowLO4yiq1gN7znGFcMAcJspytytlfYQHSczuE71E0N3RuR
W0uwzNkRxc1R3raC3dwJqPrrj803JdrSUOSzphQe1o4z5LM9KMoIRC94S2y0F2Ng
218Sn6Lt0I0G2976jDonUJZQtamxLpk1w2Erv3KeRly7L/wiGcvzcJwosDLT2q0/
F0gRzPw3xiIZ/3rozVtBG7a4FT61GkuPiWr5g0HL00GkqgYiPuE0g11LhUsk6dXJ
Rr4lmg7msHAOA3mMHPHqyJwNAVjQfuLPRdriE12Cccq0s6Pl+3GcCYo+HtlHtQR+
DJGQxwFGvfe55gLeBRRVGQYqeCv2S6nblB2QVhsgVgUzK3DAYiHgMz4lMVp2NmnV
3xUqSE10bH1ruOKSW462jVw1bDAOaeDusNwLBx8T50Tw1UhI2+fSmlALDX4IxU0S
meJbnayvsqS47G9FL1uu6u/NRRUkwXwrP6pr5a4muPX3YAKIVP3HrFdVPoa3l1db
Nw7yCJleXRo6OJFWvoiGkVmti300y33d/tWAWc5Y5ZOJP3GEGubHOyPtw3CH5Xf4
JUwdEwVMCJjHkt8pynLkBn0HrLBWukKMwsEo+GldFImOZzFJoWMcjpFtodONc6e8
GgKBj/h0VQaIc7hibEo9g093x92r/quKi5vjiWKBHxOqypGvvZT2jZDpi/R3wO/x
yihQPLTwnWejcoT8/8HDn35ONGOizivcWd6Xj5jlDXPEVo2TWjkMX2DRR6Va5421
O6E6sOcfe/BrO5UVzNw0lJsCaEgQwl871SgSQYt+W+RsPXUTqjNPLKA5qIVruGXg
T4Enspnx1OsiQ3mCf6AFurrlaM7SKnUTbtAXDN528DzKiZ0j/pCBXGY/Jui+40ZF
UcM45srsvCmZ/BtliPYYVYAQUt34kha5/RKB4PEsULrG7EwpIi2pqbPpZhbuVaUm
aH85XBCb3V3Aj0Fjv94qV5Bz7E41NcVPw/3MD8uOf9EyfaPkflIQKTsoY2GHVZhv
T0+X7xDJDBEtqsr2N80x9AuVWE/L/ActlikjKpiDsNnRewVTTL/Xu3HTw5mpIj+o
p52wXiDlYqaBl/jLbY2NuKpeIX/c+eyGVqOoLRFZSJlbAJU3K+v6y6bWoYFkIsz1
Bl6f2aM6olmo63q55mgeL0Fbqk/PPXRvs57qrrwpZorSzXY1p+6QrgUf8038CYML
+cC8m4hp3GtIJMSuhivTt18xW+g6zAi7jYEs/j2aNuH7Qfpofg1jcOz5bRSdWIRX
QkFhfOWclj7mXVKlxW/HgaeRn0fdDmp9bOj6tS24M97nAIC7MX1htqKnNAPLUIue
tv1Zgjie5AvwDksu9zMJlKZiUjwIVAQgpqxbDSxXZe9JqgqpBTD9fchkBPnSSFuk
tI8Tod/4RoFsbQW4vUb4KsK9qqqvU15jj2XGyre7WV2L6tU3rwbfuc62BTebsOdB
nN+kRdUmbO7e9A+SwgLSE9rjCWTLQgFm4HLcC3ajMzUlnKrix/9cQEKHmszUwP/W
ik77HPv99GJUBX5HNrMKhTDGuKxLZmjlZRoNMxeHrWAPVB6hHyLivQ1My5lzW6rx
vOx1SGmLtiBebZWis155Jbx8v7lNasCXpa3fiF/rcm0PBBGtO66pd5tb/oVcwWH2
QMoBZNirwNw8x6q8g+3KKEbdqS/cfr5HNBNuvIVp/ftRRMpb9zurfP2QT1DqYLnw
aWeUJfdkjGN2dWUVfwHcgM+c52GblrmCrH5bC/q2Worh3nwVD4VvMfJ1zkwQuHAM
lG9eFeaPlWl+XTx+M3AM+6zh7B5Qy6SeJ6f20b9UVv2NlGdka75F8OA0GguTK+EA
I0s9hutdstR07bh9dEoEkyFU6Qx4P07ekTroPZsSi9ZuOCfmBN7R7nn7rdyjFwMK
LQM9F9ChQbAn+nsV71u7T8cO+wVq10DebjkqjcA3ADvWh+ZsVHgJJ574H/0PnZsg
Uv/BXia3WbujMzPu9Z5W553kWVJn5wgaWH5T9kwTtPpdnwB/y0p7VKZf0SkanT3K
kLBixryr6OfuWsURTtCS+RycuGaH6WS0nD0l9c4qtNdVtbkxoNITjBaGwaY97JcE
JtH2UT3WH8Cj8H5mQftsNHdR2dlDm/s4BSlttLnBsBmSA+kW0jW2IM9IefcQiXXi
kCooOOCOaCmj/+SdkcrqhFbR7hkfooqnpz2qjNEFf6mzQ4HPmN0gpWQD/Kb8RUWl
suYXtTyTw1qOIwGg2gnhtIphOepAdkYpg4zgcKapeGTavYAf/sDuMOhv3OsAnkGr
jdel/voQoHieTUovDRh9KBEHoYDz2mR7+p9D5XVPJ7/mitvptZfqbsnilpGPnjuf
PCTXGIanXONbOyEOKODPQy5kCpaCfI7Lj1+vh2P5woS00+jWekA/3NN980TE0EaJ
VhpBZp7C7vrCavhz5cSoENs0tP/ZkE3D+DRN5ZQjHzhSlqrUrngHi776AJ4L3Dch
GrVd50jSLfXEsgml3Y4sBYlcKnR4wfbh6tCbqQ6rzrZuaT7ZUpodFEqhEVCvj+Xo
3tnU6Xxkly74QgvhQ7tBF9ydUavoJEFk5kyra83RvfA94nvsHfSlejiV/klYPfNZ
aIkNFWe3BV9szBMK10evXEN1RHgab+sVuXrHuV5Y/Jf7R02gNNFGtLl1MaP4CDqe
VieHiK2kF/eJ0d70Vn93kpP0cT7ofYTTGlh4EqhAfIRnS03umdrh5leOefBFox0Z
KzGifyCUalRn7MWWE+Zlh97R+5EzVQ5BuyXqXNEAwBltakKmlOINeOdAbDa1wQhQ
8Vf/z8HNBMcRUCfGtXE7J5xPWQPolgPloQDNvfSSw1DnzPd15kwCBN60+tgIlZA0
RZ7rS4NjA+9xRHiBLexpclCkzIjytq49cCwpns7fQGX9+jDIPDHd4Cw8HGKP2nu9
ipQvBOw8Xck7jZh2NX/2K0p1HeA4G3jOYcs4gV/Kpde7fa7ehftvvgrdYEqYsAS3
nognxVX4cQ4fSckcxYWhtwYBwOI+Ui+EzQBDEIyJo77AyHkcfMIUlcEU1+vwQ//Z
Qzxd4YW/BTdkzFWI72W0im7vcjF5Ll5Od87BAoUwUeC9zVaIZ0KfikvrrGGtsT9w
znYEjvXNo9T5OX4yuXFt+4pxu8GQYfYGP1h6kqjo+DKtKjXbSyP6dkhjzQsqd1cf
gLuU8Kn0ryqJi22txUQehCxvw6tXNC+rF9yQEOimB/VvpQzkQ2ALPOSsq54KvoRO
/QLOIHf9+xOieVa+EKUJIOUz8U5L76I+LCWT9l6DBmzfbFHLYMScHPHDhvF7Sx89
BxP1hw+TLz+mCWebId21VJD6g7/U8VSF225Vh5O7+T5wRgAZ1/axH/eJcGoQ8PEx
22KX+JIWgQhVqgwSxF7D31yMt65JgFppC/sQwUbrVJVSm8dpE2hU5yHDVz9G4QJT
sd1r66E2hg4I4fSEkZ1n/TkxTVrKZ6Evog9Gl/7IukUQXHJtaX04c1CG98Y6XXic
hkMrCHIZT9fCm+ALLNvrUIOKr4L1GYcNVlafEOjcZ0ftgah7Cuo5ADKqZrVUl0QV
jrHbAKIsBPBl/Dhio8ThdobGq8Frsb2zXE+xShdahFkSD+RzcRzGJB+7kXpCTimr
duPvCBAr4s6rGFR4xTMn/AuDyrOMEi0vGf6Q9a6C8NdBvQlpTSy24AVFr7idT+ui
vJhX5ITnZgJXSNHZuGlzIqQOrG9WSyYD7Z9SzlrQR/Ghp/uegtcWLFdGKSB6Pf7J
faNSicGJzk/VWsRyHzeYGQpCD6BdO9pxuoa7cbLugJLHzUBXo0kWrdU0pliVBncY
HnqPFKhwuWROmK47aWMQCEZv2ssDQU3UfAzHDNnNz/7qxYsJfi1fpvVJMfRLZuUY
XYrcBHYomRBzEmxLywp9lyOoh0uy86RuRxApn1C4XM+Mdt85oQGYo+/1bOIexjIV
JLSeku2LEbKukkuJf0/Ukqi5+uSu2GxJuy63AZaWNghGFog8OEbbcBrCjhAYhKQA
g+QrlYMDMMaEZMiPhJ4O5x4nXJMpjgVTm46yf7qb+MSszo1rrn1Cd7bC/ryqcr6Y
WtZTW2oQp/XkBxgRP1NcH0JB/95OAbOJMu/Y+VLfsoSqRxUx5B21qvZgs/IFIiJS
Y8yo/4xBjA8vQb3cyRQYkkP3Fd/r4caIWQw+/gROEnLuykwq58peifdy4IaHv/7O
zNHMGCI53+yzdFT8oMRJZzKD/UO/SQUtllSfyjX5JkjXHuRqSg5evA2IIvRrCP3U
QEugvj/+Fh6PIy7LyFVYVurvdUJTkCihc4mTU6oohJeAucJWs6jHdlTedDj5YwvW
ZdU+lmNYHJL7FX1yTBrUS9WlS2HhVn5JBWf1e9p3s+6kBFgV7Xrp/cWxxTSNcjoP
Do37BTpvgIRdA2lKsKC1HhRgZPl1c1eWIIJ6wpiS7Kf+UnNv54kvYgL0f+wKJ7oa
11RRHYu3Eg79TdQnMAe1e1LXMfHaNFmCWbsMwukxjIEz3mOC2Ihkya5vmVSk1JDs
rwvPvGr6YGnnil5yEJGxNSZIp4LVIVxoSvh2CCJw+uqpl5NYFoH5eXmXNIqWfmow
DTYQ5sruGans/kL7on+ErhR9f++ZMrrTgdPLTtaVQbiBHoBX2VaqMLz0iq9K4S3Q
GyBZdVecfE8NxnW80hUe/Tuuiy6X2vgkIYIq+2V8aEh744EHVxcgfMLhLg7BoSVC
kn8DM7kEfkU19UceLZ2Z2sVjmPFwgihENskyK9oBTzUiZ5KUMqiQkX39UdWfaOLa
eYlO2kjK+jTiLVH8WdqPBqPGqnt+tfzP6jNJvheVOVscUKZ3y5y6T+o/pRtqYiNP
NtPirh1vU3+JV4y03+4oNHeVp80h2MeBHGWm2Tm5LoJXFnyTZLu9tRP95c2z5as6
dtFpS7MpcEpynXfc9ZoCic86dy1SO1X1iCZNou74dgfXU17gl7GtBRFO8GjLuZ9q
aCEoZBKjzNzvtIieYe2ogqWW4w9Vf4ZlAA8SR7KWhb7SfFepiOLvyoeJZmIY6SAQ
Dea3TeCQbY6PYEhccned6O7V3fiFSUyBHsXpvxjx2CCynDC2eYtWk2p5iNQqnfVl
CIjA2MpwzXtd0QuK64C1OKt1Mj9nXHJ/bKx3U8dx68zr4Z7xClNA2FI0ClEjwpcb
yhEeS2gjeQJldkIYFKfBFHkXROYGOQl22nC9NlijDJ2zFbC4nNwpD4baRRuv44HT
GAKoDrOcL450PF3SKSQvii8ahqnWozujjKh0zDQwyRXAfnYkEWewyZzxk5CmaWTY
GQYfZEk7nCJ+bcNA/pJ3IZqWY6/K+gG46QkmQldLUXoD1wJFckQI53mX2+IVhUmP
RtEDneCIW+1QXRHEhjEkqRo7Eqcjjy84xX0jB23Zz0HahWqJdsz86+PmCLDb7j56
/KAcHmMo3GreOUnbJR9asi0/7glJlR5bYhcvYxSVCvjrz8sJ8K0LU9VLLwis526z
0oKF1vKZNenRD63ALZuusguN2V25Q8kZ66abxlQ6Xs0ZTuDXRVAh5AtC+E/s2PU+
FGjuelB/iW6AGldfDn87sGJctxIXz17aqkKUp8SrK5ukgK5ULUcCgNuJTSc+afCl
K1SChalfpXjuyVQe2E9arU8b8vw/qD/9bfkTMse+HGk9U6wUI127m6cuir8uBdzU
nQQHJyAPUbapv9XNaUXLuJm1c0ruiF2SDrlcwNfHQMfkF5ulgy50OTWXUhqGqiQN
/KvzNcBSyplTu4iObnudfstd8sg2ERd5OXTDc+Mcmf9Pq7vZyxeOHtgcW8h51dYC
A48IrCRjtiPD9eR1gYrSEg164ZMdp+W0mthkgq77SABDek0msXzrhCtb7BD7Cgzk
F2rmLO0pE/IMXTDVawM7XiZgjaO85pgX9Jj9/9lAxZyAPQtgX2f6M8RmfMWWrKVn
l7usYkoTHfzhO+ONu08mLMjDbrK6d3c/Ecj8xCuNUBbXO9AgvFhAm8e1lKeSCDic
vlLvYDZ9DqEdE8oQ0iiVfuc2ZTuU9CLgNeyscTFUt+SF3ZzcNcDCQ+iBPRTNs39l
/KgYTA/bQk40wqaMvqAGWzzVa9+32d1UlRPQRzzHLVM6UD5Rl0xraJCLrKAblCz4
9DlY5fYFIZxNEXRvVz3159pqrkeJUlPOfyfB1srDZqQ0c7vf2CxTvGxDPEJfM2l7
9HCOXcZkywgn8KwTR2e1MyZdRB9Zwu0A5sFDF6niAlhMC8CydOKLbptrv2Nj4mEv
uV9a5Ys4U/Z3hxDtKnYmujQC+A5uok+etlfOfs6AcisFPMBNtq//V7K7HUrL8ISd
qyLqltfIccqBZ4Pc6n41/Jzy6KJk1JSijMmC4IuBwJnGJXcAFFpHd1+n+SOEIAvF
QnSiA0sjFuTqu7PFl4l5WZ3xgtJf+JZGECI+x4jYk4BAJ7/TBseQUwNtAZeZJD/M
Je9iMkQPzxSctJteltIzP1RBP0RNVFNWqWvMYibtvTwcN0XBz8GlTurduoAbTeaG
NW4uGkXzpkzRVU/ulQuVmMp2O2GvuVxkS/3OIJrF/zUZxBHYQHn/3pzep1EglH6b
IKqOiz2f9q37l29DlVcdyvC3zQ+PwXgVLA5kzenS3bNIbTWUUlup9Kb4ZODkksL0
xKF0qn6EttsSqaWjWfjq0jzrhdsCYc0Q8V3Tej/Km7X7dLj3nQcWqRWshUW+vpzK
vdlEDp1EW2U6Pcl0gkw28DQQoIT8QUUxOT+lne8TzdmfQvsigo/tXO58mYx/UTNg
USj8WqywqhQpeEEjE5E7mPqqrSFUhKGOX/Y19mhRxVGXbz/wIqMUXKPlJStx99rj
sWe5Y0rN14ohXt1BAQCZSAG05V1wVLnI1EVe31KE3zmk8owBUKpwwbM2V7HUMgUD
PNp+gTwTqoRLS4igXDMkbm1vHVSY1Tea8ddm9jEuVsU6BaaZq3EDlXBQ7GfBAQ/F
2d8ZRHWKMJ9UwbsCyEEjR4X7qoBCghGlOV7gfQP96FWu7FsX9wiCw50s54lK8num
0an9lHtFxMLNAmOhtB1aJGnodErBwy+YWsxD1R7192tiYyLHjpkREuym985KIDzt
M9JtTJ3CisJ2pAGcvfHI/+jlEDpR2M4R5ATU1nji7UBk1Kb2fLN2YTaNEcza1+GC
XB6bKrH6/4XSoIUkKiUxQRXLC6FuCCouH1RJL5RhaZQ11jyhIB1rExMSttdASa3k
XlYhtNRN+z+LgSyg/m5NdWdzXJGTPFbqK690pGDlHxYdaJrS96VU0jjgFIp9urwS
L/sASNcReOQVNQZyGoGZ/raHPlB4QIUa9MLgOgIRSfGzbiVsNaVxKy0zObvDI6n6
8205DrPDnHb494DAMuC/GvIJHiNx92bYUTpBquB+gjtwrMA4Di4D6CLJc3/G4O9A
+ykuBnyPS25DjSqt2Jnh4qqP+g0NxkgLrgO3LSEDgKAz+8hqOTq4lnbekw7k/ixp
mz881uyVXEvSsFcEzYRH65vCxUVr1KeA1xfS4nIhGL8UB3+N3p6RSr8HALgcW2vz
LEq4460VZUXwa8m1oMcpqzCeJ+gXsu1tAd+oP94fhhaLxEt1xUvjTJGkTbxfa/Dl
oybFsxdi87ajASvWJZSl/TE9h6h0CDa0StAK8z0nhZ+5j6MqVq4SSbcRdNr1jQLP
HcUMjAHjNjWcu5eennahH4hAHEjwDfNmoCfl6+VA8m8NOzvj24nLQG7pNULWZCdC
tQ3YWftcXE4iU2qWv0BLK2MvvZN+2X8747Qc9lsF/5mnJmfDkipdBXT+LPm7efV8
Fe8LCUmbuK3WEG3WYpVZiwM51R9SwNi2gWjS/y7EOAXNMgusDnSXrZqpsc0uT5yd
G6DmHmyj10K5pYV2VCOn1/A82FUa+Nqsq7t/ptPxqLTdsp8P+xyIgbF3bRWtnReu
LEmNQ/mx/TGB5DB+AiJwpUNvD4NRMvuYvn3ML9auPVHT36nF0pDhT8V6YsJz27jy
9gbFzeiJwiEivhfa9+hn5a5r6q/pRfNT5xQvF0QswpYz5d1mw8FdO0cC52IBpJuw
uLDtLDuUyVT4EWEo1eDwMxytm4Um28cbIUFFCngSy60++f9rHCsLwPzuAUSDHwnR
0wB4T0F/G9oUXLLZV9casPPe2HhmrKnunIEA9ZgBdr9fHyqnn9v9efyHqQpf7aKg
Id6+eTtZaINJjagX2T8FxFKJd8FaOZIjmq2TkkV9EwxTJmY/N3LXoQOZDrTj8cZM
wUwgLWZMoiFqtzoVP31G1qlyHevmzBrXQLgU+UnRa5Y3bGfmROpS/6dmtpdXtvvn
B/zPAizuCihRqfBcU4q6ke58gkqmIX774xIwnQ40M7b7kOiglw1jmYGST2Lr+CJ9
gi3BkRF7iPyiy41yOSnhg3gS3y+3rTtcVVSpTIH25zXRXok5MAFoswjvDKlGzE4Y
EmHDglI3sJNSnNaGlZjAgTcK5Mp8YNIlbRe6G5C8pqqZrNKBf0i6jtZTnk1s1/+u
faK4OkbuS55bxbNG+wZg6IsWKYZacavBoY5zx1fRDBa0h+LuRTvVAk+ld2PHaU3J
ozsm9n/7aOIgd8YxGGrouCV7eDNgEY5HuoFREaaCi4uBa4CnWH/By7+szvXASwkj
VVX0tSKQ98uqvtSCr1WDDqL81bJG0jlTpfhhN5zKzBD8EOOslMAF1Mj0GnFvzeAS
yn/Gg67LogBEtac0XTdaR/ZdHj0//4SOwmfxjd0l8PHVKLQBfQIZW9/4yykTYC2f
X2Cshw+DCxDOwHKI02y83x7UyoqCP9iUycE9u+yhVHlie6xUucl1Vifu0y8mYQGr
zpd1estJk9oWDr+l/7aPWb7bEfg0YIFfMDSumrzvpoa8tDTS+zYsE/fDpVitUzIH
E/An8arf+NKKyGefY8odhb9QXG0sKatFEJnmu9w/bYKtJ/b9HsrlzIgVKg6bHqyP
oX+vUeWuB19bydHicCXiRIaYKO1+7zka7AlutXTBNU0U8XTs5egNLUNWSVIg/WeQ
Rv2D67q+VbiummwJrOWLoTYD15GLNzv5SJJsqCFzTZBCEe6jZS5Fe+Cp7oZcJ2wk
vqzPxEq6d0zOWOgPwjwVimC4St/4W2s5gAAV7rPqLGRi61qz6FtdZye9O/J9H995
Fkfsew10UGQiPhogs/ARTODtGJ0Z7SxlsX13jgC5jfQaF0c0E63/XUW7BkK/8x0k
Rr2F1xPX+Elq3a/4p/BI7hiHSXi5WNqkhsn3OheedOJhaGkYF/6v4S9nxL2nyGHU
bbttJKzFI25tLYga/ut3fTSp7fckSeix/E5bxjOnWo7+eSJnjN+YwWcta6E2jw9i
ONSYHOpQjy0LRWvmylNKumWmlva7ZZDC8N1wT0dMH4iM0W0pV1D0E15CKH5Nh7K6
zG9tmTwY2YLxYcHDVvsu5Y+2lZaRLDGTZSbDziWEUKwia4YyJQN614gO/dBNFm8A
p3GvKwd1WUB2b1+H/CaL//+ziQiDrbfSJ4UEuv3kltLiMEOFK11iI9eEY4Hx95A3
QAvmBhxNaL0D8tnmrLb4mUBtun/O4bRQnXQBbiQ5PEkFtR+451xYRS3K6sP+geBm
6K23yM1zamOL4ztylwp6ua74dLBF83M3k1G0maRfX0U6CM+xA2u/OoOE+F0MWeTq
lABPMCx7OinzFK/XVnhTiC6thRkYL+qRzeuIbIdb1GcTM0tpLXcXCHLxhUuma+lC
W4upQvjzuEDNbt3on81PZuKssbKiIcvYW5wUOD7J07MIjybRhkfNupW5yc6NIVY+
6KHfJoFFePqe9KPQkaqTxyItzsHLelF1WdCqN8iHI9eJMmXJbb70WrfBvpqB5vgq
+eOM7a4okw7alpj9U/OuPOzmL83uRQayE1AgcY3BJ/0o1+g2kCYoyRP7yAdwrcbO
OsKg0kEglK7bvsOP5FRAbUSI3Upi/uNxkQeEWyaVOiAp++k4auL3oas6DFLZoR/5
R+yAPtEbatF5MM3v6nDJgNQ4yuXBwBXklFjLGTVPLZ3eMgQdveFPkttEj5dTTS/G
blKulCyWf1dZSvRS4t7m2D/kDvXEB2tbDL0pV9EwoUVt4xLoVjK8TTPpmQqBCXTX
PHjqIfflRnb+aOyGYi3RmwP6ai3EyZcw6ptaKFKgDW9Oh2wbMwB22WJQJl/lwgTn
2Kv/0uSLVoYJc2SXCE516JaUAo0XLuPwJthiCIzgeKjp0JtF1NthXUDANNka8/CN
mP4/sJQVI1HjlYQmQ2l1Rynd1rsINY69KV+RB0pxuXx4r50nmFh5iqu9oaWULjuO
jPy10EwsiJFWXi2W2DFxQanYqd7G9kSXf9X8XAKjYHR/WFIaYNL55v17z0hYuGIf
DDHspVJcvjFsc7cu9gWDM1+4RLhZmZJOXku88eHzSojPoqLt8K3iSZA3v705xfvF
Q1c1j2WqYksGvK8QDZQb92vfqOTIMcWcmvSxAOPcEBhIE8YTv3MoI4oV29DJ/6jh
8RjtcOm0e6FuOAFrXIQwj96h/SHj6CmrhFk/PBt+YIeoTs+Mla2bPMDSnE4y442o
kRCt6KNJ9NWpC+vvX6+b7VEW8seZk4o6g0USsw+5f/05wFibCQBz7mHnFxinfPa+
YCqr6hFs6uPY+jBcIC2aXzkX2X1n/jAo3EM4gQxI0G/LlFXDR5a624pgS4MCsOYL
xVRTlfsdr7pjNCuM3FVhIlWb4RgKtvamT+ceILO+sswdYyg8AnBu8ze5CZ/8NVRn
PxuuPz9Xld+xgnYG5/gNKq3KtK9+pQlwEjKJKPB72BuZj998OmueG9bglTwmaLk5
f2gWcVUD7awRe2OC3C8Mt7pL7hbicXjlnadG3XaDVdRmNag647q4PK2qJ8tbfmme
yHri7NdUqt1eLbod1gmIf9ZhxURpuEj2khD8QsRK2N9HlD65fG+R4QkCHkqp2843
fP9+afbMM9guD2YwplVj4A2XbPXE/OTl0dLWcEyZa+k5eXEj46DZG/+jNs9m20Ub
lSycc1qiQKZGnmB67bsgO/zZK4+LPrIWDg5X8rTziUeiqINBrFyhUePvA2yP5GfR
WO3nXpFYqpIZcKYTh0CiW/NgDl8Dcg4etLfOgpFyklBAEcjThiSHAkotC/psXrCK
Bsvz86OoXJsZd2KTabYTM9P992yg/aV+G+hXwPI5HwSABZSSB9qxYaq095k+8xfD
nonEU2hsSNndQtTA548CFGMGlDDkqlUj9IN5D9sm083alHSO56aQzYL40GejZCGI
s+ySyU19AZpJ7n5Esc3i4an3mn+XEjUDkWyaM8FfSTfVB3ZCwvNs7bha48P7s3wq
gTM1YGO07ndu4b9riia2W4mfiFPhyCo9BvLk/oxqg+ETgLz9ZS2QFdok3WNfwMPi
HbXo+FzaB74Q5OaVlWGRbnimlkDcyMMuaXlgE5oRx0BDbjrHfr5sLaYvrBJisd9p
y5bt1O8mFYsuZNaHP6plJZs//osxvWTl7deL7jyNjZU/FmHLYgh7eym78qZVfpJh
FMxfXvipi73vGXUZpM1wW7SHkM9ZB8gI4mI8AjNXgby9h42xvRpyDh/+nYWtGugO
6SGNP1nK7Vjr+FF96MqC/rnV2I/wkC4tbPool6bNcK3RrweItOLKmRGMmshhwCm+
CTdm3sH9Rqn8o8kDqeVUgzdnLpwwJmo4/UetomqiTWY7yYWgZ2F+nbfd9TdAxlCk
NmRRRF+HyFePm+Y5lG4sIKvj/v7pg+8v7MkK8VkyDpI80S+X9C6ekeFUCMlFPW/W
dORHjKpb0rF3X3YilAE9w5VF62Qe4DrPYDyc0ESE+UQ7oWF4l32QzaiBfolA77r3
cQ0sFqU0IhnAt98eWlc6bRHedS9y/BnG9zPi/pAv5kK5SCY2YvXGw2AREY1X2nDT
`protect END_PROTECTED
