`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kMLDivLhB5tNaR1yBIZkC/Z1cOZxlwGzsSP/8obOQcGk1S//1IQaGPoSe4hO69fr
5NrZVu3L1T8whcssWQ8A09eVPSLK3SJb5DMCllb+Sj+IlO++baiLGDDRusUpwsoI
amFMc5mPsFjc/hs6cI58oIUA9x5IOn8tlWwEeD9piWzypStQXqyQGXmHNqlUS9+o
WVAbbW2A7lxPyj65d/o+kPS/XBrOvqtExgHdxgVd+ZUFvtSBHuadGP9tkLRj6M3A
bzHGunhRXjGRJF1F/0nq64bMF/hFX+j/fJUMPiiRblI6O6u8elTqKgKDvfjt4PrE
kW5wQiDvhQR/evTWzaottYQN6CbQVKUEPvVzeKmAqPlI2QmZu3yFcj7Bgvn+Z3/7
03lgFyGa4M5h3TN6iU81OfookWz4OS2eH8vedsGPJY8lNHdyGaTMmcCm5Ji5wF2h
BQwLqq4O5b9dQFZ8S5TMQUM8XLq7qbti+2bR67nEilHPypSUXThDeIY+u1lZswII
oPEsTOTm7Q4seYWTNZBNE/A9m+JZCHfOEgS8xjt+miqucl2Ywcy8mML0N/ozZLv2
V3GYuC1hd4MTnF0mf9W+JObYeQJwlxuo3yKYREckg+uwfFK2bkmqcZyKiypJOzuc
Wsc04QHj8SDmsMCsnBy01gEbL6ywrXr0F+BFNYslG5+ZZ3ol7BbJXju/9iwMd0rY
jDXHEOws/uAtWkRRqwCg7wDPztH1SqODdh/Xi5NsgVAdPqFvgvgZfsGzWcBDyRFO
j2Br4DSSsqE4bA9Y3tsOiBV19GMlWMWF+sX6xtPt5mLLqB2woWjNhhceR4fnN5Gu
TX2agpMFCiIplPzW0JCYVLLyPBdaJ60BvS2hbQHSGWq9kpbogIJTIu8Z+Xn/GB8Y
dnIKc0UAY9tZm0YpEKK30xqKsxK4khpTpJvIsmWuOqhpwEwGWiW46dv80tEZRGZu
bPNh8YTF8bMVo8pr3fFqjEojM7icatMEeYQ3iQsgxAI7pIyyXEjrjglQ8TKGvYH9
7wegKsJr/jTPrebDLGVqHxYZYtKyy8OTmIWEJLVwrAnxeDcaRVfE4t3onoQBR6R9
L7N/ozGvvtOmO+Soj/U4VFA4h54IL7Dj3RiMQgb4ZqpxlxYcDxxDYDYcbD+2RL8D
1CfJchGyAQzydILIIQTKlghheBT9Wuv8FufvOhjkJZueJnAiTSNUh8fkTtYbW/k0
o+DFD778GED8pvb2GnCafnY2a/Js/SrvNojL7b/T70fvsM1o/NSgvstTGgxgwGr4
1rpqVCZGkJtPr2MDQ69zMmx9S+p84FtYf1haZc6g18KdE10S7GkAac8GiO6f+Mfj
7RHVK9yUB8V7ZUw6pIYdB1l6+Iv/zKUvihPW3bil9q1IC22pUFK/LBwMZlcj0Xeb
vgyiaQoVjKIti8rp2C5IvekX3brI5ZdaUVpyw9IQTojRnASIN+auIb99O5eWUkpT
BmBOhmMxbMHcOQGBsPfTQRyk8GMpBEwPrsQdF4H7r/U=
`protect END_PROTECTED
