`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
seOUzr1NOLu47Dk4IxtLjv9a6xfZAewW3G1ZRuznuSBn4AWCveZAWZFZV9VAlgw8
ZeTAfr3IiIOT6Pt8BihYt9dbW29SQqvk/9rMqjZQvLW/E1IjfH0na1I9dxW7fuMC
BtCRRplMrFaDpo1szGDpzEQuRZgmnL+qiyt8eNzYMxZ166w5UgF/Hz2HLpFDlENj
shV34y1yRbBMsmhiFzdc/s4sfa/jebQuF2Fs91iDHEgQnxvflqDlsJY+d/9Xw7Pe
SFZ35pw6FDA6eCmWFH1+cfON0AqSgLVAhjGBRYimX/gHObwU/iHP2/v+jrtXgUzq
QXXBLaHzAZfWJ9fUxzKQsqjaIbdoh8OdlF0MQs7ilGnoOE5VQ/jqu5P855MiLOBs
pCr+n1P5kpRcoXr88c2XZ6KrkBRmjrAi2d4Zqgd1UxHQQuEm/Jqx2pdux7J31WA+
Eiqn/baRPie8410eBySVmRAAqswP5v6UvwL+JkwExwkUvc3U92xoA+FfxSNU8x+o
m+HblKHrmoVil/N9zBRcS0iqAJD9CyiXYnixwrSlCIUltvwiM7XptJG2qAVGNpGj
e1LDlYU0Rd5/Bq9wkGwHa7MXpECMOnBT3ViEE5+4BCkm2sCOesu9WpGK7Ua49jo5
4MAHcEU3roZJuB592VBhv+XfI+bMnviN57AN5a5aaMK5jfJBkPE01bzc6ar1bH2e
SRyiP1OV5wycO4k1rpxm7YyhrLwKQc9j7B/wuyMlEzt5oqVy4IpL/tGguynKN1MR
4iQ3lA0yzWo379WBt552U0F+ZmmMJb0s2tjqEGkMSvnYHhWpGEbbLmeSeHe6KBVP
ccO26N1Cppgy3i6qtvWsG9Q63nceN9a2GbjlP/Jmbvne/J1e1wSB3cF4pN84Mu37
pemy50FCCvy0g0GcqcJ3vzc7ts+uMMHgKgD1Tee0wwNtFJQSx5fb4EbTYLQnUDxv
PRa0qEEKe3OcYv4OVR+sF5SWZWwHtMfwmpFj0H5TJB5wpUCHKHCLFrothLLFyPSf
oK7/b9/q7KqCT/930Nt7xNWZPIZvNmP5/qoLHGriuMzpZCuPSKppT1aYaECMaFZJ
xw7eJbd0ZXnlu70iVgLEYnyqeS+kiZGAibsBxTcDZFmPBsaqJ0ZD0hABX9b1DqQr
/M09IBDrZ3vxcZxKm+vQD6f3UWZQ8uIfs9pA59gbhHN4LqMLdZ05tCFyBYsOcSQb
cok9e95D+uq6jrorJHxvvA==
`protect END_PROTECTED
