`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3vvsCJiT9tyA63+Xg/uv2aT0vXdt88ZUAGLYnyZYJQbF5cJhuvMU3iI9YKN9Co0
3V0DNdkkDhCI6k3tBbR1lWasFyrNRz+iLcBSIRPEXQdDgOGAyUA0zbB4Q5jfCgz7
WEFBamxyOiff+Wkfs95lCxzm1jl+7L05iQ9KkMWqoZ8PqoCQ/egzcegVzbaft0ws
0EoAKrulcVXesJcwatMRIf7lRAhuWUKDwKYW99Ss/IVN3ZM/b5blX2xtZdxRSU54
qstIMfYmCioZ2qZamghj/OtPfu0pXD2WK4CO9WiOzoJv0CNyHgsFb6qTTNhhm2le
xANK5N29KzwYNDKikVPiKossPFE0DhOkdMjt77bO6PtIVU/uAb+2TyiiowFH8+41
n3qcws7pl9R7N7KPsgvDFxxRsKpZ3u7JC3znM6N+5H0JmeiELQUi8GuEiSY8oCXA
FD7yD2hvL6AbiTLQGzSTL48h2gmBlu+CKLWECfVR8Qq3iKH0hocmWRWd0wWuAbeF
O9lf0c8rfSeX+ec9VvUNiEH/7ghuASRkNdZylW4hrT62jCGS825xhcCbCfAhnZx6
l+tpwiensE18Yz/KXhVHR+uJvYUaxyM6XE3cqJ3EDV4lods9hVGv9ofcqa2bepAi
LFXcP62kvJU45jkzP+l9UuIwJlsjujk7JWy16NL22kmWgggmnBpisqfvX60t1VFR
`protect END_PROTECTED
