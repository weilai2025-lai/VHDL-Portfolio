`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUg0wW3zw84wzUSWRStY1A1T1PpW/zHzou5fbkMt3TlsjymrWt9zwszalsFzqYOU
gNOz9gyUy73JR5KUiMSSllNt8T+/7IgIT6ObGqWK7uidezCZHXzIRjJNZ5B7MrKx
bDTcY+f11pvIrkoVfopsxE5Bz+dTDszMP75reOC1r5knwnLOBYEFOYsaYmWT6FOF
lge/xfcYhhNWYZgBqZKEsCfkt8tvmprpZ9ElyjK9bQBqg72R30RuQY8tmWJCe3B4
LW8Yiw7h1sSj2jHRBJ8UuIfqM/gXsg+VZHs0l3m0iyiR4JoMuTHnOFFFggadWIXH
HBpWaMLltppuh+TTX5KpWqKaLHhFsaAmwKCmmiIHgRcXWqP+T/I4K2oDknU5j+xz
bd5xU9NgJK49RdZ2jhfOdf/Au/x80wGoStpoEPRKIlu3YEmi9nPSxFCVXWXZ/goU
ToMFi8Te9AVtpSp9WtabZ8YAfF/hZh8b5dCqQTRqDcHApiVLuElpSnuAp1X/qJsp
MVV7jMUelzKEqmnoJhoxTl7YGbTiVXv/gJC3sckQ386999ZzTTf2r7BjOt5QvYCE
jJNK1E1r/tZ2ds1pIzfCBJBX37S7JoB9D5G1HxRgUMYa3hIHFluSFZb2Gp75S00k
ua9p6v3LlKMjTmsFfNhmadBNpE7CXmgnsQFDuCm3P+BS3olcuzW1PDq16bM4oL/F
Y0f/aqMXqOeV3NbQ860qbZvwVkgkRBUtmQp+y8edBnLSsL0HGqV/NXImdFlqIP5b
r81AJRAcjc5CXiDRE1knJuYTwuCoeslde3CeJivH5+a6d1UMh0dA+zZ/OhrFsJWX
KrEHFRb/Nf2kuv6GUEvqJriJ78/+I242l/N3fHjIEvD40XBz89osnLCf/8rTV1sm
z8xMRt6mLBlig/9xGUCM0MbkCW9E4Y8AocZTGvzo1zY64aOjL3QTdzRZUiK4Zhnz
gcX3Q/hxR+MWRFVO0ZKX/Zo+8tolK0nC+CNoOo+/AZZSeU5l8TihHupntwjwRa2w
RoUmMQMrc6kXkKNYj1UhJSIQFb6TZm9EngQpllHwpa9RlfG4XfI633OIenCpXn7D
nTcaQYfO6vp1Zwjtz9wDDLZYKOF1tBFJZ881D0tDpx+sFORpop81aBkdGpcKbWqC
Jfxqi4XiXe25JrfpXmWbQ4Nmfp7he9ufQJ2RrxjbuEXNke+z80mJQSbP6vbgoH93
sN/Eg1jgmU42vLd1ywZwnNRL24qal5LLdroDnYEeYJ3VIx5qZTDBmErKncv23YUu
`protect END_PROTECTED
