`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1IYWKw8wjGgGuDiFHhstW3e39wbfaw8VBQ1CeybBCbSPZruAJYvFOio3dZt7O5r0
s0+T5X+DzZZ33x1PBAIqg0pLC2Vy2W5byvKBzX868aGkoB63JwujskKoeU2j+4Ni
Qqs12Ayzh4EQc32zmkUhXhJMPtNhLjNHBejdPBxCnm/kkLS16Ja3Xdl9vQJE3ZK/
zSJvWqMnlpsOthFV4+Syt1TKGVWg+8elASNhntUWC83fIzob/7VykgNHKXhfRTAd
lMH6pSui0mqEpQuADMA6lQQpsH+yuMvWWWx/BBEzuCfFyvn+YEp09yPkBU7ZYW0g
jTvmklHlfyRlEBl8pt7zlYX29dY0E3iRSdYE0qDCkuh4dATmWZs59Rs45wsj1R1j
1K8g0OAfhyXoPAFqms5j47JtMrjQuHAw9o1ZK6A0scSSIlYCbJPPDACOGAVWCZtn
trIDT9t2ERZaYGo1J/YHtDj306HsmO3JC+q3U2gnScRo5a6wv4cSnlQLD3yybQ1a
eCyAKU7XB0met4OdWXEpmqr4QSlGgyXQY1DkuKYMXYpQXUcBVmd28Qs61JKgqpft
R9cWU7GAKdfD6X1N+0UaRH/DYLVM5I7X9BlGqmH9BcPGUN8BOuEfXVyz7f4OpMMI
8Zvg4pTY9kgoytmKOsFjtCFxwELH7m1/kf3MlD8x1j51eb7OWqgUO5Q9Z/uxbDVw
BfmLbJP77HYg6ROEyAuHQ9GaOuqWADETGSGY3Fh9cOHF5C93TJrciwUe2mvB0HEu
Y5/V7Ewo8ZUfQ44BE3TUxOWoZO/o7zXM8WaWt7D8SmW2vT+ANuAp0AV3XAaCBq3I
L1eYtigiQZh4FP+msEGaTdP6DglZT0A78L/HQcu+niyYYj2BFR8g96UUxhW97Yj6
qxHyNbXuc5ZUhNcqre+XQNFdniZ0cGnONvy81Egk3TAFOOev+94bC960j2YiUA7c
i1lsIfKkTq+KfRsgeTlm2rTaKyRAMjqpuDbxklXdPMf0Y/rEQKp6h4o0jpUPmKQW
m2Osgdb/swWerZmM9u0hyWhCePuf+6X+lJ92ieOWiRoAWiepvLs+ddXaKPdinCvJ
3vLF/kNkbkSnYDSVODvmB+ffeQDbvJsfhGcnWDgRObZWeRKlZedGSD00pd1voAS2
uYPfMG2WKGZddjt7UGWIL8hvHLckCRwo7xaskIF2/icCAWlWjxXwylWLvkj5CecS
jWEg2O439GfH3Fv5IauIbdRwh+tAodl/YaPiTjAN+pCy95goXz1Gc3i1m0GQZVOO
O23mRbRSekOy4n8A9X40qE79GY1l570Cm7qouho+BYRMpCyLxbgZSTJD+yiL+oLE
MiK6aUZdnrO0cCyaTcYIZjL9KPDccjDd/wZMR6+dLQz5zVxvAjROUmJwzSsvxf9R
x41uPreEjUvKflVn6OxiSFqYDB8GdBGQnMd3JVKDjjZqPZos+fQKVZuZFNzI9jN5
1XIfXpXQiVw9+rCjig9eZRry6CsfMuTvobdXNaKZpimrqfLjsQkQ+VXKzNWxJZYh
zdQgmeyQT8N/S5pp7VjAcDmM3TgBfvKhJhWMc1R+C34BMEzjUKILDe+srF0Qkn5Q
1WKdabPZAqjFmlyvAIyb9kjGR8JQ7qq0VA8WKhDFY2La5MaKKKGQ6d6aeVaDRnMp
iFmrj1W0yCZU3C/CB9r4eiYatDg6yfHkLCW5tNUGsx3054z9E3GksmoqvWsmZujV
lk/KA4+eXHhwgFrGkIboYOMPdT14bCaebzqXwKHW7ZDsL68EoXVrfma8Ij8DC2Rp
NNGkJyzaVvBFx3amw8smEUXxapijlISY9fIUUqJJ6aSgnqyMoGTW+5givza+NmiD
nNwqipvvH+r3RRJxqCS65401ygIM3fdGz2lv0NyvQ7ufo3409hKT4XSjWO8mK3xP
Mrv4695yS5tPJj1kHZfffID/qS1CtP7iVse3n4ZsPQR97PMuMhjYJXFXvluLhX+B
KzW0N3+O61vZ7/Li/faIcn7mdRN5CgAyH/htMqZQLS2ZpmXRGkm/pbSyoj+zlD4k
p2sJYSWsbYnjeSjRUGAJ/RUi/obn3T6uvIqX9FNQnjoPGCByXaG39Qow+TMbefQz
DtQ5ZnUeheBn4q9KloCZLMxSDepryvr7pwLHIzhRC3ea2M2gnQ3M0+NwV6usMI6Z
RWKCmDEkXko6OKAwFbOCZjkfyOeBaRnvgQJZWowd7N0PwbVHSdLzeEFJst0TiXW2
EYiL2wD9qJf3I7mEnrFI9Xsx4HGaiKPRcFq4zaUo9R8maZrAGAAKfmSXriF9k4gW
W+itLNt1J1MOB+HCjelALtAR5Y4tvuTJTLr/4Lh6Ly5aSqg3WbpB0yXUyhJyE6rj
0Uh+X+xhyyEY+kljoYfq8z7SWJbvlkGEcNEo0KfwDiDSJq8dOe4PhemX4/HhEQIA
7UFeAlCtkcAH0ux5DwbYjo85zOXEaJ+3ir6GXlVJToEFCqsMFxRPts5bamcRcQa5
ux6kGdET6doIr/uyCuJLpYFrhjwdEu2ryndElmEIoYaQnw1EuGGwfIIIC1MgxAhV
vhXqjUpZGZ4vFMxZ7/ytg3twDp33zo+Ke09/zg8HNFl0mkkYbkeWwclbFJezM3xT
YXk9tbJtrEL3Lo/EhLsoEWeihW5SHkBUeiInp4kfbQ2EJzrYdAaxubPBcBrfDxPz
3uQnwzc8164N1aeNu8at03DwojspmbasrEwo8DM3A5KYdE9suEYAOxCWQUFVk7kq
zIUbX+as4NbkK7waTt7RSbSuOcOr233UMNtR7mkCgZI72Cg9YUBiclEYRAQSMdMz
ATYCdC0sgMpmwc31aFDWNo3PpAkWvHQLoOIuuRgoJe1ODO8sonU1rEZLWaQElrdI
qLZ07rVInF5D/cXo/mhNBCIxrtH8QETzsl1tm1kjncAYB+noJREtTgxlL/tRvUA4
nQoPMCjkFoctGx5OHUobBcQglDYJWHEILg5os2lk58VyayJmImp2wUnQLh3JzA6O
BeSw5LcKAMZGg8BUVDPQ3pUDDaGAwmEQ3mRgAfCa6+Yim/7LJEBZRQaDTHm2aja+
HT2k9eXhqAxQz8oTTAqdAnLzRjgvPgJgnQg7UykFq0uHaErEqvFlITWUZh2/31Pt
a2TvWduDnwpY++25IMWC3TSNgOGuCsIEKJyn57Tw1S5kFtyWtArDpMv2tt/QVbCh
koMK/Obs+WGlHCRYxcvcHSEleMilEzYuSRaNV32eac07EMpjcoeD/NeL8MhQApMq
QjpRgonRTcbFuh4GNAmJMZ5TmbrTzSANVAtyvEClKx1m/RlqjStWrB5Y6xVXKpJ9
tWHBiTqDECmS1Pg2fZFF8KKSnDtmTaUZH3uoMFFAxa8i2144wlQnrYSuJEc9A8uG
YOphv3H2Fa6TkHUo3Ar27uDOZL1W20jAUdHX4qgPdu5hPSmVIo64mNFwVLL+Fj9t
46hHslqRnZzveQsvy1JHS8DuXF+bJ7BlTmqtJDrsxR0rtjbvLjkkTLHzpMq04Ijf
+kZ6sICcW1DScyuiu1Mxitdc4UQ49V8kVqCiT5qnTJsbw4XCb8T0kLisG5VFhzfs
nDWC6Sf4lZX6Gdcu1zMQyRr9zH1MJgWT8MKz+tt3WF6v/yZPudGULx20ci5RPBeO
kRsfT9hUprwd29RKFVlp/k9lVTPltHkqPQeyKW2STsPUl3OQRiMukr9aHOP7V01G
NlUcl5atRZQ5DyOHVyebHUrXQvSNxkbsmFxtZ118N+DEEX7/9BMLIfvtA1cESksc
WNba7aA4iRE3fK9+sApPqxyhOsJLpn/oP3vJQw7bgPl/qPalvFhUZmPC2DqKkH9K
lFz7n6ubEALJL+zReA6x1ZW+OEfT90F1FhZ7k/nnYaXorrGD2AaMwUxO/LvnIvJ5
wuwKAnu/y2bt3dDRATXclpUbJusPCeavRaPCuYE2lQqrHTNcYQ8Fc9foLQZGD8s+
aMJaYCX0jiPPhIQZdzHcuMgMofvaTl0rO3PMnJ/PqGngijhKQAUE0uYH8Vw52DE/
p/upaZzRxXF/vqu2RFsSYUNUu+xUJGQevSYxAkrjL7egCBbC0ZYpjl7AYRZYTIew
nh+MF7lD8S1Vp32TTBJVMnPautXPZ+n3w9BcffMtx2VdOyCaGE+bnsF/IOzquDXl
CLX8AupyuHMyFGRMpsE+3S8VJ1PDNVjVQHQensQLIep7yDbZadPhkKP07lW4Px2f
rL/SQ1N+q5zJ90gc6c6wyd5GMIX5CPs3MYfPki5o+TCZSgG5yWgIdXaHtPsYY+WV
QernUIt8kZotgBzlUubSfzlaicJr/JACVSs7trOzeQ+siW5P6kOw7Wk0n48B6yUi
iJxFV86nKIGW/1pnbukYioIXYykeOtZtgFCSbmQFkia7WrZX75bAJY9yUHPT2e91
+eTs4TfHeAg2yQ4UZqWvTV2cPKPxdDm30UEucLEVYgGwKGUDywmL7imFn2FBwv2s
Ya+bV4qVOp5lhXOZe3KAIMZu5jDNE4VnThq+2OZ89Zebt86LUXw3TUhrW36b+1/L
9SkSAWPhlx0R776Z28BkmVt8nLlvil2iBACFbf6++v5yJEmfT2ry57LABnvD2RHF
VpN4zCFhA4CjqNr1w7KCUWoDOrLPlxHli9D8w66rzfRcg7M3OIFiCgU/V2lZLZyK
15cfgjDAh7DOWf32AcOsl70KpjUMmc6Al4loqYkKUL45CnMrVmnSLr/DgybguuEr
/WxC1BoTE2QsdcbdRlzLef8RSffMgXZyLwikhBuq0r+jphZsb9LeePS9RcqAowhN
+bX2/ypLKnbN/16RCnAyK5YlZXw2kK/d62QLLtBuUf9l3+p23hrwzYGNj9GNxf65
jB7QIOOGRlHGn2V1DHDf9qFOqMu6FPTZawTdP98L1MoMfI8Nlg/4GPuKjJxqzIMW
Zu1KsuH/rCoGqgFyL0m2xs+g+v9FHcCUhsWBs3A33skR9zpUenzm2wfhjBXivtk8
Uo68nl3k9kL6nBvMft0ymSiqCcCJwrKe/OB56Oey+V4wzjX2M7vVg9DQrAgSQ/fM
fU+osp+V6FPK4Qf9Sok1TmwsMlQvWGat6lcxtTmKGaxoR1wbpD2TosvO8LiPTKIw
0Hea4kA+4x/Gq//6qpzCdLW6QzLULtsaKAD8ArEI3GVGAKABEnnadb9+vQqB+J+5
nSnfnSHKri77QBYBZrwobY0YBJopbgbXwxyqSdQGRJFSggB+LGOeGoedySHc/dta
ba79Lqe6f7shn9bSkPOkynCHIBm+AB66UnVTu6x80XDfo//Otg1hHYZnQln4zobq
54v6UTYNz5um0rru3YBid1H7g2hT3Dfw/WwTJRXbjRFkWbmcJVcVO+nPgqcIUjUh
/QQH8y0YjvTla4ouPZCPg7pD6ecFWJgWiKy3DB6Gz9Xg38vffjJnVUcbVpMwL6wt
L0OSXOBpTF0wcnPFK1M+G4VP8Q5/YkE4jGcPyueX5njsGthBAPZHEUkST2v2yIiM
K7cwAfTOC6oI6Cvhubiv0LHxB3EWf0LXYdmwo4EOwu9NMzQphaLAagC1bxyKdIOn
cnWsE2lNbxO8A0FFrwb3O/syPzCxrioTm1WqMxO9OcMNa9+9iYpgfpplexa1SFYv
/2UUiUNTeEHS4m8iElpP6kekdgNdMhAsZXgQomEBQ7GXez1xv6FyFT//mN6lwsSE
jUxKYCQGLy9CRhatfDKqoUb5PlXKATCbZsdxT4J0mCw3C6UGosyPavdbRI0cvHxJ
SnAQdKxCEUmkD7lMl7DM046S6IRZbdJVwQAwjgpyEph0m3qRITt7IkZrTreOGyCb
x5uYBrcH2+Mus6/iJDpRJgbSCI+eYbqiX9Diijx4vjDedyJfq+75olR+PgNbsv54
81H9owSZmLIU3j4lY/dbTIyQNDAoF/Y5sEIqFgTZ3gYS2GFaAWr3w3/PziJZb801
wrbn6Yfatg4A4wr0HtU70W5Ixi+tNY5TH3Dmtt8z3fDf+LL9fg+9FgoXGGfrGabd
wlbtBMtWp6sGYR9VzrcWtG/BICAnKVY2twK4/jaPWlgEOTUwURxWiw+FdghKqsBH
qNj2kZHsgDLTXAiRUwEC+ypCEOnp/V1hZXY1twnd86UH9iCuWVc18G41vq0H9wvE
lQBtWR5ogwGd2m0s20jLF6AMu5r7BtBB+BYnvxZwBZ2Qjbe8QZCxTAMLjSdn1lyS
ZGid9/jOP46mD6obbw+ndKCmUAGyK4AjXdZOmgS37UsLE+ml/gOjMHaD28IGHeSw
I+APVLDsgTno53AjCawuwTIIeXYIgmbCcLgKh5/nhSvn/5XUn+WTnmyxlQ1tI/hE
pHc39OAHuOG1KJgzAyYdAWlpDOI29a1+kYdBJYoHXH83xeFZa0my4CEIlAhhfzt/
vXXGWvPmVsz6jLrCSigrZII8hs8XEYVeA1Iz1SOV46HjKj7fEFnQNSyiDb8e166s
LghWJDe6PKgnrjpXjtQaMORmr13DJVRw7wi81lG/Poj6fzF2+RX8iZYTmHGRp2QD
p1L0UStlt18cNm8VpWuVbU7mcbmxTv588OVwxVfAyxUATM9zX9i6428MDdeX6AA9
GoKL+b/H6imlLyceoQ+uTOblSJIRSg7nmCkgfItknegmXviVkj7M+SMycjAuVFyA
5vE1TPRStpNUF2nBsQS8n5rboQ+b6c9AwW4V6XM5cmWBR+Lyxxqn8zB5diI9MSpZ
S9euHBclqDM75CSZmlFdcJsNmGMdgY/uYLl66E1IQtIIzMOW464D9KdMgcL2KUeu
VM88nFOowttuL97/xJbbO0Kbo2hcq3kC78mbhb6J+JyCmOTGS3pWQyR+FPO4Lt+W
s7BZ6dChPhv0rj5tEZ4bnSdHO/88Ztucfl1exAHwGTDadKt0QYHc3NEfxJOZ7oJ4
6xhxAqZOFCt6s2BbHhcL9WAB8Lz8B0rvdw9SnoXdfCGYjt/tCTJ/ljPBWfk0D4yQ
AntUdHpjBkWqMthhTRIeyTm7hvY3Ox+HEUGqruCOlLxC8PwyiUkhlAAelgwXZ7bF
3IICY/iOEaJTv8c+uFMTxkztfXyBrWs2H8KO4hhebwUe7TSSbjizIdfR2ysCpvJK
BN3BzOrYH3dyzuW4zbBR1/LGTWNivMxW6l5tFH0pJFUVun7oagv3XBlRa2yCKsn5
l/BGBgFloioYspUgKTwJWVK7ykqBqV8qx3cIDZfMA7o4jqsx2ACX3aLTmrytGR7V
N5CglO4xuzWEntZNIYnwt45mIniE5BlMMBNNIAGB/jf74mugtTAG/aN27FFtAMW3
9236BQxUIkmM47P9ecd0ixZaHdEEKZdYOZozvevu7JrDz38j26kV7zOUT7TDcc7t
8sxeZNZomg4Cbwjh0gVZtoC/Mhkk+OIs063jmq1gz2Uj42W0Q4ejphIpN7ezRJ5w
jJch1LpI2RKh2Mc8S1n2dyH8F0gQgJebxIzYNlnWLP5stZzMsbeIkZAVIM3RAWBm
1K9qy1l6gk9WPhI43B4vddBrNXzGGArDG55ENpYsI8TBw+lbfe1515INvWH/RQQf
LFhsrI8JwskMjIDR2sbQa8qw0q95z7EWTCpzerXiXu8IigfS/SvFWoKzuNJdSy+N
+mpMGSjl7rmJVSsx4qw53e1IXrxM1qYO+fa8/Jy7qmKdZkrveoV4sFy7yM0TrwMZ
nKy6MgXkvB5DiuXHQLyj1gzmv8capVCsFrGHeS05bqbsenjiBcF1jLNkJ3tGGR88
+3TH0XmNmQtyflHJ3O5NUs58Z4q63JJjZPrgaZeJAqwInDLjHjmznxvGVjbSyjK8
o3/XmT5pr4GVP4RjOebn1PWQ8ALC/8ikVy1bBs8f4JSS4yQxXULQN3XcQFNADLA4
FQC6rBkB3DMRkQMaPpOaJqVsE4H7m5d1GIb2wtDKOjcSflQ2UjVQYGmCM5oicLh0
4QSuI226558o8P1G1ZMM0ZJPRkNCvhAIWq6F69cLry2ujTqNl6hq5jd+S8THLbmN
4M4Exv81rFeHdJI2mSL/sluqfGDp2uBxyQaOAI+ESII+J3k9/TlLfQb4GUureakr
5wMyp9xrNdtGL/4kXvMnH4PvGemOgNH7287Q+FJ8PGe9QEnpWCTbp2SqVLQKQiLU
OIRlVT2NeJ6v/Yov+YXcGjItO/zj5XTFit3NjCzoKkI1RgoOBhFw+nvHqIjZonzC
zaAUfSwat4s4PwleftUdnMxNyTqrgAUcsEh9FhNko6sVvgDnMt+ufkeEyh+A+gmj
24FUnCcxRs3s8yr3foimNrgFSYTT2vIPx+odeljubT3fq7Bok1i/EOuVqnzEHXci
c8osc2E0dxNPiH3keNiddis27UQiwHqMW8/AxBq6DXT3iBrZp1Iqwv1Qeyt8BNa4
rWRhZ+nPvAR36iEgHTuV9tmbIwamM/S+8yt1o/U07hqJqI9kq0fmclQpBQM0ckbD
4jofjBZraX3RoRJInHc3FasEGKcY/Zr69EMCt8JIHir7i1qgQUlA5EVNfkcX9fnU
PS4cA53e/dIDFjEIDE/RRbMzf9CjVzHQ/XKmmaAaXIO04pNlKEwG9C3aaIpd4BA+
2hm/jKl0T+ulQ6MKyIJJ0lysX+ldgfXVnAmfuKOUo9jVhN+CmRSR7NpBafXztkyo
zbjOcfoYBAGen5A9kUo6hKWEC3/tPENnPRvKkCNSZi5SupvrxEWCrRF4gyUQZMBK
XF00EJgnX9QTu+ED8VdGu48RiI+V/bM5fGmiePgA+0A4+B6r25ehc3wQYEbkDSj6
WdgVowJfNVIxJ/2hUKgvBp9PD1bttCRvem70xHGVUP31iSglBDRRVhBGlQgdHuH+
iVoMuZOvoqy7rZkSUxmSBbbECY+ZGxrsBbqSGg1fM/hvcOLYmB1+JwSxcCJEVjdw
vaJjK7JFhbqfuRpWN4BQJCWzmkglAQSXdC6XEgClLzgbsoGt/LUxgtRblGx1yMdf
OXnxqm2g/KcKX9NmeJoiH5UZYz5JD6Zk+GQeWwL8O3asOOctWtz4wyTmwMMaMQVe
lxDqGkYvYVKGRkHEFDn2DCMUq60nLBsDalxMJcJvB5ZIoeGR1vqxowjQPGKMU1NC
Fyl0jxTsc9csXQR1kd90pnBWDgsXp9pmQyBXNYvX1rl6AzjOYHwAZAHMwptP+HHH
EB27DjRE6afUAAe7kohcHRX7ZD9gtqHOirde1elYTKkthpV5XX0XsaqJ5VXeRonM
uK+TRb0WcEak9BdozLb7d6P1sRfRThrfAn6W9nnTTYhlPONaqvNduLXCxM42exjG
bzvR+E8otxvd8iKTB/jfA79uAmlMirPd5/DKRKJTSOmzpNuL1kJq0kEAN6K9htOG
iQsvoxKOQxmfB77zOsE1i9hXmRMb0fcY7qm5nKwZmJSvg73pC0p3ie2EXe9nuPpJ
r+2+ZgeHsa1/7WfSQGOPPau2wrNAZEtVIGrODkvTmDQXDPblVCdadJj0Ho9M4e7N
I1XWh9LVkZwr0OKmw5hLxJDUtq/z3TxvOh8VlSgTkyfonI3X3ED3EgVDPExS4hXo
RcAp5uMpEGS6yOchvO00It9w8x+jM5Wo6dwwrrDm83ZtvM7FeLG5b6v7yRN7F8IN
p6JjWDlsHkfQEpcIy+aO4fY8DdpShNNFBvBqm3U6/5tWgo+UKloSlgA+T8x1lrTS
VuAtf3wmZlbdfsMoRCSa12WMTrlpoAYCfLMGFFysPXTg7X/9PavYIoecEeQsB3wp
XIOHAkGaRezx8NtMHKHH9Mp1KJTxl5oFcotKhP9vF/lCVtdUvbqO85zF+8PpvMqq
Joq6oD66unpTH+6iwhYNtHtLSGpi6JnHN8nWAVHGznxoDeWa6Qd2w7LWEbrWt5P5
po12xeFOY1VtJZiGuvAJSoe+3WJGeYCVQKqEnERo2WX86ye7P5VT+kj0p2Jj11PV
LEyOxMj1BN9C9WuYpq+B62iaOl+WRxmSjbkR/uQp5mVK9M49PLbQEky4sBuGOw/J
frJmGSCIN13c1/fLJCil2W/ZN4lyQCOlSI5MxTp3l2vADu9qzqjUAJ72b71Ikb5f
ynzt93JGWmojUSx4o8eTcEBAeQr9gKN9eqyDwAL1ZhNCMgEXkmmqzsqK7jsy5McJ
kuMJ4nt2uWWaGP69vz74HATR3oPGknQjKji85rhQi7iqUJzw/Cjr6PIE9f4Ty2Zv
/lwNtQeirZ1MJ/bZ4RQortTNnolIoyhb/Fx593/qXWGPg+UbxgbJyiGUUGtsDF4k
Thm6AcHrHodVTyKoln7kf68OI8stYD/e2Bm0m6Iy1ZcM9yyNIrQfwssejQ+j7i+a
M24GbebeCaQbOQ3pV4xgFig53rS3d+9RchOAUS+68cUh7gJPgbMNza9hMrXfVV2g
tHq0C+aXHkqk782zLdf/d2K4dzUelRYDr7Ya1v8vdRrgltxud7jFby/qk4iMH67h
caiFVidWyHeZpScAT9eOw0k3fjRvfps31Z5tkaIISzHtW8Jg7FbImuNth57QF80u
0NktR0faeJEtz40eYR6+y1nWbI1dBYAP3/iib20OU1MUPvm5ln1EiMpLrC7i8WKZ
+0tA5O1Y7PYF2DEAnUlwFWiTM9TVikRmqMbFsKlBbjlzySd6bs+XhqEtKkc4H+cT
/shSKtp4EhQ1z12k137iYNfwr8gE2dnyFVXo6fdtaSrfUeqMUC0egD4PCQX4o2rB
4xZ2aVtvAjCPF4jVljUw2arH0x8C8in9nbfXlh+GTayql0E/0n1roYqxIYLSc90e
5Us2+gG2mjDbpWm4GL+HpcR7En0Td4Vhn62tm/XH0drlRny56Ba4bq+aBuMb2Zkd
bpq8OxI/gSgggZNEbomn5AqMqE2vtSfkasXRZFH6Jb7MuJE5qR2Yj8f2YC1Gshwt
TboLqAuQVoriOFecnYYBPxDpp2fbEb6Q6foLOtOA67gXGtVgubt97yKQ3vmijmGX
fGQRy/MLQw4D5m9wwQbsuoxXDZTRm5JHGizK+ULAgChwE1R0ijur+UJamXnifAJr
5qZhtj8v0w4sb/RG6/Ti8Wm0wBM9TuIU1N1at/rQQbLi3XSE+1Bm5+qm6/HZ9rEF
l6elwhwuGGCEMDGRL6F6+2X+NtzRI17ESdHyXtNdU9ldedJzZ6j3ZLDCvuGXZIX9
muG13pisdsbI08/wjrxFzvahUFEhJRVNRqtUzTB2jgfLoYx7z1Gd/cWBVIAWyOfx
jFl46IAifaQSI/InRecueHCtHKn/zM0gDjzpoIGG6PjZp9AnjM1tHXrZiO5KEtie
KLPR8q0DGi6C2uaWeC2Xf+8SHSdqnxRoubT1iwI8C+0ap6UqH4hG+yxVHYoYu2Ui
2zh6T/IpsI2qGLY1OrtmT8JlK8in2zVV7J4zO0vqjvKQZ43uL8p7GNffF9Mn6Z+o
3gCA63jK3OSFtQFVpn8+NPe9m53QJUanrUuZbB+AgmgcgU8wwHk2QeXTZwLUvuu/
9iCfxjOlxf9uT+0kRk7/jiggsoWW0tw2SgJ0vxTub/4Pr2A9eLX4JE71fh1gfZLU
R1+PYTUsdNVbr/Bhhu8uCZDTH4r3fNqVBdJGqaZLT+SldVBWmGvlt92n6ioWwPBE
wP4FEVaC1R3he2V3bKKmWOTWVe7JZLrnJ7xisTBmU3ZZiU8pYqQgU602Y6QtIYhR
E3IymPvPxjeinnQKzyzA+NOBHDY24cl7e7voRWhgS70hidZwRxxTnyHJBgQaxe3a
vBZPUx9S2bVmk7IYze3ZFLXDIgyvRmXo1yjJftGQuOrQpzoqCegtQSjR+Gkl96KN
i+7KfyJqD1V9JlxJyuN9WWlyGUWKrdH+90WEYIiBiESS4OwXVMtY+Hc9Yx0hZnVR
yJUcXl1yDaHaX/smNwtDr79vBeqwrNGEKgeYgfzlVAVu9b1garjhWKflDG+ZM79R
ntiUorIfvCLchUO/QOIbhMgdOeMa1ujof/kmk/mc4EPDw5HrCfgQ6Er06by96KFG
0VmZFE/fjY/KZA13xpptZ4gBWYXPe4cxp9dc6NGt2PmFrjS7KPNMfhYoq1QZfL1l
j/igCsLVFwYegtQNNHLC9FyS7ywuANZDa7Teah4wYP/fWho/kfBSnc3PROkNXRZt
TIGES7icDEWZXn2fQ2wTRzPtqJFnvD9PChTWUi1QpCP9nBZS0ADdJQEMUBtw8kEi
pztI0HSP81TZPIAPVyvHUx73acwmaWDfxSgvabauRMoOBpFVDU9NNQzTQAIwxuPS
Pwk0Wd7CzD9qiXkvJmpSwH1oADzN17B5cBWfROWqOxojXlzNowkxnAIfv8AI1kng
VNAqq2HeGunjrfISmc+1G7oRDL7+/9LNXGJzIkKR00J7QtOpVM2H+EF0huIQoEIu
Hnzhh0ET/SBqcCIVzOipo0tk4+QWRdViQ4OrftzrMSliaDe5K9NFqfzldCPx8GM5
hPpoExzt+bdF6QQWOKLGA9m61w5eRB3MCn78AtLp6n6uWS8+AzKeFsmIn0bumpxb
AX8DHJhpFREs7oMMvl5XoFPyUEORtwIgfTGv36ZO1CVdsDeMQfvFx1t6vzU01xOU
TylbYKYj7KTqCaJspIE25cLwFVw8oa9x3tjlA4PLJ08UhJ3aeOI31P2x89Ec/551
e3BrdJ+iK34A5CTFHoODkaN+iPuDJhsgvJFk0W/WMFew5+dMdVgFB4WoXXRV2wqV
mLHdLQha0tfbEdGm/sQwLi33wI55DgW0nfc2Wudt/PLtgz33Y3hAx4ICtx7JK5vS
4ijY3PlevuZWhFzVGT8/Rtk2tbjVlrtWtdfMdC4etXMa8lrOjbzAiIsIMQfh12sa
MLJ/mdikScFp0zgJ/b05h1nVGb4Z6zGshScywcai+8S7CO9FmO5pOmd2JDNBqHOQ
hlg9Os3CQoeqq/rAdlKinsJtppQ/1oArILmpbqYfCzG5Fp2fVqhgdghPgA0xpGKA
EnaidtSb4U38tZYTl5m7nhVISuKvIiimO5W/rbYlSbDttIRt0ODpiGuw85ze4coJ
Ma0i4+BYrZcN/oCJHTmm3UJuhzJVdwodbGOk25X5dG3U62BSSwkyjVJRhRP4zYwd
xnAvOl5RRjXK/DG/TkPpgfFYFDbdLDEuzBUMjJGL30uARGmSVXd0dfkJ2P2PahEr
X0E8hf+ksmJNyVKfvTYb5A7l5xM7mB5I2MuNWhRy4ppFur5hX6kbYkCWTH5E6be1
GRxzb7h/lcSlnNlgpXBblubGyzbe3BE4xm5hRzMHxrEOgpabcftSdC7mdw72r+4P
hvF8oS7O1IgijUgQnn6mo0JKd0vtjUdemy65brLeFWChPx+qg3JOmOhlbpx2VIjS
o8/dTKXlM52wT3NOSrt7pWv+VHROFDTaLxuYbwK6MiZxKvWd7/ObfF0c6t9LYO4t
mG3NjpKsEhfdynMQS9HK07DpyUcteYUkI6kCEnQB0EGGxIrmmawKY0X+BnoKqxds
7uHww5H++rEod+eu0vSOX9wTSm7MAhcf+8mF27DQs6p+iDNXYeN9n6qUnQb+lJeo
nW52eYGr8Ga7Xe7g2eKdN7I2HTW1/FtLtCy4Dbqd2qcrpRlXYUzUYqOJnVC/Ngwo
jfPReX2Bc/scLorcJNwehByX48PlfsAmo7Ko72bBLYMRc7KVZN+zCj2VXlplV2fq
MZJ35TVHiWpziZl16U3dEYrFEwNRqWUHhnIj8l4oiq10buy6yoO0yvj/Q49XKKmp
8t7PtuWP2JkanucEvGVkLGNYlKv8dv8AWWxNIIQbH+XXzPr8rjlLNiVfXEioe/4d
5SO4lPEQzhSXUkgYH1O/NdY6rSQUHnhF29R9io9fVkO1NzyVD0EX4Ft0yMszUY91
u7nGdnnmpga+AHnD/Hj+odfsMGjem3JuaMNwItWDufIZPBUXIGDy2HPfJRXeBe4c
heCmnsgr3NGafjCfVhCBtPkjfw9xtIeJTLfJ+HBFhh7oewosU+5EgIlUV+LjnbV0
JgreJ1CAA1nweiQuJf26JUOJzI4HJ7CxoOSdclQsii3kOSCNzS//8o2u0E060EwL
zyCA5wh0kPFs5YGYrLQ/dYys7ftAAs+qY1Gu+K8szJEBh+n5C2De76IbpZrcjKeD
wqfrypJlwicx5c0yDBF3vVKLIsDTj8L+CzDseQ+pPGIrz7GuZubg/fkIvduyFyOr
b7EfHApRcDBgUz85ySKIEW7m8DOQCGIp7hbkP4nzNxzNbZ44Gr1TOPvbe+FvqB6y
s9ZByH2SKE3AbbMjyMJkTH8PMnCyMOOr0pBeJcpWDqmSTuHIe6sZZa8qWD75JTOf
VJL2TL2qlq5r9A7NIjjPCbAkUaYT9pDqAgp/BpjU/4XZsCB1hm1W75Z5V87h3ZoH
18WHup1J+ekBDRXsHHSkOwun990PU8Gs3DeQb1AXyLRNBcP6D1Ez4zMwrhZoDCJF
wmEp3SLqVIcecuU0bvmAiSg2dz38XlCeJUTtBHP5Qsy3CZy+MiPlNVhadllkabaK
EJt3wst6Q4hMFmQXPZPz63tK8On0eDyu/sErwdqMTf9UGyhq67dotfDc2I8E7Szi
22BIWKTsutiQil1QB2Hl9pFuG9UAIPijf4gYIolNlR1nr7CzHtlXVlHag5zf8sJs
Wkuq7lrXHSPgaL2/s+NDo3y26alWXIf7wskBA6ylNQ1a0aeOjOmepzKAfRhqqs4S
Hdj3id+3wffAjytZdLU+miXzqaWo+FFp1m4gMOxDag5txnb6Chj6mGtjeYXVdNSj
HHBAa2eun30/eb0IGhMgxfqC1BDXEbgvbWAYoCo1yD7fNuGRmRjJcLv/yAGgi9en
z/pPFbYtNM9BnL5UM7hZmwwi+MNB2Ia4zi9YXOBvGrRAw7AN6kBM2VheRi0qqHPK
YpfVtKpCU5YbC7i62tQVr8FfCMT6YurmMIEERS21+dyIYFMZAFqw7oJN8VysVIKI
Tcv1naiZIgFRnC8MbBjdZN7j1amTkc10fXav/RkI7zyC8zvMRggxB82fwdmvdARa
6rgjRFQiYHMSk3k7BHd+opPr7GcgJzQ7dATe7ri8NBQ9scjBUnoFthjFf7xUs/Y6
m+bN+Fu2jTxNAPdrwc1EmwaSY7ow9/q7k8NnWlKGSh0MYvJ9f/CoiUHaqSZ97ZQZ
hz7q6GIPvs/anU8iUVKHPNvLJS9FtvN6mFOZoFDC7q3BBJhJ6xH/1czBIjDVcQ02
M2MURLhg3zs7QtoBZ97aTC/jVSQl/8hcxY5gn+1vIhdzWlR0L2n8XqO0QcWQkrSw
lRMa5EgIpKrOeQiyGKRGqcHfqDXq3xKJcMRdbiIX5PkYh3n3CNrgMXIN/TEy4enG
auRZfuP/Giqr15YlDUpm+/3B3glnvsdamPRWhbXUQTL/DXEed5l6ayLjNefPZEkn
QxWLiM2NV8JA53S//VEcTYN+vDmZTFlvJ+aqha+0Ru0DyyztSCeh3naL2cAOJ19y
k0Fr7eFGGwItYb7ZPfQECM55/oRPm6lpOwICbTZcYbHJrYy28OgzMelnrhU046V/
q6P3GOWVZQozJOiagvhtMrJh73KWr+UJz7I5SmZlKQBJEQiFFO/914hUndQHC9Zn
oLRJL60/pHyrqXaOFuVBA9zcd0vUV9PEzhxpGdj5QNTvGp5myQT7ownNDRlcUsti
REGlOiROt0ukDMGvZKGkuulbS8ApJsvgjGZj4rFH4XsQHrFMstBwHW9z2dJnyyG1
puWxhZuUZJoVXkHevioxxaX2wOlR1gociU+wn8FSFK+W10gr2P/+0syD5EI+Vf3T
yCLBCVW3Jz94yfST9eZiSKHW29Erf19HKOhMgqbWCZbyek8ZKCG9G/w5Pimb3W1B
OZak2czVx42lKdpZ5I/UxGE7UXZR3c1Ul3G79hjL76VhoHBrjeroDP2OtR38f7VY
KGpGfV/OE+oq05HKSlOzZh+q//VNWLrOdcGFDdkj2qky9bfe7rX3wsIbBY1jkj2R
DTU55QQuy+ruNQlcxa+yDTuLDorrHQCWD5RZh2h784RKqACRtt5Pr3z6EPosVKXJ
1K/q8LshXIDBHyGRxXIDHxSANMgI1CkIZkkQuX7D/5e7VlDbXbkCm73uED4CWKwD
ohiXBzOyUgIjOZnzWP5uUTQ8LewLN8kIqVFrlMtnMSJ5ObSg3DgzmZyJKL5Jj71M
Rn9Hj0ZATzW24DIn0QgjXx0ajMfhMqzzJmMFj2PuwjDGGzhOptBeKx5QNSTzZwJu
9AGUyVsoiikF7DT1TVOhSaFdsbwDaf/5JQuLr6mhbXGqT9w8Vx368RVsopbQ6A5x
T6pKVKGCgjG43FBxUgeFcrzfZLhG9m0rDWKFllDJ46sQlI0rGC9n2mxdFA1peWDf
xmEA+9SayCqxGYeTHbdg5WCy6ZVhP1l+5MrAdTHS9NZC/mgr7FcS9bwCfXmm5hqF
7EmO5eQg9WR34KEI9p5t5NOY4sSaNfFD05a/LYOK6hX04rYZESuBfODgdy6qc7DW
nTJOoqQR97IGTOnAbVqpv/WtuyVn2R0YPFQ4Qu3Uy6i9scsrLP563dCVSOpNXwxC
ztnIPkeBTbnk3fh4F5RacZhMG5PiLZ44geBxsaMdp3ibyaiV3sqfTlwAe9p3wqjz
HIm70Tyqgib3iy8vBLxw6Ga8XOCUID7nWhAY/e1JnX2MWSinbt80L5wyFwhlqA82
pxsZW1ll1/Wfozlk7nqBT/cE4ymYiB8J5aGGEhiKuKUgIfihQpEfzeoY2oDuwgCX
hWEQ6ae7WAvI+GfwFXqTYapMPtTMdaoqQwwGaneXT79/DtRUUxgXWRyfUr6QZ0dT
eKUhIZe/WSS1LcEC6efXDgrYYe2ZiGvtsUS4nJlrXg+nR0BKw4ZizCIJLAkwvAqO
w/BuWKkmPGDwRfpjxEuoYih+V6ZzxHxpBbd9Fms2QwNv9vtDeabzkNLM4fUdIaP4
kUKlI08edojzA1As9x29bbJgil4wVAHJOBDKGPx6i6wvtgF/y5LHFMji3rDUIKud
KWcpqO8tmqtTPSQglLLe67kQIEGWONKXEcdfEyBWyzpuBW3sOprDqh6gudbrK5Um
D6HO5eP9Kofhf7D+sz7m9otAtZD4nnQ0GrseeJNA74sbcuNYUjpyM0qPWPx/VDU1
GwnS7omxhrCkTVTMI23ustU5efIDNCmjRgAuqLsYvAO5S4yeL2LrZscBqFZBRyA9
RubbJcA70dVJZbXTB3TozhR+Evv7SjoxwsiJCQeTl3pXcC1J26BWpvhK9dgStZuF
b//Fwjhr8K1NXuNGqhE/DCx3DbquIru7q3hEh3p5wdmaGk1cRmTl/LdKjx13BsHr
/cqWOAKmV4fpU93WoWZMbnLMS3DNyKR10saUQ8XX6Kavly6T1MepRa3F1Mqn8zTT
RK5HlG27UhG+gquldj8jJxn9o4j2EN46wSVjobw9wek11A+clxQkbVzNvAIiv4HJ
OE0gObCQXOhEg7zHt5aB0Ogs0rNHLWgA3csDisASXmqXnadELOV9EXEWSc1VHy/U
KoGyEhdfK46lbOFVNNAbh2YQSMG5ZgIptZIzD2SlOVCvyHKc7ygrAQa5CCcFGh8L
ds+VwZH32TlzLr005dPIon6J2wYtjrLSuJPah4zfyZOXZt3SXqizIEjRrWtNq05b
wPOmTC8XtoneSsOcOkALNuYlr3WS9tckxsyHCagWYotSlpgLUCK5kvbXMjTiqrzq
3UJqlIduuM3jYffNikQeD4XlflY/r6A9PLkAdTeMHjEqCoTHTkqPQ0ew6ZWyxI1K
sRSUphpEXvtgik6vaNrrF098LBb82jOZza3PEloxYmLGnZ9dVGp5sosOgI6utd9x
zZPlmxQ861q6JNTBsZWSVt4sn+lSMBQX5orQp2NV09x112rocC5fm7A5TqxVcyuS
SbFqgIXRaIu9G8iKSEVuaaLFI6pPjLEBry/HTBZ0gRLXJ5FB1BL3uXPlEIDZ43Ot
+f/DVqnvCWIQbZOxotQd8mNn0GKS+JN3jwMXI2WG5MXyCXgtrmTjEBelL4/54jES
zEkKUf+AbiAuJRi+XD3XZhhftlXjR65bpx9aYLMvym34l6dWkKV+E/8J4Wn9uMnM
H6lCm/u2b/SV9M9TKLEAw82+Slai6Araz8vz5vkC74tiPZ17AQp9mld/cKIt7hxL
b+uJCgNurkZyVW0CBy4N+SIgxyVnNSEy6gAVN394mmuTvGhA2mm80tO751qPJZut
bEb1+4RWADAGpc/snaY7lZbC+s1aNAH1tq5L7fS/eZvNgczAjhcsmITe+4d/30pR
ZV+PQFMTRQ35UnnRx1r+OrZPGSx5X97hRM60qsPo+TbCvTwNpZ5+XXOWM4b6ocdT
iW6BupXxwdlMBt0SYFhTec8vTbx8X52M5/Piw2ZsOqh9tkhIM3swVQMjxhfkKq+A
yQucqRqeHT8si7Lh4YcQX6tI8EWxkDYIr7ejq3c5xnqyppp6UkVM0mQ2CwG5Cg8j
86VWxxQl0XNFGB5b5Mk0PtV4+M4PEhxsB2mNJz3Un8/joNKiphtux/3kZSRvB7RJ
JN7VPC5FMEZIyUeD8rcbcxMcbZwPz4LkURiGF4GRxMKEHvL9r06l2WN43oJ9Gx3D
Qm56PivrEKleOtGhQVWtWhCFX4xaIJknaCOH8Zig4h2Y/wTauPjlCfiiD01otXhX
u72AbMkO7Ns7dyGWK90tw3leHFZaZiEZdKVZv4AQnLN3yfexC9fC2Z/VttPg0ggZ
jwBCITHwuhuuaQlJjonzEbJg0FYrvmf0lBjDJyQ7fFa4398AaOSwZccl2+5+BPGP
nS00z63VlkFHxGynQtefkWJiMzH5BWZUT6w4uWcjiaAvD1Vgsqgf+6umvZ+qFvMd
2yIEB5J50kbflrMhF4+owc+iDySBJu2j0k97W38vwhg/9Z+AFs6jH6CdGX0X6zW0
DowW1lVw/Kk6KKb6+TxBL8rWw8FkpoQbZflPHV4DshQd5r4BmfdQaF4oIA5k0L5r
Ft/e8PUaiyIHXgoeqU0u5zvFGSgDkqOOoedxBPrj/XCB+n6INe1zvOui3TNO6rk6
+fr31kIPBFVgn1Lo3Fz3bpFi9fShWXoNnYQrUwNe0HvXImLdFqkibhq7vF35Vbcv
Gk4R3tH4ovp78LNkrGZzsS8JtTujP1KjPYIKMA9bGR/j0Ehdyxzr94V9fYkbNdzM
NhsxgCsvSzJ4LnB9pYySSMm6OYwWHUqm7WKWnXZG8tb0VN4ZtuAYCEo7gSI77g4z
N3Tl++DMV4ZShn3iM7T8wDQdVRBtWJM6Zyb+RUAu8eFBLuKn8dgHVJa9erCRGiDj
aU6Ogit+JRBRRu0kMdu79Ls1+vxjYnivoIOxifupQlqEXaNLS0ZsSp4f3FHiXVKM
uBdsI+WpF94iak2j3fN3vk9x/OXVKERv/fxk0JIURBMYRGI1kf1BB9vZbHmkwozu
muTtkTLDoN+p4wB77NIRUU/e1gkVFb13sP2Y6hGGC0JbDgGYn3LMyMAoibQ+4nY7
EGeCHy+tTm7k07zS72fxQKTFVTId8U0rxctJW8otdOgrWZwOaG7ykhqGJV7VEmf8
u1hIlEFxvQaKKuxb8ohQ8br9pGZNm8ePl3n1WNFLJznVEdtmRawKNn3DgzCl8Der
yglCqVTHdKTYDuORv62dNCuHqNtyyWrpSPbwEP8EtfIEOnPl/3EanJJ4azs2f+3S
CdwyLGviP1gB7JcexxVxAcXe9Kt1CzDp5gUfPjE+mugNFNkOYUAk2FCu8Cj2yNbH
DexU8W1EaCUem4Y7fviIWLi38rMPnRhVRY0aY1zYrx4Vby5+KnK1WbQmIyPjDTZs
68+SWtEhSaTvHjHfkf5WfkrJFKmls725r21nzLa0PhId56Avq78qUmw9W1XrgBo+
1Sa1Zhx8DJWyr5bNevXAhyWo63VKk6RCubcbjZAVGutAD2rhXHLgq3qtHbP8ZOdY
jyKRbA0Pevxb0Wz9tpcXbQyGPE1BwlC/4DCiTDSgt0RgBJn6u8wZTN+OeXME0YlQ
xdDNDTbb0eZ0WnJAuTYH/K0Thgux3lsu9iCug1NavE/hp7tDeAb6zWM4uSAmiR2i
JdpvIBXNMLDSV7kxXkMhN1x1So3UHJMQOazUikzJW1mr1vWxm4Mzwi8ImoYb1P6I
Euzl6x+FZRBnIJxG3N1wEJaDwcpMT61/niUXgD50Dd1uUosRxIWWOuJym2bMKaYk
UK7QU+JaVbw076mghP1780HnHFETmfKs3exLR0OWVyghPJlXWYc7LMRGPtgWSIMI
DIwntQNT8gvOx0ABC+dM3Ql31YSNg6UTSRiOXov2abmNBgVTkvKMMAs0efReNSHL
+Ucz6tLlzsCtrS/2v+9Qh3pLvJ5Tihf0Djxvb/6B7sgl/dntrQ+LoNuAThJ/EOh0
b83eSypMGrwrhfz+xZQDi4oLn0gPdQ4ZzFpt0RZKYGAI9altKnj6Mqv1QV73L5GH
xfdK+m2nDWYAJcLd+MA+VekzpxMrTs7trv5Wac4Xqe/FBSXOmKJ4GlusERQ5pZfN
MY4DpB8Zxf9kkF1kjKDrTjf6YBtotoE95LW2JLjlaB2w6hWFgNSsJ6KEA8Si6pWE
V8RCbAR8KRa2dLIWybt5NGT3bG7gQCfzyZpW5cWeyIPwOm4npuC4j8d6EX1OApGX
6wr1WxYhSEJKIF2X6IdkkZKkqyQ+7ad3M85iWgYsXj9D0Xe6danaekbD7G3yprGH
CJ1PD2rVJeKyBioiWxbTs9deN6nyo1tTe+Aa8JK9sxHQywizBABU1QD4OQ2aWt0i
acgMBo3v95xegEx2eDMdAKgYBoyIaAut/KXreXdnmgnosgiBSjydjSOGjJNh3rJS
OsuGsDal/HlPuwzub+A7Zba7DAP6JuvOGVaJdVORO1y3vCUCDxvY19tQY0CX21NW
Ms1nhT1xBFApUDgmNk4BE4N3JtxF3w2VwLAxJ/7svOouAExGbGRmxwsWoEyuNyuS
v8PYMQkBZJjONHj7zlyA7vov/dUypT3jKtCsqls/5YSAJEDWa1fEG2QyWft4nxO2
yy6u2VzOnjNFfE9/POeVpnPO9APvCXmZHmU2KjNVKjnqZVuvEr8cGGbN4NTIazM2
Jb8J6c06iiB6681AX33XngJWpPMxxtXCEwJxbdak1modRViZ0fWxycIuhB1vwSak
nqJxv7RTW3Ea8PyXp2IjQ7t6dtj6Xqvs04LMQGAqVhVOQypx3xD1SFaO7i/YX5iV
5RY1bxD74BYM4TZfRNO2Gp6fY6/NjQDfimBQVJ34GsYJgWyfs7vnZ7KXn5g4O9Av
L9zoQxrCUfirYRfmkBQ8+aQ+YyRAhi8nBDXKP53VAqUDRIGn2oCQapqrVrnNj3Y3
7YyPrEVpFMmmJvH53X/DFQ2DZDyRS38it4Wh7AkcVnOv33+Gz6YBPsj2drqgYHqZ
EvEbscnTqNJgFS2pDVZiDNySLPAnT8V+mH840b8UDDiBr1A2czgaQRDx5LwMCj2c
Odqfbe1eBCfc1y3IRvZb+cesUnqgc10Zk0H7IF0rFt9O3IiXtsLTLY9Yv61jRAtg
q7WkyaAAYB5/Q9u0xSv0/c/uOV+hw7U5D8DkOLz/roXnZ0FCS2kXKlINdnKTjzAS
eUSGbAvE38KD+gF4hpc2dg+78XQigvhnytZdZIPT5eIK6i7AL7mSx2tzTRvBryyH
kOdvjS0NgrhISggUToOmn18uT8ClESwtGVj4fCYUqHWBBvsbguNCv+3tzpH5HthR
dRkJckV5+kt/fftarMOWMklmT+gloAk4TYQlVwArhLTFR/lziZPP7G3rnKA0IxnY
tFTYVtYM0/uXExwJwC/su9grscM0CkpE52A71JVoOqR5kd7Ri+KFbLl9fZlt1UUh
R9yiqdquWZEyBKvhraQ+ZdVKQWN2zAufICG1QK6gJma2lXUhnIxNUAK9FZA+i0D2
yC20DspZ7WjSDmUP+0lJqK4rXV9JWL/Na8uCiNk+anlTZ3f08dl+Jgn5C5BstV8w
lu1zsCzBmd0IeeaOKHsobufNCTXJ02eA4pulj1hnPrWW0ELwXeq7OYGO1KR57NV5
MgfbEUGcGD8MHM7J10GARwWoBtP164TLXUQjpchVSap3T0zGfc8SqEVzkNnCHSnF
qqZstxGofRWL1ngL2C22gfe4bnP6ZbeMbUAqDy4i6BF8vu57tc7wE3ueRrvbW6zp
HMjhaL8DltA+164G2Fn0L0DEu2JV438dbA5YCIcKCbw/9ZPcKwGupyWor69XU4Iy
x+kWl5GO2g/I69hp4CCqp1SsxTX+TRqa7To4M8ypiZsbABzZ5xlE0uC26KECI9gA
QZ5HIR9UbQ3gebTvzZ63QauLWHW3Ufveba3tj+REjZWW8dl6Z/yFrDF0bxtsG9xu
6SVh9rlYI9h1t6NqmgTZ3Re2gzFo+Rs9z6fT3xCjJkC/8xCRPPw/JZsJ4v3NK7EJ
NUqIDAHfslNJST14IB6UONAxHdFeQW5LMk5870PpLMa0Yx36/yoag3nFdAhncVnx
SDxfh/ZPOxwReE1Yi5HBcrfh1SlqlZpngVYj/OIwH7SQ3aPAcVaayPN3djZ/yc/4
VVin45ZjYwU4JPx9AQ8+fbETOXLHSLMgGENNnjzoflqVrtLkGZZwy9LIKbPd30FR
UKQhBUL0+4D1fBntK6ryAjurYWnKV3sHj/SapnPlDDWqCXRPcpOZ268xqNe2AXcR
qNtawChucJ5wMFaM6ZSjvkk8k2lBWQQvth5wQIHf2VJ5Tj7bUjJz1+wAwo8dCohT
5O2YSU1WzRbD+a8DJasWEeB8TiSIe57nl/tGrKQht6dwpvvIri6YftqXrYcuH7Zj
ptP+/bhkzCJaT4kqxYdBOmfpk/huEpcMJXeKZhReLbvLoS79YcKaFnRABv3mfHkU
tkqD93TYeKUvra3lwkG9MSe9aUsXBI7KsygMFaYofj0uFhFdeZtzilntih55MmX6
SX4mmECjp35StASwZGfHYPRmAX5EOwf1yNRRmmtptVhk5026qZjnxlhMwJpWOzBb
ESXhlWxO2c7KsKlKFJ5fjMWNKf9tPZtPItQwx9bLYE2O9IfZ0PuQRbpV6wgWmGji
nySnMaPI0R6x4YK00nYpiG0m7A5GMTUvMowv+bq3TtcATBFLhEzPKyKnu8bq0dRL
b5qjAKsYeTK/YLIWiU5rkXiQsxouelAPURXhSQleWtnFhdeVbpCzJ8Td2jWdCJLM
1Qy+OSvCAyk9QUO5dcVSoq6rBxk8QR5CFvqc21wDoSBmGWgRgWcSjs5v3u+0OReF
/IMYYPKpsxydmNhYvtpwd9hGvljI14Kpu4YMQTSVbCIHwSXt/fR0IAL252w8qM5N
dpcIpGNel6Ctlbn2mqefLowODuWRQa0h+n0ajPqWUUh/Ii6vU6s3Aw9HXM1hY3+1
xp5NQor3+q7ZKitsZRbMNwE4x+Un4foWXa8trsSf2gBgE6hnboCtQQva79fVOp2f
hddcS+Ywae7nw7o/H2micXedGqDhDe7EhyQhEDAEKJ9y5cSVrNYlPKR+GArHmRlQ
JLN+HnZGvtw6K5NXVg/Y7aUyHoqXsD3bJt50OZjWFkEVaRH81sszdemQxyVFFeWH
mvkyPvLQt/bHfaOxMzNf3oBkUbtDxvbYsGUmcQWQA1JAUDvb+bcg0cK+SLXb4Xah
RSlWeTeGl9v2V2/R6LqXbAyWadhMz7TUYjNps7IBMjQWbvde2+XbaeECRpViljMJ
l2BoxvX5xFhLum47MvdPH/ZkPStmLrDaOHyR0M51p4iQE+erv+fyP1exEitImWXt
4/dOCMdX2uHncWsjUZdVCtGu85dFFj33RTJ1fSTSpHtZJsFJhpn1pdWNBtG4hWIJ
bxA+pgD/IVCTiQZp/LbQfDOo9evIpl0gsW9p6e0uMXeUR1rZ5JSs6hXGmolMzIiA
hHuAV68EiMSztfaosXj3SQIVuDytIZ9WAiNRSAvv3MgvOLzMDjYGpqMIKQvVftS0
M65cKOdfyobL+nmR3OWpQpFUyyMtL/YPk+kFuYGtNRgPXGS7EZucSIxQsK4WH48d
JjA8FusDCx8XCt2UP7GhtJtYhLNFJ7o7lTMUZqdxkcTJB3BqyKqBVJlyNBbQChj0
Q8nNKuVxocSZrwzlkEC4N+gH0vcOaAxq3qw/mZnWUEPFjuoqVWxn8LdOnSbIB4Nz
o+pggUji8vA8tv/P+m/B6zGujcZYXXZLIu+p921HcwqAIFu+YIm/Dd0+eQl4CaUY
alY0Y98hLB6DENsgZ4WI4y7Rg+R+q2lvwBfnJAvoD1y1I+YIAATZIVUKjmtO8fZe
cY2ER3Dii5/pxUYg6G0iUPKU47kvUIO/x1o9YePGVeqLgiLmpE8k1ZvjvUhTGnmK
SyqLglyzVAUomdu2EGh+FHNkTGxuqjPmuYPORy8OQCsHQE6/7piHH70Tdpp9IMSL
dXhByyslFbCvlqCvjvZAowIZ5T1zXK+kwuJ+RF0NSy9Y2PfPYDtmXPDhGZrJ5CYJ
YttHa4U+m9rYADB9NAUbH7YUNdeZMK8scRcE7crlQT5C3iqefY1f4JYX23CR/Xa2
iXaUdW2L765sVaILFhTMxnyaHNtJ0UcuWcV4jJEROiuaOALGD+YXF1G/wKoHZTt/
SK10tsb3NMtP1KEIVFNVeMQN1X7V7aW79x5aSu+BOukHyXfzjmNdq+ue1JpFb7iE
Tt5YIwit4dYPtNXH1klBLD5Ed2nLvS2f1Auq8cjrSi93ZOolGPCu8QQm6d0yzibl
ic49hzUIb9bX4E4QNFmDomm5Lmc01I9koESZH8DREBHXMctkvRs8Rc3Ztg0qH+Gv
tHSWxgZjdRRxkWVfcSBNohbXO++TMPW/MuGeWOjF3GpU+ooduhcVvrMkyXeCnx7F
2EOgYFMDz6q7I+gHX2yRuoW2A6LzWstCAebJCB5Z7ZeIYkhcnaJXsb2SXt+XF4/y
09FFRpEfAcHWw3rRt1tiFlgnwEhYQSid97bik7aUt5Y0H129FT7CDUbJffMNfZcn
vIQDfCnyzNWOl0jI6zin1IFjCZtvRzflMJgojj0Is5TismUpQrE52/hVQ1Fm0vQt
jbKAFjREQ0IQgpq4PHt4rxB0/ML1Y+5lCssp9H33Go2o14NxfnHl39wKIbIRAyyf
S2ogiPqdnO+/6+eKCT+G7LDDWEvqB7zknBEUKXvkM0gxu6Amo9W2ctUAqmdQcPd5
CmHxAPCKyupwz+oGk57MgjfWOsZeNgFkin8ZJcF6fBHDqJ7T9nTjnykhG6HjhEQB
yS8VPl/RXmfMTWeUaT47C4Dtvh23V6yLv7/eAf3FYnQoBcDBqplpGZNi51UngH51
9nOvm48FaZH8izsyAbC19osR0GlQ4DjVkOAq4JuOSRlF5SpsReJQB3lsS4gZhf0z
AdnR5R3EcNIMzaalH2FktoCCDC4PEKhJgJI8eCnVW1wAWKkH/5R0GekLuc8y9g30
jJS5zh1Vh+tm3zbz4EdIgZF5audOnBoZUhnMC2pmUtcRAckIwGAGi8yX2E9j5U7q
Fzb2exAdWCdncern6qUBb6IDZSCIcwYd9tpz+UznCaPIcj+oTHbTrzhpgp8z+0Zs
skSx6w359GMUQ9GAvEMHcN3qQldJbjTVJoI5faCEDDNfSAC5ajtYovPuPNJB0rZx
o25SOXpotdxgaE4TFPuLm6JAqAYntUwGbgxWN6xUexiPdaaAb8Wr/VSGaz9DWdul
d/89XUXY0yaGqgbdAmeuGOAFD4O+BdTXBybj4r2M2Vy4uH8S0lQVfQPSqMOBvUAK
10uSUf9x89OSw9EI+cgbJwvJQW6ZhRl5avphN6/2lZUTKdAv43bf6wpJzs0b+mg3
NX1+5KvpBy/vuX3O8qSLitjzNZDxAolY/hcy5LaR4A+gqQ9s1ALsHNKEiv/CVqV6
qpLTaVruhPNBjEjIsh1/Lb7BuEslozo263hO5UT3OsGoVHAUqM/GowpC7kFycrg4
Ipiq7bLXH3wIXVscGumAExFwNktY213/5HkFJxCPtcnWwC5r2ZnkeMeZaPPBENgS
MdxPE9RrEtzDCPFmIZk9M2AIs2A7M/aEQJRg2SidsDZk6PlGIvTVSNlL6ywKqtTa
Ib/U1yWEaWb3tg31L5fKQ9KYJ88NzwzTNpwFhT9XtxbsEfIy6c2iB0RsHKCr1r92
9taQmTuCM+0L/zzgK8qpCUfxjvrYLWI4PH/tBDiNhPy33WoATIkFlkgNvKxfNJa2
HqjsWE8FgCj5SjAysP89uNiLTC0+jINfqi0zTk0r/hZ1+535oRlimibY53EQKJnC
JbCPbgEUUu9dgZ5E+jhAdT/dYFLqthcRz/NLDJq4gNYx+oSP4kKljQ5UawEU6zWY
lzgmHv+Aq6EFLT1bmJjUm8LY712y+Pthu5MS26atNstGmHAMZJjssqPt8Aw66oLS
mRQ7cNTdZ1vWa731bIXr+1ebinbYSOji2z+nmmkUUbincJUT9YL+CW0VrKXlorgn
4TXQ/MzLy1RuZW77n36sh368iUuL/7UxpezsEPGqMFV82BMqw+G2aGbjFaEzKBRJ
Rl/7QT32cXkbHBEnUAha4DunUklUs1Y8RItGLCBo+hzcQnAx/zTx/gl4FYhaj6AX
A0iofNoRML+i4QR8eJVEiDF6c7HLmEOPMXeps6YJBsWtwnbqJEbw3T1tpgcc4R2T
IhbqgBdVCaTu2m5dyVTBjlndsMhhMuyb+AC+BQgVacpAlauQvGwyx6WEIJQFiuzj
/qeTXOBdyzcamZZxZ9hCoScmYKB1QcpGECblvte9O+tecQyurfc3gcExrk5WgMbi
a8k8k7ryJleNMQUgRPkYlHp0ljOLb/+qjf76OiD23hPt8eUOhrCgZmGeFrhHqq5V
9mdPYrjxx9ZQhIDsmQXymXI9RgqB1XX7MTq5cjvMNZseNLBPLU3MhgyBAmSsi4eu
Actz99k1zVfxaUZ5eafoooepbYyVpQ6j2jqrtae0kB7Xj3gbJOMtBWJZJfEi9ozg
dvJQp0j+zsMNLsj6FTqSAfhBqpp2xfbhdFeEUc67VDVJO9Vx6TMxkQXp6idkiFHS
np76F9//QnhcjdAxzRH1Ugaag8TE5Sd2BaBM6dYxdV4sDoz78V7z1yhFgcJ2xoGE
6XPMyYxm02lC4ETmx9CDxIfjeq0037s/YH2J3sIcmzCbj+z7paLRGbnHTlWTEmS1
tALUay8LTcfwh/bJwxm92quYfL9i0/GYQG4Up3w4QRGfgZCr6AzfFnPpZ+mgfhdU
n3vUYLoeoe0ig4fW3ie8sd2JCSJ5S1PMiuqD+if0dPWmqE+poxXjQ9m8rLhhvcuJ
njSNOqRx0vxpHXuwhzhxx+CS8gZ28eNxpMV7munGzjfN/S5SPjKTKeEM/T7XGfpt
YPjChnb87uVLqyJkCcNs925EQC0DD+0gN+lTCNePj+Dm0336jkqDzPslvlu3JN9K
IXFHHCHO19TXqcIa4U6imBCWfF9vteghkH88V6K/K0x05LqQcYukKF/qgNUfk2Xl
JgFmmWxFwV8XpSVwG9Ff7LIiSHsB/8ZF4POEXcfBtTnfoXMI1LDQY4DvmQis6S66
6DOH7mjaJvzYPBWVefv175uxHYJx3ADv8RevZMuMfPSD6x8S8VW4scssxb192M4/
53P2AXQn5uCWb9XX/RiOIcj2+idb8b+9TnHxTZPgAbA6Ki5xj6ZpogubnigJHB53
YRwVVvSzt7RXeidZ+/8dhCXNdg1Sc+ZVYxshXgbIiFgIqwmTpqrJlJZEJSe3UBxJ
zZt7Ni0mTK2Rk5D+ilKxa/Wh8sUyBoCeiGYESCNs5i9P/RFjtkR+2Ij1SxvkOr65
/CL3PuP3UYjW7Y4ImQfimVn8DEFxxdf8qh91Ga5cUDx77OCikDfmWPxqLvSaYmvk
Lw77zl8u5Ahd9sT5u3bJAqTWvlPM5+PGuL6XZ9MFdrFw52D6vydFa0OHRGpf1h1K
+IBqOJrgx9uBATofvpYUHz7DdQRCfcWG6bWYxHTyuCr8M9f28C87xjo8WVCDjOSA
b4yo3V+bmN1S2XmmJyWzAreCjTzCrWVqEgdWo0b48kDwA8tRdPIsl2UXNgiH4dtP
/PRLY2U/fkWDXIV6vPlEIDJu8J7ifppJYS/E4NPkP7bz7fKCvKCnHbgYxxly1AXa
oIN88IOz9zjD5xBan1G7lT1xGVcMnq3qHoGpzu2oJOaadufDqHz6QzHrN0qN35PB
ZLTUor0461BvHXvpSOUGFhAaiNGshDbNepKHclK5h6RJIGaYZiN7f4FIqCxFIOWq
V+mD05p/oQtA1lG0Yig0LQoB1UBn0jACdtUW0DFHw6y7jC2Eh8kNO9WID5gx8NV1
27xvNye60NydWopkWwpA975q0XLqfKRIbu7XrGn/0JW9iHGH+yj/NqiMdivbdydT
lmb7DPx7/Wav9FyrAHDSoyq6ZsuD14oEeqPLvrYTTam0GzcJKGydG7FYl4YMSmhj
fHjFPzNG0zT2oh0eiSttEANpuNnNRgNzCMzlUTLTw79/wubpfK67IqoXGz2qNvft
90eKLSnjQO4Qelw6eB1N85krC4kjrAPkikTKW9PnFkkeeoLdMO0N8OxDOxJTWS4j
0sR3pYh3lEyV2P5C1GBE8CPAnL+XdTEceRxu2rjGJyvzlCOIF/5P6hirPwd12oXC
ScVfCmtFsKXm0iW7FP7fIyuPgI0icdZG+emqZlc59zZTf3S4OcwZRDCOBn3sME3N
3SkwpxluI3ikPVvRJbmmrb68XLrIBW0v5O6Vu5d7YElNrA3slZFAviykS4WUv2Ks
ahLwmHO7xm26nhIXUXVchokdbHGGnunmV6W6IOAgJOMB2/kcNeTleEainT6+d4sT
eANSX2oigB4QLqr5obysGj5u4zr1BNNjyq7k5ljaMLEBUu6C2stJtyS6HOvYJ4TJ
bogeC++IyTsZQv0WE0l60tcXNraLkHsTq2eh7MX8HWUKzrR+V5jfva62qnsn3SM6
4QkNK4zS/Xp8wLjOtEmxtOcAtuPFRon95GwJ+C6xEZWiY6/5G+8gq55AlCRnOd1C
BQJ9Q0R2f3mEBo0waPlljvkB2ac3gV8Yt8IkK/NWt9T+9XE5vsJ3Ba5wOQAbEGQA
eSkF9oVtD9ET08sM7nz9mi8AD1flwPgCWgpea9S+rhpb/2O+pRmK4ni0r3I+5A3H
kyfqvLslMjO9l1wsL0W24Wtxp94QaH5hviowYkEHWp+V1MtbcmqWXLemQY3Fq86/
kZdnSQtC+zIFj76sV0GCHeXtOXvSkN+n8fih83JY1K6q1snpbk4ED3h+2umiqeFr
4Uhbn+mGJorD/GBmkg1LlF9rqKaX5/Ly40aR8L+hTOgnRkZXP57ceZxs/tm/w02o
+bLAfRF68cUq1i/puIGgY8jpBDeFaoPtNbuKWYxzz1t0uNo8IpO/dQX97ANhyiJJ
erjMJ4MLthaCMKESn8/cR1B8TLNBhVmg89hFgV/Rf7kP8XkGyVwf8QLm/EQPGTOz
p53aQnhGqByljc+MX4td5gEnmZQBJdxnLZyXiwN5n9k8X3CyltBbDHP1iVWF5cXR
EI45/Bu0LkudMy3Xlf65al1V31BA1tro33o60by1toNHKnnKSiFuKZ2muskdtIVL
vNo18wvo/5HwP284Ch/lAwIS8tUZxHraWMmgKuYcmz6lWyokqPQuaZTdOxFLlH5K
YnuQq9q3HN5ZSg/fp2VSKJVq5kV40QE3FEN+rMdGKTyHXSUumIamDo64PTtFO1H3
ovdIaMmXFpb2PbpswvYyxKXkeJqTGVvRVGmENG05KTUsHkZECsx349FveuY8tesV
iUGQJXXWX+xhlIRUDhWrDoe+t1zzzYfZ+fyswvjYmYip+zzeBhakvetFjB12qdmb
Zh94d5wayI2i2Kx1fDhZ5smBRxLZ9Wcq/ggfrPA84+z4HKE4ZVGM9zlH+DrDbmmh
AoC2P4BtEkzWNW4P9PjgqsqC3XnFgU11lBIY+pzK0Yuz69jIZSq8HyA8e1u1xmlF
RMTi5zek1F6J+NaQ2eUklPvBv9ZQnEEw4/jNY29a64LYqWPOFW808IPo2DWAokbK
oSnsriOH64akjUNMJhR96poFTx3e2+ACy58qYDqn3t5kgTJkOCqJHawRSP+yAkq9
FXg50eUfON69qAIv9GVn/BPFQ+hJu0Ed/qBYGu3EIYUsKmjM/gNDW2Fdqj1wSlpv
cd33OcDpKLebm0KIvGHMjq4ItdnlGf6rYv8SQcTtJiUGGpcDupf9Fmf2G8oV2ahD
kb83qiQL2sPRGcUwwL7M+1OtEgyB8K4lGoJRj7ZMBqQrbjCL95E8Y9QqAiErXbWu
ZttrX9BmKJfudrWTFEo0hOfOQK1F7qU0r5RXrqBhWl7PNHGQjfW9UdwNbwKSiC6u
hnOLUCNePqjaAZ9EB5MBZHZUodIPmFeU8HfbymiZDog4rbunncAoNIXtDnx/vOnQ
DK3bjV8BxSsB/m5AaCd2BAy6XJZQKnWWLwItEJflHRSu/fXJGOd6y6bSjB0DWLWb
YPeSeSt4MM0W1jBiqF7Hf0M3wzk9Vcmpr+Blru+NSAhbnxeko8SP1TkilRCZQhD+
phSxsr3CrNPvlJhkisyPRLnxM2jiAXUB3yVim8ad/UyZdG1iWeMybbxj+ABw4PD3
GMW6VBdv41Sq+zrxGbjFSWY9qOrbKht3Ml4h+hSgo0DFiybeYsUk1N8PBBggZSF4
cGA1NPjBHoVTejNA+xZJRTZ4z66x9BdS5xkGG9wH3lybMFPzNKrBMKhjfdqYqtO5
A9jtv77csIwMvhoWYi3L8TrLWvjbcy0zanwSsaqKRM5a4m/8s9iLfnt0v1ASjFQH
hDNwEaxI0o85PUbFOYfsXqx2y0t78GfLsBnCJeQQxPwIKoEsOs/JbW9z6nZPqZ0s
avRw1I0EwY1LX3A2FKUixIVgE30qCukIiaIxAYzN2X4gDF+sa2tOllgCLdOtzKmH
9qazxmCZGBzDVAZrxNk52OV/tpDF8YWThzW+YnH2OmSlJt3BEEiTwhTBBTIUwc5K
e7dDAScu5FRGe4I7qeBD/gijhhxSgUo+8U9uV909T+1pd9/Z9XVozo/AGq2MM17I
wS3YroW7y+2dQPp5xkMfyfy7yaCbxhGAr8/vHkfd73MUusShBYzXxT4CGYdL4aKU
bp9ZqeIsHcssg4XJZ9HRczBimoTXdUfdr68iFzFWsG/I14nisulvOz6imK1d94wi
oZ6dGEfrFwRuLvaa3FWWPVRbCf08cIOzyO0ZrQ1FWfthYO8q/ms4Z9k+4kv3BDHq
ag3hNAFI91B6yXcpJmYOKpj+dmUp3qjt98vBHSegr4d61wbrSHFEYhuLnQaGD9N/
7IsMoBRzPT472RC/fDPsG3x18lotwseTjo0KIGj21vCLaRn8SIiemcSQRvBsWRZX
s3VncxzzXf+9pZpgZeZrFBpD7RXQ1Is/FfyTRYRSOSUIGlhvPNwQ7uJXRZIyYSx7
MewQ3LZJVPdS7IRsqTzJAt15u9JVG3N7wq0w8JtcJKE4wyCNQzd/aijxY6OOtscU
JZCwgA0WvyYCpGJoRy3QIkpfduyG4QcFNfZVfIFBPa7iQ72aiOIrVDCVm7GPSRC8
pIk3AfUlFSAKaPFL4zHZd1JvnFLfL0w+lElVVKKoOYgtUBq8u2Ge1qAeS39Irtsz
1CSoPGFseHsKq27gFs0VeHdMvRjsOHVIypmSRMOWsZvPz4v+vJTAEeJBaCj+F5Eq
y6+Yf5fJTTXUpDq35Jj650QfrRnlajJb12GzvLPnJGpDKwToEYSz0kS/yLXR9l4H
+SWrjiCaq25uhQnGpd+Au60LD7sj8UUpxAj1aGcBZW8nuOMB+GjjwcbwvoWV2+xU
PtxexzoaDKHpQWdWwQ9khGAGFWMFtej2wxBvdM5dAGJ8vJOPn83UfshcL+Bh+lrr
+gy+QTEAGZdYBizWq7S+5L5GnG0kcA4M7b8cG0ZeHG8LLz900AXju2SSZCCqCoeX
u66oMXGeTxGt7PY1EVe7shxKTFWpEXAUoJgHZtgZlgvPfDoD2WJuhRZyLp5gY3ym
CJJRl5nHrDyW8YrKReX6SvKnRiUeDbf73/Ssslie22I8cOw8gJhQ5TqoXKR7FVi3
Xz5t1zE24otdwLkJfsESb41UQGBGsWDE4gdj9ltekRlrZ0EN9W733LJiyEFrt62n
HJsuG++ObrQ3eWrUARoxIZEA/rEdy0FrOIaD4SYNHnxk1IP6OjXtlQgoBcNUScEW
ePHZ4TBho5cTedcVw4GLTStOiwyTR/lK0t9DKjw97odOcImbMkJdzLuByJkPLSPy
3G0AmB+L+tCCfNMW0yN4WUa5EpCNCImAQ+RnE+ya5xAcaixL+d3WBWE14CULBoje
ww8vdDw8eGhObg+UDOJN4lJbNwaZyg9ReFZUBTT2eZjLK+Vzq/yDDCbRFtsPBMJB
qYVnljkTRoT9P5Npvr3Z7wQIv9b2pwMIPXZq4EgQZLYPQ6hlw3nRev/9cjuKUmNP
uXpZQZ0kphcDYpRMeV838JmNJetfYqrcVup5ZvYDOfCNnPmRfonJ5z2Oy/sLp9gK
9dTJM1MFflIiQh+qBTCtQKXZbFJ7kgX3n3gqjVAHcgciWAT7UWmaY84QWyk6HuQ4
QkgMAK4l/hB8mG1RZ0KVRWfHz/tP9yTyDWZK6rjmYymCj8BdhQjemreqgHQaP7Uz
QkgdmbvomNi8VbatDnGX9f/CToTqvLD4KowaIfnIsOW7JSR9yRITTI8rfpOa0upZ
qNX/AMV25575HLzcLFMj2SuQZcuOFKwNetomYFmd+n96vxYhwhlInXDZQRSNWzLj
PgmEEnuCjtaPXMZFg/fQ02kDbOApNrJ2BFbhXMLRf3sEGKEKzMoLX4ReoQCQVzDD
O2LDXFlD8JadkWg/grkvb7f5I+bCQgi0d0Kd4r7a8kb39lTxRT6OhdLoqwhClGy9
djTKbTrt228mediXRz8GhUCRuYImO+bBAp3Q6K5MWnTgg95I18f1DcqdFyyXUBcA
HEPVgZekkEx1kSRwrD6r5Sr6FcCKFNzkU35KBSPD86ZgKCF5att+OylDkmsGeBR9
eZySH4zIfOOT9CzuTxHAvnFJTNwaWkm7bcsR75c+Q3fRW+AbNQ7usTiphigMsXWB
1g4QTh6OiEqoH4m9bJmzZNntRuFoA0shC3TdTL4TJdq+TyYaE8jrrTExdfs5BDAt
/eAguf0REsC6rplQSVkI1YhoOH3h8xojhgtVsmjlycr1SNWrot2+ZLQqy/ZibsbY
hpGGSITpUu6lNRPLKifbqfnAuFekbcoz+OrnOfJMs/xrHyz2f2SEtcGSE14sYmm1
rvtFIZzgoO6nNxdAkk49H0/LfDA8cNkOD/opN8V/r6j2Al6V9vM7NEIYF7sODUyk
Y7eHL/JCAiKZNhHHt1K+FlUVsfNh5G6Tuc2J6KWMEPjz5Klsnw9DCqptdtF8pny/
V/Yvvzn/YhQjHA08uLGgNWZyx5pwFF6nChR4KgTV4VK/vi1WbWSVB06UeRfMvj+/
bWTVuNSW22BoUYdDHnG4qWvSwPaNzMeHFN/e5VBpi4V0Ums4Cqe4PHJc8UJO3bPE
14caQe6bwHNEFA9OtWmp585ACmk4+tQYf/ySwX9+zpmYb5DcXL9N0Pxc5x39HIRF
bqalcfy32oC8nUB/Xoc159nc+3yQYJ7RtE+3iZHe1Ub4X41D5I4Jt3nJy1v5V3ay
m0YZCRtXejUfFA7VvvW+By3FxG+qrECDe2OKkFU5hWKm5vEd3rqDHHxqPMeGCV1l
PVmuSZrgCImCpd/3qH9ucEOJIb7tG9IUzQcLK95zLjHJi7Tt7OYPtJGAdBkK0gN1
ZyoU8zrqP3sVHVVVcjZq0pV+VX694eMg0GnuVuw085BJwOVE9w+uSAaYYM3Bm2PF
z/ThWAhO8LKnd2H2SOx0owIeo9KsASUJY2aWTs3UNXv1Y6p0LcbJA4ZVPyFXbV51
SZNHmCj1J7ISJyfYLCjYKvEy5Lp9fzafalNAGPxUg45jkqwyR47hcnoY2iqzUwil
zH4EuV+IafUiTh8HI15uLFGS3/7nYa/PW16uLL16PU0j/8VfKY9N2tUTesQtMQ2p
sQvHZqMKU4OE1hz7vbuDHmbLJ3BfYY5hUoJKuFRUndzn0XEp66du0Zdve33RiwWT
yry/rO7FZMEc+K99pJv+3kKFrbD9h+nBd62bO86TrLut3OOHnqbgbd+SIyyKxyoM
6dSzxC6X1VBKKfct4Q6LvCUfYG9L0WKyk7cNxFj+56F+PKP3BxLrAqjVd0vyAd+4
vjs/zN5mWEelCiuLFq9aWDptKC7IIOrdijqGJhgz46CaTj6FN2P30BSrVy4KhFuo
pOq/W+WCSSgwgeOqlMwCVtE1eny3M3+AoFgl9cTX1ONdgA7GKgtTBSVlf3GLqYs3
OBaltIHZGpgklI4kOOVkdFh5pv1806JMLTsJFVDzh9GAynhETfphQR4630rO8man
buMdZvRr+sdWUfIkbSStty3MeGaSLfGnndZtY61AGnRVg+XHrHU/HpzWcnCR0M8M
1smWeqVi//w30OR2/eQ9SN/Es92a/ZPCvtpzLi3473eRjGYgfl2ssFcfCBzCNIMT
ad0NoU/zncPb55k9qpUDMoKXkjpSXZSC+y0fJhgU0wOCVBsv0MsuWnUKIOLHbtV4
FCDQZnl8IbyQ++aku62VETOw63D+xR3cdJBFSOolDyABT6icaPLSQ1KLdesY8w7X
qUulNV+CUUi1K7v1s7XOHVztdq/1ui/EkbWyhdfmF9MZaaUr6PGnBX3ZlUjCCe9g
Jl3AZ77YA/BnL9cv0iHmbKKfmyb992oFInheUr47l+KHm4tV3JWbTI77FUw4roSA
vBAiQ9n/lsNANEccf13ta1oOnJIDpI+6x3fnDIuG+qbN2lf3Ru1yBrjDa3WHXEpi
Hh2LJxJayFXWM5fgov/5i9eykMYee/NadKFyeegTzOPah4sQVpTzLmccOQGSntc3
OGpoUYYoR7ETXa7wMdvt5c89P2Y1WtTIgk8TMMODYcZvdPVGLZBsZWAhF1/9g/Ze
qyJO1slaQ/2tfuTMA3jzlcxhiwwHDEgkxdCgiu3HRcAsUnDVs3YIEzng3AvLpRmk
YHf4uzlDzu9SPaJfo/Sope1SeZ6DtLLogkIccpBAYFz3Klf3e2XeJJfBPgGW2mOX
lOzO8pvqCFhTxU6mlYycrii7VMmDRxFGmbYgp3MqPX8TBTYZK8AwgLuan3dQnFjB
nHTtYqPQagmxl4K/AQzfMAqrMlnCtgTkiDepfYo0Af67gZzq6rGxdRSxZrkYz8zk
O3Ay8cvyCSWpu5LcIiUGn+okFlnkEy4JvODS/FlykYP4ZA0MmHm9MNm7MnlWYdbc
8ZIpn3qpEJVJjfvTwG9pskkWrt54jh+f04+qKJX7EYtghpBFjiV8elwvJ88zbR9k
ID69+1IIf8SZiVvSDYN6fudkFhN0AePRq3yXdOycUtCfURisQbwyUm94hCsTUyF+
xqLlsAWYxNFPAcsbrVJDHPh5sQA8yx/0OB0ExOcdcPjDGtYuTnhamD//M9lkwuZb
0inPhfg8/Nzrz0mg/fb5ZEIsqlvE14ezr2YJ3q/QokGurmLgx/ldefv7yWluJloY
xuhZNNHYXofF5xlwOekEVXUgmrjQPc3BPsfuJsq1qZL0hTZONZwq0TkAJscgfMFC
Y5mv2AVfIN8wVGO2fbfq0N0Kv7PRJN01BXu9CIWMBji1PZYfAI5AHxes0JKSxnud
IoakwqnVrGW6LHqF3Ke2aH16UxXHv4byzeeMwr19rdCb3J9Uy7bhtVG+U0o1ni8i
qHKfQbJXKswzovmcYjWB+GTVmKnXmpEFq1xDFwWfjdxTJ5RQ5UZuWEjQ1o2JDLDe
mLjMQphKkR9+EW6a+0Zoaqg3UqsLZ4BUiyr6YrSTXBP8T9PJFkuKeGAHOwZ+21UJ
p0k1AIeH6Jl1/0M4HdlwH8i2yaMdgRoQX35CJ7wKNfGkHS1x1kD81X7m+DprD8Xn
FNBJHibmGgpAS7w8sSxYAhqt2IKSllp2is6lUJn/gVFMwD+DKPGWljm0pRb7gHrD
tWxVuhAW5W6IHM+tfVwsy1vh/oPzuTRhMh5GTGUvRYxI/2wH1GT5ujg9A7pTTSjM
lD6xu25C89VR+0gOsgMeFOLVP/HTll8ELZcoxRUPWAtrMGlLJnFjKAeE2wonsR+X
BhDA6DHQ2yOHvCkXFB8MQFhyPwUk47UrnJ5ODNIWFwRihtFVFa93mgoPFxrggShW
/3AslT060rt2pLvQBFsGAAvcsFvEnYtDGc7mo4ZVVMmUHc7Fht16ucqAhbwfyLio
OK5/Kpn7Th52U7O2NRSrhapvtq8nWpD6sVvT+G+HPlbsK3Dy/zWwDtP0CgJAnxck
154W0ELo3lUzE6YyWof8gf9V0nzp7OJcuWFPC64PtxF1anQQnvwSnhT/pT5XrVGJ
Eb9xjdO6QXULYUYXlH31zOcgizFf4nW7zxr80UVOQfI6e4fKO/8GWkNqx4vUTZaS
yDNwLVzHF/sPAGMaIe/a3a3o59P0JVmamhK7Es8lqc5KTtgMALt+mQKI7XxoSBow
OqFyrzB1jPVIiY/OimHEM3Zme+P8ZGUObB4cOGOZ0YqbJTnFE3ZRF01gL0c1pI3n
Xdaleh5+/JclacGs5fOhA3oloRWkwKdtgTtqEfRw1F/nxuwQR5kDHzvN0D/aqXm3
qtLlXn98FgnU5hQDcgpqISh2m0ct2nXOYuBvJCIJh+QMSzuLb0xXPuqjZX57rimb
QsMAtLMYK2LzAVmfMzWB4SMOoIUVCN2uEuNL7eGWBdqBW8+7L1MjfB+r0aGhoAz7
V19ETcdyFinlj8RIHGroQUTk8/qJd9ZIwMr0DpOC7JURMWv883fxn4/JtYhktDvW
eQ0EE86to2xoovO1StpBWbUNsUF3TQZFBNvfNQ2a302cejva95h0aTo6Zgbs4R8h
0a6ljEGzWR7eD3/yAyCltj+SpoKlRH/+pDPipVKoay0pBn+5K2A4A4g15LYG+jTM
HsvTgjTfEKS+rZ3pnEXB5y/9npdQTdwntisLabT4cc/ehtGhfFfOlEFAfAS275OI
LBtUgOrazx/ii43+qzW4jxnl/X/PDneOag2IIuHPhZDqxUUStTzYAuO2+ngvZJBe
fn1ejkbipv/lpT3KRamiApm/aJX7e5w274z4Qak40Pd8NGeh6EsZ6sL1TOzP4Zra
uQZHBlKNpHL9aShlaGGfWKxR+KhcQX4T38b3I8mtRDxA+8iOn7b2oQj8lJqqlEc8
5D/+9RZqhZ0UVkbL2Ism1v+8wVLbUXZLgrSHR18YWBaf/dRqA2SxxgM6UNjiayjp
jmNaA+E1vus5fRB7fZhQxnR8A18rRdf2dPbuaFl0zN72xy0LGb/UUvhBG3DKo9d0
aWPBAcI33Vu9KM62c5ZiMKTTlY8uFuvg2OFhfrLRBPORuZABdjQtIsQ4fi/baX7Z
9slIe9K4aoZZoUElMVfJpdHbr1jJS5EwVrnajqW2PaWerUUAuLHqQqNgBVOOMT9L
qX3HGO8NrS5WxTGerlDiwyG0Jvz6a8Fys3RVhnyJwesMo5wbC2SJaCy/eQEIGByl
znbuAM44fjClkNt4GjXk1P8/7nXtsyfgrNz77tmIY7QAyXJZDUvBUAnj8uFg8C2K
bXHBXn3taoPr9h7dW1AL0aMlqY9ax6jVYtGH7IWuqve7BbEB8mKDlePEZEWdAZAj
TX7geWxUklssaKFl3HPBO6Fqm34XEy2DxXj2VV4JR7M2mOHEvHEvN1KV37KDrFCU
Ych0RvB5OVgVYMXoeAHb/8r4GEyIzYwJ6SeSe3ZEitdO4Jj2ICVd9+pSJvbMB3C1
tNf2NmSop0ojMYKVyMW6Gl1eKLLpcf9rxxnPygV0YdighcblhzPyx3WSvA4JH+XX
Amdh77K5qHRrWs9LB22PzKD8BaGgQLug2fmlK8/c8D8pj8cTNRaleX+0Ki2qzWhw
5bxXYNY6SmFmqNSj1Pxp0wuJRRXcswCr5yoap190Jl2uazSW6GtiFfunMk0sxdB6
lQUU7CgTsT16mD7QPLu6WIggY9wDzcwlW4YhHzjfhARx3e2GX5OOFL+QQe6jjqdt
BF0s/d8caSOEXDu7E2i6m6Q7Gj5KJK3zq+PkbszYo7owjeJYMrHftu+734F2hOLe
CFBd+UjAhE3kBn0ZEgJxA2rgpFPL0ySG1XaVo/IZ7N3qvBD0BO6PBfJ0CdxPSvtb
SU4J1bhcPIxojOxYM3/HYQQXYNLQ2+DWjVXfPliAxvQLPDON6O/Qx3MZvbJ1tvbO
nmWQnFx4+viTI4Uq3tlgAU0QREafzfOuaWflU/zu9zHs72jz2sxCe2OJKCterwS9
XdkP8pGONI4SnD6mSQAESaDbbQzXD5RMlOsYnI0R9CBvpoNIrfo+qlP3HMsVEWLf
UuVegyVlaNHbk7ExOS1wus7upgz8JmIx6pjjXiD+FrBpBoFUTc735QHsO5ga3W4I
4KY4rG+yBTbEYJYhD0o74YlbzMlp0lB14fgLLLLbrlNRiRkEqphf5uzp5u4wQfIu
SmddCTAS/BtOvStBQv9uItm52SzfNuz/ZC8O2rDmfZ4r3MxEb88yteOxfq/B+cG8
/pMIRATUfd6hij+MX1etZi2ZD6Sd5fnl4wLIKBrH4kiA9vt+K+auNWFN3iox+o6w
e8WPRjDJqe6pqkBq6QFS2rrGW1zE6OhQXcoo2pQjCl1Axd7RgwTpZaMvCjqFFdw4
vIWD4020T9kwKnWv/T12ZnvcPJX+m0AwgSblqGRoD9/xhc8LGvkhyPlpa+ENz/HD
z5nlj9zqY7Ln0drBulrKz7c7yQe1bJWm6YxnMZWA7LF76mKWWkep09omcqZ2b0Ly
8KWW3/JJp+6GkguqVYE+mUZd+W9zXQfwHY21Iafj8uCFDAa5noCvbuHiDO4GM3h/
+LYcZ5ma8KYpwWHUd/QV1uKJwPLMLQPbjGaA2pMUj5f5EPUO2eMYb+yPS1cMqkmj
749rKxaZVsTh97j4J3/r9JtimgBRvD48To/scgebzhQZ9+Dxa5Fivcj3Cx0a1aLS
RLsa8idv7fgrZQeHj9icaKwYBwdZ9h+vQcY1NH5tLJDdhR0xnBDt4AByv5JaOSXT
d6ay6NaIur0RNlc6OFhVyiJigMnJlQVo8iY7LYEHpCnnBCpp1Ti+NkGxcQH7gW5W
fbxfk+9uBaYaqgSf66hyMgGtEfRDLkr+rV2MFPogVVW04gWR5LYLB7BXiR2J9Jbi
ri5Su9/1F+efyx3qyqAsIYla3gyoAGWxV9Q/uGtyUhCP+hsEy5yJ4gPwiUel5NG7
M1KRvvVhqp0x7UJa2TsRwWD4PO4BcDeElxU8pzBpm0e4G3+K+ifmh0tFPx0Av5ih
DiJH2KYwNGpDcJc8JNq9+Dr8vjoHk+yInUqk7rRSrPTyO5DPC8Aq+w3itM7XPAGN
OUZhj7USsAjZGb1u/JI3o1m2esdRdD5i0vU+hRTz0qEJ5dhxcqsDZInMdUhIyGiq
TP9wi4NfQVdxJVgjSSCzapKhz9NN+tKITiRzBFp20c+FzZXn2vcYncxO1hpzwTta
WbauQWyB7tt/e1W7aJmoBhTjR514auPNfiguvRSOjmks4BAcTzCcbr3x/+z0usTr
j3dFDq8b73IRUk6Yggd3Btv4phex06i3MT/hePFdYNFz4dDw9bLtbaVcvdoFboll
Xo8GcebXb1Pz8QUw1o0rZfx7tZPUN6LwaRsewKIy7XRtYNgiPinNymSI76YfnQ0b
hRBA7z2cJXCksqJoqCkrpl9R/2yAaYIuF9NNMrpSMbZf3arxhHXYQbuF/bbEHg8q
rSEiL0zaKZaDDVsHMqLp3kAMBqCUwwxZxL5brhFBwwJ/1kxbMRImZTCRWOVmQ9sY
qlC224zFEEbO4yuV0eIFRI/rMKYDusaSYdMi2D+uq2Wx3Y64FjBkuk6m6JRIcRtD
7YEVkazTxRJf3yArCds8kT4aRGVVxVkY+w8gmyWtfeOxaDljqKEbkctX80R82fqI
TLCtG9YFdw1BwmTNnNBq3V1PsPRxMn5bBI4wScyQ9x9XTPQ/nk3GHaoEnMTnZONU
+HG7S7rKb2kUc9AvicI+SB63g2/3v4jvNR+WsAl/AVTpSeqTRkAI5CcZ1VWoKu4E
Vd/hq3CbAii4FW2dEcB05ez74g13fQkGbtKAIsexj3m2AU7Fxx/dRRkpKlp+axVr
9S3wKdp6So+15yXxqid79Evg4Sag53OVqxai8wjox0CG0iGZ2VfSfoS16FbPVOBO
4qra9tEIajOQfzwOj8CCTL8MtRq1b16KEGL4u6n3cdkeoWn+J9hNW0YyQU8NsMd8
8PHhsZDZJlMH27Ocb9kxNWQC+fNSw809z5aE61lpMctnj7bh0Bkp8nJAVvsSEUvI
cqfn5X6DPn4n+7zSvjtKaC+9RghkWpk8FfaCw/DHUx8p6SZ5v83UiwLyIjy3Fqbf
U5iBjGe/i31MhVK4o4xLQPGqBGF1OUgoB3u9LuuCsf7t77BNKL9UAzscrFEGUZot
qt+U/pYk91pELZmyyOApJ8NvGBqcAr/saZb+PXnp8Sy7K4i8LR5gSxmoK4VoFMY3
RsM4VCPgmUJtvQdbcEN+GQN1IIU0uiWiLeOhCFQPOET7ctsFTdqdWWhQRKYk5HmR
vuS9sv5KTssHH6/HXRpzjW6ck9bQI/BFn2M9OafX4G+IU+P1weozbHzH3Bpsfni7
6D6lotm07lc/jfbxlANheb1ucKnFWIxBsyIeu0lqGHJU1EBzn+jrBX0TBrRUtugP
Yv1o/XsEKyJd+5KCHP9PVCjv9RL358M70duYlsDvpBBJqoQueKpvpIgOQ2fDelwD
y5ojUq324tXUM3F1B13QLlr2EIj/p4fRPb+s0cREI5+WPLsg3tOpGyj2co+Tt/lW
0VtrmJY36ewJg8wk7r0W69AzZ5dEL8KZDXTwo8e3mD1bInETnLB3kLtSezaPMr1K
gF0bRwq+T52vRDGcELYmqA0hQQqtvQRoziuhaAyrlhbrGg6DbFeqYk45NUHLFvrD
41Yw62NAEv5M2KzkBNTLMv+26Hud5y5AKoiXbNLag4rvo7WTbcr9chmme7bAYcJe
fmDqJ2DMQ2AhM9vbelv/27cfrjTs9z3a1/IMWl8uOX2T1Na726W/OKg3kR7Ltra3
dtX/M0donO8NA08cYPwQWHLGPuU648P2JemCLeIZyF8z9TEFfTKQEVN2YZbte9Yj
Aj7s2YninuPT2nzDvlFFPSsvRV5XyhlB3tAkptMkqbBf8Dl+0EmySzcR5RrdN29J
o7nBx0Z3QlTsAccxCGFRkKDFATTHYjtoQhJWn9JuXivNBV3/f4ew8wpVhevrrIIB
DkGtk4+sXFJhxYrOQYVeW/uEqBLeaeTSopGHIDJrv1QSIhnHllY5VtjxAqUo90/S
VmiAJDseV/FkC6PD7eSbz6MRRuxz8EVDIvo6LzMIcebMWK4VPieDNS0X4YtFVKsr
5z4vT8qEvPPiANv7hTRJlHk8xIBI9dPNyST1QdsmMOteayzkIs/jThXKfJb+tv7Z
fYOL+yGu3TAVLac8x+FyW3olDAFWsuVsuANuzV1OSf4yhxj5s3kW16356df41Tsc
jEi7eHZ37LzxZ723HFpvN+ioBb1vSKrZ1rfbJRKWUxb8jdl2GNr87ZFIRxkyuNQl
TxD22Rdz+UF5s783hzyDlH+rALGakQOSKe+VWwWG6cfzcf/jhz/esx/2G/2Wa2n6
sGeX1xApb70MGcV1FntAPSCQYORddLMm62CZDl/1FV+whGVuOGi9OBllvg1Njdn0
V91xe8Pybu9Fyr7eLxoLXNB9KbPGs73LA8I1ao4l9YYBAZkw8tmp3JCd3d2WOn6q
JQSj2dxtYqokUfmtP5pnYan+rzY9rkI3WATiAIaI6wTWkOgV+2du52nE7OE1T9dG
4x6vDg9nrX46YX9vo1VmpoDvqC4CB2EMGhgJz24kOJMMchfY+/lz4pakp4/iTdlH
e/uWWNJ7oDD2s11dwAeV+p/46mJgvPWD0UlLPwlfDZF5i0s46KkyyZqtj9Q7VtI2
4pV8wjeVEOK0dW/dSOQFMz6l9ma4MVyS8qoZSU8tXXvqwbADV/1ka6qqO13olfkq
c2/Tog1hh1G2dmkZEK6Rkb0v6XFJhqnlsALOvLoaFl+fxalUMOpvXLMG/46UNBl4
eD+v0lEsDCMQ8IHBvaC4wewVNRNF+X69TeoP1gIGF4/6hhrMX94eUANTmNXhm9JO
Gg/WdINQBPzxkLK4UjsWjO97sNAON1VSgok1w0OosE/1O8NoYiUVxYPO4E6crQ1N
CQuzlEmPs4KvSoMIyvRtvUoSBfAJOnFzYK/R5GxqZXAMoIaB5isUp27vdDD06njm
X5CT9mv/hkMF0X6UgskD8Xcc9NRk1e+SuZCEbXONLSrAjGfyKV0+hr62XecrheVP
NGAwbTFeOIsIAZQT2tuSXKYUtHQtDnedOsSHPpX85TuKP4DROs3kbfV2OAvNqVyo
u1WnvSfbSlVzM5WzZFJGdGqCrJh93ZQH1+0+KSGy56bUZkinXV1WrRMykwwXeu4z
Rv9OACtXRbe3nL0IW1qfVpeCUZc3cXKSTwtt24EdQEnbABZLiSOhhYuVpAZsRn73
gxrdDUXxLQkPxoOgRSixmwuj178F3reREqFRDHElTkZP7h1YbrRcDOKCDEM2S+BX
IoRtvn/0v6ztGHo5eYsmvgdK1XrKVdJEOALZCYcwkwtyOldxU5H6t4GrEl/1HGOG
i0/YmAJdcaFRz6WcAYPdkcxySgy8ujBsotiBzZxS2cUMKeic8N506hfk8xt1nGcV
dshHJ065V7FIZyx8SbZacbiLG0lRls2ZqhHM4YwFVvkVaMjhbDTd2w8c8HTp2Ceh
wJa5elNBz36auwnRTLkh5ZGM665/FWy26ao6b6z9kMT+i/ImbkqX8ppliRkqW/6K
FZxpGjZIMMnJAKSzeBDobWzqjhlcp3TpPxbbJhU1iIWHEUv2D6d4457lIyvK0pOt
tytPqU7Vt41UVIMLBCG8Bjgik3emmOIjS1dGK+ezTXuGan9ZM/mjKpFC78mTbrI4
9CpCKzAT8wuBru88Zdflpdons8OMW7zs6+EBEcoLeefYNJTV+WVYQvfxZC9jbLwR
e4Qx+/93rzKMgzksA+8T1EhhZc5YbpDU+b9P0SC8oilCZ3H8vUi4Pq2UMvi5QruI
xjfNk+VmxlXlgLwqkQ86u3yCgPc9z1Hhtkir4hTiS+8PoD+cA5NEvAXgKuxoUaQw
v3jkCV4V55dOcrsm3ZBxtGd2iRFFOxGU7vs8yxsWTcklCGx/FGgY6pGEL+VCyylq
iE7XfwuVrxLEZgL/EGvobByT4A6CQVsOJzB8Hc9bPhetgEdvrIeGRKXUpcWokWjp
6AiQ9GdOPrF8z7FE3BrQ8vHZDHQReP+fQx83mZ+3Vde+fFUpN4UCraSFIIvPb22g
+JY6U/JzLEJGv3aNH696hY4zkp2CxFvLFMHa+WaIClxTq11E1z2TVb/UT/Mlwgyj
FGAvnyaJ4HkGCSIT9dwGFaP0kBCecpHcKi7pySu7D85aubD1pKrDIT4eIgXxFus7
+rTsrjjiJdqKHhUV8O7ekZdskRjqdbSoOPydZ6YMpOdhoDWTAXTNx0zDT8G2e/9O
Z7a3G6koURcu7tlAbiMCVGpfXjHX/DnkXCSp9QTbmueRtmmGL06tMpsifUf2wSlb
dljj7xQsvht7c+buNnY5Ilco4bBZNWYzeFzhE7i2ZmIz8XLbRetpUJ7FY5zhIqST
DgcUr02Qkx+LOd3JeCzrVFCP+KeAzC50GbL9YHHUQgSQ9QMBJZBkOezho4RY0lf9
NfLmKdYIC88T34LswRarp89F6C+oOBuvFD0clNm95TsH37JdqlS1+QAnAM3XP8uQ
j1MnwdRLuJZhI5yKi7OGHzibuCfasocAZANu3CypoU/Fr5nB1XTde8XQ6mhImsKi
EPxqX7wJ0PgIk6z0PF2HjudR9vyJlNY6iOZUZh+kS6eSnx/X+mkcAlRL1FYmUn4J
CBRrVqqIfniCmZzP2Je1Pyw3867HGw157iuiEfWM5d3fjzrtqbygHSBG8hOro6D1
S82qtl7XPWAr/9ZYnPwUd+a+THpJtykgFRzFR74STtH246fMibL/clxCp9FM7nx+
5tO6K3eTOz+ZB9eJY+qzilIVx67taOJpiog9tCb9LjNMq6ZJONRv3KorW/CYKq93
DUNuRjpsxITzD9sRiuauBQVzJYw5BO1zeFmrL3l6vRvLwP2pd3cm9Gf2uEuCA/Lt
S44sRiQCu+KJlR+S3QlcDhOdxYlH0Ka+gGAAtF6hu2HVzFp71NiXbezGuhk/bTxY
U8E3m42o9dbKfoMO+tkcRWSEH3TRnbmwdIaM7cXjFmZG2AaHZSQteIXEeY/zumQg
F/DBa/CXIskE+mLut7Wbd+WJ27/96ZEUKs9WBkE2sUNSiuQM2wBcuqMWEbQC4fiL
PzN8UUXh921JgknVwH2jM2Z31icOOH2vLZMGXfM2RyZB845c3O8okyPK3Fmc6Fuv
HuTWnxjAWHxOPkKJdDEtXDNplmgafYCoRgcKTOKXOc+TaWY4zSOeP5PbsuawXmlh
YN7LWkLJCYPOWR29LjkzjPaQiJ1e3uUYKo03WOf5AuUAqJHGXAixPxEfMjxWZX8G
xTFPUial0BdWiM8DkfzDkN0CnDzI6efuyLtGPpMSy02JadN0JewuisOGvE0h0frL
DEmwY9xDQydPdDMEyNmGVLGYjoitXYaXmg7oh7C8Q1ylg2ZwVdlr9zeCckAKqQyC
DzbcnXYz9JfrcLhUowmmiEQfNCf5JOAlRXhC+TMY50gppTVKcgaFixNFOSk0UsjU
kNOXaK9dle1wfCgY/teSIZF4KphYZzgl+lfl4ibG00Z9ia0YJiPg0ko8X/YYhgcN
2fXmIYP+dipLAH1IJMx0wCW8XgBYMG1L4Y2G1cS89XfZt9vSNHd6BdvBoxrByRfh
ZIUHH1LZkHkszahtwWE2gSPis4+sGh3C2gkALeHO4fWz7wSp80rl0O+rFg5b9U8t
OyfsUxMUgj7jxn5UgctuTCOt73XVgD5x/WeiialVsyz6xwdo0XGFGj8f4P3tXltd
inMF5fc3tAMc1JGJ8lCWptotRMRXxOja88JRjalWKhInqEyO7V5hkuICAJEWxa6J
CCTDRJrCeG0hRWmkm+1++H7RAYkPqd/tG/8eacspIJPRpAWauv1/6PfUYDW4LfDd
ZBMMrQt0boJFgabWsHsRZql7cl6Z+WiB1e3rFWAu5mbvYxT/kP1+0DEEFWXsQJ/p
woIO1GAj9s2XbXkQb+2LvWfkin//tQz6yC3GdrskGiEKw+h1RbjKrIOHE+8TgVZg
Jsp23NUqgAg4JgK5ykIlIJbj5m88VT/97XcmyrCLYS1Y5XDmxYyNr6eoCL1Y1PGu
mkS0pvKtUieXqW3p0oq+V6/4GWw/ATwY9M38nVQAemBL1nFOedsLWLZKWUUzjXcE
9dpE7ZPs6Iuj4AzgvOv3Cn2JI6YVqFrJS21KWxnRT+P8wMakrFFFiV8ecJ4TqGKw
3FAs/ZbdtSUfm2Th+f5PzfrzyKWW0P67yN6jM31aUOi7iANTjWdwYqkHNL3fUziW
WJX2HqCHVgC5vAqkdY2EyTUIyMR1J0HGa8JJzNI8nZXJkUBP1f60I5WA6NXJ0PfF
986Ze8WwQsfLkYTM/R6m0SpX5G7qJCgCv03qFGVsf+JekTAri775K+BMPn1faiuG
ebi7UycBCxF1366ME8z12O6sMbG7uPtjXojLokMSatU0h6S8jO9fUT4LqkXQNN9Z
D9zQwy0fvGl+Jfw/ozYggESacAVVsQhmXBiYjpOBseuTX/MkDVIACZoFTjYbx+cY
srXppjTgmN0dMwNX6E9aNPEPIWpAy+ZQIGgaX1r0ZnzKP600reTymXyO4u0tt6b1
0vC+guz4FM3ziZDmv+n42XdSLhTOdT8qisSf3XBdjIQ6wKdgyVN/ySbxRnf/zGUk
gPSjY948RsH/garaz76XScYkALnY/8UWNojgtnAv1VvA4Bzn5fuqyhSRbdglAi++
QTIK40JjU0xryBarmd1n3/fgV/gTNTez+KlZ/d9dZ0Wn+0g6CV3T/NHh4wO/TYa3
3MktQ1wzE4LwYb+8wlVvZFQ43Cefa03hw9w2AMdo1nP+4qd28uJMBp4GQZ7c40DN
1KuMh3EDWY4//RXFwSweGS3GJ7xOYNAV1uqUOpOWPBLnVMdzAdjRMQzGQSKPXtiL
CrHSEkrvYSBwAYBQD3+TDR9H1YN2xSWHdrYkqmoOrY8USZTnw7q97YDMhPfu4I38
EorKjp1TGXfL4F0lt+6KXR4g7FgcGfA85prUELHXLwX4Gm0L8SGN2/jSv6nkpOqQ
yUc+pcMU3S3j0gPSs2kg+48SIyewYw67QR2S/kW34g7ja8/HalLl8HUBaXQkpZKu
lPbm7TyObSs6Y+cU97fpdovfBovJrmDu68cJsaP3jQBjkWrxrNyvJMjiHd9SkGQN
Sr0YHqa880trJHPnrCw2/iPA0QK3JvIQRmBSBgDIAJvsCZtWuMNaW6X4WY+dK3tg
MDgyIYnxI+LKqQ61OPPmAArc2nt+y1EXrtk9URp7qve9e0TtLwrQig8qYQU8c4o+
34E4GtVNMVTslxWiOcGEgIdXf7hOOaSOipyIrHTlYAvTrXdGGfA0+IdCttWn1J18
Rm8gsm5EqWvls4JL4VMT+r/Mj53ySsSgbxQLCuVFCTn75asMspZ6BMiyhcHy62Jd
nNLWNRc0F9/UZXVA+9nRkevcoBZZRnN9koaMzDuXZw66/Mw3QhMhuMbRATXKcDhR
ndvQYN5UK67+pjbYsEaX/0uWmcKjV4qAjBp5il0yfP6U3hrhawzA8bUPafvckGmC
pkXMeB8Y3kwcOOr1AZl2VS9DkH1vzIbohEJIbVySGrmvlc3YxMO3eJRDd7lqtVF7
PEzFriE4Qfkg1YHVNwVlNDHedorwFQcw39HdfzxuT2zNUfuoSIjT1ACpuBJtdCx2
hjJGv1KPIJJbNRpgsWqjcqO7qaLeyY/B/MSyd5A564DD/Lwbpf8qGgOEIptfeD0L
mUjJ3hvOMP+kKoNbZmP9NmL0+3tCo+ip2zSRKzuToHGXlKxHOWegZLDj3I+ILoxQ
f3hb4dPDLbXcgcK4/kdciUE4oqnR77IOlTkpGxVEmpsOSinRmUwA0Judqas7vx9K
EI+RzUecESOMCueBxhTY5nSIsMPOC62w9A5qcqBBWNpZYEF5iCA6pGsnHycqtTVx
d946JNiOf2MC8zPF6s+F4S+UqWY/BdLd1PsTi+ln+JD9EhGazMDjHjtFfDtNVBYP
QcN5Mlaue3XXRBnNmEmxLCKmjyP6yCm0jvSviSRukdZSZlqb7RtKw0Zs8pxNHE2m
jSML25dIR9N9bEkvabUoHw47r1Gy24vXnqty0JwbJTSiFXQ/NyTeU+FB+/L0EBgy
Tq4EOLFoU+nDkfi+izXsi4qEvpay/CC5N5+V/YtYRWwcIyGsjCA+mrpyRxxDqSI7
0Zf4mdOkmf6D/G2+ADFmZ1b3eor0C4BjPWZJLXs3VvkRPo+z3FgAlxxhTN1t/xcx
1gBXtIff86/dW0mp8CcFaFxpxxbxnVnxmBt022jkxfWFiNUhsf5sEppxHFTLFdA1
u0KCLuTb+AUgo1/gkOKhPmQRQDTcrDhFk7Fmo/P74SqGWlEdJdrZ5bX4UYrmrtP2
v00agwBrribBRAAlDBkuHDa9tieNL/avg1SXBVTlnYtx0bCZdspLuSACAM+OaMZS
W9VJPgLrieK53Kt22LjrChHYeNOQ9xmFUVDjRWxq7Wmpza2IjoynUfQvLU3lzd06
2oiKM5/kNEcsPJX145oUiCIOvU4cJw3+Zd+wbJ+RJKhpOqJ3wIowC2ooLOGM0EFb
XtPyWLJ11dGO5PB3y53Tr3T/PLLgoDxC/r3iDQAMuMgt74CguH08JpqaZWRzfvwH
z4z0gxRXcfR+Wv8SyQIXHmiL49mIXfiZvz5COjKDtu0Hitap6iVFnbch/yEKuUaB
zHcAutt5YU6nnd6cH6XWqgFcGa8ArGUTslOTCI+rCliesa8ND0JIjIo00ldxh5S1
ZpEXMC+G6NbicSmEI78ZyFfj/NcDaxqiONOK3VW1tC4Y3/I3w6APHmpXEHgULEqL
KtFuAkNLrnkZSy/6eZ2bFM2AI4ChhZsrJ5IzVikNeAY9WNyYHhrdQc8Uj4qHlDah
PWkc8Y+281HrMZ4dJXat+5yy8yQ0TtH5SWcdJ3MkS9ygNX384ajH6xykVtjN0AiQ
uWLsesNFZSypOL8X3+0XUVj5jtUeMqFYu51I6ktrEGZDPo70BgYMrI2j+XJ03BNn
t9bk+FB2L6DzycZSHgBt0D+KhsaX7nCY9AfSFDctJEj+OcEyixM41I9JnJmWVELP
hR3JSUhwSveJ41wCSM3auTPCwnP4RSiELeFRVA/touRAhazXc1UuQXI7REjmM7O9
h7DnQ/frZD3e0WAA8+zKytknCARVwU/0LLRIIPtKSvqLwhHaUqudIT/5g7S/Ut13
Vr+wCv1jjjvpC14isaqh+HQ2t/6Jc2RlKLQpubvaMASySEOh5hmb6zgn5PUIf6G+
U/b8+Jn+onbC14bGtCinI7aKAIboWgrjGmT60POVWCQBLsrrretXyqJL6NO4iWri
32Jl37vu/jb4K5N9xmBPsWHUPBVBFWyotPWPyk7Rv5RwAnHJ+CBeuAa2yMYYJKqs
GI5cpWYE1XYLqC8bESWJA3IrTSltrFnMemyOjB2pyw25j2hHMYjJnlM51HOFXMLX
gheL1NIdv+TK5NrLm5yhNjBVRe2mwmV8rIF6xlkkaT6zjucUffkKgGc6n1eeSKWs
kaWdsEWj0eFbU7N82PAJsAIQaxyrrYSQb5U9SrzyrcqNsOp/3mq/4NxW9YDKw9e7
Ad9wbxII30FnpfrhyXaxAEjQEvMh9vp2HkkAJ4lDSJo80D8Z25zjLfX9V7dsLArD
A8GJ8cfdNP21q/2CXNmbwq/EfF1wLZW3R+PcNympZbI2zUyF1tOn80cupnd5fkMG
1zqlTxXdGem+1HdYi1VkrSba8fVyViHp2qqO76VaNRJTcDzabLw3QkZEKhxnfvGw
oIPUSejTLkdEJTz5HnCuvP5y8CptWFD60b3vDG8EnGQDqJ6xosFTR/4vH2ON86o8
maZf7yWfK79oRpSyA/HQ0fMmK9lxlLCbCdTwy6DHt1YZaTqk6dM55vN/fTTyEffA
CViylrIvUvibyBR5Hv1pGPYBwKJNVNWzibFyYo9DErdI9LFS/KWvvvTDnqrPDXwR
/jbQEkWClx1eltnS+2sxUR9m4KD7L/nKhqRr+us7lJPbCdZfgzeig79Juun1vjPf
alSkA34XeMJVyGBo1mzrfS6mlvzfy9uDjxaGMOlQqBGIV/yXVfNlCK2aqF/yvNnA
jVrv76MaVPgxwiQoU+4tnGCDc5TcjfsCdjkdct12g6qqt+THK16BD53azkTLYWc4
FQ2+sGwiUUKi8OPsvLflxxfNThsRGnkzQ81Uw5rPCSDvCo4uI/flhkrvqyRvAJID
3fjeOLRYyymP0X0+ukdbei1lnCxWNiYU3OFGqtzX1Ie3mfHR/2kwGiNeBF6YFk/X
NUhlUTQhrwym7uTnrFVvWfg/EVE0O1nvSik6XVGR4x6wQ6ueZNg2VueyOHOwL7JE
K4q0yJl5IFgUFSL2hHOH8ujXDvNZtqtq7lY2bMNtUGJp2RqnoySm6mG7jLzZczA1
mbtpiHtNVrigAl8UYXK2BXps3giFtPbYQzdBbtJegDcPbOjoEyJJjZUeGjTG9SBe
YlPZD9YJmTLrUXfc3t6m/39xrFmwREImpEnShvCvr+hY7M1X/uspvD0R7UvOHxej
b0Cp6iizcuCjK9uLkA/TnQLUNAEfNsFqBSdC5Na2SQ353OQHg/JaFS/Uf60bx5XH
oyPybr8qrbD5zXCSsC5XI3YvgAbOWU0teK9P+RAWeKG7MdZNlOHJNIde6hJbWJsY
U1FlEfQkmNK9bWxmQs8zD8Xo+Ca6mBLfG4+yuMkFeyx+Enoesl4lJGPvKRKyM4UQ
g8RLrPcJUePXVlJEFE1Tc8V21PtzrSidgpouZcv7NbhnAVau+O22StcNXw4ig/Vy
jUnC/J90z7oUn5in3TFsWr2TOn13Pt87FyK2SHNoAWhHV063MqvQXj0AThsPX/qQ
ShDwP1Mc4PO287Kdq2A/A7mjEb5tTQTiurdcJ3ncenLkU/IAcA54Er21jMZRRjdZ
fSov//Wa2j8Ffk3+YEfAh16yf5ReX4QfgJM4b7hxxwxzhsbW/f1JuSbekZ5zcryB
i5V8yAmAR9hQO3ZtH4TLRjmucpZYH/bY8bTrmkpyn7hYfdvHd16eLjza6pXg4RhH
8p1HNSB2ATr5yd5rRn04V8L95ao+aPfgx4LsFCfBdkoZlYtFMjWYJwXLT4nW6J2o
RfM6qL4vgTlOWTGtwzZoyIWYbglDChbFaWjAhPNagY7YztIWItKhnz//ZQg7/Cjy
nODMzuhYKD2YaEwpZaR+RsqshhSA8Br0oVxNdUsuj4o25L1g9C0zBAjObiKQpIU1
7Zt1PHEo6FgOY2YQMRvmx2FEdrS8dvlxS022/rSethv1uUIxfwCwLB1iSWuXobww
GVrEcmo9lCqVehwO6fKTM4FNBWneRNO2gTXAgEdxZ+y9OnS025O0jalsPVGgUkEE
ZH5oDXtc8N80ycHd2fH+BWi3WX0ckzUWLyqskLJ81PlCn9Dh1HBfwug58aTCCR7+
W1UZIozeDjmOGMSRhB98J9fLiauOY/BA9rp64LPH0g6l37cNaPEXga5J91T2rhiM
hKN9ERtFnBybYv6lQ/bFsODsCg54EHR4zRGGiZUsJNljbcQK+8ErXzV5g+MluWad
nsHbi+cMegZFzsUjlXHvGckdzs8ihYUY8mjkMC8roz5wWff7VjH/sY3pKvEBhEpo
4bdp2mQbllZ9ZbzW4oFxyrKEilyPriHLQi5h1xurwltmfMBL51gH3zLrcaeqAqg+
qBdZnF2YlHSdk8VdweNFye/esjfLARi2Si5yF2XLmRWE81d0AbMw9aegUDYGDKnZ
qbecT0piHrxdgf4hT9Wb/V8qZALCtOUl2+VuCVKLbYyVVItRGcqqz0MiNbLqoFbW
WhcAfF/IaqJAKCy42sEfQA+lswGQ4VJ9V/N6C4W+YsI7Ud9S2KhfS3CZQ6KJ0gtH
xjRGPVD4xyqpog7YjXXWA3vpzfrabsjcmPwcVvNKs2eaFVX2Qjz1AZDmGt1j7xtT
yXkeEnEx6XazSS/UcQCqKT3T2pI1s1zX0LPSUrNxeccC45dGagjuKrH8a8gLBTt6
vFOwnGtKEmJW6jPusBbaWg0GTJvrShd9DRUz14GuSJN8ynAXJTpsqDfp2Y+Mbgft
J/y+Q357k6BOR4Q3W7t6LRb2wagAMUmYRfIyVLwFxuBvKPQfYu4AbR52wxLcAXck
tL92GkTeZGd5CX9qLnJA06XzE1bY+ysm1Ww54pgnlytfM3Nf/u5kJu7GEqpShGfK
HAmK3Npxr+sqec/8FD00ZKGUS9fvd4ErC7wnTAKunPai4aKuxD4yyodtSNSdfzI6
giaH7BvJ/iz69j0y/hC+0PQfU3dhhjWAul5mygghqlp1yxDqNzVXTfo4cN6bUw2P
fx4Ok7PaKVMB/Yx02Eefda6aUuaC6JQ0jPnri39Bsgn3HwtJT+S/KK529dIxzAbQ
QT0H6lqirYWlYYhlWpskV2euPn2haG+HSjZjkQXegztJBENsfP3HB2uYQ/TFYNGq
xLFw7l3BbvvyJ/fCfyVUMoI9pQhgjIi8q7fOZ/xzAtgt9k8fAuBRIwDEElB7Tx2u
w2oBkYz5Pdiv2mDge0XNAwxk9r2Fg3pzsBMtPrCLhLH88oLZWS2l0h9QQB3ILVjf
VRFDc8vum99PjruUDBCqzv14kMBIGYOlT/b4UP6B3vLx7Q354pbPidWlK1SjYNVS
nmkMkJ8XPQeX479u8gvxB9Wm2TxKkMct+90HsPtC/C2gPVc6Bbe8rDvT2962fCoC
vsr+vf4d5aJsPt+HSd2WjzQDec7yI6IdHa8ZPquza3rheOpeAk+2yISuzunIb7DR
e7YOouYIcbsHyHercuCeeFlL80im1/irhhColxj2874Oq/t6q/Kf6k0ptAA2X7JC
7wFrL17oPS9HwDCmULbM9fD7JcrGIv/0Yk63MPrhmP6dJTlz45QjQVCvp/7TMB2m
Pn1cu7BqvDTU/bljziH7pYa4qsluYelpkfMy4YOKqQ1MjG/WU68MmqjTmOvPRa5M
+E2O04Tc5jAOW1VPTx9PPOWuZKkJjvanUD/y3UzPBtQnjPuS9gRw2hDeH2OU/iTd
rdIpiwrDNaSaUXcLtstafuu6Y6mN3v6eGU1AmFNgg4sv7FeY2Uc3IC+xwnq7GHLg
CiOKq7pf5Aa2tARUtfCmuN+FAiRugjPdR+R7gcmmf3TKFCFsTMGksSSpXxVnPd4F
v+g040bgfJCF5wK+yS6MZMreh2E73iJ/7RzPJ1nDXnDAnMmYNFSMdd2wbHMkVMHu
T3K4Br6bA5nT17OJqECh2Ww2LQWI2daRzLNlSw+eowHuTGQZ/wwGPovN6xFTm6MQ
ehQF1cA3x69A7JsymhdPRscOIh0N5wZctFFyBYKTvHEl6R2Ynox1GECJyPv1RWQt
rv24MWmsB/hN4w15err6UA/sDa+PZSmGX7YHJ9Zz5VDPEu86lGed1T+AfDUJqAuD
ji7k8Ovu/7lW+lriZFEE8EdV5Dnbfu6lSvts2FLHMlPYbs41fazo+3vX2Saws2wc
fIEFnYaO4BJrZSWAxuT4sZ3ccbhOgsONxkKomkO0ehMYlzUEBYrHw+cENwjCMrQ+
/jEwD9NnVdZgH5p0zi8UkFGXwLEOp588qYIyKfoubnuREfhjz/TZ07cDequxpEMi
mPxTo1xaVOA53C1xVjsiCPBRSEZCJcaQ27b2yDptasoFGmtlePXTTpGICleKmI15
cBou8DmtGeCLXiMOUHMxngqd/o02xmUPeWnQ3uCO8QEZcklbFL4n8DxF5/+qVsy9
SYqqWOiwcuQJGZrnTqiNQeHDZjsx8NVbBq6r+Pzqq8QLkKPNQOSxwnCgES9P0Ix9
2sUMES73CTwZQjIzIdg0VqFVfAQ78TKm31S4WTWD8Dp87UYKreWHK3zP83jPRT12
MDwaikZjwF2XAdZnYvfNcQ6KE/H+kRFWOVG2HzwXwTUr63aMxhVmPEAjN3rkPxlH
nt42sEYR/1cWf4lmhly+22y5H/BEjsAJL9uxuN8ZGtp4YsE6UD945yfAnvDFTrWD
HRlAY0HsRN/qCILPOcjNEnf+emZCaTmKq2yG56OYf7GyYeu8UICTAOHUNg+RqJiw
TkP4ff2Uwg8+XgBxrIu5S306eO7BZReDMaN6NJWUHZ/kJpOQZBLm97mXapRhmfnk
uTvIKvDHwJeno2bACnqkmzXHjboKUTzwtn1PXQYyUuLYBt8Vo3PXiVGIoso3QbDz
6dPiasiQ4AoTh/AK8XKiODmCXdrynNnJjxXLoZBFjQMcJqNGmQXmlJdMN8/9Zk/9
6biO0aVuzJGVVr0pKM2daYlE1Q8v9kszMru70U3MUC7mnImndYTc9GnHK+SyQF+O
+EW5xeRwbwDtgoMF6yP9QfL3mjlX/WTKGzFF9DcaJxVpykFKtixTSMen35SYBFx+
J464x24iA652cWGFikqPMy5rf0xynEksN+vbXheYbOqjHn8wOIgXOElT0SrbW8Aa
n04TX/q8TfITMmnKYEqb0OrGsBCWBfysuo3uZsl0mBQAIWiJQUdYbkQrn+6Pcfuf
oKD+229zGL6DqmdhNc2VPnRt1irWBhdUSY+E7F3Q0Qr5Dr1ugoNqyr7Hx0d3Ne+g
R3x3R4wQrcdlRGJmV7ryVUDa1jPqYqYNYdakPHLcQjqbQy8mZ+ejMfquCagcmtyM
GANPDOAzDZmcXaq+wW03lQRb9BuIDL3CbGvRhFDlwaYB/tKWJrsIGkfHc0ZbeB0Z
qFFYSv2ZcoATTlW1tCirCXjCoqT8thQPArrwR6K7Cx33nQvx0xkv7Nl2j4QrXx7k
10i9DycfTi3ZlVDK/9N9hRZUbR4+Oyx/DDaerYUky9CF9XzoYTw5ZvuTC0w/G1rx
dbVlq90PKKCbNDvzYxzoRPJKD/d9uuh9r1YPBcMRO0yKX8KwyxxEgV10eIKDIZyA
hoHdmXM7sUdUPHCYSFrnsBQz3T9ueYeyNqgL6sXC/PmiMcaOCDWVh0zPTvhp+qSM
4dxedJZwNJLavh7oiNuh9TayGJe9jA25cTcuDfzMvXKAa3qXFzQYI+RL0UAe9bNS
RGLtSgzR648TRxWF9qPTdJahfVjMB5eO2MZ9pdIEb/kzksk0DXztrCZCpgNNSbo9
G7PVX7ugj/iWCcMn5YgROeW7B00XMmlkcZ1wrNiaVRzLzfP0dPB1Qty6Ji5Bxpvg
f+TULk+Ci/rIkoTny0F8EpgSxHlgJnm2P8ER5/M1iBLLzjhl7wOOWmin+SaRZ8Id
fWcBW2c4NrzWDR7efiS4tHTSN3k9/iJMnEqhz6u3mper2Vf8r2v4NL1RB5VLSuKi
BiSR61prIZivd9MF3U9f4GuVBmxCspLqjQ+c44vXEFtJS1ZbD7u483hReF2YMH93
lZp4XgnkwL3Zdin+qXwQYrfnJHOcI+8oYqtNFzdbotwoBefq9Huv5rFacUDNkApf
H9QAQh7gx0bbRP3DJPSiJqPNSbaCrsWExqIKyOwK9cZuLKyeIydRhpYieh8+AuBK
i2pHNE5O8g1uyc5IvBaQwmvVkmucMz0czKsuR7k5ZKrTGQ4TRB953gys3hs+h4Q9
r6mGm0BvqufyA3giDXvr3lBuPrv2kcK4QPdPVHkUa3ZzOqCM441h9i4f/0rrZp1+
vSuoGawnzbeHJOa/K6xRhylYvlDXBNFpRRiHGUbiy6jx3rBTEb6FVWinIO4i6ThH
XFt+odVfkykxQI0k15SlEcM5p3pq+cUfTePdKibM/ZM3kXojqK1Ud/lfHVL9XtP5
++VkOg/GdUsthgpuERxN8835CaHBFvUmJKqKoo4R554iWEui7qwR5PEKZjLVnvmv
sPlm2wwBAyTssVP06cJ7NnM7CywIDA0F0UQbzhoytj6O5ylUNDZPnLWGZeHpviAz
YTPFXIMxBJsTeo6Mqq60PUugygBtM/hFg9IXVDwuUYHN+Qk1RTWkschTgpnbD6nW
PYWikrX1EYhgK635whPfw+rQmFvyaM6nP1X5+Jm4HaKkVsKsFG4ehRUD6EwZstzN
IkagatMCBVAFd8Oz/8KhKT6lVuYGeLeRsDeeQjP8KBgCk6sE8NVIwVicKjQCx7Dh
sKxstTRPtfYwK7fuwNvZT+2sCN9oGTNTLnIaHuSP1EnXJOc/TRyTt0NX7WJrcywc
G1BO3ObIQDdJj1rC2nRV6uTFF6nSy5tD91+t7xUqfnAqReSCAOKBiguJ+u0wav6D
tmWDW/Ru7j5GGbx4QB53QmZpo23Yv5/Sk4XQwm70/+niVv7cXgZvfhhK3ShCpRB6
SrJhKmOVyZWjenLyNelQib0vHAaBA/JxHW3n+z5qjua0w2ANrmOi2CpECF3/OCk2
1dCs+GwxKn1hK3EpDjrg9HMjPd67UEUAmQQAueb2u2u9FSMbfSVxEaQxrXpolPFr
+GguVj77X0SCb1q1G7ubYBj1v43GTI60ArFv8P+nNvW2NNd085oBoRBztxyQP4Ii
XRnHbzj4kW6hQ1mL9vxIticOwb5l6rYhjGqPFdajUMF/U3tXAscNf8e5VKKayFy4
Y+LgoMhJGW8q+Vf1YsLJTTkwhfjj9FHwjX5mmg9PheUpBJe+JT481SsVlb6P77RA
cYv2vr6l2cYlH3HFl6qa0VUnPBFgTjY7VYR+pYCCu+GPd762ZjZT4EH9SqSrpN06
3LqMrRCvtmiPkc5Zv2byjb9J8Skf9a2FNbO+eDdXUuAHlmLrd8RccSAPX6qgSfSR
Ucquk05GRV9WP3Ys95+2opl7pIgkl5iHFJFPP0j00xw+hJ/IVdb9YRBIaraDSQ9/
teh3/jZKlGuWTAN58HQtNebPtOT0GGUaQwvQw+8ZrFtqQdoyo2ozM7VTZR0fAu1A
Lznysr+n6oIM2vA/as5/yKM4xRHvYoQk05MAK6Av18EJFWCVie+sDcgD7uq72P4b
h/ABZWPQDvi/xwJZqEu+7j64YsnyEVLbOfh3paLHgQbrlgK3ARfXe02Lv8FNGhop
jTTk8V4ECOSEpJZZG6rY9owRLTzG1PE24PHEC80kbvLHKVtxY+6OHgYBjEv+xkGP
HumbzOsWM4jZZaxRH57v6dDhp8jHAmr7Qa/m1coXp1oUJGVCnc/iNEzsv94gpoac
8bXZnlH7oUKYDKM5+NeAzcBRxlsL3U0XxusiHDrIKZO6+pnsk8ah1WoBTzlX0/Xd
/TNjAKTaKicyxpS9x2jObkZN4TAtldhi9tVIDbOy2XizcUVVgbt1kDpG2I4cFz/A
cmAouRrNAl6+PDWXQw1AgtRzjO/djpVo3YFe5TdDvvWnu/VLuAuFPr4L6tqARDCa
UtMvZ+jYTxzd3vJYegmE3g0i4bbPF5X4taMuHovnMA6Ty5kTGvKaabUlVXuOqV/K
qiiTXa8raJw315VgWvUDYzX/SkiXWHEEE4EfJD6jImNWHUQ4AacypOTqbTmhhYBr
ONXpQM5qO/EKmyYGneKl14uSbHGLbX9dATPlKBUxNVVsaw8B3gSDIb1r4s3cvw/P
dfxMElRdie38xO8M0mP35ZRTbj2fiLcdG8sogrcUD1ikQxasV7dLA6HdXqzgjqZu
MLTMfO1h/snUZtjaPv0YcAP+jaXjje5xFVGbnj7ByR2so82lY2uaamSVi8KWRAjE
ywrKjUC66jH6Q7qcPikTSiALQk22a0oLJIudZ1WunMFRjksyR/BsA/HG8LtbRd7I
LOyWDLuHyYEaxU5FVo7KMFsBJ18wIkUbabdHri44tH+qQDdyULhaa0qsottutCWT
QmwCG4RaDVbsQUNAs3De8zP+TeVkW1LD12Y/aE9cqNicZlE5/0WqT7XOTawnIDrP
ijuErNxElNw8z0DT/qGVaLz14XtM3OUiN0jS0kxyWPVWZunvENQAoPruW6JLffj2
pVp8vdyu/of96/SVdxnnAAU9kcx8V9JA354tuvkr+7wE6kARDQwWDJSMkz9Yo6bZ
uxO+55MyXYFUgrPkPhkx0y7nsl50sZc5z9riTOQnxLNPQgj9ixTN1yNwY9V2FktU
r6ZkdM0TVuDElyK5d3bx4tHVpY1xejG88lSrNrvKJDbCeD+HBn4rFu+7p4YsZ2JE
o5k9O4UFyOXln37yekEgihamy6uhvTU3nqHRdhAmXXGQbxqMK2gBbqhgOof2s0Ow
u0tO+qtAUfgkg1ux7z/IaF0tS/CewaiH0OuL3OsyWUJaL6SSWvtRzV7ZLs03fVkI
nfCtyVD1wSZCVwlZsfrtv6cphxH09pE/MSfuX16reYtAHpi/m+03fc3jTcXC3NxM
bN3iykXo3100QeLekNOtw5aF471hUc5VgfPG3n9VSz2Eep80gwhLsJ8MyLnzdvWA
rbpdPTy9ywvIhj7vdK1X9Y7KFlL43si1r/kkoOfRIeeb4KZLDSPyB4jOiqhreSc8
/28NiTc4zu1TpbKa+kRxhRlJ9o5lsXsDcjy9CmGPHvXYMX4GyuwNrMXEKW7ZhgaT
2ejsayVRXpTU+xeFyXDBAMCg863KKQ+kMMGF/gWtqkB+ZC2MlwIwEdIxuuc1W+ty
m4Xx4IaWiMrIOyv96grWrK3kVY18bLWh8VKVfN258JgSEb27DhUC0UqmYcjaJ3+x
IwZYvv8jft0JO7Sm+98f1/M8UoF6XGSQaN+UoOkq2fdkDXwZc3Xe7MAXURd2Ijxq
1BT8w4mK3h3U/kjtfMaAYcKB243hsX7NQvDlLAD0Be8zzrG4tcO2AEcNxKxPrvmd
NeIiOe41yyyQMbETxDS4Gv4/rvuQMQvWy1kBKZUQtG0HmheZ29VEPd69jEqgTFhi
8GOdHC9VUp4L1X7dWdKVCTz5SBhbrUIaklAKo+QUU2BHUKuXUIsgNy5Sd3JX0gnN
tPrfhBP1X4Bkwn1kA/a0jP9GLoe0xveMHYQ4lcC59gtCsS4gfEQ5aO8IGucg3o97
/jS+Rz8rIeelcwOHoWs6tKCfE11iXJF3q4gteGG1MGwh1z/vWI85sqtYJdzl65NU
RQwf3YaMXFcnxQwXS914Kit1NmCcXd5wA4q7y248YOEnHCHbrCooYoDZFaYamjU1
Tkc2Bw+OCnmkDKncgZ3VD69FbgZoniF8wwSSctK3zZgDb0yqqFZ4Ynn8wCdf5jTQ
rXtvXHckMBpHfnXYo+x+ggEEVlQYH7hSMuVDs6c39VxJrtOrHpQvmWePipFLkO6p
vhhjABbcg0AMZpVOjnUdKR/Roc6JUkKCZRFy7onHvaro4nbw5m3PG6ONAI/5alcA
YkYhO8JNV3WQSZfOEy5uBPEYtLEAllUSMzUWvc6EMIY8u16MfbflDsXPgSeVf+v3
wuPk403/SDcFNqwXSf/CnGP04vtjafRZSD7GSG7N7rHJJvIe9pOcYPG2iia2E0TW
8UZzztnAzzlwTsXPQMTQ8gXe8CwrdOdMTglkKpOqu+LpLXvEwIRSwESqpYIKdOjr
1Fum2eFUDJb7pcTTj70tO7Kpdyu3mE3RlHDUcaVCrtvWABXl1VrBFkEHE6iqOjs6
+e0GCIKFT0r5p4CS21uvy3d4RGtYf/EFzsP19apGKMPpyEWit7w9LOUT5Ng2o/6t
IiLj/UcFIZXb8LjXJ2mm+zfhJu+ZlUQ8aHRicXGSnRscQCeEVR0+nReMlDu9Fq1g
rMrQI3UbMWy+4UtBNUvZxV7EBI+5tkRojAgizkiE6jZ/q4zmyK7go4s2md/y2VeC
fjJB0OG9eiFXh3J1nDiSw2U9qsRZ4IcGXZIYpz+fsBLIK1s3e/9q6d6/Y2rfXKOO
zGcax+X08uZpqy0Ru0dFgMycV/3FLIIAWns+nk+NDKKF83F50tifacO2xMM7jV/u
mRwAVXm0ouM+yERoxhzt/r37y6tdwL/Rb82UdU8cOasweadC3UHlAp2L5PzIY6YN
xOMoCz8hSwWj0jzI82lqvmpYqpFyVtQLH1PP5rY0k7SvGldnFwIKHxkcVGj/GuD5
F7bG247JehXcNn1yfVcV45fuuvZHmLF4H7Df5JYCL+bikFK1hb8iJlpGQwEVVxTK
1nEMcrudcfcy/nvDqxWYMGkkKGq8JRXALvILv4jp1Gg5CbbQa55tnUYx0qv1FcxY
yMX5PqGt9iyfeN9a7ALJyHQrxELWbH54vMkkuqmATLAE2FtbkHjAOLIUs6hRSQod
IznzWK4q9QIFl0oB+Ri8q5BVGNxmJXokjXuHgxq4uwsye/jpD7O/Tb9qo+ohtubv
au7OGlYtDpN6RBhzfYoBL3c+BqV+L8CtICdvXpnOXZfVi1AAuBWv7hSIkBCBGi8b
VnsDYVbjy6DTnwROMc53xQUJOXQUoRuEKlMjz5/BfPmDa8mReZv6dXk5pFvD5wAk
UOW0YJHXSE6qQsSPV6PD/PZrI1lNLy+9bRDkyxqeGxNnheEuJjS9V60ajLsfq3/l
YCeV1b+FPy1YRIFHaoS7DMp+j2w4q2aa/yj8kywfCSSWK0PH0UCYF/jtHD0yieCP
YUsCZmSOCdyICYQsKlpAxhtGbEdR5On1/PrqJjczxfymPwHLCFE/QzVzl1fKhpmt
2lsAgy0vFla0ge3OQ1T8HvxOGLWGkptxGFGxvOcUy/ekxfnhRoiD4BQQsTepzzau
AEBxadbjVKNwKzBSar1Tc5QNE4qPsrbY/gBuKVQ1qr/6ROLGGyzBas5gWhfr22KW
WjviXSP3SoNUN2b0/ZacWvFo7U4k32Z+KZaAhtz9zP+gDBeoGgMQRIcALYQ0ifec
dmhgH3BV0UInUsePKRVg5oqwrHqRqKrqq8UwcSaorkWbAy8G3Xb0v0Z7umoGM8XX
uxN1BokbO05Jy4F1JWs/C80DmCRXdV1G8Pw/xaEIleyy0gzUPeQO79bZZgmyyUSZ
bBvxTOqwkc0ZfFGNVGHLJGhHSLiqKAdQTKw1pVXZhw+RtJ24QwE5M7eGognasCcq
2DuFyPYH6qBMw3Y0mV3DH3WstUWZ4Elkc71mMLws2cLDZZN2ZWUjypGTSsALCZM4
aHN1lB38JJ1f78+8inNveaYhoKPzB089YmzWl3HEiNw/co9usz7FQ3YXTuy1hej2
bqdxdLUFr9OQUbxDgR/P+rC4px+lzMOhc1wxb9EuyJTUotNELI5QDfXSNnOxo4PR
qp2Ma54JaFU8gewUJ0/B8RPVeo5w6QhEZbOvm6AI8e5XQ7QYFZXzqoQhGlza8fz1
BKxG9qq3nHKf0f87+2+MHhoY8xucd6Q4y7XCZ32EWefA08NF7swWLMU7dJ2bHGnv
UsLRYbBe8nUuwIVtrC2WcVNdqWim+j5z4JkvcpwjZbUTeGkJprU7uEYoyDko3q9D
TFAcwIuzO0HswWLbxAUGMKuoW0iI55k2B6sQhoDlWOOF389gmlvWz+MiU61/wQpf
WBMOiXyDNjRaZsw/l8/3KBwKaEhkPa1CvUeDEiirwg2OgV7T2YiS1F6DfL7p6T38
hmmuvJ/giMSuYBvBIN5U2grlBGx4icVFJr2TxWuD43Ka3M2coEMKqw3Fa6H0MSJs
dfNHUxB24qW8xtyqIlrdOp2/XjSgHppMKUdT+hN25+hCNfnr3DDfZlJw9w/el8Id
+gpo0De3yz0vQcC+94TxuLq0r/VkZ9t4Sj2bQM8z++9oi8Morr2COPPWZgHUWVle
WAym9jy/8PnqLmmdf/nCJoYEY+CJhbnXc/GlE0gjXJJTTV5SYpWqE02/P7m2vcz8
CzDRgDi9WCbWtm9DIV3+uTOPB3EU7mvy388woZekO1NicUSGhs5y0B5q7Yl3uSxT
U9aqoc4hhvR+hAH2r5ze1TNIpBYV1HzF+zDw6/ryocykVgAh93mUzEDNK17wr9xL
4Bk05r5qBejdmAgR+3l9TX2+5iqnIfcbJPN2Z+rIJf6jtWm+6e6I7Z9JSPXBIWp5
RUu8l4okwcb/9Ly6zCVbIWHOmpmBrm/8bVQqelqA5wi1Cnum4mX/ak16eEfEk3GL
w6dp457LnGryRYvjffWfJGMb9RgbFXcci9eiCPYnDT8x+fVWNShi3noi+x3SUHIF
PI3ih1L8IKACBj5gqjZ+1vKNe+EGvAfjnafghsi14PbRRGpJ/N4zL7HZ69nSZQ3W
3vhQcCcilWbaroDrOBUDtUzbfkcnwaL6NzvgPDIv8keK8DwIYYCxm2XsF34/5fWH
UKt21UdRld0okhxBVnC7nKFFSil6VV9iZYscfDBC2ed4VVs2G8smH06Ads5ghTVc
sgfrYMydWR6AtP64hp11NNRYJ7cFY+uhvxwfyeEG1YiMUPiTX+t7SbR5kqhbceJX
2nz6H4cvmkAsBl0TCAX7aG3VbzsFRO0J/Fb7jhp9wnJtitjdc9hEtuGOxmoCRNft
oi56m15LhSCYYtpUEkec2QTrVwHNGc5cB2SWPIAfxq6KoxkYbc8iaWBU2ANhTQLn
MCa8JiO6G2OFMbILOOsIaYy5LSVNBj8gZuTCH9SPkiHRDjYuZqgpw+iMYqJ3XJx2
7ishagcnLwfYcCXeDzBHTgjO7ePUM9edThJBCl0mYhlfdHt6lFuehjETIJ2yoEgq
x3Ux11CSyzntRcgcdKmv3JjySWfbGpiIA8bA88JknK4QSWTH7t2Ac54GELzgmsrN
iMLzb475hsKzMXW6K+KHRHtTr8HWE3us2JEplxolYsSLHIhs6Yh7GXNVQ5SRmFEF
/3yWP3v3N/LD7dYDbEVSZYbtJsIDY4qLjfn77xNmocn8Z6sgdFZCf05N5QI4NkoO
6qsHm9Vv1Us93qczPP4O8uGRu02/EMmjOmDDvFyAzVpPrB/f3uD2KadhRCrqsTI5
d/T/K3p79r+rsUi6k0WDayeKv9i0lMQszenLhgVg8JOvbiyj0ecBwvDI6AIGsw5p
lq+5C0+QJAH/rK8HQTFWaCr0usnM2bqzhycWbzX9EnJ6AWui+TbDy9nEgDinaREU
PMwqF+Xzpwdy9PLE0t9HrMdqtjwYDvufKdtpXqKVY4socGSYsb77WUtTTPJAgfxv
BP8h1ezNQrhLae9voicb8O0J+ABHvoJYI1KXqHX19x5eR9dVNUji+bsDdf+Utu0l
yTn4SOb5Xu4VIZbNn+fyDAMCfl0FAcMclFnUwSFhq6nvrwZnT1VOmMeHiVWDUHxn
J8Yb1hpa1pLUoaY6GimZvPnWUIYbNtrg53GoQAfaYPHpBzuYfhyoua0vChe5S4ck
LoR0kkkxTVlLmKxwGslDDfZ5/jc0/FkEFmfn9aYLyZuIVYEu0rA8+/iFQMqSbco5
HVRMLcP/PsMfi29QfnJFeMN3vw421BtuhT4UkKMZni7TBz6fn3l/ueB8/CkiAlMp
uWZOMejvH5IPiNgk5iyGba0x+WGIQzajeGBzLpbWkdzCV9OSPqFZLXJ/4gXDjRDw
Ttwgfuq3I5q5Gmxvvt0WwtnhjCXInCen6/mou38QCk3HvulCVc21cBy/HOn//zyg
tRwEQTcpFLduc6AHgPfPp8xcPLv7FbW5+NqnoQW4mf3i236WhrxVAxzR+ZGDIHId
t6TF3vchWrabt1soOSQsS/07Ep5j/asgMOKW+cWh+GlzzFLccN63HwiVvOEWvHFv
3Gv6w6yMKr886AAukvt++rxLhszkdzPoxxm3Ai2DCNzFKpgsjITlBXdraA906CrK
NbMZeOvTNCsC2OqiPGsWXtQjZY/Z1G6KXmJZjXZCoklMdjHcAioT1Pte31C7z0hW
WAShpE9bNyKleLrGHPksFuzXSAAIgTOS+XOkGrBJZ+6TwCslxmik2kZTwKEGxu+J
7mMgsVPIYMbSVK2PeKtDTstLMarLSCmw3gSNDjPXPm8bQBFd39b3Ou+Bs5GyDKSK
SW07DOLKxYpHZdH/98SJrjt8PsF4YlQspYciopP5ASyAi6f1sgUNJSo9SK7LP0tm
VemMvcSygW2qj8nwfJ0UmXSFjav9BCwHVxzjIO1EUJDWeZwevjWH8pYM/5so1xhq
qKWmDDXd1Lm2fL1Pz1ahW0vBKn0cA/A0t+i09LpTiJgSFS9cMQ9yfkahNwIp7R1c
Q3wfhPasAFEeHXXov6oNLvupQHwuajj7pMqNVoWx5EpwBXSGTcxN5ZZRI5U6pucE
JWzGuVhFqY3aeSB70yQCSiRJJk0tNmYlkYkI8nbkUaBhDe41/h+DWLQk7Jwga9H/
7wFEfB0XVflQGAdj6sBzgoy3JJmS085VwzgVL5Q+E2tBoJvv6qS6QaGY/KO7Cwgv
Rq5lSzNfS+ViOmZqf/gxSRz14Pw9LOFhvT8sppqNPP8KGYltfSWPu8JMbFPqKCHm
TufYtRY9MfwE9QZtxOMxSfOygZiF6WdWoNYZnIhwBh0qS01YrdkflGo21ghzSOUD
hqwAE19bzH9uOprSoqhUCtva1UwDI34lsC1W//eBUzGs92MICE3Hc7YmO2pys3Fv
mjx7mur0kZWapCniw8zzkchGiOE1x8Mq+T6zAXEno7AP1oDk5qNt1/lAmVyW9wOa
hg6hfIBhNmQQUIkBzMCHykK7UbMvnFrN8WHqtS3CfLV8NhstgpL68rUPrqFCWM0Q
du5kJfYI81Q9O/rC/BiLBU3pEwhxDLSeP4n+F6Yy16OXrT1UCSNxMyEhATyW0fow
dDwWg5HWZZefSZ8mPQagIc41xXoLUU32jY87hay3cqKb1hJRzXkV2q85JokQHyrI
rs7zkNPN51sg17b/ercObo7vcCDfphPc5r0Rp3YVQUHQCWyghDd+++D3/Gd6ADez
Os30yYfN/lvbvJr+XAOqA1AIkF6DSPYqEonbyOEV8LI/13CZnfseA4FWiLlYXGK1
mu0TeXla0frdzfPQ1eHEyBXaEgCbfyU261f/wsmgWds/CnknnL5fiJ//MhhPsSif
5f1VJMi/wn2xoR1vvjZ5PNXT4kwOi9n585T0zy1QntTdPUO0aheDrEMbrsOuj0SF
AHQl+yAeNySF8BQQVMBLnieMvzVS+egUPUB9vVmlK2RBkqa7Vy9nE9BCFjA3geGs
ioBKWE2Ymp2BjTJHI7m6ucIy4IkS1TlE8m1oMomL/kbFqm2zjg6Oz+MHwsXEoDVy
zH1Dh5TMtx6wza8sQSnZI2Can49UPiETEuZvbis/qndZB63bQM9lqr4tYJXSY+/2
U9J3Gv+HwLnHgg5d16UwyVu9vBKZqcOVaSwDyW9iQ7QCGx1F+SjmvoUWJzuOewLK
k2KczmNIwOrRtNpQthzR3kcJFIT0dugiL3lPTTl0I9MjXAntd2ofdEmcBGiR5a/x
3MH0lUdqt4BSGhyuPACm1qXUJLR3y+T/EXe+Gqsjsm7BUxbPs7irsxQmper0GirB
ZtvOxhrUMa34uRQdB/3cPCkQgkAeudfXTpKRTPvqF3g6yDZ0M5GSoMwDVl4cnE1i
pGL2DvcPqcJ1rrL+mMA3mqsu/z14CUzIDysFkP+QetVKlFBqHwyj6UfUFa6D+bxH
D9TFneFh21eLJvpCritRNxITtjQP8dwCvnVzR1M9X92Gzucsx0jE+ApDRSKXYdiF
8Mkw83c6dxPaPj1PF++aG/erSnsTOKKPuXtFPgf8lO7AyMWzlUy8DLZLTFZ88rmw
BYczg6xpc8sYo7YDbwHezm/cQYGKgXXeb0CHURPa7DSeoS3L2JE/8gkumQm5KekS
l1RxYxvLdO3Ho6Ap2RRP/oSSox7ekXyDcZefmVld5ynoyyyi+bbjbjDCqz+2wuKI
Mpr7O8aDzxTr2mnxu67fZ3bXuMY+9q+IxcNgh+Xb48GKah3RiRRERs1qXY+N65Ix
0BHg3jKNn3BD4pW5H+vu9WmegJgEwusx8apwzghfiLJuodPvF1iTskVfulRNUZ+5
onsm6+d3+d+J0SKYkbOJqQrdRVIW5Z3nlsVM90DyNAV3447wfTLS89tWyn6O47JY
y5QRLZywjgZjuzjhjwhXDS9Y9PoBeSgPoBLfzjoLqr7efnce8V/EstSVr/aEHffj
5RUuCPnTCFGKyNcQMUDoC3gdo76xeUNhdWf37yCPvThK8+nzfz8YnhV3nAyplmgc
Rfk4zl2CLpfwAowbmRCZr8Eqf+XlLplGmICoxlzYn+UBqD91vs1sxF0EqfNMdgrj
gSvzSm09H6cQ7YKtWzke2CWvGEPqoyHGy6O8Ke3eKTTa7EFFrBbTGIrLRN/5K9El
k4yq85cEpod7NcziauenDlxStM+yL9tsupmXMeuHJ+esXBdGjdVh/WyzVoARR1A+
0deorxzvMTo1tJ5Ejcy4+KYLkRQy7gD9ekiGkF7BQ6VqIKvkMVC3K40D4XUHVkou
nTZvGAfGznynBgnP2TmPPKpexa25He8IN2/k5XR95qb4XfN7I4K2BePMB7ThBdXR
2hsHzXw1S8h8SiboXwlUJDWZXJEB3P95bM1xTgsVLJKG+NC9UfBe1CJn7OPb+Lp5
/oHe25G11WyWeB6LeZyjOyZWrbyHhjar2RTXmrT6zWXzQ1vSoq2tJtrcy4/Utngm
RYYULiKo2sGJtO7DUiYO8T+bIMdHBFb+4vtG0c9AKGLHv2S8PnQSJE5VqBCZXfv6
ZtjGR6ZvImvjQ4nXaTqOTzflAxgbyUaLgRx8kxaZCiJAopqP7F1Wz8xG9HLTXRZf
YimzK1DME4ppNehwH75zgrXaUXSyvJXmICtVoIobNM08gyEuXHTNsAll/YMN+xJK
GjGAUvXe9oMq8hmZ4Fn+WhopCy1SunoN2vP++z/uNFzNVvzqmV1GjPdSHfNGT/jA
w3g1ZTn9nnZEpzj2egP5UIp9XPGu/V7op8g8BIpPJgOD1FLHCHrnRoWeGXYQAvdQ
VBLaA8DBbAt94k8rfbX6UudtLCEZQBML+ICCV+MO88Ci8GRZo9JeXxCaIHbVPp1l
VN3PSVaSV9Q/XX6TUyM6f2goCrL9tAhC67068wKjAAAqv8hEzLv5n0A14AF4o/sy
OyvGKOfOWAoYfOpHdYSbjdv7sEW59oGHhT0tHFQgB5vIe5rI/sDiUZu4DJmIo6Ze
MUH9YFBNg1r78gTjj17dwxPGQu18Q47o3c2XdO2pZS6xNvztfrAyzmOthq7s28aC
P8ANyPq0zvPJLCarEmz9xHZ0LhP0DagnfkQjeaB37j1P8uhk3sbJ4XFyEaudysjQ
DCVO2t9BE7ErCiSMoYJVBrNWgmW0LLNTwKWxZqok3DKGt/WgZSpKdalEfv50CpYR
f8iXMlwWmhXxYM2i/kmHOPya4ZAWXV6/e/slVpovGbHkliC1ugG0rfAGgkbwFdyb
pOYEu5QDmwv604hIvN4ICA3Szkqg3TGr3qy++ejnxLLqzC6m3I1wGBS0xYiCwn1S
YPpkFXCcMrdv2r91+lvXQxY8pqOkE5PtzLzVba0/nGhqBshJKQvCu/SlTglkD8Cg
XF5arzjVrZzCsyK67BzT9wvPX/Ma6qPoXUPGaXJ6wH9y4Eo+Qov0zeFXXAp8+wuw
fQvNYBMfcQW1A9TnBfVHh0Fn6ayLt+e4nygeAaStixu1U/3UfVX5PKBltdC7Ai8j
Vc3Z/GPRz5OQJFs3zh4idMNn99pSkB/bwHUW9mLiRwz2QJydrFenzc3QWk4dQ2f5
uhKkTXvUz0QRXHDRfvzMKxett75Yxk6u2GE2kdHMytzuFXNo+f3hWoI8m91CVOdV
STvEYPvAQZFzNlYoz+aX769CCU6+7E1lr3kAbZ06DfDnV92cmk0HEh1uQiBh0ySq
Bxkjg7QEhZCUsHSxJQJwp1AjM9YgJ3ZvO4STFHQ9FKpQ44jLYRNa1ejlCF0LU/gH
w/lH5bo4K/9cTBC7YEFLdsKVblNs6lIIulM8AwrlzVHyhHtnoxXUI4f2p32CWkoQ
NHElBNgi8kKl/VHLU8oYmQQVMytXt6SmYiYhjXIa9Cz6l0oau+J1TS4Wf8up0yn8
hZgowT0f3f0OnwRwCqbtNOJq7c4uY09o35KdyfYSDxI6iE2M7I2KXZFoqFwWIMvg
ooQj+V2UXCxpHY/Fl3zqL1SChbOFKEksqtukQLP4dj1s+TG+losBBG6Lna2+yQW0
38bDK/YshTM2+3SqpgGNbyiEMIQxjl+DCKEbVX7wEyyO4I6TjOo9EOalre65oazO
CbtI/Pvx1+/SUlpZqUj8+nHsVvPRhPLJzC1bWUWyAPzrwxyGwtaY36FGZs9Nl4cC
P2NIDRojobsZfx2gI4+cW49DpKgznf5ihLmdQx99vRZiQy2HKKlc58G9frh+FoGN
3oCePiGu64NWyqRbm4cicvgJDmgrRu6Iq0izGsMHtacKavnCWpLv46rzQwfnpZj1
+G9WtARXRCw8TgZEXWD4i9tNsrjW8EdO1g3e+3SArPOT38gSeldKteW1Df9nvpp+
wID6ViYYLp6OLUTWPtypn3MlaIA1LlftdnaIMmTAlCARyK5K50VAMmDQtlb4Z46/
5RBPHva/yum9qhIR+gmJgrq1Mbxs0Wuh/amW2ixm1neH9uL4sZft+VcEWNRbVkHU
oJgl6P9p3X2V6qrj4jKPjlygclEMB851yRQHHBgSnDgei77An1CIaCxIQafTlQ3S
e5mNq+R868XpniCJtizPoot6mTToNJyrInYdrfvztMqBPo8YfD0Xfg1/+jUV6TmE
cpx0YS7JalWjU+TXyKVIHu/PDrnrwMu8GLAtltxAN5J09ISxI8TDv5vJI6CKhCxX
VPtECPvSxhil57/YyVWqY0VQiR0ScoQNlp49BIUKD7AIzpm2xw1ceVVngft4QaIZ
PwZYyQ3MK/YE7u++4jC84vvhCxsdt1aQUY5mKN4La77jwZdtodm5nwo4u+F+7UgB
Vl8zkmgcUu5txs4sf+KfUiOCvcbICT6c3LFXIHjUSdBSKEqmj12xPoOhqwf5YAEX
EJ8OBl2/MGpdBQevmF8i/uY19hVesiDCOPQqpTpr6e8qisTEUXoAEbUoH9/WX4hl
mJkIUHt5wgCc6dFlAzRH4MhjiRNw7IqAc2EkhssCsShzxPCU1t/So96wQXFxj/bN
eNAXPxLuH+oIglcX85A98ltfkY+kK8R4zP0uO85kQ4gmIgW5DR+zCOctvmdOnfCj
NuEkyJkCQQMWIsEWQky8Er7LFtUaikSQKBMoQ77JNkQ+ahwY0vr7rEV14Lerhk2i
naT9TtI68e/SHNAJTxyd670jXL+eW7M4CA4Dxi2ovzlIGF8//sTnRKu+BWQqRCtx
y0+SjHZdoG40JKGbVfWwBXls/hTt9KqOq1yGDvv+Km8HhTcVknnkyGIFJzeD9cRV
To/rIxtnvO9c6cH28RXNFolMF7ZbbNok9abz9eS1VMUrVQPmTcVDoyhZgKjGeC+r
Sf8V2uprVpCg6+vd7jisOdwiXGm/PHGoxeGGpcTyZzAlFfp572ZTapiZfNCXtN+m
5c5wLXH+mqaXSkwSV+qP4VkGAoB5qRyxRxmvbft/VbU4nLSd3zjZ/+Yz3232FzNB
lYLCj0a5vlwPoQqLl0Enn2SU2mztmXO2v4Ye5usSS6umav3jiIaE/PV98grsrRhL
ll/hNKMf/7LexcrdhQR2cymECpZKJtAJ8ieJcvo7oqHKev9eg9gpq2cUdnSZFuBD
HU6hOVDHRpnGSgs6rzofOc6aK20clI5yE7dId/ZoW/loQesmBSKIUx2rY2NiWC8K
F/XlG3XxwH6KwbX6gnkUlJhaxQykAZRjAvZOYgw3rzmKBAa5JC6J0mqqxFRGnceB
LpMvaNpDuicduwDxr+4zL+F3IXN+35MsBzsDU1gSbmVNYtl68ViiofZPXk+OqXxs
zKxVpNFtGeLPlYL0TuQxntpIjIwiNP45NslEcMELdJ3Q2Nohkql8uOjgm0PkdiKb
+y+QSfpJcch0fJkuUVmaJIQIEmG0ZMuCOvRcTh9roetd6HGS+4j/d6IKOdx5FvBj
ICy8oZCD7nVurkawfc1dg2MkgmRBtW3YKNUrp+W4FMyCRyuOFAAOOhZ6ujlRkc4g
EbKLyguS/muhYPr6yRm+rUjzLu5Aak6cgKAe6eB17xk7CVt+wYlcrIg15qVjaUST
bSIdRhRGc1F4s6aSwmns7myOWaPi4bn+ovBO5NbuUn/5LW2pmqdu7Ya2dldH4TIb
BAKiPSeRq29q7ibzlS0H+3nPoDTX3VeW2EESR1N2J8OSDxHL5Ctol8+bYRuUK8YZ
JPbskdp3MCFF3jmVpQ8DVfHrZhbPKlt/vMAqY094rmGjm5DyOGf8z1gxDLWZbPlD
EPyx6rZDA5C1bxGNxxB5tf2SI1SRB1KTkQ6M522j1sRyXoCJzbmOHxOLAMzSlSuG
XtcPASCjnTplpHuoteR12+MDXREqsa2bVvueahIVPJnkX8/khzLc/71pOYassOkY
uCu2zLgKL4tjy+pjMTjyTcSHuDfevRpmifhIxV0pLVti9jD+PITlNtkFQqggv7cN
XmhK4ZvbBU9oVeSMhhB6XrMMgNQo44UspEBCnLZMH1ZGBDTffFw+BhEC2eA3stL4
jDaI4pUf2Ql6Jf5Gj/bCOJxOn3kl4g3MPuf8sCWHtG4dZKN5CUt3MQMmZUlu/xYK
bhFUYilwtOfiV1NU6wzzAaLvfuRbNrcAwo+7JZLI5fcJpbpvlUO9U2tcV3IfNyqa
aJgusjCGZ57u2UDkPx79Koy4AWzI4g7mV784NQJEnknDv82NTAuOgFJgEnw9AjtM
hoLl8cprTZHvzn4kkqu1RDxT5n42YOT8qdl0i9SD+D6b0Mi4Zhq+Cch67vXkv9wC
yYDxi84wEPxTi9hAiu2XV4ZA5rUBdGI0Cs26bOk5CvreuH1+P1t84Sydd//VSxK3
2JvWDNaN0N6ZbzqTenVyc10lBBiQKStKQkSNB2Qj9e2HJ5T5KPuD/FqODBQA/0QD
mHuH11Fe0Q2pGCSiU1CavIrJ6vZMkJVeIpP+kEmC28v1iyU5c0flTYq7lm4qZ2rH
NZL9i75rZjmxN6Qoufekj0b6yLfquEfPn9Irff3jUFyGYCNvM57osYRNBdbtIxL/
h+JV89T7DR0aMVmW4nzn12V42H9escCdj7DpQggmkDf9V8u0dVEWgUN/AQpapY4c
hP+c4BpS7Iu5qvuXjtGp+GR56feiMEPi3tL2xRxSnvafqRaR6N2rutwt9zFKxX+1
kK28wLdU/7as6I8eIDTc2nwTCGZLFEPcEP9xyP+RGucV7t8MZxDzfTg81kx61npE
YIhIKyAisoTln0ByAIQJrSqt0CYT6Tm7gIf6QX8RzBo8VSn9sDv22gqnXdbX0AOV
/zvRsEkIdyxlY+Bc3+zfDKrafdMBdxaCVJLuuz93TR23ZxeNcWJegmqDZOIcqSqW
Iwn4eFvPeMkOve0yRRcOLiSFeXW3MZhbSHkjqRiIVI/fDzJga/aEjOiNkDglYyyM
pBhbBij4SLQhIL//hFqlM/X/pJ8Zbhepn5dDuH3AoaSbwJOe5I7fJt/msPXlXaB+
7jxI/K491vQG6wc5qwymkk+N++g/vgMVFqV9TTh1mWJmZQRk3zAWicA1ahECubiz
mI7LZGRiiTyMsxePDxY4uq6u3kIboYQ5Zdt8nJB9L+2bIsnJh/JITSPhnIvNugGK
+5ewHlBvyseIC5Ip2FCySGO2okrGUn3MH1vfLikc20RkKyRs6NHdfnTIB+71OxHK
RDBi2J0JLS0ajiPTITkcfbBaVI3sXfEqmtn4OicuKVLp+183FBiCxKGDMmCL+fvG
5Z8UuwkDNjYrDIzLjM8kJL+dXf0cWpvJneQExIe3kH6KQ1S3H7F++VUn+IN8pEvu
5fCp1uoEqRDuKEz4YVAAKmZKJg81psXxS7ftkO0EvpmvPdoAXs8s1mb1JWba5uQ1
AJUd3zliw/oWdpYaTo6UJLFF4AgTnZY8wrJ9AN6wrrcFxno3T3ZTAWgjdZJcxsVI
2thGTK5A8g96lejjumJQJqTEiSewCf6HoywaK6+fpAwSLJ9blM4Eq2UDofmtnVn+
0miaLSd91GBbgWVaWphI6DJRSh4opgPtDPZwANMHWYnCHkFgYbZlpsKT2mewPSpY
b/OhfzeBqXT7uVzb6gSdEjMvuAbLglnnl76ObL+nBfjqfcEvu6EtVGHIyZwVwhzI
9uM7velHW2qvUmzzTRPk2saMVzj4fCwhCnLh90zoPIpuz3lEy8OUMHkbfLCcCpKL
/D4KZJvwJJOo4W0gof2l3ZgOEf5hFInVdmfI5WehglIXULf3eG/W7z3UpGDGp/oC
W7tVSzC4X7hKaqoD5HQ3HnpvbL/auEAQkIaGNAxxshscgtFp9G+efLZ0xBIXQPD7
KejURtEKQoBizPnjwzWh7WkywEx5jyCGOi2BxDaH67RR+Vh2FAJ0JelFPMgJyUSM
P22HCHwY8XKhdLhCEgPHjH+XdbNHEuII5L9ZuMvvO6LbnvtCYfshxT41EoJ7GZfe
osxrGjJSQeE8xtyWZpGC4F3TzkGz0q7S5bdLXsc4QKjRdIf9pm8zJtGZFG9LIEtn
c9w5JInjNxT2Ad+NXeye1qmEZaDm8gsRAPfMs98dq/3Rd/LAfBxVIud6ldW0e1O+
YMRdX30im/Z0y6KBPKqm+6gPFTIfDGnltPIBFBxeX6XwNpJGiMN6dbNpGRsb1h3S
QqLVXHAcbezLXlgCvbGAXh+7iTvLMszESaIyRgG4LGm/Wv1GgA2JwztRMmVsbuqs
OB8S/bQF29UucDzdOOhe770hrAG8cQNDyv+g+IIYeudMeli5LSm6qja470Tz0ILk
Sjhy8g1ofFhbo+4DeCqXevWTv/SjupNcstgN3InYNf1Ms/p4N9K+MmD7FvrS9+jc
vusI+AbHrEa+MMPaV+CdH4PgeEc+dX0/uyWQOXk4uzJartb7ZY1VSD/J05t7TQVq
egSpkzY2ffE8K2YgyfJkM8HptqUk+niYUmYSESAezXYdHEWmj6uwt61vYvGf0Raw
LqL0dkok2qb1vZD1QN3ppYP/WXbwZ1igrYhYLDQRqszp5y4R+ziDd527jfSza9cj
W+DT9v1jk+5TTYUc7ApT8mJOvy4kNR+HintB1Ly8KNA2lyPBj0suq6kWpRBoc2LJ
ZX7zL71mISpK1sLAO4PMDHP8jNH0o0P8n3gMEchAQd5sDrDv0WffNay5e3OXqvAl
KMG8+6ijCR5Govz7dL2NzF7Y4c1M0KwV2jewxGE/CHEL4RSOl8NUVI8Vw8YQ+woD
qKb6CSMH5XQHvluHV4cKz7JAk0hBdTdxJqeGHRzD7USypsDUaVuRpgKcFuxm3uEZ
uEqSomFMV4I0hm6tP3paG2qKMZIbGCI8DXMwl0dQXYOP0HobxzlfomOMzRP6W+YX
VnjxC3t2D97zAs69bLCvh66142ENE5yaf+YlYM09ciAV9vL8B8Ma31JUAjeWFiei
coL2ozms0QAAoE5XY148zFYOaKR7V6VY8Cl+oOnN8OAtv7ylObuWjQzMzvJ7YMQS
OoPuwoZTB7sn0Em7aP2Itf1tMy6QwNOHCObDmPUwyngiO7HcHxgWif9tcr2Z17ir
YYdljlb+mbYIS+45um+n7uEq553Fh59TqWdsVwDJD00HqPiLLAPxoXugD+8Sp/8i
eb6mj3c4XMLDpd22C8cdwaC40/bJvujL7WOD0xvhu4u88lAUc1kLWSF0TE0ZUHWr
CnaMpYStaS9D5PKoUXDwN42O60ettRVMfLtcz/HvJoq9qwH/fXCqokO7EhMOOPm0
r9YivaOJ0rsZDKhDFVUFo5KizYWrLctuiZdarwn9P1YQs9IDXPWu+gzPDzD5Xbdp
LWKrOLBI90PzS33WfQY+3Y8WouDyURmiz/fQDhVfOi0UdnVpooxb6G/renWYhDhC
xoi8vl37sSVoEA21Jvmub/UAh3KpFO+acdw6Yp/j2sUenCPBxto4JP2nDy3j7/56
WA96wcpAZIz4hIwOccoLDspZzKYmctBb7JN1h48NMtatm30nHsVT3aWpBrlMR/q/
ZLN83yVQGF5voXcmFs5+ruo7IbjSOlYUWiqgWRDDcG0PGf9eZKaH3aZwp1YSZSzz
7+fBqNdCmp02t7B5HHUiqexaMLgYi48JLw5MmbQqP0WZJDIek9qLr7m/JVeDWaZL
AVEtr27wUfMmhQubk/5VKrPUAWoGg6twblTQlFNhCIXegu9d82gaJDlOtUPwHGR4
vx0GZxIKvfL3wMucoYvA8UktxmVJV8D66bUAIFlemrkmcOQ9AI4arBI7TGc9GbjZ
PkBkBPiJb3jplSJryeBTTdxgxOY1xccdSl1wFGndSNEHZT0DhEO1Ckhafu1IWJGA
XJ8SLlZA2kuPc7BHkbhPo+U65RolRWHKzRGweyLqDGY=
`protect END_PROTECTED
