`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+TujfA8jx1bfrExty+wChSaLjY5RM+pMv2waUEk5pAExLhY5VHSSgAvNtDP7Try
CnNz4F+BRFpEW2agpLnBuOm30jXvPG1U/Af1kgSo4Zm8DzRc1TXm07/Ff0FWMHk6
25nSJBsKCcBHA/KpPyTvWDqRuVxIDBdnUebIOUVxR6D9X+/aqTGePx0PwHr1BeAd
/pvEZ0t9AnSTfbvHAdlOz99lRkThLHwROWN0TJIG4ImehcGEYG92WZdE8LIVkhsQ
q4/ieOoBnnzarnVjUTHC4UsGAF+fofvMDUiXZScaDz96uzR4kTvqYoPNuhvUB9qX
0zynXVGHlOYqVdUktBZUYCDc/itqp9MJzdD0xxAmjPsZJO3SupBvhRZq3Eua/M5S
E3MEshAWZGtthvqGKgoXhF/Px4rVx3Y7DNJcRNcmB8qSHNMy5nhFL3A7xAsxhm9/
5fI3TVXxMp8ULRSs60Fa//bSJnlDWNuhiTHGavuuGHJdlUqBYYdSuJGkqOrzWdwZ
x6oihyLy5ZGoGGotUOO0Lu1ucZMz7encH8rn2YUO5ltyfJoxqRx6Pd1re+NzAFUP
fGED9byof6ClXO1/MU+VFb+h978SMnpj73+rM7dZloyJpyENrYa+A5D2D0vlJ8UE
St1Lytn/hmmMpoY/jRbFt5DkUMiBy40+PT8Yr4vkY4aKv0nxRlqbb/sbg5Bk5AQl
cqtp82OBWwoBbcCKpi9SZOuLmCdFD5FygLNOcgkKJnMpxbRGMYVo9baFy7+QSEfl
WLdaeL0Xdz3NXf9CcmfYCvBjENDHKdS8ZTtnfMwQwBqtojQ6/X3P2D3wytn/Mlqe
mgA9c+truusf/U/V21FqrEQyRfTTa5vScMcAjxnRM6JoWCp3rzPUSWU67O563Sga
JwFqtoxrK7Bg3lRL8IOGOq4pJysImWtJvoYSXkXtmTGMGZ36+rbbDt/qnWnA3l2H
qpDOIokB7VdCEVlxTxdoC9SVWvRIKwagBaIYy+myGy5QoudnMROEux5lfF9h7ugo
qTMxGNktG34enzo0pD/5CgWnQCasA0JQ9dsPdkxCAvMX/HD2c/JhZknvmk/1Vu6B
iTp8clM+P5WkoHqNuMasrG05jQI2GWa7Col67tk6bw8uXcCKBym9BcBeJcqtnGzt
PWikUYbtzMtmQQuhMORdRIBBh1Uf3YnjS+rZkRwumavDMcNNRSdEjkwNhw+skhE7
BXQq78v/yGBIKHyvVg9MZUWxS9AU7iZwxdDhxXvfX4MgMILtjh3kdRvRnzR0eETi
faN8k3g180s/PuRgK1m+8NlM/JZJpDwKsURU6V1xUN9JA2RxcTxcp++cBZWJfjJl
BZqlDqAo+wa6E7FgmzSAOqGnCcjqRuGdmhvhiYEfkvYrse8x15FQhvZJmsvsoG69
tLbLpoqY/vnXmlLyLyYbn+2K/+/RrnjBThdXSjybqpcoSOxKHFpIvtX2p8Pkj2Ub
kwRjpfZAnyTotmmCrNM83ibktYLii1XE3QS5qAWu3SgMGVFqofx7PdoAKHVkob9x
zsseVconCXSgxcFH6cejI4YjM60eYfNbXeb4ulXee9tBA92uQvHmHHJCpqOOAiOe
6YTDJb88rIwS6B0Qq5M4WBEEKsypsKkaNH4pAQxPW2Z4HFn715zOixIp7PRJZAMI
9JOGWT7SC7aJT1UVPn6ep9X4RlReWjHpgKl47faeQYTusUSt3tFe+fDp8SNHeFmt
9X3FNZ/hI0Yzi00ui9C7AkizQRBbaJccivAPQkHN0SaicMU7u4aAV8fARrb+LbIn
6zkWkZQgS3cYaYvXcMwti2Px48bJ86OGZYn37XVT4JGx6D0181+QHE76Y3ly0Yge
mqHpzAAsSFGSv4lOf0Rpyrnews+pTWcoy82Pga2pgvV7J16CJrJj6bnMGUHT6Jgz
nnYcljEdQkdlDAccZcWgb9JQr81ZXdMPx4e7mUzMzizJWSBJZSN553ORt/16vPkP
S+fLE4ohpaV1x2X1Lwr6vIMkpP5LG7V0FxfGOxNKu5c/qBQ85G+BiCtSkcvhfHtq
tH71pAr+Nh+31pHzO5VLf9DXOq2ti0zPjWuINPfxzMzF2RMteXWxWZdXAYyuSa0z
dXfLO58Si/XtRNGIvaM7vx+24PemJep9VsBbd8jWqspyHSXTNUuwWP/IP8Nz7aGl
3T3UJxxUQOQ/f1HiKoxKGyECdgTpEz2OqiC+DxF4wn9KBPljKd1tPvAgC2HenYEw
jcSmFWELqmqxyKVSX6qfvnIngvAhHL6dC2qEny1QMHQ5/hh6IMgXEK2rPHusACea
DojotGrUbiW6WAA3TD9dI/b5sZQiR9rRnhJ9CDZ/chYFC7saX7kWOSGP+uvIxq+i
OFv+w7hvQJrdPow6hld/uofFJSifPNxZL/U4Hz1IQ/QSrpNJ1GZTYZv0VQNboqOT
4gC45eHUD5mj4NNCUkg3Qgw+G3h5hu0TT+vmLSWwQIP6OmQM7wb+UQACmZWULaCj
bT0xVu+eprDUWCNu7imdSIw9Nboo2XRm7Pr4v19njT8gAvNqifKr1p9TAWLvX3JG
fUd5DGD+9YDg79Z42fwYokGW4ylsx8etvrY5Omu0ovWm8jzNUHk9RJsjc3n3l1ns
GrID9FM7h971q4BDpn5JCC9uWz0Rg9cRM0rVD84oVrIMN9U8C9KpD4uvYiMF2/1V
xJ97+StpwizqNzc6MIc5j9H6GNbGMYoJ3f+MTwAVuwXDjzMITblrf6YMB0egBSTH
YZ+zRr4CLGIetNS61GcddNaC7OWy2V9qNZujD0LdluFIQeebmfCQi8f8wvGlS6Ln
w1WCKemZUlSguJ/ldexwy3rBghmYJ95FWR66lvgqkNEVthvElSNu9VJ28tqUWfOD
xyzKJOUShj7CKx6FmN1Mcf5KskMmPF7ztm3CnaD2tYiddOQaATKD/P1KzHekBU6s
XOhmNtIv9/v036vJbkhtWLcGVUXgGTvlcb5rfjeNr2GDb3giRZvWNWCgb2Jjf2o2
bBd/LuMKPYJo+3t/mQwN3Reu08ufZFHpFp4To/U31Yduc4NT02zlQqENq8rrC0gI
3MGtaRxSFvhWdqdH//B9Xfyvb6Z03bqbFzF7bnTegbN3zk1NSEstvl81nOIyXJBq
icwQRmdADKj9upCHpl11BuR8xBpQW7WSJJ2ahJTk8ZOHwlEH8oHqiDzyuxG98qzo
tydvPz2pQH81jt5nGcZI1+3A73Kx70tp6lxy/h54qO863ykpJqydDFXLRRccE5Ra
INX0/EObi7SX46mF7Ot6Uiu0ffH9m3o4RFBYj9grBW3iAjEvZD5J9uRfhxB4AP8S
REUzfVwn31VPHSIy/aoukKDnr50SBaMgDtizFGa3dPoaxymg3v9OW1ylPm2Ut+zr
noGg2bJrlHq1qB307FJbm3n+1w2Iuzky013KN1HTam0rx91e4MTG0ypuNtvUSdYU
sqVH8klnTaGB5nrIBr2epBmBdeHyNReWHxl5a1U2qcHZ6yqbIZU5lHpv3FXrEQZx
ITN9StXJbpUEGs1pl6cHZsG3Co+39KyfGGje3XKoGnHpRxZQ6WdQ/7Eui+LWvnz5
5HYnbIU5MN/Rst4h/aqBY+esMJkSYegFAX7djbuZu60V8c+bEkXDtZMfn4JWfxm+
UiG5NOYZ+25lZCW36vF5SOblEiJnoJ5lV0GYGz7wvxgBboGSvUy7q3+CRUfMO7ba
dO/dMtZKyrMpFE/h+DnAfF6BHPNDgYmb05GX5JGMh/QHSS705dygLlw2x/2J0Exg
YxV/AXYrS0SP70372hfer+LGUXKnuGGFCh3qRH7fKiABusEcWbvLtnHcn7nRoX5Y
8mOkZZw7MXMjwjfwVQBeRcubypDG86crgEdIxpuXg/BQRPYb7ScFsm94fEJpSLWD
S/L3kTG/y4zcvhFNcIJk8KQ2WmuHlAqImj5HaDILPwaIOk5gNTVkHGhsWNeDr0Ut
dVbeuE9bJLThzrR/krIzP2usHkOB3XB5f1cW2o+2rcFq/s6xMSHVuUHcJlTnLWuZ
2UgUAYaIRJ++ac7uFWGVs9o8+lI9sPmU0eL5q35ubx/5lTYuK2xWe+DHxHs1DBv6
ybp60ijcRj4JLNc7kfkmBJZRB2m58I/yO+DrYB7LzDvyFoPzc65mIOgrUO3yenYf
Weho/dE09zsuz5vUljS2pYE60Sv+2o+S/lQHy7WJ3KeSQEgiSmtYBLfy8rt88fu/
N2OU2vJy0FXMwMglY223zNgoZdzw6+Mzcln1jgayGCSDyrpl1KOCrPrm8WWqwcOt
+UltYCDFQiou6TeknkIW0eeSmQxPCmxAdUhytGHjcvFECCYhSgAVXVvy3l7SMUSG
SpSkzaipJqTa5jNtNmcaRK6omVVf5Hf0F/kkKVQJaTtIa9MwIpEC7vngJHXEtCQy
M+aDyo5b11n9olGLYzuMN/X/rw63FDgvfuZwYyoHWJjIsrHKvbCM0SLoIJKtXVVx
9ML9wlYANZhpwswSKfw6aJ206qHorxS7T3jAMHZei83KtKSujndFrTCAZos9RMU5
m1Xf2ASiscpqDFg7yuPfjMGQo3lHhDATFeIUr/RoBwu+DwajOeVMt2kN8mIDeyBo
1nlZZVPdCdd7swckeQUdHYWDi8jRvkx7OO/XqChchyxbaNnQ2DczSKF5CjoW6hfP
YRnxLVbFRDkWdBJ6c81c7VebziHz5Z4iee/6TLZnzsTtEK0kluDkkeXkU9d3n3Tk
9EGHlGi4YrnK1RE6G810b8abacIdmVwktyov93djWuyCGPee+JPwMuLn5/BjbJfe
/RmMx7A+PiKeH9znwyFdhYDHdlThWuavrVXYAEuenaA0eBN/GcWPovUdXZVYIxvx
VXjgnN1LBw2MZUFATn+B8mkxkWGvWocIyjyPLDDj7mj9YZLJu7Hmmvmxxn3Gj2N4
oe+ZQofnhSDctS8pW7EW3lOGUEHqVaO2LRc6rJb4ExJOk0tAzyGsjnvdZj3Tf4jC
gpb4vnqIGw3ItQe24DbhNr28zpaTBSVx8uBDOt0jj7mKUEJTk2gTqwRm/wa0wlqZ
ba4u2yDdzY4RCHFBbvnPFAMFbDrgN5T6cSygB/S3ifD6dMuK+aQ3QaIeAtjqahq1
ArSlRwO4C4AE4SWzmkMyH5HeEZGeJpX8HZBOztVTRCJUSrxSKyJXwJF36tqvTpyn
AnHXGL9EjResc/SLJAVeFBQQZMnC3LLEm2gRXa7sAN9c0cVl4WX7S2OjJeLFrf3d
mMgW46XDTNAhTYxl1qERox7At+woDS6E3cBPigI7Ivt3cvKEqS/BUP11IunOBhxD
m22pqgHgh621E+a0Yd1kfiurKp2MRIMRYnpVTEApRZgLvuiF28Y4/v1wsfJ3ucDm
ckw7iJ+b5YZlRcbd5OP7O6ILIsN55mVnuEtmLB/4R63VryyYuYTBfq8ZngTUn8Zr
WPuBdtsy7qraQ3HdJ7evpTFTnZdyiegCU++NuRFHDFNGlTd3wBoqKJHFsv3Pscxo
PnvA74UejWOgrdp9HL9Rd525yYsYung1AE0jAjB0BRlq+UjJIIyDHx6X7lHguUab
mBntFYhVgI8flYo7YfyCEQr+DxGvbYT7kSc62ZiD9F+nePjD55CIoWa+E89ejfWq
7ZeJcYhj0JdmBSqPm3QWYD1g61ZXarT73iA+HybCzfjIk40focnVzmXIaPB2FcYB
lBU9ApvXwaWPdymICWf6TXdyxNBFP/UrLl2XPItCiBcRVpNJVNRxyDV3VUjy79ha
aaOPcWoX1vgjF+w69IE3TLUISyKlpVXI0OmmzVuRHCzq7DBFE7ZvIdga+/ko5nRE
SyHJPDVK7YqBPu7rlRoNy1uQZiqdURazkJWj8GlU97/15YQ4simuweEtziiOxvVL
jSRaj9Km0V5sifi0NbDgzoq9cBOkmR/adFST2+RTIm8Rbigz/y8cNlhssvZYbnrt
gvQMIMyqPz8Syb+cwIZYElLYAo/cU++inEjUTSeLDXaGoR4KPxj+fh828pKDFahb
07WKnOAybBRkdev8/zdkZesbSDl9vIP2t00XhKW0d98tNZfaScJz+se80YpH6Eov
FUl9gygIFva3FtvK6lTCwE3V6bjfOiHkNZ45+drOFC/juFDYqu3ZN/0E/9tajmd6
xMD/vpwHj+M/JpUFgWHTGQ==
`protect END_PROTECTED
