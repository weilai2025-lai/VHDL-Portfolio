`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOrkR5G5z7eiHOvSTZv1BB7mIS4C/zIKHSVQeIGmdC6NX085ti4a41fZ92GMEkqT
N1LY9v3dxmMAfwY9uQEEuwWUZopdbAc5Qz80SYYFYMrgi3wF6SbzTH2/9pvuI2NG
xrTB+c/7XKxx54EYbpoUSrXTjFrUyk+aNapAABtcKxXi8tor3lNvWgA4y0dKeebf
RclfjUzqmXho1s6tGdE4f60rg5oiRk7W7KYc/kvfUlFT742PXcij3ZY9OxRYfHP+
PXysIKitXCy+M377ZBDfKJ0jP/YP71lphUajDKfpp+ilFUZg8ur8+MaNhIXq6kpG
tFNw68fdK8NBKu6oJSLKsfd1v8BLbC5nPE0YSLarc8g6AuTLDPR7hH7dDYAw8aLc
7HQ/5gNyswA1FVHXYow1U3RBGn+O9dk6M0Bl7wZw8bf3WkpscLswH3Mpt8kK8sSk
5osIPQVB0LyqDavuhQVRfs5LLXZF9TBuvWLNaR0QPBQ5S3kkxNfFLbFmub1Y5J3Z
y7kPXFFXftK5XOyUJBkQiyFHhAzJ/SuSu40cD85QkAKPWn5hhVGifaCric4vUOEe
9vPqKp94ftbhGR0pf54WBUnVCYPQqSjMXCRUF2XN4s4Sqq0nzaPS8HC9kB044IGc
UAnWAtfuoYgprTFgZH+Fzua2ATgb44wqIMnBd/rq7fK1dgIEFybr2cc/YY7aXzKd
MOMpW7IA8SDK3YB+1luDmVg9ZjQIkcdO47V4kkV+RaRboU8lMztbDPF8/U9RtnvN
E1Y9AGtGzD8uVh3FM+PKWdUQmPdfb03/mqkKkcCIOfN31UYPf9+P/Jc6CA3O60Ur
5Dqub2DjwdAzVYB0uD/fMfvuglvbdCBCXZsyRrUIoSWk+aBLyw5As5l8I4mnjfJO
0oAqEqF7tTjM3CXlwqO6FwxmudMvE4JoddpFYF+ddh3tpYgeIiQmxmaC6P7AYowi
8EovKdPx0aHzTNFyeeyY4GHa45cO3ohaE0fGsbo6R3X5ZgZZRnHBMffJs2l+8k36
AIIdYTq0wRRp8+8SaLh29nE/ZMMdkvET1R3mK6LOycmi8Rc+TtD+SRfBf4tA24kN
7ftwqb2JHJHRVVo5C5nFlRcqspPKIUktLiY7MNCRf2kpXBNQmi1i1lJnG1XsgjU4
6/QVR2IwLHfZzKO0illJHATpWGPgwjwFdqOZJLZnlK8vaGAvy0swOZ4BWCzXPMQ3
sha8L1ZebxGwWXnyRMytP3qPoJ2TFO2aRGQGvD/Z4MMfDwqADP4Pq6lgtCiBk+qC
yG//LS85Z+20Z6Tl1dX5KBDu5eNG8H4NnBHh30PQLzHqGK1UJeQTwxCyjAmcObK6
sJSgjmSXFEh4NdtvuppG4T5wcK4H09Ogkn3iiNgBHMaDvfTrfhuBEd6d9tNvskTa
XEB7kodeUxcou8HAF0eva0GV1u+s31ERLTBQofOavWFgxfUSHzrp2BGSAhxWqdvT
JCfXewTbU2FTwgmU+rb5FpMSzefcYiQ1fJzcG6tv0Kt3YNYHieT5yWmfJT7W+pJP
b4izKZatHYaNsXwCCXf5HqC+diOtKV/lZzxluyt4dBfkN6boxUpbYsaHFp/hXAQR
68OQETJmMXNUr9QTdlpVwA==
`protect END_PROTECTED
