`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O3fD3AYABytQS6u3WsEoy2CBk0Rxx7hIkJ/dAeMoBCQJcKMMPgqdkZnjMRRAxHBe
GZKy7H5FaODkZdAEHbyO61vnSj0O4B8gXjJA3UeZ+rdDCMd0Mke8VlUo0OwizYG6
ECbKGks5BrCAoCx7mQ8LR8jC4hqojq7aXGHhoZiXz8pZ32/9BcdaT9S/WhIiN2p4
3fAcu66epg0maz5rSgmAvml9yU2hWN+JiF5a20v8JUVBItaXTdxvculpfEjB7Gsf
TnPlLbdUpKpNdsme4y3JiTruXtlWwNrOuT11LXafXmmL84/rtrMnYmnPegbXj+lt
KKFT/DXcsiiISW3oosrFcbvXGrROcjNd5IeRl23l9I1L1Kp/ew0FeydRlIoxL+x/
bYZ3/txJD3RruJH53AvRBBuEyhDb32IKUzs69CFRbE+uSiSMYOpEEKxKBE0b7BPA
`protect END_PROTECTED
