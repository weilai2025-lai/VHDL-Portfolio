`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgfaBMwunxt1DBbX1MLcJvIUmChmzu9CPKpBeVY6giXuKy+g2a2za+g1XbGbh8Eu
u/8LFV9+yNlMIF1v2VhRphpSa1AZWplqx8S2YcRC7hMjDiKjEcj9yvXwhLpTwvPf
e3C3Je9odRoIR1qID5BuhD6Bhp3PbTSw03XbBgIiZQ2RGEPM0rY726YO9qQ6kRtJ
5MwkIu2fw5suZhBm2spBzvoTRAkh4aHLhEpCiZmBIg21yXFvIW76Jvt3CiaZoHQ9
teWYwqHkdYH3DbU/dRFyCw2//sF/irlh5NAgzvGSUO+20+rIuIog29Gy5We95v2M
xppLRY9t0wJb4s/D9GFVUfcsb2et7/9MylNCIjyQz4S4ZQXzldhBgY1wjItCq3OA
RSqH9gQ2re6MwybnrAAwRUOPK6NaqXLVWafYukZ6+vM9zJ1pkkogjmTJjooglTCJ
O0vxuYkUCZAQJ++hoko3kRKpg0OGjGmKkcm2tMai+1H9iqb+gygsGtqqLGDqczsw
8KSeC1B1mJpkJMkhzn5mDVFBtx2GYEX/OeC2i91d9bmTroNz4gs8WPZDPcaWKYP6
M+Y1zKdCOPuMdActSPx+gPyGemoS8xBCvCBmKA9+SU9bPf1HSUL4Rd/2z2mmJPwo
xct2NagCEDrK6VybOQLvfZybAzzBbmN3/jjRLd4vG7EyqKC5vx0baVRcmXnXrVKA
Lel3iQu6poDI6ESnXo3X86LYpRSj+7PC3Ja8pKaKQ5x/6CkOJtWHPVWtYvEw1wj2
ix5cjbRWGqcTsiPS7qgh/K5KpIrmLLKogRRx/zWFwkw=
`protect END_PROTECTED
