`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZEbnkz0CA7QyEASD0I33SzuD4IwPg6lQJeafOG+YIid3PfQmBMsTx21cZeMPB9M
k7AeFz03VqH86ECPZKjniKARcWIrEwifnSpqnBDXAxjjGppEyCSkL0yjk1xR0Knb
ovlSl2LSLgtORFMGJL4MOvLKSTmTTzh8P+TDFtIQvMdHh0WXB5dWXEaMNqlA50QH
N8lQdzw+NovIuFed24Do+J15MD64GBp0ShYpKdeRE7THIovKsFg2cGW3PmGcQEks
Q2r0Y6TbXRdJoYXOBBF9tPDcmOrB/9MSHKMSxi3vLq8MhUZVoBhcSIixnOcAREb7
EG6lbdNlnNkZL2yMiI7PgtVeyld60GYevuelqjqJUdK87KZVGNM/0hGUuWArWh4k
i1vel3q9S5eAUODMnpjyHZG3GlG7CtEysyVse+XqbKAMoqVHnDdv0vbJVW92zfAP
EUcj8HRKutLIEi89Fs5D/BNHIP9/CE+wyxVjMTmgT5ouo1te1qGN0ACKRdOl7p/A
LCy+O+bejmAB58mS4kvNsCzs1xJxN37cH7cgeHaIJnkf7vLdLho5Xgov/Uq107IQ
AIFRTKwlCcFxzeJZH7tm2DnFhqxqFRLDxsyu6DmCTgZTXjmMBcpnhSO7oimwuSta
7PX8QhrXvZ9ymyCNwnWHnfeqpsRD5b37gUXE4LIu//CpNcpUphk4G5knHkHxysiQ
r5ZhHV6k2axB3bygpwAvggF98sxM0WCOFvvSN+3t0pwhLbM71sFYUuhBX3CupB7J
wTxhvaLfPXF2ecrVPqW+uc8AdUrAhFc0eCT6ea2VFgBCyo8Bd7f2tkJblRbRE0Xu
qFGm3pPIQRrqyH56vI2jixbLrjQdtge+IoOYlFcOlvVCHrOM8+yFSGslTCKBjcTT
EVNjXzxEAlEYeWQunQxWyz+Q8LNsXh9BD8C42HRAaoESBnhQhEHIFkJS5ktqEO9d
TWigmJXC1sHbSRNO4esOtC790sY9DNkNMubj3ojHRQWMHsBFNOPJNfoAxrYQf22y
/Lwn0VQnua/pAW5jYbP0ICrbD592HLSI+qTKn25SzX2e/Q6sGbWqTjlQZhl64RM8
3t5SAMjHhSP//FArpQYYrc7Ve+TzrKp198fOpKNOEuvqV6Q2DrRrfFe+/pC9mQ5r
rqfGqreOzZiH8iI0TPg7FBGoYyO70KrIOysSf9v+6KISuX1JA3sLcDxigiOYigAo
FTjk+epYpyF4BltLSiBFDCFSbkrykmhCabw0YH54q7DPFunqCWwSIvhvNFNiMOjO
8Pmza2sST2AaQPeWz1NbhcBLiOjiUwVsUSxmoYc/3twMe5n3eqx2xwum2DSb54KM
r1fzajFn+mDjE+nM7CGt8CVME1wflYXdCeUFYCGWD7bNwZdvivNLPgLoag1wiqOO
AvkpnmwrCnlSzrUThwLZA5S9OJz4ZcARIouGxO7swIjjLyHkNUOJVPImpX+Gwytj
I8pGFcCeQq3A4rEQUlPDirnbf5G+a3SXxbUX6GEENo9Vptgf3ufXjcFcdWPAkA3I
9l2AL4xl7K2R37LACHYmK+g9zIHpwO76AtTkuAeNhgQHnOTfDAH+f/YNZ2bdWvFh
4PQOXYwX+BQiRQFC8x3FBVA87hTBJNl6W0gjlyoz7UAZ0qp2Xu/jwv9Nzsm8F4C7
2WKsanXHwqzXeoEs6jI//34iGACiuJQNjgnA1mp16eYfgGawpD14FCu2CeLt1AiB
YrlXy5hM3I60OolEbfpgIxv1/JJgE6Ur4hT/WPMBJVahlVqZpCWNVz9xDTfX1XIu
t54+AkDPjkDIEdPH4EbJpf6U0lZnUy6mKKPkq7vDsx/37qJkYizsE2ETOODMrG4Q
nmQte/+80qpFKFhm8pYYhrvWphlxt+tMzjK++iCowO2WE8FWYzCAsqFHaSTHs65d
IjX4cLQ6Qs5oojYzBF6SkUWcAA1coTnw9JmvNis4riCc8vRC6KNP8CHjhLi1lm/4
W438+qo2t9ETc/lWnM1jJcLB6uZc1WLq1dNElmsAF4eAQtrSK2tDcBt/eOJ5sOdF
deuFDWbi1eZFOKG0+ZWO3WtUzuiq/JN5anWV/Y6qfezHwBu2k7Ld3CULhl+w/Uzf
DpV1azdC4gZtlemQiJIYW/upoNxazBfAeM3TzZ2iB0UpF7R46uvuQXInMrIoiYsS
r+0Nc6EBFjQck4iLPlVeKhqkP8s9rKCiF7Q6JA/Kan36knMKYGzrgDvA2KD19D/E
XMRZ4Odb2sVdC9SZtKzPMkMQlWES25WvamzyGdJAn525pNE9IkFNt4A9GWovm+5T
uwR0ad/S2PjrfU7RJMm/4vng2yr9vGb5Fj2xPKZf2KjSnDfUY0MK1qzlEzg0AhRP
rxgYxiijRKkUThzD/M9z4fyfi0uWrTPasKv219/lhTA29YJUVozGQNzE951O4JKp
BdNa8ECSBGbdIXlfowBXxfkVYi3eGtLnGdwRcuY+kELE/6nmHWvnKzFdV7I/SwBz
OiRfCzdQ4cbiIFvnkzfxnWjBenM8T+lOQ48Pl2CoJnkU7HpmZ//O0q4qF4wL91Pk
VevPEY7k4rDuIL3bJbvyPeSHu5wEqTzbvy+0+CL803mkBIZ2s0HhOHBpJNv3Fat8
cQ9LTfczRr1T4OUpVUD1TM6ezpblqQ1KBf6879KL9s9573do5EJMJjU2iccFBzEn
LqxbXX1T6XUqRSVq7vsTNSRDUubH/VmkoZ26KikNiuHcKiGZuiKDFHHBNiNFXB18
Po2LfHhGAeqvxQNP5uwd5rF+yHqmDJ7mF81OepBTfIqP9SArmJwY7HcPL5U6v9Hf
W1TLWoF3E0Km/FY+uaVHoj0NXdFveB77MpcohGW+/RalHkR9POHvokkE5IHbCcM8
a3VZlEixh9+zZVMiwTqPkjmTc8GnQWwtdnhwcf0PTkT1ljkCB9wGvfx9gDQbPRrf
HZofk8YWToodueLUw6jytausTtebWey6WupBXK2ub81yxvqK8+MRIcv06AOJY19B
wTVGKcRJ59nASacoYAhThHaVS33O2Oa8enUokqrTbEr3PUsSAH+RW3tC8O6Veb7t
OBjyJgdkkPCOKDFiZVbTQ+o6VKi8vzuxaSFmp/USOylKL5Kx69sl7UO0Eem/a3hE
xgb7DFUEgY8s2vnHaxRQQrT5VpflQ2k688+lYi/oz5anfzb65TMu6vSM/Mh6MSM2
IQIKSo04rf5OLNks5WAx3HFiLJSOgKrdHYd7o9csjtn3D0CuNI9+lYTGMjFdtUOt
xTYDU2a6BP9/0MbfRFveERmWcav92KIZBUTXq/89o/dvaIz9k7hS8CZxwqFR2oMI
o1WzIIUibV/P91AVIxOH2v0HGstp2FYbTj/EXd6hblicceO81ChuSIvKziQnEnn6
1ftup2sG/o7Dnt0tsEFqPy6gCXlN3hHFn2KZbSVvSevHoJs43BY7PPPEn5wAHlWW
VsvsyG0d9rBv4cRP8hxxct/NfK35egiNzVBzkeanhv7WUNtlspoGBgXgVmtxQH17
guQ8Syw7jhklE9/1zBXDmXm40cNFGJ5xyPzXB6/FhDPDIbXRyt6qek7f5NY4x3Lw
uS7wZS324hL6Feuhu5lERqs/i0jTzhHK2OHsC4GLEZPCWSeDYQgB1IlE8gcMhHbB
toenwLliRSC3n4gPmo72iYN8YPTlPXMVTdYCxpwWVghR/S/dT5lqJWSMSBLT+hzE
mHZ6bh54OhzXnm59n8cxTzNR7s5jsIgGCGioBSLQEaJsodyM7RVqY7loQsNwu8b2
EURwVsR5B8WqPd46hDHR4Vrcyl/D9mrWVL1MCWxc6V38x74AHqN8mQeuaTXZ6Q6S
SE71+Ljsg1FASNPhOV2seLBY+0D3nXfq45cev72mHzncOQzcM/w+FtJ47o/kXF6P
ZGobdiU0Ccayz9+LdDRbh5+pGwMye05+lG9dBZDSz58KqQtNzAe0ndCVq/JcFSwr
x0puFHpn6r4RsQj6hJOS/VxEsL2Fqrs51C6oJPb9P++/J9/jyRFZPRVA+9P/EBc+
BjihfKuKnGJDwxAM3U8l9A==
`protect END_PROTECTED
