`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3QBrixJkzgWTWSurNPVY3eSDU/fV2xfHw+D0IFo1cGWRkcpzUVwOvyapXIblTn2b
nDPKRGgAihpPZuFR3XLiDQq+ZXeWeT4pW1panNis8iA0pyVgCKGD1Bgdvs4UsmII
w3m7WA7EMLOSF2sSTbu8UWe94B5DzqzrhK6UfEaZ4KIMr75AqwDQ2/7r2/madxaV
S+NEa07GuFquVZ8ojDL5jmxsrGklkkYEb4WZ1ecaHW7Gl7yBp3Epm58NDr3Igg6Q
wyJ1W//ca59DObKhHb7llw+LhI0RWFAnDpVr+yXqtR/OYrV349g4rdKnDJ2CCHvd
04UATO5SIgSHLEWcwfMl6pZXZxLkQm+Q9VwYnbf4GD2gbmwAmVV3kz6dsm/I+IGq
hhqG726Wzu3u4HHzHy3Uf2ULhInuTjCyNA0h2RWFIES23kbAD5HorMGBycPfYqSb
bpBiFBlczjV5bHZPybTanTijVMf54fGQk0LaDIBQJUfBhkiVbs76mhvRuNBZ5uoh
xxt+BU7d7GwYxjCR5nEUuj51VmLzu+hFDR8ZKSNLF2VSRLl/0CR+OL0EwhJt/v3+
5qmUbFl56sqGHndCVEqifG/CZqamojU2L3qnqxj9Obv+MDaXMoA7V2l+S8Muk8VK
7ur2YYenOkTKgZaFbvstnSqp7gLHdpustcbcNH/rAEOeWifu2mA4XQYQWorFrJaW
77YmKYmX8bTtL/j6SV8gaceyRUEGY78UtOVFCfmtC4fGVM/7Z+b3iyO8WYdZlgb0
YPFnmHHwUO1J7wWnn/AiWf184WqZxfh/2rINUZ2iUV6YBsdfZlWqyJoQdDt414J1
sNwUTW8JRIHRZxwzY96VibZCQkD/fnPDIApb+4vY3M1HnTUIBGuJXs5oNheFYBiK
NqeHYbMctcZbX/2Dnq/L42ZcGPuJV7KVkxrMWSLGx3xw3LRfpGyXKWE2x8o4y8SI
VTebcwQr79Q4FR2T7kjiVjbbPB8ZCTBnOXhCCLxPD09e328uMmglm/5RzV2OQptg
EQCrBpGCBuW1RAHmJUycUt4zO1BNKGC8zeKbfwyK1HngRdxYniDQJiZv+wV6Ih1B
aqDQxwzyvTei2L2FebK7tfe88BVj27dXz/uBdu7S0FP602z9I+oH2NeovOWskmKK
JB0oKGRyY62FuVINWNrlatgyY+QL2h3rer9gySp4Nwru7GXSAoWIJ6cPP9u9mlRa
QCzFE6JRtG5dS1JeMwY3Y+sQln7Z2Bf4of6kL/G2wuDgHU/NDxqrmmTZFPimje7v
I8a0ujLoZYOECGI/EAsRWY8/wP8o0cpVBqBZmtGKnXcpgkFuNbBiNjay/tVlAkPQ
H/57Die6QIQGgprgot0DOgetNLJhNaJk5zG+OMs1FHwHPdiNeOUPOS4P5f+hOl3b
LdS/8J9u9RZhafBy/IM7+ExYZfKFlEgHZ4ALiOehY7IOT8yWhmEv97gqI9tMn+Jj
YAbEaAEVTmK8H3D3jmRPpRE/MfjIzxBVMXyAlm+fbeQw+ND4SUvg39DLS4qsERUC
EilQ2HLp5Uv+mC1sy4UsS76AKves3QVtyt9c69J1HGmqJmciVmzgI7Sfm+0x19Dl
`protect END_PROTECTED
