`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsIA6Clx0/+BNpuTXautylRygVsqL+Wy9QLug3vzOKCTqbpEtPe9kcQ0VqYYN1W1
QXX4r/6T2clJp90cP/ktiC9LiutHskqKYvTqFgUg1UHOc+CxWceKTGkzIgniO942
vN6TIPcjyjzwjOPlh7tZY0se294ib4MsgrikvlivdIcOtbFnVGozAJYueyZxkJnu
lAmHtVgeBWbxEDO9CzxplyWu57OOM5bXX+TMdJhSoc3Z+V75feSMnRz8R7+zvZWt
sgr0U4Qalmac/ZDXMMSxNGlrcgdVzn2Q0+BCKs+SRAkwtHsvTT25hAoYziIgc1it
qPF5NBkOg5EeGCgh9GLlAGQ5Bn9Ti4Fi2VFw5UgHg+J+HxVBIOxPFv7J2ZPsDUap
n6e2OnjWMmGCQrhnLlwaKWKoabww+LrVNR5ajny2NvLbwlBjcI0q/840mbOJltny
ScxS7m+9bwtQeGHdWaFPwqD95YFVelmqvPBb9pPaxKkkKO32N3OZIR+Cb3GNyQz+
vZba6t4YvH0UrFw3MZZW+HOu24XeKrdZmjDST4O1j/mmL2hORHM95jCAs2wceizK
/lgZqTI/jLgEbDBYCJVJJ46KNisvgKeH6iDKzBcxal2uHKvGoWHYodmZduJF1f+b
hyZeC/FO1p8jYt9/rV9QBQ/LYKiV1qSRjtV8emkjShsUFCP+6RjYID19SdtQzysf
f7ddxNHQuPgCSXBp+Dn8rdLlkhxcNU5AjO5ZKqJE5sqRyjP2aPaFldc+qV0quu8V
7Q09Zi2SayRuKQ+GupfH6jiBdmWRUV1txiM0+1HbhCWvcxQsCmIcEDqtaEC8hgib
6RNqUubBjHvhCyLfz7UncBeQVmze+WilJ/PwhjTGYtkgPvFL/gScNREVnvamNaMp
JdpRztrnReRMuHDnD7+lOrgPG5lgZChSYhQ/B+isgJzuS59YYWLJwJIaK3/uUxcu
1rNk41IrLbPa/FXTHXGwGfgwvnIZ32N8JJUHWp558sysY/hNc3eIkJy43Sf/Aaki
BpFuEyJEZLTVEfxtdXjp3Mr/QIIiEyEah2kYwX4mC3wpSczb0+Id6IbvcybTbvyV
Bk30hJ1+hnHdD9vkC4w38wNXTgpTXEKCqCLG6+GZ7CrjlwqhJOzkfQvw0kapIDEg
tNEpGEVOmbEzF33QOq0XWEA9a9aSKJwLJD1CoyZIINuq84DUaEx6fEwjMJYsCXm2
7TrLUUBFj1MuxgNM8XH2gIXzG98l15GSopn9QllmWLYswTubIocZPZE0AkuJzpLT
Y7ssTfVPqatRfquupCtFtKspcdNOE8bHqA+Xm/drOo8gkVizThnLI6itvq1kdUQn
Q1lTb3NZb1LtJNixyMS8yWRehomf/zShyZskz8GToaNYePy5jHFwOhm163GzJ6xI
tocO0UJpFLVze1VkvIwiwei2fvYZgG7WeTZLi2AG5UFV3zrkHMN9OSqnaYwrpwLH
gvUFmOhOTPlxqzRCK4BSt3JCZUwxAJZqlVI6Rnnz7w84OhWThidXIi2iXpixtWfz
6OpIxxd5fYR/EbvjwLW03UWkSzAvLkYugqGyL4sEZkPF0S+arfRVCgqCnX7qF0uS
rzq5ISioxrVbsvbI13U1mf40uWUCrKROcN8BLqBPF9+n402SDJZls/w6oVyefhyx
HWpjNJCRnGplNxCxcsLztVZKumQDLGAmfW8WLMnz4moesAaQ3HkXcKyBTS6OhTdr
Hp65VEaSyIWtTZoI3N9OP9bPLTMZ70H/dwA5KNLs7y0C5X/+Gxd7tgTj1CUPr5hB
qBf1869Ggf1u39Ei/ngpD+tnYg5qHESS/jnU10lyg3sFe5RK7IQ5RNRpaL5ARhhg
lHIE44cFOtI/1H/z0jEH0UttyVSEJx80DN52aFaT8Wit6axJJJRnwzHTRmlaY87/
aLu3SwUHobAFbhUdUYn9FH2NX4FulsZnSNobo8b8UVGxrbnr7JxAxKWZmSAniN2E
CLPvTMLhu1wVZ1tT2AezOa5Pxjj/QhXDqGBZC49o9wwsyBNdKZXkpiJSU42kUntR
o50RqKfOq2gUPcFsR9KVExHVC+Fo1CdHgIEMEnHYAB2UnbIVC6ZlyFaHzE16pWO2
okwr2OZq6d0Bg5FA27NLZqmgQHeRdWhgXTsBF1T0sQcEAKNJZIFC5o283jqLpuow
4LRZzcBwd30HfuSpTJXAzo9ddIHNPSDIMuC5O7JH++S5UdM907yB4Nxf8psbFHsG
hnIkyBh9ZNmmajssII2XuIaHswTMNEK4r6UU0ZNo1lEzLQ8qb0cYjSINVJSblbLW
FA92hwsztj4O3+oZgbYLNUajFCU3yj5Vf69rMO685SdiD2lfUhUNmnwVzO/hSQI+
/3/skxeraFn2WIGhvqj/IapO+oDIf/+JOaYwJau88f24hbSPmg7HyEK93YlWEL2k
y3ytI8ztMpAMayk+sUNmd57FrVaHDULuN6oc/XgJ56SF49SGP6abL0iMSoIuNRXg
aN7Td9vLqzEkRshXxR0FU2KlWA6u050Bn1tBRAoDvBWUwbocJlnE2llB30Pzpajj
gGaO7mU9bjFMfK/NY7nmzHX1O4sfZVbaixQ8hrisAbV5a4HM3yJklmzAntTfH4Vx
mJrkTIawQzS3tFbclj1IgQ==
`protect END_PROTECTED
