`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tiV5VM1D/3aZu/rgKDM8BbgYcWdX1R24QNL2Uyh24AwXsyDbgTNPYxKO3m+HpwL
gyrB1ASn7+erp56ntvwDSfmdOGDjOrKFq91IVi9Zj9wjYlVqtp3QTycDSEF/5OoY
Tw0C5ipuMd3kWKbg3vVPNzTT1LDawhtTymtwWykaKTYdh87+Viuu4tt//H//WU/T
DdrIXMmvQEoKmhikxq1DqFuzNhVmvoAuU3teQ/g5Z/hUkFuln4CxQ91kA753M/nO
yJZyujQ/Uvj9Sd7Jovp3n3nv00kJkBa6NzxcdiboQwtJ/geSCDS92+o7pXs5DvYL
5GAqKE2odU4rxMolylyEPErS2xbxyknY96Tq3AnpkpQ1TaX4H/9wtN4X5jckZa0V
R6+H0ROBX80u3UTzpBvZ3MZFINgcdzHQWIXXbpBHjSoBXfjZ1achmNA3i0JOEKeU
PlPesKWZu8MbxUXPBmRvJ7Bqbd3XhwtWp0kRmonIujp16BEie7CJs8PJzqIa5PZH
EjGD3R1UrXm7VuLPIrGsZsYeD0NH3Zxh9RMlabwzivEy2HVhNmRnFyxBtf+JRzm7
uCcTXrfUVeJKTjk0yJikFXQW8MGCN62eWlGZJuZ2BGgMUhUjLRGy09/sgf/Y5lO4
/Wc5WjcRJaHPDlG9GihtwkRg+QqHrRn80cbp7MwaNXqIXEsWO/VHYaDNrm9u0CdA
57WWe+VTOYdsSYbx8CAltKlUoEgz92Al8I+Vs0u3cXZ/6p0BoLfEct+Mt5dZYFY7
xd6Ts7a/SAiLat0L++pULqZUKeCzMDrkL/vPy7GylmQKqHWkW7vzFZDsHUwUBSQI
Iq243x+8AH5vQAmgRjQJJLw+BIBC90uQGogGTa1g8gd7yJj2OoFwfvK0cLs0yyhZ
itBSufuWCu/PgLk1t16d6vU5gyYaJzt9qucLpA4LSigL/hLocA2jmvz9FgoJO13C
XhKeFXzcrTEgm9OTlidGTBKYl4j8W5wbbMoVZlzjB6pXImjo04/4oPA1gX/t95ly
c8XHwPtX2p4X1z220CqrZmCJJUvBa2mUhNvH4FpKg4QTZz7rYSLl1oP0V/HTL45+
OSkDDxTt9TkEpWMWRSMlqkJwsGP4iGgCQQjWvDTZX2+feBym4EeBMLQqZKMebZsC
jlntPgRYbkf9zZapPDETgzocdnJjaoI6nAKFz60Xtg8Bubc+6Kt3GaisVRlugeEv
TPWx3magTo7azh9Hfn0RwHNtRGdk/Dj/jo0xkYb2O8NPj9sA+RoxR6hcoVufsLSE
OdR1Di0k+p5CiqoK/A4itvo3B8DOcpf19QQzW7iPgz3Y6D+EMk7oMQ2WcfozSMeq
kyCVwgEXjkc2NGbH0bSyusErjBVWdpZJjItL8kE8wllWbFZnmOJzOC+aMVA4DMps
dCXVYtFG1RNfDwLASDiWd6NpJ0ezZK1BiFrLT6tyu40g3Hozol5mXdmHcCSWAge8
pIKlu569n6VMpyqwk8vUzHLrsMQdqQ/rjBUbPF6J9k9dnWqaCacrnL+I7ZNwTZPx
I9DOMt9t6Ht4wk8H8FCIHNHqQLMFOoe4h4SSuunuEFIIHgXvkigpNHEA054AEm89
uY5SlVu8+enccGDJROjGq/BHSdjQSnfiuandaerCW5z/4NtlmMNeNKr/ZmySAuNj
RecTRorclOOdLD35A/Mut5Re34JWxP3itcoLSWd9pQQ7HkXCXnloHZ5XLDkaHAdI
+kccXGN/kZ+FCRd+fcYtBytcEJMdIU43sKiCerV1BsG+g4NV33fzSWg8ekdcfAO8
TccuWmsO9QYzPz4l7W3WEmgoYYwYWLgttYopN6QF1z3RPtEMnud/ncLPSczjQXbr
f7fwCICLmzrmbk1r6NnsNc9RG1eQVpdSen1f3hX+rg/33Qobe9wx/qsOmNM8eF5Y
zd5M6kEcxNAVpBxYi3PqKUGwLY5lZl1n8sVn6K0wi/tpuwZQDuQSFR9UjTcJwffB
7nbYFdUxLS9VC+0elO7bE9n3E1zXFf8gkt9AEzpbeIurqzNpa9QoVKApTZd7LJWD
I+yGa5up/kqauU3TFFkaX2H2PzBeVBSh71DEy/NMPJhq4pkNINnczaP1XdVgymeZ
Bn0KzF7t6whp/aDyw5W2AFVGG7otSuUFUMg5hhheVBlgLhZ1UI9MWU3HiN8rgBC6
YGmOCgEo4YTUqypiL9BC02RZ3x6E3irsLtvweg+xvhMgqTM2hxJoE+dSOuULw8Kj
1Kyor2PlU1FWGiho0g13eDi1V3iNSsqMG0VOB7kk4Sk99oF7yKdxEJsDtHG2hwMC
NXJ9mqnT3/Ce/IvzGUIdiPhaa5CKOMJYaHiUitwD9UiY7LlgJqXyBoqKcFkPmJ9d
Ukbqxlku1Uh8dFzH7xadEZCGi6s25GVXhkqTKuugcrCOdJPBSAaEKam374g3g2f/
kZX4kqmV4r1XN3WZ21DJbz3PwkyOev5sQeQJOe/6saVy6JmGnifoKzm/ebGojRDG
QCZ3KhPRNOPK9Csa4JvFgI5zSLYv9UZh15oTK2JgdAUo2YsBSkHpcMGXOFIdM71N
8ZlpG5AiqmH8y3B+Rx3nU0JnFNnHcphnuYxf7OL6wCLpydDg63DhhgW3VdRhWI3W
U1WMnMunuDJWUYEs2craExbfwSlS3bBuSHong3euT4yF5RvC7DpRBET3aHKEaF5g
xlDd+u1Ovvi/FCAoOlVYAR5PCwEuBPRlgogWvei7hIFFQNeSwmFp6hztnVc3CTmv
x7+p23q+/BXKxF00U64kTFWdKoOFQaRFtfc/6EZCNUVNTGlo+5hcWbxOSqd/pPmV
5yKHWsGEnM7FqGcnyUaMRp0spWOxP3NdDO8shFTfMW5vlAl8Cc4EVHHzPJm7VSPv
PPd9yzFBDL/eHQxS5t2j1v9y6F/EsEAcYGa627snKHSjZ9Dt3pm3Jl4oFy3aYSyb
fNWPLy476jye4hGg2zmJR7htuwZcgVihgl54JVfH90orPXsfBP4yA+Ijihxyfeor
ifaxcXudDXffzO9J62mIhjpF6HI0TpHJmOXKJrH9KqnNnKvvf5TzanPzxz9tKmVF
u/jkMqLO5OaUQWeMt8S+TOREQY0zhETQsVHp39sl0Mk5EZ4MbJdUJlurATnwVXJD
9vYj/2bv/Q7RSOAUfMRjQ7lZIY48I6qTKQBHdktb5sbfNP0wXzEVfHsDBunyN7Ir
wgRmH0X+ScxOMxFHppNfrMfiSXLu1FvbkbqB3tLel7TF5KOpBjDlu3DQcPyKx/fF
O+0lPTJv5Im3MwgZH98r+xvPzcfGpVPPIAGQbcokfaAEau1FX5NzFHL/LD4ggqvb
/tIWsxS3mTbtD2ZNmDzSB/+zXwB8SPrpwPW9BvfzejmqjMa8p4irv+m8Ta2n4KW3
P5MbGES0YKXI8polRFNb9d9862LRbZXeF07xdK2epFN3vCBdh23WZ+EGoeR9yzBY
mvDA8lijYyCKM3qsqHyKHmodLn00x7iyy/5L2jElKDHkXVTC9m2N56MxMEOTUHi2
j0j/hFvZbiTwY2XVBvb5ol11IVKbPua3KNIEogp1di3dQKqu0BkVqLV+shAQYoAj
XhYM3Zj8taOp143lOjeAqHTz6MVjYAS9V9AvoI5Df6HpwYXVhVfYdwd9y/Cs5T2S
2j9ukhlPq96cN0ZUcWaY+ADQQb9f8FQFD1K+ApiFbkc7STd2GIFZFsQ7B6+7P4Bs
DwMQiqS3PJHG46VAOTMcIiv0ZK+LkyjgZfRHw5+3CPYjivQhyjUlWNohOsN74JMU
pylbatduvmum4AuBTD5FIzwKf6Xp8siDvVGjCIED5W36T5A4yEnNamKztU19iuDE
6JO3dYCy/jRP9m4F6b6wLyIHSG6c0kxTVCLYqexQOaFNrEZR6l1b6WJFbL5GsC3+
JK2ApqleBuYA2OtFUfFAmU2ILa5FCz8qa3gpNNw9spgl40SgVV3CBk2fw7+TNfQe
b3UKFGH3U5xQ/tUMa6zF0DxT7TH1Ry6x7rOmDbkC9RLnSFEaPyrPWvnLtYQeY9VX
aH0BQFNwL7Ra91yJ0jOrW6tf0yg8yg1IaXXwPGU3KFEMtwQjitvEkULYWOjXVEx8
ZOYL74GGF7X6ER1BclKoV6nAkZVVR2Vr/LokVKRY/zfVq6KOBQW/hzg8bprf8Z8g
iZEGFaOFVrUaRxgZWoPkcdrP5RIjPzkd6I8Tav3aab7IvdMg6mQ+FDPctsY9FnvT
MkkbaJKhiVbpK9zDB6ieMQMSFLWWHzXyOwU9a0hLuhS/qjYYRKJsfqchDlKRlewa
s+csY11FzU66NTIIIWnIKbLjVMjohvtGnWolt0cE9LId//c9tJt8xmkGx9fRxjpH
en8WqmIvLJkE/XfrC5OVtCA09SN4fGX5PqXsQu5rzUzFRVTcvXY/rp4k+L3iRPc8
xSKUXHG7SnBhSQOG5rM2eHG0OpzNhAf8GznlfcEjvtJ01vuUeoWtMxjA+5JuY2Je
2fYObex3VWbdRVCXNvAKghQwNamAzfcykJGHaDXWMlKHjLCM6p7QRvB25x4VUL1N
KtfgcHXPdJhEI58bX0AuHwZIFl1NBviGQhdg+OIHeaQz+8pqddB3Z0o2ATYFu7Z6
jd+rfjHjpqgQauxQhgSdR1zY6A5UCzSW9RROW5CBfeqKcz1turIJFvOIARPyK27V
k19y1xlC0a9T+XSs/V72jZr/YKFvKLyrDJG1EyOHIMNIoGXgy030FbjhVlUf/V9g
w/9S7Gxi1Be/UtcfodiEBiH59idzKZJuvll4u58k42GPDbUYA5F+E6onKrQrrY8/
LpnTN249Za16U/wVpEzPjWvYTx3Z+UYQqEoFjFz3MSoQBMNKbHJNDDg0UY4qBEps
wcX5Rx+TYnFGsA3ZZd7krTXn8PCHxSI7yWEigGV5HoIUy92iaPTpph3r7HJvI6yd
qhkBTQfJz0ohm60RFNYzO0tvVeOuExbWDclAk9BvCkQdcs2gyoxl/qAbKw61INgq
QABF5bltgfvXndKFEyZPMFWV2czMTVXGoVy7HCknrD2xjHVYH4QVrmq98YgjUHe+
GCQa8YPaQfJBfnQmAueM38PplAdKu4+Bzk8AkmkO0cbijX4Tq3RmKrcXsxkGhnxv
JLvtwiral9adehyMXCzP+FVvHOXgqP/3B1eOQkUzRMcpbYYtnoghyDwKumXJpyy2
LlQM6JMBEG6V5hG1BveCwoghC4kf9/2YrSjnlBT3NKyOGioWvOpEdctWqy15xjK2
EQ99kd5n8DL8Six7COLZwtw2fgd0XAwh4w+NNrol+g4bpDSePMWxHxYBx+Lw/0RU
dCGTjeleUI22fiv/9+c6RoPG3fmwPeFucp6CVHLIMVzMm9fLWdlFBOnkl9Odg302
CbQxscMwNNYwre9SXNNE03n+gWVGZ3frKLetZnBBKfAOpUgfkQnOtAm85kPghC5i
4OBk4Gr5lrkWnADkg7Dp9T0a5081o4TsdBzCOb/+TtadNLbqxU7LC+GOIhe5rqzA
TNShjukuR9QwZ0yefHcfCk6CWHrH/yw/55hDmB7hGm19r55/Xus/1B3aRqzFAj0i
MVvcVtbWP09ff4j+pFMbLXuMTP3YBJCDbgbhhowJ12nQqHdrwh2pnsEwV3ScDvw/
V2NOX52pRhvnh0i9bsKXU05imN8W+Z8Q4dFxGuMYI9lg5ZOy+fN0BbUwQCZLFj9R
qsu9iSFqVnPpdevmxvu1Wxh79yM80+g3IThw5n2G/F/Ue9CyV1uH2I9m4NOCTFl7
VhLXdFmVjl7C9TLEEfQYMnivItOEM0ZS3815ukUpQzuf1i/shAoY7byRq8abInXk
aMrwuTvIWEAWgeBC7ZFmNthyhy4BMKan7X+oUZ3l91Xwiko6zxU47CHHBgdcyCb1
CXlLiAF1s/vCkNHFcWwrSpEwAI0BHqB3CwHKBsmbG7lEW78nqY0LVrscuNHTXdlu
+LXeemmUw93O2jy8b7NhRJv4/6QKmnNgAwKr2w8+3UKRG2/35RPvicnJbec0YdPy
Pd2mXDqPMFwsmSese5t5Q9KEZPTinSUeB2b5iVl76yleZboqTiM5UghkAxW5INF0
h3FgBj4hJ5cOtcJAL0JnknCEpJT0QsSdJSWCB9PWoD9nY269vKlQK0gs6vskBsdf
S62gjF1FJLUL9qftbLqayWrDYE+aP+oW9uWX4P6SqMrpVx4vOjKOcINlS75k6Vk0
kcEJP4UM3BmdemNnZ/pRPU/uElUuaVqN++d2dcH+InG+HwGk8vWy9IH589rRd8N6
aar6++y7h0+FL/QTedFEFjPPyZ9gtVOaqgCu/vKAp+FX3GRVMpc7c8jT1ATNDA6W
8Sczr2C0vg443xEnWhgyOm7I45xrkoleJ5FMpVMbYvx2ZeqUgQa4fQYbIqh0aSzU
43rDTg32eS0ZxoV9TEyrKdgMNep6B6vOwhzUy6WyTGEM/mmgde25PfvWRwDNMiCv
e7oqiTfZB9+MvRGx9G5NyQHUNrFsEdpsNRvS2B3iHzZZwEU2uHEIz7FTgoWY7EdF
YocOTRFh5mE68VXIVOR40LUFKSCNEOjRx8PXTmUS1fX4msJ/47RnhloKnkiDKziW
hcch5mzaqBQ4BhtRTQGzdyAFe/ZM4C22rIrdREhP4fk6JN75pRNuM/tDdNghe1EL
mjtdnzmQuIpP0VLj0QIndTu8UcB8wK+8AUIAOi+aJR4iLW2wYRv8TpZRqUfBpd2A
yNS0ocBujVtQ2QmjBSZ0HsQfvL5tlPYL1XkHBAFn9sw8xoPDKAQMGOYsTqreiXqk
a9wgZdvfeHThhnfehEQf1regqBNtOyD3pSuwjqWr8pQ3tjVwOCahE5IfU8pIEL24
Pmpr9vG8+ycPcPKSDGbPtX8O2ux5SCTwlSUO1hp5I1ullVZ+egm1WOn/dHfgf8Oo
Z3z8WxSgOoICWNI1pTA7YCIgL38Mv0re0nCiTJBVGomtfHv2UD1OybIR2OwlKItH
3j0gxX7GnKSKUo4HL0mWXzireonmC3ssq6H8boB8Xtex+T7mBv2B0Y0jvJWo9JdM
mQGeBFXngUgEkcFrSElURcMul4UxdsmPPg+6nhi/vqliCeawImMGqI9KmW+nzCGn
jceHt/RAP+xZGYTq+9ssNFoNTgwcfrmeTT5dndAikhjkEYbAQ5JvbBLfisWbBije
kC6FONDwA4BiQyloKl4QecPEpQ97LmhwaH9e/sMie2tazhyQIn9rwdajt8AreTLp
ZRGwX292ZdN1PzrqpyN+nBj3LjiYBIRTY0y49mANQiAKJCu6sMPgwFW24Ha9Dc9L
Q/2H5i3hNpNEWCoLbgD5KA==
`protect END_PROTECTED
