`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyQ16zP/72U2YjH2twv/3mU/CKov752Ek9eXHbyHmLTYYHquCIlPmnV7rzgLIY4g
aVd0ntvRIdb3YsFecEchtRzqPtrIupkzSoWwPUaOBh8br0meAxID0aVqYMS4FPWJ
ndQXETLeCw+m8WS/FowbjigDqk/+AVdH6ORTi873H8SSysOmRinf8g7uCI2Ccvi4
YJB3ww4Of9qclXK03UuogqcWO49Qg2JpSm9G/eIvs+WKRYBFbA2Q3u16pu73E1gO
NZK84yu7DDFxGwWnPIKD8nq0ZCM7YHClD0P5pPv6p2XOct4WqSsznSPp/d1a6E/I
SXEC7mR5QbeF0+2SnxwjIgID/ed79z4V9XTupsdb5rd9M2942lWBygFyD1l5GFZD
WbDhITLsJxh8j5oauejFxoPs4F11t8VxXjmIWk4EeP6HwvrzXJJh3oehsmo8Klf5
jXk2AKmw5igwBCLLCCbb3lMzNC3lVczImI7rC7uYZcv9gXePKkp328WOlSlQ8RY3
3eXQ/yjcxqdQZLqlslvP8J//TYGxS56GaXzsPi98bgqtUIzldqA9lXf7xSp56lhl
MYKom/vD5eldsibla/uzY3Xy7T869UYdJxAsHzLctksBnljw1n+8sE/t0Ckb96xB
+PCIPa1oYv74/qyLoBUWfFq1XXiFHIbxbKlzOClmgVN3L7V8EqcUBjlBN+DyKzCc
xkuODsCD7Wx/2GlpKI22lGs+pPIH8l3JICtCBl7z155IRE8txybOql/wWNGrS5Sa
03v3tkTl8RiV0zbsTnvj1FEs+4lVFYa4LF3e4Qg81yko9sBxToBAmE+iJcMJA2IA
zv/XnsQ22zWgyWAnJFDNa9D5Vx6yUd6z++p1CM0facJy5sA0JLSUsd3LwNhb/W+2
1cOSvnW0RskZ35yxj/7zwEqQLeWArdr4VyNZQxwLI20=
`protect END_PROTECTED
