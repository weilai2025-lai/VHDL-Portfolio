`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2qgN94t8FMhpMxck1wzcFll1ZK1m+pIYmbmlEiN/yX9jnqOOjX+IB2WounqNmjqj
urRR87tFsoHgdDKnz6efLu3Dc4FbKp1Wf8UOPO/cBplp7sJy+W5dKwhSNP6uZZLf
jrPyxikGPHrsNWGCXgztSVG3ZpTlwSJBrSCZgn8I1DDvFD1yU/Ribo7fErTUbob7
vMPc0HRGabKpSRBiBmm6pGZbgCEbIzBp4sy161aySCZ4quS6pbJFuUZOHgwKDE6S
mkOx9qfr0RXGgPC6s0ZS2Vnoa6fyusIRO7xkZLyv5VpDtJYGzwcelI7E/JhN1c/o
MwdT60k03VX4OpgbUVSTqQ8DoKJHrEvIaxSOHw4HqfdpbFWTZCjXtL2bnsWeSYmY
ZOUZveQMk7fn011XwBcOG2DxfkDnQv2iKAhbn5MAqVPKwwLkrMZ08I56OZRGCdkl
Wj/r1JHVphhqv/3Jz+n5EMitolTa+KfIkmFDwLC9QCFG66aIZkz6Xg9fp8ud0Cfx
hmeBk/qlJKdwCh+UlOb1TL5ruDOJp7Kh40UCC1Yu2ULjDPHwbzaZ6DYnqSPM7OrL
cGwnrLAqc7L+BVyrb+UVa88fjpPQ5taA2T0GfuIlnsrY/gYykLI04FZ0A+iFdc9r
qcPhYJJJilhPbwRaBFxo5/+lkwP8LdcRN60Kyx2H92z6yUCLsBhGJJmXmt99TZMV
DTKI6y/A1FqE34REnLFxZ1HP/xahuP6A51DoQ9qMXGYSu8rABNovSVRDEGCpIPtx
xqud8Ir7zqcAi0ND5xy9FEzAiGtCl8GN6eLbOln7JaPuoBJDCC+u3oVBCZND2iow
+XavSnuaxqMK9QyZTmJNP46YGEMKGhKkudq9Y3ejkdP8PupH/lyIDh1aHimWuvLW
5qm3Y69soMGJvN5UQQGy+mP9cCMo0Ptu9r+vJCoSsnq+JxqBnUlULzHgqCiSQjlQ
QbxHrbBZlNnbh6+6VU76rm5XD+x6iblNdKik1ATg7HibogVuS1lSuXWtpoPL2Fmh
fIskwu/q4NmAlkwLet3Y1EBaQ5XIUoZ1kxcUXNE93uRj+EDWdHH55JwBYq5F3c2F
AAJeRRiOFe6CvTqUu74IY//XcKIILm2u8UiyowmfQxwX0ePK4Mr/oUZkxuLMd6D0
DFAl6cTsEHPwyClUsGxM4YrqmQNK63w1VUFZ3SoX3IrBUpl3m9jNGxfN0x60EBss
I4sL+RBM2LEGtIAjykn5ACZo6ThXnWaVAHL4eqifm+Ch+S9gzWK70fMVy6xyUCa7
XP8hU8BiVrJUJrqY3XFHWjs3vIa7uU3pfHZ5Ih3BB94vXPFMAgUgN3uoQ+WH8DcH
T/ISazdKnueHPkygXuku7KhSsZV0ZyHQjnzRQrpB39aQz4oORz+dsX8H3gqIlyaj
LX0jBcvk9SSpC/SW/gJjczRY0ra9zrF+Vk+Xqn/s9VQmyceyzAa3jJUEWL0tnXyd
Q4aky7B//xKaQ0etOG4ImixygOANRe4V9Z8HDFCLDEdtdGp6Guc36voWyqbghe8J
4008oDNdujgDSxRGF7jcASvUygsxmgu+rCh3mHrf/uE1ygWTF6rdQhNdJaNElrXX
m3b+EqjhZ6tpY5H67nWHvlYp3FlG11/TMPzOG+W9Of1BJfxh0ITyX52z0fch3xNB
yn4jMTxntnWOhjwsXK4UNTi71X/YILMzLHGPHzSI0rRxv1XTi8ZR3KQxeDBA1EQ7
uUDR2tSuPwNNPBWQQLxEHIVeGNtpBXpvSg/u2Jcbi6x6j0u3//muRixQ60BmlI6e
yskDAe8hDRRo3tHn8Mgsrw==
`protect END_PROTECTED
