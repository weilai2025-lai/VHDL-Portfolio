`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDVx7Eev3hjOKV+n0A92vkBmM2cn61p2aKKDlZ6EtJki4noYgoVXdigJTB8pKhsK
yrtBqQIKLSR8WzTfGsLWYzglS9RX/eRz9u8TiGCobkIEWFk8ZOcfJtHV7ZeBFiYA
nDB/fnPnnju17r7i7071hjdVnmN1f6LnrlSNWbCtkDOfcROxynNNOoi6uCTp4UGA
QvYWYbngRu1JxMlq+vS3k5v+d0+1xUNgFMsrftvsEOUj4qq4nEKjJf4HCnX5Nroz
PyEoS2vwqnyp3+LRaQLx+9q5e/vEhwRw3HYkIxLdwuTxhdUJKcXlFNaiWRzdls2n
NQMOZQS5ZE2AMpTNcHodcH+l2sCvWa++gYZr2AR/fazYVZMsBV7MVyQoxv0L7wqG
F4/REMUhhfgNIofW8jEI+KiMAqOuhrr4koQ3uAH3U9QAJJDX9B3fNKjqn45KVQTv
pRdRbMq98WpIUX4aQSsvuSvn5ZVYjGPKutOvijVQmPQAhKjAYmn27h32vAqnw961
nUUDdk4sHvWogcuiMt1go84GspBPpKk7pnTm414cIohabGGIz8k7qCN/76rdF2vn
2rb9Zn/wbZ56ioS+5ASBE9RWXRb01yjo37bTnMx+rYaddpu0RAm0yTTcOAk9uO45
Oy0E0MQrdYBw0cUpUfEe46ZH/xsztvO2DhYjLnpK0chhhUUnSfO0JHRMinINlJ9E
91bZyWOofgmN6MqYpQL7t9yZy6OLQZx8rDLIR8+s46Rhj9Ea6+kUlh6OtRtewbxZ
FfoDRkUV1yHn094kGNfwoQXlVwjdrrUsHW7faguoNA99pDg62nX8HE8OpDIwjpjZ
zwsk0cDn3M5sLmEC3FN5MdpGF/SvNPkfQAdTjzoHCUDQSQgApBCHGeFZ2rMFtoBK
EveaxFgWZVZFY+4HXr4H1iAj0AeRR1xhmQSXvVErN40u7OGHbIAv3GoVrtvCqFGJ
lxbNrhmy9oYgn4qHC1IKfSPuYkqByuLN4Pp6bNYnfsHVbzm04eBPZKTdT7aV44Ci
Z0NoeXPIL6JEIFo+tJBFgM98qJUeEQ6FLCII6lT/ff8iqgRWVPuYNqaXLJzK5P/O
SNdxRbgHLnDTeJH4IZaxt+iMYSUhVqAaZmaZTveTVhBJmhxwVfDIrtydVUsxwVqh
3EyUAUHdLG5bab33YTakGYjS90LBzv4ihK4ypxv72PB3udMGODeVfwueRp0tCaBU
7XSF8lDIzDxQkYQdP119h60lryHrCAgPadVuxs/qkCRsueGF7xmGti+kS47xDlJ7
JyQcTiAPnJoOX4yzasJ13d20MHRh+pLapsYSgNMncy5n/qmUrfFlzIvEmmv93YOg
3+F7gtRTUaZS2z1xeqZ+28HsdpZIWllrEjPNznZhfaw2W/+r/QAu/f06/G4rLIls
wKr9umKvdol9KZAShik5hEg5gmDE1SdE8YdV5aeb9Yn1FAtnTJ8voNwDlf9fT/DB
3TOtIdtsWnBU3olgxv9WVPiDmaS47gUx6oeHcpH91DHUcv0A5Srn/+4uCcIiopLu
exus7hhRDQ2dpEJLiRxFZgbst8CFc2zkRY3PBr7zl+2NdoEb92pIovoOWWkY+57a
iVP8bp0BD1FPvScr9orlqy4A4vPtWtdZEJ0MrmnZfQWvnPKxysFICkRQ/JuzfMj2
tXGMmkykPuKK8SYLejwanUp5MqeR4MpBEiziJzlbhXReC5q2grM3SHnY0g8mI/Uo
OFIBedCTUduUMdfVHmsKeqLx0V0/vPar1a94Ar5mJovdWJIk9mbQAXZuF51n2U1q
/pExdSuF+Ip1Pp1RviAzeWuv1ra0iopLmLLkUNtpFWgVji8E1AmmX/9wDq1akpuS
syNDYppIhSyf2kthGPrc5Up4oUECAhfWhKJezdk0kht9kPm+VPX9F9pqUPEJUkAw
YfsxqpflS4lOGuIfJEYVt/25f+2xsD0v+aHMXgBCaGZsKbndjoYmxHW11V1/wUwb
t9fqeCuZWGp8Liqn2qRck9WYQ5glw5BLKrWtgKNMe0gII1XPwgjtxoYboiYl8Y3V
q7N5/sFjeMkiMpD8/r0U18eWk7TNzp4kXYYtuuC0rt9/YWjKsXRGf5oX1oa+2Ddf
Q4iGkaojczwD7UYid6cqZ3DH0MD9KrK2LeqpC8EN4NoL8RSR73ruEx3pkLPe32Mj
i9XuJznqwuSNGVm5uGUCAkyS7KvpTukITaLqetI1q7gSSEMxk0rkDPbRI/2+3xJ1
52IOmHr3ZUQJX1uk6nJLx3MEr14Q+B1IJFzdJJHc9CMOSDYF5tN42K6C1eoEzgsI
bUAMx56PLUU8uQUP6DkroIKdpcqeCmf+oftNi0mEiIb2Ooa4Pha+ea7njennTfwd
nZIuXEV3JeBSLfTafbNZogKRYZazC7dAvrW30kf9n3fIvOeUjLdRsm/V52/UYPtX
AZurJS35K3MOmVxdHQp+k/haj+aLRo7F4heTJ23Je/4yyiS5bQjPSCpLCFFy6gGr
KrkPiOLNzd7tyjzCfJDlFpZ4+onHF23V8cnr58qNuDlyOuFXAz1eNtOCti+uFQAQ
d5g3Qs+YW18TpaPVeGrCBTve7Lm6H4eSQhx7QYt+P9vUPWhmVgIRKPw3YaR8MVAU
XlL2prHtby0/spBHumYAB82tonhts4Oi8TVea+CC87yczejXYOHcCEY/EJynuG1X
JYguriE21j4tOCqR1vMqW07mimFTHpcsKqpsFKM1ig3ogMl9ax77BnLAzu1bYwET
gAQiTIRX33eaY56FRgVVWIB0UkqTIO5xewvl8hfJQjcpARp77aHqJBqNRTtbYNaJ
qPwnie39VpKuvmEHU24xQkuxFpIcArX70pybYzzNDJu0vhoydMaR09+giw57a8/R
CayznTjgv4s7BHlvb05zA7QT1fpj7OYUoreGZ8bNncEJJPhoHp+b+mYlGwwW4wSS
66POL/qW4NZMCvpDPfbbIQvfCGgMdCICotRStt6j+AzHwUHwx/Yiswkk9SeJHZ/u
CUJ7uZ/pQzZ14yY/6zWTN2eh9g3gHgHzuRoEWE60h97H0QR/vVwwYlps502jCj9I
zhCQbRgKuv/CPQxWJI729kBm0UruGxo9YmJ/+KMvRxpByaZ/0RIjnJMtBOA2Efep
56Mb5vFVddeaXhfvqVTHRXxJgHrk4mdudFY6yWpqQFfzetpqXTqNZmH44wXh7WIQ
+lWcyIRx4wnVubKhSEDi8chiIdzYaD/ljof5gAIeVTmff3ZX9Rf2X2cEsm7r6x7N
nmNB/Bu1PV7n52EWtF3CHQjtqn+esJPQb+p+9e302DPH7oxSR+FXg32afPD810dv
Zek9fMwOzj3IVQjsOOFDMWUKMiu8CUs0pMNIIhaK7pwj+th0JHBpkzYuSYy8oFpt
7Rdt54pCV/0oX8FQ4hk3SNJ3JZdLYuEEmyykqBF2iIfFfzZoMxaM4eBOqefxVkA/
sDa9fo99LDWt7P1waKsY3VRo+IAhMGe9jrYK+hRR3/ri+k2f/3xNOHmtYqPESv5u
8nxyhs8njf8g2S2Gj1+qacj6fK1LHQJHlwYdrEYktZ6SPJkXX6vBxsrvOoCULoEj
ZAlju3VsLbDNdcCY7bc4FjcW1e5cZESJm6vFP4YC4RgcutR2RJL8xo9zkbtWlmbf
cRxv9A37Q2Hig5ilJUvtOY3owa8NvpWpM4TKa+mj58gN+e5+6GBZLhCIgUTpngRq
wfWIcEGecVpUw5dEZwHkEpn6RyVvrDL63Ik+aX7LNZwD3TqA2kxlzCz4f3ZuJxGX
/O7DiD6z4VwYnBJT41kYubEOShFK5I/CbOi8qt98UL8y6ixWzmxzr9DZwpaupa2q
W/5SCitS2aigYA4k8+j3q0hohe+UItBDVDkqs4NEescj95XfbXS69lxlwptDPRIB
QdfPmWK+Yw57QOjFYaHLEJkBpfKi/TrXTR1sjmISWDf8hdueJDRN4ZaJb5G9xGzG
+79RWF08k5v30bvjK2A0f2tNmrDOK/OPj7r6Pd0Xjx5Vlha+7g4tKSc0celH8Jjg
6Yt+NoitMvdnotu2OZQF2P16j7Umdhq15gs2693FXbUoJxL7AMS9cc4epvp3pFrV
EjsCf9ArPX2p2Xv0TUmAsX8LEwPV3TAVuWbCnlp7HWZvNioQ13JE9LF6aLOaCVU7
I26NlQKH8qAhV361pRRXiXM5ADKxAwO33Gd1BR7uYrSpIqArBIOfbL/TRfraoEmX
VTkvkPN9aciwjOTFvkR7xn4q4l9uY3GYhA8c7b6FdH13AQv4qdt9SjeQrqAvxEFU
HFNvrlol2k8RRSE/pPKbvjIIvqlNvPZXZtVf+BYlalLQaufJ3Lv1vf4VQTAgc0CL
TI7mRHMOOp7zf3IJTFlDBJ71p7qRTBkZITapLzAgWhMngF7NZcIObEXfQKmSKomo
vE7cXt0bBVlOejicBCaYHG3Z0Gn2Y5y7LgK4RJLX/QWfTu9Z1Wo5/liMKoltg5Nb
rlHWbnmbLQeS+IdGYIUOCJpGgni9I7VXwzqiFKnWo1y14PNAp0I35zVDZSrJBKGv
e2cnee/il0im2CJkYroPYxz0GhRFjvLbM/oN6B6ViKP8OOFySNuEQq7CNODDFRiU
pdDHeBRAI+wfSKKiacdwg5UFAStdctYg3N+uW1xsoTHsqZjYXEB7OLq4d/bfNh6y
uM2cV/BIUHk5c1m/mucVScr7YuRl9CBg+5WV7epTCOaOJbGVBmM9ANGJmktMSESB
4CLtCKRyzbKZRDdH19JCtJHcbbsRNKT7lTLRV0YtZw6/4IU2vIO88+TCiz4OyhM7
TygbwjsqmvDM5uPvG4dDGiiP3XtRNRdoXo/6xNGYR2ha/iRlhuVfY409p/JB2B0m
SN4ab7AUsmLofR2uqcdy5w7bT9CRpG271p3cJ+znn10n98BhSJRFmnixAxMYzZBf
husKGFi9YnvNZz7Jt8v5oOvXgxuOsx6Sjz3MkKB6aqBroaWUzMiTTdtBqlcr+jyt
JimUb1uVLBV2zmWkzlalQ+jK9kt3kclPQ+E4UXRkC5A2kITd4XWWNZkXLYV2thGS
nOZWpkAItDa9EiNn/YLV3MoBj69c6OsqMbBhTLZF/dxjcRLwbhZV9tWnE3chEzTC
y2edGMbirJqMPTl2w2n+skUfxdxu7CGweBbqdp4rMPW5fKYl1gWR1R6Roqt45NiW
OARyOfrPjOlSwmO1B8Bwyr0dnWyMsUwn2Pr2409nHRQgguDLWwhlEMcwtb6OWKD+
/2OAjom0RsiY/Pni2OeqRHzVowoIA8l0XCGWGHPRzHU0f8EerQOOEuvTEZD3zeew
bBAI7mMtS2RlRaeg7TpW+tX8aOpJdbVfAV6TbswY9j+6AUesfFkLQE7cf1buJ0Ha
KBZ3lLFOQMU7sduc8Es/03lpB7MDLSRehxMu6vAjQfRQ6fGShPutj3FnWTL3uQdU
by4KcCjpdoLarJ4cX75ZxkEmdgcV0Jvccysl9S97MR/dD4ygQk76RZaeZT83AVuj
iN/YV7z/M+bzx5S5d6/D+GBVZSPbgHRst+1t1Ljr8u5k6X04AsLZ+mlTckDD8U5h
kCIeEGm8jtEimP4EKGPipIf6/YDGiuCvpwW48ICHauslZPrMwcJ2Rb4MBIyqtzN0
WdeXexRnfMR4wPyH6EM2BKP5AC76+gBru+KnKrVDUWz27zGhmzA41UdxSell+oVT
7fdvxflWnv+/Qm8PyZWcLIQ2REi8EF8t/3yFmr8xAJI/6OGJfAVaPPgFI09A12QB
yTV6x7QJrmreIHup/3o5G6h4vqZbYMX1QrPscDpT4pvT52H6qwiC8naGv1e4iUCC
SeJfm2zKwk9wG9J7HUrOWvEdFyc2z05mUImiJjnTZGjhjEg9YpzpCr21UMoL6o0a
jyHPnp3k8PjDca/wOO2eqIHsEDCp6Mfo5BMrmvtidrUQIdT+A4aP0Blxwzjvz7X1
UVPTE/3LxwLKex7V3qwsee2L7yGPVio9Z+reORTky/zBSImXkHNGALhhyS550GYt
7hKjut+RK1r/koCm2d0/sF8RFBtd3CfxPJttq+jjL8D7SWcKVKfoM9huPIDGjWxk
SE/JHfO2WAUL5sCIwEMP0lhuKHL2iax+kYsKhL9eNG5RdwC4Oc5xxEQzTdcDY1Lh
IJgnRRqTBwBDvrowYP1WA7t6oVgRRRy3aJcEsb/YWfOutqioUZaS4+1SSjEkuUMG
e+ExyDiT6FZ8w+XwDDQcgWsWWOPQLY+BDjEZzNsBmyRaLy5JcPjH4n4QDKO5HcKZ
AKiuIk73ELg3ACkuC1IUzSsa1xA7cbcAwe4NpSpVvyueyFEGblQMPR332AXJ6O0I
xDoftadeT9HdeHDO/0cJpCoVhguJshjy2XllEYNa2f+A3aJwQZSRQ3//NYnv/rXZ
6xIQZl1iTb8ZgjNP/iXSJ9Hyy+cXGqFkiUvUfgoJYPL1cGh6uJurGP9BY1GjartH
W0krBzBbm8UgPvUif1NKDjzVIiCLCc4k+uka2bKRbnAxXjVMkiKm43LQnZjR72XG
lVVJ8fi182plX3ClWOgrqq/477CncV2mX7zqZmUreEuLBMJEb2puvCK2yQPZpZDM
5VYFW2Rhgqv8beTZRxZ9mxhl7I3QlzApO9+jfizW8O66sreo2FGkoGWtjp7SOAjs
CJTk2mlPOz0wEoESca4EgJdW3OszsfwUcEo7DWUIrLKrNrixRZxCzX4xBEmSdoAX
ZeRPAnH0TmHWZU1rtLJ9v7z3mD4g9EaAs2iwGeT/RoK28cIy9I5qPU7ErKYcIqTF
pT3mIWeGYFiE8Axtmt0WVNngKkhTDLWWWTjo2ScZLcyW8WjeESFJdIjk4sXGzpsm
DkK9cmvy7/GzQQweYB/RutENJlpmP+zXNdJ4Sn8Bz8G2ECLXyZT3VCMlrnrggZOs
W8vn3QcbVZsMo1+OyBHize2Is7ZES0Mo2Uca4m9v+4R9HCnEEWVZgFXrF/BszF4d
Zdb4CxuvtIiyBwtww4Ul0tkoMJW9oTmzAncQkpeGNCzBxjB8qggo0O42r+YyPwgk
c9IPBGxFFRXJFdRrfZbbRHFF5BylGWPAhzUR+NneMK/1gpR2nBEyCUy2XNqzrwHG
Pzpu6Ph2KFN2FzzAgpZfDxoqsdkW9Cvrg+pzEa7IKT+yb6C86YgL2GiExVh6WvJr
hbZkQ9VPc4j+m40h0mEdv+krEwgSoZBFin9ZGaMpHWBWevlD9Envu01TD2IPT98j
7CQgm+f7nhxhWia7cBlAsf+WTOLCd6Wop5LBsqpYl5b6u+i89I0oodnKjasyzQII
fR3IwSY55t2+QedDdUlgxe83/KTA4/y+BYmoXvTWlgbXatuwYMg57HsDv3S9Uhr/
wQPnd+sGNyPan/NFAz/IubncHMB5wYwSgFsZqca5WPoKmVlsWbqC6TB50sAOZCRP
Bd4PrhQcygrEZer6mzL8CPLw6PnOJpgEtTLocMUPtJLrxpLQpyMFokwq0/QuoxD/
4tEzjUX5RysBMSytUmICaaH+VGM0vMrT8ZsIxao3vLMFEsJWdpvU8IeU/VUFuTpn
I0k1rwi6LoUxPBYRRVm35JIZPxoVRafr5hjuekWK2iR8vQ4kmBeiUghg3W+1lxUi
0v8uiGo0pVch52F5rJsmUhduHJyZimyTrHiKvpTbrRLDYbEa2ghsnsIUbuX5LJvC
sUc6xjn184sgJ/5MssXuAvTxFUtOmxKlg3r17OBEBa98bzJW5p41zGhbzy5/w/rg
A4X6ZUwAj3F+0sm5uXBWw6rIvfflp+r1tJIsOWpELis9pl5hQeI+4USQ5ArPM7oB
JOartu9aKVSAPmEKfbHq1U2+rFV+uTPEGJ4r8krev11lHRoxeWQU8Xp5BXcidQ+3
lJ0bcxwkA0+gEOT8bygOUjfhKrgmLj9GYctgmWnKsFVYlrI2uqUgKCCfeYcbUwIM
RMYUJZl8JPhyMI5M2J3m4JaoUccXi+cYHR7wpEgSVODKdUQ9w73FRGNngPDXhgNW
uUZscBNUxra2Qg7EqVYEeESaqRO8BscVvS2GWSNexDDO7mX+3iB+fpiVxN/ILTTX
vJy+VprdlGs6XyZXFNG23F59bSqL6MjcrUCmAw/md+SFI3yGroXJdtgaq+ZJ2lhI
lYuIReoL4sm9Ct6de1wCenDI9i16ynpJxWtYaFB0VSItk+l8snD22f99iLv8cqj/
8n9W6pGTwRcIYcgDMzVX5E7YxMpmALZuFuQzs3wtQn71A9D2wIgWIJEZyIt2mWEp
7i+U8zGHNoCWPdBujtrGcs1h/b05JktTqO2lSRO5QhMzKUQ+voy+vmSGb3pPctEM
sSBO80s6bqfz0fMXsq8wwqThdbL+nR/zCz0wcjifDSwhf/AWDJxK1YPAKCoN3H/A
ApwehTzxqKq93Brm8gEr4zi6rPLc6hICFsJY17T760GIKVgDQKPzg21W2NJuibrs
ulBRAFKCxGeKWg3tkzSIUKfATm3SMIyOGC4ul5ScMAk1Uv/zKxyGb5aaIbNC0BPg
O9RlINwzKgKPBcw7jmZKd0QmPtCXEAWyBDUpB8oGRfa45arBxlK5Q1DQvsKEv6Ql
FFhsuee7Qdub/M9Sl6nedsucwvLKQXYAI7WLwXU0s61Y/wnq84a+4rUSoLnbmUp+
OkPSnN+FznLmO3jiDG/Y3VjegCM5cNQ+YeeAvS7W4ufDjnmSnZv4rO43bu0dG/8x
n/6p/+xpJ+ms0dgBY7hTF2V55qQQibUT7jyujB5qxrd80Mir2iLkDW1/vAzhhRPP
y12jOpM+R0OzoRgn+tRzK4/jZtKn5miS1bjlyBUqUdINvaaEwkaFTOu1qxDkSLOQ
NnpXvhgex+u++SOv2CtDarfUVDx7dCWilskOeNHWbpcyrHce45Q3mJO/GKo0o1Mi
AfJlUizXibOE8gxM7nLNJMCFXRP/gjOOoyewN/QoNJPxZ4opIFPQG+EZZeex2i6Y
Jx6Zl/Zdk5y85EMu1+6a+kb9wSHKQ0rhi9z0F0ohBA6b0nEYTe8+rjuUMTz7RQ67
hCj27t6BkBsRMOSAVNxyhn6khz7u60wnEG95y00/1W0zbf+wb25zSuTT2vBJMOxf
EgQiiPNTFUB+ctazgPHnSXKvMAYBTqzpyvkjmbWykW6M2Vag8rJHLFgUg1INf+Z9
pFS2yjBV4sNaDn4ZjPAWnrBMMP7GGONjtQaV1w0GZlcJy7Qa5rCNRxAfbaQJuwqx
wNf0Us7RTA4ZKOGzYjpDxyWFSkDeBAHUJl9P91T/WcflMdkhoHUJJ0tlIPPBFwuD
rle/rJ301+AxVaIFunTLuN9uXdgP/5qN8tvLZX+d61vfdv2TnSzWxOtvp7NnvmrU
CEFsk5Cfaz/5JbhuujP2djwa4GbAymnhk8QhkXWqroSAsreYCFjPLFPWbdmDLuz8
FCfg8JawwaJrCMTVkbocOB6aGn1+6+RFnJnW6YXRBAfLAb0JxRlQhzb1UNMPSK9v
okPiNaaIJ+cdQigrdxAQH4KTcO5bsvn82v1e94vu2D7YTW5e59PGgVF/2tOvFTHg
89rUhyAletuSCaJclYifZ+0Ziq8kQHvjjLGYVpBKo3fy3F6A+2Ij5oVCCbO/9a7v
qvdaA8AYEfLWjt4Im5RISP00GrWLWrhDDTeWvdcrzs9u71MkoOhQX/gz2dgBgKyJ
93dzIp9+L4bBSEGnU22roOltD3uWPPEi8/+ZHRcikk0Ve3uuOU3JMYofhBVON21F
wFzZ0OG/mGmuzHRwHbZWeNdhu8Gu9Hhfrxa+b0gytFxsR+z8XeCKN4oGRLETJDb/
xhTwSuZiNoZmuY7HwZnyjkThn0WRU++eWRrHSY8wZegDL/m7HDBMRmdHCGDeSHEy
aE5NW8GkB6EzME/5ozq7gCY3+C8uIMtnybG8Zy0KAeYkIj6K/wWnu2G89ChjHyrp
vSmUcH2xcCzyfscItlA2WBtcjn1T1AUi/cu6275NOSps1Ei57ub2YNNpvYUaIlW1
v7AjNe/qT1gGzcIJAUuAdGZt+es3LDbhJlV5qHqcvdZcC4jO/2MGbawyCuxE9Y+t
/rB+zIgW7QaGu/LLuNt9vksrkvW/gE3+UHqIKIRYTwsYclTmzPLAfBVHWOszqd7l
n+o15PQm9EK727KJAyswOB0YluKuSMHR2hTAZu4qaOTiKEJObnouD/ZEodKMPByb
BxKVp4fVTaOR45lPLqCpqlrYpstm11dJY0NpQNbycN+wSH+Y0xr5JlezQYHfqe+U
P+4k54/TqtZyh7vjarZVFywkZcj2DZIKaFVMth0VjSkadDX6Xx/7Nz/QtxVeG1K6
ZDNI2sl241OLqUFcyaPY0v6Z2PbzYluaTgWcyGS3CirJTG0h4BVKrDiSla9dPvib
TSkFPqHwp4lfQr12ffaD3NfK8m/WQUEfZuSOTtQJ1PmYS2SLEV3NSGaKAJxWHRG7
FrU01Q9RfF1o0vYyLKgdN2KjsojEOMP4z46HFyJEYHr9damf4XKqvTFWwD2/KkCz
Jn/EMAkPdxx7aK/B5w/JVzj7OlBKBPNN9aaYCWTnVHZAcguaYZC7SAUrSbh8wZzn
5fpOWs1b4eKBl5YJm4JfSUecokG/yXhB1LWvrKy4WfQ04aDlx8QSGjK7FjeQVlRF
IbSIyhRsjg2HWmMhH9clwUnrx+8YB9XpQhdflnCGBYxmNZRK/itrBh9umEZkMML2
FvCvoWmDc64Ap+oukT+xEV6jjY5jxmjxV2prMKDXrn6/qkXydznfzPBWROQ8r8+z
VtKHENhex2GUL9ajOVoh7pJ6gdMFUKKTjajFu3+OFWj9Wx6mWsd+x88lj8xoRVcy
In664NJDBvUOQUDMkic6XGXYzhLCeX2Eb45UuoQn1A/xHuROM16vGJpFWIRBemP9
b5ILEgoI1wEr27Xdhm5+9o9PhyL/C9fsRQ7VAV3JxkyYRSHI77YYPfC7IlqE0/fJ
TxK4hLT+TsGA5fCcAUiaW8U1fw0NGhaOH06hEl59ghlVL0dLr8XVCfuDuCaIhMP2
uHi5026GGPS1YayhNXaCpjMQH00pFLDHdDqnCxKke0nT65AoItUU0QJ4WdnaoZaw
rEKv15Tlr7U+neBkhy4e1dloR8nZw1QR1AqeFbJhVO16q+H/eCneB5dp/LhYgRVH
AqGWRMKj4YIclj84q1gKOVYNKIOFVTwN/X9V1DBxsc9Fh85c3UqFPbWovi7mrpON
gVkgDBIIfwC1xNjSFNWvPk2QaRnwpBVBf4RM+Zkr6kAkxdjx2rF8F60TiDjxXzkK
6Qq4LVuD0msAFS7aTr2Kj9dsm3qWwQCVn4dDl+pG0NCpkVLaHLxwzYpY33dtAbSb
G6Wxfs7Pom2rLP94kB0QByUuOZGGmE06Fsj+pzY24X6cuEqKWvbDN9RdeS20fUSp
kqqrGgI04nP3rufEKYuxBYb7ifSpe/Lr8z2ikNjiP9pO6UoINyg9DOUBlFstlFUO
WCvqHahgmOI9jMq/v5lPkwjUS4h6Ud9oDc9McauYfSxifaVtkHSycghOrCF8vNAe
sJo3prXfoi320i/SKami3EucUYagqLXgQ2LCgqPNl+n7lFgcPr1vBSNFhs5zgtZw
TraQuIqmAWBl2uvkUbttpoJitoo4e3KppAYoXFKGNoEX1JWsscKX9q2H8WkWy4i/
L9rImFRhz5YhYJrWtKmRHROlUEB362HNEXbJ1uyJs0jcs2sPJ29TwZMKYYSmKqRa
ZtaaCEh9V5I2ZVWZxrouqvnb7fvv3ycYxMi8w56LrTK/Q2KUMejqI4guMH+7HQnx
itpywAhOuxomRC5zaNoG1j9LLczF+zO2FcUamexUbhz9qRcHiyN1VZMfO3WFdku/
IAPMvDtg1WoiytE7KDj6ru8LrLEdKmagO5Vsfv2mye1G6RBW+F7uOmNOkBnlF1nl
Sw3Ly/s1tBp/7sPURvuFut6FzTVv2VmWaUD+ynV/nOZzhs3ZpDEXNJaoaWkUPnu/
TAoCB7P3rnHp/o27nUBbDURs454r6aU4vbKNDShVS9cgPMLtDtRDp8R7o3wAOIS6
kdMANz4lz8fQh9qomJnaYxOXRNqql7Dn3wSPUJXY1x3jB2iUfbBbTjHaDkUhrmSj
MC4vzCwV0l8f1+ehEgDISdEJGLqFR+lUMPQmicLsWHeD4sT+UzFWlbN7ZKHHuEw+
cW+XyFPpj5j9YovFiEGetiFiJVXxcllE+f/NDdF5N0K24EYkpE1O3iDo4UDmfHA6
rInbqOzGsrBl8+YVnrliwqhg7RhxP0RcUd9tgR82LAf2t/BT/M0K+QFSwgmSuGXr
tzlSPc2TOxEJ6GDQn0UhLxW/Y4hWC3mtqTMYp1CuYXehA+Gb/yYj2pJU8bFCXidg
9UGJYH1F98pWbLsUEJ7+lw6ZKrVxfIvJuPh/6xGG8kWRwqpuscBp8D1tAGb0Xb++
4+otaKY5I4Wc+4y5OmBd8EPYn1yjIM/WCCT33xpChn/JNGuUXxqs49OO9/GTF/zq
vaTmnEi/k349lvTrcYfcE41kx0YP2SgBOea31C/ITAVAdu90cegpU9tlj8KSldIc
/OqNpII4sds88t4UcjFJb51NcE/9Wic6Hvns5uizd9KPwSXB9Xagu5bD7h2IJyrk
acYHWCtdij/dJr0+4GsIhbjap/KJXjXpAbbJyUlSDWXRXZDbVtA6C0VD3GApjHEI
YvEbYw69zaRaq0JD/woxcHdfjWto/98Sk7uUo7Goqs8JDKqmSBPqe5RjXVrMW/gs
rsfdT9biE/MTI+d78hBuFcVNobi9Md2xLUw+OiVRKblNc3j4d4Q66q5sVq9+IZkV
3DmONh4iw3jWgBySYUSduG7Siqmqm2+1qzMAdoQoLkJMCln2NRjmKQxdIg78eK0d
GiAEDqUGkIErghQ/GSqJ8rgSG+FaHOMVL1DX5OcNb6xHScwOGu/lzVMiV1KwY05v
kiqVyxdtVKwPfwGAw83NfLaaNfldCI42sgMB5A9aWT3Cx4EiFo+aRGVDf324Mvzi
wgSO7c4t3wi7M28N0ZcAiLBec3QIauhFiwHTMGZzM1J9Xjp0+y8SwN1L8jOSuXvA
omYfQ0GpLm507sW9xCtgHwN9djGteAD1GBm7qcnbWUufjspje+qZ9Dvegwzyi585
3mAWe7rhla4E1CI0vKheF93A2aigW7rGePHdKk9UerPgnfnx9YZEHjYUiQTuh8bs
JDUEn81+GP/J0sXg2eyVl6kFDIGqjX4H2eQrHKA5WWHZbA6MGqKkKZui0q67eLsc
KHhzsoSXMM1PYrl9O12wTbZT2MNVJShweTgGWvL4Wm9cxPLRUm8TiCG53m4KBOM9
MwhGKUtoelUXrQNuoQgLZTedf35ATk6TJ9CcsdYqhvRR47beBZ4x5UY9LLp0ORSs
VxdT2/ElRnL7co4zBqkuTU0ii6xc/k9HKvjH6YX/JZYv3Rxd7dajd83Tc8iLhgIF
D6ZGCiZ4noSp3sKLSc/Chj/SHZVKX9pgCVYGuyTKSmWIqYejfM7Rf+c+1etvPuYo
figBiQ3MR4fnsqMgMsP2fnVIBut1gp4SWTpDml/KxJH+t0+8xVHYfPkUwVq5AOga
MJDG0WiEkm0rF1o7AozboPsjjOiZcH95bqvW5kvphu4BAnSdvS87FwWqlRengqSK
YZqhLr2KGcUIuMQzCInQvq6/oD9jaIS0OkPF1jcKyawc04bT99HzsS1vbDMkEixI
IggfozabqcyI9ohpkHM+1H+mCX1sHTjDkco3/ju6b4GJNTBr9WSyc7+Ntwit1n9f
zOvgkmtZculNhYyJeUedAbjRrmRdFEnnv4Jz0D1jUb669h6Ml1EGRZB9R6N/dhN3
5MC5FViI4ZDclvw6JTIK2cLG+QfrbCE+6vLXBQzPqs361AFvIKB/RIZT1Y0luA1Y
cMuskfvVlm+EWLQGtg6reMqL/SqkPYFQhAGY32LDuTlhX3VrgrzNGaSxWMcbQa7u
UEXZk1D2izHAVFoGN/hujdwGKVATeWQnsZ3dlRDlx9Wg2Bg2XSIQPOF19W2BIEng
OJvtDSunMrRA2562N2Lcsux0oeR3TbY6/TYsAzA7z0ZWaDSoEvq1AwkHLm6AqCpo
C4MjC70hpOgfdmHp6HTFSEilhTXykgyp+hc9Ss4JAfNdpuThMVMWDx/FfxrjmuvL
I3SiiFpbidiy8sfHxY9uHHZDqVO79RD9lkQBvHneIHMF01KlcI8thnWMWLytXsR4
Uh/Xg5ENCNqv6bNvHtkK89pPu4j2nKgeBgBZU18bZsoLXyjKvrg/qSL4Ns4cnqGY
sUszYzEx+NzU7OQVcl2JCsEVsWE297zN8VndBzlCPGP+fWfAjlGGvk42yNP9cB8x
0eYg9c9j2ozJ0t1egPeP8fsdxDQlz4uJm6oH9v3qLHDalNMuJvAvTHwc83cCBoxU
lphFCwo7Mt91g2aiByHSSEkjbzmzJ4yCjHrNLN1e9kRG2BTzqco34n3HcqEZuNMA
7KsSb9Eah40xvsrEnmhoVaNl+GgoEuyP3iqDzbcZYhNUPec+WbSQ1oTKdctJznja
P2GYIXLdrErnl3kIeKukU5my0M5pbUV3NtCCTa9z6I+lWaypSyJDkRR0GjIvXqYW
bGw3uqAqpdzUz5o0IxNPXmtFDgngpWRpdnhJLURVf2Qhi1ZPKlcrC9dZB5od9Z8Y
LvOi1BS+Sz6fOISH7iyG/1/yHSc3w5xSFVnui9Xi6lXQGlGjSGzw8BCx64GunxMP
KcHXSD9emLjOF0B8+95/D+HZGInj3yME4lnpT0pc2ODEgd6xIsPpWeCaPBuBQuBP
TnY3ym0tXnMua40P7+dQGoH4m5Bd3UKLiNo36MR7sgrvG7/hdHM6yIrGdKMPD8IW
epwaQsHO5arw3hiuS1RXQvTJBLsCwy24ONCHzh8Y/erAATgVQBTDNwqR+rFeqMAw
qEF78ugosXRepABM8fQosUcnZ3YUWh7ikowgDgI9bsoKZ8e6GBm0t40jNtNXyDFw
ri9LhnUYcPgqWkVJTQWlNXZTL+FSXgaHkPWawC+FjP+e1A1S9LIgTW93nNVC++RT
UFsk7sHNF6gsfnrpTSXptUVRV5WbGDmXK2S7WUUGIzUeyekqBfPLihV9veowTYHP
/Kpmp9C+NJoUpiOeCRI40o6RZSp/t/sbhOwFAo8cV8QxQjEjWdFc0hGerW57vdJQ
ekTMi9JaNcXpQK3FyL5YdGa4vbQc8dgiwUrRJsgxt0SZVpAXnFUbA3FaYEWge4FJ
V8vnrIu8zjyal/gE5sfm8zCsygw+f0w3EFoSr2++uOP0ZCuPoeaemOOabhLlt1iW
/a622sX4KSSIWKsJRxoD3Sl2ZJTPAa5wVsXSlPLJlaI2Un/1Xy1BFD1BdnJiRRua
DLrU3+4du0Bl2Y5+ea4o98bvubWjSBNm3+lcedgFpe3fpvNwCl5T05Z2T0LS8/G+
U77JkNd41je64wwwo5MI7jh6mLyy/tUw5VlHEydqZizQjB3Qc/X0IzSNQc/CDxvZ
xIImdCtYSaD1gfCSJd7aJfD08BHONPWVSLg7WJdBgsT0OeAUBD7hfMaSmm6/KDgg
u69KOv0uxOCJ5PP5ycUjmVUPpKsPOmvVau2i2j5lFmBKWanyS+Lu2dGzDZu7v4uQ
bIf3tID/x0WJ831MuhntLzTFI551mC9wTR71V+zWzNm2V92ZhgJr9BIgfJHB3rSG
L5GAU/Uo3dL+JNAvIkcAcKGH9wlmEag1Luigi7hkSH852WC/RP1qkH3Mea3sBibN
tz/gX1cA8O8auQDiBPVf3a26WAcRF6DxuVazPogT+Dthqvqam3OixNXAuSiditYH
k3SYMXDSngwqusPeaYoeISrAiYUf9HNiYU4JUqoynHhnaO3F9wLXQOvl+tj2vySZ
fjddn+Y4u1QGbZkgq3J8jG/dObRNw7ZRUJ+KUVZKkJvIVqQBWQDKuwRrA8Q6AI6p
UkRdY9ZrIY70gyN28QS6E+fUXXRHqgr9pgTPDe2+dpOAVWLr5G1cdsv4R5c2++2D
2sOyg23UA0A8uPxSENDsYt19vXZdTSDeLTjls7VVEuCMri3UqM3n5gklnB6rYQAb
+jPsxYxNk+H/G48q2fdBE6peZHEcWHz9jfRtoNrcJCnIvCoekOHo5jT/+392E9Ob
gNSA6WaFhftLovfavOr199anOxiykkqxvcHrUbEWKkRW02F9pyu7reE2SGUDFQdj
9OzF7YbeS7S3DdmfAWGIIF6AbEMKC8t5+h3Hh2pUdd0rEuFCSZQEmeDPrtr68g+3
KwsAUNMftN3jl4vO0a6Qwh1VJL2Bgfw9tU5qqavTDJI9mNIYJdRS9jhNiLOJ4LrI
5jjWawPvALDdYHBYj7ujRHWJ1FOymnyOxjeN2ktqkeUHn/buHbS5/wiHhHoslhjK
gn871129TJmZSdT0wCU2Tie0Sai1fxL5XwccKvlENRkf7g+uh/kaZIiiMGPG3C0B
bK74sT/cL2Dtby0cr3+vpPM149RbuyQNTRsV0n9/RbRQUJmeU2yYDPyHsMHCAaND
IzBuD3yqPBYz17nGyT6qNV1JZEqTt+2544yfFB2StoRXwQSFDGXZ1r8X9qScKkel
3UFgcAGfS/lrLd050J03D3ZA4kRzeVr9Oi/gKvBSbXEl4+V78irM4AB80i4HrU9G
yyz3ob1MdEZGYKUFyM1RTQRWdqV70RUK/G7G2ImWiuPY/tfizbpeS22jVgga+pXW
wd2BebR9NcAUCSThhlSRZw1ssOJWXhFpkFBNOuATw5+TaBcyfXpa7gc6fYUXS4r1
5zl21rkEHssdNqS98krkrynH0iuD8J6Si0KRptNPpCnzR/iNVT/74EMkqKEXFuAM
JjNA2OwZQAaztBHNayOC3QFaIkQuSRl8aU/9d5pn3pHxl9tDCd1bMICnhpi+SomV
j21sMUp4kvZLfF8mJRD7JrVNQjqT5bKoWyu5U3b04hMvOenl1QFRbuLIJW6VaxPD
61mI8sCQCi/i5JuHX98xMoq1y3MSvxxCb6EYrelk4kIPywCgbn6CFAVt5DI+UmEL
RGG8/eSmjcWFqp821QCpmNqQoPSZLTgm2km/NIYqXluUMECjZi9/yqNa8K5gMLLE
DHvPwgAnfaZRCPZVTmP4ZI4xc/PH6UWweS05sN7o75BcVrg4mtxpj+PNprQa+GX+
EQwhnqOYSZwqYxs6k9iQaZXkptinVQjyTKr4xF9rJlpbSfOax79gzuuNVV0kyXm9
C3FvgpBe62Q4ObBcqkAOkOrqwQ87qCHCpPodzEq6pq9wFafA0OfjT+kQsvy3sDKS
z2OSz4lmW2QmX7BM7VXqTbsy4I1dTahm62Oz1rUJMi6/KVKgx/vNrpZQ0nOa/gJc
6ky7rWDX2HPrB6y9zSRD0Mvyq9qP7KpcKim176+2eL81VmsEiJIf2KU22sEzulNz
t6Y4gKjOhaTlsHxvuEfh5TZylONF+F17eVJXaiMwLkqEv++ml3Y1smmw8FweJlT8
cBb6HMt6AHJQMmoqKm/P1lgGgC/Ypy5mFjs7g9m9C8N0KRv8gDe/UhIYHlgyTZSh
pHm3i/Z8PS3dJxwUIAaLWoNv29JD+IEVd5YytpWueiX8M8mOr7ZSYq98qHdkXPB4
zQP6wTInu0+Ek1i4XUb9hWRuE6pPTml4BUOL0kqhT/9LDQ61J24v2nTDnGeY1pFy
yEMdALI7frglENGg+KKC4lI394V8diKzSQOPhlYufPsDRnRPPRQ0bLrnOVnmQ09X
0ajX0+tHjPVi5NcIDDEF1VqWGFgEFv9dDqPkO5P3FSfevkLVrVcS3e8sk3V7AnGM
+Z4ook9klFRaH0HJaCUxya2OJIPrE4cALkCfDP6oCamTiZXOCrbanJoGkS8Si1Ub
VTcMLhr3GwuzNFJU0v8WMlZzNTzSgYxv3k9F5wqsenGKSL/snjUxaNb5OAhIx6rW
Aa2zX5wGZgzb9RHIz/fLa1PRfFGLAcgF1HOGx30z9MKNAO95nSWYswOhf49s5mTg
o82rSlWosbNWWDaIy3mFDeoFEj2URFOHb1Oh2sH7McU3cuGn+80hV8PsPDuLjRvh
nvfDWYFWcwc9DdqH/+YVjaMWibr8XoW19/7C/1XVt8ieMh5lM1HCBYD1tgn9XESB
5m3ZJ7dBjsrcz7dtc7DYuiUOJlkMfZZacJASVJT96pW0wIPTVtxCGW6rCG/HE4nb
ct/qLEtjb+KnBJ4dQK1bVGS6n63u1cm3o0U4R+W7eDpAK0WbWLWoPrTH+Dcbboia
vSuVh9YhPdt7SnBAGIHe9YDMbqUzIlUO7V8NBHPZTzjg0DpggNDqLil61ionNsIP
KWocozYjoVXq1NWUPomf4SL8VI6vNjhY2s2YbLUlg6rz+t3ScEBqLNODxaagydpV
Y4vmU/2t0J4cPupw34v7jBM/opOpOtaDeETcDypjbP/w7VvaVmRLyNhswxmicCVf
grIVrqeJs39tYfMihlXBM5Vqo9US2VwDPc14mg2NwU0Fe+pVjEZjXsGrGAsbasmT
2vo/h2EiEFSYGY1WsIET5SsAC340BvZTCd9FwS/fXb1zcbYBlxbh+MWdu6ajZQRq
RRXcSgV7o9FSp1Gn8CAdvHp6XyzKjX4CeVynTp7pFWdloaI2j4LRBStO01PkuRUR
Mi+3MjI3G2i0Yn9f1jMiMKTNpCrRd4r54Cbm1MdfRwsHz2yntxujmINu3behRkLn
wXws4zWypL1Zrki4l8tnSjLAqx6E1MdGInu4mKF6WgtxhLlUiwjqxe8R1kIHs36a
k5pXWy0DHR+opuKiowAfstgYWgHeycYE777MozOtvp9H3JXQlLbcddTP2s3ezUs3
xgjNsidr/iJ/+s1kn6fXxzNRThEhjhEn6/nYDpPRJV/MXQU6unQFNJ/A1XADjSGK
a2hPuc6MM0gMMfvf+mAhLeKDKaxzLhNMK2F9IuILtdVEc93BjqbFzzJ3NOKMA2hk
TE/X4grIlTQpG0gJ0+rNaQRZ2SSrtCcHDjLLnjJ/vXJhz5QNNOi9spVgHLdcH1Hm
23YBT5lla0Ae183ElZvI+pa+pAlJ35YbyDTQbZQA5uyxRCyOgwHO+TivN2t868FO
SGFt6cGd+xBRUPxfg35TxyApQ2fFteTW/bXZs508ycld2Ty5DmRpIGHKV1lIe+gz
DwHuxXhjUxLKrb3PhuCGuo+2j1ryrnKfp27JES66j+qceaWDi3zjtGoj9N54KooH
8H3r875ppiyGMfTO48rJfZjFCpKFXpwUdaoA5uamG5inimgZ6ZERP8o90a/JyOtP
jqfPRTOOi2FKeU1V0kYn+3sIY4TwZRwBjnpTTgvoYbMu44OQYm6XHAKxVl7A2oIi
UKpSyHMEr0LRW8v5glKQXUDG7+28+THmbbUojIKvHB1BpAqVfuIohWO6CSYmsYyS
RGFGgD/8jU9bbsIhPI2VnAwlACABgUEPFxcD0ggm2bXd1+SrbNrcwt3vlk2+UF4+
xP+9Xcj0fBkjPycdPaJw/E+RmQBeCYEFKUE66Mgm87K47feivUUruayfsBO4Tlr7
3+6VSOXY8UGwegPXY940LwwrCVq+/YUYcF2zDOBGkfG/B2vD+J+BGoNkYOvKryWi
AVFIJ5mHDIH/lTYkMXini/7RLAChnSVdKjoXoxlDlwfzOgf7hRRldnhoaG13pYHf
K/NzaXyuyqFkagYI9YbyANJe7cWedtduOcqdcegRsa6H71GBwUBY/BtM2d8DFTE1
YoAbjB11fh6LyhZw2BELi3i2yRPopZFa6hHUQj43Za1l6FGDgCh348Fh1qLzwbrd
MyTLZg1R/wGByMPCUHNLqm474xqkahI28oDuSYr7v/HaOXnMTkL9f5XSaTaRWKH6
bcabXk8zbbeIbjZ+KgcNMUZz/9eDioGwWoZQJ1uGT8xWbd5+um90R5JPghrr9wSs
rWeczbMS44PU9+lKShfLs+Ibyoe1bYHunmA7gLZNyB+JKeFHorINiYQuos3b/rYp
eZbWpkWZxWRZ/IxXs4BRfhWLrV2pTGO176RGQ5OAz4qCOmRhG6OI6Ndw7d+WkAxu
0j134rSgbbg4XH/gb0QX5LWqAMCzbNZijDXvv7INBzUAasTj4I95FC2p3O115OQ6
zwNIZv2cCbqghBs3GnVzMgtnvXS0KjqUrMfWV515f1jkQXdlMY9K4J52qqUKFxYV
HueeiUQe2yr5J0GcUrioSTfJXtIzLofvmr3pkzUmJayZy4p6J0OQg3vqzbVxH9So
TxafirQCVezf5ufVbHXWHcqn4ULXc387FNQBT+g/RpxzfENG+O8+CAxaMAiBcdTF
MwKVuvtc8+AkB1B1XwnA7h0j3ETfJmS2eIj0yVg3ECBnpvau/8GxipOQQnZUPYJW
oARYbgr+KJBNIBZlh8yK0pkxOwagHf0Zxsa0aFcz6AFkqRpvZ3ze8H+UE+h3UlzL
rXVG0rOLBgUJQycWJY9JyZb66pGEtbT7p6vNSI0PDwWDtJteKLW0wNfpmWAmFDb0
CNv6mHxE44ftxZC0DQJfpBBYtLEQ7mgVdYIZN6RKJeXN95spqKbgzh8AFY+bm4hv
XnEdfwgpcMH28TPwIFVonf6nNM9FQYsRjr3xOu7L8bzj7bsA+crlRo6FODk7G3Xt
ypj/42Dt7NWYUEQI3Sb1OYEh+Q0uVOvel4t5BpPrr5mFTZi9tt029+bkVJ3P38vY
wVFoMqFZznEWzD6sjMr/Y0xq7rSHfAP5BVu26uJcP9k6U1bhG81kvC1zEUOdoKAc
N4jTSAA0vG3JdFEMH+LnkxIv9xXUgXh0U1fmWARl3rzC5BWj/GiP6/mC6VfkTBjG
O6sIMHTAjwhh68H54LlQe26LSjE5soQaS85KMA7u11StbthvCJ8Z854wUGpVdOoY
LTHTLPeZrH453lNCK5g5S8jYYluCGN1tV4KWCKe/KY2QU9AjjU0pBN+LC3IaaqJ+
RfAm98z32UdT6pI7x1p51Jzgf/KxzB+/kNsUL1qMSUgwVnPSZ9m4n0GMO3281ZbE
5cTd0m/TjG2+Rq2soJuls0RDbpud7GmsRhZVSCGsQx4xkeeLAOHGnShcPglnefl7
XVnnbo0Kp/g7KDDFThTxiiE+A1YPio3y6s7E6dZ3QpD+nwVt0EJr6X3nt19+Z1Dl
9KKp+ZLYmSc0F15HcHck1AWaQv3WjO/LWQT+wu1Grrs3NmcVtbaElMFdhOYiTnke
1sGMrRVOthuvSnhUC4jIPl/GF6VU++y0we+1YE+QrPwNoKaR8F19SrUW3/YvfR37
RVnENtDKKtcCd4AN+b1nVLEDaUhIhIJAUGZ1iJbd4ZYIABCgpEi9iJ/aUH1F+ycZ
koVEEMGcol/PsTsNk0CBB3rlrYiu6zmhcNt0b7E0oPejx8/AmHDCYgyGBmYWTqsI
zTefHDi+HKzp4oNdIfmWxUkqDd9tj978xSRiuKSAb8WOhRe1Wh22RalETPEIwRG+
bVX9l82b8eQdBo1X3sGXgFycjiww5cjen2KZLHWbsdz+BP0/ID8qXGFMs2mXh0wz
+0lzEF2NtuGyzFg+YjPDhnnwI9tzQwEHOjWARzevozBUHVgikZ/JrI3BXU7EJF7O
Yh9JqZ9uFn9RSnPwHeF/FP1Av5Cn5TJRUVogBjRlFE5L5ELdgdbRLuaSS6nurO3+
t9Fz5sikFonHJ4PGiHTe79GniTJReKjI7qX9lPLiimHBtnMUmGdBbroxAp/wBdxC
cI7kw2Aa9cbZV3NS9BwR4htaU/lJlh6yrydBkB0tHpp93ySOveshLLMfLLPVhE9u
1EWAv1W+huqs+ylZCjoeT/KxmaQ5AmntaMKxgk2LCkMTWWar2Fw8lAmPnwQnfG54
ZuBCbl+YnQs1KT+AuqK24yLC/DdhIiBQtd5X+jdE0TBS2JlDjTkJiokYabUbbHlx
1rkn5w9u6umVp3lvnJJ2nvZkmeNo5cym0OpIrhp2LOOC/B//NceWXXvskk8/stlF
K+x3egyqDda31rnmjTi1sX0u/ntkU0viKa//cczcNeIWagbIIOHJxEM6mBqP3tWr
YhMf3FufoTQ+wEupkG9nXJg9lz9IgKWQpkxP6Yin1NHu+DmISNNRQIOMxVu2eyj8
+ugEfUsv1Tkti8lDShPhLMZTRP/uNwvqBgl5E1A++5OgicQ09ymAxTAq2B5WeOhr
ILqYYGbVmbpTJBNyNiIBnxV5lr4lij5si9ffKmieN0Pm9b/ishlK+ujxmWoYshOx
LuHmgefl0EttASWrRJXy1C3H8m4z2lNYwMLZ+dj/tuR/9iTnaBT1nyPXYNNoFztd
KszED0T6/dHkq9FECnzIMtX/LeSjJ4wujm5izx1hbySEZ6p/lbrAnsOECjt66t2X
SYUKU7tZVPzFC2ukagOEjbho3scqA66BCc4+nqrUuUlVmhogK0+VqZpVX7Qq2WbG
31qrh9gU29FQQSF0MH13ebejpOX19gLZ6ma8P3CIEx9HrCyAof4oWN3mNb/Zc9nb
Nl23FBXCyBhs06JbTIVjbzMzlip1j6/mrBLt5WVAsQYvoBFG7Pf1W6vl7QkiLijj
sjrPVa2QsrodcqvVoYP8bPixsjlV5+DKB3Gtm3ky8QKLP0u/OoeP/62htvarWp1M
FpeNZjs2XwKeCWt3vxNltohrKsoKsOOe+HnbHWyoJ6occAsTrSM7mP8LiHKVEMlj
RyivQCunmoAaP/OqDyywnJcnmyHmjtWx/kQOnpV9mo5D3yLtN9IEjWVXCrqZK6o9
v8N0yNzc7WWxxKU0qi8mk7qBAx+SGqxp7p0Z1bZC8wuH/tuzK3TWhyj/gBEbwYV9
3OsxqyCAZn0a7TTjdisVzmbncWAmkhUmW+ORzbqwFUwaETtNSb/btkVXxBF4oL0H
U93RTfmSS2CMJlpBUZ9Qe6RcN82A5HkFTCSHmLYpz8dQceAcAtzlpVlXNpnJgPsn
JueUDZCZoNKM+BnrzLrtVco+H+AJ2djEe8iMjaeuXM0JQFBXHl9Nspi1DiBnPKMd
yvB6aQDn3FHeVl8rwvsgng5WSQy5NO0EeMbrsvzFeYUMG+SX2QoqLBr5znL4vWaT
bZegSiMqxHMQzd5bNNkqzfGuwp8ep/qvsqmCHoU08xhpdPTJz+pCg37S6vupfjFV
xFjb5WZMj49crm3jZtVTIpp2JYVpcNVF7DLE2EVEdw8xZHHeMp7tE3qM9b8syPLd
jvdXWe5ZkRaLUwacojsbr037vNvZTio9Gi2pJ1d9E2BBHxCHoM224vRzcieF4X5O
lLJ54joJ+oVD50Ibi7COL3bQj+ZubRuGQcERY5xGDNv3jGTYjwvnIOitMQVdCWQW
w4765IYCy4BC3htVbidE8+6VGLLiGdf8M1evRliCmS/9ghY69RLYG7ADWuDvnAzM
U8iFB+9YRAmOelZ2eyvUn3x6MnfPuKaS/YARsAah2Ud28EYyPVjNK7CnU7RESXlq
q6OgmaDg/g81ziLIGDOKfeaEme1P8EHPdrZCF499mY+LfculLsLLG54xkXbA860Q
l0Vp9eCffjyqtEiw/nnqKQBRmHejCEfPQE51Q5WAHvETVQVhojhuEyYEhgUGvTS0
20CRLVgJX9dukpIFdEevgQZFCGLG6XU27MWy0LSX4OUYS3hDIzmkYg1A4tSLlI8n
tjaabElOv05MYOD81TMv/f7F9Wp0Wm41a494tO/BOcIIZxSbBowYB3cdEK5BDvHf
IeQy7KlM+l/79hHuAhlWJ2thUyzGna7FQZmvsGUlz9TUUaZ3rcUodCBs8br30LAo
sNgb8T9AGFPQVhBx1ghftwvZU30LmPpNSOJCCye48b51V5qr2w/fQFCr6YJQG9RQ
UX9sE+VQaMxdhXBEwJLplEiKQLmE0CUpo9pfGeBRgOr8wtTvTMgzag+dGxGRTyU6
7ReiEuJYAbkwHItNf9/sIKrXAgBQjrqdndP6a5F+Ma3EJlqxQNVVhQHXSvcwVAUp
7NOoWDahzNuSswWj1hMc0V7pGL7Csla4S7wNmZQO7zsMogH0+mhwu1xGi/rk+Wnt
bB8CzWLlmEeDfIkz7+u7NQs5v9fTDYAMTHC8AcymIvCM88Q6nCda5rKBiZEC9TVs
/DQP8tlROx/wcNOZgxfoL8DF8k+3I4lrOSuzKtEDWDc3vJ7x1zDh7iqv8K1GWJTo
MiWd+4Gtf2kGNA47VX19gOnYnvR0Ath1Wb/JAQhpFNifgbtFXZbIqJQOCfzTuJ5r
L6Zy0If0OzViXQn1aY1Ov5KjKJ2gj/Z9IT5MUrkIkC7pJYSF9BJajTzK6sCC6Fdr
muYiJ+7xs1xB+xpFit0zFRKj7aYgO77f2AL/TjwqYaAqcz6qH1RIa5JdE/8C5E/3
Lm/TdTYgwXNwSbNXpF6v6cfZjnTXAjrubrBoMrvtCSFVsYA7xBoDJSRoCEo48c+H
f/RIAAZa73KhoUKyciXhD0cXyhVQDyn5Giz6rA5198bIUwlb+PQ7wymrAS6OpMKo
9/UyR+Th0DRCQLMuGJBNlILxPX84f0gVvmcFxYURXGSQc5y274lZd7Ls4nDYxO1/
z3UoLruNRxIj3/rWjK16GvrZJZqgp8MbGpjgkITDAtVbJsvMB/ywkbU1j47wcNeD
4K0ZyahSrZLcyxBp/f/vOGoliT6x9pN62DpK0DfrpqXUd3hNF9+UOODyCAUZ4c9V
uY6hF9TyivVKL4jTUtWUpg1cRFy7C4dJfIPrVONR2NTiN25rzWFGEfN9AIJmtlIk
1f6QYffJkSMrK0bVWdfEyl5zkJNU2t2dXIXHALnQZY08YB+KktDP32RZCG8NAVpq
ftnsARgGnLDSO8rylIWo/zWrdZ4x4b3p7UFBfpOAjJc4J17NTVjKUlYZkXiJC87l
apuJJzRnCO61RpAt9RJVvun3IfzHaVIc5+aDvG3Ay5SlNWvgFCgK8ZQwMKci/hY0
+lxuSfb/2EooMthCdVZyeZhSA/YmeaLqtJ+6Wr4SjROzcaSA7h2a5y6zKWZ94o2w
Fe2Vaquf5mGmbWCPsWrj07RwD8//M72lWJuCwRTuSHgzBn0zOeaPVUvbC8GaYp0y
4fA9NcYY1wcfaUP4+/E3CjWGMhjH4tv+AzXuO7P8ZkFjoYphBhRSlb7scqEaL9lo
gZlL0JgaprJpZSyGfvndMRWIZggMUk0Z5mr9OuCxUY5QWzV2Lj+a7mFfx9OtIBgw
VmtZnAS/5Ntn4uZ+nCne+xmBwYzY6h/x0MJ73dfuF1KNtABedZk9fzTwX91H7kG9
zMM+nAHGp3vKD4lVXsW9ihrpA9KspNxMAwJANzvM0i5349raPXdnVweVt9PxDaYS
fFs+YQjM1yjeZpsMmfNGj/uEmdNukAj0B2SZDnBsw8XXRKQgyU14tMLGHQzQF/W9
huxRf4Bo3JOxeh7A4DMV5+xSU5iobL7uhMnsA85vuswDBIFkOOzjJfqdq44q/ku+
zhZO3m5uWwTVDOWkLQDaiQg+NSEqW1Ux3pvswUnarjGs9wV0atfRhvRUaa3Jmx/6
pzc0oG0sN+1wOshY3nW9ub7XEKUTGHCBCdHXRNxlQ9VQjMkQ6SvrdJmsTFA2F4Gt
WZoB/vekdPzrbkrgOMwIOrps9k/MDvI6D2z7l0yhh84oXc4U2iFrKd/+/pCWfupP
mB1XsSvOcEV02Z40SaDxwXfwIu7d3xKqGNxu+/moQ7V0IHl3QLcDuMSPeC03ncxT
R6TE5CJ1Im8N6If1pL0dk6V6NuMBsAed1/A/ZxjS4P8GzDm2HDnMrCpbyqcyI2aO
vPyYIy3UkHZS9lWPbIM/vaWcfcmEq5bEsLYvkcNjCTo7/AOyvon7X5asNKmvBerY
f0b+Ux6pjAplfe5qETCMJFRPU1GV9A5ej61VKIxf+uU1j6sVyoJu4enSyKB2rTBb
iWvGXPx9uZ7jhOqrqg5O5ZXR112blSjAJrzyKqd9UKqTEO6ZdVUINplgt1EVx7K5
gLERDzvt+04ClhBf/08j7ERjkxC/QYOVTHc2KaDw0iKQSiLYXbaT5DGhtrkNSZIH
ciVvXiY82LRcoPLaD+H3UL+DI4RcQ3VPq157iwPNA+OOXguV9Pd6jdF22WlRbmoL
pVV59QOdNA8EGMtXL8i629L0dogAvvfWTACpjOwXyd0bJDMgcVRKR3kkL8z1MUIC
8TFW6R5vsehbwOCZDKsWA8sEajckiM1vqDnFeURZBiMqM0qxCr35Ajc1dCOGHbvb
3sDS3HbakBactanZ7FO/lYPvSwuG8tpdoNPPbqrskPTj3z25HFMjE0pRP0pAIxeR
FTwNiXcENwRPheF8RR1p9LDTds5lIq3gd4AN4cdC7gUKkpNAZakgxPU7FQho/x+w
0wFnFFppGnF4y4hVax5o8oQcjf0d4G4WozfxIMHFkUxbg4m/RuG28tjW0l1vNs8/
a3MWG746ZjgDUoKNZJczfW7JpYHiziw3ZMX3rcRV/ULFf+bCdqI5Mi747yD5eSJ9
+WWKq2s9bAIoNJbK7KBLMYXR+bl7PRd/GXR9gBDgoNVFUcII5evGgcort9Gcg49G
zLX5VNWhL8y4PVUAlUxorFd5/fnP2atDY5F7Tyblhv1FJz10hW4Vy6G2EmCTsBEp
Dp2suwUQwE9thYZFrPhUASq4L/Gc9MvRi9zuRn6X7kavwjFJ3mAFpyCCoqb/Xbtb
Is3UW1KTbqn5FikQ3kwWdax6l2t1hfR+dj2+6hJGQtzxwWuIM4k8nFotF6BwNU6q
wjqWa8Gmss57d7sI9AyIwDPQqvkCkVOzFHHVydKYYoDEfCHk12MJ/po4TEd5Knce
rCu2dvwIZ38teT6aOCxT86bRylnR+XyB4IiX/gz3f1SgGl1B7hvHc444ztkQE0LX
xWzkY8XaOfj/5fiE88krHkvSWq2yqa6UYwB/5b5N/6DLerX2fkjv3xSJjM3Fe8Eq
5oFrloiFaZQYhQEVOsY5D7/4o3bmnqgoxaN71Hk8dXSFSHK+tnuU/hdkH3xLC9nr
LeziFnqtgG4EWhuHQInBajbRjVOA10Bi9oiEhuilO3xltOoJqAWmqg3/Qvyoz05R
eCkRZPWhWWk1f1uzDEu5tyRp0c3MUM7dP9/XmMfFMWfVXYxdVWoSVGBwQUHh97lC
msnx9/xEzOo4XoD9OjhnEYUtdSgv6F2RtQRWPCf7D2QC9Nc690pDGu98fGlDyRWl
XaT1Q7nV+pmPi9eaInJMkMV34QO72msMTuTLFTIWKbOcEsrb8yLDy8Q8fbysKkeS
qbUWpO7JqnhKJfaqLRzg9vBEdKK28uqTJs6sQMtt0SC0jVg7TjfHbC0vtxuZcJrw
Lr757qGM2aOGH/ALLhZebtHy9tAGlxl0WC8y2uRqeIFHE6pOGTHlRaQP41/x166q
5nL1Ug9aF9sjhyiZgBu1ZRr30jouvmW03/jsTcot6f2oPSqh/pKwlkAeUXDl5rzf
F/fYgPX7Oa95Gqq6t/lwX6zU3Nk0brahmEyyawTYHmKftzOkc7iRanIkUc72jdsR
md1rqJxVKjo7JnMdFq9JHH6KsvLQSSYDLYDu2ATX1q1NX/zax2bI73BBcvioCARd
JhnG8L/vHLqTixK4vV+m4EB0dOWwU2dfZvQ0AdiBZEvTR14bqMBc4HIUf1H68bVN
ZNWoeUPpoUM/QjQfEcTskWtUv/fUtcyklA5VKMgBm/RStqD+/CbJ+k5PBiuEt6pL
1oyfWJ423q2k/2w9wNCZG+3ufdluMwsOfcScsIVvvXquNQ5BZE1E7NzxQwcZdQJD
9L+YK7ySUJZPwrIQFzqN+M58rSSZVAuHDZkWjfFV/2x6Ujg/1aO88LJU5dh5nvvR
ecwV51jypDJ/44PUeDy14K6lkwNw7EN0nkoS2dOEetzmQaFP9zNozMCOMbwt3AJZ
X26fSOIgfbqBroN4EW82gmqkZlAbFQJxrXaqMrAX5hKUxTwaqw4zMAj8cvt/haBj
p4JO7eBa8Cstt4IWBmPHfGuiTx8xOwuLYwgAMJ2mdCdm1NEJkKhlK6UOiZqSxnHy
iX3Y8VNoz76I7IapdR71DX0V8Sy6SAkaWRP6GO+jRZlYyD6XnK5JCr6mDrTcOiI+
hPlDR6UIWAuxB74iy+N43dy5QhcwqFg7q2v2bO6gWdZSfew177IFGfpDayBkgii+
bga8Jiku07dOuGNWKpdhOCWSRVdjOEdFGkYyCmgPNohDekdc5GWH32TXzIVPG0/t
CR6Q4ABi8h3hyafvvPVUiPG6CrMYsRcsp3uFzV8kCvVbZdNGjKeT2qVwBGeSIAvo
31Uqe3sUx8vNBzXF5OjkNG9WM9q4tJ/2oy/Duu4AAisqj7tSjE17Is0g9sGGufvO
HlvmpB3KtRaNf9IyGJgxbwMSAj+p07Rj4Sjc0YG0CX8Qz6vpUF96zO4VZdXVoWY1
PPQ/DyQTrcAvYpgnjOZZcKiyu6/SKHaCkC7TK5eBH31//61Y657FSqOvEfL2vLWz
1pg/d60OVj7aZfkv4XBZtKGJxDNMabT45jnC1mFXoykGREH2FqONWChrKcURFx0J
EBfWrqf2IoGCZOkX/Ss7wLpGuoaA/PQE384XXiqKh6zHtkIFxe9SC6wyyUc6LfA/
EAk2x7MgEeeTzgBKHrGQXyl1/1Y2E6SptpWa/j9T9umHGDG4n60ArTVw/Tifckeh
g7FrsfRSaOF1aKYfHkoesukrjvZg4Yb/pqEhnWU48jmiBj9gz0Y7wYgcljrN6DM2
soMkIHege3m9HevOUzDCTZkklrvSK/i2QAdJ8QtnJ/UXvCiRU0Wyfm7DRJV3Z8Wr
Jp4P+U0NRFt71+1A/3RhiAnc/NJNdg7KvOWzG5CYsYqxy77CUhpc5Zue7JK/3AZD
zbNOpNwvaxWKy4hMZNzRgmK2Vi3cBvfa7FQhAXLXT/eRxMrY+WWUJ0V3svhXeISp
yJStrZQWggKXHQ+fPYdkL9Ry26172ZSnqTB6nOnIRTAjCY8RbWv3pNruLOtW6Uzk
HKknlLxmDOX38kc6kJiZz+1v4gX2D6OP/CfKISuLJb70uupX0qj6MxB+mVjTEMFF
e3gR2K09mzTx+xVKTS/kG24oy7TtdIqKp1rzm/HqDI3R/4hQVMTzDOZRCVxdBQ4n
q1IkCB5MtuGZs+aXV/hay162mq7xhMbHXyKzTxzf6qSRP9S3qOee5GfBByQ9LH8h
X1SjGHLkS+Hqb6FsX29IVzOq0811R+0ItfLdWk7f3N+Rhx01cCwg7a//B2fbFPsJ
TaGfyGcxCeDCLSHJa77+3O65XE6STzQ6qC34hcVUPrH3z+3bimavA6kW9rb5RTpH
rnnfQS8LUbba+9BQn9iT1wtZnoDAqKd2TxZYPDgWJm3tmkbTjrKUn/QSeTELGoqw
UR5oiX+0bOujf8HrY2nuEhp7vckB5vRHL0pJr23A1MwnJcLiZtPvf/pU8B0aFqxC
jRar7Nw7euV3Hc8Ao1Wben6h2O4IbaY956DdAUEHl2KLyueLbZ8YZhp2b4MPvRc8
Lt+5EPpf0quHcuYuxOJUmlCt08PoVD3JfqLQJtprRcICPz++Ngyd16i0ICM2lpaY
Ke142/gBMqK0hze4I1qKI/QaUOF8qzwSYU8om3E3XWfnY4Fo30nR859LeXxUn11D
SUw7s8RhmEBvy3He8ZRXEsjP59+X1xnHUm3u97HMnRzhFXls2WkFI0q7MpsfQj0K
mwqgEqOto/5/cPatffHt65WitEqZ0Rs/c+OariLujZrBhu4r/JUxryiUBxXBBbPa
OS4DiKzuWYG9jGx6xi0osOwk5Hd2GvaOYOUSm7dEhYV5H/rDCV7isBycYiNy9VvW
c91hu09Derx6MiOdO0wY2RcUIOGBNqWjWOIFQ8Bau60HawQ9IxD3WhNvjTmzQTSL
iAXc5yHYV4h90VdigUMDNf0KKkQlj8PUe/7za6k+eNzQ4XjUnA1akPWAnQ2RApNZ
Q79P1QSXHGZZrbuiZgPxznQO307XmXRlZ0Pntwp4Ifbz3D7xs7FsfiVPG6WTAyVq
4zLYjgDKRFk5qujoFuhu09MeyxklsYXsuUZS2SWLbIsNSzY9th4BxaIjtfTLHcIV
sX58SptTc64UHEO7gxJoeYXoGTP03ffVxTRYUa99eMzrtjT5jGUTpwI2mFYjpAXa
ZDTZofnINmOPakScrbjHpy4EeE22fS0A+I2NEvntr2PQG3g0JRkDF5WokDgSQM9X
KYq61f9vGw/y79e2fp831Hu3f4P+WvxcmYN0Wc+TcpWx2zoHGjeiHet5fVomrPqc
NcmWVF9BsbpGKirSQI0ZsYNDeTM2PxwORBd5f9Opv8HRMSmyMT8FzjJNqwt114s1
kvPfqz1FoW/PyOe1UpdycVibeLeuxBazNJJkPIml4onJDI+LPGgarUEhiFx/WFBg
89zFfMxUsj67oiV3yckbX19Laz3LjP93dkfa3ElQZdxjahmO3GPJpwrFcooQIhfJ
Oo5QY/5H5PaXNEOGD1/2rVvXkGUQFSr3WKM1mB2hkmU7+Amzs0W/JBUpvCDv6D/u
l9HropRIfIYDOgSwvh1fS+miMBTlvkaoZQ98VcNmGUImC3WZ85DIMbOljPaCvwUl
A8oI7KpLLRTBeLIzSLPoZghc7ALE68AVOq3dyM/z0MxHli4THWNxgLGiRy4ZFLRK
fhhtqN4eifW7wgFMgLGo4ocUAZuAYXpvjQRwM/yfXTBj91YgwLGTPOnHpSgoSEnc
GesYHjJIWBvVD6kcK93oNXiwT6RJys3w1PCJv5A0AQIaxw8EmzxnFe012HUJ8w/+
eTZBp8Uv1jKvolp/BTkGvEk0xAkIqNdPTePPJNzYF7W74RVMiTRfZZeIze9+t3mw
9ui/ZAh6LlR02xbeE/MQrSk5NUOxj6ji9tbexke316ZEF/Q/vX+SG5QWqa61igEE
URGoCWnMeq3ww4xIb6K3vSB9I2CRZUNreGomjAgs72xm13C6U5NtDHnTlVGMNvKb
RUYAQLURdvsnEivILsbv1IQC3bHhRCYBgtZ57QbPcr7n+1fr4ZsWKKLVw2A/5fcV
22Y5P2HRuzRUorpZ2L9fNWehK4C+atnemD9rebhYH6gk+tbwmE3+dtMTi5402JC/
r8weN59ofE+ER/+nTZETcib8D+706iuccL0pK9gTxq8HvO3IXlMKPM/RgSFjUw4k
JnQ79cmgfuA2faJF78L4M5s9QeYQODENvYK8xcHdWgYSQ4XRGw7zIETkmi17Irfc
iYs5k8ncYCTDps9tFzrVfIJWe1x0EE9+j9wqFNhmyToC4U68m4bUAF7+ErFPAVdL
HA94a662+NZbIF6J5UmLbaGDJx4J7da3f0VTrjqc2IYqs+QftDXYee5yFZ7Vdw0l
h0f9bHYINuu8hULRsqiCbMeuUnZeRWrgmlUx6Ok/5hTjgnrsCX+lCbTvim2fRRCS
v4pqIgaj6957Z2TkMoywJGDSbw53dpJqLv3ZAbKxWIzilg+tgLAvx7MjePwk68js
YQHEzxsM6rQHExVA7Q47NFH2RyLRfwgizbXOnfzP2p5kOrl0T4usuGXt08wSr7wo
aD/MUmHujrGlk4JWNRObMkW8ei19cFP0pf7n0alh2tMhiHZn5SUPAqxlycOjD6uM
zQfxuXGgjouUzvuFXx8kEZh5k7QQw+DWVDSWjfQVaC7FbGyGcmX+orYqy2YQC9gb
xzoG5D/m5l1O71w1pqJ5iGf+1H3342znbkMo/hC0QYMrzSQS+z2/+/JyiaDnJlmk
KPoKYM4pSB1c4rIIaV+cSvx9BtAe1wdVoeVX2OFyF+NoPe4ClD56FjBdHDjXLeos
DNTzzy6opG4rcYCEMAB9vfExMbeDGKMcLN1H87T046maNfpE4r1Jrcr9PhioiW8F
5d1/HWAG+JwQLmPAIxssb/ui12dHp4OLbR6dmPMQ8vIu2Bjin9K4mQPuYATDkeNo
FIg73iDINoU+I0TesfnfFqBr4+8EzTjH/erCt3gnKCjZyJ8my8SKJgQ45JKVYlPk
JOrDO/I6gIYDx57EK/Ct9U4RjyjQcPpDu+9m9t44ZPYRpjpIqDvCWvGdkKqYUP6b
DtavbX4WwC1OQKlmjx+UMLL1BpL2+beBYH+1Fm5lVQ85iDBddnuXrgl2ozA0XZES
tqn7YxHlvd5JQq/UaUg+PejpaGzp+MSSzT7bwqgMCUazAsTA0cx2GWLniVoXmcwd
C1gZ0cy+jZVcxF2E6JV0t3KF7GNllMqy1Q4gx97x0LteB6r+7mZ1g/Lkg/18oYgm
gpGuWERyBgeML1F6ZQzHOpHWzUdExhb0RscknRcOfWrMl++4KhhIiIdJ+TMqd8uE
N8HHyRa0lAeMreFKTii6kI/VKWpzVLlk8Vqx4omAuVLqiUpZxVJ3RQaR0gBRrj4Q
gxU8I1gOCWizAj5Thhs5gbpqvEenJuVitcarMdOODIvNrNyQr8ExNldw50xnQ+ap
Vc+4r3WbD3MoNakDhZfMJQyLr+ZS0TfOdMxxjDQJBnXnpZcibPlxq1zT9Qr3jBQx
4gpWCQyHP8nZ3c/r8jeC7DDq7zqgWQPN/Mn04scOOcQqIVJ55916T4pHekoNqqgx
3cGTEkgmsj5R8ZqtYIQXuB1F7vZc+1ZYn0jeI5ANZl+0p/Nf9wP+bs0q1g6ELbfj
Ndv8IjK/GT8DUD4RNWJXRthO1JUkZ9FQBRmgysp5DZGH2VybxyyG/rxFos8NPIDs
HjHzfxXtbDe09Fiq26sfNLtwduq7XtUlhhsTtwoO/oUlCwrNIKFr2CCkgt575pDA
7J8UsJ/zXNixMwcjfMUAqTINV4eDqEiYlLesMRl5T23U1oZAYVHLLtjMgiZUG8yj
QSdJKe5pFDAsfoIBYsLwZhiBr4ObIST9O2XBPXkY2Zo/sxexF85jpje1UAEZDJxQ
tR14yHeRbXIMqu6VZGaB+0Q9Vt0LySXhgB6FtjtRnCJhE9nL/epxUQZjSxeAzZe0
sgAVPX74Mc5lMYeThSnWG99B/toWNpEmGfoR0/yjKhcvNqOGQU64Xw/FkSAPMr9U
5Fo+wX4KzjZ+vX0GKAvpTeIm6lQy27iJFKKwfGDQoPrGeLk3ag3+OESFAlVuYkx4
X+/5OOZF16OQtZqY3+9mzYyqvMQhIrc9AS0NG0bBg7h8se/T5lAjf7xtBYvvirxP
G0i5W8V8kG20t7bJZIFqizjWuD9ZB7qi17mJNCx8boMNW/4RGg+g90flWmpAus5K
3QWF/ZSd4D5AsSxTChs1a2/zA+QDkUV6Ng/9I/yfywIFB0kaupdh7ejPk+izNsxd
cPSIe45FjAopiz1FSGd6xFCLXf0cM3Gdt6z56aiibTwC4EOe+ROcT1bLJ7cmMeyx
YjfX4TX2YS7M0P1bBmOZT9sBzCRWeETTSinlmvAjyaM1twgWUNUYLoNIEk9UJ+YP
8cc5Vx4qRZXQlQY3gob08VJVbKz37hQmtVugS7wNmaOWXHbjeY1IkTu3nr+rmuVq
b05DJW/uitTYB2Ek4UPLySlGhudcGVQam3p9aqylw4ZaE5qsDa9qo8Tg5lz6q5mH
1SU6ZCxnSVfFOxv9Jhpr9CamnWq4s0VjT9NYw821alJsdTfaynOKzCpNwuEZ3tzQ
74fw+Q/7NbDWhvC8xvv5C2Ylt//ojAfnFHjCKQJM4LjnCAMnKhpWSPFVFrj9/f1L
K5oxZvLg/a9nssmyvHaiKx91iiETvu4hiUqgjdmgmUtV7l9ihdJDlSpfYC4s85d5
2EChu9T21CXp0VbUPR4FSMuJwEpfp46oVoGwX7TE7TWN2SzOQ74T8Uy1kVt8cmL1
Mkb5uCbOb4lvBZLcM9cy2fPNJQgSeWOYjg0uVEUSo1ePTZqQfAkXghLreuXQdD/c
2xQFMFnIHadFGkDBczHgxKNowtBpU6IxKeKOM6H8L1qi6omS8tGfGUJxBtFPSsgm
ejjp9g2zr/aEYhEGaehhphTC0dkMAB+zYLwkLIkUOgX/w95jJl+VfTw8gB7N2jzb
3IhJKtYnAkZFZrCrXPZBbhesGpBLD6eVRiBX/JMlpyMQ6bvcHeJXfIVGTrZb9+Gt
gG+jmB1ZkhK9+mdO4q7emF33+t8sET9mGez/J8H1C63SJviZZOcP67gqgzds84zF
V33AheMfvxtH2BB1wwC5LhI+Su4h9K6dStKcwLSkahiWEQ5SfQmx7rjyMWIBCqX2
Scto/goXoUxxJlh1FANwOAbzN9WWgDwdw62imQHWAdS+mJImh/9bJ0sA1n2Yrs9v
twsRWSUX3kvsbn2i/DekTFIcyt9Y5ThcCbs4U5GDvPz5BoSUY4TghZmmKqwHG7b/
BhtS8QkwokrRnMXGi8Z5p3zd1FDeIgXMvDEPpGm2Jq0ny21fu925Zis3Rc+ACznU
jT7GD7N5ZMqz0pSTIfmfyURw/BJjGpcjfaHfSEaOzqFsfymGUAuWUR7rmGfLNKJ/
CO3++jSSG4EzFah6BgdH+mTAhynsIzzkWAwqDmIdsQ9wT2Hm0cmg7ubqOJf7AF1o
ZKb2PqTrc/u+KvvMPkCaatgpePYi7XYmt3LGL1WXSmiN+R+c+S/M8AwJXZp7Ml6e
AZrCZY4dJexGy6cciPCxMPM+DrmfdBRn7V1vwUe/5fXc6HJg4m6+BesmNOj825a+
GNt5xmN1o8hpoBRROM4Rpo1KRN6GBNTDBhzDioDMIDuR4S1lhy/fxyfkWHqosiXP
GrC5VlcdiioWXFJHIVEbntnkBQ9tkvtUr4HZezE4cAkx3sodxp3Q3CyZi/TV9pvh
fKqU1SXMg2ZiwXNE+Grq2oFAJpA9kPqJgDMgL5ljrzU5+aUImxNfIM2nIYZBaOaA
snLmbzqEZDWAcVtjxc1siYa1zSo203GsE3Xb9KxrSdi/AXFtL0x53IfubwmqH+mY
JTrTDehfEi94s2zfDeMzYgdjadb9eb3+Jy6Vyjeqr8XQwU+F7aRWPvmBoZAKzr03
rsbuDyuMhLD8sCcsnITC8JHfZOYCkjxUWUQLofPfwJTKPEpu0KY2e3ciXuqPyoxg
lPXxgA0hDnBQv9hcyx9RNxcJ3S8BYSmyc8HViYT+XVCiFFa5YlCl/vKQ7r6ayPfp
SQKAmRSxgG+6uzVgrJUq/Yjst4s9q7Y4cHibGH6uF7cu+waJwetL5SJTTo0/h195
gwTGw20pGs8xpr5aF9VOxX53g0Mmdh7+QHq60jtTs2Tzcvin5p+e6S5h1plWEJ1J
p3KrhE7GA2aRFg8mdMVbAi1zVx8Cidem7pqRL50HlrmrH7mzvuuAb1C7e8yy7eD0
NQtgw1wirZT5kS9zuQ0pnIMzOSGAjlzR7NpKyBql8YR1QcdWbM03m+vCK8Furv1u
oxl2bBbGOPmkkvOoYN4dV3/L9A/5srPCTYouZeGq3FFlZF2RfObhfy4VKqPsQNb2
4WsokXf5i8JHwXK47wAUL8Pd6aA+oXqXQ3rCZ2ZJGcpECDPFLBfRpk6axgfuZ7lh
v9Jof+DmGtVe80M5ePv08PCw/SenQNcFu8wW3FevkaDnDIxxB8BUwwosanUzGeRl
fSluJu/R1Koz8EYd1EvdXLB9chBXLLWsp5VxgVEOH5s8Rom0ZIi27jmONRri+QTN
XxpmLa3Re+Xez5THKwBpKfl/EIfjteduLYkvO45z1IO+GpiPKYXClWvitJW4bI6Y
ZiI2nxcCX8u/G55UWXjmLo5RJ8FC9N9jmToKw0SmIqMorGOeHg7COFXjZH3BmtXt
l1fOKzXLbTztXDnJlQ1gdEOxAtkYAM0pvPprZJC6ty1r6OaFqgCTDyKDOcf1yyjk
TeMd2qvkkq+0KDpEv5rmSrtUBoKV6DjsgPmn1rEhjAEN6c7fR221Ws1M9s5dDqjH
da389Q5MsL46yxEg0Sw+tN09sKGsDQtzQs8kN/lxatpeswcKPX+UqaionDPSluUL
pb5FzARR+NI56i1IXUVdWywyGA0Af/IlVuYnAyMo1E0ziHzkmEPHJZk48DzxqpAj
Lx5OzF3JoFaUqECKvsu1AhzI6Y66XIMxxvg2+Lrma0gdpEG6zpsmfCMDw9nLdSUN
i8W61n8VbdKu4tOwl1Gi6NRDC0HOgO1uPf7JrRyEfKCqGztRNZz3RoV/zLJ4bF4E
X4T4lwpGLZX8dmI4KqgsuzzURPjGt1W/PCzWMsZP6PnarI027mlN+x8Uj7MvmETJ
vSGt+VI0iD5ldE+mxA6PQMUAWMIk/k4UCFCfzA6TTOOgJig2xxN/9Oz3gezH7WNo
YDl6pUyEE5g6ZViQAa3CvQ7WvAshzvAuEhstjsVZly/VhCNs1DVgqjReBsdDpauQ
AHWskM9l5AzKf8gIwN+sSs9yY7jwYAb9m18lscmXKsnxItHiQ2magQACnwd6GVjz
jMAa+Vn5mbtLDx0JJ+AgIfkbTNz/geIXe37BApZXY9+MGQMrlTm6r2sQ31DdlW1k
RGzVv38Yj3ykL6IJcorPi/6ipzLatpBIM+UeOui+BguYpEjE7w9baI/qPH6dJi3E
iopTHUMnhFoSxeMlgY7zEzmB1ki9LWtlKZOY3UUtWd/pXTJNYHOQE54z2+2ol2CD
VIRuK/dARQm11S7jAyuqEHKjY+3ISAjlP8ZsNDDflxXUqx/YwbwLE0kfAYUtJxxj
drG2S7IQdRa7iX0wXTmFzuweMUT19Uemm3fQh+8CMzdVZSzsUFiXPM5j1DV602pl
fAu3aaEF5SFkjNj/sMDxY1gqcxUs9B3fX73wNUElQXTX6tqOTCNK+2wRzywjpxfL
52A4hOBeCMTgIzvd9N1druIH0NtaZzuY1S7nUCsZRzaBTtba936egU2DjOJY6YLY
OCrllB+tcgjPkBhgkWFSs3F1Ly39CK7HTT+jfz5bVot9BgPBslf4JDMynzZ6C0O3
vGmdDdqIeHiNvtDjWTGscs+hVtnAyNHct8xHUabzYkFRrq2Guofq17Ddz7oQ+MCt
/vFz+LVSlv4nFLFIKC7eBKzq0J2cae1fMw/sER1doJd+diu8oI/Aurx+tRtvijV+
UpXUobvmVJIELwO5jnosLKv51Vd7Bokae0PwL9QvBhJdMxFOm3zbmBQnxKvReTes
VNF0bBgBt9caTGb4COHlsxiJJC9/F0lJMLe5DVxFPrcKXs8f6EqqWhXXU8YMXBWz
CAe9yue0mdfxvydiNLmk6qFt9IMtKO+8d76bvT5IgdMK5wB4QGzP4X6R47HcDmct
X4nCNerAiYSl+/WWhDehP7CaHtB3D82JlE9f3oUTojNjK0uZUweXAWBM1h1RVci9
6l/TXlfPQRKRC1UXr+wBFi9mqIp1yAqSQ0QBK/EaX3PR5Id+9nBZy4ED71YMGP1h
iOZuDuRqeebMF/xuJ7ZuUxM+JIkIZrCA6Hq+r0/9HNtqs5enXOaeUn+dt2iEqTGb
3yt+wZZ0At9gjVTzO2jYalG7dX78J1q34/XP+gOpWazdwH8LJum53dMjTRA8OiU+
qnZRoghEediIvGLwMlyLXSe2YPtin8spmV0CRQtM4/1jq4npblHCxPflKVb8WBAT
X2JeK7K1CIPPYFgJddOjdebaoqRYLH8leq7Ta8ACcKwU4P0aLbWRJq3hEe9Gi9+R
LY7dCL4RU4ZtSav3yU4nZP5KDVfu17xr2dybUs9BUsIr6kOlCfVSw7tUdtzP/uDM
hqoODToeKzmy2FmP/HC09DGP0RyNJ9UTXZX7EDIFTx2WwON8V5VTvROHGW4ejPuR
WnyXcrxojGeLmrBf8IqNoqeZFkzirRe2H9A8P96BiZa+3BxJxBQgjNLUvijolaZA
VKqvqOhNBnpysffA0ohvxPzqH9xYMAQJ2UePqUHOsWVgRh4SL65lqLRzmIXsKtQP
/E+PrKiidtoTpq02Lw4VKH+V9Pc8+HpeoBXHOjEtNRPiDcXDnWEPuGPXG6WunGb7
XxqJVQ4pr3f8tX3hdJ3pXK5/7ldlWUFGpVGSHnue7cDBsUpvfFvbIwPphSKPxdbr
z27e0lmnEEqxYQINvT79k0dMJFB7ijdiYU48827vV6WiaDX9295Yqomwuyblnzus
xrJA4xJ3dns0AcDe9BtEhWqJQ1JgJOrogRzGdJGUnPFAe1YGFTxqF/FaE8IPQxTn
x69nWCBc+rUVKSkeo2kuPUbOklmxbP02ERluhcNmectZssxX3x6J9Ye5dZSyKkF4
BJPWbirVdzISBfAWJhv7ia/9NZBcQVTZ6FdII1++cucx1xsCwShl/Dx50c5GUEZ2
XLwXxMLMZoDYG1h/NUR/dxpuN1GUUOnC2Rg+1bcrNK3HgDk1n3mDcI54knwnFeYm
Vp16KM+J+JNH/t5+6xPRinvTYxBTpuijPGmkM5kMCUYsrKMVNR3a83SDXUO+fy9J
yGDC/7/0pbZ7xWmDDih2VyQJWgfzvYpJLsSs75T4ysDwlmQfBvtXEbguVcpvCgC8
lb88YvD8FY+rB8kzzDmoWE/gX7WXsKQZIiKOmwqttymwzB/j00TFgBWSGonekIaW
KOTTYJ51hA1mbxqJ9ddFtWO9g7tc3PS9Rjz7g/eFeJ+74p9dGY+UbpL2YjFyoPSs
C/cd65QBs3lurZ8YAWVHbbskbAfmwE7XQVTYoNzfYxh5e/TPF1KcW4yYbrlxI7EH
TMQPmvzVleBCRBjrj0bt2On3v166rKRvqVwFbUAbe8sMAV/+BJp1p9oQRBKgQhmk
HBhvUecN82Offa/EWAi7/hvi2yzl0rYI2QECWSzk7ebH2cfUO/J1AvQVo8gZnlXs
VwXpGNkZrOzrDsm0mpQy2g0+xdbm7hctLYxSEl/W2kQ4UHTBfC0Jw7N+uekyQbk5
5rmK4lT0ZzlLIIMLPuGow29HExRAhhKjpWRU6JWfskYdv+VRo/jSACYl5NZxoe3G
7n8ogslQDU9ttU7nBQzpaEgwOxhzB7mfC85x5hOY2Do1BtF4brdq9iPHroeuw1P1
PGlbG4wjKBiCDfFDV8kmGHjDGSf/D7u7VNPITh5AsPlMKvCvroR1pENMCKCyalil
slEKoewM3i1Oxt0g5u8vy7mp7T8cueZKNCgxCBOC3W+YQmxnxEcXYpUBU1B2IsCR
j48v5FHabFsAEeZHH+VVWb/ooBj6OSovx33M9CS4R03hCG63sRvUzccfCcfkNFxy
55xf6SLakntL1pX4pia55F3vdih4Jgj5o0ZvB05yh+3285hAfAuian/zqSZ5bcvy
RPmiCkT8n1d2bOB5tder6tZGgGyCl+ll7rTi+BJsdsi9i6shswyUVgbCyw1YcEgH
jJLPrTeBPyT4+zxhpymsqG12L7sYqDQzRxDPcNb0U7AKI9wdB31yAqsFDbGRclhT
eXcd5wBgpwyLWjxo/uIOi9/DqNd9hEt1L/f6x0SJVmXUOLUL1RZWjxKoB9mzDsRd
T1sbibc5UNvOalSvD7CqH7VSt9CpwaLyWtY7xTQ0Uo/soUe6w4vYU71TIZESlrDu
FIn9/lz1jPOftbZ4d54OCaJSB5Z0T4/3jZXvLW2qDKfH8A0GolpOu1bX0Zsjl/F4
452uKELLMcfdeop8QZ9IG16zOi845PwDvCN9TNdeRBzWszI4pakQJpHcwp4TJz+9
cUlZeO0dH0H43YdFpvpxgEYNqBo2s/BFnKjwzow1hzPrGMtXT4+elIGDK4r7oOic
RMeM54C7YPY+q7td/X/CubpzHwWZjoqGPnatP/KTwny1IGOIbhKf+gRQmktdf5+W
UHG5OfWLzhS3m7nNADRxooMDZShyJuyk0avr6V1DP8rRSeI9SdSfg3DvWi6LwV2E
fKBxJE88CN25C2mdHFEoaLtiFPCzhFf0/5Ru+CawnibNNEkmyNAR5ZvuL3wfMDld
+BF0R2dyhBkcwe74prwclG6/V8C5f/ujt9pB7nkriP+lAD+KEA2eRPMfChvqBLZ8
mvTgpwKYg2EHDd3dxazPyjdHZx9gfmZVgx+j8huNaHYR1UhIpB+Md1BK/Bv7gyo6
WVgNZVtPqWOMYS0qJO9GrCj1Aol/JlV2wHZJxtSyqhPKF6+fq2Ots51tEFlE9S6r
gR6ycyTtdZ8zmGU+lKTlyoYMwRY0Pt/Za8Z7c0wzqJyoIEI/FNjLDvVfW3gqoXVP
Cf9i9j69NadP+cVebIEYdGObXIf9mVRgtKkeSr5VmfIirc6c0FihwO35I9mAzrFl
TrbMcosauLPTAIYuTeFX0S2Dd9IkLeMWl9y43Ug9S0z/hOKlroMxCLR91CVSDA8B
DG9aSNsjRlag3LQWz1tOdpAO1q2WGRGSi5g6g9Aha/2b5RytiRRcyqOyTdX0jnNo
Hg2+rE/biYOD3Y74v2jSteJftBV5e86ypTCxIGcQZkdTtY7pX6YGEe2AIxQxDPEZ
bNRk3Hujkcmq/rZlspQKr8QRYaZa6dBnxfxuRKn4QhTknd4Fz0bsET54iZJHWSiL
w8rUmalDtfLYe85crqo2Y9tb/WXO/gAPIXiJXCp++9akIji5wR3nsqKH6hl21biU
deMMGJnZFLZZlVweoPmtFPMLRGvZfQ+q5YvqYwMY6E25205dtlfBP0p/PZH69h8t
3Yesmhh9Qes3wLr/tvOfvQZY4s1epBW6HKs4OJjqS7xPqddDPEr6m3oEHb8gp/k7
+wSOc3wtkmAAFb2kanA7qn3KDHrcnQYdpj33UeV9F+Rw700wXeJIBFv8/ww/ZCwq
a+OFtHo8fryWveNtrx/1OB7jkEHMPjMN395oOgOwWLKdrgsF6dm4DAuS3If4sgEF
ZZwjrxzdhPjzQQFN4ijpooJmkGRsdFsyGEJdJjRTW+/B1U9AJ84yy18KG7+mU9F/
pT24rMhRLWDIndKeNraiftwj+OKjbK8xkd7earGW8OkZqKGGh3+YPIWoTEUeYRq1
fdEzLETtaTCV3S98WAj5WasJHvH9PeMdm7NS2JtTXUkN2z2X38w++ACAKjYcQG8e
4Iva34zglVakDZMsRECMP74Uh3Lv8k55VSM8S00uqkkZW3vzCmuq/Cbe0+0ORese
I3whwtcsfzA+8NKgA1rWW2BuU8haapjBO8XWsvFa3bEzelIaoDnQ4j3FJcn3fe5Z
RxKyUuJqcgCHXC/HsX2bmBzh00AbyOIRzyCIcksvUrQDJVUSpNR3lxvczVzFJPJn
PB7CAKTBLrWNj7v4tt5Ocp9GnAKKX3/yGklNMieJrgvBPx7VMnjqbg7lgFNz8RYD
jjZWYE+l7sdf9wMUYQf4szj/JcjRtuT0+mw7WT0XFLTZNAYJGVVhap3VEdTnWUES
6KgF+ls4RvFP3yHHhFbXg6x3VTEnjOrayEJLP4y8bC3MdYDbefmcSASrY1S/Z5CP
jlNZ6qLUQUjB6eNHYvx6r6xNLiywd1amPRBNOmMI7cX7zbjB5aq6nhwsGa71jjPw
QeNu/L8grIkUY98z7zFHH4DEgV6F2+zWdfYsjroqAniEmZisDkX/jP6LyOVZWmjM
M1C7hoLqz/hjLAmd08jcjvDSxOa8+Ka4MMp8+e2lZvmT8ATv9BIRT1wcpEOD+3H6
aXMLDRXrDsAd4TKVobDiqtRnXGfMXLsx/QKZkJN0HobGK9nS1gp0MBXUEOr/VvMQ
BZ7HkUQGxPVu7XfVGR6n5Xo1nM1O9/dkf8SDSZ4gn/Lxi1MPtT0zrMb2xiiLfmJy
3SSSaoUlF8U6uyggnLB+tmhqrc56Ic7Q2FoCXW5kNwlF1GDLrJtBKHEFE7iIaGeH
SCaZsGQZKnmqzbPo3ZkI/FH74F0imvhAs+KFj1eR9LEGPJ4Pu7/60xFUU4RkuQ6Z
yF2jyXwItuJNt5H3z0RTd4OidY3ix5NpI9srzwwO7bZD+j+wY/MAAo3JfPF5A/CH
vtlmw5ulIKQKHab9QEwK83v4wjCxA31qIW9Q5XF9dMStsq/gyKDwk6vo22neK4PO
g6EyG1KomuzDL7cOeZQBVn/OKsu7tp9MhI/j9tw3Qq0I5hzyjuSDpsx8UwBJPDWP
8eWhD0h4zpbNaZZJVf5N4fjsuKKFqPB7cW7H3d1twjtgwBNsaqkp0AXP/OiJLYvh
LhpiHjeDw7XWwkJmnC8D2W/te9tW0NkDId6mqdC6J8cXeEh6tSqmXjUkVLBSV5vi
tjIlz4/wSIgmuuaeYu3DElXA6HP3SXjCsHhe+76ABD8gIC7xA4y8f8As6njygIGh
3VDRgMrijGulazXUKJQ/YDO8uyPj7P/wrE25qol0VXqvekBQkY/fmv2P/pGzDwOR
N+44WIpsEVw4n0nooF1wYMWlIXBNGnCb0irKLPVJwFFGfNzakcpl/mzNVgpNh0wM
gK0msN3mcm/rDKEbJjPKgLJvn/Uz1HYaTRvP6GhurMhRhzXbZL4d6Lro42QbNfib
Kj1ue/dE85FWN3sC/pDk/x7dol3ZUP5xgzUQ+oCHyhiEGV1PmasrmI9lEAgEd1+g
Z56le1rsEvoa/MxCQ7awfCYlvhnc5SRFLvszmURrYOGVum1AWyfoDYAIDjzinsDv
WNfTrKRgHAQrC1Y1L00fP2+2Dt3PnL77R7BGGq9ur+cgY5AGhXXpESY4F+qob9EJ
IxUw58ASXhnutqdACe3mGL07/JEIZC11sbZ5Lu7gh6v9LKV3D9ELrqwsAMZ/myx6
CBozy+24323tmGCYBnrsh0iJkyC5+RuWx7wYHz3SH1EpsQZT11Gf3/bY/QpDn1qc
DTIHZkaVdXOBdjem4YTlqlDZ94sWWwBZ7uO21fKM7ZpGw+4sJiCSZ/zT5vIIdjVs
VUhdAkZcyJSDQWbnzjUKhpVawn2HUCGxkUpTe2brps+lsEIqm8fc5kmxucchS1nC
dQnK4rC5N76h9wePhUQbiT4IUHjrdKZ2wxiLHM6Z2xZdlf4dkybKUJhskBDldlqH
iIWRlIsFvNkcXbU5juX4TJnGAsvF3Z2kLcuy+oW1KdEL7fcvstoNaDrPkuyYWvNW
6cmAq4ACagR5RtCDHyEm0ReVTLw3FvSKlXRq71Plv4qRReHMA1p9mkLfUu1lvwWX
CLurbZh2fRgjKfbdOWcs0MmUJeqks7lJ6utZA+EuV0A1AOGUf51d0c6SgMrd1IwQ
+0Ixj9mv0uIoLR5lEbIQfBXNCHAW6ZYDTZrwv9HuoIWbeKTKUrgQLiHha007r0D1
dvMvjXFJnGbYl4Bq2NNBWRib4rZRyodMi8VCiV3k9ZbghS/oqdAsoKjnyg7dPw55
CSVMZ8rLTH7C8moI6I6fU19u4ZWYzH4Xqoc413Tka0eDfBWghwJalxsYI0Ijmp8O
YMw5Hu9DBDyoPNzS5/VUVQNZw02h/Z21a3pzqASRErwlooU5B3I6yPc2Mk0rHiK6
etcF/afQPqXoch9mC+sEtDFJWBXpmmk4A+qBfCDDPjc5anN0xJ5eDB636wjhyTdn
++n7D1MvOA3QvXyR7KPaYd9QONuIH7vcMhPQ52kVstnzm9DMzkBGCOFGpV438jhM
+NZTJpVy3wUIbOFlgY4jEHujF4VRnuBzwuhmK5TLcWhVWfePp4DfoxEr+yZIRDns
6ky8pkpqQBYy0NmtHm5bpkT1dNDgeoxszc5NIeViVdk3hXQbx9WB4WQdhDKDzbd5
7o/hJlwQK3Dcm3sDt3/spoXnq1yeOBNBwzXIUeC78E4tNzrfIGOTzwtAI0PKyY0z
UuS/LC2A7YpkoIybb0uh6EAk2qFlSYRCrr2aoEddYt4Ub75ZognUv/q1ngWPFVHN
pa5tvdkxkdUee43Qdo89IMDIL7ldCEgQtShSDkj0PuopjeQFegedYM3i+PgYLvuS
FDhs5CsnHGtiR7RBuHmDy6/QNO3R/1VCBMSKCfxx1bhMg85w2nhOUyfa6jWu3xTT
3FwbdqN/h0a+hgtUfy36dN/gcSo1d6uruAuMRoG2isvfHpEy4PVfcebxpLlmp6t4
OYAgOScE6ldzURE7HDXoLKVWaQSOWTwclYBnd58NcuGxiWj5mFaFdnaCfP24QmSn
zQeWoeOgP15pmPnzcdlr/pRPaID7gQciWSrvPpBT6Q0D+/7J+FuOiEjjxohQcpp2
9IcBU72uZSf5mFm/F98fxZ0SahmVTkq1XFvyP15YPk00i2cv7ufdqMxaUW8ykAup
AbTgb91Jn3QiM8NbmnG/OEqYHkQ9Ggw2TIj7PR+cWwZturvyWMNKiexu2mvqWgQ1
x8pLr5mdUTe953ijCgC1bd6CXY5Laq/u9ZA7jnL7vSf2N1yf8UI5WbwKvqfOgyQb
mVIU4hD4YxerB+cwNwzc4BM7Ceam6cNz7k4ql1OTKcVXJBkYmOcgskLVQmzj+5XZ
q4BSU1BPRjblszLKqTTIkQ==
`protect END_PROTECTED
