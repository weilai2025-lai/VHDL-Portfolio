`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLcJxll7o0RZAS5Wqpc0IjrIe9a3LyV7q4/R9WS0xWZDlRL0GGtCgZh7Te5dWGfI
GUck+5ZNCtpU7C+ZmkCn8JDJO+tVrvOWB44GtJjltDFG/64GhumXzhuVHuP9GKyV
plaqjgbx8jDWYzZoyLKwf8fxAXBEQAJSNZxUPEBWSaxknLcb5PJLpIpc80Y8liHT
661Mv6r2OHjvbRuM9CxBlhTIyXiScKy8AcGsjIfiX8rKmUKPU1SenRJUkCu1CM+e
tdW7irTy92G10JzQ6u2TwnmnXLb0f5Fs4jJ53jg1SNySSOkPwHOLZ13Dnyro1ba3
E+CVBWzYFdxhMvPqfDEFbQJfYi1DgUWdrxzmgV18qxoVWCcMKh5LNemqrwl5e315
77AruSbDSPdC2ptZ2eFdxRBs7aMlC8uSYAJXtQpQpsEHHtQ7t2kjRHtIH+cONzil
G/+O9GT4ZtXTSnCWZm/0LLPhqSR3hIP3RjlwsxH/Uszj5hmqKzlA4Ec7dPLmfym1
quOogWr7+Q3re1CcMJ8+vp4Z3q35EBjm1GMJxuqZXib4AFKketZ9B8O7boSeRFF7
8wJQ9GYawkyy9u2MuZeGbCZtzNc+ac+lsJ9G0TZITMI0+cIkEcfI5MJq5zFabCRC
1sq0YbSge1eiWjYJ9Nib7jrvT390M2u3uPuqVJ34E00tqJ0DUQo4R58XISUjWzPh
jNjGrsZg7ff2i+dBhYeE4ghnqYn3RzEzkfZj8oZ+DIdwNIcHMsEgIprgScoSTWiM
bh6Em2AGOr9ozanHCYhzIqfuzd3ZeJaUtzobCCTmjTxHditgCkIeP/lXfiygorLY
/fp0JE7MyRToRKJ6vtXDFvxYTtI0Z8j3ZaX4onvchW4ZSCgtVO055R1ZARR5Wanq
+bW5T3TpGU4ytUaepNvmWkelsfW87PYu5JtU5YH8tzm5bgrxvdd8YRtb3f2li6jD
o6Np4ea51tg2G7GGSz5tMQ31EmC49of7N8fl84H67em+YwnWApIHjgksuqlModnd
Wj3ALL3ZWvVbN7xvbJgL0yuEnfHDcOVQHssm/guLFDZgiWC21SOEwj1XwZXBRhDv
BIcbcZM4FIPsvJGZ9sZJh6dIWXehjxjxudLtuBHmN1IrvrXTxCx0+HYVnDZ+0cH+
FpIRZd1izLssXxqvN9Xg1yoIgcdxmTO+yTCFoubBTSn+fPd/cpm4s9vS/uWYVeF0
Tw9G9G4skYC+cB/QkgV4dSHHsDuUh7aiyK8VuW3jd7Hf1pW3Gij97XmMCfAPsUOr
Zx/SKINSatRLwe00rqiw7oVl+Y1p0iPXK7UgFh8sY6hsZBvKpJAKEGbHgtu9O5GF
SxdviBfcLcUUkAFqKKcC8Jd2ZwGsM3LcVVB60w7lZoZXRJEgcclLd8EAqCraA1we
DGm4fs5x1giaP4oxXPYH7fcmHfL1HeuC40RwoRHnL73uOmxlhIO9UUcAOGeHMUvt
HKjnQD9JO/Gg2tjdZveLIag5e9m4oMAGNXMDsqweUhdFa9Ntd0aky5s7CeqyMqyR
VWQAfRFkFlPF+9+s/YwyiTIhNJGMKb5peRg3IMrSVq9TSr9Ij4dOUl+CfSxrOmg5
oHlsXa7TsBnq/Le89YfrtsvqM+cTlykeas8H3Nr3inS0RpUuW/WzdneZSSisC0Fv
3Gq4bun0Mnyk/3+ZnXqcgQ36gJl+RAkfy0HZZciC4RqacTqj6sCurfNyAlPwCaiE
iwNMdFn8EFMxvGHh8VNlUvQJ+53NNR9Jttctpd/7/RhV+04dPnUdF6naIuJlajE4
BgT1JT1jU7gTKLFWdNNRU5FhxTP5mWaPcGWHEvQUzlL2tuhEV/ZVV7dUdKTZ7Sdu
CLN0c18NqUTfXP+mmWNcYPjNK0pZ3d9Y/a1rm3NW+jl0wly1kEpuLCF/kValubIp
PJU8j9cf4g++sOxzlF3oT2ji1l/6ZsWmI6yV95k3Ns2v4qZdvwzuwu6E1Lb3sabq
yPL6HtUQ0nJY/SOnkN+0+KgAY4irH9h2YkpinRVspondYqBa1HkiiEmb0SPWl/Mx
m4Kl2ZoeY4oVMvm0/XCU07LykN1JFi+jL6fhcMZX6AYbIYR5NvrplhjvNflnzjXU
aHla7UaJ3HuKTeYeOnEwyAFZjRhDL/5FDlHdTcnDP57J4aVh3/9s0DBKYbOKR7GM
wN67RQbk1HhU48eTU7r3DTOJlpUbhu0dZcC8CtxP9uhEJdrXpmW2laCmG2gJ1lPO
C0lx3wjdxRK7wsO/ZmSv883qhG0U7+vtoFE8MxPBJck=
`protect END_PROTECTED
