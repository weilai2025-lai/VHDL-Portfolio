`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KKw373C8BC8erDUyf+Q8z7ivp3sa73GSxukI5ifxI6vuyDclcIYF1BTy4uj3h9wZ
f7+i66Az3scxoDLYYAqbNqmrGx6VnCPQU+bk1GMGp5bgRt1+tGOPqWaP4m+TbV4n
E7N2IVu2Oun6yFQoDKQGZiFFdvnS6hWQ0J42dHNrwRfjZWnhJRuN30J0wfb+iQ5j
uhu2A+ASOBr8/rk8Uc7NAZ6Xw62rQsy2mSf/D1YOLJHIGq0fNT85GmB2h/ZdFQoT
BcYcaRY92+4kfR0lb1BQ4etEKYZMd7pBAjCgmdu82nKpkPMHznpiY3btzSAPTRmp
w4CLv7IavnJM7+llSvYXvSpyrnBURYtDTtgJGhHVvw/lCRiKm5K9d/QmaUfv9lNM
fY69H5w39PC+ZEgMgsLwJTp3kBvj99JbYjhFG7/CAvdEJjBtxmlTYmgtqd9GDq2R
2VhmqJPra4cQqushSote1o6OzbUF0lczziMxq9mz+OBGU9BJ/pFAyaOQmVsELtJn
yHPwSF/5iC2V2cmqsjmJwg==
`protect END_PROTECTED
