`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1m9t5pMKi5ICzYDUeb6HboI6NvfvYJbzYorDiJ6FZ1PF/g1Ktt09K2xmBFU0n1+2
BbG3VYng2YSjTHCyJCgh9fPhe1ilVypFxg0y2tkKc7eiNGTQXATp7VwSeGCxkQIZ
iT5qXyOBWHhwTh87QktuyMIPZDcdQQFZ4lsnHV3QfRpkdkl9YNm2G7ZI5SidLGtI
JFp3fo00Dux7K0W7Cu2Bn9FmoCiZ7DDqkkitavBTNl9Mbtp0Hu+QO1htgF6iztpf
667+jY5NydJEBeM0PdSXY10l89JG14bby9/gmpfTW5KCbRE9ozZMViJj2HRvRfDk
a34QlPSYp/Odb2E2FQLKr/ZXaXOG4ADW5S0GsLzOFFFSoD9jp63jn+oeSYXNanZf
Aetc07lW6w7k8bWlQo/ZQYeIqVTaOy3MEz24h0I32yDAPpMWzjs2n2/Fb58yADwe
IqjeemSKQUs5Z/SG88R5R6hFjVDByXxv1rGu7gLX0f0X13+Y+GlJPyQKV7aAJS7j
kcjE0VD3xr6IxV2C8kYebhJtjww1A3Ei0V8KMa1+W4nIbX4iPmDuQfE8HBezAIPj
SvY4IdKOjCxgY03mt3bYE1S78NUrwnUWpcUqcHHE9MQA699Bwa1Y3wRxwg3og58R
/vHSBoROcrP4y8Kal3t5pEAP48Uiu9p08k/qIlGLxxT9ZtjPssheZ/I9jAVIpLEo
nrEpCQfRgoo1TOf9SNbg5/s3gDeFxswbfC0M5Ow9NAevDFhWCg5yiGj1Ds69dwac
Y6B991zUMtPPRptlFOPYd9tMdPbraJ/kJ8xBlEaWbIBILfwUlv+yw0QsyHz85MXh
eC8SykIjKjCYzmVFHYVr6rDQFR3y7sGQXLU2x3OzEMrKShbYHjFNWMMboJnuyx8v
iYjP6jn2mphdHZr9umin0cCRFFvdeQJcC5pVbkbSgLtdm7WAZf2vxs8aVN8ViE/9
SGqjNGBPj78MY06Q6wmVtNJfDEPlfk5BQg4sS2tgDd4XlFMNvg1gABkur+HbCRK5
IFlfnQnTNMnEZhCBOREHZ8XBchwv7XtcHwo4kbL7xFmKXr2VJdpLJMLlGbZDToo3
r+GAiFFZlZCmMR9z+E56N4omCMIqiU3+3H2AhJ4LYXHrYGlTFB8iX0lLyJSWOGkk
V5mrlf95BAT0LuI9i1JL7kclfczSk8ZvpBjGyFspNolJEpcvx/1wNO5iOOpMh363
JQO+qT3MJGZVqA+FHduns5RvarEVkFxAYNIxsXGYJlo9HJwlY0h41hVMfs+ihZ1W
mvye1jFj7bE/78HhSK/sMkqXYwY75uY+R2fo1vhpYdWxh4782BbJn8cPDe3NiJxj
S36mHE9xsKTPaaHYL8J/KN/h2JB0YMC3kfX04c6A9D99rM63S+JhHaZc67pMSfX8
uMInAuhM0vmaVIPlFztQcCRbVOZ+BiGL3sgqn8+ZYFmQnNF1YcvKCCunDO393jI0
XPq1Fjf4eun72eeVcxwetsDT2flvXktcxy4QJC/WIHZ798k+1Wwx6NJZ3m0W2fpH
uuy7o4sR5qud0CV5uYEMK1S3LKvaExc4hEdi+i2y1Irf9qSU7cfaR2GhSp19i0Sn
Jm57ImserUf1MvWcj7bEGai8auszEdmov8Y36Cyv+pLgYHi2FsAHbJm+9gD/nVjo
2iEaluH3vrJPuQAha6UuRRuBBh9opOoEiT2D6tnj6Gi3q3d6qcxhCHbnRmWaZ/1Y
XWl+hw4RXlaiUjwBv64eamx/MNg+IncpMfsdDjmJ9XOuIowIThumOgkVpnvuvh4Z
0myk/0Cvt8ha2Q0gLaFWtrOb5rZNCuIjxfl9O3b0UhcXnTj2Ege4y74dpBVGXg78
qj8He0yCGJY9I/2VhB6NKVaj4jtjXFJqvsKtuDwKFKvvSX9eknooMsPXBlyGh9zL
QdDG4m5JXBpLD0/YuZ3y+oRTFFF98qWVDIksQXwuD8ArQ3G3e2kc6w/pxSl1Cfdn
7Kxmhl+JHmhsnbVkrr7/IiKoXmM4vkSmjVbN5jgrJvyarCSrOnCvo9Pa/5au13dv
5izF9tKHDPduOUP7Njqk5DippTfogYZk4fdkls9ZMD0ai7M9Q1tEcYJ++ii0hhsp
BqLu9XvAVB+aAHdV2TQNwrf35S7ZLG4mohNm2/fqE2Ul7RxXJRDCMQMHJBMPiGIl
bIEhxLAnpvhq/wwGtHMHAvCwbc8nmWakH5BktEtlNSr+qdMeDIhW7xj8zUKeChwc
SvTgHGNaqqU//Oz8sm1RE413h1EljYPR0MSJRcOByipHYDFQrK7jRb5G4F2fsGQW
ULXUMpaqhbYDxIFPZ49Sn+Mfs/52akFVhLGIcmPXN8OghX4p2Nnd54JH5ps67JLr
yKeZjDfgJuzWF6cQj9ZAFw==
`protect END_PROTECTED
