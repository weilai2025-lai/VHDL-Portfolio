`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
91ivSnoh7tGTvrWD2ylK9JwyI9VADFGqjOE7VErZaFCpsUNXDgQ7Xwz0lolfym+B
WIfjOaGlKVfff1rQc5jzIfQoq0PQR9V1MKFrDGC1Hv33a4Y58mRQ9ydtqW2Ak5Bi
ZeyLdMLGC5/RQIgJXcjBaSDNgkaV8a0zs/6WPX/qxxdri/V9b4eHLu2mRn2ZPB+3
bOJEntClkylnLwUoh7HdFlk/MFOczRVqBCXUlGvLRndCO0Aor7UQysLYW1pqcrON
lOxEdWkcYGc1YjmE6gfzh5EK/cI3Fr49TxhdZpiEutjkC6ny/iMrYWg20bmaBDyh
v1MF3NoF9toe7dVZsYDcKHZWVlyiSo6Q5f41wlTuMKJQDpyC3CGiLUZ4Oa1Wnk1M
m8avxnziPVGfwH8yDGAwW95i5Ce+pPNnkaSNq/JQVSTQl2wEKtyAxX9oswG4fJw/
NLSU4d7hjaZ2c/Kk8dO8cAwaiLNF6FE6z6/QptLaQriAZOqb8yKmGe1y+IkUeK0f
20FJS5RjLQ19uYHVRtei8kpyHut1CvbO/2z1hoKfxCetNI9IVlg2gsEJkO95jQb+
qIcnvyTRLVpIAmErKkMG+xGa2pNHN9dGuWkNF1e3/XvBwF2OFROJv7SB7k1A+5gG
ghpigmGFmpToOzAVT7XBspjovmSeb23nSStFiyKUN7M+URQzZ4awPBKoc92+ftQT
t5yyt7lK9AjZRgT2+6ie6/2VPSPfio3YsPDpsbw5vQfh3DERQrcU/tpb3KQe5P8T
luGOaGc3xphKXzYDzgvm/NGmAGeSSwL7esp7Uc6I2ufF2BbkASZdXkN/2F/b9AKa
jOaGLollOdQRKOrzbkU6yMOqqPyzROiG+Nf8Vm1/BZ/iKtVg2r+iY+pGPCiKz9HX
UerJtQAeQtc3sGhHUZS7P6bn86nfgR5acqrm/9XvIkhesbzOc00/2MJ+VLkCx7CH
tx41I+TSSSRc+Ld2ONzFtEc3ACyXY7EOSUmyweqTywwq2N444KYpUnJk9xS4siGO
QTn+JXoT44JtjiHz4auyiehxogarzPTf1gg2ayzvfoUG9O9fTLww1FsUm/PcMgz5
AGpHxFbF/ZEwpVdhbJt1NwyIueRWgkej4bDmr/UXBZpI0JG0OvaKkSKEi/JY6Wud
zZ2nIpSgySjGCURTPnoWyrHnPYgoNp8vu2+7o72szqvk2BwnxSXAoWMdN1whuZ9P
gwcnj5NZpB9XTrWLdegAisIP7TKY7jKSED0DzDBnTxx8ZQ1k24B0m8O8DTWdIhOE
6lzLyCfkbeqUBOdSM+Q/asRyfqtsYis9bjfLUVh/ciTYBVVfuLqw1a4QM0WBqrvl
3nP5iQ6JsEvpfNzUFrMyVmUKLb56oQNmdlDToOZE9bx1G7PX4fyS4dJLYn4qi7lN
C5LSg9+/J+mx2KmgbQfHaXddUdPmgu8iomTy4TomDYtctkLtrzvxj/qfm576f8gp
ieejg4qvvccHaS2Lfmx6OkiJdYplWrL4C2pjuQWGU5oSPavLwflFQzNVfcKgm8GD
Gnuv8kwqKzMVZu/Ox7gs21/QvHXdYc9cPf1/LECb8OBB9EuB3DZ55XayhZjKEmaB
ozSLuqiI/T/ofCpNzinVI7YQr8wq8awALuIaOOzseQkNckK645/UMFKYGwnW5kFY
szung6rrzPKWf84vnoKSmwNpkfj3gOtJrPx/4aOD/OxNeqfhi44xuPUuX6Vrneeq
aILOrc7IIhmywlaOpH5l5kdJIhMuPQgg/tmlg+6F2X4=
`protect END_PROTECTED
