`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MOXVv9VD+xQg8G/jFBp/8rxjEFjwgyig8UlSI4wnNXQuP+JXyP10IRi6n9FI3/7
3E8ADoYIDcet7+9grg3Xj/VQCFJp6RtnpLuHAXjSt0ylPMNCj0Zy7vcBxtQcGSkt
rQMEh5UGWLER4T5vGPo/FFhV9jtvQtMwWc/raj6fKVy9vQ2sG+qd4XOktbqY4Zkn
uPnMyxLJDH1IONR0Jg72fokCfMhXj+nvwi4opRgFuTBIe0xnxd2nYfT07qsNh2YZ
kVIoNoqa3QlatpOhm/jnzOPWZNi+hKo/sfufy0M/cu5wBNQs7gKW5AT3rGTXciIx
13LMK51mfmUmrSaErHO8OGC37n3KR1PHP+j2i897MJjOPEAkAwdFAvm7N/O6dzcT
UPL8Ct9Clnxm817+fFgkVOGYIuNrUdZW82j0WNxBQoUXU4aIiHNgD8bN4WhJZE4+
245imG53mxRHIiVwvXNhX9g5AYe+VvUmLP6TqbHOSSaUv3xnxoOlRWyxL67+FWjp
jOeYqp38QvmwYcEv1VzImqVyyCoJrjRiZpf0GGH0Lxn3/5lVN8HZpKiYvxfB+te9
bkDpk3RVaW2lwqIpLTHfuo65ic6Vb4+Vvv1sWSEE7svIsiS53TE2imnsGThTVKZb
XMshp9H/IrPXJxSTGahbJRy4ZA1IUuAjvMTV45EOQc5PUVYMqaDgiHryNXPZaMIk
GMiz9Se9OKrCDAgPwlP8EXYkvwQtE71jZZNYuVSDJDRN7cvCmDqG/qXYBgXqtfLH
NoMdg/Ez6EOU1cUahOBdr/CxLV7I/SG4Q6YQAkh4nQVq78X4/mDBKLf7+p+ErJjh
30us6JqUqY+4vz91JnkuVv0IsGqbIO86fIHm5n8XOY3QrSN6S+VdsEwGfpq58UYc
rcI9S7l95mcxujMF+ta/B5YJwXkvo2tvUwShl6ihTGt4+HUWR6P/2V2/DtPurGS/
sFIzkPOLCN7XKjawTTOcG1vfM/6M6DDe2tKlmWADW0OK/3wcuexURAQCR6jJA6kh
AWL3iuyxwygfPO6KF7S4MtntCDbSRuE1/zFqUFQULCsZRmLxDqk4BzWtM5xX775I
wZk5jS4q/DieJzNVEDyetL8bh6CjsmDHYG6Lh6XAswM=
`protect END_PROTECTED
