`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFs6+LQISEZwxvNf06WjHETVrIwj5TJiL4TacRyI7ZZfgeJagNT30V1MsszaFXX0
A+7V3Uun6HuVHwcrgm+WzFQqv2ta/vlrRlcEwy8iT5yhOM569RwddlpsPYHF28mS
FcXgRDqnpfFIM0vwA+Zka2B2XTSGh7pcv1TqyBjVWtOHpP5A5EFdJ7V4IIuQOGqw
ZGeQAksxXfwQe+AiCWvVsfo5ULYw9VEAM1o5kIN5LVtuPN0ekJXNkXWS6ZLsqUS6
nHCay+vvugwaM9r7u5ekCcTdyPLNRKhNX8GnJ7RVPylQfJxwrDw/OwfrwL7Y4H9X
du+/gYaGg4Wox5woQfzaecHjbE3vpue5M9lw7nRlyJXCB+1sHMqtI9Ml0vFzZuEh
Zo+I3P+E/FlCNrYtkYzMVGlLQCq4/WXXTATRXSaEjlgBPLrCuTKVY0t/pv3QpQOO
8uEeTyZXRyPhTMz7MO5Hzd0oc5U28AoOhXKavyWfgKDsB+yEjBoCDyYqZAOBnfSa
uxqnwbk2Iz8lIskaqnNT4qnjJoloY6yM/voT4P8xydK/gqEj3Oa6LggewWm5mh6l
MSTVb62yMLPrUq5dLJIw2Kbh48UogBgLXoGUw/fjr9mRUCxtFlNTxfRtU+WEvZXg
WrItA/AJ/mf4jV4UnYyIxS6F/8qCYcQ6PHLVxP46BHFfnK8F8hFbeQiAIPDLxA3/
2efKE/xKvDh8VI+f8KZaATVYSkKCSIXn567h8wvOsfbrO5KWAOtpqHW2PoA/UBhQ
QeAnCKXE1AMU3qL822FWgVcrnisU3c42zFS/+6lyC/d2PEKKpVaAuv2kx4NFh9vQ
dr2RUPVneK0u4FYnmgre6y2O+FC+8Q8bM1ox3/8JtM2pWT+tuU2yJal+W1vofY6r
TpBOgP1kRs5SaUAwMBtTmcP3ZYDMV2OiRdE22Mslp4q8ROjm9oQnaJUMrBhRiVTJ
2O0lZe5wK1XGKzn8WTGhkJpytwT4+5Pm/UFHJBgRTseCeu7k3A60HkVLiTJBkgN1
9Xkjyj0Y3f7VYClrI1vy5jimF3ddVaGJ8mFvAlmEqi62NW9dBUI8uBKKMMrC+W+2
nD48ZaSwPmOrX/aazoWgPIGoxReqIJwVhoPbKCtPiS9nyVEzI5nd/yKyMhYibk9h
7z8WtY+nfmPVRxVFVQdQdUweSrhAvx2Ge6SP9p9vsRh82Uz/aGrGtRU3dN1sOT7G
by9Q7q3gAiIGiqt+1I9c3CPz5tq9JUCR7MlEAbGULRcEf3tNZF8RBW742aqxFMFH
zdu9lSrVP5l6ps9sCZh8DUfxInEwJcLCSe31FXsKSAUNM8aliE9RU9M+JthFoSTP
xV5k32hX1HJlF5QJpYrrWl0ORKidJaVn4mk8SLjmdUaSIir0rldCRMENaQOd1BBv
DpSL8cgILKyUQIVNYq57EFnccrEf1ir1idQTA/sdX5R1fE5mJOZcTa+2KofUH2KS
lGmyzZ6thaltqbvTddOdhzihMi6f9RA7JTaDW8CED9PvIBQvkdupSLECde+//h/3
mTmwLmKTDKV2fdGgCYGrjn+t/zMECv+OzY+hgmBodEtAPhughY4skUZvKfCeaXuQ
/y82k04wyp82pnQ3Ng8DUQ23Lh/rRI8F7SDVXZCOVHytBQ4nEJv0wPY1ODOaAmGz
uiwQJYNIGqFF2HDdRKkvYb+MHY9u5hP3e2H9tloZ/L0xefH5WveR2mpLyoDmamQr
+SLfLCrDKuOsAa6YD+pjhTEuHrEJ+x105oBFqY4kIfKKbxK1O1V+21PfJbRWPX4H
bScBEgmVHa1rPX+hzwzEhSy7S5NcTDeuUPzWYE0+Cr6YRiFLxxC2k0WSTmHLG5Av
PdJTtM03MAzzBFOwvWAAXUYQ0MsfXdgldkLZZVgwF09C2bXlmgwmVF9xLwLqbEyY
rQ3jZjFoIfBWDAzstTLV6eV4FGn8P98+FqTmU0CP7/r3kle/bfAGQAU1SCGFTywR
Jm2qCNFnrqkpgObrSCjnBYbz5iR3QfTDb2rZdKs7JyR0y4XJYCfTrnPxqg2rQTwG
AKwanc0u4KRAs0TPlYhm270dIwYuGNVo3p4TBS31iRGfwlAU32t5bxAj0WWa2CU/
MewQFZTJsJd+GfKYVWado6frhTtZmjnIjblmW7hX78ld0Nts5u9tNu0XId6/DWtU
YYRGudmffe38SNOid/WgqL0JqVyQ3mTF6OJfUdYXtYY5ubS5aMuUyItZVptThaM7
L83xf6XTMa4yVAAtAzMcgtPRtZRLAHnnCQ6GxShopu15NCaBaX6rOt5rZu+43yAb
JNU7ctjvUkQEHaFu6BjIUHvDMMrRLF6ckojhL925i4abWP4yXuHaUUjXWfo2WaXD
pme8N/m5piboWW7GiNrw7my+CudxcYYrefwKPNG8jgHnkcCudRhOTHYdRdCCTppB
WTTi4Yok/pJjcP0yF8wXE/xqZdN7aJc3E1sDiiDBU/6pxs2tzbD1F8GWNVi0OqpD
ygRT1smTsUJVdR59ssVYvGlAUpwx3iaS1Md/5ZMKBtQEYkMJXJIXL6/O/BCY69sW
yT5qcK++pX5yjkzM47plRRghAFKncTf5Lg9XwW4dIkbW1CFSU4z5VUxAEEa72mzr
ZIT98iCSQOgl4gWFkOKFXWFxaLTusYXGZUmuoOcMBoTZdpQIdUxp7I76oOsOkh9r
J48yfu1vexqqzLtWbDqK2Ibx5FKFKcCvSc4ywAFfvbNfT1LqQ7P/Np8uogmP003f
qnvZXJdc9uhWGpFuXJImA0CmNZs8Pripei3bmjTwdfTtKsBoNPUGknFemXtEcMWe
fn7gSuR5kMxQtQY/+utG0rDXvd0bHTprqlpwWPvm6USr4WbZdz4gLfTZsEP0YaMH
zTrEgpJgaQCk57KhSxLG/5lSqKSm47GIEZBc5JJ264Vo8ONHEKUornn9/5Eoq0eZ
gyS1uq9gFo8I3XTlIFxLdf/xO7qO8Rb/mOiFsvLlCj8Z4vjyJIevno8C+5l0QI6F
RPMogurnK1R/rdFJ8mHaFeLFn/WDlu0iJuzdxzbqSZwxN/XaIfm8zSmIZDu4ZOxS
4XynKDgzOI8Ui/trxi8A7eTQOtU/Pe2WPWF4FLCkU3ZYmrRs6CJ90X91jjjFr4kK
d1d5unscqAae6OaDx23GY1aSAchI1L0IAHM0ZqoKrqo9W6sjEFyYHGTzaJvGKQnY
aavnbyJoZTZVmner1syR/xPQAQdOP9qP6Reg8/C6pSSDbiiWyV/OVtG9Aer2JOYs
7uElJkkeJhXy4YrXVwbuqf0RfbOefE1zCtiJOJB/qMGlOZbebLfWLC3MWQTRw/MN
4iZRPUh8qdY6q+pbimYLSibBcz51ByrPyudG+NfE85121alioMYzvfjH5hwvCpUJ
3RLhbijYcQU0c+hq9d+RYIXcYg67Ms8qxmXW208+4t0F5taFdxuDmd2hvv0ndej1
vV+MSVyt8NplKQBW90lL5vTRPrWFzwDHq8kkmGaTkCaFAqSz+eeZ58C/oCBrrOVZ
zYb4g3THCPNToLfgFjy6CqWxy8G1NOtwwDxXtPutCG3dPj+NSAjyAy3qWAVG2mcC
P/fJO84i0BtNdAufZEVCM5UT8NpbIlGUp5BKk4vHDrX1674tAsJlkRyNuRbDOT34
`protect END_PROTECTED
