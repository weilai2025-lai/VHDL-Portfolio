`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uoZrlcwvBcVOig7v47/T3LY+ray9xR+IgwcgEh0XsNaX3dP8X58tLRa7DoELP3f
YZWlTouHBD5WDTSs4N+QcGDTz/SZS3X483bJfyZIH99/dTT5heVRPe2zjcT3QO6h
YWTMwpk/j4wcVldVItdrBvqsDhY5tyXmpc+94enwckhtRfMIniN4qXuZSZoA+Dd0
rAep2wP/SLjkBpZKD+BpTx530PF4N2OFS4nWN9/rOYiBXYG2mR8z1o7EEEoPdzbt
Ka9OprXDu66yZ6z9K3Mo8ye7O7j/TdUqRmyQ1DdobeQ/njzY4Ya7uKMZRUZ37i9Z
DeAzMIz93I4uVj+HgfbrniJBcY0jZf1FAiYQ3ApUVxfS4lsySoVw6fPi2DzjPpA1
+JlLyQdeVAirCaP5WziZkURDWrCwJrlEDcv9BeDd/vR4K8lygl+7jbIGbfJEfJxL
`protect END_PROTECTED
