`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCE6mGlNrIwoXgAcjq9VXS3QddxpuK/qkBrIkDTALRPqhgSp58+Enyo+r1vAFt0c
MpLzpfmbsEL2QeUzda+KkG7U6BUMGuYNGhdd9nAiGaQRGh1+/byiABPaML/JaI/j
J5s/guAqjWFnNys/ZxsfXIFJDimnGqYkkL5oW0IZd8fYs/DXKDIvoegYos2UFqd8
ydGulP64GcZ79gaToOdURnKdzHV9aL4Ikt2JpaoGNNbqZ8ayYDgGvEJS3tHRVJK0
rYdemfpteI++zip3+Kn7HinfM20aG01BE2KUEzFBCLEtFRtXj4WFOUIcyTH0MvJP
laMqn/ULafO4f59sifCUqL7ohp7gEUgnsr8+E0rfnZ20IC0hjFUDVvo22XxjTnZe
ELToHxZOUZM47XW8jQPPLRpWY9Bw+ZBVgPLT7Bh+ekuVCSXeXOWRgfQOUNatL8QQ
qj3SL7gXMt7WAj7qIbUBGfSIvExc79l1u/rhjw/wbV+3YiSurjIXuUSZFOzo06ho
f1VAhFxehuYPcuTLab2NUuTUFzYoRSFGUZtWzDAx5pwscIewu7iCEwITyJetlv8i
IeJPC650wzFXSZBormh3OhEKnUmeY7t35kzMfzi7v7Cg6ph/OG6sM5b4uSVTT1jV
FHhGu58pw3dAnnnRNVSCtPZJjjWTyIY+qN+DJHNF3OQvp5Ppn/k7e+JzpcgABlHX
QmrLX7wacC8WadWyQ/vmsnOaLZSwhvWppeRJBKn7gM0rVUThfUtfV3dBhQY7pyv5
pJcV3sosx7iA7nixAOL20QFg8QFPBo/LL+pnOjFidb6DNSrS8jls4ml/c6kApKHM
eoOyTAuHdD5jk+QoIj7TNWTBXtrC5DKVabn8DX8Z+t2WqtuSZHGulqzj0JS3XRHB
GZhvcfwgugDSsi2+2bwGep6Dzfnyz64G2fohnxMoRzUhYgdCNcoUzDqbTNG1LL95
mE2SIhUl4zuRy6N82e/bFs682zsb1yxqO4+quGKaqQjEZUJnGMEgXFv+ql/J6xQy
VRQJGBPo5PfRHfNzJ+Lyo65o+9LKQJCN7WXszPT8Wp9D45i2BIm4CPsciW/8ZMCD
AciY28ZAAtbTrHv7sGtZMlxM/8msPSRQymU3+NdTYUMPoBdZ6F+ku5BVyRP/gtiA
xci4yqoc0Vygzpk3ou2Vl+DtZIEhC/4wNM9G8ZQt3OxcMkEyyOWhpBij6j9MnpdS
FIvRdYo7mpXHy7Jp8MP8P4q8/nZa9YkClnvdml0rIiR/evw29GafkjivdnLj4VyU
5Oh2df9HvvfNFuxpPoSKOm5uF8dbPCpWRqT7LbbFf09yqz8TJ8ISv6/mG9JnrD3Z
krf98+rqi/KJG/jLGzN9opqzeFN9UetpYKLhW8blrT6xXRaSPIv7Nwwpn+OAB7kc
w2ksur0fn2ix/sSZwL3f3dVkCcPsAJDWcjYDtaYpeZjsLApwfjh3FGD/bBJvzmJ/
jW57CpQcbIpC5+UP8zMAc4VPg/TN+yKdDce4JYDdJc2pdvbOJdWMUevRxD2g0kCs
DaKR2TumGnhqFiS8BXyt8kvgBA5hUpKZPCLBa6wmCqrwl8q36iNcfxOR/Y4q2I6H
jj1vSYoCs4sHLyaQb5vpHzCIU9e/RKLkNb2ER2KRA7aJQy2SvIbyF4MJE3rD3r0s
f7ebY8Fl71FOip4lutzvR//Uon/cqzGx2Pr24j5mFLeV4tC0L2cxY4N7Bli+HfI/
x4zCYs+ZiMWP7k0vqYq9VnliLsfh5vbb3y/Sb+cYgDSzmd+LXpOMbAxZvv9F1e4l
jlDI4TeSxGskwjRhIm820w9tqMxDHnuiZHDEmsb2I5Vk5lKYcbsTxDRV/HSoLmoR
C7ahPFOdbdys3+cXTa2e24VfM2bJcqDTyd3YTwjv0uY8kP13MGo/HptP03U5Gs6B
wxLSOlNBrllj3xxCfX5f3KrE+Sy2r3ebIfooJ3x95P0Mu1DpX/owtmmRQ9/NBrKm
fwPi099juR/CyZrxI492O4OFBX5xeOBivklimyM+CTWgLGbMxplwKxDo0xglbBTN
E/WKxVuIkW3YKPTdr2L7L7pxrgeoyvQ3wMWcR6PWPaTYQzETJEaC0ySwkQGkpWhx
Ub9wIJmfs7vVCYRgnsEAlqSSS2rzFps80snWm9yXKRl7j1wog/nMqi4M5OMy7Gpm
+XluATwLl+hyLF9o6D363Y0lrl3WgrfXSRql2LOfrVJmBvqb8tyhdgBLrBUKhsPn
py834/Ew6LKhaDSSSLKFGZlqLHhrWGq1yhV3JB8u8B/MvfFHHj1SBMznQT3fNity
57oeaClR+O0pFPsKuTkG/hPc88Uca3hxjwQ9evxlWtxSEuqqdm4at8hM40UXs04S
/j/KaFjoC0ef4ZIUI907x+aQ8jiRdFBmIkweTPwwhnjqOjZpKEP132/I9q0sxSVm
1s4Q0QuZTVcq1gS+aJCdMx6AeJPVSHaZKfjIIhVb/pGQSD/bXa4+Np9hWrMQmBpk
L7TWYfxLwt1qmOGkqBYr1NVFoagS+ENaLrEZlMnvH+rySbcAdteJbodrTABHfZlm
0F2s0o8FGo5m04o/0FjOvfmHEHGmBaGfezCJPAkdExPUoh72Ec2Bl9GqwaYpbEKC
hxSUNNog0aHyOZKdkCAjjqG02y+UDF57fxvWTyJHUuL2SGke5gu5+0RGhjDTBGZp
exZqtz578BPG1rE9cMhUeiaU75nHyyQ1v/RgfqA4idcESm819+iLLeUOI12mX4KS
rOZEL2ctudMmYYdIVFNk2oR7egOFzwDBuIXYN3xkWHwz+6ejwSqBQAz4StMKKkDD
oV4H6VC0SIEmEF272suWWFVeUPC3v4S3ppc4xqAOjugHXVN+7vKsz3OB8CW+gOw9
vXmnFQQXsVTB46M8LtztwKtrWBwMd5uka1JO9827pZslRS9FhIRnuHIKtfIi/kCr
yjP4WF2c1hQKrDRTMR5jKkXPa0iNZ3tawZLHLAXrqaiBPAKtiMjAM3xgo4fy0mlV
I/ugd93Q2bXoDDlOdhGQt725jmljHV6L0ybXg6/4oUX6BQ7GtBzhWRQ9SRzUuoNo
71RJ5eCcgey1q/sN4VEWrTq7DXTv49b+6DHcJqhaT8b+n45cNK075+imc5cE3yKi
8rgQ87/GqKdn3qAucWGNWjmU8ollHxT1dHowBHcdJRFKpm45MgKTWsSOygRe9sy3
Zk7XQ1noA6qgmD+s8+Q0ZTuO2TactN4Vg7+b0bJSdw6PQMf/V1+AnmnrIHNBTqjt
clpj3t5QxxjagSM2ynAvinZZTaRUy2yRkt5OQ/JbPuuPaC7It5CUEt8jOHacRduQ
2ZwaH1nzUy7Kc7joJVJDCkZiiavgG5Gw18Xwy11OJjQEV6cc0uYgBXWP+3ccyIXQ
380VjXkkYO4PrE6Szm4i4DrtedQov+goSSzvqjKwpHoCeuIUp7YKeSOQU+ERhbrn
DoEGujlENtmHstPbgv7pO/7WpONKJKyxAdq8768d6F7T593ViBw4CQuSTbom9veZ
re6CS/LRqe2B1OSr+cz2o2oi4l/+q/Osa7YvLS+zT8l51Vr6kgPE5tgTEwNHFYvn
nQ9wid3E6hJjN9ExvqwOYuO6eNLmv32iHCzo5tHq9FpHG5yTsGsPLxCyi4exLdeb
XwxLTVFt7SQx+2Fc5YJ9rVfv+kg4mJGI0c7ZoZqj3DLFu/h+FZPTAqUy8/tN+c5e
xdTMiP5XPM49kSMjOHyfso2POB9eqesddSE0KDIphbwnTCl2Btz7CSQObesrH/Q5
8UdOVmIQnsGZQvHk/iJUh8EkcJjNMexN5YAxSDZ3CSZ/Sr5otbxvTB415m4JAfPE
vVwTSRbCPudhWcH4hytQzNw0f/rbkRvXJ+3wQ49hnLcZtvEl+FTjeKlShxK1ahR+
rxlcGT4zedCfzwKGiP1kLOAK+OasahiZj5krI8sSt4BllPbIL2zTr5/6ToiC9iGB
JM01E36LKYfKFh+iOS2+VCUtM95xm10mVJB3kaArnoloYltlDqciPprRwp7qpi7L
n6xu4PAZnrX1ueFvDCU1sNGYiFckiB14AE7bMsIhtuMWUSWmVlNIDBw40IJ6yEV2
ZKI6wQjl/sBSJNXs99lIHX28ixME9mJ5twT5mI0SJFhIsAR5CBohiUkGULjGIIpL
Qw9QYitbQzR2HmuUqwI2IiZ5/p1dhh2uQnVRFCVzlPydjFdJ3tCtDKKP5G2gQVEP
9NQct8C/P40kD0ljTt14YSsKu+n6Wju681fbmCDOe3faw/FT6D2g4Ofd1HOqQl1l
qKGZcKuy85cb9nVvawDrw0pd3ZD/imq+8JPFiJPJCs6R3Z0+rHJeD7FAKwPK/oWv
SjIIKsXNVrwQfbBNPZracsKCdzA28tJ34ZmqrBeClauT7Ur3x+oVYJqOXW1jxxvF
VKEvd6ymuC3XlLFtO8qdMFQOUHz4idk4KmD68AFIC5yInjFBmGv9myTJt/n5y7pQ
`protect END_PROTECTED
