`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3kNScCkRlue/jnkX5xQL7SCpHlinPoomY8Oq5GJuzfWgyWaGYDmwHeXjH7W7MSC
TYrfFJt/AZCg1xfA9MUnT2mRhf2wB3kqQk0SJB8JEjA9pPZjaeOP6Rh+KvnvAJUZ
R5uEzz/PJ5aJE74GuAkbV1LR7ElgrPx22gYE8VLLRFh4cWTmU8o4E3Bhc/X9CCsH
P3nmlFZgQO2HrgFKKbDYUP0vwhMxKE8LX+2hPl9LIjTp0ASpRBzmexoqdQH4SjSx
fbV2BNqPrE0ucUfReUPhsnELs239BaRxlLiwfGJEVZbaPwGeb1adV+yIHnLlhWst
4VRiYJFqV8FO3GGZjh7k6SG756VqykWSHooSfP/dAhgukt3VmBrd9HPeCKs/TQo0
TwDuh4vYYq0sH6ID+6WF/JUog58IVmbuY9WIkQzjVQ1ESKJqxv+sgMVC4FWJ2PA2
j8/7Y+ZKNhjlUpsew1pFadz6rcq9IUSAbI37yH3TnLRYUnfFb1wfPWFI1vR4vZNE
jp3kvdbReta9tCvO/Lk1O0OEGuQi7ozLgJQqJhIUxQ5iWA2zFirF0XS8evOsdDK5
nE2cpmrOMWnVQR9lqyosfycvSTN+KZAuFWVOEhu4GusRxYfug5IR+e/RmAtrla+W
dDj1TWIhPhpGJ1mdrt+WAwiLGtCyhPeJdyj1oYQVsj05JOVgCwMQeeFKSzNfsWTc
9JflTmsyHOjE8ahYLSAUxtELkWcgREQKGLrvl/IJkqQOnxfAIf7BcaN6P/1ewGmW
jogvU5tLxOS1lIUVASln9ut+jwczCjMFsTThiAI5Hn4NDCdeCVeF3CUHm78QxX2Y
OwsLQv0PR5I34xUTJqI0p2hfMfpe7XhMHL7wiZGL8YWB5YY5bzyp76roas5/QpWu
iCn9V+hGK7zRAiyb6RlAZBJOouuQxUXwNLM6wOEzil7rCPC39FBRwXkyybf3mtGw
p5UphElFDyyL3axV/T0dMQSq7Stb1Q+LfW5azCngQ7zrhZuglzWgJXQAOcEvhncd
b/dxx5LhHkw9pcJ0iLEeQqmFsUicPLBs6u0/nD1HkbwwObjOM6j6k+/65xvjDdxS
8Lxhd1z5o4Qg1jRoK8Ty7EK0OsdO8rKs7x983lsCTFlwqf6Uy2FY3VIneMTZIWzH
XkrO4Ow/BgZTBQsvzyGEQREMdnI7ZpiGsIPGaj0v+otepRCIjcGpFQYw7eRGapEK
u+cAdjAjDNMGXxxkxHClFGc/X/+ZceeDEJkW/xWkc8oziZ+Z/Mcq5v5yZXavvbco
+Ny75JeitHYm/VuNa+RT7/lkgiPTEm5Vj/CbWpf3/Gu/IeT3Eh4gkTnNqcXA2NdV
jtEUJgYWM8MFvdmm72H4ZaB1bXdwZg5+lT5QcrtjVOGUsvQe7JJedc4DJr275XO7
11HOg9ylfDjJg7axQd/yhA3EFcP4aySZeSbTGzeWYf64YbJ/TLnJUDGHBzvY7Jpz
TH6bRf03OLQzcjzH6Z9obQoC9qhdG5KSWRaM2XeV9N+krKsNBZxrUTrfxQyZEWVI
qPegRIDtvcmbkEatFY841rEkqAj3ceEYIcc/mQeEE0KlIFOLrsTtvcv4QdU6bttH
1iH0cm4EZQsGfgD/b3JFNopXsSA1GUVRblODSjF6D+UZzVT2UWvCs5fCWsM5Dfur
XLVHsSjvmCWNvWgt9beASq4LFYSkKtGheZ1iqkPbPvEwSkGlW9DCXK8iN9eGrU2A
tqQy49wBeR5f/MpQ0n1c/pdS7u/kQ4FJaA+f6PXbLa0RzeXJac7MdlllC4Nv3EKR
uUbpeDn2qSEhkmhgoxMCVj0X1fnIAg1qeR2cV0BFwcQ9bf3NwMqD+bDNvBj7lgnT
k42iIABQJak2BvjBTw9pJK2MTLAjY0tjP1S8saj7A8Lxxmv7CmCiJiOFvuZor6c8
RsAxv4W1zb4hqWkH+xbJb5QDRylS7Oss0k07RGeeAxYLqvVHtPhBP67wQoDf+fgg
2aFMuHDV0RJ3LY5X9bYivGFNiKv5YNR/YV9qF49F4BuvScqHHxYev8c1mhyMlH77
miWt+mCdOWJTaBJt0Wy3ygaac2Nqv+P3mtGNGMBXbTl9X8qQmZuIXZHm6sZYMU/E
inU4Ql8hGqrBIMEkXM1md4fslQPaPNUUCM0tTKJE+XKrBe7EjcJK5TT9gUju6Ff6
n1S9MreaOjUjzPb1pqXSwrLXE1AXl55avKcJgR7I0PBUA40+qeYF90ATfuPgcPbV
VmwZSSy4X74USGvWrrc1vEW6giG3Zw9CCWvxY4ewPK5D2PCLf+2W4p6dQ4JX5eM4
6QkXoI6Z85oeIZw4A1QnaMtzVFFA1acaVZKxnXsz9PzW/6ngMgiM4PwckM2zQYxI
wq56HSEbhJ0WKLM5Yj5BuRfrPHDxJQNwdMaRFZGKZgbfHINXEwciH5zIJj4PpE9y
Ulsu1U1vB7wJBKMdSXO5QNCMG2Vf4y5Vi1Kcq9xjn728i1wpuTrCEZtVksyM1k/I
GcO+17hZvm8NNN+VLMW3QeqIURlYdN0nh8wdIUwSPCXdCdTLYnukLT/eoesSBMwU
XnIkBgXkNFMfDNYOLEEFKW9JRY0XqzynggaJHm4r86x8xqu5+54Q5RaSbcFhSDpz
tntpMKqeDrWQEK3kAyVmg2Ex9VUSaOK6DtfQN9yB0b0LrBZpqFPCnwIf8Ensd1c5
WcWWCP7OghcWUTuYR1G9XXtf9dMUqfPq7u0zx4eI3LtCJ7qIG30DnWz+O5/ox1Tm
T9+azqxbr04IhhaJfJJbMEYGMdlRlvmqActwulcL3VgZlVfhmTouxNxEpx026lpk
Ue36AyLWoE5TKc8q7eLnc/ZFFzuGCwkP4t/5bdlxPG2NW9WIHnGaEcUZKkuLKLVr
TWXgxS3pEYFhYVCpFNJBh30afONr+W2PGMlwSzKgetz2GHk02SSdfXdOrGZUk87R
PVd9S0J1Iv7a359QpOF40HU1Tmy3K/mnuhGBZBDyDL3R6FQKWIqWlFHaCUs68v2S
Ot1hlhIobOT7cRCs0p8brKVP+QdDwms1C1eLvdh0jYFT8IASHO8PvfVCfUTzEnS5
26p5nJsfr3o8njcaEfs0BYeOc6MpRT5pENoCHAwWmzYmXSHkXHevth7POHVgDyZu
81YnssOS2BTaO+IQBG+TEEd9s6qQwI+O6a0fQNf7hWuZY7++bKLdNnAzmHULYnQV
eNvNvwOxtSRFFVQaVJ1571kvBZS1L0dTan2g4KMhDLUe+4pj9WSc1BjuPq0rtkuo
606/cKmlr9Zq++VNwvI7zZuA/QCKKq28/xNkXJZxS1hjV0LLEUo7yoPcEwD1hgUh
E43N3ooPNWAVf2dIbG3gtfzB1mf7b/40dKcSXXChvOIodFaPeyqtCm9eV0+ZDulQ
jiyrL7Ml+6DEBVIrft/tcCfJGQH+IWgH6Oeyz76Qg51NlkMOLlPHY68vQ8iiRXRL
kpyFucXRgiv5cp1BRZMyWWNVGY6cs7FQXNnEQTARYcCtmMMuOmifCFCuDQzh1f3K
Czr+BxuszbasgWQp01tS6B5jd8Ca6ew8SvZT08RchDezX0hV7ldJDg1qOd3rxnd+
kc/4EsI1K4qG1rKUy4w71voAqElxEN6X7FAj3H/dTZmd28iZFe5cQfD6n7HKvz6K
/zbz9xIvOgZRY6sIHl7w6Fti44kpzcvHrTMquQazFod124dLLMbMLjFDVa3DUVMm
2dkxMTEcqqZvLWoSE6oVwI2pEE82hbQtHEy8QxZ6thQUhCnxpTzmY4PCG+PJm/GA
0PZuAEoM1a63N3KDy6ha+3s2fy1rq5T8ijQi8K96Bvd94blXPcS8c3WnVpsY0J4l
KiRoDpirn0i9HQXloDtdVJvsUSdD3hrqaStgWkJ4Lw5b/4DFTny6A2qSj7OJJ3U2
UiRtFAlCdcBEjfMyKPIoSrJ/Kv2RUDH2EXSIv4LzYU5ArMCKtiR0Bk2NTKjEUVe4
xrQeiv4xK6P/7qt8p22vJ5DMCAPhGcdNvuafNGrGWjlqKh03fRfcKdataY8S9YEK
OzzdFVdVumzX+g19d4at4hBQ8Ja3ewLYSA9b0ueHzQKeDqKKGw3wweYEfyh3G+X8
WEqCkXJg3wVivjqWRxVZyvvnpKmrgzMorEippKtgNNBRx9WzMaCAdUaq5587nS6P
p9Pye1EBD3IpBnskannOl4URmijE+H7KJUqQaAH+RxQ4H7YXaJDo7ATVfoe2j59s
7OTquQq0d42LttZh8J3k2+WE2MKMUi4oE3GeRtEh0WRtU2iLxtQfwvOU3Bi5utyb
cPh8/HjPi1E3eRpuopy1PwaQGuMpbQ8W2dB156612gjGbarPFVZsWinhCb4r8jGO
S3ycqCmzcJb1BA0WaHnCa+NBdAqhRGkG/Gpmr+5K/EI3DJIiVsQpQHr01qEOW1kR
PyFlyVifQkcw5t8jqSfFlP1oPmadTYL2Bv9auhgWFjYKk/WJ/LUdmJHUa5XV5lyp
D6VIPIfPiYynOTnkYz7COUBDDs7/WAzM5RjubUkcsNTGZ9tHbjisYKi3z+GK+eoG
+v1/AEKSwQkNSWbh+OziuOXGoTu3f0mPB91DUiQDHwZshAK+JNilIi0ShdEehw82
X0L8Y14UcRq4HOIH64yqjj7FsIo2DGgRPw7k8u1w9IxqbsMQKoeeaaeRVzxB2qGV
QChkd3OzKguOtNF9zzZxoYpj9EQfCqCJwMlx77ndqzTQexnnf/cZJKOCcDBIo9Qd
1z8U8YO+C5HOtriDyISqTVaDYMTR/L4QYi2mVlv8iOwnZauo2tLwTU5vi32scQaB
Jgu1ZA4cKGwXVVaYldJjkbe7Y/KTDFyeiq3fAoDG/FEQD5BISs5Ja8exGR1Cg+UA
LP0+E824JyXvnXSq6S/OmcA6e9KgTfPJ4XJouYJhtUrYLmcKMLqoAQmgzYwLZE1/
FWVw0Cx1XOr3eGHS8Vu3wXH86wA7uHU7G7oZ+7fH8zMrIKaKW3nnH6HQm6HrYpGu
PmleXm8frrWfrH55nQ/fANnUJ0aLIi1b8gKN7e9QoAZdyrIRILOIpP/L7rLstzj0
cvM12rbVC18aR5HWMfuQDOljl5F4nFJR8O56YiVYwhggEX5mFgrJSHGAaJeBzNb5
keznXVb8JW3cw4tPs3cGH03ZC2IcpA7wks282bGQ4RvJkbLdasq0Wozy21m9Q0Zx
DcF+zOaolT9S0opAr/ISqplMFz4ZGw5cDR9priCMaA80Ro5PxSf9noawTOut7RaC
BSCntWJpbNpA2Gkebzd92B3YKubO+ziIx5rm3VyOo1dnM3+pbt1FHWNFc7dWLfdo
kQtXTb5YoW30zxgy830xduY5hmqHeQ+v+UJCXl4+N5h8G/Yb6J259nkMYnExh2Zu
fkSMAa+xHMLdReusZQhNISNP3sNejoYObvNB1mUel77wexG0NIX/BlElXdFZy4Mk
EaTQuPNaPHLL8D2DQCPgYqtl77hGW+uu4y6Zh9AALrnDZxmSOl38PbfYpvZ6sv7I
s5SuRAMCGcEsesiKuhGYBDsZTtoeEbOPQH5U0YP4J8ieDZ/glR1vWYFmdtDPgUUK
M+z4EIN8mXh6wgdf/8yQr5nXfrYI4OirAbAEjUb1Q1n8y4XleZgADpdLJptKGV3I
bmB1BmkdyjNhS7X8bqbr5eZxCdl5Aoosf2k0G2Gkzw/T5ykV0T8BLpkFOqCCaqBG
o7497niPshwlk+KWxNxOfkPSLv4E8MdF/9tU2pZmOLoeb8rfFjJexGxm7qjBr0c2
H+JsBt2dVEzD5fgDvqx16D4pxXgD71tDL+YF5LUNBSoUjSS5YSXdsayq+Zn0MeDF
JhfRPaJfdbUXQPgVQsCeyhsHO0oT0pBBM1zKajobaLC1hUG6OJ5Q0uDQcIFI05pJ
LVF2htp0jkjtpMaW7S+8aqS8QxBk4O4riTez3aNE/i/bXflnxDxo2CFIHFPkxzAl
RR9Kle12oHmGlpTOhif8eQVSp4huuWpQIxiKgEatqvUpjJVw18XhdFMTHOqfxnM2
d8+byK63duF3jXE1q0aKxgmVbAXRAHhVMmtyQ/tidoGVnvK5OrznVwTbJ4VHgYXd
tELXS88r4YpcPcstx6yIb0QtIlzEyd7XaLdFa47Vdt9KzSazPP1aLYxoOpizvoi5
UO0JC6yVGveOL5u8elFPteNP+EXzJvbH5OvJe8NFnk3NcxIuQzEexbgQSR4QLPvN
bMBZVdiiWKnCCH3CAFWhBj8dyNnc+Wzhi20eBoxzNvdmfRRr4arX9Hf1c6uodQf5
8oPH48qz0P7UetcwDZeTxFC/BSvKCcFGV6zTMqvAnvxQw5HNoDfPla0mmkoRRV+/
IMrt60BalW4ctqhmIiCd21qim8T2rBQVA33EmOW2tc1I4nlRHH5ZgKkeSrmS9wPi
6Wpv7BuTMkXgsqyJnjONOJXOHYcBy8+TEN9sDoEyVe3Bd5iL2sXWgSPc78Txpslx
diQekuNu1HcZ8fe1q/19+qVlXJYMacJytC+BXw+7dbYznihomeRk8TEr10riI7Qs
5iNB4Awk2bQS52y8pXIKV7QluCVvWaeJFg6W8raHRPCgPJf/S2q/BXaKb1Bpl1pA
AchOrgHUCqGx3hcVZ/cRVnhoE/PB04AxzvyUbObGf4hP7rAJ44kmE6lT3marbTPv
rZuOQkgjh40i2gFX1pF0IiXoiQXaOU8HVK3e1HQUQjd3bTEioE6iPpTJ3aaGapde
+aoa2gSbGRMZGfiCHyYvlKecR+hCTwh3ZY7rXqzADXdfSHaP+VTKsrI6jqiRveMk
O8vnLCMBd18MPzWX6MjQuon4bnOrg0HcSUgnUG1lFFge5HPCzsSsJbSOV5aE4h9I
R5DtysEinr1WWIXHr7DwyYzniqSJqCIZ2NKS96YTGlfCa6UhQKpTZWkx3xoT8JhP
uozhFtaFVKy3L+6lJOQL4UrjU11k2mlOP/LRgk5zwzRrJOkwRTzaxGfW5crTD3Bu
1FAtsxp+zsf6+ihyTErFRDR/PltMdZfj8nFF+jqF856yTdrNzDFGONXNRckeF0yq
32WLPvbGBo7lgK+g9Seq13OeJ4TRDfzFPr+KcEC+4nx+3etPSO41PDsSxoC6Z1Qg
pNsXMEE64SfnaBbeL9yOT91xa9uFc2mXyrHIhwGUaejwMO+fYCGRhYSxKXKeJYGR
NhgH7okS49RhMrMFX/P8v3qglCKpuW/QmzO8IpO3GXLBkuxxfsrJR3X/v8v1W3C8
Omz/YLBcDh4N/bw6Tex73O7aAngxeYom5L64JTuyfDnR4jWHrVFJhQcgIZogrqUc
WCB7gXLzVp+MctHIjO/yB4iuLL0Dw7T9TpCdBcWpkCtWPtwWyRzVdSGY2KlaKTbN
LUU3corj9h2v2gZPoF2d8cBrCytcnBMdmEsXaSzNBPQKbCtCyJFAmngZfNnQPqiH
BM6fCfZvxma3qNpz5GmwwuTNBELzI+pHTPM6schQMvyaWfuFJcR2I/8uiteeqrrm
inhJp+pIvesG48dtmFBxYs65wYeqvvrlDOU8t121ol1GC+SIF5p9sNeRUphQd2vg
jNhU/97Iio5JdHiI4Og4CTvWgubVSKFuAJ6lfQ4llZAQ2UstJP+mu3hA4pBGVaDv
7MZBCzDooHEDmTvPAHAu73+J0gtREe5GJAn6E02948ta2M6y136t9MtzqOEKR75Z
nla015IY1jv4YUUeDt1WNQdDPV10Ioft6HFE4M2cZir2K2ytHWHjAcJHBkML5QwV
ZBPIpt/g/ZbSfpDbJ+iY8Bf/aWPp3ujGjC1KbihhMCd8ggZhw/bLGAew/5y80JSw
yhp+eVPm9rvTsLAabgY0ZBVtFvr5wTp1d+1yl9iylYiTHC7jf9T19Pd/H15DE/9Q
Uj+gXPpzJqTm8qohx1QgThlQZCt+o4n+KYgKpXyUq4DMstIAPq7apAO9wH4gksLM
YyNt3xozMGruVb8CAABJhMbVVqM40I05o8F2GkZ0hKJPe7sGpxEJdnbqHZgYs3x4
BkNlXIxA5dfi8ua82E61vrwatbMtmwZ/dqcZgR5ptJ0sMZUIw+5AS7+xI1+jkNb6
2g/rbWkWuj0GaqdcimfL9Ak5VdQhsbwnTZejbz9kC0WT60zsBVj5L9UNluU6eIri
gMSUEsiXkp74FtxaHYzeBK2qij1yxuDvbB66BUtHgaN9V5FnTvqpeGNy0vUKAij/
IgqMPeO+hCW2RA+PnGr0zW35ysCee0mOpiunWmcU6y3L2hx6qUSKf4GafVKhWMDD
9cwP1eWrgUmX5tOsEvaLQ+03QDQNXp+VINlX8xKL1EDpfG/ycpALnpkXhm6qTrPK
XYAfy5Rd+/zOjdvcwy90DZhVaB4K/ItEB0dpuILLkdgE4GUvr+fBoqN7gf+NulM7
QzpY18nN5EHbN79WyfiQHWbxGN5j6JZY9r22AT89QnQSuU1KNBfxuDjzEJYDdvHZ
deUC7gLKnW7fOEAHrvQBHuO2/fwHt6CnO5XPoXgl9J6eEoDHoM5gkZKUICMZoFvB
THxSSwYo9TgOjMN8C6eJ53QtkAB4CrGBM8zLKtxGxKKPIg+8puCw3oaQGVpN0d5s
nL1cG6Mas3ShIkpsgYYBAgb0uamRP8kKWq/6RbsbsUISql0cv/s+vYEliVR1SjH7
pbyKwfL0jE3jOlfnnT0d+KqNH/HbQOdcNZNMp8h0SWHPbHhx+D240Tx1x5ACK05o
uHe8VvNNz/czA4Qk5I+BlQQBK6qocyHb8EjHQXbXYWJTqGvyMDIXDMLZnPtBVouF
esovwVRD0HQ/ARYGfTDa5JmGNV++cAG/lFDfKOi9Me7votkm9pJWUQ4pOqXaw5mC
i+Zud6zSNTFViTyH+8vddDbFpOiaIdKAMFT1Jc8d57ezRHgBFm7eciOdA2SfzCVA
k5pKr4GGaRFwkXWhyjyD3/e5r0MaaQ/BHM0+b1L3upzTyfYW7DP/MjqIQly5iyx5
EtaXTH98qJgvK9/Gyd4j3t2ldM5K24oakX+wpzS2M0SmWGsiXO+kwR5VN1utVwYw
amTsjnHi5MF21cqMLLC9hF7dNO4vN8k7+JdNtUSzi49A9fviQYKqX3ZXBcOJcW92
kxkBwfycrGisU9aAbIyF7eOVje+6xMCwQqpaCYfzhbUF71AP2Gilob1XStcd2X7o
Rsr8sPjKB9G6xK6HFUwqWAHdTY24vYRkhxnETVwZT2VWaimeNRv3xzZp8Q+sPbRe
E1OOpmaf6TFWU7bSPpbfFu2LM9XuNv8bvxO6yXQ3eqsRsxosY4vHCGscLJ+ciJKf
l/UAZTmw0i0TzUMSe/mHtdWhZAMoRpIvcb9/TILMTn2PRTPe84pxNCppLO5kSiCy
J9eaBSFau8d+jE3GD6mGrGP0c+AsBTBJhkoEd7I0o3yZhCOOAP10kZZlJ0cx3Z24
mGdJFgGhZl0JfuTCG1xqddzzFas0q1nIQntHC6NxjkWrEI4FzPVj5ZuqdzQTCHF4
gP73Fd9k1XOP0w3GDgzNLZeWBjeabEQhyyOsNJ5SID+5ejnUGC/teyOnZE1enw4a
Jd7vFCF4AuNQYj72cI9MB61jSFcbKT86jFyi4lE9mNwb67PVa+pCqpTTEnlWKAnI
6+H8gZZyIxdq6z7/Q0lQCdYozhtc9TYXftxQ5RW7XRS+FKz86EOuWHOg1Q7n78m2
+b6NA+a3ABdoqhL3G0mlATl9o2C8ay46pvRF2SH71DBHIjpsR2FpwJmN7PiKCvl9
hEQyXnKWKXCQW4ryXTQ6qxrQX7sQK3ecS9dpjyHbjvIP9yEodPUwAN1fbJA5U4DX
TKICkJ49VE7w+hXZNkgCYlVc1rlAz+fiRzAgTPMgiY0nu2jCqk8G91w31qBOwxE3
zgSIwXssGVSdtLridZEUk0QY2izVPJQjHgnUMhtF0lSfMeig+Fg04h1PTA683Mue
isxIPCQeC3fJ2LavC4Vt8V5AanDGKGf9VhddtadKXT9ZUZ4CM8ktfMFxTQ9iIT+C
qYCMHkyZIOysKYSDLm+Uif2TH9Ud1pjMFVNmc7uyieu1J021PSZxu6iSIJuB03DP
Pl0GWJykli0TKB0htuFnuUzsA6xlCqodpu9nW5gnVfnZSCoGLBp/Pfc/VvFkRucm
0SUIyVR/1AFEVoNG+E82RbL+W8wGyFU2AQ9PixQ62j8bR8cdYeYPvpDwMtdradHK
RoYEwB6lSa0RlRJJb7ZxCfOT89MFghJtidTyeP+sSkFNC63YYmUDh/djmj73t58X
syKkNi6jHuiIJsSmjGoE9K6a4FP5JvpN8MyyO6oh4bTjythBWB6QlxOyMkeSo5f0
Yfp5o/qdp2W6WCU56zXfMkBRp/0WdbXICPtVs4swkN6DvBVZKQpddx02bqUU4+6q
EouFHGsex/H/x2Jy0p6MIt7dCaE3/uhNQ1XozucZeuNCy6nQNV3NtJht0acVTTa1
FgXVr+lI1tpsdxBONZYwN1XO7aFpE+m/XuMx1xJJihLrZyGnGft4zxyaHaiPgPh3
SQTUyG2FjvRCEpwoY7Jj4JLw2GerP6LoSF5lHryYg6TAgn8yqvXJVO5tqlcQIeMW
vS9XTpackJ8QbVA7/qs36zW/HzsQAZO2pvtLCyBPwcoVAOWOu8+Kv5C/KM15PIR+
nrAGbP0rZLg1FczX1FFzsWikP9r37AOWk+iNp3eKySRH+WiPFVvT15EwQBGdtCUB
3apSo96oc3KkXsBwuSpWCQTlo2DyNuc4a9ggo5JaqsIGDLOe82zY7gGyCE+ks4Vl
KnwH9kBnVd7Ja6Hyo/T+qHIORv0kOL8vOtbgImigYa71QxRfU/QozDMVypBhxpsQ
/MRn93RUdFSGVyvlUGz2XTFzKLKKvSPI17nPi1rz4ro=
`protect END_PROTECTED
