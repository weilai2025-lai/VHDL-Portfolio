`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FHL9R56jIa6R7pWImu/M9WJLuG23ciT/biEsmWcZHwfYJ6egSzpUa1tdrkbgGLG
pSq3xe4ApaKG3wK3aMz4jSLf6WaPs7Go5bjzftZV8MB4jWKkfKastURNYZVTLgsg
yff+LmPNgRUZ1hTWaoRKHh/Cs7X5CPQKr404nDfi1PpFxofzuFPyAZT8KuWo2Edb
sAReKfhJKRNI65MqpzxV7plsXFM8R+WDuc7muk68KCS1erOADCpHt7xPHXMMjK/H
iFji9zK77hkOvixbf7Uo6PuN0a04igr/cToEH7YgXgLmAZCr7G80jJiZ3iYSNSdR
Zbx79QFDI2PDfDCThIJAVH3moSZtc52Vycw6L/C74SOz7mn4zh15RyUSSw2IqIZ2
ttCvL4s519VS5Mpdt1o661ziscrw9j9pWZw389Zz0uI7iNiTaQeiaqU7+cn6yE4A
gZu3ZBxAAPFei686BQwye6oH9nVGjC4sVW8Uzcpkm2DVbg8YfivIUmyOmW9RLCek
rKT5wQxlc362ENw+Po/+nIwa1ur17CEm2LuQ8iMwB3eIPZ39l2Ln0jE9i64A8aOK
keItXaSaDrJkOWEWuW1SLe9ZcP4hTaZ1Mrf1dqt2Sd2vvqZcccB10mvQ9OXGan4N
peyg0TZdU0E+4PLjEeUnGcgpfbPqI1MvZCpUVrynExIwyjjOLSL+dkAPdv0VrBf4
cUTgC4JRj7LXxCWkc+ITncBOLyEvYra/Tac23pX1BDAS1SWObw4miONgHEuvPxsf
j4kqN/Fxwy18NmFbT+/eA7aW6D7SmmiKotrdAHGen4UA8cQncHVCPyg6qupOAjgf
2HSzJeHeytqxtcJl2+reZ2eu0kBkmf4cBXT7VUiSixnpneofUWLXPeJMzx5jX7ko
pNNLDkTrDZ+ojiLyeTQQ23UN49tKNfb1ICLkLAqXKiWpYidcoQUsdYh37XLvPwqy
NpYsG/7+ZFfG15PYhMbU/Vhqsu3DpSZYRInuG6X43NfPuFUxu2EDIl4Hua1rPW91
m/v2hMIyWPYRLobp7ej2RBC+uA5YDcVUh22Z6fX/JJ2+mJI+zW0EpSLLX+DIQa6V
IZLzbRZpT7ceHhjDVKSVMyWMKgx3PoLZULnRtSib51z+R+KSyo/oiQB5WRjkSwtM
mCkjDpWsInCMFqxRoIp9dCFwZarR9/LU3LXNzi4ioxoA7wxiV6EwqIjdICEb8rKo
8LRoGUH16e6Ti6nX7InG+mnzYkh0IKJlo3Z3FjqygF/Q3S33Gc4HNBq51D2AERhL
YZaxqH42de8k24D8mwwsRmW6GH5+4gI/lgFucoC+kTH/rKYb4rWk7blYFBLGM8+2
t0acnhKhIswpA8OawXEJNXyizBxbp5FJIUIvjmsKVLNUTd2WtUmwZmQamfDxiWjJ
5UzJniWDNCno9F+gHCl97jQhdBjAw/lwOxAXSKg07XxCNv1oM2R4D5Q+Dh3oERsE
cvjM7KaqAMbOtSy2L45rZJTgsm4dExOb9WTVD4R8LOmwVzIcAuiLjmpyCtq9K7p6
BYZJzMzGtGULqw4dB6kZJ1NVcPqK+O199dALKvDPw2ZojSu+bIshWyfiXvtXPOWW
XnvOSfVdVKpUtzgyL0knWFh+gHT5S7fq+T9W00EDwt2Y8IO/CLiptXl6uQXbuEby
iDRJO6/ZVvVw0A5XXYvTzB9km6ixa4YIzBKYlnO3jAVTgNBdrIn9uoWcgB8EDww8
R5AKbTRrd8K9KRskRh/e/hnvj241KveEmcZj9iCM62wpulW+EthQvARJ6OLnqApS
`protect END_PROTECTED
