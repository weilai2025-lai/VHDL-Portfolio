`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKc/7Cwx1LWb5h5zg6v/M33KTCiNNQA3egfpSYp7M0VH3xxPhWl6w7TTq2olVf1n
eDl1NK8MQKl6JZ/BCUnDd6iWmljqW9XhipIKiTAwUamR+aVqU8QK/MLIpZzRMPh9
dgqkyZ9NG6CSOnSCjDkVYUSEt+5Ei8m18Ss/3jvteFonZeoAMaYoxMbmrNUrOJ+Z
e0O6rljy+3zcNhspsjvEVxPnecNlcPDIVoThlBlX3dM3iJaQjodtWbJJLpkjpBGu
0kCY7QK87kqfgyQF9R503NXxr4EtWVlBvlxBDaXrehShDRZKiWJxuNKbeFlWOsLr
tGkZCQuYY1fLX48sj+IQZ3WiroSzT07sUzwk6jOlvWpN4beHu6DJSfmErQ9Y5j6y
D2fzuIpq+8AhlRp2nmw9JpEVW7Y1EmuzUvjvu4Pu86rubr1qICO4WqZhTOlI+Aif
vtZO7+wSTsetAWX9n8bCFU8nI5nr/zTapjIN23lLGABKm2kCrsXaG5cOZfX9Zmfu
lsEhAEdP0ofFZqMY2tlq4Mvii6/XDUVa3ZRxC+zQ5uTD4cJQCiuKZ48NG9vwqtoS
l776Qzt/cCjrCVGCFNU2cFygOhvxPR05xiNiXzM6mLJbvmuXPcbmDwPPZreAB1RK
fN9J+6LQ0WaaJ+7M1kDGHZ16ZncEsFBEmRv8Z6U7kQxE5aqeIU/9y1bK5DXy/q3m
+Qg89uVkuAKWgcKPuEJeyXREzHM83gQxbfa+UWjYpbk=
`protect END_PROTECTED
