`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PcERSm6n+zBb/q2sH7lCb0h5xJ6XTBwS/4b258lBVW4tTjwqjVPcTKE638LGYV6U
jtAhm9/jxec+XXwJdgcmkqdkakIGn7ylEHglBR5FUd0CkltKQwsnhfqPLogQ5IPb
raqy4iOPJcu3vzvBvWM3nT6F/46MQUxRFbYWQdgni9c8rJvfdj1pUMqyf9uFcYVe
mKD1AZYZPh3lC6Z0sNc+dKHIM51SrwI+rQXLskUEHIKXxu934XtAHOBkW08KoOt6
BJSuxu/LQ+075pEJGJJVvGl84D1OK5u+aUzcP0F/t7/V+LGBc71Q747B69oSG6ok
y2wvqIDFv1ZA5QTE7LKt3wLts8tYcC+t/Fo7HMpVyAZRsLQKmvN1fm3dyv+n1EZl
bvHw7OC2VPY4rL7YBJG+us6dy+kSGPM/yp2iujiUAGfU09DlhyFtZCCKyGvNWZyk
fC7yE9O00aJ0AV4aRMCPqtIZCbnePTjL2XCXyCoqbw7NAvdbte1LIwg5GJRUvrtw
KwxxHNZaIApH/GfHC03c9IJba/aUS9vy0rBovBKf7eKleffwTDUlfpC6Zx4JcSrN
NgX9SLTKPL0UhXb5/Mp557ExXjCGfOweKkMxG9wMr28DOhx1BsTJgQT+5Bd0fvGd
ctBaml7khzH1L9AnkBzDl33nyIzJ1gH17sDRfeCOn/TDlXWb/yWobmwdlHvFuAvq
3nWnfYaEq+ZbVyrlHp0wT+wsYBffNMXHfsd4uGeQymCqxwJgz+cTrz9tIDpeyqqi
QzYp8BqyBbENrU2LgUFnuU1PJCKP7rBEkG54pHL7Uqwz4lw82OEZLjbNj4G2xYI2
+Cj9p1kQlltI3vEK1dw7ebjV3pRgY0oO0lNteskQ07geJi11coEv8ZuXODacdhY8
9EaN6auOXYMWOXBV03sa3x0lxxiYCSCEJyAAfYsl4ZzV3XxqLS7hIrGdJ2oZAV4e
cWKIdJrMeq14552YX5wlWlmqMmQI2FjtO4vuBcN5mQZZPHTkLJO1iY7CVtpv/1wG
rK5/FXj5DgJArIgmTIFxC6XTUmHemE/Nz/oSNAscNg2zIpUKJw/2cUUsh4UJyuXO
ir1ESyaFM28Eu1pROT/B3xWMfBp4XzwaeZ0H3CUk+fbRctLoslcTPHmM47sr2d9Z
USG6kom0oMtIDYCkhWu8qDIfuykVzgiXbdloM78195BG+bXQrHWDxP0KSBDv3tn0
qoeSmRXY4JUhyYb7Dk1GzncO24S9j8DRMEribN98moqmBtt0WlXbaJOCudBtwuLq
zM4sgdhUaAJ4rgKKleMuZU6Vc+IEwzL6lXftRsrHpy+nkqhXs9GTtdZL+RNnbyDe
PtsAy55FHqajDWvTmefmYVlQQhRV22hJ7iO/RVA2oka2SUsbbztWm/TP8EMPwvW2
HlsxuJeUIEJQcDAYzmgr6O+RyzbbzS9d1SiIbjDDaoV0oBZpUTk5nacY2gEdqUp5
QhfJI9mj6aqjUhxtAT3g0BEmcvnn6vd7UOXRHowcIJ8UNIEBN4YCqIK4gEENtlB4
rMUfNv9HAVpiafyUp30PWYmIfDvMQ1qqvuQ48Bt+V78pkBMvu2VtplMYRmJzZ85l
zG6F9ZuAzZVyu18PSfxI0kkW/UeIIXR0ep7CeugOXycMFmeRNkzBiOPaJ0p2o373
5ka3U7PAt6lol8IjSrysfNmZeDOJPqBh0+Pf1vnJDHaFxt5VYWjRHRn8n+yq46dX
N6yfHwcW+34lyPeuuJ5hDw==
`protect END_PROTECTED
