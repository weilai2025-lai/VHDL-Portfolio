`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHDiiNvumkvgDHVIuC3VzkuuINzqYAOGTkAiIFytXeMnVD+2VfzsvQLN6m8aUksM
c5V4KQEV5G+oo3qBzyOPIC//OyWRP12zqYVDudH+NOb50NGNv9u6f1zPxqTx0hFM
K93vHIMhe8I7Tk62KfOtgED4TuJNMZ5G3nC0YpnM/FYSKm0itncc8Urji4yI8dE2
hh9fRPTBBweddN3Xc4I0w4H+t0ZFaE9l6DUQhtqGfg7SqwQVSaVRV6GzWS13xHtS
aA1lUoF+x49H03oD8gm0CsQaKHrqayaHvOKx+x6EJ831d2oU/P4ihiAJzbH+P+Gn
oSaGa81ajrIOjDi2Mql/ArPFM7SkI0grLIl11nC7T4mPIgQGZiH9Oj5MuNzYzr+H
/gBikVgfEmiV/HyqL/M4Kn+XkQzMRUOCJAPxY/05ESB/eNxB3NAHwILIYa0FboTS
OEgtX5GR+RiacedwPxkpu6zCNqK8rB61ve8Bj3ZY/uGmEdL+Yz4279LuZY5vG7hj
H/Ts9lElF7f3LgCgGkS15PCOqn6otomcQY7vtTjTn/DC7NGc+YvIUdUXR9L+JvYf
o90R16su3pO/Rsl6KZjKFGD8S8nDpNi5XiZJ956dSA6UaeuibXKCoink4ppDbzJe
2cWAmi7fGjrGaywOFe4j6orrchP8irf3p/yqsiEg+6yfhXogicUSHiqObf8+UOBv
DisFK8RkKjzsSCuwTru8BJhlOrpqlxKGbpLsfgcpmm7fnlBcp+5yPtneH5JbNvC4
WwgljBM0bqF7ocGC0Jy6WL0HzTvE58Gq0gRnIEN3PM1tB6wcpE1P1HtPN0vIGFCz
3sQwZKlV3BATlwhsqM4uaa2XHRNSfvcDqpug2krnFLFep74SdKaOT38Lz6HuY3Ve
ZZVvt29l7PyxsPAF9hN31rqWMHVH3y6EstHtMQi46D/cATPix8t/cIcbU1mCHtLi
8hyxCgp2y0++TaeBsI8DwF3ejidZu7O2taKNuh0ODQQPLen+pUXBA2nF1U17Who0
fbscNwjr0I+dlQLNrtC84ODevAatqrQOZg77zg/52wZMuvwT9/7emxkSXtV7TSE2
CLFp/52ovhwEiXzUlREz4B/GWP2Cxkp1qfsg9j53kMsypT/mT3U2/LrMkSm6cK1g
C83mB4d344KFN+QoWoTTyYRe4ChWrG7E6HswYPiniVvoxDjVCTURJ0ecr8ZFuQT/
FkEIFlVe8hC7hfS3tKeKAl+iu1awUue/9Ul8k66FHug9Ipu+i1Utu7yKYUsqMO+B
m4OZGBzmV8nnD+0zFKjlWGI0dwSky2lkrql0/ONQT2VQD4qx4HDGL+Cj9GfFuyAH
Qgt65q3ZAFnLvmvHxn57OH7GRiG0eM+9AJr7hiazKT61KMPvP0Feojvr6bdiJHx9
V/FZlZBNWKCNCgdOBDRWB2sZUrndUzqn6WOsFQZgL8wsqcmuXv9AW4plHvb9sGGd
whkLNt1i8tyARTqdOfoLS14nzqKwBkT3FMgLchV6+0F7Z4/w1zVOKygJEFL3hqkr
F2QOQftRlwLK48HYP+5C5yLiJTJadieYNIUNtVYV3LwHMYIN1SXEySPjkdSm4aQI
nuyTnpaAhBwLiQQJaFXUzfl8S8pz/XC070RHCqqw712YwhOcOOWM1moTAl/eollf
PJ4lyVizFYfCulR+6MgA9H8EHYh6syG152dxp0kanNu1/04FK4ioFgDlEmoY5sMV
wIGLNtBCVrJ+Phnlgjb5f8tlofyUdklkTDvbBpA9AjIwkg4bF51mQ6E4jvX76xmX
0+zOnuwLcOqxmCOapLt0FGvQ1PAf7sGPbM0qV+05VJTUeFLmlwicRAmcAwnUEDzQ
dZTkSmemPeQ9N0kzZQAOpmY6pnlMJQfR+ubF+hNmx5sy97PnuCtHmn4r7SqHjpH4
F2GEDEq7HcpijmzgwgTrjIkbE2bMse/342dEHhaNnQVWe5bYG8gkI5NA3jZRMGvn
D9hiYDKhAwD6yaKU915Eu0PaMyQ1hk6l1J/QvLxoCDAzMmi8Kretnu38IazZH7TW
vjvAo2NTDUt8/Gm0uYwS8mtYS3ZcYlcUQvYV5iRy15jJ+2RdK3jmHUPAdu/XJfZF
qCSfLMnGkZ30WWlwPw/DlaVwCs5FNHcwze8qpUlWtWe4C/j/2fdrINjO1Ikt1ca2
Qlz5k6MNz0hPkV1JHonrH7H2+A2guRlzGFJdp5rkNjBPwsRC7dgwmoTtOyQRANah
+t0qJ3KaV0cIkuRK707ocEjioPquUno3+/gTPDWi4DMxAvSbaIWYth4mwKxd3iyv
BDHvowjZPPYfg9vC4F0jBxqZKIreVvBDelLG7tgpbr702ijR3iaDf0sCX3dqEvmV
HmhQYmS8sLeQ4DJ9vsu/Ghl1V0jI/XIhXGMKeGOfJubnULfo0CrX954W2t/E0+ru
PZ70E+5z7XBwSpbY1DHsl4pTVh8W3xFM6+Yf/BdyT3+rIm1hagbWY0B94+Z7gE3x
2GAJL2iaFeU+kvN7dF0tQXCsgVadaDZvNa3QsbZasH2ytYrKPmvMD3Vvri+RkFKv
DMtUzgy6c0Cp6GrZEmWi/r8At6jhVFvlbnYfLrAFZJS2oPsaYvSbz99sdXxJz1Dy
+Q/miWRPzoQXLsU06TlUaJt/ML9oZRrIvKYs0istelUniV0HzjgtdHN2/JJ6MmOa
uv4bLMX3F7HFhJjGHN/QWuCagSQchiR5Jz0+gM9Wy7s63oLEXZDMZTpxrTXdq7Pv
mT69b9G6evzd710gd575j97G9n0Vc60VXjfCFmmK6qYFZgZdU8HoKG+Oa2FHs/SD
lD3mCK3MKAHdqRpjfoRuzXi83flxqJFiheY9z/AaUYlfDaK6LPlmAC2JjkUGkBaz
kg5A8KyBJQq1LSRCYmqY7ZX84geFfxnvaTPS4PuWmRFifPWJ5M6C8b5Vbq3IeIa3
BK4eW8OTM/92rhIKCckO7BkBOFr/xplRf/CscFKuLNOEIiDG2/q7AJpyLZSvts56
iQVzg1ylg6J4QjMngdcF8F3RVfH17eePZY3HgmrLJGmhQABjC9NsdgWlKKvPgrBv
1CK1usl+59za1Kg4dhq1WQasT8G04E7gmBx5OoE9P6M3i4yGaxgWCXDI7Fuo2yFf
RVofETrhhY0FF/SLDbqESIKmlX8SO/ULTFHP8kx4Gsj+/evOV5YvHiCv5xhtyUuI
w3twgI5fm04en6zSeG5w6meAFlw+qYmkx4qEHR3CouToomvYBjcH1E+YrnUUD1UZ
PU6wo40CJVof+Zl4D6gkHZbFau1Ohltdd1xP5h0SFW7a1HDQil33s5vylLO+OWTR
UpAtKQGsPxnUkQDG/HJ5FN1hUwlxzTo2vaVdlgwsbhax65TGbZ1m8zq14MGW5kB/
dOT5osMG/XC0P2RgMqbjncXmw4wu91ASYM6BvrS3zNhp/DAJ66/aqEsPAD8L92UE
XGPiySJ//ULUOLY2TNhrKhbTyIq75WZyumhevqpeplm4Nx1AsCYlVvpvOuMqRjpQ
rMo8BdSGGb3RwpniVdFqVbk25qIVTy/lpHd0S6u6PmWKLRVrd9RRePpG8Zm2rGIt
x0Sexnsg8UQ8XrkcQp35sm6xVYcwIZdEJWiWknuPDWQ2LyZ0fUynnJCuzJl4DNzR
jaFY3J3c0Uz1XKKCFy1UZX6dkGhOQL2Tsz0FNaJcHdHh1WRPHNV8+bulXN1ZDMa8
gd6TH1/TNP8/U6NHiJX/0zlbFg5AAZIXJYhcQyh1Y+5XJqggoUavb8JAp12eSdC7
Rv1pjgG5wdtTA+qhmRuCpqvy6jLPJWtV9Iwr/1UzRHvm2uCz+KA36Ep6HBDxs7JY
zd6Lnd0IeVuLQq17sMtDjsC0SIhw7ezwaFmUtx9g73ufesP1J8s1kyqFdFzrNr6w
BNUhhC+ohCIaQah6lhP1Ywfx3t1f47SKd9Il848yQBNRB+TzP0nTZJ89BvgJq4cF
rRaOmYZHbjBFeoo/Z13xMS+m0OZXEhfvqmRxux2fSPqDmoIh3gu53A0l4lr9zJFi
Mofiv7BDBJshW1xVb6QQlU16vR9bl3HZZuh3MLlgIsxyKpQzZM6eZi3rxtSRyiSN
mjXyCPTedqnBLqxZSQA7D94fdKBo3EvGQaODmGiC0CVXONiYoxEeB5fXFF3Ug/rF
6qNlpHoAtxmy5uzkPiiv5jkAuj9fr/tj0yTKK3iqwxTe7MSmTYG89kcWbf4311G+
6JNhCgJCx+ungO7AUpdR+/zw8+1DHvgTVWA3ErZ26v1gaCrO4fMAGcAs5pmFFUQT
PgrhVtP1XlWQ/Dk3HHVfCgak27j2kwSD8QSeppECV7xddyItWiRtcn11gucLVUSi
Md6Naz3tgLiealamxtT9/Z7582UzgPRpl8F31shry92Mm2dqBKAC4tcwqpF5kWtU
SX7Ct5tCJDfkhTS6AtwaRnc+I674w0m0QIqo9R3JfYV32hnvWRCSwpI7N4wtzKSx
gak2m6kH02GwfQ07clgjtWv98tVDlJcZVOHJrKNLoBc5UkOdFOFfy+/a9BHd27+G
FY+JeHD6Dh+CBmLFH3pCBQ9GZMBW4M9m0p1TJhJJnq2B85Cqj3rt1YHhmdZFHFV6
GQVTxrywk3bnOqf19/NnHsylpA7o1SJ/5c/kmAKEZE3aUyZlP566Br2ZVxWHPmKK
XEtvtc/TiiBUOC8IGtmiJr5CTq/olCwTeajYqYnjKxTHZhotoutFxc5bTB4eGZEq
L3yserkWOIraaqnp2gDprVi/TnBLspoZVXXOUkeeBYKerpNKqgTPgx+7N4iuVvfu
CG7GuehFhZBfs2VajtMTvvIX6N9a4kQYbq8wpxsXJdX0MMB6e9rT5PVvUjOfqTjO
Y9B4jNA1dxyVMgERSCLSLvoJluxzY17kLkE5EidP7TGEBdv7dZ0MtBIT8ma9jHUN
oeT/tiOLkqyJgpZBdYw7XPr8zTy6fBMBz7Q3YOv2E+ZxH+YrxSGx/BLEp4yL46Bt
0zSxjl5FG8Xmg54HSMOZMooOb7mW4mQ+nHg1kRHVURN8CZQveTTFNS2MMKVdLNf3
4wrVuhW0Lq5tGyJJfnuLRzH0xPyWLwDdITzfyExGfuvDuh2zRUEFukjfC5uC6w8F
+ewBVCFiTxHBAOl7P+AQe9oFlu2/Dx6gozaOcF2DKO/+IV28ZZlS/yE95hqLjJxI
fWg00dZn95p0CEuKERAswRAHvc95sVBH1hPSAXCrrelLZZOvx57BLjMZE/asTNxm
3LCiTXX2g1/oFEr2+kees4nZRuZhxJbNVx64UEw4BZX4JhElmw/k+4KTGKJvszVk
5SYH7tAC7SIFSUyl7M5kUJvmTbbkOQV6AQIUzf6xB1q98BipxcdsWY/GZ+qsyXLi
AIPDC10LSOVuLzzNui7GD9cTaemfoD1WpP3Scb+LGZGtUyX/YHbgrQFYs1z1NR+J
xil3FB59iFSzzoPYjf96KQi/lsYwVbM8MJiZ23fhKIwjh9g4tAgitAOm/+ZOcIcV
yRcaLiJtsy3uDgUqF8P9BAD0jzRHMsXvmgjOhmQ1G33Ycfs+tzY4+5ejxeh7Asqf
pDWIIitFqPQ6TLcwmwI8xPXX7suqlxvECOLic3Yn/hS8TNiBwi2RzOqeT2mG9AY6
8bK3DVEKkErhMrPFWvlYyYFEBkYsOTnBmHfuzob/24a8qp1Rl4chDU0mvsTiShRZ
4q8YMXYV6Wm8phdS0e1P/+apGaG9Da5qLf5mjsKVDawRSuu4zJpKMtzTsh1vxnWL
uw3hSvj3p8ORNhd06n/gNoSuaxDslkv7sy08xF0Xcm/9SEnCYnfRWOmAqFeqdepJ
4+6oJWNbm0RUdYmIV9YAdNhvUHbGv99ahE61c30J8W8dx3fINfbfYEsyXNrT1XXh
a2QCESTlUPjkvirPQkFuJp/B2te4/Gzo7hf+NDcMIAvikUK9n4q7zoMHKtWaU1Tp
yNCUgka+NFg5Zuz6jgJdqVIQHxprsIOTB+sDdEgQTOvXnVPwL2I/gP8Ry/c79XMq
EGoKOEeiNCWlkjdTlFCsOXvlsw4MCfQEP77Qa2TFI3ZkqiKVBRnZYPCq57eBs0zJ
iSuBs/Q3WCm0YM37oMA/U3dzTuFCj4MZUAh7RoK6O1tjGObBKrotGoSVG2zv//DH
W0BeYaGhxutVzxb0q4XUJP1a2onIJHbkTeZ0I7GocDOUzuxUfc8JS3fUiZdBz7gn
nCRi3QdSZkcFK0CMRKEeHFMy03omG9o15Q4HpoRtNfXtvyWMLcHLVt1tR1A823dE
zxymxn8X5XERslnePxgbIArJ7nVzX3Wq9fgKCpcb/M3R3NSHwfsxQBRNda/zYpPr
FTHfShsPSxPvXkBkx/0TsqrIXOv9Qm0acpANglR75iOLNgNZfeyjKdGioPO3qDcl
Qu9lqlShCJg2uv7SxJ/4AVaTY6jsIqauPsOqvjGuTzUQinB/YdmffjUjW7M2i2BI
Jz2KZgv7JZHYpjLDHoqStQ/BAz6njMdfX4fyDnsYnPongfL/bQiLxQONkYdiRA4t
hO138akRWT8l3HPOBMbvIWYzmq5jrms6Hu6Mp9l/CxRrqtg+fiRTdx9q7oVc0PbP
WtveVQ1sCwd8CF7FjvmYcRibtgrfBxdxh4bYjMxqXcL37j+vj5/7428e1EO+EfsR
UAYqreou4AIPlxw8u/yTbnTXDF5YmFnB72O34H9qZ8GOmqlI8G2TawjkI8WCDtsR
xS0JSlX/CWckQnHn8JUD9r3a8XXc2N7MqvLUPY/fO7gJKIvqceNNiwJuLmpxo88Z
YAxMI1RrcVNTqpgjk2xTy/sBvbMWrTdAOtV2HAEJecAZnG8T7x/oWVghfZ+YgjZf
IBZ1d6koKeWQ2WqHEu1iCDP1S0DvcMtDyv4m4+wYSkPf+SwLgECG1QMVAzgXRsuA
TUOidVRAUxXReke8YGOu5HSquZCRwqq3DEJxQANl9LCIbEMbuIiZD4FVM9P8QQ3d
erCJOuvYhahkHqbNTGfMOjPdxUtVQUYbOuak0b/r/2SYN8b/BuEKLs1csZgdJOEJ
WsjcBEF515l7jLItd/ZMXLmRGHW26GIdQNk72my8KEFtpPjRt8FgTvDvKaVng6cC
XPGRduBA9/7NwYUa94exdOl9k4XNclt15fRJaTMX4On8CjdVYRWbIpWdjA9Dx5FW
uVs21I65W2BtU92xAJkkSAXuKHqibKN5nAmxO5TT9mYX3d9QsWAC8zg5X7AM7Hmf
ondNcNdaRRMUrr26eqrzAGP8IkyA6u25QxCAOH/NodY61EBRj8km6hxv+LTbCtC/
ijptlEOByHMhOgt6LaVHo31x+EZ9znLVhrt6o7ePzKO95DwzT+MfMaJ6ZQ9O3jUF
gkGWivdrxnP+C20zmDXxUePBamjLbhnPseq/Y1uTDdgVLTTmzO36aOIafgdLP5zb
s5rqSqH5cORJwMyXBQVu6e5hDV0EkWkYCBcbx44QdkxnWc+PgEDo8mvVSSvWv/Tb
FobXkVwo9OGcVAXIg1VsLmlITOTGTKSDoDM4DEzbvUpqzulDkqO2aAlXRkTN1T57
rSNk1tOYmLNYenCO2IW+MMbaY5YxCe8I4M/x+AgQUwFmXAP0Ts+SCcykiqsFi5p4
FSXeY3I6Kj2gZwFKbxAXwTMdZF1wHfgd1R8Kqwp5WKhvZhPzkO7yrZ3aZn3wMlBy
TY8Jvk7m7tFv5rn/cB7CL+ZxEb+grlX3uPL/R3DmzU1vCuk2fyNHyB5RO5AKRDDS
3qp6+M5Dl5BSbcA4TfgzFZcrDo6/hcclX0vaS23aKNQLrgE6vIRMaQ1unqn9fhg8
qz1DioGOiiM+4EKgQACKOv0rwOqiXzrlP0/XEUuqbmpDyHszUNCjw345jm0y8V7r
NcBAydDSIUkCEK4Gz5qT5Ib1B/vLkRSEB3rOxfm5P36LkRr9Ir/8urH8/92zAU/R
Ui+559fPc16mZ4usfXQT+ecBSDLIWgj0irRHuFdvX3Zfl2j45XRrER73GmHm+/6Y
z0GsmHLqhMEy8ykKkpOijxVYzJKR995IJO7Z3XAEG57q27EgcTmpZ5CcmgBbuBj8
DCfS5qmMfrt8hHtcKAJifA6F/eYPgKuKc4xZb6QmHbRsr0E4+ctS8E9M2r1YVKGZ
NZ51xA7xD7HxkzspF4uoWu3GAkb4gxFIBwSYRo0l24QFDpmdDbd0Lmr2x6mlgSBC
5zlGqz95wS5LN+HTN+8cGLIkLs71cuWBIxuAA28c7R21R2jcSUe2KKtEW+PcdPgS
bwsBAO3DWhrZhGlmnqo1lUuValndfJ1Ba7qSxkc56QkOvO2enKLXMQhvHwmrM57D
lUAW7lEefEi3izr/KWi67RpG0QQKthylzWKzKIcauWqhY1LPqfaebRDU4sRqbkGs
xBhnqruSLszulnH2WvAYYO1H/MRHouKLdGj83RVJLlB7BB7gOqANrIrXdDsRKiH0
8kWdyvldvY+eYyV/p/87uZLcC3zlXWnS7SRMmMnqMZ9Wum0OjsTdc2xmHV55t5nA
yIVbVWQxIMg/SKRnvP32F+SHyKYx9cZOR7CvwVZOq7cm+85FgmiNHNLk6l1Edxiw
9jP/LeAwAssewTP9xoPqlQwuC6b0zaNZG0Q2waDK9kNR/GlwFjtBdNI/TqRMDGWq
OgLR+//yRPWy/7OVr8znpRXWFCqbMrbsARarvPjzAM1GeZs1z5GRXiaSArINaPuM
nL5toRkTQFEzhZnOEo/PYu4DCu+rmHKOLlqr7KBxivdO2f/MKJSVgyZlFpMedKcE
QEL1SRlnj1gG1hupDvWlCpzHucdwM6H72SzIwIhQPFklwvGRWNoo2jnXdBHeMtqa
usy+ZjiL2yEinjIN21ArnAkcdWzqzYc/BVQqL6w5yTcoeqyuC4v5ZdqNN+b0wuLK
Iw6vAc0a0Ux/QFZSbkDpVS5KXXk35vxXV16f12HaeZx5wj2botr7+8aD95A0FTqw
qX6xl7vIUEbW5fHcNtzONjqq6ALRA0A6FJgSnk4WFpdC24DW5UFYT3pF9WNsEqTq
003MRdMQXqWmvbumgpLkDx3AzM1p50yTXkg2CTZuPgSwv5MgAbzSQwjEaEB4a5Wj
xOn8JntZnHZXxtV1yDGAL1CPP0A5aPLS3lBIlkyzePHhhqppBDzaSsYYHp7yCqtq
LyrxJXzd9NwFodI57XtVmTr2eYNFCBRPw9r2yRqQO63OASIkJeg0KM6qGJcrAVUl
uo08KLqblOxB5zeVd6pFRtHc6n/pojQbF4xHj8i/UmEOe0wBevpnABQq1QEusse8
xNL1cJGl7+GlV5IwM++ju3qfbh0J2eq8DO0jjIBafeK674qiML/gZkY9ciFU+9QK
+fL9d2OVbUArnMQZNAQJ+7RWjry52gRhe3rx8b8cqwtXSJVGTFNfpY1eTmpqg5HO
ZxgdzpeHUOkhGxOiJkpAjg0WBlRto2EC0/drfNYJF0lnKLVw96XHUerrhTpbq5HO
K+QCSA00blodKw/3COT/uFb+cmn69H2ZYz96GuThTDdrW3nYtWfEFInPUIuAA41l
eiliB50euwSh4wY1pNhxsBQyip0d2uR+yghJIqsz9g6+Lx03ihDgKFzZhtCk2b+x
N7lRFXwnamN7PpcACn7hmUfRWK170MXLzq0/vRmdjWM84YyNKY+lz8r9AXl7Oum9
j/r2NveQUxByysTnvM9SK/BckBkZCOoV7V5yM7p2of6Cg1QPySMxMiWPjTzArzhF
epyFNrJl1nkrHSAcy7/elvj6LiTUpEKNGCD5e+Xvp1If8jLkbHWc2smRgV7ti48K
dCkVErAjtLFx3K7zGEHnX2Ur3qDUU/CEETTBsqqEDZ4mtbWKCSfBlwE5KUjLAWUH
09ZYCBaY6bEqyxWyJqeXuUFr5OV49fVca/rPL2U60by8MChXnd5+/2sUP6F1VxvZ
ON+pmOToJzerLACFRT9odt7iql9pT2e/nqrpwe2sl7a3gk1J90vbvrLQlg8mJKG7
rZQwlz9R6D3ZVi2tDPshk2SNxHG5VJc0jW5vvVrWieY39+jBNHjQ/0i0ShxWOlR8
6F1EL+vUiI6w0lS+op+/e1CS51AoNBLKaiWuve1gF7WC0VKpum9eX+r9PpmGo1+U
PCbwGGhsJFXmvbPJsEYnqv1utPhcCBs/zq9n0WIvBrqut04qv9bvsk5Kwk8kwrop
XtjHuE1YqQTQV3zuMyy+xJNS1BqaD8cz1NLnka0NIhdACxNkg8zGwGnNkj4sdVNy
eb3DObQd0mefH7y6h/8bY+kssaJAwEcmiimO1WGADItkZROIMiCynlIMGW7Jcs4/
eirvKqT+22GSDHaDjOmext4cWlVy0w/WicBVfCGlY1F/8szudHNvUmSxcZbGfzIY
ZPR4zV+g1wPysk1dEQ4xcEvkaq442b5A+sNekm5RyYU70f2ZKeMtAgDWdaWiUxIL
vSxxXTPslnXH9cNZsarTQVb58Jc3EdX8OmGjUr8IGNVA6uJ2uJpLqUBEXQxPd2eB
U9SicZojLNpMEE1fMsqYPGdYGK4Qj1jtCgrMRz+UuGAeO2kv7g4cOn2FfUXxqsfY
m1Xmv89V9JYryv4oPKo8yBdcxgHC8AThxnWjJzVSJ7pHVs0vgJe2vHZBr7FRmepl
3XzbJ32Sb0y7ViG1xrxisYiDaEQ9IF8ycKaJeTZFJq8LdxOCWXLTWp6grVfmU1Dc
qp1Y6HqM7vyXb8eWcR0gpFlbXULpzF0WT9Sa2g2Dx7U8NUBKQgd8OM2FYcr7mOHU
5kQoxOUDxQ4wywRY+x+vvxZR0jyh0+43DV4u6/XE+uGDQuVHOhbsfgEL8jXwD9XT
nKpB6eW7+ZznSww6no3MdHh+S2OJH43q8F6zSF/ELYWnNqq67zopyjzGz09TWWL7
T0DJ24A/MbGGt5f5iV9aFvhxEItaisY2OmSQq16Ox0MQdout3oVi2fWKdai4UFDQ
flHbwwJHcOswaSGsY6IX0QTRPjUmSc2qa0/Tz2Bw33ZLj7EbXNybYrp+76u0zkub
H7NmYNSERKc8gp6t3t5d9SNdMYU4V8lCO4KjRneQFFLCLU1hQs9MXMsbgVg3Cvj8
ZehIV4n1WnlTwdOFADBosYaL1TrnyyFAxb7ENl7U5ptSrqEDpMzTgQo2ZAGdSj2L
PCi2tl/EuyCknLSBN2SEQW+ISyGiEZgfqf1HvKUzfGVgkGExZQcdFpbEH95JFuXC
8ObPqEzJTDqYieQBtBcRF2Kqa+bdGrlyGZxEpvuIny+jtjb+cU5wKDWgibN82w18
winWv2cjzAkzvrYfyM3Rmm0wSMFM2dE+j6W9Kv8DAbYixLlvoo0vBD4b/zO8lzWx
o5kfgBRynY7DSwllymTxsZ/z64l7G8yXyQCAoW+lI+uWBNBYkzyZoSXU6ajacJb+
nQEyMxVf/JOFUEkWZbtjvrln9cEw+AkAFl82///wNmlquJ294eUbmUP3EAYbJSnZ
cR/S3i/WJtke/BV24kWUKAAfwP8nH/4BVfMo7tSnZTzub0/kekMawuUhV9snTxA2
q7F/yt998gif0iaOHIesIHOnnOgAxy5gCLtGHod0GNwb9aDMYcYD3ZdMiSpTjUTm
k88kiRU7esDo85IoY0criJGjW9wRByz4gjHdtVzbkEZlebSd0zuO2RDb1R9d64TC
Fx8op/yqYnKs/eRl/MhPItyeueU8h7JIYawlKw810NcNRYTqrH+zsWkCPUWPM77G
zZZz1C2fBGRBACaTGvbYdqxDV0qfD7BfANw33PjETawIJ4EL03vj9Rv1wJarKp4H
AXZR8VbIrA4+VcDy/jVWAPYNj/7PCu8UTDvVgJSXbztjVf9xrYUafGN7oCskoPKP
+tNwi3yf2jut9EtbcbsBt1TKVl5giSt/pEEd5l7KDbZLM9/V+0+liMYIb8vL5BiT
hviWvapja77JsbXq9CMWugmUqfAoI3m0VMWEqpv+Qxi3nWp49fUi6+cTLhX0LTP4
LZXTAfBOPigkjsmlDsBod2Qsjx2nZGkJkc/9XRs2HV1H5uGiC2+vRUuOGb6Szau3
FfbvLlqRYpm2ECE6Vmh3rGbm5NV90OVi29zX/wX3PVZPFyJBoxrJhSzD9Dt8okky
wUdDMWJtaHJrRN6wuQz0N9Qwj6zxYDnjXSE2q2XcMSTYPuutnz45L6mqjDt9VYxc
M8LTLgXpGmGU8kDSdSB79q0xApzOdIJUXjSe/EW4CD8TvJsepftFhJhST3eAQmo0
X74LL2XLR1qqcvCx3pbT3FGFEcTY5+iZ71WJTF0rUwgWk+tWmB2yt9gA6tvaYT9E
nTW+ysmu+o/24wkkfIyt6GhbheJ/sZUNxP6GvTBIBa6S3cXzQpjqL0iJuTnembaK
KIz33L5rWxSK5qxjKSOLZ28XRcIDQkQmwpxQItdZhm3HuYLn33mDJeZJ9ZxRHFV5
y1eK1/ypOixhVYWhJtCRm7aSWpuVxgL3n5IBJqvLFRXmRfSbrbvpwYsJQzGHYMlD
ATf0i2M1IC1C22XvV8N9ZKNYgmqqBTLoJBygv01xERa0fYHB3F3dgK8ce41733Uv
JBtCRxdH6ZRdoJhcBLX813lkGtKZMBg0jjDcTNXTQCDgHKzVQy6s/vOWcFahvZmX
svj1zLRjq9KjhSstFm7TJESDqpbk8W0idWeK/vagWlLfqZY1eodAD8m3cO7PloSj
Hrvf+uoBDmjT/z65t2MLadbofg3Yhy+ZKoXAL/d4Ad0N4ptMsCpSkXXwqs/JfTBy
ldybkCJ8wlaQL6/yrGu0rMtdqhntGeVoZlFLrX9MsfZBVLbysaCOLnnaXMQQQ4wC
NHEUw6l/z3CY/t2ciBwBYnIpCz3aKTx+fSxEhs8W6N81+MTr/FYHg3ZvezmbDKgw
x3O3zIjg2Fjg89OiBHf90pjEDt7hfNqKJ+YaoFFqY7MYYsz6pUtbqVAGH1hZQQbh
+PcC/IeuGOTpH//zc5Kq1ZM09Jb27DAY70ezHHM0fUYXU24Vl+5NtRy9F7lOt+sX
QHoSh6mv7zda43dEPCdgNo6kIrd08t9E5ICy56rSyx0PG/jR7HJ6MZEPoL1dvdTS
ulk2LWs4q2WcvOJb3TEORRl5+oWqwzBUHMo2wzR2sW+f3sd3idFrunUiFB61VLn5
JKKg9IRt6GwH+Lbz9FTwISNBgj8R8H36qolVt+VRIFFNg+mcfr1vtm9NCR6TNyx9
AMMn/3rmLUlqZOyhvC5EzBLcgN/pga0+ROVc9xEvl/USwZNqzYP5hqdbQxKlpCu7
HmPLp6VKU5ndQuqg+aBgNxhuXL44o5rIQtuKBiUFYuG8gP9SGC7Ki8QYk8U8ym4X
kLZZTY7eviS9hrbAUQTmNTe1AixIjlFLRT+ryqy6sYE6WslShapSXZ45OYD+DLuW
myrCbMjPMb2W7/iEHq7ub0Xz/OvZyRDxxu5RXOFeo6CllNtgP8tqqEKgRxvNXmPO
I+gPKDIMXc7d6+DLuJJ0c++pG1N53awupORZav9Afwpk31jw8N6nQABrrgBFL2Sx
HTf3XgvXNVnt17Ysml/iJDzPHh3BbkbWlhFMevdi/L7A9QnGXaU17IJbGPYlxytV
o45O2x+/lJDWUW5ip//x6hRDxwzlC++WnSWXSs8XvLT0BNfiiMZhAuAeMMh2ul7Y
g9V4q0nFIkwTb43nGB+MExmKYt4aGWzh16GLMqM3kuj9MRAbLjxaXtAVaLyUe/mg
uFo3S7LvYVeCTT9Rb68xA89JkR41xQ7ZsE+A0FLYHrHdEzYW42AkrbqdtsZfkZdP
DVPJtSzoAKEjrehwol1qwRkhOiwFlCSSNmv6adWJv9uI6UdSYzpr1C+wxc/QDP4V
t1ouBG0I87r2JLnSygt2zl1fVVWfpV/s48NRhNfz0n725GhofLhpxpfFR0j8lmHo
jARyCnd2VuhRhrzmpAqVckD8cjrfj1LLUkRHMFzr9kUyyZEe7l1W6pGAx/wFMuaM
061BgGF0y/osKjF1RaQiWjcHB0XoK6wFESEfTcdcCMvE105T9V/Ape/SIHJMqz9/
FSQlg3aXCuqr2CPdkhcsP2i7unU8ekDE4thx/7zDGRQAp0VRoPq9xgl0O5tWvrVM
ZPL9cE9Aj9nXyIYt8wjYHgZF8eyVEMEfUpWNhHpbg4kp7IpTBdt87ieOl0HOokSh
g+Ht7So+ojWu4QDZ3rMXkL2LlXgbZHHIb4xGqPHKoWIgPkvwqgOx+uxqde6HzQ8L
dHbNYPsr447TxB1lNWOmFancv31LgN+piH3oz5bQIox1oXBwWTKGwgyPvxFiujrP
063vikV5LMnUPlsYAPbt2CMWboI3FcwbGoU8Bu5P5pQzOBnUt4Sbvxj5LOHBF4+c
KgwkT93WD0xIRh4titgHCK4avEjvQ8ULRI5ICVTvhVRU1knGug1RzY/k7FmY9ZcM
Sch9HsBqzdMiVghHOmT4c7eeIh8xID/P/X7soXIz9C3xDxkXLgEbYf6sl2fWYLWS
kvtRTwz5nH20pGlTGGXH/SxWCo/A1QQ/eQ5sCDNl7Kees8NWuoVdPEvyT7jtSCni
ivpHU6MzJriuEaXiIknBm1+ns+MQilM61bGVM8Aw3glOQPOVPfvPTQ+oRke2anfR
EoLuHlpAmlvLsBZhM3KSn8nb6dETeY7TbhF45+2zCozeNB5c3i+eCC3UaYfGh7eh
ZUCScB9quvZr36XnYs7I1rHW/Q23vt+i8LDADDEU++URnx8TazzPubHGaSE6CoV1
3W3XkF7jd4H+EkiJR2zEa6dGWdnsD68BEw43JYJxtixYjiy4hXn/9ba6RVMgqCVT
PyzHTqGUFarxy2NSIq+lQUMyk5hdacVqdUfHa7Q8ZFwwYnYlzNiNCPdXimpfYkBP
9XMCHRyZhLDPg9Pm7Rn+oUKeaduwKuEnyeAN+Qz0biRIdC8MxQiQYzMwdyueSJjy
4I0IdAzuuCYPTpywT6OxS58RAyjHv+ZS6J4tAIsXNtIzcMYoegcfq+M4RR1ng08d
nnAU0Ao4RCd8iaNgUdaQ4QgAI6LcnKZ/84rCN9fLZSVCTVjDCufCCYQer6o2MDQZ
jyCw/cB3GzuSlrlsvxGgHS6sb229qcFJ3zfNtLlnuZYT1jTikvkUv0gCwxJJCU6I
e1nTqT1+bxhWxvjNoLoqSaP4V5sV7FGHYnkow4RO4y4ARP93PhEt13UYdfvRG1YE
oxUzLaVV0u3cfK4vnjJxSTzYvEAkK5T0pqj7wuvjK/F2pNozTnLvy/ClZNi3ZvqM
GEAQjiZgHF4rUl5V0Ah+znuNDIMMBeALNyHhwr0Ap/WMiJ1kpzBH2vjPLvR8VvBq
6mV8L70holeGtKk3IikQuvCTKMVscCY2A2Sh4bzw2KjZZngXTztFQwg9v8FU4fCV
2FElN5Pm/CMgWduz/orD96p2wKe+Dy04HQptulOti34xhmHPBBH1U09u1W2Th+k5
1/mlUzdK9NuvBNc/pe8RgKqdvFRJS3Y1llx6fX0NfdLKipHBAnH6uvt4NaV+EN4n
DtZQTSzj7eXUxGdH7xBAhvhf3AfuXBVQeTcnxR3141fCMPfm2to+4nx8M3NulQhG
7Rss94lTlcAX0fnG8aIhtDtHzwlTXzCXALXgmsRlhIuPGGYNoYRPj1q6p38+sUIm
Z75P5N1SXxO3iXVdPsLRGX5i2HbZN+7gShsTcQENW290pqr+PdaTh0gFai3R0VfM
Xg4IiHS3pMmL6c8mOAu8QL82/7rc+sVoTDm8qNbyk+enaqWb2z230WvsRtq/4leE
hcKqdSHQW9zbnQ4zO7AgGRSDPDzHFFw/03va9QC9e/E7CAoC9vo8vqQww5ZwYPG1
9E+sDTvgzbVj8NUFVjOZCYz36dDdpc8ED0MzFHlBUUPggsiJ8D8WKdRm0vgI822c
n0mtuaXfWTYB4oRCgZ8hUouiZDnsEz1GbBgz/Y4lYR8t3x214J184DPhGgzRTXSJ
TKKfoNYLZH1nVKhry1/T4R4RoLqk/HMvSXDkjtXrJT8oy/ezAWim0exBirFad+eR
USvx93BbpwFVgNBh2drns6JnasQRfV1I6GJrj5vq7Nnh4tZNimdZoVnJ0S+WVR4n
NXd1OUpxDShz/+FqO4BcRYuToUxerm47jIe8Ad4XCnlNxU3Ub3u7ZNrPJj9aD5Va
wtQ40k/EPDv77I0NkseBfuuFjoEpyNtsdkwe2nluLMhEFU2Q2GQzHeT17dQL09na
vIGqNXE6s3QkKPovblPxeQYMJjKqXrTzxJDB1WlMWuCgHIgg+HX61s4AakmC7t0s
mnNrth+F2vlExLBJLMXGTj6vNt8znzqEWIy8h1q+CNEV+bAAiA7QMCwN08mT3dX7
11M7xkBN4puMJV4fYIuFJC5wtlQ49OefQV53PdEpSl5Jd/a9OlU71+Surw4XvWNR
zH9+FEppYilkUuwA106FS+NMFsUx7RUyf/W8SZt8oHVGM2l2xx3RXCQyC4O68I3n
iMhlnq1MnlDFPdCegNVGOiNmRJxmKAZWl0rpK8yOxDRlA+YR7Ls2FhCgf3LDSnO5
FZddoAxQjKiWAJ/I6mui+U6reD0PiDfmLfRtO9kRk4eOau+lRXXdvwcA4iCBXxkq
SN2Q0The5ZHy83bVjAzD8XWACoa6xrkQcZxlECrzteTm4qXHCjCImuwbf5UbJZ8n
Vyu1hdCPKNqoGYuHoHJXwHJl2Pzzjk2KPn9Sh1nT+nL6UB7rg2lL4TXF8icgS4HA
i9Bo6/WI81QItwJViEEB0LYi9gUu/TizS5Cxb7+vtAEpNrs0pp4yoxetm006E3OY
PZcgy3yqGJn361Jdjpq2cez9FBvumx75+2eBfu1Ovn1e4iR4zt+dEhV7O1RN8lC4
0uTLokYeZIKfFHHPJ7Ey0AOvw2dUKc9Iv+2PjWjm19BFJPP1lXzy1g9zYdty8E4Y
3k8N3CMENbHYTOmiwgpxnwGkATwwrR0BtlnYg/sD4iGTljRWqIyWfo4+WljBk3MI
I/MiZ8M06Et3aw/wDHduaQp3jabjwYSVtqzb8JhoApKXXbE2xdvayapgCASUBVZT
kbBMwgx80AmR5MN4UQ965C8chhVuCudlUz0iRCQhayrjqTaHsjp08g46LlUHQKid
3q4K3fou9psLKi7mw0pO9p0Cn7MWC23G4Asuk8WXuW4ZOMXMONhd2MI2GbEu3zq2
ASFI1QfPy44VWZjIRiDd2OyWIAfeqeHGsDllQJ9N2EFPxGewS+fpc73EtET/8ag5
jIMKNnHEqdX31njnW2BVgS9W6CYlOP/bkXowu211sdStDzSN0inDZTZhCP+dGz/q
ATVaGPRl43A9tHhTvVrz07WwlqSWSktAVYqGIcMsccm3wXOIMRjEFcq9GYS7jsYI
adDx2kg8kga0L6d8p/RYAAdEwWaPp3c/r345myjBFOOTsl72aaQAC/4V2QDLvXJF
J1hBtinERL3+9qPF2pZBvn79mYEGTfSXwJScWni2VfpzjH0HkGxY9A/y3sGzEN+c
2DRYmMDgclARMRlVDMx3tvQLSh/qGn9IA3BJIlOXD20mcHhep7UwGWvAcMwWtUL3
6sYY/JAKgSKLbwpYb3Rg64YL4hGcDyZsNMpPKNNVOGpdjp0lr8JZCQ8DPVu7z2gk
PZIUJFuXy6zhFun4qSzkf0yZd06FH5u4peOvSRpKfdMNAm6L5oHOk2QdmPP/gaPc
3ajJVxu2SIjKsug9eZu02Di4oTyUiB5+/DPJ93A0nXhc1Zm8UNCkM8Sb/5BTzyAr
WxcnVIOQ+i9ymiLKeBsdECSobugEVu+onuYwLrkN02lajMLx3QYJhQQlPzURSHww
RBstO1Tz46vYsjiOuFZkNt3/YeB7wXDb5s1PJdYnWJz+fSEJFQKYqDseYEABlgUX
CX5VaGbFLvcjYODQYp8m9HSA9pxGbOrH/lLOEPqFAi760c7gtpPakPNkUerBfVcm
IRDdFDHDl7WIS5k0nhLGnfWbusFbZV26aLNvNYNeJCbtZifj3cFmlovO7zBeLYwM
JfGQ1/tvvYHr7SZ01WoPIc+V+btjLoPRkN0YLVYq5wa7lXJF2N+bpkEN7vQSwOSd
LNKtCSOJJCeZhfh7N77iOEhXSRv/0H3sCnIQrQ6v4O49lywO/q9Ra7PQ6ZySdsXQ
43LR1Lb7rnVJzfflPQjc7hRN0i6M3GlNf/x+OzmsUVtfoiKLhk7jDKdxYr94zHwJ
lLVu/yOpSDgVUe2ZJ6S6Wj07ON7pmnY8kkClwBN/n7xmBcOTen0fz3t9Jp8CZTqT
q2X73746qbj027A2tulFqHFRqRTuiuaTx2vLjAR9ACPCHBv3an2NlqrHIru5BBjP
nZZw7hDiI1zQPADbVCctKIovLy+SP0baKmaHhA/1sBsgNUn8KtbfZPC3SdiAdEDo
thmHevR0cXj+HLAHUSRzGogXz/N0KDtIWT7h/hsIygLflBveJBWiXf4UL4UJaBGz
9QJi+yXAHQHsmgmOgcKiHXvIOgPBpLA7HrjgmdhzNbejHFqJ9Bu5uDjKXmbU7QqS
vvhfPXbI+I7WM8siSDezafYaMq/4VJep4JtLoz2feh+MN57GV/tR6lwAVr7RxSrY
TfWJ3PbmG7LsjvkD8WQknPmoyWF9bRGyUG9w+etORTf0+W6cQrRy48WGCky0ZEDI
KTfshLlTHAu6VDnwoFPOLuDry1F7C9V6YMIyHOs/F0YJOPaj8vfbqEDw5qDL7xGr
Kr6uFP72MuFm0s6qTKaXpO+hoJ/XA/yT6wI0hnZXTqln95AUa2fCrG9aBRkS0tG3
sCOoc+KEx5JQod48rgjT6r4ovQYNfeMia6VuGJ+SXoJMuheRHdlabpkgZSBnuguu
wiw9Vx0b4NxhASD51GSNNDmwLjH/TJqVt+0+leu9Eeda9tQWlbs8hhZ3XH7/EYqi
y4fcmAxmlAMLB/CY9laGSaRmo/OwiLflS4q9XPUcBvmik8Wdqqdoem+SeHeyPByp
r1msE6LVPcZyKtVh/6WcRKTmKmxgKvpaYj86sg1ztoVIn+JeEH9ocjCqxbqAczvB
8B6JIfsY00QMtVzoLQEvPjgSQgcUgHGO5MVqyCseNcSbHDC76FAGYlU0EJCejVrg
z8bISj4h4qZx4JiVkTwd7ZBfO505tamQ7AhVitKIdlhfnMEjBCKmls71WRYn25AT
EDVISPq75jkiYV+tZrqWnBFoHNj2XDiDTw6jo1kj2L/iNuaxBIFJNFE8MVSnBe2g
e/QmO6mjN3Yiya/GGul1GjfkOG8HFPAtBjK4nMzx+p8nIAPAueA3puZHdpDpJFH5
AbRCXRkUagrjr9I1xnwZ0Bln2oUAOK+iWYvORMRKUZaRXLPYsETNplgSIS1dIu2m
0Aay6zlOXNJ+HbJmYg+h3CAVJdCJt2EXvFU3y1+G0gbK3MRZMqkFvTeCSsXDgvav
IraqmpR0oXPQNwaOnlpDgzFVJBMgdO4h47KoP38kiIJiABVViyHMt7BAXjQgPKDs
IU+n9YCqCIhZUs6BUtfnQP0jnVtxfpgTbe47Ae1voi80R9keP8X7KY5psZd0e2CJ
El1teaVXvHGOGP1dtp9P0DmlWfPJiycXh8v8r4QivxtOCpcq3N3693+A12SXlqce
Cpw8D9kXQTVtR/1b925mmSc5WMkZRlF4bJ0NfQwtgQHT2q0GPZACdbmhmeEuwfbJ
DVKDl7oCKF2FSleRFmmK/L4fPsem7RBwzrQrLCKjR6eV/UOahziSp5kS54t9YEoO
bTjgPoM1+u2i/AG8CXkkNIj9t6di1vaggvBh1dGfBE/7tNd6apJIjGW6UB46C4BE
8yg1of7HmpuWD7iOYVHoPSH4JgzEv+9Wl7Gynt2vM4pCvSIes7fsaHdMT9evO87J
DGMfoCOpgtQOvPrHEP7H7lebdRflE7ThiePEHG12ut6P3moV0l5+camDYjBsc1aD
kVIRcM3lj4yLEBik831qtdSyPf+lPxhfb1OwvOLwpriKtQHbHRtE1tZ2qOuoqavI
6Qrl8aZpxS7IOFwDrNw/LGcTPfYmJWtA2563PQXgzmNi/23UqGjKtihl8bdhaNXT
rsPHkFaq9pKi23N8TTsU/UkhIN9AVYfxYvDBF9TuuyMtWmhtV+aLbI+54eFY26fY
mfO24i2qyM/t5i9bxIcvg36iaezKMRr4cCg5suuaYVYVJQnMzkV+FZgjj7Pa6exg
clXDRdSaK1i1GtCHTe+LErL0LVnd+q4fE5jUKILhw110A1/B/tnk3ahc3qHSDFlX
BMYEc0Jl4cM+6ZIiTNnOiK3SxgB27cJriYnP6E6F8jpERQZ45H9F1q+hDXnxOi/f
XBBGq6Hi/dJj1ZNQp/BlhsaHKG3Uj6CmmyDI6F58wu9404DMkfdQQU2lXT32wc5u
y38Y5rSxwPZXgrgmSZmhoFLhgAeX34pyI9UFuPFg/wrV6DOdSHdvNNycPPPMx2or
4U6Mdnnp/K0M5wL5q/APt6o0WHDd86jjAzhGfxPuZ23ixTXvnTOk/PZjy84LfLLJ
7gslL+t5Nt3jI0HZAAgK15POnk5a04E1W18OAnwIj19mu+YXauXdV3D1OncO+z8e
mA4skgQVXvMofzOsqxs99lIqt5AihZ91NbOKTiRCotV/aOvgX6n1hwplkdVIsF7Q
OSKPVCoPGdf6Ggc0pwGFP/aLRn6xlxiOGCXokn/zhgNLNF7UnT6mRH8/LVaZUb0d
gyA6GiIHZBFA6+u6LAwolxED0RP6eYzFvBAGZ5I6ZgrSQkg1opTRbA//GMmIwuKK
KRfTxW2Uworj/SFn7oBWGwtIR6HLhPZN8NqrzTUJh0j3kA7y9GJPCDHky1qWOQGm
NjIVhHnzaW4jZbtdUzLNCyiLeqmPD3YsjmnL2wxDOKpFiiEBkFgCrPgfKicndvkq
qIZcWYck4VS2Dnz72P2wpDyIcL3aUT1vIKb3MAQFEWeLoszw1IVaYuyyexJu+hLW
RiZAN0aod4aGDDe6lv44hVfmc6YDYV7SbNAE08TUrXY5404v+y5GMUU/YEtchhF/
ugaogZnNMZZ6cpKd0CNEY30sFxI7eLD37mmMvi6Dm2Nbm4HOmeYCLMQfCYK2xVF/
wRJb05mq5ZxvApjyywiPszVDPA+W2J93k5GOTwbhqUIvlJwjrPVPjneHM1ni6gam
OqZNFUTxJWWMZyANMZFID2U15LgAGIAhJgz7pmuBVVU=
`protect END_PROTECTED
