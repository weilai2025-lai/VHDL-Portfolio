`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YuD6Rk9XYZCIXO3DlKXv6Ljgn+TqKfp3yzSTV7NU19ibF7rr3uSpj4ZiZl/7/j4f
mlRfkiXKMT3fZ9kCkOBFtDEhyCXz2/y7pPFPBe2BSYRt8tIIQpm6mQDYNAlwBm0I
bqUWBaPHegNvaiA8DKCD+5XavtNwNpYCPpLcCZb0K0YLKLCLHRJZ3aI4yW/pr97o
GaHqNt6IPAGS3SVOUX1k+84ch1AjRRHy5AQ4Itkos2AurdnsNrHDMKhkYw3ijUMM
zZ2bt6i4cNMBsDYniMw4UDBAdyqp5eZItjoi+1/mshXG1Cqf4wD/E+C/dh58SlIj
TuMjzpz7UpRbmrmwbHOI1arEPGAICiZq1AF2pHfhYAjDb7QMdNW6grdWjwuiv5CN
zjx4+mEnm1U87B8CJ3bqaHK/hdrsXh8YCUDENuCgBu4TV5NswvR9lE6cxr+2pE5z
7VM8uK05o+SKxu5HBQbeapjgk6HXxIJ02J0bIvBHRbzrFNAEV0+5O+2GusslHeXj
OtkJ6/KV1FyUgS19GMw2cfnJRKQ+bsZuT+23BvRoHHtGNlAtZzqBp0SiP3R2Jhhq
pn3vRdv3if3iDZu/bq8A+4yUg+yVvFvitA5wIONC+87ylddJmE54kL0SNjB3gX0i
8iPbL4f13fasfLxBhYQt4Ub+qAPX19fRW0xEC+HTUqhH0BaPWXxS+MMc8uUXUZov
+2Dqj1eMe5LIeISYIZR5/4qZa1u7Umm99lqdFyAcqsHucQ5O4M26I+xuaY7ysppl
YA5aIJe/j4CyDE+zksOSDqK9Jm7bxD58VTw/aGENvWkAZsdjFhdNswzPiJFfT8iR
lEnN6enf7xdU3M4XVU7r7C3zQ8NE5rnzDcx7sQ5wrNpD730OdHg1Xv1yniVO5S70
fgae0R6BzBZgZRinS4uJr/EjuU2SBAqvOTc2TG5K+5DSvwSqBLtpLSyvhd/ifT+e
mQwpnbCCN+yTu7soPr3Q4YAsUIJedCbmVB1DEllMF94=
`protect END_PROTECTED
