`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cq3hvU3evRoGJrzEFxXOYsey4MCvuu9HpOYIAr4EZsyWSHzk8IR9uTN4Lp3YX+wi
bnUgzCM3jP1o6x343BXm5QhT681G3BUdoeSlOZvBtLMBLnc32ufP032IvmYHSHXd
f1qgDbOGxiUlnJXZtIYDILDztL2ObPPkESt5neUSI5s/sAeECgfq/vinPBKeyueN
/mS278mVspgkGZc8UNglIP97cBw2ngkPxqDpjcyWp76rdxrV89NdXJqVkBrxClm7
3dH4lfIIcoBFDCh2tF5WRhv4UltKcYJX3HpGTv/VgXBNeDaUMHWLhrrbzHnsZghQ
xGRLBHcZCueMpTYlRtbwY+w8EIaqM3VLxbjKJgB7sakXHAuwkc21YrnoTqg2ivas
PqCmuNgzpRWDIef1Bx4pQmnvPSxN+03zWzhuYZwtFpXE2iCTCoU1shjZQNrUqvpt
Bl3LDN8lgcdPGZ+3u2ITk58fbWcC8EoDAbB37zSAT7Cz3kDs4Yev1GogzmSE+6Q4
Mlq6zKof+L7Jrfql95zoDky4xxSNs2O7lMtONt7P2eQ3iNHXSNolHDk/nDOZJc1c
DH6/0pSX354WV4eMSaAdB80U+ywmMfE7NRdRo2fFECk2cJm8+zIQ7rIyF3CZqyFK
GsS+jdxYZwJmEEdtuWRKK/t99PGp2o98+Af8sj75Qb27i75N4rVAmpHYK/bJ3LfN
V+adNmEzVFRf/2tALarxPXx2miRs0T08CbhkaEvrOdZ7kDVHsyuQTKWiVLnTVNML
xB/23RzMcMzjArXJpy9hcXfknbvSxwhFZfeWA9Occ+GgH0xbeUJWbx6V79QSXfoo
Jhj+3NslehOHjqq7uCV26LtysJHU++SWLlxoVmyc9xp4z808lnE1Gcr4cF4xBDnA
neWD3D4qFu1UeX5P3XgTMbyIXgmBYichgZZ6q6aMm/fqKHnZVkL0Kx95qfTJwfV4
Q0mPILpxEbQL/EfC1/lnidkTmVdoS9nu0CXIpjy0lJeYBThk0coOwWqCWymsrd8y
e5/Teu5Hzb/FSCsZBfcUkoHkrzox5VfcgusM9aLAq1qAL1ub30GuP8gMVOhgAUwR
I9vszmkdiPEfbS5KLixrbiBTZDVG5UuCYG9zKeGEOgLp/ykPQFaJ8atn3j+FZk4o
MGZI0KfgkO6BTMNn8Hx44/7VbF4SkIZIEQMB+ja+rMl8TXQ5QiTRdHdJZjS9WOpw
iXyHebjpTdzpU+2WslmnI98jt1E3SJohrDoPVot4Ux3/0NdB+XZ0u21xK9v24L1P
uQhWpc08l+/hWXy4cGyc+S7Ng+AnzFrrgg+qL5iFN+BxggWuQm93toKsWN0uOKIY
wMf04+tgzULEaoHRn+nIF5lsIEmZ8LemBMEj6SKkAqmQ8o/Ie7YtE/zdqO0zphXe
Mo4yyRdvqfmQgoKBCh2jvu4mj+vURKpWfV6usy/3kbPa+FSgkIohNsYCeR2oQkjb
zHgD58mvt/FOZ/SPGsnbcjcX30Vl6LQ5adQbJ7QBHGGiHMFfqLDrKuGRKVJZUgYn
MTd1fIH4KsaMiW4V25YXSahWwQtTx+3JjGme8ksLJjUC7q0Y+hu/F0wiHJmToZmr
jFUcU8i6X0Jutto1DY1ryBxrYj6MihQ5i42cLO9v65xFvU8323Z5z+Cfv8Ob/w0l
uVm2dDKtyJZeLd8Xa/sLjLup2vRa8ZG5zL1kJ9sIcyY9awqfWRLzt7wrO3zAyWBe
Ga2WMALGQCRl9G/rIWvfThnTE9ghddgcwI6eDWNXE/+bzMQbnV0QxHntJG4HOEpY
Vsz7kp/LuTgswUkVXs0lRVmJTov1krguP6/C+XUI8Rst976oqrYlc/9gxVfxbtEZ
61AYK6XZj3Amny+07Xp0GYA3gtCgv5qonoYpsrkGbXLK93Qog/Uly50otY/p5jCj
RASh0+/ymGNerlr0+2+2agaLfFh2uEeb4XuXxw2B+cWSfTeDFAlBVI335BAUcZXu
sL8SOoUZc1g1R22b5euuSzZHCJQXt1ejMVx4+frbkMMIOdV5lC9YsQ+QNbXLg/w9
Pbm5GnPquYTEjDDSPZLSEgNE7EQ9l2hq4jsAtH8bFOqnZxzLRZIHw/7a42lcizIH
VxnfKdIyqBMpuZdDJuGDLmllVnmp1I1UPhB3eo3EbdaXwdvq3PUUHSp1/KUHFAH+
dy6A8nvUrJ4f/94UGYpan8DUypE0rIXNlw6eWdQnlM1mTwJ5QzJ7m8fOBFScsi1x
x7yIglnJ+lcZDuBjJlj7vHra1+cVe2DTD+5BLnECt/4UP90OxfculFP24ZuReAWJ
qsHN02kTy9OBswdXNBlsXnTOb/JoqkNRi2PNB0Ht/Uv0F1R2vKpm4B2JQC0C3L7Z
hyKHhT7J2TTytMN1ZOvx1zf/KDa1wwfDl+gsx/15Cqz/RwFyDC0QsXYNuxrcbD+R
TMdb13nIUjVYTwJ7OytlMPNyylHCZaKKTOjA/Wkam9EOpTC57u0JplqP/xX5Z9Qz
/Dxs+SuailcRBrQq6Cigc8lNEBJgXFOpJkCj7rWj+2MHg3Y8CWhFF2NEWxnSzvOd
nLokifXourNqvkO88i3r6lnIAM7eniuowA3QwbJ1EWbzC3Y/FQlA1/ZLtCmOC3ql
9CO74/RaZfvqwWmuW4aLJAm5erdIgeovpUyUfQ6IvFjsG2Ee+BHkZ3cgsYM3PxMD
7ozfp86k0B8XniY2WudxtDFufLogbLQ2cKc92ti/Xjd+lB6DATHFlytoDwPvkFcB
6jk2UjBAALCv4WyWS7gQFg==
`protect END_PROTECTED
