`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uwv6IgWenXTDYksmflz/oxX6JkOxq7upbCx294laG8pbG39yVKwj0lZsx84lcHye
ACxmtH/1ZEUQwxZ70JEMlgxdTwVGS2AFqjo4bEtTc+ElOmul3rkvfFWdSLcpl1/D
x84iNoUxdEIInbFAMzi3keWiCOY7tTc3Bekxi5LYLxYu2plCDwcSqXVLRqtQF6GL
PSW1RNYS+y2KLR18RjfZK5FVFqat+5VNQgyC3zcb37fFS0nNbjCrzMXZJ9aRk4bf
j7On49mP+qy5nX04l/yiLR7INSaCswgd0nzYPeHZSKCzbp+CsAQ5eCh1SZ5j4cO/
MQIMh/ZNRdzAXokfO3mRL44EUvPVee5wUU3oAzRM99FQ9uVDcn15HUGVPBL8Jfif
yAVnGfMEli9IHyBweHziMji0/zd8uWso8m7Kf/2Jcsp/hrS5fDEK87zedIB8oBlP
a9QLxpQUY7miYvcHVCHXPtyj0u8Cl1DAfU8eKkyiswyCv/22AACz6zDRL971xjvP
1a/eUHRBphP4sDYRZutIa/3/PvNGnp58uA30OE/QX4LkwfmjeFCGSVC0Txchccpg
AbI2RXLMyZorViok1KuH+UZy9NHLtM9qUqobaFu54DL4iDSLo/NCMKkMbn+frg6Y
jbdJcVuPlR+wAw59SFCKp225PqjXfmUWwOldyNjqs3dPLAciDakuG66hd1nR3Km/
VALGhhAEzYrfuKHgcmuTcodYFUDsm+5lKlR19GYsmYWDIAODk+XtOcbxSOS+f4bO
DUo4dfjTxoMlBMW5xNwoeVCOcUc3VIymTmnPJOdNvU3L0se0sHnGMDFlg6UpVos8
ECs9ErJiLesjl6UwIWXk+dwzxt0SaJOHy7UPUOo1DdJGzCewcKDRX9EeBvobOeLR
8iR1zqz+nI/mAZl/oFuyxEVD1e2tU6lMgIx4T17ATRfVV2eM8WSAEdDWX3SvzjaF
o8d4L744PaUWEZ7U3cVR/cVdSwx65/RrFtXntHbB6QK7FoKZ48HusYEgoffBj6Hk
GhDcHvq6A3bBP2mwnxArEw2xCAjRg82erpfnacDRGY2eQDQ1ueyYQvq4e+Ol0H5Y
W8A4ceXceVpnWUtvm0Cg8r9W5g32D3ErDTnSwRHRZ87sDzu56mugiCCPlwrF+Gzd
QKSudfy3bleh3s7lhYwX+wXc4JIgPuwe1wsspzb24PBk/RdFDZ10B/sf823R4+g7
q8RC4JKxwDoZ1MJr0G/YiFqm+NF8KEg7AvE1Az+IoNTehwoZMfIQQ88mcog6W2N8
ue2Xn0F+EJouqcoFEc8iDcTdnXGsEv98BSwdkANSB8MKJm+DzEP7z0c2EqLBlFhi
l7tL37HMS/k+hecgEw6hf5CFTkFk04rlvPCvUR7q4QV9ocb1HJjQnJ/U4j3E2ww6
y/vbfc3piUzGZ0z3h0rMSTZBAZATy0CL2ml/snMNplRWaNDlB55nZN5Cb+hFI+/9
8AwB9PeHolkjPMk9uWeEwXNtu2XO6mfcYeC0azvSxfaq975py3E+1icFJehQZoGp
2TElMzUIyifLNq+wbh117P0QNcOznV9PHqapn5L1rEmwBWMVtGrwF/KtOwYh5OP7
ykrvUcO1mfCMs28D5Y9tKb1MDew0HGPVYfjwIyiQUKPZxG+25NysfvlRTFrNCMIh
MAZ6hivlK0YyUTj9HfTCj2VLzXAoHff3Zk1ponjAuSKOilo7UzkiTD/3+qLcmgQh
Q4DKd6cKe8rFpljRi2ZAnTT2EKBq2vZXnLRej+QmT2ToCp8RALq2IhdAUKvww+nS
qEL/T1uVEyntKKcpupyKbLMIQQw4R2Ymd6NWUq5/d7uO+CqAQ2ql0v22Zy1iURxe
ghDdQedYsF2vAcCbsxYqRAlfNa57jGtLfkPAyneablg0iH85hcfKgEX422drkI25
szEf3EB2hxHO6hnbzHQf4M4IbstKcDW6WoH1zIfX111iQTSBcAa1CfS1HrsxdiOK
pjF26+t66uPLoNFfzMlpAcEfLNFuJuhgvsPrtzsSMa33+XqL2JQ6OhKJJ3gwjOl4
71T44wBAJsTt7u8svXt8eXaV70JaMdVt4R/tJoD4/YS2LFwSgAIHnCljmgJgetHz
Ays/PBI9OkCb+iRCs0AWZ44t8C+IwfMXbR4p09Qqp0+2sEu2o/18UCWxj8luqPsw
6JMbxIrbO4v4lHGfxgJYhAf04K1XDQRB4XMv0ZHc5GDMnIncVLVsHWfmWFSf1egw
3XboaDrhEVewE9sY9RMXeC+NTpt5Q7viQYw+jbwKWAYmh89QxU3SJuVFXgwTtpc7
rehgUUtsF/HH4IdjY/TK6xJdwO+pSqrLxQq8tReF6BoF/BQldAzwTjhv9CiUn5P5
0E4FfB1eWi6BdGxNH4MNKBx1i3T2B7Vkwk81x1R1kh+kCPLEuynZPT08avxZq5gI
4wMP3R9hi5Q7tuLJwSGUhNY25Mqppv3KpPnbBs9cnRthanj4FMFNsPwT04uk8DxI
xyoJdoJLRtHT48XgTKXLC7cxeHUT3+zqpvhbZra4q8dlr8lkIAnkzkQGLDDefOUt
Z0JUWtBquC5Zp/L6+uinl60VlwCVbgkkaV9CGafkEzMuOmDQKt02hwp/NEkmTVW4
F8eK37eBR8JtPCl9rIbQTxPjnDoKv4QpGiqaRLxxK+ZQvM8uQa9TeD+gtN0gfKlf
VKd5aWSJvXGNn6U6N9Xd8oUZPeydZCPjrajrtBRrNE8gOPxnwS/k+oU/cIu86oTU
ECZFkwptlZYnf8RAj8C816TQFwbPk6QhYGWHk1veXRQ69iSSAuXG0HJxGIvRR6qw
NH0JEvYr/4pba5cIUM2686mebiB3jQxZSWlGhIHlwd9VKMVcih2rTHjo1gBYZkLC
laZHLNPcWOPXQXXiR7J7AwvMQHIH4Itab5hxaVil64a2bAWQ7K2LBGYrVylxxL1f
Ahax3oNEUdDnro3NpIK3F7HdKD4smlk26LE6WB+mmCS6S8d5JRn+EA1NVNUyLQtJ
/JJz/e+Z5J2WdJjPJlOV8dZupnm9DKZ5T1delsO+IYN63YJLEMoMuxTSFs8f5Zxq
45neBhaBY3SLYR61sWt2JzY2vhBBmoPdh1wneRhGEM2sO2Kh+rKt6YCBsnfcgi/i
G54hSkShQOtKg8bJoCHBADGEb0vOvC8vJNN3aeId4TBlXDOj2gmEpNXWLDHg3V2Y
f74ARnI4YT9gtZNe46J9ldUkuklF05Ku+AhSxWKoOz+ji6spAg/lsv4uoHenbKot
kS/6yir8rM5w1Oi3R84YZGhI78x7IWWMLLjNdNPMbmmrXuvo2d8rJvn/dERDrgI9
iNEhBZizF1f/zY6Esjoht5DX4IMBjdNzrmsYoAIIeYIxksDPV6Mg1Bd1LNmxtHt5
yezVVEOz5ztSOOJKuUBzzoyK1KB9CGhmSZLmRrjyuydUezu8ZaTkhNPXNUX56Tio
eKbVny5FItYcaY9lh5XV6nSa+v3fpv46hwrJoqrEZK69xHHTF0bP1z7qYvlDaydj
oLS10TVLMRVwKkboNLDmIDjJZnoSiayVaXOPxeL8MLSSYJlatRSC4Spxwq2H1ari
xMwInAybLvjAYElCT8PjUDvftxwpV5n9Vz6pGFxTBYK45gwbi7ZnhLgUWc7/oXKM
/biD5/kWq9Upsc99hrDinFGClZm0DbYUL5hWnWlnyg8W2iWXzwj73v0FSmVhWo/7
+IiwV4Pa78OpLIWvctK+uz7Ds+vi8ebRpYChlgwp7mVFKsq/RpSm4wKDqw6mH3iU
LJ6sunl8hBEyZuCTJ4Z5tekzsw1W7Juil2yJADy+NvFlRZkJMrZxMo6AaQVqZFVF
Uf9Bph/uoJfv6sSGPB97br0ZG0cJ7R3kWnexePppjruPSzYM+FWdPngXT2D0q+Vd
UBrX0RPPRybRgh+54ZcxHbi28Y/EppnqfJIV5fq6hcKZUJSxVd7MIjaD/0/ELeAY
OK2hhaw9ZkFwn93BAt49LM0yfFqW0vbh80IJdJvqhRTBJrcIa2OmBRs09vSfcdR8
boO4HwY8ZgINZlRQW6tRdHaqQF7UEabwIdXo/yX9Vm1n/misVGA3ABGSAdX8d82e
GtNL1kqSZ7gau5OtVt2aCK09oD2NGUj/SOg3WWrEngqVvkSTyAmkkwkA/oeSdu9s
JIuVY+9wORX+hh2rcaQrMp5NZZ1fBbvjmYMYUUn54mEzcyl8yYL07YdHTzkfhn1t
UnU+6Mt/JeJZ7m2z6xBRmsDX9iw2WUifkcmzTOi/fZ+GVP73738mel3EGLQmyyM1
yms8ghaHfzLQByWXuXJntVNdYm2MFqJ/cWfqqj271qcxbpcrnjnd1ApJRTQc2OJp
FEGVC2JlMgbnTkXVF+QZyyRKRhDyj5P4M3qEYn/dxCUYkTN/Ctfoj21Iu1fUsNnt
n0uzIjmH68wD0Vwk1M8ktIdsB1NH8r9FcUCJLCWMQul6Mwz+lUSNE+wf8GKBpcn0
54JbAIiljqK9hrQz+lne/VtJ/ca6BzooezYZe/DI5etp6uZOOl/OSssl045/+Znv
JMnxeZftEjPsLy689SqJ0RseWamIfjs/XNvf/Odzl/gYd7yeqWI+cZyqoXBaVFTS
meJpDqsntaMM76vOQHV8QsXexZl+mBgI8DFKJ8I7iTwzyjqYG+G1qIrJ9Wvqo6Gy
M6tiwZdQUnP1PX1boYmAWRfrBPFFhI0D1L0Md/YdDHaRH/2jkgKTobcpvGtt39Vj
D7gBgA9SB6ws+dXX4bwSDh0oNslIYblyrOms6yQUWqfnagYlp8FlVacpof8n0Sfd
m7ZElALBlHhjw3MpkOC4Wt1lx65BHK8ppUMqMbP3dMyjWAge8E7SjDevb0d9l0ly
1J2XX0H3h8elDiLkdf/hh+nunBTGnkJ8xUz0BbnXBkPsMawd58ja2kojnt66oXzL
AZWx2M/QBZyk05jR6HKfFYDiB2rDMf2ECaHSfjAb5wO9AWvowq6RVcMfZkfW5wn/
lM9kKYEVg2dP9lF1KC68WY/ckGrOfQov4UAwE6IsELKT5htsYrJviRwV7RajFguL
1Wc44Uta0henpUKBtm07SCvHefDiKnhmuuPhpxnBXx6MrVBHhswD+r60Mf46bwZP
jTBzxnXD4UvfrkA7ct0+BPsoYUp2Bda+GbOdabBGGPWepyLrTxhOmc4B4br3rzE9
oq8aQpD35vjsF4oXmkBWAedM8ptF1u17/DVOA9zrawDJqgYMVjNH5e8aMSmVQ+NZ
s7PH65XMIOtn3qF707CJYAEHvwiq1D/MBsnZ/CdbTuL+r1TTwGk0XRw8nfSJtZAo
ILx9JRWFJ4h4XVRMUEmX1ApDP4NTBQmG6Hkt5PxoUmV0qDch158sZQuybFBtgo7+
WoW1omvAxaxG481YdzVmHdQWM8wVEVX1KaKS6KL2Pu75Lf5UrLnrrFeRaQWwRpwH
iRil0u4H00152IpucNeVF8U+OsQm0HB42a4QQIksbQ75E/JjYHATd5liD+Uh9hN7
Y6hOGmKALUDWhMjZ7bCw2+n/pfj7jviJEMTtFI6/S0tgrWr/bzCyJr81s13SAzW/
Yo+yyHZu46ogo2jgtPS/grmDk4/coLNnSNBp7Ut1hbz1nHYW8Q9ip/oZxTpDdrW0
gGLgXq5iBusz6IOv1/4SNhTIKbvu57kIzGTcFa+66zcIu8iboQEC1jHukXA82NwB
bVHGwrDjydN6F6lSSadgs/Sh1g1BXjPi9UWKplAknMFJMgInF8J0PMqhdg1QiSP5
drpaRmlX7LCObltFcIJTB5NFsHldohE3YKhDfGmo1TsYuNZO2eHqRKQDSjxibMH8
dgxniQiM/o9kPozGwpoWAV2vUn4EqfA/hxNNrT5Sn+K+8L5KOj4xRfAWjWZwISxT
+p0if6jHV0x6PdTfgdmGMAT+sr39BVEarGd2JYmIIRlAkS3i3Tv+MkRKnt9BP7Pi
3LayENwoPqlkKWdgZPz8H5JNG3L+SmRs2ZWReL6+u4UMcoSeLdga3BoRVXYlQZ9X
w7pB83NXBAUoL12eyXqKxRS9tDgGmLyM/91g+nb73Duj3ge5bwSKy3vh6yfP/sb9
ehnJNZdwWpSv6Bs3r9wi1C6KzVwDh3RUdQvoekPy0t1e6rCyWdWiMIJUrSae1+Lw
qpa7Fx41aAspr+ofaB9oL2lcVozgqJCZkrGfaYc1wrVRN6nuA1UEI7BU/tsGu07j
C+zshTPJZVMD60n2+8VRu0yD93b7oaxqHgIBdpHq5cGP4XXeW8gHnIldw6ANabqj
Og5y611iqioNLCiSEHAQ9wGedTrSODQG1VuJJWLnL8WQfISdKkeHR8ipURPtE6PT
uxGbb42cBCZU97yM6VB9wbeT7yL8fFoem9GwIto2yfrWtLF0YUf6Yy72Lu9HXQ/3
cKe6za3YIpEh8rq3RnioRQagBHSpofQvpR43L1imZ5c2vmU8PlsQJPwfKKPB7UU8
SJj4lVUJmlKLusqWP5vrdLgAa8jGDTVdVCu2uT+Htp2/HmSUNaygdA1D38rhZkaZ
cHVoytYnODm4VdlS1gRPiSe56jbU7NQzEoiUYBLcchg8//RGEwt7rfEX+iWsOe9G
gh0+cjDQ+0RE0nhhZ/kqldHjzw0XVMk7+qb7jxe5vo8qVqNt+E6hrlZJl2w4nbCQ
UR4N9+JFTj+ky7FJgxdzIC6CPBZq1lwoB9uw4DOjOgeaZHfRXFFwYmnii4SjRDO3
oR6dCl/XyAPjvSqFm2pJiY7KZJsNk/gV7N3cSgw2xfylu3W/XhLU7/haJmcY5y2b
QM0yOn5Ehi/n0IalqoCOz1JYBMfUyWQD8HjWJ+waCVRE0BBxrFHxkdS2kc8QHqC5
Ejjpi/Tm3zM3Sld6+JNKr/Mis9UrgLPpGOuKWqyxyOJpfOXsZejQJTi9o6ALZY2t
fyRwiJM07a6qQ+tyfy8RI5LZzVrEM+Emxx/78xhSAC5ngeEN3KhuPXhEvwBznhoj
IABiykGWFvSV3fMoe5+vJwH7z/WSJZwHenxrjZp7XLdSaf9XJKWhz9DY/wYDjLYM
cRV19lkyjtVoqYfDrGDbpcZuEdE0CAamzQwU1X9ivWcXUcXlkfPwvdUjp4GdKhR7
0HZdbjkoIpzGmAKFNeOOWieUF7p4kE/0yGDjn4ACgHiFTu2JDcmJdXAMjzUNUmF6
XMz0qmJiai+V8IvnJlcVctHlvUANcYjbLjkHLiszvkPqjigw6Wjr+02WPr7r4+UI
Afx2ac6i+/6eaF0lcCV3uV1CCH0XUGNQk8GJJnW70MoNkZRKePzZKCz1kN98KROq
Nx6TV/b7D2gN0T0SfHoZ1vEEKd/ucs2Mytr3io2hrGDgQUNp0LNd4xhd+x8KDNzr
nN2w1BPayfpnb8XoeZ+VNA1Uh2OKP4MC+rjxnseIuUZnPu/fpNNyDLBKKMD6cvqp
KnIx/4YpntIWJKykDi/Qz6+8FgyJHPKWZ4uIaUXs+uLC5mjZ7NfB941U6F4IYGlY
GQWnGS92YqRZuRnZzZlexXx1tzklXFmNHgObQeDrTgPuzOnsL02E0PLG1Agvt1u1
ux2xAQ6+oAwDYPrCrNmjcxDxeo+4ZlIbo+uvSHQjdILZ6zxIparv4Wj5kMJVWPNm
chmdn0vprawJtvU9wq/6kz25PXaxbnvNm+tuVmPUl14v8kR4Txxrx4K2CMRB/kqs
6RXss26oLUsVuGpMwxgKwPofPO+tBxRmj0QnS4N9k9YFFwqxTParF9bnFZtJtIho
y/9dlAk/cgS4FWnI1b6ZKoYepnvkEH2P0SKBfLBtGdnKnYf4dYkL5buNv/xxX5+z
cAG7zqKjPhDb1i883LVD52hrit8EYusQwyRXYMuupuee/mqg6wZjP4yEYS8CTdOl
0Zv+0ce8Nq9r3pOhIjs44QyoYoGR/en/H3AwDtKxU4f9TalkfHou66ZiutKqo+1o
FOMlR95h7ZhqoCPN3kMIO3fgNL2dE1eQA5EUjiHVQ2YRrYlKDToE28mnnh+C8xt2
f8vPxcrjDuhawrpW3+ivnxfwx/YP96ZU/wS3Y/yHNI4=
`protect END_PROTECTED
