`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNnM6hLKGJ9HF4El5t1WfkVbJD1y5sP9XOBSyD87te79NMq0Ws8iM7eTEXZ0MRuh
6vBi/SU9D5d0W9jcz95qGewoG6GitBkAzG70XwPWXJWJ3FYPh2UjGIta1cJtTjeO
qA1gQcyIv5kSYnq2lPK/dqHo+XmHKJ4ZKTNJz68oo+b2BZebPS8SxYiPXRThT+dd
bwfek7E3pWnWONroPxz/MHfk83su99GZmasIPhI2W0V/ggEtfK7G/9L/pRlmSKue
Ck1WPOtL1Yad6KSckIw25gUM7692cSNCK4rnsOaYT91heuntEuY4PdHP8Q9WbN9E
YEPQ+J7ZZ3qwyIw8oKpIHiNT4nAgCyw+j/sphlMj/Ql8TMkCGpQGfmQnMfRwj/XH
RVnTLKqfqahGzm/oiUjTCYvufbJpRF0ykNlouASedjcr/ie6QdUC28QNKEbztr35
VYsBSCe3CBkPapp98XUA5bs1S3rbwSt8nj6QnmSDa9eUVphuYlZEEt76nyjPot/i
Ix0Y/nzRCQPfEoCGs7N1NxD3JjaY3vYfiz5I4x6IFwb1a1voFhpVmRO1buZ8F7i5
dtixkNBKiYiwyTkP7uGY4GP3XV/dG6KHdfhRuc0M5/W4oN4Vx5q/sOVgQH8EG4lL
PaoGb7hHJ/LYZjs4FfWr3A0eLzEgg4y7IiFVAJ/0Cp1leDT5d0pUpq3R4dyscjJ0
WucFTwMmYVm/Nd6n9886yjeQVWIy5Jbmfwv+7xuN4faiDE1Lu9wMSTQ/VCJuCxhZ
zU1xHtPT8Wz1yhAfI/nm9ExkjmrEEBpYCmZPx1tilMWVIomfxRx7O5V0rcvvoVKb
`protect END_PROTECTED
