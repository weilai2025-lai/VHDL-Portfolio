`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PbXo48XaeaK8CePyut4fbBB+Bw6eRpRUKNgPD4tK6wqCjUzQ3GapEGeG1tv8Gaau
mYglHyD5pQxYsYQsd479e3kNXxC0caJOv74NHpbg9miyn1OHwcMJQrzkbayUZzB7
MLkuw4kOV6ErheOZk/ewy7xVYSx8B4edLnIO0gNtfOCpPzHMYQi1TAY2TGcZ1z6X
U8yTqI6d+vN/ONBr6BWvn5XWmEr+MbL6eZm2Epk2fGaCdHwBaozy3MDzsmGdmIEP
5/VLSVUIlpgN+P8vNVv87+ff1bXhFknGsyuQ9kEpei5+RVjBk5T/vrJPDFR9UlSy
OhOHrDMmsahEMkMOAK4NZ08l+bXQYKyg6NC30bvv9qth3NW+evCJnEskDcCQybqo
pCycc/v+x3bKtPV339OmwD/TU/h8CAlA2SRCpynBlsuSpgs3BQZaUkzRx35DLeUF
4P9ygV/hqX8j4Z9N6Cr3mGgjNVsgFQ1BEorSGUKQi8RyvTJepm7lKs5umpWNo2NX
NgnMNAjPDnFTUrpJv7nwx9iRgVgDSktT63mTiHupbBww6EjGOeYgTRtYC+JZ3sKI
LMK0HrDD8Q41cHT9pMB81A==
`protect END_PROTECTED
