library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity fulladd is
	port(a :in std_logic;
	     b :in std_logic;
		  cin :in std_logic;
		  g :out std_logic;
		  p :out std_logic;
		  s :out std_logic
		  );
end entity fulladd;

architecture gate of fulladd is
begin
	g <= a and b;
	p <= a or b;
	s <= a xor b xor cin;

end architecture gate;