`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVxRni5ET7uZ/n6X/MxB/uNxqVwwKwTpg8Q18/Q4GDVDnUe7oNFNURXKzkjqLScW
EiaLCrNXOGUYRT4ydbc/DVRFfgwblBxPnQK4PuiWfT8o4EeGEuazbJ0uCDDwO08v
L0OUnYeAFVn4tcYZJwPk3A9/Iysv60bnX6bja6pg1YVPxW2KMTKK2Gj0RItmvCjH
GnsRcsgajlsCzqWIgKeRmBYmsq6BWhqfPaplKSUdCM35ZqlFOgnqKSNMoeS0fFWW
GvEYloZJ5+F5EyPFBtvsj0PFKZcWnNwyBrCZaF8QyU1q9WY2AnHWJm1VkB1IDU2z
JY2M8/UwFGgw0qGmpNXMKI+jpvJTYYb5PPFDagGI7SNTGhcnqoH08s4nXjhZ/yDF
x2h2kaR62O1Iqy8/BkAFIClAsYi9KjB8jsDdwTOB0mrCp/Jy53bLE29OakNx42Zu
v7uDamzx5PM0zvbJgrQ2rOyW2cqHNXgke3sKUEw2vtOklTwISnf12YYpHm4GH7eA
R5PNmqpC57HRGDMxwP/dQ/FRsfkh3k2cmPNkTUHoMlo28E1qMMVtMWrF4MbeWiwj
0UQcLHovRYFQGATwX6H8BxbFHkxHCFxH5vUb14SvFXaVS4+YxDWho1GB9RT/7643
QftELw6sme7piI+BofHblmdoZj7sd8FniaiasgAjGRUtH/FLkYzcciysmDE3hUGO
Y9FDGVojmTg/Qi/55LM22WunS+oYW41bmpmH344T45MnHMDtJnXz6kl117+LstPs
VJkH7kJe8xt/CyM4sSI8ZCL/0j3l0DTmfhSsnJhy4mHKi+oks3aYJ25KVZEz/kVM
Q974nK80RnQ7ERcDV5FajQ3U5QZj/umwIEmDg8FRb3Ao7PukZVvB9tCV7u2Ft8bC
hVm+uLOxNjEHaJTH+phjJWHRBFndsodx9QgLlzMX04kGRtSjbpxjDVmznyECqGxv
`protect END_PROTECTED
