`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzdISuD1FgUYOrGAhIko1ID4YyUf4r96nQBCy6mF1u4i1efd3HAHPOL2uXHwdsTm
zcvKodaqrDkNgeg89hRWqlBEvZUXKBb5D3P51FieVpWE21hmIvnxYuA8+2Ca8ef7
tcyFE6bmNX9o2n5FmmavEgcAdZB/S3qpVs4va0n3IkiyGqUwvUm0TxBoeXbARzVo
tBAEjbLGsh9LL5Sk5l8XpBQuNiBMkCToVTpDpW/zRo6ohXePHzTpUDHqBpB+jZ1O
+zV2djnTWd+AePikkxcbCmE5OPJWWFXCmL+2Boka2YreDFZ9d6weBlMtDIg/EtvO
rKBvCENHw+9O1ywkJBz/bjcn57cOWzwagZRvEdG144yRqkFmxAzfCbCEAQYVQyjq
e3rer5wbcBoUCV91EA8rezEcvjGCZyN8JmQrY/4fi5slfCrbRRtK+vfBE/t5Dbit
zlMbns89VCd6WKQYYHlo+S9qzsCCq9262R8262HJwedmLGaKwRyn4bKny2lj+7Xd
iVXCrG4/2kMGImld3ylFfTBwxyV1d3GZJ1JxlvhQo2rGMdv2xM/KJXPBS0TO2Nc8
KGgcibPocghZV/9iTl9f4/dxc++J8GhhBqicrcyOjVQwQvWJcbXPMg3nLEiaG+i7
iJjoGrWRLhN6RfwpZ9IKFxYpzGjuL1IRq1AOPkeLzK5imazgC3vGQ6rKSu8KzqzS
T7RGSq8o2rbDrZ2JiSCH8JKdRhceKo3xs2lffJj7wxE3FjR3dQ3VC0jK3Ijt7H/q
JLw9hD9MZ24x8mh4YY7huijhA4mnt8aWgceC64l9VTIryXjvbOUDKqj9zywpiKTD
M7JQ96/mv4HyZ2U4Ia8omTdiGfGSWzAz3kG7YcBKtvVI63ti3rGIeeaSife2adgF
5YA5uSYBH5NNeBq+8SijlLt10HGiOOfyYyrNEIIBPh0KK7bI+UhaMTVtI6zJA2m9
T+J8k8/0lpA94orcOCjiggR1trs2iz1Ut3LkXefEA3iInUG74bOcboe8SiWr7dgH
gotrWvP2pVdrB/ZimTCxLdMcmPd8TGQdnqCwVVvv4haYK35eHPOpWzEYHe5k22jg
+JJzwdRZmKWN6xeKni3qPVCsBe4d+2oS6q1//oz8L6trkIvOh/lZX7hnvU9kQvHt
HZhksH17X3xLflHqQKyluIt4X1SL9dXkwloVLkIy9nvjtseIrBmPUVOkpfQcTmkd
Y4r4L+qakmXQV14YA3AtO/4C4T4fhoBxORhGJ0C/tnTnnsUnrCougl8vuV3Wms5+
kwB8fSESNaZL6mehDwO+7m1Ti9yqYcv8JvHOrdXnZcyNS+ETWGOyIPUiMwabrbyz
6img4jgTCv4qr47jQFIC7XoWxOVa0Way1f4ZNbCq01bqNYknEO2zm+MFiU3mRXfM
P9aFWO9ifNzGKHWi+pZ4eAkmsBHzYlM8bC6/9wEv7i+eEpW9oMaH4bPv+o3H2Dqo
JeXFB6RDdbNC0/R27Q0HPQ==
`protect END_PROTECTED
