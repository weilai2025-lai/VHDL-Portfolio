`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A5IlSuOaBrTc5nXB2KhdWqJAz8rmfiAa5VnSpyvTPc/88FEYS9rIILtkPISRNOI/
nBEeJhUf8WeqDVmNyxzckRQAVht+l/u+7+SyRtBbzj7ckagwJmrXUuIN1y7/ryd4
myu8a0SHCBo+qPWZneA5JpPkIa22RitJdx3lEG81zUOs2vpGf/+d/QFsMEU5y2+H
G9veOQclmcvB7Hr+5Dg3EwOC54i6lZQBJ4H1QqsnufMt6xCkf6VKsIv0DI1sCnnc
NsXxCOzfkhCHoo5EyMzfkMoHVJ06k3+pdkyx2X4IwXgULhbbSuJ5190UAc5cAumw
ROlVoqX4OacS/fqmQQwaF4gYdHu2Kp1cAHGMrMnorUzydN3nEcdI8EZ1RPmwbhUe
fgDmpJ/0p+GYlNBlSz9RO5kp6JbLMLp8/Mo1p7xOyTmiGSojpw3mI6HyjeyOO/bX
1NfS/OJDOxQwy839sNrCOmu7niFfHsEO6wDRaV3WxrthlqWTL8E7fi9ScCjWb2ve
JQEIq6ZAartqOZPCJ3nD1TUXfFixuZMNf+YrRyzgutoFFp1BlirUO2BxHiHgToyZ
4LAGqUkvL//BONpB9Sh2Y6jqZPoCe94EtCkz8uGpQd5dIY+k1uQ/5G/i4sKaEPc4
1y8CuLNNo2TMia5F8LwBsHXYcXDQA6wpaJVZfAi+SU8VJ4S1p6Yi348iYWuZALh3
CQP5LusNds981qty69CFLzK/0i5lcQjWjpJbSJeaZOEdv+sKrCWYfPOMj84VUSdx
evLmKYqbLbsHQ6Rsp9D3PA==
`protect END_PROTECTED
