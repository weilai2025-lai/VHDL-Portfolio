`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkZTiqkJWaI3bdK/SZAGTf+s5u6BqoLvDgqA0AFZZj3gRJLCS9uOFxp2cMIj6MUA
BTvxJRxN4nY4Ya+Ao9wbdohJtktgEZ6wj09IULGNBawfYGEVGRNcifnMXsmrUBU+
ujDn44o0Lqf2OQhevT55R/NnM5IxEiWLqJ0P2flcEyxk9zrdcuuazTj7IB74pvss
X4Mfrg13+axnL2zUyqZhI6JskVo95C+gKROWGKqbT3K+6fUDX9gRUajHNE/R9A6/
Sk5hjKHX4u/+wWtN8fOQxQqwalS3WJaNjh6xnsVJnwCSqMT73NfpF7M7pIbDdDcg
C8OeltRmh/LLHbF1iJS3ESTHKHQktcHYlmMFHMLpNybzb4AIzH+v2MtmYIjC6Xjl
TAicgZozj9tTg5+l/x+YgqdyXW4yfCYrr3AZD5QFi8MGzIhY9+ZZMQBQUW6ddA/r
TjXYkSuhWUhh47hxIMJRUb3nh3gYlLy5YfVXc5jknz47SfAPQ1WhB/GFa5WrilD1
MhgAwFUSYOYXltrGAkVqwknXnxbpXYXzcFq8RCvZyCDm7G/jzHKhpnn4qJ0/43BH
LHYnR6Cc08U5y4kpTm4tKkgbXM6O0CSOXUS+RpSqGlw+f1GjBsr25vgxhMD9J/0R
oPw2elDKLFYgy3YvGD5VFMx9pdsolHFBcFxOw8tZd9qmPSLwJHVQZS5Mani9d86z
e8LNbCjhNfoM1Oiq9DNa4lzjD0r2hvDgC/Bpe3ChrfHB3d0Icd0h8jIA1bSnEk1d
RXA8xbxAFfcQv3a28cNa4wGeZmHKB5MZqJfGizgTwRTg6XzY5dBLnvN7ieCCg4Kr
HfJP0PJ3DVaKF/YBM2f4nna2Ltj2PGVy/rtcnQSfpPm7705t9EGCc12mdnfvuNjO
2G5Yr6Ug3AlB0V/fBj+9S9NWwkm4nC4e7x6BjK59eKYc08BBSkMAMHEk/EjjyEPY
nhGpBUVA5SkxQcXD2W0FLD5MnqdO2MBGMEHfuyHJUVvqVnOvt9fZ/2fo4r0G/Uj8
9rQWurrMYUuvGKfYv+YCQm38dHnema3Jo+FSr0BfGHn6ZyyaVFxOKDBe3r8EsNqE
2ZPsNWX6i75h5sqb2svxGJmTgntaC2m7303ZB8R/jA773TNO/UVLQPE+heChuF7g
6H7272WEltMi3kJMtkVy+M2JB9L8pBhR2fQsISvnG4nscCqig9NixNRifXsY3Gu9
0hS0BtgnykQBHilTzpQflNVp4HHR6nW+ne8LHcnSiCOd2WKk7uCi3fVZpli29I1l
oow1wqDzD3IUt1jxScUKEDP3d3gQeOdABjwd7oo3cIqSKcilnYUpvZKxVUQPprd9
OG5JahsYCm05ZkChnFLvYIaEyFt9/e/H/bucbIvXDAB10kJfNE2Sd4ec1tlPrMJm
hZCDXrReYJcm5nfmx0KuFqgJ3EnQi0QEyX8nSQtzijh1cNUyt0OsZyUolmzBqt6I
0OyNIr3m8Phu6JdyYr3YfY074jdhojZi0tl+fdqRs9fhZiIHfUvtg18rX5+kLfhr
x/47CHwCfnVhUvQul7SwzKMj7w//N02yyRDfdpiSaq+W0gBDbpCK7YUGwY6w0IEy
jijx3dA1XKK3OD1NILhjgcZYWsj2GYzUT4sXHsgABnOXeKUJBGZ1rSWYnlbolGUM
JNjddOw368sJvvkUIe80neEHyvAcwc0fk2RKUbjL5RHs7CBWF0aTtbcr/LN+HbOy
2x1YRL2c5cEEg5qaGxTqlu8bPsYGc5qeXCF0JMlMNXeVMjC+RJJxZnNE6PhiDC3W
+c4O7vPRkh7bAvbmgPTne3om3nkvGb6IjrL5YBtM0umwYtg2/B5EXZL1JNt6Et5l
4NUpMQcQcUdWw+Cz2YgfviLg5ULpc0lStjbnJCWH7ZK+aH8+9g1Fw2YrSCVEf+iD
FiHUuM8Tzh39YvVLIflKZuqwifzcrMf/hW2UZCyo3bnPOzGKErkxeigGxxpnc0kj
iCnogc8M7068euAil8uypymxs+NMnYCj0DCJfCzuCXg4z6BS60r6NM6uWslK2Btb
sw2pF4RF7olmKKHQ7Pd+GKWloAjNuVjUcOwickdG4ZXy8tLoJHVb90Z9wyQEH52q
EqaaQELCjquwOMTLZgBi12FaKk//yGsRlAM41Ka0gw06cWsCuxptJGW7W8k9h/Bp
oNt5RVg0/U/h1SETWlZ6J0yD8LyCF3wIO7cWhD6XHf6crdjAa65o7GA6XhFD23HI
sw3ZY9WgP3wy/vPA74ggAkEgIt1WFTOUHpw0cvZKoaaMlnfSRuZ7aJHQo9x/1tJ+
0ALhFli29EdpUo6hXfrD6UFxZf0CRWdQ0hLYosYEbw9F7UaFqYUYcNc1zEDlgK8x
RuRfvAMp2SEhtgLwa11evlWehPGHE7+bAfawq+7gJVKUqFkmgMhLopU2TBxbt+qs
C3rS8PXQT85MnRC9+6/6nLWUY23525EvcqsrBEuYoHUVQ1Xzjd1UsTW0zqv8o+jN
yRC3Je5wXIsqWB/OJ+vaUlJWn8hYk3ZFYzGxbS3IW3yfPB8QA6STUI3uK2+8M1gu
8zNMm/Sizs3psjflP1v58Gpwk592KNYSMr1Mydw7W9+JPjhPUnchGIhhpEvKr/rC
Wa1x7NVoKh1JfwxXpYMQ4Qq0SnUf4hQXGLTOFdRoDdPVWlT5lQJAzoq2kbzRMYDl
mnBlZlOIsaFvzOZkNaPszZxLSNhNBpCpViczqjTkBP7kDwy8zgIytqIpU/+QWLnc
P0im+dKYrL5fQqLQ3bnAglloCrTvfU59qM8Z1ucFyrB02/UCPN4lff/B/UQqAl3E
hGrpluAB2Gnv9gojJOVk+v3OzEMrwTrwrc9ph9/s+Wzosf3nN/FXBHxxvxUr+eoK
Osi4NefUUccZVLHspPQXPzoW6tD7PRtZ4mMTYJJtctm7eFsRddu85POilYlzabgN
hwE8oMiXKYuGlWYRAesFDyDYv30hbnm5nuGbeyu7hPTJCr5S3Qkor5dK2Gox5rSr
/IBXd27kpxWdFStB+et9H19QSJNXmLedLtJlcoWEY4bnzFBAyKetnsZ221rC5Sd9
JHQBqq7kpA12Arb3yGRc31TiYJ/iQpLB5FvqlfahNvEnNGwxkZdNrtzEw7dBLF9f
RIHG0wV8r3kG1U6HX+8BYqiI8LbCmpin4XOVwgozPEC3m1AC4fsxXD/6+VdbE63V
OkAKt8pwGEPYBqnliFSjnH/F94GlA5r9tN+X7ZosUBqZJ4PF124IxpIRbzJNWvLk
Xz04GsJpeql+fmD6nX8fr4SzN5J27vxdVziQV5fxN6qA1f/KUZ6cSd+hJaPSHh17
RmAsEDfw+qR6z626Vmzx0AlMd/GNMmsGYZFd9RieMT+pMqLpPtfi/hIPMk8KsgJn
z7CBH4GYzNrNKb3i4NOptaHhW6z7T/ylDWL+S2T4UhvYe+ctt8GrMWy2ZWrJLhVy
uBx2R3N5O2D3speLCH1sd8nEa/FvYU+K4O/pq9GcnCDb7k5MEiEg4as/lty0aX39
6fV3i0N/RLo1LSiLmY0EUEniCaLxRLhCWxUPy4KTcGdU5UrunXasoRAGHwXSHOGW
cstO+rsGOIpy+614ZJsJj3QugD9upapIWiZx9tM/Q2k/tI2mJd4iLelwU4MOvKEz
wqg1PHJLyFQAWHy0aLfF1E46X4wXSbBVLbkuND7u4RfLcn5m54MrAdat52M5wwu4
0EJFooMxfheUud08KDYbBwzIaV8kRa2bU2uXb6broHygywo6sXf0TuLL2nVDz67x
ooxAgmPeU2kef9ewYqFe3KYhXo3da1z4CuwpSCMtF36A6fmmvcS/voTfuSsT3sqm
UK0UIgqLqRZwwbMlrSCUqhy1jB2cKvx6mPB10NZnBoIMzUhFCQxrpkIOpc/uQTW6
hgFxAiyAxIn+NSSk++DQFWMJHta/9TzrlT4ojqrm9nwB1EufnIeybve+3Lt6hxZw
QRxxqZF7EgTFWCfZBRZsKCGwn7a9fH5ubMHAQfTSoy3/ra1cfYiK1AIPfWSBj2cg
BMaWOdBuk8UfmeXY6qrvee+HB+heKMFaSDoaSIItDeJwJtT4kMo1JO1NfZNe5Hfy
GpiDZtw8D+zr4CB2dD2+HSQ5aEayyT+hvy7oh4V7+Dztp2OdbO5LRFfJ2vGQbNJy
wumVtv2KrvFXqTDzVSnE6LknJ0Q+lsTLXtkU+KIRQDKi3wggNDFv3noCMfi3L1u9
QD1hl3ZdN12hAcoBolL6jNQfyU2q+h5qnklL/8YnL/egRs1P6Vm5biQr8jDgyWxt
9dSNSit67IQDSzriAphtKZ1INAANzZM59mFx3XQQ2+SH7n2KsLMiWdmJNApfQH1a
514cEz56LsixQy4fDUZrYWVXnUKuQixpXftBHMQJbDD0kB9HTmkYkVoCwpxx+Orn
Txux0A7B3xZ8b2j5ef3eyAB8ZN5wf6ug3ozaG6eYW0+kEaGhljOnSsVJoyhSOb9D
mCTDqUlELSjXHxWzy1vn4UqxU5dShH+ogITYZGX6/rOxWn09uAJOL5e/C1MyS6w4
4gg4B32jVXxPTbgv17Vy3VBEuv0Z2zNMZ//Niym01Lykg/OTlSgDhKJ8G5wxj8kZ
xcB1RCUULtGtZcmMFnA4LX0yNRspVB7YXj0xQq1P6WarNoDjevYBxAWkh/zzVxtA
JxRqAg5ya0Gf8ZfteMWg+oeim68efy4NrMy9cbt6Ia1x5/AGrNhhC+9IgWSeOveA
bQzNkK1lJzUL5DXtukawS2kIsfKA4xG0NJDw0HIeI92Xg7rZBXbqcU5SPpU+RDrh
jmJZgXD2u1o7tebfcJu7wUxcmjTMs5qgMOpLf+5H2EaaVuK3luxK7UuismKfiqkP
VjlnsqhbTamswEx5E7RjLFmudl+FYmPLu7wD/yPDorcTE/x8wvgpfhk+BFgq9uCp
NqiOUduOqcVQ9UwG8p3mYBh74Hqp76kA9wDrkGg6QEfNiLGQoVdUK5uVyX+/h9+f
VXZ2lI2xfl64DIbYkvjuEK21qv+0/x52KaMIcND0swQzy1MJTcIp6D4HPlnt1QJe
1NVZTBL89MZfggv9VO0irj5xR1/0BXzR6b/AqiRyf57kIcmWiNheQ1TOoeeK5M2J
7hDnDE+sgFHY8hDsphYJed49S1wo3TWaJ4lz+wbIJidPRn/aGRFdmf3y9V8MiKW1
HyWCJY/PmWDFYzbu8HoW+IZiFOV85Kb8cqLxVaq7q+9bCzmMkYn4Hp/ISEYSJHBU
PFtXdIO+MLUhJdHLzAy4KJoaR7m1L5mQ//ialkGWV43UI0I9oZKrt0C1cfOPHSPp
cDVRBG1xqdsiQyk0PtGG29n4We5n/SEBXwSIOy55ZKr4wZsLp5gwxB0QeGm7zIHr
syw2YrViZpWvSPlAEjJTkKdyi4WdhIBdecwIlpRXxjPJSzpuuloPkX3fgiTIz1wr
FH9g1e2hm3LgGgI9QET4vxcNcsvVx6Mjr3KezgsHbtPaHr8YLOes8WJOMkD00ndB
505zuxqYPrPXPSJY5UutUynIkqZFFTulXI1WCV3Lufv5hbNTpNE6TYlwJdSzZ9Ln
W1Z/KUYHk7ZbcjmD9gxPoTNZKiSu0MGLbhyhAqcSsKMZnYbf/8tG/aByCCMLROoX
A6GwSE8zX51fgWhKtcFi12uii8ulJmXw7iwKgztwvyU/syIaQOZif10wUfb7eXFX
MjpT8x/suJjitRhcESe/RQqobizQXKNI5Jpwkm6PDnAnZMFKFzM2gC8rp/jCXM5P
lQiDyxxgqNNqIkA0YlEZ4yNRMVVVXxfxe+YpVUroKvqFnLARONxm8H5v6OVl3ix6
0Vu3t0KjygZVugicIWX/JScbPdplrgKD7dT8YbKjz68Cajo2YS02h+07+0qrqppc
RlcfYFtoVaRVRjn/9P/bnvIBlbwDZBClXHJuFFnN6OOWx5VKCQLRmgWRE2O/cola
b/9ocfTficodjHDk6GpuMELmPq5DAYiZiCmYNKnd9UiJzN4tQI+iV/+73YTUtKFU
cUkjOasXD0oGXxyI9b2PMQlqTqoEQ6Y5frMxvC8TQgtuYS4jl+NW7Qo42IEZcamt
yjgN6XT8OdbB9i/49cXfUJSI9jsUpzkOIe25fYnBZrQ/pNSz1xU8sP3jFBdDD0/0
/QzREp101NBDbHhQvGO4MRCQX5Gja3YdV89ztmfsQ6vK9IR44BcZrbJMhoHCqsL8
JIm3hwlGTYMDRehNfkzCEvzP++bu+T61HYe034ybW4g4furmorctsSI7v7jKaNI2
aBoqIGAXA+gKCsFA/e/4J1lgcvZ3DS/wS9lIX2TjQtu2BxQXCyXO9dUTfTeQ4QFO
+lF5e125/q5i0ogz0uRLfoqQCYjIJ9IgqEBOtnqWyvpJmW9YDuHp/+7ygVDv2uNe
ajCnMLjiNYnxm2/QVUYth2xVrHgTrhG29Q6nh/RgQFEy2s286dQztHLKiPan/nbh
F1CxR5oni04aqr56/mEm2bCFMfCIJIx9ChTSgcSaHMaqoahjSGoS0y6gIuRNXK78
9RfB/RnXpmFbfb2K5gRe7HTMxjeDSR+VaFcNGNqRZgrNFdsGsbyJec8BP9T04X/E
nmhxjrvG2WhRbVSH0iUE8IruqCnvECSb/mu+GplOrI9W2Un0D1nDKRq6wLT5pXgS
9pbgznF/MlWN7nxxOeJ6y5zx9DM8tdtsgHjPmoJkVeppLH97yPPcmCISawJPWyI4
u/Fqurm0hoOMmD27/BMcnaYm60HGeK8Sg11COHuWBegT2wAewe2EuM+Pg3Qac/hf
4u2l3A1hUNUyW0RkGeiR4OXMhmjW6ZoD8DXZ0wun3DwshTf5a+6Aq3cNNSQkTvGE
`protect END_PROTECTED
