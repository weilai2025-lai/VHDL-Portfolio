`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P82TNweCrZeK5tofOrga1Jn2dtDdMJs1A24HXvDPrxtWvWBTWS7x8kpn0RgyyQd8
5FYvQXFYF93Rw8WGAf+6Fhv4vnFb7PY4c1HmqDNH0AKS66PAQiFHAKWDGdaQjQfN
drBmNCA/2OHHQygR9LKGeqaVN+4T2RZdfgGnPzXJxgfpJZjGxfCGnYnsA9FW6J1R
S9O188VBSxPVY3SnEtCbnBQTTIDauD6ylxpf03dRDamk0b9REXB1ZZy3SjluYndY
n18H9wzqtSFJKkVSd+Q6X7CfnCQA+7d6BF45O00Nmj12n+fKQhT7aPH+vv9VJ2re
JKdrRW/eRL4TdqfqBqyd7eMgK2XJG7H5OoW2tG5s6Y9B+V8Wa6Ke5HaMBxllX3ZE
A6F8+on83SrE+S+fR71rQ+O/jZA20aFzGXmGNXakMNn6diJzhEpMF9gQjRV13upQ
LJaeeh+VfnewJqZu1JBRPxbBrlsU2DzcTBORclgqVEk3H3e/2MDxj03GWS3BSgLZ
jnql3HpG9iAsCrJwR/G5aiwjDO+HjPvdye/BUFwRgaOh1YNt8eOPhnlXsOW7y595
MkkCvTPRTqjPdTpLNiEJ4s7BHBB7RQHPirR++pweVXbE1zVPCLRLYOoVzKo26XuY
oebPTh4VEV5HMZJSi/sSgmjgCJlbGOG45xyb28xmWPofU4PMip7AjvupbVT1bPCD
ndDvSFgGZ5cBCN8si0WH0qbT3yYfVIc3ztNaBIjUNPSnZm2SPKTv1bibxN5TEdPk
2bdtZm9uwHH8yb6S5RKAsSab0AjYd22gIc+D8CKBpXXnmceTvh2G/6G1kue+6gAY
Qf26Rqi5RMgpRPeBit97zJ1OPQtLclnphiTg4VSKT6xFHKg2LQJBJkofGnOQfc36
gE88lAGWMiUkSrrd7SmVldTJ8IoS6wEawVtK4QEKrOvZTtmd1gqUPHsnPbbd80qp
EeUL6EbAmfgtPD1yxEg9X+J8c4QPGp8SkAcJbL6F4c5M2rsm1GiYZLJqlqvj6b15
bK3rE7yioqmwkJgDGIDKkHtNPMuFtfKukuc2pXnj4lVvnAr2962NwtAeh+qzpxfA
jpxBA0u1eUJOhOxAQSewyMNqtB0va9pU8Fj+YsWSXP5iQZc972EdY0FYJrxVyjpj
Fiw4AnOn+JO6QW/TAiuOKy3ZptDq72kr/2FqJEolN6pJ1IQ55LAy2fmDJ4nhwPX/
ZuFaTjjBohC1Gp16Dev/l6m1FknLEQMWrfbJkARar6Feyfs4NR44R2/92Vxarhzd
12Ki1xReXldudgtdqnq/WA==
`protect END_PROTECTED
