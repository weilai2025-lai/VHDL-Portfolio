`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljgCmmYMo7quaePyokH/10G5bBKbMJuAOYisjGU0Qdws73FbeeGAzf/rymr6DNtJ
kyauok7CcTNx0zVeyGYrJG6NYd/lvFoGOCAAcvxRzPlNNtcqksQ+juGmPxiXEpgP
61KOKAOtBv5vLi4A5fYokyFEJXM1hfq6OLq8VRH5m8hUVuMfnbQA2FNILw1bTakX
0svL5YM14IVRYCcBc0YCc+PwRas4H1vvp1muy9yIYs4k6MAW/nj8faJCb1qzd4bY
5uHpWwsB9U5VUSnMoEGfFhnvAn9ZozGOqKVwzI9kXYe0rCAygNayjk/6OiD3hUer
u5QJzPW8rUfx4pTLGNxZ1C20ENj/slz+XSiZPwSXjSwPm19b6Szf9nJJQ/nRWx6Z
/ancm5P3gGW6PXHZQrh/oEDUCZDn17VIy5UsWLfpeFMM02Oe2b10bpd5pbmkqdos
hSuXN7IlaZDNi17ocZu153VSK4gHNTGbQhxU+Em9O2rLU+LseU85BKM2Gh+fpKBI
NQWpXZstISZ6w0VJvLEMee/Nq0QWBnutG0qjVGch5x4d/+1wUwR5GIfH3mX9dwRL
iYoARBS+cvsHudtDbLCr/HHaqUOSkODaqHVMKTyRlRRMy1IQQgQNd9sUf4kAbFgx
do4G1vhhEi8QZZhG8lfi/AxRA4iqnxotTiGVc7PWvTPzmWvZt8V3y/N1mJvWPSx+
KTAE+mFrZ5UdcjKgsymGZY7v8xcVZpyiPUg8hD+Db3BtllwnxMDBgOcI5DW7aOUT
5JRIvfBO0OgegLSleBc/dEj10FgFWM//NipwZd8a1SZ4+b5OVIDAwZf/VfmZcl4Q
pY6tSiQGLmS2HkWp7WI2CqzWizIFuy9FWIys9aL0X7ERA9UFmCEGxV2LRdkOCZ3Z
TesbdKkWaJ62j1qobYrZ54dtZjcspdL4fpAC33CvlmP5iaeaWMnbwyDc4QTczIQl
AONJplovmOBAZmtJA4MooRvzX/PlqOBlUk+2BrjwR4YFOZN7tcasAMMwMaWTs7O6
Uk563O2q85TLt/zSPfiNH7ah0YPVUPfaqK+d+D4zrkhf7nfczDZzPUjVCAaSMxRj
vdRP0OyCOc0v2nGNMq/2GxfRlR0YdVLKS8tDbg/764PgQkVbzPnv7/hwzvbzD9E8
Yjb1dJa2Oeipl3QrznK9KeGQT33Fc0hP7nTWYpEHQD/9R7yJKbq+Ow3Fs5CnT3cg
`protect END_PROTECTED
