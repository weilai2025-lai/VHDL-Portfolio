`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pe5Ki3sqZHhmUywosHVN6jp54w8lboquTiS2wdQ0ov5q6YuH3lBr8qIaNVKCWg6a
XIqG0Sprlz7r/zdzM+95SVslc4BNefwtDMg3E6ZeUXgSummq9gG7G3Y805CcTIln
+9wqud3p01T2ig2CJpnRksao7FTs2hf1GprPI1lnabCINwVUHH9dkC8Ub5RIbYRO
6PlcKOAmnD8EtEDs56i2QkCkEXlEVRJM0HC4CjGG2skOk1ZMDt5jCJYCGZ67+E8V
SHpwu+EsG79HVvQEAJRIJH3R/lKvFs7xd30Ct3pYt3rwadc72J9u8SXVzGOc2aQw
6cPtOFfruB25mgITjhTRymoi/MkZ6m/QiTj3bNzJi7zE1HakxE4f85P4J0kxq4LD
8UMBV9RHK6a5UsfnrnU6GYSRlKfOm4nobuvppS7YxsjveaMoyi3JcQgt19yYMyHN
Xkn9Juw15U6Nl/ZM3L/vPigAdgMtcyfGHOqcWszpl1gUUcjzsqJYpb0HkQh6+rJa
/C+dwoJi5twUNXu3WPu4mcmHZvgu/vvbnmOk4L/wBaazOTvalY6EOEuyFKto9dnS
rzQoYr43Ytndnp3v7SMQGnKPk75s9leGOPqhymxgF4ym81Kk9h0BAZG/ci3HWBpJ
iGjQLyZsfZTgaR75QEUyGIXrLM9lz/wtHk/tv98BG/ArOz6MhpKhR4B56b13U3Md
AH9mJp04r/WuEDEQGZR4SKuUPgK26tMX9KWdlSkFp8Gy7B2f3CJOE63q/tI8SaOU
AlC/h2CfpX1BXiT4eGyi26TbYevReMVV0VQbr50DUI8GCi46tHXoEqW3FuCtgNdu
Bvm43k0sg+3qhI3oemUjsVea1u426rjiiGRZUHKP5ziLgdwhC+43Gru1xOkwqwN6
nF3W6LP69cHVbhTSsTEsXlp+gTzIFoAavOnoKt8kqqEGG3Y8PpvCEFH+hMB/ONWn
mAOLUJ/9/zbBDf+STMRlDAgeQNBt/4G6E3cz2cTFy2+FBuCpGXEzwlUz+yrRAN2+
PXxPUQIdozTuJEu7PMhRsLnoTTPtTIHn+v1ttBOLlx4mQKkqRXOZMvC7HNjCK6f+
JsWt29c8esMdd49vpJtYFxde6gLwbBKdG4nOm/ljX2bgyh8CnQXaAW85K4A64Jf2
n21ko+ClZLWR8+qsz1btULyUXQ5MyGy3R0xGghKZDX/N2IBkjydlLM97LBsAESqo
f/3lJfWKwJYHouCyPkP2siQBaX/ZbRRx9qgi6KQdTmIz9LZ5mL5wBgL1A6/yJZIk
AUmwfgEQQ09p+su5i5kCw6H8IS9RBUH4JcOrqX1ir7z3+qRNaflnHJ8IYALOeFFO
AYdsypFzAoew1/zY4k2W0nFpla6ew9cEEunLgXQcdDOtZg2uSMJTne6SNiGU1OyY
lMSfw9qFpkhXbg/Iv+zYQBslcCoyTk90qGzuC6pOJbnENxDg9Ihwk8odADmKT+fT
D2BU5Qjin7wbXCGyage02z5T9VOCWDiI7s8MU8w8DJTHBx4ceaPFsowWlsJGRm7t
iQu+tSNcgErn9NPBiOyGlAoEThJg7MqtB+8zaGcEpG7DMi5+ca7HGa5VNq5FrcSZ
4ReJpjjaPNZkjMs51YTVXE04VuyWCCk7F/ENe5jtYzXEbpqw+dXVDv4xTxoia/8S
S/Alt2fcZwjEYb3mFystan/O4q4lVxhB07QU/lsKInLRfI+m5/IaWuqzzm/eUo4c
Q6GD6xyFWxuFncaRHS+rS5RJPJt6zcL0R5jQIiKgh//DRLJ2q90TLbZwMXaOv9N0
H3t+jwiS4jrM7yndTkJYzQCpPcIDXg8HpD+UEnfRumSv3oKOjAoYsW6eJdZaMklq
f1rE73HlLsVdVFtkDJq0fQ0NOT2AcFllDlM8o8mADZS7Ejlsxg4h26pZUyT7ZSa4
4mjfeKHHvQKY7E7fSVfbHoHtNnKJPycGADUtqbwc5C0uV849+WHEsPEeUOsJ6ghX
HE5Byt5zAh5gPjVS4TyaAzQNIpWiLKuwIMO/Sf3DqrC1v11qTu43S6q7JmhMJN/H
lFZLaVeM+6mqx8wTOpK3zU4zTHHk+aj50HAU4fmh7XEhCogPHE9Gejoq/LLiPPYA
FC0Z5Wv/QcWzRXSo7HeWfjNmench+W5/MU4di9JplAy1E1kE1RgocetSEsyYXjjs
c0UcElh8nMUnYcWY7yuQy2lMcJsZvRu1aw5d5AzfZ8A1W7KUFVtAP5nGAzP/69J2
VUjqomX31EHBkuBA8xGi5WeFx2/1jodbOoiVRujmYHYxnHb6nvcQIyMMiIzL3CvA
SSWkvQUTBVzP6JiK6qWacNhUqpVOLCIE4qlkGsB1516tVtPnw9UiRlFzEnfiw8W9
3Oeoyz7AyKzdugTSZCeFDbu9UVLGMuW3ygflrqbjloCcoFhW5K5ilAfTAvqfcOvz
xgp+YZa4O773FomQwaL22RH2tngMovdHebV98LexJ7UxOiV8ledWl1tngbbh728N
fW/rGpNhQw2HYwfnTfoTuOyMjCTZLT6dcC90JkGigQU8CuVrA3/h63orqZnYaRsM
2qEJcJkfycUp49rm/2g0vnCfgoKMyvuQXIO4+363a4t2UMMbbGCUFDFW520afqT/
XowbjixzunjN2SF6W6jgdAycJqgi8Dj12pMf2WWX5FH3EjygZayrozPvFnz+vUF7
prW7xbcUlaFPSzk0kEHTED4Kyizcpeuwi4twZwVo5VDBG5tI5BZSBX/A2+npmYDe
2WpNuFeSiV+EnEb0zpQ8d7qfXpBreUx39IJXjlalnmWI535q3mDaigcw5bU3fEUA
p7PXAIOHBPvLuDy6JbbfRAtL4YnLghaRW38JQAdhlXbe3kGxr715MzQOK9z6C2r4
kj6ihQmZgRgpThh42PSfbN2jvIGzFQeK8dMvm6kUTSmYFNma78ocYLZvxOj2USfF
+vLTEdgoqKNG3PvAejN2VaJ8oElmLw9mYK1D2zvrJF5TbAsrvTSarzCz7ZNXpv9f
3MVRQSc8hPvVVEStE3SZhsDl/u3cYYAIIVWIw2lM0KM8EWyNtRJgGXs+BndRSf97
d1SU6w2MPpR+1HEKUaRfrQTP753/NyB2j0Tievs5KiUXJxvZdcles9XZ/r2eJFdo
gzIyg55Ypz25ndy+9KYwfkmdi63fKajm6rxJG+oeyz4lAqD5v6ob2iFfr+GMhOZR
6t8pZPuh1OyV3tQ9zglC4M+aHLqTNljK0xvkyEMsozj1PSegEJd0tCOz2Mz5yZ6W
TtxCmLiHrDwsl846luTTCL7aPfdGLw4p34+nhDVSGigySldTGnv91V9ODyjUURas
IA8h8KEp8F7zdKKu5Kbn5jos2efxJswPRLpWeiQPKquHe+T0ZD7r1DFeL4AxekjH
iOvytAyThopowmPjacH/7AGZdm/SwLzWvoBszriQOkk3uWYUFkzlkb6mwbPTX92q
vjjmfL0TNNmEmj4tXWjxWdZbRp6Ccu5AdUa3Iyn5dQmh+zHC9o8i+5tKDZPn1GWP
OgYnOa58/anN8G3QWN1gzNuYYjnARXDlrY7+9a5fQAakM9qKvIxBjRrvBeOMWatq
K48HqhJS+h4ScGvLnPRLnGL2+7/YUKZH66YUNfUe9Fcchqg7w7CAn3Mn05ElgmQB
AhQbjHNc4v3EdcaxVF3b0BWnrCe/MlcTwE7zJf+Va9ekjCmfUQI1MX8+/hQcOHzW
x1yq611swOh+M6rr7lc0XZO8Ks418RIejCClalEcNlgsL+uTK37+1cqBAv0PuJsT
clfXe4tUtdFBc8kujIJVjoTpHz9RJosUx/52vu+e4tjbCqaWTszEyfTOyqvv5Zxv
pnqV+kjYqXTXK352r5F48rk71UZdNJIohwgFkLxuT7lpVih4FCN8JEatCpgX6PQ6
wisVLGsiYkwx7v64K3KJFIf8+slwJEPbMTVIEbvvir61nuirPZfKXLx9zpSluT+K
NCcCJ9HphgkbN98nalQ9qE2uhdK3HGTmLuokGwN0DR3kMd/NBcTD+/5v+YVPtoBT
QmP+f/5hf64YZlMo21897gZP6S5HrAaoNGZs8TRfvCHHcJr4aK3OIVAd0g6A8kiV
1zXwXDxrbRxaWUVBdHbsFGeLHH5zWQDqOLc529F/M4InpVMhicTQ/PPUpndRcpOY
mmCbbXNwlf1/Vw1FedaQU1mNPd+7IQ9CH0A4R+3DrRlOzsHZSyagPMxyHO6xVCwZ
0jdaLWGa8VC+KKZ+07eDZLheFVlhzdvv7oQbfLcPIPFr9JD7SdJvHRLddysjq4M5
QIeYb6X4LIGdytC8aTECR7KOZDXuIb+kJDZzCvRDkrnMTd0Gso/siIETW8K1HZbw
1xO0YVYY/eaA4dnD9R1Mw1/9dJCSH2zuaTj/wAhohP/RRf+PT7xz3D/PB2h1E7r5
PFbX8xxxqgCU0FCWKUPuU5UTpeQXa0KbO8airZJfX50ru7qe1/vsXDho9r1vHX2r
Sk15+zVZoox/cQ/bd+j9SGZNyELF1uKw3SC6zYxeWKpHhEi3N9JQlxmhX3427c+A
r8PRM5iyQKPG3LMkI0FoRD/dIAC6vNeT/ZXSeyW0h7h1YaH9cZX+PVMxdGK/tl3n
eGzRuBSt7I7rVoTmGfj+tP3CSBYiVKQKwrW+cA3EIMhOII7u04dk6cy5v1A/Tro3
V3G5KwBsbRsCBY2ex8FV82gJzUAemBDEFZmTLRvtPRM+3G8JuyzCEjm6PpVmQl7L
3MHACuhIPB3j0HQRZxRDEU8Wod/ECV6JF9Xy4W8l+Y2zihCBMX0ahDPrLMOa4u/S
KURn4wysLSEP6nYqvWUC0ITtIq7A0ILvQlsCtvJ9GQRfM4V3DhSjwGzv//MkzILt
feGV4bSXPS+sManj9g7ubEnCgZv1bG6FBVk6RNduS7Sv/siQf8Ot3OVo0YlMggJY
psSqKC5CM25A49mSmYXe+ABUPmkQXruXkY2syb3VHovi1yiHk8iAQOWt6LHCDmMQ
fs5KoLQy638E3NeMRxl+f4PhtvmQK0apUjYLkqbTiyzwVAI4gfl22+yRb5+KEHKp
vq1wzaMFvlgK3W7GvxXkDARiNfGPjEf1j7RB3J6cNF9Uw0hjlIxApX27hHxjSB9Z
Un3bHMAGrO+5q7Jd33Hx5/8h+2+UDNSZIFxGyUgnwYb98aeBd/9CFmkU7BIdCG7c
uuxPClo88uSa5d5zuTGtvQlXwoTWxC1pLBmK1DQieRn7REczg0HWgbMeeGq56gKY
/kHvNtHZ5tY3My/sC+x0u1CCrRpUJuXPK3oZKU1YWEExu+agxHB+VIQ6e/6PkRqO
qUJR51YzdsdngyuH28YD8+PIn8xQXi6DuOuqxBsRFSL5ks69gJQtjpoMplovpz9g
h/szSDt7XQqZGqbzZXwAZXsE+Nxi7gJxcnRaavmeWVoUfxtudzkB5KVDQUMi3aAx
NoEO6vo5PIxQTJ/+md37mJPqxMqKpy9ldPKSByJM081a0wwy9Jg8gONQ9AijCMjX
qaLsvJzMOJzmPsEcXEWq+eLGJCC6+XU2EUX0wljU1aUBNLUefZhA1zVsg7huBkPa
6OQkSM9cVKvmExFAUI31krU1+fzO7hizWyXuAIG3+tLzCz/yeVub+kGTD1/CkljL
lXaceGiZTM/LiK6JV9J68IaY/tEwUylDKoO7waHjtmkyyzWdlmPvkdufVD3IZv/1
EYUJ9t3DRyZbvrxz82D9Kzap9MXbWO2ZR13uXgXsCFLCzFdZtMUwMMESVAbQ+2Tf
zDMpT4s+b8pcOvFsL9knhvAn/DDaeVBp57lbNH5Ojk/SqB10eQMW8SLdVV2L70Pg
JFKij97NtyPT2l33Kej6RQghPeVReYmKUIVzCgYL73qtShZVo/v4/LtzHxkvu35X
MBJxvpg8qCUc7etZIG9H0gttzA7rJlbdMP9e62PTjLixDkSM5RQFIpvb2DeLv++z
jmeOC1kk1n1LpYdaqQvx1G/Y4jDrQqjHAoUXyB7YH/wPcPNiz2Z4Fd3aUzgZmzpf
AlR7N3hm6x3sFyeOOdqgFxllogfpyg0XoFo8a96QKQC02dG/R8/Ph7MOtfoGFAPf
IV8UgjkGLj5rMuvDya1xlRj4h/a9c3cRbOKJ8c8/Y1JF7V8fjWLy4BQomJ+zjmot
G7LpyIbuIS5nw5CkVW5jNRzl9qp99abS4pIvBQ6enrE8jIhWKPaTq4O0hgLFHuoZ
Uin536zZBY+lSFSz4QR5DcVP67FVd7zh6J6cYL/akJqLWMjIGNCHpGgv/rABYP92
n4/oZ37VqMaF9DnticOL3s2F+z/f508mEsNlC//9QHuWYxp9e4c3RLJNqlVZxnWg
CNWJ8sSd64hR53jSFXBvcWbRW+INdqV8eBa3V+IsnsD4EuYVn1uuLQfhLYXK16Xd
jwUXtHeAHt8xqJUOJRge9YkVRvicGGzSCreYz5tuqEEAEofM1IEeyMOHtIpyod4v
NyrjuNzh9j8FwjeXkrCi6ID7zXFwSnV+fk6s8p0/OQee9u8Gx4Jt/XLuqPmH/P9F
rVeUXtvecHdkSFvtXcx2lMezs+sRqYi5/Vpb9QVZqRE5Q1Nk4CbFfetH5mMOvdh/
JfOq3h/STWc9DPI9VRm/ZB1BSpdaHj7ki50VqfP0dG5zErL1RMwes7mMM9ofqH3V
QfLb6fJpAmuy8LGsgUbjimdgBSTmfwRD6STgs0wkumOYbf2DOJlaLU3viTNxc9OA
3SwYcs07EBPfu/rLqMHXgFzAeWVXa4InXXH2fjrdSHS05O611B/wfgBwxqt3wV3I
D1bwk3fqfZOpZiOZJbh75tNYOQ+kHKp2+0wjKbAPJMQP0vyQykNCRzFvcAWNY3Lx
qZj4tYd/trj91y+gpXApjtUFafmJoMxXbanwQ6ZwylW45BAqGFyzDoGf2TNLKQuJ
HZRnaHafA9gK2tADLKtTqgm5jZOGSRS/obh/AEy2k0CQTZiXmkhFowo/WZ/uzu67
CW6ZF2vjgGABBX8spfYHqeOpHaznEw/ttboGvdlUjb5OgJ/qber92UrLFtAJL7TA
XDlhihiUlSolfMCKrB0JjKRC9+ZEz1VYZXv58FXT6EUsvPaVCXM8OfjZQ4GPp4z6
kzLgkmAv3vJ/RZHdD2nEfhyeTN9bxkC4PxGJxcnLmO8rtj+u6kn0ZVu09E4MC68i
/Dk20KQQ/XxRKknTLd5JPUnqs+huxJZk6QicJYvaRou93x5bVaf555AJ++KpiYUz
drhWwUIbQy1bKJExe2Mk59tKsvvlNp+rbGIkJyNeoyeNJzW9OJAVZYLb0vyEStvq
/dMhbEEDo2ViOMlG9Ab2BNdAjUwL4xRKrxWU0r86wWFYrSb+0WHuIDzECSHH2JLM
X7vqo+ZTd+euxMlf04NLI10zNGWmbYyQE3I1A/WipXV+zFF5xSKXDu8HfpcbASY1
llAiTVVxRnIZoXBYGvIzonuUibLOpBs08K9mraPxVbgQ//r0Eo0BQBdj/E7eVSFD
vA3Tj/pWuwVKJKe/YSL2rLnILGlX114j/jbeNuwDxI2gEgwLqu/TH1rDfhvMphrs
IL+02W70xfv1gaucA7XmL4XdetbpSEs21n970H6sRfGtnhFmBKBQS/QaMpA3LKIh
GB3Btflx996vUeReCzOaj/yN4rbbtLjnkDRazZ24gzfTFmrvXXGNNC1Rpzak+4B6
U5QDa75qx8I18b36wblMDzo+jJKqdQzWttZYWRUf5AKR3o5zy8ZX8krgY9ZLYjx+
QdiQRzPqcl99Wtj7pIiKDkfJNmT5WlpEBXJr8/AfCZSbPMKMVPNu2szfssFrSBbr
rU+lrQ7AlT5rvCcSGlWVu2mW+PrLY8/FlgnmSsfiz+wGKiJ7Ipul/8T/h6vAXJL+
jqvJf2HmHyzYlN7UMJYYIGUeco268VP9XyzSiKW8oPXar4rL5+huuGPFaWtv4IEs
7RX8YPIwhd7KOOGMrnvulkAzbnTJ+qBFS/ZByJ1s63roEgCuqFTOd68jTwqGx3uc
JqPNmHlSH4+eFJsV/dCxq2QDLtOzdmdrz92iCKNoE8HK0gzc7Bfhs3FAvnHl1p34
waHjf4cRdQhP+JjRZKUR9avMvPSFDAVPRHNw0F/3BIv4NyhoY82ryqoYpcdrwS0M
8RfA3dwr4nr+S7vEQjPyMdutdNZ0pWBGbwzcutMKk98jQuDt4NeIT9jyUS8OImSA
y4dDDheDdM2YxielcaqpniNJHCOoEn+SfhhUgA9NcmGYHKzFym6sBqQ5Qy4u0KJB
YIXoneJAsmz5uQDod7zKhu7JHVw1rAb5hT/n1i8Ndwq9Xc436KFLoospTZMU6enW
6sG1/v4vtnBmmzs4EJxzoQmzyRiQNPk6ygxxubDxOxw/+V6Gosi4uUItZaPRBKKl
7NIXv+6sGoml8X2OF9tl73AUywFT9rhXhpc/0dsm3gVF9yfqKKjUgyzmJRE5C6dr
nZ1tjx9sNQ+bPDl6btsmC9RyLNt74kS/UkHh/x+bQbPNp85rP0R/XAQPRoDM/Mvu
67akjq7sAs4yBF97nzWZLDstk5LxJH1rwJZ2hkxU75YUn4x7vqPB99PDlKN+E0Zm
t4Tk/dEF01/x4UD9zY6bjlLkXiX+3LsGrey3QHfZPvsZp3+5b7AgQv5Y5hnjdSOi
6nyk51Y5itcg0ob7bRKt1nE9f4S48yjL5FsNd4ZKcRBu7nonXjDungblci1UneQH
muQESfxppXpHwELEy81Qkjmz1aLsPanKcOrhHXpArb1zK6GoMC5PszOD1dwO5Mk5
l2tthGAwOnWg6r/IyXGUJxfuRsyM1ofgndhml9ohqNxMotvCIgNdrzNol8pjIb0m
OnWQ+m2f6ds0Epz3labzJ4kCtXA94HAqMTENo270kzbAjPR1D+GIEuBCHkVI7RQw
oWeHWjDjhRa3n5hPiZjXs0TytmlFJXNsk76KhpDNXCLvX/FpMW2zf6IA3VZqcYjX
PnS3uc4Nw7kWFWp8yiOEyZl4xwhauwy0vcCmCFL48/gCRQQbI6OmoPe07FqZSFUU
zRX5xtbqNR501kJv5IjND11RPXr9Re3JiYwIK1LGHtKGXmt7tTMQzDOiSazRUYIC
RFWOZO5Oe++3O3Jpcj/pRnsU6ZB7l6CDcfpyNtAalNO74jtI1E19MKtmIwJacev5
L9lNxMeiME0oLh+D/FJ+gp3YLunRa2jrKJX5ybRjQHofTbJhTNJYjPnDJwe3muDS
QgBLh3Zp7GXIp3pMe914Ss3ncHYFQCorY+CEdAr45gPzqlYcRPl4jSrCaNicUqzE
0bhMCf7pr6KyXzBug4R9KOXuKc62Qxug0zpMI/kACOeV6weQArok74NAez9BCPry
msDDIHhk62vNm8q8c28T5NpNYF5Nl7nHXYVX5XtzPqF+2dofLEf2P4QtQmDUogXG
YqK1z4dOLpjWQWWa7WL9fL5FbggqCY1JB6lFSySwP4PHZTYjjO+Vgkp7cwGxuv6e
M38jh2oYIAgzdinc4ZE4WuKIQISG2xbmdBrfnwVxX4hAfC+o/4zFJ7iA/owmd603
UwfN8/6+BmpLIZw8dBj0fAckUSztwYlZ9hBSIQIQnbs4g3GmTnUmko2q8lIqxuXW
VyIXpeeiOilgmCHzFdZOOKUwdIPhiXBYG6XObRslW+em4AE+13lbbQJ4Om6IuquY
qpBtq0sCeEPVBN5qEsF5pnVabPPJrMYoKRXkgd3SeIZFXghtsNP7VyR1NirHaVtI
dhMu8Dq/BmyVPQNDEA/nLIXO0URvnt9NwOWLh3B5cLqifb0soz4Jyi/zFALI1sH4
H2y/7t3bch/qxSeC2Ws3m/2uxCS71bMwiDbxhpeXtrcXqpTuFMa8e80ilNoJqhNv
F2GRCnDhB/7n+qq7d7HZgPq8YTj/bc78e4t5esV1WOVJ3G/gc+c8q22Ur/c/syi6
RV3JFzS3+pSaaUqpOCYmgPtk34/U/ARAKmWWIfmo5VDXyvHMN9UO3bAnPH78evzn
dX+o+gS5wx3iyU9kfIp09P1JdJNlt4kgYlIsrIYCA02jplb7RrAyN7NMOycpQP/1
7ppPYwhrMJ09w0Btn6UxdLvlQoLI7UN+RYdA1Wp/DutB9qbNDuVtoNH9A1Fuuz4Y
LTfnZEZZr6PLyylpKSlYZ8G8Gk4Dr+y/zv+u2rcz4zlJ6evAG7hMoWmw+VoBUyHc
DQvosiDDkfMjg3Z4UExm7V7vuE9IEjTbwpL37bR7rlQqbpZvoX0YSTxQTuToc5Bv
au+U1UUWzohsHJR1hRuLo8bLSc8TcJdaP4OpGIHEq90ra0H0zQYgMid95C9O1ZEv
gk9MQkfaMma952CwI+iH2rWCAb7Oq3+43W+DBYyADS17+CIPhjoj9lK1klAlT4Ej
TKJg6WpnNWXJ02ALBqSynLqH+XVD4t3D90CzJGEhb9Qq4p0W4AIaEZDnk2TcfP9a
reX9o5xmTyzm2MmMDPdBLpupNZNReH3MvdvRRV56dkOR57UUjW6BF2pCKOPGpuiO
9QCB6/gsGRw1HWLXBgGW9uA1FgmB7yURjSuCPEUhwRHYMOXLqXbBCgw9zoOeQWHv
J0Eh1tOOF82PgEFyYco/pR6iYPfxKTDgP0IL9Ew+60P6zz+NkM9g2/mlvpW5No++
cHGFmU53gi5+SuywuACiigKyh0XU7h+uOFoHqw7Z1zTl12INzxs4ylhN57l5F9uD
an/ZaMrmktCadwbaxpL8Mdd93APD68L6BMeTod9TQ/h45i80w5xcm1jSqs2vUPjT
0TNejYmG8V4woQ7MDKpdn7Ek3KwrBajxMN9U7s9xqyTrrQrY7zMhPQz5z/5CMHCo
Y9e2UoXBz2WdPFu73aPDGZmdpH0RTOHnoxeEOq/uNLamtvTG6FBXQaLsfYRp/MM9
pzHoFyqAD+Mg6olCr2xWyA+j6eaBUYred8cg3QHYs6aPrboJEcFBbYoDZts5xMKH
xvWWVuNMJ1V8knpV/qvhW3vMetDR+VWomJo3Q+IoFTz8yEk+AG6RnohDJ7BCIhNw
BbTPb+DUW2UfVz7UtXg2sh6l+VKF+aaUGExBx1pXSO7IlO1XmQSvzsg3xqgm2Kga
BYF3mOemkr12ebM5cSA7Ksp72caSlhri95ycTT1+Zh9YrAUV9mz9G9kRhZkEOw2o
+hv2ObSd6DVA1q+GsD3xkk1A4RAA23uduWJoPWKfsIapfsfvNGguG1wCkjb2SQqK
HV9O94V3LqaAAoOodRLDOKh67jp2RFwVa1J7HzYXzOvj88EMcCPkBw4jRckMxY1q
C7/VJwMjdX5V/jBWl/w/HgXziu3C+uHuvWFAfNJbZEf9QEov6pONK2yhFz2D9iLb
SIUWIY555wfmLeO41w7SziW5fSP5fTnYv48GuxXcZOF02sad1WZAnPcnOBkBhrP8
0a69zN9S8DhL/WuoP1qO7iT+tqVhbE7etxh9YCUQms1fINWY3W9Yr9Na/I/5fvIe
MvdVb/Emp95zem4sy5oFr+gOTlNzRBMduVg+gOb5JphL7/lXfxSwugxpmJsEiBT3
Iez55hJy4/K7H++eQ/hxtxEufGjQHe0GETMzQFOcNjOTyexsPFanxR+GC+mEkPvD
HcLcvGIlV/P+556CkkkCJ5Dz8qpGF1A9CDfVBi0SJ2sVeg3mKMLe5qgYQnu+d+i2
04H6HsndyJcEtYZf9VS/gLV+TD4RR6Yhf/l3z1Zm/ZOJCSnvuHx9O4aP16/8zr0t
dmBbQ074p0mPeOHKUeCyCx3aennuYsanzQ/5Dl9YOu+nE7MBx2M1wKTUZw8/5Cfn
8EHzHpOg5TmGb8tTU+FofLUZURUPB0beBRjMnXAquRfWx05nf2h3FWWfavV1oUgu
+a8ibO3F8JynndxDIrmNmAfRHgmMiedtGlLAqbe1Y0s0Tq+5SlLccMtzrFox8t0j
l8nWDOxhcHNm9i7uMXDR0o7FQJ+s0q6GcNQjsMjFPmpfovUHVbn8JVGGJGuEeAND
AGFnpXmzaK/1Bpln9xxpS0a12PljHu+o15jLxZedTH11ctPsQg1ZAw8e+vKCTA9F
uxQGEhrkZl7ksV4eGx7+WUgOXk6WmXqpxiWx/VuCCb2/FVvRtPKDsUSouoGUKIuT
rWlSF7N88RgokvOzG9zmqcKdRjQZ6maJLfFOSZtV09UkeN8Ydi0ezq+IbuWLtqqI
fs1xupVpGmy/KPkoQfPGoTjTnthhkicPvXHZTkDQQK+dnDkdk9WpIbdjcWsnbi7o
Z+7LV8FJD1zMvlaD/UyAk3rauHcl+hl6JY2gxDxTpp1Thom79B2gwlDISn9nbamd
GQXBztg8MmQ8owmNCs35U9aWtfYv9N3mYdHWRpJwY078KN4AdkbviXMghWwuENIk
9gTrGM9Qri2yiO7uIR7Nj7CdaD7OymiDk7sjAGcsB0sfQkED+Bwj7NfrijTPznl7
vRWV5InkErO23jqJ7l3gdlj6PBmvLQENHCFkA6rF+1viUyrG+VYY54sf9JOiU3zF
1liGgfg7U5Lb5hgAhScs56dS4slMQAy7vPBoV+eon41zhExpIhoEFD0MIPVh9bEM
Egk43NWHFbcRMLDeEaFAg01YxVPMKfcr0/nhL2GiKRYviyo9m9iI7LRx0kDTtp10
HeuhZpKyNCrtuevVFGLiLxljt5PM0CPQf8TcTf6Tp/qJJjHOXhddgM4vUJ4fNb5Y
P4A5Hmmzow2vWBEUKEYUK6glizIS1jBWdzNm0l5C202Wvx5TeY9vmasT+Yzk1j+5
ZwYFYsrLPdc3v98MZHz9JwbO4/KPQ/VaC8zKqcjb1j2nEpwMp34XQPj1LWdggNzm
QFROP7lP4DFFj7PSY88vV4JCeGmwJT802RNECYYtu8509Pktloy5mjUgAzsCB8L7
Bul1Lt4slqvBYHqpFQaCNktcLXIuFprsMgckAYNwsFqqUX0IXnpd42IH2kyMHcCp
IgOVVVaGRdA6sJF09mFLF9hd2Z+dgEFUFeAAveNtC65sM4HkSCvJikx/mbx9ppyV
vtu5EAUMBVekH2uWYEbxVUpw2I+XkOJnKKiAIvk85kKZlguz1Sb44HhvubA0GAje
aSa3RQ6ITcu3ibX8pEpwjM/vy3/GdvTrr9Tq9AoxUhjPsDmZQ8PmFqKeUyuxJuOW
kM4VBl0p9bo8tHNeTvZ0hXJzFXqnC7VWWezBn8xtC6smaeL+FF7uccnwVrXvAn59
F3+SPYvw5b0MevX5eMwPKmEq9s8/HQSSwuQn4IOw85mQfx9rVYBRKk15aFOutmKu
7NFzMiFFZL15SJ+9jOUYtEsm6/3WOBT3u8b9+ad+xNvRt3PZWEV7JkRWI14rtyhS
PnlUXGyhM8BWzMINk4Zgs2BxBd8iOqBQKU+YPQdp56oMbfBk8BEXo7I8DZnllAL0
bmQKTnTqh9gozBlA8e0bql1KPtZ27sbPtAPIqVmTuoADnnXbX2NH8POIjnGFlXKw
U8zSHenn6+EzayGF4jom02CeElFcLojSl6aLpupnbpQk5xHVCuIiBqYCV7tguDK/
KplHdx//3VvSmTCJAQWkWIcMpevMO1RMcPPLPnMHJKD3Szadc8Xg4Sm76Z1MfFRd
FeXWGVFvwIx6dqBSkURRQPavP4mO1r8O9sHrZbkMkWz66+7R1yaxv7qCPStI54Ee
DzzPX0vcWDM7cpc7vTaDGfp1rYkZNYzIHGRVfd+N4rzLu8DPwIPw/lLv8Xw9N3q9
jw82kUPFd0pei/rOyxAri+He2Qat0mp+qcEVAnMGqh7pv+/oIE7M/r64EJEQmIlI
uISSAqIQAwxF6dalv8Mli7INeDWq56ADKD6yHNWLGSplcAt+7hYzBMX/KYABxIuZ
OSeyhcZr1qNBVQsbVI4mysKUzYgX5ywfdYY1EE8131vjvDoA4g25xXm4btXDCjlG
PHZTu/FTiV5nj2DWdomy74TpRFqfgwG6ig3DlhOuk7ObOwSY/PjNIxcmj0GbmbjP
+qs9fJWrtZWYei7Wf/HrCCSgEBkiN+hdMrM4a0uEukkx/+wmhy8bkuFbKqI27/pi
0c6c5pcaG/lNB2z+6ZEZPOY0vYTDNT+lxg+GQ0tXHcicjAZq1VA6xxaYsmVxoJeb
ZEfBODk/sg+7gp6RQ/r1VzJ/ILXrKmR5235DVDsQdXI7KQXnNkK2IORgNjKWZ/xJ
mzhHgonux6wLNLYaYPc5irlVf34QyRD/D9+zV5w2P88ojjiOKa54+hyw/pe52jEC
jLJRgJrmGm5G428llIUB9Li/2rdQxyS9IcXwqaAm5RoJBvYkKAIbCy3GtQbfj3+t
Rkxl6e/vNi4+txlmNbWy04YPHdS4JBHNouZ8WVXWitECt5zVRKLqSJUaub+iNaiA
xx8gIXo0oQFDf73Eiyhp5QiGxzmyfD6an1+Kj8HBCOB92hcO6QlUFjEKuL08qAzQ
wOBLeozsaSfSwk63/ouhvI/BY+FsBzZRlOGdfjAIC7wRzfiDh3osaalXsCBc9lzd
c4eKhly+PP3SMRgixMcr3PUpaHtmqE5FIIlTLG2aIbmyJLctpS2n1rqbUxc3F3He
/+UxhTLEgkz/r6fFCVbT+UtOBRissm5nNHf+QfoEzPLfKv3f4KOGc47WUcKbctdn
cGZi/a+ohAH0Z4ZalQ9c6LqSVgxzc6tBojbYlptvNSSvd+cVo9LD+dyqtxIF3JLA
DgjMc0aBCF2faCdr68oy8eOpw17/4JzBRccbfUEpv0s9e1bD9Q1FPqDpaC8SWSS1
c6oOZVbFVUnPIpyTHyZskQSbtfOZG2WdqHcA2okKf6OVUswQYFfJV6XYCP9OunUu
KiweVhIvJUmCvKyCjnweD8IpKB/i61uaEJIbtLnQbrO89Tb3FWODcP16380VHK/0
1KeBIbIj8CY7m1y9E2lb9kUSxa9bjLtaQJM7RzSny/pun6jiBYSFnKAn9eXe6TAo
Khh7LPJAxWQUXJPVv1YMa8ceC1iLRf04PxNZuGmHIpwDTJAO0QIPk6Ow0+w3erLZ
oIc/2ErZDcZLyRd7pE4VSp3ksQ2356m+Qu17+ba0EwJvDJGHxHtuRbA1NSUgEJhu
FQxhldovtvCuo4tLO5WT5VaGPQJ6uqc7oh4MRgaeXYUOXpfDr1rV+AvInB1MlLAH
mhG/cdLDsfDHh7k49bWREKLXpr33Q5KE40l8uBEeiCgS/FCtUAJXm/11/7+LJZU2
8ksm95ygOj0yI36YLC+M4WFY7sWSP8q2/Tyd/BGt2mcSZV1SszMo9+6rBAz2cnyj
nWqHnXW1gnca8EvG12W+8CCXlUqacmEps5tIKZjsjXu0ZONJIEkVP7bvwodwAvIj
CPkx8VtUGYYYxN181aGAU3wdWeYkaUtI1fnkO2gBbRP42svO9HCTeennfVPRvdlK
qC1AKdcoUie7FSCUw57wwnnunQlDMr4XuNx9DbxgEB0FompS0dddfJUXR4MWAWXD
oBG8cgS169wGxX96cX21K1NL9rJuRoLmfkE5sJIKuk6fpZpR+Shq1+klFMSAjP9t
sRSTj/gwMiKLzhY20SVFbghouTGZJxSCHjVWFxQLauq/bMkMIgO2r//JG6gKs9aX
wLnZUgm9lTNVk8YYFJN+rcYNl1gfq4kZjHRXohhDjQFVLdUuHfEQkc0kxpa/XME5
SpI9T7ueQvZmZGKr4yPSA70iOAFEdUf5h6ciHa8bqS9M+J23SreChrbNKJJK4Gr1
RGnIyVo4Homy2sm1YH5aCtjqowFBWVwZYq7TYV68vW1T2xb7o/h90PyT1xYm/xmW
FO7tqHsrZc3Z2kQZnBSXUOT8WRaMXrsrbLlxvkDPTKqSHZD3ZAmYByAP9GbUPHer
HAQU86CXLfB607Xp4N2dFYhR8YamE0z6xRfQNJsb6mWg3bLeefYUEW1azPUgs/JV
B3MEuCvIXa+6pnzWWQ3kpDRpKQRDDYEo4Kp/HsUAzIdQiu1ZBx4k/z4c7Ugvme2y
yGYBLYGZh3PFUo7OrHuJrfPQSaCJ2IDDEaqC9TDd+ZETrDDmhmPIGajDjsnCOkW9
XoCAf0ZuF/JRfN85hxuz3CFrUffcYrT1KP595tCTtOjuChki6/IWuR0Z1CUldjHI
S5h0fqrbO/tdN8kSLWbHhOOcdUFKMnTJb4JDMvny82FfIRQmO0rjpjmbveDoVOQd
ZIPLf0g+Kcv8kZ30DN+b8iKSVBvj+a9dM7RBBaxXaqdpISaN05iuWSbBARMSgR3c
nMnsXRhhBfCk35aNE+iPq8gK+AMoOBfd0D4fkcGH768iM/waqGyZ+ul98RXZ1In2
s6J1WKctNKlX9bAikZH1CObYGXTqFBXzs+++nZiSAmjtCSoI5wjAmm0Ew4HbcP6E
Iogvc/AKmKVkZzd6qlQRsrNeLHFNJ057ra9TPf68Wrix2X6s2+T7v8mrnr4ECDlF
8ceU/QxWTyXDna/2PRN71GlhCcVjL5b61J3NiURJ10DwiW7R4dCdHpQRrASFqC3y
0PA2TRbKYDhBktHS7zfu38a+E4J03Lcf62+rHGEY6c6pfhit3JvYiNahXxSmJQlm
JoiEwQvCRNX4t6eTjaSv1auCiHi6OMXLWXxrF3AqyFBlvq/8eGoGn2H6dI/yGzNO
Ce24prpt19u/TFAJgPYT2VKtAfOdWvb4UULHh+jIt+Kb8e3UMyyj6y0XgkDJUwGE
xjd6hhh7vmrlD+Y2068AfQ1buzSX07VQNh35PXCDTR/5qCYTpJ19X74sT0rRt8Wd
ab2nl6BCNMkMA5HQshz2hY/8HByjjLkO66c6Kxad3XDX461VDlxw9c8TV4Rn1Zig
PveaWRTf7tiqRnxKec3r8hGX6O54OqNOHW5z8D5Pqf4L+xnvERzbheZSUm1xJ91j
kBjZta/I4KH7RUCKVbK62kib0yWU9UGA7ZZsnANll9ID0odxNGdyqMyIQ5CTs0ii
6/sYiRt9vteBMYWtM8L2PHNTT0aw6Yw6OCxJ7U8he2fNojPyfcDhODqowUcH3Bgq
ZtKqbml01g3lW2E1EEwhYPa3kPW9/es5ApmRkBk7Eje6TMrzkGxpciWZF1y4Mil9
1wyiTbY0kIhXJzzD8dsfSenEH3zf787ASk6XJEs7F8Exg7bOIn33Fj0i4Hd44ZTr
MjST62/X25+tZgGdY18QeGcMpPKOsp19rb7m22xcb8uYaOzPfUylDbdnJYQk9Reg
xY7aB+D8lVGjbCAVO5cZMh6gQe4nKpKLXQ6P/01YBOgyAB7kWTTgVOcJZGXDrfwe
fBrUsuW0V81h40yFyQm1s5tOuH1aNKfJVE/MAcNe8QU20ikq29PRXmOv/j7ua38y
lCNXmiRt0FKWLjYSM0okOg0Eh26gfGZhsbFF5BPtbz3JHua/AicOvFUFzAi2C4BY
a/fKL6qPfx3kRvWns2a++7spxa2WIN/wtlRo0hLahg7yVKh6ZnTtXITU+mvdcuep
bIELNLR5CL//Pz9g1BVjex3fEpnrjcnB9WDcAxxUNMN5jOpg83p0/g4QKbYDXmju
y9ASeKXRAq7viXPmyxXRdsFHOHY8ECnnx4KtL3WYHjL7nqnSprhKsEuSS63hVw/y
mkski7djN2U7kA+adcVWn6iUAXlLRCKt7Xk9+mHgWspIwa1yCDGoCTeD53LMYzz9
ryTt0KiGs7vc1fqPrOBPno1y1NXHribE05u7wF16OoxN/GAgUxNkysUhdySBM/VF
wwigaK0W8t4I0favq7oRMx5rAaQ0LTcFT9EsWU+rd/GTNwK9rCGz8+sF5u9DYMc6
dhwNdRd0vThzgmZj/KPhzwmR4vmpom3k+aB0Ixv2XGnBwaWM/g5Qjbw88KOW8eaf
291fIOh2ryKLNDliHnFUXYIXG2NcnwNSwJnmLVuIucXNNwISwji2sAqpmzMhejGV
F41tfd0ynPtIcjJLuou6UZ59idInQ1oyN7+gyDfRaW9VS0mtmzkycVXETJn+9eCe
EYo14KOPaRhGYtplisyVxaLlNqMpY4YCkk5MW/0Dsj/mb4Zs+t9NuJST7vmydTq6
7Qa7W8gwvOwSrbgmfrUYXLjkTjLpqoy3UyYPfsQKPMx3SQX9k115g0CvZxfL7dY7
sWzCRbS1CzMXzXYh+k8m9SfYvfYzznMVk8hZvj7lHiEZirBRyPlTrCeYzN4zt8/h
cCDfXlhYTMxo/A4YcAsl6Mn0pnW2HMe5C36RTRvjZD2N3Eu6P9nHJOL1pFHp8Nsw
ieSPgDg6DvjTEWNo4HecW4NHmAdb+Sggfv4ZQRP9HiarevoFdl0osYzWQ8CHiaDG
T8hhYPqML8FLn69CcdTlOJawNi4lks+dlzCspSG03jkJKAkaktPcqoHG0d25s0Fh
0yYvvpif25XZmkKWicvaaanaxtzb9iT4I929nz4NVhSgoeHoiRjt3yenS1iDSwmx
8dwAEGPXJ2uT4Y/wP5nVeA3O2QbrRtFXGmIB+40KmccgrwMg202VgltA7M8nh9Jw
jV44IYXxj7A20XRAbmbtrgxuqEoctF/OaSyLGS86y87+Bcvt05XLKoFXjljLiN41
Ts/fNaoPABapetibAw0ylVaxyA2yK2hvY0xzumb+SXc3ImTpkZ/5W3mgSEF5oxOK
+WAjJu2Qt+9Mq9stfTb6jnSH941780rOFC7I0F7eB82lgfnrAwcmaV8uegttNK7v
b+Rq3U1UMBerBlICYz3gYCGC+JHFSDNp/M5kGg6/rsbuiF6C3Rf3VNgkA79GJYNa
wZieJiQzB9BQbEoDJHlha2b+iCdL9Hbo4xdK9odYt8ifoIuSbaqo8sbh0C31PKCk
nqADtKLf+Vg1f4dw4T6nfmVZ+g7HEvIPivP/K3DZR5BxxvCVnJ6pEyk/KvVTz1a1
i7BT5Lus3xzjwjT5tUbYIDhHC5ZyScfhKTkrm1BAZfXl1kJVPY2WGq4o8WGjsh05
mHvNkzwgQc8VtQReWTtG0LHCiW2+7yLEJOwgPMrvvvNJOrrIZe27eJxdLJ2HtO0G
vzybvPrRUwMF4PYLA6RglvzE6QQ0fFg/uS+ZSrbKweOPMv4b9F3dlRJU+/zEjirT
7/xqC6Ab3P/j8k2r53ic8lu/HQRsQZZqZQkPGtVmtXWsTpa0VgE+WBDBajzeV8GN
UVYmgtSFEaDJCA5a9MgMe3ufJmknjX3C7R4lywgCFKoVHkOe3zyKEBgRS/lOiYan
oOCNN1F9Uw2udIHK/WOdKS6IrHwUfX7bmAbJsiBKDRz25TaKWfF4owQWD+4KvGGa
QNG6J7IbuPpilcO+Z4nZ3jA2BedVSM/yPcvG3jI9AqqBWoETF3drrLES+5jbSNdA
gj5sxMVLvMJJKknlwWCUnrxhZDm4AjSfYqd0XQ/0hl/MUnsbN8U6AUHGQxDQ01HC
yFkcnXbK/Rkdaz3RgU5NUpGDky66PTHp1v1270+xwvV/rhV9iTelpWbWYhbwti0w
/JjmSLB6VhZUVts7YyvIYq9Nq1mBXDptNixEuJabF4y8TRFYGlO/FHENezzzgrEz
p959aJQZlxWgL3OKHcrxTiUHfBjHFS6l7DdVRE5wdvGqRmhK4mUiITfOEe0kGbi2
0X5cNHA9tGUsnSKyKXInco+tMS52tRDqBv9xEw6bxKrrk3m++uFuvCBfeHSLGxjt
XeEs2pWPgssUNoH45pz9rRfEr61J0CiCkj2agyMtLa6vtHIoO9I/EV51w77TTIcx
VzOILtxWJq4D7BvBLfVvF9XUKTeHxA6w9PX3uFAfC0f89VJ+5MaB4Y1Pm88dEyni
u1v82CFBXk0Wx+XQJYkKgGs1mlodP13dnQla13PP/7MTUp8ejY6VBl6ukGEvGOAP
/BLR2WoFM6Mzl9eyLf5UkW4/hCMO1yq2rp1j/lPu6idR1FdxQvSo+8WabDLuVItm
R7bCrIfLMMjbXCFKOqGKQ+2NVAcZeJ0qaa4jsQBlW1o+uAyGPeN3dW56f/SV17pA
T1FJnwrx+d68IPLCZNuT4FQ25P7er3bK2VbCjdvJdg75WPTLQ7ZvKJ9s6yFQICls
fw6Sb5HPZfjl8q8/o+PgHizgoQZl6QMyAhUj/iHiOzID5+4k7qzFsWaNuFA+pvBC
iZ+l7tGGFvgljPLFTLQ9hx9AtdX6MzviasGM7CwH6xrspkf94B6KBpuK+f5yME1b
oe7Bks+dqqgCNonPFhKOI6D+WbDDMcFsiVn5JyuZ8v+tZUKohUQNR87Sl9DkIkId
aZRuBfqiAY63Zyi6VFERNmweZvPpR+8+f+V1nizUb6NNdEpl3GDbkWmYq8ouqcrA
vIL/DpAqNBOCUGuh5Qym7n4hL2lE/jOcLtI8U6QzYj7hcnYNLDiva7Gx8wK5iV0M
5uagzv8mjAAv+Ygl6Y/PXpvupP82kjtZ6omMyM54H9tv/0RCQojp9U8yARZDHdjZ
uhhmORhb8D4Us8a0Ho3i+BJlgITqTtXxY0t5ap8ZVFPmHBPaIB2Da0qcO0qPOqrY
2dZlf3vr/cz/Reu8kJILqFJ8iYGBwpiJztR0XvZ+ARu3kbRjHj4C7T4h7WmplxxM
NmZiBsF2vyigSPuz/zZpoDw5NlWvqH1ZfdKGL6J42k/lOq66UUnzMujk+PEigZqy
e4L2vu0DFtHxig4dDhm1NqQnFVDOdLBcTg19fJ71wJ0VSMX/G26VbIM9cAyb4fYN
Lq/XDULHtm5rvbz+GkeJifWhXjQmW9qVItKg1l43aBgYKaIHgRGjJ+Pa/yfXs4rX
NR/C3prah0mBFKzSej6ExVFY56TvadeXzyhojFEJ3fQQgNf9GI3jMfb8okYZ5bxV
dbuVYCLkBL5Rl/uplA1almb3o6C1G6eK/6b0a4JuDTWkH1ixItYVsZ98jmqpFF7H
d77Yl8FNcihJbFwRDdCayRHLDRPLnat0qi+hugutbNNRkojNnyp2mE9ssIDF0qxn
2BOIk3ZE7xEC5q491PMqH0Hncs/APHLVvVxzIj9/eaBTtU6lItoZdr0A+OK0GysA
WfcOMNilj+5yDawylgKH26khC6ayEtbuA+s1FyWQZly+hH9koWUVSTKblQUc86z4
RKuXJaGS4+yT2TmqpvAjvYvxe3D+BltNm5d1AkMdm7SP6JKuUD/VkfrjQ6Ags1eP
S+KLqGK3yzkn2UJLPDB1Qo74kkOBMsKbInkKaz1sxGzznIr4RRJbShs0561DsLSF
5B8ZXrR20+QdziWUFchZP3AN+gziiASY/a89NZsRgJJSNc11+sKVE1yo8Bd8RzJM
nO69ybHURY9QpcLmC4AymKJ5BOvHmJcGCgGOn4GuH5ECGlnm0bKjf0/brAkXd8EM
velZOI+KyoeGYbV9bplWGD3Vu2WvfXQ1EgnrMorlVvOT3avlLwfvem6gIIICRf+G
RrY2VyD/nSP2PhYDPwB80CEV3uY52s1paJuFtuDRmICr2FwxEGDD038KJpWXEyfk
DeQlk9+Ovo+NmdDSgbcILrY43rImcck3wDHwfl3pifVZn0vAzvkr+0JoLKufP6IV
kCPjeZHJGyJeDbkNZXqnJXqHwPFOHuoktUgJrRa9Lw1fBVecdejdAklLvZm6UWAh
PeoBdwsIFjTdFkkLg7hGWxYVEjcxiB82pyrhPAuKAWYR94ihf8i5Y81Ehpv6ZKPe
HwOFoPvUi3v/VKMq1ZLAZMEC95sQ5Q3oeLj/h1/KykCxBiGJDOkytorLEhs1URW4
iZ9EnfKRcpZ04jxc1wHQnRcZZlXGo7T5dfJk3DTPdAZXMxY/VJxlVR+2o/y7waMj
sgMMrA4ZC73pXPCLPFYPvMi1EurQnysH3dVNZ7iYxOspDSh/UJD2keBKEWOjA9wl
zwyFsHQxwy7eNo0B+JelKPxE8UYwGEcknNJcbb9vfQAz22GNRCPkYQPoyAN/60Am
i/KsCY66nNfhD82OiltKrPtbpZK3+F5I/ov4euPfZ7xg9QVefboiBIsk5D8sGOYa
1w6m0Zr9ya8FAsOeAv61rvpATv44bO+vawPj6STlMOmYsqshMdHGs9fgYI2tPL6N
3mlxcEJbbddSGChMqgDPxUgrnlJFT3uWDDL7SuL6p1kfvCf4/diWY2QSARuRgU7r
s5tgnoWdfDQ/XYYYc/1tpoPAe13+ArCowIUfo5KmlyqV+uzx4fezQr6VW17A6a7L
lMD2VUUfW8IWlo13BzQ5Jwqxc76j55hVlf2r+maCvEAYTng83mhzaGLb7GV/oltK
DRsJ79NnMHWMXbOdgZEyxRaZlfNJNjJ9yH9zu/cKIAxFXAJEzbTKqqTDf9aTgIhq
k3DUCTMoQXrq1ZwiNkpuADiw8+iFp+ksMGC67ld45r0tRuPEiW5hxSxmPUJTJGmw
sVVrY8TUBJmuw3kKOPw6EgfLH0rSpovwU88932VooGGf9zXXV/W3zAoMg+LfKKJd
GdnHlVv0jU57A9IM2CW37yGVxYT4GwoGsbsv4jdkRGpmB4SRLfoiR5JLryiRGyuu
gZpHqRpqFUlu+F8c6ubzR1FH3ss7sQt3oWos+Qj0BRYQkvIepkkXtbjtr1AY8nqt
YIrbJ59zKFp1yunEpqvwxHL2Yxijo+2nsz+IqRjBJ4j5FUIDiHkaGm9QvzKELV8g
nEoOMoVOmg5c654sPUheY7+Rw8V9jjDg4qkn6FgrDHrgHjIbDjmlyraFyJbr/JI8
kTDVfzYHTMwfwFXNRnIfYwJDhcoIe+F18bIpEP9upLKkIsQflBJ5aWU8mNELfkNv
eqm64i59fqrGonHv4hBHT+ozZBScEI8gZ7iryNcADxvJVyyaKIzMb/8bn0EHOjkg
RJVckOYr5wWybziXs2LDfhdy9RTap23cO+HtTm1LFJSpX0on+Q+69fJRlFmSG1y4
kktuAdQaAllMYDw2BM7uweCixbGdIudQXBSj4Zwv9mo/j0ftR5KBvqDaK5MvC9E0
kPxnEEXcIdofwkJlOr8Fi/BK8LM6hubLV38xCT09f8eDP+fBvh/6yEKuRLAnUYSL
ooynBVqpGl2K3HBruoz6ylaHLR3mZIbYjut7XaXCAqLD9eRx8XM62x/TMmbiggv3
mlDbou3z63UbnWDtsBxyRiTJO5JaKo6k7YPdmhrExJ+3S+4X9NAJ8Q0JacIn83VO
IW0tNqnot14fMlkMoZQzUZEzQsIOpb7TnlYI93fbz51UbHMImJG8zZcVX1TFQ0Tq
sniWek7Yqzdd7BUtqaFbPjFvcugTY6++zdRm4gCozdDyNJFqrPXwSw7OXd4n28ff
9UPXEED6IebL/QUXZFkvBdDcE0y2Mbb12Ba+t6pfAtfbGpOXrvoNovTCM+wdXjeL
FweOHnLJ9WMAWSLB/gqFboo4qKXY0aXUb+z++Z5AWRdf1/d61P9wSMaRQzbQL396
9bIGWl+hDEFrs8BlArp3Pf2bl3YJcghI1WbYffSO82re/iuBMemhchS2IH7s0iea
WCRGYQenvPD7s7o8Lyo+pjpCpdGnqR6ZV681n83QLfEfCVKtK52uVtTWxSx6tiGH
6H32Rv7oTZ4lfx4QDy4lFoV5fwWPQVdSpLmVsuSEuo3zqpEGVjPpy03Dv9anP6f/
L4JL1YEqGPVrOiPx7/jOLssPYK7J7gMT5RViMzhw96BHWhxsWDhCCHebtiPeDf/t
03bXE2k8O6t0Ydlj1ozB5kAwXLXYTeRgfhAJda6eCqho5XLtGapZR0fPQps96c5B
uPu/K+dm9XX1jKihlw0wU1IDrpropq1txknF0LTt9kPmiEJkwdgnJXZ3+aTcUvLn
AQtKMCMFERQgrveb57TyoAUA8hGfwXqlTeoRwzSge1X6xS2d/PoYQGS7EM5Jehx0
asOgp4wgeHyW2JOcN+kHYnygQ4Ai3DUWggUrYY5KefuZ9tTqb4Dq1VOffpKd5WkB
a9PjgMctPU2Rg3aBl50VWzIOf9oJTL2SLr86SZUeGl7vQw3CpPKwsp7ngzT/uTJN
jJhGj4EiscnvU4S3So8j50brNrY8nVdHaohsZWiEkX/2J228msf4/ex/EcIQDsox
A0L0wrDn1HzJLdzvgLT4Ig+5p/uq0lMKYYCEoVkN/keT5+AhRIho2NsLH4nWnw1D
2Ha/gERsVZleH4q7bGvzSwSGxEY2c5Ylki5M32qsEcOiWyPG+ExhfCuU8tZism/q
KG+WP61qc1U7PJ5Bvxvbyg1JvJy3Gtd0gVUBpR1DnA2Mnm3m4MO7zCXlHDyn2+I5
dz1OGLEpIkgOmZHc94jAycpFxO/jGaSdGPJkX/7xGuQ/fxjqFLsP+UNVgZrtOVze
6y/ULxs4QV4ERNGchNwJRkxr3MgHB8KaOdd5q/lvjpYQWSNCVO9Ev14dIc3Wcs/k
eKcy4mBAN771IUqaH3LdCs+q55JYanoUn4F571bH3NlLU9j2bZ2UNoiGY5hta3O4
sMKz0tvyR78eYQ8KfH2q1NUmfJ3Oth5FdVPgZDPTCA/Zosor314r5SH44JSmgEMc
gZdE4HaeamKLIMYSzcIr/N4R/fqzpnpSaI1rfSFTdConesuaJTkYRnJ/OCcOK9wu
Ak7cT/fTWppaBKwfyLeY3rk60Xz+r2CT+N+jmJVgXJFU3iJZa0lvsxQxGoYhmgmP
CZQaTQMmH0CAzCkkP8kxXV+4J0lwlkfpAsLlGTYWz2Y=
`protect END_PROTECTED
