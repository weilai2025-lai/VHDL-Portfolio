`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/zthzL9qs870AUI84wtAhJElTx1B75R4au6nHQxjnevPuHTfPi2A+gTHcyhjOpL
7PTy876jZM2xmKya1VR3CG9I4xfroIpjWagoqivxNb1ICh9lB8F4QtpnGX8Jba03
+c3DvV0jAQ/7sCKUsA1GXQ9opRK1Y10aXQSBXYhOlweMufwHfc+RjoJv2RRU2SZp
rP4pZ4Sr1qtOmzrJMKLoqwIZP2jYvmNVU3ZCI1QdWH5+jZDz3+QKVQqY4bpwfyUr
tT4JVcqJwI/QTgacxGcKLr/zMNvpCp0FodKaLuYiMpu85p99oBmRLm3pHRqe/1cF
boFMjI9H18bmJI8gxdQQTlokQsP3FGQgUVm5InOpF8FaQm+qUimWRK/pOzlQ26Ag
6L1T8aeLKqcPYd9BXbMdojcVOly0mXYLL3j4/q1cbipaDn1K9XSJHPOb1d8ET23l
y49dXWw6zknRUCs4oA+2MSSeqaKgjONfH+li4X7Z/zFx9fkOcNrvab24o0aX12MJ
VVIKjoGT8RisBWQN2QSfMG5IL3sluxJC6DMLBmjKn/ke2np85/r500vU/l0lRshc
SBemKhIKw70/nQyxLiCxnUwG511iqNu76jRPhD+kTADpd5CmZHe7FV4X66TSwFTz
GqmfyEsRgeCVq5clzyPVCAVY2q8Rj/aZFZgoFai6ukl18A8N5zphdPp8+yIxYvbw
qyrw4NqSbDC0Ari+7yWModsfaSuhdUR43Qc2xwEnh5rsDL8fkmujDESYlqwfPzJi
uBgw1asSGlbB+fzkh887EMt7w7PKAmXyEV51GQLwvEeFEQ2slcaVyjUFFS7q/wXY
Kp5Mzz4EnInRec0kP1ElThlktxEQi9KG6YaNnJiRIFoVNRtqDBz7PDdrAx15GMtU
ECCgs4VlVY+KNePgIaHH/uUbRHESbWNaNo9Cod74gn98T+8HoOUduNwya+1QEb4L
OjOndlwxCMzmw2/x8T7BI1SURPOXbXuV6zlybklHxy3FpKzxx/BJ7C+rZpZh0AI1
QJTA3V5ubBeIubaFGlENbgijceRe1e6rYn/9hKqhQAgCufZLRzGDechTFizQUqYV
GnVOIYEE6lA2/M5T6wkA7sNVeAn4AsVrixBNvPpDDC18RrriAkopo9FxKzwsDmML
ar1YBqsPg/QwoY/OQRU9bDUCkNfP7e1lDxpz6GGDiSFHlVA02uMkpJWSj05s2oct
d/cG7oHjIaSwm8+LXvzVH/5TgETXCJle48WwQmN3pyBc5JKEL/E7R4V7nWBg++Tc
imLt29UsqGny2tTYD2UhOjowvOfaLWb7rAfPW89zbp0Ei/wihdrSR2t4kFsMny22
UCHThmvNDRHjHce6lHR5AaZoSzmxFFGJC0kFTDG2diDhBq6QD6HDRZkCfoBWaHBP
pWYC+G8P9oOmpES7rGP29AQMtXedMnY5NggKH5AjymScSgKatooB6V40SSEmgoyP
VixG4DRPhN8nL0Hry0R4Yt0di30a6zSb1dr9xmchBEFU5Hz9GfRgjLtBUSp7j5rj
cyagofRijvRSu5dqj/snt1DKZ9rEX9aZ1CL14GB7dug2ZyaKDB7iEkKMvgTsQBhj
IGDWZ/NTj1Z9gFs0sabfkQPXCosBH6uDWfj03ks6oJBPkhxku/5/oWIjTTLIVVf4
k0QIuQUhy9Jdj8CoGF3TMurMUP6G7aRB46STkU2/mIASXIYyvh+gqNB4VKi9qRw+
cQbgYeFfwSKOzFpeKIwUBK7LLxK/xKOz6dmnJiSCe7oEB3W9SU2EbW3b9GAGoGJf
+oie50igpZGt3gyJeiAeJOPpoqE+SxAe4wP3uwUDEcVkp7BfBy90tUy11CAr1Bj1
45gKBlHY3027A0YplD62SPQjq9Q6yEWjIsNiCs8LZbvjtm3d3MrBS2WjVE+ausgR
eYUVoYQoBSJ+MHmUfl/VhmeA5kMEuFxufNYDf3bqu6o0F0vKAFZ5yudidVDqG1i9
czDAX4kAGFQnAesc/M3ilvOMlg470zJLTgJ5SSOANF4DCDxm84M0AHLApPNKGh14
HxLr1ldWsSXRhfylvt3tTQtNRv8UpOHnxK2KJRWD+sJ1RsHYPIJ42S+x8PeHM8D0
Jo1o7iHRpx6aANRPIngFe97Flf5ArdWThmPfIovFkrM/kWYKC/9PhT+GXpyhd4iE
Gpn2jOJhj63MkA3pfAT7o01Ex0sZ+WX+97pTLjyZeFUDc5ZDQLUorCUlTRL8DDqs
sKmGM5/Ol0T6wayRL2zK4nGGNhFb/8vQNcEL3JrSG7aojKqpcvaqy1NGlogkiqjb
CLGUWkMbPbTzwNjgX6Wed/jyecHito3U76dbCqmhYLbQDm9jwMBaCC4EmVf/t7ux
ddbHEMh1rgi2r5eIjKhDeOk8sDonbkBG+GteU1tXzBxFc8HBSa+Hd70nHjNVw9Qf
vtLL69uo7lNO79Sg3WkFhsqDlT2sRthNog9a3VudjUrAytanpVn7Bkg7vOeZM8Dk
ZXWw5loZOJtXaZzbQ7xlD3TFj+jD704dNJe8tFeolbRSiGlKLXDBKqNZbRCjBJ08
DmZqmcELU00Qajuut45fRs2y7rvFOsNQknbKoY0vH0LHK7WypfJWZn1Fssfm59Td
PZ9vTcMxXGqjA6DxlfwffISVxih+DK65KqLpSxUzHnf+5cSAia4CeNlVz8kb6mou
e27uD8a/y5Imf6RkLWB/xpDjjgrrxSx+j1CeG3JLK4Uw4ZXs0egcrvjgTDNYWHnc
/x7wBqZuWmfHRRoL4jh8IGuY0bd28I6ImiTb7qb4AdIUwuNLMRdMCvpyCJ4sKVV3
RoYAroZcqTZA1Bu6BHtgdOdo0WRkA97Qb/Ng88xqGJUanGHWb/hzrNh5TpqgnERQ
W+4NBTgsFooowHHzZwVkAZOMSEEp3r2kIHJf8lBJYbqqYrvEBvdkRP/8LrL/i79M
FS8qmxVsR86/FJsdmY5KM8wzd0jO6gBtfBkULQCbf+B7EogS/uEeWJ4shv1vUI2O
kCMQocR7rUJW+TelC2rFW+nUS4OUPaqAmULo5QImX1jGzqizgobDCNupgTng4REp
u/g4iwV1sLdaCwr0xl1rqRBEoOAVgCeu+iawkBrW65PAlZYhFDF/QlwUrfLzHzzy
oqz5fMKxPsBkg97uAPS1AQbd6akRhFm20nEc27vJN2IGkzBtiXgVwm3rwHJAfw0z
Y6GpCXqQuoaavLBR7N01zc6CyYq5sbXu0Tb3pS4XnKYzZTR+D9Vil4lSsEwEOnju
ctOATV4V1v+MnTp7q/QuMhtOVstDQSPn/E52cxWxcF+mmsRlmM1lxwAtZCwoZ92q
1kmBNl4Uoh4ZbWPF3x3izrKxqxT1MEOQ2k2ygKxJGV/ppsCutKRrhFv8ENryobJ4
EtLSNs6mXYc0AZdnWIY65MgVyUC5B7Q49AtBAW/KmwEjNSs1KiNxjvjpuroj+YLH
MPzhrQ/21TLh77v0E0U3Uu89W5GksVPJ+IHeNjjG9jwA+3RUtAyRBbX2cXbW3OMO
HxFVE4t8c2wbgyP5MUNadcGybC12NLDMkUsLLQymJwHoIkGnr88OwX1b69Yqytqy
SgcNDV4XXDLjY8oTHe8u+qT4ZH1OOBkJras6e805wX4ixW22rK3zSIwHOTDxwR64
chNUM3rjdsIuvtBmKdUtHVIgFwgDX8/Yy/ONy79TAFvI/cJVJwWyK7vH1WvTgow/
jpE+GHHk41PDjrV1KlsSLsNICIWgdVlnxds5wFBl/KAULosfLxoXAI0GDlbXJXEG
AaoHeJl+vy780u38tcfXis7SSgZUBK1/SZcYic83R6xapTVH/kXOa5JFaWrG0Ujo
yPSrMCM0ymNaDPzUtx5Uv5GZ4vEUA5jiXXEDKPpfKqfQ+v3YKORzNRug5shGAULP
2Nk6XnClxkxiq3EKXR5H+WUnhi2XeB8W6iKQY+Q0IOkZ1HetzwfjOq9mkkZYIOGf
ZqH0ubwuZEnrqdy1N840S73rkTQMXjPnJ0UzXuBNgHyZJxp83OOUkDcC4yvJb1y1
/vJXCxw6TpvMwUZ/+71e3+s8+vshvhL8L49E+enofpsisk92fgdDkoiLNVdE9YAO
/C6xTaQNui72QIYK8URDf+asry1z2hSpkuuzwSg/QSaO/+yH3fz5nDR6G+MDZxmS
+asakA1uVUkwlLeNIglQE7HH2/dtWnO3AQnkNcuNZJxlWkshbiGNkEp4MKU42gM8
8/kOGdVQbIR7MmobH08pmAJ+9bCsDmRRA5f0IL1WQ0+1EFiZvDnCcI0fq07SBBuK
+1WDzwn48xmdhPzgYN7jz2CDAImE9N8Q1zlGvbngO4JrEBhFI90Adc8wt4BrTGrq
OrVqy0DSfrLsR1ZlbNragonjKQcFv89Crp5OKzlUwbkl1/EsITon/bJZS68U/ZjF
40z4xGFRAfDBTyhI2Bd+9eSnAsUOlaQArEyTK6oYrpEqp1Wt0JH9FU0ZAftuoyWq
/IdYLKeHyMgxrXUNTY8dDuLPweutFaU9voXdHRbY9eeVLlmwfAAnDS9Zq9TK6Nc4
dv9gM+stdFDWkBDknbfCUOteJRoXqCGw5AoZVCngksbxJuM3myFlOxcxBNqCplbm
nalaNnz35vGXnZshgTZbX9ieMQcvb4BwgyDXCQoufCgUyhql4ZKocJTIdwFo52ia
yvBb25SFH0QbhlLUnDfxKhM2Z+/1y84IO7mcWTyVJKmigvOXG+pGrRJqMJK/EKhp
n/9EkQ8YPut4/99v8rwjXjislqYzRvR5qzgn7SUbfGpIxKYumCH2FnrdzSLfT4pm
rhFrwzRUIvPX4o+S5dx8uAFyV4f5TcDcgP0pXhxRFiXUqcBwAJJY4pTKCUL/iBQu
5B1GSfzYHwWdajfelWVInwlcBVSW7Y23eio/c3c68DhLmx/lbX371ag7W/BTlwtH
yHm10QUcW0N669xZLiHqw1394yq9YDCDpQBPOre9p+nNwPpEWGpJfsFR+jbL0rQR
sa3bYrVqQCx0FDlAwH9pgJVjlOC60olHY5OcweUlP3ix0SAxu4Oyd9Im3H3xOijv
5JDz0OUfBRV4AK8LTB4WaFh+LzqmqN7nE9mCRhgv8FI/iJ1iXwdO0o5kl5VanLbL
TOaOJRO7UtCJVoagt1vgPTdFDYyaLhYj38HqWEaESJQCHj8Haljlxl1UPqZZuOK3
u/3Qv3XHdHawWqUfe7f+9eGcGTZH40JFHudRXbWPDeJ3LicO87EW77dahKBD/lC3
ivffdPYDK0uspIpUHSj2eRUrwPWYLlapGAUp557oP+0/f7xBnhqDIe+Tl+pPrW8X
HVq0jt7VHLIKbQeM3/MfJdutW3wnT+9lKZNxhiPJcm31FYNKMtfPwwER2YB1cpHU
8zqkbH0K6N8+JYFvYEo0D2vS8Bf8qLLq6Di7LZtMoz8gjqr8lseA41QVnNk2XDpt
0BTEP4BHvuYD98LR6L+W+z9bTFnl5gXj8dP4YlA0O0TuuA7Z3n4IdolumyNVfact
7eb5pUeKpb03eDuQDhZEytQ6Nd3LsCysGAnXsGYYTyHgnPvSRF0ViqIJF3qa4ApO
7Z1BRhaGJBt06RtumrlBUnUO2OSr7lalHD+xxEAgqJeLjuWPQBQuybLFxnhZ7VBF
5UwByxSv4DGKs6mxP/HYUs6SXLsareEkWLMKsQLO0HwuT/hy7My+a5zKR9R0NeL3
YxkaA2eqvWUjSjGFbeJAMdWGKwBvh4fptuHlJwOZ/O8h+6+pRd+2/Tu+eyzKaA4l
Cr0whjEo71EXc+yz/iqNfjhJQHKUEZ/HZ6IkvlaEfd0bEKPIDFbgNWJA1lj4dBC3
Z4U9GjbDbv/r6tgw/tpDfd0aSp1f0x1dpBBPobQD9D7IA44+Ld8g2W/RBu7W8PlD
/Wg07p17FmRY2U63tZT/VrCRbWLbSqJ8jdVnx0BY7zNIDVZZH1fIjkDr/lhRbe5g
pD4TZieeTchTtnwTcO6v9REL1ozZsMOi9PlaiTZn7VV/xbnGVcXmq/Qquup4C7ee
xamHL2C1sJ4GZ5lnuFsAjA9AwS337/Q1d1D5QDx65OCuPFH6pI9jgMvnu1DqiJQl
9aCny5CcLjRaXzKQGMHZ8KYO4X9tnoY3AcrMVwMu9kVDOok/rv2aUhp1zmT+vfpg
3bRkZpCV7n54yEIIU/LXISCU1bgAfEELsjugqEa5m6Dy41ziLhEW8WLL6NxxgW2F
eOe0eyYaCF8+9o0LUqLgPWTJVcELKrwWA0dzDGYMMAIvwhvuzvAkLcr353f14Ru8
Q6VWySeDxWL0D6d0NdhwOgzW2fmwRRePxXFTHa1HlwAjw7IucRX7TvEOrYCBCePf
aWDi5mFrOJnZ7UwrxsGx5tJpEy7HBzespLx/Vvav9ZCJn/qDA+TNfT+y3xELm6iQ
7h52/ETb3bKzM1musn/tQ8HPvgpl94+SpnnXgD7AuV8cLQQE0cZQ5VQ/pEQleLK+
dTI9HWA05ZI7G7OpXCJWsIX0JfWRN41Vt8L/QBZJM86FWxGKMHeenjM3MO7S+N0V
hFHChpgHNJzqUPh52fR4nXUqUBbljLpRoaDzVZx0zs3Bci4cJe5LMssZFMdnbxpr
KM7YKHEI1YARzfIFCjpPtrQTWszlIXzn+Npe7t3rginGmfHRUINmWZK/qYq/UArq
H0ZxW/RPuoyBMZg44GRiDGikEjaVon+VBqp/vUii9AOcaNPGytfK3UWjHaMfdB6v
vyyPf3p+3vb5t7XZapyqdjqywRNctziKA3tU0cdfkZMcq1VxYbUaQgGh0BN88Qyg
oZ+fDgNJHcv+RhSUrlcg0qvKb+C5Gsm3LUHoDb9eUyvZ4jXB5Fav/YyoxjoypvLm
6ocpyxaPHmn9a4+MAHdecYAWlNeBq3kxJsmXvcGpYJGsEMHZ1aP3g69LHK58lQ88
2xpBk+g+PnV8XR37r/AFT1Ft/ChHO0vncmFrxUZcAvWQl4hFeZVJHsDb0hCOmUk6
3Brp6YzukFmsjADxjl+qnE/2P17EW58A4gG6cQzeHUqGZhLSLFHfNsNMjsBDBYEX
Eyyv+M7vKdKwKCA0OMX48tfrtFWj1TpsWQ66/nXkBQ7zuUi1bNTIlj8WKS4bnQ/d
/SiytpaNAJMLpXFazANFklMfwPol0q5HGLv5DgiXyehyhZOqyw0wOqlMG+hxFS0G
rSX2z7VfwtdET/EjmGS1F4G8JAtxm/vW5M7so+PH7mWbPmiHPfetTu6V/Ophv6Je
dgnW6EEHaVJxTD8T/NavbtI5B1/T/4UwZM+A7j/2aPVp6RSz2SCOBAZGaJSiTNTr
ABvnTG7HkgREzFeSiEVdd/0BowfmotviXJhVjZUJOGXO1Swj61itwskJN69OBKaw
TheBeCG9afsNHXcCoeLPXCHJzZF2LRPXsCTcV/ogSlxZcx1j5XQ8YRhmeZmWmlMm
PIbs/TOaq/39Cdu3G2UO0r6wRLRXFd8XztyQn/aGEn0JpRSBj4BgJdFbGnulntKz
U9cQ+iOtDebFlywXcBE+4E58DIKgCUulHnxi8iTlSxSMMHv/GGWJYe1jE3Xsvst/
z6CJ4ywK/0cqj7tm9/rnFxYsaBOTIkGyTYlrS7fVzscSYT/wKyAVMlCRuqKgvpsR
c7x0QGfzsVdasH4kIALR/KSn5qGumWPpd+TPBqAuRqFdkiySs+rlH1ikkaToXVLS
LePZTtgAU6/Vwty+SmFTMwWhHWWCcY3Fz/Eng58h4Y4UmWzAJU2e083WgevMthU0
2crX394l6iI7ZlreQ4eJrss5xF60aUNdso0h3gW2zXJTkC7EXmfgknJdQWQxZMjE
f6pQE31tUrqEBn3ZNmyvZXUr0SrnsujbqPcp+C6jPEEF3vHXGVPwaVtLcjjeEhCd
ifAQChZ9IKVHnZYkXyLvZRGOHjUOvEmtAw67wu1AiN8uiXEUA8tB+SjgnVUjX6qC
RnZ8FdrbnnDfBaYss+I3OS40vc3kE4i7YjPiYdV8SB+l1g9Q7JH9AggwDJirSl6o
so2IcIdNt7KtV/KwmBcl7/GZVJTlrDPJPYnV/oRrJRD/LWbFDEIM1heQc+HmNE++
k+c1cwim8VBWYZPW4izvkeeQ73LqYSDkd8nG+OKo4Afl/n2FpJIXTvguCNVk20J9
zEoKV6KLyC/zSUqTA6ac/a7IMx/v0TaN1xyMEEHlbG6EPn35sTYRQb92tuo7thjv
StHK2L22YgyvjILDMaGhBxlFWOKSj/IzbQPvMiS8x36diwWzZL0NeJL/SXeXQ1ws
l8/ZSIS2ZYbGqdQ6UGLcShgdgoSg12v5iVJBzr1v1uEcaMI8AptOPpSgRQGbC/y/
PgWnqiHf3Xs8DlL0eWQRckPm5ps70+qVcC4MrfEBrovvwSzsnejKUMVgLwK3wJz0
VhVf9CqooqyVIuvGhyvWMtIuhUgF1MIcCncxIvJt5rznQQ+cmxJBJb4z6WAt8zQA
SihucT1L8vdHxyqgMlTJGJyBHNGerCVFQVV++rWLILUMlQ9alNXyrc44MbZ5mL9E
asmeXfcVrgNzjqsUJifRb21gF8DtAPyIipCqLDNLzMQ6UBFKPDektEGa4q5eRRrZ
TEdAbIEKTYDdDwsktj9hwoo4pqETHGRmjTIF0iNbp/L/5HyaYCmH2tWf5rsEoQy9
Qwaq5dLv84nZGRXhA7t+MVkob7LGkgL8NHtd3nxvs4/Z74cPjj+9vLRQavGdlbbz
3AgZRLkSs9zkEFRufNxfaCUUaUj5Tg9vsEsaOD5MiFe5cqCdnfPm4KvMg7AW4EhN
qaoUeyvzfxva6gwvvL4rhZ56qfaSFFSnUrdQ3hQHuAuVt/WdYDRu/Dwi/Bjpxx81
wdY8CP0peTbh7I/zPU3Nr/0/DXWEJMfsqHGp3Y9g8SCPrfpOLJxW9rWQoO5mwFX9
+AV1TLsIpeP/zlR/UpLaWmwEnnjGrdn+mJKhNl4STucHHS65xK1xrZyljkF52ADd
1WWoIR3fexxaH6pSR+lBahIZSD74MYfpS83qxAYqjCpUclUCYDMOfV/dNuf26Tlq
+mD7tjsLJgj74mSk5WotnBnVJx2HjbaUdiUpLZ9oYv0Xx0kPEIHz/Bw++Mo32Yjz
n7HvqNcwmv2mc4hy5OXUi7t2Styd8rVODU+IUn1ZG8udllMiQEOtCcYVjx+1uKX6
8gzvvXk+e1YWXF8xbQQ8M+FaPQMo/fbvfXC9q16Sy8VxsITD8HPUL//dxdFiHQ15
XIs8Vm1E71JXjJw6IAhPnVUJZcSN4bBNvXITY84N8LMH7/l1N6WTIteEg4wgWUgj
rwST7iZq7x6gZppzMqWXn/Or74BXxA50qcfZfPi2Rf3v7vg6424etj9MmpuLRzYV
y957jMPeJnkEYGHET5lkL0lw7yt8z2L2gIVI3Sn/eSboqWYVea8PytOmKOzFepg4
AxN362YbKcLO81rw50plcKuOzh5RX1pTq/Q7EfBhyMpqBP5oPdXcWAG/wnmfnrYZ
LPeRRIBks0F272lOMH1SK1UGym39bPBk0fEOmKpme22p3/y63E0lVL2Oi0FdnSYX
iZ/pMESpYxMtoIsP0JZXDteu5OTd3HmOkfppFaYZ+sA9C7dlHlupPXWycfqqkvk1
dPnrmZNuc1NPotpVSNARe3/buw1mTQCFqMzKyg0PqZdG6HLu/Cz9tl4z8sUfwRvk
zj5wckkFP8Yx2QosAEgaxNKpJYoMKli6bsBulpL1WByYWxz67I2zQwYJI91kjnIt
sFeKuVTwbkO0GbeDueiP7lOCLufCnaIm4KVyCdNc+ULGehUCo3zBLUmerOn2fBcG
kTeBzGMsXr7DftxKbwSfLHSsEIQSoi9cHKs7px5t6mTCNbpp7x+zvKgvVw8eyYP7
PIso7MRvd1a8p5UMu5pr0arZZGK/hULeKThSoi0bU3qggArCXIOv0NXsrnV0E5kH
BARTJqD7RIE/l6J4gecGxj3XMsDQB1TuwOpwl5HkS6W+pzZyOIBOOksFWc8pkvYT
e2ulIzhadDbIbgBniSrDqnpF7PLPms81jl5tO5H5XIJzntW8BS5TLLa2X2S6e3WK
70wGReYPGavFs3wa97OSkPtlTQLekcxM5OL2aDowNns8RkC8zO82c6oI5n5Px/TZ
tIKRX3gDSDT/TpqY6bWue7NiPrm7dHp1l7hr+qJIuu1EbZ5LR+8EKr3zf/z0OZ6l
lcfJAKEfb/d7TQOQrrsjNJ/C6K4nmQNAKbZ0DKA5EqivIs7ob4w2nt8yC8N2Ba91
3DkS0nPb1reEF0/75dT2bMZGPTlFvTvJ28Vqk2M3OapxHA7vSmJLC3qzKxJV6BKy
Q8z4lttpzmbOaYMBOIot0HmN+6e/kK8AFk3yysoYzUdk9uvldB/6441eWCSv+F8D
1vmxowRb/d2GlJHMRdbYSRPPrqGHoOdW/9UcLHObfdontGCPJkw2Ci8rZN80cx++
rWgDr7Amkk1EULp+q2hfWXY9HKCZqXI6WbabyowHAWTHozew+RA6VG1xKkoJHjDN
B32MVte/FrJcSRLzjFyDcF7V7O38Izn8ud677YaxwtR+4064Tgsce9teIoOd8akW
/+V4zBl9iBMWlUwjy9ZMRIRCCMC60dbu89fUvXR5i/QSeMUtBFb+gBy1RSWwYXhI
CsHQMx25SvoLZWf4hTQ/JIt75pkS9zAFlAA30XIyPmYDWbzXLqxKjwnOPIPif2xf
E4rXHUpO8nJVfAgMRHSGy2dWO+QJsWH5g6ofMpKzIUSqTC/nmkg4BNzStyfkzD/d
NNOYlR2BXjkRFdBeMqJNvZF9dNudJsKZr28jGMADR/qhhgBeF2NFIwNGPwS0SbJT
N1BDg7KGr9+CZm+++h4NUWq3bOKhQnKhpOtIigE8aQtcyvFCO1TlgdTWckkpRjiz
t5Dxx0hH8Zq2MQ7b06qoosGe5uvBQPWOPMEAOA5LrTlWuMDNYnn18M2In7MIek47
TM7B2C/5DgwLaV02foMqqQzdBzUM/guogwg3jBDFBn7rwVWFyzKIhmEl9fKOgl9x
H/gYapttVHC889AaWfxKa4S68JVVYVeE7IarouUcpuvyvnbDvDmFcdmUPTMTI0fV
M1TmnzMFGiDSAZMCfA+Q0LsvqgIpliE00wquobPtKpyHpx3wl9NZJxpVrQdn9mu5
lSWh0+Q5QwzA2GpDpuj/ge4jBsoxG8/bCRNH4NdCkwPciM6HaJZovWLC6Yy986G2
AoAGSUs8YbDS+jhWFFBikw0+cC09WF7UxXxwmXBCmhjaDc1HmAZiKKbddZWz0CXe
sHi/39dqq9/ZCNpa93U7NBrBYocl16Bntvx33kQySBYEh6TSfIVm8LTeCq7j4e/4
bFHlPCv5eiQXWg56BIj7VLMt9jtRs51GM6hYVaCbLieYL67gbfIqX+9TlMTcQE7N
oLhLofjaCSKtVg086CpNK7GAMYLuCoEoEgcU5OiXotnZQmz08hP3Cm63npPimoIs
ExQXIumSkWWgBuHM5qTNJW0yneWEOwwLSLImOgVqOw8dxTYbP7Ph9AcIGNcyy3z2
iHnZ+Xj/BBXH3sURSTP8GXl2HhZcoudI+EI1EGVz0wyxlWGjvfg2shWAJDgL/m8y
w4LOGutBC8ljII6Oi+1O9jkq2zcucmdzqorUa7diw/vtE4oUoP+jLa/0p1kurHEK
EL47C/Tfqepv6x1rWJvn9FMrV1C+CYYKmwBDeZklOSST9g7DTJ8isIWVHGOXt1U1
9IEf88jURdXxrs5RdCGuiZgqmOCL9EwbCl8KUOKi6UhekYkyiUL63pDPGEVX1euq
licorX0Gt3mEEy6FwX4LQeEyzGt1BRCenr1UadD30bDQpOpj6IkS+cUIC1FFpShI
dzuT0k+BO982pahJsXeEBCgHFkr36ds5i0PepzteBrjlp4bUvVEG/5Aq/Y1dWASn
DPooBZNPF9o+h97sDRmFHwD0sAKwFnUdJ6PtJesC5w4N/geyCBIDDhjRSJXXYy9y
Q5XRa0DIoPE+74CX+qRtNi3dxrpgUAJMZLRLSn6G/Ypu1A/cmnFfGItveqAjsO3t
lQf2gnL7VM7DhM7HKHSEJdA3xbYWsKtZT+54uyysv1q/YwgHEzdEpKZWR76EUvkg
k/xePVTM0c1hXiN/+mawy2hmNIjx0PeoyTn/iW+gHbdRLxQL/uL7GzCtLVh7OTWd
vUku+Bb3UtU0LvKNxfWzJEatjMtQMqv40GdOj+eYBC1GaYVsjoxrcrwCJZOm6oGE
wN19LBAaNnAdH03rWX/ZpAcTmvLsAQj9cRkY3Jawi6Z6m16D19gbHYRYkpot4l7r
6CIiQ8a5s9wYS4KYqL99hV5hOgI2y7H5i4eMj1bzWWHZKaQdMq8jksdo9sy/QrpO
8YDIQU++8+/UNqfNuG1Ny15qsIJiHtzDZcHzMX/N8kZ9UzCoRlcRPG+wJNWZcwsj
ccmAdIeo9IvlK5kP2hFe5Q/9Qebe/L5pWqbtXVN/cC750cAgR10/KDFIEB2D9oEF
Unq9V9eX2i/NVY3mISYiq43v5Cyu5dKM0l8JFFB6NbGei6kgbd1aiN7FpSJbpJZ2
hShMyaIZzofCAqjAAbfWOIjeqvvzZAmWD31iyz86UZtN1mfRRPcDCwJ4t94HE+YP
iaqc1Fut8YY0iE0Rh5w6IbEDt4t5aR2BKlKWTKwaa6gEQ3N43T8t9KBnIDafGSJP
uwk70OBTQh2EYJJ5sdkwpthOfiwPJvF+CieSfJ1kUdnHK2zB3gvEe+V+X8+HWDai
AB3NckFH/idOzmoofp5Dvz5SK0EVYyqrhJdiE1xnh3kawgMfqeJ6qm11lx00328N
spSQbpr3uUEUCjlmR6hpgw6jdsFp6xzMrvpKOrEtvWGIwdSmpxqjFBN2HoSdOj0H
re2cVBibFkNf18FwdKOx4QGixEN45LvC6ZsMOZZzuQ2QE8VwOTLBRCAjG4KtibWX
XxWNknC6/HQDCpEyubTE/nZZsYdpEaKlqS6xuV6J81Cu3pDmJLE6QKpb3N4kkbLG
l4k5a5mXWpIpbKb2ErGQeWvam/qfEKNFZCPVOsUEa1PjkB1AYkxWVgnis95NVoPw
MlMb6+JlWhAS5NseGSnSyKHUqIDWgIaR+Tzuqpnfhsy4oeJr+o/3hYdBVLEuWPGM
kcEWpeQF1h+wstLdTiFaLQHsTQ4gdgZ90wqxOtvcA3AKta95wLKxtYbz02/Kj+V6
SkRUyMhHdgINUpbwr8pJbfke/DqJipBknmTrQkEQ35r0q3HCJXlneM80qdPR++u6
xsLKgAQU+TFv/y6abxQwTxkHpP4Ov4dRcK0cLEKiKyBlvUwU6N9ojj47F213/3aw
lSwx3aSVhFPc3CptM6VfDCTDOFSYb9r7bpvRzPclIf09Vv65S+yxDdGHmRvsKpVO
cF7CUYDV4ncF4v16WarKz+dOxCu9SU8JvSGioMi0rDYahEiJ2gtt9VD7UzKcl15y
/fAGBm5QGeMZsmnpBhjomS5Ce7X8G3e4f/9qi0ZZ+yMoUd7H2xYlC0NOJ8nsOXMg
hQlVvMuPHXap7w3ZjLbIDFPuzszWqRa0Gq/Gj8Wody+Zlw0sOSVZ3lbYSqm3/xud
lBNbWBa9mrXs6VQcPsK7flHvrNNGLwH1PvaA51YIhzkJ/E5EqeukwurXg+MDvZvD
0QyoepqWPglXfsZq8TJSgZZd5ypON7M5VJlOHzUa10osWDspzX+anVeEn2uWKY8g
Qs2ePlnWB+TLRg2WmjYEL3eGX/AB/5/ltyuVeXtC4nEABjZfZi4yXcKhX3z1ZVbM
acU6TnrDhqas6ph95sq9hS+JoSJB1NjRr1+U1/nlVotB47tw9IB9uW+3TWDgjQTm
TtUCtGC6uPelGtk7IB7rS6cmLHOKxRONemzecLfj4Hz+ALoBMOHezvMdMfTP6g4D
CA/6bo8DbQHOhOM8gKawET6L3eRqeNan9UGXFT3a3LOgVxdrfPQhJgJGMpJCK1+4
09oDcR3n1wA7j+39hxZXjX/8I7QEkqovlpKMbfR2ErnkVqBhE0stAlndB7+f5ij8
lnZBQEVQyemFe+ILaUh15rUMcL7To3G0Rmhg9IaOFk19wLMhah76Jum5JcCmQJml
cfhit9Ueyx9BoHrkDftNZlTVslFZyyNKyMuO1DoT86Z4bKt5qTI3VqT39nHM4ROb
0FCJ5Oi2O1iWJJyH+PxDKnSnern/QomeecNCWDPLfsEztRUxXXSaNOr1pnAKPz14
DhoPhvtlpSVsi+cp2wyU65yD5DYw/osdANqMKwvOeUbT5BdDT4ndqV7UTlGtN2lY
mX9NVjEAQj/idhv8PE1h/2wQskBc6rHgq6oZjsUevqi7FmXg9eWXK7j+NPhV+1Et
p6/cq5MCaw5vxoiMBt0pc8f6JEO8U2wjnae24DV6I7INm3i0/PVGv8E6U7RyEua3
schA0y5Kl9XsmEcA3ZRlXtTu6fHetM6sATvaHjpxUtYBYakQSYVV8tEk905IX4fS
4PqVWVyrwErSmjdlVJ1+dIDKuKm4amNgnVoUwpTGZwawnNZUCzhSH8Aprvd58qld
xoqgk/JXM1JiEbfGgwFBEhqzdzb6n7wkTI3/pL9zDytpMssXF8TtgEDx39hrb7Rz
MLgUw8hW/1QwkRUU4Ui6iRVUrTrBztEjc3MyOpcc/uk0hLv8Bzq8X17OkhI7+LWM
3bWLMnjymAHp/5sF7zMj7GmnfxuYRxO6XKIz84THRAW8hYrsCwnd6YpH1ayHpYEt
OYPNluRKJ8jT7NuV6I4QxEPgll+rORR+dLMcGkL1C9XtBuxQUh4wPDGsfbvMRyyf
tDdD/NLyM+/ItfmRrHrx7oVliCxKypx0wZgqzF3NZkRYeTdSNBWk1OlPK/CYtTE7
uOuRlBHvJ3h+XpzoAlshAD9dickUK5smFXe7HtrMejlVX8N1ub8UwsMDA+IqOhMw
myMhOS6Afudqg0PXpQDDQoS1/4+Duzr/G52q7kee1tgXFU+84F1eV4q9hlWAkGoT
jiVvJQh/ijRBxv1uwg2QLmIF2cFlBxHzOuHRsF3V8oMdMApyXJsZi6Y+ZNjJ/7fb
3VNyYp1Dyz0C06yMzAezJA/3yAwYUbvA2C1cnJHJWQQF3Feaw4rmc7pRFE0ti1Ej
HKGC/g5e1/Sd6G/3Tgq6RFQC2HpRxJDVa2F2LrhMUuLZKNiSM5ObehbUMdS8whq/
AzSvRrdlWYRKhTWq/ebe3HqtgmtKsOmEHecG7lxiEp+E4dgDGOrkPn1R2jaPAHUW
x69DniaTnrCKn7zN7CmzOBbgoF+unbr0MAIX+XQAB+xXcb3lLj3Xv1pxWolyAX2J
BWYrv6lxVfMjQTGfeFth32a/knkQkKL3/0ryvrzn7RwXTrKkF7Lxi1y4OAYVzhz4
1KrKeMorfJZfx+6EPHA6pDCIUSSGmDU0qYvZNXFgM+gbf6kCS68J0sr8VFsHzc9V
AOt7NpQB8/4zBonmKDPC1U59qmVjlNTm0LwZ0j9+pitAEEsjG0y8YcrTUdcDKams
DNyTmudrcPtNc3nfWPdymo9V/iJqU19gOarXEzgkbdwSCa0lKMXucGToGD97XFxz
WF/NUnjfpatOoi+rSe0/xFBj/M2iJ0vRJwlP3B0qhD9vCZO+cjJEs9RZKs1jWA4t
juzeOTggADTnmWl+HSZvm72TULxnGJ2MjvBF2uJ7f69uf3OKG8zqGyY1wNTvMxvf
T5w/4rD+lKyfZGGODBEP1o3gOOEzGMOdHdIvCBMsB3R2dHwyJP/IOgBaaGtDMPjn
/K2KUFvOA5WeYt6luYgBGSVK19smj6ZspA4CkkXHm0QvhSoiW+kRMsCL4SLzdqLu
188YZ6rPYfkOZo7eGqk28TtyooLP2Sw2NcTSc9aP2JqMsOcHrRIXo5YXykZKXPg2
YXtWYtgdyNpxfaDz50b4q8eUUWlzAJtj7dBpj6X0TeTq3YmWUHxT4lW6tyXJMv2i
pIve8Rjfir7SPMIdI9io5WqInb5UEPm0mSwDhoUFQK1odbpoUygo3EkfrAs9RX29
5XmGxJYEGOv/u7iKqrPltDFlUzHx13Np4aiUooqTlXAznTq/wl1UqiIqLXJGQ1IG
7iJNlJtUZnZwYFr3lKFCgHhu4anrRPrHEVvN74qiDhEAJoI8LQHeJOfc9Hgy3UdD
q3N8D3SzgUX284YzIxSxs2aJw/Xamt2UFvVIiQ+sK2bwYGPu0SlzY1OqbxQzQgW/
UU/y7xq8sc8Ro66Ii1uMG9iW8wwOkBS4kmN+g8e2Ne5jjko3oOF7Y0nlX1f48k3n
+OelvE4EcKeJtJcX3A8PHxQP78ZZM/5NiPzNFqb+DM4eTuEG6oy9IosvkzDX+xIM
blMhb9eRzWP2RRb7bQmJiL7QP7AGwUQwdZ1TzH5K3dELfFlTDa2vhNJBOGnhxzde
P8qIvSBENt7a9tqp67IAy55aGm3AiVGtbe2ZnRZ2Ezil+wKK1f0wczRpY+DTfNWH
sFOBACb90OJP9savA1ug34jBfsEqEvozU/DGfztB0cuq9cmQPfuPSUTQBbzpgMiM
e9v/oflEoFqxvRMushP6NVY9/ULn55bxS5sVVL+wuMaySriCPQOvjF5qgh/7s11O
3L5g+zFGqXxq7J1zEYWRBeq+3CJtcc5kn32LhKUE4KH2xqIbh4GYnLR8AVyZLiOC
sFUDo+ELQCijaQv0iu1t/8fPbcrTzaMNgklF305FYrn9WasszzN3vUc/BGVkggbk
UDOQzrBE49SwYtQo5lC5E3WCvtV8r9VxG5iD42xE8gVZOZK94MzuqyKwBx08S9Uq
joETHNMEaTDv/7p+FZLd6TdA7LxeM3AiZCGd/8/oVX/gLMZcfBuGayleXKMl9TXs
1gfmIHLZ86Oua4Kmg6Hqa1rKdHZmpQrwQgosTnuTDeUXpBf5sHQv7IuPwHhmmIid
Ft7trigZr3sl+EKPsIyffAHO9cJcWDaZ5ltEkgnuF7fswYIkXuPChsWklhqqFH9e
J9B8FxGS5/PMad8MoghHyPj6sK1My9QGU1rOKiA4sgry8ANFigOpGp/1V02HXdg/
yuh/ytq5vdxqgceo/cLM79uo8Qhnf+YL7GuCbQDWFc1wT+Et+shNr+XmY2Rf/SAC
uZRZFdFIeLUeyEaSz+c0BSwW2blu3NIKH41X9CknpGwmWUhTov3E5wK+Zgi/CRwN
d2MuTFVdyv/OBQHN4mjluW4BDfRCAQ0oXCzWtHz+7r9XoFMkRo0eaS6/QsVcaVpb
URjo6PJp6soJVRlNRLClSS+vgatAanEEymfz4J6XsWwUybq/LoxQ+wsYKuMQfeOv
8CCe9qt7aE3TNSKTE09Wksz2amsIue5Xh3DG5B8ZSUBIgzvDEZfGcMgF5+38KpYy
8yZ09Xl+ZugzO0nqbRIAxo9pl64q3Fdri6Q5CkAxGuB1D5ogWdi7H6vYa4PeVQOt
lfCuYHl8rmqHLfrFl9e6o64lsSBlvDrYC13u06gpe4iMxXXvOTe6OlOHRz/yt4rZ
vzDPfCgXb+Pl5epheJmgcTm8UZNU7yr7N79BF8lQSB7nrPJSia9HoRGf5h5UqsnI
9BteS3dzF2JULgcuS5TQ1Cisj1apisVp/2787Ey6YffreMg73PrC2p4Q6Apdjm0Q
457YbeS4gS78jvexD44TZmdmwi6PR26d4XOhHkdrinGuGoRyKhwaOspqK3uYS4Ja
12LTsxyE5wlJQdGC+NATXqJwYAIZPgUvz75C498kOxW3NDBm+0pjpHra0zxG7Opk
THKQKa+jVfkYoul5dr1LcDvJ730nWdisSJLcgNUDn+gEKrnB1+90GqD7G15ojUP+
DTWIrwOAJZOOa8O2T7PDm0avUrmPV/crSkmSOtdaoxuRik/zjM3OlJ03eBIrNZmK
B60J6ONdeWCbmxDvI/MIYls4jzTBiN+RNjXToWQd85hBuC7FubdBMB2UDHYfqoxO
EZwznOOarwK6xlEsuGm+VLNrhYziP/lrWuCd9S1xRdrxh7qCyJi+SLPxR+Kyv5KY
V10Vat8BEWDzgSNwf2IxPt2RLZrtEFvvAH0Vf/Azh8vihDlIUkh0CeCbFkUZi4Ue
S5Y5ERlq1WWz8RuM7U4r/sm6FxspTancFX1VNr8RxODaBtZa0tHQZfNXH9AYD0WE
QrfWE4HmuZcTbwxD/4bRogKLhXX2s2zHfYkJQtHkwxDwEn25HLLaQmgQyV8klkne
PWCdouZfXQrLTznoMcVofRmUmIk3zocIsl2Ft5TPDrmoBhfLidOSBrY5BnrMmKbr
FiOnLbCqvxqu15ewqEiMyS39CE0zJYNli9+EuwzmyEJ8pvvY3Bbj6A13Yakmh4hA
m+0PRKhxlzjW8NAy0ADEGRDtsVQ4yqxi/GBAskRWb7c82yl1FdKZNl3Z0qPAFfa6
XVlyMpcB74gW3xGBDAq/Y+vfHOfwT8je/z5yaQE7PkpSjMQ4HQRO0BudgYmGcWKx
4EitDhgYQuwKfXhuscKodrDY3AhUv+f+tzFtLW86u0SmPKq6XwtHXOIGbGhQYqkJ
Il4Iz0IZ8ipE8mXXpCgYesNEjNLa3+XRt0R4FcO5X0Qj4y2i6Rlk68Au98jUcMvN
lDLgsKGesnwtrE3aYLGXun8GnKAv/lBTFCV5vBthFFN6esVlSRmj5S9WhOEqFaWd
B1RJQ6+rqYIUtLzUwRs3w4mV+DGxRjcuU7LMULZmPL5jRHPuaphddoq0Mgf8FKKk
xwX4Eex/oK0vP/6DzNhlBfh7+UiNltCLPNEpNSRDpJap0W+lgaJLebzrE/dVD5UF
ggVh1/N5bKf+oFuKoq3zo4i/h2g3RBQBxO8OESMPYUtZZTkclZAC5UryNDnci5in
0q7UWkTQ96DXx0Tfp+SBS73Ko2U90vzi08LzJR02Epyirwx6lpJMY99kYxHd7CXn
CivLwoFzaoQoDUN7EO5i9eaU2rdNvwB/JJNs9iZ1tP887Ll12CUCD8WfGk0jigAB
yoiq7A1NkNrL2AXVAt64l4cC/2RzevdZRCaCU0GWweFPPSBOy5Zgam14K6cSXaA6
FHOKtJNVY/9RcNSTWOROdEYh0bMfm3I4NG70RZwJWKcvuQPJTtgUBVmM3xKenHXp
mrflRUEdn/mHMSHWBV1YoBBcGA0MIhwhcVzY+Xrx2gXNQWQuMv7XsodgtzXVy8dl
W9jZagCfUV9yepCzY0mOpr4lQWd4BuabJJTMLTAvCqax5/TJ9lSp748Yg7r02QDT
0ERx87lfOBhg9QfxhwaARe2RLccYXVntmuU6pj2quAuK8QV5MAGnqg6bOCRv3IzQ
0N8IpUnEu9XTabkSglqB9bSH2zEzS9oAH1cwqGj/dKS0LmDOEajY7f5OK/yELDhv
Cvu6lKpy3f+cIoLKzYl92axC4lbQquUKAwgg+eDlHawv1C0bYT+uw3EVrUH/3sJG
EiMb8JZhYtfvWcPRIVsI+0BauHLLuxJanCqkyHuKboPlntjzKWh2QtnKopg0qh0t
Y8nNTvWs+flTpNi/9dZLMwmGnpL+gddkuSYTxDhq0Bm01ZHnEucX+T/KDhxw5Pvu
TYmyG6OINZBqpTKhfkl7lqAcbkx7dLmYEpN2h8d7AVnz63jve3xLgRCsaeIrP0iu
zuBMMsxEfJ4rgTGJ0htKohSlGwdtXhHFsJa5qH+zxWNPf7x/guTpqJIdR13L9fjW
BzoHUw3/9gLz6zBhbIBeH/ck7PQHuLRfHtQVs0UyygL6M2PiqLdy5JwJ170oVPqq
8c/sr4VDo30I4XQD+Ya5/jMuCzxgECqgiYW8og+5THCb/LrRDvr4/MEQsxS+Mteu
io5Y3JStFWbyl5PNNGRwVgZca31QxmlenpyFDgHIDBZbMuLwG9Jf7xVxfaaxsAI5
UncJFBLOvj70wgE9OCz1us2cn888IKAoo0ZiN1mskwKNKhoBKh/At2/36daevIoI
8bUrmpNQME/M+7c41AfwQgRd8gj3FlveO2BpItOI+FRHDJYGfOm4cRjuNlIVZtOl
+iAMQZlb48tOOtBz4yX3NIk2wd80RjgGKv5cx0if9+ei5KB/RekRPdqV+SwCgj4k
8xSdHg9CzazqNrrasc9D9z783kLcTKwdIv6q2Rru/q9UHCDRqmkGgl84lxvDs6Yn
8klAriUSEudwED5mpiL+rq4PQC5JBtmoFp2pA+pUqL5JHcKhpjlCuww/f7OSiOHh
9rDvdwroBWYc5aWQqqU9kffOrMEuQ/3zykZv7oN08gRNiHnkxNFoL9tzHL674c94
3n45zRFKW2D/m0mwQFXEbU9oeLnxOP3+w8kgUffG/mHjzdlNOvd7dURMeimorr7J
um/XCB7tW+DsT4PVS4+PSDO6Pl28BQG61g/GWY+BIN/5mh8p3FL0kBRXtToIOAr4
sUqUxe688Zypf3C5hDU5gyP1zLEaUr8oaTzCDftpxMIGZ+9WYQfftDaS4oR9y9Vm
1iXxKQk3JTwwumx5iugRElnYOG4NnZ/BP5AbRjJKY9wBciB6HdAFNvtEQVxjwHeN
l8BTlWmqXGR9eN0FwdlhtpG1mlUwgtcB/GPlS1XtP6bx1ju5tXG35WKbjiaY8LQh
EQU2IZTppaaPJiZEdeN9cLnwH0s0fX8Zt9L/zaXZ+dUBdwh+5xAuYFqDfnR007N7
n0vBW7T3IDd83zwbENbtVBtBgTIgQXflR2lPSqz1Q/7cvfKQYfujf6bVzy5EZtcb
yLOWX6iLj3zzcle0JmEvQNTtOHYlYQN2r/XUgh+UQ9dHO5RZUhZbdk7ZWdQ7Iq4Q
KMcZaQK06M126On841R9DRWVOpopbnZ6QZ5lYQ8nBlJJg0UXDs8SMPzNOupFYUhE
44xhHPGrbdNVz/OXuVgPk8IpMhGCY0rYvUFW/O+1INp1IZX0l7nV9I7A4QqzwWBe
ji+7ooHAO9GwiB2qmkkJq72SRluyZ9SyKzVgkZ8GFogQJEXFb8kyYhwNhlAguGeG
nPi3ORWroSuPbZiWcmkzZUAtb7PylxS91NMf/0FPAOLBqnpa3u7VbU0CmsLVELJI
C16IB44lOVqm/rowf6Ody3hmyaxUysd4vaX9qb8Oo8NUWn41BxjwMzLjU7iEJ2o1
wB6mAieHXCycQTuWzOpZRqZxYPc97ACJnmkAq6xbMd3voj046tjLMSgRhhih72vW
MLV7OgrZVYnQH9ZnQS3Vgg6E7txcm6vQnqAA0K467fAsLQfhRI6WadU3WpTCJ2GO
OaeLkuUNVHUpHTS9tw76Y/TNf3zabHLJurrZiHeO1/4+oreLFeceXMU+aoGjaTht
isi9+Hk+KF6fDBgGIjgupW3SFfUNfX0fyLD/ayoLfyw4n7NAE5B3r4T3CU6LIjYi
ATb/g7KsxqLOoQz40PdCzhMLipXVHarzgiY+GTaybustnIgQb7QHP4ZBaC1WsNw5
5yedNsMbhQoXWledt1PPObCZxTIaDOJSrWM7tUTkJG3nfh0tFqjZZv0gI9ZcNT3Q
57zf6kOvBU8xYyRmZn2NDQ+FCVs6nFo9hIKw0V7w21kvgk1InAcQABu9rWhvn/G2
XC+JR06pWr9STG+HxkmQaLvL3/PoEmNOAsVkOMbqQsYsCw/5I7Q7dUYptGZNDgt8
+smaSRvCvOIqw+Z28pJqoWh08ePUph/2JPzSHg69l98kbI5FVt3+fgHcfVd3PIgk
RUjI9tuHt2zlDHyIVb/j+1UWMKE/bxm1LmOZsWpWXebm7sr5BRwsdenORlyfe69W
7tk1jm/0x9+vQe+qfSdm4DfTOF/dLcBCJiYCuyuXWljUVegs+xhe24TYL7CIhDcU
pQLsXLzy4RonzlcMqy2BNz0b7ow7oYRw8TACly9brx/sDQhNwJF8+yy0peIRHngA
3pL8g6gj2fMQuaGvY58Rxf9QIDK9pds5uQYzXbbBorDYNZosU6cJ3LHDcgXEIRcD
X5j9/7GpodELKEEvS2DgwM17rL0od/B9xgOJqqIkFoYN/jTr/2WNlV28fHzYJSNM
3wEIZS9pca0DkJSyqkKi6aCscV/lvNkWN3rU6/Wt0dAA+YZyj0gUofMbARo4IOTO
VLGVSaWLVHCMrNmnHBRUm55taOJQLOLTgwuUjagDTO6w7f0JC6mxBzo9yOX6PEXD
cXZvRXamc+l5K/9XM8GslPaX0pZbm+QL6BQmiePGxi9gIF9YP9raEjdUY/c14EQ6
XmFK0bRr96UrzIMqFeXUJ3wCFaxfxR+3PPHq3IKvaJDbQjYsXC0kph/8xICyxekB
Ypx9hrniNf3v5sfD86v+thajP9rvVrEauyZN58dfXl8TQsf3GIvLpGIGoRKeQ5Ik
4daGVwryPzPmSzohJ5elDJymBcdCxMzgkdRaON4edPPOvVHK2nwdhq9c05jYQv9K
BacAKGElsp4tQkKcBqDpODq3rquUkz1P+j5Vd5WrE3vlYFYm+xTDIoyFvEoP5xM2
w78n/UIuJ5bPpApIqaCSo54+bwKTkdn1pNNgSThHfImZP4YogBPWnH8PF4vXEhn1
caOUKAnK2bKrV0qmXGNP903p5OUUK5zAbjGaq5dL2fM/lrNAlKuIJhGI1x9RRHNa
jF8dukghtgcbN0sANxEh65oaSg5n3VwbKnqH7rZRouBkHEoLD7UUGLvVocwKvUGu
p9DcS1BF3jDcx9mdFaJcjU3RiWgGhLOUgSwnGgXbHTiyDtlpBX2o4ycACAQBnhTv
bnS9DoZu9sp7Ht5cMZxNexJbEBY7C63BMHzqylPNt8M8X5IENSLuPX5ZQ/wYSq02
2kjmtqje2K3R2/lkV3F2mTES7TZP1qMJ4RIymAdvNTaFpOuRbjUJlmJLF/J8v4K6
hoCaWnrm0YH+lzMLkmAPwFIy3Dbq62pvJupngXNehwZP6tDKsy7OUAQMbftsKY1S
jJBt4vveCxWo48UGA86+oyJMZes4mwRZMOLj3yunlgmZjWbPXa0526jxja8hM9bm
qm13TQ1UMh61LuaSZ3EVh+M8F7X0dAm4OioJz7L4HVmDfEv2aadUEmeFsuZJNAj1
vhHBFDnbhmd8UztVVy4+RFxLcx6WluyYZCcmzP/az90YeLDwhHHXXThEpH2SfluL
DiDfe4s8PNh4ACbc0YbhNkOCjYphP6E3T+6yTg3kYkEoJ/xQtdE0ag4MZzFlEHhI
CIU81ru6bjol7XShTsHU3Z9RTJNCFB1e7IoRu8xirnwG0r+pkA4hcNMq1I4T18xU
4Cd2F5t4ubArc0MgUpjNQQJsMgPEb6o2EfvJuCP8lgglPNeFPjVn/GoYVGLKfGC1
AhB5ucF6myJ/MfEoaDp3PoqGR0XrWgEfYcYvjn1IlAtsk2Sxg8Hx5sEMW4u1cvX2
PMWSZ0SGbNg3LXsKnCre0/ObsHXDK7wcPn8WW7JhXBAJspLTDh98Z1HMNmtku/qS
DZSYovZKQCtBwEBVzXnb1SBPZUnmKYgvhJ5GDU/kCY+67yaEIGbhghTHWqbH8JJ3
kMu+KP7NJ6v5LH4S81d8UsWdEaOXfpN9vP4aDHm745EnTLbUQcFAoMRg9yj12LIy
qNhA5Bdt9kg6obz9ARxTPOSs8JadrLNNa4O3ENITYnqGIU5WTCrD2KNp0aQFCWfn
NtHDlgUbN5hhwPk7qOLXLKzJb+tiqf3rt1fy6BJTN3dpC1K8aGVPnrdBKTLfZk1b
/HB1k0BWeSzervZCZ5oEjyLROtzqoRMeC6yUU3Otpy8jHjhsOgRWCIRdfXlaeg8k
gBfHAef6plPNtgGmnt4FhsGzy8+CruYfMJpF+L9EZQ/9foQPliWXTnMQWgWekMa1
9nbmrhnHKnY+2SU070nPfVA2r8KD6LPs7sx9bnqiJzWvfI7PLa55hG/y4rgmLWL6
bRHIBljF6LeT8X757W3tZpcEFd926ku9mZ5XYXyMVcVJeveUEqOk9VcaEVY3GO3p
hM9w8/H5dneTAzDBNW6Ko0sMqmgGBzlAEM8tU6Dx+hvfa165F/XB//KeE6svj5ZK
H7J/g9P2heY9D0fGOsLv8HxLZcGk6EDZPJVFk8ozqIa7OZxGssq5pj5kdoFSmK8e
oxL4wad+TFb+oRIZ7VhHdXmyL/vhDsvgx8ZcvWuP62/QnMz4KzYy4HmRrhxRtHrM
Tx+boKFubhk9rf5zBlAxmVZ7AQXfVDqvx0KSjL2kn94a2wQz2lsJUq2n8pTRKUlT
5yoryUYSYhAQ3RaVMeX30u6f1IxltDDJ/v81DEoWDHat9V+9/bm5f+L+ksGZwr+h
r6NASNfJEd1UhdnvemHjf3mV4jEsrL4ICs79wfYU/mAOgJyPY48PqCQY01U0wiv0
I3tcbFoKK4NDrgcxlb62HArxWDjyUbWvcVbTmt0+17e48wU+7u9PGxsHqeHcJVl5
zTyRSgKnSzn8g72Ajx3JnZddn1whKfu/FCKnhMIEaWkETf7NqneAfTVfWJn68TZJ
0r0mdoX3abZrHauU1aoHvmfLnwB4s+BVLW7E0zUa1w+FCrELeHpNI3NAaUg7vKY8
UMyltbHhqjUvwiNpmShccaLMWoHGdzgqlsK1cEQTsfusKBcZVveJ7CtNQGHBGAwC
82g+zKp5040zoPQXourIyI9QSUch4opJw7nlBQ743joC3zRUzLUZ2jQOOmPR2Fro
E9ow3fxNQW2P++8FVqQ3ZYiuh5fXkKRA1BCDSmbA4PAign7txYYFOUI2kp8du1hd
iMcld+Fi3dRDWsfbcnAzM9HDFhMhmOLfomUw0bDxWSwcoMlJMri+QW56Zf+q0UCo
VUiW5fzy/OMnz9JL2QwEcLsx0orQU6nuaYFlv++GWbPYX+bjLd1Lsp1fNg96ct40
gtRxfy9uhopfQUDJy851t29HZEkFib1QTxjw/8WBGNqIWdgqJAh0sYsCjc6CLz5m
yQUYE6WKSyF7CQMv0t692n6yGV3iZ/wDfpua7lgrIAG4N0ZymQlvg5Hsax/fVvTe
huI89uxq8eajaAUfzGzsKPGDggw/k2m756BrXPMSm+aOYwiBjYAaXBh2vFcsWT5E
PJqbI6G8l7Ln/yd3iRPGk6/1lSF0z28SGrYWIYf+prSKlnJ6VnVsudafiikOnMcO
dKPtXRRnIjAJfl2e6T5HPLLQHDG4eoi4ElKvr4o5xe9PB0VVhCkCqrmm/qQ3Tlve
VD2her9LZZkcE9HMOE2Gj+tgYV5MfvS3qAcTvcmQXFRs9qpo0U7qvvuz//Exzj7n
s+Xjt3ofGmF/6aTXzmakE7YP7yU+S5d8+MhpBFqZKeKY5VDk5Kv5GBmqRGEb+nRH
QYbBggF95J1lig7/g9+1NpgPQO4yTTqKbeAdV+9P5zNCG7Ig1h2+JRq5XtEl7q2F
e95SyCiXD+bQZqSiiKrjlR33OhwemvHAUgfOJYctV3gx8wvCT56qWGSZuSM8u0sS
PlUSdKKDNFwB3p/GvtiRxqjzztQut5mTY8WdGdUuAcIoUuzs/zYLyZSm3kgIDJT7
sWuk4agAa+46PsnFDemucdqDEZL8sYcIpOsUOFEaLlYNZusK4JMGUzGglo+WlUtc
IYyIDFgEpOA1v4Klo2Bt4xgVJVpHH+jejWMtNw3eAIbadEIUCEShkpryk6zD8nSa
qtXdb8kEjU7h8zNW/XsBGQMOxCbifO2F4lD2nttobnorsr6B1z09m8HHKdp0y1Qx
007ue1q6JOmbwt8juK4QM0xr0+sPtbFCzwF0hk+V8iI0kM3acBbEXd41Q4JhASMY
eIB4brw6LG4bwuZK6vILQqPjcEAgMPQnj4FMMoCn7rLf3LuWtGOZFUK2pO3RLv8z
KpOMDkT4qebyRd531pyxU4zILv5ICreNJyaq6ySWzxMnDC//DSIXtuiysBasYOy/
XSQoVHKDFEygzAlHXXg4gyrUC8AVO1AGyY+evOr/D/DvZluhZiaXNGScV4XI4I/P
++Wl4sOTHQj7X6OlOPdxevZpmbC7cJGwdjKyxeY28MFLu4rfZoQ/1ZFcwrak+OrQ
2SzVTMWgmqcOv6p8/0ySq/2bCExMAPjy47qovblxZqJ5ddt7eeTHs4Pocfx/y1Jy
Mw/HTQ+JGOQVJahXw1DyJT74yCvy6SQsygyClyYLgVuYvaj6UxbWz5t6jwqSa/Hd
NEFXVe6r8b/yLWfHCyRF5+0cyzuLYhU94kY0lqASZuAmGxN5F93yOUcM/2ezTjiw
JH4YFQIexVA2523PUpd9eDpJWJpl5l24hMZpC4gPtFB79kwnCQXY24A1d2rtx89c
lOixr3i4CdaxmPLMrN0cbyouwadRpBmNGZhm0T0O/Vnk+UbuLZ5C4YyWdx1rwOrj
cnHnh4bsbCrWS0jY7rNkcJexeQRRf7XNwB1l1+UaKJHC2KBIhurDg27TM69SPw6l
b0mlokkbyk2OvQJdtY8Zy3TAY3AtZCR3U2QRdgrHrjvM8l+B6SlfoazFNM5hWNrZ
SmXx/yAh2a25hCcv410GMJKCIjFMiJ2lgUgXpf05FpQKg4pn//9BN8KroFlJBrJp
T38Z0BcIAFG0GKStiow62UBeTEJSzi9sBXkm/g1A7X+1r2a41gMCk5vovVwZYTYo
JHssrZwSCybLfVsvvRO7HaAWgsykvNXlgsDIpQUkucIdN6LzrtpGuL5M0YYHSbtu
9wEoBsiOFgAghfzZeXIeU7gYtjbeDlyr7uCYuKDnTuAv9qN7/YhErXW2GoJeR0CS
+ziCKXsJsFglv2tLDtK82eXTrCI7a9FWsbmUmnxqnJ3Zz/XtO+ye0OQGdA3dyOwb
C0z+fZpnJ93LvgV2Ju1Xwppz7wx86Kfn8uTnb460Rgd3q6TVeU5fRUdN9s8ZkSVU
KpLgqgTDObWVTAUK+oyYYllZ60+nx0ewQAPHy2pxWfXqG8ibcpzFLtXziogA5bZN
ERbEls0qNBwoTdBPCu07BJj8mqErPO6I6yHD8+RNe/Q9QR4zsEv5nV0gxeasOsGh
2WTJzqupe3GvT0KOrKNkzGAfQsDu/QkXZss77y8yQGDuHUpw7HnqG/VJytuEz+3K
9ig0DIdAhz7vKmSmp3pcym1sfH1pPZeZ2pktM1rJ+67vKRDWeTnnviJIe8WZemm5
4AY8LHas67y2gLjzd2BdESmpquuqquZdRDtPMlj8xIDftItBdPPjG9YMuMSWkV4Q
yYWFAnjImkr0pzWqdrvOqUU5ZQPRN0qFc/WCv3fNDZWfLTx8xNydwJaxaI7HRYVt
XLyFxA8Db8UIbWVT6phyRQXBw2FWBS8ZWMdUHg1G8r5m+NCuRpH8yecWwmQnB19e
dEW+B+vG/byum3Wuky/SMPkeQ1Do9uKz6eSFuKKu9o02Lfbznfphj0TuSaDTJRja
XyNn+eyLbPFsYn4Z81/UpasK0LeBb+ocdoekr+CIk4F4TOQneAJkRQNP8OzwsmHy
4r1qvxzcCqHetQvl293PD6bmB9cnFSE7/lFXhnSMpTP8NMm6kyZb5qKvXhkr7ESf
n8dGYyzi1heg/t7wyR240eHS8pPWh9ErRgdCGS2say+vO2SbumNfX0XyLlz8vFIZ
IkDB/zNNjNBKHUwqel05BaPk7Y8RpU3uWsUEm4i2Qz4WqNiKX4hVvjM1gN63Mlql
h/nBfsYIescUHIWG57dYyQc9BcZw/ajqeLCP0BgwODLzvWHOlz5K5u+sRqlwO99p
HGSm9n58m9mZ2tOH7ei+UaX5HB2ITFfWBkIvKOoWgPP/7B3PmIe2ukrCa79R3jw6
yJsSgUhgZo2emx7fugcRCeoC52hFYHM6cyDfEW2NMlzStYGimU0lkZrQlCEJtvF5
A3yUBaJllVUWgh3O49+CGlMayXJvEe6RXWW1VAQFXP5bg5LgawqWnIKEX0W9pvv1
qJOVBpTvdHuwbjJxVKhoM3PyFX7L8zRVp3koIMPa2tGmgy87oFOe+2aUOyibLIof
2YojOSWqBVPNHM3epbSsYJ8y9iTV1ljfONDQ/LNDBqClETkFLqQBi+V1wlVGxIdN
4Ae3wwk1q4e8/vY3JRT3GleUspZIAksR7Hgz13l9vxO5iMLjMKtLj3ZZIr5jfb4Z
Z6Aar/QLemvMtSUq7YWAoQtx9mg+pMKTceLbvD7waVcG56oY9Ylc9ZAyNKjpl7us
5AGiZwzXzVPwHxAbXk4/drLl3u2YSuV7NJfyXujjMK76qfup3M7DblOhRWIGWR3k
u0scLQ1gqd0RSNsvzTSbfdkCEOEO26PYnN8bpNO1ZUUcHRofrAN2UXhfsaVlmv41
ZgQUCAfmrr4R5At4ws/QsHPSq/DNc9lfo9kV9NsrZAjW1V1KmgFZnv4ZlRXteccd
D1Qe3PVy+gHeI70saTtLUzETjCLvEAtP+w9A7wwqnPFUtxhB9lJICPwlODoFZCEg
RTjnlM6NBhPfPk7yE1Yjp1r4hjaePOEN7KjnS5F0XAIjp9uJgdunACQ5+QfCTMSU
NWqbwn9lQv3bLS1RfR0zOL2rncKmb75mBLDiyx/B38V60GLA1q+wyrQImg3CUQfy
qG6FEGdEnLxqJs04/gxNzb+PFOjLdg68ODtj3pXEeuBMZcD8gNJJgxnRrIOKlbS2
7ggaPu/hVG2X8sIVdbLkcqkaRTnFkkeFFSTA3KDI2LtjWd/9eH86Y82SVTfMQUF2
/aw9/ZPbNSL7td06y+Gnl01hIN0mmNlgE04jvG3D9msskGKYPjMx0vXtHScn/ew5
3+K3PFipCfC/3vDtph0dPWU0p89Bz3IXDFEly8ytJiUvp4i4GfWi2op62EY24h8j
VWqvib1fXbLIzZ97u/JqPHBS08UCYa/26No41gJQb384ufcspE/seIu36IbSqOp9
CQMnfXm3AL48e33NN43/oDHwY00dy64FqEqBzbt65G86Oo0e4bycXAjVLKPrbJrC
OmBxm/d9AOKfs57uuc+dlLZSSDRz1P32Zusc2Wwq1Jrai70QWELjkADGSjwzUTCc
cc+1/PnqdEn0suQySZQ1VgfCQr3K8dQ9/i/2DFnePRLYWOXooFbKpaqoURsuwQtN
EJg67RalKL3RncwIbyR/uZfDFuNsh0v5ndUoSFoV9Oxc5B/gxy0+CIJhCaHyal6K
YF2JypGlekp2VqcRbganVirb3a2s2J7DjNexkeUB/9qM/aTGJ50tTEW5Qyqsq4fH
QVBVZQpGYHZWOHDLnatl4zFLIRFRNeLpy1d72SvHcv/aRRWGbIDVqvccybtL0Vuo
IB7NCGIAmlVhMOdRM49qk0qz+xw58kgQbBRVUftNLH4MZkaD6sHfMn4N6AaS5eNn
R05Ymji8KQ9wuGKOfyI+MhxUxxLLXvG2WmD6em0Vb+jQuf5Ta/qa/3wubI0lePCM
A/VIRBXaQUf4E+NGw/Kv2SiCOzsKEOQ0V8CqRSlZ6yQc5wI8w9mqdWIXLL1KrA1e
ESjFVmo7YPRsCL5VmOVyKunusS4MLAXArPu9rfyHZBJO3KvH3Z1fA0pgMrFRIWq6
8ZMxqiIPzeuun60DHL8f86Gp49t2+TC3UHudv8JEYq8aFI/RzkODHMEDI83UREnf
UlvX4EzcI0B0ABqEQiiEDSO7dhBeuL4GOHTBMUAbY49Ph3UpDIPW/xlWNMtybJ79
0skpXU9LEJvUsgbIRhoFMHxpKrG6EehLo9ReJ1+7Ik6W/4omHEfHOWKj3hyTbnsp
GdDsuc0+GBH8z6AZSDsf3co2RIwmlHOjDND/4u3ymjV+otLxq8cCeBZTHbsTZH2J
Hx3u5goXZZ3xfYlVzIkeM8SWLQgavaiTrhKH33sPgn81ANuqfLJU4Zxth1Pf+KR/
/G6PYV3lPeN0IqiUuo6anW+p6v8FVah9PCgp9qWVzuSDu0crvBaFlnDiiyw1qkog
k5BCOmiyg/tgl9JRtEFsAwbeGprdPS7MostY1FGlsyF4PDUI0+wrqOjf28Ohhlx3
sE0XghQw3u6qOcb2B3+jcX9UiLILRhNMrNaQGEg0Yj3W8exa9ZL7cVYJ0sUjqKTO
Jnqh1PSBlFepM9COrgB5+96CgQqNXJSC6ZnY0I8D2QDszC3ilvUOHx6x5QbnJeb4
EZrdb4DuamqiGJ0e9kEFOtjSfWDzR/wR3w+Ud8V56ve3CkB74QbRhCjFq6dIwkmb
opdVRtwqljGQQZVGaLPAD5luqAjjDEkc2x4bDYvLiRVm89WijOZwLmh6WrOW4gw8
bPiNUV18mpod4epJvXwTcthi+Wt6NltrAUsDCr3/XgfFdR7hAMSL++dgQuV4EP5q
lNfhsJ4ZraTHgKSmfkxSoDp4nVvl+NYGc22TLCSf8+HZpX5K/QH2gH7+PsRKc0tO
5zRegiXM0LSI3gk5Hfbo4g9dE4eTsqrTrlyjGrmRO6qv9gf8rItiMSNMdj06E/33
KX96JLQCEGhy2E/711Bkryn7RIOm7rxzqGZNZCvXPvtXaYn2YzeuvzLQmhW5v9jw
fRR2JEr6OrcGz2xxDd8wCu0+I1A6aeT3QL//YthwVXRJr7GPvdcZ/JFfsuvyhYI4
yK9Cgs8K/wK2GQIwOiekVo9TXsVzDgvsufVnKvFO7UVHyur9tqcSJ/bEX7a3Gak7
+Q+WiRDITMQIX1xDKzCPs0e5jMfY9BhEmVOgVZjyIFv4qc7CaMPtxZEo7gc5fpKo
tsfso+puS+KqaIqZB/bLqAVOT3aYE8NTE5j3M3Z24mVTLNQ1KWuospIRu8cUWGUu
uyKKhcmjrR5dWHOfE82xcumc4hYHHGuFBFhjjfyKIii59IrnNf+1di8fhaNSBkTv
dJNw2loP12y9BsCOFPsD30bQBJg3JXgQjjmAlploCdmFIndy3ZIOGVLoW0751n11
0vJ/sNHCxo5JQeKoNt1Wr1zfYBGOBufFeK1gz1N8RiuT5yMt1I1u5lIernlF1gUV
QtI8SwoMriapLUYDSZeUQ8YB48xzMEMhicxalsyL3e9RzpIgG+6zfPV42G6mlLje
C130bSSirl7wZvbVRG7GWt0EO7Vuk6F6Re4RfKKlthihFJCSieun8IgyAxC+7Hwt
33H4DwtPRJKgLcmgwmgtmJ2x2rFb/USQl3YovOio8er3gLWvJeVdFcYjnxr6TQ9J
RP+ym/ySEA/oF4HNJLzdcA47tUFGxhRoMrOrwDyCfHjx3hEWRmrI6eHCMCzSnDP3
IJ8xUZz28e17mzpeXcENUnUoB9SrnWE6s1h+p0CMQ+V473d28LwWb5e1pj2ykTK2
5mwQ0Dqmt9XTcVfbcFt+nqkLCTxsAFRYrdwO68hBsxLbiEfyGLMkir4ARvvRHv8Y
f1adBOPyGZQ4Kzha06DwV/ZoRRz1Cy49jI9mHEkM0FIwChm+kRx/zzkzRJgi5svm
WsYHwwAzghrhQ/fu0frkSNzkGcnYZu+RqDXWfG6BXG5R76d3VUPTn3xPgtTRclM2
I3yQmnDTqE9YyjbZ99/JiwEEf3Oli7BQCC0+n9jJfI9wTmf8qQpOzY9gSVO2AsT6
V26ZL8C2CBgCZIiI5rsZbev4RO60LQPnh4p5qyjNmsbwknqi/GIaw+HFjPeiwJfV
pMQzxleP4qnyxyF0ZcVeeNd6/bNQE+9P3ixAYJ3itcmb3elFhIdr9HNWrqYqo972
guIqd7nsEdSfLVvrRgJaB7rITf2AYTekk+fN+vPW27LcyIkCBHugS+bJmJ7ejrSC
tS+SDO1Xp0hbSs5o06dcEa101lXy2EraMSZogeZgMqUCTNW6Ti3Z+xzsomy2U8a6
g8J4hEu/4dKgrFKy/ex0dAdLJ/icgVIc55WWVvQEBSXNB0x9fGeXgWFiikzXwCm7
HSlEL6cPwa5/l6lGYMpB7UJ2cMMss08E8Bi6NsTUCT5DwxnEOs23mcxwkQhiZIYt
6oYbD43rE3g2wy4qFGpDEE7n2OBwnf4uB/fFvjfxDAwgMcfJ6xfiwH9G0ZOstbYU
ZEApWjZ2N4gd11+g6A6Zo/JMOKDYzqFer29z3cYVk7NaeKA6g7h24u0aX8LmvjX4
vUTW/mp/vL1miSlr9BdVOkxhyXRrohlFUPOlNAyFSLDkRYvyCZpy3P54MMR0ARVh
pL5OiHj8fHuBYpwL57Laek3TtchlpSbX/Q3KwvlCyNVAltPFGGYuIMETnePMy9O7
jdDK1CapNsMgQ8aGC/pX2uRHMPkOYYuZwr8UiecYyj5sI0PYIfV9h6yYlDPQ6fpm
/CojB7mn0uNjM+66GLXNIHG7OQHGMaKG5zX+0uEoqBQAsNQ3USx8mN9IdiYwjwJC
Fm2Zqy5w5JhY5zkWFv+7vHgYP8rxtIEF6vl1SXHVeOdXxnWJbYsK4fD2bExFO4EL
PLxSadTmS5eLpUbVNND/txHf6um5l3QLbSsvQ+21rJdyPk8DJ6vmpdmmROXp8aOJ
ROfxugYORn5NO6ZrA7mkDXaJz4v7t32TdthV3uluzSFNMaMpmoMLiij7afRhIQOs
BScMSRHta7f2Vd9AKR0aFI9njHyBr/OzSmd66Y7UD+InU36iag04Nd7PeHIV+3LR
R7B14ZLf5K4rxDaciys3aexcqh+GU4T8M18rwlcLBVSsnO8b3Vqv8y0qFm/tUJn2
dl93uDwLafhgc3xYVifI4pWgs4XLgH187H8faQIVhTG6cTdUjBDh587+DDWUpwha
tYQVRNdHbZ+eQKXs79add58RFnlPAH8dzfPeL/zM0TqrjEd0UQsaR72R4tyPOrYF
FAgwhDPAj1Ct4Aq1QIQLy+G++ec/EV8++LvLAb1oOGfEYkMuE61ODhfZupKBBLfJ
ccn3o05uNUJZbGMOHqvBWMc4x79oiWHZV1jYH8lemmsoH0H7/VssXf3GQb69UKsN
+OubT/ZJ1+cKHoqES0OjFZlEo9Gv3Rwr+ApNCBzyuJwoKhAevbqBr8HGMzGW9a23
QY6oWKSG6zmALSlu+IkfOVsV2a1OCJSCQtHGlDZ1ZwrtFA+Jmq1AfY0okfePd14K
ELZIipwmVnE2m/koE4lnmz88xDKXvrnse8P0/ExP2cIOo/Kvvzw52tHk9vnQVd4M
K184rLLvf8M7hjmcOOOQmJK7yHtBDkkeazY2ZOmGXsTbwNV0sSkN0E47yBvrIWzG
jdW/P3c1R04q80yEfsNEpSIILbh4zJoORmJFsHYw84cfZRul/xXVBibOmXqj9nKF
1S6FvLxtVGikM4ivrbgurJoVvzhYO2gKAdhqI4SYOuflikx+zdAM/CPbFmggqXrC
EzTh54fvU7wzznyPQf693f/soZuDxX7TeJQJcRRJFENj93gKU721eLUc/advMlGJ
TyC1yxyR9/s5kZ3hqhEtFFAfQCf60irJEGhcasZnCW8o2wJrk+MshqXMqWLk37kk
wcpKPZOIKyo8BR8qsPgp+SKsPrffz/acQwvCCEuSp/M0vT3wb/SGAK6Xm2LgTyi4
aZXAIftLOb8xV+RgTsc+G06zqjDJOBzmM17KuxCzcoH3CocCGUTcdUEGZZOjcvKa
AQI9Pd1zQAtOhyFg8Cx94ukYAS2n2kL+X3zBoZUrrdU7BfagsoOs5aiDrXVNUDRj
hhZXn8NqyaZiIVtKUEoOSD2g4x4rUYUyXxCy8UCMnOsznoEwp6v6QTcNXoMZKmbS
62w7F+uDs9pPF3bP1F83pyJPbaTIYzdRTxv2T9rAs5GGiswOjuBrU4/8uNM2LHPp
CcZAfBboCwq6XuLT1tgnKQpOEgvZOrqhMo4QQTrq9GmhUAdbgVv0HxF2s/PJamOf
No2ba+VxDekEh71CRaNOR6ebjs6WNBDZeS2vkR/44Jout48RF/g79ngjVZyM9902
fOSdNeluPlG13VWHUzG53Rr2SQlwRx9/hiJb5iDo+EXpDZgMOShw0t1Eb6ZY76f8
ylA9vo7noh0+fhrMjyn+Buc5uMCMiABcBKpAy4VVPx9EEfRcMcTQApwBQvz7qdpU
8tFrUp54gI1ZM6pzdEoIwNOoALrb1iwXgUqqd8rScAqoD/aORun6R1ZXIONJrHB8
YPRyD/yQi+xiyFI9nFvd0GHZEbA696xjgyGEt09udh1fxnT+a+CvELkHjWzG8btm
2dFjRGfSv8fpd2reEHo5te7RsBJ0BUHOg9G4puEXbZTSDeJyYwq0Dy8uPFwqEfP4
H16HXlAY326HA8p+zBzzF9HYqOr8iFME7Mwu6QRvl7807hEn5He5xnoXjhDBTu1n
+FpZmOtGhzKtm3kn7MBVikvjp71+FHP6pQAZXMqoTwvm3eUuM2I8G0rhOsC389/u
OoOx9U5G29lwnq6cYVAe64HPYISIsSCz5pldaayd0ANX5SLF4lonXjPVmKmbAwFx
QInBXbQxFx+j7mOzSNXmgF+oYe/bshEOwf3/6XZAskHwsbRDtbtFNhHRVnaPEQfv
3wFCe8wz1VDqzmsvFOCx3pZRTNVin3NUnaEr6OAkwtysNVeI3fJrSIHcAmCNqBti
vqrdqPublUuYbmFJCyLJA0p1j3cDjsh+usSiESCR9ZJ9RsFSU4jGeB5+tlJLu1iP
0JYgH70SisnQIukV1FUD0NmA4SM0vNbLzeZb9tzhQhm0WHAdRlWUDY7Wgtu5vv1K
AQsmL+LY6h5jXmeX4oiE/0jSHho/1GjhZwbDNqCXmhxeoOEq3yea4oLrmrZazI67
jTi0gm2TEk1wPVosqutaByo/0uI87cdM4B1L0TubqxgYo3Ve64Aokv/+JZFMruW3
VWqfmDh5+lutcniJJeacp6Q8ju3zeiNfnho7vZaf3PsD2WUBEFcGxrDBjZC7fGj0
QtcyCvJsdUfMnAa2fS5vBt7gfDPP2eQYcatX6hZEOqtr0SI3QOX9xvvLJVGLWgVw
nuFeWxnVo7/YKbkuLLlVMrr3DPmh7cH09KshE0LIb0CeZxog+JAoYDH2BP5iKe01
asJHeQbVt7JrE1oLp5AkWSZichn4n350rruCnUnJLGdFwecesAnx7ytZLzky+h28
c4+N0bobwv8g2/xjUYTrqDOtZQ+LeZgMgc07X7Fqnm2vLQdD7zFt8Zft/7s+35xh
BQkje1UjPpG5XLubcuDLe3ZA+sIyVx0wDBfg8E/tnly7gFs0Fn7J6WZGhvlsV+EY
JT3MG/qt5RGQLWGD5nP2Ka1lUzpIAKnQaO8K7zHPLsJvMsNHHXSvgwHZt4cwrJNQ
CnYVRlx6ZJiYu1gvuT7POvE/eYOGkEP5lZ+UxD9D2iSOZjNhm6DKl0wR2simT83Z
73kwavhefDj4gHuboWZGKz6ZaAlDChUGua2rkmo/1nqTfPTqHuUJ3n244RWeq9Sl
domclKF1IqCjtN7I5hqxfxxkQOuSf40x3slTLt2XYZ53uakKwRIEyYuj/Li/f0K0
ywG195XlUBJX4EUE7w7H1LqJ+hAVmBsdgVEzWewV6EfUd2QtroIEcGO/3rmuCFVw
fu6dYljIw8dZ9yQZonzIbdqkycgzsciN4d0VqzzqTrJVE509jp58qrxLAgWexc0h
yOQqlXLLkPhsr9MOHLqbl1HNP4TekaCc9Ipraw9HlRTP1jAQG9vd6oUUzCp4fu4Z
tHXJmmHnQecJLiJXsmF/zlYgFsNrHCwuwlRXAPa77vf5PkP0jf5v0hKyQ3ahOQSA
9wYiWLNTK7fbBNECTbmwSMNUjW75GYg9fEDj8dmRZZVSZAeIqGLz1LEZuUYKLg2H
f9MRJfNlozecrtdYCrtgFmlyn3Y0lovXkTwxfB3nsLhAGEOvxZzKVCgYB+mRPHpk
PCFDV8lI4bCO91zbemA/RkOrzDID4I738iYbu0gvZHU5TC4NN08IpsSPhGU9Z0Ib
j71H5FVIOL/r8vxtug3/QtbWFo5cYnKjz5Hg1JEjA/2q9rkzQTvunS0IXW/0OC39
/hcB/FHqhIZr7P1RTpjfqKKfPjkDHEHXNoxybumpdcvAc0EQN0Ut+O+i8z2mT17E
UtVXGBXiDMdnU32XKO00svyBqLydFY941FU0p60D84qXah2sjvOlwkLKNGjt8YKe
m9J9brWWdOt0oB5T77ObqckWY6dEp/y0Iv8RivriIP7Fy7tBsKhm19y0WWTyOjh5
px8PSvyXYf/ctR6UwmCG1ZNCIFCwL1amSvhyuyI2OfOCLoS1XHuRiqKFNgaJaHCi
k4jFAtwT3O2DIpNJagWtmGkjKdYca7FIHwHd930T+2yXIlG0c5yCufV/kEjXov27
uz3cQeWTD1ePTiedEpADprWTeabJLkczdLgVZDowBuTKgriijc/GuBiLIL0t7Tpo
HhQWsFCEHTNexkG4MfJizsCMSK2/AfhGfDHxfjed0hyUvBEkvcIuwLCwj2RRWhLR
NcskazSnxlOlgPtnlcj62vIutl0SbVLU9K50TgSKDs2UawR6mKUS96xCIPFWRyrN
FX67N/2GrGRBT2vOgzu1OLXh15ynyHkVBKKAPvokvxGMT58p/t74tX42kifvkWBV
CzWEzaD7k8tR3n9yzr9Ef1HyGiG5tM9MoJd2A7pXYMiRQzOx7G60kSKkELTHRAt4
Ztww69YHilMCggGjwe6sAX4FclZtHq2tjzn9Kmx97ORBSMmpw5a69rfzCRc4tx8c
sCIJ20iVp8gXT9ppIczkSPui46v8YWiykhblIqubDYPQXtv8dnnaCiGq+UtGv7pE
HZL26PsBP7s40HkjDS1VqTjoza+bP0oqE6UER0+qW5xS4m27Pkt7nzZKpOuJUtr4
39Y3qF6SGljB6qYqfsTEQQGU1AwUOC1YGb3ZDilOwgf79kuQ5H1ky1msYfhbDxqq
v/FuZQq2rloGUZ+J4H+iDGLthbDu3QuTl0fU6fK3wk99yU1xeZ1YNVSz9ojk55OH
+UpFgqz9AWQ6riNLhRXS112j3OBppXqo8/y+kKmij44MuES/YplkgcZEO657HSkd
w8fCsSFotHVJeSgUnaRAdo1JyBhGDQZ1z2gOZTa1aGhukBaAuTYQZso6eJlNrq0h
KVyezYczegIKx1GHsxGrIUEfJ+xpH5iL1QagOkmntlE3tpGSMP37cB41rGXE6o4M
xL2pddafiSW1fsUQEletTFJSi9uSxjEbalsm6nh0dnUoyGNG1OlQ/WDXHgkHZihP
LFMGbHpWMhHHCn4JIuT/OsVjXSPiYgaKFzeXU/0rlvdGYlrMKCpWZ0n98a/w53Hj
rFAUbPS28mvkAd9sL9munAly9oQajuf6xo+EaQqZCCZg8skbr0XTWhESqeu8tGqx
nfMSO9neDjn+b4fzmCvcpWBZaUq2D8+gUt2/UBq8Lkuc0DlLjhCnLXt0Y3KmulBg
dSY1AVBuxN4ESw/eNFaJ5Oty6f6w8lVgkoF1gMi+b+xZO8hS9O4DNQl8Q/u6SRKG
SdePxylTFk7sBIL8fzsxXG6c6Y7M7UMUWAPnrT/DXVrI8mePzLZgU0rn5F1yCdtF
3H5ELBsEsPMzHkZKiw5p8vKHA7ZbvaY96kL6YajKQ6IQIO+zxGKt0Xat6G2en+Vb
t6T9FuulMcHSZRe5W/xRzzX/UOrYPTq3K6Beo22kTuSKUwFrw2b2ZLaSMi8LUBYI
VobRMNRyCwRz6xYXkaseA6VvNXYGRI2S+Tlvd3pj1obizVWKNWDAAW1kZr2pp4xs
//W5AQxFe8BFQOHMvreo+woD7+m5fQZp0e+yXCYDZPEDzbvP/eyLO0lgebyvX9kH
58BdyCmSuKfO1rXwbQS7xO+J8VMxF+NzsBk3LPc32U00RQXAHrUII+29yDRxc33T
72MrJwV+nJXH2SmzDw8iCpbeK2y1SjwM3XxgAcC1JBOncqYuLVXzNEbrfyAD+g2+
RgiGgjlMXRZdS2uRnnIJlYJl5sQyA7Gp9Hl+rs51G3m5o3JEAuNtZPZd55Ixf3Mf
eurjP/xbBXHeCqYfgAAvz9LqNu6YH7Nw8/et/hH84og5sFc9u4qe3qMMtLdVxcgD
bAR+qmaMW2O2URBJeWNexnXnZZpnwI5O1/T/YiXzeMipPFAza6j4kc5TwcE0oWjA
j8i2WZ6pzkHazXvZ4ERhZC9GIkcGjlRtNyQ7+6SDSeJfMsIz63Pi/oo8TZktZwRK
kqt2tpqZ3Yo5nmZ3gZ86FbpKvKIlT3XC784DfKBQ3XFTdQZdxj+R5qyh/vSwlitP
LqEDAcGu2UjMAQT8yakVy/HoYhW/YSyQD1nZQR86egW6jOyJd/d368fTomMLa4Jb
JLLIpncBHayTK56JTtvIG+DiE8FLfH4C04z04qui/BPzl0nOvgBhHsOosyhmrS0v
UYSSWEtK/De8Jxdjq1NiIW2wHCC1yM62myIl6umBaXxD5Vpm4m/Ii/n7w57/mbIb
QBkm6w3WnAQAWSB3QuVdowpe9GdaN0SokyABzMdQrpdNm395t0B1RBYJIUGTUkfp
q/RReHROP4rL7b+UHMSqMZ1vs9Deuxl3+re8f/hA33rgCi97pa2ThKOWwsOn80VX
kuF8uaCGyV+NG8v2Q4ggFlNWBPLx83bCh0yMHzS0Jb1R9Z4zvjpMdQ6E8hYbpen+
JzcfiCGIw4IN4TrUbEwXvrBXj0fE7P6o577MYClWXqdFNWu3eEmx04uFXH/iKF/O
JfaUJyQ8gfxunDKiuVnMPZjX2yIJtwbHD/MG54laHJCORK4rG9PeIaZGf7q+oOaG
q/JD5yIEzEwErGeeRVfwcEh/ot/fJyqiGdIqfJQEdNLv0/8pYMrvzxGQ+WQObm3H
B8iG4Byyl6lSZMVD3loNT8vfc3OaP3sfwtJBb6lM0fE9slr7mFCmDjCLbbBXOauA
FpXJmy7B5t8b3sKD8sLY6/C6nrdL9yBESizeDkKEsL11A8fXeephMlQE42nhSOr8
iYoW8gK/X/IW0Rq3cxH7fowjZahEzPSdahct9i6Z0BJnXIaVTdipVRLytONTjBxf
6bcX7ywWLkof3WaTnVmDOEmwgyHQQiXx9gSQCl5l9mbUvk3AoGBNYw0W19z0EbGi
Vp6EMHdT20/2GQE0U9eECkSDqROJC4NVfSHPwp425IoyJSLsJD9NFXCLmmyi0eCY
rMSeQaLoLyHj+qU8nL54HvdeVSU2Rxlp3pZaeWhAag7PlYQnHi1C56Fqs/Mjj46b
3SgVytkEUSzOVkFNDrjcw+IbPOHNWzDM0xtom7OUrezZain0UfCgzjC2JEa6ui4A
0CjtEky5yruPJt5GfmcPEIdnWjorGq4dGx0pU2JhB9OSdxn8/2HKH87/Mfj57pYi
+8lfvE+5tCP56JpjBjDY7wAylSgrkRptcEc+vbxX4l6XKqE5B8fPrzPR+gkfKHw5
SjTfTFaPtR6zmrLkv+nLKhipS/2gK4vZC2fukYE1TKrONUZZ3xz7AWf0i84TYyIk
WrQrV2j7fYxlLJ7JDZMcEyq40kG/ELx4hR13aI4NXfzRW69FB580NbFIwn38FqdS
OpwgUSEqnFC2GgxToB24VrslY11lrb78AlXAE4bFxEaiZhHpZshAfero2GW0Osc+
Yqkgc13Wjak/aBZZEPE9h05MXLwSIxJyIqeeirfUMCxVrmx+RmX24hIAY27TVkJn
/RR2Vz2P8ETp5t9EPhbRwrOdCE7yqhqvEwaaX/+2K9GO0tu023uBFK/6Dp9951TM
4GvJm1+6GG868tTFtcwOf3LE7UIW0L+tPGTj65hH1+uAqFuTlCe51T9n6hphmmz9
SrrJbV8+IH3wiE9d4xplvNfCIF4q6r7XyXbWOKT/3iILXGwwFhveebSUIOhUcJ8S
FVdcB53Q7oYewYNPv8mHsZs+c7FHiJHBdbpt+mIEbX+AkWfMaml6mynEuxJtt3bW
Gd6DXv1kGcLrrtsKwe6WHunY5VDu6LVtTKKka6HaQW+n2BVBuMLQunVetXFpOIUG
WkvB63TDiyVGVVziht3j9CTy3U8DwDlQcjWr/iupTo6FwOzqNaz/71l/6Msqm6mO
+InVMmBPwsXrokstpTFRyUzM3m5U4uZ30SN87b2F7XzfckdgiX/tr3ESIfZtluTA
l+tabqp+wWutKYKEBL7eaMhrPrZgKTR1siPLC0bnipfdi6M+pVzB/jYGNSV4MOQ6
gh+eTxfgysP5QYoOIzyaFMqmc3mbiKQ9sfdjucbsshkD86FcDk6Q3vqRzSJUpPdb
EpuCIkPrJvMxHG42PADgPmE8T0fFY2USE+Sx7AEiKyhBiiRqsTsHhB4KdT75qerk
NUUzpvfwmrzU6uRkLuSX2P8K/yquYp8GG0qLVNePGzx9QpyUssj6aRDFb9QgSXXy
t3JlgkOKVkZ2g7QFD90Ww/7KM884IEBml0Wt1HyCnlFZ+gPivb3tinBN2fxXy6TD
R+3jaOrHsHdVHyt5sJeyV/LzHLeVs+krryufRRMBpAudIPsjPTFMgzkHQVupB0ve
G74viJ5366dIbFPNbzSFvN63k3nMet30hnwvbQf/x6Igw0rz+QGZUa4e6xf6oZzD
xXSasazSbJk1avS0kFzI5QNM5tqiY3uZ0TjnHdABowwGNx5aHYsWvQN/kW832v9N
47DDhaTwHY8G3Bh090W3d4iwY6So2CDBkOs8z4b5hGphL6N9OVTrcrrkaW37W3TQ
7/I00D3sMz0BwsAWMNzTvwPP/FsDfsAf+5mJ5qbbYrExooF1A4o22rfZMmPbMf6A
1EWUUwBmHvqykakqDh/jDQ4sGmbEUCtxQRgcQjMre/J5Wp8ylOuB6tlXybsdekvi
89RHQfkDFm7jEBpWNNp7zPaiiCYsg/Fu5ZU3GeK51R8uB7TKZutrCjWZ+Nqp7N7B
XleW1y0h7dP0nI9JwmeRscrvIcRja5qetF74iVauL+OtT8e0+isayoGKPjOEAVC9
u8pzbJGhiqGXukQqaTnkyeqV/Bfv8IIijsfQvhXrYmLKXmWPTHg4g7rlJUiuYWVP
AcSfE/ufMeGml+2MIrnrTCNFPQ7zRrhYsAu1Ny76ZHfZ3rYo+NR9Q6p2nAfWvUio
M39fzkvLBNMkIg+1jVSVJfceRy1BcAml+UXFlU4zW9F3HkdC+kIhekkTtnbjhiUR
1G5elz5bfcdD7afVD3RLGYQDUl17RgYfRkUlxVDM5CFhRR9kYLNZ5CkjFLgSJW/u
kHkSTcE5B7hUROWAZFoGmms5OTb9sSAWWoevFQ63Qy6xjtZJ5tFuEouidZyJ6VfJ
cZhZJKHO9MRn2wytLSzvVzjsUvDm8oj4A90JsNd/0XNZtz9A2mV/2/KM+cIZRBNj
vm2aEQiAZ0OMHTHwgQ5uKiADOohAwig0xL0ceHznF/6RkVlQS5QzLR9jvM3E+Abf
l15xv+K8vc/cJD0VwW6EkHgVgt/WG0l54+KuMBjLgKpqkd6dtNb8jDWrvb8IxT5w
zg+/BylMYx5n0upEpnhDAf5x+V8Fz3y2I0YEYswbsuAycgyQiHz8x3qRozAagRds
2ZMt/zt3alxGQsKTDpsKRDZgt0H15sW+L0oCV58UjhCSxAZIt5ZBVyDdIqVa1gAa
ugO5KN10+hxX80BmvHZ6VSWKj0UvJWFHUpMATli/ThzkZpZPL0GnxxwGalBDT+S1
ozsyTDGKsybz+9tiNNZPIvI2/XQaO0ZfOGAS1esoA1Ag3zul4iwk2vSlxZHIEqUN
f17jBmHU1b5qhfKyDPFOZZNzmI/wFEKTr5Ty0lF2CuYw5IbTAtVsANDXoGbwlwBu
yFZK8p+/AGq9Lt66VOTXWX9JYVu9RQDQSd4ZTA6a1jhCQRdeuKNihjeRPgXJ3NgE
QL2AFIxc8o/sxLOmCN7WLZzrRzCQ7du4knUW4ouzSw9SOsAwTo7JKjUNfjpMtIIw
hQYx9RB66ZbsAxsqSIK86RMVAsIdhZ3o5AZmWBaoE4T4hORS/XUrgds4g5x/MhCi
GsAaRZ34nGbUDbTeGDDuPAmzoCCGY1L9NiyT5Z+jI4ga6lG6xpH+QXaK1dMEqKg1
J8jXUCllP9gUO+wXY6V02teMapUSh0qQFp55JCRkgb1YyXm9lrEBH2SbYU+daM1N
u0qVpYvQP6kpJjS0AQnjTh73DbnkQqdxaQcQiiTlBWtVpqpkgOgQejYDyYfqMYaK
3jxBA8gnpT6tM/tM7w/L5cHEu3d0UN8eFkykDU4Dr6d5QBw4eXtNkZWzPepJ2l8Z
tLqFk6WPRcH8EYe0bd4LKvx+jedI/NU1PPaMuxzWd/AbL9WOVpQF5OU1NH6lI0iP
nZPHke3HrtDG0SoOYKMLXRJbVxWRz8u198iajnuhB4IfnLFrT1FplJUSQu+AExtO
e5V7vWWxzvoGLtrjSFwmnoxqDurS46GtAgO8grQsFpPJVI5gM/qst053U3FPX6UM
160M9XIdil7qP6MG96LUMYnxet51qPf5Aje1whlpZ510UVzR9igKdz82vKgicpmI
aX2C7UzGVh7Eruow7u5xIxMq0DdrmdcFeBqYrrmFfSBnBUQ85+IqO0KdhrB982pl
29h0Mib/qX1zWk0Gnu6aGhdcY3mQu0nJUCLVBjxgDwLcbRX+p91Y2dUB7X1ilnFT
3sz9CgMEsHzY7ZlhE/qDh8kyKRKYqMRH9v0kzEgki3zmU9kSFlAP2RF3uylBA7dp
tiJSHEXIFu+JEuSxrgMQiJ6Hshyu9yJad4T5bYio5GTo5YH3625s7SOZF8qKPC1V
tFolkvDphEzP8XddZ8ogVtaHFSXPX5ObDRnegUFGYY+xVPmW+WZU6yOhWXA8F29V
ANHWqekhRQ5qvIJGBn+fBf28qTz5VxdhzsCoRSolXLIC7iUgCo9p9XlfMSPenfiK
LRLGlc/9xBiBg+B4YOmh+j3smm5IATLRW+NhypN7rEaRUCu52dl5YntqbD7PGXF5
tLD0e6NLiVBRfilSXKLx1qs07k1S2TBMckLAz2e0PeDuSi9QhyUqcTtkgtSrWnw2
0yGWXFe0xfvOD9wmK7A3nSDVMwmb0bDHDTy140K7f3zKSAasSJpJfyKYIizt8Nt9
xK/KWXR+emV0WPsAhMsojLGW7678p2I7DNqhT7gjmKzB9PL1HS+fiBew/R2+VPuq
QWMpuNsVitq6TgiHR2S0w+fauET2ZKSsFFBQ8Squ8SzUlcLPTz/lHZtivBNwmMu8
8lDZYKQx/qkipqCJWygx1utora9ht8+6GbrfY3uhiuTRMoh8LkaRLEeb2l3ehhKH
MdICe6UMjKsgAMLOf1xkBofkB3GQHgh6uZTAp6KLo+azofyYygpV9wCd6DhNbuP1
jAWMpsWLTOnr6YG0NxCfHcHkUvCxBZlQb3cW6YSnQzKf1QDEc5HFwSGNzA4cOmDs
Icis/SSgd1Fe8ibV92jvRtSDey0ZSNfdffz9SOmJ/wHxhPbD/6+BzUS9LJ4hr6ij
DlKSfDCugRNf+EdGExYhY5pVlTLq0j3/vpQHJQjIhxlqRFyI31f7ezOR0fSvWG8L
SEPXHQBGeMfVMU5HQ9oBGGjpzlHqQvmPjOTnBxcvZV9Je6g336rAIintNahf6w9X
nxGoA1qOaMkMc3Iyiu0ZCNtj3ZCcuNtOkDbOBvhGpteNk/A+fPDOpU/VPoUBE07R
uSfj8FMdfKHdty5hXAxWwBTfwQVy0EHE+jxy8aoUMBsQhLobhUQkfhSEv3cPV9jH
uDY9geK7hCz8mS3jbvSr6Xmin+rqfr5QYIEAOT2AHpM8hx551NAAcEx/VF8BAD0g
cnWpLPTQR9RJscnMImQ8rsOAhLVKtrrjyw1PfT+3EOEK8PUh6kCvYAjlRutGH/QN
LfS7JQ9x1X6cANCNzeYVpY3H1Zc6jaxIFfh0SkwNjJMYNnjaGxUKOROHf6rPtq0v
eBH9cMT7efkfHPjLAn0WlwaO3gHbQIO7R4iLVVRz5bI7xikvh3Ck2wT4QBLflehG
nLP4bIO+gby4DNBGRwsipn4xDLXfEQn+wPglyYTmqhTWIICRFZYUxSz3MLWiltop
qzBik+8GDenoA/PiSE7AQqPpWIqeRteCsAKSdfQUbhuRRc9uruyBBun0WOsOfe6r
EH8ZUVNzMjBnsla8CqGoMYaYFMeMsampwxqzRKc1W3m1i6pGeabLvjquFNDXYqNY
143TIUmQbhftmB5peuZrqnOA7BIIgYfxxsk8TBajvZcOSEzBUVijpJqzqPryigMq
35+5Hwcydt7LQsHnwoIG8BOWe4JHMcxiQihCDSf9E72EhXAhgy2xMjo5NL2BvZqO
KhWpwdqDqbqRqShjNl3Cd+5nc1oqOXe/2aXah0exdbv7V0tUfCQ+TWRNNIxNVaqQ
Rjl5ZALHO0GckdlWqLKdDV1eO57Ydz7RnpZHDo6DgivId39SmCwX4qJmUYVH3uHM
OjWZrG9ede/TKpM4eEay/qwzAq/pt/SZmRuM3MTcQWIRHQ1YsceqbJkrrDqbVNzh
Re4oYmRqD5QzwDYsqvIkxywgZWTv8yWwTti2Ebel3fk4HVjeFtcJ+Kur35AHUZhM
7SNE0LNL/YYasBMI0aEPtGqxAfakVc+zTRMtZl8xfRmtDP6kBIk/VjbGoP85I9Lx
yt89zdNEmRhElJkxXvVaH8LBG9AHfpzAhsvGpYgESItihtBzg1sC6fwnwXSgzNRS
fItfLbazFFprCxxvtg5jWUQ7QL+ZyylBobpvGzaGzHqfSF1yG755IBBQEnXoF+6U
RHkN7r9d9PgYIKdfsiPkzFkcL/BEx17Q4Q6giZY509zdRroqaEkFAIGBsBa+2/MH
2WVl90OMfgIO/8/wxciJlETr+I+ZZ50n5K35q+5Kl3gZt+GAbw/kibIbJl/NqD6M
CsSUHNo6A6AE2GAM3XvfFGgOfqFRpX+r3G2Kl19nB5cwBg/g4HI0GdbYxMkNQD/J
in+4xAVeQZSIkTIVuwZscqbuLwogQDBuZMesQLC3EmKWYYQzlEdQ+B/42FKHaFXm
0jfGUhhU02a+1Moi/CtPn8VcINjlJIOSg2GqQL5ZqyXNjjRFW7AbWjBVoMSWHiSw
boSfiT4TJZVSQmXhkrKPhjzbWRD21L32Aa1boqif1WiJanQTGYf2rfJSqq7jH5MT
mJ6vEaHZVqSAkm31/uk9m4zrWsIVemgpoYdP32TGu/h+j1j57jRJKa5BRt8KsZnz
ZE2FazxggTXjOddaLgpXAvgpuWsTRtHs1wdCGQulMlCulo1GLD3L38gg7sr+riIt
X0m2jR7jxQvc3LDFLwv10CvjgpkX4Xc9v09y7LABRJEgV9v0N+q+fGr0eptFcqUW
Iidz1zejNybz+6Gu0PtUQfvn1043BSdssEC2NQazckIKCZgRGM0krkf0F2Yf/YDd
pBC6zzcMULm3dTBkiIoXD8Yc3cTMS61Ez1Q6XrfgHlZEMgHr58nNkTFF+1pKcVbJ
S1c61lWfLhrobTMF7cNi0U6NkM78+K1lWwWzxJfA0zwtGXWBwmDqlut8V9bABZRE
kyeh/s7lxI840UPiBYttHrf/tf5ltY+l2Tp/kiSZBYjpBdzk7X5O4W6mM9FsKrDu
7Gz/BnZ9z+AeOKhj7jQfkDPTmMM3HL7uvoBIh+JUZSI1bcB2s6/vg/VNZ6VxOOuD
3F0Quiczn4ykafQ5NN0703dvW75QBe1jy8T9qxSJnEIGnhExibJVWkxWpOrbar2t
stG2HoBxVZBO63knDessk/eWZZsrFMv+XxTGz6shWgGtL1lg78VE+SuXXLemdPF+
VS78I0WneQX8R5uZma0FU49RIiRUav7YNIxOixdzUVMhhIaV4mH5sGwHUxo/znpo
kFnhwWjoGeu3cV3DIY033jC7oMhIAjfx9Aax09mz7Czzt8NLHp1wI6TIL/VsPRr0
pjH4vclXNEmtAjV5EpUAN4RT37+L96vsBT7+r6jd2V1CIuU6QWzxdlXxkV8Bw31w
qtosnAXo/0nPZW9bUfIFU0EWlpssggkNwBqbVzvlsRaCJibdoSUQFTkUXwlJgb6p
k+WbDJisKt3KJwRdcimhjOf/gS+qUIV1Z1YlTOwcI120VpriQw0xD0ouqNH5ho7m
d0mVV34iZ5Zq2r1SVQkMnT2cObkRwkuoMx8a8/pSnfFzY40FExBkkvZYk7dSG03S
bfwdUmXTqoxV1xdZYcGs6LGDl/22F5MiA9tZp3GjoFoqhDctXb2O+uJzBc/Pj8F/
Xct9Ag2zuUyiJ2wlW9RGqEYw9Ag7ppwwz3VCfvWyJUhmey5odwMLdlUBK20TkZIg
Hu/0+wq68FaCOU1uck9W2YqAewpHoJi+SSYtpFmVYPbOou1Egy7ytqxFlAtaT2fR
47mxCxJDW59sy8HZqGco50t5t050yrrd1HIY9FKi53rdQWgcre1d+Q0HyDi8cTFG
TbNo571s+Ge+EUpJVHuBnJjVMv0PiOz3vBOdZldTTJU400Voec6FwdxSLN0vJLtR
EphKmFeV3Nz9qAcC+9BTQqM6LTp4f3aDrrjpUhNthsX64Mbu6iDspxhivU5EoW0N
O2kqv+FAFd3CyAei5voUsvBeMyDES9E01ID9MXdKz9ovNCvELTE1S7pr/v5Q8kFX
Ao/l1JH7/9HbIutpLq6A7tXKLKHo8L51X5aGbadvKPqq5t7VsHbeXsrdkpNenhrP
ydbYt7CB1i4q5dZR45u+MBdhwsv2E443LfBWmeHqJ2Bo80TYaCxkFpkuJNOq9/c/
vOWyv9PIRQK16qEuxFv5u78dVvoO8tBkuiwq5SZxUm+HFx6yDzRqNRHzCU8QUIpR
pzEhxS2hlhTn/f50BgMVm8UeadvN8NFCvevv4wuEao65NnCQMHuW2ZycYCnjiLt6
2X0LCNqfQnSawUeePoqCCF8Tm/osown3GekMbuZgkykKXYzfNEUnMFtA/oRtRan2
TnmjwVCVcj5M+Puaqa+onhROvP6VE7CntfA1MJ9Cl+CKxRTuLeV+J3+KXQ0uGp05
iHkzpEgVMaWbiJsrrl7BFHMWTzqoEgVvbKjWZHdb8AFEQQ4kvqBF59ar7UdjOpip
yYDQjZ1ZO5uHEpgBvukX4IlkcUKnNrd2JVBxSAQSx1t/uxAaJw4hveVxz8Q4vrPH
7vbKVklPZ4JWAlAtj3Bidi4S6x5Nk10/NMKWl1b3wtHw0CIbrfdlYhHfFm2uktaW
bCCt0Jf4uYWWiXimUHB8S602GhlBKcm4Ul64gFXXpbL/AtzNZGreqUkiHMLLPeA/
COa2+X1BXHsAWU2PN6zP7EUvtPegywOnewp+F886VQ1A29flhRbBhEHfcpGZsHx5
UdYE8F9Yuf5FNxvAeCB9+8kuBQXYDVMDLF4qM3QpW39TAhZbYM3p+OlFmfkKny9A
MQjLOpi41T2MceYenCjy+QDu7dpq9TxCqhmJ1CqU5PBPJ5+L77nu4/AO+wvYCjIb
cDYxTYR5cutw+sdv8nhg13H8+gsf+uRbSOPOMZh7Mk47178QJYzXZYARwr8DfVpp
rRUAdvsFV/CYPlIqdp0STITVgjPJ5Aisw7281EGzvnZhBkdgcRrN1jZYm8xjik8I
La5ZET6gcgvgyI+tgb18o+e2Yxb1Joteebwdbf39YBpVJaz5Qf1ue1d1CdPChxoX
PF0sBisY8ywX9VJtCgKCj+MBjJX3zzoAUUfvZ3uxUp2ZLVFFV8IXllYOVMemJWCF
HOdSjUpCkIVmAgl4QDIV3S1F0HU7eRvIsQ7vX/ulh7kShdJv+QSIuZc2t+IpgnuX
uzIwusknlDW4Gr/mcf2bOVkFu40Cr6GVT/9naj1zWdFTMnWw7hectAXtnRGOzZ4v
oU4k1PdDuXZfjFsH7ZUlqAvKFQj3+xhG30dEULOw8NhC7Mg8etKMJIbNxtwW9nhg
t4yWzB+pEE/PcOi4xOyVbmfBJViXoSk7l0+kjb1LYOmxmbsTvmHQJkmfZ/dW8el2
/fVNnom0Hiz+i4FM94yEC94+hh4/4xA1PVNkkNzC3i4bL2+vEnhbOtQ8NaaSoT60
M7Kynszx6ApJlH3rSDDK2xbsOb4yXr3i6KaNJJZZc5UCCskDJ5dh5DKw9VCkbogA
3PD+XftBlGYpovlHLWWpLFU+H+jJlS416sUxGxviLFcyuujifUMYuimRvzYs+hDf
3S+GDJ8BBnxdKZuKJYrHfMft0JwkVupbeib1SFPlJmKNcPT5Yz1f3eWiDVl5Y/3I
9vxltPfnVARyBz5vzshaX2xmARBAC1UuFetGMtQ21COHUhfciScTJSrgGSbcHha1
fAX/SFkbbuFs9uu/hagsAgXv7K1rYs0uxh1nQUHUTtpBTusMe1RAgat4uYInq+6Q
HGE4Txhb1bnBKsxI9CP8K9O5qfrg9ZcYgdBCBfGphUCvpU+dJgz1Gkigcx8jJdyT
a6E4qkjzHEHbIZTkZ0QguqsmgswY43mkcD7RDYgx+7Swu+Ccm8SMkDMrTyjuvHwY
M1aTb+vcwOtCmWVQODxho2ql+7TlCF5iu51Jiy+zW93oiPAc50mY2slklR3wzUVg
YtVk+jU0Y5kaJczm3ZXlVlTifQIvW/b6d7uYSIKizL0nNuKVyZ0zpxIwLk14yoNJ
d6BDvbMRzOhD1aP07aJu/aZdLCdsNDmiNvvirw68hJtaGKForb+miMPtnrmytCzL
z0XpeyTHOCUmPQTSELqoYWHv3ccXnCsN1Lmgh8jY/lXPK0iHPXQwnuSpOO4PZhom
1OgELIn1KrLg4GAvL0CNIyKm8gQFJ4LK62nPV140roVMRwkCHIpGSalyTaznc3ln
El8ySTvaLiBpg02XN1PVCVnWdnR6SKio9ZX/XMHL6Vhv7ZsRi/32X/fwdvmITT4U
9j/sE/VdKBfDL7fqvsUCnfmdbymTBzmXBoeA2qox7XszGKo9auwYnVMHCMdytN8V
NdwMVbvvH0QEJJ9yY4u+rv6wm81Lb8KvwWyIjo8edqNwXQ/BwjKhh2ilyjlSNDvX
E6gDr8CWhnULEV/UUt8fOGetcCiP61uE/HnrV0gC6wH4tew5S0kUaV30qRGGdTJ4
6ziue5hvC4wyDDCgymysljV9sWGvU9Lj1RmobplqxQCkSsqIEd/+fo5d0Cnc5JND
A3mUUuEIakme/Gwvelfq4xaEg+zD7yth6lHPsRObFWlEKWfY2s6b7pgdSlZTvFt8
Q3FcnPTzUlZcYZISYdN+F1anurIrIq8j1uY8cAIOzAP8NYqUg1NnvmHRcNQaRLex
6yzaodQUbDelf0+2z7B05XzovU5rU+ClBXLWiUtoqiBfnStzZZZVTlA6l+yssJUv
ZAcdwdh6y+IfpyCju4MSc1I7/V++bEBjfxHcUnPoAe/wzPP3djbSw+30XVVOj1qy
pW2L45UswFEH6jfne2sbGWkUiPf3WsAeRBZhHlYoHc7j/iUCShcoj62/olVwU3nP
jfL59EBXw1dDhOloC0NBZjh2S0iwlBIghijD0Hdi/tSdeJ1SH/DIhgp6/xf5DEM/
rqfcwf8LdMsXrZXyNPJ4KZ5nFOQMfPNMn85Q5dSwPh+3IXUCciZVU/DBYFBmpL/4
T2AUu/ftleELahMiY3xerbwIBiYkQp1d4YAGPK/ld/5VqrQG3fWdMAGn3hh9DgaJ
0G/OqUJydJKxlVsyxT8fCxAKOUgzDHOpnOfPzMopEgBoybmiDerBpj9jAWN4xL0+
u246htsvsn+RDaClhT3vKRa3o0vUoiPdA5aBLMjQEygtowqHPHNEO1etuZ4+eLhA
MqlpuFpw3WCB3+cUb8YMm/+pS2dFhg9L46xKfmyg2GzMiNo89oB/Q9Wz6f9b1Uor
B9+DIGQGHeLsj4XrIWxWej2gSem6PEEcp7dX4zsIoIzssMrTwka0aZCfGqHhT9+v
9EgifJv1TrBMcuj0RgJCjJyMGeAxHZH6TTr1tB5YjTaNtJdP+zc1JUsJI5mZwSqG
OavDKdC8kxSJD9KuXJlGPnTghn8NFDTp5MF5k0I9qeemcXFIgBR2TB9zhfsGcex2
i8N5royI8lOUkQmm5N+lX4auXOOj4OU4vyGqaKjq3BpXDH3g3/RtgI9V4bgF7bDQ
CYmzRTwBUz/p/miEbQG+A7oOdF3GfXYWU1Mb5hxfEKGimIDkXClij905WJ7xyVsI
iX9uvHPu5MtfmC8fa5WBhT+C8zUP8bydS1Zwy1N9C3ILmXYTM3gZG1Btbk94retw
oz5UyopUJRn4vdQhWZV41xjs/P9xDPQQrHuAdEFOnYfEVYQ6lBUHVaAuDPcwAVd8
D8NnySqLSQX1+sd0NV4grQOyzzoDIhJ3fZ70+ffFwxWFYpPo8thEPARVuV4Z/J8D
+au5+s3tEYT835MqmEQndvvDtjiu4tEDAxixU5KAnQnCBBWesDQlW1CCzlJ4zf8i
8+kZ13GqzQ4hjzlbuUjzddP+pVYxM3nmMrn+1Dg3ZLDGZANRaE8EEGVqpjPNYSY9
ED68IictpU31Bb1/TZlzrPsGnSrp6gCmcmBYDLQNm+2XwGyMxp203RlaJZLpL7Kr
Uq8J9CP2hAkD+OxM8vcFqkolRR9+pDVQ6AG2G08Q3fIQL6X3ztUHTe1XGT4af0pb
jpl7Y3YvyVx5TUrmgmdP0aws8dg7IjS59dz+6K9qpG8MzIAsM9E6VAUWj3e+76xk
yUAxFGkAKTR9WcfunqDavBVMTN9CqSxwyTgSFH0+DiLfnaDxVP7Kvi16uO9ssXBe
U20nh1BvoG3WqWKnicgZ/3ZhMC4OFXqk7COAJhDqwpUMKFa65OWneGWXHTjX5GYa
zkK3dkFZlgS+Pm2coXxDg7O2f+zbt5ai9dVn2ZXBmWnh2HVZr9oSNe5W0fr1FPiv
LM74ExMqcDOCqnkP1TotuB96pm++oBqP44y6tYjTF+BKr8DoZsWmzSgrGMRSdZUr
6yxk0VfDv8HVL1UPB+vq8fm2uwAxF8w5d7BkOPcJ8n8r62OXNIGVlCKegBLICEKK
U3ui9VB9Lihq9F2lzlYlCWpHweXtz+TnB16Q+F0Sz27f6+pJ/hgySTwVLbTNupUr
q37CHANV/zdnqzBdZpXR36XmwsYz09LDJ9AuTGKwr8h6CT8sR4NzMSUG9Op92LLL
l3SniFHz57qvD119pSyI7+c5kOqdT5dLq7wBFhWUHCYdcVGcsnXd55wnrrFrILXK
Wz9G/Yhm43BevaNT5S/r/mDPRrJEfquVjzOdE8F5ynd5fsc0Pz6rIf88pemyVMNe
57FUdkJ131VOyG/8RuCgeK64kacphKldztmCjN2JOo98Ec3iU+3xM8x4Dvw/bSAp
+oyj1YhT/huhWj5lLbj+X4PayaWMHsuN5tNQvaU4hOz/ZwsYW+3uER3rJIVWXk8o
e8UVtcP6jXOR1BvcYKWIgARlxU9YdIHWN9EuQ+9+MrBR5rS+Be+HX+mwcaUCHlDa
vObrktHeCivLp4uCIGGrk+HYAQbgGJV+DZ52THbLaXH0YDnLGdi37DzMrD2sp0JQ
+WIgtoPncdejvQ9eyRy+UJQ55UT+2TyTNp0vQomymUOOBTosKQ8eSJ9+0PzjF9E4
qaaK2L8GbJQv7NDS9j/mKRvAu1zhPDp9ygTUV1ia1Zp2IwLK8H/rN6oOSqw7ySG1
NECV8mBGHV5R8slr1EbnQUuNQoONynhrHihVBZCq/2FqYjg7zasn8IAU/iA/CyVX
VGNg+si6GdAy9W4SdXo5mt9Tp3pzlViu+jwDarGzzWI8c60ICPo94psHwyq42VZi
iCXBODy9JhoN+ww0X1EzZgMVvBu/LtKhJxiS7fC+Ml/he0AjfNyNf4H3DycgEt8G
b+nWqPGr5IO/niAuy9pf3mQt5eM84NSGWXUxOZ8N8Epk+W/8hYIWrEcagNXUsP6h
WUATbkmirbAZBTV+LjIfj+jxm+o1pkzrbaOiLg2cO0kE0P62squZIvz0BkPBoV6i
A6/6cBTb8khegtaNNJwrnewmldHvYgabrA426aNvGQnmxCyHcUo9oW7ep4CinPdG
Ud6SA0Nhy0WcHy5+4eNeIuE1JxH9NVbg+eAM7EPwAhfG6iaW+qYhqaffYemuKuF0
ojjXps6WqE2/aCCbuq828pm2/19puQ8hiQgK3XOLaOCoGncdZou8BGz8jpaaRQiA
T+L/eCcbqf2TRryPGZ1jqOFLnra2ktpVDDqRLV6NU09I4BTWXPn6ElR/tj7AqxrK
fTcWP5z4Ln8+IXl9Gp81Sdg+TnsmKoSk3UNFqiJ92ylHHn2vcetl1VVxa4b8Z4La
mLp0wratNMqTkBAmQBd0r8oaACrY7vpv2jDYDaEDdFVlA0UwqG/RpFQtk2vgAWus
51KNHC7DGDyHDPT9cpoI6yBrimPg1g7pX5CJ6sgmPXUAASr4GfddEjvzEFaR5jCo
NNHd2w02MoU4q6NCgztCUMa24qjgd3D+3mUqOT0xBttZLqkDkbeCTiFdnBR84Vbd
zQlbLX6TkV6/MAJz6lbQHIuzAdWn6tq0nIAf5x4wF4hzU+O+8QhPc70iY9/rCE0j
ppGilDu3CBKqHbFHyoWNmJFIThHlJHOfp8ncGZ5EG4rl42rFJai5CBt5LH+nI0bT
7hux/koLUCj9gWqVKtb8aR7MMR9Qut+W1SMjL31C6n5QyCeJ93JqNfxDY8aCIhuH
5QYPrizMA+WOKA0/HNdRXYVNIHL+4sBqQKbFcMn/CCZkXUvMdlNchfSl47c7Y2jS
yFf9+ieDdmargRhpOUNVQ8XRabkqvTJEbgVkNT2C9ajPdt0SrjFv4USrE/nGO929
I0TJnxmtpA+C64wSVg5EuDU2aNagK/P7GT/91jl+ga0Vj4OuSBLR+ZhTIewhVYSC
kv/W+J7O8tpWW8chgRFs8IZaZOmmHsMIetM4GAoXCLdgAphyDLcTFoZ4RsRsZDbi
zz5UTmBjWdR6YqN+Yurc6RpB9caGF/ww2PKnDaE8ehzztHYW1kGB3huBrA5Ppj7f
sdHPvRCCIOL0nYhLmXa3SvwhfHIMUeL+ZgkLyiLZwTey+2movcut4HF9icL0sVMs
03n9o8D06DqZ4RKgJmxYj+Jm2F1M8emDGBIS8K7mrX56ghWN3IC+cG3hXq+JdpqP
Emsvh7udrdnRfCRbmJ5dP2auqN5pkPTFSOl1QUWg2La6DMqOX+8MEODvrKs7QEwh
Kv9ekI+kNoM9tMUtQACe/4j4hI3Q0+t8VLMGx87iaFY/QNt3Mye7ZVxqHjVjQuJf
24D+6dL0yaeDu/vWnQShCKWVq3FOuSkCd9TJAQ1AtZ9sNYPLm/D3EvTGhBftXfHx
gBLQwtL0Zbyj9Td5FS/a7IG5+9wguW4oVPXykDTetLgVzC5a5optGihE3KZBGE3n
wUted8hcgy/BAKqTo5eqeJcF2qNk5wKgFbiBUCigcWulOnANfmDCRQEkCy7ylCZD
wTcbqDR4ZBNkSzxxgqbt58k0hcsuBxl5+60Kwj4rLT6/nGeJW+b2ljK3haFVIGio
bLKuxEr96uMW485d1+JpsnOG+yepmJukyeXFD/3P1tyTK2jsh9EZYG2/MV02D6wG
XZiBVgD6420nqWl1BDj/8DjcRczXCswGaT57uT5tFaUJLoPJPO0+dvhL4yc9gj8C
Iedp3C4iQF5J4kwtTYVssGu4Q+czz0CAERNaIChFdb2yQPZuYjwu6naHFrpJV6p9
nlEl/WtpX/99PlxfA4RV+pmipR78yEpgFx0AtTwwjy/DXdy96m8aamkKvaS00Vmy
UWKaLieElL4n2fHcs1vQmKB3XBv61RHdYouxDlSQyryxEwEcq1ZTaRiYSOjiYoMw
Ndpv4T0fdU6/ehrrBomJ1GtQY0KzgT86qL2vTfOInsWN02Xl+3t2yN+8uq4Ospx9
WZzlF8CVYXzlHgfQq6YD8O5vfXKANnNNm2EwIfTrd0VGe/kqtsTW6IKBm388USEc
iBpzA9bpfeaekjkCLDK2GBDN1heByjCxgz+o4jIYkGGvZQa8tbJcr1LgAeca156o
W7XGd/Ye2sm++/4BCCJrCJ7zIofG7hAFzE3GSkw3SE4ocBfN/viq2RynHT4No0dd
U8Vx3xSmpT/Vzc2qEqMsf/oxknITgeaTsW7Ep1ukMajl9+njO3ASJxoaHjLa8Z06
nMiNdFtjkS9DhbTz/LsCdkEYjO+sZXab6S7RVF2jFap+SRG8T/mpu18PnczxV9ww
HzNYE7pdIPL71TTP9K2Bc846pp39SQcBZ9OkaZBWLOHeTtPiwTSGmH9sJlHkcQVN
BrEFd3UvzQTlqQ0rFfjRwhFsarzq0TymJ27YM8YbQrseDazJ+fEHnlcayQjfZ326
9BiGnEZUl/f2vGRVKCfcqwH73zrvoPHXLAiEIkQ91H3hfLE/6Ogn42LVqTcBxhpn
0Fos3/ZRqR1hwpfkVDxNkTNw/6RC11BF7TZiPOH0evSi9K9KHObTotXEsoDT9dpx
yq0uUdI9qfAqL9mlRyw5Oc9cQBLpmuGO/VaQh5BmqGYNQBu5IL9tlWVwwI9Pz/je
1aXGuqOOeKXlqyL4g60XWy68qRfTpcwN++sOPWEA2vC/j45qGEZsJQV8KdKxxkBb
QnNLwreXDszl8F9n9/yRA8Ct6aqQXIrA6yQS7Q4OKH6ufJy+R+uIyLQZyBSMgyoB
dAYZsbhajVbTcZ2TnXWt1RhjZQJ7/KPA32RRGZLOHx/Cf90hLo0vzrELvcUMyoXi
ek1oyIZlH9J3we9Xs7JGmOQAc1bnsm2G8vKJquiJ29Q02LPspvGcNk0kx7DtOyqx
8KqHYP6wxcUvrRqOqJ37qblsF0wxiyqV8SfN585AQgFEWhkXuMUZBCZTqImj4CZD
lm9zgfeu5U2V8hLArHEvans5Jf1OXCnAvy4wcJONkIudXJtw0upYyiDTejjERswk
uPNIdeUykuI9y4JiXBuT5SX2zZ1uv/ZnFh2BICovOaSKGnNeMDHSAs+eAoKOW+so
pEB/73c8UldFN0kcGWS3aQnJ1ncgvS8OoWb658joDBBLgtmai6NwQdZCcDS/XKHf
FRlhjBbFMmiXwXOg1R3PPd9KK5K75CFbwJvAzDrDEM6b5jI8bAyCfA+yVc8sd5Nk
svg19s+kQKGe6+PMOYBXyiVI4oz/VkpYsL6TJlu4nPUGV4CRAzEtPbLayABL7waC
zn9NZvysxrylV4MWpcGM+BsiWEa4Mz3ctfx17NbfDgFBw+tNXs8lMTye0LnckFhX
KRQr3R9HgMLGVzHKrzUgoW5iLLWAjOuKM7O1CYIQdfo828IW32UqkvI7YnjxwEqr
sv71Aq7jYrvnSJLlQU1zzu/D0TRuplc7TwpwpBqYMoS5Q7mEMWti/UO1GM61vQBX
hfe6EkRDrA0F6WYVFRMdQBxkrG+A4ax5P5VsYq2DxkgdBl/7Z/1sEUPBhfI2ufTI
Y+Xd2497sRTELPWTT+957LsFg8vj0X0n7XLs3BBCchhP0GuRO7B/RpfsgAG/79yu
QkjVOqfp5SYK0qOfoF6BdvOgXEqy21amX1H8aV5pvm2TUpFOymV0w+sAw5vpf0xt
+tnTVyGBqRZ8pXcwlPTv+ZzMs/b9dQa6LIDsTPVnyJZtboxYSGYqC0t5VtrZheYG
gT7LBc6711517oBZFxBc4VCb2vyu6wjY5D104ovW/aZhH9QZ40iur/Et+xw0jtr3
uuBLCnHW6qFX2y/1SlKUI8q0TcHi8LOXob6ZKspudrDeIPq5RIjg9VZQMiPefcJE
r53f8yrWhzC/tMeR6OKlLrnryMAN0uQgCiPB+1cA9zFHlq3IrIzMmDlTX1ZwE9BC
vwgjgWwj1e3lPTCSnjtC6TrB9mULt3r+oIPnT/ykkRZseSUTf7qWW/UtXJG/HWjO
I2mvKm/j1ozZAHUSX1CRXhC6+4SArw4g/1g2Ww5+TPlXh/9t0CPJ/eKBaFTfDYYH
I9zg4uHbBEjJ+5t6tkQlEHjuSEwxVceFicE0VnjbtMEVL2gd7tVwsII1dKcx7+I7
ZeNpn+Ukk+2Qw78yFDbXYMBk80z3dvkvsEVyZLpCpHN/iHnCUj6huaKYXbMerHjd
Vm+DVUP8PvUTq4RFVF7O4AFvWxyRTcRDLIr1x1Cg1osgy1LA9AzH/ngQDOXpZ0d5
giSjTEbfZXHdO0vlTH2gNMOWHOChW/ICbq7EswYyCu+a1zoW+vXAp8+forFy0uh3
HIBKKuenIa7qWgtC5CSXfJP1d6WXE9uvGFB0gbW6r7CvwjZjX1d3SkIEdOosvEwn
pYPDsknqethrylEFLWExXQkIVLj12GeOPe2z7wteWM8zaqF7O4m0zTi2NUAkqv6P
l05mXed6JgWDbs9cofc3q84M5AW62c0FLb9MmQK+ZzESXMJhl9DE3MBA7xJofCFC
LUbjvSnmv2I/hIKJOFJEtOHr6oHmC1TWyazBNxBGSuJCNimi+4Dp6i1Vpv/uEeG8
GWtZQumlFlbYl2pOtVGKDBo/ovL+oJUBpm+rwAtB4zy8d3IbJYGwuZV4vCDcZijk
/dXm/qs1YVE/0cZ5vPqEr53NfoWwe4kmrmkDL3pqTlqIWETOT6pi2u2dqROFpad5
eyQAnuxInoGb5n3D7Tg0wDepx5YI56YErUkwx3YbUWUNldtw+ZMoDDJheII0ZSdo
YrOJuqju1FVCWwOl4mXXhSQwQD5f1HjOp3ver4BvXoaoIC7Sg1OS3N5NuS37odL+
oYTdN1yY+VMhgxpMloXwSfO8enju9+vAuo9Zc05i9yulVFWtBgh4CyqFvh94rvWS
Kc0nSlnoD4wq3GSkEXCMtIAZ95mbSZKEW/t3nN82bQQjIuAobEJdRtBiNwiIoSq2
k0Yl+Uk6nPFUPS+LQfkoBFh2Jt3Rbx8so1rCy/dyJrM31szC8p1xP/nU73YvHxLo
spvtcFmIbR89LGG/rnumak5lHfTLwSCrHiKvzGaV5zihqH39sdhZzhOJ0sCX0b0L
l0fesiLkCNeLOzURqXZYK3wPivgg0kw4V4O2PQGziXR3hdayKH3Xkcm75aFipF8t
AZMG8LN4Rd9wcJKFhvNNcw/hZZyOR4AxRLkSjyz5+lyzAGsaJZYNNtr8Y99G5FEO
PSWqcSHJssTt4A3ljtVXzaHosyz1PpaGF4BTGGAJY1JcEUNUvOViF3/w6m0VWGIp
50v+qLe8Tba2LgO7y/72b4a3ldhkSU/SIb2SBmvNQDFPzoEFtzgQ5WRBz5pLmM8o
ZM4az1okz0zBDPdRSiT2L+BIrrYn/4fcTfHOvVaytoXp9Sy8L/VTJEdKn8GJbp2s
wPJX9GiykCTe/WtTncY1coG9N01PDU6oO8WRlBl7bakp4b6QWzdD5P2mpikWRDls
eUVY5yamn66D3WUWNkiVXT3NUDZAx6kwnhNY8CIgYwm49WIfBT/qCaa02zo3Pjve
VzDh9DwLsBeEsV4mFSddsPQ6yFIQIJkW0RGFBkBFynuraEhA3dp9h8RXP3rlKrD4
mh/aqx7sqJhVXn2AI19MdT6Y12NmVS205X+7iUERTnMS06ldsUHcT7zLj8l7LKq/
Vun2DF1wApZKI+trG4h9dm9KYMzjoyCex9mTKsOPSu8Sxovm72O0gOIyOquO0Jh8
OkgnSw02ooUAcu5zdOV2DiGrnAEvsWcZzO7/HbZ7YSGQTgvJRrP/l2NSWIIq9fIw
/YYOr6HiRWUcY4A1VfrtX8xNSGeNa3SFP7jbnv+ITrZyGH3oLm7jPEU+JGe/UK0j
5r+EeDOLV0IYZbGYkMbdCUJDvg6ZdkZ8Uk7HYw6YMt8joJ2IVjx7fRdvdMQewjIJ
zOU3nbS/EeeaYAqKn3uDeNhekHsGIAvJ803OA58O8qHsWddtmzJQDPpCtWHvIuXV
Vs9BNcw56OC/x/YYtbdOoeeWUOg77HRYL4dx9wgQeqGNhmCJIKdgQOTXTTmye+NV
xaDuEL2nmCOU5wAOF4scndK9inVMMPDcFPyjza3aUDEnaJkunptRIUZ2dr49+U2I
Lp7grIvYsK6u9j5NFESBeyxUUkiAoRidaB1nFR1LnjXsJOR2b6BtOFiJU61sGzFF
CrUR3V4/AQsCwBg6YLfYOfT0S1s2H0jN4D/BK8Zfy0j3cmPwvl+pL5cAx2hxPCkD
R7z4mO53d0ASxs74wYhsDadqYbqCqVZZog+0ubZ70sx59FV0LJWFJXAC/W3fOxlE
Q1lsifGCqpJC3GHbkFpbtETwJPi1+yeHEZNjtoP8PawqZHubNnvPz/ccNXnQ3oqV
l57TYlGEJgR7VChxvg+HnC6eelOgpXQ18lhYtgaNwOtLdu6TBdH8JXNJ4GHEABTm
nsHq4YH4OLC4HsuSuDE1lUyICAZHew68Yy9vt9ziZs5ye1dPID6oihY34kEJftTj
iY5qoYqoPE8j95ghhztFoFZw/Ij0mC8UmhczNqDbMn0Di6VlzruQ5txlzzo3tWlM
XAZdsn+mLhi3S0Tj9NY++Q0s1lHWhUDGsUx2usQbvPFxH7hnIxR+tNXUTtR490XA
YZe9ArUrU2MYWn9x/v9AZeqSdjXP+JrKoR6K2lolgyoQZODJuloY5KELropbMJcq
u8HBNEsE3ph1tWCpYgLKuDviZyjoaUWuVF/EGHAHrJYPWYVihICUhv69u1hdYTMG
eY/fF/MA8qTtknCSzxoJVfu+L6dBKuLVIqkMZ6MXv2HZc/UqV6kIF1O1jNAK2MZ6
3SMW/WGGJ6xq8itiwEbDo11ZOiAtw7q52V+eUYIr5mgb+rZEps46uL+41ha7qeKe
4c20oV9plusomMzpGhtcnrKnK0MwhEWA/Im2dwCDCg2JcYINZtRma8j1sNO+9ZBD
dkAhgQLRA6f0q+tEDEnGGCLoKv0rgebUqGfENH6I7COvnKIwSGsK0S4P1xQFiM8w
uXNsDm42TpqmzKZS8WNdO1voUC1fjXTSA8IUfvoNB2+OpZGnNN8ZKSHbgkBP7LHk
pvFHUyepF7OKBGo55GQxQpzPmkrqnZhRXgrrGONoQv2oE7tDvIlLEyD05p2bunof
BXlREOlsNmlv8eoXN6o+U1AXHSGuBuWx8VyetHShy22vF590AccilZr+NJDn8Bpi
szEBabW5nCcN6DjYd9dlv14Gy/NLaYCrr1oOWH7Vip/YiP67QkK8rIllXd3wYzrY
jRMvGBP/TQDQgAofs2Abr3GLMyeUBkrtEC3awSETZnFjFHiG1tHedw2UuCE8lXFY
m4etAKf+Mc4n9htbyRXwqh16NM9l8TSZlv4yb6dDUURzJ8clCB0glXICIYCqI3XZ
uy13llzFjR0yJ57dV4/Pw1rdNPQirhmI5gnBzL5vCqOuiiIP1VY1Rgnn7qzTERlE
Vnii/tPGUgipHYAWMdReh9b33vJF1N7BCCtMv/zMNuFgAvrUEd6Ke3SfyWMidAOL
jVgXtbA0P4Vr/kQ2GpyBWWX68pAtdEwjRt/xLsnMgxh8qPmWm3md5gDx3YKgA42L
dSW6wyzG5XMVwWfBdoduv5lCa8l4n9Xa+IWPBfngSiDV0EciVPhjVFU9X3ZTr0Vv
rHmBfEMczhLZwy7tPOrS4t66zxZbnR12EB/MS0cFchQE8EHWkyAHD7wdNNwkYh3t
s7OWq59t/WKBCP/69PxCZEBLi0+ftp9Gpn+Q0r09iIK9m4q/L+6PG/IjYDfa75Dn
Pb4Yb8CoMxSCMnEjLT7VsaioSGDIqDuL27atEJHhYmZDrP4DuTpTRqF/Hy6B9uw1
2uVboxqtKxcjjC1L4apataNd7hAaqI7H7cMXLCYJIjv7aeZMIEiwr6iMZirEAIYt
XqtSxiOEQfjUeGTCGJEvzaNtT81Aa7SuwbfMutKe8CmLZwtDZ3gMESmasiNbTKCg
VKIZgPjYy5nelwizOrlmn92uKbAf1WYcb4oFXOurl5roAEnPc2P8Nu+2PBiw0HK/
pXdJ5sf6bmYkt+MsuSej5EH/TFmYIJTN/1J+38Cq2HewXPwviQbpLzjlkQ4GtotS
h0xNhHps/7KNRzCxzu6EzmYClJiLQFpGJtemvkOEdoyP20dgENKZ0dKgoBYFZhOD
bJuBxQfASOe8S+xdSc7p/dJHGpRPrIpABpZOJW9m4yd+z92vZMPNdRlKvvxL7zzS
K2wOa4RmRfUW3C+1XDWvfGXWrMaz3HZuQopgFZUDsChZpVuzl/ZOhzstUHK9Dhzz
C5BIkxkgAd9D+AFPGysLh6C84+GqhjakvqUCQ7MeGovx3vZhn9p4weXVWPZvyH3y
9+1QLc904WEVazgGy/CDnsY0r8GOEwYsLrVcMlIx95jE9JRhmT8qlXW+gXPIiJVc
b1PomNwVRfqdoj8cxH3Caru+a3qrF+NNKouUZVqtt/SsWKM3XxKx7nH18QISDugn
ZudBXGIVS+RBiJSZ/JbkYTuV2ycWLPg/Gusgj32QvRmrTslbAkOjfcBkn1z+qi+p
+8q/gzw0sSkHSwPvCauwBpWORnYSyxSg4pAQLHbi/V7a2x2jZewMXM7Hg5STjZTD
vemngOYVv9yylcuIRQbGqR2d339IMdpfkVy32qC9mqwJvZ+WHeWhvw0uWN76dgMx
tK4mSaNDGcULCYKpg+SQe1J4CfCLNK+RZdL58RpVl8IqeMZES4fhXdYvpkaB2qg2
4SU0YOmKcWatI6zvVR7fTqnoSeShpXwJ+H0VF7Gd/JbrfFRrBW/UUyDXPeyFoRYX
GhAUxMC3eU4ff+B592MIr3IMoiI7upzYaeTMBRR4QzCnZzRd7TPQAEa70+H/1uDC
f+iEgxx9iYEEHsesI+ZAxZNlqFPI/SwLufoN4TdIGw1qaKniJ83iPHLBMf5c1PHw
MixMK6EhqqIfqpgvsBXe53ddOY0aX+BiMElBw4zjqy3ReO6ex2G1Zcm/tSDPOjY5
H6Duo/FdZnHLx0z3URes6QmFyqCrZ1XBqBPP4ei6uYYtHGBvULeOoV5dATtPOKNx
ePWpLrLT578FGb0phBIp+Hgo7AzPksVndL1Dq37oR0Xx/KnGk5PVhRZYxFHFn1bC
23Ak3eA1G2jETM1zS/PRv+Jxbae7lEB91c5zJMkzg/5cZ2xjJoqdTmvdqp3U3VOK
FiE3oqXcZln45794tQtFOJ+SmiEmvhoSN2KKEF3hVmB7V76NK5JkqL7ZJgqha4Ea
/PiagkaiOz8mEwtxwIyGlnr7jenHW3P8umdgkd4pgCvG/QCt4oQGkaZblmTnIvFy
NkEVeTajNU0GfNiBBgDnxsNzj16nbJE92YrRtAoDBy/njHULptwrYsTev5NBfLr7
0ef3uA76eTxWrKzntSIgGcrFEoNB/pnKSuHgqFmXYH8vq3QpJI2habuGxzYLtmxX
umhg9vdEDwrOgC4WBuIavKT6sUSS/UlWKgKEiA5qMG4eOVSGfPwPxPjHmQ4HCI8a
quM1n85qjYxkgH3e67uwk7broCcuyyNWtS4txYWREuzzFRJwAkbBCwzCzNgRXwNO
oMbOCKx8d85lMFYbp4JAyIhJ9v0lRx7P4YV4G2zmO6Vf6uUQuNU+2ZUQc+9ONIpV
Lt0cyEMtkX1FcglULxdCBj97/jeiZ5flHhrWtSRmrIzY3Q+C4+iWB3j3+nF274IN
NevXfNVdx+oIY2d8Grdahch9UPKASoha2pHYDPIPHks47iO4mlXiKKyIk16sfO/V
/cJ+8QETzASSGdolwDb9TseZD2A23wcTics1Sg7TzjQNtQ6WDFcgWv7CoIRFQ2cz
FwPlQgiyk4lAG3R6ztup2X6tg0DyWXjnCrYkqeAIpelQYeWYdTRKS7R9h0PbjdZe
xoDFtGMIA+K++NEDm7qflwSuSrI6JiP4hMC/CD/HDdK/nKRD5pjxWixGbiVQ7TrB
n51cQQ7g/7j4fDwMViT6Pm0SGFbSJTEsSKYzu6J5vtzM/Smg8ilR3X5lAeaMO7r+
ikdE9n5/mUADzNI3rYU71EGofmcJi6oFJJc7Km/V7FReoheE9uUakr1yPquFZ5e/
JlBx36QyZyWEql9wzWOk8mnZV/bRLf76J+FT+LQEIx9p4zxlsT7Fu5FUSRyEXk1l
tvgZ4Gldc0jeI9UKDbhkAmDLzqeCKL2CTJVcrhGdl11tzOdHCDs4ELx6C2Sdw6IZ
EKSFRy9qxlN70RqlMeN97wCiFt2JWVN/xlLxfKgvfShhj5Dhglw8SQwqkHP7jx1a
TyE4ON5+6YZN6u9MXYVzu2Oagc0TdDMciejzfWcVUGpicP48NMc0YhbKMgZ4X7Vw
4qDHuHtOoCJi7FnEBAxOSOC4h/6XViI3ubGgIyy8BSkvonCfbusMvsP9zkYT3OxR
NMhCETTmeqahmcrDYqEu9yHYs2HOy4EjnU3V/SEIiP0U4crIJ1DCoHPh7giLJrjf
m9DYjQrtMwrqhmQRYGSWbGXVOR+3ybeecrrFjHTlKlF1UB9Rt6nJEVxJlFoykHzA
ZCK688BGKcjOFhVkd5OW3HKHyyVa8UvesWZHy4ic7X61hFUs0Y6RCBJg3493LZ/3
8HSYGao9QyED4Ojs46PWVnocsMcf+sVCWey2VKuSbvidsMCiH48jbKv2mer7Mdzz
bVTeGf28XLAkM79BLLOu4HPuSILaBRuBmS6a1lWWNkOV4ySsBQBuLVQWm7Cd/0nn
3iuZkISzQx8MxIf287mAMb3+5OAhWntFapYXSOyWDzdLiBAhYzj9REvA606Plr3X
LJup/7W1r1Hh3PFolQZZZexjRpNkZ4QVHABksg+XYJDEWQuTGZd4AFAI8CtONjcB
EH7ucZ4AR2eB/dtTY3WBoyIoyL+7h3VWRvHPq0z4/jyyJYLjUcVqy9sh+9W/of0r
B4XGnrN/kcbely9cGFcdkiBXa7d9CNSLW96dHUZRcX4loWShghdJHVIDrnCPj/18
R2dbkLjfrfdkXV7KbFf2BUEyUuzxAXYHCaR1xcTdCjayGGeqlzSk+KCF9xmWsuya
4xC4FTYITc0NAuH6DnZw27Aq4E2FR3Dh9h9XGsUF9HJ6L0Yf6/rHq45X1D2dCDe6
fseV6EXgwilR+GVbYPrLAUoXpvKXd+JH4hCxkbiEVMbZb5pZmmC3bdXqcV0r0AEG
6FScQrbpM+h/TBl6WO342Z55hLI/q9pMWnDtlK1pcJZrW7RhK1W2i5Fqh52uAz/T
avBbgToM9aL3raKy462F3enN6igk1D/0/SIc2Axt1+meIMBQ8bi6D1MHbWJG4kwn
meS9LHoS8rrofg7VBo3OtbdOdE6bOF0McuEFuK3zveh+4u7H2uWB9brDlrKnAlHr
/LC+phpVk4SBTwbxnwesTKA5P2DEIJMvqr13gr5Biac12MeiPqz5duzZiZk/yqiY
v707LhZEv2GkCKmjlnV/Nn+0kfSBcU9fsZWxOo7+IJnN3Iu5cKmiMh3K3yUpd06Y
604jpTjzmh9rfcSatCq6gA7ANGCwZe85f4LPGkLfCysAkk+6kDG8DCprUy8PDXyk
cGu3g1O5oGkvg8AIjoyTeldf0NhKBHqbyf5ElarybaaPXVnh8Zj4bA2bocT/tTJm
yEtj0PS5raSx2aTVWT4Rd/9Z0rDBixH6ItL66SXSiZXvGkr/1OsebGQuCKsab/uO
ieWyMvSXsJOTMrUIQz053ijMl9hprpFCChVgk/NRYK5LHAjPSdCviDhoDQhsUm8L
zlt5f67aX89sQbdIXYp1N221438LTV2pN/I1V/Sj7v3aE6OgBkwCwHxDcAECWnA0
2wfGA024O7BfVLaLefsBN4l/ieYh6/+LvPjszwmQ45mnPPedWlTPCx03RBlLwR8P
yU9SYsty4ol5T4HuTEU8dmzBoX/qk75z2E1r5LQj6guPu05wfNowR/3djR2mKzkn
jnBhN8GQCB59r5XW+V1SkkIDRqvk3pAWC4FvKKOceiNX0BazzXYZrjmIA+l9Pfbh
U7SfJdghrt6dvfqxGaYK4G+Tv6PBELuCVHt4olufvTRmXRMGKxrlaOPmvfZ11pSn
sI9sncXciBYeTmU3IdYnuv/B6/xp+QTnFMrOYEARvrtrvrpxOiBovnTPmnnjf/0D
szAMveofOihg1iSN+XtFmb5YWr2kflq9G8n9TT3L8uNdECG2Mdk1dfRQKvfhZu64
Vsk6mQCOXJH29UHI7+YBAFm/b3MN/BwBBADgEB2a1o3nxrwYb0v1KDhZNV7SHxcr
o+T0zIIidaDrgNyUODs3+3RG7ytnwLujYNz/z8pwroFbajwF9GT0nysOKLUiA+Rw
Hz0N1bwqOQL8LNMKluXn3QOgtU9p1o+MFwuwsSV5NXlIiNcrhK300/WRFpWUkEt3
brr6Om9InzIfemw8vnjlgyPtk5qUhXVHt/6ZeTJKj+c1ajw8futN07sEK74xAqtv
T1uXcNgnzBlTd4ljF0rMNsRALoDf4JGSLFl/JlHkROFf6U7z3HEjnzOI+K5bkwJS
P3Ljl0tbKA0aAExQQ+3rhuCYGko8U8nulJpbTguaJ0YbtlXm8GCtBSjzysFd2rlX
/nPVmyNVaTgpJ048bp0JX3DT9vtaZ/tAF83GDAiaUgBpR8ulSwkmxcm1wv7cwbPw
/ybPLfQ7DGh2++/YdkfJ8LaDYEpHnkvRDaWDMpQH88RZa+a9Cmu7uYGEs93mQkPh
ccJqJPLDrWxrbIakcStStObKZqyQpdvWue1F772HNoSPwqOqcqBQzdrJKFzVa17a
+2T8benhZFaRGIUssa5uuZFVlXUE5Zaew3Tf3n856TvGD2bAuJmHXjKsCHR1ko7E
nZVSFZs0XNf91GqxbwCU16qo5qkTdvs1oBd5mX9vuqF28NXmtiFarQi199HK2hUd
Nfk5YVjPot49xsFJtQ3Oxq/7icLcBrWXQtjl30VHtd9irUlQ4MKHJvoIgMK8VDoO
8KChAy1aRbAqskdkM8FElXQKngusM89Pg2YggOk8m6tcZm6AdRAPEui2sef5CEI3
6zqcQd4iiyAfUT5oltscSK7S5SXC5IsVqBL3jQ3Fs41oMXhvW97rfYhDuJN30h/y
I5K+QaJ/MZ7+DsZsbmNMLW646u9BEfblb+4QQ+LPVOQ82afUUfN1whJdgPTwerF+
G/ll0OoNLFtLWH9MuzxUZ/SD3xfKTgVEgq5S2aQV6wxLeBOlk9nGdnKelrfi3QlP
L0d8Q/JK0xO4E0l4zbQQOk85FLT24+8cVha/7ug+iE0a52CgU7xpr8PVNhwooq3M
JFX2xHznHwYAp+Soi0vbKnUe125R3UChT7tD0nDej36GbI48QKu1rDdq7gvcP7y3
7HTWEDLy6bVGWVszBHjoIxBqfn8vxP0oPRdQgeEKG4U5rexO9VVe/3i6jlDH9Q7F
R40AM7MzArGqE61W9UlWiVOSd+N2oyl8mfXfTpPDG+i8DohfF4yu346os059abUG
d71qqPtzCB6Ohex1ZCsqffEakSdo96pjkLH9s/ZuiyFTs8qrXUOyZ33qu1IB47C2
9jX155Y1ZRzJ2/ghlnD/rbGBA5xZ3MZ7Xfg8TiyjV5aNJqrAyzjo7CMI+YpZUlGy
gTo9ob2FE/nj25j2prrjTzUg71X99k9WfsOpYzoBPeU7DthUjnlE44WDXQeTobww
ypja//YkA6CJPuStRTxQHtxVrHFFaRMBuMCJhDrr6uvVyKiwQgmxBCmGH1VJGXaQ
seLAbzAgZIQBE+Kzmrvy+dNAmjc+045dKn+PBZMmUpIWBtpRmwbcvdmrmU41DRcr
EODTgeDv1abv+VNXAZvjjmvsxmXu1mjyhANU3diwWfhjCJ4vEhAkQCUMKOO2S8HI
XMeQv7VD07XbZFc3A/qTyCSPLWDFoYgj6B9W/0qThyZSDXlnHfe+7UjRwtsHyqcf
1+WlZKda6jR1aetuaBxvhRZpS1B89BzPHjFGLlynfo0xNqxyD9K+vTrRltQ5E5IM
oyZUDM2BeRX0CuMsgBvQwOf51HW3wVxKD0dB28fQxL5QzlfrenDiD41YHKzxyZYj
/OXxNq+ACQfwTMqoneuTWEmKrJz+jw0q73AfZUxnZyT/bsE5jRMOQJhBxn7O1fgs
CvNGmKNyJ1m9wCcEEhH+xTU2jYyFfFnMTLUiNYfTu9xdPoiPhrwv/7sHN+QhtKF+
98/tLBRp6A8P5CnohpPXeDAQ2f1i28NtzAHOnu04qFWVbASRizyAA9+tFn8AE/ZZ
rCixoKFzezdwhhR+3hcLpJzzzJzFxCvnmEkrSeFF9CsqYFw9rKsuLcQSpsZ26Iid
DYcUA/EotAPTGLxQ+NaUGP9QwF75och3ehKgw+Axd53ydQa/V7NGtFVVdv8cmYeH
AY9MptW/ZUSbLl6d1heCf6A97eUOQe/QuP3/Bo5hxmXpih58M2p8rFQ464wpnNDn
RS/V+YHm4XX4hNqhMgFu3Deq346JKnld7Lylsy0IcvUAnbg8ETi99w04hzP1GBs/
bIVjI2OC2ncYWtLZtoqH3M2W2W13JPgrn/gmlF68ugNwUQPxrSBVSZ42k0j5+MAA
UFAMECzfHdstH7Uv56UCmo93qtFGwguiBrXjD3FoxrLFTQrQmxJbRG7dcZ+y2DZr
fieLWyI9/vPGeMnQA9IJXvBmXKLugMBwr7OyxrVMSbxqPGW3woNLbKctlvrh0Kt9
gI6W5dtKoNZWPS3fo3DUJ6dnTdO3uR23i3WaVlAhwIpLMf8SUM5WdYR6G+Wq/dhR
I0jhOqQHoJ36LAxLeK/gwwi5IJGzZ6fRt8WK9eoyI0cE+Naj22vQsmMRMaYhLJXG
t5/DeQOe0Ylgru8jYEq+/iik+vwrp1Br3g0FUYTjO76uocpC9McNOGIN3QEezR5A
SMWigwrwr/i0x8pqT6Hm0NfjzCuiFETiIkA50ryKoLG/+luGUL00Ix7DY4NAar67
Z6xkTXGLOABVrbT17MyJBc4k41rS0DH7engC0AzDYVHdO8Ce0PDX3+7weFRKpsym
Tnm2l0xLsHnwlK4CBIj7qRN84mclmYgE9+lFo3zX0Mt5BGMGmIsa+2YsnTx3fV19
V84C1hRfioBP+A7tasqheEiXUjWXcsTX39QMV4h56m7Tdj+0vzZO2FckC3aMjwUh
KY+ZzRbObT1KOKm3zw2jRX0pX1avJJZGkVgw2VUjsdZCVDpltKsUvxzKMpb/wp8t
hsadl475+4WrenzhXzgE+848jKGKpsTcc7yQW+snyVPoknnCNP2P38NR/GuBHOiQ
AxrcqJiYHaXXBOxR8ZxTyomW/X4SZHDIGIy/2gR3gKtoMmw18NzyMgrJhOKKWuFN
0jw7vOjA4a5eg/geUk/jbBKkh64xBs0jbBG4lF5/aCpCll5nfsbfhQmCWFdTOCsH
TsaodqgHJVexA7aWoAeyXvrCh1ZvBJXicStW2h/WEYARhyyS+Km7zF/v1yG+zjwi
SrIn07jHklsDHf6Jc5+gBss7OqjX8qvkoEmSTxB57UjMtkUi08nRlMw+XLWVQMCV
w+2E5azUvy1vids3t3Q+b2LtfwGNS1dnaHreesHEZxsRHdnb9oM7raAFui7oRqZW
M69tTHKTbQL9RvLPhHQUUNxsJCTu1dd7Igxq3U/fTg97AI0MSoVuKP6nNkNlYWk6
1AuzanNarO7nldVWJM8YAgVHNbdnVhUTXKHy/u/p9cao4eSBGc2ZrsP+m74tccQq
f8ZKw8h4rfVV+Rz8Cy7YJmvB384HpNQPNzNgJ2+1cce/OR6kNH0FHmH+xijb96z1
CqfF9ZSTJDIKb9a36ta3tUbN+IjIVCx903dBE2533mTsm6rjLONS4swg65pmDUbU
t7Vx7JjXcMJ0Z8tryq/FNCQICW0LS3OUNuVJ3CjHuNK7LXVCR+vD8T0C51Fv6Iua
ltXp4TU9DOMiM9zCCpZFpgCfc36B1eJjFirGIjWE5TJRvweJA9/B7EucBMDM3NIm
t3v/SEqFP5wQ9ygyRRyjArYvz4RSRO3oaBwMAtH9vuV3z8M6JGFHq9n3Vm6AC18J
PzhbRHUgBs+bNJ/nUkHBu7NdwGvxsbwOquC8epbsBtHwdto6JTYJ5T9ZkCHPdbm9
1S0lUxFZrVNZcf+EE1mWPMR9BvT8Y84ZwHZnS83b+0LbidjnbQCGXATWP6r0LjKs
4MdU84i/igPi1AsXU7S+fH+VEgUgGkaxCJ9iz+MKPRsxANMdoGRe4XjDsWWDDX/q
sgras8+pQAViuDpLJkfIXl/0G7l3AgmRw/rxPaBmP9rkuEnYILxZdZpx0+PfdxL3
kMeJDXWJfQnS7i90v4tt58xTk9xUteW6YzGRav47hU44+oMD3BxNCKs2I4pfi38E
mh+ldiVk4QKre2lOTytM2cbZuNWRa5cf+1dMj7a6rcG9oqXAmS2BlIIln9k1iMjw
d2NZ7kZZOqYQEo+q4iFdc/7Md6HsuJotKAHAMx7hN2GqLZ801LRJbhs7pFeWnreB
du2V+NOF0aUgXLfomtizdP55mHl3aLUbEdn8bleGY2l0CUdiCfqMje35Ql80akfL
pLEMD/p4J48Av52R3Az0jo7IQn7jgy3eME+OEj52vhMxS9RUPZuVnUX9Px5Rldyh
S2OBYWKrvbbsFI3tDIbn04HdDr64dLMbSV4Zcj/fbx7sKNDFd+OZ9mgtvXKpMr7Q
5FSLue9afPFZ3GSEDtHOV48BQvt4jwGlTD+NoNe2hGK++sZlufnPW36suYzbPWdY
LNBr5Djlw/EC3YdkCEy4MuDWhWvbfnovyFnhbTn6gFbrHd5ZoWfoU7bbFViPW0YJ
kDqqnQzzHeUVreaa+F+xGzIta5gDjGoOKpmiVP2o5mxxGqBcJQRCKp8Ys/tJHrP/
KoOa94FEespmJyjDS5ZcHhOH/2wSb9ZMUe+bh8S4WDEzmOQW6GissKdToHhjLebm
Q1YgqF72LoRzVSwHbKMEHFWdPuu6MK94rBxrLvkYaFUrQGbKAhx1e9oQm9O0zxYA
sUabU1ZcXox8HZ77CRqo+Nb0Pnyz+P/s33XD3qVqQig0GEunKqLvdmUBJHShm5KN
BbqoaYb8Wr/LptFEfGOWLAlUkA3Q2gLe4F+6q8tqRlFC8JW9xu7DgltQ3T9pHvbn
zXwPgGIMWGwJrG/08KwzH8wGksJcGrjTEiF9FBPDtvpXJreG0Za1ycfZ5L+qwnKo
N9T8xLAC87GL6ixShz4Hvh0Psc9nZwD/KTF2caEzgQr78hUu423eDucVDnDqqa1G
maW3j4SphMLxpXdNPXQ3teeH0H2Hu6M6YxAleHCcBX7rHLa7f0PEftWxSRcZVk4m
/GteVkSsiOrV4WgxXCOfPMi82Mvx7hBVfQbSTO2AEQgULcOr/dcIDnZO+hPMtchm
j+5ke4dX+8/FLsVJC3aYa32n1HJfcR5HDJPY1eFKKvaDfdLuxshAY/Dzq1Ey5ere
mvQSYigQUHTCuOOLVBvJImx+bUDuYIKH6at5/cW2+Rv5T1tr9ax/rrGqRadRKJOy
5wIZ0ITrZEqNBNNCvGyE10zXL3+LTc9zK5wMjjFz6Psw974XyQwaONdamtJLedXg
gy/tfqaChCk8xqfynOuFsIBFh4h/vBu89iJ88FRJwCmwNPI2h4p9nn+3Tu5s+vRZ
+zPHwaeI93oLfmOwTTZAZW47dn4cLekI5fDYhLzGTB7UWIYzCMiCUagZY8gRTUfR
nnTzjv30CASiDBPDYHvye12u2jcWMHMjsPe1RPK3nV1xSaDXv7zFAFleusFIuM+i
eJuD8QsLI17h6cwRrVxhnApkpPrx7yJmIPzR1V5noWh/teYtdGiK+4lzLtJJgqLV
j5yjxsBPfahWl7I8IsH+NSOTVvuC17g+77a/ceM+2WLeO2z/MZRBIJQtqSOxKhzs
mjtTkZLenghL5HI9OBYZZPX8SiePjnVx9/0kOpn+RQSVTGBoFZ/Z2kVJfkhSxrD9
DeelzrlPMMRMRVdQXob7wyX2JPImCgUiW0336jhDKkZ5SEZW0fbh66FcLSTzsw6R
j5w/EKTxk1GnsO9r/PWEtZ2BkW1wwTjC6b1TQTyAwdeZ3CeHvKKorv1Kfii8tWvz
zGAXoxpihzAH8bwxUJZTFkGbI22z8sqPZKe8tZmRElgg3n5LXSpplu1wXg0nm7NI
sGnFoNp75uBu9AsbPZmYofzmRqr/TyQf4rMi9Gx7+L7ig7sl5ACP4B85IPq29qL7
nARI3fJ1H5aD3sfxCnUFGhMD7GkQdWH57+7kAk+047bZcJQztvMRQJ8D3pekMYvY
J3Xd/bw/29DAS0rEmrOzbXrGnYvT9LHk3lmCnpYBxyuNwdEgtp2qwYqZfqb6vCPo
eEaJd8QTMI7/opVgbfjF1zhkMm1nliUoi34IEesSIED50Gw0aAJnstd9+Wl132Gr
RcaLRatLSL0P5+05kRn+6DjCj+/f77vTHF5y4h3Pm/ALbuQHgGxmllS2YHPg46UN
Y0h6uXHmQ8gc5tgyOtZhlBqaUysItlQEr5hM80uMezztUlfUPEYetujudMGdKnLB
QL3aLZYpZkE43IwaVYYqLKVQRIqGbtCfenCNST5s1vEZ84TVCtPsj8rqpqPrfN3c
x0sOrQ/hDfdvRWWm9MMxzc13GTg3Fp/U5pBylXAXIgovCN33myzX6AGYliPSidgj
nWy/bWBRlEmXJVh5C9my2Wz10VbYb0W1cYWPvcPV3dHz5d3xh/Yale0L1MFMzjmN
sXuc6Lp91tQ/WnczA/rDpUm0EfuQcB6V2vFY2rbsl4kLf2tBKo0sy8sAsvduJIaN
43km9y7NhiwzaBhyfud1qaLmc7go2s8Mld8w610AVIWoRSxPQC9eIEDTugeNXIT1
q/2lDoelcwBGAweGNjN5sLforDz9lIUIm1QhwzxoSmX3QRSiA1tz88bpf0mYA3zI
cGeW96BPA6+s1AQcbKDYIL4nUIxiazs+eL8GDlAIC54TPqVeO3LTiy9O2JuVwSbA
O8+ojIIZouB+EYj1k7TOvHlLBUmFBVf/BaP9eNShHqf2asMpSZwV/Xt2GWJ/vrfV
+lKWPS+XxGSKdHRN+uSfPqu5vdrE3OuH/LFO7+gmDAQ/Zvv6phaOCJLSrDd/Eazd
dhw0k/CqKABBQBB6EMBBnnXRTP8zOd5QqPUQsWSJbs7yluw2CqWf1sByc4ouMdMa
C/0O+7PHZnZwRqoTQiW+CfwFcUW1oE8JzcIhGoqnzY9T3T3/xgIQSpNrcEOatBQu
bMgk+8fmtN+GDMV4GPQREuf6+H3G81cqyWP3S5efmmXDn18dFMA8VQZfCdgnx980
IBsnGGH/IwFIQ01IOvAsDDLOZxFtcDWQmJQo9IQKLfbNQgC475Hea6sU3CcdN81C
/uyA9AIjP5HHcJc2L0zbRPhM3JpmQd4/jS27aHHKiF2uvNgs5Oe9MbZ8G3f7bBOf
UNPK8sUIUJWr7vtcGeblPZVYR95Duz6T2KfurplaTZOhP9p6ytCqxezBve7nTmWV
83hPaXzLutOChaOlkFf8xI7iuc0140nICIfWMpsxqMg4hbFlD0G+96wWBVOeX9Sn
nEnv36RCWvdKHwcxvEsY1Y9Cl+PCjDut3obwsgFLXGp6lErl4eK0UONjPZ2LKJCn
P1/CZ+xVOgSr8r8XHVm48LIBObzHrVJi4LXigAEzRmNwERROykHlc7j6OgpU5Lui
6zSPPaT7tHpMFpvAhe/d/z8hUvLUqjZq/lfpikK0iJiKy/UB/loZm6/+xKZngkmb
JDTyWlY59jfjCy6yOqzjHbdmuzqZ3f6nLm1ENNBwWGCQBcHHjmPmNWUjw8Xv34tD
ccUJlNhGizhFQpSHQKORTTa00U73q9uak3fkoLATvqEEhZYqJM5cnCmeTQejMfn7
f6FawM5zRZXbuXZDTOIpQN1NZzy8w9TGF3ij5LFRFp9Dq9x5jwbHaRLlHOcDYKJl
v4R0HXU2QNqeCc5W1F5+23Cn/noCL9P3Bi+tj3oRlut5NkABiquld0F+CrpOaKL8
mP+HPy9cN7dcRVOLBPfKbCm5uyyTwpyWHsdSIPzua8wvyns5hKM7s7PzIeMGezil
rzlDoBnv87399v1LfVQ5UxxAMbRsQJ57RutkVyw5RGz61eBMV+NoeNtDAYbAXbuJ
qroO1Gm+fPPmmMpM9pp1Oq6WTFCaRPJe1JC1PKcTtwAPeRzGYXX/BicUqC/JP6IS
gOOMeGz5HFfCvw0JlZ38PVv2NsDriTslVJEJyb/HlEn4+QKbkmRyG3voPjI9UgQm
FGxEPN43CecYRvk0IvQSCY7lPIgJtc64fgyBk3H3/xCI8tYOL4bUaXB4uT6FXIKb
UpvrgcbCJYXMXm+FmQTg1rO/ROLWSR2pJeInLTKbf3/GYq5VtOZtw/sgPqukSkmx
jnSLGROMX4Vcn4rT9A7oWAVpS3DPB+VMNHRfvvWj7QStTIFdVMHPL9x7sdHOAw6I
ALH0iOH2aQTPT0lxk9rFtbA5AeJ2Dp8lxv5g2KlxuTwMo/Ft7QPnrCs0Ymmuur1h
euPYU3KwpXjUgv5gD9za1qDhogSlrpq9DoISCEhJiH812Lk4Ms19SH7+AwKys54o
837faSvmDHA7L/NXKQODpnWTBfJ5DaWwfMSoaaOOO5owbY2/0TuUVAlDkwKKZuig
tEhOHjucs3TA/JcP1RdbO9SqfBX16A7ekzbwNO7puMiQ6mz3wI2/bG+nMm3ucBHG
GHIP8eaHek6VlCOV/uU6NhJx6etxA6ZotJ9VHg/6nR5YsK9y9XTPvcwKqGTMx9dP
rHTVNsn9axnoosHbJD4qvoFfwk1sy0lEr2D4v2Q2irzQijhPHBINPqHYoTZfrk12
dOSpgeNWpOHfIu3wDo24Oiaa854wLSieubKuQg+NF/3W+2t/ndRL1jI5oA8vVXBc
xmHRLlY58KHi6mi/JlH6e/OQB38N5hMPU6+HuEoRcnZUNhlqj8HCRrMWiduG+7pR
8ZBaqHCYos4Xr+d5lH3ZQinpkNuzaqLVtUT2DX9jQW8k5ZNlddkKtblTgNVaob6p
y995hgxoUSJrPAnVXlHynFR6PAqQXAhdhrGjmhSA50nX5LPoeqAiTIPdM2/g7w//
bJ4/S+xB8R+8q9Lird4Kp+xaxOjKqekCSFjYrUrHs30Yy6Hp387EYAqxzaFsc693
awjH9NfdoEgDZmeviHltIGBeM8Ou93x9+9rELYYjTIvDXzXGAw9w+weSTwFIyoKi
V/hneaaNd15U6/pXA2RMk6jB1DAXcsMnpMP2G16lY0rU5iN5v4Ip8Vg/qcm+jplB
YTBKZ+3Ss9jsESYNGM/76106mCL2OanBf6Y9TQpwXhPRSNUgxC1YYqUz9Ht1/KXi
HQhDSPp/txLfklZbmnWTsuiVBxitsUYGsDvL/jsVWKWQdRT5XzdfF+dk+ulS+vyS
7YqYWS9rdJQveymRC/0ajHKNsdrnhgbgJ52SxQqYRzvfnhLelsoe5pb0CgwT7xGm
zcu8pG158+bVowRsa6TBOQEM+/OPHZwk/KOXKN7oZfqt8cz9zvKLn54L1UaWVsr+
mZ22Uk5kh2gdwu42YUqFL+4wIs3u2MkEh8ieOjFkH4uModMQ+56HDVdpiob4MRg2
LUmI2NMoTI5qtgrovUpGKmJJrDmzIv0hVFqIbPDeu4bV8cUc5P76iZtH3itSOABY
IR7zD1kO48gka85/yYDIVhgGYROjm/nfVvf7ea7T+axoV/osuWaPsiAowExCL3Pe
FEIRqhAeLyZAu87yJxR8Y6rLpA84iJ+UhfOgj9rRjJoppVcpuh/+GnEDdWQ8ww01
tl4j6rLsA5n37NmALYVIw1bwjA2e5gVt9V5a5iInU/fmkqgzFbHOyOhnXkrgUYzT
0mhPgJU5zeVOTRZXYx6E9ajP2kFq1eiPnrFrkNh5iSegTmzNe0OU9rHVVX8fsgIe
ffYbOZQEThpxqRVT9sTf7g+9/PBc6UlssbKg/CVbLsMuuktZuXuwkaEYvxlFZ53W
zH+USFC7aDTaeY6LXZas0DkB33Gtx+Dmm4UCMDQ5dorBdoSUhmfyuE+XiJVGDHm7
in09l+kkvLANgD7Ykw0//+rIjofMKYRkUrQ6czXTXErWXsmdMU7S4oNh24gcf/68
W46Rtpa3bjr0ls41iYCtIyJqojMO3UtRZfk63T8JQ515oE2+T5pj/jXsqRZbI2sP
meHQBTs856HLWEqFUWYaTzZNAZORWm7bKh9uiHCIXoaHp3+F/qIwjzXa55h9gctc
RU/6te1a4y7DCyeNf80JtWoGajaOClhu1ZmQUnsqoUmuF7uRiaEWRoYZvVxRhMx9
MG4cF9fHNCsy6mlHjWiezaZibGGTdkyz7SGYZIrXM6ONDxVkkSiH7019HXi3Ut04
Pe2XRXsT8snJlsXTb1TdZGlTYCH4bap/QYN9tzfscUCk4a1sYqKKFMrna0rY2jwD
/34jXYQFC85Wd98g9BJsmS3jtxIAdno6zjG0pDAiOzFobVF7FR0vnqwz+JTHpNjx
lkuLGaKEAtQbTvSPUOzEhJr91q+03uTr4FP7uifkOTjMsAX/BWPYQDWC9RlK+8ww
QRPcB+O2KN11gpasHf04+daPtDQPWxwiODKGCKzWAR1OP+vchnyUtwXP+QyzNjqE
nBBbcFohDAy2tam2ATryRZVB6jvPcWQm/YhVCdab1HTl4PAIUvy9gsU5SMSTFj75
DcF/azCqF2U0Z3PHKOHHXQiCSlpJXFLOW7+Up7OVYW+MnBMQy6ZXFpbJtnQh2QVD
Rv4MdL+irx5fNkqNXE4a6c6xZ1McI3rDv9WPQkIDFxXxg1VMVb1+9lbUtmzuAw+q
LXacNDZK8jLgpYAudqJDQUlMCwOx0HtT81bMj7knr1f6/yUSw0yQNljIM4E8j7y4
57iMG7hzfnSHiCWQMElt7Us9vpUPZdivqmgco4HxEwnjv+PezSvU6Qxrzm+mBBZS
8Gl4Jw8mp3O6rpLW2S6AinVkRmUmygxRrX+6TxdNjsyVZm3kw/2dquVSji02HK8Y
dpvOz3+GzkgmCj0f2TceXitrm6CZH3FegQOL3VAJmjEDAfZUnSap443F04pEfdR5
O6yhCMSunPXI29uUpT+WYIS5boUSVZGlOc/crN25c75EakEkvtfmIkU1wy+222uF
wUKsJtYzb5TCOxPHaGGr38WCyItpRccKbUpdGGvIW4MLVKi14D5SesMqxZ+zPCgL
Jm26LEei9SspsENJ8jmfZXZmc3amoELv8IJ9m8+4t51mTfxJ+Fn21hLZtJ6PXdya
L1SSKGUFywRGdqdbRjjuRVE1+N4aBpKCYRKGcIf4IYdJdhTBlDaCS9LGyB/v2yXY
yIhFI3bDNBCF+it055J6BJ+Kxw/Q0qsWEBgnZ7t6xKWx5jtnEIW1ey7BccGwdacY
4+hEkScXkrJAWWUqO0QZTI5zUuYW3ev54OgUiYRI1UV6iYCnayJ7ZjJpdzz6jrCH
38sdQHdEXiVzoaDVQaopa+1LVgo2XbK3FMBaB+/imeP/ei3yGvXRKCojEn8RTkNk
L6T4seQ/OCoYgzTVI0ife3OL+OGRCBSMuo0zoMNnmv3jQtwRBCEtaqF5Vk1CN0gW
lhsI1022fdzUiXV93wt8QR/6TjacCexo18mFD8ukEtiThJdyMTcj60sL2ygvaIJ/
gMCJkjCIkxcccAOABCYqBAaLn8vRaCveysGlh+5RlbJVfuP7LwR+SU7BjlYLh1P5
2TashtbUFSSUXQ07zY/cg2XY/ujXmX77oqylAr5YPoBxpQlmf6U6FvAn7HunQqHJ
zJweY7PUYWs4eKpLsV4uOsUn1xoWThjIiGtAl3wenprwFfsZ8sc1nmT9BPI9dlYD
Jitl2eD7jtfV8gMgTHYWI0SukXvC7q27kVbT5cIqVWqCsETr5sjlpxHEE4OzQr2i
jG8wtkvz/VBjZawh8pxrWL1u+XLZh9/6IQdAxrFxQ8zvxfMOJhyOjceGOcD9T6Hv
kTFFI9wP3FQwiM4mGE7xfyzzJZHQFQrgnoCv7tu9qTtPqZTsQG1W86gn10mjQ8Cg
5eoVwgftewAqEmn5d2/U8rYILV1s/VXITljkiEbQ4PEuIBhGb+Im/w/y0qxzTjSo
GMtlWoyBGSGumQLTOkYnUOkE2iT/Y1I15JKURYpJzV3vzULkKLcMupZPm6eSyEbd
0nVeOOjRdmPUesjHPTSagYTPqPbVdZ/Vi9JqZkbKr0mXniXcy8ex2N71rDvvN8Au
bifUAd2wbK59Ig+EnKYtjc1/SVX80i0vf//LequYoyOCzEtP4op8NG8Mz//3adH8
Urom/6+hnuCx0yOyZP+wRmyXmDVkTB/GlKUKAtgGEJcdhtZu2SpezU5frp9+eNr6
h5B1ZS5jstcoRK+JP+XooJgYzKqQUxjZBxDVVeYNd6KHd7tceEX21803dDg5HRfs
uwgVA5P5tYAxCoP48OOKwZP299J3/2OYY/W7nUPu58QcEBXJ8DStCBV7QUUNq/dM
y4qWuNQo8al3c6STV1+7hCG9gbq1sc49YwwNJua08kyH+1GQYTA1Ouc1xta6hjQC
AIpP8hl4gEECZK88r2Y8s8zHf7GN7nqeVmKyzGf0zAPDF4d+QRaThhM4PkyqdvjJ
sXzlN2WZRY5aPDpToA+qrRxS/es6lJLc453ycCaElEMxosOHfL0dAW0G0FYmY7tH
hZyUgfZCPVAMc3mmN3aP+hEx26F5z4ewT/fNTXvadCmw8TRTYS5PGFhq0hF64Tn7
gVfGvtxIXhaM0J7L2UNmK3vxNB2q5vdZHGNrkRW74SFdPoJzh5rIxUVtB90zs+Iu
MtH97kLJcH73Tqg3LpQlfHWshPRwRJF3d/RluDeaLsA6M+N5fbKxbpBzG2JL3/fM
wZyfnQ0YIY9otth7R9Ym/Hetkuu9uFkGfGkG5SIxBEwE0k0Bh1d2WaU7KqPWb9Pb
clmMC8edyL6qQIXci86DU+owYU7Z5VwnQRqJs8TcOoJMSn/KTwz9434tUxJpytC1
aVUO9DjkfiGNQzWdKR1PiJZN8BoxYZslqyOYYUv3SicoKNVC7Gryxn0eJ3R6Ii4V
Hrs2jkqvXlF1djcePJQJwBQ/swixGn5uKYafYxjRllVOLfC/tU+aE7jIGsiNCd2I
kXRZYJNJDrCBee+pnmWDN8XR56fdMF4MolVHEPJt8tpJVnepnCZePscf9663pHvG
nvYdgmLf5vYQghG/6nXALwKNoX8DtFqqJ/x5zvXlwUAduyfvjSuwt8StHoxyeJZZ
rDP/8tglvlTu0+zFOeYT1m3/SW3imGhFlAwuvOJTFDeos1eXkMv1MFXKcEYv+/Vl
AzhVKZjSjUW8NlXiuAYXHyGo2JpAHYIz9hjQ0c6eRoQurdsmTyxY1wDMY3BbC0Nt
DdSypubg3rvnxsX32co7Kie7sExGd69D2gRk3DVvYfeNvdY+zE2ZExP2vWdgmC8n
jevtO6sgiQ9/oQPjTnrfzWYdkh1hVl9N6P3oPDlCYIHtoFaUqMGsph6pQSpSRJgL
+9jCUQMCskdMbaLddWJQptXd5MoOhm8uXDaqZHGpC3pwADHfaCHJN7lIT2xdj5ci
TDkInfMJY5pL5fmRjur8GrUHVcpJqyxoZuvRmtXf2WhDjZlQSgcB3hkpqbIixmDV
+ATlFgqHNL5TbDatYVA8WSmU2W7mYcF1I7IiLECSAXxHyDxvoozP4GLy/mOFkaRt
EN8kD8/sXfOnNjx8Ol8Ya7G+xBb2GMZmWAkmGMEvG5mSDwQ86AmRGhbYgywVjRkG
EUSRoQab68ielYdk98JTjoICqGHoPGFJHz6vumGKiBv5mjaiiIcE6J6m+iOF87rv
vg3AE4Jxng95PqsQK7s/JgOSRcB6JdafTgdBYCGZP6J+1/NF+AitgHzbFcschOu/
THC5isyGt7Eo1MjMPMgxugAP2UQFdVxG8ckqVD1pFs+cOw89MTduvPGs+AufjmrJ
U6l7WIiztonysbuEiVlpggxyl11a1Pql3gjT1cTaA9pc1P0zjjnq798EAjVmd++s
XW6Qu6entAeWzwslbF440EqNCvoKeSjy6/bHBTk6INHt1xjg1ZjECJGDn3Qo5fEe
KBBx/GX+YqJ0jKiKgM6sqsmzb1LZR+GLro5vRF+pdAVbkcpdnMOjWTHnLWTGKVjX
TExtmS/h5EGJLa8SaSscTeEefGxl7HurK0hUlRB6EHdpFB+XLIPIqqXtMRMmzLj+
9swxt33jUe25AeJNhaQx08Tzr7mRlMdlkoziqQm73uyQ00WIBVBs8rn7hn9x5DU4
ZP7Fa5x24GYJ6vUSMjQDcPsvnrJx+56l4eZy4viNhFfALOxOYPJPRWRKtjCpd0HC
MkcY1NSR7m0ps3T/p5LAcyqcnK3UuTPl4lc1RsA15EO8jORu+Cd/c5mFSh+8FZut
1F7GQt2Frsj3uD6p/qugzYikKTuBb1HDxdT2Gaq/WoLoFGrEe8IsU/PgFbhU0bMx
b6XhF3K/XEEKJBhzoGBh7vL5IIFWn7KUZPuJFBja+KErtX9RdXOEQ8rWwL4UXpnv
HjuWXHMA+aBcKkhHWKbQTO66DZyvpPF7qTwiXsm7My0J70i7hJYtf/4qpKy+tsC0
VfINFRXVDwZ1dY8UhJCaydt4f3O5Z4oNGxAK5V9cI3Pz8rIoLQz+BBSMCK7UAOo0
OIzy2jQJYk0imOV9m5pneyuI8Ht5lk7DL0os36rztqsF15VzE6ODhPWZbEj2G+Ff
bLu8xOsFx7uSyAty5ASr9GhlRX3E0mtYXvFWDnE1RQPRbSD1i2I5x3XXpQSejjDl
jXZiBqwmofJZbNBP2XgKIfc4PoAE7+BI9Laxb9ryfKywl1igARPrz5Vi5j1AkN3W
3QHTMPFYxsx372dCIsbqQd12ITWy4equmBZpcU139dOkoh/YcE/ZOyM+kTXH1vUE
VfK8z7jcp/jFvy+xKSAGCZOFeSWUJO+XH78cDAoMG7UXlsfW4Xg0XDkP692hSTl4
PrM6SGQPPQENA4gpQlwJOm19mExPTuW/toR+F6JYDupB2zesbftlzJoCYOHfKSAF
PwVhuU3IWF3yzCNSI9eIrH3FWhpPZHEgf0W2HBIAn0qZezFuzlm+vzASqS5mgnVT
UAV1V24lP4xqLn2sAK7yNtrVcNWDT2pzEOApgJR6696tvKKoef3sb9PDKG9zbWx5
6MVnGSXyzaV6PqCwYLIjv0BdgAa/NT383Gm+CXpbdB2nhLms9gYZyt8EDfvhF/N7
gMl7Qu9T8SJc2tOVYypsf5PTsF1GeL48RAl8AOYX9FNCt5IXre7JOG2CtY2sNKOr
koynUJkKGZ0+eyCBsdDknaSknumb65i62P/4h5NX2KRAGnmDcFjChv8vMdfXXt3C
VFWS5RhizF56SoX4YwALV9m0tqnAnLviFHnZY+oIaDJkmLrdEzMQ7fuxtUByOcML
PsS0DH5Hh1WXhY+wmCKYvQY/cuwj8yuFuymg8Oj94QRPJruaNRfCfvEoIt/1Cq8l
zKz5D/o/YOkvvhvtZHWq8NctHcYigK3tfAW7q/0ENZOsJ3oQTKm17uvgZ9Y3IVBZ
P0yObpHHiEI/AKZ+cV3WjtsFIHXAf8mkJ4DXACpYJxYa210cb6eI8fPcpZIyHQmK
LvmvlL7Y1iwCQdrLiNbSXN3peScNAgUfOsqj3k8xnZekUApx/sEHu1XUqUgr132o
55Q5lNgq77pWf3R37Do8LVSGOxsdIA3h3bQtYJFtcgN2yzXDwLWPlXo0RAIlG/ka
Q+17KjjXph8uMfsf3+shI3am3z0dNQJOZ+zwIFStf7ccM+ewIyhvwCbRnB4lFMPo
xkTcocU7p/dukNEZxTDVUleHR5GPMzMLmw+a5WueFaoAOcFN2rEb4CANfW7yNQeM
F8o0ky4Aks7PK4f/NaChcHyP42RrFUJ4cPV35i1dHmmXc9MhE4KLZ7K0D0OKIilQ
e5ohNKCpQkfasIS86YpvICLN0ohk3ajl1zeIiyVEYGLWmm6KFxIDAMaCj62C7u4d
QKWZjzgnDzteuL+BrJYwxWjvWsZ6ejKoYiIIo0oUvf3vLcejl18aiG42/S5oJ/4e
iNuNrQmRKHlJCOji6mW3bpQEJmO6aOOcOhd9cXf7e39n07AvgG24lE7GWr3jzaop
Ssf5IaHtDmJMk08LnvaONavVo5TAhtTKBhFvJ5RNf/LLZZ7bYmu4nosegTPMXYE4
Jr1AG4GcnKm3b+nsu4yTilU1OHBnBt6hX04/43kZnz4daFGSYyMivBUEVJfaplM4
tD64fANfFM1p5x29TZkymomjRujuIiHQLtHG6XhGlxqngo2mrcoXYXcvNBRJGVu6
5yzYjm3WRi6xDsPM4eXyMV8QfpXWrnFGu8+vm81u8yTDlxx+PZpiBXLo2P8DBKBO
M/hO1G7AKMzbUtafg71Ib5LF8oxurGMCCVl2ligqQD+xpYRsNyXuPIMDdbEFWzgE
O1GfUIk+R00KxNk176iJ097uwN94F1bPqHou8tYYqRB4saTnbPmrgmuOzzt5EdQp
VCMMtSVpXINbYXGe7VHjCgADUQWjX7nKHEWyNeYZh8lnRX1uJd52ID8u7cmtcEDX
P6POgOYD3fmbvq8Q2sorRWWfiHu/66U2qtHpy1VosiivWJ/tGaetQVMIPgIxDTIe
e0lm6viPqg842G9vNvZZjTHXDUkLRSZ3BUQGhXbBO42sd9j+YIRJf+TYas+pILmb
/wXff8r3y2eP9abDzb1Lvr4yAGuFkwlERSmtl7IpvDAIglvZChdbzLYUmqqKaAFO
rnL4sDqIcei1pwFxzbC0/wrRdaPX5N9bc3KC3NqtDbYCP6a00E/Fk/yM7mQeKcDD
d4dO6M4wWN1lqq10VBpkET1lprlxCtlnibsrr9KN70Iu+0IidGLXpVFqeXTtmUiW
bD7OLb2grZ2qfUOaUYHdc3LCrnuduQ3ysrxj/D3SrdWv4UidrMzJ2x6cRdz+WY8Z
udFvXwLNLOUtlb0+dLqw1MLuP6B/gLhsuoBy5GX6+sN+3zItBgi5nSLA3SonsbWn
gjB5xoWc8yCsD0Iqk20dAfy30hcS8fq6hqSltP2MWBXxYViafQLXw1WSSxQN7g1P
SS2zp9IqYn2prSNhdfq2p+UeLj6ybf/SFSgjobGmZaF6Q7A48UKyTGMTw7eaPUjP
lXENje8zUBaih91oZZ6Q1WX43LRIEv5p+gPEIRtH1XY3MDwy2wPPqS2UqVPhWMU7
ghbkh3xitvQUKaicj+j7PLa5VJ9LIy/PRD+PgtH1rDfvihGov9/uTAUTWDlNYrx4
LQNRAGcnFx4xWPIQlBv39im935WomzExHFBXY+aQU0qH5LgCwNn+sw57aF+IpgmJ
yHiEXjXrl0m4gQkA23CI/UM4XjjlUwaE67t78OO2ORHpC55v2UmdF/PxI2Lq5gvf
fBSZcT7xZwszAx2gji9S277faOpUYKYVU5RcXXiTIwUOkMoUhUWTwSKUkiNtzav8
LAECHWdGqHtMbOub47EwvgU9/QDYHZojOzxSzde2n7zxXYei+BrPCf4aGpXLTr/b
8yujDZ21QfgMPuWUFmnph3NUCjPuEQHoHWw8mei4m0bpbyixuSnj+W6Hqn7n/8pf
R+snN9zw3sITOomA/Qf9C0XBeO+kPz+299h/DoWjp39QSjWKHp8r080tHDNxpIUJ
J1MlbYicO6yg9fmlX4qwhSWaOMtPn74mkVEluP8VyHy2JvJEWjh1iYL3O1hmp5gF
QpvxjZC3hi2FVBPa4+8FT/qNgYlXNB6ikjuKCbz9p7IOTpRDf0mJAMIcMHxxxCoq
Qbx5QAdafULdCqdB9n5zdgykgrb4ittSKfSjEsfQSkj4TpfbwwuqKuyriGuhiylU
Pv8mR24Y/17eRHAhi01MvwLSLcS5ufCKQILJPNgZ/gDcpDzSpq2Rvc3YFM+bXfvU
SVYHgPMJJyMehAK9uIX5N5JLy32YSznfVfj3RT+9H/JKsh/nVBj96gWDTDoHJXWT
OyUdanYAWK5smCbnSySiNlvrJl4FJM+1xocMMEguOVjc/TVXUMZzF6IjZ/YhMdmc
i03avKBx+pCz1/asMBc1fvi9OMSbIPLclAEXhe51WxuSLgq03eXdnFX5FT6m0WhH
wOZOtsWLg/pkP+weLieU9do+8GX36rKjyol0qGTD+HWuGOGKJBFnaBIGJCqt0uXN
904WJjR3XCKl0jSRI9woO6X6par5zMqV4GwZfIDHecWVs/geiG5DlsOvf+04Q6Pk
L54xaWDqYIV451nVWz6SpyFwwnlU9EBmyFhjUcIefLeT60TwL/lWCZtfMEaBZdo/
xF4+5Y3tZRT89epbqZmFqSuEzYnmMG28qmGcyrkEPgrhlDqE7n4J/CealODrHa5u
touQMrSQAb/NJPZtuVF7Zxb1KdwFdVN/oi39XWxxrm2P1nzrFNSm7LyFf8d3uuD6
B4UqXOaCzbptkt+D0oFcff5TA03/EF0Wiz50muAjGZouVNgPZXZQUNWgMsPatGm7
0AdE3jTk9XJpgWM7AMOi/ee5mqzPTbL20HXHrkUwq7KKPH/eNcMB0K5Xv0jBK69c
k3NQ2ckCv3Fq8UeZh2HXebQYKuB7hILxMZUGx4J6FS8Ft/QlxzHo/0ZCo302KiSb
Y/uKeOWH54eIuE+Axs4loFqtvqqIUJltOJo7hFfvMCaF5TJhSEaFnYDum7YwGqrj
sjLDiv0qOuv0ntL7dd7g10qj0Huy5UVVo/EtaXunwQNbLyiOjrZLXyvsuNNMzdss
JUTJTPrvlhMRFUVsjFS+a3ElOXvIXCZTlAGBxcaUVQufaX7yXDfORwm1Nx2l0b/u
OOizCQ7OhW3zZ+i9fWeVkynIr9hZandQCYQ2yZb8IabR515DAEeIFgOCol9rdVLb
EEYRqsnKT9s+dChgf1HBPDN3w5xvhseSImOyNQXf47RxxdjfDWivjly8zMfQXC4S
54N8N640ox7qc5ey3f3lHf4IJlYshXMkt7q/zKS/CKyGKQuCLWFzWBUzA8kIMwmu
iyojHXsRo+xPdvhPfAZB/pAVUovFC6DL5F9mHrPkUqtu2/PfGqnszZds1Q/5pA5w
w1/QbjM7Il4Fims7fxPZoNyR4vHuiwtT8wqGECkJzkt5QuSWxrVRUKb0gVoyYA/P
ZckXV7aOCgWKGXO0/cNzjafyATXWb+NTBOxs358b57kiYo1F5rC+2+d8DRvv+Om4
Z+B/jpJGMhJJ+zX9GnVDZf5GCruyuGJ/xUSnrqWqBfoAjVHiGAEkvOp+6Zlbhftt
wBRoMdMG9HZ89uyh8T51MXZuZ89+Nq33yMU+2n9IfIJuWLUvxHJ9FDGM/wLHUbEc
AMRgXT+BxuVLcXq8xyfkNw8C5JW50h78V8qJsdthP1zL3OTmJFYSVmjklmuJ8xYE
84bzptcqAhLyIq5hvqXk78eyH1Ex+Oyn98bTcMAOYqqOpPkLeVZMghWwxRveaTP0
61F7L7VYPDGlFPB3nvxJJ3asiGEcAnc3l3E7DX+tbrtMGF5aGmwXNzOthGLKgFr2
fvL5OAvgWvA00c9+Hgbc+3EoulWPkMLuI9qXwAWBZw5uY4pEUgsWDMqoD9kcH+jZ
17DckNe5E4h5IG3/bNFLAbhFjbBJVbsluRGN9ZNsLCbl5JTfB4d55FrdOFmjosE1
bpwIF5PQ0mCzrkfDwKT4wImhulK52xrTAsojd72oWfDsZbCtEhlwk7j7mEwCcp0X
8CWOLlZyRkgTBnKPSYUKWl+naBoO/nn2trKe4PtRJvoid9GbaWBSM29cQkfSE4P3
ue2IMnIR+5CFJBOf6JWsRywvW6Sle03tX8WjDqueIVnTU3c6OhFgflP8E0KBCf19
hU0FcH/G4nOfAXRTlzSAXN1Uc5RPD1bOBY8lQ1WMIlrg/xCa27y0KBALLqZ682vs
UINaZWWMOtxE1VPLXtpXKq23zGwN+AoT8s1hb0e+f/zUIrLtDQO9jznw5kdlPx7E
iczfws4FXAIpVF6ElWOwv4S9BPOW3l5p56Fva27Y1i1d1dTraADNKqMb3VqC/7Y0
PrYf33Fjq6BOn2wLnUrJa8y9tFPhv+XWgLNCEtLuvWtKXvz/elUe2VyXTsXSOmtE
N3JFvjyfhudDi3kmNEA/2DksQYdpGw8/WE4xcG+tEsVeXzl+fJI9xKRhZ+gwkRHP
JuCH9E6L831Z6UWKCd1LIg4V18xGH78jo0W+tNP2eVDlmL/tKcDA4k+DfrsdtVSj
dQjGJTiUNwbxyBuPVXZHfipDuZ/kx5yO/CWnJTIpCeW0EP3YpHIHEzUCshLaANGC
Qpx0t3pB3C2K/r+tnk9puatUFGsq2qVZFZx0mEZc4D4/ZvyMnQgCOZk0aVW3pShi
rg2207ruR7oBbdo03CTZGHHK9O3JhMGaflb66buQIOTxOlZZrPTFqtCdL4U8X5wc
QoTz2T19ZeB09eP54EzeUkcdbmMrPyGA8TWtJlixE+RMWw22F1N5+Ira4L9JESVv
g11t+YR76qQ0xog9S1xoTHSW+yMOaGRl5RUh2bXSpLzdJhHRK9QlVRKFos8wcBua
qOBmhb0ZFlPGpDgSDw4XT+iWi3zIXOIJ+wMl8HUDc17gGAU+ZIhTxgAvwGIEWFe5
oC8qOpCpuZoImJIDsd+2csd0WSZ3JMqRY88/q2fb/ryLZv4z7zVfjTVYS8XfgeWJ
HG3yFSa5vkPqIY29mtJx6urR4u6RHArQVx04x1xwutDXPi0bEmmvW1JFC7romGqk
IqFlrhANXAjsEyJNvfEt76sCq5p3/AaPDvaPcQWrJIYtKenSqqB0YKN/zGp7EUm+
wCukBZGy/Oj8+XnFvTxFBcOUkGPuIP+U32p63ujjno5mDrvRB+tQR9fsU8NFiaip
C3J1TvUe9/117z7onDFKyO0o61nXrC3csd8OByvg+YDBIJvSaZmaP40uQZFHVGZe
2PW+BBDyAVm69tcZLZKClzk0S5PxlbtZTJWiQfvStM7uZ74kwH7cmaWOK4ZC9fG3
OrGGI92BAZvDBxd01AgOUWJAn+XEgAPP2ha4cHmvKXJo+A/1iZW9eC2HGs8Uy3D9
AtH8FRh43m5PATMlccTAQ3SnM/EJrNJvbFKIzzF9EbNpdiIJFO+B0n6IPlK74TWt
FX8bTEAtUOBzsmrJoU8OJ0Wg+lEhG4Q/EGqKkeu35yFD2CdHRBnOBV5Nad5XlGQD
L1u97RZPu0NR0C1iuRYNCQfvc23bCyoqBqWVbDIZjZAYipVDSoELcE1JuE8l4OkS
CW/QZcsmRQbEEm8RkT8OeYd7+OKfY62WisH6hulKgb51N25+EhuXaEKI8eLg7pFl
GhI71OAAsyJyDh+/krY131RwslPs7WxMzMEQ7+kH9hSXL1DcEmRm+SCX/1jtwXx1
rilngzSsoCiXXsXnyPzjx4bZK+jFm4VU58iM1YVf1lUbE4RWhjKwZKcIlcunvtVf
I0Iy4CPWWrG5uKE7b+PPUmEhiGckmJ9kvhuIfAX7OxP2Px6ZeX2xi8rZgH1seg/Z
zDseQPbfwBGUva/PCow0rZ9MnovTpWzMV4Y+AGc0zOeG9iYZGMFGa/wgDyu0HZNI
zLqT2WhSU7iJj+ym2RV8Tr/e2zaQ7sZbuypAjTcWUIbOMNcZV0/ehKt4YK32KRHL
6zXZkdtmBfOFC2JRX7DQZ3unA0kqikraXP90Lu6mQs3wOQRn9e6lS3t7lov8rX24
mOLoMttP33EYvhqg2CTIPup33GUsDj0S9wW4QKKni/hDlllMtSoJtNqGhPJLbWUB
sK9FOvlfL+rNFl4CcdFcZOrpKNLoXYoawTkuinPXv5k1hks4imL/rl55GVOT27nj
1X9jeBXof1GASMCHL2CF6KP7g6pvyGivnqYy6Ym/8DjIU3chXzkm/iA0n4XfU6HW
BaQ9oMrgkLX+Sksy/9tEN281XOWQiqFFmngr9okFEoIaJa99mh7c3f++kMr+Hxwh
8thB1M0TH3tlmNHKCgPVFsKjIAidiSscLxCRHwj79MKOIpQqkttc1Op7hkPN/71B
pjh7KfB56rQqdsvC4blvYlBcCEhiGMNeys88c11h+PdrnlzPnfPasZJvQn5jDyjX
/+Q6FxqfruRu+86pL5hsuZg54YtvBJ3T5nQF67gr7YKfuBmJaAqFNu+h7s4Kp9te
g1NuMIfs3tWx5v5Xm+v3rRXwfOgahFUjlvZrTx5KbVMDGDZdwqVQSvoRWLzDirfG
QdLITnXu/g/1XXMgoBU5ebAkme0bWY+1mK0vT8jAZqiYTIKZfa60kOtkc+Sc0QQQ
o6wkPvaNqNrpNpOlUiae2n5DW1R1ONav+sz0w7yTA3G25/s+S/WPRboYJEVNgNko
T9LR1wn2AtBPYLiUS8kkPvpNGLG+CqK2aISiBcRMYu38K1YFbF/qFh2Fp4MmWyr+
XO4rL1Ss6IYmaHD3K+9sGcTxJpwpiu773QEQnUGaoDoOPWWbOGSp6lsqmhgXiMIa
ZGZig1kb1TxG8s1CWHil/hbQYOQWDhPheFtyrxhvUqRpX7w1MrGUra50VhVfKXf7
De8joXz3DZUzR9sz+XSR2UU7Cs+kNf32e5+girnw4W/0e8jdjk0FGQT33RQqiuxH
XO6OB0lRl2CpF1/Pb2TSufu7jtX7tTXesSzdbmgMRfA6Zbkfy/6w8+BdaC+CiGk3
Bl5BJ0/pBAz74nMvLptXglF00Tc9crJ4b8xXjjmWDff1MIkItye/lxbR6IrOX2PW
En8+/QMZfscEoLukbLBiS9ywdFR17gvkHis/xzzA3eaQeg9j0gpUYk8oWGJbdZ9A
+VXFBLLx/sjNXO7ucRwW60B68sdW5NiQ5DyD+zDiZKZ/X4XVscBxonQc3AKvFwcF
6FCAHxtwms+swwpq/1QKVAPsR1zADl3Cy+daLa34B+6sjNPf/mPsoDBK/k/ORdXF
/mKmmJyU+r1LWibLfEPKbFkDT0fGz82KQatwP1DMAUpoRaVh7pR4sbj1mI8CANMo
kL5AxwTPoBwvUdUIbHus0wShkjuF7hpvmYQ7+/n6BQ7Mv5DM4r1JoJj0W/eRIQVc
vPtlQu6701/dga5aXV7+ZPnd86kbrgGXerKF6mAjWqaFZsobdH47wbwYYU/gv2qa
cz95v3JpprUEstlQUJk53fEXOSKOcOHMtWbRMp/vARsDEvYot5EkzHyNWJPQCLM+
Opu1Z/Qkdh8oNilAkVXZCLLBQ5DkgSzZz83mrLdO05Rg9KJIMBDeOZvPxEMKsWo+
u37aR6sdEQBarxyJ6MVyxjwcGaK59iwSBo9OAu9tdIcsxIi9IulIZJ36gPDHp3c5
VyqHVxUQJQjSs7I4m6jNLu2P5MFinqsJiy2WsVqjotdlj/AANwgmLD8dETUjeksh
mZBZTA3gxOt2hkAV7Wep+xELBbg7OdjtbuBYSno7NU/JhPDC9lAOsYZYBmoHVMPZ
eICZSGOhEAk3FOGDykYY6+P6Rbd30E98CY27pGP9Vn/Yhd1GhmP5JrPRpbZVyMH3
SfKr/UYSLufGtwz/Z6DHo4upk8Q4qjQB9E/mqC/Leru7AqZ1lGd9PcTJuvsVVem6
22V0a+XR2+hMyY2FF1F0jxacF/qKTbZPipfnSsIxfhVw9jzRYnaocak15nDNxuvc
rNbfp53dnVYoyC4IR7bxN01MrkTiwTg6Fti9F52JhcfAxlZVRMt2a9yH6G4BlG6H
6L0+BvSvgEaMQHcb0Ucvkxho+qyxbJwmN9mWql/D0kprYiau60b53KKLu8kX6PMd
ZXbcC6oGnYmaMdWEakBj9e2mF56/Cth+qAQgDj+jKPqu9VBMpPIAr8FvSjiLuSaN
JQMTljJXzOVfpDoVFQBEfvEv5N9AMT19SeHXzQwfqMzUNGh7kBTeHyLkTYDqcN4x
i81dWyawWUi54Gtd4nhlCniuBSi6TlRx33QKZqfH/caRCOvGuIP3wzPbndr0lA73
Vcs5+nIaBq2S7OxGUUNw4KrTrcPIENzXg1DYJ8ffOQlZHR3UiFZWwiuZjn/CZvSb
3KGfKVPSueX9UOW5NQr+RJOgMsiJ7ENCPTu3KFubSX+8ncoJ1tUV+srUqcg3Jx75
GCEZToHaEmUuFN5P39fhZ0xe8jUnHshhSvJBih4a5j+8SQItXKuzgc+H9B8ngnJO
scejSXLdp9Fo8GIJ6hhkxmdEnx8Ux4WVK3aW7O1FFU22VWl5HS+rsQZIZD9YOxZu
A9ZPVMvfDT83BUnMJM7X/vmRfqfhC4mYNwGex7GBObntm5t6Z1/3MJLNTRo0rWO+
7jgbdJyZnXKzHzSaITQscn4Zmua83JowzSJtNR9TM5/CCQoourC4476MhrzzAHdc
xkWuFMUoRyZ2cluvlMihyzZgLYCTKXHfaKHkzU+Ia4Yc3vL2w1SxKRwhtj9OOaKU
UQQXpUvBzd+qlEzl+Bh0dcbn+AIW0Vmy+cVEMTPi/sH6ddwhINX10chFkT6EwoLM
o5hwoPs7kZdkJArk/mS3QM3KEvCLSFV1qLpq1tqWcSh7yGb5+Sso+7GGTpvJBIGP
BqKKb3cS9C/7J3TQ/Y0aQI/wH66q/pETUQ6m2HL2T+jdRXWuzT6TAUPkG5Rw4b8K
Qi1iDh2vi5UYqZ2Vk2ejIGOyYIoakyltPqSjH5dBqOElo7fZMojsMKOEd73H+NoM
JpMY3n/J/bi4IZ+9AH5bPXaIqC94ZngVW2KXFgfXLLU5dNfcc+XF5z22/jCOpmpr
vV8cLWO2PaqKOARP13DpGbyMAU4GRu++6nWrTWPJz5deXAfUPgCoMxo2PM1SE8ek
q7dwPG3YK7b0e0mpO8KSxYjCuPi4+V0MfNLU9HiAPFitgqcu9CmK5ZajYzPVSHg7
+tH2/5jvQ2OboCJHhx/Y24zHUawEyFcTCcn2D05cBpBLfbxcR01Q2NYQlX8Qhk7S
QQrNMbJdY5TiPkfj3kefwK56B0X4xbupBMe4ZpSCQkGf2X0iYw6MYNxHKamzwDMQ
PKVU5FpYXozP3Wwzi/KECsDYIMJsUS4y96vzckThxeWTYrqVbRfuwhfPr7cIGix1
hBLWSuEQeW1PcrtLGPZsYZ0wHNSL0Kp0U5oSMyakhstYJF39k/BNNtynrTiWsGgp
GYvY1dKhKm6lAPSM/e38KdWo/pDw9pC2RrCmD2sI15ew3CB/AM6e34fBKUEWEMLL
y4JsX2vaWkmeeGrGC2UX60lpDF5GoK2HfPlJlUMbPtwbi8BPJOZ+3TyPBMloUNKG
Vmvr0VOrTfFVGq6f3JGkM/XdRLAxC3uf9oAAK4tRP77zAFtXJzdz1EvKp4Odiqqj
zf4vbZLjaP36J3suqvKsiJzPzq6Su7sinb4K4XqrSHuntGz9wHEiMv+MIFp9WoNL
Dn6G8EnjTmERSxJgX5deJ1BhITvueWdU6uZBN6wzDcLXKR7FsuSFmnW37v22BkYp
WUu/OAO7h9naJXBa/9g2B7B52KQT4Z9B5iaScRHBUSezO4SM3xITQSzj5O9jrMPM
cUHRjQdDOHyJrvYqsJ2+orgynBAScuGSLq87NO6OImSLSJbQfHVavp8yEdMK2hCy
lGBjZmge66daGKN4+f0GMMuC/hWFEEknm4EPPnbFKOght8X6f2CURP7dJ1PtIrpD
C9X71jbomFInWUnTin98fXT+vWq5qxDpInlYhXCP0W2oW8hgL3ekSR2IiN3f2hhr
yDVPj1XzPr1duB79kiAFBCNUwnSlgSbWK6/2V4+pcNHqr5TxJhJMpk9hygVSmAwN
SqnWh8Key4glaGJj4yCOC5W6vE5OmoS8zneWh3pHuV+k7i3RTLEUmR+I1OU7pBd8
VD8gr0rgrlr7fN54ALGJQs1bXTk61sgMtuH6SGWiTpwPgS3bNn7/HhGXtZ3BTVdY
Vt3W2JA7vBd3jRHQ7xAq8J3Qyy5AbyRhiQ40QbS11R2OLVGrQp0108mw16lwk5Ie
77VluDpqIUbjiuYiM//m0NG4naYeqCF7tPfNA5h2a79Mi3FoM5gK/nHmhdD9GHXi
YvRCjXcPufqNPgzKlegt4h9HEI5xd4+3JiVv59t9y0kKyAiNWKz9lPyD0VG8c/kg
KEXOOJ46Azj1r0RTYLhiwHC6yHYUK4TZALSoTRDRCyRKU8dt3VyHg74TCbksZ2fL
lnizAjd1a3sUYqgIpnD9flcTqzvw/XWU5SMxXms7a1eSXYFxWjxgBFtv3zjboAs5
XegQLcrx/WvA5nSS+Z0D97E/fOPM5hRkfTn38acYpaWTCjZCXK0FCOQKYqiXVqUs
2xUNm3b9RtR7XrYUmFfRVXFH7hs+9oyqCFtVN8Ml1XpOgPqxLknJmgN7NYqfh7fG
nUt0UkClo9TOysRmMAQe/vlmZ1VMQsz/7RVecU0q1gY3YS/pWJxVUxY6eHHVG+YM
XTCY+infV9nI+DB6QR6J7g2DOEr44dZWewWUlSWCt+MOcM9EMnOkOhELvbgd7jBh
K+40F6Ty3aWsE90s9+KMl9105rrAne7bvrPHn0XJ6ZDqsrwFgge1Y6gK9uXQT1Y/
hCVCt66qcGEwWXvGuLt+ayLZ6z78x8YhWqNAZRYIA2XFeEAv4CoQzPJB6SeN7BDI
sKWxLy8N43Pluqkeg3iPFcRtnfw4smNFjaZcTuWrUq0RPRxdsq6nFEaiqCrNvEwF
QxWIWIvsAPc1ryztyyElqEiUn7RpdtAga8suHgGNJtejf/mIM1DeqWn+Aveur+++
0IQps7ABNaS13As64a3vGsI8smk7kaxfIDk5nkXfNUox4SsNNFe/ntnvF41t6BSA
EGcxEFEMl75ejrDfmU1EQ97Ug25zJM7DM8hEes9f5bBKj1u+bzqavRQ5MP7RSFAv
f4C++nZrUD6KhoOJusUH23nngGAFwkkSU4FL4wFx9j7FrchLdztcMiAsOjp3qJEv
v5pEpVBejhg8ADWXBtNcxFZjrP1FB6/QK3wx7EMJyuz9ka/cNT59WU7Up1B0e8/f
BAkJU+fA5okwhiriiK9KXv0U9MOJVOo5QD98tFRc4rPugdyETbe20EuWz1yqPz1i
KYWUQada7hpNI6l2FL/dhfXotrOufhm6y8N8tdTYNidiaPLuMeBddyTNvs17PMWf
CrxPQQOb3IljcBHlDXP2YI+6alKdmPDoRYLXFk8HtI8sgCWbl5Ll35Cc3mY4ja1/
aRrNJrkHLtRjNgYVT8BRIXxV95Fy5nq3R+xXyvPPvlcjjjMnVDXpYsCYDTXxhV6j
Yb3EBI+8k8Ap/+sQQtu73cu+70nePVdqQetgZqSkihJa8HFG9xHm8aDilbYhEs5E
0WRkIV80e1L2AHSn6e05X1nMwijhNwcob0Dv8l5HCvmj3oGpKOX+OCtgG/HPl5n7
55ggcq/2/6uVCRWJVeDjng+K0llwME0X66ohNKrNPYjIbCiVAER8+9v6wx4907eS
vSLzRbUvets0+vSReyN7Of4qNRpERXo/Ha2xgm9z1Q1HLJ2L7D3yBFYxR//obhhv
xPokNscTdAZfkB6heB2YFHuoX8O0XDR0LV4EuEsTKMu0OOT2SQxWelEDDNGd0ODX
uPhYZxA3lgFy3f5SACEK+R8XpHrzVcYUrRhZ7/7xrGkvvY3lc+Ky7cPmvQ1/WszK
SYf2zt+b+yRvrS0+pkoURzNSk/A7OmiviIdDhRrM6HIgv+hsSvjZeGCpb8boAMzN
fmkR25GIFTVxGyo9uuCLTgqO7T//ogPjldSC3YlOwxikeZQ9+fok4sEWShl7D8fC
iediY3L6Ol0t9axjxsMAq5v9djoa6yXjIAykHAcitYIhUnfbi4RrhWaZJfCEIsN5
1l9MjPy9Ho338xj005zFMpEATsxSpzSbLwamZ4MnaECHvoiOTmkO/KrZPzAto9MU
7t6ZrdnM/VKgruXqTl49A1m+7Hi+4XTuVdP7hwwAVE5UbfkF2ojrDLf3Wwu3VSMc
TyCMuFqvWYZKz6oft5No05VFpRk8iXy31L2YU4Ts37C93PfvFvi6yYkwGydCrB2z
LN8FBQw89Ix5y4DpdQKI2Ek3Ye2rgLSD99o4RkcUiNV/Rr8TYcjJYV19blvqIInV
56qbddK8PuxewlRbynhhhqksWRD9v1pBvX9AMjkwQI2vNJVKXKyDPQ/eZqHBqotO
Fhrl0sGy/zAngoNwFUKicGKgkib3bnayChPImadKb03LzNge5VpDeYx8brHaG3wT
kUSKoQkMgAEGIwqwspiv1dJeIcgVuCINdUYu0BP7w2HclcnrGYcy/edNhZ6co/bW
Vo+dxaGKuxigMIZN8zUWorIWkY9LZUrTrumFqtgaSg/353OUWejX+CTyrosT+y66
NYe9F5njsLaK/cMtR9LYkujHgWQFfrOq0+v0yeVu7WmH1/lIs2lR6a3yqn2/sglQ
Talx5fRcpOT17sgIH7Jz8U/DUn1WY479WDSGJ2qq6SDgNu0Yur0m8LXuXqWthWfj
f7vv2q1xqA1ESZw67EHWPvxSHsD0xiyPEWLLGyWosMDjpEmq8vxhMLET068xY6XQ
56b6s28KYM0wZkjxWO3FsRErTr/ChcCJdQTQseT6eiQMalHB6sj2qNLBcGjc3O2g
zLbZ87eXBQvE6/XNYnsLYFQvpQcGiUR7ewXEOZQigCQelFyCZmFb4W0UNsnPwtos
pX4n+JDcEVS5u7tog1ddRq0xzy4YfTmcziGx4wj4c/SQM9qA9M7ZyHwZnWxkf0a/
h84ryhzKTWkHkHMninyyiBqWN94DpZhreE5HUr10H5lkWP1XqXCgn0lzZTb3nGjt
ejh8xO+UcwtoltkP5/gO9ttZhaMQtkcJckbICuDwN59zGs/S8WKzFZ9ovJblYjrP
4I8/ZE7FGR8ToGg+873yv9FhFGGXS1bgIz3UiF1J+9HTC2k2sQnaXE9qbVj5Vj98
UPcm/EuuEypfXF8kxEOKsgoDqu/gT2eURjN4RguRl7GgJbZJL9InB34md8ygjcl7
S0gZeiEkVq7aAd4M6Zd+WBCaPkGoUXaRwMstG5BEygEEKKBVc75E5qGhtSh9dMrM
1JT6dNa3WnU9qjTducZACmuTdAwhx+mFxcm0FouqXZNOyCM6rCYe1Gqwsn9FCL7x
kfuGM4yJ85LYQJ4EPm4c8/pGBqpWDhfulQWlkhzp+AfYRa/ABRlFenkLcQbcGfSG
sJwVFk/dtdilNkezErcBZJwpD20FS3Yh9hV6C29xOWpy1KufQSeZfSDxBPp7MS+T
2xf7iLrypI5lhCoV7zIsNKofdPBBW3WCHukP92qbtRDta1y8028PwZVC0ksafBlx
EwRzVS6PvvyEiDPMlJiAVDB1sqeVmp39zf5+bi/M6i32/+yPq1CeYVATKIeORlhF
QJkvuvtjzgDcBJM8gZYOeYtHQckN5rhJWnd40o6pZ5T7qibNY9fgcGMRT/QcWJ7S
kH/aFqlXEqi8VzqDyUBVWDdsGJ6KtVgkOwsJyB5BHOqF4+4GSaUfB1SY1F/ylbEu
6uhCFgWiwgA74TDZOB5dWGd08DBWvvz5NdiEmF+IYY1VGkuqD9UfnICKjPqA/G8a
zIkCM4I+oOOfl6jWGTmhWf1N3tf8vTdFBdarFz4KzZKW2z60ZbR1xmYqC/jdDKgT
QmUZXciatYvzGKTicidopFZBMV0ETKhwiPXeyZ4wRk9SFKEtdNKAAO47ii0xT95R
ppqYSyAFA7EFSr9b//3uM/aqKFbeF4yniA4EtP5BqjbyFid4zjCjKbapwyypbHno
EbpT6En7PWaxBZgSpsHMPcIzL1VSZzUBudGT1E5SlBuecQ2GzynIp2x327bUpRVo
n7VW7mDjvm4wL1EFjIoOyeFnkZ3lBr+2v6E4YAE60CuteVmuyhuwKWe4ClNp3AQ+
ECmvxc0I4OBnmcORdk2pJTRErPJvNwwZqJOj6zbUwCESFBE7LxF0lbAfq7r+HaaR
jypJo626yf82onqft6gFMcn4CZfL9Z6PDxRjV2xzX8Rtf6TylZC5D4HCzjKqumQj
JxGaIjy+wfrwO4LlnwpCHZCu6+77xJt1HJDG6MA7uig3RzkvJYX/dVD6lUfMpkuD
B+gMAtWVDlfpsJ8rA1RceM+ISCedomzYP9yYtAFeHgn+vDz8SKV9jZvkQ/I4Tm0l
H1lmzgC2rpIwNfVouMsVz1YF9sxHSOwHDlj1zAFEQrfvzm4hnBPYPh9iQdE9KZr7
dAq3nruTh40Dxb4xD5Vt3lSUdS59eeG2gKIA9N5+ctohRxrQUyMsUdKSaVg2d5ab
nwIk9nExIKir1j5Dy6Bvo4edETNmd1Y6Unt5X0DVMtzw43o7yc8WQKDL3YAH0EN8
`protect END_PROTECTED
