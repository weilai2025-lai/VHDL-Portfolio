`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljWBhWMpUL5Rd8C3AGo+flhYFRnAZFC6X2qbXA70uG6P8Z/ve1STnf1mz6PDXRJc
/ljuntQ1mcHMZF1oNG80uom3g4wvERAIqPZN7sqq91nfBYhSTYH+Xzg3PS+7SSy5
tNIL3LIS3HJ4OpxeZ5IpX7zxDJ3eBAh4G60GuyAM1lApuGMdKQw6uG169aX8clK5
2pTnn9MPD+Q+ifnX7zK6KKTKbawJzqv4XkZK4EracvSfKlUjO60tIdWnLNFtvx8o
mQ9jDCXOjtAQKDZqxQzZgaW39ypcB/50hGnrSQGXHN8DneOrDyimEQR45S9rbtUe
ljyqDwbStT06geD1xvC1Ud3vt77r4ijVJd6gqSRF8rLOnFKzJCE8+bf+s/KAoGai
mJzT8BQZ0SmwLRqTAqIJ6bxBMGT44Tx2iqHzPC/61XQAU3GQ5RZ0GAvxDd013Hkv
V7aHeu6pEFTmIfO6CFMZG1wJi/kielTkrDC4za+gsMb1puoti2eqgexhjMiXcwur
0mLSs715YRF+RGCCBdcR3cQxAwzjh8S5OcDpWu3bfXp2+kY4UoUpZhCWRLelKx3c
4vKFGprkQuJLcnOJAzwYPor5wB6zjvWpujD58B9krrYRZ6cHVg99q66/SCRu1gUg
9zmxzr2Ytjp3WiMCKWKBCaldICE9n6ZfX2evcQJBwDnX+nsbADpvcFu74wFfXJhA
31L+jnh7UD55go3JLh3CIl2bbFNRIBmUgXOzhZyiaiwddrP6Fc9KGUzWhw/W2yPn
ZPhMkcsmucNsor8U7Is89+bAoP3wpkHZ3STPb0jEKll67fhPZcd4QW81WuZlNSbU
bpm2GYQ8v2CmLrMAtZmx43jxFvVA7FeVYB78CWzuyaaK4PiaLc20gAUVYHhlHIjY
ZUyddB4vRvQCPQU86z/sHeAkh/svQ3tOKPmWn75fEnzkWWgXFSEexG8oxWxk4vu8
Fwu6Y/q0rphahpS2CEcVv3OYeXNnIHRNMCvHAPqT2CQTUPSX7X3uKiHuXtnskQ9F
J+r4lZm476QP6+svh7qPHTTELcu9w3Zhf4yWs/XiacrhnoJq0EOJyg+n3M+Sxvhy
kYHUbc4p0Up5vxgkBaWRgOo4lVV8eDss5i76XfHIVrwvQUJzyFi/NFXJZ8h3m0lY
h7H9JfUuHTwJjb/nAHM9S+kjeUiqLscGt7TVevm+SfCavSuQJfNNF2HwAbNYrEtA
J/ZCKz+s1jZFaGw8Wy1kSTo8HfF4emY92gqIcyKtIzkgkfwKZpm7ALq0fxBOUTK0
R2d6NALmEsWa74SDB4miq1L6qvllnvV9k3ig7fB5abpMzSeWO4VuirN2HqkbFvz0
XBdlL3VinU4P2xmM+fUEJL9cdn36ltpgDr6WzJakoMb5+xE/uxR4YLbqCFZDeNOe
TKR/94O18nluTxkWWL1Lh4RNf50TYyAYg2xo6zyGIEJgeQ0g5qMEQGkXNOqQR2zV
ZW4Kyv9yScoTc+4QemdhKUMzlVeI92J5/Gv3r1WEHmI56th9InGMT0f9YnujZMAB
ae4XuGCA3CDA05tRbooIsv40dbmnvWC2RrRcz3p04/3oYYRpTBhiITWTCykm53vC
1/7J5MNSUlGwwSS+ywqKh12w69CLyfkR3zF0k/eK7gJM8qqTk12eLWAhVPvwWyMH
TEE6aBKvC4y1XKs1TEy1I/SQKcrTpskT8236xoo00OKS9S+HDhv1+UFKQbWqVskl
yi+PEU4UmISiKvtfNwPZGFs4GGSQ3T526w0B4v61OzFeOIrYuwKDACrD/Tvw0ASV
C8xupzzdG/NaneBihBiFgmq6wRWmCC/I90FjT3L0ddUYzwEKhRqKHiKA12J6KHPK
+/z4cQgkblq4E/3/Db/wDRuQdBeBngn8IFRfGa830QZ57CvlrW4Odb8rxUljy/h2
MHczYWHekZRiEqFR6suoq3ZvsxmIrcVfd+FhRPg0ZbI74JdX9Xa9DMPM7r6oKrfj
NoBjQ2jwxK53dWOgZsPqw5yVzLpgmyPkOg/uF4Rrb0cmsrBUdcbYUXHkvSVESHbJ
0n3oaX8UgikjHwyeJ6/FfTJWJE++BNa6cXFAZw+Pz9U1ZazqwVFa6jiAFc/sVbJ6
e22keDAvK4inwO7424xji+7TXfl3nQ/B+X+/FCUCaUQ/DsakQmvr4CET0QDqWZzu
K0lSmu5ElGj4vabMy5RTftz18ClWRpwBYjt+FXHJWV79KGK/Rxjlp0qNhFNIQefU
LYKO8FcdnYC9rH6WMvap9J/IGIvcOWIeh80W00tXLB2Z3dlsuHuWGfPcxyuGfxSN
r8DmjcAiW2gndHc92mqxDf4K1X9ybUqzqi8no7mBVBXsHwMLrcDFi+rqHLCqxQI1
jF2cGIpj+eQUYpjhjJZQ9ejPo7uqzGXR5096i87mjo/ygCOgYqRaBevy0kz+3Za9
ZuJ5UldQgxCsEdnJq+NYOj+VbqjRURiZvD0AfFMUU17oxnCB1cGQN+z1rfXPk73l
or5EXwZvc7ZNLwdYOvDD7et3hThvh1O2+y5pERDwpe0nzAOpcGdlxVC33PiH4Z2l
N04RSQjyup8cqw4a4kjzYmhnP+F7j8Clu/6xtAt7JXvyod4ucdRj8AS416YzgqZo
afP5mEOFpmifJ+JpW2ioM93VbeeRC19XNzGGHlS+7fu+dcW4oOAvSQii0szwEQuW
kbVXTy4YIeFjGZGoP9DAy4869vGR+Dc0eMOs2oLd7XBewrsVQI9oZyhFsuXlqmeK
UujhGkv7V7AyCBOG8kEz+POX9Tw0u8l8LhkinJ438jsCQJw5egde4ZWc48utYeLZ
qoBsOgJdJ4IH/Fs/IdWx942/LFA/DphXM9OITmX+VMWUB7CFwGZsPmG5SKR6STld
PupNOsVGvCGHNtP4JnX2gmmI08HtqrG3fz3xswOr+qOvW4+PSCBSCziG/cFkfwum
tBGmNVrlA7BgWfaqbfoOajWAsTGebksyPOZ2+CB4C5PdoXiyOA/dt1xge0BLx2gW
C6YGABpFL9p8JS2br5W+OgP0C2QyqnCEcdUswbT0X89tiXH87PAoGikuKH2AW+hL
tpY08ZFmFG8qUndmmUxxj9qJH95EcMpHO31Co564gHGbtPDV4j0kv3WWiKclHGX7
rzXRqnEUQxGE1R3R0swqBUF3ln0jml++a3Zf38C4xSVkd20Kg5XpS57qookYjnum
Y2Ye0a5D5AwqGmsygPoN3WiuK/sbDNMySoiPfi5KsfPvMWcn1pNUBOMCmjF3Ttwt
1dVEgcQN8VJ6v5rVogKeud+uxrx1zbSY8iMluHocchq0tWt0NQuzl+rjUAngfoop
nZghG1fo/rKsglnRO0P37BGS9ouHXZ5X4s6oxanmJe30LuGub/fmB9iUfIaTIICo
mrWT6yxkjQR9FHF9i4IkyuhWALM/YMcHHnl5cwbTEhfd60na24RwUJzBiHXR2Fm7
1ZhF0gcq8u/7SB3ihz0AxMsLq6wZrxdWnZyqE1RPy8K7bsMZqFnvsu7r4RZaAkA6
rsam/VaU7PiX9sipzZ1m8vlrBBR4TvxlfPieF+XpZIU6TwfGOc+0BDiNcLoh2cO6
K6x69dVWHQOdOWLzwq4HixkDllAUSa7b7Xy/okrjrBD2ZKfQv0zCkagJqS42DfTE
lpa6Q/oJkiIO6iOFKdP3/I4ZTFRu9p13xyIQgXCjsdQJidrhRJKU9bU40fgdyfzZ
8RH1sD3DU/DohMNEm2JvFlZJHV1i5XMcPqHC/Qj5VyJGB3fXdk0kyTwVvlD7E0ZZ
WdQsUtp5v/qoP8fnLf71Dt6N2gQGs8NgVDRJYi0QNV2lOsBF29uVFwW3XpQJU1Xv
Q3IQuWoBWw91z9bd6/kZGCzx8zHyol9WBRX+cGFFQda5sPaUMrmy4xdKPJCsQYOw
N/QEQgZVpZJej09UMbPpZ9cZujWQwow5PT7bKsA852THMaoAMUZBxHcAZssCV/UP
`protect END_PROTECTED
