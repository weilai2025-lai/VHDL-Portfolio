`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAyo5rUOHeKI3C6/w6ekbmU4oiLQHB3ufdMRmA4uMUgjOImTfvbyZzdTT/80irKO
8ZmrCX3C+orFlOZA0ybXZZ2PXWBe8qFZetEVM3Cwg0Jdtmsv8WnwajxhlVjsBaud
I3ZSioh1vrSut9JXb3ESxD7xLavQ3cdOjFjMd3vaFlgs4djkYvUrsJjpgtCLWK7X
kptEO9Cm5Wj6cmtKT72FVibMAVsdK4FAcYQ5IzrYW0U10bxwIiewocU2w/ObXg20
pH8IuG6dCtI0kTJo4koS1GxLigPZKk/xKe1X+ZAkgEhbzoQSryAmHLHgCijXbEbS
/4+y12Kdsn9ymJOYB0CGwHaMT6+oh4cMrxTSmxNYjzF5ThqtPfw3Hbitn8aL79Ek
5Y5JTaUM6x7sX0KN2EoYsDAhPSSeyZTNgiVTEtjbTu5eiNKSt68P0qkJh4vn8y8D
UGoASne7BcY0Qk0L8uTd9yUKJ8MISGb+vNtbc282eU2XrXUSZERBD3utrlBHzr1r
KQmrYVgTKndknlpftqm21QcTLwNTaebcNqDMrGdZfApJ8SYdH/G5MBSTDjRwoBaO
5iTouhJizsKzQhn9eASzSGMspYcqdbZLmfIBfg3nxp2kMl/hZ2SddbWX42CiMRwu
83VKIcOqWDIMtloEWY0SJJoL68xJ+T73Z1c5j3FCxvfjpJDSrjWpphhS74j9pQvn
vGcRCpZkFqU5GEOVJSEMMO+KxpoWXXJ1AvSq8MOLPkOtK9sCBba9DmjMMFS/qDaQ
AtUpd0Fl2kqL92zUiiTFC1QeC1lZWphBuXJDbvOXBRR0+bnTWxkJqIOeCc53Lja1
zkR6vdevCY9SrQ7OUm2HdAuTT587NGXcugEbtLRsjMLR29j6H54SQwK0LVl/nAC6
fJGn/gfDWdlrLrfJ2cO7p3oahlciSLNTg0D2xMhbPiTdeq4hSxX5lIsPfuzT1NO3
aay1blXUDl5wSWCDsheWkmGoUKxR4RmNNtsEgZLAsyUtiGIransT+E8Wckub30Mc
cAS38GhopyUjkLK5xXpsdvrjOWcJiCnxJl669ISxY9qnyLhO5cCefg5zpoYF8n9l
ZhzeVoLF7AMqj0Cf+PlVBFRIzx/LMn5I5Ykg9sxoIoxQwKEJA9G4o5SSHpMPwoug
FsBWDHCfx8ZALVKqeSPe0PSO2dCN5BAuktUg7W83qW06sxbEY/GtwR3KPzghP8UD
Xs1CtPNyhedEd4EcEbzaq8YPhy34B9FfyL+E+ccDsS0BDSvz1b7dxkUhGq1Rb44z
Uak9bh2cJReNHv/saPiKyf5eZKFULd1KYloew4w2wLxafpgfHgzt8PIsZJsItBiO
reHMUCIdbJiomUsgBl2joMXD9f7sy8S9tIm10gckmGM=
`protect END_PROTECTED
