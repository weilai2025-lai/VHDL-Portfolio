`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4STEDeukNd/vLjpO5wwePPhMdhg+NwMQGh5Wt8xU+b0EmRhzs2o2zauPh1FoEbZW
k9zAiZB0zrjGk5NIUBtO9yVVbK55Llyg/7TZOu5E89pd6twaEecTTaKojR220ZqF
JWwOuQqWlwvRMsFRz6siJarkJRc5CqjPsmUHlmkE6N1tgT8uqXR1jxJ90HlDtoId
WosvoV2jnji+AW2E7yTtukOqrK3a6HOy9ZEjecoAo9KcBNs6p4QLUCzkPc6P3MqX
jSuWHkILFIKsDFoYlIIuo/w235T9Gg7Nemx3LveWBhpDCkdm3EqAA2Vy3+tEQIma
77O9IPLES2WhPycizBsifZ1ptg5g9eDkxjuDh9Ofoe3882/2H0zcqa/4sxksjgmU
IfvXGmXREAvNiC4alx8U41qwKlY5PJ+EmM33sZgYchN6UEfWXnSQGuIpUNquY3bw
Y8NaQArSY/A3vqaxLmN6vnx1iuZDYLMQrdcooMY6e/3jqS+H4XnIPs4mjFsAerZM
XlGo8pqBii+sJ04E/7r7bR6Inc7ZuMMBzBTaRUPGCX38SGVAtdWtge9b2yIGGX7J
SSFkMANO+1KnyFk8yRid6prHYVIU8ccCRqCS5MSTrZLEloe0rqFIVD1pdNdBl6BZ
D8pJUxiE730T3eWAcP5FqyMkTXQNpirBDd5bO1dE8Hn4GyxAa4k3EbopLT6uE23w
G2p0V2vvmGHIWUTva7JTtdElr5U5leUaNUgFQiZsGOljUuF2ay33nF65XHAMhwaQ
r7S6PN4u3Wj1SMgqW5qaQQTy4r3Qh5XXUs1MvEB+Ft+fIAjqlbBWBulnCtPa0Xsr
mc8kzZSfr/4712RCN2R5gQc7M2ibZcEzriCSTH4cz2Av7AMUx7MgEok0OFWlwxKe
xAOOZDMvwuWP4u/m/TubONahit364N+7YOvb/J2EeFzF3rFIC/NqLf4CSP0I26Gk
r/7mnt6nv0aUJi+JpFjFkbn6IbjX+xjmqvdDUM1O70HbFZiqQv+TU1EKjg6eaBke
WdE0ao03Ga4bKZID0BhzpPVRYaIbUNqS6/sjtngpiFpfh2dooXdXS4XhDmQL2213
kC1nMWkTZ0NUVdoWQgOlj03UoZZS2xMfvEyZRYHqV62gt0hHxrSTFVWsG+GXQE0U
7VGhd1kLuSm0OH+aFtat/Hm7FP5AIok1z+7HUI2dynboZaG7gKHokG7JGyjQSs8l
9Lr6a7/wf3RtLiogdhQNxBQ5YlHrbJsojJ7JoV4Sfx+UgJOkp+sjzRZA7IlR+vvk
2V+J72gRfO9LJsEPGIaJTZInYlNgKg2IAxzwFBfKZB/U5iG1eMaNyEHNbEFx0x1U
K0A1EwaDD7R03bmN4nknjvcSCcyWzRW10xo9U8m4heiFQBjnh42yA3TiEBxPGSBx
HOyDWg1f9A5l+WQmlBeQWoitacNzwJiFnC7fAbs5/vOR70spBg3pdVsj6qmbt6D8
hqDeeoe28kbIFVKS04ueaJqNf0YPpCYuzUJ5mxNQm6bXPRONWrPJG4c5vObgcYrS
3viFz/cAVMLl+1czGiksmdb8X+OlkuKIjTwhu5/Tp8L4G0t5RQkfWBgduObXXUfE
JzoxqlAsF/2vhwQ/9CpsaoyDRaNVqqPQ17rUyqTY8FKv+Pqzz3sXfjvYNJ55nNDJ
ad1ldoxETJqOs8omxKH9wKrXt/2bAFnirdLty0B5d+0+v/X0nfuFqVFunPfOZc4K
akHwIMHHU5z85xBjqkhfyukwcGSzZEWRFAZ1ofht6ehmMOh1xy+lpOkkp14gdj/Q
wMfovq3OM6glO99JGKoY331msxstjKDAqNpKfTVK0J0vimnoUwDnfjL41oWhG2DI
FRHaiAIReOQak+UtTLiYIT0t+hJI16SVdRHMDTB4/rfVckGHcfFaVrivBybimVEK
sYAL7ZPDh5yR7/yzYZoSyu31ywv4ZNa3bNE9hADkpmKuwl/Ijx60djyfKdTjiNce
gdLnOZNas7bGYctu9DuDJKBJNczksdfFWTdxXieqsdju/cVNHM1nuOSQNIaAkPYa
A86rtgNa9FfkVN3+WVJYgwJiTH9vLAsX5uk+ZzLrZlqq4rLNccAX3UHYPh0H8rPn
jlGCchEwZLv5AObOg6YgZqXlWteeBgXiYglIfTecpKPS8vhFdhFKgyCIlsJbiXAw
vioDtW1BihsQzRIHGOtp8ebF+0f1xVcNrKLje+60mp3O92Bgvfnm87HzbqWzRKt1
7XyN887hu6ZDMDaYPyW4TmQtSfFyKejyWRBQW6DkgywH4hIZBokUWETgNevGcYih
NBRgeZK6y1o5f43lzV5QOe2OaV7uOekIYiSPWw18aM4LWq3FUDyDVZLbxLYH7Ggo
tepmAeDkyKY9SyWnuDhzqpL0b5EY8zhztvZAoyPRMJ1dAjTSDr+RAoJZBiL2h2Dg
hJOoRDSHslCu4lXwJE3dw3CiqNdjIe9Pq3LXRY6wyqRHqqHrJSkrWk/NCp8yB0pz
m/ZPpNennFQ7Vve+0e9QhhEzD3Ym9k1PrAAb9zdju805u4VtvijyKXWsgTV6AeS6
A4sGJ+s9tNK7JzLtQEQwwcMgSvIthZbcI8hiScU+6jZ3ves6ALd3kX/7yVV5JUUv
GxZ70+5WktvBvCd5Yy7Fi1WSu51GpnHmEJOwL14B2mOBLd4hkWhtDimprdusfXm1
fP/1ZbnEAfMMAc/+IqLpfKgxd1NSHTTDTydBTykRuN8YxL83LHzeDl+p7B23kMu2
6b3S+1dK6mi0DMnY2gzTQkMZe3PP437PsRge7/+K+HFdthmUKZWGUCZlTntgo1/A
GCEE2KsLhz8LvWbVYb4fc5IwIcrFu816XT/1KY4BxwlHxKokWrw8ZOOB4FC3PDM3
W7Dw3g+lkvdJoiRk8XKZW1qfawUUrNfZPfvxUC8QMoTaeZSVu2UwzyeUieH3Ub2a
/CsyS0Zg0aXlUVLSO/PclRIeiZpej7eEk27ljq4ydV+1YYqUnGa8qaA2qubuQUMn
VtwpnPPeABu0cQePUv818aVNDqzV20WamhF/lLux6/746tB62v/uRNzJDQuImzsa
ndEqs6jAnnA9x29+zIEZ4UC8oyz6kV3JIBfdreXg5I808YRoRNneRgGh81//bIiY
T4+M0KadAHxrh5fNJZ8TpDl56IYXY/C/Y4z44Bmw142EZCDnGmVgcO1/b0QbDU0J
uSxTxo8c0SIQMsH2+TYCiNf6K4otvZ0WxvmPFaEL9Lxu34Z3THjjCnbjkMqQKKic
SCz4mkAJHd8noqDgExhbBvqVuaoVe5RnbsHCI2hrXtYBrg+xucv+93bPGyd2AMyT
RDteIPRmgl5ZfNSw5M10YYdaOneU57hnJ0k1UFvu8VZ9JYii+AVTGzKD4nnSTkFE
Ao6plKKeTsDcxfBLO20ENwyu9uefFv5baMtdEQ/UrhxRR426h7NfrUZETY/EeGuP
xg8asdSLUmH8QJbdiS8iQMUBoKCQ+3jVD7V4WSYfhxzjvLvkmG4/FLb2W3PQH4eM
vwXV0r7yk4QDuysTPPzoVZTsYS/Ky3Pwn4na8FYDW6g6BDQJPXCncwvLw7AnYdtK
30lYgbhF0HTWyxrwESnVFuZkC0BY53vPkgZpCj3xqnvLmcId3P2ITD77fAFY+Evc
3Tmw4jYEkNgvSHT8v0RfzJHjNFpgf64ZGpCvJHYDTRP+W3KcWE7jQgw+NG/wydmO
WgiLByluPgQphr5TVQg0OXUepBhgwPmeZupIGmOpsri14vVdUFfimgAO2H5YZ+O/
wHChEsriMLPXpGWg4YsLBL2Xb8advHkbEiY6Ruo1hO4GhUcAsELOY5YtogkIJouS
zzqYR5BAbijEUdcOYX+dbXU7IHSHS1GaKDUJ3q7UiUszyhRRJSdHiaG8rnpQzVx5
XRvCyiu01o7wNG6OuqLV57FpppzhNNhRioBksI13Q9IlLdivxbayqgBf4hEENfAh
759YvFqqweyBDIJkhBisC2UCMZe0WQuhw9IyiG5ISJlqCfsh1GjoiXipSYHW7t0l
Fyvk5mUu9YdbgpupPouUA05AkZyRhrZ1/5eLX4wgWESIcUerukFUBojx2ofD86VQ
k9jL/rDXcxCUAlMHq4Onr2pF/975C7p3umxuHDalo7Ca6ZizQHuu+UJpB5gX0efE
KV1sz2EA2r44U89sbc6Y3DvjOJqsHsoEoPd3kJKKXUytdNrNJBPBptYquT/mVJq+
QyO3dxm3gZ7UqgnrdcCwVTPdaxz8siTfkMHwNnnWsAhOCLo179lLU7ooQ4aM0u4b
K4SF0KN/Vlum4wqjQU661ax+BInQB0tQ4c4FqXsgkrejIcNdZkJem116+X1qRG9O
emrbsvozDe5HI1+vGz3ZI7qD4Mp8nkh69G/ZJlC0ThdYV5zRPfAvlpSo8si9noUV
di2FMclItQSth5q1kHEuP1ufWpR5dk1lM2z/Rsq5XNnqgkHfxlNUrepM3nrescZ/
cakF7wqoals/KqyYW+PcLwTCm8q6FExiPO6SpIdi+5FreYcpRogp2hGL6AsSsgEf
vSCkVg90Zdvc5HBb/XW7Vz7wC30Uz1wNOhQHp64v20KEqZpPxrXbnsLhvyHk9Xd+
iXwrCoCfwBMC+2NoCztxNF6BfuxVwv9W6bUefisb84ka0zzPn7ePgwuHofHv9eKU
4Nnuyfpb5tvkdwsL07r/Q1QxoviCAJiT77otslzvY5r8oGgEpxssnTxWVImg6OPQ
4pTeN7fLVhVx92N0LosbqBSkTn4RQ0VfjqhnxByF3I1QORUczfbbKZ4D1GdGImaI
nddM7AxqPkt1pfetZ+kyfocIpiVK0RmIPJAyfp9Yb6/cape0QxtlZXXR/yQUwNUc
tl1fbujFyHFiClA1aXA6b46inbvMv6JGUs/+5GnfGNy4SiwjC4UT32rzFnNXwE8I
noWdk8T0aXGJ5aNoibJSnitptK4vk/C6oAiUc+cAw1htdnQ0tjkxRM8Pou7dlmOD
xUxd2mSsBb0ZYBrpJRO/94Ws8c3hED1cL24PgFDqN6P1pGAtGVq77abaB2fdOsDs
tvT002Fvn7li6NL1bbK2bP2ZsPnt/T2yWjAUWY9Pf7hzfrDzI/jR66cQ5f/cIjmF
/H7iGERa6Clb0jnHkX1a+idvy4B4zeVqNa+j1f2C/ANFkU8qKaZ/9bIMB7jZWllB
8x6NV+RoTI+hMBaPmQuHQRWhHechf0nr/uamiucqRXB17F3XTryIruoOJuFvS05R
DqZxMyWfdSxQCHxefRCSQ7uG+BiZ6o8OAXLYWmPDWF8LhU7AblZTt/nSIkAIDV2c
15h8fqj+ZYlPbu801UOVBX1q5tNeWpxKOu3tsjVc9EDO3WQewUuFJcy/Mz8cD+i7
v8QLuVJjdq/bp6QEQ7Wo9oJNIqQ0XAdtlCyw42AAKyUY6Ae2/+jVETm464Vf+CPv
KKLWGc1infRmRMRa3K72cYsGMVMNniPXsY6MbkB+JUH3XJ7pIZpgbMRaQ+FSK9ck
B+6jxkweEB1/p3jINSJk+Qw+sulKYYc3hFGXQM/8lLVBtmRE2fm+c4dZHsrrqmjz
P4VqYGRd1QMUpqr21UCZrk0hzppbFEczA9C0DBr8VoS2qnEiGjTzJ8LL3YQwRoVm
Ch+TPihKbyGOqiykCHMKrJ7rEGSJ4FYc3e7auF01meepaj9bf+EEOUN9uemIMNrx
8ddf5k/zpPBjDlYmLnRIyL7FyEohsPuHIyWW84OYCgY6820cZpVDgaQLtoKNDo1N
sY6Oo6yM7aTJ/zCyJeNDX1XwXGTJyYFNOrY1W7t3cUjRSzXXKzBXOptGGBuKgyX6
jcQViFvxaXozgFIVaeI25i1o8flGgYnedAd/EX8aD9Flsx5lEaSdAmNa36/LPEZo
ldfGtUvqRkGWa37wopWYEB7mgGbcNAZwlqQfzlff6uiFrvsazBXY5GBSxG6ssAGA
X/EJa/a/DidoxD4QCnADRLjQPmjQ3t4BleIuPV49a/NERtgN48MFLcI7A1UUjuMh
2yovQ+iGmlQabW68MnIhrI42CvenUCTnw0P0hug+Y0COWHr1j8tqtQRaucvQMwZg
H2j52XE/Ubu40nGCewW/7oQyeaD6D9VaARxJrpIeeXbT+ABc5ubER9eQvHuIcckG
X6bmHTz17+8t1NawS5AVHtT3n6v+KPSs6gT61B/mHfOzgIXwIZPBFdGtBAi0K7Bg
M7b4L/HUuxpWnlBui+ZOnS9fkYxMUi2KeG9XZNnfh4EjcChasiHGQQqjemRdfpDX
BW2D4IkU2kTV7Ja4GD/sX7nPyxftapLaUpVUYnjM9FnfLtM9f0+Wt+GrKpLdB/2A
oN+0YVTmWP7Jq74EzixH87rppOn8d1/17ezMNsT40ExC24M6mxGKmERjEZZel41G
7I2+a78qOyVrjUd8CxClnddCEEjWfurJPly1APJnUpKB85Bj3nlY323+cVWBRSEq
a+gAA/1Zmr8+tlTgfg1EZDY/B2y83potCLISjqfs5VVUOPTmkGIMqvRY0xfoVc6o
+U3DOIg4R95ATJZ9yKNKjy0njdNT8ocqLD3wO/Qa6YejdhgTMf2Pjp2Qs+eJ3qeR
F+6U/1oq+GnHAngyWttxnSEmHBa9pRahIMwIetwyi39ZYlpA4Kc2c/sVUnwO4ukg
kUtfwjV/8aitQlAfdHaEwDWUlFJst/8cK+0uKX55MMPmV+zufNeVMTfBidozVOpH
N3GDCAQF0GQtKPh3WzqN3P6SRz1MA96nDaePq4A/KmdE2KJSg5q+fn2gWdkbnI8G
qO/W8HObU0M1vnkm/oxWp9cM6YuAQ3ZMbpbn/4bT3jup5lf3UYAVbdWMBrJ8Z0TQ
dUxfIm2l0Kx15cUXmx2cY28bc9WISTLUFmoV6k6yUyv5kY5xZ0pSOdOfL+oMG+3+
KqixIL7J2cT7KjShKqkHGJolRrkuiHxnjFy7aHu+FdtACR7PyMAlwdvp06DQtq5m
SAEl3rW7wudmgml4TtnkU8xSlREIJMet4Ycqvm2wY7ebhvhDE4epVmMWgj9mNFfY
WgjcNzavxGM+1e8sGA0gVtS/X7d4HaLMx/l520nt1btmrB/hLT4/80XH5LTZeON6
qZRPSN4nJeU8jwEjL30MCRuSnXQw5UEE4niFWU/51UPTBjfdvdWrv3WThrvDBD/O
EiUY0kMz3vAsYer8II0nQZ+WgC0jmaVYZeDJVB2BydmTSEyjT3zP8eaDYXM4o7xO
77PP0Y3VvtFdNtKsG1Ajvye0DXVLkzEkBnPKxo6aXNKyWb3pFseTzE+QnlPT2mcO
FTnoUucflMe2amAVE+V2mhfcTlADIqGoXqKzUs9HnKCMJmQEmFYzQnlhzXMKq0ZX
xNlbit9xjHKfspT+DqYzKSBoXAEQ03a1z6AP6r72iVzmocgIEoUpEI3Vti8KlTXf
iRwRVSw2XWAEmwPZp+3OeeLxSQIJaN03Jc+72TMeNuUmzmMhH6ya64uHW5MOu4mP
ku4uo2QlH9HtNssTbV3go/df6jw9w+qD8WgaLZtER27bcO2RCKlu5raGX6vdxF/s
IQPjlfv0uOMhPBOzYYqVQ0zLFe8tMbTWRZx1BLXapa+60gTwxz81QkL39TPkWd3C
DGAjkBH2FlqA3K/h4IUpjmaVRBBMgrnS80mPiZqlXZVdQpXWlyTpeCS5cdI8QquG
7fxgZsN2WHvl3Vu0ImUIL//NNz2iXmHFhOJJEAH4oMxolwCOMBDyIBMtkC9HRoE2
4KEP+2c3qCG34vcqL2I581LIwBxC1simAZJui+msvI3EoH2dzAxZ5fvbhyJOxVN/
UkUlUZqqvphMMNQMLDmbZUSzbD6Bgy/He9hBztFuv7zqCwPGDNDCvpnfY/o6zCMy
c40cjSID8lK/wzvUZFy/Fqw3D4uyZi4DsKMe0tQiNYdH09Z135DbPV8r3u6vWnrT
7u3AirkmBjL96dDsFACBX6bOMmXR3TW87JlCm/0M8KsdNg2+G22BbhdQkI89DNAr
aHmaMEkRLA2/CLLMrIRP5oz2wU1N4NloWO7zcfgWJWRX5oeGXv3DaZo4k8865nnx
+OckYiZTW8V8JkEaoBHjrvRExpsEvMg0S+AEcxYBn7fBmNgcGWo9SMxhoYXG7lyO
hYvzAde6x9ozwVkyzRM6+Owx2oBpEQiOn+w8mDbz/vcir0/hvnwCI3nFbEwcjgGC
0v/RW4jtMAPNPOh1j2nvCgBhzJMMk2F65sLVdfsB0cra2VtSG5I9MHCoyVV5/dVS
kIOydumaYk9jJeva4MVjxlBZDPlUMYtmW26V65MZZKW3jxjjKHjU4PHNY7VcHNsv
CGGN1RT+TwEx+omDTp9vjZSJZFSzDD79Myidp+zDQ6O9Jlzt4CkDmNlKxzImx1UL
iy+/7KrQQZhevq2tuNUR8q11HtL9UjIEKW8bUwblpTP1Bsi0InLeTvFHaefyhTaM
iunlr34Fk+SExrqYqp+4gmHYXIkbxhZmNdH0a2oiRwRjHsEd8mOxFAi1ay/IVw1O
xJj8BUb16KBEALY+JDz0hvTozzIq6EKcLcTiv3eEbO6a4F7+Ufd10p+SemTyBeib
AWWiexRLWp6FzqLB67UfFXjCdXyL/CcHKH/8qq5FAYYTzMAiJRQhbKYAjj8btjtA
3f0AR4nAk7jqubyR/pjT5rcGuEwm+zYJ0xjM58Yn+UG3IrPfKt8N9t7kV32XOEhS
5rK9EeVuGBhFaw3G5yU3WycR2R6wDEAYURzmGkiOjPvb5hhiBBcRTN0qKrLT7xMd
daEqRsKQjxYdPS8cAh10i8vfl307g4xwOpyejeqIH0O4cgxd+EI8jHn7gzmZJ6Ea
bF3n8P870O0h85qyS4MZaLkO3dbT/B91ybCQzMds//nPMMjC311OlbM3v3cyr4cU
/c9u73HAdOGO4o9ByvQlEDPxdki5eUAYH+ZTVQrB8C52sM8u/JOx4QU9+c4h8WZK
v2gw2o6g+UM9gn0rkehA8UUd7yAXnuzeCmbeG4+bF3rK8pk0qnE0J7QNl1oBd4FZ
cl+rDls4Vp4P2UwxJqFjrEZtpfEQ5wVlnQQO7Gdcilt8GC2vLSnvSpryyKiNmyoz
0cQyHytjWySOf+6H6etyHPseTMDRUWpBzVaLKomRd87gzvbhwiaZzBsZVgFTog3n
I4hijHb3EPzCWXhong9tv7D4uiWMWxdduuAlLQ4ZFIk+A/3Y95AEiSwK/tZBEZCv
datyAvuU5YaVbO7ZND6C9LVNaKfz8Y+w66zEnD+QF+ejkikfBVPOjw26j0It0P2Z
34zPyZtkUDVZGjCz5wOqv/7/u3y2byqBJO0uaO43LkzGkPxGkJ98NeI/3GTvGVVB
jaAJ49bFILwBhepafZabiZbPCeQ919UTre5ye0POPKH7aLyDLKkvISU/jaHjfW87
LSUKr1pRVOq9zHEeBe91nbgj0vHZaPhvwBKB4W6BFfyyd7BqRnsySuCyQUueJmo6
mKZH4rfE2PlXtDC7Uns3o90bkhVH2TVZD0c6g2LEPK/aBw3gnoHMw9wQOioh5E8V
vqeVptaNiThyhaPxkJ5NnadEeieHxECahXKXJ0+jV4FsktNU9fTcvNoqBcvXFyAs
FcK4kEYhEuwTrbomrMRsfHt71RypREV6LI9riTpgfWETB9hyzFSTk80OM2pOmOSF
LCJpK/j8Pdv6v1HadQPkuMOzPYFidTo1o6eGrDkJJJJH9fTLZcMRswNI9FWmcxm8
Xjx0iwgKcRw1PKFWM69hgDRmSs1UWIYFad7eWUiEXLwTA5NrYAcXwObP8gOt9QXC
UngTIaNysQyFGjW4mXKllDMhtOowZP5Kw+ZKx16d/MOsd+sb6nA7/PQgT/T5Wlaq
qzRJIUIyfNIlR9t6sqKznaFWSllxFoSiRpEpl8XX0bvCzGme62zhyxpyYXUAS1BZ
Uf9kslzjvTkk6sRUQ3XbVUngqrkabxfdBFoOQ3rU0hV7e2mpgtE1tvqIF8lEty6H
j3TBUYLNfhZ4RwOe48Hqo+Ijq/fsqY9yqNOSQ41e7VkLTd1CZkrUpgaJEBCGCSR9
HTbB2iR9QxdcJy/bHu4QkIM01WtNgVKzCAq//EdPyjW8QvcfUWYxlCCakA/xZiuY
axRsfDCoutpIwBzHpzCRQpjteBM5CRlu3/BNjMEew6hazzI/weVBeDrDWmlzWWoo
DXXUh9jBWVXUcmXGZq73RG5JZgqXnvv3J5t1iL6NpN2zslOPkO7qQCAFWUCG4NjF
I8jCfeP8W4blNljA1L8IzU1TOkHfHm5RPC/V2IoQgYNaYVljhcs5U4P2PWkl7L7N
sSaEsoyc8YZDEFoCj4zAQTb6ZFa+jSfyAvn4nSQyIN/884AHhzDY4NdZsqU7XK0B
Kw2jr2Lqc+CPu3TJJAm58Rk2E91e2KRCLqYf9PiVmZDb136uEAa60zw4WqT7en1/
j0fSycbEnuEv5uUDHunxWLQj2+CZtPgBXstQx04I48wOMzsG3WS9ampHvCHICXWt
OQOH+58Pd1i98cjZpLRnCr/pPqo6DXVpGUf6H9nCYa1GX0z/M7AmmWUkPaSDdEQ3
lEAUgKLQhS+NoJXyuLJy1h8kaabjLiEdnnkI74pdkVQO2vSawkqzZhgaVkObKOBw
HhOXryyE632R8sLRVjdGMy9O2nRawq1n7Qsmz2St64y1cpl1YnyFY6r+Y+IJ1QYV
+Kg2Mg1sAoNUi8ILHXzjMmy/HI+UxaK0GDW8IfDOUpgrdintv/38VzTAsrndvEjo
Chi9yPd3v5YCgVyijEcXMXDWSuOtBw+bxaqcjzSq/jILKqeAq2PdT+LJJsQjqaDI
9oHYpzc4p15GZO6+Pa5sElDlRA1O1JDISi49GA6XooUOp+R1+oDcjq0ul61d8dKF
FXtpdq7KVbBIAy6eF0h7+t8X/ASS9VkQ+Ckg3ciOGVmihxN0MPTv7LmTadmdQe7V
hZZjIvwdXe3JWeUCotNIEKWOMBarOM09LiktrJNMBu4VCrG05d6QaHyaVI8I8ylU
1LIecSsKZvhKt6NROTKdpEXQp+gUCNOtgvN91Cs4EC2mz7GNrDehBa1nRaxm/vhz
Z4OQID8l0ZXO1TOnjouygX68CRHJqeIPzrbuf1SjvIYhXbVmz2VGTcz79jwtwz6/
isPXmpokCq3j+8lp6kGb1jrDcJn9CWrJZwHsAECFyDke1fdpv9WtFFJwX6hGDRXq
nfYMBGuR7PSzRIUUtYhO79OmVgVE2w3L+iD3FilsjpNpLk1sym7OVRd65u1K3ATs
dAx7i8KfuveNC+9ARO5qaJh2USwtZz/pN1nDvZ1wjf1pZrbE9c9z8uU3N38lsoLJ
MRELei1iXgtCv3Uvo4eX3EFZ/hFUTNSXbsVAjz96uIHYkeqi60HgiIm043MdD3Py
x6x5V8GGD9ckfG5tUmZx46zBwc4F8WnAABvLd9poFCUS4h8dGukLxWCc4rry14Ss
aJKeY1g2TeQ31IfIoVOhCgd0cWtZWpyfq80ZjK37cqY0RRQxWe7PC2/Uy6HQ8VmD
UdpTzhHtFkIHAHnLeNEH1MhJN8yazJoBS7pkgc+RwdzBPsPm/gQ89SStAsoIx+DD
jxgsfuJYdljoGJ1uBFyrYVhMwv9OYpYvX8HEusWIBu7YnqOpukP1a6McLAAwf375
efh3Zs67EhPagXSQpSAf70iTaVzI4ba4EI/NOsL9W6I0As5dRuCjK5O9Hq1b0XEd
hMuyTalu+JoCJ0fYCRi0stONcz5tHKAzggEpE9mfSerCKAlbB/2tq8Vr9MtMfXw1
lsRjDQtK/uwMcdBrmdjNXRRb//HxbqWUvZhdjOz8q4CzqsrMgaTrQ0lVbEBU/u/m
fFVNpT6PUfFFMTvLsciZ6SAFtEKwRiw2pIn/H/rwRofy27snLnACaBJ6lEAFmD6Z
BkFi8DC/U4pTj87VxJWgLte3YkNE+oCFeyoinBGQFnc4+yVNJiyLXXnUHaq2sump
pq4VtS5Oam/OI8PZvtPFSsmFGSY08+Lme53NT3sU0ufZCiCNhioiKn3TsUpvx6WA
mldVkq5H0NtCjNOP8JwY8pi+6JbXLJxvZkLCzaQODi/EcX5yxebd2iK0KaU8BNHz
5ZZVSVSXdmx2/79NOSq4BCeOR6dtnF9fl8XTkxkeNyvsn6PcFYh4IcJyFdqaehEm
oVMcGV2RfG/Jj7C0pEz0zAgahibF8xagT5+VnKUS6SIOExgPpJBEqTHALhooaiEj
hP3/CXHLMUyfJfv/+7yOeIfqkaiz9M7bmHWGWdrcCe+BuM1r9E+qWQFNWRZSL2Qf
RYMOAGcWlbaLLOxIpxrMT9VjBRokNUlH1iAKg3tUclyyYnahmrEtic3XP+yK6NYl
sMg3IyOU+QwCRIVOqCvW4y+sjmLV902nCzkJg2qsu+vAb102xauvxvuHX0ezne2x
jrB41D0c6sAmRklNpnuFhAMKOshbJxNtfzCHVB//htsu5Y8svkjPj7IMhSSXnfty
B0z6HrTVtXVl8Rx9ob0nfCSOg/ASyvzE/Xexf319ID0=
`protect END_PROTECTED
