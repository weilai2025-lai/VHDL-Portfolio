`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJPDkq80ekY0d9V4TeZX6UDwWwCs2yswTtECcs6/K3Op5ETUO3HOoGA/wk7J1UO2
zQsx5e7sPzJGsu1SkzGZsK5uDIL7xB0tZ+CQPHdx8rr8rGtmF1gt6ATmLrMoeInx
0OgZcK8oJOCVpXhUMxN+9qj1G7fWWjK6hjrQDcSvDjo6MGCC6Z/kKE0ZW1fZJnS6
NAT1lELolt777gf+6UJfhkWujZQAf96tq5v1tcl5mYSlQQCdXv0o+61gdFqGGKSn
sSduNZK6q9mTNV1Jt/in2ZNcw4cPge6CFp+NEclzzegsqRkyWHccqciCyAeTJejs
R3KGeAN4GvHhbni3C+2zsj9GE3bEgfc6jJWx1nMsLe1cGGIbRdgix8/Xdm6ys1Fk
KdLYDroXBLIlF77KQonq5pqSHqRvJzyoqcpmagB2aJOTNvVfL9P8ATP+EeG8Jx3d
eFgZ92UmsBxQbRTW49a4GQFgw58NUpdEpUffAHzSR9YHUFug8JfzFa6QNSkGvPZG
`protect END_PROTECTED
