`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hiLW92KI/EAHOKG2t8YU/ZZMI8a5IlvIRn/7hs1PP155k5e+wTQGs0Nw6MGarMy
wNWQ/R/DBPq334HG33xsZW8FBxErgf3lZ2r5U9uRF33kqnrrHcOs76xSynPu4rTT
90SSTAsVrDBcW7rb8J0hneKmsdatARb8OLi8phuKi6NUz47dPIJmfFBT2DLFvwy4
KFBR1uCSpQ72PrY9Wg8+j5ySjzaOfi+pXJy1kpGDyJrTyLuWCRByW8ulI1w4zb2h
1YFiOXnUTd6MeFiKw9PLFBk4cp7NnaGIXLY361Cwe37p097iuGFLaC8qoRE46/kG
9jzUjZm0WtMDEcRcGtSmMrCP4EzaCp0haQYeMFoD4NDKPIm+4vYWm9ViMMErJVlE
tIpnhdu7Ij0Zaoa/xhHkMHTM3tzwvzHKu1uo5Y3nwMBnR82B2GOZqp4mw7ODuw8i
tdAsoICyVG98yl8LYFKcYiFG22ek86zYXHN368fBcfz0tlKccjPtBqwHgvYwS+Lf
wgdATwwtuBpkeCwbbE6C0dp1Qcl0lqPqF1EocYAOtBlB9uWQJCJcZLoRnju0vkbo
8ubGGUQkpIfOu8OIeJYOqr2tsanHobMVhOsY2Do8xrVL3ivNGh5cenrICRQb0z/W
hzw14tqMsDN/HGDQPAuqdRxOaqcbmM1UXTbOu82Y/YF+bxv70id0DLOT0ieIKg4b
msVSetZDI6fN+Enu8DM3I8Nm0p1v37LLxIokKt4xK0Rm9AQk5zVfRgjd4LT7A7JT
lyuF5QcstpHEnoLcpwRb9BsqR3CHaof4anbLY7SbmXjEIBOVQhvQhyTSjXfx/kUF
UE9ijLjRnawUR2aNODZs3Uas3PaHyndrtKvgj2WVDzlSGb0ZhLE+h+VwzUwjjGNE
NLlh20wwjxxLpw0IMjQTDnmcmgepLpNfvj26YbNcEkTl+/Qbk6q5F2GjNo68DLHo
7DeZ0XuSxKemkQFypJjYlG9YOF9W0d4O0gZGCMg0Uj3mYmCNv2Gp4B5WrXuv8H+O
76y7Ey8EWGGh8/iCnIutgXffeT+nk5w7xYfERgT8EpXncRIXmBp/CmSdQfjUYc9o
1g10/pTNdT9l6y8qYlkkHGE0gwrqhPt4jyBLlOJ4aYfkMQWkZfYQ4n+m9xI2rY9W
SDLTQYxECtZg4Ut57V2w15X8RMnXr6wX3jwlq/g5n+IRLDouf4lQyt4oUTzZydhZ
zf8bH4uQ1VwE7ZqhqzsFSZ0dq8XK7pYpAqEDrcXB0YBBsu3XejozAjm4y5eXWd9q
6LKgVVIj9zuWrni2n2Sfa9RwIWwQc7cVVYRAgHb3efCJ4qpm9JlH4oGyAGcht1IM
twgr/jPor0qPc32pGFVIX2X7riW02lnKv/KUZO6wrfelb/Fgxp0qwVicWZa2p4DB
YM/k6CJUf0qVCvnwbriZi28hQwtSEmRGpoSQ4fmYaSK9QTN4yUbUbkDkFZa9+veR
EJ0dcRIqnKpw54Vy2SofmUIpE6VwI3+c5TJJFJIc98T9QOGoHnW1Ip6kCRVGrxSE
GM4cthJzYMC3DGQjZQrlxs3+WDeiXA02ouD0Zouaz/ObcX2L2iQWt7+2JV23QksW
+HMXoF2K74eqaKl1nEdQKfhDlRxNgIHdKrWdvHRBDrMLHaQfBSDXTsgKk9Mfw+2u
QG/3q9p/ShHHFPAfrfCALXAIilkQC9zeE+YpBHbQdIJnmitoOluYepMYypbukCbI
ZeXr/mmWHGsWDBUUgSVB9azXwIJ3WE4+7VH9N2WokevQRKdKtYt1su251Iuz56zc
pxe4CkG1HTUYzKy/LKuRoya0MGa+igFHyy+bA3wW8kh8T6YAJdrHgMW8/p3ciQ9D
71Qx5tvlIVPnuLGhbeQHk+Rjkln4K9QT8uaRRDtvxvrI5o4sYLmspoZ1nPj7XP5u
tbrQeaiSfuuHSjxONCq3u49L6ma2FEIFiOZhgnsrNbc+paXy1PPvoUk94FklKkHW
A8m0lJ9Q03o7GThrCAl76CDlCeBzzFHCHpyGvL2ulqe+ife7EBWgknovwhEMa2mY
FZKazKvbo3jC0fZ0JaBF2s5zYB8QID1B1xAbg09KkVZqDABca57AOSUMnCXe6iwB
n5vKMzc262lNTXoNbWAfDq1HnAdRlKQ/adpBjWXIWDSgKowk9opnVJR84f7QllTN
T7ksHlwIzviPQpRg98VdcgDuzAKz060ZFkuFjpsQGI+hQq01F7cHxw5pjmgmH9Sr
NLQMbMotP4j2gM08iW5XPYTlAfaEox8LC46pWUwbn+H2g47t8Pz8VuJTuJs3fj3k
KAMt2KRwtjTgdr/grK12v4rpavjFjD33CZyY+RwNrO31ClcmsYBsStdxvK2xsC09
Yy0Eiem69DdUXxsi1JmT6+V+6bQGZnqenTQSa2DoYZQsZXmnjGnJZ3gycuFai+ON
+D6VhPv3WSuexUAJl9UxClSzBvQAyIYURdiyya3Xso1dpZs4lfy9XZaHrJpQQkto
ttLwhtp2b1FE9783OaCaTcgCXTf2yff2xlrF6gf719mq87efPiQKWZHYb2Ljhf0u
Nex2oqrGPo0w7IyoLkrvW7U/Oer62C/SzXH5oCrYvMHlRfjhjRZ0Unzq+oiUP2cx
VaKNIv6ldaY4f98yTy/I9qwIS0KaTJ37iMcfrtxxJj40PTrjQQIP3ZJ+2a6iyYq9
CZDgweU4oRT1SOkdvLFUu5YAMJSWHUsFyizym+rXWiFFKYSzcbyrwE+I+iZ6+ZFT
CZGJ87W7pz254MNHiqVp4dXAOn8YPZRgh95+vSWzexvv73vg5Oi+V3j3f7Min7r+
ONJI17pNv2LYlux4X+m6DWjTAJKBiiAcSboAtWHEkayd7YYKrhgA6ADPW0icoPUT
Y+hpFkJ7WQ6MTYUir2oJM3YBjeLkjuOvBff505wx/2nNKm4jmB2JLdrWQkqP7rxV
LRNP7IvOFvgduwl52DkVGFMaDv+j8eJHkk12RuZLx2aVA8TJgtfKzJ9AKBgf611l
l4a6FLFmPiM3cMpRBJ4w+f4Gd/DtYQ4Sfusgxm/FM6+vkKTfVhjv0QeJRBmTyw/p
BReTkXyjjvMiUT7LQoU8jfgVdoOUVp6XslSG0H3VfMM59ZFoswWfvEgWXGQciex0
acpyDevOcZwMRuGso+UpeAnZ8dUZGB+KPFXY9YiiVKAL8JbuAEoY/iPwUDax+soC
7OFELbozwvdQrxCTdDUXZ0/N0DsIMeJoYeXOGC/GQsdbzwSV5wZ5x7xYUxqIUSil
vT6QrVdRQpGm0aobkFtpnfJqXssaW2LHX1hyBiuSV+KuwsRS9h9kCAVr+shLc3is
ECAtBTIkyzzWPxt8rGBBOgAsm5cb117eWCdGL/lr3e1lfTGM1xM6ppXrMPV9xNF4
HFrDIXtlMwsDmx4K5gMx8zMfOQAkJNaN572jCmQ3QpjVBKFGxc7i4Ueg20kH0Mgs
GIi1adCNB4siyCUkIxHCWhN2NAKJ8evH8aZXRH4Nl3INd2e0iihLkgWIlPZHM8ph
npviDVvSXvXfccM9gRpl8GPvM3t+TbJIsLwL/xBezH3VNFTxUCWbrfzzKNvzM99S
PH5LH5C9FucVqqYBKVUwiXrUMTsiN/jdWfAhNkuVrSf+SnpDxTw9v7pIoaCvDMqz
5KPUnsq3xCtHgFJfggOC9L5h47bfgg1aWLyrMmwUEL1BZThZrvXzp+pPBsSaopQJ
OAGdQU0JjM7KxJu9B5Yyv2znChHo1b7mxJmxH63FmoJOsEIBZR24Ns031E+k/Ba/
dzH9APEalHJAJCyYmnB3qOMQuFg0sSdR6XrzeCI/b44BOMDfabO9LxZYWg9MoGXT
0JqG40m7Jwv6bfUNEG72uIujMY6w6TeuP1URBmnGz3AmEtXD7zja1l7DidmEwuiF
060svWBzd5t39ruh+z0cGBp4a2mAIIoa7CVvm2SEnEabQV/rAD9DSSiSziIm0bEJ
q22o5UzGQfRBNmNp4p4GsnV/AlRfpVyVxRJeHprbzPYfY/tz9QzdAFlFGFEdwHB+
DYiMtJrNHQnoB5I6GWz/pqrwucPmeJXOkNiQ9cyNr7MmyZw2LZCqSrddi8H6YIGB
p+jp08Zc7jYtXAIR1A79roZx5QwJ52Mub0+sI7twKF38muZoyIjD3Ypmj2mpZhHx
SHi3gHgG5EpKvmsDenxO+Q5RVZRu+zkD66+CZ0sDnBvPDg286qwgonYyZRjooe1H
eZOYKVLAqWt39bViD2kTzd7bWSPLI/Wvrr4RF8rk3I69Bm3KE/NfOZzuGy/ETMgU
Ib0LHX+syokOk7JZg0+nsjoAKeKOhQItWtTyHsYj+DZ8ywyMEzdPeWAm96Xv/Fxx
ZGRDEo93rOffBX1BD/6I7Npkd1hJVCEj+ioEf9e7NLzDv8qAkyVVOOJ+km9ri+x5
4c8UYNiHUEdhKWum6R3w0pBHcTwKkkC6wBh7C7FZZVafWTFkGf6WEgtbHN6+pdaj
JgI9tHVB6P/47YrDQPJKop77hPLMpaLxeRxzf5ZVlPNrIV7PdyfCbNawgJY4LQw7
9YY+0u1NMT1iqtMzXrrvfK1EN3A81NWVbXUksQn8XR5y4EQ8ienntAdWaxgYIrsN
wJWvo6CjYSwmnza2UdfMDmgeNjyIC0j5sMMTdAmDN9FIKM6a4zAy1yvDGBXoTlEk
OeQyJ1WR70Bjw/lifujMHNq+aVy2yfrRflOG3qdPLsgO+GzAAKjYJfu1OIYOVNMA
rdX4ZLZkSwip7dIde1aNspsw9U3HXPrrRdyNMxNUqj7RETFezD9DBrpIuJpvDZxB
OIfs6FsJx/DJegdMKWOkjFE8c9HYB7paWwA/d8QardcgQinYkbqYTv1LsMcCXveR
gmyUqju9+2h7g4BGFf0q/6XYcYQGUs8DQ3Jh2cIjuDkTL7iGMKshXQZHp4oUBC+y
arCOxcBoUccMNeLf3y3vgHlP24fZRXTwswy7PxMPR31fpoQKLVcTOwZ09Q+rENJJ
Hr2Zhf5mLq5FmiAOxdn6CmOBa6JGzFIExc9FdqRO1ten7YKTmKrpjXFvuZup4iYh
xND3SRt3npM8kH73yUb02DSeWOqvtb4VS0n8NVL2TcwP+H6MH8/VhTHRoClgZLOt
Ni4nmzPa/qmdEIZVon/yzPvUSeyAN12zoAqHlckN++NUB8i0ZTvisK3c2hCExUUj
3NdUFTqMwaMCdJzHCDbjO5FYK1RbdJ+Dvn4N9FE0NwFsQ5fVMaz2qjanTpErYDkr
pMF6FKKmwZrCdIwq3HTq/+GZA7BNoWJ4+vFwYa892s794TXknl2aCa4cx8ejCKg7
KEF5423dPHmc/1Cmsc39eUnUeLYXnArGc55bdTmEeYqWYGR0F26O/sU5aLmzHlI/
5q7WMMrCbdxwKiSrWh64cRiC4m1FbSFNIYaELk4fFDuo6YLqwB0vdUGwtDyfj5Gj
iZggdDOYgQr24uMN5W3d0uhy3KIBkAZloEFgWcKTHYAOkxcCkmq4/1NfG5cUGsTi
0kjh0aXQKHRmd1h0GDomVmBrrUDo0BnGUJw9aPdC9MlYJY3PDoeoJmOu6gcGgn8F
eX3abH2SR5H6zbwxurLN98bWXyHZAWDhygYcxT0hjG1XvbuSTxWgeI/Gv4ZbsG8o
DlK0JO6Ez5Lo7xfTmKNhZnKkJ7jljxDxj9KuDauIEoPtOgL7VNf0g/WsA4b5ajoD
nlE3fQRP7/lHewz9hfbBHobmGPJwwGVZ1DadtPdg8c7Xj2Rgep1sXGO5EygPS3kT
fC2OqEVnvhTtyCPqhbBU5oCDZQ0e7So4PX+uUHCtxtPCQyZvhXF4xhps6sddQGlb
ltYK5ZhnJpJ48Lax/Su0Y7srE/GySzMHnv415Lx8v27oqpRRhu+7QKZk8aqp2oFe
u9QIx9u57O9UylXBXkar4DElP3scnm1ahsAFt7HUuEYNelboJktMEmMZkBnJsJYs
dSoHvueN3YnC6ZR+SadUakqNoK1O6RQh911u/3090A7m8oEhhk5v+m5l3mYoR2tq
zBnh+L46XgItrp2V40+5dUSFXv4JMg6G0y3V5rs8cQR6JqYOe8O/H4yMg4g7NxKP
18dKHtA4IHeItNlr6FvZIVvEZIFptZZaye85LJVIKpBC4z+fYSXbsHqlPdXfdsZl
Zr1v4ihVir8optTGms0rH95lagjalotv5SqtZTz7jMRVRGLnDS+7Zyy1d2hsdaYp
PUh8EFZO/uKfd3lcAcqsE+UbUD8J9G+gUf74y1pS8gJuHAKQz7v8QRnoD44xPABO
QQYqYDNs3XGLJmKG/UY7n5K5laHy+AlQryD3OKTmFrOl42dPVG9O3Uugg4jFUPXJ
gnJex3fJqCVuAaaYlQ4F1kFTrhbAlFhzaEGyBgw0TuGPtMbRuTsXCsH4R50I+kfh
3ITplVuglV3EqctD71IL+OPBDdOMAjvU2enyIY+RpPTjljDhTH3e9KWq/CBRzTXg
FilrnTi4/u4SUIpI1fHSf/GB9xnb2DWN68l9ca6FmmAULH775r7rNynC2G7248xi
owW1ZX+TAKkD477sU8igwBfDkRSLRjhKSK0b64K6HwEzZKZFT3J31nHXxsXxqO2i
q7lUrT8JlqNMZXC97U7MY4gYrmDqMgezUMRytkkzJ8QhxD2uDN9HUjCGGunSHZHa
RXPbqxhljKrKeWI1Fc/e1fAJD6Lu9lIjGLgVK0m23umRY2Y0B6BSMMlZAEWdZwRq
nxmdh6XjB+SukyOAKkVVsxQGV9SB7z1hh9NkwHQHYld3ekurgJseeRM3CAdcgj0n
yNMYNL5mhMATLaSJUg4AK+LxF99VAydK8XOzdYJQXEbb+gcSgvGsFbGgT3Bkvx0V
JiQpbDbp/0wwt1UHipnyDg+/voRe5T/cZ8GkAmFJL10XAr+Ks036KhHY5fT4Piga
qvCp+BLrScDbDofVinNtBqyNT1letrUCrimCO3N6OneSvUz/8S/bjMfg68zLycYm
GRp8mLpn4kdn/quYy+Ce77xiUgJ3oIelI8cWberaoqAKla9Pcp9xpQx37l0OCm36
qTOtV5ZVciAa9p40RR94/AAslBVIFv5didOwofVATsSQBlIqfaKukx/Iv+3nx3C+
mF/K5khn5kLEscLML2FvK8SBbEVFfZxRNyJ7OEv608RXVWtcbYICNhu/Qksyp3KP
1XBbOC8fwPA4oTdeXhBDThTWFirWQc8wD9igID1eK13lkQQGZhHDWxNA6VXj5+L3
UL4drvY3dyfF5awuBv4LqPDnCA95mzTX/Qrf8Ds7K75Bfn8Ot4yjaKMfT//4xj45
zXsrTAgxcuvVMtMtJkaBE47X8qQBMgJ5oKaH3yJKwJ2dz+CAA9RZ7YNNS57rB7SM
K2f+nKvnn2YsOspYH9p6ziVgS8xKKFyX/U7Ub2rzj2IaoqJbPye6QdeZ5zUnrEQy
9urjbyv+WeeXwdL6zTCO1KPEHsCJZrl1r22d53sZbUB8Nbh+pcPIyKhuEj6NRRMA
g5aAliM0ejTkb3pyD4uXWwUp15wZVFYHUnroq/B7qSrlOZt3NaVwtaf0Pe8JODit
fPmLefQW8etJUb4Dov9RYYkMwMoEofCknL9DKbfP/bcQg5ahqQcbO1D4Q0/VKjTF
IFxW0qUWQ7GZ59i9/7MXyMADswo9PoTOmyegqj+FnKffUCIaaMzUstrNFZlIwEVZ
T6HZFWT2jRPg3G27RZUI1SC/Mv7yPQEXrj74uiAdj+cdA8zz1COTRRFZbewLeqlO
+rYIJCsyXBYJg4MYWg2oIggXErHmE0fhOWZtqYSCWDVBUsle28qENF03GXnc77ys
EN7KYpxglwt1RWPJPGCPJ7jCerbkdrOpUu6hPLNVPnO9VavxWVoKS/14PWHK3NYx
NIsfNRb+dgE2cie8yRjftoGmiO+HkTlhCvLryVrKFiDCIusZ7M50e16bkS771wMf
paLglVQ0XquIjCLRK1BjPIX5p7nWDOLGrbfNkB+DJb1cQ+7danrpKmO34ZTn0J4u
E2EVgl3ASSlrT2GNJ5FVqcr83W3TTbhIArg33Fb2Yw7AjJpvrtBDyv1T/hbSNOEE
gD5spzOH8Xuv+0AK73CjSHkzFXa10LfT9E1niM2kzAVZ0kzHc+g+8DkDYz0MNb3N
JUGOImkqQQP6PIjiYyoacfWU/+O7XJ+JPWvWDTi8L0aAWT7tBcdVFyXEAWo8pa+y
5SfN27bxU3eWM4iX5GfdQ/fJcWFSauX2bYqaPL2ycPaLqulVqDEpVk7KvaJm71mb
e4Q/CTwkJYf80HxBndd7fdDhU0fZKtWxMaAx5BASVLLWPPM1pcbzdBNVXu53o/H7
Wn+nXSSwGFaIkkzzj/qQ0S8ygxdoWDvmWRsPPY+E75M8QwPRSDywFSf4jFxL7nFJ
JVBSq9gJMPf/isBgAblg/GMEcweFfrL+kVYJc/TTZZufSe8rV80lyNB+NrdlaMkJ
sKtjxwcUX+j1Ae7lJdyWB1N8G9X6CxsW3027oNEI0p08c0WLDrhkIKWgrK700diS
KkYaudX1MFZBd1f7UI0pvJJvbFp2dEcZdJFWNERvRPB1CHqJT8MG6WJ/6aIcTcwB
HUE4FnIzo2J0laYeSoArI3pyPDq5pqyZBMQ/IGeIJmMXQ8mBdYaU5zkHKJk07tXS
wJhCb1fd2N8KTlJlNi1Zscv00ceHV82QAnZiU4l6rc3JK4dAyrEetO5PvoL7NpgW
DaDEGoAooxxV3ZrZtMCW6wJglKNRx9CnyqxPRl1AC6ipSoOM+OzdRl6NaWMqLRZN
A3OB2JloP8hk4oTn759CTOPqG701f2BAEbGjMmqsCT+viDM8uic6pgCsHzzO6fhV
YldKeefFil7rmTzKH8u5pTSG76NzfdB2UP/RfLml8SdkNevkgovpTZFb7b+UyDCp
PhaKERynJvajNKJ5UcepxQnNk6xQmBar/0hRL3AsQX859oJwE3sxhdFViQzC1W1u
4YkZE/EpzHBSCBAkIOwvPraizTw7SW/I3Tm3XWfUtAARNqDuYQTeYbzNmBL+I1fq
MSIrs93xqr8VjGu5AzzVyy/oK16/CtoNm9JPXT+A+ft0UrbAC/6t8XmrfjZ7rZ3G
km5ob8vjWmZJczoxlndZgXY30fTT05M5wE1GwTq++QF99Mxa4SsBQ1cLowCCi5Tl
L64/TYFNoEA3p+9w95VkBFcveu8BqxpJ9d7byesmKvZB7Fg+/kCNZrsjZGdIKWZS
UHITVUN8BzhQz2tzACe9gjOMyGdQTWJyph1OlCvq5daRuIcv5Q2StIBCBlywH6ma
x2pNx269vs6NIwxlnrHXDPlzxaJhxt035dOskFjg6aSjNLRHGYwnuRzvLUCer6oQ
aKnlYJPn3iquppFKl/LejAEZ4BXf0LHJX3Ahd4x46FiOP17uq5+z1wEbTpxgqrgv
plrlNZWcC3gCfmDglYV0TV3eeCSzZXHxB8poF9668rrU0D4Bn7yHhwuN4Pr0n4Xg
YSkssdZSKfrz/KmSP4djthepDIt6Tf/TuMnGD6OpThAw0IXqO2CAIVMGX/TOOxrf
Ml5ICgATFUzbBGgdMjEn8EC7YEduNnEew4BBICnCyaoxzhunmVzmOmUkt5PKuYr3
SR7XYo19v2vPYrLzpPvDZOJSqEbkgbjq8epZcJx/Aw66YhhYlPBwUaIalNs44ZPX
+ABvcYVDEi/dShuUaBL/5sirzOmLg/wIzyJGCj5mMcvEdoQ/uOCxJHjDWwuhxCzZ
aqmqi+Z8qH/XWP+v/Z5/odwgLdre7JXHYUTBUmnEHrXrrY+kZXJUOI6GuLAaWm1+
xyK8TDFvfl6Etr8CAYB3nrGm4zrNYWwm/WxDKSTmiuRrtYMcGYwVoIaO9aTiDliR
DiOyFFLKer8gMMsyoiySsS+FHb6uhU54HmryrLRRhzB4hZvGhoJKiOZRAOjPCRhN
IuIN6Q0kdS0T9bkye517Km4hESHjaaGy1GlRCxd82OXxjHdxFez1ztd+Ou4Imqov
fHejH5OX6m8r6kwrlvjC2zFiVQ2oTHqRrG1VIXXTmjiisa97fKeD5nJO6MNFp44E
N4fVWcC86kVRdrdQV4qMQtIKfexKmV2hLXohyjZLILnHu/n212Klk+Tv/U6jF6pp
r/jeekiNvSPbn5eH96qKK3WajX0miEiLYifkoT5d3K4w1Z+Aq+QUPiAsLmQtOtAM
284d+xQvgmvbm6PPjjmZ22cMHD4DMBOTdtak6n5Z44XeZ8DBBxlMdnxKAowqON6c
js1XYqRFGNtVbmHCd/DaV+HletUNKZIEtslAEWHWJn0=
`protect END_PROTECTED
