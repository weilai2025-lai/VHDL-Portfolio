`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmZS4/BQnABuZLdQHshAr7bozMaUAR+1dUBNZhdei81hyjBjjE+Nm3ofDF1Cvu7A
0GFGDuKoljhNs58UTF6WAdMgKj4Ck8Xbak1nQkulOxYDoA0Rv7JMcf6w2mhbJ4To
fuxG2vTYvTwcAaOE7d8XBIITzWrISCtp09IbMHBQZkjTAjB2hIhCnkt9YCWg348D
HrTo2fYFCM5Dudm6usabKv/YlVqSZFs8sW1NXi2wBwc1RtWnW0UCKaM1RJYYcYTw
zm2dMfa6KiQzgmDAvwoS8vLTXZSCSJZ4rkpoBckarXEbJqUDYk0ywT+SQLAT+tzD
mZk7/Pyo56SbtQqvLey1likzUg2gfHcNBYEbRng9NOgQIWPkvR8EQVOaY4knhV2S
lWZZqaWkowhNFdqX1UI3lw==
`protect END_PROTECTED
