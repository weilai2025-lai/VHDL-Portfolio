`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1/zWcf7b7QZN7KVbyCZd5XyxMCnJo6p+XYrWHPVFLnNWR6a7lWaESJqEF0tAYah
VolS4stAqJX7bYxD82lHgK9KLoGBDNhlfWKMdjgxaDXebdO4MQeVNAGXFg1iAQbi
+63tK8geQFhKb/UFnO14xV+bSzclIdWZvLZvRkHAkbEyPxlSV72HMOVTsKFW5HSa
HES9K5afw/IXGHmUKKB/DcpaVyjkqwPc0tYG/jeyaJkB8wO0feR3zPHMVdMRsmqo
UeMNgpHshtVtTVoD4AN+pBlTEamnIwJCJZa4H1vHUQpn2DYWshspPm/EHozYq0q0
pxh0TgubjANh5UzhZEZo+kKIeokO5d8/2JV1Lt51nqEX+euk8yOpNeZ7Yo/PsoWE
SYkqp0L2lZrha9vYgPS3s1bRp9jbqHudK0imp3c3L3+65Wv3c9YRS9gCIp7Bhuyn
IwLqkjjk8YtX1akFayFeOCFH2p2hWIZYztMzhSL9y/KISVf4I4OThhjLM02SNN+o
46KG2WKe8c44UeEuMjNgNuWcTQ6VcS8sg3AZ36ODn1Hx+xYkNOik1qo9yYiiiKY9
o7xcGuXIFVTQWMd2dVmrq79GRATuCwE+dJe2nYdvotcaKrQcXH2VSNzAmMylAhkI
7L9NP0JY3I3Zi01VDGKzSoAyQy+Za5Qhz9ipxi1GwY7plqlgEtf9lXTAx7nV9OAM
P6DX+3Kcg77LxR0gJwJ/iqM4S7yH6pXMCN11NXyqSD1XYheezP/d5KI3pNPLQrFZ
E4ERmebYGyPKtp6YdP6Rl06sbwHeXIpzIiUGLDo8Rx0s6Gxd+/X3rrfvvPUkbIh/
p8E1W3YNS+/ELFp9CzK/z+jh9iwl1OH5GWld9tZhq92dEvlOUHpZqf79p951cxJx
Dl2/7fMgSGAJ0sdvtkJmDIDi+teUHtS8rK/lq06imRoKRlAvu7c4JlYBju9N9Zt9
/perpfFgz4Jen1TEKpI7GQZE6OO3c1QhTo8l5h94HWkyYVE99dmaucLCobEGOxSH
EldMaqkPEP+pD6lRKbvZiWqps1JbIWZP0H15kmcTGr3mEEv8J/9GKjjkeehshDa3
IC6mO+A13zNaqxl5ytqvXHg86j14F9iAHxfrgdpObwqr21ht7/1hmJ7gYGmXV3LS
dET4CvkB+2T8t93U8sooz5kCym2iv2WTrM/h7BHH+Qa4kF3aPFw4FOuvUHUbKKxe
HwYtm36rnBeij5BEF78GaIsbocmOUqbwAos7ojds9JHbynb9PpPb2T0ASs866cd9
UiM8cLTPYqMoJEALEfQ0kqqCcbBbaBxhm+N6e5fjzVNZtDLSeiIpQNISrtbwe4zl
XC2Is75MnTQpocvHaXer6M/hn1mjQqae7RDKBWuKi6xnXNbTHq452NZ21+WBPYK4
nVHMLzZoGYVHVtN3LlsgFYiXzegxthJn1dcDdlZ0/xKVG2SaZsYwk6p9UdjO+AH7
x97kwQCLrJmaiwtRpQu2z+D5NIEvVeBJuncXZ01Q4pTjedWkBLEEbQ2hmVkTVNfH
a33CUsWZvFT5CgFVQM5/9EAPrEqZy3VwlEM6tO1WIqKGpiYOzKnCTMhh9tKrUsBb
3oQFY0Qux3UVWHebIwY6C2MpO1mJGehLuA/d5fqIXvE+VJbQS6MVBSwVdetwNX2C
lGO8Jz1u9YunQK2VB3+Xvk4EKIL4JiP3yWuga0jFxX+jh1uFLIkhYLetPLS/CLEn
T79vbNJJ/W3PMoQ2NBzthg==
`protect END_PROTECTED
