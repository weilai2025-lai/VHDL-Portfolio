`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pw/7pIJ5fiwate3fEc0kkMPF3hugvzTRahEYSdJi4q0ZN8F0/UxVSDZu8FOkndFF
PsshC2/1Y7HlRjkf0CEf0q26XAXrYGsniPbTRrvAdxZ3h9yiwMpwQDU7hIVb5LxV
5h4ZTvASRM6cGNf4ve/u11V6SJ6eEAlCakHwIXStRhrvmHXm7vJQTVqIG8yms/SF
GhNpx8Xqvj0/9Hnzxr1+0IKVGKhZ7vAx5XSgEbPjG6nhdExiv/0x3vC/u1zMH0yU
5n/vCd6rdDW6sEZSMT9EIxWK0lzqouk3rQzQBaVRg5mNb4laNWeadO7F/KjlYCmP
AD+Eop2o3i25922VrV3bTuwItgvrH/8E+o+CpV5ZCzZffisD1YyxXaeyMs9aGFGs
eycmgG8eZWmSBVS1JCA/6AUfOVfDqs3lOLIiEukh6bygP39XunSayMZb62OwmO8U
AhMfco4+Vbyhh/ztsH2h8VnoMT/LULMxr52hSwCUIp1cnla9bjl+9nVAzCJP/Xe2
G03FBq6GsdQN1YN5zI/SE4McD2KMF1kTGXqUV/ydyOeJTT6A/aDWjaWvHMuRkpbz
Kj0sZtXTWmFUaH4Kxd4TjZ0mEUubOFM+WVKyPaQxyZFPUC7laoJIJK4vq90+zJvG
79cofg/ttaclpO/tpiTwI9uB6rZZyen1ZtitH8iteip0irENeTRDa7tKTitMY+QP
k4m86nE4CpGrzccK0AN9hQ26G9i632fYYnW5cyDLYRwBfYFqvjiBy7FAsQSMnt7Y
xSYqaUS/jWJ/UBS8a/j4CUFiPUC9LW6VvbaF1Ulv5SsCktogpkTfYDTfW5MPvrSE
raqFDzuI+QXxB5TUaU9bfplFP+md3LnKs4qHuGDFPG3VIdlW/NGtumE5cKvYQN1G
mFhITobERNa8Vw+AYvo0iIZO3KDl4Qrx1jO/oq3vuORNsqTooOqbFU0WMNwVr8gx
fkmdMY6qSTrWSkb2A4tZ2j4sDT5Uw4xdSIOLrH8HTW8ut7g5q8zwhHfkjgiyBvHi
lFw30FK/0LwPqF9I+Lx2Qp23DyBZlbFPqbp0la+kjYnYF+WxCoEbJQvULREiRi1d
7tNcZnw2OjzYnUMhr9DOiOsaoqPNSgKg07LuU259vMdU7e5Qu5d2Ka0CyNJeQSa7
jMNsle8NIX2TB/miTxRHDIHd4cotN6FT1/JKDhAcVkNRYz2piaZn0pOs4e0xn0VH
TmhIMJd60VaB+s1p3504tykegJuLF1ueR8W0LyPM0CdFcJwzTfH5z6ezHxbVaVzt
gZ7CJdU27xXN6nYZ04VV4fT7FtpVa24cZhxI5cW8unClPyIb7zbjkdqkXxp6I21H
D/eAH/Js4qIodnwuqzhM6hfEnb2tACKqdXc2qqQ9el/H5G7hHbwYhchcelfM3JNR
z71bACD0/YiwR0tzoBm5qzVjldzMaqfm/PW5T/7p2e08qg5b01ByRnvldNyCwr75
KPvUv+9X4ad8pMYQwbRiVfankxu/1ZYUYltnzMVpejQllmI8jbCPjSPymkxoA2NS
6i8NPEXZKWDA46EZw/8ZMY1EVh/yL/lhZp/yXYvRZukGajdckgdISYEDZVUjE/7A
k9FhwH2Eu3pK5xJlqwGypJb+jv/l1r9zMdB2Iu7gzDznAgWaJpmVr4fkXVAT5GUQ
02vMzRR2BN6dERi76aoFAJj3w++vChx7dGeymDAI+XMcRYSD6Ke3xqZQ1R/xI7tC
6EeZCsNhEvWBcPWvhLXuO29GsuqIF1iL8eNfeOO5JWjFMRg6WRdZyy2i680fwwWY
exAOAAFVWVutqAyjXkg0YlGL2aBbwVC0NuZMdrvKQ3EfQIJF/0A4/qupblMEQ9WB
LrBN2J+6gGCf1YKP8aMDpeVHlGU56SizBboVrfjxnaLmctP6Ajmy6rwhYljYAsJX
XmkQPAtK+pEf0L5OnJEwoojHbvZ5mnGq//gchGp4SQiirZGnnorqF3ccWjccXcbO
dM/PR3YNuH2gaUZuE1U399O/PxKe/0FXKyLiqGXCy1KDCvEVLHERurpxG1O6ol0Y
JaeyFBgOXgZ0ZsA2A14Yu0wgIb7MgruDAOjZpFXP7SjWtIFgHJrdhkNO3uBMqlrp
aCHANBQ27prjF8giXDeZwvtFaWH/lgmbPGdH6IwNYbnkH4ITdoviSFpRlZ4vaNdI
hgREKtU8HZBdf3lAy5WGVSOPAzhmpFSm6IC5kYZfO9/4Yz9xh8Dy39mw1r/KMgL+
Y1osx2FP6KjhR4/AzqenkM6Tt/hsgFMjJjI3WF4iC8qf/EVh152MPFlWhjNRKd1N
qXCkwWlQvRqeKKUmZvPv/+yUACuv+cTI3zTDjkd4j9L6vEa9bfVOPo8AH70iHEBt
Urb1GAuBXF6fQbft4p722hRKUO21A4RFjB5APnBBzoJh1rh2UvlJqztbj3/MyvYD
pJ+RWFLjIEudNlVMlc4FD06KaBQ94XqsfCbyka8Yxc1j5o+tFN2u7uNCXzDkqx1a
SxwQIc/benSn4GNjbzMUu9aoVJsap1DJQBtG78+Zf4kPKzcwl4E6nREH032o9U3v
pu2r/JmZr2DCw0ZYC9t2Lnxo4aqUU6lvbfVUUd5GarQ/syAqN9TdRT1d6tVdMHn2
TAu19ztXI52xMppZMpBY+4a/oIs1xW3jtwah7RxCmfq/jLdEH62SfonGm3kNOmt/
/HO1SQzq6mPpgPx9PelFqrSBmWQkxfIOpVeDWWNxdgyy0K2vN0qRRnToHl5NLhzO
vvFQK3S50ABFiQwT1P4U3D07uUOKS4UXMXx7AEhwhsuthHp3clfkxApFTsE1rpyP
EYZeTwmgpFfkFRk4STq6PA+fKsYgfpIS8loiPNjT6pirGl46iQCIgs8h//Kz755Q
a5ytnQk59Pv8QAvKmg5dwyx43ADj8OAqLIbNrpC/b/GfRhCWgZOGfSU8/q3Mvcy2
ylZQl2Gz9QLM0mY2w30fDMyW7mWOzJrSFENrRAS/e0apIwakF2HDjQLIsM9zfaCh
LYMoOhtkUHp3F03GSSGz+K51bleHtYtTmyGMIVoomXPRWZWA/EkhNXxReyedWfNn
g0qvOCQ5zZ3F0Nbq4ajgzO3m1y+dHLYaKYyqPPV8vwy2AMuAm7Acaj7h8MMi3Lcp
1Rw56XxccGFaaPri/Ia02phu+FEBsDV0FcOTjbOhR2edDZs1I7xJtN1j8Elt9qJl
N6TBuLjHD+L1gtYh/Z1SxCF8oXD/l5NIcpCyiTi+6vB1eNm0Exve8U9M0leD02VG
qZm5WnODsXBdUqmHnwXuC75m7054azcPHnfN/mLZHsaQO7c2xLYcQ52DqGcu9E3s
yGZHnkpciXoJNB+ft4vK9fgUykuzd+ew0EiApVp/G1AoGgeiIxwbh5iE47ef1SQy
4w5W33urK5F9dXplLYxlVyRRiIoCHXC/c+81UB2fvqK7yb6XOUqWdNhtEjnn95FV
c/FvN4pND1EyepZSCHJD560YAsUrfIYXGTh+yMuxGOVffr81Q9CyzZzxF86XNc7E
83eLy24r2dVC5TyXHwZxCPVi9igu9yUErjya5pxgkhUm4bor6rD0M+vyAUxALAjb
ZchiZA+ivFPXTceZ7lf6mvycd3rmo0r19Q2nfMZBsSMRu0Gw1N0/YerIbjJYACnJ
kLIzlI/N4x9We9ZowdEIKUMdVxMQN/59/fE5kvroR/rkc7/lqdQY4nfLjSOf8fAM
mamx3hOR6GnPO4BkiSEFRYbkHqiROUZK9GELBZ4grtlU0+rYtymc4Szzi1YlnKR3
NvWsP4bZFg7Nex5YKoe55XxXi9tT/6bo5/zhWfOVvGr/ursFn/BXbSDX4vc3UMq4
Qak3/evTweiv7G90NorOtVtpO37U+xXLnrCd0mJ8jl1IhoYzIf3/sDl6IDVunQ6p
tk39fyJKeLh5LoEFBjo4TKcTHNNuL9FB+XgSJFfmx1m5NC5n3g3pL2/GxqGV5Z5C
47Ix15Qt3hfZfm0Mrk3VbTCgVd7SUce64j9o94CgLgWGzpDAP8GWn2fLyIR2F13C
UhpdcU20wP+e2WVFBzPfht6pmZHFr0oc8Lc0pwRaMY0ogyqT7irF2A5myEZoGopB
CZeaI6pmyR7m07l5CKvNAZLXlolkKSzU1/Br5Fw4XBhtGzrafhb+Wkwbl5qarlSN
67USXs8tpvVazw5AVZ2WonxjtBLgY1EY80j4IS1p+11pqoQ7+AdQuMMHxz6w0BGT
sD0q4qJ/2/YQpyD6GveTGRWfvnvXZtZ+m32FMiWqcZ+1H+dd60zofDaowe6u0onI
rae1InH/LuVA+oTArHpcw+uywqjuLgdiQWSDsFkr/PBLgCzw91u7VWxgaZyPt/xo
KL5u2vu5iDePMigh6L5ojyT5YKTgo9heLgiwVnuMNSJ/q8uWEBrhmi+EmiuxcOZj
TW1KWARUuZdR8sW64dXuPE61WxmgY2EEmhvTujM95pUVcip8d0lJB+AMhw8ILOBC
1iA9mRI9IDgGw5rFQfU2OSvKRt/Z11GD9y8qXi0W/faeEnSxhuB5nsAUn1jpOl61
qotjKcoR1p/bcjmsEKHUNmr2zoPvNYNZW8+5fWNeMXUOi4Xrsy6q2mTGNpRkV06D
QvBJuuCMTHLlaHT4ckWSdFZZRs0S7Fg4S+jZSYr9xSsg/79AopyUtivymM2GMzld
7MSSo7qngdZed8yP0o4xNwvsDTEDG3K9FyaiMN1U0c4Qt5647XaRqVrcyI/A/C0p
iQlEUWajh3U3lsanP3w/e1krGHnXpG4CQdE0q/l6OvCa019DXKR16Ref5Sd8o6u/
dKmGZG9nte7R/X9AMPkcdRDyuZYQrPd+g6URckq+jfGzaiU+FBToFCCuGYl732QM
gnEWU3SFcneUb2JcjOAuhI96ZnK8OY6+UhWxK8pjWwQtB6gXqV0kwPrFxYhZd9z8
sJ2GAKpBkJBEBVWpbqTtqL9daL6+Pc75THGQFYbB30nN+uzXlYMV4T/NYhBPpEKy
6VUR8WoAlJvPfgFyiynIe8JO2u6cJd66+c/pQvE1Nm3z7lvtVuJ95hCewaFQq5m+
ujTvP8/xWkieVj8bM3yIc6mubrKRZu41Yf/HIMGfbXhwy/nkhoxvNvLRx8SvzCei
NJ3Kx2aqix1EQ/Cw4ELET248uFwUgPBhmRd3zjMK0BdIC42JpvElWhmZThrasBWQ
bPwCxBTgkTu3uoGHsQ3malCZLw/2j98CUe5lihed+f5jrlynUUWSE+qRcB0grAAp
SQ+Iyinngv0/WS3d9VQqn0cnNScVv8q4GznMrfqeEOff65QIWcvZ3aafnIU/UFMb
5LE7QchXILhT6gUcIQWkOWfd4l22ChwKK+2fVl5IJ3Uf3NRqSp/8+ZrgLRRFpmra
MqbsriAMtkKahlrEUepLdmZi7qrWVpteqB/YaklQ37FVk9t4YkZID+oVigu5wsFU
TMPp5+gURMpH3o2yTKpEQEqTGhdxbgbrq8VUEHmpSRgL47Z82ZhsFWtvHuRUfJy5
opaW2QQ7XFVgliruTu1EJjXPstjO5ZkY8P/HQUIFm3kq74anrwBOeD4NGJC+Zrif
u/ka9FnlDrdKDjomJpH++GrvbbJXrJIJv8ZWp8rSWzyHty3mvaXP0Yxb7KKuS+mV
kFK8pK8k1aJ8lVhCEZlXb8lqPPnBHrULoHF09x/7d0EnR8B2QaA0Pf+DBzUvKw5K
Uu5CdJoCyrWrVPSGsglbijQOBLG2Cl/ZcHLWc9/nONAbCZxha17GKc1RU4Cf1sQ8
vY9Y+7Tm3Ow3d43z7wdVhdwCXkbwhWR6kU7F8wf4fKSqAutfmV+xBnNWX9d2PtdF
NJRJ0HgfUpS9yyOQvvI6FMycmSUsHIhBkF2m3qDumYjx8Rj+E+uD7+tF7HM8511C
Ztn9H29rc2AxqlGaYBxVziSmBDG19DVt9psUrxhwAxbV8IsO6SAqXGBo4ntY4LCy
aJ32apkqoSm+0GEZp6yuPPzzwuXX16Hz7S6zXk2XHQ5OjoFM74phGHJjYAY/ZDv7
3A5aqdlgI+ueePcPNjMNuwctt0MhIsE9wdVWd6RDYz9lNf6/PkVOXfv+oeKsnOfl
+F8lcHHwDgybw/bB/3w9UfYpUhVeV3u4dMBRr/fLeTY3vAhgY9ldlQOOlHWXfIHk
YYNowRRl+Fj4WnORh+4tJJUAdGuiFl5I1m/I1hBdXn17w32HzOxEO8V7nIuBQr9g
HvRDFF7jN2wIk2Fy+P94yvT+in51DQj+TVe1OhXc5g/liH+zYb/CCO8OKx9s4O4t
R1Vo/ZsurQI/6iY6yjix5s0nlqeJp+mt3QrCeshX5KefRwn4N2/NKIj+/EpdNeQD
8qRkbYKjSPF6gPBV83ODow1EZxO7IQM7RwqueYmaqFWMKlFEvh+k0Mc1fqWXy1T/
pB1NMAmtakkF/eLpZSTVw4dQXdSpow0ItJjajq/MdQjzzFS8a7OkEErjV4stPERt
7wEeGvvzhTvQBl/mC4xlc4GuU4LiLz+SlCdrEorRLF14u2aT/Kyt0Fr7GNnBhM2a
9/IkZ4K2jtnN7VM6rm5Yl+zi737U8AIkxfA/8R6iQJOJMuAkc3577MF7LU44N0ku
Q3o40yGyAZLPBjFoW85eEUXW7xqVse6BjfC1l9KXqfITVCVd8v4JyD/sdudONL3G
CerzcH8WVIznWANCvJ24QQmlTTZhQ9uen2mB7DSa9j/XrXdM91h+s8CImeQzULqf
0NKf91TUuafEGwXaMja+vc/iT3JP15iodcuMCIVjsrWXaklpKUBR6l4u8jEkTnrh
TVvsOUdP0AZ8kH6J4HTjsAYTxPbruw1UbwZhA3tX1pM+V4OfmN8Qrl4arKcBoUlp
hWqZdfCRCM22o+yo6WSl72P/LeOCSua/ydFQeBvPDD7eHyZi4Y89QAbzbc1r28HF
jmYfpH4mP1p06iD865OySQ2/J24X5bIzN8jixZdb20cF91GhmI45c13uQoADdPtN
HkocF1xyuTwsjfBuvnU6Tz5UZcjmwDEYWZLaTUUtksLmWAFT52tscUrVnJRKhk4E
GjnjAvdB7pl4D2y+Bbol1J4gfjTaMp8DTPDBq37XbnCcB4bV+GGTVyBdbtgPBnXm
tI5BXbEyXS0iYLK/HMxi1IU8vFviyWQ83nHpuTstvxuvQhw5Q6burFndmSpp3wro
XNg4FQDW0UQcgA/an4YeOl5aNyGjZjvRgwZiF+FqnwAM7dOYPF1e/rOqbt6buZ3c
Vd7vb7F7BhQhYXZiDbnSgUELHzfnHXPKKHYo5olre9Gk8Y410EInrnw6GBTZC8MF
ZXZuifWxc+OoGYP8IGRuLF3xKNdxd33c+eWSRbypD04qu87wYUvKYMuLXAZKMDSH
Qpr/+IiLkVtzTJ5zGiFfCMDdgml36G0UIxa/exheF6AJvGO6GZxu8u1bqk6lglb5
aNMrX5f0Jzuf3eyua2eqDX6U8Y5UkG6xRqGTWjigJApyn22CJyQHCrIizGlrN6hh
uETs9elAxl+YgTmVJHQn9ESgyGX6BZc79zSLSOZ06fzu5pWJZs3uCgtPo1FGdk3K
3Auh4pfeNttQavPxQc2nhvdsuZPO8K8ZoIj6i7ubcFdvTkt5mE1oRkfwf4Ol3zXy
HYpKDYkLcpp+JtXHZG9SzQG8yjXuVmU1wbaZcyETAJRMcsTiFeZLFXVf2yj7jd/U
omERJieUdCocuOpG+vZ/HjnCDW3kpl41HmGQiBaxtxrblOOIzY7ipso8VN5R7j8q
nDXkCLN+6hAq7/cKGTw+aN/WyYK0DXHCZboD1x0LASreIrXbbtJupfV7SjPUc4ZT
mLrX8W1B+r2rWkiuhwLsxDCJhwnN458C9ANXdVP9Lx4BdzhjQJ60yXyl7v1Y3NjJ
Jl6REsirzHLu0uQzFP+5YI8nUN8iX7oavXSVURX4I5CYmqaEzSgpidB6Y2RdyMHL
IStCSZj6h+DcNxXulfp3ms9QlpOQ6ZpVMVdiMf6BbjvcYvZ06a6PruRmytlMr458
y6/H/negrUEpx6woClXTxIUZfPEQ2KuwelIjrzYK64JmbqZrv2Yu+TBsLDnyiOxm
EGmVTbNH/iahz4pKb0e8WVDEAZ5xjdv2ZadFc4r+I6AiTCMXeh/wfW9ufZtIZP3Y
ELCeE03lQLyVvzFIuW140gpjDQjOS9gAzuo63MLL6e46netZa6wSgpwz8CNC+wpO
gXW4MGOAnXd4XuXxkTA7Dx4HE17zQusTT4CfWhtww2GQbfhGy4dVTbDQeN3NpBf2
xLWcxAb78AJgvF0r46URAyGNRaF051T7bl73kUZXz81ZQ8zZ3E3XdvPzvvjxgsPN
CbX4v+9JuAig2/Y5llsUHAtyUzqy9CdAAoO6Dn5QtC44y1SbeFBVcgvQgIXs8QUg
Jz9bi7VtvyyQT4//d7vJjfirftJVtanUV7DGmJpc2hBz0LaVb/s+rDcMVJ8H63cj
MSGlu90Dofr4ogCwKyVbgfzxGpgfWeL6juLa1V3q2QiMrpRxoC23ThXF01Q3Y56U
6VNF2Yqvv/1vGnwRmSYn4DApgYw3TF3FY+/EzM14Y/OloZvir4QEsiWJSc6JjyZA
cu6MC2oqTF/gNQQAcyhUxHBnIZJxfEWPoDHziWuF15pqonOds2PzJLHFJG5I8R1W
3vSDlCjWOdqpOnjMvajj1WuB9S9SsUOk22gmepFhKaicQ1skSsWdkQ1k4P2Lq6x+
ADY7+qcDSZKCF+XS26nS5X4m1uHFkKHRKyMNsmXZHdiFa/yNWwPW/KvfJENIGB+b
PEAF/VV3ypdLa/SuLG5WanN02t6PP4GmD+Y2qVIGVR5OgNa77MKWDEEIm6+Y7dr5
4p/7lcMo4Vtnjswmmzpl0VOdbDzaHW6Ni8F6Y/z6KWhr4PB8qN8UB74MQ5dJ+34/
ek+Ni7E9nXJZNzRwM5d+ks47PeUrKYQYt+OznW0Q4eawCUeP8TTWv96RP+MHsPvc
vzozrYT6RNdbMCX7NzD+HESTnM132NZtDiOVtppsnEOeAbVIpnAf3/l/CE2Ia/F1
4ID55M2tLjsCXq/JrWU8wfRYGFuvsXHHvftY9w+j2+NdZnRNr2Pxtyx6XmoxdXY3
EajwmAOsgExfbX6GwRKWLUhzk5leg7LRU1pPBdPkZ5jWK4vewEkGR1n4d/TaPCGi
ZdcEJkRVqlaQ9rPjEEgvVfDWG76HGUL7xU0nmm7+v6S009cTrNj/jhBWNKlF7eaV
GbFoVbtdzRa0qSWrfsdkKsQTSWum23r5Hau71xtb9XXjYCi8Vh1SWfqKv2AoacPZ
P+2wM3YppDuJ0j7yrnPrFRuylJHWmiL/hSnHQLXJwXj3NNN6OKRnuCznFTHMgV4/
rwNlVEYzkLOfr/IEQaarmJwkPhg2if7EEEhZT4fk2l47MESsh06bLsAlysgzv+AR
TIKAPazsuszmr6O19t63JcOzHhDdbYBOwrIKrIBMnmC2sFCQ3A4M9tqJdtOJOOaK
f+TCHweH7tS7uAhRZjyB9k/HxUsJw6pxAaXFNKIjmIUAqbEgzz+hrOLZ3Z8Wj8re
WbJxkLCAKYzUjBhi/vJs5PrsmHvN6P/Q3tD7j8JZGzDLwmpFpXyQYA0fW01Erhhm
FQ46hHhwEYSQF8SYM8NbJNyepHM814fdcQYxmO8bq9XqhutUxfSIYA6oiL4TspD8
UWfTrjG3ngvbOEsJZP4a44uXcCl+AqBwNL4heChwWwd4RggbK/6J6jM3R0ZQaajX
n7/rW3mnu3V8USCPMlP+3pIP0CihiROSXIBEXP4H/dTwm3IY/LrOQ0+B80A/TrQe
sk80SwNeEnINC7QIeaUHpV9qdN6lXrg3Nqa/AF448N7wOzkAfKqJvWNQ1xIH0EV2
X0mJvVEvfB8fIQhB3VWCBozwRXRXWVyRCgg4HesFWv89eTUI9v7oznxcfaoX6YJz
I1K44N9J7LtzdxsDac4h2uR8pfJSNd5HPV/PMRBFnj1m9+P4BdjzXxAoUQWJIGlL
mk1sHJ8H83W5kOYaghBZinL3kJdv7Ss8SNIMVkPRVxkutzj+2AYyZShiDpNsCVyb
fGoROf478BK0C3zIZwUEqh2YL6wSi6XvPRKYgpPhAfZb1dtTTGGHWDf0m/iRi1Y2
xCA4lVrJ+Yd9hpgUKesm2FRhD1HyD6spUdB+sOiimFDhm8Ims4bHjvRqyZlCZoBp
i5GTh66qcDOjTLOjvmy3q4zBvaKol/sQZF29Kz1RKpXAPhxRqjqwMw6C4aYQCvqv
MSQeZS78jZRpHspHYn3ofRkX2PXdDr8seJXtfIQPjwfHLFvx7ZHfVmSg7lFzZ6jK
NIkYI+8aji9Oe3SMzGi53yaSYo0btz/JBCVUGEqFK39F10gq3GOzNjVO2qG7ljpq
zWKvNhzDHvyWYQdYJs8c7GwUv2pSZ9fkUwcUK4syCeSeg68S2AjgTNYSmRtkITW1
PKd0PJHiBWF32jFEoiuNI98gjMLbd1tKUwqFjU06DJ5Yq0KCCgL1g900azRsRAlM
0hkTHgwGJsKmr6x/MmcQ5gZAUG1TK9aKqOEGqyV52oAOXL771VS/GYcOXZaHbOZY
pQDPuSX36eqUszKKYLvU2XYet//H6INvdzw7K/pAGRxofvAJEFkFz6AOz674LXUG
NbSoaq8xPYiS5JSiZ/hFROH1S817mCL1hUz8y5KDA4Ff0jASXryPPAgSrXeclpWl
i04QUWTyQsqPmORYXfygoKQZ+QMQsVPZTOid3Hdz5B4MhuIEcarHhQV+E647LpUd
dQN3am9xsCGIr13gF3ZLqIHJKhyEvj5sHS6zePBir5lAxWvGeNLtcJrGYRxArCrn
o16svM7sR6JC0QlqbU8D/3coYcvrnRL7cFIyk9j8nRv6E5W/Dk9Pr0VOgA9gulN0
ihxX4UIn6Et4dIezIqulII7xAYkK+1iGQ7udJlBweD+xkoJ2iqKtbmvEIPkukdST
qwrYVp71rCpFkN6gMAKrDsqC0ebJmYjGs4QhAGPfamiVDe0YxG76I03yOxK506HK
ghJCB+cW2pSYaOi7V9wWVHxoL5J/h+oVXd+2S0oakK1BrFe2zI7vJFS1HLqWI5CR
9QErwhJbHzAT2iude36EWNh8BUB/l1H4KdS7rnnpka5K/OxK5LAwJpIbbWE/VLsW
aWOWGqiK+ghoi5afEK420bx4pACbA/q8Lqrq2tQ3RfLSd188cLJBxABXqknBjjJG
DgY9GxBAQ/lopA2AAZGbdG4qNAkdPdb9vNktmsuEh3204+lX1gLj9IyaGmz2vZ6j
fbWjd8Sjzb+GYTZ61dHAkJSSqwU7iZRMJikyNvUvyIa4rNMVpIlIUs+A03DUxcNc
Y+F1tenUaV+M4idNh/K8G6MTT/xzBc1K/4hm1VQ5m2yS8iXn4S4k+IFBanHAUKZw
9lJyU9rxvMeLPf6a3bKiGq8r8sJmKZ+X7EdAM3pL0Qi19rrBraWRXWSD3tKUzMai
uuuLmz8geFypvtTv4eYq7tXPE3Z2JUiHdl8D01rSZfwouDcL/i1P72Z/HaFRY/8z
WSCPL4GQe8u0q62XdgSQeNb4Q7aNTQiD3ORayggutXYLeYriaw4vGCuFjUmt3wsA
i1s7znr2ZutUo4MKBb0mThbF1dVZieXd9kUtgjNIyRb9y90ZaOAeLNUsq/Zyds23
FyGaVJvrY5Mzbh66qkBKM2AL/XauGldd25vb95UngtSTdGlXoVc0NAOACacZPx/5
TTxmd75ky7p9eXKVlyHZyyuABkCYQvWzqWe7Oikg0gL3vEpL0bBOKGF76aX8TZe0
ohPJ5kN9IhY0Ukyq1Ce8R6gJ4Gb7IGWqtI4aUSRLPoro+lXxevohEYs8KFpDkmc5
WugBfzsrDRK7jQO2mVh7abO+WMs8U/WxgynC1ZfKhTFSj6GCCOpnGRkNqANKNcRK
0cS0Zs6XEBwDNwb3SEliQou3YNArZM/1KuHoGOkHos7IcBzB0BNiPl29S+fJ4mHI
v5MwDxAicW6uGu70ul1WWtfCJRTS7zUz0hFaogRSj/TEzes8n98FFjinRpW6rocf
dTnmBMOZzAjJ73i0uRs/cDD77KZF+exKvqr2hz6YNwoNG9kpGhaI0ZFneen50d/S
HdVimZf/MsD7kpsNze8xRulRC10LSf/5z6uhbzVCab/uaxvtG6d+SMTnO6NyyL4O
FuzFC3G+2eKzk8grePBxdcG+uOy8hs8eyxjmOkxoP1ChWToCFMhBnmFd261XCl3O
Nm0isvJsOqj9fUCSgL6Y9uM96rYpMZSDqYXGz1rxJRyGg9WZuKZI4wIelm8ldjZp
czLnm/ZmbFs/4KLm42I/WiTNvblDTEpCbHjm0YCAlzIyBJh/A2TB94w/EfsU/YPW
cXJnULxuzye1JeOaU0sBkJb7HSWWDbl6of5/PhawRp7dXvXVw0PHdR5LIgNJ8YkS
eCPBUZ6mjdKwJmS8BMmfABpc+Xy6oe8Pmk8vQF4fJ/iOdkNZIVmrA9kVzdU8Ysmk
ltI73xwJ2GJE1ssFTWAqlV9TC2blIF/Q2jyYByjGWjHOrUhXxnJXtf82FBg7v6Vn
jgpGpWr7Yp/0+3t5w/QkuPcYxMGbyFoZp0490UijUwSpRXRX/zRH5dGdLzYawhQy
jFLEHu5DXUhANf094Q4SKMmEq90pS0oT1nwZzj5B3IzKraMsaO4oIc18KUdLFRlo
L9JJPjOBew+E0lGI0Z6TqSgv4RHTOfZMz6yi4ncfpsME96VtSsKGHDEQ9HEC1Wkh
B3haKdQv1Kd28wJFCGt6MuwgaXbyx8eyEDK8n1/K0poa1XfQ+5FKTJrzh3dZhmFI
J9zclK8QN0rTm/+V0bks7pWFndNP+kjKUXkmw+oS7Q5hhx9jI2/nrUbVkbEvgSOO
LfJ6QazU9dmn0RUlNsd+FMLldlHoF9sm/p/alC9tTCRh2B2HYr7Uh3Q/WFv431Bi
mbh+Qrkk3Isscb018rsKNUwrp5gqFr6K65yTvR4SeRpLRUlqQ5oajOIIKmBTJuc0
vlEShuTo45hDIKUdwX/85Qihcz0K1Oxz/f51TZZZehug5pjVENNmYt2A1uLK+Bzm
cWvHbpGSxHoFwJMLiVWlQMA0Q1mpqp/E14gokcqTRpItwxWc/nwSOlh3JB1sswFO
gk2GsnmGzaogh7OVufkw9WIYYHM3qfMyyflhEMOlDMqdP96O9i6u8j0uZEAYzUlg
ptbsa4JpognDBU6OSc4ciNz8vkKo62U4FoMoVeJP2zxTt+lqF79GclF9v5CPQJ/l
Eqd4slhP3hIIKVREbgI4JtgQeoZIQkQ28JqWW55vFbw6ND9BefSW7QaYFk9E9YSt
P1Q18hR/jmFmg7zXYXOubA==
`protect END_PROTECTED
