`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJ5l+tWFAHqEcaCMQPf8n2h3GZL76X12GZBkvRM6fToIH7mbSloKhTJYtBaAf+Xc
t/yDyvEe4KI4wAKK8BwKEpcE38C5a+6M4n+foSOxThlOT49GFj59zC5UozxJbTNk
aQhdqfYZc2xB5nOZjLNFckta2D56TjGxgGcaWE3uHldHw3pYniq6WPR9sWgA6VC9
qj+vYpYUepabEKAx6gEMOyUyZwTJnOXHOkBjZYO3nu6TspOIpUICrBdgqmvliOku
QZgRVtqk/sRTUB4HCICEVjKRm12KrV3g6blhsB5ce7tCVkLMArN2I0EVK80YBP+s
NYED9bEo27oV/YkaLw2w626x3ddovBR/g2PKD5cIuWJIky+oVpWaV9MZ4rlNc+A+
WtMFVIMPExLyD8Ye6Q8ZDzTwiw59irSaIVhwirv96Hm+ATgarHo9/g87qcmvaBJf
wU46QBPpU3zBwWYqQZr5BfZ1dVosWYzjp71PKGpwzUat6qN4Yj+o6L6wH0SabxLp
bfXQr123qHjpaKcNe6CD9fplcruEGj4UN3GotzWu24jzldOPRBlLLC0qZmruoi8Y
MRYSafCjS8PVXEgB12ElZbHz1bFkbM8+5P2WZIegooJbBMH3e+sYRRZVcjHoukvI
raR2JYQbrBTJQ6mhZ7PfkduUgSJnEdFoynaGuAU1oeO1Ujp/WwaLC9dzCmtFVd6M
kgxJYJ4YL92KD2f1uAbivwVpbeO5ZvEgsJvJ7jEu1W6EJRQDex3Ic9ummUIWXmeH
VBoDXuTlZeRZEEvnT7xeRhNVqYrWFzf4a55Zrb5mv1/s0LhU4Dx1Rg4PGIZoniSU
psK1MQZmqgEYQl/pVhePQVtDEdkGKk1fmR9cVHEAJFbVzcxQNfirQdUWgaLCYZ7k
/awJVaKZvtv1C8LKBvENB4+6mVM7GgC7kg3vWTmRTBoy0u0Vj4/W17piVFpw7aV1
i+gMWsEsCsTSY/EpUEWEaaR6/IAFYx9A/4sbpa6VUuNUPaN0jnay6ETxYjx4uDDR
mhx4TEL5ox1Egtahia62cz5q9IWJ/nrHv3alC/pBsoHZk2rcDMDjxWIdaMj08kvq
had1W/umEbbFU/DKqwGinqXjrr31KFdItAyAwRQ/E7C8mOguZizHdyIsutwv/70R
kn5xzuE1e7sPhFN6YumJHE8LhqNPmg8jp5z4IqH9bHNMLKmVEpE91+7VZFwFmRnF
QoPNlqnKxSLmIypC/el8q/sjX6GJvJwxWYKEyESrboSvDYLgBSdWJPB01fg5PgDW
xsgIRBANQb7btNRVENGXXikmL3kKJyVkbO1H8TQS0xn6cpmV9Rs/1QjhfNyItDLc
ItY6MyO2GDeNMeHsh2RBaaf28e83fstMQIthF1uWMG9dk0VZS8/Zm4+mz/UoxFif
hyuag06RBWigxjZNduIWWRkgA7F4mGulLaWb7rrcW77VeYrET7Ru4/DrnWjyftO/
E+NSFvm2B9dHVhq1B/g+x8qKJAogj+hf4MhAMc3k6vYv6863bcyyIq6TPkoen78g
cn8INDuFrcYDo87uMqURCLoBMxCuk3dVjYN363K99cH3g13JiZiFzKX0ayColwJ+
fik5VfdwuEvRGtHEn7KrpJHts+80o4x0hiyq0Th4n5n4P5ug3ytqAtJotor+gFdy
+IPio0HkZ2F6/+pJMCb+DV/7Oj4QcI4q/zHQWQsf01wLDfgf1ztrdGASOv4L6gOC
r/lPCnKsG3ZDtHS+lM6Blwaaz8jbjCQjpeDT6GTQmsDianx0Pvw7B05lCmdTqWkp
2K8Ihb9Apwm+nWCWD3BwA3hqze1y8DYlXd0P/r5aq+U+M4pvo/mFDSV//oCStx4N
7DbqWUm+Nu0XqUcZNJcpeVoC+Lyion/bjjrd4Tjr8/E/BVWdwrv/WFAoUK+lD/MZ
YPWuWspt5sqaU3LO4uvkkvmsEQ06iHGdmSW1bFvTploV25A6/umNlc1WXf9NET2u
G6NMb1jJl3VNpcGaQb8YAkib6IIBxtU14EXhj4OCNkr/WJM4pD5xyeOHSDs8sHPb
2ZDryXVNLmS2XxoeoQwK6CYReUmiiD7KZXrWSAC0tVKsOr+ptU6o6+Ry+QcXlMn+
H5D+W0gCDTUxqMCMHZQpUS2bVCxwHXgx78L8yddb3o8OYpbgqiQzrTg19fcyQQbH
QmhN5bbnyo083/WsNynxQWoxAeRN8TIY4nCa+LmJQaOqrcmOc7PKc7SxahpG3Xlu
4cHP7itfVaYUoFWp1zkSm6qG3J7eUydCdHruoarZGEBb/LhAvVtk0aA4L2QGjO7n
8NO0a+qadauaOYdjzZyZ6+Tl1StPcULYa4W+Dh7TjcwMnfXflojdm6+iBy8lTFHd
vL7RtTdnXlHCV2BR01506XAFqua+LU621cBj1x7EuQ97rhP23EhrWaX8ZwSQFo+K
esLj5EWe28gVFFXZioWXJ0QFU3bzZzvtqcZE8sTHRUAJ1yj3MJ7Vqsq7w0Uopmea
Ze1xj/dqxyA+2nLbFGtGz8knatfFFi3sOHXKfpEQeLbAyxNBS1t0cHt1O/TkSwDS
TakmGqhFL55x4l6pGe6VXr9kh7fKXV9ecaqU6E+BBPFUSbSywEj56Vk/k6CMQ1BF
WbfqHsk5zS5rnd8wsYR61wWu84CwYsPyBSTp9BcUNQmXmTnQR8ppS7oIn6jscHgC
B63uqJR6u+grX29pL0NzBskyPdLmmEX5rsLfVontMBEHBPFD8ctE6Ah7zlwsazsj
/UjwkWJ6qyv0Pa8ybcPxINoS6jvtlyecVqg2tOvSiVSHoLsR4LQLNqNlugT2Ncdi
/YUScShfaRC9f37aRBTssIC4TtooZESXgv+dc5X9aeoSOPEKT0MUfbjVr7AHNphk
xBwTIlY6GHGC4GPkkm+KIHVDXyQIpOOKak740EreJqnFu+mk+gf/uC9onJGcy+QG
lroCFc9Ao3ep2jRqmXR5tDTsnZO18Y0/V25IB0MVQwk7hiSyMT2bTqFLPxArXKX7
4Cwqxl8/jTkHImMUGGuQsFVpTWhU+pLcFIAhU1Pertpf4RlzSsWI+hGlxm/+XXhx
FuuuvgR3w4BlilOpuFfbjdW0fjXQ84vKFVTohAEYc6sP3B/QI0yA0+b0Ai4zeHFY
frVF+uT2KGKK9ywCpXPxt5zspxbqoPIR3JpEIfPcp16CX1DlMVol3HNmtmRs9P46
YzkyCQ2Bw/ocJoVdVznWlOcR6eg7wsqnpeWSkvJc2BsPE30fSqTrZN2uQCEy0wo3
1b1E0EsQYG2rCZk2HmaiPqvOi+zz5idCWw/ljUl27VraSMVLy0m269Zqg6qqazqz
JxUviSOFMujJJlqjf+PNa6tCGMGyAa22/ude9h+YlY/e+jl9EBtwpSJjL/QhFGFC
79Vt/QCQ4oWfmasO9cZL0bNj0T734mYWUj0F9tyYUF+OmbKZdhtFSW3hFzEdfy1A
DDc/VYaLZUpm/PPZt/m7yPBRCeQZN4yzXmz2A4Udmkr3ZhAUQcXHwwCLNj2Q+M76
`protect END_PROTECTED
