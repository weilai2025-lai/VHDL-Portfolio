`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLQUZkN3XYzrBWJ+FL91wF5lP2EubX0BUu8OIpeH7EdHjSPwDKn8LoIZw98lw4eT
D7RZYPQlBQ5XV/ZJYxJASj5hWZdz1ApmLLmh/guuHRsMEUXynUjAqd+W7cUoa7LJ
AQIvicyti4E+2MZg5jtkmHqz6jbVL5mwogTYNoUSFhNbidYtkogBs58S6XH7pod2
WgtSfGjy2H/zHW5XGreNZDc1sg+zozZMv6KPAxQRS+DPz3+cPTRUvbhHZIhYN2mn
G3Mi1RMtKsw9Rp5Bbh2tBZpqYGry4sNAEMr/rB9j3QROA/WdDKRqUGuSfWIjN1Ic
8thD1A/yLXp3qx8HKhIeSZTdwZSptMzx2bInYXNiZKQ6smVPCjBTtwoBX5ZqiED0
1uBpsH467U1PB4+N+NqkIiO7GrGSsbnRvRN9HvH0B3Jg5+I5GZyWY6qzqac0VENb
vMEzNEHttCneIbuK+rsrNh87ls4naiqdjT5uhfdqMZ9NSnJMtxcbw2CPfhfIDhJC
XUgSHPcdNiPpZ5wxDUjWQ871/r50aylqlc3M27I+Re+hv/+yjrVdfkyYxXQtFbwG
n/UIKxpoglO6ksJOHHkf019RbAr9Sg4isUTVwYscRqYRR2sX/GaNPEIiKoCP2s4v
MtmmEcRqfeNgHriqmaJS95lUcoXR/Bi3mrf12vg1HvcIKbDXXBQ4sRNo13JpSp19
8EfLsqFbLaXNj555cGksUmjBtuE+gt+fdNwPdR8kCMMMBft2dgejq7uIj0NNHjme
NMCn4i/3BD9iL+PznUdNtaX0HOCwyw3GhEZLRyZrEKtj5VSGTj/mckGsK05QmYYv
Q87q2Dh50FitowAVtlCWZg52GH3M36oXJ2CsiU9uxtYbnV3zLoYZ4bjvWaY+nAMr
OS9Ic6amCoyTcTiqU2j19BpZZGwUSAD2Bl84AeL/640NvI2qYe6DR+al3TmlCiiO
73VkmtISEeuktoEv0SCYeNtKAdDLwt8uEfVLVDOsSONhEQ1Zs5JIwDoBj4gJVhoZ
sZGue8Kih340+zf/SzWxo5tAe2eVdsJLHNLDuYCbHDiU2XiK+zETez8ateBFw8SK
wxIb7g08Dl4doLUUDgMpTMKM49SIyRjtPR4s/6aCyfFK+yc+GFRcsstPL7zC2dt0
cN5OkrK1k0qS+k0ibSIoMXX4aFTC5VuHucLpMfsvRsUlx4AicQ7hZvB9B9D8rJuL
Zu5jXjPqiC6v9I5jUMIabgnTwEeI2JtsJYepHhE0Hvp+3pUz5ufu4UB+TzYO1Shc
7jx9zE6ibz3btl7XxsB01bt764NODh5ohGWo7/V27HNsIrmdqpxUq1qF3J19T4Ta
JUwIbQoYomFRgW/kR3zuPjwe9kCp4INUv9PXl09FviLJSMBe9vvTkD0sfZcaa8+Q
VoFQIIkmT1HeM2ngx3IOkzSuH3S4AgBa3Zesj1Au7wa5CcNXy9V+oNQr7A1zNslu
aQzjQeP5neNWNg45ASN5p3PAZOXRLU0ss7k6hRgCBFrACxTtq8Zjcls/Y3kOVC6O
92LLjPrJ8ZT8MaD82bAamnAgIauLWWLfr04zd0IOcKJuiN2WU31c4BaLrMzYOXof
Slvp4wPbs3zx1QkYjaWN64XOqKOe/2agnqF0NuHagTW+c62wLDEMONwseu65ZnGV
ruekNAN4EXZ83N8LpPqQdasVHZcGiO8iZ+/VGOabhjTt8KifsEkADsg1IYANci8E
xues33dc86tSbkFanDJmncls4Dl4WaPrnf61imhMrraTBqPqqRmdystyGr34Tysb
NFKcBBKyIvB8E3yWFjO8geyxk8WAgDGL6nkF6daV7H2ezsP0xYYNXY8+lt0aWDaZ
dLaFyDBAUt7njQGx87a283CIVGTIWHSZQtPQsF0tKN8z/IuejkTHzG1FnszzPogm
KA7sTZPsiV95PB9ABZn/EVmDU8tyKJmpZNG4cdjB6BrdXmJQ1xH+swq2dBwv2UzB
YoGy+Kgz6nh9kniYSxAc8dL5wvW86oJrImg35ayUijibWMrvBARZKfzGN72y/VGR
Rsof0FzNL8EAL6Qd19NiiA==
`protect END_PROTECTED
