`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fo3yFhsbBzecVnRG6HUglr42z40qsWsuhRf09HlYSHFgOhvQm/Kv7I3UfX+z8/Ne
sxqOXSwDCSLm3pgADJjcCR1Mua6FQ9skNxJNPueWGIdTd6cWNyxvZ0xgIlJ916pP
poHabyIcrjv2sLNV5C4AiZpwMIyW/hN1NQAQP7bQu9h6DzWz1TffTjRNLn27XNbK
TWzFbDt3UI7VYxF60OnTefncVEaabZoBMww0s8uTU+ocsEoLwU4DZwpnxOzgiQ/R
s6qjyBsGPN5KBv3v/4CCI1Nc5LtHyrlKBg18DRswDKYBFnpfu5Qw70duXXvNoptm
/rj7Ml5xLeB9osascQDYJawTUUgoBJw5sQZ1I/KKS4MOIVC8cgxgIvYRC4yi0ln8
Pvo3QTNHeqIiMLznojX9mg==
`protect END_PROTECTED
