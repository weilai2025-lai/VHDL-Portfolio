library verilog;
use verilog.vl_types.all;
entity multiply_4bit_vlg_vec_tst is
end multiply_4bit_vlg_vec_tst;
