`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MNWE1wAq5h3OchCN3q4kWs+jNmZTxzvowIlFROKnWYMCpRlXuCuTjey5KDtSOLQ
9v8po97ziYrb0v2dBF9oI2J6OOZjZWtKNl0gmdaw94kXjCSfrKkW0EubUBxBRf+m
hTq4h2sUw5NVekAwKuq5X5rJefFvyVx0DEl6vssCjGgivosL7lolJtjiXLvnOYSU
GPy7pAVauz8hFyxgr0LuK/sgc9xrxKCGoRNQI7ZVSp8CZqN5+wdlHUJPHiwC/sqD
864CVKR0OyOwMfxNJyfBg7QORjD+F5L0eIX9ma7PnR1KDhbQrDxfaLtCDh1/V/6V
bYTzsuvvft/UlAcrjL0ZEhXQEPaN4w5yfbwUA+BELwYfzM0n/gChpdWLlJVG2TDQ
S6QKgd/9Ebm+38EIy2B/EKnYJGllIxt3Sctu2gz6JB8T8N4AJyPl+8B2npz/aYAW
Q1U5ZzALbX+7ndZ/SoNHnt4pjqOlHYPizTjg/wvq7q1xBo2CJs/zelR94A3qs5eb
0CV93p6WAoy/gU9DjA4HumSQssop+twt/zDlddCGqnWhaKniwCQPMlUiRKo4jb9E
+yIAh+pEltgHQgdDOFeh2e1THJYi+26EuwyW90W9NHp7rl4QdgTlnXPlS1FMUTm4
w+JY9nEPX3KooiX9jiSy81NGpBdolcW6es8nl6f0QD8j1/S/TFTtHlEOt2PcRv/M
dBOwmHACJoNl1WzRVV+P4eTg4egXAOteA4zM4CG7JQ/5O1cP0Vfbe+BrDsV69JMT
BirlPcDa1ee9AWSzDfpB8rC1fkaofDxbQAn7fHTb5RxO0gAf7pInuDp4vDlKZDoY
wtHXblPdXFOXai9U58lTHKKkAWa0TK9yLSAmIwCaDHYSV1LwyPI2Ur/UnB8dlOec
YEwSON06oKJFf0bXhp7MFs7YKAw77+06IcCdMHNWJf+vTql32RH1lzJutAeZhcfX
G4MWc4ejSflgqESN1N4GDCI3MaB5q3o2Ly79gXfUpKj/V5HxT/Dng2PYu93b0wSd
bw1N92k1KznNhK7tcKZOckJg2ZAw8B4JOGUggqnh6EqKtrLQ0UNot4KVhUNrAGpV
`protect END_PROTECTED
