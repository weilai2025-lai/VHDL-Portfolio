`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBWlxp2vG92gs1heGmEGwCaoQrebaEBeBgbUF4rSZcWMGxL6cukSCqM57ifGSEiU
a5c9ANNOzWn1mVIIA+mC7UY0tyboIiODdtHvIprVJpowzZV+cl7YqBdhvPB6Vfxr
tp1jrORmcV8+S9WhYXfGOFS8FXcI6H9zld8+ppLHE5wE5eSGEeGVe9mdXuXRgupz
ICqWrSvSNY1xMYf7/blcL48PLnQ/g6606CYp/OQvc9KjJpEg2m8VoFxsAI8NZCtp
tOzj72kR3B1/qK2iTB9Vd5DXkgenUsvg2rJW9HDPPqSlTG/Yn8BKX+PdPy7g/SW+
66EeT01uciURYJE4dg+gnWs2uFRRBtmai7TVTTUCTykJqBZge23PemDoEKAAUMFz
3SBVaVb119APGSj4qZLpygYTG1dalNGZU2qicICXAQR1Z/5k1zuxKaatYT/G4FFP
LLUb/x/5cXR8r7DK9Kr+QBNVQVUrLA1ZKpJ+bAtstdlOInKJoiy2vEIzQMaqnFSY
WBQD6lwgkRfFsUt/v0uT45Zn16h7u/V+wK1mI1v49RJh07/3sG59wvPlfS6NS6Td
bN8Sx18Hc+y66L0BdzjLlHWRusVg3FpebVk1j8bTU1ss389QhgsnBPLhd51bQ8ee
Ql+4eSOVYYxBFhbkdo5nRAA9iHaiW6Y/f3cb1wKuPvZPyPqWscyExtSfXo+0Dp+1
QIJ0PhvznxHqdP4jfuXGmLisRB+VFQdbFqY9+tIMRYQBptfAUYV9LLlnLzMzC5gK
UAlG2xFwvuODqEzgyQwGM7bohNXvkgscFho3+KKP8B1qzWBudvPxHOX/8ugwgXvP
kzzBtYl+sF/Gp03SNsWR0g==
`protect END_PROTECTED
