`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTtwM5JxLboqIumekBA7rmNXkG8fAj7KrfpvJINv7XKY7UnfPDpqv9l4hdvjPHtp
YThR2r4SSOc9LHM5dzKxSVItFW8YNKk0aL2YS/nEKKQeIg2qWyudtmen+im9xTDv
9aCSNDw1AhBC1dDFrF9Lyb2cSeG3CiPTuHIlx+yLTtHayH7l9SynjLslr8zvT2sY
QYBw+/0v6D6T5hoD1p8xHOJIjeeruMIBtkLjN1KIrSXK6Xya1n1aNyZt5OLbstsl
+DgDcfP9q8BTGxXdgB0DPO84zSt7xcQcdLCRT7VG2LI5Hea5PgjsFXdA/ES99Sjp
evljaWnG6n6k5YX0NAwpa8VX+Iz77G2Bm+FNxvGmQlMO4pY90221MV1mj1+ZGETF
xWLrwXvciNcBm8gkRSL6LGppxI8wZLMpMuanpwULcZ0Zrd5Z5c9OjGwM1tHlPEWA
yS/JtmvYUp762SnK9onsMKgo8y18eZuZxgi4ri7kggBhoM9Waswe2fKxVWpnKX/8
1m3YkFGyMqD1h0hudilOk2OFZN1r8SWEY9rmbD36m/Z6/BXEkcdkGoltjEOlVzH4
/yxmBjtNb1hz9BJ0K8gvX9MGGfc447HnnF57j3nyYKRfAW7Us7WmZuUq/VlED1Mj
NTy+MX+6mvIMtkc7HE9CoUk0ixn/INCd9KY96r3OUkFlRamZF51agLYOmuB0yB2k
3TSxhOa9SHiiDIyc/bZNswWljCxcXUc74h12voPEYR7od/OuTRRW6J30bwCny85z
1zvg69wSIXu1xLh8dOO6uoerOByfmL7F7QCEJSVN4/BUmfBVQ7K/QUPes+gQbMZg
5yvwM0fVHAnWnMYDEp/xDDoC21+p1TsQrEcwzifMuoHgDKOoe4LLA3IgHj/9WPTl
ZmMGESCSewTk24LIIqUq6Au9VE/fkX7BqyyuIi1fRMiPJUqnD3EK+henI2gliQz5
r4wYDNthB7f2ZMvMMcYNSObAMgOOhSAoPBERqu3p/OT7v8qjgJu/WU+HWRRArXs7
ijU58tCUfDJLFVLqgMU/9YC6LJX4UXP43ha/F3UqE2NnQ7zCUcHZrz3KaGh8P5X/
8uRGBnNozUkee/3Qn19BYhhcDl0rVS0pd9mrElxVYZfuYvn2sTVACDO2r6m7F/iY
/Ss1NNsbEAqyqQiJPsQRAHmNpVmrTPjcX6K4rMrPOPJCbKXig4pbRsHQHlNaazVr
dNqe2kd5LvEuxBzGtU3EhYY4rFtorcBoOI4xgSSQUb78M5FS+p5e8C9j12zZsqs7
m9ftT9DAek0CArIQgWEAIjfYh+ZYzPfikw1l5saht1N/Q6bjbp6XeZl42Fa3/rRj
9xIcgpuj2xG483SPtJ/l1xQ82UkIHUhSLv3zrzO5WSavSYxUacKU7XvJItVSznbN
YVj+GllhZZHNUnXjh7NOmCtuTDxJdYioFPtEGou5KD8dnCcRaORXdIxhMqWTT56E
BMlH2fBOc+x9lQUsXZuwBIsZxygPnaLFKjNvGOrFTeFI9sTDnLK3UdiB8K1cSuh2
8CCH44pbyU+3v4l6eCcnIfXPx236FWn/SkEcKNoDOpE4KOZubfa9PcL7y6VfPMNo
d6dagA5KzhvSaPS47mrd9Lf5T+RBvPwLJFd+ONJr7XZKFaCZ4aj+Z1qBy5efvKJP
Zk+dxf/FyJUU7ExjBBAKKhhjLCcAux094Ji9ZrlFBmTJy19Vidr3BFpoYPc3phnc
2QIoT4rQciJ+/SR6WTgtpD3K+hgbBJ4jA6f0thSiglTOUY1nH1QU05guTbGhGo4f
OG233sa+PNFZQUE03mlZ4d42efvp2OS3kLUKLuX+4YJrAMNngSvF9FCVQdVKqzJW
aUxXmxutYtJMw2mxqQR0A72Xrci1rbFvlstJ+did8PwajkJAFFKIyq0Tc503dmvq
uhkBhGsOky4kOaPX6UIYSqWC3a0ZCfrR9UyZjpU0KuzKiHdLoQu8+AbJzRMOsQ/c
5nXYzTcFH2JclsVJnwvsQlc87uSJl306nMtuN9RmBHOo7B/oZ6NVMwcF4sqETiQT
RnIoIiG3OJDb8q3963l96QonxQEuihogHPjSzkkLQD+iTEmjPpHGI+leLll+Y1bT
7bgwIZmr8nUUEUPvqmF81zCL8yY9GuOOeLBJRy3YG2DElML7a+d+ScPdr6XryKf8
yOJkMUYu1F7YgvV5r/KAqIIKfeTmlteXXeJxVKB8iLzIP7noRtCUB7A9dgioK0LM
2dTqHfp3MzqnfnxyFzqPdC1g4i+SjKdKWSoA/wbSVM6kdVhDjmvhlpXlNRineqDG
rstIm21asWxVpk5lubMhiKAI4ZvfBl892fXdg1WhJG1JbIOFRT9pMnHSCF6gJdPe
OKnWomAoUSBcsL1mDL5qy2G2q+AAZf1uBDTIlvmtnip5EjBHuGa6o9dcIj6tAGIZ
MqMz5Zlnz32DYBV+cVKzhXU4+izyIoWtte3JYZrK5UtxvjLtg5NyNaZuEyrOlQxD
npXquXAjBnRZoy1T4+vRuMnXfMIoh3y/IzXJjm8LIVvEFf25K75dSK3n1qxgM6or
QMSYhHAezV0s6tS8QeAKJsCJmSwRP2khklpxC+bHE3VKA0L7og7ZCiT39LSecQUb
pvFmo/vLEx558PWP7iwEB6KsZf7btEleRKohGOlfM4xOPEJ4SvF/G8bV2y/mbTgg
4nVa0I3FKVL+1/T/3fn1yL99FkzWbZVmBARRZ01bBJMPfKjAIwBrvL6p3UVpHAGl
Yk8eRz5e/WFJcrCg/1sRZSTmSCeEtTfWgAoUg4sFTLeWNJe2/4HBSENaBCfq9zmp
CEyy1leadklYT0ApsyCD9D84g7G5r2W4DCSZeZxYFIetifLJuhaD7w1Bi2lsOI3O
YvO4o32cfB0VA4tac4tvz7Ty0SGXe1Y+CaoI+52WGoUgB/8AXhBQWXdDnqjC6P6K
p32rGx/EXP/dn96VhD+Zfva7TWGUY5CU8l6tUJArCArW0gS6d+o8+5xUtpxb9Gh4
aOgwT6eYIXy9/HaOTwAdMy6mjZUUIpoJ6Jgv/jqSaHmd8hOOfV4xjNu+95Dt5pJS
+QOsCfhErV+pMPIz5jeWj689dDzP5dCJsufgl7Huow9UXDePKcPVAHGPUBPT96DJ
r4RMA9pVg/mPIdX/rdlkPZblBLLmzB48cO47lps/XLh5UB59VrEADP/bh91WGI7w
60YWOc6zh4Mm1x59tgb4V05tDLwAGmhkaKVSjARqGwxrLKRuYx9XVb8g8xn5C05J
x82dFq+6cS+/iWMmVvs/wO0xPlXUxg8KkJg7VdFdCM3opzsq3Cv4Y/lp1G0dhWA2
idxhu5iiXVMMncbiu/UcIAKY0dkmHu3xbTwV4tvOYOi9euTNX/tXYMmXQ40NF1Vu
zve7g1gBtn8jIbrSOD0f1u+WKjSIj7SR5hvCxDbt0l4EISCZHV0hgoX30UOK77Ah
bWyIvU25pS/HKzGRIfxGS8N9i9lH+GpjjiT8qcp/RXMhvZJYO5l/6EW2KMtAwn1H
nAiNIyUaulryv8bD1k8qz1yA/0APZJBP8/e8XKFCiSon0CkuZiEzFU4GLm4jM8/W
4e6VqAqTC+q8JA9oGxuNwj5vtboy8WIZQQN3oWAh4FNNIO29as0F+O5ObC3fwGNx
ug075eeDQeL8tQeBTcfWxWuNPSA5wL0Gw4KWKbs8jcCtDQ28DcQJf9fB2OtTpTJS
WhMPHOYp+hF9s3ueAQAdgL6vPiwGUEkMsUAwN+qqQeSSoBPh0bwR+wQnLz4N80ab
4wFDNS0eUERwKTWfr+PDW048N4S6HWpFqmrRvTbgHTvh37NFWhWtE0/jmnLz7epu
EgSyxxR4UKRGhxDeoiEuSBimP5Vk5ge9Q+aBw7aR+aqa2PpomOKfjGJ/iyMM1gq3
tpGwZRfVmd0w8NHhbXADyfQ4vltUpvK/JyvfxenIuym3YFxlsEvGVGVWzaTzqfFj
8zBVSy1Awp7xhYUSPgT+y24XpFAGLvablpsQXwN7huHG2qbDWGtNdZIYyrsNDxYa
BAgBgDfwpYfxPrW1pA7e9r6OpiAGpHqUVq5KMT+nf/q09Lng7VVBaP4v264Q43UX
LMDZshgqkOPCGMqMKAfpLqmwyDv9dm0qlqEhYRn8ifPovndZbNRqAefuKjDcuqcP
hisgMy+u7CkT8sz2g9bLapGopkhpeZ7NRRzH6OhVQtVNRbj4C1AleXdqhcJoLOxJ
sOdhgjGOMyDpYr1b5sqTQzNasT9NxR+gSZ7YUIAWcB1GS6XoI9F5F7z2rdPVgzhJ
ax3jZqmOpbFQ3DHabqPSga1efw3LnH8CF2GXD2ueZc60lOh8XkQRQqAYcNEf/bqF
3cRElGKj+7b8yf7FGIDS1OI4CsBhY0Lmdm1zBIVYMeAMVzueqXwDnaIGUB6he5km
jBilygc1HYyvKZHuqTIJ3QaER1deI0a3aJaTsuOTXuCxAC4Haol43g0x2YBcBOqG
qIwsoxn9K+9gm19Z5zqNSUY2qoL8xCeB5/b+uH73Ey07eOCPrVRXzwQDfHAMc9ef
Ec1W3Bnw/OJdc0RHz5jykvNtSRg1unH3aZHQsUY5KiOyQDi8J4POxmb1bMMWkdTQ
DjIBW7i7PsUJL3u4AAZWuC6qlicFXagtrAVVb2CQW8W7lr7A8173xc7/sMzSXNqA
DbPgNzqEjzwyGzRbCmjVU8dBi41GnUkySqAU2xdaJykn4QsaqewM6LrWbLF2Z8Cx
d0wKMvB7eVpwvBSYy6G+p9oGnXRUXG6FaEs0t6U0aSN/pgLTP0M/JG6t8IZhXwwS
EaPpCd4yfEKFErg/Iqimx1+3Rp0/DM12CQ1OOI7R2l4DahnJ6T8f9gNC+sF/vpb1
YdnrnSyjKksBb9xmwWfJZKOaTGIFNH8mtL5DCtYGHq5aAEAuQXwSN8ucXsIfBrWF
+DHGUR50R4I8DSrbOdc/jIfZdtVxLN2Iov1Udy4gtI2taT2xnJyU78XZOyPdwkKz
F/r5RKlVkNmPLOTZ9lBZ+520swZj15N7bsxWNzCW/mnmqMziSxEvmt4SZWLHHctK
hxa3eqq5IaGSE/5XI+sjSees3B+WAa/OMFzbGnxlN42eo/JolFP0hikqwvbKsgaG
nx7O/7LQHGZZtq5R+OgF606hwjydve0K+y3b6J7xYFaXgIXsasNdic+reqsrOqc8
vijukHE1NXx/hqTmhw0hMPodOZEjgevHZivmLd5TrVPU11jCzqFoQbiPx/OvG3c3
6HUXWFE8Wjhl8FocvQNfZ8dL67wKe+sZu/twvziYNFGfMYTdBi4BhviIsfq+kB+w
tS9rFFP+8XLs1iMP8h9JO9X5xOC1SNb6pYt+/Nwq/NPxSbGrmnZIR3ocPWdY3RC5
aiKTZT8UySTOhUVcjAgf+8BYO8NVeviYg8qXk+OxLILUNztCO5rVWs35MVyXxbiq
XASKIJvJma/+hGRzqg1n+a94UQ9gZDNKDrXtc1shrbaaGbOumgdp/pG/KFfEQsCY
5z3ZrkGTHPUxLdxYuzOgUD7fRai28dWTdOGsMqncCK3nj2P3NdeygfLtz96CEAER
rrt8H7FkltkqZc/T28lnOHNTC9kdf+laRpHv8+aTmRXDrMMwROU/O5Wonp+n5tcn
oqefz2gmvU51Nh70Is8LxWjMDYANk6QnxhEsCAXnjzcJEWSuWIgHdNPcpW+z2ofr
oYbP6SWO/F86gTisThkhRCJMTxehomU2Hwm2g8ha5lGzIHk6sRSSEbzfxMk4b7nU
GUUZEOZmACwjZkJJlBOd/XS+SHoJtcfGKiuZy7kFhU41Qk4tVpXwsaS/OolDyDY+
5Ujta9KjF04G6NzproVPVjEKathnA9YUU4kTQxaZXE/TO1LD0NCs9ujF8gmDlV5t
A9g3JP1a3rKuID04F3scwI8r/MjnK34oZSebrH94BEAwPULwdZ0WfonDo8A+Nz85
x9FpsrmTpATP+3Hhlwj/1gun3cOqcA+OAKm7wRjM0ekSpJtKIRYB/joFcyjzQxoF
DdWJWZFSMKlYzGeWRelflih0YS59EhD016IcHSaaKX2pS3bEa05kM7ZPh8y11eZo
IOZg96DafpS3NP08zJ42Vu2n8N3mQDweeEFR1QI8vefXMTogjtL4VDqlKe3BJzR+
4mNDtAx8/PaHFubBSOavnAU+k3a2f1JyGaJ2VAIJTv2DFwSrZYNrTyJM9dnSeEwu
1Fa+qeowlw76wR9iNZcccE3zIdeiayTCOUVSDoB83M4GlNWMaKcOEcqt35VsT7kQ
EVGbdElJ4GxDeZkzgaHEh50RPzZUv29UG3NxY+JZp2agoRNUb9dDtjfCTR1369Xq
8bJhZPSSIzXJ+RhFdoslW9mrDFih811K1ELCFRkfohb6xFvkw7bYnivaDivBXGZY
F5hJ7Ph/sfc/AzCM+DadxwlS++5Oeb8jyieu2GWZdoR4gsU/SQHu+vZqhMfBpG4Z
AWSv1dWm2d1IiL8PsT65/wmbhTC6yrj1k7BmSGn7YsQgsbEP3XYBYgmpL1IHLOJx
od30PwNYo/ull1maNIlZjg/l0EirYHibl2Rv/z4yuvjX7lGIsgJExcxbwEiJ3iUq
60fcWwuBkGxz+rNMW0OW/z/gXtW8stnV+lA0Us+jw6FugM7h2P8XNv611s57of9J
553D0LWc2GYdzrvB5HZpTrwuiXTt+moVBc0Mb9LWjW35wxWJx/ryYqVm8oTkEz9T
+ITaXdVBjDPxnaoNjGW5nu9wgo/eqnjd1C7s6yrmpQqY4ptdykxLyxE63TLT+t6J
kb4rBy2n5DtdDP8JqgV3vHYMV7Y9ZS/YP4QQpvYLT1VzV1X3T2K1n5Z/ONj1RLXw
A8owM8pciaPBLrm6GievG/BL7lOdQg7IJx/FcIBRKg0eVFnAPgIeOMTtOY9RjlzI
4gEjlQD7n0zbSf9AiOyIqauINpIffsU4pKlwLYn8nrXGqjiMeyWMkKq5maUdAk92
RMwQB0UCYqIrIKEu3Fqnw+GP10w8CmCcuDHJlIHH+IydhJPYe9GBZjSbv0MqSAf1
EtQ+h3FIokRunejHQmny+Ke8FG4ptRw9i020g5DsWFY3KsR27ykWz0AGvDM5tp0v
pY2f3PH6tApUgOUh5vjQRqQqFFLuvSTr1hXE/eRZ8EL02KFHP8PuvavqJQ3aZC4y
w4vd+BbyD8d1sNirU7zwP4hzcdJp5QxoL5hIyf/zG4bWZ5J7scuGOnRChsIhMDux
jp05Iga0zz01l635sqRGvIRHgucYuCY/vFT/7ciwGlOkUPEOTTAUaxbQNwFKfhk6
X+QjgPW6j0G5F324vNnnAiagCwe8HQkLfM23Gltdg8xXz6g405qjxli7yodcS7Z5
CkSOVhPD8SxcrMX4kr+MDkmDU8igLuRkcWIU/5luGCX8Z6RuhPN1Rsr+QiDbMwe+
fWxUNreHpe+8dt9WQo2xjnojcQsWfmR5jJ2Wo0s0kJP2nYZ9wZpRXaiIX2kZCjfz
G2Ghk7OCFOEVHfgmeVkMIg4pVNjpCvbLMpdA4KuchlR990WJujrYe34a0wqVwiK/
2hNd5gqCfmIGgAdZ0/5nxuBDy/gQifSVHJuXNUfy1cTUDyE8b8xzDxI6xcFDMKrA
5i1LUM1pFtJ9bfMsTSh5xHMpVbAQIymhH5Dm1XLdG5rjUC/4Lie9HYBIiP4R626p
ObyeWya5n4qJrJDZvB4xGAdnSG7Tf68LK5XlO5RF+n1fCE1nSjyibUzNB0358H6x
a4tbSZqIpuXn+aKe2vFUW4GC0duMzEKTCrKCZQM41qdu+dIHBu0+Bb3557i4pXJ/
sYnnGJPta++9q1AMQJF3jmzBM2m1yjiv0cpwFzDbek+jpblX3y+JmIDtcMzQwp+G
PCTH6e1nSOzxzX10NtQkMNvLqKDbKV3yYTFCIRJM0AAl6Ey6TMj+4udlqkR37WGZ
kAETXUeX3mAsSf2Q4/cYQBYR3+MPZxw7JPRzwmdBre7Y2pDzkDkKhRFxZJ5KJagI
Hxd6Hi0owqoxT71X64IqAkRpmIHBWo8Ga01MhWbdbRfpgXdHd2Gw74V0vE7zxKcr
+HSYY9Zh2EI9TzACZ8lWE+T2ae5ZPWP/iQyymQWGGwzvQj8ZKy3qEqzSf5rVCuPp
E1wyHNxsJAlREhfRKBM8h9zjWeJoscD9JQe24+87s3KRVvln6R3JAoIL3umecqKU
rQXH3RxlRLOGNcmGUtfsXDc0ahQ4tlmndxOLkuHNtOQbOv/Pc61+Gn8ZowSvxAZU
FiXcYmWqcYbRptyXSOgji+onkFa25rl7EVqwpj7K3Gx+XYu72tRABV7tW9/I0ST+
BOWRzM63Vuc0/bRFcnb3R/Ii3SyL15/BzZ+IEE5M32FaOvjBQRIuwqF5aVGOX19h
qQwhTnRX4SxXOWAZ7ObBCCj2EKXh3+IQB7aj+lAb/AFlWXEGqm1jIpetr43N68ea
iEvLa4EmorviPFLUM24httEJUTUWQ+t/zwTfrs49w1f19bXxH/oA2HzRQOPUvbq3
sKAHhtGw06/fcjbynXYgTnE2p5/dqgAY7PeKmT9ys0b2Q8uc/NrBme01lUf1/O7M
LA47rdOaEfBSVOtTQhVRnOc1Gal8Vn+AlhLRHZqxGvwib30tpKfw43EV9JIH5Wjz
CQBqGvyI1IuXdIDUuj8l982W/Jgu7E+wZwMg4o75Kj/+dmN2uy928+OsK69J/EMm
Yk/seDkxkVSptMETGaaiY3ln7Rr31m/4Vj+f8eC5aJNUrDh/yXXJ5MyUTk3a3QC3
eViNK7oJFz60+9lmsvUOxaMwbBFlc92xXB7rCNVRBFiuUoVSQIzeuo03fHx8/bMJ
VoCyCBEZnTVJvMkkYt12qgetWm7r6JISSrhQwEQdWwVdeAm3xqUZBQ9afF5oG/24
gpyPFz+Ulw6SquImyr7kqFAe4i86Ia/qqzYDz7Z4lEFMW2pMVq4UhFfjT7JVJXym
AQm54iJBUjIsdOz9LPIHmmIFZlNGxyZ7+pnVM+gPXvaze+d1vdJh357oOd4iyqdP
TjPmlzLynHgJhBQAuyWZcbb2RyKJP3xp4vBJLT3GUSLRkzH84yAqriega/JHpVJY
J8ALreQgS9ynJicwjU0je7QXLb7GoEqDT3PAZ4J9Baz/qKxOH55W58K1uemMe4nY
M5CLso1dnG9KuQsDzsPMJ0d62g7kLoTgGuuQtTM6+ULaUwDgPAggDGJCGjzsvw50
ONUW33ZlQKm90In4bVm3KDM+LAJBqjWSJP2GNi5ZjLGlwaqML0fnvjU0kYcNDB01
C4UUZS6BpiBVeo+N54EKIniTUeKoqlEcgzi0Reh4ubgGwJKVzgJhAe9lpf7XKB8Z
3gvtRRbAdItcZkUClLLc1Bn0m4hhFgGFrIynKxBbKIWbn9wY9MELqpWQcCH7c33d
CujLTE2DFsQyVm1h24jVI830UA5ZCt1lQe0EhIDZ8eMWACgGjUgWNHNhVq1PbFPW
JIzQ+ZmBa+DWSWv7mid61HRgUjofMNhiYO5sFfBvh5mDRL1cS5FqQVGyDpc4CcVB
AgBwLEyiJGO5HpfMhJoBm5e7nA97RyN04lFeC5aZ3fGYNRxJ+Rjn8xlVYPa1amVX
hWPgdSptTeH1GD3X/ErX/scpnXjrx5mjAAvWKHn+F75bHpbrCoq3fGOAS29IXBbS
08vKs9gAedYiciYcLcG30/H8hBMDXumcxxnq0nndJxXBpHCDPQycXTqnlnxgsvH9
3qAoGx8a3og/mq1tJFPJcT+uTQm1+peLhvoNVkgJLvJGtgk//yTH/P7QUlWfkZAE
T6rt0GX48Hiz5rmlg7mo4NIaqFPgu7lvH/61Pyd70zceZd0ybv1maI751R6+YYrC
gEBhAmuTxGoY4xfQ393AVmizfycz02Q56s9WtVsmC4FrSc4kaAL1+djBxqW6egGY
VtwmP7io+q4zppsQN5vFfcvCltZtUzB1Z3bbSk+uc1vndube0p3ZgUkoS8IHrYyL
CGPpFiVt7TfyUYeSMLV48x1CjFfpJN0VhBTGQlGbqgMX6Q0Ein1+rqGu67ECQGAn
FWoGyM61Z0Sb0IJi/ZQj0Ww1NnVgpYMS1Rv9ZKCNchg2qDmy363gcEVl/EwCARzi
jlSOBXGwKSe2RzgIC5cruN2fsmfYaz2Ts+/B7eITkLVdtYGeQ4vrcxNG+9pQdpwZ
h26TCwz42Pw2ntX9bVb4iu/EQ7lEmmTIvgAE37rkxPwncTyIBYy0fhA1JM983v6z
+k9Aqh2K9V3A8Scwtu6UiKZJgChaQTXhreezpXIVUsKsPObZsycEuwlLnBM/zdjw
UURloIIztoAf1Kl3fJqkz9MzGBfCdhe4HGkIeZcZPdpyiNaF1KSdzm8dGaoNkuLf
WNsnA+j/GeijBOUOE1WmrHSpJeMsXfKwYxtSXkNe0LIsR4fhyOX65RuAFE52R4fU
8RJ2+E9mQrJMzOwl/yHqZStOxSi5GybMGrLKlilRdVgx0N+x7OzfZ7AQXyyvm3cI
MYkFqFgkSZ5VuFkIc0lCh/4PsA01xcO1bfLvFr51L8CvFN8ZuGcJ0woSwg22IUBQ
+DQ6hWOlpFy+JG55FNY6do47nON9ADgUNahEHQguXDTQSWjvr1xH4O4RYJiIdFyj
hz+xvwb9gwGqNJ+h/UufAf6Dzoeb/i1Qng2nD35PiA9MTuf9x4sLY1md0ti8GS//
Mnlz2ZRDN1PZVsZrSLDEMctzy1YbwURrhnLK7UOJYkUJFn6V52iUt5nRnJg5fzMn
gw7g7rtc4WbVuubHfSFueihGbD7f3D9kqo1Wafd7ACvaIDltyRO0mAIAw5jr7+md
sMyQGFodYuJOjp/6VIh2P22XIdyigtyOLl8h7rny8JwRCkCiHSHBVjCOT0PxmxeL
mzSBDf7dgaZCjhBnlTSkQ/NyL+owHhUEPk8K042HhdRblYXBMLb3RRfsm0A67vKU
PXUlHiGS755jlZN5cUW2fl3wkGpKtfODYQ/Jrl+FV0qOc/lox5/cVx1LGFoeiSV5
/09ZHy0eA8f0/S8kNUJVN+V0Q0oi4wvUQMNwhtZ3b6MitB8oY3SBdZlFAl4xY3Hh
ivlAN58dmh1UxjL2/xq0LFv35EC8D5Lb+9YQ5yHuEmApcBgCPw5mwjYlutt+BlU1
lFOeIhDdZK3f3xxg8ps9hcd50U5VMqTAS+4ZUcABzDwLTt9y+T9OiOJQ7np4KC9P
Kb8KmDhYwjhCH12EJd6vncVMeqiQFIv7cJQoVGxWlA7asx+fu7GAe/WYSpBMhyWu
dvCZdIFad3Z5f8NiRIl2XtfwsMa6v4ehtHGIKQcoxqJTLBacenK5gHzvAzGVYgN9
qoOHU6azvW7P5cP61IJ/1wMsI+zFmCceBdjc8F4+B1RN70IeLAaOFkUKBPzvedv2
CzF1io5JLRA+DGcBknCmli2G1GV0FqnLhunMl054Qcz32mXDIlwkhkjFjDADftDu
CqG6LD6We7Cd2XJn/GJXZT8zZ1dsMI5wXOFNsLdwaAjYjPplrzs0zQH/tWa9LlTt
xRUh1zvRwlNkT/TBK2eXoXre2qtSsWgg7UsXBcPLJhKqr3ZX+g7vkIgIyZ9JNpDg
eOHfQwO7e+2xvFpjANur+B3ZoRsFS6qxobrKRtfCVSYENsWqjQT1aE7EJ7guWqW/
wEy8B8CoEcshpdaCW81qO+omRwHwAEwLCVT1wMwRYk02HS4o/2ie/Hu5TSM5vtSe
5aK8AppNW/1zOPfwRQ0Mk954ofyMMD7PB+CKiET3Pp+LZqBOG1/HoYijmtmBQpxz
cb5NpwUnIZ6j2BFhX4en86TSjXkh9On2lSFQj9Rok1tesGJQ6Q7nVQjvZe+fBKas
ItaLLSxyHCa1ukmDzF8cPZvaopsThhhDpL6cDP4EF0nucJqEJxo4v/b3R0XzHjqi
7VDJgsGxjojtwZV6erp9OQbHFe2LRx6IJ42qvJ59ocgAqfuHnuRSuJnnZ1SGORM5
tQq4LUp6zMKfmku+9C0G+ggapRzs6ckYjT6VemykLOPp5KPfJsNGYIJ9ItnhZKe4
22OiTS+G8rRJhs2e3FNgFIfNquFZo3MBFZKW8qbMTp+QTt8XLrqFqCbU1ss5yeUl
7Tc/U9UNVF2fKfKPx1j8HNRzb1QCYQ8Ny0LK3tkd9sBoJvQGW9PC5oOj7iRXNCds
mKmWMqc57dIUZ1PADvqsj178iN+vo8W3p3SVYhc+OQ0b5PqLMrtioBpk5pholMKI
x71IdFm7PvAJSD6rqb+oeJtzo8I/CEWbtzVV8WS6mwd5yt/ZzDkxulpJhV9lPPDx
hZ7UCdelsXW6WOlFpdAMD+TkW/7YABHW6AuJ9miejHZDKH5/VvaP4tYZetD00kRm
wiEIP+fOWBbvIoP9OEX8az0Omn41VMHZQcMiooSQZaXiE9Ca5Y2qbsKDHG4MOaaW
sxBnBssjBeTySp5yEdtuN1zg9stce1oIaXF+vKLgK8qS3BPtzz6nKNL2LTnRIMis
hmWjdyZRn9OXHZUUoyoaeQ7XRbFLjdnffbiBzn7Fk7LLWQjyVAHXb2aD/BVrRRl5
wA+DAaCbVoZ3FIP8oD1jsRAxCfy0Jc7eexvmNB0x0T7EmdIuGeYqxxr5KdErrUob
ZdTUfe0krWEletr/9VPlby2SSqA9o1BnKAEZwOdoFLmNmWIgRq5CzaNsXdMOubsY
wUVIUCScL+cZ/XQJhKLnik6VU8LxyG5XxbH3SAyZfBhncQhYmmJE2ULhmM/FgquE
l+wWHX0BlqomkWw2Dmh3HHRkIubbEJegadojAtdEr8OSVYn2DVeAuZETcbDVb9K8
+Hx4R4qtRvc6kRcUm4o7nvZm52Axrib2lQapamSBHDLgY/03UMLz+zLLjUNwx9//
ENny+0ERnGvIepkYVItNRXJS9UHkZFuvit+dMozYkOxNu2+jJmj6aLNa9ISIilpN
ngO5fQwZwirNUaH2RHn/3WueRxcnRptjvsAuK6H4CRuUiRidC0AOdSRdinvr3sHt
UrVboXu/A4zON93RC5UOh8uE04Nm1Wu8PAjW35QCJqR7T+UvXUaC+xAuTmgSfZ9b
8HTs4rTXg5B86+DXck22e4dhB1n5WRKEx2j/YUTSFguJNow8lFPUj34KFP1zJZNF
RkaLcIcEQ/1qAdpLLtmMCZsGelskN+Z6VOKzDGMUXeSiX27NgQSW2cyEJf6AvxXs
bJhOrCMdJkXtoHrMuwnYMNhqS1cRrNdo9x2CjA7of+wMDBwqR4m8ioJ/GQ/HXMLu
giKecpCnbP77aqagHx1v4xeJDZQ43kIb0+4/z5zhPYyz+VbI4/vb6Dm1zYbOzdD3
w0r4tlyY9G9LyK7DzXUV/YSbtvKKrxnkgPervwycmwD33iRkfUWSVusKDQffewEo
bUQNkr86q7cVfZIJPmkiwS3Qlh3CKm07KXsjXRGziQuSSfftV4m25Z58+/3XTc89
3yPkQciNPVjdrWQ9uVW4KBQWB0XLCZrHQu7L2XweMsPsi9MQDdyla0Cbr/F3B+gq
8HPfjbp1qtauAlBToLWmt4/+tHcqDL0AHk2l37whgvC5XRGMrDk59lGgI7UzUZX7
JYHIXwUntuTcnANgBQ8DmVqLJALS3yeiDL71o7gpfPlfycTRAQh7LNFIk7v37VBD
OxeIUwWL4sK34YlsO5Vj/l2Rz4IlWs9bY3CzbnfaIbLzg9nU+Nk6R4Oi/H+BhEEV
w5UpSHIEygWi4xny5WdFGIAnjneN2Ltxz10XewKUSq0wiB3AsrzwKmROnaxmNJGm
M0mwjQwiVxnyquV1YpHU71lKHxchMIJlkXDZ7B7hWGjTjEJ630RGwXi8INL1uXpd
GJHgtcSQo30n8jLLJ+inZx1ke6/3UDK1tw/6/PuNb3KSxNLWtHZNKtdnKdeeV+2e
m9gGoZ53LGGG2PX/Ntdgldbc9PPoALCKyuPX4jzbLs9XNI/aOm2INdo2VQxNVXo3
P1G++8PGLndWbRRdlkldqn7B+DK0CGNEbU933Pkm2KyLQnBzsbjtHV1vT7sKrDEV
2OcGdD5mjYZ0Rw70LbTx/JqCYxrblcnejHo07GOwL/aj+24JNa47TLquieGRc3bv
xAUFIH2FOWpwKLabocBFo7DUvb/B3Qy0q9B43QzTV1wPn4nLZeRR79eNXRllia28
9l4VlYP7FJEyPdbZeBoY52F6lbb5gOBSiKgt2gsJIWOA3yAtCvW25jW56PAWlc3/
0clxhASrubQhpUaCrrZ/GcLIxyDWZikM6oDw2EuKUoUGuCGg0XMWCI9djBhzRHkM
OHGgIrz100EKhmiNQhhPgdbk6z+wHfdXobuPU+LqzDb8dW5VWbRNTe+ULZA9ol7S
xxa6e+fl7Elb47pmhQsT98x3emYMh4yt2fghQKMWwbwioKAFg14P5ohfRBBf64rX
9lvM3L7Idm3qpDiPyefTNGiXS8/K46ctq/tggJUxMnyfR1R4xFCUryne3BC58PwZ
fTYkuqcZgY1dFjmnZoNVHJ9iR07I3DMr2Qs5MtPuqvWrt0y81QsrZlF2d4y+5Nt4
8WvF9q1PW5jeEW7+z/CATwuqNN3YeYzNATR9tEHkj8lpPYmkZvR4nq06T9Vb3pYb
cvVMtFYYVlVaJYJxQDp37EgcmqKUc+GGCiFWYggr7Y8JY7xK6mQkxky2xaZPiNxf
VI3D6JJ/UqcGM1NdsHG9z2SpMFAnUV6kfdROG5Ykft4JKadD3FStc4ty28L9zkpg
+NahAzfaoC95wxwYQRKkxDowhS77oY30aH1AYyl83QhEyYJCsjhcOItyyUS8NL93
UtBIGJ/lCCBIwFEypQZL+iSxfNzSMf7akEgZiwBiBVnfIRt9vG3jXOAOG9ttpUpy
SRapf0tgl6dkepza1qHWxIMiSre7u0aNRvOi+89Yf5t8K8RzrTLwKSsuYAj6EF4A
VrTgNTfomBrBAkc8QNA+HoszzClpXf7jBA69z84myUkBTguflWNLbtRL0H41tqDd
7VVQu532rKPp91i9hiU/4ZyczMHEIwtsrSNOU1S4lNZWf3c+/d+zg0Q76W7HyrIp
mMLHi9ajTI6LtFsI/m4p/YI161SPExscyDEaDA0Oa/8W/0Sdt/V7zRifbYtgJlaO
4UgJ9ySckMGQTUciCNygbNrtH626QxTyb3Vaea+Dn8lp/jct85NEeJBV/EIzuaO0
o4PHMEaNgc+p8+lTcjg69L65PvJqSZvMp4k6yvMoOqvM9TAci22e6OkQCgjzZvGg
Z++tBZkSQg95mIHR3izOn2Z2Xzbjn3zAVsMcAkfaeEZ0FGb+1ChBO4CeIR2xGIw7
2HQxf9mzCLe5/QMZn6TYSFukFJ5fZaurJwizpHh7QKeR1e4TZDfzHb0mqjtmZnR2
ppFF2KXGM4ZLxK06GpF5ZBvlfeIVZEQitm6x23r3ZD3i1StbdR0IIqSXsu0GXfu9
h9/cpZbSAK7aG4j9Nw5DQCyoSgHp7qCR8tZuyM+8+EB5Dlb7phNK/wnlNLsqpLvn
WLfukQAqa4i7PWUBXwB68TmgZbaYQSYjv0S+stmRUrSQ1pu83sc83euJrB5wUi67
BeXW2EuW0Q+9DOJAAvfmWLsgwHWdicWc+0NxuYtajxQ11Xt6FvHtJLrLgyncCRIp
ffdZcYoA60iZGy4gCnI7AHr4VloAmZPFB95Iz646yHp/5tRPQxY1RyWANiW2VSyy
57O+PWnkAYfXYVwKJ4iG7SX/hrSufmsriyekTlWV+w9S0mobuYg7v4e6MKs8YM/Z
uTOr8i5DvmGyL+t7thNQNTL1prxdRanreNqy9VjE3JMT+rUe3+cq9CrjZI6S/K1j
fP7DAVQK/kfNGO+5cpYtV7WcrUmgpeg658wx9OGoCnvnkNWEa+TcbMkMVryAEYvA
TKTCll0WHvtKJWmZWwsIRqjghL5P54DeuQ7JbCTfON5jPBomQYVKO5PyBLrjvGTN
bHaj+zcjgTVJ5V6N1qtwA6VOamLabD+t+HhiqlbB1JTz+jyf/ZxDQoH13vM9mhUI
tvea67xK1bAge/OY3jhjfNLczbwBBtWI9clV8Kg1yhZsUJP7xEngfg88Zc8tfAaZ
0t48biKFSN2WiFqV4xNXIWpwQb3zRHqKlahM06tKJCM9u4lZcoRh7W9XqMq/gyNI
fPWJPWRr/WK/dNYgVaYZOKf1ZabdqD+WC9Afi0SVyrYQ2Mu0eCy4cGoSXmLkKbNt
QEEhZ6soRQo8P7GvGDN/m0Tk5SI16KNHtZoLSQpX5yiHcQPFV5ekKjlTzfIjalIQ
sTeptCo5/KTX87d9/sRX3yrVu/CG5DrJ1dxWgGLOfmnS+m7BSP1VCGMozaYFLqx1
Dmy7rq1qpiTwGI99lzW9W/UjmE3C54CuFbM6z+txgc03Sw384AqWKAphemmDcV/b
zqLvABa2zXEH3hTp6f9NzXszBGmi3OxGfyScoTxwsianJYZFfCJTd5fAOdGruIEN
TBCiLa2aYqPRdUeZkjjtc3w6/TvDjKCzg4PEWxjKuQZYdnKHhkfbrziaR4Tc1/0G
Yizs/SCp1PqSZ+6lnB5uWbqTTYz2AgC0nlnA9M5bpBDdsIAiqDrQofj7TtNobCow
9n4jol/dTpirr2y5Xnl4iwTv77APCn86aqayGMwSFySCrd34klZo2uJlw6hEHlRM
B0BQrvZR9N/sez9iBYSmQzKM6aD8L2EiyME7QA0/NNebwa+iGuWtFgm4DEN1gUFu
jX2dWUgvxXXgizUlix/bV1+A3zFFKhHREUbelDeKKmszUD1fyhnt1QcuBv67sqhJ
VciJy/vsJnUhMxDF+2QR8+Xs1QQPROk0wiX0zXpq9+2FyOSaNIjKOUrfbC85FTbi
iLxsVta6PqgOjdFpaK5GQ+l/D3AtcM9LOyhDM984keCn7/3JEo8n24nbugP4vYNF
6b8er9GV7hnb4CoJ62MXxUtWsF91lzLQT3xb2xOEuLN87Wxhn8jnyUlmo6uD5v0R
kAND7RHCuARQSyqlNzhvKUeBVOPsO36tkMnD5YJLXfvIkBF4nU3nKIXNd1FWPobr
mnrtjTcX/1Zq+GRsN/CE13mNq8WM2nFO7OIQ7SM4hw2bQN+u+Qp0UlS0sk/lKT+U
KpXdkyKqqGSiCDfvX4Oiz7mwhk1TSv3y/pYFrTvE6FX70/I2lBYN/PUykMPjvVz9
4tR8LujfcpgOU5KNECKZP3QD3Oe5d85QOgeb6da1qSdxoeZVYaT4vghY1zIUaMdD
HIQs9/Lo3l1zFi6PhRedQX8kT4Hk7g/EZyzFUja7VpjrEakwYlBTPoYGlPngsSw/
X/dEuUR7VPOnFcIYzAoCyEKkp4cgR8ZLkVnGlpTabr1A8+OUZNIeVsHcuZwA8Cpx
1xw+76W5cHEdnS0LkXaT6VlQdvYLEFjs/iaWX3I0YWoAYl1FccNy2O867mehtPY9
4EiYX6PH5SRw1s4Y6eOOvzTDw2OiWy556mgVzOmcQHHR/S+3mC+40OIaRZ8iedZ1
AnJKxjSGQKnhljwvxqlMcURXXSINODVcQfWy2+TytfJIXK5aCZ7bV00jKVm+XhJ5
dGfU93CNXlwWD4XrUr+PGiu/4pJFAPVaeuiX+8j5t3f07u1zPCaiBFqTfdykk+Vl
nS13q465fg8gdpp6JRB7QTSVy7W29ewTlmzhNR2Zu6/lvn8vKzYHdwaSzgVQhcDn
vSECYSY4CQIQAG+PbPSShU9RzoCPbs1EGofrPvQjRZe/Baw8DhFtI4ipw+sa9wFs
yYkHuHEZFHUiRlX3cMLW860YDkoWc11ZcNpkGI2hDT+Ecn7N4IQClw42V7+nooZg
1EHCW24IT0C26UJ1S790T6rj6EFBGYo3XTYXlwmVWCrMORs44bo/APM7lJVv4ipR
tf137jqspGMG1K7hptE6wHc1bPaumcoXRqo7PDPhyP2m0l9kRK1GJqzoEoDBPXIe
MoUEqyiABDQpeBhCyeAe4fJ/K69HuZ6r6t6QK0G3Pbnv48UsnBqRVWJJCJJmbeIb
1KtTUseoKfQw+rP4zQZ2ofm0Q24g0lfSlRh+Ht2OVwCXRhc71vIgDTB1rVeUU7CN
P3xBYm5Ofhr/pFAjmyPtqpFzrbjW19nPiCcTxy+1wDYp0/x7EUbq7v96Ihq3UMGd
ltC2jB1sxIBt5A69TRg9vJlZolMzcv9aqYbarmLGBmBZtSfqnnmGWUxwoR15/Q5S
FBPTrZf/1mW22FGvp71K2A0FbPDKd+8x4J6IHHiM9cPWtc2ph4d3lWcWkM7X4Gge
wKBYWmF7MzUP6MJmZFjk7yEBgHVdUoAO8RI24Dmk0BeXeEmZ572lCLYpI0GoCK+r
QSzwdwZNsB8BHRhN1nfZgMMZQp2xsCbHKUdctFEl3slHVi/J1p0NYnjxpai3sV/d
B3QCNF5ATgciwN35nezPA+ZPdSbNoRi9BzCsKqPe+s4Xv2KZ61sROUfMahNBFgL+
9MTIrpxDmD6YaDv/tztiQnpldu+XkgRkQnAnkwvJmtzeePIH9EfDjBIGY/jYumvg
9oM+1E1pzmIzY9hmC5ZDTkeKIYAY6pmRywdZi78KeplzWxCMTVW8qEUup5nSp0xT
ysZPfO0ant+l4YYa2osED6dfcSgTgQWtifcsVUB4rJ217OtFPlE3roBu0GNpfEj7
hzt0JSM6XSog7pBMy4hhrz+WbAaW2AOQAh31p5E0nUqTrGOWFpNzGL9PQdz9Fqax
f9mYZhAjgorz4J6KxEmB/wNNj6wK7RsCPHEFOnQUDb1sDDJDnULJYgJkPq7olLFS
nU4Yee/H3AiLfzmXXExUHFK7DJRRssQEC/BlvEwxbanfzG3b2lZK0ObESFDdudye
yvwkAI1VDYnsGyVJiRE/9nzPg72/qAjQUL4CP5rdoGHm3eRqS0IjmwwZBLACYkAk
8dOrxX19BMgQErYv7Dz+jtrQAeZyaEYIBpMeU6WbwSPag7u6qd8V2eea+OAOiym+
tqyzQkGPXsKOvR8zBrjBHTw1BIlb8e+nEEUXY523tkmcdpUy7G4waOrp42CKhF8N
zYQ48RtT/ws2w+ouRauC0cROTPnqbDU77LrfAhR4B2lpK7uo0lBMYKkKlHsdJ4OZ
d8TBwOqrFp3AOl7DWL4uPeDsEP0CshRpTItfoffj/MjWRFfI8x2QDrKKXHtx/zFb
t0gFpC8ZpdAaCMpxNkFwhkcAh1umY5GVwNjQDZqU0th5PqBMkn00zba2JYNhssrs
vWPK7ctvDO5/yhPo2YjjNQGxsbck/1GWVnIckHlExQRzKaifRuJxYdLrXV1XnNcL
EVkbL9czALN+KgoCy1QMyg7Y5hhPTTdZdBjd9TTwHZniAaIF/tBtH6Yc6rT7Wpdn
wt4WJxTbX/IV5j1THS/6/SR72Ppyn+Pf9ymap446C/IBo5sARMkQKm7wk6MdEUC3
MGw8tfUEZRJjcal2/MxO8v7SIF/qQZ5ln8/cH984Wwc29WWZyRvv83gCb0edPyOa
DIDJYnGU51aeJ6860a+8vBKJ68c4fQ7hXkKbktTXjDE6HBAFJaaEfife4y/RbjlM
F+qTMi/udon4WnpWSZyUvQij/k8osVsTZC4ZYfRDawravsQbjJTxtILwQvo+IXqn
Jfz7WCFeoh7V1kBK73D4BVo71J7zIJ33jsSiwnM3Uc/wM27tW3hWACs0zb0WADNu
8olaexvgCIs3v9mVLtFN4Lh45MUDQpQrP3OVb27ZB7WwoWbkpdIyXRQH0UMv222r
XTW39Yxs9g7sdQNw3FJapM1lRPgCT9j7Z84GCNvitojz4v4acspZl15lkA9w0ysF
fV0uJiS9lk8FgMKM/FxM/hPf3MJuXq5Q9bhoXNcsoJLzelk/atNCqdayGk+eSCi4
8XS1xMxnX6WSpQ+TPU6UjgE0nPifI2TShJsGoOeJXh5I4u7WHOYdl5l7I9Gn4HON
C1YR1LDL6sdrn7nxeW+AXBzYMdRdZehmMgX6yEJIk5twqQpzxSyt8DU76NZ15Kav
HS7TAgQeNic6+NpxkKkGtCA1Nu8zJImdXLADpzUN+dxoPNyVbuH6sl4QFj5Fc8lT
AGm/dRN+vmGbX7zPmtBcucFvpU+z0AKCNG9msropZkpV6dCv5UyDpLRkDTv4HSiu
Q+LtI+QjQsalG3Y9m+kI6LsmyYUITUjQ7UKrd+8O17H7oWD5U7IIBEARveLhfXRr
iCxFyLtHAeSv1ThMPT08We92FddjQfaiARPZZD6lUJQYkJmEOFKqeUxiFu8EjBUI
WpeOF2shpwHxWMzYhBgdmZGe2C/XI1FlGt5lDXncRYfi5WruOiKtofYJ7ADaWerO
sBCihRhAaBFZrQxzgupbKFr4Apj9FoZ3zCHuiiHoue/gRVs44u+hprUgnHPkbAym
Hzv1j8ZddHcOyLWXjj1wM06PpwexZNq3TloVe1enVh7fbRUx2cQdGT7l1xliCm6I
CtRtwpa6ZToODfkB+M68/Te3oUmtWgprLo5tmGZWR9F5BOR99MdVqwS2gFnmhDmW
2CTOaZcV3DMQdBg9IjE7hA+SYD3pnigEH+lQaEPfTtlFVHZfeDoxACk6L+qtLO34
hNwxUAsVESRvW3uP9/IqOGs5ERhIxCs/TsFF2s4Ib75IMVzXuzWhaKdd0tu6rzse
kUi8ZcTU4FzTV+rU0VWTHC7IkqgVdxLE9flpLAdCKSyzVE7NcF3P3RDFAIrak1qA
c1p/w+0D+aUlF6Ot497S7P9t4nDJmbUdVdW3BfdTxyz53wpBtb/KSB1Hz5cPzeMn
v3IUobUHizdJ6oDIqCmef7iMGpPVNfsacNURVxv5kMSdj7aAKzjPKS/Ieg3VYSDa
Pavyie8Hy9Sx40fcz01u/6vnriQv14+hlCXQyPNmnUY6h1/AtleH7SrWLXgWTT2+
6HxsGxHxJsOraZiI+i/0w1Do7PELk0i/3lf17kWmWuU7IqsTy01YY2yauZWFgT7b
6rVZMO10jubXxkSvP3C7xoyCYAbBAQDSXkScwrJFT6CtlwhI/WNCCneRP4DxgV2p
dIF/Ig0XhLqEDza894ivuDPQRAQohZyL/wRCeHziwcBdK5p+BonJZJ2OaZXVgPc5
GZ0m4RhHTLZS85Ozatm/AKAdiFMx7kLUUaFfhXb/B7KaP74NX5Iog6coyWK7R+rM
JWTM1TuCIiyv+NlOwug6tKPvKEZkTYyqlnREENH7XWJjCY4hcrVKS6c4InUCUz9B
YSo6y9rG+d03yjDR0Cr1K1dgKSknEEUSL8h/Sz15mDZnub/LPZgdeT8KzOo9JPUD
Emp25YcgTclphMimS5mZwTITDoa73vWl8qwpW8WFzpHpYizW3beWm6ZMetor2Bq4
+FMbHufeY3Du4l1Wmimk04LxmulcRUGVQzBah9xLu5xRqjBH5ewKynfi3NF5oaqM
SDUoKFlNJkg+yWxsglnFAjMSGXVeWYoiBb5T0LqTOHzEF8dnFBfV19jThrN85t6C
6VP1e6gujjV41bzBj5q6k4x8zeGXeHDJJUWyb1iLDAz/GYnL7Q8znA+7dnyi1zYx
dimu3PPLcss2yBw/YZMWHNhDl/tYKYtgOjFMl6gTyA8we9j2f2tDrVecj+nErdOE
apy51Eb80YFrebIXU5W5PGtR4dSIMv4PvZ0LE5KKKjB+lGNLLtiQ2YpBgq5qwTar
/q7hYGdQZyTzrv8uRp1KDDlzqMcOa8co5m/Fbuh0quLiKiEKo0sVdJbEV2mj41PS
kwD/QuPvSvc62+zML1zX6V7JFzmUk+g70CZ3jvzJi7BlFsPQ3UhJ7c1uU6Kyzy/i
0NyvoCyMlfP5x+XFs01w++mmnlTr84aupcfxrDjMVuhgdL+7GrnhlYo9ZdcW2sdg
ehUks9KtwMluuyP4wQ5VGdMYddKpX7ld/W0lgPYXkkH2jztOmUq9McvWpcTuuFrr
0VWtFXfhmVfPR06CZ0zLx6dkTOTU9uq0V3XegYbxkfbK3GHI6p3Iu6QKtR3/bZdM
pHTYFMFwbicisEpRGvDuUMjgLIv26O66MNf/albEqMMWvUh/EbLzjtX6c4cxj2uG
m7rOXPISKDi0eivclCZCdmeUubrFT81JE+goyBLYUJ/s9ec8U4yZsZtAQ1hhajKg
JmCzG+8r402i6YqFP9lZpXB12pxUl3IC7z89ZnLFXYJS1nD1LGlpqJdYswCjN/VD
6d3D2TtrLe9zOPDmYLOicxVo2mPoXt/++6k6XKFNkyda9UG/kYL70hfDtam/Dd4/
FXkyExpD7SryDraCiC9sun6qx2C/0JnRgq229k+hIPSQkFLgVlYlGBD0Rh4/aKS6
Vaf0WlAFMbMeQ0UPDJAjloFPc3/1pGTvLxPBrCXkz8asn2dkO1hfmLG6T0++QeVy
+99II0SqhznslFafXYqvujGg8gVgNZImyUjcqo5PfAdzq5JKbyOq3aeUShDyrDKZ
V7zG8KEoV0w7nFDlZl2xlMw0hwaxDGwa4dFGdPZymwBB47h3ML825Kgz8e5u7HlA
VdHL0t1X/buZ7V8wa+dcUajZyLyZX5ulWG8OuqGkffLY1f3HYBqp0//8VoDevmIb
DVEKxD5DgR3LSaVTMaUpOVuZYmJ2BOlS5ETDVJ5rYRj5BKsm6pwTJX/Mzk4KBa2Y
oFileeIurVlBPStMokFhEooePo61Yn8iLIRZWPiQteRq5Oc+2ix6mS0aiSRQhoIv
EqlqREqvJMbBzie2JSD6EnKArm4FnrHRWPlBZvMhIX6ej70JDQJt53jiluR9I0zk
argCq4jAzXncW3q4TYi/ZQmSNUbmKSiVslXrP+RtfhNmmGShS68QdM5cD7W6Vxn9
XqYuTmk3S+NP8DvPtdJqbRY1hUsMbYCj/KVk9jNlpfuabZsa8R2ktrcaf3CS6SaP
zj/0utnb2ANwYSNnqGAIFXYlgx4wCQSElpWQiB+ye9O4B8oQHFW4rupS4qdpF3+l
ARfGhc4CA3HjGr0xkv6YXn76T48kVXS0BuVrQe1seT+1g6WOFa5xMQOjzinychBg
xpH7+xg5Dl87Ig44mzIdYwF0LMrcqfmB2+NZTm3YbpvpEluV47gWn/xAqV4NFZ8u
o8aepKQGDV20i8PfbqFdJHN2yjnzTgXF4Uu3bsfKjuIRyafU1g40nr5944/GTEwy
ATloOagqo74TnLm7nTHhMhw3u1zh92wyXkf+tFDRd03SMxkSC2lOndvLVbtP+mLS
OjnQLQ3Jk3UA7gBkUvkNSDc9CfvzmYCf6u0fSQUe4Y0Y4X5ozadU1hAsH9s+2dWd
yjt0LQ1BvVbJ7boya+kg+/JcBXmJPnmkM6IddaeThkA51nX+YZZk8pVgCHbqiBYA
h43Tp+gFfNtg6nmsp0og5Glq3POeMj76ggrUOaw+b2PiWLUJmERTAG5/s2+SyL50
ngmdDv7v1T+WMFmLRTOR963pUavZGf4419uMqPmLhcycXq7MpRVsUmT2SJEeklto
X9LfgH+F623yXUQtmkplTnZkPJnL3vDM25LB2qzpiWHYNCKoQdgIFmo9Vw+GN3AC
tJBEVAFnTcx/VsAvSaadxyyv5VfzwezXGJ2Uj8yQNfUZs0cSQy5w5hhdTaywhPYq
bHmdlYUFfScbdg0je7Y5bPDLcQmQtESpijmzTLtJjYbPxuAPAGlFELaLgopOG0Y2
I6zEfjo22QzKNYhSs3uro47lMknYfzMkf++74+D342DYOBJH2QlD7dl/f+JRvbMe
s3vJ4BfjI3STy3wB8hJkMkVTAh3cyOELhNPVN5cEKbB6Tjmp7eoMfMOktK73g7Be
/XrlWywv10IbLuXKZBMRW8eQKGStitk5y71LjSUcGUdD+EaoWwyf/9dRPgHvHksG
Chtagy47AUa9bxme9duInTFBFoaiaGtCGASRSJR8DefQXABw9Xgd0/hPJl54k1C5
HL6SyTWTc6HSo0yKDfIGQFVd/3FDrZ8Wou5Hp4MfLRo5l5uiz5p3JOkady7UmWCA
ySfEK1UWBEoahLi0vohV0bdFYPVyptkxqqWncNbpj5cTZuBAgAyFZZrE7Wlh6yIQ
HCJCwD9mYM35povMGzHhtoQktnxbdLZKJCiMNj8aL3ONIXTmNjcxf7Eyqj2g7oT7
GMSvLANrYdPBJ58dht521cXMBT8iszic6LS/2akDM1X2zin4vA9jesoQbP8UJ7RC
chKkegVgY0zEak3xWhjkZcZXfqBMsO2Ph8vv9kxSMR1mi6O4LWAxoU8wmmqeyDb9
dm48bMJ3++jOPQ0Wi/bkJ7zmgicOD799Wg9mZh7FX+K0ABsarNOTSLtE5dGE1B1v
yJ0GaKYor83zFpK2JU0h/KPD9k7giGltnVgrQlBShYRkZmXkZRoUXY5W0pAJdMIb
sApRo8wk1GUmNfqmeNshuF/7VtqfvygKb0/0UmDSAq1phle20ft9u5HPRyiYkQqw
gJ95Xcl/y2BBpbwxLz8IiPQ+8fHV3Zs+qOWSS2j2XQJbRN1BB+i5q4rda66sDwRj
N04UlBGC5c8GXMx9sGsRBm9ChqVgd6tMRAqWieYE9WH7V52VyooV2Vn55thjY/T+
2UeaTZWDePx1Z0FsDhaESer1Iq53M5EwuYVi5Zcl3qW4vIwpy3OPAdvLfpsDDl41
wBysJXOs+gjRyUTbf+7f+PmDUoe0Qcw2B2cRJG/n/YPGxT9/JBf/BreTPbiHaBt/
/VzPOwnVOG41zRJcJqIwImwZIFY5rTP1sp5T517ikphucdqH8efgcstWpiVYe0yx
g4T6l+R/+jO8n027eB9l4rBTx6IE5Xd0wRO7O/uZXaYRrzqE8l4tfsuAhl1jUFGa
ZoKGkaBfhGIc7ABuCbNZdhe5U1YJcauSCAqX+c6st7n4RviiqmVkNp+D0AtwoJk4
RdeYlLgGaB0KJfDUZHWpdf1gpieuMy9gAFzDZjbsOH6PEeRm2NHq7i5JMyCUUkOV
CAF67McGseWgwBOyJIs1PSsm/jY/BKFgLijRQPM5WkeMBteXoW3RSTjR+VtEhqZ0
HluHbRQu5B1EC6SXCBIUwdWZXSvMZWjkkfE5WoUZQiH3T1LRxvtNRYa3jUYIzjlQ
TezVU7YZz2I8l0o+nnvvrh1BlnmxPy0XptvY5hqqf2+k9bs2g8cBSQKfuVjl1IiA
0gE/Keet704mst6MTY77HQHhxLTI2MWlznSY/EYGWCu2qhgvuC2owP7XonFFxAcq
Xv8dSae6iS2U8bWdU5ZunCit+EjhO9rnuRqgzv2VUgwuICfEfjJyvpSR8ACKaOXB
AX28iDpT4yeIDDww1ol2CCVwZRTXEg+ltXwwF9yh8beIu1jZxvymnsk7DC9lwCAq
qMqB9QC1PYcL4aByX4Q/Vfo6Zgsr3w8ktwlgVbb/0xvvX/b9ppUJAZmC6BMyEQoN
WcYveKWRdwewy5gx/8ZeL8e3OpxQMw3h8hlCtud6Qh2CEohmoDilsEkgLY67a9EI
8KhSqhWs/heYN8iJIvo2eff+1QKI3BJQXL99JQYH0god5PHhawnLO2/NTp0w9odB
YlGd1o7XkUGc5/UPilxWMKLIxfG0+WlUgviu1sTakFVKNzYnETvsg91X0tCPb5K7
mqFzzvf1Setyp7BcRRkqvGUr0CaVFicn1oUUdNJLxGNrYD6NN1H1v1iEAIQuQOH2
gSdL3fX+vcAT7BFRGqYMwBafnYd1+EcpLeUwQYpPmAiM5FTpU8/oz0HCU/ifrItx
qPh7wOu4YvHsC1V+qBnSMXN9q2GKNtU0xw6V/w4MAw0MTRWwVcoK9Lc/IY05HlM7
b+CLI+EyV2LHoyWkvVXO11szZK2BbAaSFFRLtB6PKp5t+4zvM08/2/oVVvg+Vg/e
UYzPfegaRR9/PjB9MzV2PgwWA5Lee3Mu1+A2/tpRUIScV6ootrdKbUv74jCB0ET7
6Je+bqfDsysXdQvEgwzFs4nr5cquA/GVGk7+aBByi885YjWtf03fFVcZXBYrMasI
vwkZVc5nJNyVf01qZhJki4/g1FvFmk4rwE1IIxD2MRlEC0eMoM0TIIY/GyKZft0H
5KEzKhlU7rAbLeiSQvgxRovV9/kIHus/A6VEEKKnYjPF/IMEvPSsJx0RLTlhJSWg
6WR3NqdK8g1KD8Jlo7z8DlFrGa/ZLx1DGXIfkCRfyv8W74Pbo5kyQXQu9hkIQ1dC
Tld0aN7AJ2pEhkfM/rdBjcM9vzaOPifVBSFbXMsFfsynyvTQk0YiytIjsol1baLv
7JpWQQw9dioTfWHb7TCKZjfkvbT8OI1jzBJTMY27aa5IhNaj5V0LTHtHmlZqhijf
YzW89JSPv8pLljsZkHIjGeQjIvoPzo2vRk6n26GbSeddQEenTaOOZosB+hIY/gAP
vtvR4eRnR7Qx3euw8yruo8xuQFhf3nGDvcVDerVPrAIIcc8AjRQWO8c2LgoxfPRH
9DJdf+VI/Rf0lx0eQRzsGqChsBaLEb8SPookr+ohemoS+35wDWTQccNLrdwfqbQN
habqgVQ+4F5JFPxGs8ojTLjDf2i43kqUnbdammrfOe8g5+lee76w3Ud12LzKQuTW
7BCfVqTcUO3nUpDWe3FMmt/JwGiDLqUbF4MMPGCask7I44IE7KgrpKGm0FyOjcOd
2rUduHcpsTWQ3+7+6S1LC1ZajNK1g04ZBnBtOc6x4cVNYo/ALH63NjfHMgMiH3Me
nyFhtlhsdDjEW633xqbCGWVgumZR8HB7Ncla7LXxuKarxAYXIZgW2ieTso0Hzwzx
EK4gBhwbfALFgjJjLa5Pm01M2B4qhuYTo7f+ccJyq77NfE4ixX1SkFr6IyKeeqKW
HHpxNlr3dTvI3K2M0oAe6uZTqvTwijbzo43l6mGMyupGmyr8ITDKHl+5Msj3R9mw
QavkatSO1HMTFXtNDeFfcm/aVP5ehYac1IEa2OeM5kkau+g0RT4KlxvJjVF91maU
CtxR1xf5N7551h7yu0XhZjEsq08KxuujjrVM+CMkP4vG34p1ahWSuv3kAI59kcji
M/98YYYnkqP4+Xjd9W+b+RJ0MyIjq75Ge8IKeoTRAEiJj6BTH8ne687y2NJClqHQ
4Y/zIsbHv+XJmUB/I24RXejd14qYBK/JPYU0V01fh3cj4JimRMRUp+g5fWVNUde5
uTLxhxk8TibDc2a/LMBR2aTlMNmeu52OfUSqYQ+5C0Pu4mrFBIAyURtKZBowubyQ
SPie2g+no22qvjMIX2Yw4aJn+xho/znsjmM7+FwnFYeqRKnme7G2rryg2M47lZj8
TpHY6HFP4X0Vr2C2V/Agd4+4UqZmbuBraBPOVce7ia/daDV1Jt8oPZnCB2WCgVL5
6VxU/aN2Dcje9vpX1Z9AuytaLTOqrT+f0THHjz2BNMpztNHUxCh39IoNEPmuFOf0
xe939rXOQorVcjAGMMKKJEG//ZoOonXwNkv1i2GiexSXqL5cWlJnZ5mRcqWVLym1
I0gWwEmLdg11aMWiH260qu/fUYA7xQyeEY8Fu9OXpakN2Jab16gH9CiAwzigNyCr
U/IAoyoksJxz2/iG23tIuAj3o5KyYdfM/roO9Wep8nQijQftK/DAQaMkmPja76y9
QoVqFUCV7eBTi62KCPgLAV705gmaJEvOvD2X8PwQrm2WgEsX+1blBPeahzRWuOtU
aIS83CX9bha60qNO5EzKRsw9Ks7aD3SS+newVvhWACkC5+xRqgF1d7T0C55iQnlc
4pdqhk+SOx43fG3N8bgvDN1oO7mRKIRnSIWGBel5EUwx2b96q8ubQz6cRAI5uNVd
0WOlGXXUEUBeahKocrBtjUL1HbBZ3V15uaduDeOia9Fvpy0f0FUK6zevz2AFbMv0
rx8FdwOwMJx6SrJtYXhzwPMIYNOmfHM1sqt7M6ZFdhhwbzkvznfoLXcdjzEuQayU
XMUDoREIxlye8bJEypXMi4bQVTpMH57QaUIEiWs7eaXYUSWHKqJJLm+vItytzFNG
c8rb7FZrU2iJ6BmiWWkv5I5QOoXgF/FJgJcy35AkeTAJqn0dWasyErWy67IStyc9
9bE8gXTxNV/DArCXSbgYzaEvlMJL1Lwgt5QM3iO48opKb/dSAhxB+ilSBgaP6NP6
7SX7phsaaodb+VvX6vEjLnQx8wlppRF4ZTuAFyfO4igHpVDVTTQao473j0daercr
UZHgC4cdX2wpYLaVZ0m27p9/EYH6CpeHHib2OGRNOU7ag5canjSjSGkYB5YlCkXJ
+AaqzLdCkdmhSEZtbW0+fnK6Zy+oC8ed2OmU8wXaVIKioLwvsQXIZzFXwzc/6LSs
N22jniL1+duzYvhAi61vwhD8N6nVwoxLIkSVpzHTMODCo3HkhHiz30ycfU13fPpW
ipk0KBZUYMUjKeUaSiujTvRjf44mDtSTNKR21ZlweAnvxAVNh6WH75BhPtaw9Op+
lklm+21vxFmkk0GmeVWLoKxvufL2J14HlrcC+i2DhssQDpZSqRBxxTb44X0EUOPF
fm3+vYIVE63B2lFXqq40NKSzHopb8UXZh7dXqGSkt+lX7BjOVVgGtcHwZqJhM79L
rf9AQoXsrugthee7go6QZBi0YlfjOo9Awe0KhGzkpJfKPLcRw6G0wrZJSS1l5yaI
QaJfDb09LkImqDUrUh6vuayU6Fqll7j7qdgd2vLQvcCK2kz1VjlgoshQs8QZ7WRy
7gSNrnQbvuVL+ZBTI8dIWFSrU8+Xt2Gm1r17ekQk8Ypt+xqbuTRBtmjunoybiezW
6DQrYPB5YMeL+bMcfBxBY2icnbfIGp9IVeajdX4jW2uyiuUbr5TNzUaLtQ5eJ7jV
gGun97Nk16UjWbWB+Q0XOAxcwUWvYlNXzzDQlenC2v6miqaD+K4IoQVWKpQK7Sn5
qamYuf+xS5S5cA4IxvE2yVkweqROetBuggJwBjW1s5/fhHVursfHeSxqhWKJM6zA
bTZavQwTxgQvAp37omvA7YwsSnENzoXQ9RscKXYo/giWyvaVLqpGh2rrWkDQxzs+
PcMlCI6g4QjNoQbh+G47o67t5X5bqDQxuOKmcAH3J39sTMpdwu0PHQdlUMOO3GAO
0xa/UCoxoVvhEOVhton4k2Y5hrB2UPasTSdNroxbia1RM0R1qdQyEw1x5JTTiKhM
gk6S78CZmf3BBCEXoLER4BpcKY/o8Oo+m+OJv/17R8GzwGwyjtAd6NV08fcJNddV
VGCZffiCZxEVtZsnZ78l2Vd9R1jR6tWtrcBALDlvhLIRbcsEts0VFHkiR1MEV3oU
rxrMpK6Ut5xSQrv18gJFgxs80VMPX6rEFJ8bZHRZTCBI28MM9On3kdnCIpzdVAPX
QL1JXV/5AdRofXQcb2eaRlfUzYs0c/wqZ0P3JwMu/Zujwv9Sc+iztXzulyVn01cA
Y4lKu08dFH96ojzQoJbH9yH6TANxiYNchhzvNoGk2eK7eEubwRmFkDD4U5cOwGBZ
f7vk5nxtrNmbnJxDTaYSSknhAVLx9r0hwmnTL30jwaPmCYMjs5VzjlxmRdhwshgs
giOPnbrrWD8m+XQ4Ni3b6FcXYGMzf7Lh7+lCSuNJdRrq3KLo9BNZfkeyclLPqZod
C+KEkMV5sYDTSC+DMG2xp2xTlGjAjLyUdKT7v4qtgUcEnvAxCVFxFfQOWaa1fRSs
3yyzrhkn59XAyJEiqBF2RqBknYSGPpbd5k/Seyn8sI3zK8mNVo9VCoOcfAak7s7R
qlUlk0FcN6o/1vOw+0HmtWVgjU9cyr8vRjX/t8vZ3iOYCarkNSzSmNAr8p+cGE9b
EhNWRK/k1XbzHlnWXQBNznuiK2JRF7DYlbdVg4gp9L4O/9VR0zfJHi/UznkLDPm7
TWX6d3nBUrQ/en868kE/cRGrUbe/Ooniouf1XSIuSWV9GC/M9CZSECootbzqwhXQ
t3anPFmUScN5iXuo3Nn6k97HopGH+EJ0wkZxTBkPG9DjZy4O3AlDiodI4EHTXze4
fGIoAbCNo1sX+ysM0R+dbkg69R5qYr/4jVG/T1KlaPq59GqWrMECD9acU1HPp6nm
62GcJLJHuy8rmCvER5bzlbM+Mm4MBmnmQTPnfYMp8RfUtOsdWP61tV2q9wJY3/JK
PPA1NiKOgixP5QTj19DGIk8sZfxeY9LhwZdyzRYRsmV9Ael6eNXY7riMYw73SJAQ
HL24evpy4iJSZjPcZzL+ASlXDTKjfbFyjrVVCiqkNoeKPD7Afnga0PQPMgm6N7sF
hdFGD2DLXjdY2dPv30deMOQITf3V5y2/rTAqpZ8x5T3e0SS1aGhiMTf07HEyup9g
E3bJYbjSdJi6s28TyiaXxIVX4XAOACEMqZ/OUvYx7oGc/wgHHAQHcJ2hLP2LwL7d
Ucmm89qDjpp+ha6RgV7vsXCG1CmqvaqxMCOU40y1XWcC824urxtAH2Ai1k8v5MEC
IdajGkGwlX1IsQFUt19SYrfVaD7SKoVl8aD6p9mru3a35P2WyB143qQMWT5YZHVn
tzUg+xarFQCIQSGquz/7Jgr9oNqQ6vd5um1R2dDb00k7vtnopHFx03nbJJDYq6Tp
k+O7niz9jp4RFxGE+UxDjwpCKSmJcClO4EfF497f42/mPG4fMnjYRARor89154K5
Dq3mXM4mWpi8APYktnv5E/9tiMHFUGd6rksKzPDWnSex8cKp/mInOejK1OkQKtkt
cehK2JronvQsCqx1wergS5zS8rYHzbn8boh/YKV/YKsjHyRiwaOSxeYX+CuU1KJq
lVJ3sP4TXq/KNIqIe/wobnD/W2qk7UtuoNqzX2H31FnYwf+GVu8qPheQyOKQsOQc
HADdYNw9NPdZ1DLkNVQI/VWeDv5RaD5R2lNoWMO7UbjWXp/Ocan4bcisoVNAiTUp
VEg3opEwXj/59bazfCQzLl6/FMtfe18T1ot3Rx/WorrdswC34c2Iteoqt12WsaDy
GjNGmoaY0faWiGzP7xJSoWAe2Pvy9CieEU2m6OctW8fIKa2EElRmkYod+vRE0eJf
I8mb9zxvL5jcOLwAS/VzYDooslHm65rgb7i3CdMPlyrzDfIJokSLxQF2bHSqJZ1Q
S5ALJWSLdLNKoZ3XqqTA7T3QSo56ov1WhS4sQbkwIQWLPZBGtVYtrdWHTghxOVyw
K3SrTtmcIukMLZqqhixPpHcQODGMjR+KlmNgMmsVncAyWVXcYArgY6D1e6vO8DUr
jkyDo2G5uSIBIsGXmKQlLnsCZkI9k55TG4v/lJsvjpkMgICnV1Zk/0HrmWlyeRdt
NDuaBQ45QAY7eaIvzO4nIhyz/1Rdr9yRmPkTeE77s37Kz5gCue98rfSbd6VjFvQ3
fNVPZlEJM+Nwv23UoCNIR/VqPNRs/0XQZ31LnNq6fHUF0lZDb/lqvchr4V4BbVUe
B6V223Zm1x27BXIU74VFiezVlbWajv5/GbpxzD09LfRCW74n49HS79X64sxFO+2v
9hR4Bu10lOC4GjGw8U1UgKM0u74umwGX1fNH7lCGzfe1bYUC212Ypv1PBCHVlumV
lbvNqTY7+/F3ApB4ReRZLAHszwyFeEliV5YJH+PSKTBecvpFOOCZRtP2VQThoV++
9ImTj729ooZN5n6+iALKfKDJ+NbmQjFOURIHHinZL88kpTWjqOgyZuCn3SU+cqMy
kD/lxrtBbpXOUl1/mGCoyFbxRM5jObEMU5U7R8QNHjYmqCHaV1KQRqB1LQD1N3XH
fdMrPeGyRr+V7fiqL+2th0+Uofy2QRQiCJ4LMdPlFlmuMJydeSB70cu6tGQIhn+0
W8QLbndUz4ZLV444J12zBR1T5Bx8UX1E0fXPR8/yrAuYpZFZDugdmAmrOA9nwqqK
MN/r4cInZ1w4Qh78/ih+hMwi7PnU9f0f9jAvNM4QxhXU6QWPG+4Jo7mTJwiI0Rr0
us1qMHllIYvI1xcK1j7ll4R9SqGu/gX0fUS1noUYC2DULLfoznPw6sTlygdCVrwI
buxzttlTaTBsobIgoIQJ0Sgur96eOnpMvPLMaCZoE2y2+T8uI9iS9VtAu+gzn3/N
UWwi4rIrWfJUWBsJpbaLc7kf1cAoI2uUxXA7LWvg/w6gOWyt0chfLcuaVCneudBj
pTYYzjT8fBjXonf3b8i7nWsXcK72NQHxP3AqZ5G9HUnytkttSQcu9GnjLw3QYvz6
E2q9P/182IPgvZexxFHgGpqPfaiX1EFyNgT7xg96Ia4o6h7wWMXwNfssJisGYr8B
cUteVd567UTUORWUoq1dYAMpN7oRF9uyP9HQEaPfDAm5Np142JGDI32p1o5AO64L
XpE99WRJgupnrDisbWMRIQVoxTD0JyegNOsTHCJdL9Bgketxp+Z1E50nCt1DoYBk
Wx7CqwpEtSOGHYouDhxDc7zbObufK8XYd8Imrg548b4RSmJZTN51p8d6hMAUBtdm
lgh1C/WKgR+UpPP2JkHyn+3O8uThGdDzfCPyhqPhJqsOMTlcWlJV75oHfGnecc+0
zXBRoMY8MUo/eXVDAPqRzkoi/7tQHj3SMitcMsPy1Ep/kLfY78IQQlhfNkKAkyzD
uetNhrOK0hhyu2nJ1mvjZ2LQd4zc8RCESnx9tvkOAwmVXfsTVysifnUyojFWDWpo
PeVWmS4chC6Xw3i1LI+rOm8KdeFXyHjOlDrYmcDIDU18Hst0swu6Lg/S60slcBA4
jR26MnZT+2xZjk2qIA71YQWHdzcTr1QYdvXBg/yEYnvuj5Thidn1VDJtlYGnMw1w
Mo4D8896yXkcpWNT1krAQ3S3MgB2T+WfSdRLgxNVoYiXBUkEVB1rmX9gPIe3BTKx
e2euVeP7//p7/OgyVNiF2K3hsWQhrlcPLTr7KCGDcfmpwexLuJHHQDlE3ITU62AT
KES63JzYsrEl810c0d8Uh2cW4/7sgQzD0+a6dV81t/R7vzFe6ydQMruVVnCyWCUZ
jkJntbffbVabMMFP9TX2P8XaybmRoQqe6DR4XdZZdtkVQaV/2Vq2zlRAIEv4pBcj
Gdpu43kZVxuxufYPs1gBX6ca8xCwpCCe4w4Umo1exA6wybFzRWf77TbGS6hHGs9V
Qxlb9kgYJUvNSoUBnH2NY8CEuQLKTzSmG6H5OZaZjEdPtGq6msbL1V59uzVQdjO0
LbJUrjuIBBBftcP/sShzAKq7QHyiruBRZCVvWk6mJ/0qPkKDjMg1JGYXygDVtpig
UfBIMfkuh/h0qRF7CzNdAbTJdV2sKsKCVEeWBlgH20zH6nx3TSMfVY123s86co2X
7WFsyzvMxXDPmrJpsfjanC+Eg1nHkMIxgu/ryJwDc3n2ewkjYiI1mpbn1/UNCWzy
Wfgp3fmMTILcFylzielxj4uAmnM6UFJlI4SMic8MMm5R4MdTmPCrsAOhQlJy6BrA
5MCrNk6WO4rncLg+Bo25LHLKJr2zYw6sNXVK1nKFL07VPhsmMOaPleqtA9UH9Uie
KSCVw/02tGk19Z+Bqhb0Tt06zd3yAjg31rlqgKso0+xmqIq3g8gTdaAUwGy2GOzl
maVu1n/wm4DvvaNc+0as0pDi2eFrMz7o9qoBpKGds4SyVd0mikI5VWbgYrJor/ON
hat/22IX8vTsqmvrdkNNLLf3///2x4hXpV95Jr88czIXs8XtTo/pkRwr4CoO6q1N
h6phRz7NaU+p/I6T3b59gjJuaBGxF8DqpW9HvcQkpxbqRjRI88Luc6PZY9BppT2Z
9mnnaqHLs8/2Ug2b8k7cJCLtTON3tpGjgpDIa0W3gjb+V3cZRMRHH2uua4vUQ2nW
WSETuihe+7IbSmOlObql5rSseWOuMKaiSQUOPu7LkNnndnWZlcjgqIS5Dhr1Feh4
83c2Y4y1KkZ9NwsdvH11isc2C9Kw2cHB46e6JrOGr+XlpQUqsTEIe59eAw/VzSl7
Mh/I/NnQljKsxyFpV7uOjnQNo+8Dhcb3UYuwmHAkqY8nn5VedYrWhh1y82HdyJeB
/XH4E6qpMDWqLgNGhMQ6EnxNUHbsrXv8Fq8gztyeM50Mgok4JgMWuXvPvtOtomRN
VQ/Mtwe3WKA6ALdmjR2Z9DF3D4F1LZWWq8r8pZhyMF7aVn443S8iV0+ToOjdx2Ia
o+d552UGLiYPPIot2Z4JwV+LC8k53Bf6m4zlKh93jqJZrO3CbavCpzo6Anfhu564
9tV4ckqfCr0W8loRah7IIOKFgXOE/fS47DYNCJ1JZfqjh85dkuucTOhGEQQ+rtp3
tKYt+AuofAf8X/ne4AWFILS3+mkRD5y3xMoCWf3z3ZER550qSAwHo2T4889Ie2gH
+Hp67+7J6t9zqp0TDtTkY3v2wZ+Bn0Awfav4m+ohQvgsJpOya+GpwKjMJ9fUvA4e
jJSfB9NIJthjzdgihyXVcX7vWZreV9OJ2g0vdsOX4sGlq275SXN0MRIyBvzLSKKQ
UWqrLSNBj3R5VxeW3IZ1gyAoCfKLkiAULLmrZ6ahfnDAPF+wzmAsbup2QsL+/JHK
dAMR/5w5/xWw/Xk3QuAQ/G6zu4dmjsxtPjMwKijz8XIuOCX2uYW6jD98BcRmAx58
x53CieduS06svqwZioJt69BTDQm/dwm8Ng4VZSNwRr8fRq4bK7Ew+jj6pSBC9odX
ElylZaHRPO0PEvp+ST54hgXzHRTWcp15hhMaae1ZTw5/wIY8Ev1QFltp9MMNkxEj
2q2VuQAsJic1B6YH0YnzlzMQM2J8LTf/fzYCdHxF4e+OjqQ4IAMXT2MGyWdV8lm3
eDpAZnIoDNU2obzOKRxU/p5M63UaTs1I4prCP96eK2AJd7FGj6TLmTDR10p9VDJJ
QVATfTsqjaqAlEw91uf0ML3QoWzQxCAlrOJ7DofjEsB+q9AK/ZS+QsPxkbhIzPFa
/L1GZgJ3t7d0yYyay+vPOcX2Mau98GTzttXvxkHyGSibU4r+4U7ZqKKTYUKXz4xl
nr4hYvTgO8hZWbKW9iyoYmNFk+0+RxnHQ/N3n9VeviOfBBb7bdtqATEF6q41SP8x
KQCtS6Jpwnd68O9bX7/H0Cgr5+oPooZP5Jutiowsv8Lqe+SLGJpiU8xWyK3W7SEP
ifjvDCssYajrZsO1b4tSCBlAVTQ2GGWfxZ5d+Am0bkOOa6r+jGjmGC1UI0c6SNq0
qrv82ZTfKtqNFzGvaLJtpvQG+IF5iHVooDKDTt7zcAnOVEgQk/N43/bntC4Z5Upb
sYpnqHIhMPEckaakGHxuM0Q1ykIxtzDuoV86sJyuM9Ep7UDE8bBPYMJgQwQyCZ3D
lUSrEGg64OdNk/zxvpSZyMGrJZHEFrDwZseXacltJMxr3k7wPKkQVHqFnUbxBEoY
RHsypDKpq/iw3Rx5FoQCOgKC/3bB3I45IHGfQ/M7Xe12fVPWiPq8JwB8ehJg9QVH
s00yucqfy3QgcAH4fposG8w9Xpl3Ibys8u8ofAH8ELc6MMWcIDPPniO1WaETqU4s
5CnacWEuacTb/oDIyeLoYnlTstkQV20ADiJyqlJD0VbEbNM6s5THVIihGRGbWQcp
ATyw0wXKBOyKL949powqGOiqS8zsxv+18M/+x7KFyDzx55qTlGTtTDXED2is1AlJ
gr2QC7JUvSzFNcQHG4mR37bjWluHS632K6aa/nyxIAwidR4fsKPhnQHJTIaHSbXp
Eu0Kr1m3jO7HkPguLFi/jpxyZV4gtaKnea/keyTrYvmb0pv8Y6NUK9vAemISzY+c
+cfwLgHh37kwlloSRzan6Aqzut4SYHqTSuvm88ktaP8cDK6PficXM+L7kjDydzlD
i2BCtE24v/f9p/aRvy5eRm0G4j6h1UcuTibJ1/PsrCGY+19bR7QOr1bAjNZB567F
oSxGfvFb0kkVuZDrXZ8fX16k2de5h0x7Erzbd2s2dKXpD6JSTdsGPrnHhuVWDLXl
QtfevqcmgKMvukPCz6Xf7O3iJiX6T7lQA6ME8hRw6HG1qvIgpol9jSxt2HcytKXE
7j3tntcwmo/ULYqVHwrdfgpLPQeIzKe4wpxU2LWcZ2IPIZSKL3AHUotXn2dwvD68
OBxiJPy/evoowZXT/Hss6kuL2bdqZp2+G+DkVUwkzFOQh49FTa3jlsJDRc9QJIbC
wQQKflGA4Hyuda/yebQzNPHR3YD0O4X3g/jeC2EvOYKw1e1OtBUPK1j4RKx5eNM+
mhdkOQF7Es9aGM3XcAmU1/Zq3qOdNOAl+kmR++SDAuLHZcbZ920qx8tS+p6rBu2J
UCpiN95eMf4kW71MSYwv16Ie8+pb8ViE2VQmbhYChVESE3XNQdNirRmFQ15kcHhJ
OLz8pltlEYfkgFkOXVU7Aoc3VFkwOnlJYlHJTnspRVQsVvHr7DRHymCGS0INEQS9
r1KqPx6DOBlZcqomn+B95Nsz6Uv+JXHLx4QNETUwpEsx60A/JuQ2q9nC1BspfpQZ
5cXThH44FJR3GHAyW2ZSfQ7vCBbyB87wW+ULysjU5OTJcSea1P0y5emTLTC+X/TX
Nua2vapZmu4TLHkW0UuIqBCWJNNKOJwlGtxHCamXxhZK6Id5E1O86/wpJyh1Ve16
F6P2JHSIXQJHzEKjTAcZ8BWy3l8DMLlXekyvEYiMv0kGgjd/DdP6lhwzF+87Te4u
l2LEjr0VYcOpJK56SzH2M8Nq6HOkMVyLjNKcrg0Hcb5Edu+R5umuch4B87qmVGDL
upRaGA0cMGEQzK2VR8wfq0fWAqSoyHsIzWjHUeifydxJppFl1y7HjeSLClVBIfk/
8yAtMUxap+bwEc8vdDM/v1Q4+Zd33iQQbL+3xEx3kWPMO5GL5KIgHZPS4j1Ha6Il
XlIO1d89V1GYoeidCHmk8d4wiah1UmMFwAk9pSkhjcVX6RoQLZicSOn4bdKyw7zC
L/6ewlELQIj+EOp6JMHHGmoqOMzWh0zg13LFGgTnVrBzWaJmHjB2TkzmqaJB5Mep
NTJQxyDdL4QHJlOJaToYtbXujwkFnGQltiDSTy7QzXiCewUPm8x108oAcvRMoJoM
+hKSuYygxDx/vAv3UdclkWo/QR2p90WUGbSpKotg5O36MDct+V4xcpnyqrnJjYzH
go4Cmven0MJLHBr+OOgRFDf1WUQqDhHHQL23JaPg8DHF/Qt4km3xunRQRgtcn3Ly
7G00nWKfrYYO2UYIVLRSkk7H3KpuKtfWpdNZsqa1HUksP0pIEKHLLlrZ8LqILJik
LJwomwVRDbqAs+33eFu7txYqRKs9t2PQsLda1IGsLn6MBVrM92jXFIzKuHIDpSDV
QsIJCE20B3wzheY/e9v4+bNm/U8ZOuLH24F3Q79xB0iODl0WbMkIvY3PAp7PKNqt
PIsA2i3jawnG+awZE9unW2uAuX7a1GWS0horqzdvfsPLVpiWzvQYFkvnnvR1V+gX
Al+iP3uzWF3GWEc39L6rF9Rj8scDYtaCb8eBZ+eNPa/TCrz1VrIY9TyTlE5FTYBC
C/Ho1kcOgjyetlAzRMKGgsh3xH61spwlof+HmCiFSUDl8450b+53lvxUamO21fvZ
DylDVRYWmwfbpM8vH7CZfWaGsBKCsbc5UNlJLVhxlDuyn9sRjxFUJlHAcdiWO50B
ri3USL0MpwJnxTnj4L0jWQ1iJWA9tjTeMmCzBpI15ce6fO2OHwWW6lzTIIaPHqWo
eXnnFnvRfuoCkDCaucjDl5DSLtb2l3hvFADb2KpPffdScNEvaBt/S5nI9YwK+rEu
0vZb+iSpsRaMobLVBQ4SB+PHXNeWYncgUue2khEDxrrIaB6baGDJq9MPQO1Cjt8z
obv9Ljb13CGU4OUYG9415I1QZzOrS9o6Adsc55U52x18Q+1KEwwbpMQ6IA2FCb+q
/za4K1TTMDpVt6OzhuZpoyZFT8GXNawIwrRDSOpYQrPYsjmf+Tw5v6VJ77dZkBzS
pjjP86xNvFcGHDiD9DjMGPhFcHyoDKBvCcFitRg32eKFCO1BR/E54/rQMVa8TY5N
tFgqu03DJCRYe8xuyT2NhP/5DbNdxpfyc4C+ReoFV4Lw0EIKR0yS4GE22b2NGPPF
ayokh7GmQSiRtjD2l714pS1HxmVfJiNrhRahkALLpLvIRvdC6AjObMf1qKg9w/9G
nXZ8AScV6zBzqtEc1riDzubirWVnqF4UlkqTiAfJV6bmva2j/ThQ7LZvh7zQTYzq
mUrBk5a1xC6u1TfBmd9MSWIBXoCaFUb9hkPLz4xVorWbN3Pnl9U3C2Eb3qgUUEhZ
KedF7qm7/4dNwpTdg0YhSlRtlEvsEWmGyKcAtIlvc3fv1owmpkgaEN+Bfd4Awv8J
G07/kd3OEbqPh9JD2Q9z9gO5op5gNxUzGmfvNgWoMIHRFUhoiE3JttYR1RxafSfw
Ndh4h3hcAWoG86FxiGmeCz2QkmaOzU1gEbN7AraZ38yn8ZOvcn369l5YTquCIFMg
irZDUGNb5/cIrDpymhluopohKbQsheT9b5Bl7ffqUHAIg4o1k9t+FwrwlSmfQmse
EZzSkqC6fIM2iYOZ3qoyL283AYhoCYIIp+U/SLAWJayS+v6bizNs1hSW+3TJ8Fsj
+w31IAe4qI9isD7JSzSyFNt7aB/dnLC4uq7hwAH/up2zNdKv8O4tXMkqDazlP+bE
wayLPww0k5IKylnlw5ppaxRwkS2kaIhRWov1I+08nAP3v8XXCGB1rds4Izwy4UY5
9jHWp8QJTaxuFR6pdMMXd3zzTD3BwY7uyG94CA4HO6wEKsRDnECEAyu5B28NUi7b
szi4F273DAeossd/ee/eizMYtPn9T7CC+Uad4BMuEt8+xuHO5hZFLWIj5cOWldj/
gVYXlINNSB/5+pesae4I4WWwa7KIdkNEdvjzb+AOmEGamrhTLONgR4+4WxnsPNxd
Q/psJqfvE5xb9UDHpBFpA9lChAqzHlE5ApYUWK3hG+NAFmBzIQeP47hM+JJs/H67
K3VDuKKXzKOqXpAzp09HcH0shjIAL67rIERWti+OP4mqMHbECgDKr4pETt1Wzr+4
yEoTCBU3Z61SPaMPY9P/5pEZVtIMT1pIwRJ3n9DJsMlNdHntaPRG3uaTK2Wsn8HA
zrv9iAhDHDGyoRSQ5tFJMmM+b4mbRz7brWjnAHpAjr5uql3VUQWMnW7YXRMB3KPo
7CgL6RkzMNBsGSQ1ndu0VfApCaq6V17xNH/tQk/oEjODal9CN9JCFQVgyiU4vaX5
womN1bLNPwq+sxp9S0jZllp4AyyV37IRqucpLJYgFEHJUlfizvHl5dVnEiUnGvLe
iEZiVN8fSpEGgfs2uBdOIZb+LA5fx40OHAAjlzZotdSxfQz2v2sz7n3lqSJjDgBJ
Hyp7e3dR06AopF6mYLnts4IejsQj/0Al/Ue/Y4gq4Oc0jNd4bfbYkwGd2eOkw1j2
8sJN2+o5tF+SAOOa9wX15yUSDg9x7LQEEX5EKGKMJuarO1U0amRyzpOBj2Tr6eP8
nYeeoPp4expttPgj+b3weS+RvNl9ap+KEzFszZ7+Jejuwai4dObOHMVxqKk6Q+nb
NLwWT7fe+2xAFME0KS292CN5hOMxXdp7lL/3BNAvWgnjvuneCeaTry0ITcJHjI8Y
nNnNeN6GZE/unZl7C75OHog8QKeGkyjpzWvn8/g5wYcRQMC8jpR3OC0omualMtbz
lZG308jAEOuXXCxOVgW+GvQIj/TxWgUafQnyDLuQSwI6233tcEGU5pQlZ8dBMmmT
GnPqhOEEIJPDBj77FIsK+NkkAhOhMtSY3GN+hTQZ4a1Vq0kETbb5k2kG6SDLKJD4
/0DGgxhmBJ/H/e/uPoYt1ZBSGzhVCEeFQ6RLlxfXDAasLXgYb9TcsB45J2RpXq2y
Zf0mx7BGw5tDvrLbmgkgTvslFaIX2tGI5sxyEIYnylVyBpcVhJV0GY8wJyVVbocB
QC7nEkuzzgv44K2Emj+SkU0kSlNAKN9qZshzkn5msm7Sc+QY4MUEEbzmqT8Dd3az
IypuSW8sALrCHR8gKRIub841IIzHaO69kox/JtrKi3nuwW+jhf0OLKAs8lcrnJT3
KqkeiDBQwFkQlHfCBBTL8czVTkKaOox8ERz4GxlxrFdMQ0jkd0RfHs301/yu9odP
ai0J24FSAMmW5/eny+2ia9eTF0PR1KPxeiBm5xDXb4dHrhF7HPJ1BqOC8Q8eHPyp
2BTUc6ng2D0aou9/WlrGyT/GN5KAFVrYzW+DAUS2LNxwpmjKjNFGd0uSkgikhFys
T0elshyDBhSzVjujpnlJCRcX8/tQEG7+2M6yoJYUWV8fUNjPbZ2EcJ+DLleo+g9G
ZExGoMf9XUEgRViR3OaOhrM3K0kArTJNkz7i1Q3bxtKXP1IbfWhnVCXpF/QXRbVL
eVfAMw6jegWC/a4mYDaWneTQZyMh+MyP20hTAmb6vu0EoiUFiurn4MD3fsKfO78g
FfUniZHsl5x18VlL2mQUl6d+U4okiA2vgPf8ru1e+4eEc2lZvjiGC2gpb6A82eQA
FeQoRmA7kBeZehOrOG2J/4xvZZmUI5O7jLdgkbJnrgAQEoEQatC4DMHjhw05D/Dc
KXbb5zFZgBwoVkJst+F0Ha4oldQAWGUZB5bs7ATG8CLiUj+wG0RjxYQKv+CEfnMG
PIQtsuTiS0oc0RNTLUmuP+T3mHypofgfVXPN/dKkZXqJ8cU7zqe0MYry5jbnJzFr
xYlpLZcvGUln0fO+Y+qiU7JqK23OeaV7gZg6hvq629zj+tL0pWo63qd46C/5OZ/x
SiyuEZUlDU3YmFEZS4zVJhHgQFSBKUGz6MUCeYe0J++f8Nx9l5D9OTjnZ+cFyjBI
pKFBbAn6+ddyr5UKTOybdPA2gLyFS5zHJSZDLJbnvxinti67Q87sU+NKSWtcOcr5
VE2rDNP1FVo8ODNH4HHLsQzJqrBiUcT6CFHv1yl5f8I+dYmHUALXslJ/FEvG4jmx
at6wp6x+4RIW4iCNcLXCdZoB8opJaNm1k61RM/z92T+3kmUe2+vokwHBe7aVBdG6
PPxizL+FDXZjLEuIXqHYR2dMa4W74EGzanQRDlzS/B3EbxCp0ezszuNqurwgaHbH
/T/pzcX95VQAjYC6J9JVpp2sJztwSKp2idmLjWtfK4dhV4mBvTYyJNgKKfQMi2T4
01JhcyaeayI+QVMFiP5JqoRC91ahD1z4wBHm6YSEEGZ3a/Ay/S3ZgdKPB5CZsDEb
+2+PEG8qjBtHqREKQBG6RSdHfWQ8NJ6ZsajZCqXTqH5d6LGbefuhszKX9DGHJBvP
CRe67Dv4AZ0Jw/evx4yI6OYl4I8u0+AQdQ3MH38y2ks+3TKMGLRrzUqqwB9gEYay
MtMBKb20Z9Kx3OHW2t/gQXfpA2wJCJep2XlqXCjt3N3X894PVB2b5HaBL2zOmvyO
lgr4yPC/qTHBzWOmb6XzUXiOs6lOcEwNI0BCa3uzaAINN5ALqeUOB1JO3WTwn6ki
tnXhzsuAx1kVTEaL+DzoQFxOEP2HKeZ32sGscdh1B5L3AxW9Zi6pVEkBbFDzRD+i
NkWoHfYXBgZldgHF7Ha2SITwXzRoGLWmo5ZhCKZuP6tJu5jSYDGsFKRkfVlLHVOf
NXtgdZggTjfG3r+saEfxqm/xaI/141ioaTCS3XAmGW2jAhtftBRNSh6hTrBxGneR
iMaRapAMl5PueWyyEoNEt/0QYQ300+7ZVuC+zZqOqcFw06NsT/dQ83T5P36pi/Uq
OTd1YNj3PIeDcCRNWoSke0iBjlTnbtBl2kLhD5K3MVvGM7kmDZ1Bl6s5fCEQpdGt
SKnxaaPX2dAbPMurGSfeoVgctpIFE40HdLnwaCvzR1tPK9IUqIbe/nsl2mt+6TLe
0idNNtg1yEisEnTNj5hq+E0vIEOaGZMwElikP5NOp9sae744llpGFNuT8bQ+0UHJ
sxx2fHFO1pBuG3XWy8BYLyA+29rNAOBRHCKrJb32HSXUNITsCGnUi7owxz9DeByG
vBKufhNrJQNXNzxHERlJg0+RrVHIMiIiYq2Z8rSoCXlm0waUgrDhipWlwGD+jYRo
WL9f9TDrAAv+uIBapod1RI+RbD1HU/JvlF3kvzn+6NESBK/Eev+0TstDvFRK2DlD
gEdwI1E8Re0zZrQ+1FbzscK3MWyVeeUcYH2sDm+vx7ZY7Q+zguOewkSvvwJb9AKd
eFqPm61na1hpF1vZ8qxbm4MBdkigEsXxWsAFz0GCOCa1buFKal7CxxcWhLP0YPut
grSEifMibcb6nmW7aNfvE/wKbSxwS6yGjd1Q+aQMHnHKx5nSqFufZ5XpnMuoQhCC
3yDez1h3jGTpWnZ4fYZ6wsmchzJ4A3wznPAP0aCaOr8eCrUAHDbO0twGkUsKvaZ+
XzMTpn2qS8D4nuPHmO4mE0CY5C4uqHRODNPtbGyJo+yy0p9S28dzL64+4knQ9RF5
ryzRSZUvbs6LmWvuujT95LzI5IV1FQyFwwojthDoC7nqhMGsY/fBLpAe7qHP4sT2
jljcYV2gbyVyK1k+QUZ7GAHQCFtJCUy4YG1GyGQyHg6qqKH3X8r3pXHlq1RkYg/Y
TowGRtqDkgLqqdbF/RzUtlVfhIXy6lfoViZ3VR1iOWDu+Evsc+M6V6b/Xs54m8WL
Czd9MGioPM569V6kQ0pZ2HvohS4x4sSWl0PQ6cJ5nBxtK7u/AruB/p8gVKjJu4/q
3Bt/XTQ/ieGICOgbaRI1JsI1iiAAerfohKYrvj6pbe/qTzbenzqleLyB9jePu/k/
vq9DJQt8FhDBYvarPrM+espfRuv+I+0D2902AiNGpLUQT9PNqrGCu7piKNcVKCT7
Pbk7qG6EyqhRnvlx0wiZZtfDo7MXiESVfEcpwIqmd7suhA0JeKGcUzOtjI+8kofL
I/dKJ9EaNxdHwkzgkjzZPBVTU1LIPzlZs5KoV7CqewAGJ/Hkg5QMbNM8B401bg2Y
CkKQn9n3WVuRFzFR70cfCipgt1ovfv0gMtlUh7YuLdwdh/ySssbntaOdfDTz0Qhx
KjD/zbqHx+hsczWVp+bMPO+BcE+ytxH8iRfRHNq7cpzeLMRMfUmwQy1K1bMHBx+s
lbsBcYca8V5uYljq5GoiAOPYegaK1ByhOWhsCvPzA5HBEq3JRdCkt6WlNtqLXYVH
KDL/4YYcHc0I+1AZzNu1tAridhF8Zy4Zc2jWzX4l9wsOzY0gCACrNbCa5193Z7BR
Au1ztioNHhdI2PI5s//7cZ4xoDLjRai66tEbAJHkqk0qbwG479/lNWB6B/O+cLsr
6g7il0AQcNBDXJEiKeUTVA7pjxRobDDTrxVfUjlf/9gNwT90dLdj4fPF6yM0TdAm
k0Znp6eyv6CGhXggCdDe03FfQkqHYGBvYlpcxy3ZiRVU6Ax6C3ERDeNUG/XD2PNK
7wQcJSod7pKEqRkG/EZg1NP5T++gnlg7oxNVQpyCY+AvUqYNiCUuh94gF0Az/Coo
4pC3gkQ1Z9SHBZagvo4OMWBdfi0IaDnn3PBjsnzRYLCDUjLxTS7miVZIuydIK85B
8h1bgc2FkJLB/sciMJrEIiViKLHPZOz/6Or2MHD987DpHEf061V9bGUeTPAPtjO5
bxGGGhO24rWY3wNesgFE+MIYe0tpYPTxFoRit5q4WDY8kj1WimmPH+g9PFBmaWYt
/UkiASYwlJO3s5vcv5D0LzQT+6TYGtE2pGCebzIpR+r5BI/4tiVnyoT5gtR9L3ny
r5V8a292ELdbclrrvUuyut9maeCYQcRbt6AECQ7r/buwe+nK2vUJCPnpN1MJ0EUv
HbjY5dOsM3vJNoMKShYbLZLLcmykn7HKnEpIV69yIhlXcWrECob63pBHCL31Lan3
NnHBEkK71JSQSX8G0fz+oGdFM2Ahg3c/CWaLE1StLr8HbuzgHDQRA5qXYkOEXEP5
p1AFkw9+vnqOoFEX7c76EynuZitEjIz4GhQFO/KSj9qO66M4y7Q/t4ugIiprm3AK
Wn1h3ZxZmTaKs/zStdwIM0x4R9583nhb5/q4XVZqin9lHx+lPcDm/lzaUZ5VUfCh
4bGgaMY5QaYx0H6G2ygWVbufOoBnll2GOCOnG27/0lQFU7sMXFACFwQIWsEBQR7D
YPSshVajZ4qzWf4a9z5xPXPZktgRCg0QEYyuvHv0GOCqWDcfxAcrsCxHeiYNWSz0
YXsEemmvwLKQY72jbr5+LO40kYchi28/mzyfmy3pY7IboHJEfSFILEG0o+bzJgOj
f3KcQAME8din6obpY0TXIpF7VQ8kcJq4xsxOgK/EFpiWHfBwkqZ1Hu5NPQnDBXBr
91Ghw43O1wIO09XDsPyhaAg59GLw42wn+IFMZ/LIICnv8Wdkr85/UI51Lmjdv/LQ
Bx0NKlceVG2PvzuSZ2Ua2mCHyNdnXCLOXF0ZSmW7kcfndv6P17RDooXUHxxjTdDW
/xV6I9zNcrwoNUrnSRw6oVaJJws1o1FHhiweX3e3eC6pA+NAHZXLzTspC4SLUiYK
gSo3Hu86njmWTSXBNY1ahwHzxSEfgq7rw4LUu6A6KlNTO98ApL5W6BYmyKKSm/8Q
8detkeS2TWRa8NOt5vApJWLcxGiJqJEzIbLp9JIPUVwCN58W/PTTqDbrDOtOe8uq
kLaA28gojsmyE+PePKjONy+H7c/VrHKTISGSCNoYoEbpoQ+oWvqg4nK9ABpd5C3r
FduwtN0QbxLLK/xrkuiuCLXwT1Qy1zuBNMiXiZheQGgtgiZdnPZaIrwP0It3ju2r
eknhbgq6vorYs6onotSOyFKKS9SswPwWRqv1Yrw834+JFBG6DNKWslW4MTePwwCS
HNeRC+d3jyq/6ASqBdxeogygLqhghVs7yHT6TP3lDUWcqKWK3OkiHfP+FI81cVjr
jKBiQnb0p1Bxbxx8V3/an7Aysm/qHHDGR4CeqZQXMrLJEkBeCdPHVLgaAbRuEo8o
A8NmvHtO7iAoYWeGajIvJm4vUSRolZK81rMXVVzJvjPVQgVD3QpJiNXPnq8bEXiX
O9ZBgVS89MrFTVaeb4uVyMC16p756vceBysl7FwppQJ9lA21sIJoHBTWZCAkGX8w
+UxjjoKoc9jnzJsCXw4Db2Hje7rVCTnZMQc7cxygyj9qHaID275G7ZJ31pJzBMmE
NdvBd3Dy6jUPGXOY9W5ACFowRKtZEHBFlv5/yVty86Gm8/AxN6EtC8/jajUNu13M
C2NyPGOr1g2ykTjW5A7fTtxdWVgxZ8yHym9rLDDZULEDLErKkCGplFhSoajDGN6z
oo7I769No7+mkrCSLQQMV3d+3jMvL8Jt47hLihRb1YK3gP4CU3QavuZ3BIP7Ulw4
Pma7DhaG/6hKaahIB1vw52624dcA8GCeTYrFYGkz+mBF1Kid88+OXhpc6hbzIjkf
M48mN9xBk1bRiyilXoFm4aXWIn8azkEodiFlyyzXclwMmmsJV8cBUg0Qfa1YqXjA
PZoSlnVR0+kax1H7XUPE/SG6406+zdSobM/K7QDkQFTS4N7hVXkwSoT8G1+pQPD1
Dk7RzgESGgDFQVZ7YhBlIUaYknVW6mUaf511mbq5yWeBUe299dCoTsJ38Q84zb0l
5mK5pa899xw/vev4xWrLdGQQWNBYpvC2J0XSINaKlWiMDyqmX36zZcYhJSmaxXTq
39TuLF6Jm8VnXT316h1tJizCAg6JhVtQdzSpl0DXqb/p1ZcDref7yIfhVk4SX1Mt
83NPu6eMsLglAjjDC9LWEnhBkVHKgpcp0+QXajMwPARPRBW93rAuQ3eQxyXFkCg2
7wV3nL/G3mcxSBhSnrxPbMAnEi+lF/oRyu3aI9vkRgbTlS1MZsD83DqsEYoYXVj7
VXgMiyRPJx5RHj0UGP/p7zPeg6SPqNEnrJyXx41BwP7DwHf7r/2/RL74ng8MFAss
FP4dsp3xUOO/wL+ghqyCal3n+6/uKo+OpPaQcxPqtFraaUVZPSdBln9jN8v3ryfp
CQ0V2y+KUpGEctaaRzUEWPD7kfi9FCSpFEWqxLiqV6sMOQ/c2pl9hXolxid2/pl7
XpUiZjR+vW81U5B4AieBF+kjeSspB2/jK9Ic7ATFZe52y6a86T47m6JKu3TJxEHh
mk6RGNCSpA1cULsWcD+X67talRAo+X6m0q/ni9I2a7zeFVf3EjTq3qjHW9ZY79qb
V5SOpb0pCaRLkOH4BPxLNjS9lsDo0ItXqr4bAoX++1Gnnn/m2dvv6TRgXynRBD0D
qt3kbJ9KyeoJAzam2CapvT+TFy/98jqZBWKkpZzNfKexU5j70nmNWe6ggwR2Rq95
nPgxD24EDU0vRIe0FX0PRq9Ee7UI1GFpPyi+RiDm+x4OwQE5OcsOJdMBsQ/fO0Sd
xE1z1xpUZpkPEzD05HiHJMa4gpItSdWOPfLUjI3ANtS3NEDVoyCkix7DGu3SxNIo
xuDwNv/U3O9eXfV4WpUdCNZgERcFGd5BxjStumYNPcWCSJvgp/W9pEi/aw40SojP
41/SRKgcyfJDHtXzUcg2CiqUPMD25AkuTdupF9Z8Ezsrqm3kJ4QMgqBkh9aRdMoM
5hfEefGzBTD8j7rERTDbJ2UiFdWc66VHA0LDTiQdRndIDvTIzcNrAOkF2m7e8VvK
o2EWzvDcC/50kuEDSLy6Ts8cMAqdmfAfEFh8hsIz5qoWCXxMz7/fobC22tP1dKCP
ILHQfM4Pd6x7hpDhx3+1YXLzageUwjeLMsTH/iUSZtpChb5+lD1zcG1vr6G8mZX3
pryxCoTQzNo0OxBXiz7MLavLdnyk2N/j+H5k1GkfmvvaARmpHFo5WaUJ+ZPeCWa7
jw5jPoq5PsRASOncyTEIN9VWcTveHBImhZm7PzovFw/nAmY3JU1hdmqHS1vtomcR
md+8MbUABtRPhy0GQ7MGaJckKHnA/s/KkUrvM3chPDd5jvWh6S+IToMeoTtmoGcj
xTp6ycaXy+Vgw8kb8ncpc1Q/MAInpWZK4mS7iZRgNmSuTrl2NUMLy6j6OHXi6wHp
rcXft1kKpCCXjfq9mgy4dH1r07thFeaIse1bdimUwZ+TkAR8hMPVOatOiWe6SV4K
utwNkTq9lSYYJp0Ga8NBvOfP1iAIC0bWp89IlnGN/kzugvIYkVX2v9Za1onr0iMA
rJl6QTbLt+lOpvzvvM4R2NXGixXANVkLW4hKQS4p1jFFuV7sMz7S57k07L+XH7zH
0Hlj6YB84TN+n0DezOvQOrQxAkzwCgAjrNM/P7Fi2UHUcIEBrvlgbM8poleCAbdI
f+RTqFk+Oe0qtGqkouFZ/CkAA0Lb1bUfOK+vT3gT149RNW1Z+Yk8JuafERv1fS97
oQM4pUreZ4Tl0NMajC1qcGZJAGxqQ1j7mE0wZRqjgZhEXVMHJCWjylbv1amNcQ3J
ZhTsLv3sy/vitlgNqovpwBp+CJ5uUkfFdQhu1/Agt6lFiHAFYDiMYzbcTJQ6f2o8
pUT8E8d9IN4Xd/UeqGSVc4fY6j/yqHYNQkRBkUuN6tDnwC1k9njd3fP6uGEXcuCm
nkXUGzxLxuJuPvOEQkuK2uUSdfhzWcGSP7t/gtZP1XZHtYxtmX5W5kCSKMy8yici
bYCY3idMBiLl191gOcyhsIyo/Xx1XwwdmdiiNqxfzSid0Kf6jVlcFqcsjmQTXHaY
re6V2UTILqOUkSWphYifMld6dVjIM6QNs3mdVK7zWN0duPvLAiMqFv6z+tGKoIOh
6Q8cO8MIKO2m+7heu6PU9Gkx7OTCxuLQ7zvB93sWJkFa3HEXOz7Smnsdf7bnkqiX
4Dh3PuZFcmRJqzwb9ZVyMG3w0CJcBLnVIpEdrjZkOFkgl1CgpsbEz+PU17ICg/V0
h0uQ69T5IgJB/wx+N+aLpQH7ZRuoEe7ed06jIYqaPNCTAFVsv3QO3LdbcuduEa96
f/WKJLnXAasJD3/8vjk7mPzVrTv4+BDt4vDNwGvUEAu9vtr507dBmgDMQ0T5B7Bu
KeVKcQQWMGEBUN0997ShjF3ZIGBW9S2jeqOqdiXZMTagz56e2OBLRkB5TaOvZjg5
1TPzBTU6cgkKVSCsgdXZR3y64ma1YRo7CdLymaeZUdf9LN0ORr2aJtabSa3WAG02
FrmvLiBEqN39LExfDj35kQYXNRsp9ZVGr2/HBVdz6bAFXuhJoJVnJLiuRqr+h8VN
/eCj4zB9MzCkvhTFH0rQJwKZtQCfRd26X1QJumIhaGWTodU6DywmKBir+iYd5ORD
z+e6KTauvej8Tv5krro42cbGN0lzjI2QYWlAxVV2PIj5kRlnwFRotGprMpmbUJQ7
+TYb5g6JzudDjamegemlra5xItuJ1Q2S/HQPS5ddajBkO12Qgi5sGYMRmWplsUmA
+od2OPbLqmGQKF/TaYnzxMNeEd0w8LDE1aO4drFRRPV/1GiI37mrx/PFWA5Tj7GL
wUx5ArsiGpIu1a9poRC1rqsBfVbhmPzv50sZxaEq55iR4i2PXnXeFO9Y+w2Wavuw
dqQgPMESebWZXx+cK8YHXusC07RXaPgnMIBay82TgAqJi/67YSGuFVlBFD13x8DW
MjjNWeZbKEH3ps86uUliuQCH1Kac82mfbCru3ItoI5dAIs8xpdbjp/BkfTtuhI8q
2Xc0YflEdqAuxLgzthDQf1TNt1BThIrwsJgUc20aNNgrwPDjBTyd9Axb56GURlg9
u2Zh2/y2hcya5814FhcZY8jurFT/zfUcyOMpw4Y27ngWecf79TgYkhutlgzinvYt
FcZbIpMBKnTnP1HP+cPMCYfVm5eNHrPIXm8QNg/t2sY0kdpWMRmTTnQIpZF/xoD8
jLUOZEXRT636ugog0HXqz9NiA1nnRQGVOYiEnVXEM/dr29QU2L5trRm7SzJ542ko
zL8M8/c1Inb7bCGQEq5uVOca8sJvEPCNC21+DQNDn3jv2xi9MI+0BPX+5hNgTR4b
exS+fEGw0EJqN8w/buKv8tIIaJH6lCUXR01WhNtudC6mKl9gB4E89WGEqpKXqmiv
C8zV2cK5bp+jBLWIdV+0GjUrPkd4sEy7cc0/C9QSljtLFCrXtadH55Yc3kWd14qd
QW6lR0kaxfQjzw+3pXKxiO5LWcP6Gcag/AWF4q2L/spsZweSaUHZW8JrORb96WKS
wGs5a1ndry77KKrMat5K2cC+Zl3YMc5HypUjGPEXXNlOWSLej0bbUZ2PH8pwT3Zd
thEUGymTQA27TebQ3XKl/BeNLVa4NwLqKmT7Aa3Dmjj6ZLm7qBmwtGQqNNPxQBf+
N9g6HEbSjegQlGLfnzRz6aV8dye7A483pb0odnyoGCu5epq34a/1cVL9p+2veP0l
LZRk9vhCWQ6ZCkNXxVsrls1wXa9g9eb2LNeacazE8B9lKjqFLePadft/JDM2SQru
WEyYIhjfBGo0Kp1yq4e2cnYMwpG6N2rKFu+WxN16n1O6cHRgzl0U7jua9qZ65Fuk
ash4rXUs60D06apZRP9OahFygZuaUIdRjUqxXSrSBS+0EC4zLWLIvWBNUTkfPnbU
kD27qUiKKHXSUhSN5VTiRbpWO92q2RWDl9WAV6p7FAGFXSTq2RLJa/BHI82anPqg
oyRjLQCjLQ0GcJPhajLpsyYl2JIG0GK9sSg6rOj094asyECmG6/RKT4n8CZEAOZR
ir3wMT9QjqmLKpifcMQmCWcLBi8SkXPs/GxscG8eHiLb5WC7lPJ4k7V3sBRbhNh9
SIh28Dn95EzNsueH5yVpaez7ezDPnmw15WGges5fEJ2SGdD+htL0Hyop1hZkzBry
OYIvqiaWVum5OcNXT2QdWQfA0AIVnjfI066BWbUcksRp+IUOkNgpEH3T2RAYPCu9
VrOeLke8I6ebFfJdr+OBnck8Y+Wetk2505HwKaS8gRd6lH3sBgE8hpxnGk+1JGQw
7uV+PLXbVqakG5E+QLbnOsSgiaAkWAjmhpQ9AQNw++lsoiMhLeSIK0FGKGxpivEW
Hl0uA9BIQamApzFJBc/8S8Dw0+o9UOGB0G4vzzZTiXlblyuPy/BSCVd+XSUCtlGd
HfX+5V+zoesnL48Z0IE/lzYAZJG1/I8vqv5cAMRlKaLOGxGRxnR17oxMbcmW3psS
LDB4UomYdmsut4TGfNL0WgWGd0+7ZexpuZk+jWv5r5lw8Fekm3OD9U+1rfANrRJt
j0nDd4TJIvqUZiX2OwTGKAx1qxZeN63c9Cjg0h28362mURLpXXSVXobFDujnOWjv
Qnx4xAS04n6epWOwaqq+f9iyC+ve3gkLBKQSvGQa7AfUId94PENHPPlhthe3pcjw
1RSV6EXsVKtiMssXfn0MMipfhEre7knSOm/ZlNhSLZCFoJelm8k67mYgnNvDQGHS
yLQ16hngUiAxjQkY73AVuYNNXUV2k6eClyZM7XJYtRnK20vf9vvsQQvrJHmn/Hpg
7CMwBdESsCt6wejdHrBxXgvHzbZlNJwIe3zZjWCSfK6Yk/bF7AECdm9HbOiIG5y3
+EFFGvjuPXbCSlHDPdl9NWGSf3u8ZWo6fQMJ+OOT9CP0bCb3U32Uyyi4pEpWt5mx
5QskY0berK6jjArhXt4UwBfZs5XYcLXbd12AHFGnhXcY8FR7VFAFZLBqP7F9eIb/
V/bttR5+SfCU1SxdWPdo1swnwhDajRzY5C3fmijggdIwSF13eZvDoeANkO3KhQMT
8WZLsS2baG8uiGdE/ChLLgdqzCVyHOYd/gFDTl0m+A/Pd2+OFPanqsEa+wysLuh+
zO7L6P5E+XCHU89/kXNwqLAAYULhNsPk/0hMhWxLXd3oYC1zupdLYaOVCqIxnKG0
/kdf2vt2024LRlH3cG8Xqgb9rEUF3FA5eBchAvlrTyQPqboCYWGOE+hQoIvbQ+l6
g3Nt4xc/ONSP4OKESSFcj5bXLqNu1ie9+MD5frZunexBwf946gvG5j0XRloASP8j
YHSKiEVFtdb65+0567qlQAuUcT09+azCF0jnJqIZLZRjQXEAYh0wQadP29S29O3R
42WX5SWBq5ydjaf8XURhBVGnBpbjxfJaGjhZPqWW6bhx/K36ntTYjQAb53qF2YNx
9ErDhh2E51Xzg5eOxMbuySiv1n4OkSo5qdMyoviYfBvWIQ8ECxRfT6B1ykzvMd5F
T/KaOuEJCWq+Fss+OJbz19OK4cBI9t1vbiMe7WIGffuz9I/UKKrvucY2INyV0TQT
HZdlS3b5cNdg6WEKEv/b/jq73Spy53nDy+g3yR4jrftt4N9BEC21ciE05iveXAsI
GCR1f7xP3spAkJT4j1j1fSPfIBCK3BIv7S+Ulsn8bjSsNrSf00coYtXp6VZ6NXMm
zs4BjxImuF5yLzRuuVu46Y0vqYD0Pu3dRzAlF0sokAHO3UloQC8p5t81M1XcOQvB
R9z7SUwBGPzRb+UDtdBaw0DTRRfC+Y1Bz9OsceCiXsY6L038dByfJJKXoV8VgoS9
zhJOyMU/drlitQvyd1AXSJUVHjecLGwRJWj33jwvW8LeN/Padcc0kUy49shiRYkL
HufdbvzJLvp29cLYVfC/Yv2axfYp82QSQ6QFRFAZ2rfZVWbBBVZvJJGfLVfUSow2
serYhg73Ug3RoRD+bnYngWEb1SQ3KXAHGk+RA4J9x71qmA4sPydGdfyZ6doDLlqw
x06M4FNlXP9gDBMIQhD4UpIEWKoQXPp6Wa7bGZqB+6qv9aM9NmSh+vdp54GeWdM0
6Q+0MVRA1HfZJCn6dgooHYnO8ZIweF269BHWd9iMWA+oCZHm5WYf2h1TXMtWgeGw
wcrhus1qeBxV21jxuQanA/QNRVrGyleM2Xbdqm5JwKY9b+EL8c3QevaR48Kkb/DR
dZti6F0o0xKBm0YFJJjipJtlHfeMynkGZ2WXoMz4VhhgTtNZxm0+3X3akDogx14I
u8Zk9IU+QDzm92EJTtyj0OcbCXrB6QVmc8MiESaMLCOE997HKQVFuKuCqmWlcB0j
kUeAM5Gi1EjUrf2oZbNYhwpKOOOTQOv95EuBlK76/8OUR6bfoAGtleWJILwE88S1
0g2A2CRI/7eK9lr/pUASckqT12C19cwOZM5lYOMK9T9qRv5UoZsOfHLl49kebBEO
YZkkRRrYN4x1vfiy9njo+K/ASuDVEgqOSNJAN1sj6BoQZcMR55oSoUARd37U0d0Q
FktnP/c4nO0nYo0W3UqJlfQbE8CQFOpGKaK+fjADGkHWFei+HNGpKmPS7QrakkWy
DKTAFvuRNY9efRgtpZyOU9TmpVTAIwXruHTmeM68ifRVYYMjEOtBLBH4mWmT9Ex3
L/h3FLxzVm0Fa0tQf+Ak3auucbR1qiyQpIPM8AdjbmzL6DKQX6sGnyY76Injfdpd
9auzmszcUKcyRoxpgAyK7FwgfAS4M+0Yredm1jgKiTlABmfcBPQKQ28D0AXeF281
C7mA82A0zQspP/3G11kkNZIvqpOE17iusJFn2tTBlMHzdjtPcxcQcnLRdxIa56Lu
/PE3a5wNtjg2b6X3t4b4sKNHxQP7LLZ5cGiO/icH3oHPSRu41qlVdYLHx0/PLCbG
1J6uFMMeDepmrw6ENxjfTeR1qoZwWk7oJdchgqdwrqBEWCsxbAWOl2kl0Xi5i7S1
KaUBcD8N7Yf//P/n+Qy5xm4I0F8JDpF8eIfb4ClzPusXT/W7AL6Cmvh2NlPcTKe6
p7FWsnorNdVrCzVTRmuQu7JlleM+xTfeHkMUmHcj4MboquJob/rH6kcxPBuyqmY3
L2catw10cBsYZI3DuDAKhXJ81btK9aL5EaSyVhw+pWz3YHN3PWD07nQqPT16jm6A
FNYmFwbR19DkB3KLqxEUVe5zuywL31cmkxXMSL+Hs+fBbeJILwdxtS4Ay0GDG73p
L8WP3TXnaTWiQer60IiERvo8rP3gYcmjw2zyth/cOVwxDhAztNgc2ruoAHolr4Wq
6sUBWQ1Sj3dS+Be2rC2ZujS8c3HNY3/dkPpWebei2s6F4A7witB3yb4aWSeF1Zcf
7/jkZQUDWUhisogeblTGnkrawViwsFjT4SPHQr0Phliwmhj9b6hGl9i5ASI3eRFe
6odTuYQzk/Q2Hj4cJLTuzgJeGWKBZ8NW+efhCGLpgZbOocOANr0YxDZpQQF4sLa2
XEkjr/tjuOF5R+9REdPMvxmFob8TxiX4Lbsi4q5+Avl0sSmXL/wag0Un2FAIZWl8
ahW/NMWE07sj/9axpwRgpn4Bain0gUvufivOMOulDXU41ZZlPsA5bfBYJ8hlJrn4
ua+4mJ2sVaN4rRT5ULX+WO1wlhwQKzee0rcSYCg2ejo71rZDsW0+UkHFs1f7THws
0FNp4YZSRoN9JSulpi6Db9ZQD2jj6IoZljoli2St7DEMN0cs17QYxvB8yng6N1WN
DIGaA0mcwC3sZC3NHTJE51KAukHc640jcfZbzuydgx3LYxxYAj20CLzDtjTpuhn2
e1ICcfVDl0i1VNcIX7N/sK3VxFuI1TpyE/wzFJpVBf+GGPLFhfO2sn1BzaqsHx5Y
4xCXeOGLkEX6g9hof1MxEMD/A6XodultyHnWGCRKdRAPgDa9z4d18uHgMVypstTU
kctlVIaImEy0CP2/DZuHw1iTTjEnyRzeH2raX5DbPvWavO5r8lBXProMAEGgcZxF
m/WSdjtgYEVN9F0hSyv/nA55vr75a4LXIBfszrcvvki4seOKLBnMH08GIVJcn+ag
jdRx4N2G9jG3qmQR4B/uPefyG34OILugp6IiFzRa6QH7NaMN3sLhgk5IVogaYvy9
4kLUwnfYkIOq/+XQ3SmHo/uK3R9CNId3gf0mT0z0Uakm/x7k84UPTJyek6kOBRB2
mYBN0pyVgMsaRd8jI3BvqVu/Y3olQaU3usGD9xXUGMoLFpNMbmF76orVVj3Wbqp8
cZVBHDJ0EuAWRTJc6LaTS/eWLY+dNYiNsEkdRVRrCajtupbi1KBJcmp6BlRQaCR4
jpZykfXVr1vuezEfiymsJLJipCOccJL3scjw/1fBWgzRxqNK+yJ21EacTDFT1z/s
XKI0qSvnBXyd9p8Cl3DLpf1ThuV6kyVMMbkMF3oxvQ87Go2aJ+d2Ja0a5HuY1x3K
Y2c7Lv1QPR58Nu6V6FBQba8ZyAk6QzyOmbwZjqOnbFtny080kbKTEK7D86sir5KQ
t//NLDBb3MLDvrE7av+BF/CMlho/tc1GWcuEgTuf/B2+fNGVdhjEs1irmRkG+4Yb
3M85zyudgXrQlYoWl9RZJceoqEsOOAFOI5FaVDnec8M7VFZAWHel6ZvLevcJ3QPx
DphGaws+GDqLzJhomnYXB3Y/72WFBPgKYxGczUojdZovkzxZRyt4g694qBmcUUWv
nMmHGWtovGe8oFbMELc7CSqvlNyaxHiYLVXG/baFwswNP91KSGeSgOup9bWwPB9m
exPS+rlzpf+RLPOZjNlj5PDodXVwlZ80mTkZMIdegwYfHgK1UBR5+xsHE7jhTWiX
WH/YI5a6QjrJTn4hUp4YiXAVZJvAl08QcrsITinvCzm6Zisbe0OsGFSzhNQWjyYE
il6NcrTIpMFEPkUrF3aJEW3xbXUyT7964Ikugx06vyXb6sioNSLAA767isiDNhwJ
`protect END_PROTECTED
