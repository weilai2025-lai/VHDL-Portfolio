`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZSyY/juzUdvvIjuZaL1pDywByu8WDMCiA3iY0nHTjUBXVuECknCPa1AvN2NfWjf
GOP0vPcuEog1izI4Hs7OWvAdfLXzxApaG84RJOey1eEkBU5jXXaxmhz+JkKSuydF
Z+NSKBPLTX0oxZAyu/BEGwIScrZfur7oMypVS1wsjYuI7eMA/e67WncNxMvkKhMW
4SFNLDMqzmS+5/CcxHrp/A1aGp5xNCNu0sElBaZNBmiKeSZ0v9fh9lPn/nXJh/cj
E3tlmw8sU6vgfFwDi7f+6As27vxqlvgKD55Rr0IMMIp/zScmrtcAmioviUrj81B0
X70SwaUdQ+rEZlF/kCND0Rxjo3KJQd8bFxQ/h6vwoU/kcx/6mz3CTHYHK7HqQPDS
swo6rNiC7hOLaRMHZGKKCKYSpU65VAi0rkthnNGX/FR0n/sdCskZL7XoNBbKsUQO
jrU+XoIUcFzhEq6IGVtAhHhpLFm7byCROEArx1JmnQOnueDYInrYKIEzmzhmSy8o
D/ynmla1bK+7nyLBelDZq8OLedtxwC5XSVw3l1VsvuvyMgBsJx9mKEPzKrAIf9gS
ZD1CD4u2M4+MvmP9ahkteSRNpRxDXmtGS2Z5RNVLx/8yb27KvtdivKxelaL0LNXS
BK4VttopNNBLX1OGK3npJ3+O/wl+L+jO2BYFwdHQvCEAhPzRboitukbRFqOrX8ew
Ni4C9QLtczsYiDuPeu3tW2obfBJe/XMTmPU8Op0vsbXcd+4rfq6hj6OKdAc2Shxs
nds/gJSueoy53EB3ctuLw81MUdz2G7i/vi/wXHpJSYPS8K+NPA3YggmKGXk0uatT
g02blDNCtbVY7aw3xeZUWspQaU6oJA1VdcNCw81LZUMrV7VMYhBLr54iV3idumbv
7Hk9qeGS8ll6XYFBv/4Ps501Unpk6xm0fozTrc0YfdzY7netckfmG/zH6S/MmffT
mLoXSGWRr18U2im/Leygl/Ete6lJIdBdiRYH1bbyfMv4V84kMeq509eNYKwiPMUU
7xFqYbHDBFsGlOrTRwhoOMYjduGdmAJwKBgE8jHSWbgGayJI5uGvw/hB1uhoKXgC
XUYt7unhyHfR4I0JFqJTpYtMdXLV/yKYmYm89PdVh/Fa8wnp0DD1WbTMeonLhTvg
f9zPXh8c5Y4o2Md+8B2EBda+E9HxD1/OkF27B/gNkFSh3+b2tfvepqVjeJAGC0KA
H/ynagugg6IlUu9BAfUyeNFV7NEdoRAaNvbhWyD/fkwW9/3Ri9wbF99zEh28NVoo
bZO51T7F2u2VVbm7VEm/f/vcvE7sJ5uilLfBwNxe5/57lkwL+RIVaw4m1rEsPV7u
f9R3s5sBCg3ROcWlu7R8T/ZILa+tVo7Ci6stollC3fh3SmuDdzoDnLH13JTQjirQ
XT3U89Zc7/coV+eGStL6T2H7iJhVzRBHjZWamnSsz9y3D6aUnv7njBnj/KzJBy1u
xXgD5b9EA0VamZaRfQHV/czBYVy0opTNctlKOa0d1/PepnlS/1jTaVHoII7imZBA
9LphIJ9X9Mgc3fyvuDQCaaWSLMC31tYD7F+IdJB1I4kDqW4FdWnLAILsjn7Wq5wJ
fsezchD6PhIZXtmsuwTM89J8TLtu2jPAwuGrTcq9mslDjGE8iy+rfkG2qjs3Pdq2
BR6/k98KUf0a63bJnOuJjCIWzcwUhk1Ct57zCU7DJ14DFZfyKTzSJzv6Lg64yVMK
q7dhO1Zj2q/gvfACtYsKy4rbMnHWLIeEB/n6D7D8SEoprvHVWOiGmK7uamEugqGt
tzo4AtYtpyOCeZC6Saa0ugcNOCFTvOOr0H1L0vByu70cyGI7kZ49+tx5X7AoYvAQ
Lim64AJGIFRo1/mXQ4SR/rHsv4o6vbe5xrmGk24nrDYnF/ZT/Wxi1/6XI+dF9mhI
6z/rpMxSyW91d3DCxoLpkaXjiJlFemmfPvQvhjR56QkbLOS6QiMNsrxFT4rxuPen
q1jOd6V0UDzRVvXKjHEqoukvcWK/PVrI16jGdFhZ+59jZqDe0EV7KpvjhSsDWbWG
35WO+S+z63vyeB6lQlGDQPTbJuYNka3T9L8X+GPb7c2Pc1TAUuFzVzEX/3uoggmM
w7xIIg9z+3JBQCB5uBZtbOxi+rTm/8bDUUHXrSyT39Wv0MarOcTqemxcZ0/twQmJ
BqudnNXaodX5e3arNg5EpZX/nIxJQXafemk7AUfEH1WYfJueS3LO5OAYgOciZoDW
R1jFZwRpE7BHEoOe9LhhsCvXeCs9AKfSzhVcmo72asCauz6YmeJbYvfvbzb13wia
12W1ftewSLSRxH0q+ggbokJynM2Wrgws6iMyaMDoawOrzXLD8bj9fCX6Og7Z5bo6
86l2RkxIhVz1t3RExYaEVbPh29Za1qSIwKIWU5DR4CGMuLxTEwToJomy14SUXe0v
CL9X93siyqk5wWBfbAq0sEdYqZx9wxw5jKgWbNu7l9F5I6+k5Nv//HNDCqiK1hRS
Z6eTPogjCGMFiWZdSrvYTIXQqu8gk5Gyut4lCtNFjdULE0pZzRqqPQTYfr5AOJr2
uPy1RzshR2hIIjYNYZvplZHEHMEQ0R6kg6FsP3FG55nGrf83DieeHxWXbt6Ws7yS
3fFdByMdeVwYpN6BrwO+9pvUxXV/nQDKoWUJNJCJX8FOPc4xOnnwmLbWDrxNMEMO
Ckk7x83D22Ppxr2wkyx+YnGfLG5GPc2TNomuFtmliPNorqpPz8TetwKbm+88H2Ms
V5PDTEjHs9q+yfKFbDsfGwTKmFDIexenNy35WtPPh6PWzj6YQ/jDejJPzQIGp3De
qawtgX9DI6xlWhZ099ELTk8X1HfDLXs/YFjcwxj6c9LszyDiq3LTwws4j6ZueVUj
+JgDckv4WnBbdKc8GcJ6L5zU7LFNZQ2msQM1sfq+OIMjPikb+D6p0ujRUY+uFqHC
kU0g6IbBmMny8LEbsLjAmPcsYKZpr4DsoLNTVZM6D8RUxx0uAkQE1PDooV/A9CvY
vx4+UG3Nqm1wnOVnOC2q6Czgf8ZFseDpb8sAdBqj3XK2o9ixJXoN7qZ1MoVHvTgq
iVPzGStpEVBj8wB1Oh8z2TjMygP5i3mLuwtSwuegWGa8DWKiA02S1BHk4NTZBC7d
HfFyGsMIIkDkJjEwCX/sbz6DjrwNTqewQcMNT36TlUzVv7ZDsD1R7ASNePt3jKYo
a2JjBkklzoRBNvemWsMgOP0XIuEhopbrUO8S+AjKrz1xpZsdfO9Em6HWmogtkkMR
MRVCBzyUPlLmR+4vanQ8C/titwNo9bW0mvaPsxNm9rxog9O26jfOzOiV9feBTEPy
1QimuEFvdWeKBqqZNVNEwI+6qDHtjgjiJTCzTuqHS0jPT5Ky7Qfq8kYLZiMDSnte
Bv/NNwnsHQjz7D7vhk+yAOeMnTb3M5tiq/Gq5innpUpB0gu+v/dnT/eozf6mz6jr
2m+kzL2Q6TjcYujCou6Kxg1YnxmyAzF+UyzrhTCcznziZmTsYtzzMD73TiUiIAdV
1KBsF5eSV7RB28ctTCacbV4vHoE/UKTRp3M3BuB7X6A1y//5y3MxL4PumyfXgAh0
S8Sl/Tbp7atK+ZPIYbotcdBECURAbySInvW5XLAF3VlMWvklznWKJmPdymfW13Xq
rEccpLx4zmQfzbPNhR0Up8bO6B133Q05Bj16qfCVr/t0bpSQIZijNFR521Ao8Dpw
PS5X9pRljub0Xm0vaHC/CS/SG623oQdrH+Oq4yGfFdgeS4xvXoNnZWpYS7uZ6jFF
MC8AXqHWD3eRCuK3iYubS2hb37Lv6qJIYVDFA7+47juA4CgFxXkptaCqlCzlGBp5
QRSZSwzS04I3xoNnHk3TABuIQgkMxo21WJCJBC8eHrjxG0bASXZ4dfUGcOIFDMQV
twLSp+BNe/VAELZlXujBx1AFG0e3QK1HJXEjf0WvE1zVLOBMUh9raDSfWie565ql
9OarpDgF0C7/+5FNmUxSs6HCHR2uvH5xEMW27djMuEc5IEf57JF2o3YkuuYyWIZU
EsUmKqOwii+gQk/eq6D44AWXx/tJD+pPLZR+/7rzeBCCKVPq/dA1/aosjoeBOJEH
le0DNVsE3QTYCa5XNEw5mpLXEh7PhLfAKaRI4PY0uuf5uErQ7yO85hQRxAPXKodg
JoK+gBiE00I2jHSbKs/mi0rN1HcW8Uf62G8SBAII2CUfLHaE7DbECbCXzQmeKcGH
5ErhVrF/tysSFHM9ViXNFsCHhDn/JKIGAdxDRPOWmsjAKaC4rCSb5e+wSVZCB1S9
tZb7/gqbBR3vrbiZSqMV2MDMPbQX4sVpf5CUnmCo1o7xjuJFC2XpM8IQESE334w/
DwaaK4PPRl4oQKpEd94u+/meDR7iD25GeIQPJntIOFnD6I6xK60P54RhULtLP/sb
ftz1HznpCpYiaNGBqH78MLZBYZ1QUf17+upWhKqbWHIrGx8MESOPkT/eSd/7/fX2
ZJgHe2DRyemkCdqz3XLfxbnjV55OpMxTYrwgW8Z9zuuOXVm0HG2vSWDGy/V0TeF7
1dnveXIvEQbHy0aP0KHy7UQRff2/djH1ipq688BUvqxawbKvMHwXqbnthY86dzAK
P+TWUKhvenacga9DiBSn8wZrh50Z9V3J7NmUI9cFtK34SfqshHrHpnb2ZBD2zoUd
12znzRIvq3M2k84tlBro7P3q3Qt+dd2P31b+3dw4lT6GBdqfvSrUq/asMMceEqyq
TIscGpLhcaZjyqIPh67Ylfx6lWXwhVKekUK1U34CQxX6LPmvCoSjXSWxjqEwY3Rw
MuqUPcC9uJf09BNfIkSMjp85oGvdzCSXJD9bzji6N2Guc29JNsvFavfhSiRqGPAF
CONndDIjP0xqRZcbt6gRt4zXw4sr7s5m5+WLQTai1LYdZIsqhRNfv/hCXE5zYyxg
qKJekv3QjDgWvoJPqIeqBXcYM3mLkDrQ7G4mRcs1daiDuRT7pGOV/ymcf1gRzfnQ
rZbdjD9JU99Q3WwMWt/83ft89JgvGl46BgrB0YZszeuHHnx8l/388q4I08bo+hk7
t1zEFfj4nIWU6E/QRugjXUhliCmi2tqkkmmKPOz+tD5bdZ2E5uCkvv/0Y3RRf7Zl
a03RZQQXlgGqm26bld9LpeaoMATXDiFQDBCujNlz8vb/tqKsLV28wXsYrCquBgnS
TCKCirTPos0/BrBydThWtCgq2KDpcAugNlznUpxkyTIC4aNexreQmPhGQcOxJhWq
HL+GdW8HFHijPNu5xxrdaM0uT+GtFjKYc73p3h2SlYcGTvYBZo8n1NaKFIgl6hpd
VJ3CMEMYbeygQsw42KGS9o04nMmak1mmAvjFEYQUghA9H1AKA627a7N2kMLW7ZBr
rK+m+ydivmkVWItJWmRYDz2rFGrLzm1Xp8rA445TP49epJAspyPiyDHFK8xa/rcC
Wd1Hv5/z0oecdUgNHXF00gnUKT5Ul2iwr6B2aJoensPJFIFksJtZcv7p5974PMZx
fAZEtNawdUiJ3l7nA3dY6Y6olY1NTZYwT2WL8pPypKVE8X0MARdK4v0oC4iKWVTz
JQw60lgN6vogm49Zorsx/kwPMJWQm1+rOuoqtsLQlzcdKT3jaEa9ABkyNwW+NsQC
KKxcKlM91DEA4LkS/QY7+xySfBfX/r6N+i9AclUS51xy5qDHnDm7qGHEak9rcmNB
DEVEH3y0b5LI/Zjj7zJx+3n+IiC1h0jWmgZNO4KuazOmczTNwgmEpSTBWntsI+4m
HOpd4irxKs0t0lx1N8w5qpNpCmLhAMVcY4gnYns6ZvI7F2ZiWgRORlPwtsdvT2v3
JZ5CVFu7ET5BnkgGx7wlJc8jpNrgJuUqOkLkKVUTQgRt4jwpBmtLON2/NC8QTO5u
Sn86F/LBLOBrYGF3jfE2dJeQIdobC8rHVCbGT7pv4lLZ/JzufsYzBE52qdUkKiQs
co6SoI7TD/cAP+jXQQhk5QuOmpKDPUlf2jmy8QljzNLQ7ttw3YcjNZkNN5MRg8GD
Ni/NNiJAWu0hWR79wg0bBIbUh+0rtKfNEdC6UhxzE4FIzlobunA663/Pczrx9Nxr
O+XQWa0c+oMhEq1HpsVep9AC5MlsVx+qKCIxh2BtJCB8BpeTn090LBgbdcmf6isB
F1rFkFtzcfnwbIOwcXTjlg==
`protect END_PROTECTED
