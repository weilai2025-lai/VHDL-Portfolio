`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBl4ganOWAby1J/5UfoHvSWUG54KjiHbIfrmke81RQmEjOmpJhGz4jaJv6nGw4Ck
jH143ptx8/SRaY3cRZ74wYVQ9p9wv5JVDL+np2K6dZr54U2sg7XUf/IFlC6Ur8eN
pLX2jBAO5Z1PYf0BP1z09P6xfUMOCWduVM0DZXqwOY1X+tIYR8JhSSMuMJvSXdEk
SUIn85qJ3ul+oUA9TTB9g09voPnXuVl9h00s/wYT6RN4ubq7WDKJyADkd0XicTD4
9ewQQ7QioDDaH9WJFtUrz8wMquWjVjDEwAZ6FE419MI1Gown7gdMsys/sjjHL25z
FBf8wjnAie17e7sNgUjVLLq9NyfsrgO4EJnvtjvNYlLc40cY/uEpZQfmXM28/JQm
Q6ruZYwd8g87Lc79m4qVt7h7xQRDHpIhNhXWj/pHA4gtSfHDoK5Rl0Nevwf8mR48
TkXPvD7uLe7+7IqVY53bRSvVVagJTA+F59m2Q19Cejp8Hg2+8wsOq+raC6Ny1cNU
SEgeia1DTeL7Q6hT8V8ndDE90ARC0Cz/bTSfd256vcrU/QracrukyiZDmINiioea
MuOrKzGbzaBovZu9k6EN+g==
`protect END_PROTECTED
