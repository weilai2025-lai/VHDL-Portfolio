`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YdKY0/9cLTMfSfJp7KZ2V2Mbunu9vy4IRhjW5F0RBSpD5O5uyth8vpyQxxaItUk5
+aarpvtogoW+sRy3F2iOxRRfFBLSM8JAebpUlwEYRIibsyyORuJB0+6zOCw/hj0n
iMzCdMQRAAnKV2g7Dchpe1Hj0UdDl2q9rLDUPBi+TMF2Y4mWsDKLpzz0h7du3qcY
LTEBvTdz8Mylkq/j0UW+vDqcE82F4pIlWq6w27mfx1cnKQH1ywoLpxjQSaCTJsU6
9zlOtEEYfYTlHdYYlvIYUpzBI6iSdQx0hlfUy04HPXyeqE8LBO+VWFxod0O3Zgvn
8XCs5IPo/fb2naPBozxC8XlWQ5Dakgm4M88/Q4Y6jexZd58/2dyFdaTY1O+rD0au
IpOtDfc5w30PswN/Eghwc/T3GBUFCItmFr+FkSPyN/wgkocq3X4l9vsD0JAB0Ae3
sA38dKkVXLAlUpQj1Z8R+a1YEd+y4DwzkMZqusC1UQYaLLDYCyHHaCsAEGABMSIn
zeChXZw3iQtzg0VPESIJ6w3bw7kGc4NeJLujfPOSg5RcP2M/cC/W+D8+pwfnr1+e
prl40Ah5Cve1/pTxCkXKuNR3u8sFbTifju467FjpbCmCBN3erEL4PQ0C8ZbUWzLP
Wq0FvMeZRHemirdKnFiK0oJ40f5PMvHyHT0I+ij67+OzjTLpVs2ZXIgWaq14y0f9
f0eWAvoFTuh5AAatvMUBzo69VDtTyetsRoPT7/JDmR745NZ/Cg34NIg3q/6DQczL
J0MVKHxogdhHrP9ZMJXpnNAp4BqcYBAdUWxR/tVIt99xkB450pTamvzX+/LHaGiC
UpNdzackxS7kcnDK7HN9o0+KRgrqK0KtaTXdvemOvPqQqV29SvwtHbgwKF75JYMX
hJ/m0r7OeZQ7jKpi5whu7W8owbmEtwxC//ZezG+AM0GXNk8/C7Lo8mMWP9sCxd3L
ruPhLTZvzKgDzo5sePN3VQEcy5djpXhGZX02PxwXiHTRHDxn5Vd5pR49AB30/idG
MW6y57oVoBYoPvkLc2ijx+rMB0Ikz4n0uSiGhE8UBZnWU/HMZ9EuXkPTWoKzXjjp
eNXNroPP/1cB71jGWZt2VbhZrmzddRP5de5JJcLRiNNXpu6mxOCwcs5kmnNwwH4o
uPEsnZ41EbNZLdPPhrcqaVtSRSGMwmxwrhVJacVXwb6bY09+9CtJoJ3oUMvmHywc
Bapns6ua1y3ypKM66JbJS86Uj/GljTIvjz46Vm5eiRb94MT6YTgEYjGqOP30g0eJ
6OHgsDQgQ4IsV4vAmQkVb8nRTF0dTF4eH6L3cPOkyjHPA0vT8at01qHOntQTHt7Y
dfMU9fGIVUucC61kPmZgZBW038THFTZoCHxrHeuqONJ5XlyMfvxDai9Fo29MBdjM
7JJE+M9eCCzQ7gfbfYY3yhqC0ADUJkFykeOKxoDsIcymWpe4KoxpGm272Is4f1j8
VAip9jeVqS7aiaujApGPYw5REDVTZv5+SGrE+oWv3lsu6S6MctxMlu7oIbLdlgF9
CghqhOuDzee/TqfWCoVeKOkPAKpWbZH7+KWV3K2zSSWT2bcU2yaFxem7D+5d6eWE
bcQ3DcVXGPBr/21OumGENPY3QsS4Zpn5calcHRgvKzZHwITCiv+GSNPviVCGU26l
RKm44fXzbkw/YL/yasyLqjWQWko8x6bdk/esGVoAgB6Rh/jKuITxJ7eQbG3zPVns
SiI/P4sPDvyos/y63g8vqzxzZO3H7yb8IWmb+N7V3CoPelMi8sqgOdsw+8Q/6KvS
4Bvm5aEAfzf9k+GgdWXd578saYuhRVBbkPZoAjFvcr9Csot5fRCCBaaPFApKRRqq
ggpjIuhOFiNc88DC4YSnFfGY1l4aeQB20cFc5I7HVWD6kWeOjjX9tyhQtKJfZEUC
wkQ+ZOfNoYfoUPCdgWCWjRIjcaIKdd3f5tnyz8BOl/ydNsajR5NMcGgLIBRA2Z2x
mf3+b7hfQd2aZjIzjCGBHOxqrK38Ahu2vQFR/PwktjamdESqKM4OVQzCz2aPtmDJ
qgTwv4jEmPPnvYlNzp/fl5AjtxXmr/qd6AgUsLa5zrpQ2VPaf4v4IUEv3CzpkvGs
E+ICEEoeCZsT5X0oXK5Px9terHIhz+yIuX6wv97sRWKSOAghIXwQNaBFoFBbBMUY
IPEnmQ8AS+RDaHjf35steBg1B3YqVt/76M5r+D1WgfYTghVQgJRlEmq79rOq1JmH
cY3yhG0djIiu0kjGfY/10m54caIdWQ884rbVKrQU6ew5QLA+PHQVJ0MP/zw/RkV9
9KkNg9vF1ga2BVK9IbemSeS9RpcnTyNeUkuTQ21Iy4VGKskhuQmgKuGM97GMGQ8W
xWg3LjaqSw0Fp0Ml+v33F8UE5MTP5gSWKMc09Cowzok3GGQSXyBLH2UWQv/e1sgv
U5uz53eIuSM70cJB1fVNCPqvpdCwz2L2ezM6f/ci0Sxq7vDLMf2nJahE9HGX5r0h
rOOlM0ScT2RiH62vYJjakQ==
`protect END_PROTECTED
