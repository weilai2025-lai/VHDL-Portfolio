`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bV/9wi/WT8c1B7h2CoQVeJWvG47K12xBcjGN+0qcJmczQtetTu++qDjVHKUz9QDD
PAKLpPEVlkHwlhCIqMGwte/UF8ZPXlLuBWJbQZFiBnRvkFW60HNfc99LfEmbD3io
4Eq8MuZj7W1r5XinHlPQhNf9AQ+ZQw2LzKRgw04d/J2yr+FvxcKJELe4MzCO1zrL
QHsVSqNgk1Lo/oavJDTyAy49HoyKqAT08DNUXX4WzgrP1tHdaREFEoZVs4j8TY4W
q+r3mVdXdgxwVajWgqQvyGkHvhbux2DBjTCsDEt0xaFwTEyWSmAnSkdoR8aVmrUf
zL8bnoGCRESy7mEYkT1MQeCAnxffNdEFQVJRUfKM3kmVcyiWq0XrwVMLodfTzH5g
2DqctyV9tzWka77lcJhEof2x8XFyOoh85gLyqUqMF2WBBaKPOPWtOTos9YIkY3XF
VAyjuuRJ2A+lsZg9PvkE2OMrLl93QZfrYAV/RUUCAv+VwcEx8P9bF3Z+od0aEVfr
yrl3rdfC+bd2FYcZBo8cTvGtRnmPZAbXKHzOPPowpZK9MKAFvSTC3HPVupisrRWX
d822NmZRKbDeIU2QgHhKZmjNwaZudKC8+cywG9czuQ5rpxBpOq2nOhjytrZTD6cx
/EW1AEUu05MAHIsZbn9Jw/XBvXFi5JM+j8pEGMESm91zOQMLLX9hwbXfScf6lB/O
djIRRB0MJa/8pyzxFaLjwOw2+Wge7VqbcNXx0N6V8ZfrsfX12rBrykyN3BdItlOh
MxyKPmg59h3i/UlViYdLR5QuWBiud3T9i7LBJd2ve/r0ImOCKyNfgRscDYTM5Gwn
rHcbmaJH6sn1NquemHJlu41eZlS50Bf//PzucKTipJnmgmMli8yF1IexLiK8eu7G
rx7GJ1lUrnpxIGfQQ9FQPDTO20cBOe6lxi3Od4dz5c21mk2pDDvH8zWlfF3GEjbU
QmS3kwJdGTV3yY6GAYO9mGa1kewOqQzLgNaAUpUlOtncoMqwvaIKuEc2j+3TxPPJ
MmAEg8Fg8INlfRgyRhBVjSjyjgzx8fzZaqYVe1ScKaKR/xUmvkGyIznMWFD//zHj
Yx0J62ENbKA4iiF9PhBGMTvlQ6z1kNBykC5/OYuoksMTtkXHf/UoaBtxe1/dNE/+
WXDCAT2nlbITYbT7AatDyu3XcJgydSvHlZ8NpseNNX/AatLhLTORr/iG1DAZQJGt
R09P6k10LNQoqHZCcjSzSyjv7v118AqMG9tgT9s8IaXc2G8FE3bY9e5rE/jYchIu
zb5n6/RUzF0TTbDXVy5DOFr6UQsddGPM/M4lcKaTbXUp9WqtzIumOlwDMsiOfUBE
3hyn1ByyZqm7THW2lSFo0BBzm/AUNCeFUusYlu+lk594Ux9mOxnLLzl6gxWU3suT
Ivy4Oxc4PzZ2/xsm05VA28/fHWmfRd8MV0vwHZLBiEyAd/IPVD/vDfE5iCbnI8FH
6NDQhFe4LUMk1iYDV9gIqIqrsTwV6q84DHLvlWNjOnKN/opjmA01uqWTMx7s1qHI
j9DCymr0DAJ6S69pREcJV1jG+DDKGs3pK/6zoSdIEyGa8y4Vr55WrdLTqFS3l51I
Uz5RMcLi1ig8n/HG5O2I77KnmOy4afOx/gtY2afemokDs9/PUBZR4Wn+Nhpyun0d
noqqcIRfea2obbLiGQuehpleSh825+2d8okJpkfjcarRsu3CCrZ4uvEYJdx/zDyd
IbCazxXMt+4uo5EwZqk9jP850Bk+1BUDqmnIRMruxZQVhg1rgFdrGxW0ETZ5lS//
H+CUgvFh37ZyGDp2L9F8Iq7PO52zAzZvF86Hj0s/FhT/cPgDAUj0LpZrX4idhzX8
3ycABLEFLHRlHpVH6FVu4RcbPho8/9oDUX+q3FBb5GROKpKgdpEN7MDv6FQQABPp
/P2RnzUkBXQt/gh/ExubXGnHWbEVMQZvIoCpginKkfX+i6Qkg94NWDOXmOu+ADrZ
f80bZ2QZnheRFD2hoVQm5XLyNNKyhoejnPGixiyMHeJJsk1tpNKuZfflNRKIvNZJ
u7+PeBvodtTgtxsJIzL9bfemukINXpssSQkAkD4IAG31gJd9itja4crcmfE1TSU1
7/ijxOdrLspqJ6177iyw2XnlqLw2uYk3h9fn5JIsc+l9gFriYiWfkYO7KMhOftI3
HyOybGK9RockMKJzT36nEFA51GrOLFNcGqaYZgie5IlvCjCCiCfLM4rvc7c854ZM
wQJG10h1mmGF37freoUYoZRrtUnyOv3EEm/C6kiWNlXLJtb4nLvEc5oJvjLqPl/l
0mHpAK1KO3jQjWu3xrPnnuqMxEVEKbgjTTytkuEy3UKYPEVpjp6Lc7GjlNvtWVm2
/DPgFsQY+jPZe3Xmw8O7Fel+GGALJA3KifH+ts+41g3VfwQWAlXkwcMNrnpQViPh
d70rasAeTOydvVye/beG5Q==
`protect END_PROTECTED
