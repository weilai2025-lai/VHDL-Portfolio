`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzxlPq6emDd3NrbJZ3Jrs4/5Zqq8FxunWYKi5it/CS6MekInkJsq0uoYCoMGSI3Z
M4kS3KanuSSwx/V8/yRdvUUIHb5SbwSZGEYpBJoARAHRvUjDf1BrR5au0jJVn5hm
nSanLx1qSqm/X9JR/ePQ6Q1mZoRRbQ6UqBWbe0TDctdJKYYcfM4xkiBSaEinmc+s
jXL+hIC+05kro3qRbz4bO2ZRL4CM2XQacx/t+6wF4tOIJrSSN+YEdJGqYP6d8Wjl
JbFv1gxnc5ta9FLV8/Cpk/zJCTUaXcj4iFT3+96gsh4P5B2uuzcxuck8b3/zaQqB
W5QtlGCBCodgzHAxMX6y21f/bj2wdy6JmCuOC+0UtMswDO0860RggLHj8h1g1R8u
5T/LW9tHqeliKtPmgDWoI9lIJ63XTmVboSVTyZB08BGoJw4HmG4jVTAMxrJvGfQu
ybq9vjk/5AEW5qG1IefghgBopjsbTl/fMz7WoZbI/TWcdBvFaW0nyjnMmtcK6ETb
fJADQId0mFdYLfg2+IX+KHinDNZ2+f9I7kJ1IYLysOymXj7NBw01gzlDjxcrls1/
cB1bRVB/FPLu5CaVzePhjzak024VJKX2oCEBE9hTqiIfbFwqsUs5dYlQDPsC5bVG
SeSG6b4t8vZLs9PyhxBKLFMMOVQeW0XcBRwimgL2wxgT7tDb0gDRhUUtrTOPwwsc
47yIQpY/RYw42XoEpqoXxWXP5Yih3zVXpLYmvouA3jlngFVbO/X18ury9OBxGIhP
8XLMjA83GfXJD7wU7SoWwRG6XqGFNQe8bBORUGugviOWejtQHVcC7YujHYezq4yK
vwJrKqlZVACWt7YmFs6px/1uNh2I/qIXDudyDcPJnOa1TUMk2QrcrexO5xHpILi2
nLK26ZrSVdZPh7iaQgjkBC45Ok0LKNZNDYK1+KF7bV0FCOx67NEbQ7Rg5/R+F9kV
mS7lm0qsZrVTu6z9ITZtSMvk2myA4kR7bNs6XW3xKdamAmLIrj5HPHlN2ctNZ8rs
Ji7z0azMMuJCqhOzCSm3gta0EaUM0IN6D+GHcbB1TF4DOXposPyLbnRa5h8OVNvm
2sf4SPGyIQoRHVVbBEb3OIDYC1J8oV9W05pAKoWieWfRBkdKzPKmZao+RZrxUebe
Mnk7NGSzQEMcqDsIxJ/BhW2YxFHoKK5Fc8Qixyh7Hmh/r4yILA8yGPRe6zQ92BKI
7crHGNyvyUKU0HIwZZOanyWOG2czAUGVerGOW2uokQBXn7BIlLBloNC7+SkxapaI
t3sBs2IWhATqecogexAbyW7vSg+kW6qdDOeFbG2CjN27JqtA1Ijr6vuoQvRiJMtO
McZSN0UnkmPCciLcQhO0G+nrb7Lv++1cwZzOOyP2q46f7a/6qkVwH39MSIDnuBOz
lXn52Fw9WUR1uHmaMfFCKMNwkzZvJRtGA7uwLqUDnxpMNWLa8mx4hwlYp7vSqi34
YmBOo77PXT4xhg+oqEDv9piIy0nA8T0mk/9tMtF+3y0DgKVCiCTIckPwFINvWxyt
qs3kluvMDcWa+rBwRTxA/QExkrFpj34md7043G1q3DtMWEsDhVWtNRe/07bkG5mK
0YCapsBdPg9LxyagHg1ayX1GHo3znxc7n8arJa/r3gG4AsgiTV9LsRorvBu8F/ay
+zG+ObrDVDSHMS8JoG/ryNVlFh9B/K+vQvSuIt74vTYUqS/7lSzCkHUyL1Ex+5M8
4trUopCKmw1xwwMe9odUEWkKWjtfZ2RayohmcUVGcbWCk83DoGOXja1ieC4JSfEN
Eavn9YNLBP8nCUQpq+yoEacFuj1zMCmnmAc7NJw2kHWMNAUMc/OQYpR0zkPB+/yJ
aeY26TpiOMhZSxw0rlLUiZs4ZdiESv0Z0RRWtx1uX2K7xWrABWU4ZGV8lRfoRsWk
4Gks6PDLZ2UJHz2RXdJjxrWezM0HT3+JhXmRSM+Fc2FhchIvcQ5LbUerM+T5coII
6u3dIaPG9mRIYbyRpXyCEQ8LHNLaNVAp8Bv62ojDHEfhMI9A611o9jKWeIK/Bi58
BP7BZMKif2pvAUiC16kJjAORSUNzfQAUwl+ZXiw1Vo+Q66zkF/74gKK4AVIxk7o4
CXQggmGY5nG3ScPAQDmG3JMWrvzssXGf7GgpCXgmq5aiO+pjjaALSSl5gBYKl1SG
zrpvHPsf0Hm5hSHgSztzcbfYqdwdlw5rU6gSENtHGlwd2Fiz7fvkpoNnK/bXHG+/
DKkPkxK/OyFpA4mQbtrI3XoSPWso+oDeeCvnHZT47Cfmfk9sLLF166w0lVmDTr+N
hAeJmZgjBot0VjwKfx/IegepFMucaTHLSkQF6szIg2ibP4dynZTtUx1j44wtryKd
1CCOYGO38mHyduz4plgFeap1CFt3sdkNKFG1/ydiD1FRiHxEQ+vEAW1ZWblwGN7L
TQ6am+9mEfwWEbbDWUB9ibYYRkxrPxX+nQ0wvjRmsL2qTQ23ybSKTRihB/4Vqj9s
3DeMz4MxhTLP8sMvlQR3zB3Dj9qQDGXx6HodF7tlJNxJ8gMoxGyDnwoZEcLqnbDp
J4YQ+MYOXUzwYjOEQazkFxHcnX6Oz98shnMll65xaIFrSGaq7sXGDQScC0BCyAZi
/J4bBLCgrEzEmlPOvK5oAIa2dgLOv6pkC0sSD7oEdAl9MlbVAl2y6usslPQSrZrT
BPDQn+5dcpfIoVrz+ZPwRJcJe6mo+WlQmAjSz4LSEJvQ/HFMK8N+qPoq4eCU3eBA
M29uLBEdENjKM2h0c3uTZe8XemKehWAZUe1Vp51URMthvDYiFTd78jodTq6urVvb
rGbNAlaH/km+ILUQCVtnMsNBNwUdjLzCIczBgI3oluJlBoaTOk2PsAogvlNJ5c8O
Ln284HrvmhqI1HJgvGRAPCXRc+wOO1+EYmL8+Ke3nvYdxwy6JG352dZWSfp9pBIQ
CR0KXhYzk9g/Ax3rBufkhgZmP1mrd/2pQqIuVAyN6owcx/9+ypckhUpXddB/iXPA
JCWIELVTy5QDuiShatnmIaRGUch9fSLk1QVSXEr5df18fSULkG+ceYFOVcJm2ZDR
rTKZ+b8C/jbWTY4AbdjmzpCeLvrDpJv6lJbv9Zbx1lPhaWdjjFBPnUrptqOv5ex6
EBeSqP1CLwn+j3j4yXmi/XqLyrm7+XdGWfX7o8iZAIijQ/9ZHoFLPEWMYB0BoHpz
CDZPvoIUfXoRlFv0ioT+n+4ayQ+7J3do7zoHGqFQubfPmy9OCVhonQ28+x9GzyPf
WuWDJayR/XrSn/CX1ZWEWugr/nI8QIw6IwoR/tVraPeRI3owI7Z50q2Yq3wZTDua
XtzNsMEUWvUm9pZTjN+zbtYyUSMLyWluMscqumZHhrb0GmAxvDKCs0z3VAgYXeIJ
rnl0nZb1v9Y8yLZDriuiyMyW5xeoaRm4zVrbqaDIyYUVB1Oqree0NFyIUuDq/LAY
K7UwvisYFm5sdRWDqVDM9C+UoJYqvv9J5OU+8Z7D0tFZBPIibk5C8mOVipGC30wn
QaOPNjU170+xSqUpp9J9jsg8gN+/6NWTAUba7iJCGVx7poGBBtZnKAwWSfNBliKf
jR9oDko1PZOA+5ru126kWIJoIU64F9YjvmcWyK7A3o8+IeXi6YirjNzf6c/uJ2aM
oOCU8Yi6UqQfhmnxlYgsPInSS51af3bzQWbf5qQQaHaxTidEAYlz1qVHs/wzc/b4
pPXKtRIz6mYoN3FMMaWEkS80NM37HCcMuvNpT7Zqc24oHOCVUIdCjgIJDLVPtW1p
LMl1BgIZRkb0j9JzXCExneG/3wfDtSXA00YEFTucVUEAG8DQTFThpBM5XsB1nea4
F/yO3TkxtF0sp2i9FmPv71Um3yUVcYCDo9be09GrSup8i1/esj7IGEepODMcQV5s
ibLizwkWQlrNNDX+dvDDFblf4OgsJWXRzNBir9j/ybut96pbWPaSQHA7gvuqWySd
4eYB5cmaLAA1ZsqmjW7+J0gKLIz66m2gI2yfxBh+cJi2LUFPm2MFFbzmKZsnxZ1d
JOm3h5mdSMjxWx2169VfjM3JYSv5KeLqpXWC5faxbD1ijPVKrdScXmu6pj11fGJk
ipLfTf+6/IwiNpl0rc10xa6ZUGgZAbO4d8JjfYsRZH/wqf8u77rAsTUeLHId1B8n
yH2JTIQy6XcMG/ej8wq1N+XO1+f0/GVa2bSfJkdOWM1o+rbNsEuVtHT2NuHdb+U0
KGeI/mZydqijoc/hy7HbCzRZjgP7ODlv4S8STPRpBtoXBnV0dfK38FytrPYO1uJp
k3UwsUIXYTF2YT+/xaC0cAXbZC+ykIBPp2bxknoZWiZUyrOezXbzati2p3AwcSG5
66rkTqXKeuyTYhwCAwh7UAsVAGmf0ubc4knIRgUh/7UOLK9v+yIwZ46xZxIfDmQs
GkaqG0tMndqOHDFgLZnewyvnUnDt6bGgE1BHTcsy3PpZBwvTCqtmSyGSZ4j0/pvt
UKcgURd1C6Sab+eNUmFxpXLpoTuxVIlzCeQVbDVew425kwBO7C9u14mxVOrVQJqp
HWUsOi2/GmOdu6x2dTQrO4WoWpUaHxMSg3poshPOvXYstJD+PKRGfhk4alsYoPLl
`protect END_PROTECTED
