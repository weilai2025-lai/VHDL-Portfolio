`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZCNtcmEwkXKcJEPffjVDLh4CaquUGi3isq7fDH+QvUhMhZn3R3ZcSVaTnpvmJ6KP
mF4S16aTABCwDrbknIXnHjmDBeM2JgwyQJ8WvOqL2fVbaCKO4qTxn5plRyFOwqGf
QpP/wbhLmnYZfzj44iVKgYlOFAxP8Xsh8V8liRcV9XMgOgj8umVTiWyjxUguSkBS
lxzzwGov3+ieC/pmjhQLA6e/frKEdXvx9OjP3bXy1DFsFAYZBj5kRG9WVL4PXtOW
XYdBKHXxrdKvez70l+oR4koTjwBz5WIUSyw2upNFNjCnZcNRHLzz+JKxXDsf5EDY
13bBzNfr7UVRfb/N+cFZW3q/de4XPMimW2hG9kP90ivs9IMhxZnI44kjNGUKhccR
fD5qp1E38DWndau1NtupfCEilV3/gLB7q7anOkni8/hr20ijPaRZX/yv/hsUsRws
a8YucXhvEcgO4e5gF+AcAVe8g3aD/72jlf6NIiIOXCOeyExAvnNGxIXRrT+XM3Vr
VMeDea09g92Jd0QcnoZypDtuDzRkNqW5pgqPrigkopusOTCkFaZwSzxkZiQTQ8J4
HcZQjjRqpH8MYMHXqD+b9gi4kZwQbAWAO9zfKE24U1hUZXEbAjBWGgt3ZVgTrgT7
QtSJKbIXqsNfgu+22saJdXUNVyB/xYLEGflZ9uUXlK762EQOkBupmKTtXFICB8Op
APH7XY+7096Iki1ixStxgpNYLHvQ+CATGw56gstEGHhtstfUdIw2zVYwHcf5vt33
V+HEFh8Ws25FSVVFHrd7WElzXYAxxHB8dZtbFn2+3lBzKbY2Dn5IFKlW/hr4YYt4
W86K3A+aECTIRF4HIhphxl5rcQK2mA9JlO0BbHl+Uqe9xAQcqOzRSoGYHNNVMLQ7
y2CfkMoemBfvGnqWK9LScQKw7DO2pmNpD4IkHR+3uv/ekTUvE+Q3IXLDf7lApkmE
lpQuKu6kDj7tTejvvj6WmYqzu+FgDHB4JDIL/ckVv0xs8ctzC4UKsUk9snDMSUUU
gbyCSb/+K/C2ZCwKLzIWEt1IQwt/CqFOYuycrnKCPT8Bu+OHPIhsesZzRoBlD5SK
BpX5Xn/8WjpFVbCTeZPhV2vEgY6DgBdR9TTPodBHfOTLJ2y0A/wuB1dAU6tSaClb
TlYrZyVe7DZtsPXmfiYFULIFf5jEps6xXxwEVPVQwmep1nqL6sc8tA7BO1B7oMaJ
hd1DtqXfRboXnf+l4Y/87sXS/Jg3TkGZz4/wCrAXIlQ5/VGwJ1MpSmY0C9VX48dP
ZH8w0PYVGKC4fSZeqTdy/Hv2YrPgw6HpjZFqWigasE8PxhpIgQwKE7sLris97tVX
wF0Sl+Awx0bMh8OPY/PzJq3IjtDWmUDW/mhw2hnhamL2gB8wy3mKSCqbIqdIM6B7
bRLVfmYiQy/Lid8hYMjgo2qcY6nq6bWU/kU0I7tAFeEnuSQnQ4AtsPRcE/MsZr4Z
Ali4SlhzsjeD1h8bYcej0CPnj+BzTb4AZUBVpMVy3vs1quCtV/tYw80F0XiIYkKQ
yAmncREV+u9zQy4AqXEU9kC0LX+kjDpnBqFg9vbG5nnAvt5AmhBdbojit0jMJOza
lGfkBPye4sraQZTzD1YYWzM9nsaLNI+s4qR1Q2jZWnIailZ4WSybUZvVSSd7OroV
lA/ik9YT7Xv97c5LNR3QHLBYbE10OwZ0O2S5ADLLhSvhsdAye3K4RvjMtJZw9lBS
PqIxxGLgmqbiHxhKUm/mS5xY+LQIxV1WQsXcpgfOc0x3Az//3hClSkhYSPULtsgB
tshgUhEWmNMhfeAAL+YWfrbwcQuI9uSaQEBzVsKwixntP+pQwTnO4fPeLaWutEls
qU7pq/Mlh3MjHwqhh0GyyBHL1vkefxRw0EdulfXUqrztHgQMM5NWxLyDwdX1P2vA
02aUfqe3qqHHz6D/eC9dtsDy76aPmSe94RVnMNuoZpW+BXNU8b03xNRDD6kyAqBZ
Pmcgt74pG6F2vfAGjDvELCHz89MCCpKTwcS1bhYqtQl4bEf963KwgbMDsWhfvjZZ
0NrxOQvv+roA7joPx8IhBWgGV/pnRB998+7dwR0YF7NSzSIsE2dB788pWaaGjlNg
LNiZjURhrD7NfIzadvGZV1RIOJTaUt5xf0qic7sTJbc=
`protect END_PROTECTED
