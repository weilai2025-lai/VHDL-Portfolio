`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8JXvFoaBizLeHCvCCcmxnJcarZrnW498rI4J60dY1T947mYvtHapXl0BxUCiDkb
0cl0opcfVbUgeQkRUwushcdb5xUGd500I31g2Fak9cYG1JxqWQUtscjb2jnL0xc0
b146Jy2HjP6Q6PzAdnU0HQdVmsne450MC6y7jlbhbO/5ibYdfVIAPQuDjXlYPmbb
Zd9T+jygcIbLzNILGplIi6/kQu94Ae/tOg2mXJqt/WtqWhRu2xT6S6JTe+pzNOnb
9RNMCNs/tdff0Asd00ceMYhIb8ZdyEoXq35Ar0Zef0xFn4IZdAMA4uDbojp/x6aS
xBhmwiKGxVTuLW0XSnorGsTOEwt+DcKgEsxL3zgWWEH5LE7Iq0x6OuEGxtXctcoA
Is3ybxF0zab5fw8zYxhwg7jfgDgK7uyAsqp+lzLfHQrhGL/4Jv+trHL4lNZUMxVX
OENiSSYMQkxxmomXJkDU/hOFFODBsgDavrkaNWhWiz2ci9UF8nSGyFpPX+lzcNVC
0qB4QSZscoIH2RoAI1F+zHoinO2i96/asTAzoZhMziXnTo7aKub18Zc7ZoetZ4yC
oqk0s3rKpj5Wc+fIn7AXfNztZIzWF3/J8PlYlJ4uXQYuyfXbbiU0s8WHodHrILie
DyTpY9wEO5JZkL6+n/dtSXUS6PTa+ig0vdJb9tgaw3D+Q0gUzP+A/FfM/pybe1vw
w1INTETyNvOZiPEh0WQGKOJW8TUEHlSx71vANrtKKRkLv5wUozuKFmICzex8sFYN
nO/V+5FsvgiFNXJaukgINtZChMxEi/y7EoRp+ifLTLkknaN3UvjuTsnvIREqCaPP
IO6cxdZlMdAkX3bGUKWap0xNWqST8KXk3F3JOiZCvU0yUzLjU1uwjqLr/DqRiufK
lwkvHFoHJ6kb2/05Xrj+80kdLJ2+iP514nUCvpvf3BwavjXuleha6zFqQ/2BrWUy
W0TulKROJCqivcOVK2y1s9ayPt7glI5+YiVvN5jS9fRvDpiocSin2AuYmxy681qq
Mg8SeliKX8QyP4I+jPkLdJQuLc/cs59re8BBA5mHcjHqtfGtFpR63KNXr+Ydyo4T
IimZzDylam773Hwsj1k8tIkQpFhYNtxpfXhR5+oxVLm1cGsVx8S9DSUtC9QNRkhj
LMLP/4mJIgjE4uVPgIduvlEsDrrOo+yQ7jGlV4cxPW+x97xWytco/Yli4dgNwmoQ
SBwcsG6skEGye3DScn+6w+4CBmFgTlrXsWfdK0M4VqOFFjyh6qztkmStBNI7ykNr
93zIkEpbGLB8cNB61zO0mI6cBBh77hCadVuXYIwohOah2/w0AB9sV3ECxLSrPfWG
4WaVGUnWucRsqaedKoq/Gij3EgBDFLbcLYS/l3du69c11EBQO6BO/ezWCaVTwAih
A9ex4qMDOteVa/scLsNV2HL/+L/XDJ3n/ujMT8/ieiH6CQMyeZZaV2Ndq8Qp4k05
sg02kiZuZuJnr01cBXaUliDLthkpZGDUZ1bfK1OVEo39tXah8lgvPIIyjeDpC7J3
`protect END_PROTECTED
