`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
psRf6C7/3Mu2zhhusMp/vO3gD4CjltetSlrZ/Wj4aazJjxr3rcv6AdaMOfu/oPLd
yg4+VcUBX209KP9HtRv+l+Z/+8CCLH2cgPrx8C/NAuxRIoaoALsy5MxjV9134FeC
J+sOHZOr1iHuviy5vNLPJZhKTY9yHdkP+9OrDAFyQ9ewxYDTWOnRdk1l6LrqOnxc
c0rCn5euE2PxwTv0cNzyg+/z0BHp46WTZhj7sJUYHtjTwHQbdMMjRny83N3sFjdW
AEdoZ+sgUK8PHXOyq1ukYwhR52TsALcRAQQHx4ajnaAN7q4UHvP8MjqJwAMEtpeB
xFpOimBM0r7iDjjWfsrOPY9OxQFoHgyk8Oml0cm3C7VeeE6/7YZCBAWSi8P7BVtz
YZmv2Igzb2N2IN8O2D3mnI+r4SN7oUt+Ii+U3JgTlyhJuZeRpIkVcLH+mIEZQcBj
o5/svGI+xc7ODw8AFCwFKyqQ7UpZa36Qc3kfwqAZN1Nwy42hCVQwT3VxSZ0mXttA
7bverhSgYUBPPbpj1RUsgGOQLWF0VRd1Ws1BfdBBStmGaa+1JJQb+TXy14oyie3C
0sYP8+qmfRi2byB1yT/GBnGJrb0f4o8WGevZabe7rvbNiWp0glffBXYDWs1Ag1EJ
6xsu9r1KHdjXS03TY7c7DA==
`protect END_PROTECTED
