`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CK5SZEyB2vwOqVgZ8RbBUz5UWDPZQrSl+BR+Hbp5AbeX+zY96B2tcqcoyLqNHBDJ
+H19/2Hog/wfitSQ/VvSmhRPBcRDU26gWwO0yFxpNlCOEm1T70T8O74vE3GBxRpG
akGNCY1NA3pkRc/qJ1FI+TEsP3VDQ/I7JZg/zdBvJBIzHuOQ7A9aWo9urWwZDRiu
zF+At3NiFpsK1G7Jj1Q6khva4ToDtXkQj5Aps1HkJiST7cNZ42NPjRHe1GHBzg/+
gOyrsgr4R9vBm5fWAMBiioCLgCqMrQdrJrp3mMUOUTd2ekjo9ggkbyykL0C64iag
JIBw50FDHvHMgNBSZYsDv4mPJzM2W+aPn4JLJEgjlJufg1Iqm3rXxwTwSm9CI9Fd
N2+Ey8XkJshRLrMRJ4ayp0UwORLO4IB0h36vRnlYMmZPawuFmeI7tP4mM9tXjJeJ
cTw+27ryDAH9aSfVwzmq1LQAkGLOtUzR8ePfRv+Cy7ZNxYS+jMJVwh4+P00GylyU
4RLJjKH74Iv1vnwJTjrZf794AJHD3J65tny+aUM61HZnutg1x/AbSkE/6gm/XfNO
M1dW9Ls4stgZcbmBeO4UlJ/bR54R/ZoGKgMxbToxNUHg+yHIYpoXcbxDbTNsY7jm
FkFVQNLfGgAgjxxXYmiZfRIKmj/yUhSPMjLX2TWuSI33frH6OUANU+KJFtHD4SMp
KuY3BTH0vlhBs+T4S5VdixIiHr6OFGHNmTeqbfFKMw0sfU8xd7gFH54MGVnSIJ03
hkSf0fyxg9bbccG09JrNmlfjM+uQo3dKzD+HMmEaaQFwMVbkc+MpL6cIawCk6G9L
md+9czSaqn4laa7ZcNCUTq99TB7MxXozZuztmzDD9tGtIkGdL5sCTm5b48P0E4Ev
ahpqDX5+IITxstiNrRidCqEbosBG/sTdINllnbBDL7RUrg7SySqwgeLI5NZR/33q
mr+nXV6THqx8nNPZOCKESVff5CjEXIIQPH1DcbuJwdJ7A+/AuU20GA/zE2nj8zX0
4L0KKkoxbu27bxrO8SafLAJYfLMdxjyTAYSJwWOqKtxIM6HXWoCdxoTLvJ0rdF1w
KqsVQa3zA3FgejvwXrSAQ8qZW0l0dJoGPYzCVzeq1nShFpW02caMjdasqK8XvnQI
432g2RzbH0NaHZ/Z5wEA1s1iiUI5sm+1xr9bN3ECtUT8ffnBPqv3Tn9eNmIkZPHG
D1VcMrCsPBKNedmZV45q64FNWRoEH+f8JLZ4XXHT+alhJjhpiSH3I8pziPN2sOsV
Yd4G7HVKmgl8ICYdT1tJS8Rs8B+LaKQqbDm8yQoshmbzOYHUXp3iEls0m5t6I/QZ
yYBmyoVS1x6ybH/gb3G1HVzJtY9Uz58pSB2xofnGFsW/btDtjAGsSpxDfLbRmMLQ
R9+9bVGmSJIVKgFuPipicwBZgjO6bCyCK7iGh/ivU7uQQhoGwE5uh6ubA7h5HMJj
2kAvTFwrYdJNhzU4LFX0qQrlwPwpKYuFBO+n4QNk7z8cAvVnMYYRLwYemdr31j5k
47MlVKFHJlDB3XD1zYxBMA==
`protect END_PROTECTED
