`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bO5LR19vrRHadls8JWW9GOffA9KwaeagWwxESlco3HDM3cBAtJb8UkTioK6UtOGp
9fMOFfRZCHSq5fbFFwVQ0cw7NK3icEsyfewmuqlVx8Jpu7lnI1L4plfGbK3MOS90
qNbx07wUAxUsmlM5Rf58ErG+w19vMCAxF3sWe5jbYOIV+AJKhcFpL+ocaBHlTVIl
RZK8M8QM5mQsj6+PIqq8VCiQcblO/HJTIodECvs8DR/YZIefvhLlrPVoSV+OPGXi
hfeaJ9FSwPa3+qBDjAKs/FX/7f/RRC5Vp6yGu3QurFsEnjA/eBv55A3PwoCygZBU
8iWL4cWicva5Bcw2WvpWnVFyXKWloxyVKp0oQAlFXl9u1XnhWR8+rkE26ZX4Rszw
j355R7DCevRBxNTKMob3PsCSp5eOgIbzS4lpn7qd0QyNlSbhCprixkueL4vylqM7
hhuWpm0RYg84iD4kho/WgSz1pGB3/NQ3ssFefnTbkHtTslvPwcOZVttF4LPIrGF0
JjOhJ0XqJYrFMIgzeESt+k5xCv8zWPJMEX/J7UYbBx20Ne2G1sQmfllRRgf0C4Q0
Zi1LLtNL05adNzkleFoaGqSU13bP12ERmfWZid3V5dMIBxKWUR2hXF2nsoFXCEUT
GCnUHtGOD3cemihS7gbueAKyWB+t0xNolBLlsedohu/Q/gtrIKMGIGFwKjzZc59O
85Qr50FOhqbGKIYTzmbaFWYsjtnwQAgWuEoeG+Ch+zOhCw1f6hKxyIjGFhuZk+/6
WJa5ns2RxUdfcbc/VRTdNJ0EkQEZEKy029gFhDrggV/c5Qc1cyiQVU1pntnVxRFh
FXQ/FE3ErI1xby5QmVewPEPJ98heFhXEkJtWzSK249PzPIGp1N/3V2aApgWRsJ6J
FvKqdyIrc+de7diDKTvZ/rLrWlLS+sKIADvJtcV0KjRNsl9q1Qj/qEBA439HGfsr
/Rq2YK1fmg+WkPePh1kxpblbVvIEkJVpRIJ3TJUvhsnnv/T2mgD3BehGeQ4OEbVj
PxfrlS3bK/CZ8ZVkl1m6COeIbkFMH557a5Y5KytX+WbSQHw14Wvnb3uIwSVm5//d
leVWDhTKJCLziPbQSqjmnml01OXF1YBIkz5M/N1SXo/YX1j34g0k2B/tA8QtJ61F
NU2NyLwFh4Ls/PfgZV/ouISr1RJUx7k6T4m4a+oDk2H65fjOtvNGzQX1Kj/QqG3Z
1xDr1b9YdA9sLyfXYd7Pz3A4q4eX32aQqzcLHW9bcgCAwy3zyaBxgpBEz1q5LrhE
TNYA69KP5yiSYznoXuEJ9taaOGlZtCxNrN6J5H+Mb8LrJp1Vdz4wCkk1PQLRttyv
zO3KoI4h3Wom2W9VcqWtVjXUoj84eQA/vj8qA33qUcHcg9rgVsirzzxOFLe2jqAy
g0k0hTf99u+YfUxq6FIM3dMQx2tYkhK2eGyCoPywRwYpOthYyHoMojuBHSfT536O
vfPVLOZ+VuDnf79/DIEuN+ncDA/lHG8N5vxJDQS9Shv+RDugDtZPct8Ax9CEP27N
796I7ayrjEr+d6k1W8/0aUPu2eCia0r4ELbLN3ae5jnerrVdJHqx+hWop2gK2Hu4
07QpefhgXg8XpK6s0X3+qlo0pWDhOqS4A+XvKW4by2wfcnD3+O67fXQhpuQnM0Kg
qvM8UflapDUa5/pbE5Rk4SCDAR2+SAx6pqfUyD3NpwQ=
`protect END_PROTECTED
