`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eubloaoR5/rQPeO5jCFXEPB8E23TUj9HLfcXFcKihqjzF+GPXrhWe8PKre/sAikl
pco432kSBE7rm4x52Fx2mJE2t01cz4zuOLimn5y6Gtgwr1gXx6GyYAUHPncPPw/t
s8/CyJ14Z9nh3wbHeQaZ2ykMM0lclLJ0G7m/nYM9kevKXns2/bnpvMUqpheBtFG4
0ItZGGucM1xKPdXfXCTB4U1nq5+AQgpEDu2idrwZ0JlFYhXXMwcBwhtm1LkeaRHr
/waMnZJxFyhu0hWGAAu0+F0lu1McBaYmF/OOm6naD0dRTOdyH/1zHqPGSvbIl+Kc
a88C3iqItv8WIPW5YbrlNYWqhFVhbeX4LJvOU7grl+5L8cl7KrZxH1J/6wjRg9pO
nKBu1OrPe6qQ1zzQywq6Zlagaqfgg67lFoLZHIErpm7qXlz/Y6IzG3CadmCNiX8z
i6od7Tkp4bAV/BojkZ7H5Ftl6ytm0Zh1Sf8hr6LIRmhmQWmKrtz4P4wmTt626fwi
mH8ezpnpUQunjJEJN4rzBL/byq09zIe8VbqDoAqOmWMXzVwUgKErA456FuRC4jya
GNpNghl1kP3/0f9NylRbXLSyvgDITDRFZcEP3SkTqMBG4QijrVxhkI7I4PtgOU8U
5bxZ1aWqbr7/IfZwSZbPwXXXdF3lN4HSh8Q8i33gAYmWmpnbjxVy2l9D5ovBPOUi
K+FYmdQHCm4KxWTSBkhBEvn2d1bh7SHdvczyjoImeUo6eGIbZWb5jGDxziDWbYJH
JV2uD9UO2uFwK8BcBWCgBcJfIZWOaOiD5QHJNWSL8xcfpzXM0ECkmfUrn2WY1C0E
G3TbTkPCrHS9GgbpuZyAIL63iZOJMJAEdsM47hHrDav9o1aR225qoJ6kzSntuNih
PKQP6wUvqed7cjFsWPpB9UWWONs9XDEXs+fe3WbNiBq78UDqTneiZWZ8Uc665nnw
h36zojvLfPxdjq2C/ADVEfBTVsRZ7xNki/508BMCHEbOAwdRjw8ishKmiOLptUjo
oydH9eHw1W/BvRfZuLJbE3a2rVfAveTwM1mIijCN/+p5fhXJVfw+iKVIXUGUSovv
fMFFkJKZ0Jfs9ZkECFVc9Zg7dxbeknZf3prBW1H9BlC2H3ZCZRiYIs/rzvKuoi37
lAsftu+i2KI/4BGHeuOkiXu+MhREtd9pqjIgcxnkYIf5O68ql509b+9g04VvSZtH
y1ZtLU8fzWFxgs8j8k2iMgkUmK73ebRjmltPngDh56TDFt0Zb4NyfZItxtHDAJId
jp+MnihDLPnvlTLwl18KYVTwA3Jz9h7IqNrikWMrM1F9CyykQGVz0P/63/Hlr5y9
toW8xzwvw0wsZBHDEAGOjDl+XpYgf8fHFR3vl5828IUvmUC57yS+NOL0szjgg9es
1Nrsj9tjCUupgsHMauUZaSQfhexYuTXwmBrGLIyAtw/ZfOGAaYAWu2pfPEAxecUF
IfN7uJ9tTqRqakzERdNwAUH/kQbEbLo+6oeaFuCkP8tx+M/3buQiBRxmXblnrinU
A0KoZto6fBw6sTwMOXkZNwg8aUnRF1wur/Ag1inmDmo/eDd+dHDsyXrF2Cvte8Oo
GQsor3yZ8HaFi2DzDl973EiOIka28d0wu7uYV4tIpWMtufs5tIhaYR40mN0ArnCQ
lKosvOWeeGxenZta1jn8DJtqQFJbIqXa80dB7RxKNf3PcLqo7/hYWCk4Upq5MPnN
IDOBj7rOGoKvaE3s5Nkzjswli321d1by+nRtAGDnCWLSOl1I9jYPMZXPOuC/QhTg
QZ6WQrpu9lGrc9ecoRiuBjfkYiwSmIZt/sjSWElk01YQULdYglUsaNFbFTBfWQC8
XeN0jfUu/3/UKMDkyGXo2WLQenOoez6MLaJWneWMM0bX32arJ31nVCWhXrALRfTl
+vWb1zMLKYMkxLif4/yEYwODjnKy4TSPEST61Spy5BTEUT/lIQ27+Gh3hvcqZuAU
NK6YZ5BzfDPzbxrgAJJ5TbMEBn4voNIUuYeWiSsiaKJy//wFHGM4OQUvYiJZ6DSO
srrFyil6+T/7qt25TiwCgztX+OLoCFdXfYUOynO09h2TFNGLMVbbCqWY0vOIOBHk
47qH+B6uXNjtA7gwd9UcoD25AxHIddQZBCPAZTaNRPavwu331bZEXtfyvnwxKe04
4a0X6L7xatT1jGMw3BBQqgkqULcocoQ32W82tFhgXviVKqvGx3Ln4Z7+LMyRHNcm
CuHLdaPE7dfmvKw6O/7wQxjq59Y/VWkQXt7/y1YgUGhj6BbszW9/29BDdGOJfiO4
iqQl5kQ221ujynb6CO65osX8SyaCSHneBqGUpY2sWAti61wcwFBLeHiy8Y9e7zq3
rs+WUB/1f+i+zEJxFCnCubFX+NKJw7EkZeazNOIdYO72z2k4YoYOICxFtGGHz3Vz
hiVNQfNAkZLxEhvrgYUhP7+Um+wVLTPkh5izKf9y0U2Ek01ruSDunyGIVaDsRypn
nxsEhEwKPUSqVy4NWgsno3Od6HkEga5f/G6mXbngvIWIDj6950R3PlHBMQlPDSck
DYpwc7EVc33HqDqTtu6JnPm9Obcr7EyA+G1hWhr5JIq5QIIAq7g45JnuKQ5oG6xl
4RC/xepLQFAjJrppoRFstrfcZKRVE8LydnMrWu4Gj7O6MNvMlTDy3iX4QWYziuQg
zEHLrWGVfuKW2PGQuTJ6bM8IomSa0d7DwvxGIiLCX3J1nldinyjDRkI9XM4zdzvT
jChhB3W0zLb+KQ6vRFc+JY4vH2S0YzMx6CtGp5W8K3/VeTtnqtgRmi1BjD0105O2
biHpGxzleYLXqHxbpHlUZH4KgEnojA940S0NUoFnZ2r0l7Yj0cVCgruSn5sgneka
O/m5uxQ2Mb8Besf/wEX9vrA/ikK0XKMZTWUEN7SSt6OknstX9egdxzrrw6iZIwnt
xiI1g+44GKg5i0tGoBTC5kLrBRxHu2JISi0Jyv735ii8hMY9I3C2CEiItT3xoHWM
zLHz97+wfmqr3E+1KjkUAtDqlZYrUqe6m5R3fBfFAonUYNiyB9nGm8gYQPZUF3jD
tmP3u+hD1oIpPNG+BT4qJ8x3rx5fIFg2MVfN7x09B+T9DSnpQx8eCbFfaGYMZrti
ngtxUWx09OGSeL8vbEtujAZS4Yn8fR2UFuK2otgkmC2Jf5n0xj4FrmMGcBfrc+7K
t3wNck7L13nxv1JW1O7IixuCpqhTdgpF+5U8hYOkt6TFMUQzhLYKc+C+vWLBUsdt
Fcrc7Cc8oCYZt+K9RGHxX1LzEBItzsFyym+cXEf4tKc1ZJz1Z7Di5/k2JMItT36e
plv2K/zg0Hf8CfbrfeKi6lSJzEU7e0+jpTHe4dVLOs8r91ktj+EtghMX5GqwvbJr
nTjnZAVGf9vXyQ8SBt2jywRM8zYZwqlHEpUT0+ixmmXvKyMjecx4YdJqcq343JN7
3nbQbQKWmuzY97//t/bCeDElBpkHCZId17mP9RlF39HGc4gk1H20fTox4+4K+2tP
IqS4j4NxaT03s+MEFvOBw0yp0W3d8Kp/9cNddvXUcPLcisQX4lE6NjOnx6bGC0yH
klbvBsNnzYPWXjjyA2ALUHhVzWzNF4aQcLTSVdIDot6S4v/xtTQ1QPWqsqKYTBxc
RWSypnHMR9Vk2Cdzi4gCC12WeB5eB5GMtki1QcUesbiJL2c3Pyfeul6YBK1V4hs3
AwiFL8A99F+43H43Ipk1B9bn8c+50pzAvYLXtz0sKgWsbFYpwBgCzJWypmuzxbMN
sYkip39+T4YOB4Rm09TglWZlLxy4QktOwA+t2HOEzAanPVkNwIWBFhu37IAc5uWn
Ws0JMoGisGkYtczFdaVqXIz2cAmzRpwcXI4rxXxvv/xY9mQ/rXMhOEJKRhdinPqx
fyF1HEz2k39EiTozA4OLsAA8HZvvY2rVJChsu3QCvvtAHapWo2GzQyqTUWhU5bs8
eQa21wKwv150on/Q8SU3pbqy7gyuBtSItxTLpNMf8i7ZVgEfYf6u6T7bIMyyyQ76
jpJ56cm6Xq5C/m3bHtpVrQOOQJ3J7uvlUgO3Lec15gyigRZ7pcOA8qBnxU1/RIHg
q+k3M7U3/8nspPdM6BYNbg4myeJN7nNpA1Hj35XYZfL+luKQO/kOQZTYz6UzjhxM
+Cah3fccR4x+4rytXM6VKbizS9hQp/FGj/9rLqGuKmWnejJWPTQam4dpwfjnjSVJ
tKPQCuBZZzCoZ39RRPVy9hLhFsY9oQrjw2N6EK4jK2X1PnNsur+U02BwoDdLSa5H
+dlGQHnV1aXrxH6TgGBnx5xjTjRsS8LTcsbgalO1CbQyf1mziibcuhrhTF0EJU5D
1X3xg7d8QTQjzANBfng8yyOmvv75k7/XaZxgGMyhaC3NjgdLiKF+Ee5kbFO9Gk94
z36Ax8oyNHlVb9qcpmc5R7verAlRA69NMEaKA4skFqeZ4eWDulrBISXmLZBo5MsZ
tbinRGKXA1UOpO2+g1C3cW391siLZ28z+HVrUV1/2mjIRYvJP4T7to24ndge9Idb
OvAjG9pk5b31E4B60vhfKjOX1SEqxPozNug7YjMcQYe6mB5TRlr/gJfs6VRLDXJg
+zMuotCNVwJ8Ndg+EHaAC3ylv3rKm7gsqpqGyDrnFKxm8xYwvJas6DDDXFU/lT8O
ZRfGqLw6V31BA+V/KHA5qSo2RSdpP8YcEHsxyxDajFLN20sV7uAvpUS60Qkn1TDs
A2hZhRucTcBg1sZa3oXXG4c5aQfDBvz2PA/4Rv7eP6G7l3+hagmpT312kYAlhPIp
xxn/FmKyqAFy3tiPpcl9o1QdzDqw6KK7eZfXgBLk7G89bNav0VH0WJtympEu4hRK
BYVBSBTA7M4zbCE2++osM8s1EKHmcbz9lAaRTKPPMrcBk0DYY0WornRH3ImVMhix
o9lV3/bNW4IL/CcCmmoOrsZYnOI8YzuWNqaE6TgUE5IiucBYhY8YdtTRGuSEx0Hi
pV3N+hZvwrEVkLU9xN4US5B8+avcRFKPrrjLgzAFNIxm8oh7Uok2ALflw0LJNlNl
4L7gtN+UlMYUx2h/F5X/C9wPOb7QAeklcSY6yk8nhmgbIr57FlyGTOzuH1XbcIVa
x1J2tcholRk+wd+DNBO+v+cyrxXPjH1JymR18SKRlRf83lcOx/8vaHICwrg5XYKi
g20uaNlGQKiPJh0UhMaiwObfTsUC0CCSnvlo81bYTHIMqdkdmMUqjJNQULCSKnMF
1r+ryyNUk+8TjzMhhn3vA+sO80Onx5mrBvYCETa+9Viw3DakiHoB0EYeiTgHAqTo
ebBNEPzFNKn2ALOg9ETRSesWnHwa8g866rPuZpH2gC02yEvFhPrjGvbaJiS+HFoM
fvYY1AeXjzWspEeXaZ9rqJxVBcJKfIln/FF8spexW4+C/Tez8OrJFpFrrtDZFBlt
cLzFu/Q1g9CdYNepejo8ju2ObSq7MDHBRUrPjyF8huwgIdB91D/R0tAqSa6JqqzZ
33eKVvZ5qRzLFSudAbTGSFxUL+kEfiZVy0a/FsK2MS24sCyGBOuHdQQUsy1HUUkV
rjuDyHSLRPad/yvOn3ld/QHafL3ibiM+WhnkVDltF/5Ae5WMgkgjyH79wrLwgok8
6fohiT8pY+24toLntNppHrtophGJyxldRXIkALw1kVTEpjjDbD4M7Mlz+8k9TSpp
mRi6vvVSaEm3x7AQZq0uMtD5IFZgg3o9Kew4SzuaCigURVQQsWsQnStcsULArS8G
Rmz9TvrhKisFZBQZpnUnwvCF69XT4Hv+rMNuWO7R8CB/HGR5oCHidtmUjS4N9+7Y
s1txpO2cH8YLYqfoLPNO3lFWncZ3b5+07zsTUfNnJdiO+4or21X0FBtb1zMwaeni
mO5QK++E1wOm5s5mRafK2affTn+WASupPUPny5KifRw0JpCree/guz6t+Bb1Hq7J
ovXk772sqVolZDTYjOwNQR5zkPk+dYqS2f1B9VlPHHrLPc+omkqV2bIXQjAi+pRA
MRg4AaWx63WzDAigqUAOqX7+eWPepMk1SRlLE1xpxBIax5nUl5Dp2MZTaqVs9nT9
o1L9VaiDe34DpMeUCJMkL8wM1Hxt8d7b3hPBWof+s0yXOKJlpmnxBeA/We/M7/aN
KtLCIuIQHSQm5xIDsyczTXR79vjjXG6cPfDzIa9ruNhbaWTT1tAlIg6c5gsTKokG
bpYrk3ZXS4h0RJD+QLWSIdYOgv6/qMZcyu0RatfpQDsoq4ukgFqADpihqkaFNFFi
LP2Ye3wGQuC6XAZKsy0Qq0A44t0VDlr3AF4jxRjHgeXtapQXVS4Lac8Bre5v60sy
Bnc24XhQvJbIH+A+UaVEIPDXai/bbVL9CR2qMdnDnFqVSnFBEVWN0vtzMLnMHgDs
lFYDoUML2hsKUKrpiLpaloqvlZICK83Yd/uOIuJ+roOHmrtZE1hSUTA3e6fQt1Na
N4fmfngop8hjSJQEIHPvR1xwK7qtZqIl/8uY7rUx6KHpOZd3iET0ZfFu53z1qZ4L
DSjfvW9fzfcNBwpn7Jj/gEl/d07CM5clQTW3nYFAtNkEcebbYMcZJn+vqUTWek/6
xUb6VTMSmbXgbjnLJG4+zlBvxUMBAHaJbaZtsqPP4h9kIAXwTvrJcXZ83tUWJrtx
dDHAX9EuAKVhKO54Q3zQvHG0WtBBshddiIFHkoCdVI21tDds5aWS9dKsT956JqWu
PWpYO5CMpI5xXlzolxRAKywp3euNMrzdr8AbtCXls/597TC9ULtwT8/MUUe8N/TG
sULUZOpZWVo/929B9wF0hzHE24fFhzoOV1QGwfy0RFtpeBXG+wZtADHuboobCtiw
cb67kHHMoQO/zfqVMH2FOjxNEiDWeiDQ6mqhCExdh54kWlW6pYUeqOx87umYl/B8
4sQUdKYHfOFDAz9LkGOkwSc1rP2hPY8alAaY+lRL9hT5JHPWy/9fLOjoKv+4CK4p
+6RGfkqMCDLdCLBoICs5/9ajpBBFguEcpsYxHViF+lLT4DSHxQ/ZPGtRfYv4c5b4
KOL/XliGM3Y4vJxhuXOA/OS88W1SMH7eRVkxMc4S+l6Y91IkE/6vzqvdF5Ee2pyz
FElgrg2GOyjUjz+EGMWs9lsuFTwia60E9DmZULMAMl9puYGhS73zr0XhcgvNicbB
6N1yN4VI0/pyWEFFBmJVvhL0fB5PknbhNPst2EloL/dITnIfJauu5iI8gq1oi1jc
qXK3VNAHswE57dScIlGxb6jLWMTeRZu8aT+0ucLo++kkBW+cJB4XyLYvAPaDZF+J
hPzxBEy8BKy4sS/4DlguOSoC4HFJJgeBjsWBhV9KsFI3+PLrk4pW73yET+HjaRXe
eikzbpZDic2bhVssjLMVGqFqo5DjufHjXtsqYdUJYfMFjGzePqeTMDo9QAu1TNCz
6JnjQYj08nrGzUnSp6KvDqrR/pojnq/cbTZsZNQtSwD0xJ5hyCcNV87xtY2K1kFD
YrglxlNU6Hd3xueIz3nh7xthbZHxWfBWmNYw6vYfgkZhskfoUrzyW3C/TizW7chd
iVoioJc0GIbZK//EVhV2qOsrDacldxxReh/0/wXWRSuDviRgMqiAATm5soWZGM/s
xBer43U+8+23Z7gc+jGO1C1yccYuHwf3FWgw/SewHWjzzMpb5wkwrDf6AqcRtr7H
Z8gLB57FzukFpk1dJ84n3vQwzL5lq5e1O66+y3okRIZikr9KuTWAsUn4nZiGh6aE
UyHeLs5clpTrQn+xweOaAWMLB3q0oRyxl7F/LgcsRrYn3yI1t8T03SkoP/l9nUmG
V3lHPTCXFKIpGrxI4CagBnpQr03wDV/SF4xiHdVFnpgkdYf0/wyEyTFfQN6jLKjz
D0qeMa0l2EN/wz3huVAshMBnbWKdx9GdgQEVJJJHeTLK3rq40wHnSmXoIpCX7uIy
VaZHDNER8r8qt2ruEy+pA2a2Q1aIVGuepsy3YSUNlWO+LNrz6vBEOKJLek2uxHKT
RQIszxXMbP92V/1VR4psQJzPN1FkgA2zyfXoZGUUvyuR82IwULfofra14gsrVpRI
FDAi1eSgBfcNaPRiGWNGUEBll8MRNYY7KM0/kVFt83Ju9grFxyMczBsHEzkqqa07
tGaBAzsXnO1thSJcQLetT/o/AkaMKcI9Is944rKqbH56P1uXPDoXGxjh1ZvF6sHg
EY4lW/iQ7yLisbJ01PEdvGWL4am3Oue03UzT7SPnht8PhY+rF3LStgtfx/+oVVOy
cTWxoRFf+h8TIGe/Z3HhewC+c8skxYev4eBQ+zQBSEgq56J8wIFTF2bZbhMbVrtG
7ei7gJyONPI5BePZ2+DDxYZhJFLxidmBL2q38tz+9ja3lgmIJ9MDEIRojz9OxfYB
r+VTrzZ55u52pssFl9Rr2CpZFhM1lcxv5zX3a+nBO6Y6siLL4omN8OYs3ZlesQdd
+Ikk5p37YG9TvcABUm1Q3WsfRKLECDjRYCUklpzP9u73yM/NXNsWiQy3WBb3eEEm
+5c2kb8FsJuNkq2zkknJGwspDOOXPjcsCnhfxHPCUZgfIk3pqEn+IuzfoJQI1BE5
eOLp5GKvO2Wi1OLaaoegtOyU+/kMAYpNjxm30GCdipsE4MgUBa0nk76qRPsYEqo2
1IqFer6dNEuHV/GtoM1aBt+zfNbtz8PJ8PrFDb2EPon5FOPcD50qNZTV/GetZBkC
VuK15CRAQ2Pfs2SNr3xjt5X4fwEhlE5wxwwAog2pw2LXW7g9R01EftPa8Eyp3UmH
ZxFFCS8WQueu+HNz0/1IWVOPJk2WfGXeAdtePYZfjDQvd200Do4KPmGC+H3vW99B
Nnikpft3ABIndjWSpvs3K72wpiFvXapmmy/Rrsv5lDe1f0S1vIyPHZdJyh2WXml9
mpFck7Eb770M8daOFWTJ+f+nn8l2ckW5Q7eNTXoUWr7dZ2eYicOrx6lEQuaUFJ3u
+p6X5rItSCA4e73hfMUKlyIqtSwpSF7G39gzKlkj9JfMLuWJ1ha39cNFjCWRYeN/
UVVjTonKSAYkFw5tI79Ic7dhj6WQULq00Sd+ITf6ARhHEXBMJP5enQqyAOiVodnK
EticU/oi9lC6qAE09OjfLJJuT3Ch2SkbjxXj2occ1c5K4lHNFT1qlli57rY5YV7b
cix+k/sb4KQG+qPZO6qSAUF2JZQqNwDTmviy8yWR8wLtosgaJ9DS5DIDDkl8veJW
DzkIM/5uqGAMeXNubp3E4er8yFAoABFceGJ3XLVko2+dkPzr+RNCL0ORQzypC+hh
rK0GNIBmEKtYDlgrjs3CEzGfPntJdlonFEVmhHLTbnmgFI1aUuxRAm5RtRxIp7Lg
Rn8mIS8rXS90Qv0/SGrxQU9oNOf4v+vUap0KrxBFhRiYXm41tVN/QzxVWBuVLjgE
CKv8Yyd+ZpuvcqZOLah3jwX7NlHzRVa+NiOIpm3P1UG/I31Dt2vNBbXD6QofBg8v
KyYxnzdeVZAng9Qjo0aB4t33XoKwdyhVgxEGtIPJyOMps3Siaa6jMWgoaD47jC/Y
3q8riC+Ood7n3vl/VEircAZugwfEdSPkVejgfR6YO34YFUJbPTzmg3VibhGDoAnb
fs7fz17oB+Dl5X3EBElazzLyUt0WBh6BZDC4VOtxEux2hFoTazZGTC2CyKLx8LYh
KG8ql64DeP1K2z9XewOccEwcaGa6qJTMsfy186J72BV3rgBo/rciEsqKvM1/Ojud
p74CQjIxpedDdgxIURzOiSbAevecXmb7ipw8nF7XsHuZkyfxzA7V7Mgocjqw1iEZ
N1+JJ+cn536skmwR2AIFHYXBfOxQ5s+LNsNwkHL5C1jH+/lATkOnImNmZwN5b951
Ry7zEKET32TwMrIfSXcZURiEAz85Z3Ttd+LC3e0a/5qstiQDjunBNhkaEpjLeDby
Z7sCayzc4CyCRBPmxZY/wSq6Cj6wEM2T5lXts8baCLt0Qew2xIMQvudJBFiAQoAM
j0UHBT/nCanKGkMy936xTERSeqqtbepDgyrfw4dy1J+DzTIEx+FMN6wLpHDH7BOK
szbGIFOYp1b0mBahvRR62oH469lIzbCoVLoJrDwQppCUOJ//E8lDcm4aYEvjvOiE
2wNCrjGQzTibcNiVhKAYWG6uMuQ0FhX7qPrlXbLlrdRR8xpA+tW/GRCQJokipIiZ
QGdeieMDvC3ePSMcqZEF4yuW5ZwPx/8rw0or10zNDyCUSXdWsgr5dsYPMvNoQr+w
nKNSerCboUUxZ9RUA5Tu0hCbxRj4Zz1/vXMXruWvElc=
`protect END_PROTECTED
