`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E9hBrTwzgXwY0i+K2Ez9rLE0FLO5uq1cRLTlfNlpvpzhFAo4JqO8ZgS8mc1suNu6
+5OyQEBloZTbOlZFrga+V9e++BcExqfCguwnSZvk0T3tPi/694h/rJKGU7neiOhD
LNhn88M+mXaGiC0t7beN2qLFyiqOCneJL6coxI2YLt7v9RL4Sxdrr92OMCneOZ0G
+/MGBVIFs+4WD6/tsNnlRhBUG8HG6jhZVdsPFEWa7ANkCRerVTdfC9qBvHjEPE7D
R/k7jzBrMSp/FYCr0zJsYg==
`protect END_PROTECTED
