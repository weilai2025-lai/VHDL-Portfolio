`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g19F7BZQrqQ7iHO2y/ndtg87iJDJXOs209sJdZGlA0taJ7clmBERPMX3oZQk1oD9
UAyyUylBbyIxeWsLFxGye+Q1LkLgMmfWHUx09XR/Mve8ODIG8EW/5xHUBN34l20z
Sn66Wg7ui0gReJJGM8gGz6UZFRpXFc6MzCdgQYI5cUFjWnc6ZpiKIzvOxtCBo0ey
W/gtZW0eGBxvrHZSri4N1q7YIEgONt/2FojcU6wMhXxd016AQZbY/EiSmWQuONt2
iKwS+K6/egKD8bO1XKon73W3FivrvhoRxhTWJJhk35PhW/4ZD/6yECAgd4WRyzGO
1065iYVjQTEfGBtGBNh2wewIkFczkhGjlRI11wIOmehkJLeznZR9SXOFMDRG3enE
2TSB+YRyLmxuuxnNCo1evL1rW3X8GpjTfooMJQFkw065JnDcO/W/D/uBa/F4i9k+
UCUlVz4GW5UN6/SdfPmJNdwzYkZHF8KUbKoAvAoq9cogkyX2R10G532uOIRhqWhJ
h4m1UV6YIsk7nB5ZdDkDDw48snc9oqDGrGyBFdfUBT1UnaKXo+gGsfwLkTb3oi8d
IuYrmbHm25nvdNfZIAuHFUVqWUUbi7AtNVfsTUsmNALEIYvnnhFOBnCFxqIvGG50
xTetTtQiNRDP7RLH7b6n0cPL+/MjGJExb3A2rUVHtEIe8WEby9xN8IhNe4/vHdf3
3hLG1ND1cjnaJRZF0Xc0lgAdAZOeM4GkyHa9H1Qd5K/yuiqMnwQeVxXxtPBRWqB9
N7Q8x6XAPamKs4UtzSbVSVpfiElLIGWzEAOcPpHzXjO9Xf5qegGV/q0Qwbko1y6d
`protect END_PROTECTED
