`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGOqFuG7xors6rnDYeSBvHCBk5SG6R7ST5kIVVr2J7eVkSXNCOqT8phR+JX/pJuG
Y0+tvIUK70IDYZ8ORRjlMntZHY5mZjO3XPyod9ufe+W9KEu7rrHi4V47wQYtEcfG
8V7k2OtgCYi07efrrvAQQ6fXLc9nCx35MxfGTNxXNDm1y36zxD/aV0qBrJEjcCV1
CSMee13gIjin3UGJ2DYdJWTCeZYED9P0j7CEgJWBlW09oTUU1ItM0Mz4rl0P4tXK
LSaFCcLhRfbB81hWmgxhHdbL/cwReMfqhmGk3bZDjxu2id2tKj1FgF4gg4Am3eJx
BrYgIPf1iip5dULerY/favgH8sLXxJPWLequbTaOviJzwqf45sQ6OA0KjgFJz+XX
TOcRsx+a/G2Wmswn+J79h6AxzHoS6BgRomTyz/T2U5aQa2MxKb/X5Y6Mi5B3L9qc
xg56DqLBUevFhCXa3Noh5EjsKv0pviE3NUVfDhUVVZ4y3g0Pk66AjmgPB4ZtYDMg
+5UnujFoZEYE8sSOqI6qYRga4RIyP3kHY59dR6MErQHbD/Kuaj6iCk29deQdBSO6
EUD+dRW2jFFUUi1hSahv1UfjlsPmuOa3QTcZ0QXHTsS7rnE+OsdWorgZHby1RFtC
AX9dfY7CD7EuuA9iAkmq6ZNBszEGOIntBRSY7pWiY4yNM5nrLjn1IoOTYokXPwGN
YsnueW7yjBIAiXPV6ahAhQIAhspwYbmPOrkz1aDhOI5GME2k10J4VeM9oZuQ1HwO
hmM6ff1sAS6XsuPMywBCltQ6NPj5af4aVe95FDCaQhTUQvjX71Gwf7gToTlWY/F8
Y2Be6JyG1CAyMYB9556H/1Z/4HyQ7kMXURLRH7K+zAbYLU1gOiGNEKI8eZ1gALzA
bpQ0RwZRuHV4AHvIXey/K6x7wdMPGD7H6KuD+u0CbW/fqwj9EIdQhyOlNfGq3ZTH
x7/Uis2zSNcrgenFJPcRQKiiFid+SN8ITRllBc2LpS75YJLtjI0UQMySXLsYcYwu
45SafdaMAtAygEKe9FX2NPIK/fjqOyjcOeXlKOyvnCNQxiCNlGqQ0PO0FlFPd5mj
r8OxMtU9nRW2e2pTP+ssra+dWQBYlEX77vMquCcGKUXygm4UBzt0qe2+whIt9gvT
po+sOAA5oCrlM1jjdFtt3v+s3+lg0V88pbHcJ7t7ltFhHpeU1Ig/3WEuuuVtxZbt
4S7Zhcm8r00mlWBlOBhjHX7fZq8KtqHcBUx7jXyI8I84RG9WsBAwi70tWgT6H8+U
v4ImdlMuF2E48Mtnt94c9kyLvwuCLrpOT8DifJzRIkjgIhXXMgN4tM8LT8UE+qOf
hSyOpP6ckNRjoNNJNa85gSFRciYbe2+1gAXYCKHMqa8wXfAAPjA1o4XwreZShQiX
G6P5Y5lusC4bZKgxxVgSivwWbzb1dXV8iRyWWDMuak8zLUiIKAVNppc4mjTOt0lF
afvOwMOmAlwrHz9DNycXmUVGfvEMz/m7NVaXK1PheBCRVfl+Eqj/Gj+EGV3v7eGy
hn4radaV1cfRdb02zSp927YKrlEdTZAIpQQWxqPiPBW3a9f+8ahPF3mUyUNIv4+s
J3lvnWGGzoMvZvkfuB92p6OfxjY19Q1oX2QNYiUk3xXKz5hYv28x6xZjeSMSJPT0
1xYofU89GVi0y/EqHc96EIJVl4wyR1qDpT5qoCYUJDkLoNyjQWgk9aNVH8Vpqvpy
HiXbSy08ALc9qzTWnnrlZKcJjvgVNz3/nDp764GKpDLYegLhHwDsSTtpySR5Y8iO
g6n3YmrjsZy4QsG+ZEwxBfEaiFaIzGIu3eJQBS+TIUtqKTVlgIwKWv6FRHS0ICJ/
XGxwxg3dRv5SFkihptug1klINYZghNsRykZ5SSKy4cUhRYPZXgg0brn81k0+ifQe
/+VBKfQMN886HYR/q5qofyQ6PWdrd7w99dyYdfsUfxAXlxich2GiMcxHcVhLKQA7
h5FTj3CrbOapU0Kh6BSblM7muRwOxqAW74NM1efGN4+MKPVPj6CttWLTPxxHYjrn
cvOrgyMutL+engwBCHVcuO0ixbnl/VIknME5Vx1o9xghUTtUb3GrpkT2Rm+UrPBt
fUx763ouiXysdyEX0ewApapUNGPMI8TsTn5r71HMRu/7UM9WQvDdXBf1zv+Qw7vc
IOJ0CIC5M8UJb0BBn2a5qt0EX74WosJDDL/wQX/iAF2cW3Tlty/K/BJujC01Esuo
pjPi2qtvhUFv8xjIIyw/tE4BwXwmpyPbEWRhxhkaFfBOmAT0BuFLeEEdIx2BKtlo
XuTO97tjf3wk4fXXh/rdouDo40ZsK+RNTeQJ8RtiNJDJsPc9u8cSImvLOHNNB2XX
lTteEHZoGuKoc0kngdLzs6AO5SclOR7KUkP4bMn/Vy/oTMipZYSPyOa0HBodAAvM
SrcA5WejRJOHABWOQpEZDaVLtf9CqdjT0nSq+rFs4sObHTH/rtF9D8rXRhJ2Mtat
qRiJuZ/LVTMcAY00OVz29X5pzlQbpCvuVyZZfQ8xPGD7fEBp+NDBE87IjpOojBao
zf4RwkCvwV8GzdwjNY07cko7vL/uTxpNYYh8+DOBc8PKIGXRNMBjvAuKEv3iEpdj
8ZH1tYJGI5KkPrjUrswtP0EBD9Vr1TRAPKFEEU+RO2NxqTKDIU6pOCFX/MpmZ8fq
Jr79MVkqAbSeN+ZfNSHyd24PNT1tdapq0pH64obSQc34FuYoDfgwrESr1oUCJ/Xs
sPU+1jTnvkXNukWg/vPxbLqbvcxVhtvqrchZx23+yEus6Ty8YbD/ClrqYRH74yuB
+Ch53mz7B3NNl8iGD4vgQZfLXCYfKgxDxxO86J4GgncMXQKPn/VbuGKo07cyxPjM
B3qALc8XghHvPKDCAgTnLTZMwwL5ErKUMUKEfaitg0sNtphW6mMhI7o9pD7FLZIz
A9q5GJ90QYF0jKtPq4u8bwuj+r2NGxL7oP5vF5qkSw4upUXcyqZhpa6wcoe08ito
agVDdPVnJLDzgB3PrpADJ0lJ1Zz5yL2uE3UvxOmHjxJGsdajX0DnTzYMJRMsHP/Y
V3Swk5zyCIfzGQa6blXPuCMkE3Dsgrw1HKD5W4HExMsK42xBDqd8Y46nKqoLsVVh
vHZBfdCqL2zabByez5TFcU7HauFUu/VSbcg4RTedkzy+3jkYQWJSMeHoXazWD3C8
ehLZEvOq8H79f0qAWCj/if6CsNsZiU8NZ0WPYvazb+yDpPem3li84+P4PdWXmCL+
cwPEoV9nTCxgUlWBaRi++JqTgpR7nFgIhxph4AbPUXimgPQYJLLzJAAuJXM5ca/V
eZzSMNtrpYmM9/75WLTiGs2f0byBx5fCJXxqcJUcVWpg9YE14C81qR4Hse8vv/Et
Bch6x6zyu8AU3aIS/oMp0QenEw4q07PgmstuA6M+txq18HdHHcFoZkihJdwU1yOK
c4SO9nzpz92MVaLyo5kzToQg7zr2jmoKRUTvJIzwkiTL5RliZusJLCxl/+Ii9LJZ
MTH64w9GK/o8/rypht862Il5z4SPb717LIkznwW/Kb7xLVQnhhDSlcl9w81+UgQD
3+Xx9+MdxNFw7kKzgDYH7j92jpqg2tCqqf2tI9EkzxKl2+shLCPPwZC9gB1EJRni
VKhQb2pN6snmJvECkk8Mp6rxg5rbiRq5yyHZEtudub7NuXf5+sRknJiD8+PvKuam
Lqfge8wtRv1VItyEqpFtxJ3mdNrEgEWuLbaWp13C/uvMypJNGoELfbt8hBtsNGH1
oG5YGUDnr1+HGFmDb2xN55sc4GsGAElCnwX9zL1v6zve/AvMqt8l1XTDOAHKVN+5
q2a4PtdpVjzK/3q8EMOX/kxPgLTOHRvzgA1y4RibCZhupgCuKysJ494tYct5AirY
mUrRBGVCiq9sitkt1I+Cwfs0DtYBU0dkHqOPUUXQWu1j1lXgyWtBVcXa4MmhLT1F
b4DfKn5Db7Fz0s/jUA78Nrlh+EOCJrnlyaIEcZ9tBiUNRflGfeLbu3R1yhlhGT0A
6cFl+mJEYa05rxvwXHpgmRoG++VtOLdIvP0YSF42zOKxeBC8W2tJKEmrpoH3+kq9
6Lt3nq7F/uqq1z9OIXAiilbGR+rtYtj97sF7HUwApo/bm5dkZjv1knTE/59xVEON
q0+bJ2I62FIHkjgSeSaurXwpxOa17hv7POPEZHBrrmaBKt43Jxebo9nn5S1bTK9z
/Cl9hFZ0hDAJ3Y0Ypf0vBfwjU9ewMJvGZa2Ozh1S5ifXaMh1+EO8hRkwgjHEzP1a
KcFihBojzxvPoyGY4epQc2zwdDL1ueDCux1YSjzTgmaWfylXsLgLv7LJc+BKKWkL
HwOsMLaIIQhN66mOhbH5JofitKV7qk2r0goiktt2SwWS4VSSzAWsnQubrKs9DuyT
ujnoShZCuqchor+D4+7Vrp6reAdQVZg5QSIvl2KuGkZoSRzBqHXgOesbDnIn3Bfc
TGW7keA593wR/b3M1+ZttYwFsbCeUYXgg5kNt3UJzNHomYobcNnELilfiIGeZdLK
THmXB71ScMcll+YaG0hVZJIz3XZ17OHswLC7U889Capw+BUtFYCgZI06NuSLR8YD
O8s0ZoEn5Xu0r1O7COnxq/MXQR5GW03RyuXGWZWOeBa6wD7HNoahT0g4CeIrCCNd
+xYMB9L2xcjazzrOwc8x8tyqLMvVKw9OzEmoUCtsxfWS26+68ePmJBaa42tBMaM9
BpNJGXWdqmThHmRTJqhgvxfaNjzq08xfd8orvcVa8f/sA+5BmWALpxg2IEGk6Jb7
e9Yk3hy1l9bOI+ib069ReGdOKjk9Q5QiMYSA/kXXXq7BYzx1w5jIRO8nwY+dBxhj
xKEJEPgL4lCNKciRgF7kYrBBE1Lin3eml/QzdDr7Jdr+y6a9E0Sr4nhC28HXfuD8
UKbbjVP95PJg2ZE2QCV61GslL0MxfgsNu3iZBOC34Mx89ZZqazJVR3nkGeBmmLXy
nMtEdLUXNgbaLITd6qEE4tuSL+RdnacVFzlBFQqckZYUe+BK0F8akHykdr4GYFjx
6t98chPhg0ecWLVEDA9k8R0GaKqa8DT2iNRGDAI2KvlV8M0+NYQmN+qzpVTnXoBw
KOuz0fuh8nMUtfFwKvQP7I73Q1WMgiFnSmwfUOiiBoxovXK74nACvaYHngmRrM8P
Mmqms8JmjQUSCq01okyJbtkkbV6FbSyFjAlOTYB21W/FD2skfq0IEunDBbeFCKXV
Sx8IDOsx/Q+tqcZIaBQ3Y6zv8haQhKPGbSIG7guFteMzVzbAMlFOye6GpX0uVAhX
LA2B91+vMyws9D7HJ/UXwCcAkH96Act4P3iTw7Dz2xK6nBx+2amzpG8ctdsCUfCr
Of3wIv8DpO4kvutIpY7pGAr0QYVrugRZBdUqwKwYDfx/J/pLA5qdpV3rB2UamVTd
bqU7TAyVJIrJIz0mAQDlIBGfUXf8PnfH4OfTcEVAFA5hYWQY8yXwIWMXEevxhf4O
XURs8knr8lVs2byTnoUCaRVyOW4Fvmq10B2buOIP48KN+gzyVMcGJnjs97yz3Quj
qb1oUNx11sYfdm2YWcFscCsainsHENG3AvX+rUsXMfqmb3qncyT8pHWE2ykYLX/X
HX3D6rbsEiAuwV6soWEvcFA7LCuawr9uptbuDKV6kz+B0eCYreKUnTSM75umNN5v
dkvgek/HZDcfGxEQfFRkn5UxmOFCQdekeaQplRx4G8NOn8zVXfjfC0ibtqcWYuwE
HwtcOlX3xXmA2MBxhxxZIsx10FNL2ySQZYiXOLAeA8RStJnnJSeBMPlWyj622Of6
tL6gS0C5O7Zbm70XppCq6AwDP9v7OKwj+o9HK7DLz5WFmx1HAOLZnYVXGBIYaDYQ
B98u1MB7lRYNqklQnH+oVGGvwh+Ze0VWSDrM6wP8lms2HNZ74eHAoKQE/7y7o9zs
/wcpxHma9gOIgCHiBle0HHkHg/Q0/GzuRgnCyXlMFyauz+tB2l7I9rXW5vg6Ia+P
T1ou8bB2RBYcWhi8DDhF0AWKJRFQLwviOHiEP09Pj9t1dEbqLQA7eIsMVtdCwvSC
4GtA4VDHnO5tb/GowDeg0r5aM+dCPxUNYl3UW942x9RysS8XfmeUPzi4vYgTnzZ6
Zmls5LtPSDh8eeUAGgQb7h+O530gwkotIM+6l0nI8XmGw7QtBUE9JXUu2oHs8IaU
8VQbM3Rbh7egkhURdpFG57GsDD8XHdHmpXUaqCZsnYeTKMOHO+MNl0ZLfIdLBCnb
XcX6jMSBIUv61IuXc0n7YHIDRtrph8KqsQS6w0bFj+EqaLpNSaA4UFyIGweOzWgo
tSu+W3PtqypL9uQDwsfOQxVBmLETCqiC3WaSYKjQyX/dLb5rBBKZnT7tdw1+a+ZE
EovTuqKZ3LTqClvZr6JmjO3CHN33b3H0G8KjJgLy3xUAVH5dT2KNEGsl7yoj5yuy
AGCCreo4SDNJp5knQeyQHEbTjPSS0oav3ud4PikE6YYbsFbmFkGjRjpBpXAxag4L
h2J3nI+UeOU7w8hqpjpvEs5FR3l/LNwY4FrxQuCG6s+xPk8pUP4uKJm6UvGPKG5G
aaka3RZX6f5sjArtq1aY9FmNW5T0+lZ3KLRLVBufI9uFTtWWGq8E+8w0xovJJHXn
iUz/Jf/NfcSD1kctoOf6d7jCK6GDTZWYPm3ogxkTw3lnrTSv9Mh01OCQEUQQr1hP
kMRnwoFtf32VQMm9tz650v2qgq7zEpI0xcs6BHWJhC7NnsC25UMHNZhHXWwIkk8s
WcoA6d9KdMxlIBROkbWZscwxWT5wPpHDyUhyGJNnRNJhXbOt/BwY07yBj4rgLLug
aEM3PzqFduH46deQpKxHh4vNwqtpBU03U7B8Tzyi4M5zOQO6lTbfyBGRmTCUGAYU
zb+NxVhc/8G0FufykaitAMLoJJLc1hQDItR/MhBSeE7Z/kxKx3AxFozOIRkAsas0
PAR69X4kr9UISORnyApahiuUe9URFczy0W8lxANndfv9PC76rdOX5lu8JDU0J2ia
QlHtGgr9J2YfQEKIpMDzWpspI7U+ix2sO2fdZNptecyRVvW8pEC7cNBkN17SVWhM
mBwtjeJ5TpXop4PY6Eo2eSltq0WVZqp+FfWxvEhxKF+xB8CsvNI8EEHEtwllx/4m
GLKlCspN5y3H7PazYFGyk6PNZQTb/u1WKwut58yuwQp1yvGLQtMIDAk8tmIWEx1t
9OqdexPZNlm4u9qnckRvw1FrCkPaoH3sVaWx5RPMFn6O5/PBxqFcIzlVWgAn7fbv
54s1QyQTHSoBTrMY9ZBFOXiyZxktxXkZpfAlOrDFe+Aajkw4A59xueJFsZf1CBPY
5AtlTFevJYGw6OzLLIKl1zMBJ2bXjQ5miVUQcw9faRWCH1EoDy58482Gjay5+4h3
H37Ycmz3mROiBS+pBQ/npiC5hgM+a4Zr8bTB0lp7p+RKdQkv6H8rVQUgm9pOnT34
xhSka2JwzKl7Dr84LPP7Yzu4cPA1+xkjFbh+RyfIgST2OdXVhpTotey1syV6o6oF
uICetl0pW0+6MTZpxihTMfi39o/IL4GWkk/5r2XZN+YEuS9sLCDr4O18al4fus8g
N/X0Xt9BcgvoIhjKVvL67chW1UbnNL6iVNP4VhM/442bHQ14N7sp7cGPWLPUcaFE
O3NyaR978WoY8kmEfHUzp7iN4ixtzrqDCdmIq+/ifjMJagxQkOGf02nW1xQsis2i
i3otWKO8nF1PMaxAa7vXsuXwtn9uFX4EqpQG483ULtmHo5FTKvV/hmkJBL/OGGt/
OdTJcHMcKZ5z2FF4EIYnb9EfoiVIpTynkKHMWMpCaZrrUnQ3OamC6cRVqp9AcjgA
HlyNcFckAfvcAwOCDY5j8LnJSJUZUNSSm3AFgzn6tK6vZ2XWkzwvhJtUYecBg4Si
dwDOj7spaHCoRx9S/uqGDuhtolU3HfeyMmUVaL/gwI+pH2pjN9nmlOZLvSZXFICn
MH9tsjhLQFn5Y8uiRL/n7vx/VioWwBhbUQeUpl5+ujDEKYR7QgiGTr/MaklmmCLC
udVFsfwecO5U+lul4A2ck8WV+8HuhVpbE8wQP5xR9NjagrWlhdHpu6OprqKC+AGN
XcEqbP8sqn8hQqPZpvn568Y6f8s87ojaFUuJD537Ydm1uG5AWfjAJFdUr2iRr1SA
vzAPjts8aqoPbLvDthVhbqSoS+ZbhuIdsz40wnLk+BNdoaWHQuIizmkd92PzbCwW
lLuB8l75maTZO5ouQs6Re1l+jkOMfPn0yBwS+kOmhe4jlhDUWZsU/pgG3Cc1TLbu
zCdNbd0hUrJGHDVwYXgKAK4Zpg0pI1LcAmtrOzKGYUWZCn6NDW9D1qZXHvSp5vxW
JfJaTcppawM1J4eiMJHqv6zYB2f//3YdNipFIZeNAhqwnLGqH0q7MaKe8Q/a6RjE
QlXOQgI5SL+XX48THDX/hDBHadMZwKLp6ockmJvmzjUdV2uEhWYuyH9Ds6YvfD4w
+Gmva5k9Am0nAcbIkbcA6EV/Qx4LP6ywCQIrmucZMeN6yhIllJQDwwxkdNBGkEbr
iORfykKC1JeOkHABkvY+m1i+N4AzhNBE8kxnjdApbgnU6IsgecaH4tKSSuaigO2x
2VXZGa5CImKc5lHM6WoqK8yHSsKQ4n6Fuavf8x6tDxvSKmSHUhkoBkfkKcZCi34q
5cKEuswNS1ZTW6c2ngBlDCo2TehmTmYSRnTD7yyWA0bS8Ywz34yOQwQ+uHUACA3X
VoBHp5hfR1kdTfThoye4jA1BNIXFG7a+pReR3Rx2KBlxKfGqYI87tISYlMRpsPL5
Bpx2cbLJzz+2xRASpw8szgmaxZ9qB8JmVWcNsFMP5MCH7qlkD2ffJEVsyxsYm6VI
6TgPxAfi02Un8ZtXlhG5EEiTdShQKJ1a05gUb6/d6tOYnOrpIBJEBG6FLCUWJ5Zd
07cWXt4cEjg18Hbl5sYNPPC1WeMSiEIezttBrOR/NVTJvuhSuka7UFhVuIsx2wsO
kj7f/yZL+4Q5yMqVVA0qY2RyVRXuFwnfSGqfIYOsroz5dES0xZTXJbbpcmH+Gu1+
CecQtD4f83RI3NBWui4ubztUDztXgb9fJcbvplsA7c3AC9ZrvEdPnh3jxK+BUPbz
4oWnOyR6WwoKjdWMl6sHqXTvMb5XSRUwIOyTVUv/+Nok7iTh7vxeM0sJ8lJNAd24
cNNTX8aBPWGiM0XJzODdboY+M7QsVjQ5humzNpTgyhF6eyCR/DghuMspFeNXgI5m
WPx/mfHpLsUJhQEeuqBf0/LMMVNun6cSTSm6KFraB1Xl0l2JL4ClzIm0xnaZFGCY
oyu0PfZ3JjxhPUKvRhfulAYxy1nY8uWDNnynSNnuuAjDeq2w1RefFKBIQHnkFl7q
4WDFjmLPcXqkkuwqtlEezA7ib47lyADD3lOLBjtOYiAdl0WX5Mq2DGhkJ08PWxk2
CH+gUF00jU8M5LSQVhtGzAhB//pNffHZ14tFuhcLabOzLGxG7enCsggOMmh60Tk2
25cFJMcSSzlU5maBPgjjalZkK9g0sSmTkbAB87w8Q7LDCCYDsL4lqBILTEkWMl9G
YVmVB/Uf9FUSrSLYFXOAhK7rWQNGltMKo5kNXGXbHj0uTxcQ2CYzzAM4bB/WKzzg
4hnDiNxp2giV8CBdVBZs1kxzBaP7Ox3Tf3sLufektCQ+TtB7k0Qp1WX/E/ItHQmD
4aqcoQphHm89VfcoyjErpCpGued1noj0OrDDZzpVyqo2JSlzRwoG33/NiuAXJZlF
lney9IcXC8ctLuGKhnUks50cikA1Knv7QuxVsMfzpsRkZ2XL+QSi8KBL0TZzxA7M
fZ7xC0HCWKkM7C+C0PptpQd3IXPLj10a5QehcaIFd+5m0AUEFXDUlfHcB0/3GlUE
t699zAkJD5Wxu8kPlHCocgufkdSi7tshfvbYLey9xvoqBKa0MDXjhWR4UYyILv53
fNJof80k9z9XgBQyxgKUc2q0xmwnfD9p/2ZuTc0HdkMzGCTRQhOkCD/miowEk+DA
8pVhacVSg7+dCzyYuV8mq+0aogQ4657aqMkq+4Dj8+iaig2aoC52LCujaFtO2w3S
oqLmnfKdOA9UoIQSkmK4970Qs4XxyV9vmWI5yb2PVjRL8Z7w/56r6Pk1Q9B3TpFW
a8phCnrZJmLX0iAwxZbqOyzUqVTWPcWLNqplUH0hOR6RryH80UlueXl96kWaj53o
Qd3IjPhDPZlEIM1Dzxwj7yOMtpTQNXSpRQa4JzD11kbTj1yXr+Dm2649+zSPAwlX
Qj0N9Qg02MzTXqY0fF20MXBI+gzvsEyGvrQcj3Ys4sqG3UhyA53N/n06RRWr66em
P1PHDCfBogFBQHmP5lxevTZRIKD16BFMkRXEUHNiNbDDL8U+4yd8gNikPKluGGkg
BwsMS/qwgvl8aicXXRlFRsfKjnDDthA5hKekNQ0aYJikooOT/mhQsCE6Pgd2CFJZ
qAhglzrBfcO6ONmvY+yw2PVZouRdGmUyjuyydRoN7jJrlecFGoKCrhn47H2+DT6S
QdHOohBd3KaQalsQSFNXKGRQTuaTaN4IyN5uWf/6YDOzYrt0hBmg9dmOP+AC7eBA
+d0f8W0btLcbFknukaiFBcYmtptt/qGu9lOzNtETeaih1FrOrBoYRkoPqH7loCg0
gO1D5fAwv2erwg437Xm328nVXzmKUOS0VGQVc4hQC8G2WWPMaQredx3ayll7ORtX
fawTDqTVEblMqmQc3Q5Cw9LmQZDzsGrgr0RJQYzYS7shVpAwEhSSzIo+b1c/vl1W
bDbiI5l4hqSQNcC1T8DSTi9MNO/O7e2Q3XvRI0tzMKluLthI/nUnhyRLYdGTdFOZ
3cIBrtJEsMj1NTo/lT2wzYyTY2BJL1jYJQlVKw2k7j1bAxoNAHBRO6SMgO+O823s
FgJBkPL96jQ3/7it31BOsuObfcynuTXFvtW6lXWzmBaz6XiyDsb/wYxV51vyvfAB
y4ceqwCVxeiMiIpsypQQV2vNmVNkHFvhpEMYX+z/MTH4F+mGKM0O7o7CIvOPl7kt
cATNerkgHN0ERpj+VsQ/1yN5TBsBZAPVZy3QEU4DDmaqD6eKztqLLmEeYJ9d/bSD
kLdr5Q2wzr7gJ87tTofNQXyERPxLmmuyeRuohnIagcetoeMkRlKsmVQw9a1cuOuk
Ht89nMN6if3zSIjn4db14u0TfQuao8u8HMeh9JG8CsgV6dGhydEH3Uha3o3SQGc4
WLhlfp+JSFK8Y19X5zOoOwJM1C1XRa7K8fw/svHPO+vSrhbV5uOt+EvBk8IiiELL
x0gCoF/ykL+BTN63D6gUT8xeV2Jeop8HSRXxuSPoIy/RwGlfUv4uW1YldBQTzLi7
fsGtzOKfrcgArAQiZAfhRtQ35yz7zJGMPFZudn7UJBsckRPVr5fHUR6gdoU0MBbW
KC8g/dypo0IC+6H6QO/hb7qO4jH7HkxE7j/I2t181wKU2WF4006VsKB2diy4AT/u
KeIlgy6YEcYAUNUXpk2oi82GBRnmykG8J7t+CfVIryHXZelVwFBi/Gdw34WGoieO
N3Pe1YKZNhFEQrSuzHvyFo+Pe/O8IYxNtUsCdd3KAgGM0+r1Y0ASiG2ctHh2b1GB
GOWbVh7rY/oQISfmukHu4wJ6yC/UmNiemF7s3bWeuXwnskVGSg09gfIqNTusEvmQ
vgr6TZh5LAk0rcl3uZITQ2E8PKV7A1igCbM3yiCr+rFjflafAXnFwju4jBBw99gg
ISVMjtDmCIzwuieVhK4N34zt3fEYL5/N18K9csTT+cbUCtH2MIlynVCx91F9pUE2
9hxLG+wYgp1AHsILXhZDe0lGcX/B5qrSHsWDroldG3IDwsU5pmmYHsujy4pup6E5
ZTAKmClzHz3C7yCt0TNiINGsz4tcGwBj0NdrLRI/EqEq+suKS7xZ15xHBWgIUMyR
J7HS6GhJuJN5vj4zmX9nP9BandtAqXyyDQq9jiq+vI2RLokwsX3g5bXgohMhqUs8
FsbSiv7h9JZFJ1JnAM4jvBJGP/EGuLQi6cI4pTW4OuwvIzgGah4lE12kGtO1ExMz
6CgdQNshrlXX4T8bxMoPAU+hgvGORRjYAm41g1ZqjyZ9RkxjFJj5rAjNSqusBaxH
Ly2KdwkLdyU6AKk6hg2jz7xBLbCtdg31HytJEDLHQiXyul/UzUT0umX7ZnlOW7o6
lN7i1mYcdltXD0la6uOe4hS/1sfrRYd1JNbS3Mrq7MagKaygdFhHKQqTqql3Uj/d
fYpmSBVUR+QS4WM6RCokRt1tWSki3ERghULGtnLiI+kxQWwET84FyInVXacUN78x
fAQIl8mKidJ770QLyCTBd+6jk52KFgx/4hdUwfR/eNFQHF/SAYr5Pyq69HgRbA4o
ntBFNdog46BQQ1GrtYvwyOHINVicNXYDaqN/bHzO1taew700lxy9agYHV6tmXwo3
SW88/c5noAaRhdbg4Rmf7AwaZfQ5ygQh2Cr4+uoyvqoKKWLbs76xmuy+DsDXd0AF
sodbUI8hUP6IdypLf7kQa5YG0zNpYfyUL5pa/hvJMX/7h4klHeiJWr/s6Zrwlmi0
giDE+OPT9tHm49ag8soOgbUUKR69Avr0ewypk6TGdTaXoGx6hXuzWlcpvr1o+V/p
3yTqnNM3tQQYKR3VaoxKHWZo+zKDLQXs0yR0KwTrfQOKiJjekSqdGTzIvbw7exk3
Pl37ilOBQQ5FCNUr5T7a1PIAgFpbhMhAgtNNnX/6CZGFm5nUmM/myHc0Z6+dicZg
mWRlrvwOOgfuxxrY+QHqVpnKGsM6+xdfXeVUK5Q5Znc3mNuHO1oicFlPVu8Psu6U
wJk6PQLydThXFCAMI93kXDahXPZT0NSShAb+cbyIv8gUtfR0fGtz7HpJ4/Qrlugr
1LEd9JxkID/xtBOQjJrw8+aVAjC7bzAAWF22DeuGJeoJz3F3185J8YNouB/SE5Bk
F3K6744WKb1QcI19CwSoUFF8cjKktF9B3JvTxQGWw7StCUwSnH5EQVahl8vBXeeu
Pj9RFkt2MhQ5R0DAVNs0uiCJXuwHCDSkkOXC2VRKqrdXwypuMyKqlXowDB7Y2gF4
2rQ4qaqMvCV+8SwvospBb42Uyz6GPGiUz7vrjReE+rPYLJnW6oCJnswdbXhfMMiy
iTFq4qXAWFu4v5SR253Fbo3OoI2euv0nyuOuI7LiHfSfg5T8Gl5ZH2s9BRbLHM7t
Gm3jFm8ctjmYTIfXVrNYkZrOd2oXxl5nK91cMGvGet8K/GAR0St6NeLcyreyP81C
7mGL180R9+yM9fXOqUp16ZlfpaFsr/V9XP32KUOBd3C9UMo6KiG1WQL4RYIRQoFJ
GvT/Xrg0WachqXKuUM1bSmNm+VLDZIAlU3TEQYMxnycHhnrSGetq46ktu2up18qq
rV8/EyDzdIYCzS174ksP5g+Kk9dWgjCM6ycAVeVy5z6ZqKfwcmyE6FiB9KJdne2F
iNttWHnwJMRias2aH/fywsOS/u1j3a03xLyoKV6bb1csL9ri21yLYZEM5EfvH9sF
hStC+aydiJsdDN1q2SiNBMWAoqehGOxDXPUSFAx/KDAAkU4kjsGNEf/dfbsRPP21
0Dyy8awOWSQmaLJSQ1yBqzuWsvxdLTN2wWh3RHXviSJrVE/8daIUtoWx3XesObEQ
sLuh5Pw9gtzFPfFWNhJmh9vZzM9bqcs05SrW1XadD5bqpih8aMevbdTGG7t5kn1E
4Img+KbEvXbsoXq+ekRRJM9Jqikq6xPgkh83YnwI6RaWc7o4ENSuscoSYjvZsTjL
eQpiyE1gZSk++d9PvICzLNSU0m1bYYBkkobAwr/iHTOgX7rRWOj6rBm+RzqPf2AQ
7OwhUZ5YIeagQ3QjKrN6iPptlH8nn9QoN13xcIPXlyKIS7+DYF25zluvAcpHEbP8
h802SUMyqOcizqQ+3U99IFfCs6Nu2msAZH363Z9Xg9zKEBtWzYEVnjNoQKJKOqRW
5UsVT4wxYN/Y6reD8OeGS5HJxyqXsK7kdXRbw0wnMKYCcCj1D5/UZJSlJj4xCaT+
u2TKyk0oNi1d7QEv29O3aPPW7NehcC+SHdsg1q8vdnRuLfJxR45aewOykXhFcwTU
ozv1gh9GnHfR7AdCp3J5LaJKyTzAkhjus8l8tp3VUuu5HNL/uw3TBWVth2pzCojp
a5+kLmdL/mdIxI40eCCInkla8qskk03rRSByAf0CTG3Zydim118qnYv4WkUy5NpX
JXbx6BxfFaGCsUQKONTg30FrijiDJ+89LLV13MywL+3J7DrjpMcDn+teRCgpHDL3
v9x8wHAmXfJoxJlW94JJ1ccZNxzGsWcVLxQGyi+S604zsHA3VFtzgeHVJICocgUR
mJvZlir3abcB+xFS/C9thIErmtUtM4apcR7wNHf478O2T6DnXpIMc6cSb4kI0kxE
bdCwH9GodFVnAW2IrcW4b45qBnsXvK86iVY6rpdePdIdfoC7QSpdkiCPXucaYzSO
VVghWZSCd5z9npbHaVVB35CZyz5u+O4kWpQLVypk6D0rtXFntFHGiKxs/2Q/D4hU
TIlJoP81514aIWrOOcJUO2LGSABAuVDPl1I8rlIUoHSQy5ZbE3s9NHK655sS95gW
mtSjkGHI5AfyRiP6nK8VXptMyBFd7jcPI1JewKWwVyotLDFjXFlBeW7ptmg7Py31
RI0OIlTZIbs9/Ecq2TBi/GennVJuF4+GtBjJVXMfaFOZOcnxKIBwE4wqV/aou61a
jz/NE2gu6So+uLZUlV9gzOP9d4Qk2S2/bL2LbnqXvEOW+nQdd+8N4USCNZrn46T/
2Z45ucDKx1Z7hgM3S6PpER7tZUcerTmAKxIenOltkUYzfmmIC0lcGoOxN+MWHZoM
lykdTtXrMonkzaK+MaJL6NshdORlWFNGeRcBS3TzLY8HgCwFns+5aSjSsbw8/s/S
+8hY3MkiNJ2J4CSMQ4QCSEQ7twMY8FjfiqgGwNjgKhkJhFiv73uJNtTIyo3+VhqU
4GPZzGZPdYF70ItdqkHUF4erHyf+96DN07GPQP/C9ODQbm87IoKvRe46Rc2P+0om
/hMBMjiNrvFAA7fY9ab5kL78CTKefd+cCjIsB0wiBFYiAmR8Hg7qYOhlkoX1n9DA
91Kejn1dMPhjZZYLiTHDtLSW234QLfPDNKDBJ73gh+ZEwvCIppquRTQ4EPOylkkZ
FDTzJzz74eRkaHskXeUD2y6w0u1HGJghbmkO6aJcGY4vR0FIfbgLcyeEYlUNcI8j
1J7+IsnP1gWvbR8H8ElRsKSawJJw+hVw8LKm+8khobELAXXK7I0dAHp+iPtjS/wE
mSvR6k/vbJa6LkzTiS2zKN1wcr3r/pFrLLazrOavbdLXJKH7rI6N2Jt0CxQA1/e4
Wkj/U/N9mo5n7MZWQgMcIBZJEoAXHMGkht1JUq5RwkanR0NI1KbKz1OsJY0VERDR
1e3hgci6Rg9lCAjBN5zJ7qksTtjzEhfKvKvMvVe+kYITcLeWJT9Ccdpv0l8Tjx10
4vdtF1qDVRk+o8wdZ3Wi987N+1TzOmQdNSYvml2IqDzPRJ+8hNXSo52kUYJ1GpCk
TH6ZiUmiUNCjkJLeoiPFOzlBsYLL+5SrSHs2KZ5TfGu4fcbdOka0O2esT3Ck2kxz
drXccHa/VZUiTwBU/Wz1aBr2NoMw6Itsh1hv4fSay9I3o3r/Ik5sHVJ83o9uP0vL
Z8Q5wb53zUjdFYClzU758W4mUT+V27JVjds83cncTln+z6otWWbxOiFwrqU8KQ0g
dZ+vnvhnXDl1pWqnrii8xGARSA4//nAazOIMQ5TgvouuXpTFr2C3UdOZ8tekpYBO
AYBZxXwCTl9aGen8thTN+zTh3e/RqwVTe6y69LVAEYRJBEFk0Z7km0OTZn0jZa6n
yDO75GtZf12/3ne+zGnycqahDmpkOOIPDDsqSrjXh/DM8ynx+MVj1CYyVP7px/Un
TiGg4y8vDwCCynO5vSukPvy5reUBPFoSAoNhc7rAoJXvONvATPy9EoUeygQhILqR
6VHBk0vcMc85qGazEh1xJjBjlzT5Jby9Op5MM6mwvg0KIV4/AUx/HaeaiHXOS0m9
SmTEFtau2HSLoor6TeeX+GbHEzQTlU24GhHHz9jSVH8rz4zwRiUfaCTHono75T0Z
L07fRX2/+1o8fs/h4As9SOhA7GstRYcHZYXZVdr0jDRbuC3s+srBFu1BAaa/1Jll
BZqGiXA5pMBp14cV53V2xsr2g8m3kZYPkxNU5ttHszZ+uT3j7Y7HGfA1zZiIFJEc
8lv5MiRtrOjeeN4nz62zBVPK/rvnadOn2NgSunHAe4/FIeR+b77Lq8jjz59LEWWS
o4xC2jwrREJKqqHQl9iCBP3eK5ZE+x50o7Wfer4VU+EHbpXWmSjG7eKu+46c9SzE
tYcOei9yB/cGkIf2ZjFuujsjEmMfkSUhC2v9tAFzNlazAwDj9fxf1Wc9Hix4hg5J
ZQWKBtnFBNYt2w8/lvWnSOXLL9V3D1PSaQ4FBbChs6T7H7ZmUixcpqjWZVPaWSj5
cE9cBeQEpghcB5K/AZtcoD73PIy8qGG6KYVb+obGZbtvKDmzvu7d8/tSOMYTVmie
g+XpNeF0uxKrrM+FVfkfJa1/cvehcKT4KmbcX03zYuwdOkuEk+3Vk3+9JVA9WZ9y
NHSJkDdawtVDeqZFuwwkreX3NHhteIr1ipnbszwPhvAU8vRRu4sx+XzKvR2xuE61
qOPhPeqdrdri43eu9a/Trzc795Smy1JIKaLqok4l3JLvrU3uavPAq5Nc+vxIwFzt
zvpV+x16H77O+E4hafZote7JIpHpWIRBb71QNA180tIcOFgfbGp1iEzr25i1RKFF
nLq7ggm9rke7DhPoLoFGZavwxneZmWF97HRrWix5fqHNBG+X9wk5PjkrBeQ49RZw
rAM05vqzpsETa7CurirPz8DPFbVF0qpnW6nnTwPFtU3ltDEwZ0g4Ghnkt2Z41Y7t
1+cSUhvHEjbq895yoPo9W8ktVUT3ReLKbrkzphvuHRGjJb5qGAyQfoRYfFW4upzW
7QHWskZJ7zW4566wvSAnpXdGd0N4er1kK6uFYZne5H4BoQOVup/4IPsBIORbyuSy
K1GD5HtOeFnyzWRHeFwYJJJ7x59rzpwxdks37dzAvAhxvu/1B8xhVW6yIs4OTmZz
UFVH2lJGqy6GHT4LcbdPgwMEJXn1v0nS/ebbQW//HXd7gwLTyLmi7G/TYbQZ588C
lUFoCptnTzWd6L1eQl+5j35P+m233kC/eO1D3xPlPeKpy2S7peNiP3d35grvMpJf
VSurFPDyiNcRdFc8YFxZdAvPBfTDUPPzGGeJtlfL1E5GGVgP4zpqYywXnb2kP081
rz1SnyNCWaHEmrLJwkVZfhs8omTrhNv04db2i0YT93yN/C0yU5niPSJhyT80ynIP
FE1dWkNy6ugPPuHCQ3Yl6R5OTGztkcAZ+gslEaZEMR5xC4/yuHssKweel460LU1L
YsxQB3jfQ2IHYJ2Ks21Wey6j8WW6v0vc+W/wjhUBtdwCQVkysQocn+6ITscNgO3i
ru0bjn7M1x/xyNCrAP52t0q4TJMPV1tObzPxmyXbw7j8fEdQhJWbS8b7eRg4UQpg
oTe/vOdOCJ3WPtctHPV6T7FPx1KlQXrn5i5nJL+g1cBX4qQ5rlJT49ZCQrIpuohQ
8EId1eJNGrKHyKQHL782ymjjmARdl0mKrvClvGSpRAECLniZ/3pULCLgTjQqnU3O
hqB4q7rikM4dURS3NwDMla/oVelddQ7ZRmSX9Xlf6khk+2HmpG5R++00Ccb8ECbR
an85jZnI9tLHf7q7STV8Y+rktSrpAoIaDWHiF5WzJzYQ8KU1aLN4jtgbH4cGz9zc
/kc5tbeZH0dKEChd5nGN7JuB8VAj0SsyxSBnUeQZEqtkbrypiYKjDB178JiIDrVa
rrelkK3yVM59gT2WE4eaIBMk8OSaUcXQg9uLFwvatVqeMBgeux5os61UX8OKGIeK
fkH4kMTqwAx/cIVEvFH0TWyP/teZ3F3JS+clADtWgZDtI4RsHZ1RrIs3SdphRCrK
yaY8v6fxcd9dNDdDFoHFAfNJLH2WdND75LHZusewdVIYCvcT8cIq3WNFZDwREb41
futs36nzl9USDlhCwKY5bhxcz+KIZcz6PQk7soPKBewBhWxDQYBF+xAP4SzzrvAY
QSf873DTbKNTeRzlw/eR95sgu00qHv3h2feCEsqOGlH8i5wIXUedFz2UMnP4KVQX
vtv0vCw17WHtcUHdxHz3QWC4nAYzAnyF3VnOzK0zSQ0WRdFh+m4OUYbwG7JwFUDk
wddFTP7oJC9227NlUagyEGe36uR1UcmKTWiNBTj0gYwnPfCr2JCzxj3POZoub6CV
1s6AESUrzcOYi6ziUjz4Yxn1DhQ4HPzCl6tbLsn3whnGrYERKuGeyKzUdQkAi6bE
RjA63kcok7PSH04SWmI6/ykYxTEBlhhNYqS3qU6yIM6Ac4ge9e/A/7tBFSRYoix6
P02zSAVo5lVdOQbRZH/tX8sq1M4u9HuDaGfg5zlPq0/nBdOtEK72X+EUg7qYIWdF
lDFIKyPgw8+Kpr/pBanNyewZ4lYsqc5SUfDXzPY8ymDsN3Enp1/irlU8pmqFNffZ
UDm3gp067+N8X65urUqoKKNFqNINdOh2OW8pV45QfCDNE3pzOK10WLQ2KV6yQJJV
OtzKCS0DHuiu0LfFolchrc8OVFVG8JUkj1ETEwuYsIq+4h6UDRb0xEmumV8as8FQ
xuFBrDEn6nMzt1I9IVC7ujCJhx5tE1z+QsR6v99Bzosycf9DxJJ36rQhci8c0+8B
IzyHQzoenql/SUWe20Hko5HdZemMUrBZB4gZCUqfa7Ehn2D77XdP/jEqlU+pYcBO
dgmBcWlbjglbd5p6FFQs1D6d1/5hplTMfxOkzu4h0feYnMFMBh3HbOijQPUm1d/6
Zm9JOw91CwZ0qo33Dck29NaAkzKWXA/sn1uBEaIgnu/Q5rLl2sDRhxQvJqKKjtqQ
PS4azTBfiR+h7L9oinCq5NL/XkBjdxFeqojv4HpoVD5lfFqJ9vseS3H63Vvcp4LX
ZCjSsnZAZ4ctvrmxfXlZv9QDnE4jfnj1wxJ5rmq6hKpBe4C+tUptAbjJ8TsN7IBW
ZSZqrHF1rzEDgLS3/DEfGoD/hTG6dmbHlOkvAXiRGIBorJcB/9FC2PVF6dxwky1g
M3CpUeMcp0Is0yiCM5j45GK04NzjxYIgYsg0LoFZxVS9rOWXpk8NdZriac8Xs8Jz
cClbFrNcLVj9ZG956/MuJlm0ge0bb9ZlmF7hfJol0Op7BnTbFgD0/g/xzBzCcdZy
6iQd1/7z135wNj5sTsLtGbtKhOrpbM6/q/nY9px74QzK/FKPCj1D4UcKRrXom7pQ
2Lw1xJYC92fA9ZJ3v2GNS84MghzKJ+jNLYM/A7CZp6K3ql3jnd/PFBGViuNpGp+S
+Ors6RGbhrLHJSxUlPvTu3Z4e3oYYamtiiWOiU0KpBmDE/ceHaEoaaakCZYH1UYX
M++nQ4vzQXbrI+G2K7b70Cwi1obPf7570/uUuF0vGM4ha+2oMiB1SEaPCNfQ5bGG
WPhCO94qnFHUyq5zlrL0TAdEI8MFjvkLC03rjZz8rnUgPDXFD+AIaEsR5g51h8Is
saSUuagnJlo6S+InYg5sgpYYJArmL0XiasEK23zBhb8hYQe67LUuZaSeMNpdgnwW
+jNZBtiAraQ5THT5NZKtMUFrJLzS2xnz2Evd95D4+I0FOLXMN4uc/UYa4wKQGEWu
Twon1IjDeKcHdXviKj+vKCdS11nEjcqfDUAn0kLJptQO1O8QE3aJvNphsp9KQ2xf
Sr4lwvzBqTh6gJMEa0AMgVmt3yY8durWwjHs1EOZxzs+BAHPyy02q8mw8TrvCISF
vqNyH4kwcTcqGOvfRm55YREyZ4WaTseTNQr7kLdtzg7oizriBcQQSi26jf5GkPAy
2jKdrUPfwQx2kR/E/xrDUEZN23KTgPal5tJdcZC/irlcjkegR54qZnSmA5t+56p3
3gfd6f7fC9sIXsLK1dQnzNAMQXcGIzqX9T3WffcqqlEAYOr6yBG0e+Bt6hEGEyzG
rXjvwd3/M1q0mQj2AafT9RYChtcKFSvuWr+WDVhkHHAvJlJ8SUymLl/5ZheHUR6H
bHv2ysq+DPPn8SESOySWqibzC+VZeC8+hl3ntMZlVYHX+dSZ+Z7GnuWT4Bi+N0qW
gWN2sFkzfSsY/K8VFtK9rP8e3/SyXwOqToWLXCQBxQaN2lsZ/yXYa2hMcZOPR1oE
pbNuJcvAw8IsAZGhA2J4UtkvtP4tC7M5darvDhXXsaP9Zv9Q3mWsXstqDCBsPQ8q
CRYsRZD7L5KbRVlKhTHSIDjCUG1oghk+4eNxeJSB/XZUVwO7wk0jI22CgxN+QH3I
7aCl+WfPofCTfR+gvS+2rv/qaLDEp6mnj8OqXgGMfc6xe/Vj+aJnpzZ1WAxFpLOf
BHYcypX/VTK2wc5nGZ45vDox2UY2trKoy7LN6i+tyoe3uYLJi2jeLooyzvkCwesD
P69m4YakYbUgjgjrwczZcS++QoG+1fuYEgS1mNwoN6b+Hqfu0QNl/ROmzf2JC8nJ
CJvOjaxUmH6J+7HkXfSxi9SMbrkB2OI3hZFDkkHAJU1aPY++pb8k+M8NG64ZuZab
NJfDD6QCd9LUPqu2WSwAITqz+BHVKyKWF9PnGQcNrrYEYvemub3JoPRycMFoZc6M
hTiDOC+dA4mbXc3/464pNuPFI5HHwNMHVt8DCu1oUR6P32xc7LQzo7sKzrg+wAPQ
/ahQs1N4i+dNqGUUAbD7izt+sPQwXIccjZjTd8NvCFtX1ZKPJjt4V620YQmDc0ZU
OyuoDmPjo63aMwe3qhsRnjz2drHoi80jMBP6BEyf2Pl9gLzfhgp5Ykv9slkke5aJ
5rFaa5LtyVDU6mb5VmYUCVuXB7T8/ItGNIare+J2/OM4MLOaarlr0KxcBYceUV9j
WitKzKPqveY5imobLR/mNn3boOyUZBEW0KiDC+Ljzlb2BOSD4UV9eKHxkuXgWOBI
khgD1xoDQ/xeMIrSuACsfHIRlx64nK8pxbtOM6OQEp/fzncO2skfofJt6B0R+Xn+
Y4szJbQyDiw0sSI1iPwPfUXJbZgU/LuIAmo8NDq/r4dVz8KbUQmhFswVJFMVrduW
PDrnGpLns1aDNAUfC08mDWKa8Z/EVUEuEfTg6KxEWoZNkzyu1VEOBEhv2zuZ9H8e
X/QkKQYJWRii1WYrcjgWl4/FSYggDZBoFBo7gagSP7niMOfPPAehqFvNoCNqxT5P
fAXWhnAmCqpZbLhNAZJrdi3lLSJGr9cDYO2d/Pm+WzoVZrU/ZY/hKGPksVxLAqRs
5nHyo31U2LzkywT8l8xf9eaoPtTFY/4evzvgZwD8E0SkmrLqwI4p+CzsBbV8xRDg
x2dF+IEzo7aguwtM38QKN3HAEJ2fHEndKgfK2EqTGjBUZePUYB/qQZflBreQjJQp
2QycEXHslYpx+9AqVraMoealSdC83hUH+jQrXhwkBaISp3CXYHvW1yr73Wxnb1c1
Lw6hhhPMehdtWdKLsuToYmadEa3upZK7t3hJfTg+5SBpwwJcXS1M/V+B6zuLZI6o
2hoebO0lXEOJdraNDO8zuhTr7WB+d5auC/qUPN4PemtR6HGr8TV8zinhFjgZPqls
T32yYX6ftE0Nd8myHYyPkjqdblTlh59PbTI5S9dir9YPSo5mgBwVezR8+kRjPh1n
LZLQVa4D5gGoUbi7pS26dIDhwLq6J/XnmCvX4ukSjiqnsrLLqRdTv6qt29Dz5s4Y
nZW7+MOYCvh3vCbEIkN5fYTJbZyTW5CVRkRm7jQqu8jvAvkrKDODZTlrBh68AN/W
Vbwcd2NS9jrZrhYf6IkYXcJqWuIYXXMCdhSl+/szrRgK2BfLtpqA3KT+FAHs52cm
eRJcwp4ThRZAuL0L2arUoSk57LhJBSjsZTBBY4dx0WajEq6Qe10e+/nUbBj64TBF
ypzjXS/3m3BJdDC5iHLVolHTU9Vqg+xsDxE2fnTSf0VnhqUX0TXg6Wk7Ec0T2U60
7oIA36yVFsEEKZ0yaq0cdJFx66nxvtEScG7QrToK84nLzbvq2BmHEuz/piCD5PkT
hYSlvWPTaBtLXmDa7E0xNOXnEvhAmO1BrWeoXOUbogcyqek8YdfTJSw4j/1KsrkR
Dz3y8F7NJPt+Dt5NIUG4Ot0jlRQHIQUvBR0hgxrua44I7R5al2cNGc1RvjjF/4PA
wdNhExhngd++yfaF18WNzDiVHxH/naWmfGYKR+qyKhaxfd2qkkkfBZvJ8k7HQr38
MfC70IZfQas64rNBU2rgXYN3ew+9+H+CAbjVwFc8M+SzFXejut1ZCzjTpm4ZbYZK
fo2ssK1fX+axL88AlCe2GvqQe2Iw6iQl3ppeLmAANnZX9f0STHdsBate0AONEa8s
TWTOIA1HRkfSS7OCkuFwF8x7H6zLK/VGg7frQd1KXTNTmFM9Sf6ovvFBaE++aDui
98+UcAOPo3O6SmyZaTSQjd2L0yed5E0Rk6E7rWxe7sBGvEfn45slpOBw2k+H732O
+AYm9VkfJqPt/WEa24gcfrJ56YJgD3igORc2FwROG8MVNmy2aPzB0hcqgn+01O8d
YjHw5xNTdorIxuZg7JA6SdWI0RpddW5QpbLl/ckxJ17rvp2kWKHnXd4RAPoVAf4w
WOaY16w51MECXDDulVb0xrmFj1Q6FtX4aTA3VgJTquF5DBL/P8dQZlEVstw5UkzC
6ay3vt2nOgpsyr5Z3uAgYXj1mG6OWw1q4GBhuLhTduNre3LJ//pBQHPsRHUcG3VK
UvCiFEVKdgZCqMoqP1Tfh+kaNzFObvMIhAYMKL7UZ2wXXKMjGOMBtwn62Xhxawq+
KbXUmeewRj/nw6CoWUjxNeC/TVLyTzVbO3ermUx4qNTeSKT1y+XnI4zJtYem7Tin
l/TkDJN5BRsJ2dxcuzShRmZ9KTh/NJPL1RWWfSNxx37DZoukRvoKXofJckCxhAKo
mMxXXnJ96g3j3PDESVLYG/ovtbvjUZc9L4kMwglihpWfChB65GtAigOhkud6xOtb
pmpiK2CO+m3BQcW/4TyVpOUwLWce2lAVlplvIq6yrcYWhAUWkwKqzfi9ryKbEAhr
CougR8oOetgoPu3ZzF7URVRvBcV0nQimnw5t4/afAP3hskLbP+MEiHzgLhrArPe7
Ug9tVJkar4u7tsLuFt5/rEP6kcKZRnnlUwEZ2NFvyYHRS4Wpv1ZuAwcNJtHuKcTF
ee/HOLxZNNLT0O1IltcHUmjbe0pvMPCNxWYFEH/eLrsgVLj4wDyZc/hL0/2sj4mN
IQtAX0Xu2XpOTbnNnZyeg1aOlq40dsQmB0dbSzDtZc8NKCTDWV2WQEUYxdijGcEi
0zMMy3bqNzTmoE01+yHTbmnt0TBfTtX0YZWEzrWii2NAmxNr5DQDePlUlamIvKB4
AeU4yuw7gGHG9a2jiY6QBdehqEyb310gjU1OChnMo7Ska+kvTzkXadVq8v+HiQbA
WUnQdRC3j5J2HzpiOlI6TiB0qdtskHUcLwsjkNDj9O0wBMaF85wDLjVHlPS6/ybF
RYaexF3bTKCh1jzKyIVBmSzpNQ5EGGp2ZsAPgvh5x0RS3Ia5XQ78x/qkbDWXfGaH
5AJyCScAATIn4p4DPdPB+bzp05V+YGJiDnZ5KspiZeZ1skXj511KzjwNArHh+9dV
RGQnG5zuMRpHdNsK6CpTt9ROyNyWBGCy9RvOnciDznPQPtMTARcQLPi1x5GOYJTj
t+OZEL7zA768mJxNd19dJaT/J0BruUVBdejBBJ0FhzLg9rFgiOYwRp6I/rATUsQ9
ZIRj7OsumnvVsC/BaA0+U8hDMhdoxKcMgXyPZHfnx8wKdi5MQ+GiqwGLRnmuOgSz
N9yVkp+n6NL4UHMeQXmAKvrtG3sJebTR2RJg/HV6vsv4WO/CvBWJQsf3BGODtE2K
iDxim8Q2Nwg4ME+ZEzVJ+YGE3sDQ7+Z5hnWXdUxUbwuPi3A1F1FFSuufFbCZ8A/9
QKVWeQ588RGzLbOeihAabUVOM6/X2rW0rI1NZ6ZUmVW83MMNgLFU7asjRjCnggeS
Xu6ChWEMDu1n985SdbpukLbXzP5vp/aa4zr1/OhM3SgE2j/sDuKdQ8Ka4QRP/WT4
bC4e5y0eKCMojNkwLL2CHiCZVHseimReVIqYs4osLjLsgNl8zXvlEkDEiT+oCzNl
2FB885VlgDEkhSPfV+xo8drleRlt7L9tLa+sbHOuGHKXmI3OV+9jThbNkIQiDytU
7CEf4qK/bdupwQVbrw0U4smEl+OCt3iWoJcs8WrHGHdg5Dc0fWhNiZuSe1U93Oak
qv1tfUXi2eE03V5vQUHhOaFNpFCh3A6+IGiSsFnUkNfDyNxZ1W3J6vLnevSXHDEB
WSdywlJI9ooMw0cuwazmrNZ+OETpJOSVqLmWBRMzDVy86+NlGo1MdLtPUzVkoFA3
xLngwCg1Hl6lZz1cfoEvdO+LxUuwLgkZos3mT0D4LwRDpxrrStCDktdEbxsOOoyS
xZfZndzKklxzf26zZTrDXHfw9meQOovhQIdkxBiZ/f941SD0V6BUSc5NCCUOYHC6
jOQ61qwJNikIlXIJic8Xbc2I/l90ynGwj8QTFkCwRz5QT1ZVVDPrJ25xyOeJ8s2M
oH6wX555eN6dW33575PSQOgNW96DP4s8n8uhdOGBbm2O+MNCFkgxTSle5qHqt8tk
fJzhHDxqaaywbHWHxw1h9FLYPYbNlU4+X/VIAKyhA57WDsr08vDCh7Lvz5OoZcso
Qitb2LsOet0CGRcyV7KiI2OMuZKDiPcXt/dhCdbcsuC0Mjg3AkqG5bGvhlPLvn2K
R48DGQFu12BDkkCsotxuQnswnehGoh+fb+KwCUiYjbOapO80yBXf2ICqWgPgr83K
mm6YnBn8WmeCVFZkd8avp1Mm/tnaskmV/+hPJB4ASvHnJCBWhmZKNRsPo8YgSEo3
IaeuY4PDnTDKbbtZC9NNJQjWoLnzWpcHLislHOMBEwXmou0dEo8lI6uQ0E2o/lsp
GM5JEmk7Yz2LlB5wI9c3G00cyMVKWZMgJYHC5KC/nKwlfAVjJUjpqqDqY/ERybMu
d/b5CYgx6b9lxaQ9ZXAMr60FeK8yPFlkiaY+CrD3rgxNDhTAQyq3AAV+H6qdULwg
pyggMp7eUNW+WGyx+ytIWD+MfnjUkiaDeD7Yzni8HQuNdAD+sexceryUmsj7Dx3x
HTAdjTCAHQ+M00UyXmV7F/OHV/Jlkvmc668v+EvdTS9A0R5SJopYq8oP9G/dh1Pf
yaMnWSF37EkmYQVd4D28GqruFC+TUh6ZiIZDTIXwxPeWRf34NorFVk8fSjRrX/Jp
Hmgu5MjJ61G30RnZ+tKHw+RUInTcv2zSx9as/UIgGqKGibhCKbwmQGVwVagUo87z
WpQL/vIAOFJHhfepNOqfAkO1NYMUDrM4j45RV53WNZ7VJ7iFFsRKzUeCj5cqwV+L
hq7M6pA72ol6qNHloy+Hsr7kRWRo+pQat72/h3UuxNw/HMlNfDeeE542jMRJqXnh
jxSGhSBpbBe4f4gcDeS0nzXvhRgoNG7T5GMWcqZIIHU1TGKcuOwSP2aErSD9KrF8
u1BoF/8MVdXPkVwN7aappld+t4HbKWsMrmaLw0e2iR8RDmW0W3OuVpINzeej4OFZ
NgapRTwFWEFfYSbeop19FaQeQ/cTjmWAnftrCHdQYiRdFSa7IIfOXFFer5lVQ2xk
50qlqRh/BUbUmdHx1IZSdrSA3eBUo/G3NDD4CBniPe8+VScmPgty5feESUyrgU/H
jXbr2CqNXLG/PKXydc6EgilGiPog1gFG2UfOOegtX2gLiD/37w+YSjNHQ+EmT+1M
qoEAWq+aLc717XvsJcABRVs3Imut5HIjYoelwSFV/ZkuivHTCCijtcFytYdzZyOL
VdLAlKHGGv51LSrvBMim9OYJQkyS+PnKnnyfR6lAYB13uNmAT/94m8OpaqvdnBcf
nn6jTLhz0Cwud8k/98UhWZ8XdTKQfiexvDlri/B6W+bxPThn4rJ9Ab5I3kuE/NRB
yLSjc7M+8cTaiMGJyFhwNlZsSZcS/zSGoekmtSzrUTxn0esfwNXSoKtrp+fppeLZ
G1zAwj0f+Ha13VicTyAY1GQWm7bxkdSDTeCCCY2Nuat1Hhp9LyW0mCZCxsl/4fTE
sacC1wqHbOZuM/rmcbT66WSN87KtUxRBtpb2RJlsTO/dfxwjvcadNIYRGXLFqrGw
MJbYBfHRniD46gh0Uq83mbyd3c4PCdkqbPSuAbm1rHTwfPAUpGnuPjYn2UFe404J
UJwTELqGSVJ/kr4iKXvEfeJ0YrQ5ApnDmCugmkmxmujCO9Ou+h5X1PVoi9cMNMuc
mPKCvc+T4XmtQJQSqohDZ/wQa6qO4V4nhNomqDhgEjzoxuFVNjo8qW+87K6l6dRo
GesJsqhwFlsy/OHewffGuU+BiZekBSh9Og09St4E33oU5bRUyuYp2EC5Jnsn99bq
bCa/WSE+uiOrG9HQAXa+7Gtu11Wzvt3NgzEmAsSbZev6IxztZt5HzjU4PU9CjvXy
WRRQv4SILdS1q4QM2vHzJdB0tI5cqNWGLniQoWpHlPOdAo5UVN4RvLim7lz6YyyI
0hcIWEr1o6Qna/FoBlE3utYsZd+vWsMNwEI7B5GElUG0+p2xWCMusp+LgAzYCebT
b/0k9uJp81otawanewszyHnjDUIRzoKz9DiK6IRqeHYOozanXdbjm7sG77huLn7c
7Vw4tBJcD/S9vqSK+/CkeOyjOdmfrYi0H5bIVtbgdKj10dnjE4wi4/RrW0pNFyMW
ec4l8qBeBvjsBjocxsRD//3reZs5lrprT/TQQ6k0iP5GCr3hV/5E+ITOCnoIOedj
1RCXIS+R5fbd1ZjtNeiXfZUpXxgK2dYQbsL2fG+LtoDGtUpDqtIwg/t24zx2aZ+j
2QNLZBctWufxRCoFvyOydKADN/swUeRvV8rN7i5ICCdbmmIMklPiRQH6nCY2JjcW
4UbxThitxnrsoXZXh/u68k+TAeIy/kQPaEyo1yXOZVoisJpLyJwMb2B0z3DsJ2gc
T0+mzKG9wts758Uvv1l2xXHOdcgc0gXxBB4o7W7h8blztHDiybENUu2hqywWFeyO
jo2gg6JTpLm/UG7Z4zyC/5ngOVJU0YGZ8KrhTf8IfRedpzVPhKJmT4RYdJzq91Fj
uIsh3U0/2Gy3Ph+ArRdTTzrx2XRSXcGmukyLyT2YMDRmofXcHM6Sb/JZV26O2bkj
AuOSTnSDSbDAWScRbehiSTCPpavc7djF1+lbVMHYiK1ad9SB8sn+0MmnYngxbdyi
XFMGLIdQ1Wt++XsvwxpJOdnMk6Sb5QSk/eFI/p23D/aQ51EvQXRpQrYJAkfgKXDd
xgKllbsjyJnErum57ejC0SASCxJ/vxznqDpOuP2GbzFkNvJOSPyPbhf51TICeXtH
mG1ULinb8e0XkPv42T0s8rslTY97xA3y7AhN6djODHKEGNRjnJWBgXBp+Gr0ulEt
/n7nYBMRRFyBKJoyckPMCK2i0Fj6zFCtTDoEh6hz+oP7EEnEKOrgkX6C7tj3hmtq
Xrv8+3cc5ye9PcWGiqSO27ra8I7E2OrDs3bkZmBd6jz5uY7yMlBdY0EPI4gQ9Zjq
tpSpGIPBAlBYV8PMiaEcE75v7MHFYWd0uX6QEXOGnLDPK0kyZNgV/oLySwcvoyKN
u867lZNm2Pg9IV42vh4QHwUnaxbYwJ6stcUTiUqe8umRsO/fty6kca9Izibjd14P
sEKgLVxe63pSJVkKc2wYhuTCcbHisyuFEM447PX7+3doH8yIWe0TCgQvKAfiCHNX
HVBf0b9GAjRrdTuYNe7uuvFuxxQMmnyubnfZMuODf4XN28nVgYJGkCIkV2ZtSiOq
vyosb5vclqmux8v1CJ26srJ9pyLK+gRAQ4luy1S+cuOAxgRQCpSVoqmlGbhw0yKX
je3/ns5lDkg3xRGgQXhZT+wZEfk8lyMK4ROqt7vRDpvzrbpMoM2ckLCFn6xcFsck
CFfkwU0e7rFgTD5tfO2QxiOcqKU8QBGL4IeQ1Re0TCG90uifEESPn26GTO7BEgf+
TUcCl5d8YhFUbVipIYzLtQJ9nHZwXaYVXPQD+QypFNpe84ZvbAEvkbsrFUTNy7zS
gMPbb+QJ0JPfaiOCDMGsviq+ukdRiTX/8tOUBRDb8DwlE7Qs6XCV6IU55kDUdBjK
8ZBD05Oicp+aRahliiTmV0U/KxeJwXmyi5WQHal3aamYkrKPR3G6Q6DqXPIEIYyO
sKDXPMntpFxE6dkxQm3AZjWHZsn75AA7664WVb+IQbgO6qmWyznBX0z+50EuRfFH
XOrs+zhAMoI4wF/ET9rmw1B2ph6eF0MHNt4FSd0ajsLq7irtmNXRvaTQxfTEQasM
NoTQZvM5uG4+Pwp3KSUlQmUmj1f/Y8B4Pg5g9NkbHwBacaLHXQ4FtVCKDqVTHvjG
GBZzD5/vx0YS39J3Z1xVMVegJFk8nJ5cpFWssHRh57nJbbIcvwD7/qwLvqr6O1T6
lt+r2NXCJeDa9Eu9AbyULIBFs615H2MK/rwz+qz7GHePLYhNvx+mOPuVRLTuZain
OXGIVmBjNWIM/lU5nph45pz7b4IXc58O/UcIFKSEniznPlUPn1fDT0L1PwqROZ5L
3u9mvpohiOircfamOt5Gh8gcdYVkaRlBYou8jrCarmT8Y1Cn4B5r5T2ykHL8H0+g
ldaJddIncI75NOm28JujnixkdukrMBx5STwHngOxRat81WjJdMvFqwNLpXuPBDAn
mtjgPQ1FtcVOvBaTF/TXmWN0KLJIkUyGmYVB5EOl+sFxXE4B3muIxjTa10+UKxfy
I6Ep+uE0tcWMDNN78m6uEhCJ7P8J1vbuF5w/K3emp1fQ0pdEt+xq8dWq8et6rp7P
z0TM2hg2qnG+CleuMbZ+nvrQYxfavfU7kOG5sq03HJ/cAZqfXKQiqmf8z6/gAKYG
XWiOQ0x9/zqJbQlLrXr1oL4x3pYD/rgh2fgPOWOKJ497nHK2YbQfkRCJ0ecSogEl
8KWNOi6yfgD7e4152EHOo02ckzQC4j5zlv56UZdcmIJXRduwiTL0hu/kwoJpsktU
h+HwrmUi7xr0iSpp+0TZm/x03iPfovWTYy7GDJsMaYHrXHIOEtgx76sjqY9yhHV/
8CKT4cutRJALZhANrUy/sDPDKUNVaTaqHLjayOIJXI2HYaSYwXQLw/Zfzg6tT8sR
8dVbI2V/e0NRc2SMEkX7B+BrNsFcptfbkPtfGG3lakk8utc4y+emAAelOeRSbDET
HDYs0yeptG52Hl/i0O4DJY7tOwv54eZSTz9/JQ8Y4Yybc92cW59YDu7pAVHR8aMz
R5P8fq/UdZaVuSW3D5UV5PfY9i03Om2MTrHr75HRExPPnaIOZfqJI52qqF7KqdRp
kWQADSvg0OpBkq9K5YuS3aKgZ7uEoh0cO7QRkZ7ae9vRcBgfAVd3wmLv+ISgs5K2
8sNeAnbDJVYKm7ZVcDU9wG9C9ku7n3at86V4gCuYuC5UVhIm5pBy70E4Q1YsZzYz
QhPoepr/h2n2mG1OWgabzQxG/MzsrcYEGvHVxuzsBMYPUAaiSZngSOAIpmMZ40lr
BOrXaUFAUqhMRdOmPjwp91j9pfz0BCwfuVsU0jWQA38PqVFbtIAQnGvqa3JMn1B4
FDvzU+GvzPAmUgjIKDyFf2NOPwu5a1cunNFxqHBVgc3sK5LRTALo5jXjzq3KUZux
2B0L3ZEdHe4t6dAvg3+I5yZmoa2GgWU1XoiL5T4j1kQX0fp6yxwF/b3rfre/38z4
CX42++V1yD+WaHO5j7jLa5j3VYZ4deTXkaipnTW65ANtwL6AzOLfIuot2EW00DZf
6fAo6K1R2G1viNp2VcWxuoSo6u8DGP317DzSeKwm/uv5LbI0R26bT+lR0i70L2R6
Y5C8GVkrnaBBI7nx+pTwEihjS3R978Zs2WTDseNyZRk8xF1AbrqjL+ukPgjnIso0
XhTtQCL/K7yceRnqG8hFGk/xsplMupm8dJHLhH8KZ9/mSw/ZaQwVD2JF4ulWPFhz
r1+JxGbvfsQ6BsZI7kjjitCSa0OmqWLPXwimjh/2+6zANAKvuFNL0H3egcezLah2
7ZATtD1IYiSii9xl7nUPl0091iu3ysE5BESVn2p7CwapJjwSRWYSwo/3UVX79AnG
DieQLDWqJO1/Hjf3w3+Ca5t5pvXuV5KajFj5+ZQm2tqsKwZ/aYTLOLHPW8UEWb8S
26YwSJfxxKV15IEL7pN+iQMQKazxPPwT/tmUaXguZPfDQU7UHT8+LyDbfpfMO7GF
wQITKdRnczmuIotpwAJkz70XkoWjY6+z6zCdlQfMpx8J1rtXB3aINSDiUdN2VjqW
MSs36bE7H8jhg6DLYcqTWRrB5L4MuRUxoDKRX3zRUtxemws8oRT+XjZC5iK0vcxf
ZUOhG+pZxkdsh2qblq+2kFI361vZJSHJm0n5kZSTaUkPBZdrK/8Dncw9TRBs/5Zs
9S7BNtl7HqWDLO0/WmxYe0BlBXZI9pyqWMhJvSi6LIb6f6UtCna1Wh1Zyc4gwfAS
LOxCEqLASWAN6havbKFoG2bx6HXqA18FSFIGqIcrCVieMJYowZB3jMQERd8bYnUB
qtw+/Bh0N3o3YLwz0eY76lKTX4sLOSDl2aqD9BH1S+s2H3Q5FJ/66VjgBAlgywTk
/+1Ln4uF+GhbNHS74jtqF3bsniLlf1zSvYl1PImpdh1wI59cuoyClZrSkl70hOgm
db2MODnvx2DSigD+9wvzasjlfRMDpAqcJRiW5sjyOm/4KfYUM1HhYXDEt0ALXRYj
tdCm8hQVP1T8CkwDGfZj6OcVT6hFkGcY2AAk+LK9oxiG5nQpn3JjQPmk+CClxgHL
nTHyoN6SDOeAhf+K/eBpiIc62TCAq1quRm47h08jabm9SxzOwGy/AAuVudrQq1np
wpliSJzEnXHZJnypVEXiCG345msS/aWWt6GKbXnbQ+Pqoa7BPukZOxA/nsU0Ha+l
oGj+gBM0Yx8M+Nc0LD3tPBn1RsDkpaqYnhAwonT7wjh27iTWIiZnmJQey9qDIJ7G
7v1W5kIyyQr+9unoSOx4xOT4JmVg7HBqTQU1FoLCCyB+/aWBdwKYw5Zh4SWJOY1k
3PWrXpVOo2UdqtLknYF0Ptl89s1P/pHAYtgjtkslbnCO1ZGi8aFEiZynxhg/PQP8
+CxtuAgRxQqoIm/KI1b3QDbHJI3qfqHoE0ELWYptfLCwiekvGp2gbJuH1g71Oab6
3D7fHZTSPxu8RwPX9OtuA7Ed60gFhKtTZWqa7PXC6MMZJtmlWup5kC79lkY2oPgG
deUAFPbZgEtNKu+lf4s/TxpqWkFMCg7z9cLMPNfwhdCm9Y48YlOrPkJP8ko7SqWb
pZ0WOBWf1buYbfgF3ERJBqnSOKoC2fx8W/nHZDgvbkIVS1R23tiou2xIMWMeG1kh
c94HYAma6y94mC/L5OXFGOgBN0H1//wGGydJg6/cNOGFxon0J5fNvF1fDI6yc76c
7f9BrPFwfw1I7I0mHalsZJDEA8OnNzj5+Kq3cf/SBvw20nJ40G2avMYkKxQDyPKn
/LfjjNu2qCW3Zi6G+qHg56bqAvxcmp0UcZCznpW6qFj2qzTX6ySUNPON53xq+m4E
Vl5KtPY8rwdh/YlTlSyoMpB2iz/6oB2lwCG07itlXxRByAyty7Dt+RUj56Ocsonz
sQCNPGrqWvdCF68dkkAmoD0P8a98pxsWeIenDprbY4yr1yIApGociysgW1MDPn6G
YYaSL0QZfmDAbEVwVxqaalRTQnhuM+Fiub7LWBpOliDTia5xcIwc1xbKmaCbrJjG
wM7ab3ZMPTaPFrAnE+0V3YoNiQKyeJLMmbwoBGnJTN+2JQ6iAe/i2R9Kh798rJv7
pDEqnX84IBUiTmS/F2edw308emjw+pKlBL3a0o9uqtBeOcZg3rTtD4AFZ1JXYGdQ
bvNxNrSTGbTR9rAPSpF0QJANKraR9VUY0xrRXXcfpODzF6YFkp/dfSalgbWf5BL3
m5fovzWwQrzya4BpO/32X4ZEeFbtnDOPxwDRjBf7qdzl31EsB+77aOJM8Arby54E
/++gMkMYnaeIV+q5frE03C9QKuDN+9Cq2h45dsgDM1DjlO6E6e7oRXrmnn0Ysf+A
0A1JNg+tCdq5MCSUSuMLI/ELqMxZBIfK6ORM1SkyuLdAIJqg5abINiAQYQzmTSy3
nFapzMZlXrMYD+IwKlmKlPR2Qf8/JTn/V59OSVOHY1v5PPjLJ8mzuduGAeeEasnt
7KZm5bj4zaOI3M8vycOCSl+KTLD100d3ewL8DVxbDBisTEsMbvxarOQfWdATu5Rg
K45ajklhdy+3SqO2cErO6l6ay3H92HfKZy3WkKzXzQ0lmyxNy2bueEKWrz4cBde8
OnLzmVQylMoPrjVLdAADKihm1UjqywzUbPh4egtGkzzHgY77xkYuI6TWBGex+Pjc
4e01+Uvil2+lg0R5blzg9Ks0q2ol41Hg3w6OGn0Ekr2YFeA736q28tWGB0/jBX4U
wMLnI9FuojojIrdJKz5CSI+UOoJwYvvqFKO/FynYu/itMMYIA1cmoJwZP/om0RKg
HzqNg6bWbf/yZcn4FL0HORUuFsVYWb1CmGjbd79f/RE06gekop/oUK3+8vyOQpfj
gcR1iYRaitkuCpTpsSerVIBaMqnzm2r38zZMy3gZ52sjR8SUc1B31fWNaiYlYLH/
+9586BwFM6sAbDWU5nmGLUsKRxqRy6i1A+NGXlYj4YFLld500gj2RbiIkeB9Izw9
q/iNOLmpyUYD70Yr31Fny/ts6CVKl+s8S/9QnOZpGMseYuitsSo2G0wEWHrBt2Bq
EUsLxacvsNCF80SfEKDEXy8W4StCxcw3PxehnLgHT7aYaJGMoY8CnKuCswUMtGfs
T5UHpO5VR8fbvU9Jarqhdud5jeuNgMeBK9lmIICOS6uc8lr4C5io2RB1qIuLoxNJ
qkRx2fJ+BgB9xJxp4R/kLsDyqXeyX0w7U0CsqshTx+sE4GXiQiqhVpc8EJURs7K0
I8OdJbnnfaF94CaNJ50wVzPgWOAt4iuAfNmcXWRhqF5gE29OMLx+/nkAPUzx5NGK
XcVCOkhO3gtGaNG8f5jJXtZQ/Q+iFXRiJdCncU679eWPEE2ZSyqjZKYp5xLCeomC
N5z8Tsf93ozxh1lb95DUB6/vrDvQqyiaxKui12cv4bfIeyjzhnsqDOHoV0MZXxbp
p3UCT/ElIstmsze/nJwdXGbZlSxOJYVGkK7r2p8Hu7z22uBAFRuNRqNeRJtOMEDg
YzP0+m2HvR5UE8XSQUseSvRq1FLDsN1S+J1kK85fH8WhyOz3Odvzg/6hqxT5paih
3nmfZYtIdrqYBtDTziRti3KvZGasdd2NYiVDzaiyVL8d2WuBQuBJ7I6tPK7t707k
qh0HDTu1ECvtAbWmtdREKXz5O9OYPOHlh1/Msvdfj8ogaZWfrPCjFku4Vx7SqJ2/
fQCyzBkhtB7lStcu7oBQCpbJsG6P3u/MoBMK1Hbk/HrYonFauytVNTLP3/1eYH8H
FvCK0P8RpdHiWS8tQnfqa9LJSDy8GTRv7Vcdaqtf/H7TWHnPOnC6q4RFpsFIyQjz
csPK9pbK8ByFTQFx0kCAKQX/4Y4ZK8IvBxS/TPeObxYO9btGAZ/tRHbJJvmiuIVI
hvlo9QjSEECFah4aHZqsn2PBSsZKd3D8nhjdtmj31Q5t1z4s+IIfmBi32SL+0lad
F7c+3YN/05RaFcsFdJsedXs7Bkl7kChQmyu5jZC/WgHVGTjFjNAm1j+uJuPa9iP+
0DYqkf/aMJDSIjNzOpSr55orB7NEm9fu36BYuyRc9XLnL5uUJb+bkWxR2M+Yts8N
j73p3b6bUQP3/mcmv5kgcP/qBpcZ1WpMWa5hNqcjbZkaS7Yg0kQZhA1FLoYCUD8F
zs01ogIyacr4yF4yaMTb6Oage+xNkaK9mkZLZj32pKvQH2txVH/j9RoBAagKKx0n
lSRkOLcqnDBtLq9tOSoArwp1gPDv6Idh4TR+umckj9wsLtsbLaUV5k4z/Rqm1YpU
qO9pUZ2BZCWgQ9IiOeui1jNdeisdyyf2veNfAVeFG6x3Mjvh2OF6u/9Rs6oBewo5
JCSop6Stsi4sIEE6SKB4MB8kOECXjXy1k5IbRQuiE3hyGshQl5Hc+/r4TYh+acIe
ui/eBoUxnBmjn4BJBIKlHYcFYna7YlWZbXKPjgfgNFPPy8IAjP576b8Df6XF6y+6
DW60Bu9SwOWhymDxVE0qN1Wp2j1eQseC5ezB800hqCGNC6AeBykpiywcWxR0Ajy7
rtUBqxBXcYCHOukRg/2D7f9uIW4HIEMhrCoctVUOaL9T29G6we//IUvZ8I/5A/HC
AD/wh2sNVQfY9DRvuSrTclVMJ/iYmn67G4p72T3Ok2K/xICg+E0P2h5389AGedSQ
IhzMQ7KzdxKQ8Siczhw8ExgTWfEUqGplceO+CemfOwSHw/NuNPthPUr4sHIVlEwp
QWwziu7dSb2NgHFXkNVp2d4PvaMRFN6NA4tpEkHM5vflqbd0B6Gy2yxHNJLryqEQ
4lJuI9Ps91Kp5NeZVIDUO7Vpvaj0EyTdWCR34SLfeKjimujEUN4+dEAdL8sDndyv
oPWu/b+iorZWT4ocIJrE+h65qjiBURG8XUiAms3OLWqFvN/3et5sWyBYhQJkyQTZ
uxDZU7dnaWPSjfwttGtdvDheVp+RHFlrvKAilgie0C93IPvbHpm3M9QZsAV8BPOn
r8nqM54yFfTwvfUUpmurHyB5+UT0MWLf72idxnKXZGL2a0P2t4Ivz0U9QWJIkcxi
DMaVRwXPgrAJbiqw/VCgf59cu/rw7S/KV9MLOU+EcFnvSx5vPUD1oHnQOVC42iRD
ozb2K2SljOI0Pa2FAXslWpzPvvpFJLHf3Z38OQfuMQ+rJcksJCkoN15XvW+rjxT/
zKIfq6OoFyl1uamp4BW1XM/pA5bw4pNz4gnw8S6jui8GzJekGkxAMa6Fv6r8LtYt
MAGZQ7VpNT5vNg0l3cFpytyJthpYoekUplJjD76bpyAiCOa3rWa5L4DZOn8j2S2j
1KAwePJjZ50LwW6exNlrswQ7Ed/ngfD6vhfFjPBP7wQf/mUYVMuNGZclKW+pz+PX
QO45A3sErQtinHoQjWT8Ds3yLE6w3KMBgqdN9pazucgWy+4WBEJf9ssEJQ/SDp0a
HOK78ON2ppruVBxtes8ghoqJGWcF9jkJbjWGPtHMXrcor+u7xUOPQjWZC5nBXO2O
m2RhbjY7f32OOw+6FAgCo9zkemfaa/ED1cVcv126/Hn2klKxkbI0fjUptAVP3IYK
9o+tw3D81Y25Z7HkEaKeiKx6EnOOiw2C/shh8hh97lPoioZGW7wfqwQf/98laLJI
hiWrpJN6huE2ojYp0Ogm4DfpsjwPZR7SjWSO8AHcmeVbSlzfRdxjLhLcgggTbgF+
9HhlzS0eMGhjWVCsYODJ2/eQXHdqsaR0YGXwpHN5KAu/5Ji3Suh+6KQXttwIrcSW
naenDdRochrJmhWxpBF3XJZxrE+/4ixNZbX69LstAmtgyFhqDrpmoc0me0hVpnOw
AAC5bQN9sptIvMgz37o+ToUXJ+yWkOyrZ17ipsJ4YLR1or+6PS73+1zv8Td1gnB5
O2AnBjzgwfs6vhWR2uO7xgSaP6tTxbkq/IKP0p5nHbSGVQbcNNEMEuHSBD77ET4G
ipAYjqPTK4igK1mQjqppE1796ivqIzukGo5+LAfvkUhBmBAKd7/41LKAU+HFiUtV
ZZoCaufIpKVG/8qcXvpj6/ndr56tWIogvQHzrPXeUEV/SXTCdjy0K3rURonkywRl
p2HqR+2Lv1N0SoleGMME9TL6V/YViF6qR2jK8inqXpfcA7sYaEL5nfyr/v7otTrj
jl32tf1efnQmGxVglfny8UMhIE2AkyeWm64WYZNL/IgwcDPQjHHNd60sXOxYVcWo
q7gV7Ksj6yPdM/qU1NBi4acT28pHh3jRbIRcLVCvNIlOxQySP6vzA40YdfXHQNSS
57NyoznatbmHYUwvimkKc035YeksKuUY2JHZA0xGiU0XaJB3Hz8sloBcjmYkKe9C
p0bbe3uqycWC1BpwgPO+rkDrs5PE92D9UQRrMTkgo3K+9rdB/vJWs0Zrym1U4YBt
i6vLYadVodObmyZydC3n43LBhmnjZ80dNQ65eIh2DAouFl6ch+a5QUip+4OAkdzP
B3EHBnD3mOUM6IPopef32SWQnyo3tYqXLVQKbYZL05nLsCRN/uUwznxpnS7sym12
MVNGV1HBegvW18YrnqurSkjkzLmJljKjRbf5PCdQIFA1vwX0yLzRSpqEndyruT2e
lIRvzC9bTUXyZak+kMjGzgum1gqcpLbfN0aTuVvpkf53BAe8E/Q++V5aHzddnagm
CfNQB0U+a0XA/Tz2SS76XTpwMGr584o8ApASLgXrqCX86+Y+SoxR/fk/JreEcmMH
JZ3paDny+AE656dpKfx4ws24iu44/4+UHVrw3MPNnREPk707Mf9HwqbnFV9PoJgJ
QhbpmEXqFSX8AZ1+pDuVK+WxGt+aq9yGOSfo0IY059912h8uOeNH9DU4w0A+Jltx
iqB8Dn1EOxNHrR13C95AG/qiIizy++tjtLbo7WNqnN+lVc8Pb2jAqzusyoDOgieK
WM3asRdA6qUzQLMeUmPWmbEkMhBdB64NnIvbmVA3ZtNb/lcIbuJmsdP+D0JiP/l1
a0N4pVbti+fRBhIz019U7mfcWJKrUY56vbt6cm6+LHWq+Gi5riAQ0NUESFyWTfkf
REQQEr13sBXEmbqGRuoWgY6kHL9Eh0fVilt9iv7XogGiWLuwcvn01ErK7zESYQi8
cl8Axs4KCfVLG9spzM+argslQsWdfIheCEVqOKNzlpzQHUxy052tX3MPX8F+rNJs
MNRY28EwtaVzXZPycdk0f3cig3wQoTSS4jyVBQzU0383pazDTb0jUpi5zc056Yym
YiIIBMy+6LJKLG5I+X8wO06QQXDAW7Dvcg5FciOgLp+40pbFzUGO/7Ndnf+XXeQZ
Gh77AQeo9ZDdURYyV2uZtL+UFDV404W0tVLYQDHV1ci7cWJSV2BgY7X1hnRxtjbs
tGfo39hweFIyBs8XCAOC9A6fB23U9PkJIHuXO395chiNLiA6FOnG7j1DqCkG6R/+
OGi0HPU6LdIBEJsncm+URB9xPn8lWxOcvrI+3+j+meP8KgDbVhUfKzrWgwwDimQ3
5W35bW8HAIevRtAFG3gYZhBlJL3v7HVnDeBFnUd925rOMIyurwa3KS56uVR61OGG
MspR0vEX8G9k3Qn7sII8nt8yOMwZpf95kTDNppyltPCM1uV1Of8rff/qgV6Wa4zY
55Ov3u0cZxlTjFpee3B0EcK0RG4W+zzBNIZ5auK3wz/t3CayI9lmJdsqEMCmCedY
CAADL7WO/rNgwVnTBUG22bFuMWFDB2DPWkOQ85Yh7Z42bqxSC07zcNlG3xpTEcGX
QDInRhr5DE84F59Z0BtGFw7F2AkGfincQPxv298S7kJdgYODAoOKLvwJRZYBF+Td
dxb/VVVcwUUvcfCljcRVOdYsj1Y1J1wOfXkKPFaZEyDAO7ma2g375tY36oLt1aUP
BEdp1ZC1s2DJEv9pG+wgpo7bpJ1jBox7Zz2K+9F7Wd+7D7ycoay7jWJgBL2tYSpM
DbQO2AuvxlfwVJTxxQ+FhU6ZgUBHnP8WqbWZqIRBRiEz1SF28uoGAtPEHfgvyjBm
ggEfeJ1u02TBx89lcetYVwqEWMsWRGS6d6vx6tf1gsOr9+bH2zk0J8qQcoQI9zyg
8qzkp7AGnrOynErM/3tX2nCIho6ipXV6gF+obr+ujnRMo+TZDhCZwO5Agx6orFrE
wxyplFNqAzsY/qgAJH9cvoF00pH986OcE0IcPSfqyV6oBDf8r6rfYzcXq4+zG36E
06UhbTKs7SxqpDf9T0y749F2w1EQw6aCF5egXaEQwTX7oBCiPl+vg+OIFm1C5h6v
HwWI8m+DQZksEnss4IYTYq64EQkp9yQEZcQ00KbtD5tR5R5tkLqQ6FZrXRJoC8el
OqgecCNKXVKSlc3ejNNsbPPg0OpMNR36um+vJTGctPCXMWPapvVR3n5uT687AQ2t
K9ggEwkG58Z9+V8idjIGy3FBmAMoiPp37DgrW2hg3+ehLvKLFH2skTGl+zdIgNrI
mONYLWhr4fvS6ziOsIlkAnO8ATGYfNP4a9hOp/pLwxrs9AdmjBu65hszogkGKHfR
NMvowqJPtH3d7YwNmdm2InqVZO1kgA0oTcKGJRvCTGPzskcGLfOZlrbyFifSHBBe
zR5MLJW/cvDL0/IKI+g2977Gx85ikCMonYWo0fS/bsfmgzswSpklY5mZCP6sK+//
rsQDGJbQMoxFI9La2XOQBJkzfhTQxZ4blqVH1O0ncuEBnXpx++wt2ns47eKP70q0
JGYvgaCGU2ymbq5XVCbtIrzUS2xg8mnR7qwdUdrBoyG3rIoQALZ5d6x6ShW413uL
sJhL81QZzdxbCwSGKsybl/pCoYElo8NvXR2RAnyKNrhbuxFFZlSaqPAYMC4riD26
lShW0lBD47V+bYSXOorFKrogD/a9GLO434/2IIQgUKP+2540CQln6f7kP5zS1dsF
WJQxKirzF7jv775w1qNyPw5byC3xBzwmS1Z8gPONT8md6LRo5v9jBahtijgZEy2M
NYlPTDCLQMtWwhWr1jrpIaNWbhJ3YoKfio4feXu6EvrcSncrc1w1FVtd+TXS9R/X
zObT+RqigB9gl5VDglso+G/0hxpu64uVPGKRY+oIn5kNMt1HlgiCaRfHYxCzKj+P
F3z5IArAYZ465dHUnDf+Ym+PwUMoP0fDU9zLs1rzluxd3pdeXotoK31QpbfZeQPB
04MW2KaSGssAYhVQ8Lfskhh3bjcOX/gxX1chiubMMNHSQXzLy4Bl9UnHnaRxaIlu
83/KMU+K3Lt60DM0i5dtMUe5e+yWvBrVrk/hNmj2YdqvcAuLgjSfLTMVR+jYazmh
aJtPI8n8s3uNnVd5i+FTLO1Ivbug2rJfnYinCnJbcbZUVFUDZ876y2OU8Qw+O1w2
QAO37uZ4xOCeDXV6ykBeoFeXAThWbjWSy7cvWj82nB1uJmWbM9jBIAlaSAtzw3HZ
xVJgxYOFOSx20/cYdV3YgayZGlN9HlVhoSQXO74rGgVA6mw8ECgPUBpVNlDh1TNr
87E52T1FE6Ye/IGaD9gG0IohJzWYiJEHzhK6wCZrrizOk01p9WX6jGRQgqMGscE5
JLO6WoK4I8pKfb1yq29aFm5bKv8576NQBaG4EwgYyZcpidzBulMa6fTh4njIZhFx
oeHSXSa484JJxMTodq9Q53HagOiqOBR9X07ykVglg0HRgKubCsPykfhD6CGn8j7o
Jol8e88gOkB4wwPwL7zx4lBYmIl5FZQtoFCgORcra2Lf4ZwxXgjpOQ4m/TMVfLwv
1Th8Qj5jeoCF8+cEvbgFebs2vqNWoyWbl26ZgeCgvTOc0A449rLx1UQ4lpgXm6iS
QLq6TYydO4iNIkeOKcqvNR8FvY4C3mHZJwS607S4FigWt6Xr7SRsHroEsOmArRc0
CRfjIA5wSBJ4cUljSjIamtxkuR+Opc5f5lg7rbPj5oueoPhZ5grI4vQQzqL/GmMV
mtLFSgwHhN1A3Mj+rShDg1NaXOvY/EMB9xdeYSX8yC4Yk3Gw+jbA2K7UfRek1IBr
wsRxeSerUjgxEIOVSzgXcP5Yc/HZ6mkLZajiUYOotazScmsY5h/+KHF0SKUk70Wp
zQBwE12W8uORP6pFYZgrkKA3g5qpQ4Vxs5uGay173xI7ElD8PmaDg9NX0Cb+z7Jq
Fgdq2f8sIya1RHU8lFPeovTZNsnbst/u9ijLmuZYqO2UJouv8LfHZsAZhDg5ySJH
rBRAtL6HRM3CTH+rRRkoqMeeyDzPfckY0SY6FZ1kvWG4FAWUx5gtl/xMJI/nK7Mz
gOq8Joxhy8nDycM1rVC0K6sjKQ+4Dulo2tGFkBtsYeSHpS445guN4KcsdlkA93lR
wwG5ozZmw2z674JtCL/9i8Dnz8d26TZ4iGFx8ytvmdfd3ArbhwlO4fuHKpLG3BS9
aHCD32HYjYW2/zjFDf/JLwYfOj7+8CwL5ohRofSIwemNxS76Ce4M4el+AtwLothC
mDxfrcjrXKSv938T5p8RkIa8dxxARUuMjMmJsQyvvjf6yFsltYR6ab0kpzAOMJtH
lslLszP3TzX6Fy5GpEahNW3Ldeym+LwoC9ZM0ap1yAOXMi2L9Y59p2ENyVJOrjLf
A/e89fbAdOiLX+Ftv2xv+/ipfGm9j0Bfvt2oQKT8Nuiy0ugftr2t/H+y2obUGz+P
Xtn9VU+MU4ZxFBUIObvc5o4kD6P4Dg+tEnMt6s8Gz7V58RNu4O4YDnWXKq9EMk5C
1DEEiVHlZFUePyIe510dTEztFJnajFc5QPCAbkquCxXpNYNOYaXsE/BKMLPM4BWj
rwLQkps9RVl1ao8qVGy9qP7B2ugbTocWQD2MurwsDkgprXaPqMh1FdE7gyDns14B
NsOkekOgSySsq6U3B3gEcJEwarANBFUEebQBJm4umSdYYF/i2QzJ1hNH9RbBOZIz
lhPEDgN0Vx03iGO4EpRPfMKj4zbPg2X8shVJEQg3pG9MmEie+F3Uyi6ySb5rO6sd
Hf2Q4ay/hiNzaDsrheNeZgD1LAt5yMbOT71aiqG5krZScK7Zwx5xwIz/pkXv1+ej
APvNFCEvaM/z3qsDIUuJkj4sO7+PvcH7IvD2wZFw3/Je444rlbFZ2Jm4PELygzIh
AfHL1CVcLH5+WGcaLfsGAuaPZ4sqvLQQ94SXyJuhLsoWRNa6Q3VBVkAnUZGg40oN
2tpda6THyzxr0BDK2oujmf9hQS01qxyrwPlP1IU2n/pCoHf+kQMLm0MgBpx+maDi
sH5FVcDrzcct3p6Nuuq3/f5koONvjozFes5jW+Ovw7/Tk9dEudWkmNsf0QnvOAeC
8fnWGZW5ZIVjCmlW5lNa6A1GepRRQAXpF1PykkA4RubVwlKLAP988xKXn0gQMftd
6G94rkh6/Dd/6PUZmT3NsgxeH3AZ1LCanorsBU2N2qtQwd+hf/Chupv7+zLh3TMM
abG5neCXgUiuA88LRa1IMFDAkyZxj2nXhaPB/AOUD4khBOwlbdfcrAMbaNTMSqVe
UonB1c9oQe2wwFUbg50WMQdjTUuwNBQvd3z6excqUaswYLjpbS7KfSbb/2J2+13L
ITVPeixt8FrnacRVGw9gWZa9+fGdtn14xnmVAtEwZ4e80bSx58JrWfYI08dJw50P
hV0W0+ZqpjS6pD69P3QOs+xsqyc2WHhJRQEhKkBOZJjPGij69UESHMO4iLD1ZMGg
GvuJnq46ELl6PlXts8cSYc/DuWlS8Eo8hjBjaOAyuvOZfHduH/JkEtZmqAyU6GEG
BwyZyJv5cXznLaFEpsjaS0m7Bqurf1Rq8Gf2Thd/+DtSOjsyqYY3iCZAJIBQPjQs
UhffDIuoFLii5e+A5TWU0blQqa+5B7bz3TQhJUgswBWTEMDyZ7AYvB193uZuImYj
vM7QLv/8lgTLPPWq8gCemDBK7boA8/gEXdMqGbyC0Z4BuzwLL0VHSIOTGpFoHyuk
mVle0ZmCgILSvRnnn+PnsE0Jb9nQh/1/KXH5+zBqosQpKoLpyllvcTxQ8doJoNmD
QPYsjqh7zItxpM3MWmQOJnRL5sQ5++Z5VcEp3/deMSYiLsnfImvMTHgzETsAVbFJ
71BFXI9PeQgbS+67KBhOYL7x3BSlZ31rC+Zv20LWfb85/HeHZBRaVK0Zjt2ABDr9
QhIy7wNumVt6fORqEJMcdnXJlUX3o7/Cii9Mg4DED1LQttfr9eHYZnIPcz5X3kCE
yf0/sBwfg9rlFceiAWazmdOzQdUw3yq2cwFQXRAwlk9M+DP2FEmn3NSHVzfSECCl
dLxuzDrzKsYhJMrtRqePi70sTieCVkmf5kKy/HZ3pQsoOYovQkmKRZOJmyp1RAkl
VjkcoEbc6xyaZ42moUE9bXL2JIUj+W3C06bIrnWB64VsaB1Gl7ypF/AVut/yIRbf
RklYzcKmtJkN7RlDCmoxRh0tfFbhGlv42LSioyA8gcmx6DocRDdioigYlbV55zXX
GYPGKCaAnW7CSr0nqDRZvcpGtNhvFbmXWRt0keA5qPtmSfqp7tP9bCD+OKirJo9q
aAjFr+dCTNFSm+MlipI9XMG0RzdQYKuJoCc0onjpIcXOvPfe0wLM+Nbq/lqpZcN6
yhklVdFUe/MlL83+hYmdENi7oE8V8USEkk5ZoKamZ/qcPsX4HoWkHhSUabajMF4c
ABhCaapD2c0MOy3jCU70w7zL/0kKcx8LJj3GedBnk24AkJsaNes3wt/gHQl0cz3g
ukVLm4N6I1SNIfdUdqV+hjceZ4U6sDmgPMWaLfT3tK8W+StubNOWwm4/R0L46vNP
muIa2plVpf/iNXhu96UBxBH4iVsSKyXx/Z4ihZHXhugJHjZjKDQKmCqRfnGN4zWZ
S1lh6N1NFKR20l9QcC3Ur6P1z1Pgnbt6P5cF3IKOhuOAusFovW2IBNssH2Xd8/VN
VdSfN1gpjJXHU5SbxWTOnyZnEBUlt8vFDnZRQQv4Ywk9gPEL/nPfwUMPh4TwExGD
mGq1xYjTVAzm7F17xlT0aFdJ0DLHzKQysTNcId/ddewX6v1/jz/sMO5g3T4253Y8
TJ3umsB865Uc9UpRaq9M+cdU3acGK/gkmVN07ZBtYRovsrOXC+/UTMDF769n6uRd
nE0CDxvPdC6s1rZPB7FcgWzC9y0qFbWSQo26LEchnBO7Z/cEtQ5Ba45vWrmMZ7cS
IHLLxD3jTi2vGTez5dJvzc030DkBIqozLQXnV9VZ5akV7jvZYn7kYDNzf8w8Omf+
+8MW/W5OUt2Y6Cu+qys+1WNyoSu00Eg2c7UFXNElhz7VgdjLEti5c4tJZcaLxSwx
IzcYTm0WmGaDMm39bbvCMXuVKxT4nFa90cC5djKaiqLtcfYNMa7eCfyyKRBzZGOn
kWsoPukTY0SxGT9OKzUJUOxDd3fw/z+PRx6SyxqvEwV9GSeMxYUHlhdiJz5x5vME
79muoBHcoVw1l5rA0/kaVqO+2/2z7nc0WrNyMGQ0199rtTpgMTawGWjqhh/5Ir1n
EcLSnnyGmDp/pvLPjRscPK9C7B9hW7TEcV1pqywtqRzqD6DsFJTZXF0TFnVNxvAq
6zqh+vMrDRexA7w6M3cQ74IAIreXjlffByrI00sxpjaLugiFZ0325hdvU6YO/tcN
+3xgWMrYCm68I34HKe5iJRc2siToJ3JC70sLHtQ6Y2R+j7wGD3q4QZa3TpZqG4Ph
g697f/qhubMniJDCJIjbm/flBt5M0OmyfZxxgqBGXTxABvng/NOHs3SBrky6djUj
MXVU9OqZZGMYBtjo1vcIHRL8crGrFp+Maias91f7inBZH4LbA5GAwSeMxcvuZ9VV
mbmgnT97JUjHXYASnX6r9Ri6jydNI+urONfv+uBogc7EZqQyLPt22wArISgasTwB
O04MpeNgMWro9L7ABXE6BOnFedrotKh/6unFs8iSd85z/6F9H8JW4djCGCDMyzuo
SKyPfOVsURFebDZx7C4dbnzGGGlrcEjopB2ahEndM4QS9g8IXAP+UvM0sdOaweBL
C7GCnq74qPRoZcWeeRDL0MV1sHLELFhfM0D1nlGValqQ1OEAFf6qbW2rzxwSmlAv
oJr79pGVpwxgfMNly3Dpa3TI49kxjg4i37dlaIDI7yw8KRKe1WP8sTxzVKf58+Vg
Ubhu7VcS3b0O3a/LUprd/1+YJgtRY9lyabdl5xi1rSLGRJxbEe/gyzxwt2mHtDmW
ixWdng09VrhRCgS+PICfhXWdTw8ng0IAdaRusAIkei5LV3rfO0+tbX0uXOIaJvnj
oXRIFrEQUbOMny7BWMrtPRaPtKmOdfCcEzuJY3MksVrA42widC3gt6pTR/359bc+
oU1d5xeD4biLrbAfxIhgrJ6vX52sb0om+gJcA3Kg10OZIcHS9DKAv1Csw1NaMqlV
9EG7KQvowIc6VFOR5bJTc/0sPBTEu2L+DXRuse20I3T4glOBZPO+uQFrpCahcOyJ
gCQx8LjCJqEaX/mPqjKk00NQsUdoLJBO/Gb8e14UH2KXJZyU9W+4NULHW+RT1isq
Ba+RO1jwe8ph7LhkDpaIub4+DVhhZFjsp2jYS1UWTQs2RMZNDcvrqebGXDrvqoOr
3fKa7tFJalqaZ/mRu80adsTEkwfw/CdMBcUgkXQ/1R1CAmbelj0w+8eYpC00pdhC
otsVvRg2AdCLDZcRmuybKgSq4xfErdw+dOoyImpJssfuMrU+wVxHiiZeKASXgq7N
DsSzT2ikfruJjAfhbz6DJnuu7yyfNBHeEigfjuE5bmfmGaHrKcaBt4ks5a7uAsYx
iRTmGe6XCITLMXp2kiOHwtPnK24mLhnnAFmD90E3ZHf9szl8kbgrhZngnSu3rd3o
bCRQVsyHUxcTrCzGfKFfzbm+QA0HDCMb/ccihHjPSNTTE5JM00I2JctDJ0YQaoEs
CNZawtH+vlIHvnR7vshSuT8xlFn/gzF3fbUukDik9aSUxH99MD6fuBeTOm5CZRw2
KTsrPeYtgcLjq47QemAtzihmWJMzmQCNxyNeWZEzmXah7kl2xHq3xWKjl21W3dPi
bDzIowyGGlLjQ6HHcJhU/QI2JMXSI0QFFkqPDjoAywlZEA9ro9FxwST3oZYr/lHy
vxj2UR56VX2q0UR1ZwXlmHJL8YULrt4o754mS0bzuKLvcj8mrpeTZatR3DUYKCEr
g8zZmnMIn4r/DNtlpa6tHkUboqRMbdX+o4TZ5C8AtRcbKDhJV5tC4LK2DbKyjRj6
SKunnVP+NMUVTJBPoSrUyGvuIwOkDCqetV05B1UqTkUlkWwBsSZbO1FljcGuotIa
qR0Qhdg7wbOzIOwBYvtDa+VDWHV/ak3GF0Zecf3d0/b1LrY52MBw5nTGigtWybuu
CRdpfSTe7/WdgdfkbgEqVjaxigTZIGYG0ycMaUTgQEECcltdauNzoEqFtAwzZcfC
6NwDXBupuJebpIZcjDF6ssdtyf8NosVA2wqLF8kpAwH44GctmjbeFAYjnrCPJKWa
BmhwvWKX6zQzaK9Pzjxpny012XFnWOiDeHwdNGYqn5IViOKjIZ6ovAp1KRPqFeun
k7Fq/yIGKYNvUpd9+K1gMixU7Qmb3Air+L8R7NtZs5fl+5hRwpPA44OGHzxkiON0
2K3BwuA6pk5cOWwCbzpRxLt++u+aMkZNT3zI/8szuO4Fnbk5vJKKPCjEtDWJ2Hze
so4uxj/ffTadDtimzYrbNuT3cgD2b8XCxYHnC4iSNCluhbN3mb2w75pMkzhGqles
KyrvJ6uU3wSCUTSTAfoFiAaIJUDhHLlSyriV7zdxsj/EOAbUDT5DlRjy1L7qPvFD
gWiRJ3Zzfeqovrx9uutIUt40VXCRpfeRu8/krQbecDqZjNfQnvAjBoXXFBBKqUtu
22cjr4OPFPvemQ2ykuFy/b6iWXVfBzFfKiC6N2jKVD2GPPis3QbYh+gW9bWep49k
GXlbv/UNmOScuW6VPTTkEVZmSMhJn1QbDRaj8r9lWPD0GUSbgEJyYmnsKvxD+7AI
nXmnLSDRNT+dqDVU4BnHJEq/KjUjNB1hlX1fuDtuPZ5HTy+imP6LAcwAOx7DSTtP
v+em5aWG8DaeDLVEBiX3pTAAGWKOHvlOnICCOZSNFaf6jejMSoZD1MG+hUs8g4mr
vO+co3Yzk3TAwNSlU+rgwjtPIta5ajCfbIq7WFs9NLek9FCuf6frJnpjvHEFRrfO
9UNI9HPH/Ka+fajv4HSIpTM07pOdFmKXUvXLMbm1yyfTjv40A5BNHZQmj4QhxniS
9NpjCtiHJwHpcHWy6j+7VvHoXueee8qyjT/fA9vwQjIWmtJQnAovwSEPUfj5LZ3z
w3r50lu9P1xwLopWRVcR/Gk6bUbtI4KxyygQ1wBuXJjvyYm0aIPn3fKNejaj5T5/
aF8FNcRDJc5GsEDLNXCF7GCBSQU/Yu+wdBC/wbHpkMJXgeHjaFch1wlpkY9zP9e8
Ca3tyjVSzL0cVB8m/sRdYBEYTcPXBqG8+pkq14dns9kt5SDJCM/l47i+vPMih0YJ
cbS/aanQPfEOCvlvME845H/Ypr0LyzISbGThn1UwpGc6Q6JIiiLEvtQJN3buycxa
5LsLOzjUL7W7DKL002pTfNqKjsnLWOwi+fNiLXMRmu0ecDRAsCnjzUjQ7sFl47LI
jUn8Q4ytSo8/fBzDTyp8go+hCMlrb33ThU9Q2Di6H5jCmfXWYLQRMfzEmz4kqvj0
xGLu5EL2cdlKLUNbFTDRaX1MaF7W8JuWnQJMJEDG6RUZ2yoG7x85U4Sp7ypeiAxH
hHml+f1FfBKNV9p/JMJjeppAp+ET1S0zu4A9/fG9OGy25wBsDIlQhhCkbPuwpaN6
pcMzATWfUNZPvOH+AaMJVVEHebyyFYHR3o2O1FDYMyAd8CgOimkn4dBYrzUYfiTm
KIIO0UMW3A7mDEEAmwDcqottXPbJoh7b/rlcRuQiEyywLL4kCh5nmgp5g5H1a5Ha
vmvsePtEWIQNSIkJFoc9nKZTKszBtsZy5gGxjxGQ3p1p0cm+eQzGIEEoYW8v4rP/
r/grJfFH8FaSlHnbJqkf/u5NFww+0YW2i7eSIBG34JeeJy7C8z5FOkxfh4ZE32qM
8ygnkm+Xy9kOxNLI2KSORJgPdWgJjl59IZIZZZm+8RkTy+H+zlDJH10wsh+tiZ4P
HT0t75JvUUEhBZ8jUQ/9VeCI/l2LhZcJbPLtU3QX3d7ZZvrGO+qysDZgZvtwqQ1P
FK81lvuKwwBkOOkFTYhbWv7e+yKnD7FtRRLtKr1BucpkFAb502ii0lT67MmL427Y
OgJ8V/1KZEWxe32LrEwTnz1KAlSfaDxzysduavBXy/Hc2NKT66WAnlXLnUmX7cuW
9yw5qzoIfFOmy0DWMfyE8Vw1EBuioi6zlx2MJrR/mCcs0Qsadb5eC/jyd5RhuFfR
PVvwnPdkFL5tARL6k8jqH5NWxbMSnCMfNjsyQq2Ug/5yzTmH9YunmyqHhsIczw+N
pHXxPJoGIZ2lDbN88cLkbwazp81PBsakctKi9Cfeh+gzpFUCfl4sW8/W45B+2oTU
+F19Bm1hk0v94iSf0qTpnJDBJ8pYcNdwJrChsxk36FlPyfopr2N7g9Fhmh2GAQfz
7Y05YtsM82TPIruKMhVc9huzU0fu00Ifgn+1v4HniJcRoZ/5m/g59vYxYFs6Gb7G
zYRpFcGvSW1R5+hMdrqIfRl0vuWSheEhoppZT5r2H/c9wYVjRwECdC6CyCfOpR0u
kH52rVaTdZ8CBwPs+ZQQqsYcb2PZ5Shx8S4oLXL5ToTQQRm4plPAPJceAsiT40bw
x7Le0OXBpOanPJS5bYVybmjYTDfe1SUZXAAgYkds47BWDuHUkY3bZkcw3gPIBsY6
WPZ70gY2bhYdKzsFpziU4WZKvrVqTLvBCxpeCpZ/4ql38De159LSMd8oUHhAOHMa
4CULkUKqYjOPXGMic3BrJGrc9qaUjwDs49I8SVcb0HXYJX2CGbB91X4ZL6SQVIhk
ffl20SVndB212f+5ApOCICzjhL0w+WWOVth1HPQDfgfxXnlks948l9OtvzPkpr8C
Jl2xNGGsQ0vks5s+nHhr1uDaiLiNSk42dtAp8d2gIOJBzMH2Z/Um/n9D4EDcgs1J
wFFd7smnB0w07YME5VovW9/gVE1bTMOFnBZp/70bBs8OpiwPCn0or12+kA8m32PP
ZXVXuNF6TPnUwjaufpZL2sqPTLAhvwZDe1BWtTkY7MZu/pzsMtcNBp8Au7FoOExf
bXwlbg2qdaaLMHgiOhmEh0uS4oPW2A+0V93394ezY56DBQL7QS95eJcmyCNAvrGu
AhXpwbZFwVx/mc0l93G/q7sdk0uo0YZ92Q4t3JzSI9X51hEnP8yoklhFE8oyt462
02lvcDm5um4BBhtXS7W3DU1m7Z6pQNLfsKe//nHxPKJo1h5uw2jslsmi3pTUm739
fXmwrnXLOXz+ctaDF/vmIL7qpJpoem4K1lNUeqyaC4qy21oA9oh7llI+pIFjMRdG
bq8krowmzJVi8tSgxpOy1BqpISJf1xeZV0kfs6ZxvNdcyn5mE84hcJ2hSAppqPvm
9auj+FTCjmXi0xw7LOyb4azJjis7HNMo32lE88wPgWsJh6SRz+IY0SUkQ+2nCjFK
6mF04hdgydVZu04+W+d1ICYxfuFtyU3FmLA9pdlk++p+7l1MEZpMPV7m7wV2EPS7
m/wzXTMpLUabPR6IBNyS9xJIAw/lEkFEhOzIXKGb2d4mwS8fPKeMEWIm5cHglOZ9
jJKC+syVpGQBUD1zkRoVpcGLjEJiQASrczU6awKIimi52V/jjogIDCMorSA7gdlS
QcfokP1PR2GSC3XtdBiCj6jg6ZaEyCI0YDwMPFcWHTUfFFbwpcpnWgXo6XP6v/YG
N550cZBpki7yQSxZAde4AqawCiw2QTQFNn+uit7J35+ZcfCjdfqdTlanmv915s0C
IPFSEX1jIGmzy2D+ppcL8zqSxPxHvbJ5XWi8XalcmIAr8niMR72L+utlGQ1bog2o
l6bCCHGKCzqkDznbY9ZKhpDTQwaqvPO2jEu44gwWP3/z/1CiCLZ/5Ia1IGok1yl3
WmrEwHzCc2FQkeDGD1GOtw2LAgMsNQjkBymPQF/M6hfURMM/WjTPn1Mh0AcTw6mJ
NSuEuQy3k/v3BfrPgHdidMneAr5OSR5pK6d4wOfxQKf3fWBIVdvhFuJGxuKjQFER
c/MZAh6fiLy4o7ze4jZH3rI1ZWgGSfzU56Lub6YaqhDrmOhmfpH07P9wONZvkm6K
6puFDJv48UGoZN5CGelWj5VkcrhXwbeitKm8Oc3URisTbmM/jYH53pxDt0BDfPsJ
ZGnj8LvdOPkaX4eRGiWiClDlBF0ofd77d+p9kldx5qo2KJiiULjce7Q+jdClLb2M
XG8fpAtAklCcQerb8gbG+vVH4pD+5rWWvASF1m0idpRNOBe9/vhhCSZJufOXMkwU
zAPVcQ/WIXsLf75g5GivmbCa7guJcA6lXdkQBtEt7p+zj1rMuO1sK7k4taGnkeOX
q+gCzxrn0Y7+MoXpmtj7SbTHYdsMKzJpM7JWqE1LOg4GW/fLs6/0dtnejwAJ8A49
s3BxacuVCwwqx6R6V+YEUN58vJqfrNrmoTAVWrdS2pOkwcL16aLE6TKwUCwW2xJc
zMowFrQDsyr9iy7Es8B1TJkt1DZmfoxtodhpdYla1bZyLUsG/uZXywCTzICp7XPb
2uk5D6jLN+w8pq/HbfCeAhRk1l174PFX2BTyYHqGzpLrSKtHzTP5jL5j1/6uU2E1
7LwGnVaOIDwveqJRzWXztroQ6Eh0jFjgNI8RElVLegyJ2OlkGoWtchOKISsoAyYo
UINvGQaSSnwt/Eh+/T69Xrf2l82BdweelgdkBpJRBYn4omc+CYp1X3vHApKMntQN
u+BsXH64H+yZhpVjsgZf9VI1cOvUFVbiTYZiY2OV/AIr1yyiA4BSbdLMsZrwoRUY
WV4tKCM/xAvI0cvU3ki74Ho73GrrlTsvwDJhyjQWBxbYcVsBqddeXC/JT/He1E8D
UOeNAvvoxJGDTmYkgyoFjvcwvGsvpkCik/CM/SPULQMYQ+B6l4q3fBehM9Wygto1
rXV/p4ZEXeUKKVCg+yIOV80zf25ujRMPSNYQb1pS3dDL+7YlzvZ/bkDxWY7PpHIq
WPzaFGQ4skqbkA8aIYN/DN+KLxpdgFSjjO7SW46rDHHkp4Y/QzqY47Z5mS4oHe1W
5UAAMygCpOQD0u/eJgpTKksAJ9GHV0P+sN37vCnu8eaDPshOg9eXtycT1bN1028J
yYbBdzmjaB+5wsy26m7iOKKRREueODoJRvFj4To1EoTqIrYpyEUcvnNVq1wKSrZ0
oZWnHwqab0ntOkiMCaF1e/F5G7dqKZBbznZ1tcsd/UKbG9uw80rN+jKO5u9vxSoc
Y5If4igJ63U5D6pAcIZfnNs/6flHe1xYf1IFMj+J2kC8kVO+Vgg17bKDhA1UyG2o
JFfTlx00xuaKyZY+Z9AiIj1e1w5R9AnjlSO8ncYZPLzftqEGQpVUys92KYef/rkg
mCFwRD1ToiPUzTrlJwcU8ubAphmDV7ztG41iBLvpzrqPXhdSiUBLKxuOr+3gRS3m
W8x+8oR2ahetztqWw0mFZQv/yGFXfJ3USER5x+sAAaXgKSSTl3fBKyJ5e6ctcfjz
vVzOazzpe7liAu4mEcDAnp3XfRjgI8IBze0X77w1/1Ud9riEJAux5dQRw/u1qXGG
X1VqKf6Z+w+1KWlbefivBSYBBVrHSCHWXc5wgiDjmzf4/bFyQwnMNppnsCW+cX3Q
RvLSqCVFDtH9CbvnfsqUONcYDfFQzKv9j8q7VvHEgrITYakMc23U6Cqa+cEYnpzT
hNMDO/PBPbDyNHnWbM61JS5MfK1ExtimzSoE07TZh7qkipUUeFGO1L5l3GKbAeUM
AZTDkJqtwwQImA+HL7P5cWEvgQd/gAjWMtADJfUh8UDLSp6zpTXODXrfDcFmr9jo
kx/sDAyAaN74/Bk1Hr5UOKNF0rdQw+h4LU1x7paGE0weF6m4yYwFp57w1OD1MyZr
gxad+5q2f0ePrRJ2M4NaUF8YNkW5lbw+jAyAUEu1Z5XydPZKf0WGPG/dU2OPmF+/
R3sofvpc3+dqmUctyJKyJnMCq6I8gJEg4aMY6D0Y0l1LpuvkL9jEjZiwvpHPLXur
2mrPesZ7yZHFLgCK1x/hhAktU3XnJJWLqMMnGOi+sabNyV/8glmEtmRl+FWW6gRG
MtOUstbjtWmbduof3090leLi07iCyN90a+bMnFXVdTpvJ+zpRzCcFaCwZtvDNJHT
yVMlQEiLvlbAHHDH6DWYzTWkQMKfBa0VipnDGqP8ceRLByhFEa1UI1QjgvkRClvl
e6dC2drNxI8FpmtyGkBrFoc1gqmdgWJiNwbe/44rbfhlM2n44hqpTyNAHDT2YgO5
/liIR/XaBTSnnU4AOhjHTKr7uh/ivQa2Ugl/ldp2ReTGPsYX4p+3dkK7BIHQWDNN
QvwPBg3IhfDgpbSURGZIrRFANkw3QQ285cVm4YgsYNYNMSeQ6GsJWYGaXoowzT1C
GDPqpfWbApPw1jVj3sKD5C2rAqmlE3Rt/g/pbopOwsPCipT90KUPcnpjruXRIY7L
GJibdjgUc/mH3R1lsqcx3R4rn0f7HflmiSN8xNuVqPfU3zmC+68eHNiy50PYu14l
Wmpo4aQIGDs0H1kJIeTMt9z9S8UDDNC48AKXMswf7unV5sIjCsQC2/PYRRB3fAfz
2qhUePsnHK+PhmTU/K9Eap6XTJQuH7dMrR1m7ODfax5dOI72Firvo5mIivGbvQ50
KbN0IfRnb6zApeLxXswPX8zO7BZ5jG/aZYrn4gcnGi/afMBFGxCr3ervN5iWNxw6
PgI09tN3nJdQSiKB398I+yUgfinLb44A+K5CgcIQw7Q03rH2ZiyWqBXWAbCmCF/+
POZuBEHcHM6HyGnsKTkO+3ujZv/oKT28Cpn08riMGNIoK5GXt8mcXesrOPYqkJIr
yEOVprVKnGsiZBKYWyoxTl4aoNjDX9RmxmXOE0cLbeOITGprIfdeYqi1FOMPh12V
24GlHVm99rN3gsjgaCwzEPKQIYnNbz1adey1n2V5pmDZr9DMuvs2Ozj1+sMxz8UZ
WTggQxoRCriO+t6dZ+bvCEr2/d5M8wgUFmrvqpDpU0q/PVSthsVWAbeBt7A1vgya
/MeahhTrDR9R4LV9okViORhdK/lhBHMYhReFHwJH74RJwFEH7lsxu4f24DwsM+yu
fUId7p/fCJGpedmrlV9xTiGxzQuLS4ITkTl0JsTib59PqLBKSRQIMdT8bzemAqNC
cLqYInumD4UcAP705u4FiCGUpC/MBGDTrkWAOIdSXiH0MOwVlBEdNci++TCveD3+
TtgRVuTeXZPlUuChWvSzL5naHGY/l5kGQIDZymloRuvxMgtATm5KIaJTLdO+51xW
kZDVh4f4s3N4zBJjPx0ysQCi0o0rScmUdtnhqmLteiAv4wJk4skCqTvXWgiar2p0
jAg0uRJg+2O9w0JrQQ0KyQXbVzbwS9mGrVryubKiWWUjbSlMbElMZV/bG9DYapen
1FJYSsZnEPZCC6FSLxCqtljf0w6m8UrDRPctECGf+ycOZ1cA0lGZG2e8X58eTVK5
6UgJ74OLXfYtz77LnvHwLWgnwl2BQ0K710ZXXTOPLd56m/kPUQ0d10sygk8gPAux
lFz+sYbRIBMLWtoqOL/AHOrKtO8FVfgB66Jc8lzKMZnwqwzH93wYMkT1FSQQHD0m
qpJyBOkFcigK/kn9oZYFQmzbzo50qPnMBbWJTWqko5xpgaQK/9Um+0b34JNHaLZb
yJm+CBTkYS4SZUDmVhH22Hxpqf/7Jr4sQLrFm91nfaKCKTgW0Wc7v2mQgqIRnOPB
NxYCw36ruAvP9zmh0tZD7RTIynCAQACi/jtKBqPGfs9fzKnqoPsx+em3ktxXJA4m
qbLup1dxm6wPbiSMIrFrIikAp+lxAnwTJLDXVac2aaDlNhNkjuZehJGb52kfgxoO
JUcFTDfBoc5ljJMuUtk2FO6GyxeSCYQ/WmhmVi0VEjKKvNyu8+4l8t9MzQpW2rgk
OE70LsCQfrMh3zEMpRou8TPuGnJAp+5G6Kpq3hw/Jv/0mAd9r/psK8UtYKXaYCZP
aFo11Ueu7zjWAuw5ZbuGyt9ZkY6UGDfXtK+wa0oHeYbaxDL0V6f0IcpytwyZ8bgf
+akjicVjsENz9QQ1vBzZFV4Ze4E2IPGWndwaFM4KiP26jAChQ/4pf5vjacKs/xX5
tZeJAgoLkcYUELnn5tpsHrYbUKvXEpL96M23gFo/gb9WhLzKY7LIX7XJNOMb+R5c
1h9WdUWllTGzyxD0Ka6ghubsVO8c4j7KJ6c4xqqX3lvoXUA5SEarRP3ht+gO8SEn
MOQyqemQKhiBGqidkxxhTwbwF21LFgeKGI75HyBVKgfS8A+HXNUc3p4GxJUwbqwq
g9qeyZk3Gqw46oo36sQ8xPrrmli3FXk2h//3QilvcjdqzrW/aCp0yWftdW5yBzqN
ZnwGQj6cZ1JtjKKh9dDzrRI15v8bIfv7QqTKdYq+9tP8HU5F6wDCcfp+SVjkYTgZ
E6kS/V3RZCbhFw5F8zlCbNMLSvVvDNXBAp2ln92LbFhF2RxN0VKorqNB6k19yiVh
2TahzUxHacHfrwYYu4inb+gud7CSNAw1Tko5IO7Nj09Zo+0E0RqkICGDSpuCz/iy
RnKVWou6EjPIYgvYUtm5BoPXH/EvtD409+csluNhdxQ4msOPF3FBp6Q0tzfunZ/C
nXGRwH+v4CgAG+MVpm4XXjnI/r6j03fECmhNDgZIWIRp3iIL4SfH3nSURa9DrYHf
3MAuWOllCSlBRw9Fh/mK9y+VhbuzW9l+A9rFafdUji6sENQyr2H7utecPTCgmPR9
oQLtgRIRbBqBoyk6mcfl69FuQ7SLL8pQKpKRaLH1BGGgr/bGLCaJee1ILM75rz6H
7MLEd2B3rF0W/f0j9wtYm/+7mni5uh+AW0GZdxzrrn7c9GQeNEbfyIMfiFm77MKu
WqwCZzFCp0zfSZR+EzLtItS1jBdq/qzgO8PFTJqBOCyou2r5cBLDRLpNlFf7ypQ7
gvkJfOPInOafsi4Y0yHNOJ3dnPqUsvBo5yy6Uc4oc2K8Ew6RTKMRFT3ahXWgGDmt
qJBTnKeyEHLfOGwz48Wx2Yrw0u633ctV0GBfGfxIzP1BCHMkHj0gX/J+TYbTdFm8
6IJm15KqANPAPI3o0wjf5SYmS6Yn3e1/QjGzKudBJXHFbnDriJl0EJK1NEN9stc2
GWcR79EaL/wnN9gK7gRgZUHT9dR8RnP2P7aFDZBSsYYVqiIqikqv8N/sRjCykC/t
cyJE5MXZJTtpsyrEY4mE/O3pTM44ghB4/HE27NM5BUqBwNjco03ZpdQRqF9dEYTm
2UnYptWryYjXhSWpq48Jm6CWdA4MlnAZrwW+Q7ZTTqy5fvQ0XpYYZlWdS5qDfQFU
ZWENyDV3Q9BLAKcgPrNkoWHQ3yGG64dY01hjiyVvv9WhBkrJYaWPTlpExGUzdmCg
beP+FVQaKugRhRUHP/PtFcxKcv7CzbgZEkwik3fo0dAfVAVWiwN2+Z//0OH8u8r7
pQT5jc7iHpLYkBSPRYh2gC257fwq+wWpsmYmJlupTE2HhJZlmE0bzrjN+nINiVQG
CZENc6kWK275S25sip6ARliGy9kZAjnDKTr/1GzQSIbqr649nPBDZHXQaNn9zHSZ
lJ3/v2NDQOt/xUs4DIjVmbyEvzsmjSZjuJYiqpSkgyuDwx7duVdThHJQK63jURRO
S3FEVF9AlMpUq2pxpimOZ8bHm3vlASgRJklQwFwsjgMmm1OaE7WJqGem/onccNkh
e9YdHy6pkxnXuNM47kQxilUH42Fj5Wil1C7pK6Vj77yZEdKjqDvK9lbJgU2xTa+K
Y+DRfVA3k7TnvcWCbgaegZNW1pY+s1VghJzA+P6b1b1ccX0ves21aRcI4uPVQoNG
7vKdpA2zV8EcMiavLg1AgOWyZN+kO/LSQZ+hXs9jWLJpDMtrLH4wngvUaZi0u7EQ
9GUqM5Ck4MRsmfLKMY7reCuFEXq+0d63+BBTakYlaRPLkoZ1hyMgNBRPwsYHOF6R
9XKktDTydrF0+/+ftxnd3sgd8sv4XqqfAG38Y8A7PmDYWg8hMyIwZ2jjxnuZY8Ea
SuK9o2UwReAmVPOAhAvIWkW6VdIASABKfzNpYgZsyPlMt7BBAJfK/Z7159SOl0+2
knDmgR5aWDuldIMNZVCWOiykdizWMREnuJ0qsBPQbP3/0wHp6lQk+WDAAGd7qpYh
klR9uXwzQqdwvOwPifeHDUAL0HE0YVFULYFjjqXdCl4l+zC/RQUKeCkHIVSqY1NX
Ez+/HIfBNuxzo47l+VTGpXUkXBhjdS7TBEY5jLimUhGQOfYQOpJPqm6fADp/rpg7
LSYv3kVn2EKmimV83Q7u4SA95vOOpiWBhznNHjw+//4LBk+2yHutU3PXog6WIi2g
AzNgy+6g1iootWZcL8YapnnwDqMyBGCOPskrE9eCpT9j4gzkJkNfjCPXkrYxLUuN
Upx2q6aoY/m55k/3oRITS3vjQSFnj0+WqHwuyZ9KS1cFqFHY7er5nhtBQZsB+T6Q
r24ijNmaV5/dIZYDpXk69WvzNknHeGZgvn46qe9811r9ZA/XZfxvPwAPFKWjpDos
AoE+Jb4Wim5n06T2bFbf+1bhA7EUuwO3Vqz3bZ9A2pJlce9V+Y95Bz0PeMPm06O4
++4cs87ZZWly8RUbch2J4xUn0MAwdstfbRnWkRvHt04aNH+FCJgLpga+jO05fmmO
G3KI0E1MlQH7HlCeodESPFoc+m5EeSugeXmnGs7Va275gr5sP0+lL3jXRIZPpfT1
wXFuHcdnY7jyTZW131JnQ7mv7Ol6ligud+Pc+BTXeBxoyOkAic+UK13IpGBYiweq
7OuY1T7zAdPQOMpT/eXfOsUKQTaGQJltQZqVQ20prPXd0VvNZc4mrAFbvxd/VJHU
1UHI23pfXf/lCitvBxVmu2PeIEbSrGpz4o2HM5bcOyxgeyIJIhrFJQtWSgjJ2Aqk
ghher02OLD17YCYpvTtaxx7uYZ/TeBb0vLDZ+aon0UyBq9TwUY0Au2Pu2mFAoS/i
ER6LDTgkTg5RrXZCa5PtJplSBsbOIP+Ql5K7/w3K6rkzCuPicAvepxK85K+9WsQd
GgBtUGmnghj5hhjuBOcCBd382pWWIt9DcJPfT6/PZGleoZxmvYk5J4fxrZpHOgiD
y79ACD/bQjBIa/fwnl0dcrFMBvvSSHyj3cikrEbRFfzyeVV4xPAW2Hs1LMST5SEq
R5NNI6IhmO5IL0nu5eknBaDmra50iTbVkP+Duegnd5MJMzSvO/5UKICtH0V7ESr0
d0/FLUSYD0mFFweLbKX943USVyTQK6I9dk7GWOv1RxVTBcMf3Hiuj8UnhApmlLNB
cx9kDS4rpdEDQl6zEseOHr5biBelY5ZR5Zg1nqVc9dfhmpmmwnGhb+cmYO0ncnZ0
oireo07hamI07O5wLRVBqZCIYIZYNRtkWpYsgJQ/yOcRhY3xTyKAJXX4S4I1caTh
V0lMPzfKY+wQ7I/IALGuFF4W6YmYtsYt72pPd34dopdfAh4CJa4nZhwZWI4Qv3CU
C/0EW+NE9tGHAaa70NFAMHnJY4djyinEIMro9j2KN0HMSfbpZWXEsjlQF4nOD8cp
7umVEEYvIpOhd45QtWbqcAUp0vwsYOPvyAoVSaPap0gttfOPMXaNNEnQS1hnljbX
Vp+bwF53109+m3Oaof2NLgIfDFBfL1spD3VlZR2pWuBy8PoSRDMXrO5GQXQ2cXup
SiIn2CNffOPketleB/eji7P2E0bJ2EMif7MjC9CuejuWgEtHoip5d68eH7HaRxO5
8oZ4KJAxMMSewFEECsIuciAGTimezFipGKBdU9IzFK50UsdssPwwMxjikhoVNO2/
B/QZpHze2DlsINfRp9K0e+gJRcVMKJkHBdOqhg6kHjANj0DmUnexRA4q3Oqhy96S
hW4n3x53DvVvtpO7+9mNxCC7zzsSGSFEN2ZWKYXRQFQinmrNPtOiKIn9mPPCtr4L
nbgimxv1Fa+zpJmBljNfQd1tgz44+vCAxAGbPEkMY+61caaR1ChasIivWqHoGnLI
EPWYu7ZnUzC8A3QKMhB6K3AdSnC+7su2rWGsIN80jju12ExxdrLdkgfw7ZucAOuj
O9ijF4JQSDiOFaHkXmxBHz2lI44yxr43TdU+naRMd2OmsBSsvT8eFFlJDErd8xAv
yeyFvdaTCwbNK78mNlqVC/RSCbKmW2y8uzK9n17ryHcYoclbsC1t5JR2sux1Tm86
5/DzpDtMyvYimpz06GVUvxAOEJA05v0MD+SqCnHqyVwgoXC5oanlc/eaSgf7YPiR
pqQbJjcNkxV2IrNcEK0Ye5D2x6IlOeSY6CZklxU9D04mf54UfICGlKMLuCrEOt8+
g2gGLvqY+m4TMbJa3+BwChHX4EQ8eY42gmubqcJHH4dUYZXfpRw0sF3rItrqPRKX
Ala5r4SK4RKsrjCsjmUh2vAxa9IPBE781XuZEFVwRT4+yDrNQNID58dx/zBALh8T
4zId9c0A+Wc55zqmRYoMf66HAdm6mgSdQ0JNf3ye8obREe0n6BM3NtlfOkhe5vgM
fRpsFFUpueyarwTTQdCcIfbcIUP7DwZJIAz5lwbs0IjaII5jvycSIG/+aeM4xg/j
aGkWpQD1IIcfI2B8Vo28dJygtOioy54xrmWy/uAzR9DqwKP1nhlRZDVBaD7mRXsK
4V+Y6q/Pp3YRPxxX3N1xQ2HfWuwP9E3hhgJJHjkES6EMGtQzviNvtclSLtrbE+bM
6PZ5ZlljL+HjjXlyUH4+4OxgtxiCgG9fbOqbLLHQXtEsKkkNiCYoQ1XM/deYSEmq
D8gHTF4ReVJXSQyvoAqkTvIxU9Dk9IRBdaFCik69pjAVnUzNWiZTQI5mn2GeP8M0
coTRa4S7fmQz8DJ8h0mU8ujMiRDc+eswoH0WfKqclBO0ICTjpJfxeEUijcUAJHYk
xQYf54ebW3lDUfDHmn1gygswOn3/txa3YqQs7UBTzuiqJv7bXMMi2q/VBc4Xu4at
FitNcA+awCasyB8HScdqtanirBlC+qmFGo2AOtKgaIkyuHm/buJL1ay8tB0lIZl8
qsdkmlin0w7XktYA9ojPE1c/8qEdld9vKboUCZeAzjAxjG2Z5qT5wrNx+XTs48Zb
3yAz7qq12+WbhVOLxFIt9WtMrfRAcjZHgA8S+nwZTW3o88NCHoQcrrkeeJ5IGTpL
TvG22VtGtjSYlBT6cH9ABRxS4Z6yg2AXaTl2vMohRHh09JHiQbZo61hta48ERNw8
DuadxQa/uqFXcvWyEbe9lGnmO7VGU0HhzWB4T9TxHJ1h8D+E17lVVPO7Tbjb7IWW
bovcwy7ZhJbV604uT+TgFEjTZF4LVWpUCx29ppXAYQP5J7AnJZpmjeRdLzkjTbMN
s6YCWeLU26MGi1IMIe8FgSOobhxDreloxhs8MVaiYHf3lxEUi73eSMfI54Wsknzp
z0fLMN47dmDfAOj1kAzKmP/usEY0snJq5uqbfGTPJGcAaKNpx6qX+vcsUg5AyJgf
TatDguQFJAjOV56VTqw8FtYbhsISH3qqKxaUUKknBEpHnEit/V+sDWODpoV7KVGc
r8Q6WX0ReV2YuUYAZfE58z3pTY/XAYoSYomGJxHaB+SRvzv2tqljDsQAu0FZWWs+
G0q6Hil9qOw6vIdO6Ki6TzsQMvTtYLQrSsDr7NX6ic7NbpJk59X4cEyMGxfTVz1s
4YXh861Z3kdEn8RI6waoLbmTz5MsIMPegIzMwm0wgOGUylnyrxj8LJmLbxUhhtpI
bOweYqIx2CCVnpdeT8L+MJpALuCPBigNMR/nhEX1huUIAcmUH+ZcZwRXsMY37aSa
maVn0FclvJ2JB1+xMvrHtA/ONVpwxfd1GpqE95e4TR2o5L6aOzM4sr/voeofpr7r
nw56dlSkpGBQzni1i78c7U+VWs6oGm+5RmLvVnwdhUetqvedIxH0d//m4mQpONcJ
os5f2V2Eng/EzVrhT/occ+PgP9BU0fS3TBJ1lfQXLe2+DLgKNCrdejbJeVh7t5ca
Z0gZVM1fjIMpiBIk+PyyKvWK7ioG/j90M6gqTzCfmJ1x8tAMcw673CqZiu/3krOG
P7Z8F9bXsr+Po8G1AmjLay1WmJu6Jhf/HsQ4pDJ7GqwvPXFtvfileZ5/HniRoMa9
v2K2A2Dtq8IMZ3BBycwFyQOnk8NA2P+NAj+F1gQ4ydK+JRvfa0Eo3ko+g3HDRaf8
fV+ZBaHkVJ6q9uURpFNzGqrAHPTFjd20bNWzEDH7RubiRmkB4Gub5gHHkMlIorcv
G5/GrK9x9jetNtS5xJ9jUGPmSE7SLOVHT+zEU0rzFkhermGV/9h8Vc2u1V2QLdKa
to5WcUSYvd15QkQH779+WbIxFFOOhqjZ1hMoWHABulfGKoT+C8GDxilcxnu559Hm
AjpIsnWy9sFDZRtj2yT0F5LsaLuILevNLC1vpyBHRStgCDUoCseOQvNWasO9/A9u
k2ZWh/wNfMwsO1beJlMaCINIeIGJrn/o1QbWGSYeu3meyMPY5UBebnbAzUTomqVt
i0XT6cMnKoTvmOYxqqVzLUnffrOnI2q0MFlo8e8neObBik8G62KfNBUYCkXj75er
UO5GolSITb0wQMzZXNpXice7Ree3aTUiY+/Lr0M151JUDeM6CSB9Ukrty/Vp2DqI
tSUx2OhhzUy0rDUtCHZ0SgCCQWgCEHu0KI7Fl63yG7U+f9BVPdR9Hw3Gz389b0cU
YiugZP8Eai6UMYdO/pTXPYLHohDjXxlJMPP97nEi7CUj1NXYlSwTihuEhQR3SlU5
4zV6k7bc2KyQh0dUZ4RIfiIyw4QopqgpVhVIPGPDaxvNrzu9zxVRxQQW+Y0gAxYD
Jq9R5la1KRoLAi26jhOOUZ8xSfBhAjeKd+oNHXXmSzuATBVHoA0iAOGe0AsVDsTk
P2MfZ+FzJ2qvWo6U63qEX2oxtP19lbfesJI0nSVe6+nFmtBAmuR0rD5Su3OmybD3
5tEbhDQJRTCOZTH8SOHCQ+Mx4IALRutFIGF4z7X1toQ4IvGAeIk9HpykeVLqphba
QKFOPD/4Tu3DxAq1XCmG7zhQaLWRhSK9Nqpn+hZNxZ9yDY4OQDCImvwoTanbBa74
UMRw+qVwx165gP4zXI3OARLyPlE5zHodXQGCp2/jk4Q0o+aXkJ3U3/1WujXA4EdI
1ZJaauTvSq0rC5I//HqFZVQQ/Y+/CeUWTg48Ix+POfAFYPpgoKkCV2oJT6VjDMOV
xlwInrh2Ehp22lkf67lOYHe7c8hDNNfPSmn4vgQqO+qHdUSVHAQdwcABmZMuD2SB
ZDfqKI927TiyC79BN8N8lh72tFzmHuw35KM31lUGj4sUZXHY2CUJnGaKHWn/Uq9P
rWWIL6OJXUziB1U1mh2S2sFg7d0Y8Ixt8BA0l2BWTO+ukXB9fnQv4XvFK/KW/6j5
KTMszWbLTTgBHJ/FrsEUvRJ2kNNf67KVj8jpNMl0cN8pM7HphwClbiJI9FApSi4P
bNhPTbvuBUe6FxDkrPvzmM6y9lEr92NNy4VXchcZMWFoFHM93xenXWDD3YpgaJgo
eJ16Kedt4bXgIfx56PrRC83jf1Q+/KqTAHwzVOR3wQAUsHSyrNQZSazvQoTcBmki
ygASH2bhZxYrq/kEd+Tw0BTQhgdaPLzcXZl7ASFxVnpIZxLzhrj2hfHwc1mJYtdS
WSqiIvcjWuYdGRAhCYypRmyicTU8dS2qTxgPwI6VVQjBMakFotwxBmb7xGca2F3+
bysboPH5TyLa+LCxB4ls+VDOKVuLVG3eur4MculBSasPRCNSttFywqj6xf/n/G0e
Yo2OpN+Nc8BvWbQJNoq1oW1XA8PGz1jSV0FRhUE1iUCNr3Rv4OOMCkqhVE7EqHdn
UM9XyHtQDS5vcVvpIe/zVXj+KbsAn6dNTKh9ZWP/AFvvJkB3sx+D3Pg5oI/DPiND
VTWE9aGLR/6gJ1eS5GsqhMoT72Y0ZvtnZZygExcKuAcb8etuuhkcqyN9v7tAyJAb
KZEanF6C+QaQz0OG8sQoo8/vYtWkpF9WLmfDHEI7rMdDYylzxx0vNRF5se+nyg7s
/rR9uNSWDMWD8H82b9JVHz3Xnn3uFNK1lWMYlONbB6xFJZjcSJmUnen6crSmDhI7
MHJjRavKxe7rHdHbOpqMKPiN9ZBlMBoOO8AAGSOSF5qKXvCfWAgjYgDOJzx1BN1e
GtQP61hf7m5lLdT3wP2gcn75X0SlaY02VzK5hWJ+yxi6wIctA34Sl0jXB8sXoQo8
tZHyohwwC7FP2ZO1K+RbViyUxdVnvE+2jMImhyy9HtTFHlm/kDduB1WqQjbcI+K8
K9lo6aQtsuT641hkm1RhjUJB0x/tAAS2WUWKuF15FnlMsWG7QE5R9zUyO0I4vyFS
fQsmVEJjN+4LbYwxnXeyHRDsGXqdryOddOhmA7IdT91OBWap5xaNbZZIvzzFnih1
Q8T1ZkZOELvy/5SGzgVmVEZiouAHBKgcUjbst4APuoGV21LRaxibgFx22jHI8A3U
2i+lkkCMI/vKu9N84xpBX4jpTBQ90T+ngq2uzQfWa+RGymDC3pra50Ze3lV0HjyS
PWa5bzMrHPr6wkk7xOn/FSBCJa6t2NYq687ZVrmhjw5tuMLCVrKWTH+pUUsIHQdx
zRCJkSaC5WhFz1JAUSkxdNVfrZdn6DgisHQbohsb2PLgZp7e85OqgSpM5xwnoQwp
pnc8DVYoEOz4PmF3eECDTqB28qZSxCDgMfWRsbHgq5XfMfw1dfy3tBU9WnRrQLGM
LkJPo1Hrfr4Abmss5uvAsMO5yNYGa4E0eswGP6VYsoPAF9vlg3JUT1tR+3TGNsmh
Zcxw/kD7pu7lHF+bzPxzutIDyqkfTsQZ5OIgYcCSGbYeh0pYRTi4vitrrL7ifEqo
FO2b9g9Ou/lHw8rVEq/iEAKpX70sNNhhOttFpQpdmgp+ii39mBtjej4ygSHLL41P
KPL9drhSNMVmli10QOhv3XHNZxAk9u4ebAkYYsgy97HQRsvXpSuP6aE2R9C8jNx9
+DdoPgG7BKnv2+JWceTBz0yaTUU5TnAHmUFW6o7DMXOkM5Z0Eh9p1gWHkqiZhjYO
xwrQhe8LfRN7lM9Ses9ztEQT8qU5/qkumHr6rxmi1CAlv9UW3R+iY1PE3VLgIgdA
e1lajkoDvw10NkkDqWznKx9XA2qqgV3FXl1t5Li+ZGL4wLhyKdwD/r/zaFTsv/Yz
cr9N07BoksWIxABEp+Xc+MCmuvRwsO7FPXNPqpxDhzpZ9c2ZfuZQnMVCT4SsAQBi
17AokBoShvHnmu1IajVnivdRPh5AgKW3wLRQ6q/39F842735REKYJGJZgvcxRs8i
DyMXfTZ5xkQxNpfxO7UzFZJvvM/3P2Mx+KQOsr8CCIMLGJ4h7lJqwcon2ufe/Z/2
1Aj0mS9kpu1zPgFWffYzBCJbhONehe598gJFDjEALske97ci1KQj7RtGIMM2zoN+
S5W2IepcUzQPprrLZmDFUM+4kZCyvs4unMJcMxlS+W3nQ9VyFsn+cNoKU/SLpLSj
k4DaaHMQx2nCCpwtPAHyLIbDEPbgBBgEKsfONrzdadD6wRYSY4WtBdVKLVgqm1td
dXWiDHpDSnX8xBfyYUAZW4/haDXkWR4iChMl9ZI4HQgHS4SWzx3pgUC8H8SjZbot
M8hXKcgX7e89MKuXDndk+RhNJMKPx9kt1f8gkscrBKtto5OvCuAFfGlpnCR0RxZ1
13dJWivQjRpsp8OnllM/6E6Lpp7Yg03EYxjWa7WoKubz8sjYguVjPCPPB7vrp+71
rI6dSrg+orD+yE1dzflO7nw/TpDSxq8rUors4IGGnfCCC41WSX12e2hwFb3s+d5X
Gu/Zq4Gt10VSbYRF6osGbkxORJ2CBq9hJkZywtzH8Pptbtkd4HbXxcl4tKYrSEFc
pCL3zwZNjvYF+tF2auircPFHO9agyE6yw9KTwvu7EOU7SIXzucLQL3Ed1Z67H333
ycTutaL4WZB6G6mj5wlh0HSBxpxsbBpZx3QxYKymmle/g1mvVVcK2spAlI0Dfdrs
TChIsgKJ9dfsNfNC3E1oYFZuRPGHGx1heHX3w+/DmPB6+O10Un/6LTmqm9bFoCu4
gzfETTqQ3cKsQcMxFRzU7J/ysxIpKNLP6K2W3Cwk/78G7yzg90sP5AXeNgy3TphK
1eN/jTXOXD689czzZxK9mTJCx8gmsp4yz9PAtaV77KIJQaeWp2BinYLjehzTVXj7
CwMdT57XmdyjQz/xkeIMHdZ9hARf39s9x59WWFStehoLIT93s/GK+eG92VIjKJmN
v5EZgaqBvmXQfoVoGxVEZKa9I1yAWPduH3Ub+GG9KpbObufFL3EhQWZOZuxX6nbI
1yyJFSx7iam7ID0Y4OFxtgIQDRCqyBunSZv02Cri/cfUhO5xy4nKNtbwVCehISQ0
AzWA0a8yG2UlZUPLrHD2YedTVxTiTZZMIH4lOsM5WV0v7YjpUIGHy303do/XJSRD
mUcihz5KnFYZJZYD/ZSUIdgYW0SldAZuNHv6rIRZ9vR21QrXH6T2jfaUuvDPQliU
5wu6Lk/khIdz5sMy7W0j2QT8wwl8S7nWEmAvYXOQjpV0ZUKbEzBxRm73TAzSK8m0
UAeSSz396qp329OJV0Aq2dX3tcOX0TiIHU41N8f34YET20FXvSGqnHn7x0PNjD1d
NvikwKLP0I/5T9S7dtcZMW+2oJHbc7GUnRtowtoAa1AaVUobcv08xstP6ChZX3UN
wloRyO+oyntfZn9PX+2CzRYzvDQzNNQta6PcjYjI5BNwSHER1j9CpTZTyMu07/qn
mtW+tXAf3JwirvQxyRPtvqXec+Ms9ulMqizGStviEIaaUlYTF4twXCDEILAvBJm1
XJj+FJi/q4mMAZB0Q69KjLEm5mPvkDIUBRqtztJajrLad2C0n3x2VZV77ipkt5Vj
EDK/qXGmNCZXGd5IuJTKlQAr3I3xuYPKIxjT3gyGhzOk7UNAgHJegImI/iHsvuQ9
VUdnMiCUH5MpTlBBnr2QogMdGaUHv91aJzlQEm/Wz1580xZzSYnKy+7S5C1LYDYa
FmdZkClwIQ8lDB9CR0pIrxOThzXIjgt7B9etkKgn+0BoOqMcn6fI+jObeC1Qe1Ob
NoEy38euuqqvYy+EgadPsiqdLQY+xJmx2smNRcaBgTuYRbkREJfFEORk0fTs0QBu
fe4V711upiYB5/MrWASSAdy8QOD2nr73cNoX+PF1brHv6vYBlz9ug1q8sJullHOZ
QidBFLDi9MrYDsPGRkKuogqDHD7pmQvis1TTU9y9y+2TY7filoG1kxsgm7z0H8U7
2vgSQCqy2gyGtnaGbwubbc0CWuC4J6fDxmXAnT0e2VujUcpPB01PgDva0kgliPhB
KuAkPQbyJcLpe+jLfwaN7kGYQEqlPQXFxdn8QMZBoJH6mldXeRA5+FPxqiiCgzlj
X1BqnTqq1burk1gwLrNGVN9lGqwbzxxT4r0H1Gr+ORKYvaspG7NsC7DLnovm4bPO
YUHT7q9HEt/wbqx67blp+H9ZUvm+aefipJWgREZ9vqyUKNHqSoziAXHphcESWwKg
V5VynGVK8DkSc0Fj62RCMtqNsq9Hk33TxwEdV9KuyIQCzmCVL56D/UsgL5nqyIj5
8jlKUDy9WHBF5rk6UiWBIjUPNgScX0mhGY+T5jHeKut2ji0beuRwEtyr0qoxF9sI
O1XFqHZcUjvjeLMQXRHj8gSA+WzMguEfNdj/E4GsJv0fOoQ5xSrBjC/L7K+1BuoV
yVHn1DrPF+NwCfpwkuWPQ5df1XXUygJkbNrtch0tt8MD6IUrPVvPL6i9ASkwkxzd
IGkd6hhytPHYLkD9dcp9kKo9AVFyRi4ICZZ+YyqG5Fh7zoJLH1aEt+nMnZTkdwPZ
T5minMDGsGt6aVNCjcZXULJZ1aPdsh4KFesMcZn/bJRNMjIm92h7JFyByPjN0gLa
8CLGEBMsBCTPgR8VuWRV4QKWOrRkEV7TU5QSmR50lxOfT6LOvIj5e+LFvRrGyhtI
1ZbUslzQEd0pGIxGGWfX7M3eL73Ftdk4Ed6PYlVYIJiAds47XrnCE1wVYGzGQ54I
A+sUf95id4qDaoYxW/W0qOgzzWpEVlRIjDJ8fpxSTehadF2qciZ3K9cRMOyhTqOZ
2CrPrOgDKPUQKXRsJefZdvA35zs4pqeB2SVYbSyMaORrOAcRSJOBd85dB2oXrOVU
L05HQWTJz4vtOTaBSoabY48+iw8vxOoFEM+1EozCv+eAtfMmF5M40EpFKvaAaMoe
0l/buw2h+TaP1CsDgJSkc4MGv7OlvAlZEY1pUdMYD6Bay2x2DzyDUIoVexKo1cBt
Rk6HASOI7iKBrNVBE9kRnHk9UvU4kWJf+c3Ea2Y4PEUV1CjEPCLXG2StfCQdTGJD
DUXKstVI/ugQMsWOuY48YA64KbyUwpO96DJp9eGodoIxm9ckk07x1f22OhVTJ5KW
S0nI7JJZr1G9kF2jakTqBZlA/SRFAVF8blgW1AfOJoU4iP09daR/y+WmORL27ClE
5RMz10Ohc+o8eytL1Z10pccKceHDyKIHv3yE92yFpRKLMWIzw+kAwHAtRD7uL72e
tAMZmqv5r7J+M/x8YfsS/F0I3WTRAG1Qm711YRw1RumH5Way0Kz9gid9xD2+FeUG
oEIK8/Mn6ryQyXGNiM/1fSOTlKt0OLCEioQZfaS47HaOGasojg1Dvn6kkVo8XIKm
tNp+Is6t0g93MkFHY5zEl5mowqVK8G7LKvKw9w+kpz8kRtxI30Cv0z9B1C3kVXjb
UXU0DPYKUZ2VBiJhDN9bF6ta4iY+RvDc1uR+ATG1fZ0FZIhLOQyC2Unt1IlmLyPu
4i+OmKMXOObHjE1t2srKEmHSkZUWUmvq0a7QdEhTQ7cYznh/T5cNc4A4uRA1e1UD
uwY/MxlTsXjSyc+uI0pUjXLlUIFI0uvVSEauYfICQJGTIdgJRn/LABhE/jBY/4yz
3IJuGWkpb3hlIVqX1mZ+p9hsWt47PKD96TJZWMFKIfQA2hwQ5jjG/6LgafGAMT10
ZbGkZkYhMixcKp2hkuOjKnVZ3YZ4hPNIAVgeaC4iaWHRyKRjt2Rd8xvxstKAJNBC
m6xy9q95A3nHqEjD46QV/54DCewGSgIFWFdX5k/eaLYfJ611qCxxpApAQES84cSs
qjnc1e6zcao55E8P3qsAwveQ1aKz0U8YnR/LdYPJIvgdAmn8tRAPQeGtyZOx531c
1Vtp7FIKDE8xciBjQsvTprr0FE8rTNfYkqeNLpbaFESed6DDNLnPpFs5zRGcVToN
Ruaq7q7ak8x9GoDpxyT2BxZYi0Hc8rWJOOBe9eNWh2ashnX7EozRzBwzen3ELXnX
ZtH/m5fTMEbz/gPSyBDAmxtlPrbNF5XN+4RjWwAuSlu3Hg2aOzhT2MsmpshOd9CC
f/sm1dj6dMoTY1Zb+EhHoX6E37zYy0DktNobK0c3aoQeuFBz2zeOP3HDImwBx7tX
wNAIAwqomDe2vSLd5Md55jrRxzoENcLWWHwmhlP9rnpN+3kMexB2+qc0RSZLINo4
Dkl4COQD9J98vS2Oo84gOcRZFBWuCQN4NoIGMiYUT53kCs8j76A16o5wisH42NcD
860MMbOobWUTksYY8R42DAiuTje3As/T/nYkMb4d+2gtNKGlEO1F3opd/erTU25W
17SnLfQbOx1+ugUa5PZSRyTRz3UzxtKhJfpdGNZnSasYs6kpwJzdZvg5XWwdVZc0
B9/IWNrR9uRY+bsyyodVX7LATAODnSfu0zk+aKdRQI3/cImY0EY3yDUa9ZmJ33fe
e0pb+lkEBD/bBzHqHZmZEO3TZT2sZJJ8YNzbvMi9jrKuzxPsHTNF/ZYvjLRf7z07
ePn5+MwfhpVhVzf+IpPvtJr6Tc8nvsH9ompDHsWRNn3pvMSXAnsI/I5LC+gVrAn6
e2pC/rKt43dzrKUvUW62DI+FncHiEQh6ovkjPdOqBaqiIly3BffhOSAgMUaPu9Jx
fANJe2Ca8mgRs+bSFLUvY/ivvHFclaMZanJRd9WTHdCM1WfDHbFQlNcp0FwlAjE5
/4/+pYkEZLsKrnNY+SfUBGUAIQswsou3z6Tdmzljb3kcjqJQ7yQRguVphuup8Gai
KaWzzgOYytOgpVpXZAFn87Nl6iWfmdP1S5ePdm5y/edgcRxqndB+ux0Rs8mriRzo
4JRl5oHVpbo4ztJF98AVAA6fRjcZhVPQxfvQz3rw0YYun93EGvhWHayXZJdAhV57
nTL2K800ozUeSO7Od7cf1rm1AUCx1Rp4bqbasWuagGFiDQv8UMIPlN3lCklKh08w
saYfds4Y2CPYfRysItgEbTCvHospcgCDF0pzzs5V2ZMBOJacVUJ+pOB6L1vDfGWh
ttxqVFCFfltWJC1Zm6X/hJTgTkoqe/hgO0nH0naaVrHqHvlt2jVKDW5+0GrSAy9v
sCdKjbzEM2JH8tvv9XGMKhVdRYC2owKr3iV5cramib1eyTUae468nFQzL87iSSH2
F9X5SRluib170tZoROdD3E22jgnI079N5q5ypm6LZrRdtfUdRyKQzVI1gemWwhdw
AJeGCxgKCs2Ok3lHA7vpPU0YzbYRaD1jnMJIjeaDVM+O/XcsRBBRW4muHolOAsRl
XmmBOaojnTHKjDLrQZy9jc+gLwtqSMJGZ2p090u6AsI0qusVUGYns40EKlMyDmBg
uliCf0CkXew/sZOsAmKskPjjPpg3w6NSaTi4o+mJT8JgqoKoE8V0Q5gCH/9qojXP
iGoCwOFlMz8gCny2q2MiT9Cy5WRviEsgJMIYMi1nvkvP3gPjCmshJZvxfAsmc2/B
IMGc+dtZ6ltNo5MElUhj3EmcWM6nMsVtHWhioG0XNv8FX+nTZnZHxYaVSEsSdPaD
V1GKDQHK9nrfq14Fsrr3ahj5hk7jz6WDJkLjxQ9SzgiaK9mKGuusfnStfeTLoAtU
Q91r4q9QcwXAjWhOlFN8kCNj9Iro7L7pwJcZOikHz9vKI4rUQuZF0R2Uccfpb0da
MdGwJume4Nq+HCikv5zhL+ym1msyBnXReN8gRhmFLA4F3NMBfLhtBsperLfHdxo2
hoRh1UwsiSJXHEXknlICXvSs4LWzLqvaSE2to3y6ALnL0rd1wttUC0YNDocEUtA9
kQ3+PmRXGzA3LdQH5Knuz+oeAwoMXedIWkmDyZfA9OwFIiwJ+mP0CnyaefK/N7wm
8nT4TRNG7U8T9TqVNXd+npiA+8mXw6ssGyZ/UZtE3OJ7tcRT8fkuaez6tkx12ecn
V+Hi52EX+Ojg5Nm5ajYBaVOp4k/6fOvmdafrCwWHFRd8KIibGcL1uDduooOzSSIA
IbDBUDUtUMMZunryK0u/+yWQP2eTlaQlqTjso+GRBVYfo24884NDYK4Zl4CGMqcj
Hs8OAyyEx/42t89hqu2ZooQZWJKA6S23oaUdvgm6ceLoe+6pw5Lq5EDSbmi9gL+7
deHLUYY5Bpb1N8otsFIjXTQPfkOGTMKV95bYer4gP/LkanYdHbGj1uNhqoyUieWw
kjRO9KZBfN7hU6Udpx0ZWBN10HwnaTIQCNW5aMs6SHJKC4fyY7SV3V/cj86phlAX
oozhNlTA3S6E66Ex/r/04wfPJFnL2QWNAkMoc20Gd/xgG7HE0RMJM0z/YsMaoYPk
M5kBssKc3TbCCItNjf3589EHrTZzQ2bCFil7ddfX4XPgee79o3lj2mtAKBDHVTDt
x22yYafDyOeLEN7mkQGWsgZ6ZNWrPyRErdJO9tXJk4u9DxrPASKjMGHbIrlbsq82
lSqveFbzUrhO/GqHRjIWJPZts7BQM91Xk/AJ2iLfzV3Cp6Akz3bBc5KzBLV7JTaP
rBrg5kEkSEle2++a3dy+YJt61ZihjEN5b3LgwwjCpHSUsFNr37Qn+dDGE5fZI5+j
sJsZLHq0v/w2jEtJj8IIuky1BkqxsfbahF6ZJgUM4CxDq/8ZzqrJOxuhDcNs0q6j
J5n/ikHxWSxa3TJvYObE7fo7bmVF7THloXSqfj0gq8yFSa8CGGJg7qL+NIGzeHnB
d9kL29oaHulP/MP71ztYsS7qqWtD9R4yBrmX2C2vLxT3BfT/WFRy4lQwwWrRbLCf
5McqPytyc6BAU/n0SvcSY5mgNA7UafBA7QMe+FF37lwWvQwdV3DZBgLuYPHpGxt2
12g3jpLF/JB9g3bWrPmMzI6BrAnEKRDqLJg70KSKDDGwGeNeYNVTKmlPAbvPKrzO
gzmgcUwVDBAcA/xUb55k0i60x+rnVTHUf6Mvhr3XxMeuBDgF5uFdlz5dSVpNBw14
IfDtVUF3opZMOW2ty11xirFAENdMjpRu/em6/3uOsSCReVOSaHtzs/H8hj01IdlM
kE+5vMi16wweTHiI0062TI5Gr1ueIdLXYbkyz7Xd++Hq5669ZveYKi+spRpKqh0t
ItXOm8pvHUCJmy4Lzp40ncegU07i/0ydV5bnvZEmf9VRdq4F1wttAge+HeMgjddz
jbGbS8DktZYSuG/7aKOh2dgNbgEx0zmlZmmJc7x8UpiLgkaDvgeQFL/6/W2bIAvg
l05PEeOPkVRixXyHbKJj4hp17Urwnn7mpE9vbLfJ/IJHvw8zyKO6Dhdw2vW+3FTr
RPbvjcNHRQf/D87HtPUC639/I+0n1oCQiM44+46ESjpeTUIQW+d9LpFXJT4kERK9
Vc7GJ99g6Kue12MrUCzRqrd61egK6EB5i9a3H6w1bgBvb82cp0McohwPJ+QnuiBi
JgC1++dzcUeyv8OPQ5lJzQUdoWzBcBhSgISxIQ/C6tN/BvCIxdfMLjMCinO5KTey
04FvWQ5E7h3M6OuzJPsqoeI1F4rt+RUIvgbdEgvqXdhldy2t+9gYdtqGMtU5XPJV
Fh+VtElYsoDwrfsYRJiZZaohvZXM8tOc0X+nmINKEz7y7MBgEZGzLJVRg+hbUHYE
U5c6YkBZXbuSTJyUkMPW7kSo9isSF7FDGlITvEhHi45bHSq5pRsy6L07LWqxeUBx
xJzxSBFAsp8xu+PuOCrhn6sVxexceRwDR6Lzr7IDf9KVbeVu2iGFyWqoFFeQXWJe
+uUZHriglhbA8u+JU+lR2qIuueGvFs/NuKiTwZAOZ0hEq0jeNu9TNKb1a5cm9A7c
SGljrnowc4eLQ2Y7QU7kt8Zh3qLVgpWbLt+Y88kgIkKx9s0627kQaMD70rchCfj5
aA3iW9X1IMMkJsxOKoRSEG0J1WP8F2opbrMaO8ufPl8Fo9zTOlEc7E7XjvWUu5DE
xKHkxGu31ju5tywJKvO8UAGx1TRTCjnm+gEYMiFDwcaZlpcMe7jF/yiw5ZDJDVR/
RZ0SHEgmW76WbHr5FlaU3aW9zfdC5arsairKlOMQ3tL968v78GxRo85sJXQvmCbL
/+MS7OAJGRJz8gYvjaISAu1lldqBtxiZeZVFKIuf7W5eHklbGL2ccMHnEOBWA2ZX
aKpv2aEPzLeuO0rnOzm2jCF0ndMBBfuAmi5e3N5YDrutTA9jAgeI6un1RPBODxYl
49ugIS0qKqiqBy/JXQJzIQDfhBmq4I1XhJFfG6Bx7VfC09rAIiG/Wx5TDs9ieSSt
gyxgqemRB1tqH8xcmOKpcbJJb1fd1FBU9wbxHsDcWGnfOPCF3NaC5aNucIgz7YJL
yrCVEjB70l/A67X6kGhHQGeO50UhgxC+q/vAAfnQuF9eON1c0l8IuxNKgk6XV57t
1BIW0ClOWFJMOvACdUeAgCHvzLoDUTvT0dljxoNVaMi7gkzaJqKCvH/ybD/22n57
uru1TwvIPjWiXhdIrRfVYeTvL6IbMkN7/tPzrUvPmrHstw7sMc6Gd7LXkCf+/Kt8
QBPfjmALDbve8UqVceG9vasXPExxTni77wqfs4d5AM3rVqKL/hbRQnKrFBXqekv5
cvD/wPfOC235qqur8SIaIDxMt1pBwAVL2VMKwIEmPYvBjLnCKUmI/D9toKH4bk9n
DBBo9xdPLyX+ufK0q/wUeWC6R2yvq3jhaHfb2I5plkzlG9eP6YhknnTYlQbwTptW
TWqzsv4TcSNkrZi1xRQzmxqhyQgzYFH6+MRnI2AAD85LhuxLOwu/OZpkbtZkZ511
G+BRnxLj0uPCoj2ZicpMYTXfyfpQqXa1+EahOHaEb6eQdP2sPeXsVr17Gt54Pbrn
627Eb6mocJ/JJd5ijjak6F+eGit4pdAcfVx0X7w8q2rtXwu4EoNa29gKBEePxbW+
w8LkXAevezuIwA5W3saW9EnTU9gwRy/3o4dADEmEIyvPPjSv0/h/o0lsJPiBrfXs
26hvwUFGGb3cAkxX5VeBQQfRoLdrGGBmCMQbSt5zKY4YNN4JpE4+C/ICEEN1nv3i
TmQT85XnNEuhTIfQxzY1LhaKByNHzdbJBZKvvKk0iW9x6uYf9KtHRiIO8DmvSwFc
qG/IZ3f3dGdiCdNPmibLUVDKsfhE9TiWpWhgGx9KvEr6x+exjPMFE2M2Y7RUwy24
ub6uvGkK8fUDh1wir4MibUDWZYcJ7FPQo0Ba9KZB1dtg+oz3ldKKYBLlnGo/F73t
MAeCOn54XQLcp8samt9je2KA8ZzOHQ+vHeoLYYXCzRPXtZnumm606IEDmYI7iBDL
yArO6lhfaFJSKD+uJasmcIep0CsUTRUhKlKu7manpJiGdZwtpsI4JFRU8KlEVGpw
FoE0apa+j2Osst51aJDo0xZ+K8PB0GYLcX7NWKAG6S77lOf7eZNIu56SpgTCd//B
HTr/4glnnJlw+uUok/G+WxYZt6oLGihKavQ/S9aP1so2PdTp6N7fdB2LPjtftbXs
VU2zTWrs8Q1i03JHsix/ytMpX9Yqn89C2vY6reip7SM2zbNLY/um893LL9PRBJ4k
nO64aoHOlS30OZ0PeDIEgO8U1InnKdJGIZK5RgNtE3h+GJKcIb4Kh/3Bx09FPawn
nQRP/C21UuUuSdNwNvkMAvMhYcTgzkoZud9xGc2uTAR8qh1l5G66tuM590FofszU
VTnoU4cxzG+7Tp9pbYlZNPyOe+KG1hMw5zqx9ievs+SK4HIX0QBPKMYCZAxi0eC7
GHaGmh3Csf0/MO12tecCu6rhEAWqKs2UWriEl7ydfdQE/n4YdrgdVOfDFVkJY+QA
bYBsO5WYdJvBvHEmcv/mnQ/5wD5te2sfsgNSh0vYrMDWwIkxjBal7WK6RNGQCLE6
IFilJG+vZcvoP9A65VdLHkovzgW4GOUPTHCFGk/HhrX/NgaqkRlU3Izqk9GnHxLv
JMy88mewA6wUKJNDx2zEMaizdBnE0IRBnly282vcg1sCh/2NMnXrFHaESUwQYJFc
E5ZYXLhoyw915Ce0kuulsXf/MFOR16DqltAEZIlKqf/mGwYE2npCNZAS6S5cg1nn
yvYdVgmvpdQHork+lvnf2otVtNfBNcq8ZX/MO/n15L9lVL9Riq2nT9LIXeMVXfKn
W9NqD6hwVxySiuTKq5rsU91BafAEgvk7a8Telru2qDIO+QsjZNNHwPcBeYXow9Wc
EGGz29scSleDfSGiK6fQZhwHksGTdttt6YcEx7RoZfE1a83w+JhxVpgHEg0eni0T
W6XSCDyrvcv58caIAHi80LPx4JW3UuONZBDEke1i/BLw7TQFUXQtLEfUP/wYcZTq
MzaUWNkHQy1TUvvLyHpHjSri/enRwjlHtSS1EGhrYHGXCjl9YtAdhDU3QtiBTt5F
RCMbc2Y4u5b5uWuvg3NPbjTIcoADhAFzNunMShHTL2+fx1oz/YbfHHBCBXgl3Hcj
MkxB3aoIrX6Cm4AnLCcreQ8obu6/ge9SZnI7qCGt/VLA5bhBLPlaJn/+X3/wcN0+
z0qVyEbkU6DB58S3pd0v3mS66to70yEbsLH+e/jNeU7SRq1bAuLLCt6TCnqg8Q3V
tOOG7kmBFISKyEekoxy1HphtI6uzmZBGoSyrBj9nBuWjpH1LiguGAeyZfE2k8RYo
3c+gISAVec5JfApk9raV/lOJRwu8av01z2x/B0bZIjL3KT7Se4nZeUipMLZWqJwD
Awba7T7AuaEaxfYY7GOzUZSzEPxNwp4GsdineQ3adlPKT1RZFpnZNbv+Jdw6UhmM
t+PKTh8BicbqzX0ZA2ofQthO0qaK2YtRoxhckWUFRKZzeFZGxYjxL38fpfc/KdEI
SNatKSfdkXhQ4QxBfpvHYQVrpeUKYtCKEusQr5MhB9JqYuiMU5MC6JPdwjYT+3S0
aOtc2mlgsCx5DB+Cm0aLmfa71m2f5YVqbK6mYJXSiMOp+DNPfaIg3AdjZwpCBU1i
dzAbxi4/ogrdbZ6paakgVDApAXszQIR2fFP6xmFL816oLUVPgOHbrwoHpiTR8C+z
dWPsRAf8rNnOo2f5Mxa6jXtAbx3zrcZKsqa8Ms9C88Pg9YS7bA8EfGwtXOBRyNzw
ivQP7KqnX4ad5meRNJqcWq3InOjkJ7b/ON1LY2qj4PE=
`protect END_PROTECTED
