`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4e5YlyrqLT3B5Yi1/q3VfRLcuYDvJ6m6ChNsKm7Q7BHS20uYA3KJBs07yI4YhaxI
zoTMaeJBVLdPcD2gTonAID3S5a3KP/t4REuLOdbluqi7bxIMtwk4kAIdf8mUmAet
sPZA7tzXE8HH1v9C6hZrESzj4xCKbhRztnMAd0192Xb3Vc7D/EWdha0VR3CRFwDf
zQY0LabSgHj9oMmcOqtALWSjzIF067kv8Lg7NVZ98t1V7ATiKNy7o5x6HY22vZf7
FOkX7ztae1Ql/3oAK51JSAXS7zom9CVU4y7jOpH2Jvw392pYE7SV1swvbOTmNPnZ
7E44wE3yRWb85UoI3Fa5ZiwFGypnAww/Y+y70RdsmXOB9fFOuyw5KCflGfpt4Hgv
`protect END_PROTECTED
