`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpNKZbB7sNXQrU5xXGC1lnMhTH5fuD5A8kq3BgSVmdMgiZ4GNDLCMhs9kDjxXYgf
Bu1wNbKkwdHz7bbTfA29l8asm9Lam5+OVt6TG3f2/gaI/GraowHmuCqKwcnVTJoV
nheRJfzragWH/ry4IehZxckTO1rVqhz8FY93DyU9u4Qe6uPUfOaBS4zh+BAeb4k0
/MWvB/mRK8FN+2+O4Sm1LLTrmLEYDmQ9x9AHvnnCyf270c1RYiDEn7CKKHw7vLMM
J2gapc4x85+OlftEAZ5moSwi4rY/Z00x+mYPxQqjJP9KjFAlognAicH5Ts3bJn7m
t1/GtvxFCmEPmNUxpz5IrO9rID4/ah/qba210UT3/H7b822WyuB5pGuvx+3+jLH6
yw4iDNjCp9cv+ktZQoNra+5q3YvQ8o3KWG4BWhizG9FKfDeWr+tOja9TBTElXW44
N0CRgJrCPic31PKg2/dFQXyLYQlcpdn/rhTCgXAR5JPSEVfVNJNZeocdtw3Se8BH
oSMnXWSG6Qsw7uhKrWkywG+r99WuOn2sYXz8yqeNqyAKfNd7z/T+RhyYlvijlUQ+
ya1fRMAJ6dZ9nut+ZnvXZ4MLvjdjQynikAx4PwbgV4edRTGRs1G/brbovY4yzm+i
fNbrfVSvUP9P7jj4l12IkSVqZTdvIKGKd2wxVYVM/aBvvXFE4ypfcl8ba2XYiOcv
`protect END_PROTECTED
