`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8u+998rgm4lyv40VKab5EY+bxxpLHLW4L0Jvf2ByXvT4E8M0NThmJCNUS8jlWKEW
MlFxvVRKMM5I9VBPe+CQAzr1N9SCJdZZIK/1s/yS96uhDZIJdXwTu2QmuCLMeB7G
vzg6xkYOkTKuIIA7DdeV2m0A+tfIs6siNOMiHa6pqfz5kmY2ommVTcfflFh/Tt+s
d6awT15dDS7PDfzEbXGeargxNCcIRn7+716JhYcEPIKx2BwUrhVrzafrxuarIBEd
nL4dasW9pZ2I3Py6qoXtT/1JfTWC/zPusb2iGVj1oYN8e89Pm72TxYgK3Uzw1YeM
woEfGIQXYYtToHaFNAYqIkS36IeOwQpgYIZUuIYSlY3g51XPdS7raJiGm2dWiZTo
9f4JXBWLnwyNejrhu1jdt1QFF6FEaMr0a8DviGDr0WnAu+ohWDbK23pNuCTkRFhM
FGdLGomp09Rak9tp3+aS5hgm3y/QZZMxqWy0cfNXlbvLyHDVugHsl//+TV3Q2IuQ
2lv6cTzrvAjCZDYDSkMWgzlm/Ql9kcueJMappUPO+ABbSnR57Fw2cVHgOhraLuLY
iN85yYnKL+SZxw+V1b4gcitDqr5gLIWUyKF4AiKaYZGorUKhMbIctpvaeNtVray0
j/6zFQv/UunVRxltYXizUykIt0AJ28kIFbcofFMIAS8UHE/nfV/zNd7AyYSuIaVE
vX+b+Vmhbxo3885t9QC4DCXsSW36vUGB53PnzEQBuUcMrowOuY6VBfCN7SkCFAbt
KQhXfwlmEK3vJ5iFsWvCk5l9g4AqdynIx3XnMdGHUq7actEeIMWimdKomfowKscI
K38MGdtpN7YFInFgc0Kp6Bfubue7hXx43tCwi87VD1do0PknHJhmwH0/NQVrC5++
3A0uMMSG76axLcDh1y5aK7Kk6YwCvZNt6jRYcjODneQJgeikSbfH9v7Z/eGPbRKQ
54r47aYhXjsuh2PxOupyPdPoIRWsC6VLgYrlPHc6Hg/2GS3PiQJNmjIaz9uWZG7T
l/HtAj38d4JxzA0PrDzcqLfA6k6fWCRDJcyPMrTfy6kU8C7JIjsmxUYsUYaLZygj
5Z6FeE0XFVV11PAYU3Pwf9ID7+FCFXZ/Nx312bF/0XiRWAET7DdAwBlzXgaa/ZR+
PNlBH9eBYRadIv3fd/BWVC8KHIdvyRqSmPlDaCU8y/hwCRsBGwJ2MRO1lmA2j4MX
GkQnFPsBzREeJYqmHxzNseOmLtpmOZ+/wm9w2IE6pv7OC/FQsdY8guAZOi+z2vZi
imfwnJaCMaSUbBtcPG6BA+0QcrhsRUlKnJF5zNFCslaG1KYfa86QY7cLkJpemI5V
Ysy+cBGMuS/Iy4Kjx7CfLoOp8VwdKOxVku7nDo5sy+K4jv5B711mPQ65mxKLhJkK
njqHirrl2vuAootV8Ut2JuLEWjMnH1M6RLFBtESnjXB/7+J6Tbo7lPn4IfjYGvdE
OULOcli3rAJviBSoWQrTVKuQu1g+ZlfXbQ8sFIaGKhrrBVsTgw/gWX9enVHR72nc
kiaV9jhM+H/0v5P0fWykxw==
`protect END_PROTECTED
