`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3ZJYkuyNoGXNdV1AUBvyTiJ4NdRSTKxGRuoXD5Ub11BeuX36ZaPMSbUUO5V5wrd
+IuM6Fa6k3HhSQ/DfFAg7TnuWc8l6AQoT8W30b5G1N4tttXcA9o2pMwk+1JQsdYE
H4Z0woI0FwO3baXYSTd4ieGQelvhlnL+hPJvF+ffyEilKGBvUvMfJ5o8j0Mhqkp4
+sjfopJZVklEDi3wO1HirYgWbv/e/abBmWI2oDY9OcAs2D63lgCD+i+Z0aYUDl13
hJL9kP9nXImU69h++DKk3vDyy3WJVbdLO7BKToTGYA1dO0F93HV4S1bViwfXRJ5t
/mxll0l84PDKLVaENVDsfZvLW9xD7ErP+fDpMk2r3xoh1Gq+D4lHS72NsxhGFNEc
cc0faqn5sun/CpKjzOKDt2yx9m14P8AG+covF12V6GWe61D/Yq9sw8oDgn4j1GfB
Jzo+AZ0bQN/KwmOdsmXTEqnLe8Fqu4xeZLUzQtcNB/yi3DtDq2lvyqVDQFPoid5w
kj+drr/JU2oWFNQN6tKNxouYc50C1/aKUo8cbc+hvCru6+70P+H2uROWAw9V9COI
WJWfZ+Vxz6F/4FgJf0YYxeOvJu4P8lf+n4Rhkpf/3ehOUuK2cvKBxRfa6A8rTsX0
reAwBZB5C21B7hWQ6B1kh69RTQvqoROzyyLapALmzUXvUZ1mPT8jrbZkU5MnDML9
hO0rk6O2EJtKEIcTKQ1jVAozJmW3Ulh3ayKna8gLIJov0+mWfZ6yoSbGxyiGuQNR
AiY1fwou2MM7dtn6EOCNvXChN5ctt1BYKFaBLSTzQSj5j2nBPrEIiSBkdAGGu9jO
a6xcuvz8UfU6d26Z7JQATu0+zyG+dppXAVVuZqCDqBTlUatGADIjYhbtRRvkSz16
N62+dt5w74fX3TEBjgKGlZubKhZemaHGYL+4Ms0SaqLTavYWGsGKj4S4UciW35WY
djVQVIVgLWfyyW3xQkjnzyCZF6ljezJo2wWTEhqfPu70tO25dDPMzCV1bKhkNFqm
dFrR9v6Wt0EQ83NAGRbFp0Hjri+73kE7c+HWoP8aGv9wDpPH2HJQNkDlDddL8oRD
lyv2fX/jyhfckhP7/+nzwC+1xpJwkwb1vE/7+lEqSnnpHH6p3RjL8oMfXVGCexjS
7QMc1ShQiSbgIuLCgF2/5xfcKzSnVQvlIHC3i9LjkMvpdDLwl8fmjf61C9/B69JR
zcdkye94DZrvBW91vvFpVlgntkvmQccyt1io6yfXy1Mv97MbXq7/LQGyEgRQtkFl
kUbfIHnc2yAD8OIv6+PUOPTDFseo58pq+ACUOTlFigQLSUir2enNNK+2U165TQcg
334WDADLX+JMjbU9wFSUO0U4xPn6xcLwub59gFTrzOiDuOcr4PpjJ4sjnJbHuh1T
UuLV52IErHHsLG/ERzzUDsYeYnj7GxzbCD0s/4PKXJ8SLwfwgal74uWUR58+9+x0
qGtsUG4dZuWZLlChxpFDFGakEll0az/LQeUnEbOKbbmtmwOEf3FptVQJFgykaMBa
QLlOWG8ZoUjh7aBMZcBS6NwFwCJ2f4tACkgmzVY3DjjuHiwb4kmUryqUmA6Zi+zP
9mZ9iJZ8hB3CbFHc5Pas3nNHC9Fh6F2YRBG2Y0d8Gm9i50xXGnDJoxxqXtx34VRE
rm3OwxXI8HQErqL5gjO/Kx4orvWkKof3+86XG7O3Ao6EnCnH/gjZfFwSj5TGj5Eu
CYDgpQNrMBSCRq8mk0o4OwppIUqrTLJAMoqn/R/VdIYIO737BPDHG0caZlECXdMq
KEvRjlRjhacs3ba4QxWMMgrMJT2jeMi3xXtE8FU5WHQrb+bnAzRhdgO07voR980A
wf6KlcrnqpbwHIpFlBFc1PKwy6U34JXqfhL9N87kUAA3uvVIE0q/B41ja2AoamFi
aHiWJ4G1KnFkOYLz6If4/nqllSZZ4wjlKVi0/EnRLjYCXThIIAz4ilFz4R3MH+7g
UXPCxKyf3CrpcVtv2M3cYaHEWBiN5qbNKXVS1qO5gKHX93ImKLD9HpNcwjInXORB
RmPZ+t0SxGAjQ9TsVRU1MnuTGPhZD1wut+ow+jBfsED/WMrjT8CahaR/Ci9++dBG
02uyu7gUnx4zYSmlIrmjDvOpggzxuDInAwf2GuqXZ9NdRDay14SmwN+S6bXOZqlY
Zsz4pdCvG5KDDiyFv7itO84C+ji3jsamZb8/laPZ7b3+serceO409DO+0FDLvPer
s5spVPi3t21Z9BxzAGZT+PIupqBL6bih65iabwFAFWMRud7c75wCdBg3zClvXOwB
Pn0TFrtURLEVzMwURBou5tCAfNpPXRb6sc3Fa3H1bb48Ki1jF9UZS5wVH1IexqyU
IFwB48oGDKmFhIx/W1U1eU87HpMt11uiKgJCHYgUMCYERYmUmvFmAGptvIfgt0Io
P2yl9s9LwWVATm4gwXJojdBajzB1tqojt2fJpM8Wdeia/7WgTseKnNgCyE9qmFqk
kgoe7qJLZS+pKe7f0QTM/CLMmwpp6FTSvmeLfAQvsLNkhA+/uH1oM+YuSpKzGECk
lVMMlCTMxfORfqmgPAh2/hxUWh5hE40/EysvVLyfgYCg1DH459uny0iRkyw6o/Rw
cJlJ41oGGrBc4Gv7s+9eun6kaQ9SUu5W4X07supTFQGAL28+QOUZ/vRxlxaaUZzs
BmwyZcNgTx84fm015xGV986Jdx6bNEMQwWhvfwFJDnoKP9tQn0+WiMYba7/rqnnF
KrppB4vHwY2oGwKqijMxQb7PdUwvE4T6k3wNpKg1822GYSLFakkZUMzYyyHTjCI3
bSTXtsxdrjLI7FW5AtzHzErmEd+6qtzofOwTJgdRpxLEpOF+CAyNM7DXjr6TZBeo
iL8Hh/GRM32aBGMEGkXV5EC4enXUuDsBftwUE/X+7BmlRuiTkx1Op25KAAeyB3/Y
KXMx9dNSDdxNpQU1KPbMHYj7KFwZP4GOWsib81Ptc53izvkfvTkKdG9X0QuO0CD/
dhTQluoHHYrjo/OCmK2h6lJJVy2ggNN1V+z6f6xAR4XvT6GUMazvksfsu5jho1pu
vFtqH+b+5MqapHmuE/38hyRqV+7bqTypkjkVfxwUBp2MM7xAdCuNGRbs4R+lAOWd
0a3Q9Pihxmy6xIQRRovkb1HwXV8JVHP3YjSntlh4+gP1t0GNaMDjxtwQ5TC4M3ue
nU2lPwdGpdC5Z69z9knBTkvax5BgXxLC03SP5mepCVo6UVVRzcNT+F8rFZKoHdN5
Az8AsDOffKSlpmN7Qb2LuCRNUmDcU5y2oUFWvZNW55OxfVkTW0UgE7s3JUkl/fj8
y4RNQcGApyeCb8K4qAVKDTY6TL0D5uOd93IHgK1UEEOTdXXfQOzW6yEqu+f35ViN
1c51h37QXoIKrMfaXEij+xcXiFBJ+Cg2QQJUp1UB89BYw6FZocuLR+JNHq32Fdma
6ZS+FTMgAugsggvH1j9XJd4AHgHst2uxoYafyrbem9ilPbYz1Y06/i3ng4U5Q/y9
W0qAavROYrmec9EMDqENM/QqPRBPkFBHqsAZyESfKt/ljlIbGOnfwIDcBPyg1lBU
aBQqGHJkJ3RCtaZxuLMGq7Bxx8hzpsTXOKqpSD4C84TcH+ORXMyY1ifaP/iBlpQZ
61nx4ZlZrgN4YwC/EwrK5t1icU6HqRtJd6SmQzm9Lm4BCVvXZevQdk5LnAzU3QKj
+RWWRYs5N0dS6+dTVv0x6JMDdEdezNu0x36OAqsOac9+MqKwwpWhfTWcQs+NNyIY
2gtbr/8BO5iBAJQem19Z8ddaOOWaFy06RenFX5BibmnuuvDG4JYegcV7Sk0oNIN2
7O9s0DWnpj8H1maxZQ29cj1hKbwuRGhNvGrQAWYWPq+lyZsX3BxzCp7KYikydaUJ
d43s+S8OjRxhqf86jEW5NNFmBRXuISbW4nfBCzkaciHL61MMTWhvSPOAPw3xw48C
sx5cnif5v49TrNZx0eqabc/LpJPTq07tMpj2/EmzOFk=
`protect END_PROTECTED
