`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3iVppwy29TrxUkWGTRgq53mtStv80jCiRSFDE1mWoWhxMoLPg7zuHtv23HNGfar
AUVptfR3nzMfLFzDOukY6t9SKACFj4BdZDaKt1GNlYU2qmH59oQztZMl5f/wxO78
3DKHSHluEXsXvYkLdOiVh/gSQi+bq6dcik+Sjl17TKLZR7po3cQqe7LZsQG+rQHP
s/VsqKHTjEDf92mCGG+ovyqE2+1RF0gxM7QCmqEMCy3tnDx8ZZvE2ugqYNcxL3TR
TJWTwH21wqiYCp1zL+AqPEFS7EAU3KQbPs7ZjW0WntirYXXh/KLCjMDn04+O+uhf
7klwO9iqqgISK8JaY1MVl+r1iPNgJlUltkrEG85QBEfd/e6+Ir0rZEd6qXIqeiJX
eNa6wmIkmxSwIUDNBON1I7FUF/RFSmglHUTOiT9EYXnhrBNe48JfCPk+9/flH9zj
4DmygOeqc49t8f/fU89Uk5abUQ8mkfzmX6Cnp+CTT58=
`protect END_PROTECTED
