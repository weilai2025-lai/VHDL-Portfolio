`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GnI+OP2LhPjga8kqza3dmg8SF2K2HM0mEkGzbjVYmm3+qcp/ATy4JGs5fLJK4dBC
aU5pWkiqc0etRzMx4Wh5SjdGYEKZJRUaoAdc+OUabe+YvPfokVtLgZUNp4Qc5Ixu
ssu4XZJIoeX+eoe5leJY22zjxpf47W6VkL540JB7b7t9CYi0PNYzz8yuCdd068I6
kjX8SJGL8E4Dj37GpSyO//Y0ElvLObNq1PTpGFF08bLGvaScoC1pqH5xDe0SJ256
w0yixTRbF3/lnDPbXKiKDXhtJJTIEMR/5YoikoIPJN0LKERS+PvCiLHvMs7+1xKb
uQAT6o2B7W02T3kvWSeGKYP4rOA15YAPSmROnreJ8c6/W95BAVQvHSdcTJe+Fc5U
buwMPwUb9pkpiN1t7aEpx+kSInHdS+taYTtmv0IQc7aQgiuUz9swQ2wyWzKKENYw
sX5Z3ndt9bX9XaWVq6r6pUFgPVcmvEq/q8KIzvc4dlnBhT6v/6R5xO5iGN1yDFRQ
lTGIDgNB/5wyWvVnZhH6yktYEk0bRddamcpGq2mEAmiLXYXDWyUpM/zkj/lwK5wM
+ZWkeMI4U3OmLwyS8YA9PL40aKcmxRrzahF706FBGETXf6Vk+SmoLqKovNXqYQ6M
EaYRHQKTodKY7sLrmNqN7xZroPFNQB7cTCtPSO7jNXdm1KUMq9oKcltdA23NDJnW
HZ0sWxrx0aFQjtto5TV/p8jcNByd9owF0wCEkaibgiGqQx0Cz4KoOoan8XYnYdTc
2JEnBOsZB05ufUkMmd/r5wbuKavoppY4HZ1D6P6uIt8LE4WQ2sf6AINJ04jOP6sE
75mZhJ+a8qQXw4guS3MHRYMZn2yPT08ak1kYHIVCa4u7fOSXEtAJOe9+x3IlBQl3
FnENoum7LqIWYeh0nR7mcQd25jaGLRHpD2FiA8O04I01QSYmxgBo2UKLbrMpIfAh
UbYlGriMTqlYjgU99YJ6nBqQwVN76TVXm7Tczom2thtepum9Y2ojkdWYBhKeiv5w
JVwMKEq3eWS6H0pCZ+RZPAlc4vIgslsSvf4yRy5HfKUPfJw8gwHcH0fjyAkUXnZh
XJzhdkGkROoNiUzuzU1z7Ch4vneAWiP/SvPRbw8+SbUUuIIDufobMS1k0LOlySAH
6nz9krpAqfb+QsEI0600dGXrzh8xZBPte+UneoZyx2lIfjkOu+USr2BIFtcAXrnu
Jihmrm8rbNxoZjvrO+4Na88JxB5dsDcjPFPlF8Wy/u8a/7qC1ZE7NJZiwQX1Hnua
3U54BmMTuX8DnqS1jaDdwFfyAAQZkVB1TFRt2duchMSkZqIy8hsVNUvHjRyf4cR9
2epygdscBpPIsgtMA1KOT9DAOqnsUKCvkSH9HeS5z6EO9oAjEjkFBJ2SADdDpbGU
nzJW3e8piRpxJoBVNpBnHGSRg1BoK7v+3wUX2rlCde3S5xX0f+BTHmW7lTibaCBc
qDtkYxbCFnvYTTo4B4aoKBREgrXNuiRQuyp1JrkCdg0TPx3AJSVmUVy+gax7LG07
x2/H+7Z5usdK8j3se1u+Q9pbyclAZ48DQKbR4FPunPUyCqrAa6J9MpcRVZ5Lh3wr
3aebarVbrXeWIWkQGL4sIZNwxHEw6wTrQ/1x29D5zwEnJRF3Zp5D3jDEIKfoC963
Ons8Lx8tPwMYO2ho/xqrQivJQtlsHJpuLvUosZWvp0wGHDHVaSx6jFpGqpkh1Ul0
8Cyzeew8sOxNs4txRdmG5cKTjTKx7FyKXgo/pSFDVG9oyZB8YUO0X+Q2YGXIFmwl
EGh85yelBCwznIjK/fMYEPueQ45Aj0F7Ep3/G833lpDnMWbBlG12/YCZ4yWTMKhE
h6HUiMTU3oheydHoDFjojob/c5XX0RkeO8dcvtSOtbqJk5gI5br+3FcX6R/iyrJ2
R7EoZwNRyV2FbEIFqaQbUyz0NRQFkQ3+vv26YfLQ0KkK5sHgiUcN4BQTLX74BWxB
n5IRXhDq2DcXm5PjyBJlQQOlgwkhsIOl2FJGVZGVAB8oNRqeG45j08sfWwCUv4/1
BAxdnMrNyX1Z4Xm96OY2+aMOKmutOwXjj/+y8UC8zcaoEZx1siOMXUqHlL3Tkit9
3SQAFn3ngSjy9BLWc4Z1SQOHYxNfjNRlas4XXjYSrZPSmjLtZR+TYaXqi2h5Pxlp
zuY4ngEsqzePERLrnEV2kQo/hsVxY8qWl5me6IvJGs9OcAHxTWDRsBxJM0wcKnO0
laU4L1kgsBbD5SLWy6/01+WXfv5etTg5mIouDbSqglVjmN/EK9wj9eh4QfBfKFGP
UES7CU4gUH7oqVFMnxkH+7KeHyRc7uQXQZW0Uepzv6yQid4+WDa176e7UWAmzTyj
lAviA8akk/m7GFe3XDF8XYGzAVzuY5W0sle37FMFPRmKSGR7yguNfXhBvzx0u25I
eEIdSzNUb7O2aV1RqmMQ9W+wl/yTt0U8p53q0fPYvrSVqIXUMQ2NwrUOeNCyD4Go
roJ5yjmxt98udG7/22tT4VfuWP1ISLNpxkKnlkPuf3LrcPgYqGJeOnvt0FVZ7d35
/zGR/fPUTikbSAcuC5vcFrFtJ1RAaegn89620OmzlJo=
`protect END_PROTECTED
