`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eTApqFvR5MASdeB/hX7msG9TpD4pSgUc+dOPHluZPrp0TKSNiwTkyc9b+A845nip
G0NVY1dhgvQS/18daoh8WU00Xsuh0vUSZo7MKCzD8RqKyyQxJnJGoxuIiGg0LXn6
wptDOTg7HdWingGn/9Bwbv52g94ZPtkBIyZ44dYgFNzC760vOqhUPdmbg230Yy4w
Rh9t5OMqV16nDo2HRZ4+f7OH1mWo9+cGdXUmUwX29TJ8jQQ42my1cukDNZYo7L+1
CVw/r3ZDIed+BXYMTjKzcpco6pfkA3TVYt3BUabDEaxldUwB36z92BlVyUE4oMHC
XxuHlYf54ndYAcCEqnDcBx7tyzpCx/gAe7Es0UdG4ABpORHRQNMo1uCSl+2FA3lc
3QVImTgyKreY0YqEDXBx16TAgzPyL+QTK431Gm6pL89pr7Xdjcf8k0Bv0fV8G4Ml
WqI/hgQK9lbRO51aW+YgxHG+oV64q4QqoB1zDrhvIJeYIH8SUqBWf2ByPTVWjGGx
cLlRDg/iupuqhngkz5LDSVZ8CTEhZXEjs7wPBxCvvsi15bNb7yAkgAuHUJ3k7d6C
r9Abpn4SD/kMpyfrplgHUi56Rsf1wPCViZeYkGk31wLm/zf5dUw8sSc3w/yf+NqV
TMzPNZ2HfI46o6i0LuWvC+6UmsTaHkdStEBiAs04KbjER+RbD/Rdg2SN8DHgKUH5
Hzibz5kIfNR60yUrTKbLIy1Lri8ArljKYutaKuI8JEQHcSOhm3OzfqWtWPa3VSX9
SNbcs7oGMHYLeQdKL+8dGdhSXSAuOS6aOLKbzUaaSfWHDPbNw3jxwe9oVmMUPW8F
Y/JVsBm6o3IQ0X1pKuSzBVLxZiHN5mvWG7/RCU6HCLWkqyQizzjc1dWtVV1aZe+G
aiLhfqPdwDbkSHA1LkWuysEeHXYYjukmfrXkbLEGPmFf2e2kNsK60F91eqmXg2tX
iJHEVK+ZGnqP3z1NgEqkjcEnCNSo410Di0p+eqfEdJhyOQVIvfGHJFy8OCEcM2HL
3A6oP9SSUZEwwFtrkhgk5VKNj/w4nnj27jZ8Z0CoGtl2uID5vPWCiBMQdT4E86/l
959tvROtONGY9PrBnFiGxr/g8dmGY/+/ZVUtH5nLdVmQwmq0ZYCNppmyYkaqq5ZR
QHUgao5er/+pcVIX600toUIc0Rvkwm+IoktxT+Ca44E2/sYxc5QYXc3WX9Y0wamN
C7VJjo+fOwnm3fyzkwjfHbymHaMG59PQHvPPiQPQkXJ9SBj91YZPg2nEGGN1zoOG
3+ibqC9nF97EOy8o+uxrnCgAr+KSWuDvYPOkydr63cjqk5QaZr/f3Rb1ZnqmzIxN
jUHYU2oUfROjVcA7PzehNPOwp7SgJ5wI2Er/zco3im53+mrlalISr8fIOtLLmZ1A
7bCTfncPGvXx6Q6SP2twXm2FyVLqKcBx5qSN0jPGitXy8Psqy1U4HKRUFCdVwhDz
2ca5A/Czs1zKo6YaL9OViV3PlCYZ49tzS15jRPvieQrJV9tkPC92VsV4u0+Fhg+f
W3YppCTHfGBFyLZtHWV3dCx3tCOptAoGsQWwNqix8LutLczopkkw7ZAYoEKP4KRq
/oScHOVVbrabHslWFWTG2+vQmiV8oN+X3TaS+sq2HLeasFPFvHThq6/ifQHi+lcP
fQFxMe1gcR08oKOiVkNulXt0RmkMkmI6ONEb3bUZouoejS9Ai/UjvlztyOmCUw+Y
4Emo1XEXkNsqE3jAi3RYEZR9VKI54QxpsyuFe2+t62c+5iIKLwWejXRK+N+BYOTY
mp+k5k3olUkwbaBvuGUP/jm6L4z19wluTkGSKJdROnzTaJc5YgASYRPm/k7bIlz5
NUoPNHGcfShjOy4cc7o5YkNrZ4DthvVgEuioV+Nis7mfZPm6TtVZGyRVjKH4p9tN
QCw/T2WtxDI/3vCMfF7aSUcSdWUW1MxIZGul7ObU/x8XSr8n+6OJ++NevwB/tcog
bFTAEZlcYIwOjjb9oUs7wvW1tRJjg0YOskMCN6eeUvGfNPYBAwEm/syANPBFJ6fi
ae+7QA9ESDe2LSO7jXmVyAd5hHmA66lD5JaPOoV9TraeaDBbLMGivJLkMoGJqVzT
KL4rTrq+kyuEBzrzJfhrVbvkp0EPJjTs8EZEGHk5NM4yh0ZIIhSWmVFJpkmQdKE5
UDsa1MEAT4GvZ7VI0w7Zyx82sbWpIQ4JNCocZslFIVL7bGnLOnVbbQCouWDupCq9
dQVuR5gex4Xa7wo7PDCcBSh5tCv3KH2jnP4mn8DU+JMRJV2lhBzO8BCgMCph64TT
29rf4w/Y4Ig7PUtNwzZLDbT4LOCchWAVejrYTyS0IADRHLTlv4ln13P/fQaN87Rm
SaYxj7BUN4kC5lf21gq8PK/EmOYaU8dELJiWUdO1SdO5IfYludy5Fzkxz+qhPm9x
+cjnznFA6LKYDjzokwWZT3ZHgrrVsn+tfmy4U23pqzS5nXtTFXFB+P1U3sNw/zGX
IxtIfjBDMs4IE+4Qq9pCEqmD523WzvdaE3f5Ma9RW8IPKEvlZNAHwZopgqFSy+pL
vGLde3C5tOD5bug1oqyDt+l0MeAZdOeA8uzTm/5sF+J4gx2OcTicI5TFZ5XE+XYX
RG9wHLWtFDfhO9THBqh6+YefAQXEW6XsKeKW8wmt5QZxH5WqI/2ZaEreJYZ3nxnh
GTicEtqCVP7Ns1RVMmJn0c5anh2HTu5RYTtuNlc6jx0HmU6AbyZJFh3gybqAaZzY
U3QVk24WKg9ZfggyMpD0SUaMQOMSPvonOi067jnDjTc/QMna7HebRORU0Nc7/59z
oych1phhtBO8kCg9DYwz7YZahKfC3yQh+Y2qGqAmkvgYK3EgCoVA1RvzHCNqBdu6
kOgyFkU83slFF1+WPL8B0PEunCZo5HMzxipb898LvFTjItFP1nNmGy3+pvSye2dm
iFsIBxcwk2bOxxzKDBRYqjrtxBVt65lZURjeDrqU9QW3C9fD84OJBWiYZV3k674f
GaPge83k9W6RnJmAZBHmInoSANm9Qrd0b2H2DDKIVFWWUonHzS+WJg65Ov78mGSR
mpTG5Mk6tNUv0YhoYcmgFy1OspYa9u685ET6iKeoZTKkqMXrypAZ0W9gbxcwZJ5x
gut4rG2jrI6oTlUCHU+y3ZXkqTvEqPnxiRC9VN0MUzdqp5V/tetUcSKN+1A2HX/o
hNoNLKc4Vd7fn7zc7oBBr+uZJczgNXsApCgaRJb0DauzWHFss3AIjQlMvaESzOXK
TPqaTwdfkBylfRsgY+35cYj7rQCwzCljxFe8VMLV74R2weB+bqoZzeUqa68np1HK
1kHahqxcMjmVQFN7n2+xgkP3+zriFBbKh+nYr4aiaW5T56yqpYfk6+vvZAdn/i/N
7LKQY7T7yyZpTD0P4rtOdSDcMdCxrsk/oMMGlJQaKlyYgVMuW698GVRm0IsGwq9e
LJ01pYRRy4Wmc87G1t4d+fuuDANLuKtZNyy/f/yP5i24dhXdtivqExxaEODUrYwN
RMsZmnsv0fcPfhyKGJVsjFHlLVkoF5elJNVk3zqv8iqRu3x6E8ZHCjQc4QahyoQF
vZ0F7tqx3lxyw/uWnnTfAUUI4Y4SP4nS24O2CA/nRnll8J77bbzghf92j/6beW9n
BgLXfp4AeDpPsosHlYgAmYrkTuLZqQZhaFJOSYLg/bQqW9h7deawH2XN6FaT4L30
LIet2XdcBuDFm4jCStgUc96UDx60BfLc9/Jsq7vvT2mrKzY8EQc2WkVP4tF6UDan
RSu2Z0fusxtCZ6gZ7io9nYQpa8WX89lyIIYFZ//v89BehhHwq3JikjCaTSktpaJe
f64pcgSrNGtN9YWnyL8i2f6Zt+M2aC0LYf3vHyE3FCn0NbuPE+0Z5UtQHaoR1xqR
dQhHA5onKRiLcFgsuS8m1mkJynzaRgNUNvCJAwA671MwYdJV3O760iiApsUtUy2x
a30jdf5I/IZuR7h8mtIGnv1dS+k9F28IBoCjoeG8KZAXWH6tP7YI+l1nP078nOLa
/XvJTgumekxleX9Hd1b6D/bllCfo83KXzE28prq3mO9252+tFJbvz8N/Y3UJk4vy
lTU6bdEad3PGE7r0V01CqUjXzlG8at2guTvcAUg2BtOJszrs2UddE1asEdutuTVm
LH17nFT9Zkf9fs2TAzeHLLubykwTgYJtfEh/Q3N1iMJP/n4SakoW08vBA1e6SEhh
wa2jXNaIdjAxKUOSbrA9eFyto7OliPqHjoMzdVSAnKXyqETyaqQtzvwlz5fw3umC
8w9w98wzshGWSF+INcWkMso3jq31fcBuZxxhlbS2smfeYxNoTXqqucjaP0qqJ7xg
bNFKMO8p62uoEtBZy9Tfv13xEuUIqVXtELh+IKAGXXqoOTA5KGdLsB3DgpsetLcl
4IbR+ybjTTEj8IuKtHRoGPecQvgICU+dZvubzdxJ8DV7DEJfpjfOmPMXXNBou/aZ
ZCmOgVWh5zI/sMnwnP9QUJkjqlANOmcd5IncyqYYnP2J/cw+RiUji011sTnyGGD0
KthqDE+ZqTJMRtgwNbhTs8hs3H8buqWY5VSe5tTgCYG7d6shW8j4jO7RhOgvxwY8
TQGJZTjx/dvhnYgcbjOFVHJWPRGbVyk0x1kV+3QCfsaE50VqJA32XC00xPGHJ5Di
gl8DisFMyBwrfAAQMqRthvj4xr9Yahx2hP2cUBdKhnkFo9VxG1/rCC5pOqzm1pgR
Gn5tMHHXncwmSmftBbMj7BeoT4THf8w5LugB5oRPIzIBHpB6SI6f5OIt0EopviWo
a+98p4Cm6DiihRkydV3ehQpwFYgIROy/Y7OpPZRoCxHwtt3TLKW7fPMMIg/mkcOJ
LL41yiVnjwmT0rnbfdC02pwQlAFXUuOI6+bvBL3vyU2j20F9Fkreo6iSA4gz0p+5
Mld21RyitA6uC9a49nY4drjXf2fAUS0HsB8biRftm1mXl07jxNsEw0rv0JZlbEKP
VRJCCcqHGroJ7kKUPCuaM99oYOIbsGERNSQzSkCDeIWTgFdYV66jFB3f+Z0dhZ+R
GP4XpGHp7XF/acJZ5vNqILV7Z/lZ5eqzM8ODS0DTtapE0+r51ldhVusWJr3sci8J
AwwOfggUwpbhi1JPPqjseqMVObGNdPF6cRWOfuFJ2bcLTaeIJRaOA/GfWjHwYYVt
d2+zqaTOivTtfAH4GDkjJiH7zPpVEIFBpaxCmbiey8LGRQ03AwRMrYF7UsMruMU0
0JAQzzCNYFRFswuMJi5PNRETJ5MvDXBZGCkMABtC5RNM4EjCjLIa2owl15Q/aVj9
l7S971QsuFGRK6or2oF8e2e8HG2t/UleitjDve9WGt8+P328TZ9ZPySnJdqDtnkI
h/Ag5+csX85UTj805REEcDkDpBYXdIbPaIn1cLZz0j7hOLNBHOtsCJ5fyPGKOkoy
PUoJesJAPQ6sXutADDTkksmvLaRVBx3YjYrouF3NjC3wWylxIKnitku9bqXvF1KM
2TJbV3dgsqoBdZmhw7njC5lfWERwGYRUAYywOs4+OxvBzxS+chFWIn5tZWqr9gpq
JmhSD9Epj+2yySreXHdGgPgfj/f1pRrBS2OYT/HE9TxGVrAHyty6VWsvgq8I2PkY
nV2YSR+oF2tPx50GrDr6QQked5JerXhWCb0InXsrJibpKZ8S/AB9xMzSZOPXf+Io
XsYrP3XTDRsja2bpImw3WidAy/9OaQE5tYv8zvLV2ASFxFjma+BhtwM0iJq6feC7
r0dt/1gNrQ0mGhvHrLWWyKfVwd+aiX3mXADwZssKYLvpezXmTPEEbxucAyaPscI/
eBB7MlSc5p4GcFet8tMQ8ODHF9imeSYNNF4mwsB/i6QwlDC7p1X5f0m2TEvzH3x2
RomcFnQGJNYgtUeAz1Pga33ViodigIFmhNPyHmoVi5JvpqZOtH2eFYrmS/UeCwS7
/36lTL6zSo2Y8yFqzXgme53SntFWYxzCK9OAxPBgHvGSdcdRXJmbYwgOnnt9s7Dy
fXwDAoZM9XuOA9XjNHW31xUdhlmWKb0jxIvp8woKinVdr7TqoY/sSgnxaZPglV7h
ajBaPUT53ZrAW6s6kv6OUm+om9/PoXOtANmf4ydNU4x3q4/D7/mBtIitSdmW5m80
bmWrKMnBmHZ4NCbvNND2erBzlBf3uq02hEBwm3LM5QnCPSTa12prROtmXtHl4JZr
jmZEDhb3WPOTSaL6JeJfafCqby6MsK8SHmDeY3yFB7i2hB7TR0/i4a3YCrf63ckI
aoZNicj6OFh4JFu/TmdTDwJQ9zG3E0MfXlxMM0JgSVj64+q/ZLfA9Gh6nIHsineZ
hDV27EHAuKPB979wWWbMmjuFSz6E1VFiJocuHT3KQudZIob32Z4CqxxK8f/dzzci
g7eksyB//+ayYsvAn5GXCiKjdiWk36Tt7c8IhTV0RLTSIEmNTwJs2A7T8aufudAv
opOU2WqdL/yUW0fipNxOR2GYLrLuxRGxEUhaBjABzukt80GBekdVXPDnAYzEtSxb
0NJHw0tmbJgVZhwbknWLs0T305RA3s4GxoGmCxGUzvFx+oHARuX0JIMep1b3i9fp
rrd94G88R+y/02xngmxzCTX7aHdKqp4QmqhKarD+31w5+sxl5TD87hITZO+NeoqN
4VDSBRF/+j4uC2UGEB+YXbWIuip7XfMIIxp1mY837KVzkz2Xz+feq1VlTvodocMf
9uc8sceHfL3FTegkpruTwB3/8Xyp63KD3ABcnf5Zw9PPZ84wA0DxFDh1znHSuNGZ
9gGelywUeEB8ZaqeG4oaT4LPt3D3ZH/vU5u2exFjOyZ+HFVBsW1OzDDAcnr3kxrz
SPdLvFGAvSMmr9/oRyr0454xl63GFLFezZm4VVIh8Ik53VeWv/YQb9p/0XzIJvep
74SY8f+Q7Np9mLPCz7VNwgJ1B2CCOkRxIXMVVdCm37TlbOfmcyg2PaiIeoZU2Qq+
gqyBn0U79OJ25iB7/AIeItxPO9Q3cSxQxmu/QQkKPr90VhD7VR8J03+iVOxK1uXn
duaME4SBjqnN7JulRqs/2q8jyywA+mC4hAt5Dfq7RpXxGeDUN3jpPmcPJc7rr+R2
sGEzlaZOTmHSW/RcHelILscytK26WZyhlSgmyLRZqwSsSKUZ+ls63je8+dpMseb6
PtIJUR3eWrUfu92vsFMOgIj0eIU8wAha9s+sdhDaiT2+Aj4yToAltbGSDAOU/q+n
mm3iSyqDlYXhS4IhZ8fGumr5slL1IjWzYKN0nJFcNuqYvWNQ94aZDaPF25U8O2CZ
zvzMEW8yrbI2NqrTwKSUy6VTBBuyQgMIrdykK+ra24K68PkZLBwWbXm4E62ECQrW
1+yFP1lb3Vi0PeUejEQQxY1w9bwFCFT6iWc8vCEG/dsHkxVFZ3Xu6mrtPQbKVYlz
mTee3friKh13OWaq8l5Glrj7uc/tNE4pI+RSbt5+DTYTQr4JWbEVNMdULRhuq01M
eIMI3mg9irWROTJEI+EMHboxyH28+SqI0VAyEaeb/LsXRmJHpVRGzv+kKI3qcm4d
h91BDYs091q50mUC+7uAXwEcnFkJk377ihWsd2rq4F1OgCgPazvrb9PQrrgOL9vG
9vOsRiUvPjomfwLoI0Qchr8d3vuuR+S7h3DXS/g8Ymp+6pynFr/hWj79fjXGdVao
YP/AnY7XeDukQX+Y9HiQoGeCYwW8WJzNxdMcicTaTEtjahGUQ/tjAcQeYK3k46v2
tgiAhlsktm7nuHBlEkzBnFVlhh1Sauxw0XRX+TMjBYrgrx2+qBsp68KhK2buFi8H
ckUMPgjs8l64/7BbsN0HdpoOuzT8aH0a9Uk4v9YxTFPF6M/BQYIn4tRdQived2xJ
aGRvX7gTp0kCs1F4weGHc36mMEFzGmkKbxtHH3MNp3TFIpKThgue3qBg+QL4/0WE
4CL2cDHwKzn15e85aunT9tL0E6oQaeNZLYZDTuLu09kKEDiFTLsWVFgk3Ush34Dn
R7KYn+uSr7ka6J7DYrAIpMPpnjzvjeGPiNAcPtkQDWKvGQz15keKej+GiFTxb7Su
K6MVA+68Kkx7pfEWFE+eOpJCgd2K+BjB4AhsPPj9/AGrzm77048acDKybfmXC6qh
1Xo1XO8FMuDwicEgTzqrc057y5W5OMEQTIp300/ZrH4f/vhD6I11ZGCGcypS5hDU
zLI1yK4apVe+Uos6jZ7Ld1l1Pt40mrEgoowMZhnT+5KyjlsNqzTBdy82kv00g/tm
/qRT0kFN2HMiZ3dB4CtM3O1Mkw66IcMYWUHdOHxOXg0SOZhn38pZEfyhVFCqI3X2
ddMgoOpnEO7c+Uy18fLodlcSE39wa/XWaCipSH8/bcmbzlHC13ZuEPMVULWVa6Ph
x8Prv9mbhJ/5/ehCC9SYZxzfYX7X2Dd6FSvT3WK0VOXirbpgTpBOW7C+iKfD2wp5
oCw3W8ZTpX2n6oK6p/N+8yiACoNtRzAbnNn+WwZNGNR+laHfSUXF6qjrzUsjUGsf
WTPhbeWkEFfAjQ0ywJBLXOthp1MkRhhbUf0V9fUnjhH1qsvGp7U8+oHuJsuzeMde
etOBGhtqoHYhbHDjFHovZ1f2QPPZiCCfiuSl8mmWMEWMWVufMOEpvpkJ6yncgSOk
q6gG+p7ka9XpMcDyIaOopdJEf9neCD24V0+Z0cmn8nwRQOqwbmdEehnK97UAAL/o
tkGyPdCfhWhBVvcd/55RYpejql50d0laCfma3vBMwbXHaPJExtkmT02UG/Vk4E6U
PZW8EdcZDUzdX6yH5q4V5oNyGMAg8qRKEJH8RagpNGUw6TksxgX9dsmFv21ieuIt
PRg4AO39WQK8vAowtPWwbnLeY8ECKMy6ls3iYjSSf8Z41mCGkvmijoVOS8WgISrY
nSdSql95ou38BjJrXDsed/WzyzNGyK+E5h0uoUxK9I9GMrvY1ODev6VdzYm6dF6q
z6+M5jTDaVg+QoU8uSkNu+YRCGzTDELzHgvJ1dLwi85hq+9vhkQzHp4fRpA+Sj62
hkNldLGzUDNGhij0kjADUB78rh4xzy6ZYak9Wwp9/0MGhGu3Sgrw7IvXQaz8Pl+4
WyYmcfaKthXlmjPPy6uRF1rIyclziejNO8+XdcjCQIzMUDl0pwF2zP+utrYMkV3+
os4pNnyrpCMwVA8bhwFze5p18CiJGZPvSjvGuVNfzGT0txPCpHlvLbvomF2uowdC
P9z/PlPiSoL7u5gTXTOuTZ9PXtATmxKP1dFPf1sI3OWU+cZQ7u2v0KZLBXczH2E1
WrXneWGjvXM7+wgY7c067o1AW5N3bnPI3RvrsURBH6SxxMdOnM+iaEJf7R+RsdT8
S8Wr8olY0ubNiuXvlPDzYq1eTEfB6XAyJdaTag6mkzxARM20qrZwmB8pC59m4VfJ
MXh07MW3NU9F+nK+n2zFGiESTW2ieCB039BLWqVfXZH7mwpwTy53+EHlUL/ABicI
HB9LluDiAzNwKxgbspfmFNPkqZcKsVkMKzaYj+3NeRrh0SJmHjns2Q/NUMkKLCcZ
ieERj35DQElDb1n0wPUW/wDsPLurjECorQ6q8/ztywI3nJ5rSrPy0Sw/DTiHPlo2
4o5i/RofWwLuzSNNrzW/8TkfsF0NZYulwX7B0FNO4TccIReEe6ClJthiMd03t8hy
+fZ2Skar9H5jqJh1wxsMHBEVSBHW7SaIAjJ+gJpLpnUva2xoWLE0i86JQMkLzUUf
se4mGYgQ0fw8fQ1NCYUJ+Dz+imra2mZJpalYUAVkSF3Q9VmiBO5LeX2kQTmi7upN
2B51WYKq+kiBMMUmvPUtPxrKwtTt1SxcrPK3qJbaYEdlfkb/oB5eNHtLAtZs2LtI
8HKuCZaUw8qccEWl/RoxpTiYot/K2q5mXA65Ay6uKASam5QHY3zfhDY36jSa6KRf
x+9ZJn5JTVKCivwJOQvtLHSnxHMtP5s9inq3LZWzhYTxiZGlt9wfXuV9cJ7BY8O8
8C2SasKluEZLiTUrIifPDLcRFzw/fPL1nEV7OTEdqfQ62KO8o5epGBg4iALmmYpQ
0B+51oCuCTUu9kp3HfVv61dnH+GPSpI067xtfypGo0b95UcHnhtKUG91XQ8zbU7i
/PefBZ3oeJQKDlm2t4vaj25wuJd/Nkmh683G/0gFHAmUgUpdtyAQNoxb+ANRWUCj
ZFFgIuagllP1yPlG2VkL+On+Jp/1vO7Co8VdaIUjZ6iaZRdy7ogOR5upgAkdX0Hx
ujB2bfVcoGF4T30CEpCbd+VskdKAlRS+ICIXKUtkSkqhmbyaOYO0BaqPIgam5R0S
xUVY8OUfH5WI/ltLtZ1aLme53hLV23KnifCQGAsw24EVc8oQWgNc/q/F4JY54qBq
cyYPqPH5y3J+Z2HP73vdcQqyPSpLij//f/esSjlbMI2t7sTkYJbMJspaMFltN9OE
Uzd0GplNqSzNYgdxZOU9PjzhQFtAc0tMrjjxCX0rczqVupBhcSPvp1OqL62pNOSk
9mgdn194sP2Kj9zzkqLwRPMxq3ktrCTEOmjktDH2Fa9ke82kb+81+pV+UAj4UHtJ
KgRW7G2H9gTYo3eYBK93ep/xir6oyhHShPL0YA29D42jdI2x6MSrk+VTFEgY0dij
6S3E8y8nOKXccMuMOxoMs59F7nGgFpY+FTpHEi6EzilC2osf/fLGCueHkLMJIrVs
uABQ7y30liTVJC8q0VwuRlV68hJ9VuqGV/8N4qsXZgNaSNWcRFWJbQ/eWMKo+pC5
z5dlj7Nj6dJuYONsi1fofW/55Ps6b+//Gi/LNYARhYXN6H7BB9Rp2lZA2CNpBamY
p8mNu1UDReozLEMFz8OedtB+Uj/LIUtM7XaJJUcs8gAINcrMp7uUUkmdyXN62F96
Ib8BPohq8dexsaxyEyfac87znFk+90Jh/ZUQVTeXysPBtdL7PRwKLZ8YdllZBxh1
XnXL7lHKMDvDlwDTmgVfzlVPuVJOlTy8o07oV/cU5A7hebOUHrd8Xj8JKlAzkTyZ
NaTbfOPzivnZnpkx2zd8otqdCXauDbO/Oig0YUeAl9NNKQ+wwDkloMmG4+nKHu8W
WlGC/b7x4mVm3Amt6OOkwWqFVmLJ8bWlCKyiy9/B4YQtRtRPkEeEUg8xNO7HKVV5
D/HUx0KRoQxgoa9V7fe26dcea4Ak/YsUMX56aEQ7TRTtgd52izmPbVVuEmqj9MnH
/vg7q8+0ztmSOI/QobZ7iQXGIfk/fA5wLbLcplSj1Pt6Ea+QQvNhegy2x3qy/Hnl
aHM6bTHRnmQGtBhh5nQWcmySlh2eEwZmvK/8IGKpduRK1ePjhc+yDnX4MwhTj2vW
Cm11EK3bHsThecRYYY5KU2GfXsBie0vnUGIVnUCgmEhoTEqi2o1gJjUmbvzHxiEh
hR/Xh2UXEOSakl/yX8OLx066kiS5YDK59ighuqbsT4srh2jh1o5U0kKN9tRHc81L
h1VUoTNxfGQlWdR7kfVv9njqsQ232uWxPwIdM8iSZfa7VdPptYb9k2v0DbGjYCrg
KyZ0xiAnBzSGPGRO+1zemLe4gF4b/63COJW/rZ2c4qzLe8wlS6KBdUYJNPNLCeVN
ArsoS0TdbkWqf0On3WDYNXh8WRYZB/UsCrjOjMM2oJKCmZ1KiUwL/5xjjSr5Bjgt
XpMmc4LiDL2DI/ewyNZwjs6Y5M7x7wlqgJHw7M0mJb4bDYUjw4FQQxkbdMzLBxQd
mpbn/0d+aHZO+d+nKBSD6q2onhveH5ljFWY0jLxZRQAsN+BuOAKnsa1YSqL4NAJq
90qyuskiumZiXilyy5w4QrMQW6X3n6jzCjN30MRiArQ0UMnxNU5sZbJddedduCtu
eC0nQxUmhi9fbOjwZfaZjAY2PP/wUTuHqpwv20HPQkIcF91cFaDgilybS6QjVZC/
zfL0XRf9hy+dn6SC/BeNNlUDqUXrzkqZ5HQVnzwVfIrOy/uFPKw+fY9NJYO8Wk8P
RsWIGweOlg5r/xNNQvYQGWOWPf2QgyzJdVlNH0Ne0ggIAJeTehjxqAZzvKoUEix/
73jBMNlfwFwY14x2pi3am+2MUM3G10PFJ6wrg1W4gZdugoB1vsXf30JGC4byWfG8
K8mNtVaJEJtFf5K1+2Kcc/zSGJ4p9LPw42/S7A/unPhm5FrFPnh888lUPcrIQcFk
8Qbcxpie02J3BWibYXHPoHIyY6U+l7WU7l0gGcC+/VZJ3IMI8n4MDW7WXjiVjwwg
RS2n52czGN4IUtNp+1rVQlI56LuipCQx4c5WZ+ZxjH83dMjQmWmV7ysqKIA9sZYa
2k+ur5r1p25EkZI2RVTpbaf9974WPvl+bD1fma5AbHQkc5t7aU3ThqASGuBw/aCy
Q9rdYf/EBb1p+E/opH9CiAq7BGwFfzjOODFDREV8h0FWprBhNnPBYT440m4G7nLj
RvQJIPQ87DIFlr6Rep9/3Vmv48B/FghOB+WDhPF+STqM1+zS4IjnSb9Srx5NDhHa
ghuTjjcuorSfFbTvU+Ga9BboWFAeae7YqvtBDXIWGsxQVBi3bDNEbDsibw3C/rSs
Al5/PbvvKS9WvGTLCuSahTDdUBGKCAyzM7Xqgx4kMRQSGMYne5cs/+hl3duTVdOO
H7bnnKh0mHVhRi71fJwuk2LSPMvfx2CHY3v95wNugzsmrlBN79k6tUvAJLB5aYkj
lIkHsbGLo4bQg5xrtmz5QWLuZ0y4tATKUeeCxTtFDaCepqBDdTS5jd5aarwZktI6
VBM/jQw1kLZy1HphLcQl0d0hrulMEJvR737eb8t0vAAQgrH6MqM1WKBpwZ6Y6+ev
FYCxw2Mz9iyRPsPQaZ27NqNNHRQ/raUYqh94+6tHvSEx38ft8dbb0t+UAG8TZhzT
YP/LOgy3Ry0sMetcl3GaZ9GYPZA6UhqySplafS8ZQmhDygZL445huzf80ZIFiLye
90wffYpKIsKGUyUy4pjgfIMefxpNRSRWBpZ2hkZJ0n+jj1VwuIKWK8wiwHKKfkEX
LElWoODPdA45i16yV78IhNvnEvP81yKmZz37y0SZwRnxjBIrYpTh8YR81soXf6ea
p1Wnl6eJjB65Zic5qPly0XrmOVHwZCvkJNn1jAtJCI2ZkP6DidVcqE6gRwXi02rD
IIIzqQdLtzCH2rgLL5tH9XEWlOIinqyDcnGa2gRikuwu/7SlWxIjVAuph14ShqZW
8CfHR6GNB9bpEs9H4SuUC8gKjRC4g0nhkoPjX8WAAdtJXFGqPoZUnlosjch1dR3l
KlxaEqDqoqLAHmMZ+w+AGw7Gn01iF1MfLz8fDjlrv8EP3siMf6AyRu01A1u2wp1B
hTHYH8SQAQOh82iR5yUyHiIBmUUcjaKJ6Lo3rl3nVNXCXTPotmPp982V6qoUtNdB
aMEE5PB6IGLXmpD1Q0n0V6foqoMorlKnRzdDba7Jkkff94SWUAyovUf58G955aWi
7fJ3nPuy7s7CYVQY6c1oyAPo5m3JTsFsWoNzkrf4C1VeNU58nNsKRVgaircmybgK
EKN+067EdUw4X4VN0u2/SPrL+iJk5Y+YpC3Ql8HN7NoZ9Cd5QE1mnmGJiL4mRvg2
NMSYMzUZ21QsVLnEMkC1kk7KjKVrtcV9l9ZR33/POXKX+F1prxLgNoOC4AB9JH+8
OPq3NP1knDujVgzopBYzrz502mWqpzCVU9TWbt3GKCfG9tsrzvyqjRYwh63XX8yG
g5LbyBrfJKqXmzpuoDG5Lh8a+BHRCrxAkD8l7TZVu6bpvrw4bzY+mnUzK1bNjdT8
D5VV2GhY/8ePrTxj/mx+Dmn9khCQcNHBLr2793TDMeQRW1jqHcHHZWFEL9OnEKdp
q7mfqnLwiV+jK6SNR9N+ny+51h4iIuHglbuY9MXq1abhvAO+icqqTcfXJDkdyMXZ
CKmIpyz7NXYDUP1c1yCj2SUIrv4adgBDxi9g6VxdqpSLa0DJUrYgbtcDnNU+01jG
YzlpT5CYDqOOORjRGyf2Ttj5KkHXL6UcBCx56W4AgA7rABhnGjKwFp7+IDkxGPs3
TfYq/F1Yhf88B5pSBv+llfb3tRKgOp0lapliQTsBIRYSpHCAKHG8fepKUR1oe7dS
E7octI35gPz5bdCpFN2ndR/SzIQOTJ0FIVo7jgys3RZ8ZyALEDNdh7UUrXOY3XEA
kzMRwZOw+GuR5CS6wfN0cJMv2kCEKYvsnV0ApiPVBB5cbaMEpCvs2RHIebk5e/Ag
CrZ5Y+2fSgtLogFd0QKyjqaObCOBC0xDShVg9FxwPGZemkDSwJX8PedbDsSHZGko
WF8WYn0N/gUp+6918fNNyCv0rVNCfIQtbPj7gpu92hS8II6DXHXwQusB960uaX7N
2kZntvRkgOkAA6ZeF9+yGoXMY/vleza+l6johsmpTDPFQs85Rs6Ee/6GLdhpmtYL
BmOdhkTdoOvBytMVAuS7itOHMrHQOfx+7VbmYpu131d1sU8lZckUNQ82JdH/rU1C
FgtTZhBl68mtXsEC/KrAmTI49YETedi1uRnfRWbw2td7Fh8rERMnyzYH04ICL03h
JdQAFw5sM9wrhSxnqv8N8yEPowdTO2BHUc6Y52aqpxcoFpp30GzvmVTLlsTmMpsd
K1RyPFl8fb8X9uhd+CUgfYplOeWm8w28Qr4roszdy35Omz12W+JawWUdF+Nbb4VU
tiyBDUW5lJ20vdtdmVqT4yNnKAifjkhJ3VNIqhqvu9Yfqm4yM3ArWs7j/rcatkQW
x4QSCirFcjLIynps1sOGBvse0d8tJK949b+vyKn/PwZ/My1YBY1rCXUWKgdqLUhC
rJ6lJg2q1qR6gTuXVQj0h5EPuKlKX9H/tcCQ/h/6vlBZATD+IqhXYZLI/mZR0kPe
wbdlfvNtNB4a+rLbIjI+JYS/FF4vNMUMquUlrfVK8b/vtaxZt1E/qbdA6wd80iu/
yh4swlspjpFWYWgD0YCrISdWW+4TEJSUK4tX4OQK2ee4dct/j52ezt6kpG+GWy0y
xWIff4faO4tO4PeEbxrbWjCaDCqv1P1XHHNK+skgZO1zFzHutGNUqzf8MjYurHVp
UBqlChZdBBsAw2CjRfgdM+Cmb7h2SF6lTNrZRKGkDfAU5YK3HPQHEUpscNjX8iPe
KqlT2Oa1kRUpySkfknMCkSv8qN9DiM+Wh8CObHHyIYxR1tQ7wOnsHdgLdLKdjt3b
IukyL/ugHFPjft2MiGBB1D8KX70kgjTFcf6AFsE8cBnrH9maNVo0tiJC+fHT/z0H
MpVCvTOetBGT2Ig9HmXJn+Tqd8cHsYMh4kPjw5MFF8pW6VD9NMCjrevJLGQU2jRa
EGmKt9u3A7Fia+YPO3HAq7eLS4zZYjDLsVbv3zqseLlezyA+4dIRU85/L/TufGLd
uqlHTSmv2cSnGP5USnsIwIT3hTLki0ozvFd2yN2m2+3VsMEqFkbIb/oKBSTWGGVM
a+itKmtAD8714Fhi+ererh/02B9tXIRDVQ/UGrIlg1/phlGK6KBOLL6RKWH/pHy1
hclWS5x8mWNUcnCKwLKodMHdr8eJ+c3aa07sfwXxou8RdXMsiap/tI3cpoNQtHyK
55U3wv6i0GpDSvV8a39KXoeq6NeH+fexWm9We1k749b0Ex298SUgtITMT6wAq9Hd
xtIzGpaebfDaLZbWfV9wrS6SqUS4ZsZqCsopeUSZTIRTSS9YMBQmgBpMm45VRmYc
qpLC+hv4FBhWuoSAdD7Jskl0vdX5xqsxY4sHS+LIFhQpfsI+i7N1YlAgUVo1O3gy
G9dxwsv9vyZtpjXBTpaMmw8VYX2n7pf1chXSku0o2LNMH4+DgqsLAZsznz3ICplH
wAx/1QgbvbTuuS7ZFKcvrmtKatYjSFwdmu6UkBzOubrAkgLCwKwnmgd8Gs0rbE3J
a3gz5sELqhPcjQF6sBUEyhWTWLXQj/lHpkoGQ+eM2tk+TbLdidbSgS7PhGU8/noq
kDddhNITilJaRLZDZp/z4xzAnav4Uc/KpZb5MvyvAljyqM/+8l+98DUS4v/4rhXI
roH08g8HcdGHf5RtaigJBfNs8oMnQ3Q1iSx0ffqyOawF2aOAtwt8L/9TT+nE6Ysu
VYyHkMYlAsqvUhk/RutoJK7P5RQfgyuSK2tmTrJwJ4Sc63Lt2J9SzwP0ZQTgbw+H
rCgegfEJ+ZRod9g8drnFkH7RWAaM0cYI+062WLIrH37/bWx4bHdjoBAsHVS5W38q
sE0OojDmrQEjmGaMeODeo2640itx3pih5LQu9oADQFj5pZNo52/+KfX7H+9E3S4s
Eaf24VwM8TujLC4g2iJ2vXvi938o+jaxYwlQBJqTQeFSJwNcPBX8bVqmJUzno4N6
MOF9f5xrD+Gmu1if7Z5faY9wG5baMsbyfIFbZRZ//gzh+d8npGm1/3BsPWjjiGQt
Yy4RdLuXVmtp6bHCKNxbbFiyMnJJ8t4JWVm6r0/5WkbMmU8+CGibJmNdD8m7SnRu
XzKClzmb3z7YWaiK5I8vFJIckOc1kGZgfoZmErdmfmU5Z0H/2785xCW+IXHbE+O7
ScuDxpdHYF1Y8DAWwWgnDZMrr6TldytEilJRS/l39L5I7qSSRbx554fmUG6M/Xsf
tXdItR9Pl2lPLI4QGRc2QCXjqcV4S8VxJgM2PZJvr69tttxor1KV9RZ6vQ5NVeCu
6LLKGzO4PZFXtxr4JqVAd/oZ5owC33oJsxJfTnXqxph0v2F/7/L9nB14IKpM4RJY
wuQ+IToBvEaHIEfHCwqyjsnm2yVwSDNJfS3nbCDq21nQ4vtshv/CnfGmeFuKlGAd
CTFDGLe6y/CKpcFHXHZ4yLa6sYyVv/+ba8oVf+I8OSQMdZjXgFdvl8HgBly1guu4
c2hjbAFU9HomFDctwIiPRmIlT9Ldv08AyiuElXgFm0DqGurx/OgcO0SDMNqCAc7v
y3WKwt4lGFB4fNWHMHGKVorNWE8MNABmXSQlSZUik7d4dobAVsd/E7+/QqnRhzXI
JmV8vyR+eTrdyySXvKFIIrw/3fos3rqHI5VVxFBivCYBO51K+cPOs/35hKG1dkJL
VLiEYm7jZQ667RE8iLUOtvKaS561xtTjPG8Xzn4eJ3QTrwvk5bdjdW6t4/VyHiwY
L51p5rYjpRmgF96Q3CKE2sCTBGXq3Xj4b0R4rxbnXvD1S8SBVneXf9gB4/a9HA1b
GUoEdlyDHfcjXQ9OP72NUXrjFsZu6vmZQGjb92tGbpgaMQBBeT/0Os8DWAkYGaFK
zJBII3GStUy2RaHrSJ3kg7IkEGGS6A7AKB1QeBuMqJKUn+x5tEGDub/khaEMmzYb
FuE+/sClpNJeCPDFoPDbolUAm0J142wcYNys9bTmGavhef5dtSxhg7WhU8UxMahS
JZXXzL7TMW3dyrazUK68yKXLsWy05cc5hkbsacFzvcHliPSfxf8NKamGXpSwoDT7
MtfvUqHAHlvfbNmRcQrEjO7tr+2FaPwLUJNiCHkG+VaJE6a0geUQ+h0iyEMAFxZ+
f2VJLIms0bG1aA4lUXgQ/U9z/EwotUMqKE56dnoGw/cbVuwsX1gxgBhVaxX9ioQv
bz6LkhoWZEyLlqxs2NZS/KRgyTYCGlMiR7V3dK0fbRw3wylrk/FsB1QtaETh5xW+
AusfCJjnPKdTK3V8XOPr+LhrS62UGXur9AAe319fpiaRZsu2dYArLb+CR6pZn/HZ
7AwO+ag/dyvaDk/968kYPuYWQJuSjeN5tfZ60Eyp/KffHDXtQ9kk8eLLZfaShzs5
f+FRkGnqRlZF3OcjmaFPgpO3ncnQ10c1qnSKgeHldLpyn2l3QJU2vWL/bfGzLx6F
17E97nTk9/Nlk6KNqXwofG8yhIfOm722rdWxzYlOsMe/MCq1vU0enfQxl/mQD+ST
7Hf9fuzlrnq7lSyap/an2hlHF5n8rub42Z+5WQuterT4mkFMnIV5JeW7VIVPqDZR
L1Ks1z2nEGiNl/VWsXRf3kJCRbsGLeov8CXDHgbW+5ZQx2idU7A6iiO0WccdhqQP
DlE3ALIo/aK+GY5WLthY98eRg7kJuzDmwE3wkGIY204YAeOpx5rygpq6dnboQ/ha
aMyy//yp4G6vzk6v2vt2m0Fh2U9AJova1gPLMXRvEjuEHRGQZgw+N3sKkJGFqFlU
+u1CFzwi4R+/W1UtuGyLwk0iRX3l40GAN95SMkupixBD3SzgXSst6QSEkAAq/JFE
vrLoQL8qK7/iNrPj8cM5Q/ms+Kz0xVtbicPcVMNejilf4cresKAcoE8oRX8Iw2FA
Lx/7uMnlBoJtxgMKiRcFY8SmcSCs/oNkpds+B2lZatcadZdP/ydIy2oGRM4LFg4r
6kTC5hgnKP6XpzUal4ViEG6h43/tnGQJk3hC/nHJ72GZ6ta+Fx59uMVhW+ztqsaJ
tVMgO+B8khISBHuivsupic4bX1qIKd3dYCUFHR3JuWxiDFfJFYi8OjNnOU1DJAWh
IsK5lJ/Edq3JRXdHQRM9KMOxbBm9LPhF/G9b4cZzSfedHh/rmpoW+Rn9UeHDIqWX
fZSxOCYxDy/JVmen9Nw9ukqOvSi9AZEHDVYsMWrQUdB98+cD1F9huv8N7SNRDIk6
lWfsrqP1CJZdQTD/ou5Z7sTClJiKRSoX82a4Kp5Zs4pPM/6ZCkMvEFcVOvyA5s8O
yEsxa5Tz4UiLGbaWT7IgbvOmV7GotIgZteZKlYIpG/uqqyl3hCgif8jeAjkOydSu
cnTFLA6zHc5sgHX9yc1NCVPTDZ4HSI8Ix7igJwvF7a/X5ljuFJ8ySvYMHkqwVFVa
cSnOT6y9+vjklUaXv/YC5bxS012PUStN/f1nKIGyvNEcCx3+ScIyOaD9ulzME2bT
GGMa+bvy7wVdLYEaAIe+LkoqgUyzIDeRxTzP/apjt5hcaBLnBddnUYJU1a8Ne+ZC
9oJkY7NQc0ifChISN77/ir/qLzDIwTqlOebp/2A4yaT0XBMohEIy64Py+udpuxdO
Kq2TWwloQqHmyWIPYmwDfh+0wzy1UdchTZlamBWOPcWv8w/SPjx4iqRm0gPXeovs
e5vNc725aA5CLBwtxJddaHQ4jFz5bqanD72jGQUkZOTObMTw8yFtmweMyCJKNxbj
fIRs7a2o9dA/uUy/SZwA0pIuUVII9Tlehz8o2L557F18/ZtnqGO7FPEp7i3QIozj
4FWOPTAVUf/CqlXgwoFYdVZM41f3XLqPXtUHsc2tHDpSVzw4XOMAwAk5hD1iBVUl
5kvPGGXbB4VZqBg4JeJD3knL1J8KZkxy2dByuxCq/sDGOV5yXVuoLIdJ7ieTJOpH
G69rOfuvuu+I8PtIUVKLs+i548dpLpDtUUPTVIo/EH9eolpNbjntnAP/8/TdE1+1
inDsvFWZj7McEFhTvqbRG2wvHd6MfIQJO/8UQ+b/QQ+fPWWs2rF0vGrpNLk3BJrw
RDuIVC4kgTtEG276CypyhPWBpT52++0eU1Z//cBnz6RghhyK4b+o2Q8Ns6nBMsiN
7vaKxSzG9ymoYVd0QQifnDsOZyqrlNfONFm+kDDeNMsAEshRuG3gRb0mjtFXO5z+
9Gx4c9WHMtrNVkvJz+8U9TRqD/l9mBRyu7d1bfP2wRPajv3Wpa3bkqLmhu6QX07W
9txcH+LnUNrPxFkC9NpCBKCYZd3eBBJCcpE+BoV/YPRs+LdxfzgCv/qiKfyzmULe
R4MsuPlPs5XIdqCEQDkYOj2JXsOT2Qb4ceCdLlMm75RLcYOty8OhHT60gVGslrfX
URPxDdOh3kqUAiZJM+fhRJoCwbLgZMQtYKYEYfleEdjpKlXAaIeZDYgRxZ1QEpU9
b0lm3jLACSQK2ExyrGvmyFZKReAFFRAAHKDB3lfuneDOAjzBZifgXq7fPslK3xbp
8Cgg5JAlDyr7qQk6tBoofSXXmG9/M86uhBwxIIMrLFlD1gaOXkfF8pnX12WbEdbs
1YHZ10Sv9WAU0NssGNo0+c5U+2dANxUg9CWxagcZtPd64AyRlPhznWbFyXWZTxan
oe5t8XAa5si36kUOPtTn7gYKC/2eFIru6BjgkxWb/tXiomWusQT6zAtD9/xvIpwh
iV1wxpLK5vFEQsEdsyR2IZ0+uSXlDPDQIx3+AVQlOHwGoCbPwj/5I842krvquQXj
5CvvicacPXnSUsZl4T9/g1mHjtXy9HpmzHNFRWeLA0+y95Svya0QXFGCTyL60tzu
Qa/7+QCqDGbfnjwaX6XGOV2CgCsk5DDRkblVDb/tsztB6EHPW2dGgGoVJcFxsKYx
O8WgIObRmpdHULDLAV1sNm0o91HlDTRk7F3v84VfQcOwkR7QUrc5kK0ivPziJB8c
lf70dhInUn25HSPf4NGEjKkklvYTHtJNI0qYKxvCtcAO5u1ytKdUxB8LRqoo9VVe
bM4wc7ubMwV/MifEs2RtE9PuIR4Aj8Z6aheNDVBtN3wgidDuJNuo7phTfmQBBiiO
dneAGglsyJwz+j7gJnqSHJRdDA8g/GKxOzNreXm7BMVD0cgDwJRQA8SFGxB6gYFK
C3mROM7LfcSfxB6S7BM/fajhEeEun2yx8Ka6zahIzzWgkR2Qo2Sq/rELSnUmE8WG
WhBGWqHPp9Nn/mtgZcMPyxvvLreZTPdZgJPS8Cqe15IWd2eINjsaVkhM7SLCrzTc
/sN0h4O9pMgOf7ioHBMQ8v3AHBtyB3y4T1IGZWMKlL008yooLZHCFjWRXIFbhq3K
moVFZj6o/QKB4yQtWwPOF5MQuYAg1+rA2S2eRMbSs5Bg6YOd40+WcBet6g9AlWBQ
NPYXIkQpm6E4BeQionvxgmpmZGqNhhxcaZTnXzY2J8v8csx5jtS0v92VZjGoMjPw
pUjJiJ2actYj29QNoGyxBBZr0bdgy+2y7pkapOrtQlze9W4sd+ErNs62+3Hn5GgJ
wc/kCpDW3Q0k3OllhONwrbqbtQ4N6tM+Fw5nf6WthM7GwRCUH/eczzQpMsTQITwh
cYuZo0zqVpEFP0zXbopaBBk11csA3ukkwvBWNSv4LgMbcL5RO5gS3pdJqMNdfZ1h
ukfDT4FOOiFbOZ5uUfYe4TurTts2nEgGzxma5cRrrZb/Rmqr6G0wAPezk6Nh//d8
QCgHbmjUy58cwvCqRn38harHSXF3xwscZMnQneHWAZb9CHa5JuMcvrSCyUlnDzNT
rIGsuTwdreHF5NhCADsuUpM0r3hfNzfXmCDqw1swJSU/NIVU3tpTMirDfIvNcf92
FlgpTAkVyBlMGGdTlbcUGM3RLC1ofTmlRj4TlwRVb71bKGTC3Q5zfzlshyg8/OsB
d6MTu6CXFTKpP+LtEtMurmbbsU+EK7ttVJlDCpGDP24jf3xrKyP4+yQKHa+oSFYa
qbpSv5AzA0L1+iPiQUu8duWPAJSPAM7Nr65dj3a/4h1gSRpzZEujDkrR0acr0BgF
XgIdLiKyHScd3hE/raDqk4TkZ1bGjucA64khYeEJQnJ1Jf39dfqlH639HRdRZLiL
DYNIcsinFAxOlRVysKWtVa7XZsOlLEBulJBA/vqKC/+Bdx5f8bLJLz0py5v1PII0
bzWa50yb99N01Gn60Q+xckAdf6/l4BCfBuvJH+5gwvrXt7ZXxe1fklrjFpelg3A2
vTTBb01GjjsY3hlFXebKZ5ibqX5mzW1xRoX0p1UzbOpjY3u8HjjjlHcaXeec7r1S
sgVc2nKrGMKvjmmZyv1/B9JhVr5SxkOYWa7B5tP40GWjDWrg/zmGiRW2g0PevqRI
VDrgyRYkVHDFdQVuL4F+I8VVk7A3GO7N0mM2j9OsC6/zrY9jApE79pxtHkEEf4ht
CzHKcX6mJnSH7g0oXzMWr5913CYh4yhotZd7uoRffIYgq4MjpvBW4i72uT1qZXpX
xkiyJ2uvXLctuwC0cjRHxsIV8yhQw7bfsTKrji7pdNS+5qum5KgjN/Mlo/ROuIVv
XLsHWDIl1ksg4msW4VepVlaRvBzhJnQygPDODRXr21TnVMzdo3lgMunBUkXO9bCA
pI2Mm2Cqak+JoZWGdkbu2LnRqmrowh3WabXT9uSMgjOc7hLSmNsRihvSGmI1x12L
cvWZH0Sy76mSdDpDQ8dGEXZdI9/aiRW12EUEr8dR8xhRdMm4Y/YurGU5T0kSuaK5
jdMLBUDwJYG+JySyri7QOikzNoksUT+V1IhAwUB42cFZn+96IiW85Uy60XDK54BE
7QSfRHL0m1372UVMWDmv0cxflYd8ry8UUZQNuVW/AghcMnP9EMRegvQUbnVDA5Mz
Lx9yVXL+jms+Ok6oC9+2HKy1nM+s7fNZWz7oCf3jMKSuQU89BosIa5fvK5GG1H9G
/55En7tuowUCEJ/cyLQntKACwMkSGV/y3QXrn1SjUcBBaFf7PXAp1m7be+EpUMjN
hGoC5PEUVzarlRQ04RnZkBnCP0mxzhWGNvZEWZmndoK4orcVrb9GxYtRSf0USuNv
yh9g7YbcpcVhvByZJO1bnOARqEvpkYhLqx++7GU+5zSeFiWsiXQM97D3EYDeLvi7
JkKD2SH3Bq1sZOK6yZuaj28Rd6h76hWEtXGmo/AHUKZHwM7Vs1r+ZW2emtmaah8T
sG5i4jKcAAoZYZ7DckZvyX64vhHOYwi+TUWtKsmfXIkEMew4ZQObpTC9WjPjSaUY
ffZj7UGrMaPYT6ZIHCZUATA6lBTFjcePqcq0M8VOloDEcf62zfMV1/++nPKwMIVQ
1S/+HXQ40F1PT6YCnmTkw6egqnUep6ms7Eb7vI2LxokB4YdGtPTaUdA53fSE7QOe
Vm9mTd+PEKkXS3Q9L/3/IiBpJ9tbHoGuO5fNnhukseOeND/NYRuf0lJ4E/oc1QOH
fnRxmX/FxJNczLVxZXZO9u1YBoBzRvcaclOHhDvkrWoNeGk45/AX5TGMuBH0Q1B1
MMOv5dtdsgdrP0RaURXzuEoH7sXvTFmFMvSu7YRVAM3QT5PNn1lRYJt4LjqYopMG
UQCgPUJ6NUoqgYnuvcedWLhLJEZdExbpxTNM2q6rCSpnmTT6lhAmq/1VEy/oA3OB
+hUWAuUlMn5YAXYpRdTPVlz/VpCywtTIpIUb+nMU9M1TJoCKO3QQrOxi8CZit8r+
4ll0Jw8mGUbhYIhsXLm0gYKxNAmlNAG2IkX/rWLEzstSXZnBNATePmShGf/3P0D6
4YJgEwoIZuO/uYwu0I4H0ThcmY0UGmhJ47WSXU9Y3RFXC64HVpNy8m7fDLms0Ce3
+dSaW3AJkZi7a+w+uQK8ScMGhN/xI1Qqi/MqnxbrNf/c3cx/FmqWyFUyyYIqCBsr
SbRud4nw5wYdkwUdWiAnLOmGrh+fvm8mBpKMm6SoJxPYrIARRlwVcucK9KRzJhEt
hFS+bXNEuzINHgLvtqRC33RwTpa7CZnqiqUAMZFJLql7LUNsVMVW7M4h5beEz0AX
c/vC5sU211Edo2lTztx6BHMRCdEeJG44C3iLfovaKUWddXyAT3hAFw9heszo7Qe0
Ndit8mUPBu+PfAEhltsVo+hE4yrH1dneW3rgbzeS7US0UIvVWrUtp0reahLbzB81
JwMGG1rGP2eQf9zegXQpDnzmJZacydfPFBNNDcY4dx2D73VZve/skyU7p5J5TDh8
smPAMtYBtyZPJBX10HEzsjn/2hwlci6iW7EEd9NbYo0+F53n+BExeaQ/h/JbV7wn
/vPOvQcI9M+UZS7nLNZdN/eoW9kv11AFq/4S8EUvnF56AUH3rQ7JP/J0ppRGG+H5
0ux0d9EvTfMBLNFZ9OzEOx8bnXdpmXDd+yjtHXCsZ3PiGNluuJYoTGFwZ62u1QME
VCBS0xQV0HuAo6tteLzVdsnPEvp08cgg2G++/I+pev6t6Yx2hJBgVT22CaimA+6I
bqOnhbe7SHl9TWVJMK+2UA2far1j2meWu4BbJ7209m6rg3CZ8G5DDuUeAxFeib+8
E/qC5dRNFPgN4pPvbjJgydiYhhvVLe8lpWplx/on7wctirGCjnajtQ5HtocTNDAs
wNiX55kE4w/9lz0LqYPteMpwDFlpTOtsUus2dlpiLHXPV1MMnSoESJHxotBvrxjP
kLt4XklEqv7V7uim8s5TiiDKBuKsMzCoWeyYdrcrLQW5KRkhqEpP92N9hIx3Y2KR
Vy+kV1fwqEp6ElVDlG/Gr9MDyJnWXASEl/M6aMCuzmIBS4OtELwoG2xJ+I+CHT0Z
qoso2TqyRPk70BGH7G/b7YQpN0hYnOFWwVZ5hiDQEQpcI3r7Akws3bQTevFLcWVl
nP3kJPt+eSISeIjLt87lyy9fJ9gaLsSYqFqvfZk0JE4Htbo8L7O7wbVrLppGk0Ah
9+URALEjidnFiTpWqXxngPYY4rDcLuJHFU/qSFalA33i0OYTUQ2sUuly67avVzNX
jNbOpk/ei2U9Swsq7/x3fMlRWkMk+UD3aqjkBv9zrrXoLzwM8DKQkgozI/JFA85B
DBA+w2j2hJMfDKWNXlb36VYHJRbSj9eb7yzsQUYqVdGkGGr7zl+8GzVh/866znJ+
EZf10Uiw87bN9V0zhxc5esmZ8/e5swR+cHqjh7vSQUd2t4CFKx42kn/Lt7Njg7Fc
uPNG+AVT3h5JLMYfx7RtZpakTH3Mhw6EmtwKmDKdkWawPgn4osNAFZ7tyk4kNFpv
swXubVZss68G2mCDmJreCcA2RUeKR+19Ek+tuXy1lOBt8+8z3L/22AP6jUm1PIpe
ZBoFLtpx6fdrPycnR7EgQLWvwEBrDWMzMg3l0rpuwojl+aTeIP2vA+INOneU4E2g
nbyHQSI3H1FLsXNHu1oieAXU5Rbhr8MnmACN0XnHzTi1WMHpGpjvj5364H85aQ07
6Dh/NZwKPSj5S7rAbDmI/d54ERG2tY+Vbd5ZC14eeZhUHid3gRE3DDRWI4E8Yd5Q
VsjzIbamypi7F0CQtpo66wn4g79rrt3WE+583d5XzOnpUgxccT79UyTiconOB1hq
dsiR0iPBKZ0IBLnlMTwiZypwXWXGXO+qwyRhb6by/bT7WAx+MJuk4rkBNag23WIE
khRQ3L7OSo9/+FUFU2W3NBa0KzNjvRalkZYq1/wOqqRpTfXj5XW5YyYEUmGneNoN
LyT6JLVZbkYgJhllOhHtrDM9oUgpn+AP+QiZItqUcA+Aufq3//iPVeDdUmMMCiwt
VtsLcCmDmeWD2zPABzXX02zn67KgTK9OfjdQPKWOQVyp4cnkexzBzSnRuuTqtcpq
GFeqEaNGfAsK8mA/TGdjZXa9vFWoPYkFCwI5uR4PrcDpDZSmqxhne5MRZDepoRAx
PTfQK1ZuBjE+r1FWCnPBEkrol3fHN+CIEe1sGPFTIRLjyfHkZVMUTLVD44aCkqSF
2fhrZ+NpbPBMMD0phwV8UnLCXO8VANF5gGwXSGjVnoLudjFiBEEViCkLuKGlLOd6
591WUKVqO2ZcMm+2ht1s3TDPCscRYwWN1XwvON4vjFUFxRVO2q0hw2ZfE2okGegN
YDTkEdR+BEfrFpKvTmCsjIZ9TaV89jxzRo/R6d4j+86Pmg5tpL1ij1/A8/LvkYAU
8zXonHSUSxbzh/zX4DQ/OudtvD1kWvq0p8C80PX3Ueq1Djr5EV/S1ISVljZEvAaq
J3UQbFZzY17Yd6J3yXTIaWmBXvOaMWaCIzI6graH4gc+Kzzaxd4vG6W1PtsU5lHc
1ZDswNdxAOIMv+zBd2c/dgdspd7J1ixCvxeAORZxfo+vjQnV02TJcHdNK/vd/N1U
K5RU7z52U709CR5mKb+LXgL/5ef6dz6V6ga8ahryir11jFFn2rK/Y4WNQyQbXL5V
yFeTfn8QO0Ort0HGA3EhxdpbmqAZ47ArTIroWUofZCvewOs0c2VD5KnbIta+2cMd
heIEBHwGt1p65sq5BSr3HMKp/4KbiDMVF/uZCdo++gWbgNFwP9Nb1CmHrESfRdci
gTII3Avy6C2S/RFZnHlIrz9BFo6wCzLweVSDmYnRYm1EOzKOkXkp8ivli6ykjzl/
W5HsLBQ5ydRW9HDX9v5WIrDoRaO2qTQhPy3RFBcdnyG5YDP07Hpq561uVxxZ50Sf
GBsvIqbEOcOYv+NatWm1pTSUPGlHaatqpMJHEOMn4FAWF2qlSnnDdts5Hy/PL8mr
XKUvpR8pFNfUzu4dhEtpjuXnJoNUVWgYMupSM/T1hkxJ6RaDdhN6pio15Zi7lEhR
rzm6JsS+UMdRt41jOAtaImXG1hpw4ZwkMzHjctXFRiQ5WTN9bWcHsAIIt84fyp4e
Oc3sEh7LmwuVhd+3TX9cujGHJiq/C7c8TIde9bu5eC7wCtJMUlXsOVZg1RR53taR
iwnXEDIsHpvwZLYHXaTAlRWv/Bd4TeH550041KcM8o7k3qW1IMSKFqnVCUxW6GbO
r8PYxit5bPuO1SYdgNK8PuktW1Fx5CRbMo2QrLNLcbQmHi0mPo2bqEP40kScSUu/
L/En6Sk3SBoUC+m3JZGiMfIq9W4b36S9yjlzcMJBmo+UB5CPGjXau5j9gf688PY+
q+1H00W1LcIVm0KhNuSGGzA0WzYP0ZW6tZsL228rLYwi2f5aOCoeXVH8zU1dylBJ
M74K8eilXvBm3eOYqPY65rHnMCvne8JTuQ7Insd2/aiX9crUSA41wmqaAqjIRljd
AcVoV9inTwOJCSRFQ+ReV9D0QooE5HWoaWRuThz/EbGyQ7qaKRM6tgRLQ5n9TaK1
qilzk+tULEUVcNwLipd55x1DC4FACJu6woPBVK0iEiB7qkgQAoQOn0wpDIqRWV02
imWumDQDjMjCTt6M2GosjInLeCNk8FGysGMhMrFiGY71NMdq/ylwlhEwamQStW3l
U4UyhEgrlCr+3VGLJHnkL353lkiCcCyAuK765PUlkj6HSK97D48ftTsDirDRDSb7
UXN2yKvBwpWM7/68Gago7RYvzwEXQzPSEwS3donRjQu7gKeVyPhOE6AqbIfWaA4S
gQiZzLeK9+nOK6dYft+Wl8a9vC9BReHpJxWYb5vEpaztbprGlfnAaf4yuQxY28/4
sRJBh2Edpqhda7ZUQ2Jfb9pSjf3pGusXZ0+R8RJLvxq3WFO2qYEhTD2J32GyT3hy
t+Y+CSjDfZbYy2R7QGMd0dRxGp3Iepz0FO0GtYO7l/FprrQY71ppH74Zbv3dDIVM
Xj+GQWtcTAjs8D6t1BqZ8udaMdLeG2sN+akbBQZSvAXWGv1ZbZD+WwFYnJp3BGI1
dy1yDNEY7GMgAgJcjbeQDx8HXw9wzSj08pUD8wEZtwpLdeQiO9tyUj/GpHgBf/Q2
5Kzq/V2XWrYSZXRDipDTYjFWtn4qCZQHnOeSm7TnlOo3RH8+euXFlLBIQNSvW9JQ
wncnahAtWQ5/EOW3Zml8wktw93x1MGXW0jY391djZEaNizLUPXuf+2QyodBw61vZ
kCTjq9itEQ6NjhdryIS0OEGTAt93IIrU+6a3TB7PCwkCuM3uwxdDb8xjwDVKeh3x
15HXinC2UPCgsyGWCGLaECxOdFfyoE4UKoIag1OPKydC7bjj5Q0/66X7cA9+5duL
Jn0DwjrjdkS9o4VkbJXMlz04YkG7B5SrKNyx2JGsoiDh1M+WtrbpeJ0oHB0Rzi6X
yEckr0rsxYUW8qDZE8/7+J4111iPEDEPzNhScusAhJPMn5VO4it8YM0MUikiSFYi
+3RI1IjUY01EPc5cF1gpczbbYZPn3b+uW1ZaIaqC3wbdy3lNmbLGWPvwEd9VNDzc
SnE9aj6iZGB+QSXUtNPY2mKvKL98WkIByalAcePVDVK8BpCnIlXazizNZGxtNbO7
TLed73Tm4WHQaPwwGHBIYzt+44g5v9FTPV00mD/dsfezjiS9gZHeX4v8dQqkzflJ
HHsiiFKVQkrBubxmcYLAnunZ6PrBkMWLoMKZzUf+8LQIa8xUbwKe2JlOFWCK1LqO
te0LZj5BFNBsb3qbPP1ZjLJCMsP6zFfaO+acw4qn6FQ/prbVEkoDhHImYzAqdrod
GZOuDcsS340O6CcqWhLO+ATly9zZPQiYNgwWlWmA7pv+1ex60BeNgeJDdOjkVw5S
kXaSVX4nVKNMkncwIgc4w80fC056sVZKKNPpT2FJT2ePn03VBb+EjIZD1uiEvlQe
23NETUliRDb6U0uTAuiWlQvTnG06EwbF0882R2Av2l7H7AIS1ABZbDDuaTOerf9/
7KFPF6OL4yL/b3plvFh/asXPrZ8aF0ip/NzeOPdshRJ48cKLeMEZ/ldOM2RQW31/
bY3daWsBMOpVZ2CgXhuAXlGP1BiVndAw453T+c0NYbIpEKVjP3Ln8IjeuJCEyqx6
Hceu9IH3ayPmQQue486DNgHRGirVMOG5F0i+w/zXhvXuzx/ZbVv2SXbpS5w+wCQp
bJuYwLa97sd/4ThpxVIxlFJpxlR32bUKCs8Kd6s/yPh5x2PuKxFQQ+OhZAw9MshK
ADrbp3rTx5yrRbybxCCNWDGRx5JrhwlX7LyhSRnjIBtS8ZhmOUDIXd7Y7BkRkRDC
DKJpyQEWryr/nCIhSf8+AcFecOzPScsBlKmah1bLsgSxb5n4J952AXswxrEs6a5P
lOXcUcbtbCEtJBGGJZaSpXU04D18DlfS3n9Wogm0/jQnubUXXRzFdHYADS4tY2c4
RNFaoi9hR2ACfXeUyRcjbcAoKbQBUB9qi+vKlsQlpmmvhxuSw8hxUcI42gjyKpjn
OWogy8CGEtBusga/00zo1Zpbnq0SgXFLuDY9tqe7vgOl6Ba3R/2roRsEzjYk+SC1
xQO1/7mnbDr2VgGrZgoce9iV0BCy9QHgTmoX8pWShQYjbvmEmYadg2QJsc/u2lCQ
5YcTtmbiHQibFS5d4TrOIyU9EFma4PgtqtZfHRJJU1SCKugNV0Xfl+1ttCGCv+ZY
A3yTJE3h1m+zfmdVSKX13SdRxDBR12TFjxm9jd8TXtz5MlooXUngAimt9NTzKuWy
V7qWsdudM8T8qWxybR7M7rBpcH7XimdKmr3wafmVrCE062L4qQJiJcuHRekLCdyZ
5mri7HU41ov854Vc0fXy32IoL3Hpho4P0IyJ6jAINj3u++JXkscUtcnK/9gp/wIq
VpR1SZcfy1cL3Ll9zjpWNiNDBKvavMz0kl+r9tjg4fJEWzt3s5fFTOAyyrE5rlxI
gWdL9QZg+jnCQMOqSBLY8Irobyb3fFfHLEsJKS7Z81WBve84hJxbF3Cu8xxk+HYB
HkW/psJOK+lmfZw672AZMz64HoN17qLYy/Y18D3BzlNakRq1tXc/GorIyoChVM+0
9gguzNDRknxJJTHiV9hhhx5YcjBnuurcPlKw64aivRUoNjPmcGuZfu3jgbaNTeBb
TOGx6NrGyed5z6M8xWfVj3D+43POnlXt9I9JPEnyJYFrJnxpyAkD9I/I+HPgeAhc
j+qPL4k/LaeM97UokwsUrN6hudusBKDZnUpJjnVC5Dnt6Oyxy0jpGE26RTFRhxP6
F06fCpsqlLV5aF3XZYJzMYGuFyxFiUh8x+ZEj/i408u2i2Jo5LS62KEJ/YCIzq+3
WE9PTaEfLPclpCKr7dOGrg4KRX9jvTXjHXRG2y+JIOkV89N2VDDf8drYS9xI+x3G
tS/BwA4b946q5F6L8K7MMK7NMfJnT1Nbr5vfQvqVgsLFi8R0ys9do4fW8M+wg77u
RT9Ue94fdyKsW2yGNgJCIL/nXzF/4yeH8luJRIZ2+sBQy4/MckIgebSLw659p3WC
/HsGWabyzusk1SC1b9KTMnZJtYZCoFZBysBQRUL1WTh12yzpy6tle/NY6cWZMQTc
c+GlNAjR6HIShTloY5zxIn42Z/pzqjTtnvZuLtRjLNWsYvQjeEUX3joXi1iBj6/H
0STLGuzgNdACdwDEPQ0hZSR5ffv3cSWAwQQGKIHpt9Ss2ljDFmbHHyqGxIpuIxcA
I8MFm4uVqJpt7Zs51SDVI55dpB3Tl17Nail3zzP3fWowegCeBbS6sdkl+xW8APe4
F7u25ZOEy+6OrQKQ3uGZyITawmnByu4OpidNxh866lJYzygjhMpoTp3xHUyvOQBN
kyKNqNdFQm1Pux1jhyHxxIYBNfrVW8xIbfUNBKeskDlmcR5e4KyJesbxWYe0qYv+
7AZbC9K+rRSh3u157JIUv9xUw9oRJ6wEwVukwVJJ17rMDov7hBwcjM3eXSO2UHnf
38BxFYxSRSQYW7MCiofObwGGuQwNWIoeVFewTbqSdwEs5CDw4ll1nCG1cQq3nE9l
M+G4l6lfNoSIGcfeI+/Keo1/xNvPHeGpsXgVlD4NVoaZ9iyCgnYdPVLgijLMMpH2
qvz4zQOFdB940DWp1eMeJSd7sgB9jpcBiwXhlBT3mF/UENsNzUiWbghQmt8VYNMX
VyGcEc8kpluS9WO7s2uWeidljYC73W/tTzvwNgMda5+bplsgRitwViaGlbfy/AdQ
1ZqbxMNZgwSv6Bg9CpI7BHpKf3dr+itIzgGEKeD85mJMDTKMUlXIxZNSwpYM5tyK
yJi+r4YWJ/KZKeP4UMjyv3RMCz4Dy/Plqb7W6DO/kY5hz59DtijwHbC5Yo+34Drk
QwxUC0EFHVqbiyJIuSkQJiIzmRCzr86wu155WDUnfzsyao21HN+/BoHSdzKeccXj
AvnsxQQfv2y8XWI6c3kfSLI7YqVhwlONov/vmcONXir2rMdlJNtpcVd8q8XwO2S9
ReXzoohCJ9I+ojZ+NWHOT1CE/lTXdtVe+jCHUkgIDiWsXesGmoFiXSGSKxoBeAIM
guI7HhIre6F/ZaxYS7LYkT4Rx/GI6gJnOWs2P1NWx/rQd0KM0ZvoVveuBzcDbapv
uu6GJdLm0BPUWjuaKRKspJjVrDDKJfVNCJjadFZ+LgB4g4040nZODgKL0xv0Bakp
J1wgc7oCxV8UVeAxSIJ5C1w6LI0mlfXU4x0k/d0dTTiIuSDl8Bxb20Y853KoiR28
KZ2JF/armb8BsMtuI4FeA81hj4UlFcjN+5+grZN8eY+2T2s4eAIA1OpMX9Ci6Pr/
5AqGY3DC1R8YGXg+ZKDbRwsetOceXDwzIrb71kYfN8S7pFCZiaaGkEau+CFaQjil
ELownDisUr8rEcEmjjOCv2jyxoHWyrl88P4YLGdqH8fs+rnxHm0brc9C1YZwLScA
61ITVl8J14FzusjJKfHPebtm/1tvGsPuoMB5wHlqgHYt81Jvf7GE3YwrKKTA5O/A
8i9i2PdKq7sH9Fley9eSzu0Puu4FmW3jbgAvbbi7ZApRX0RDylwCqon4o6gFnNFg
h9dhBCCRyegfmEzgiQvfmEKWPQhj6iO/UP5N5K0Chgai0A+8PYXOV2YplvmGPMk8
m3kVlwZNbuk+e4BVTeYtvKG3t6c5Vpz+vlS6HLlsVWDlzGQxvOd/tCFz5aQyd9/y
PhtZ3h4n6nsCC+afmCkodqtpg+8FPZ4CgGI9/CzShAp8GOgRSk14NeVhB6nMWdb0
uw5cF1+7UFUSczGA5n7l9WRaqpKJxFeRjUqCvImK2jqaMXcEPOFx3nf/aXnZYj+O
lawk4w5ttMlBZ3DU4dzhyBW3w69U3LyFSMQm03h9CrPQSVZj9NGiDER/tzYNAeBI
9rWzvPRDJyBJzuLdtkkovDyd5T+4gkie++wbI4/6qr0JuMfc8AqOgEfgPskGBaRG
BaqnaLFUX3TNs1lwou0e3+jKlM+VHqIdgAKPgiO6Od6lf9nrFHT2eYh9yL2nWgwb
fuIaAbjDEfRZDD0eiLcguwuwIo4eHK7Mw+w0mKMA/lgVMH1TKHhjbsTJtmeH41wY
Y3MOO3AgndvbDXq5N4e78khMSJNtYv7WfdJgh+aKAZ/n9tECsAX504tzmLorYykI
lV2UKSmc2PWf0O5kt3xcdceCz1SGpyaCpNYrLXfrvcFu/VbAoKf4NYvPyd5qwqdz
U6xn/HLYELo3g9fPvlEAGX+VPh52BPbXRa3keDE0804z2bxAVA7k7c6XguL8bT/y
9MGD8yydxFe09p0mjvqxNuDMahMa1Gm1g293doemCDKpY43fNpuGaUR/O9BMffLl
bBUGH9Igt1pEf9OEe04XoPja8qkrSjZEOi8VuEX6MNN5i42pqjthxcLVvyw6FChX
g/UChaxXYJy9zWzdhl1Jmj581xFQ3tUXfb8ULcKEp57Rjjz9F0vvhwfotCMQAr/X
xKRhiP622xshFG2hyiFk3zzbsn1MEO7BgC8Cgt3WgqT04dSUYh/MmS2Ba+FyDKn1
plS63HSMrSHXanHHeGuZK9Da1wEEI7O2ZrjHZnBA57znvz7T7aW/baMrNEvXqpuU
n6VX0zpIPGTA2O9tFsdVdw5Cuk32BfU1Cs4WLoJc8MEY1p9bBhZGKPL3HwP+STCK
U+G+xtHBtuCUBMGRmL9qw9AKYACPyi4H11Hnjb0yoUnsKqOHrDymUKJEXQxD5C2h
0wfB6Wzwdawjx8aQOAxyEE/oyKFjaNu/JsJ4EXbk7T8PWV5wh/+WO6rOcD2iyyqy
O1xX6aPPSPC6Y5Cpcwd34JgmLs8HE+ldgyWWyVKfWGjTezPNErOhaRCNBAt76mcV
G+CWrtumUJztMNF7JmSCT0rfU/2x15RqK4cmXOKRUuqkRZ6bfcODQf5Oq9NyenEv
VJAGfT0lJC1dCxOFT1wVyek7EPRPxKyHbt8ROScsvn6iRq8lZtqlQDdZxJqB61+O
/oTWk0MFQsPKEqlNlSqZrYUHP0tIz6srG2TcTubqvFeVspSmyP6sjpCoF/Ws33RG
Q3Yl644FNtsim+vff2IixJ5MgqpOgVFLDBUTcjSj2EYf6dC4mR2O1ivIHSm8wv59
XVRz04cyz1X0cMXTZkr9CizQwQKmAouuMWSFb1bDScESbRV7XGsKjLK95pyKh2ht
5rXv/l4hpK7dDceMgalYbsL6dYcx502Aw0Ppny7k3gcjxIhylM8muXKE2XkMrEYd
cswO/QWB+SKnPrpneX18AGaxHZY15XpRo/gS1r5PzmENOxMDiKYPmWn0E+8nE5fy
ygM0sGfNVw5JYreDkuxVzKuqG7T8mjYACPvq8BEawF80/BnE90WLL1hhMDiviyBP
p0rKhOILreGQTPGpu1zuvCOI/rTppb2FxZ/zrEryjF+doHAXNcXBk2qceAAFyUzW
yj5SXVfz5zqyeROcgnTcfRitncOSLVqCTRJIf1rxyttf0vUDW0Y0UF4d9YufaJo0
uDp7COZqMMuSxp2M/GRrDfd5KxBhjcMXBjGcl2aLahESzcKvKl0+rjWVYHcu2HE7
v24Fze53O11hDU6V8tfgrjN+FOMUarwYGzlBxI5/p3MeJnbJVbtCcAPIiARQOi0O
1eCfpxeYmeA01zZYgHEMZW2QdQ2BsLg1FOvlbZiD8+pG9oNRYOOvWcoNclAKbRP+
rDQrmyPLoohL9pxp92AH+Y+ca1It5Dw01PdqgJMpmJGO07goLRCgqFdbQUQRpGGA
oEWufY7YUNODz10xChjNlr6kmDVbwnh5NnL0Vf7rP1OTZu4qCpS69+qJYd8x5LRL
+dtFLtMovx6/RYofq34Vun8apcrjCQhfk6vwsYlx9VdHvJGWel0NfNLO9uhYKaib
avN9RWU112mmaLjU8X5Mvx+2TbBRdQwvx8fT5U4L6eWvXfqvXOsCPX5HkrYE95ey
NdW0rfPUku6luD15oAoXfq4cuRxb8SNHRn+ZnggHi9kmsZjt1HoVcSiw7Y6bNX3q
TdHJbbz2oyFh+Ex3whwkZCQrEVLlqHakM4F/l4ZwxLtJa6yRhOX5O2UNSUeO/jjF
zt4hf3Nozhl0wrZX9CLJWRzSdUUGn4MpNmDufe0vuM2XUvCV0wxLZTV8kqIDqNNg
2/t5Ok3BavHVZczBf0w8m06wJJkrZ8e5ccJWmLgK5zuCLcWS0CofHivZOq7ZNcG/
MoYmaYGINdYSvdrL3bOAanGf50PDmYJtInHGIdkGJp3UaPacgw4/MQaBsz67qgLu
uZrGt++52tore5tcdFNa4lK4bY1o+VsJ8Zat8WiS4QwrCvtdgNPDyj78h6ybpOuX
iX0Jcm5c/7L0h/RBkzytrrareU9LKVA2Ab5LzsmpejF44ayDXfMN+sVmn/zuUAey
VtPdFu7RaZEcMIOkJjeh32KGEbT+Q/RqwlUKal3GjWoUm8leUwx3kq25VxXJeiIJ
fMM8gw/pRJ8srnyhZhNPFBEVAciBArOvv5yGb4ihebxPTDWmkXiEKNi15yQmsm0R
M/jfamAzWMeU0LQzTFDANE+JLADEYaKV3hOEqKSCSnON82PAMgeEIPiJw+gQ2bly
mV6wfBRdwqY5BNUdg294B9Z94/wzOFojahtQt+N7jHuvACwo7ZV0f2fsWYbZp4ou
aVypcFb7xwfBxHzR61+IJzQM637ZSu/ZwOaJjXbjHyHuznGbM0ebZlHr7FN003Iu
ZXqa683mxAHqJ/TlLLIsly27+FxHTQ1F86T5UOy0zAdOjouC+nnOAw6TidxJ7J2t
cNctqzlD9wLWZYyct6l2QKlShaRB2twOe8tY/P1lyBca82USQRMIKgjmTfL6zFbF
ayNKxlStc5Bg4UiunkzjUoMuxJd7jLrnFY9UJ2xwyuCXe4qn5P2++zQz12pRexCI
gWuS2YG2zCZUSVOroT6FtBjlvZ7A+JuRhJg4LbZgeRSBTQRcMqvmgTH2D015D4P6
/R8wSF451Mn6/gO1Kpj9UpGuhNoA70GTsrkjFvHqrzWv0xEV+ETNUMrnxbmRCGan
RsSa4r+Vu0rqDDSg5h7gPXPdjphSpqU6ZjiHSWVA83TEmHb1SHgZp5XnMdok0xEm
5ePiTi8TJFYROHk13Ru8IXDdHSoDSWu0VPSiN7Ar5csnFZf6aoNbj4kOUuuIpazu
SAZgZXC28XzWXcsB5QkbrY15agXMcsoPRBQn1IOFC9c1ZS4bgL7u9rlrkeETFJbc
zIVUH5XJFjc4q/HQJJaEZKa2GNXKZPatWB3QTtvqhQ5+BPtDvp9VPJnPH/zWXgm3
saAjhYcDxTkRoVf8Yu1idPS/EW8B+PMN0NGfVENpxkXLW5mBnhoc5UmM7j7fkjH8
2/dGJX7/zbCGuEAjU84yvufFTdngF6R949O1Jus1tZsIyUXZ3ky/7PqNTr30TOtF
vAjZrbV2vyU6F39LUEBxVAOhSJDzMgHE2uE4XU8SJzzkzbtFu7OWFBOKgn0nlVXh
Zroi8ddxSqzmTnZmwFPs6pZ+MJm/l5R/QTG9K+dc9yw3lFaZxzs354F4TKXkIbCD
01CUeHkbkEmVNxct7CYCJhKgmSNrpGzxgfrXmuOYG2ayGQ3j9D6C6nfKzDJ8Z7Hx
xUPjwgjrKL/Aa+c4nqLpAfjixu9+gNtHpvMxjJCOThtJnvjS9ogPdavmcq1Eu2fa
iH57xuTTUCjT8YfOEbO2QL7BYPPO+VeQ27PzOhg7ujth7heEjTZVOfJ5cizF67CP
LsgB9fA3jbRLF3ZWfPBK5feHKmrG9i+QwTq9YoStAmFZtK2J/dmteFwMKIdF8xHK
os3LVPooErCpceSL+EKCbqX69BPFXpsa8SHcnFEbWDjbHr1aecbFIjkPv/Ghbbq9
/mtwBTceTzGiPSe57EKbH0HQjjYT58/y0qz8QajhXwF3kO2BtwjbLHrKvUeecXHq
wRkMLYY45Y8m/02lvu4hGxTm+kZYxKToaCv5CU3MOKypktU5VEVFf5xM0uRanZW6
RV8g4ggu9zbnerLc5vj7LfIr7XImXz92vCcbV3BdTDtWZ9TgmCauaMXpuO5KUVMQ
qLFdZt/IYHts1Tbw5bkt6LrwnUfcBYxEEWQX0H5FAwdx5naadjM1XbiKdxrmTEnv
K5JUKRtgEGR3HGqgKnfQLZ2mwBhYIkeDW0w+/FAoWqOiynYeZvsYuhso6KklDn9R
2ZFFp0ZCo8wRad1IxEIcu9iCiGWmEQy1LqQVi8PKjKf3L9fqRQJXBkcJwD9CdO03
/IASN8oN5nj3msGGyy9nxW6KcZGN9DpPttOsQyqoNXQhpBn+6piw8XY5CjH3KJep
UCAnVHd8Oygcwh+b6ETrKRxx0YTsmB7hFfUsgdCX9Q3WSG2ta6wpuBMKCP477o2G
uUhXplRuNYjmiuCQ4k2CucN31e01S41mIZv+oEHPWt37MtuSKAjtJ8zH4y4+ZBAc
aElvMcCnVAG23kV2rY6FDhGsFJ3YC5hES6sBOT1DitSc2kO8U0ZFDWPMyhVIujRs
giQSi6iTVv7XZLyTijcwiu3g43+OkJZ8ra3uWovdllnVhfAc2X0G7eJrhdllj16E
RNOXnFpjn9v683D6f4bMjmmZlnC07AqIG73Fa43dhgfifi8XWznctu1Mar1oVuCA
CmwjtJJhMzJKGDH6AP5N8nhyPvwj5TDDxceLaWz9hAgwXiv/86fupsJjyE1J7I7p
yfQxTfQfccJTTQ12HC3t/EMAxg5Qqylhbn6kjkoMJkVNMW8XwGWfPw/KSxz6M+Lk
+oVIeyb+zQicnJbfQevnCnVhW6R3HaTdBvdgsEUnszBacY2At9Ho7AP7yeXdoC+F
S0fc2C4qjOCBVq+verrbw+ectpVGgS0jDbXIidH81eH2Y0pCjCendtmQy0vRGQoH
Jj0Lqa0tcJACGxMsgjrFrUAPPjr0MFy9gTYdnwC1ga175OlLwVs8WtdW3SkilWy6
WwOSbBd+Id5KayJ9n8vPRg6dWK99Uyn/WjQqBEJSwGyznxIMc3x95lfsR29jo2DA
Bg069N2+/FpMyhOpnfFPiOfr0/dYyVDyqemCcB2ppR9NH/kTscIjUFg+DcqNZDyf
ToXSywOkYTeJ3cPwpnwzxarEX2EESwZwPrK3Ibzt9zP/AEA+Ya/QOvcrBPPY/O2U
N4AIrKBDsGpvGMX+hDuJEIpxfge1GYLfKZEQBYhgx/ia/QsTjjJu+rq1SmaUSFZ6
2G1wzUy2/O1YqqGGiW4amHq9WF3xBHy7bAGGnI9kc9vFrzOOCwETiYxSc1bsA+pS
cP9fhCrpp+snWDXjmvFyPj9BsOreeupePwb7hto4L9HLzZpg07PjucNO1IkM/3nZ
Pg2cZ274Xrq7+UgTdUTw3LRmAbOqpf5XHjYIvcAibvn2X066WGpYsLEQrE1jC/ir
OkTozZ0rcKFlnPlTEHP9XMEg7bM1hYKjehaRkMoVfU2PUXXQRp3exA9GBzD9JvUw
HcIJojKBrI+dyV7pOfyzNsR7BNawAkH4yJs2mKO4hf/L4X6GDAqj+DG9OSb4HMx7
VMFuOU+jAI91kLyLUnYEl+6EVJTP0/eKQCAwv/7M/nGoaodAGPxHI7tOVNy7MfU1
HpDWPCNm24cH2U7JbTS49y1u/YuMT2bYvaOQyZzFaul4dvw3fvcLDax2HJ/VTLQU
UQPpQQUiV7g0xgvpJDbI28rWd0ycjSPOu57Mu6m5Oc5wZVCUa56fjGrZ9KJH6sSj
MUJdxFegHPRvyut0115c3wPuRu/gifrajBVkB6VK0SZKFHUafEIF8p7PiNWkh3/v
F9F+sk+jHGrJLUQ2QXhfLBt+Wplanvoc3YLnIhA2zL5i/cI4mCihLu3Tem2ArB5K
VqNsUlbSsFQX+1k6H7Cy6I43G3oj0hOcka4Dwo1YpkDZPEhbCIgQpC2tv/Sm4kWx
O3tkJhxtBB6uQfDuD+2cNf9d1TGhOILw+vcmZLrRtHA1b62E/OWrtki2Yv6vZf80
227xi4+Qo7HbTSCxjO4kCbfKNPhZAeguqwesYeV1N3Lg2QfUN7D7Iod5Yed+gjqK
OxZrv/UeQLIBZNvgLZ4SRZjtV5gt1g1b6vUeRVht5PPn3kD4KPuLpZiUSv5ZSvZ1
/RvQYetcwaN6hm7F94VPdlXUkBv9ONB8bDg8CF3ZUvqblqVkrYnvrbSqv1czRFE8
v854YchcoWrdflWCauZ42tjkFiSRTsQsU2czEZ0Bl+G/gHfQgFkN1UAWhorEqhTu
QKX2lr5PGxNDkTgjIeRG0k/p/UJMkStgKr6oQsp5MwlsvB4YVbR5SOQZJTXPSFnh
+yf/zFzWEJgUz5GCqj6rbwL2JPe44XLFgKOYGnLIcxMDsR2ugrnH99TAGlVQU7P/
6lzUCGyrSTmJUA0KcKDT8f5C40y65knG6BMFir5Qb8P5zTvz9FuiFxHojTkTJshc
samVym8Q+njvTxoiC0lz9Dw5hdiaoa6jAD2HIEJI0ZjvzZ0/qAkS5Yw2joB/V6U2
ymHipWfVak8D1xd++Sc+mzfLWMtaVJUdlYrTAl/h/SqLFa6d+iD2EcxWi2Xm4ulF
ctxoI/9eeqLfkGU/t85Ee2RJeKt0tGsiY1UIGYL6QUZnPN3AHU8peO4+YRNeFYof
2bGlEF+qrqk+8kwxWem8KzEcDjhP0UDVwbekjTDykweZANNGeuvABdG+y8sBjcvZ
JFQJAWAZmMPIJJ7kkyv3xMJZrZvucIhiYDETYOcMMvckmFm59EuBuv7lA0oHA7VL
iwR6SQqEECedyNVY0c/j32Lvciq8E8tULlODaa9aAS0pxTIyDSQ9uPbAvgtkYEUj
+7M1+VzHN3c4ZE6LVz25j1NtdpFagYHvMKOyarDPnaZfN3Ri9GvOEZZ90HFepyht
zFNVmnNKpOe2+0VLmbT+RIoeT37CicvqN9ojuKifLdz8nXJ8rwWVuUX4XA5QG5tz
CvhgyZpm7sw+MbIgSZMV7Sbc+v5yM3tVXQIYLwTxb5Izme8WnDWqZ84zi09V3wff
Ffv1AiRChU0e6yFNQWISzkUkomu3NLg/Nxes9ke1wLFdlKVhluD1difMQ2at1YFB
006OfYmxxrgPKfM6H9UpG1DDkSSxJOo2BLSQztVuQMTG1Qs1jmIwfemtTjIVZHm6
/Y6sSvTFAE98M26oaPMbnEi6QQ47Jo6wN9TMaeXik8oAWPyu37fI43M6QlDvoZsf
fGscIN7w4jNLhYJNZT1HXTuJ5hYHxxT4Droxaf0Uwz1sULo+4tVJEk0QrR0QGC1R
qw3ACVGCOYQBSo11MWvXqp8t47xAAyKW8sChU2PPMz6p7Hj10aIdcgc/V1kjdSTX
0ZchFKDb3HuGtNavKzS/kx/rGnKhRwWCS2qQQKiv6Bn0breuFX3lxrJWNgOiECj1
1oWZChLu8g/BLwB4iH15tyc9vL/4YHfsYF8win9wY5jLQe/djM4gDxu9ynC5K2LZ
EwGrkuDEo2KU5CBLFS1sqm9Xba2OY7Z6LlGlO/vFQCROxAilUVkbwiWQLXrzIdR0
rVEQ7MJgaKlH52gN9NnH2Uc9jO7Mev93RjpE1sZtWlu4LIAh4F3qKuZt5fJj0Hxr
jTRFSVvc8vLFdUIoXhtLcDmru9PQPmfkYOdjUIdW5+oRfXzm1SDrrkG42Bde+Q6J
aW6VvksBIwdtiV1jW1aKnIetb+0Y0mNv4axSg7FdONgDvVJDmp4UYAeZkYcVj179
oK4N0JgLrGboa/kTSosdoYQfNNzSks1AdoxBKrDYAH/FP1YKk3LdJOKNqFfhDRw0
l0JmI2PXVhkdH44Hej8qaSQE5WeeJQbDDEYahg7yndhdFrKUiWMfxkHPlGiZ84yT
oqimmhHySMhVKRkfKOYUq0+iE9Jnlipm2C+RQZcFuYSy9q9PU1ykD7Koh3OPSLAs
pXti7GzEubvDHlfvqGlqPlpjQIzkZDBI8yhvs5h+v+ZbzNved/TQcBZ/A2tyL14c
wFC+hlY70QkrywDeKeIMr+vu9O6pXm9bVcL1+GJtJJH5W0GeK4lKghDjE6UpMm54
X6YJwehgcdwUcAVMXnoFGe3xzfyYhTFMqxCCe2+UVmfVBxvjThHENQVUd6KGOsKL
oZhc8xO4Sm6JbNJ+o6Bj6g8/eBNFqJ0DXymNnMrif8FhhKeYEjv194W2mbh6w9XM
lbZGLZ2UWlIf91Obn7DPcG8fmZVUXAX/M8d3vFv2b7D6m6G8EyMiJh/k2YzQtTy8
LnxxvVs7IU23COjuCEG+UxyyPSC5ppXq+PPZt+zhWPX5oKd7vnzbRHe4GTFuv9iB
Mmo6pr7WNI+ZBe5PSQa88IHmGxjuBQAJdpYMSN+8NkqfY6gPOL6qgXdGbDnfnXeK
u9JE3tGQwXUrH8gP+cpshgN1FoFgO3YvV9Cn3eijF1brE1KeRQUczPoCcMQHQMY6
r+oOHV/2k9FGdwrc+GxTWFvHNN2NhUXYq8ZhY1rEL/zeaOSJ0EbOaJ1mb6Hm7FrK
4Jwzi7kqHkB4/tuiG7CVtVvY04S9AeQ7dL1cmjsgtsp8+8RJsFpSxbhl32H8Ww8U
UweJRmDhS8Phf/UjwsBSNwosFYYE6+l1Ed/Ejg0buGFPylvl4Bipk2Hz9zaeVsal
AXHKOuq3DCNFZobmL+06aL8iJyh822B6NPuEYSblVtwedR20nPi42L8AxrPDfcTZ
cjxBycVIn2ya1NEAoGmpBHzb51BDL24G+OJI8pzJAzQZ+SliCRFFNpNfeh8th1wH
DEGGXtQ7n0scoMNQl9cm5aE7lwplzBLYxL1ZBq2t65vu6pma1yGND6uQocaNa42Q
wjSxKCqxzTskmX0RSR4E9/E3iRjTACcu97Qga5pofxoRMv5MoAzDHg2keQpPZmHQ
YwljMj0+YxSkowsu4E6U3qWAmHkVoJ9KwN4PxA5NP2FLaHGIrMPKbH4aPYn5aLjH
UwIvQPj1Y8zaUeCFUbFkTltLPeNWApO1UIFDw0pIM+AlCBVMgeThag+yElvUQ7pR
4+sFspcQOESmZR+r+P/EEhzvBtrjv5pL55M1WknDEYWBlojAdrJfL0j0NKAwwW7x
Jkj/CXemf3FAGykcSXLkeqDXPddJfW8I5QglSLQeAcIjILNLCm8wJwbDvyaXkwLP
miVbCqT7UA61ydramszSsvd2gqOClLU7kXa6xuPQsBOwrA4lO9q0QvHPZBn65NCm
x9y/XzG/l8fUZ7P/bT+1LaOscyXqcQmNvs5uBppLKqebAFLcPZAjezNpbBQoNoqn
DUf5YhcRsOi6C5WjX7aMI0j+amCSSguX3za0lD+U9306N+m7Zso45KGbxGx8XO7y
PkHrrXtLbIKdT2CWqUu2+mBiyElF8l8RzPpblTM0F6vVBZdd313hsqY385QeYb8R
+mdXeHzgiJESclWv4HG33nFgoze/gkCniVVIgdlUSuvunf7ld5Q719lnmyNEiPaj
l1qimJeJviuPDksNfQ3+MGlNA8AMpzouXthpGwNsAEliu312VZ1010fr/izDLxg3
UZ+KZv0WMl6YAoKvTCcW35/eC68+WP36peISqcxSEUC8Y5tSyH3mQPDn074PzosZ
ai5jPVyDJHpA+3vcNLJOGjySFY64WgcqWdLzzhLC2BTcSGnfuEeAsL1iuSNsaxnw
FBFpWE+cwe/CsfZHeCSd/51gBGRrEaEnuBqw7uwvXS1laG7AGMJM/wC5A3822FOz
LzWsMSmkfF4HVrWBLLnUQ8RtoinFjTkvtW0Zk/DRV66PIdiSk2HQa9sCfPqvipXw
NVEjmeRzgjsDB4rB8MBTSuY6wRklLhmFYROgdbgtgT46XBTqQHfpkQf9j3LwAEFb
plVKdvzAyK3nTSihPZMPD5SIz+HhbbdN0imco8LU0hwwcTXTV2fZnGA/x4uhKrw8
SDJW/rxYQuv167dtX+UuoyZAHMpPSlD1nc50h1hwfBTImyWEjcUmqMKz7p7Vwt71
2ovocN+g6tHb19tdQQsuXEbgLWTLnr9UZz9Od7QdaiMVdzaeHbSAiB4dZmreccaU
lDTxN9Ao74WbP+EIg2jwL+HdAd+UfMNuaR3018xaNe8y8a6BPvHdhP3e6JUyDHPe
l3XRyYv9tdGPCFwqLeaFhuuXd11Y6pn9uYqWdH0e5PrkPrKiEMKoDg3U2ZgvVJxH
Hbi19raXCyzF94eSvBuS/fr0FneDmc1R8SQWOIXgN5jE2ha00nQAPUK9RMuU5kCp
BPsLbsSDfsdf1tjDJLDmarFcMsSH/FIeA7bYAJ+2wViKMbyQs+wvIJUnIJeyPpir
lxZVFI8X3X7Tn6AyKf/ga7vcquw/kja6KTw1MbXZlwySFUodVWyFTeK0OyQAiEeA
f3tPYV+5RzC212rpytheEBSuHmJeOsDd+tq3ym851+O8ydGxDTMSSQmB/Cl/r1qA
9sy+C2/QxivQwe7aqG0NVu2kpl8VwiqAKxPWaSAxfLV4PjGUmRRD40joe4/FTDtL
+oAYP/QsmWVcx9blEcwqyL6KZFyEyjcfqiu4gADQml2r85MXu44eE8WlizfJ2Eqs
FE4w7B0p3C6xysu4siO84WhQ/UskYnEKVmugs76m8VLQNYjuBSL9ypMUzn97v5+t
6uBWGcovcSA2fdQoVvonsl6GMFtF36MQRtFL5LZ2vHfQDZ85PfKRE0Kzx6dT3Qcz
rt2ez5GO/DE8gaN60UO9m2R6YdEaBWFhKbmd9+lueXlyAe8jslHxZKRh3mHCs9+w
xz1en63E1qFI186E6xmi3PWKB5UHk1g8oaNM1ske1pUWZTHt1Qcb5U28zNt0QMXo
n/uazRbiqnRIMlguRN9SpfjmWVSsSPhpbL1AouulOZhpjb5wxqmclznfPpp7xLIl
XWl5lnCxrvJble0joA49+q3owTpwBzt1D9IKRlrdU2o2KlkIuiyUA4Wa7C5XVeAc
22tCcqdikNLzBKCvynSXSC1Jk2P0A6WUE4igm3t/o2ne+KIbboeWQndKcY166LDp
5ADfJGwtBBCrP3OBeVc0Dw7AX4ba/XKMfU9+TL4Dg230p1EJu8PCC/xEoxx3mhP6
5xNiWHCj9YkksiVCCLcn6S1E2Yv0BWtDPh/zJSS265z01rnVTQRhqugTuvAps1I/
ttWicRcrlMvjs6LNlIfQO+MKygZPB7jJ7XELelryejYsW2N9hnu1WZQbVAhsraM0
21LG5ytD/MawswbF28DWGpUUm8BzTyAGYeO/Xq7HskjkrJJVSYXKNUgRA18lm9Sd
l0O+wVVE6LHdSwS6pa6wEq0IuGHcLa3Z3+w5QeHJHwh43QzHAjAf8xvURISN8z+e
UMemHpUBENyDuoiZOroLoZkHUXddxCLXi59h2H88bVhF/7z9n57tagamS8ImCMDf
mk7BXSeYgNrmiagHarbq/XwvDLB+r3Y0An5/cbU4nM/KqOA3pFt64wK4xEmI8Ucw
tz7La+Gf6ZMHejxMq03OLU17M929yn+FJHPq78TImG3mqhd0PVxwie28Wkcgt3FT
NyUhV3VI5+beOBNdItSJ+mOVsCtMqWAFu8CjMSrrOX/qimG6Un0upibfoVtSlgQo
cpCOllntAvmhJsqIphijQAe5gaKC+TPYu30xXoXwYOjUKLjH22DHJ9rIll6peqPi
DI1XlQ2QCEODaq99FGvgA0jxeAED7I2Rn4mQ4cOka3MOJeX6FKikj2AYf3wC6DqP
wyDIIBFey95aJHO+vBXiYuRbx7qpIrUggcMi0x04c6zyqJ/RImrEgEiRtfqI6zgn
hSYlDK7OcgXpk+fptJAmSG5jkF34LQEvXvKm/Uno82ZHoARb8zylxNMFaeUm+cok
mpR9hBMhXCx/GF/8uZoH68KQIZhHXrGCpaPpUeK2yJGjyKPQIQHF85PXn1Mx13j9
zV8D+iWVOojUdimXNfcnfLqBV+WXEcRNBuq/R1AoUGQDw/cvNXkdMWfWsZmYorVC
LGveJA9X/HVV+v2SxlaUETA/lmcoeXi+jR2ZRhbLjgn2YlLgqbu4bPH36v8etO45
Vi4xuDAtezJ3kn+CyWjvNQjtwAWiETs/uzf8Q6PjwcjBlSmOVG9coIlnaeI3FMcN
PoaAPM6Phqt2xRTc9wUd09Idp7h/uMaWVPSvfWrtGBGOm1FRHC/vRbjE05KxD04q
3rTbxTIinHJAvbxqyNF5bxAd92rxRF4QybRoKzxYDrnxYjIAQc94Q4Rl2xB8SWJX
4yeMFm9/ryZy5HWrpoG8X/5+D8BhvnnltMbZim7Ofk86stBbnItxWvMWN/xtitho
zxP8sswqRbuhWuYY9ddyPuNBTmwHfij7Rs1UZIYVJgUBtUf5iV+u0A30RsT5vtTH
hw3UY8w6GNYcim4TD1ZmQVjba1YEwWanrPrCKPm2ttbrRKHbrwCqizVvzpFDdom2
mzNrjMhI+nXkc0VhxYqU5uVa8utRaE3JGXrlYBUmDAZ9/ZpQIApKfIYk6pwK1Ohu
B7mSg0IDVtCYqfgUuFPq09leyFl3CENdWmiQg6M1dZqvkxf8FZMm9+VzKzX5RhXs
ozTuSTXv6/8I4XjwnYExzzMNp6hPCOX4fYX4ts+EFjZ3+ysO7bI/Fx24ISQOnKbf
3c9MIpClazbeGvJ1jMPYerJ4D9y65bjAUbLLza1CqDgMg2rj38o8PYzl3UA+bUK1
lBFrKD8w2TR/ofWMSyqmjP+8+ROCJl4w3lDLcKbxpWqnejXaafiAIpra/Xa7KAMs
+RoreM+n0+3bsrYBCTP5NzJVPJROhP23BiA6YWsChvFkZ+kocAqMmmR4n2sMA+ZF
6Lq3ykmpRpExiamX1kma9Z6De8XoNhdxW8obGIlv8DdxTWd69l7YEh82Rm8YKp1I
Rz14wv0EtO+/6DY8DhQ0tzmsoEDdl/whcTeTyyNyvtKr/U94v9bTrzgyWpiuoG7r
o/o8XHAwb4i/LCtlFyNqH0jZSIYQs7CT0MeJwPzAtHVep/k0hiXTlEIuJXWpKy0J
Ri5TvD61veFhzK/3jvui9N/snnbYMLnHeCEh+sU8ZdwFBeIhxDnsNG8z4hDVtQze
wnsM8SWKi49YvxGM1CULLo9b2IH9D8Mz7uhfSsNp0/ncRdKvk6sWnHN6IhjJkpwC
sjJZIBYopywwlW1h959fB65Ntr2RRHFhhmstdp1ZGeR3VRhWJRSYKEsS/8JbrIND
VP+NV0ySghl5NTeMxmLJoE9g3I6H4ZmJwsqRiFR5uBzQw4LTt9l5IFeEMJuAR2mD
1hv0hmw2Ahawz8Tem6UIVAEzAvfoWelLKlxbt5B9SIlI6Dxt13+nmnSOJYSYOwna
10mnA8iQtiTcDcIkIk03RDxWBh5k47kyLATOHlBxgZzT6dSbFMMQXuXcyE4KLGLm
e1jr92/mBqMfZIJlErxGHIlsohG1nbUurss0LuwNWynN56uQXleJc0jMaBeZwkO3
sRWIGOr/ENyUyrVyxXO7LnhtQibd8KmzD/BNInZ5zlbUJelS2tKcCoUxQKwxNhqS
KrYo8EABBYEMIOUHkPqH1YImAhVi847PwIxppLupu37a8UPM07khfp7WHcJxL6z0
kvtFEreNF1LdWbYvmkzxt26syY9pXPck6n5/A//9KidwW7alva2/Bf2hyZkhx8U0
GHoEnpVuBcRY7cBDcO4Q9eRTrwOfizpqQvDTqDnoMlKcB0g4puSmP38ObxhcgOfL
X1gYIKeNhp+kNQDmlIVFMM0yW7QJKq8m1ytNediB9E8hgFskswNPnlI4IS8eyDF9
2SJwLcbZDU/tLZvceAEpqS/pLIpmgojAEHM3Pp09Z0S1q0HKnNn24fCJXBn4rX+J
UUz9whXcwp8r2xoQbI3NzVrgjiPX5PbGTsCLGS9/G6ea0YDfDAvp/VPgkQVUOPur
WNb9B4xk0rI2YkB1KcIDouVECHSyOtRFZRbJMeFB6G2Ij3zSRCp4R5fmTPMtXQCP
AtYAU/uvPhdXQiEfnAEq0+Hy1kddR2qTI+z1MDu8Y2N/XNOff5Czvnfwx+cRehos
XAMHGsv+79TS8Gts5f/N/AG5cejo2YRqzleYM8yE9GCihnkHc1l6mn5zW4dcfPhp
xW1Daj6njqXDuMj1SLLVL1BHfLjzES40DTHOCQBFJfWnW7aX23fBGCOSKqCQPMN5
8aXaY+DX4exczBBrOvg+lPdGCBbZrzde1IOYaz7Ta8JCHvDqB5NubREfEz/4tMfl
J3XPPOpokUCsolm5i3lZm/ILzydJCjuoYyo+orUd6gIL9rsMbWAvJtYQeejf+eAF
N6CvoeRkYfsmD7LV6uLxpJCtzwGjzWTUbKob0Cp4Lhifn2BQvPBVg9seW8NrhZu0
VnJYOiiwY4px/UaRH0l7boFN7ju0xMGIH0mlADJlzC5JAecXDzzY79kyR7Pcc72w
GBdeetaLW8On36FRlMkV05CmXyUQmTigIlfpd4N5Vht4ZkqOL31NKnF2obVvQTqy
WkwbH7JrN0Tiqcxpv29tpcMAOayioRYvzx9llM2uWRdEr4ptdAv5Ufmg3AYP1JMx
POXitOn3DkRJL2QotrxRvYRTHLLYqdOwQNy0CXeV9Jhu5Wa1RWDNVTSt4oY7b0R7
tdnHA8lK4+pnq6Sb8gszbVtP5j1tHUCnuvvLdphtYP4TCT3FDo9+FOEKvYk3Pivj
CCpAu65c2tchxykF0xwba8ZgEYLBiJDKeQXpfFCz57rY+GBpRZohfqgLcgvDPkf5
mHNq22tTx5b5soiMqRiVeuwbSmQ8s7m1syx4sisive8J+BHBO+4gZ511HBWKPH+K
SS1ROKxCPWwNb0AJavcPk2BcfqL7jZExYorHr46YCu+wNZYlue6xsC30ObsfIl3R
ojC1ofRlddDvb3QRES1nlJB3W1ZuYwVU/EFX0ZAsJJ7oE0zRkd6+YEg7hmJitpRU
5j4hbiO+ylT+FPYQKnf/CthpnVIZh5UdhwgWAqwzUyyqqrt3vHXaSGL1iOzuhnCc
19rToPadUOsLUrrjcY8gI07j4Y2dZxDsRlslTXTU9aEeiF4OCQgfCjJawyTrPYSr
KZg8nOWVrXAGyUC4n31q210piNt68lvDXfAUPVLkxx0HQVIIv2DM2nUCC4+MSb71
Cni4AJm4wU/rpzj029RuJRGpEPKv6wgXgdycJrwWqXXqQGFj9dex0E+2iUb8oQVa
pH1jAB+eXTwWKuUIc/5Wl3Hn8jF89QjKGBQJN3TPQAgRkmLqkaM9S9EzbFB+MxcB
qMPVAKYAkZXUTu1JV9540E7jiASMVLYo5bgKPpMxUEc3YSUT/xdvaGvw8+dnBUG+
uAGGjmVgvyLvantML5GrUnEJkycwlcQiB4dSmSGKe+sJaKjkzk25Bhlw9pLWslfS
6lzl57mJ96Xn29xHNLPtPVoViG37TVg9dbj6Ezh/VslaPVcvXgMdofTEUNa8wFMA
Yu+T6Ub8NL9lPEJvp0VZOk95cGoXdREt+81u3VgQ7v5ZTMBdqn3MfUp6rf7ZDnYs
PGQhwQIAkvzvA0Oe9ILtS2zywe/f4pG0VaXEzpCEyhqjH8Wh/SAnw1gaNIubtZ5L
8A6trlFe6F0ne3wo3PajAKk8SDbOYSHJhwk5T0YAjhNMZc/bpiEI9pO6eMAWwW2P
REsGpX7idTvF87czIZZWvwuH2rSQF2l8Ls0WTTSWp6sx7k3VDXYdVbNSvjokbVCK
7a07trv7BgxNBkIbRHnTNkm9HWXOtAjmPxzr+IY0ab1Gep8QSLIcz03i9YzaLb5E
77KFmZ9NHaTBSl8epgEz5JnZsoYDJu+O2av+63V1HF2d8+wzv2tVsqtp6EY/5Gsm
6LibIrNfv5eO8r88W49sV+wEmArHneIAgTxesKMse4fXENlRRilZWOZQOybOD1Te
Q8n0O3l/z4qbjgBPhSNrnlPN5es8ngiWBgr84PEvcEQmVr+2YcpJShisaV6a+O6x
3CGynanw4pH6PQEgfo8PLpje0aCS+QjaipAKqRfIJKF16ojLkr96Cb3AkGDXEWMN
LW8rPZ6nTtI/x91/FaPdRZ5JMk2lnI6TFjawCynKC7lxxh3urkMra+o7LQfS+6HL
zXP8JfwYpVfy1T2XIRws7r58uYK+yE/uuRv1Hfw8aK9gKDLcHmZTosvgPxdx1v4B
jjA5uSAzKfllwuqjfuPjje/3vUlgNOPo2qnbWfhMMnJIgvLdw9g7bPBVLPD2SSTG
7kfTD8krELAizi5LQoDM4i363bLnJ3b6aCiSUFChAQublwWM209xIMey/SDm0pM6
W+V/f9RssSmElS/HE8ZJF5kiuWCIkxxhaLpBwnvj0jU4sHazM4HLwk9A+jFHgnOL
uLZLchDILAv9HVPktOkoXAE7L32zIYEBESaZmLpVpgWpDiFhrIwu3NRbFXZ5Gxsc
AdqgjqqH6GSfiPQmFoibjLPypHw5efgn3NA798roLTJ5BiWQXCvZzb5IQRYr1E/T
sV1utCAN1i6C5SMHQ07soWFjhk0/6ubSojOb9UXg8AvBFin1JMCJZMdHOPpBOuQI
BOtBLa1gPIljtkCNd23bEeMQIveiHOOu6DSGHU7/qAnpA8Rqp98a3IsYKjoA3KAp
dZp7L/h3uviyynBW7kKWQUUGNLd2r6IUYBvGzVOSoCT00FbaRLGOI8WVoENu15kC
bspQ2COOKGQminv/PLmFrW9GL7Vbulr1bJk1DyT9IgFvOwq9PELGSL0pRWgXFk3U
tQ87VRMguZSBNnUt5GKC0Wrwz07IosTyD52xh+aMvKsyVYPvmRLQnPxq4RhDYwmZ
xR42yuQkOZjrSII2HyiNZ0RNZWFN2aFzEVe95ZDgalDGWMNXzVFlOnndxAfo/9tg
0QoRgbIEd4vUMjhA0Yx463RkO9unrddT2vuZscSndGru1ttV1jukwtiudC8fUDDJ
2gMz7PaLBOvXxGH5dpxnfOYF8xROeWJXZxsu+XZwT9puEUm4ouoiJwi7B4J2NH55
Qji3r1n9flubBbydrGIkjtNxPMGePJXt2Af3wWxLNjxI6d8IdlxiR9D5fXD9UwIz
d2JlwobPwG1bjOGFAixLtV8q09EpIbmtmpYGDm/6WOF77e4+KJ7G9LPBhPVyJvYb
eC5vYcub+zCRq5hEMEBBQ/GgyAArodaI3kHRGtjAEjLv0vulgMN+gXydV0Wje2TC
610q2AhDZJZpBMW3tJwxgE2Gof51bFXzsNUIT5U2CZK6C4XIDhq7AqM9Tcb1uswm
CNJnAVEDdPtdhNfZV6DVnoWUlFAT+Fo4LA9V0LO1jETDW5T29zmM/Xo2sQBIghIC
IbOHwpFdk6OIHpVWfXcwFPgGmNtWjwGGwKw97r9F4a1cfNY8lg3Laxr0oRjkL1HT
UtyQwWDXr7OplADqI6kcDdDfwOXzpKfpeCL+rQZqE+twzckAmVWBVEsplvtMMcnL
PPWUJP8Gbef+h6GJGy1Vi9ua6AX3vCAVt4j0UFStsXKece/NFMk5SoBl2QKtJ6YJ
jlnAXmQIhYq8rXkF9eyTyRq+nNS9/V9JfmxJ/ojtW6bPGZ9y6VaySKsBJsOxinN/
osLV9Ex53+eIUIDKVLMx+t6wBbS0+ugA+nWrHcjA6wVaqGOxW81EBwVmYwi9CgaO
MzVsDWfw7rhOS3IBm7euToWY1M1l8H5omQEYyfwGL/Cw3hRu+J0tOwiTaQgw0zQH
DBaYhNu3ZmLzQe06CHFlPTfx8GEC1awU3BDgXvOPJMhZ4nSaIw6qgjT0dqiGnL9f
WbvbDxZHwL2VnmDlpZ2LDfYnOKn9O8vGHrIbQKKszjSfqo4JqNpgb3GG/Xy5mx6x
sPh0TuHSLEn7xBqPQ0HQ6ZAQgaAK5bOIPFDZcaz1bBpRbMlxSuriR+3YBe1cZeRG
Mc5vl4mwtCrQwfHEZ2KMS/4glzTK4SYsgz2dPQN/L+QxCf6Hv0IKfrmWCl5Vjg1o
gcn8xihUpfURuFf+iIDSlRFljctu6Ik08QrWAMPEzQMY1IHTq1Ua5ZepOTJv8s7p
vmNKNy74jGWeO8yUcE0KKS92B4Op15oPK0wGmrIluLgqRQXFeIag1ZpR0TPTE8jf
Qkum5miZvcwpQElSYBMvr0E12eV+QleFqYp1tCLhUAvrp+ggnY4sOVaqpYsKCqGw
+JRqOn1pUztcxBxXfVsMadhAWVtlyVxpjg83TtIe0MG+zrm1+U+FlAsR5iFa2zPv
etwz9pqWGUBjxD1DMHR6qU8NhqrFvQBOG3UNNoZJl7NlHBBYAjQ/dFncfZy94EMI
nRMuYTP0mgD9VMEk8XCfGTQUmb86/UmGjUK+NQXLHHc3GkLV48pl23R0LZLA4nyc
i6ZSl8UagH/mn765tpzCjG9eT44lggKvXRETo5MWn0xMoRmqbLKJPuj5YEX4/luQ
QTK2Fw5DkPtzZVmTcBuoGNYrss9P6NKdnkvC/mgXqEFeRwpMFwgdAo8RdpbbQyGu
kff5BMxRmc0ozksn5poy4tx6ePuP2yXyKt9xcqSa/hIdE2+wRrAFLjtoq1JygRLC
AyQxvV3Po4wSIb/x1L9dLs1lW8Nfw2SZJWTNK7kTj74Q1rtAhtaDmTeREz5jw7yd
iTmDY9RcUFssHIKx2CDfqZKIMsjU+fj4VBM+GdqacSpb+DFZNLrUFGHbyL55r3Qv
L6HKLp6eq2g+C9qqoZE+Yj+jOINLSFQpEHIJ5FCdRXbLdauuT2qUgN+uFd2AbSdI
EgWhhaZ6UyWvng5nabxWZDnvBgDXYgd8fqfyDUQizNuFWcquLPU35JRXrZyzAMbu
uYthslZpAZeobxv9HtWJ0XoA2pd+o/673K0sux14IVgMQO63efiZDoIQzEL7tgOf
G4Fyz4ZLRPrKbpkw3Y9pSGHzA5VUctUyHiHIDzhAi6huf4y2XhLaSvLJSneP15Jm
O8CVshbxEYFqAkhrKcwRkreaM3wkHYG/xLwObuezUYEx2CYL9N3K/2zvwPnRN0PW
2R7FEQ+1E0V3tlc6eNjQ4t1OS/9s9l3kRjrtri9Sq6Cmy/4exm5quyICTUOydcw1
MYuHoajwPBccjHfP8njMP9adY0Qgvno4yMFlIOiu17GQlV+DpNbIpT7Wi0K/yYLB
DZBGw97Sfa5AJmx4PprkYH1ejDpQ2XWESbP8+psq/CWCTU3L18fbOL46bJKDJ+C7
iuztrYcvEziXwcjp9ts2x1tRpmnw5+gGMxcCqgbp93M5aVs8ocEA/Y4L0yOH+VFH
zmh/zKOh47FnvgOwqdfJDgkahuY0RG3U2Nfr38jMO2eOP/Q+yK/5Tuirdopy+THt
XjdUREHEEiTLsskJVHDAQuxKGCNTuTWNJ5StFlR1ujQGCuiV7Zwa8CzI1GUg5E7f
1RD6Qcl59e8ItQ09fJS3u8HXcWQJqkPNaANOQyXBqTKfbOfIH2zYWLwJVMwRIy7D
a1MORDRweSfALJ9S1FMUQGgbU2B6UaWC2bAqf8guTxizPETW/ya6SjvpCg+uDBPI
xN4bcqD0qpXJvMm0/a7pCmRNjscK/lBVsGrb0NPLdLrjDq0xaeQZrRi2gjSH2Fzo
ppG5vax6Dyggl9SWrnpXUCoQZHGYQYyigWaypvX8mYdDjs09PUCP5rDAjq3u7Hoy
pPFkwIuGvi6TZnkxjqC9OXN2a+w/ZrkNbAcx1agwu9N3gjVNp4MNY2qNdPwhcsBM
nCp2lQcwSWvPP30I1k3ZUeZVs1hF2RL0I5gywhxgXFCnoZEoHqcsMpEkeqGs3RYd
EaN36yrOXU/Dtmnl8vZ6lShtmTgYpYSxn+czPV5WKUALyYZ1Hq4ev9iCX5evYftg
FHcMJNXRCByYTn0A0F+0MtMMsjVraOmBLNjh/lvvERJ4nXIYkm9JG4tWCn67Ox3F
Bq9laS3w56Awm9gJ6oRQDpcXva+I9IsGcql30nBVBgP+EMVy27VFCcx1qKhpYo6X
YNEI1i77lD9tjFh+lW+Lt2qBfR9LM28bZuvWPIsy1Efy84w8QrTkLchfvRHCU0CX
J6cRj6WORHo73F0+eRYe0DntRj9QRxOZ7kjZzdDyJ/0zmnEat1N18Y0QOCU1iU7i
8xwP9FZAWqol8AiXUXkCrnqHHC9aRLWpMA2xowT0bGS7iwhiiINin5g77DnaD1+L
s2EXO0LcCjwirtZI4BeFPKzZq1/Cmhaq7eA0+aa55i2QQXSv4RWZGLademJLoZMw
IbdmDuCZnIKiO2rCUqRrDqMy03JPVfUfU8zwknIgVXvtU+xaw/brvpZr6EInCdlj
YQ4EG/25rIM7FUVBd+nOHprorXRbceDFKVhAChF/lNPBczLk8zYzQKxI6fKj3cF5
nnLqzRmtSqyB8qEEw/CrcdC7rgNusTV+SLt5jh8FHV3jzfT0HJaz0EvOTsdJrq14
CHeVBhnFIl2tK/m51kT91ZZwytIkryUjVDT10K2E1Y6ltMCp/OBW3BGp102GIHtX
cMew9pF4yEkSHd6CQKV6D178iX2fVfjqiIzv0ccyiGDdWvFR6E5Vk4ItE/qmQ/jG
1xNRr9N+RwXCc6TBzbkgEvZsBqMA4OxrKxO5uhKcCvt9MpV3g4W1e0rAkJS0Uzfd
jb5P8HZwr2Tlo3hNNENivpiJJgGS9FJXDVpFC76wsIK/ZeM0nJkBo0YYc8PwNbyF
2XSFri1VrwPiXyhra/T3wOYRQAc2aW6FDWcIPla3msL7cZWLNItVYrtMC/bYge9g
MOqHL3KFkipyKRbWdjtjnOBLmqqiQHEPbpyABFW6N0tmHVgQSHUGqXMd/CZZsNeA
kZu4f+i3NnkzfTA1usD3fGu0lBP6fwH+cwVCmv6I+yoAfMEkIja9IrBpnhz8Iiez
X5POSU3wEdfTsi9vhd2lJxJgC4ywSJvGIj3waGlkrIW0EkJE0aZEi/GP18xE1xX4
Snn2Qj1O4EeWQpPlH8vcF6BIwSa8mCacB7mbiYnsbwkMtPyCNFBmMzivL4SiTI6e
LfCSyptaTa9fQnYAx18Ircy+m+AoIgQD3yl1MGjBXr44CxuUlZcQT1yOb5TTZLyx
DZoE6THDLb0C+rcpLHgNhisi0356ouYBIysiluEzzxSb36F1rR0M6Nf5hcL1d6q4
l4hMImx+a/EJpJ1Ja0hz9iIT/907gF5Iuw2a7UoRCzFHDHt6761ZeYYaLiLI9fKq
KOM/vUBpypAB7A7sK3gGkDgymqIfOoBmsvbNNtZG29MY2Of/cYLRz78FwLUpmD/E
+fxV1QgjvLSyNM/nulaHrL5ukVari6ZkEB+4x9cV7y8q9y6wUb0m6GcwFFT5Y3ce
xUCF4Zt61NE46VSxqpvAOwlwwpsIK0f6L44AGV5F/WbCr1Nk8aPxr397kLoP3zts
MGDUOBL7zYuKkxgUsfJezVW+JSh/VV40kj+ecyDL5xa34Wsf8Ss3n8vek3MRN4Ob
2ugrMsFMKm1J/NALghd4W7PlmIhoVAt5qiTRrx46s8oKjZ6U0ic36vTvm16s9p3y
GD8QArvrgzkDHxyJzyaogsNwgO8HuqhkCfkaj7JAtA5grao4snBBqgSL0ebxn2W8
q74k8xEnWxz5aFrlW5FhJFxIuxL0+w2zQOVWeyuAqFN3Q6apnPwIXlCumICqQUhI
lHQX5KUNx0GGi+yPivfQstr139c5Xb3si7X0SlzGZCeEpWw1nPX47MRllj6FKd0a
/KdPBDlSzL1a0Uheqqf7wqPE6NsNvG+UV9tLEacyK8cYc5BV2pX8MTZbcq7vIVnq
Yi7ztYISN0hdIoBC0LiqEy1in7Nv1g3IS3JQfjPPm6qUAvXX+jFPl9GSzMDzpgnv
+UBZAI71Vpu4688yn+Gzg3YdHnvAqpssqRN/sHM76izzCVsCj2rUuQhQoEsztIuU
iNsqfuzLTl81fE7nmLt1ZT3VNhHnMbPmIPNyBVcDomycF795wDVChTmt1qbrFqP3
BAoj73RQzcFM6KLuuIJqhd2xuOqiYEcYgZRTCgWBWWsD/bw+g36u7q7lv/+N4SBz
z84iQzxJTtsFJ2fUbAVD4N2tuSkI4vcKduisg+s1feSRiuj/O7zMCN+Ey9r5M9hc
mEGP/eKH6VLIYQ5tZB0oRJp7vN59oiA9Pm+ybP42HFRnCDAybg7Yzwvr938mTW6s
8Jcj+rJhA8nL/ojLYCTzyRvFUUyhEKmC5S28YhBpv0zG2GE167Jd2tdLojpGbmdI
DTzus1Bhpm66BTdjXDkCNuXcRBqJrPTIScHWXSwq8/IRpHMKMdvOEu+BkeAukIQC
yXJYe3bdfd/R/4fw4RZjgaMYFegZs2FP0/xp4cBd75fa2Mr9NVftTMfh80nY7QoB
u+M90DYaWM0Y6o2gjD3t+lgtrqmQBIoOp162aJHvb+A2lDa2/k39woc6MoPn0KaQ
Kgw/sJxZ0urPlmNuy6esl8c/5UJriPRrNJonXFZ0bJyGXd/ywaYKlzAhH/uMJ4PP
iyBECxDulI/zDOqo1ZNIJei8eeVJTnAeEc35ay6pqJ57nWxmE8W7hBZH0ppLFbEe
ZzVtz9SgmHT91IWNrqiWI8VGCT8KQ9DmBSi684+NBvPkIzXddadyksIXEzkuyNwy
7VkYiRGwRh/WMozsFWuUA02X3v/WpxYaXJVZpuu5AwIFrby2CZrE3wNnj56zEZxn
lKG9RiJ1Fw460ouO8fAahwjCm2iPAMxgO2V4zlnaZSDIhhOcYCS9zAegSlAPbXYJ
g2VirQAxNWEwo9J+bZuJFL+GRZX4xR7vJCcBTGaSB4cQ75dvx8SPZnGL2B1BSUFV
GoYWP1Uzuzb/P180vj29LhupzbfGMuIC7a+m3LT/Jb04LHMmLfjUUJU7ELU5CPVh
`protect END_PROTECTED
