`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9XM/vZY/VX8oz9fUkSAYi5NWtJsGAF2jQLsH+HcvBHco3gc+Bj5GZ7NXypuA9RNK
lhnh1z+ygL2zUs4fC0WGfILJ9PWKqLxG/cbL86aPhEG/pcNUsfHS2Zi0xlvmsaK9
mJ7Rz1IzDNs2qXjKzW3acpI6wTORd7XHOU3MVw7KRtuu45oyVxWWeGRWhgRWt32b
Z3KFzSQ7RjSeeAS7keCbPD2DNiep8bdpMPRmI2pzwci3AAqS7yK6hgMFRIYex+ve
RoPko+x5OSiXjE589X5abM0/fkWjXZ50It/0Nhif0W3nQPkWNMQTKj3DinMipENs
9kT0kgHY6Zx8DJ8abp3Of4dew44AupYqjLdCVURYSRO/NaFPAv8lJl9VOxjZ6I/o
vIYFmJP3XnlptvKyz8cTIL48cSKWZdNI/HG01hXvuy5B/9LI2u8/f8WOVLwr1g2l
5TcYm8fxHTaFKypGobz23OB/c+9AjutSBwNw+PwZMZmJQ2TNuzJQn52t58ij+sy0
UOn8HtLYlsXVuepnVU+oyqEefYHjOHykyqvXrW+zZ8yjiHZ7C+iXbXLdSrRtXUjy
AOCPhP7iZR3MoxzIR4RSZXiB90x90+2mnD3EagNUW+S88z4Pxuv6zKR9csYMpy+J
QCmUqr6FjBsL+Ya48Dc1Ui+J4OhZtUY1hElH9ASgznkKq8rUQnZJRIQHp70PY16i
dnwMBx8YURPucKRS/+ZgBL274sDoHKe2l7pxG3hPrJ0jmeJZbGL7LniAuYXY/Sv/
WMk9UtJq2TsAoasrccEUMbjOPBdAGMalfyqOYMacsZbfLkIu1PNOvsTzlvVskVVk
wHCZGG8C3utfhQYG92mmJxceFlcI4yX5TXoOikiy8KgH0mv97sdlROCljV07c2Om
Z4+NDm7qQ59uXs9tliPz7A84I/f6BJ1cG2JOpjteC9MVQsab7zDYgR4x2eHgcc4S
zcxgs1GFvCltmi8M46DZLrqRG/+SJjxOy0LP3diruv3q54u7lDDH2C2FmOVF0jao
oleYnhLLk7XMfSytjpdGbm91qBnPMm28o5W4HktMRQo+8Y7iNvKyZTi/kraosSan
70JsmphO+Bq30ssliMqnsh6H1QZ2YB7ZenPWu4QXNkOVsmgGmQesTsONPGI9JCdX
9Iy8UPF9stzpIrSjQj/jhQPppYnh5slSghjRfe+5xEBV3NraKKZIG649S8mUYsHL
+Mql9505x6IPAUm826fRbOYPcjrk7ZL26/n/u9sRPlUI2qqHA9r49tOiXW6mDe+G
PvCmwKF4NDK0RBvGk03AmQuDbQfVk2ILzhRHPze5ABc/44t1q0+kHfXSBzwbbSA0
y172bIQVfhJe6J30NA9xKj7ZUVMz50Fv3hUcVwtxuysZtF5RlAtzFjhh2u2jYo5N
fnUVxFYZqFobtfLeFgTAXILfwsJtZG5c9FTWce4W8X1lrSB4EI9o7gUBN/67/Hay
zTHRZTl2DT0xtWtp9vKOEpe6ON3VKaG/n2ulMMwWQAgoDajbJ66pawezABk1geHj
al0rraMsvLQPqpoOwt/hWSxfqdWTBCFyliaDblKIlf+GPwHsVdmONQ/m6ytyPTkA
/l/gVFlWA5ua8i+0SbTNePmHIPmoesJGoZKBGneANl5z3MSkohPcNJjrl5u3o+ct
5qjmnykXhGpjkdaZnYtx+PAbh/xUZDM1T8/oIc8gv+IgzzqeWETh9Zdg14i8pcch
3L82WUlIDT1XNOPqh3+RHYUVmV3d4mO5nzHXpyR1PHNx87Fa89xFBP1MFGgzrGFP
WN3hTQXFxxdTMOI3sp4Uu5HdXJDSOSrZilSDeeKwj1+9KkdqFz2Qz5kdsQfae5H/
tFex0zfNV26BalvMr2TLwn8YMpkHqXPdrcx6+5N/qKTk4B+KMmDK4G7b9hxY6ipC
iYXbvwZjqRXBcvLpQIyf3r3gTDH5rpy/O4MLu01vUUVLEtORC0O78uKiaS3n1Tlq
mYR1L5dSV6nG+md1DDEGHX/0WoGbg+JC1hM7OfQl1LsgzgDcJ40JDlu/zQjxe3PL
S9jJoy3yHb99QM7wg7ShtHH5C/pJLGUa5P9/RaSDC0nmD2Bhdrv9XQuwIk47RauA
6tH9KJKuEWTBNrEvF/4XH+TslNCxuorb0caww2ew79skbETNPHvFQSPdNAwmpOET
i5QZs6/6yK0kUGwC6sSE8t7Ue99qPFjJrjd7MHvJB17dEuAgBMLo3WzXDtksoFdU
ECTzGOAeSCijwVZQKpjwEXedYaKK/7sXk7N3lJbI1EOt7MclEL2BkZpvkD9NSjYo
AjomjZdcKvEEkCXOrFbdUpsWdk7aojIHNOH35uA8CSQoMzUtfnK588JWTQrHpzWI
BYEw5ML4B/8RK74HEUnLekQmrPOaCd72NTUvNYilVItxminl2WKyWxSBL3VswOpV
GJLOmTfy8+gXSAvQIVDqTx94ZU2JQDennJgGRJkLmPZlbY5lgZLmf8LrvW8SnPbm
d7Kr93QZzHcmzRkFaj+N5/yppayjfC/8aqZRju0vpQPfXqabvdEdTHmtpw2hyB8R
lfJow7BtakecLV9g1SNtFaTL5tADM1SfqfD21o8886aW0W2NFABU450N+WefqfqG
JkPKaNEFaDrSeQGeyQwOPy32stKPzu0EgoKTiYiMlYmZ6hHdpuIbwp42MU+26CvW
bEvH6eVCUA2t9Y+eVqENfytMygrwkCW5sBgwhGkZi6lhDZZeiAITDsFdphm4TCh+
tvM2KZzO2L1yMTzCVQM5hfuf5WfERvkR4WVXl879JxOgKDB95G64JeWoQZki70VB
3/bGiHtn3+3ixoqNjUt391zw4ij8P4B3sCszKymFozkjqeITFBgpcM2L/lM4mYwh
3MYBAAIc+BRAuRu9THDhXo+h/tpe3qnDnUO+ARlx7tRWEG6YgN88oDmuhXrtgHoi
jAoqxGeI1uDTMzmSL3ECcrs21xF73IQ1v33uized8Aip5+7wBThL5okwIRYCtjuY
rlLcMKgW8iddns3tjKTyljvxYqu0kfpYJsIz0T179+MwuGDSRMNMyAmlgykz+d68
OlClnEfZaZ5sgC0ir5cA2AeKmn4Mw/olp6QvtLNtys0foxsFY7KdOUsqZM1BczH+
v4m6+qQHxhA2VULziUtHZko6jVHUFNfEHN6RTkOi6qEI6d2GKEg/K3NK3wOMvJCM
ARybBwT8OFwATS9z3JBPZKWbdEZRspZ+mvqCFJHd8hboKKQiDlBM3QVrhdrz2aHI
KtTHRfF0fkf2qYudMbmphJv4G2FoLCDSHzYnLguA3GFK4K8piQMM2oWKv3FdjnN6
nAnFmB1fMSyd1kf2EhJ3k0WwxRpxUWmNDpP1sKJCD92zymakSFOK9ylgO1fa8HSc
yr9Wj2Ay1tNaQ5vSJynPJRyT8TfLibm+ysGY1EJuX6FODLzR6SYfw3yw1LgV+Io5
siaJxDW8z6Lek6rpsKJ2EP73sJFe58ILgZ12d80/9mb/0bBZruzcGT11H6B4jEAF
hsj/n4kCntzxj648wQD5Aawj4Oq0VeLjs66F4n6/OJCdRJDKh3DzqrghycxXNwtP
OPehLjfV0tTfreWZ9NMVIIEVw4u+q6gFYbRD9KfKCmazV4gw/xbNM7hFRvuKgD9I
R1DYZSBcitpF3MUtuVeCUeD5dPfTVSydpzaH+7+mbOYCw8QZQEi1QWrGsqRxUnZ/
qbGoqFvLhj1HFQVko4Ax44E0Al4IEzHKFMYP2PYWi/aAeKLs/XCyiwI4AEa0Cn/X
Vqfmy7KZUop3G2rW/t24bvQoA3h+u3dxR0Wy/Lf/+2kpm9+Ou+eRc0w9gcGGp94h
no/t22kTz8QDegk4auYE3dAXo1kWyozzOJdkt/cyHvrhKH37MVKfXA3f22+c0+XL
XQjQ6hb3LM99l0QQvYtV3UJ2Rwap9hVdlyPZbnkf6OL1ugaOYs33MrRSCnhJxaRB
F/GhI9tGf7yu7bVATfwlRc/DP9d7r6j05b36RZiAR/RWPqxET1ipyQQrGqTTEkSB
1TzPA0IOGlnBJbOsEXyYP1aENMPLIJHDQhXE4ue6UCOuBnVSbRkgcb3FfZ/uU0N/
SqZEZ+zIJXxjHP20zJFr7T06npFMPNDADmBXCDO0BABytUOHYt1gYRspr8KQZ658
C2JnqqZpexIdSH4fUKgW7djC8BitwjvKnCKd3Aj1B1OCCt/YPYtpau+4MqDXTuUI
1KW9CN5h6YXNmiZPgdJhSusgiQIzVqk0dgeLXNrxr8NRdtQCfLlCy/ZO4L6KBYD4
glItvpR34+ozm1F7fwMDJ/nvWDApaK4Kh69pvfqtN0T4m/Bl17VSpW2686JPWkFQ
jAQyuzdKNwxFn395qZlWPeXDHXTUfG1BNwdLw7qbK2TLjNpEauzeGxUr/n+kW4BX
Flg7fQk1yPkzrbOCeShqQ88auuLERQjYCnpL8tZBAhujUO/JdVMaOYGotrg2tUcD
B+KdARuTkQVmfBzGRCADSxYzb1ukfUAdsrcXRVKIbrHlWUVRWdT7V6+LAK5ITuWk
JgMmFJxQi1PvIyBYn49CcyJteixZtN41fWXkqhSBtlQKR/3z24gohTSXdGFFZQTE
0ygInH677njA8uYsIgRkxNTAcaOBpahP+vaC57HWOcfV3TPZgTBRUbtOwuhuuhIL
LL3+qDh/PmJSTc9aR3C+ogtAqJ/T+NLFlYFhJe38Cbymsq8igwX4RXN4xphBjdMa
FqvkwkUa8O1nOp5Lsn42Jxc0lPYEvxulIVmb56QkDe4M0tpQ0ZoEikBUIozDekbY
XJsu5P31BRTm1myBICbHZimW3J+F264rYtR/jnP2aboAb0a/Bfu0bN7G7OSWvoGC
IGuIRybNVuMfHQrcWzBlIWeDtNEiJkljZ5Z6htxNnBfP4xeiDT/XF9C1W40qGAuG
jcXPFdzvva9Ehz7vzyhZ65cGxNvZGDO3KQQZJVuqAI/6PGU/ErLuLw9VQ16NNxnY
nbL6nnmmmjYoEmvgw4R2eR5qK3X4GmEijqELKBm6jKlfd/k2F4C3OXZPb+3+/Jm/
W+sqFM7hJDhdAudwUz7zTVhQNN/h8sC8fqUoH4y3sTQN2uakZGnkM5/98HxETULi
vJbHRbr4al+Q22wwyPRuwnYPL2kHfA2nWYiw9s/c+ZA6rJgL4ST3GSJyfPKKZGLe
ivyqWP1DCmH93BSklmmFqF+do/BJNZjjC93prPp1j2Vaauf0zqyIUxEYCHa25NAv
0PhIzOhp/UN18l21H/SwdQn5XSS3HKc1rF7BA2bOFNLdnptUmSunVwk3XssQbfwx
/JyiQgHqNOmWBzr7CvBApp9wnfy/MQkDgQIFgxyJDLvAk29zKMr3QciRL/kwDmLJ
WsGVDVXwi2iyAMpaTu9Byc2xP3jJv7AgrF9jDW2q2HhP7YRLG/3SyJEk2okdbobK
CN7z9v0Wp17G+mFzYNciqs0kYV20kTUjco75QHzh7Co+75jubwQNbqZhb/0NbY/o
C11pRTtDjoKJxfpOCiO9oXo6ECcDd7w7U04jrZoK4yXNvob3Tega4aAz4ZkkbTiB
YY/LC/Lqp5Q+Mb9H1lKVSy6CMoHQOikztCxJfRCQBw4T0JEpRgHwYNKnSXl8bjZM
xx9Pmzb6O3bT91XInNpcw1UV45KPRqG11MsJFXReZqGi2hjEUHkIQgCqfuDUxzV6
Pm9a8lzSHJnzlveOa+TFxpFFsk3pZimHlnYJV3r4zAIxyG3ZNjruHgolmUWtlOZM
bHCijlCqMRFGVxa8D5m07IlyK2/bN8gNemNUqYKyaXLVLTyEgfqmRMjbJreDZxs/
YohNF7SkomcDAyU1Q8jiadZVSeDNAunR/FHmUrHCG+3prJIqkez0O0jHYRh93QMu
fuvoV3o/DYGlqUkJOhXtXOVGIqhKo4Jv2Vkmsosxk3JScz7xslxlxQtApGfnRZaN
2DB97reEAvLyej+WDklFSsl7h8SSjxIDtzpZ0zp9ycdcPLDa7hr52YUuZ3scIdYo
2Zaiy6k6WykVvBLvAnmCYvVD5P6f9vVjJOvMSD6mKCKBN3NnjEHRNoLoI093+Go1
aifAFyuwb+XE4ZeWhIiIAlptqbTKt8jUDU21DbHc/DpB4i5MhX/ExbOiiEiXfkNh
cnCS213P52D4Kbj2SZBRYFDRPdCV1v8q9wIUY/ZfSKPZz9UqxNyN8zOVo2/I1rUs
7dnaCJMyhUCKtUf416ZwW8VCWihipIZgsTC/e1QpUPYg/ahOMsfsRgEwRyQz2Fn5
r/n2hjX32ew9OTvgG0xKHmxBCUWNWVbKKt2zkS3K1S+S+AWBpiK/JFt0Zr6bLwVo
r95H89HTa48+8i3dvZdEBoSdK0j7PLu8x8Rg82YCQcEF7xYQFJ6WxDeo3eL2Ig+y
CrzBs76w9i4jpyv89iytIAecGCVQPsEMDRpbga4voG4jpFDKLBZym/VwLCdcdtiZ
C4hjR7mteX6qV2CZzCsdiyaCZ9DoZwUW5VBKstpirczNlGH2aWq5rsJB8xrf7aJ3
nvMcmGZL/+Svy8sBDqq0HECO8S0GlvrU/UNqXtyQCcxSY8ChArd+snzpZLZR7pb1
1PZQFxZmDc9VhiDV8Fjf5PncHLbeiNk1E+olClwDtLgO6QCZC1RsAmXJTX5MXbXE
2KwxRwVDBYMZ7+Gr5EEoF2OLb5jgHdvrB8YDlryEi8EI+idE90ABoim6gMSHXix4
yDgsBZg7DsG5iVbRHpkNfM/DkrqAVdj4uISMf7pBw6BP1MRr1ZvMBLRTTch1H44w
HhKeNKa/rqbQzIs4yS12aZtW2zVYl0QCg5KcYDKDuV7w8vW8b9fw0ouOot7dWxt4
v6l8kdurQ4lmkr5KZhx/cf4zJzt9QrnA89qRt1WLzgUwdULqwZjfGf7stMCBfMka
r8dNKqslgD7Jm2+OgCXSTk2xlXuGwWwZKfWr50AhqKrI2aY2FK8z47ERhQuJNSSE
0vbGLzDWTTwOycJMMipPwrptvYUdVDpPy/9yshTPV8f1rvGLTbYZ2zzXy6wIT1FS
TaaGZiebru8kFpwJeFOzPPYOfanXPpEKOGH70v+PUmBbvD/+LdBZAr2hsilOaox8
rVPkTkCoL0mOZ+zlAwkC54M4gKeHnyZ5HK1MuOhWB1mB0UfQwug5Txagak+YSnG4
/IKVo2yYL7ggwhG6F/geMcEO9cbexXZBuPWC09Re/VnfMPsYxnq4nOKVwY8pEpHi
7TGa0hsYWxxPAUXkARN2fvz13N9yxDP8TCrBYskiZADWH9OuqCF1vDPubuDFE6yN
GDmWcsQQ4k50S4SvP77p2s6CI8AWASOj+mXMd4fQCPEVPTA6qhaxN+hMGAP0RVbl
L9pvqbMPm7maDTBJf+1SHw1XwglqXpJCpV+okB30Y8/sTstBh8WkG7Z+P8LVd8Mu
LOInWdY6wXp+/KOybQ5w2MakhGBa0DegMkCpeIxO2CrSyniSbae0czbR94bpJWUt
QuGTbSu2ySq9KRnMPuEII0Fa6L0a0uKbYyl7NLbFDoYVqvBbmQJKYbIVHXO9amsi
6jbTOpInZL1vnZAEUJsuhFLuUd5AQmxtlAZbNO7yTSCUSiyhSqMW1TSPs/S9zeC/
RRdo9bkOdtFHzJxKIdCSZUNZAm4xHosR0/j0IKdnXRQBX/4pxzrMefEhn9zk5oqW
Q/Usi1m46qY2UXrAxWqx+1wkeIGSHLF7DwUWX1kHcWS9CCBiaxTJAkU/30kkInfJ
3fEsW9r+dzvJzBHs3C2ZPc1QAEv80Vs1DcRyYOIdD3536pKTz9rVb9Q/W7pzf2AC
HriAyxE9g9yI8T3wRrrZLJGWtwbUdFis4ybcmn0ymIRzUlSluoOOEyHG5vI7CDEd
MhBNEA02mdRDFT4o9zfjla6/mF8althxGAK9NiIJMh5j4dGDNm4cL0VR7BEMrN+w
YTyoEemf2fqG1Z3fvfBbXuijBiiZ385pinW8a886Uv0X17LmULND5VXza2i2XLQ4
mjLNwHki6PmZSW68SOqqVs+f2GvmP70mYEXXb+QhwZQPCGHXdajZ4JeYXzle323V
dDuNOJ3MXoJjGAs6Eq6RM2Nl40bYIi9NPbSpog5XkHtfcLstvqe3PuFG+9aXgBJ+
BQtr48USl+psImH/Z57tLDxCvAIs+ZEcFo0cTJpCYQ9otKfXXdIGr+3QxdZ3kqIV
7/j1YI3WnTgmhS+NhkMo4IWxU+oWbtYUL2/yzR5U/bfJt4nT3BqEy4tDQq3LBBwe
IDV9d0r1NuyqwOy++97lHgSy0vQHmsJtN6cO0ADucBe/wO0FRI6pwq/feY930Es/
+NiXfnuc49ZoggcArIteLK3BCPuRtp1Eg3Ey9GUQaVyNzjSeM5YNKRWW9e6O08sH
YkwlvccNvaZnoms9JuwfNuecPxGldz9zERLFeTKcfeeasCviAiLh1IcDDb40xT/L
NxqTa47hjR4oCSbJf1oPTrLnVJDHkK+xDO9GngHkLPoX1DlGtJ2I4lYA03MMHy2w
EhLLTr+/RovNQTLxTcYquCK+deshuIuu0YHS7CpwlShQYF51shzPto8+6G4PPXAj
88IOFD05VymEd5+wF8DMo0Yi4+kQlidwBABjlc5dJ3PcEiSqh1C/p9zuufSFa+WB
vYTgSi/8A5GjJbGc9ZY9WAc2OuVfxzvqlPEUcAmvDnjhE8W3v1/gggH/XwVmly+p
BZxPW1vi1cVu0XKnI4jZRWYvuGWTPD5MmzZofkpm0JpzRbPtdREkF8P7wkUWhMg/
yyqiRdf6UA3QqcMdV6qdFnGRCY8yYHTfKberUXglcyyBhVva7S31ke48LilUJOsE
3nQ9+ZlVEWP/N4uA9RHXeU1vqdBpcrOgigQ7bm1v1UQxfrzHmPthORhnPQxb7W0Y
gNSCx4/axns4CxZ3lCrFZ9EdF0fSQwdbkFxgkGwPZX+Uu8Aa9VwQRrWESP01M5cN
thyhYsAkevvvm71EcTCgXkpd6jpw8xR8pWyhWXb05OOb9UEhj9WS+8RqmgVAB1UM
acFrG2Nv+YxCcsK69+0CgqLS13tPJDvKRHT3MHe1ipKtTBgOJ/DTKkn6lrKsepxK
8ylpNMTg9IjT4KBz01OBCC3yqgLmi1KxJVyLQVDqBMbr/ZuI2sQpC/xRPrJnwqC4
eomOOM9qAdbWiPZ5CKm4ZS7GJDkgbRCRCrS5Na9UMU3DST8vIhNMfFtjxZv2i8Pg
XuYjtxA5MGUV6cMmspq7xVTIXfBR4wBCdLrEIgLFQ0cyPENr58H+s5TkIjMyvqyp
bPqO7kjcID3mtHv1y3mQN69NqCla3FNWvX+lT9RD+hnfO7bzBSPOWWIsfp2l2r2M
5SvpNgXgw8F0+azk15vYq2wjzhzRhwsfsk1X4KQfvnwwtCPxdVI34YInRSYw2DB2
bVK7xcpxWzWsml9ayuP3q2mV/MsbUyf3gWoefrOwcY2756JaluXdo2tRh90Rj3S7
vDe5ech8cVpFSuEnek6VS8kSxZz0oWCeIHo30DtBgSEPRd4gn3i/50cPSdo7sfxB
4f4/QeJ5QMGc9vyVNVv19r0BnUslJu4aOas2wAg1lNJISD0xh8Rk0eE5YhwIhzsx
knBdYk5Vy/RsRm3nfbmbi82ccfySwLMYRvNgsx5xlfkz3rmt2Q+rV1b4N8w2Rd3D
yKLZ4iE6UVQnI9gYi6GLs/nK6MUgr3WqYgpxLyDYikatoquq/+gU3iT6LXDW0QFu
FuNLH1uhHwJkVuTHUQa0aHJY3I7gPYeEFLmF/mAVHI3I1s3dWNKZH6P7+MmmCrV7
u1O0IprSg9LzOBb0as2xVU8eDX05+zbLD++WhShJZbk=
`protect END_PROTECTED
