`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TuOQQfcJX2DXIWKrjpcj0ApI/gC/nctqe4aKtHfnkCTjQy+nAU3C0ldD6lG57A79
EUOD+9k4eyTi+upk/DYc864Z++Udc1PsLt+9mvotC0F1QnEDXzl+TfTjjqwemtGa
UyBlFFkFHWgfzaGj1njwOwcJ+oWFuS8tGvjXxWdxLcilVKlMaoRmaxMB44EqQ69q
lUnr/it5HpdzV70Ws/JaqxTpcgFCNoEh0bCRg0XPau0GaBxKyGFxZYGsQ3pdQ5kM
4uY5mEbWYI+jWoV25vBmasGfzhzzayBaGezX/19fAdxoddAu+CXw6aWlCoZeRCuy
/SXG5ia5qSE2UIxe7lDsuECy2mAL8RurVx4xy4oB+glhn1KejRV9pJmo/yJEGFmX
p/6OUkhZvnzqJuSLOOuuMqscg7BMOyBhIx7w/+qC4+EQtIpQyXrSKqMf9ALo6KM5
RxJPYusn9Vh/6iYcGQ3k68APcGOZbR5jwPG7o3LQBUEJzI4k0jwl2q1weo04V9eO
WOi4wqcEWaPwaLPnJ9NBl/cNtXCfW3y1Ueczmch3xhyboF217LCsUyQsLNhs1qqK
EOwkK2BvW1sKbNu/meoAHOViCyXGU3nWieIp2pdVdklL2b+9tKmrAse3SEnmu2BC
2S1Lnf1cD7ir2MaHcAjh4LSm5mOxbqc6lzd/u6n+PgIRClcQsmPcWDF6g9wF9k30
p26zMErA/7TrhI2myRYgi4+Th0buuyUelkreeYYsteGTqTn3TvibqDdNbRTEjo6u
7YroP8Ks0AXOhilmreM7n9mK2bZGtLTKI5/6Qa7aZZGqEwWCP/Gqo7yEojpvgHiU
VVzQA8R280e8zB3wFjByRxoQ63wudfAfHWY+8Dnoovt5tduhWVx2l4DybPKqxCAZ
KoA1D+O67VngO4qLxBUFLaB3JUGnnuMA7XU8TlGZjlgQep9UPAcoO9v/eLOHOus3
mAuArjDvW0LGI5WmwRN8gyjlYzlehbMHC2YKyeUq/XGVQA0ZueYM7ybHwTft/iQJ
9NYC6vF5exwsG6DzxUbpmkt3ZXlxh09kx5CqjPN2VH4exD0RApMnVHugNVFvCwyV
W+exmJR8FIZn4uLL6phJbrPNdn8ePs2/lfaaiUEANwdyjwHSBOkLn6Te//TDmMao
ym5WS/NoDGk8uEfdBuG6td08GdSmDRBC+8wFRR3z75Qjs7Hk9ajZ/VcpUDE2m4B5
24VyBywoPQ44qhdLF/+ulgBHMM77r8ed+YmcQmbsvbKEOHwsvGCa+nqvtYdajOgY
WhYPdHRmkU1BB60btyBEGQFBlotTsD5KS99j/6EyvxZfHFsOGddG5nIjlGyUDc7I
E12jPH1uTSVJtrRl3xquKmofAl1J7vt2nscjD2aIcIwwDLEiI8iQ5QPgJ6zB4hv7
q28OBH6y7VVxPLlLHZkvMA==
`protect END_PROTECTED
