`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kug/Qbg+nDCVhV0t9wXck4AciP0ZlQoHy8q85Y9aj5gnGTUKVVpFyrREVnCdV6X0
8QsdOUd95e/VtU4lh3AWyFLe5aUBMoWHJfh1GnGC0/xrXy+42qxZKGcsfvNHfU/1
opf9v2ncAu26ILFw6SfdeZ4KcyrMr8mJgMnUug852BCNoXaRNSXMHMzvNlwQspJz
igtLotWCYqzixBjU8iOJpsdI9kwxe+0DUZ3Vspf/Ds1TSg1FiA7A+lqAjcTfBGC2
98Fajy9L8p+o01st9FMP8ECzDnOa2FSJ9bAEwxSOWm1mPn96eVIGJ1FHXkn9rX5W
9MQz20DLr4ighGaJns75exzTh30U9m3LISMUo+yjdbgu0foXaUa8D/xXkFrg8t5a
exwgFiIL6wG4SMR6O+JBEK296m9CdeYgdkN9EPHFmdP1S/sjb/PKtHqCV2T34S1l
puzaDK2PUJjKeaeqiUe7U1JSuHZhlI+3WylZm57m+VriUSWiCENPGMHhIU8QfflA
EeNGzAbMtSMCPSTNWX22K5CJqeFzd+StTaHDS3sxQ5CNPD+xJf2yz3OM4PXOqDob
k3ULfbGnsVrVj9EVkT8YBTfwKrSAqH65hRC1wrJ+euTvBLRnJTzDxVksKz32GzYd
KycaeAqGujM+faXGXvldqZYeMHkc66OGkwmpCKYImVLB+4L3QexZDXH+M48Hdv8o
KgapVMDM2dR/jmA3dBH/iTVLiPcnxMltw4MTb52M8m1M2XmnAkz40WSINFTh5C82
XpAzE1hVEjOSlu5bjhX9SNedH8TKahe5qNuCZmvrPsDRzBRlk0VdjNlMOKYKC1pE
mI2WisAFbV6wBs2Puib3WqB3PmgrUq9o6GFPAdblTpGus/fDt7sEdjTBqpGLq00G
BSLx/1xarDwSDfchn0Z6u0rlfkIbcpe2/TVZ6c01fCmZ70UWz+Ac7sRU0WuiHqHf
LT+NVqUMyvU0CVIU31/e/pOxpP+ESh57gVUc1zvaRFN2+KRWgNgoLxDSopNuS3Jj
4QftavqUeRLIVWz3QUcxQmy+Rzx1DqbSG8rtFWamhZ7rxqObadQRPmEtQdgBYhd0
Onc/frpkE0OCwWspK98Llxju9wu/+IkVaixJGQl7AqB47OSw0LvgsJYbtnDbUztW
Z7jianepzMuuBehJx0uBCTgqKI8ty5XF8bg/cCaG7VykOO3kOpGPcuAZIYRKtlHQ
HidIvx+Y4vhrt8fdlMt5X781nkY32Iy3GNailkJ1WjzNspSZt40duMQ+5IyFi/vI
8znI1mJvWnG3PTntGy82TlYxi/MdhIIYKrzcmCax9TwnjRp1gGmVqOoAMfSpe94V
TJCCvOz/SIyxQaCBsK+34+lVoyZxnVeYIipRUWBsQ+HPCRsd7aVWNBlu/cQ3KEEE
oWmra8u9+BNUjA785vZozQgz4GZQuv6pxs6j/UYJhe/rkXap1fy9ekuAwWH1/pLk
fcEblj9joCj8bDtvX+t1kKQsvAUf1vKNbFcTXMKnDzYWvYC/KnavFSeXRb+ph9dZ
JMqQf+KvclBg5sgvddrTb05JaaJ/Qkg20KWJGBX6lN8=
`protect END_PROTECTED
