`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8bGm+ic/MRH/S5tNkMQoM5WBZ9VFr60UF5A/MHXfyPEB8cf4U6MMMnJG1LKvZwwv
oP1zNAkhtqnQUlnbIYiqhFBKnZoCiYtPgF0Q2tgu/fA2lhO05+RSkAwcrFXc8FB7
2Ln9EySP+jiO8q6r47Lu9/Jk0HWjh3UOSed5tTHUgxA55+owYyVaiBg6KXReLTGA
2V/TSZN+ql07aJ2i5Rp5KF2ziqLVC6zcZcbABDJ0mO1MNRMmhAE17EbkQUQX68ku
AtUc8fv5zF72114jtMwuTslJM9qRoM/x7khyPpw/7uJ9xP+529d73CRdN6kJkIE8
IBJ9It5RoSBfjauDK3g0yjC/QxYLuhFFClQUDgkY+4CXLoNRX1TWp/0OzPAn7AWa
/Gv/Icz2Ae+3rW0RriL3K8xwvpxNcT7IVX5NnTGzBtSGCxzn0uYfGRTNDnYDS9aq
y3v0QxzSXrMxXOj206nc455SgfbdZLNibbT5tzmR0LJlJw4nu2Fax/BKZh+ZiUxq
wckzim6ScTdMp9jKdBQduqnO2hF0rjE2M/GT1DohtBzC1lfQGK/JbMeRhNUL57g/
KbrGS1EomRnH6JADqxKVvtk7qxii5tGlmofOfq8OD2WpFKzl+mnnQKqXkm8exoSA
AcVGKna37s1bMaWivu3WoH+Mu/O6TqT9mPG44r0NEigrAPgMZgzx3r2pKb6Favqj
yvwPwO93CMPAhFkvklvbmlV9BpzyYuCSv4yOCqUtOo/r97rUbPcrbJEnJTx4fT+6
WioutA8N3XblY2EQ3Nwc7X20xgakNCHvVGKK6zqQ6Y8ofWWq8/g+hPTcDwae4KDx
E9c34X32zDo5BXvnlT3cf0RA8iyF44G1BaO72QwjgqEzEVtRfwn6gyVmvFX7l3eu
Foc2llY/+nLN/65TcbzQ9n2nv1oBmFw6H3hKeJq64cG4lHtpl6AvEloNUDGG5p48
drOAEGOdQGTFOYHOGFG3LrJumKgHehy+RanBVhkFOc7miFQcer0dnUgKZJTANwC1
VCfF4VJlLWdA+KCWtlPhmggJknK+W82e0TVzyCbBdrYi8iiRQdHJfIdf8V4pxhHh
OoC04VWhbLOwuHV3+sBlSG9sDJguNB2ssQdZ1he2ePkglayIuhI+biGXtXWuKh3t
iuSlwwdqjs1BKDMdYK8+Bv7rCn0cmjuB//CcZ8kG7RURHgUE/JYeypZPa50iYqih
4qXlluBdI1G+NGm5jl1Kn6mcBxIPU8WZIItuJJgQTMjbq6ShZxINDekMqYbzIilW
1s6R7e34TJ0bRCQ4MoFgs/vplXzlGZsaMBVcxqIjKf8HPLF9sIfcj4la1oZ96kQ9
4RCuIsx4Ce0DMmVp3XVWMLERXnKtmdA9dUtbFFbSi6l1cBTNm0uNtGuRi2qg1Btb
kQuVyvn3vvPt/sTYoRWva8/Kf1mLnhrgH9o4rZN7jjsZAxf4h42eMEf/byKH/vEt
9C+WwJkvfsjeRJSFTFQfXxOsRiukNDwY2hbNinj8TQnsVSNxHKuZuNQUJmgBp/M7
jUH2qzE+Vlj28UJQ9TnVLK1e//FmRQ7NjtDPufEoWryONrRKiygr+wTlrRn8LMIl
B07lJC9qmr1N2iPTB5H9fIqxjP5PO6FiFXpY8mdg3yENBGLTSxQC902yLEBWZXm+
c5KPBq2n00lDdD6BfqmIW+GgDl+YrvMfTxL5sq5xQjvAzmJ2X76UG6CHZmRwhzBs
+ZrxtPHHcyQyaYq9bI1hcXMzTp5iHTRgXa7kiPdoxsgMY9lrEwlXj+K26RECNMGY
cvWi5zp0k7a7s21xZnNWQ0vI+SDRhM/8xf0HZt9z8/xt7zKfz8rxLOR+NVwk3pah
8gR2qCGEKl/O1Ks4QfjHrRsJbh7XhDA4BZe0QclGbRzZYIOTNyV6f0h+f79JB878
I5zdZ34a1xNFothY1gXfdQ2dWI7ZfcAxjPat1yyLMPWDpi9Tg0ed+m1phn4FMimh
5UntSDe4tQ4rSJUviLBTflHuOZuxgmKlg7cOqavzAtZRE0LTZ7EZ7sNST6a0kn+r
LEfXHvm0QqmGrho5LRqEvgktqzVxHE3q2sLk0PLZ62I9FscnazkuyshBxuR5AYoH
lGW+swXLwm6zYc6+GiaZEQTpG/ssjxtlqv90n8/SM4Oi3PMoQ2aPzT+/EL8bdgNb
vWDa5IDFJTF5TWmYTj5DzbBrP4z87g1AF+i4P7w0eOy2ZBi08xlWviyHF+eWa9Gc
xAKwAy2WTjDJnORW3jZ8EJcPoH+BfphLFDq5P5HC/EOrRnbSIXgbtu/cmzwE6o+3
JlNVu6+JoLIEcZp6SCvXwBTtbKajc/uCJsELWR/7goA5NvG7JFVq0Ef1BcwOucCm
t63/f8MoSyjtAcLGR/F3DuJa8qzEkoTEAeBhlhYJi665Mo2J1hkqTXP8SmCTTnEQ
jpkMTEfObIbWXTq3sDLhwY23DQzr1+EYYsibXieatUsGLSakIKq6EBlck3dzVkHq
DS8vV7ysEzcUdLxj49mtkZw0k+Jm6Pz3tlrZpijMvakLOeWEMu/lyXnMtBmcOUJw
O6/7+lXZ+/25HKqUxemaOddhmMPrNm4r/bQJ9GXNeKiMnybFI1czMJH+niOKyBoD
fuMcIPVQWVTU2m2xFd8zU2ark/XCyayd1j6NZmbRYeULvZh5Lq1KBHwqBkgrIUWb
DvSkf8f4Bmx6T/H+6iGH6m2SNHMl61aa+ULUxedjoLw0fY0UbXoNs1gQcntf6ZOE
iZG38mqIaOgfGfGCBv3QcTFDaMrxVhcBXbOj9KDETfTj/jpVeqAlSP+TNxyOFMKk
AoN80F9XwMd2Nex2c32iyJXrtTYVYwdC4q1utRoKESnHUY3LwMjn/nnOPgWe5/Qk
adc3GxiuByGgHsiWt/6TRtKfAyJHBhVpigj1b/NPcwYtatuycrb4EAf4rkVYP4a4
Mek4iJRPWXJOFzXwBWzU/7EjDUoWKiKTC25QHRAEecZ2F4BGHgloF2dXrQU/ngQB
8Y5bbrUNkPkPnVNoGJz5cOVbm2+brJ+DZtaB/cC8RBPzw4Qn0LUKuK0q2ouarYuQ
HoePFZirH39xaaCRGfWA/Xq+W9qImdgict7uukix/IIRwEg4qP64QX3KVO9O9/KD
EZJWJb4PbmNH8s4/DKqAjne9jL9kRt/dbCYhQhWIdDXb6/RZnBC9PVPCg1bv+U5R
UDFatMQXDF+7q78CY6ZtKW3V/n4ClUNZ/PLWnIIblw4rZQX0wDKGdlJ8R4czV1Qv
NbevlIQmYmmpEepydPhR0aU8QAYRKnkx1r0Qbk0uXGdXSZJpS/m+oowhfn020ETo
qhiulLKsmWj23S0e9OBhs0P66a7tjzaOs0iifat2CWAij/5n4Fj7hwlkMZ2ghj2z
Cg8jWQgxP4ASSqzw8bEDzaR4TAaSxmfXXJKr1WmRETfubLu0ZJjH8Z4J5xW2lloc
b2dwxjVB7OKYnCswLo10baH9sbGEcfLEUfwf7vAVQVLKh1z8oN13NSfaV088r79D
uCTtYF7R5Ro6bAHxZaF2PcmSsmrxgOdmt6yiIOzAGltv7sb/guKvLH91ULfLHqLp
uDJPGBd1MkwW08Fzkw+pWlWWqI9l/p4g5mAjbdxT4moWTdAR7qVXEk11qqHiRLys
bpdFw+HxDMYrO2TtIDdPjqqJJPGBSXh4J0NOXjBha4TO3+sra4o/A/EI2NOSZ6fc
4rbe1eGTPnfvUhKvKMYgaftIn83yeQYtz9mx0vOZkhFgDSVaeYcPS8nokDCgR+3N
xGMCfVBmf0W4q/7sQBPobqed8p5JvdAwrvGMBZf1mewoq/TnBluQRygl9JBLQjck
p9ODnTpg/edtSQ8BZIfWMZtQ3xfiKdrBjavk0QML/IjqM24UtFmOK3pvNRS/SfVE
pw1HsR5PTtfvQid72UQ1V3S2b8VTtt6DoE9NW3N2LT9bXhT4fRln1SbJwO7cx1/8
DZlZ1ByTTR+EgvzBBjQTZEXdFyP3Bp4PF6yaJN4jaCPHk22EpKe6wX5hwbZNxXWO
YJDBtRAdXdFbQpNCGbMrTn1neLck8GHACNdA5QByTcHaVhDCGxsWAxBe0iTtNXHT
P/5yQ9wWEQ2JJwZ3g/vcW5YGOxuQVrTJXvccoOvl+Lvym+kYhSIZNmfg9LLBrfwz
g9VV24Ht5UO3ZCsd81d1I1ZMqGKYZ9BRcr3wiKyeZ9JAA6QwFab5zNyaXceC/ksC
OfEaiEqKf+B7HzgZP+f1Wg7jKxbUuJi5IDzyGnjFGdT12OoDfW4e0smtkg+4hBOu
9GTR2Q61J4rFWYebd7Ihp9uqK6bN3tv+UujIt2iHqIFVMF0idWmEeioLg9i1isVb
mMKBio7YZYnMi4v1N8ZeJDipS58ZXw9azlUhxp6u8AhsWCir+V5Op18QXoiy/+su
/ys7SCRxB0zdsGMPjdeYxIm1t1GKZMsNcoCsSWdqTtCRe7ciwJK1lKzEbce2r9Wp
LNAu7ReZuMpch+gA6DraWPGWwOHbL8nVdoqZQliw8FHiDSOn5h9coWu4fzMHMNBa
I2AFbiXWHF/X1Gxw6rDItQ==
`protect END_PROTECTED
