`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKq1b14XNbq1XcYYQuymNFp9i6JhvIQ7YW0OZgfQutMRkYtOW+CrDyAS1idfLj5j
EPodoJvRGpqQ84QnKJntBuAsZ7npiYTGx65ZOvDoHFosi2Z55A5v5IANVxhGA86G
b5bJH41mR7/DHHQG5AmkROX7wwObpgopdL5MYn/GAWXlNmxET0znBHOQsiVmWMqA
Cv8qAZ5+/Wqo1RKJsllvzAOlmuQoTkfWwrsSCxKHweO4EzPKeVgt+WDi9gGRWq/D
SK/vID+dDlyKU9Ko8k5DoJ6tJVni9JaWRh1ButgvhxCGgVNc6nMEM3BrfhPhyvqo
UhRc7EFClGKokV3rgRpOO8dTNgFj6qiTmbzrsxj1ff1T/mX5NefvonliIN0qazva
Rfjv6rPP5N3g8wJr0mSM706l5LB2MHq48G4+47ia9mmmK5fqZxVE8cBwf4xx2ijp
JPdXgY5K5eSYmd0rnLEQ7dWe9DICwEYJZXn+G76uHI0jJgGXm9/i5dAcJi/XfDZ2
wd3Hue4+9fswWmk2ZZn8HcywRO4EqYnfVzr0gCmXO3gjF94rmxpSiZGPo3f/TWiW
AU2tuO2d5yZeoA+yoI08retOQehRaI9F+3xppWJJwTpda12/MaM8ahosTLaGLGLQ
dRacjjFKr9LPVGhvtAX1/9GkGONDTGllR1yItGPZUtCe/oRP2shdT6erdu/S1ReB
ATfknNevGY1TU2sMIgKbmrsLCsOmAPS2B6EhuEKb3hyOD+rqxDNHaduTwl6u6/Zp
S8ZOXwg5Hj5ysXyozLXFTQ6goNduTypW2pi8/DjeFOePn0oX2OI7rzo2jV5s3KTs
yA8dzJR0U3oWBCfBv+4lMINAhPnCCjNcwtUOiRZZKCpNGKnsydZAGqWRmI5Rk4/0
iPWNGq2G13O6e0XGW9Uv1oi0fi0QGR2TrvTXrsKdM/vZooP1izFG5boOGjJwZ+sQ
`protect END_PROTECTED
