`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIZox1rsl46dfRspSpevKU0b1RWZXBkk+wdtLr+KO+kuE0pUsWc+v5g9E0KiIAjN
rKZlmezcjOOBiQYICbYoHRS4vzmrziG46WML9RFvciI1Pq2MnGTDchjcT9ufq1FL
p2S+oH7Kt6s9ESuDSMmJ2z6MW6jpQCPBT3bNO3gUs4ngNH72yZpLiEN/zOQRWs8k
gwCP+Y1R4kuCrho37GukqY8Z28wexEexa8zuY7P2IhzN0O5JyTUC4ST6iV/fNVOb
abAlR1FlqvkkcUCmC224BD0Q3CiR9Ql89UHd8Is9hqBUfUdfFtvFZ8Pr8US4Wg4k
tj/O7obv0coWwLQqxny0EgbLDqKOsFb4kpIpeEXRL+2Px4wDAnz8WgAIKdP5PuSQ
/hjPH4pQ7kcdU5Cj349ta7wbtABd7s5NtT+fhnYkBwHSM5Ek80ufFpQzRpzaTmwg
D440en06QlH+t9eqyzBLhVW8CHETKWC8Y+AxcH1o7w38RKPe6R8WRdLWk2CAlBil
zmc/bR3m3tX68fLM3A4DZTEs6Nas+ZWfT3RQ4er0uxQvweTjWEXaPZ299PKEFcLK
BZJmQHnRsJkF9oLi/yPbKegfVb65zOy9P6twQeAWDfmBu/MxiJ2vSIoG8ohUlvZ9
5ZtlrsFYfRJjiDqHDSKbXuR/PpSo3eXtuHeWAFQPkenyKjH8YyjmtcMAMqoM0Wxt
s1DjlfI4ArufJQINfTmB7XMvUTXsvMonKnUPxAorGCoYrvJQtA5t8o8tjKBRRCAV
nz3ootN0q2ymfNWW7KfYe6CmK7rQhnwl4kySGe3jp3WAOiuohd7ypQxor7z+o8Qx
Yioyge7XYTWaXIzCCO2wNcgoFi0sCNxZLJd/2WnpIPe78zmmvKW5iGmHYASATl2W
zRBa9dtKy2qIA61QNcZxNqEivpesZbxYEAfN0mz1u7ueAYfYJhMCjD3rQnkL96Dc
Eh4lSDE5T7pgakD1KtoIpp/Qtlix8IHP4qZJ9LzgbfNOqHUfLvi8NpuY6x7FKvUU
WCJRTMjkIBjpUl2XYXSpiBMYqs9yaTCbzrcpTGUE9hj5gnrqqL9zjxi5Uj4xoDjS
1lBvUyfGdyTgCGKs4WOd7ztciC/HikcDfqlKbP+BtBhpXEAIyIUkC+zpD164j9iO
ukoednrm9OkMNb6qlF9FQ2wxqay4vRiTWmhZdeWdTcOToRZ0fCV/gXEJweLx4/kD
zoiECaaSQ/yMa1ty9Vaz94avgiJilIND6xxpPn0E5N6JMswVkKEFD4eZzvWLgXFO
mfrnF1XC+AQCqLuUnnDjvI7qTO0ZuEnLw8ey650YmHXwNzmPx2/FXJHrktYcCxX1
nzj9W+FGQZoCz2uc21BZjt4iz3cWsG6MpS136Hfw8P4Dryr7lstfMAS/M4uQqbux
2EW6q938dqHTe5/JQPTqVVHoiPDlS5syOCtEP+0jP8S18yLo6+qzqb46DA8HS289
4eYH9yIg7HxeSg2tGaFicrQxJYAj2wYP1dIEzaeJoG+13ivlNm/ZMVZQBOw/Z1bJ
68yt05Sz9e09k/u754VFRZwSjEkivVWp4XRXni9CtKWUYIu7NZ8cBRuc399UAPvO
a9gh1tHsoTsAz6KcpqDNr89UpSxlKM8UnbeSeEXe8wHOkeTU1XybLoxKYbg8Tf09
rU9XVxs2rya/jByUabzAFj+/MOuo3hJdvidEBCeXj1tVV3CXKRBvsskKYHgG9OlA
S+rrfPmnmb8yMnTPtnu8fSso4Pow/e5PhDA327aHCMeyNr48ZZSYM3+E4ez7xAIb
8WxHwrPUGIYGkBdz5z3V49FofsV8kjgrj4ETH6v70ou4TT/FdNfUnFLeozIWfAeo
yX+GLJEKAw3xCV3EvZZONVvsvVPONKu8FUuzuzIDWuArCoRrMfAmQ8c0kz9RcJl+
ZPotlmsb/twoR5W81L4UtRm1DnnAV7ECW0TY3Ykrhf6l/DngYAwoWpFC6F6WsPMf
K6H3OC2d++yuOPlX7g5fNIDqajuuy0k3JfBJ8Pep/nafNCfIp7X8VVxq1egIVLoM
mh7HrwjUx/bvUFqZi6fLzs4eAR/GczcM3zVlLSReYU2Mwj3nxRLASIFSWyddqafF
dB/jGgcex8WSMeJxD3hpgx6/toEDenJfuPMh5aH7/E3a47afezycXA0AU4bgqm+K
sEnrmIq+DHnLU+dvVqiXD9QkIEUFB0KSt2IiecA2HmBdm1ncthbCBkBctETg2+23
yaCj7fWNMQE4T83X2eI0e/y08ftK7jYOuJMfnnKC5xBfq4thaID16+sDuokxZTNg
vU64eIYNlGXVWstI2paROW1ITgHIf7uSm1mQ41LM7LXa7b2bGWlPj0NTVrXfm57s
WR+Lzc6d9qK5la7QBqA31rokhxb1Dt3nFN5Zp4BCPCjeXBc9m8xsvlMO+7TuXSnj
SEMle4ZSzG9dROSLXr/uwyELY1EyYH6RlOoYZQR4O7gDwn7PuI9tUMlTrj9cT9qC
8cQsybY/ovFiP4THdmwMYPkTF/jtUjcR5Ai/EkLtXjtf34F74gUO059tZGSFedHI
7g+mvAur+dzmToiJSXid5UMBcU2L+ofWlmpikUjdIuiwbfG9o8iTJNg9IhCB10hh
yi6EhvKDMaMVEwYPcrpVEzraOL+A/FKCO8eGApOAwXQMaEy8wHVhysWHmzvJiblC
McYdXuBSqWxKWGwzzCsmKZAVvYEcm+95YXVbe42BgawDy9TGA7kF+TX1/A5FNBVu
WPiRnKdKXCJaruo8rOkvH9BQGRdr3Puz2IMk9HlZYN9eqcW+lW9vJWO2G0uN0oLH
kOdllPYHXWLQJ+D4XcBZGHvgAqHil5MlBpB/KOkN59MfvoqKZF76JWEs3OKOsCaO
xhnFFQNASt0L1t49vvI9BIaTskJ6qMNp+P6gFrQKPLJGMKxRK7vfu74H5Qj8brOx
rtIFzxmuBlmlCOrWiMp2PMwzCfhrP+oFBFA+decFJX4weP4hSQ9H03oDFohnzidR
f7jgfooUu2RjplB/9rYViUgnVKbVaQBsQmJqenpzGVyh47pXToq06raOeeCBLXcM
GM24+dOJEi7VlTspsqVayISKlCz+WZvnkphOc1cJZjXzVflcGkH5Md5YXP4vgnsP
eZTonaJEouzcUovwRqqa63IyLrCp6nfXiV2scYQLuYrnwa0PADNEda1W4SQ6vFZ2
Iga1dn2qZ6mJk4fn2L059Ghuu8yKk+mx/IMqiWBYgkQlaIiIpHCsARdHocOLn4hJ
qO0Byy2MT0fmrEP/PXkEBnbeCeXk3ggH/qqwKVanckjl6bMq0Q2YgPeHMTGO4Z0T
DsSBsaRJZHGWfv18+MTzMzsuKwS8Laf88So9iVf8OVCM/QOiU0Epm85EpiZdlevP
mokXfMRCEYus1fyUz+HLsVKbf445ytMwxQqM4AwkopNdluhymalmUsteHLCmYGI3
X0+CbQjpACIEjHcMRKTbIyGeRl9yCX3Np6SR7Idvvw6u3Za5AfRPX1at+c1o8hl2
mnG6nBhGwbFbK3cTz7u+D6x660iHR49n+ONUDUYMqOLtETOWjF6HtYK0Xd29l/oq
KNQT2X8Z9PhgJ0kdoz3TjC+AIDxEA3zHidgkYoCyckoKdyc3tb61gSthB3D+NJ86
cntQoSt2KNW3ZlKAuKRTrl7n/qd51MYbfl+xtYq4gl7MK5jqZuuWCFbNBIXQmYbn
PyWVQwA6pg41WycLfvBUqJSBAZLfRNqUZh2/vmA/MA5AqyBuSizEOz0GNZylf8LW
x811Wn3vjdhePtrhDx71Km+x0xqcw1sdHT+WB/wShHrmyyJR62lO/A7hAgt4Hn4m
XZKrdK8Rmp68K2Ojk0R7iIg72voSlvvNPGD2g67c8yUnpg+50Dh5sLXq8X+PFbvZ
dwr/fJUu9wBycmYEbIUSEBcycazaFFoHX5HbKtvzBuanqEGNOWAG4ZOsnku13upK
sga5v1z4CmzcqmVgDskyFiSLkhTopg+0lA4t4nPv5m+KJtsB2vb7FQWFRDqH5Jg6
xgxDVUXVRFwM1aVApL64yyb/fAFO8S809V86vTqLJQXq/XYNQVT6zcE12Obe+vnG
Y/upkiPJXDEwhrgHo+JgmPkkPnrPlt6zTpIJBTE8Vs7cfV8F9pcrO7+FEhOa7JRH
T4g8+EiCPrFzdWDFkx0ZYoHsXb2ycj/ac/UBfWAp+LMPk5RW35iJlW14yw1ee18K
5R3KRXArDWxxJ0BdGeSLvf86PUBJGBWG9a+sB0qxaW7m9aRKvuA/myFnebybM+1n
36xNn2NTDwqK8H7ZNqqMxkX2stH41jX8JQWEicdDDFP46tcSVoTtLZ8LUCyqJGYW
PjyzI5n4kv9ByHBnGlZpV+kZO/XAfGQvIEU4Mim6EQ1YzFeZtKbr5ksYHqdGH6jc
SbT2ntWRKy6+KYifUS9B3523vlfwfdpR1WEM+olgg4gfa6+zovVmbM5yoUII+63F
EJaFbL9cAQ1vo/6A1oBIGZJmiwEziVWbex/g4mGUjGXiXMDMrELm4ikpoCSmbS4D
3IIs9SQ/hrGhNXIqTQ/f8gnCJrqouwH++A6vrir30dN8W331RtZ6DYT9eT/k8vm2
iSyVXc/56LtiYgxe7ETdJXthCUlGuhzfhYZpANKzCGDZz5h9UZp1acdG48PaYek9
Jx7rZQQhsjJ8BJzBMUSKepC5y3w7wmYwiviYADDmHsU8/tHHSeG8yL6fMlFuh0XY
mHbh6ibWXTK3j0uKLs0H/U33fX7QMT7aAO+9a2sB8cSekrZ1ZYNtFJPxthV5hkwt
Ulu5/+iq0BtkBtvQ8+hUtpR/7YW2M5EMqv6zkDnBdYFkmByD6qalFwdv4/BGDtPt
Fo4Jh24yLtMInI5ufSMUNXykuCUD4x/SPYYMfctYQeWiwIYBF1qiLu158NJzqZga
RbbADu0ZIlPf9+/vbsTHqT6SaoNoTGOtRmX2IriLQmd7L7fK+y46tNFxXulP+ILv
O8vYSDynbjTOfR71iQGjQbrgeM4tJmi6ZeAdwpJmjUSc0Z5os6UWynfQr/ljQt3D
HYanFzklPmnFAjPiuTponWyzGMAX+cKnio/awvC371mQ4KETBh/Bq+6lgidBj5UC
wVwSAqd+YAOCUeHpRX0WNYn+2BYht42uZOVZ1R9dKD33KbXuLOEtn4pJfkotV2uG
NGzjaqzy+E2JN6lRKRu2GZ0jJj0u74Lbz6nzF+8lLK1Xsij/TF0+Eqd4P/lN+ljO
ma8eBxD0NUqn3bFigjWMYAZoZeJ0Z36DGANZvuSUjwqSVvfQVM0Ht4NyLjejNcC+
wRwK/A9vpWV9bESsi9/orVDIs0c7SiGuXZ+4xQRoqP3ZPfEDcDvWM5XqL+kqx00Q
qM/Xl88ZhF+P1YXiusaOFP5SL7WroxcrdzwcewC7Cc9h1jKK1T26lHdbJ7D6dZMd
TgHRPshuR098Zwm033PoBeddtrjv6EB1UtnFbit9+d9UHZWyCmF2oFQVR/CNX5Yl
idsPc+v+h+wXVS+b0QfeVJvrjZnxyU4C51XHAd1FC5z1L0R4dWABNDLNsZY3Dm7C
IfX56iru/LXDDEGq3y0SWU+gr7OtO24Tej4I6BY1e1F3g3tWKuqAjMrA5CrE50ub
+dcDDmbQzAI7OoW+BjS4l08VxUhvBqub8TzkbokyztvyKjh4mTlQegK9vl8AHbss
VybKrVyYuJtvJq0vj1LjQ1kMVtZ7ujhhSwF7Tg3wCJu9VVKQiI+N0l/tWhi3nvmb
PZLUdafLk2tJXTkTZqrSr8wUibS9tLQDmFj8O2xuuCtYKhOcbOX9snOqQ+Wsdqt9
vQRvT9wUb0YV36P/4BH/2tnMP8UMGQF94h8eO3/7D6wQzcpKLNCaVS/RW3pA0cOA
tcxEUeweKo+j8uBHJTS0fXaXLPANOxtTKLw/qfMQFdF8urzal1w6No2SIFJLDzib
DgM+du1XTi00VRBt5UiLGPltzl/JZLJ5NciKAuIHn9/HWY+z8K4bglJnKlLLk3Mv
mWP7vGdUNvdIdDLLfJD2hGTSJT182zJ1ySvLiiNp8XE9vyBjP1BVsSzqHK7I37/c
kgjNy1YRLW36nLJe08HnIxhxzpRniiYULuz4nmwcb2l+GIop+zRU67tEMqRjqfZP
27gYcE9Y2dnwefBbH0x3t2LwmntJHkg8uBg/q71BFYmrMYWPedHf4SCAfFzdjQq3
WHjnuA3zQiC+DfMlOShiF/F2FlQuw/mri8L1DEveJe5ktBCXwAG9rrz0tpaLkNZD
reZQmoRBc741+xZGKxGDyIz2L7FT0zxtCTuG85+TEGlrD0cd12XUGDxtUXBc4MZ2
A7ekdhU4Vj38+xQz1a156j88S+lfuL62HRuLUCz1PiieI9DwADtJIXXcmxNzPJP2
mTjLDyWeQ1Gptnyg2g2za7PO5pVELGXz1fMU09L0lbt+FjCv4DbswBzbRK3Os3qz
MrQXljZNePyvtDx4SK5htPArdU8TPEMDFyGAh4BYxOpJ+iU3e+/65bsS5BV5YU4P
zX79jRCC7wshO83mK0PoXwj70vqsrA6cxbj4LqKzK4b078Jq5fA66alAxak47fud
FK7RMrb2xryndlerzxFzGisXvrD+LsIqxm5SwpIvpR5Rh/TDosH+CW1zL6a6EhW/
bXIoBmqD5788kyBe4yktll16ixiu49iR4Jb0wyROiZ/IvE7bfXxyKA8dQ6Ndv+/E
u1brnVvERS9sScF4m3fw91tdUNF7FtUp3KY+2AuwKNDXxZSkLO23FlVXuKZ/pb7A
CWJ3nos3inDC/8MTWKb1WpV8qs9JVd6qrJV5ev+J5LocJ1M0U7qfeWXTNL247wSH
RlQ29JyGRMRAjYJ0c89yk/dZeQ6OxLxbdV4ldUVD3k3d/x0CZDYpkB1xrTgr3mR1
D0XzIPWo6T67hDo7EDvCAXQ1B25dMup+Blz4v4TK5ku00nOLxDwc0Hclxinql7fe
DohePnFGruELlIKiWqu9J+gxk92rMdY3he12dzTVskRW0jeu9pR++bbSQR8QRyTN
hhih6elsa6j5zxlJlSWcJKxyZJJtM4rH+9B32+D7mJx6K5Mc3hU8YuXhfrCwXqoJ
dsHJzlPVH2WHH7Dr89Z1wAwX6+WZ8Hu6s5yUeLT18BuO2oPQofi7elP8ULFTxTcy
JYt8CXyB0ZKidR5l4Wv7CW7odBFC8y2IOlevdxfwcA0v8V1nhOTxLIC3hk+8f4Ge
hZHZ0nIQN+20YSj1QDqz7OjQ4xs3fBfD/a2RCOIxfvly1SwCZu3EOfvUogz83kX2
HPyrplq7K+oQ1GOXSBLOoIE/hYVcviQk835/kc3RQL+xpbCPAOhzXUyNNZh9tUzR
V5CN1UqHyHnw/z7EUU+rYptl6qbQo1fvsje0IuI/50vbh+LRkmxlUgjeXBv7HuXU
QfcfWhdkr6PNx39125W7xgeN1mlam7OHOhzNkkr4iBdXFAhJRul6veuRfJJS5Um5
qX9iyE8VH3t3Y8MsYoZ9YXKPBm5B03Br/wj+riT1EI+7hvyjZz1MD3tk/V8KTe/V
9FimdMY8wvPd+hTXAfgtFFmCt/MH0VftFIK3arliQFwboK+3aBl7OHHVERMUUFAW
RLTz45c/z0M2Rn6XRsVcVuvXS1gPPsbf3k7FmeQrfMAEzmTfEMGlGGMBVy831UT1
0V+pGw+TyCnA0UpKNm3plPRGxQYc2mjlihvKK8v53DqqtMbenmF2Ho/UMKErd10W
ZO8jYHw4ekc0B+BVq95vV3tXeUmzIFZhuHuLcUBN7M0wtQGNJWW9Gk1hoV1Y5J0W
Rgx2AAuqntb2y0oT2dR+rbhxQra7n7Jwf/3hz1E1T5ivI7JZEGTuvgolrrRdDl56
2Pv374PrZcG7v06X8ePUj4JH3w3K/jv0vtjtKpegbKw5pOovUROdcJpEz71un4yv
AySXem8aH1c68Cbq4+35MHBFgb7ktrqFMgFJF8RbfklT+pbbVbk7xV8YJ0lrjB2Z
juZ2ehgmKziVqTFOCwaTT377dAR8XlgpsP4XgzrZYBSJv7oTGEhl7Em238X22N68
kWKQ4ndljKgQqsaZVzms9sl/uBqq+6tFvaY4CcDEhKd17FY0y3ZQwwFti/PcBlaN
ihKQLjXIbMR0i193aIXoLqxnH9iAljKuVerJvkzGhvWqzXUJloY3Ykf/xwQnlHi6
ggDCNhxvGZCvhM0INpL7HhD1HMRAoHEA7YM0lg2f40xnzqgHsDwDDjVagFkCm70r
eKsO3Rw92+xcC72xK42eQwUpuOKp18WPrcj10wg6Vet/JNKXDnpME6Gb+JuIz9Je
ztN/TUWzkUt98eYu7eHRJG/daA5eFGi8K47LtiIHfbKkoquTD30DZcZka8TVdCCE
V/jvTBIX/N6Nod8n020gk31uYqoCTmuExhIJp+UDnWd3iAZWMrERSnUxC3kN40py
M0mfOyT7oxYVjcCqaAT6TF2MdJSQ17S+W0pgXXgGE1s+/6in3ZBc9a+Cw2OrrFeN
bDxvZ08PcNNwSJRGr/jCuQ8abGWeOcRRoU2m//ofEMOcA9uwmJGrmNtpWoF19Ca3
5TbfntIrxvqKmt29EpoiCtbrbYTLpQVqKSAEWvM4+Mv7h1WjGdVazXjYbwc05hcs
GI5F75vgW/4whXLMeWOU1vj2FyW8j96pBntCMj6UtgmhodNPO1DCdqg4j4CENJrL
j5FhhkyumK6LHeVetiHF/hkH7rCBJOjVzc1wp4r2SJmIGRMPrzD+Kr2JAaMNuyY3
JaxRivD5tien1btpR2Sl7GNIGBPx7BUG+q/zKG0vk5NVVYnc9mbTBlXe+clMmgPI
AuUePGGxjQj7NVU1SoL4Ap7CXh++3WKX2NAPle+hpimhNMouWj2Z8kT9WBBLtTZq
WCLlog0o7wsIUirdKpAhi+BR0iDpTaXBQWt+4+zgE2cUoUAHC9FFXwT3zEI4Ri1x
/7H7gdIh2rRFXCo43h+rNulppvWOW6ieXEx0V2Nuif9rt5senFZvA93CJ19UY0VC
RWBLKxjewkU9TRuNqJzIIcm1D1w6fzN1FINIV4vJJCQ7xMrNSepia3cFBCYWORWg
iJiBxYkPeMklTZQdi5hkPC5XNxxz3jO/3lnKVNqaNhQ4hN79QpeIruO5DiE6dfL7
DeKZxyW3R3Cvld8x/DaP4VQg8Q7Cm7xh14HMvNmDK6gUOuDK6+7bKyexMUUwgN/O
3MYvVTtwxXW6Z3sLBdhkAeGrNNVIeEg1Ac+w3Ei39KxVdKa7IdETx/nw6BHw+I1l
RaLS42GhZ5J42pRHhB/JbxtOMJY8TmVu0Z44og+W0Hh6RJkTg0oYkKWJgfXZBR2T
YS2zenkSXAYtpxTtmzCR5Zh5H/hBkaPDephKemPvMSQgTKhY4nuUfrYpc0nYb9Nb
5j3k+fnY+Yi/6y7JmaW87yQY9STUtXuCfZ6L2L4R0Aos0+N37HyUAXpx9WUjbYgW
O6GIgUlwffG16M4t2I07c2kWWEBrH7EZuWfC07+9tj4XXN2jAC1p+Cn9NNkYAb4/
qME43KlZyvuSMUXDjg0VYo2GNue+db2oq1pWyJnbTdbiYORPj66M/aK5joys8B11
DIESmaj7d76huCmT4ASo67l8aTesE08mCoSD4HYaMI2dTxxZDOEwrGMtZjbzQuil
NaE8wESQIBFaJaIL2cHjN07a2OKbelvyEOuPIqhUfME5kpFsGSiKEVjk4Ley3D1e
p8NGCieMS0DBKh3BaGgOF97AqJ3i2L5zNJFMtbVqBIjkX2yFiVc86cE96BqSWbP7
fDSVrEc0O4dP5RcmdRCturgGFtADZzq9SkbE4Ivubr3yst6cW65dXuBCmlkzb2pm
14dTSmCcy7SEbkDdNdoOMhhHbKrhbTfCHeSxz9CmBB8serjtm19evLvp38XmbDPS
ZgYVF+lDmm0w8dtUfqcZMS0lSj1GGG7DGJXdjbihySsplzLMi5/rQVX388NtfYCd
as+bz80U9LsmeTQAYhLwlesmv2uaFJxRevQIoA/FDKpD58sdWnauMajPg6KPvnJT
1Zkbt2ADziGIoAMIsSVRzUjmACqB8RChvOnkdhBkqoQM9VQRGnVp08C1i4UUebjH
PvsJpislTK0pkKvxUugB8S9s+PSQaR+K4GjvAmymfvCHKaMgMGU8lqBREqvqRDXS
vYQ4x17KX+vSR8IqeJKn8NdaDEaJCkoALm6FyOupag9V7Fw1Tp2V77ILhcUYccQq
Nwf1lQGU55eswfhMxgR+f6ToAE3zRjVuvBIR1UpNbvhkRQp/3P45QOqvnKt1aD1S
tPNBSI2/r0oibUqMAH+vTz+kS53PNeCXfcbd/Z1LGKTM/4lKTjm1Bvd8InaKqrqL
6/OQO56sAn2Y3Skc7eBkka7b7GBeyOHNE25xtF3doXkbwwrBnf3aEdkdDOwdre3A
uP1kXsPClLN7eMFrvzkgocPw/baOYa9lUZt1jMpJPwXpbi2ujpXjE5Ms6TAg3uJv
bdoE72kjePpb8xnbt0/KM0u8t76aCQS2PEuL6rc0NtZtpjXlQ2e+EwBXwmZjdLpH
mZStN+Q1Bal3lRBLTKQjqfQqtrKa8Ss0N5fbCcwzw4zZpjo9WY3wgYKlel0ZWGLi
hF6fiGCKfqLtOs7rttJQY2Y0GQwcZ69IGGjbGs11tH0NUuyuZbZePLf0i1Q+9r5C
Wzt49/R58Ft55BxCTm/1wqT5CwNmGl708IrfZceSN4KY2dGjyTQTts33Lk9r5DUi
8lMHe1vMyKvEoPaVfvHtGyKSEEoRze2K9Kv6QBWT7mU66pdzJGS4hh6X3NI5XbE1
PEb7NW1yslIZv1o4arANEIs4FPqGdCyD+7hwjn0yCZGCZ7pVbHM3CP8rW+aq1ZVU
K/r8ah/O2Q6J5HZJAzEGoyRiQAAc6FcWpwv2hUQYPng/83zD1/UIKRLTITjgB+xx
dG/rLR3q8xX5fjblai2WfOcMsaLbplH0+mgSS2/MBgVpsqtkH67Tt6ybJ1LlpF5V
UeQ0hTF76QYq+VktQRiUa+Ao3HnpPektQzMiCcW1znMUg5uYARoUF80VYzwWyIBx
y9cz32P4PicdMkbD7oxKwwCoRpCV3CtcTi6tMctEZ+Tn+IScBC+gYW0drDOzootK
hJrE8EUqrpdbcjg8YXAbda/i+O/OL0z+9SKaXAiixL9wCGZCERueX+akeWlvytQS
fMhjE5hGikyAEbVS79nl7undJcJ06Znp1h6qUrGltoT2Dug7OqzTRVLGzKaNZg8Q
S0kdqYJVrGs/og0ZsGNP3toytDqhPTzMPDB48JNNAQ+4YiNbrISgpDwvM2tby+rH
G0dhG6gz53Qaoj+3F3lmVz1wJSLQViu+b1Sqyc25UF68lttOypfwNSYEDs8rXrJD
i7AkUGF33V59Q96xKGyERCTIBGko2YjLrpg0haWtLM8FM8glOH/AKs6vGs06BxYa
BDmtvMo+W/Xu6QBIBnvJDy9Hd6NnNdojnOdziZXGWdLoV7zrg8STt5uior38g5XX
NjQxa+eOxGZDkMBQU38MpPBXRJ2gKfY0ZA8PBJiw05PGQ5HhQ5/vA0k11WiIa+4h
kaTXz0LBaVeQRWtegvhakF0SmCnXfejG1mksAdvIw2GfPU7LsnWKv4ughhQjU5WB
ADI5pBuvO7lbWqMk49aVfl6lo13KS0mv4HUiZRkj1QCm5W/AnUoQ+juSmQuoIVQq
GJDyGnUAi0C1LdyrPrQwfQ1RxO8/3PUT+dJ6gWyEj4j+vcvhW8Y8rqzclbwkYf6R
lHdRvBZhVDT3bCjiOn8AhxnbFS8X/L0+KByrAYyIvGn2LmaPNTVgEMuWU5GdFw/T
P8q7ftcbYYNr0A1ZtwIXA6aoUn2y/zfOKbJkxdFnK5qIb0giV/J4Kj4vgZV62SY8
K9zZ/Ht9ez+9w4F0EX8EmaD1/z7I1npDNo4ZxF5oAqgs7EaN9ovqgNOqSstm0Eom
3LcD+0UHitrnpdFJnnJu2bBxek5lWMjPwczA5H7BuD/P9tYgLKn7GRTCu2SgJQyi
WLGJY1f4pKosx4BNV8RxErr8gUNYCd7puuQ27RTgg/fBNEmixD4R/nhO9i0/UoBE
/MjNwlZ06Y6SFtpClFeKUrvl5+tJ8Tr2tPDngbOBx0W/iKrp3uuWyxr8WVYP51MJ
TciR1vRXdoQy9itIMSr0I7IQueqRs01ccNslGVmunzKoRethlmHHtySFmj5SBmgC
n6bYR/UWI0uhXc0ejwubiojiJ1BLk/0cFCvQNKpCjFcinxIeJfo8EnWY6/8bvK1f
Ub9quBXkylBwkvbqAyDOO8cXDqLF2L3avqQ1D3nO5d4DSLpCJx8whewmJRkWlZE0
Gm8K9Z/Pf5Mfp8jNvkB03tu1wr3D/Ip4hYqSdz/+sYkP6x2Rswo4EcVhzCkDEnN1
30vJSTq2IPn56uN4QPX2+3jNleA6JRoorOzRKoyREgn9mLwpQJaCkb7QwllqJUMi
RhLgMnAMG39SV+AAipPeVzdMPYCbKCAR3+0Yq/Rb/OoY6viWj6iD2qoyn4iKhuE7
f9yI6uoPg+Hr9Jwt4buK/A3/MsIjXEK5gbEXtSrOB3aqBtNDb51w40H/TUuLCXGw
BpcQj2ICEasp/zv4ddPbvPMw03OFYLkIBN281md/P8qVAGjrHCWDYEmjPygepBac
5a5KfSHsOuPL6hHeUrrUXg==
`protect END_PROTECTED
