`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AMiGCDvg4i/xt+EwrAtoo3XtwzPcjXKkhrlA2N1BHG762M5A03zAu9cg1482vQtC
GpQVEipxcVxxg5d33urmgS5Axs9bRe2cMaxQ8lyExkwwV/sNBLGuOzPaQwygqBZF
K+7eGekmEf2Kra2TBEsV+6jAz9hgGGA3UxLlNTQ6FOJVv+w5HF50irEctQQ738Gz
Poy9fdRR0gLLkNn07MclodROz4B5P5Fbnth6WSjUKd3G8sdTLqq5Cr86K5t+ue4I
lWb4X8zN41FN29M9mlNJMWFVUgR7x8yLqqpHzUPxojtn0RqB97Hk2gPDfqh/HPRx
5MqhBEMNGQ/OrNYjaZ2XaZUjAVePPYdPj7LK/jgQhp4adnrr8F959K/DZQjmP2fi
VPB4TiCJOtvumjmac9f0k5SOtuKtVaTI/89xayDuCG33aVHGNbsZ484bwu5yX21+
TKAt/QDNE0yVy33DteDodk/f7nOcvy+LbmsOCM8JEOawhybKx6c3B0e78SKUxd8i
GIyHvkvgpzulFqbH2He0VONO1had9qtpnMSEjslJceYNz+QmBESbVKbMap0ru/d3
WE2MacnO1VVzyAkW0y4YCzstprd6BLP0CWvEYFHtWl3NJe2rqlpse8b2bparJEnd
SEzAa+yJKHUCRxK+Dw8xjzi641SAEIGKNxhTPie2BiQKcT4l8DU0FMWNjnBjJ9sq
l1tk0KQW8Ro0ltZBzJ9CmfDHoORjOmnZBQtroxc6BaARiw/UX9Aku23gG1ae+WTo
olMH8/tHHeqhoKPhDvcC8R5FSu1j3EMGSXsaFvjk9UWCZBT5AjjI711C71EkjXq8
UKXUmW4GptNp7bClHFJaTonjohpjvv2Nf5zHZxsfPZvSnH8++e2nsklWl4mf/BED
CnhzP3ZTRC023ENeDro/dYxPVRPugteIL6+yWXgX7KWGLgNLBRD6y96ClvowQd25
YBv62XlJUCBAibn9It3uWsTxXJehHrtUUGb4UNaBL1y6E+LHm1pD2O5Dhm2U9j9R
ncYtGklxRZIog/Zj0EVh7+OGBU719t8gSiNWr8D+XWkXn70fGv7iO0UdGp7YyANP
n2w6OP0Tz3Ysj217VDUheHoCUdu+1z62mmhw8gnhsKREum+HdsxbLyy7aFR6kYfi
imvwdTCvwW7fXZCAOu/4weJW/rRmFVvQXg3Ndr+56mc62vF57Zn0r/dGkFxL2UOX
T+hS8Yg2xu75mUXcZ74+uGfm4EIDfE6SS06qJQruXH9ZiFJpDA5kDSGjZJ2QrNlu
62b7/346WAWmVMfokzxhl8gN/gjK8jgdOIjb0VxRyAbxB4KOOTrugzw7Zh20mSYL
hfUjxw3rgrlMo3ty64YOp56jlgvLZoDi67NcMaq6QdOKIWfgM3YLqKNKBx6c4GoN
mDH4GUjTqOCm5AKmT0+3a2WU+84nwCHlsbv8s0/40KjRodVUZY0/Ygrt4DdjdbEA
eHgY3deKyjwQw4PifFnwViutmnqCrxGX+6E8GFvdmTvwX2PYfHAaazjDbtd4qVFm
QbRYqy3aLshiwQrpGVT+8JEhMSwBHE1lVo50k/dcQnzHjoUzK+GEqLf4oFTBpUWW
Mp4tUFEKOSQSSMOvr6zvD1n01T4j2PwSHnH//flPxGz1leC7U43T0NtMTs172sX9
iEcqDuxG8sKD2qPnCjI5UB4nuwo78ym9G5HEiY/8pMOlrIo7IvO4KzWz7PHQrKU4
nhXRuxB3LuV+DGcedP5TJ1ewy/0RRzwMBP47rR31M+EYMRrdaazcjVJMb0mOlswp
C+8mhS8B3IcE3AFLLL3s5a4YYxr2ANOPiDnpOYsqD8/orNK+oJtHIujeqLAUNNMQ
Nj5iEtufkPO74XImDO8m19tIy8s27203AnngKNiALB+gmB4+EqzFU+SRcFIngccO
5xxdXoWG1HquwwBlQFzb4siSjmSsDJ8rKvkYdn9ME38BmVZlfXYYTdv0t5/ThZGi
FDAPJwYAivEyAE8aayQfqsaKUU9r+C+O+tHu0w2LWknURNzx5b1Edpt/J+tUmRII
TPu0MlbUEzcGFTVYIezoPIm1+3Zr3uTgpej37q9As/S3Duqa+38KYxXSH+29N+F1
LcKT2epg4GcWCvXCzA4w7/40tKdfiIPBEi/58HrVOD1nNZwg3pups3EzwPzWJj6+
mbUGrSXXCVQ2dzYMAtU42xZ29Xo35+wrLlcO8EiMAKLW1DWEeywuawop93PNqPZg
P6vlKWa4xZYhcyhwE8O4TW7m/QOfi+PEFZ1Uj69qATD/kRL5wal8asPVYPAbVXfU
KBaM4k06ukgk/HSVB4Q8YEw0Mx/eFTetcZkt4PwKElNOOKOKrdo/Qy32LG88qlvt
anjj4JGECb20UOFxvIoeHt6mT5RX/bXvQ0n1pYL6ZigO72AGz7IGpVXzWu0EjRxz
aN9i1OGGBr67TRKbmh2kdDbpPLyXqQo46QM6XyIjqimKMGZppH/mVg7ppDRuU+kn
HBQ3texLfSlK+uQeBljIl9uc10KDrymh3YfPa1xjFkXoKYfSCdHP57aDKNAbGmqF
AuMx+o915JTcwb6MxmfOdw50jJoic1Lvvaw0OEsshD8u1xDqzj5rphieWGHsla9M
szGBEguQJfKFpL5c+lShpvmItGr0rfjGyb/DvHvusGc0tlyDdQg+qzEA8OA4fB1r
sohHwCdbecaveityQBIOEI8KOeoZpbxtcaerX09KhdryK9guRf6FD+h1bJNPYHUx
Ni4yi6cu98GXAo87naY2sH8+vv88gEVmqJzTOVYyP3lAt1IG8Eeg9EkPaVj2MydC
yjYpg/zYzoLXzsxqHD59y++MnUHMtpZjJIJ34YIC6nyI28xqUL9wNjiEKSV38HOl
NFSb/KHL7RvAGR9J6H7zTQwVCUYr/x//hQ8/bRQp33uMV3WXrwUBs6N6zB8hfF4O
WkxBTXlII7EQJACd4+knNj/AY4CRs93TY6jpfE9ITcNinOrYzjuCuAt/Y3cWzkfG
wBK69kgIcWV0ch3J1M5jqQtv3s/kXw2/9dTfA4ruzDDaxNtlp3+fPq+6hbToSkZU
AvQg6/MeAcP0sPrPK5TW1iVKu1639Z7Ua5QvJgUexxOMKndxLvD6i3rvKRaBPwtr
MnC0C3hZQcvD+wsDienSP6XHq2L6v1oJSvCOnXk4y9LVR/HA4S3PoSZVVlbd252P
4As8ugLi/1TFvf147MT1MRFaubp/FmOjhXilIywa1k4A5VVmCE4s2kvgcbx2vm4h
i/ozyZROr5xruOkAMxi35mNpfYaqtWUuD2sR7kUcUainZ+6IGsn/YKCotARrbZ8t
CwI2sHRzP0KFzaomiMstszYm2GXaLQ6XuSJnF0paV0FbkaKF8Kb/zzLdZzb1NcQd
UrMVM4NtFFhQRgXohURnHxyGoSJMWcfFETYfJfijlLXQM+q1KbwvRooNMgnaABWk
nuksPr/dJgDK6pMf5x3e21MU6tyaCrCKvz5AIEzE4bjjHJGcFKvrYK/xztTdRbTI
dza10jHSHDd9rp9zhZnYYndq7BcsPQgif6NaIV+jxenfifTW/d55ceu4hKJb1VNz
Qb4S+hQcYAUgijl9gsniud+DHDBzEGrFH/tpGRRQiktCx8yB04O4WI6lKy+iZqbL
DtlUds9VEJ7T975xqnbXXrn5rcv3gvo5/UnUJp9D1XlOU26ZDxJIjRYDXPjqvPuR
Tl1ChhOyCY4qynJGQc3pt13oZWmSrGoRVSz+vUVM62BwyGPjZnR/QJ2332r4zBRe
A5CoKO5alWZRlGLavwcxsrZIDZugGKH+z9MaT/GGbTl6BIJpKrFI2OZ7D5hNfKtO
W+xz/YY9KN07D8oAX/MSoolT26EQGYW6AAjHAZHOOM2EUS1Y77c5skasVIHmWKR1
AMjUd2KBB9yBBoHoDDYXPH26R2lpKiyVVg8I2+ebcAfus0Qle/w0iJMtLAUyKcck
nLe8LZnYBZlcXvvRaiXJVcvgDdKBuEmME9hKXIptYr4ku5D3wXphDSm5CIbIe3gY
45lH2tguyzHYOkTl6Uyk/CBEpWQMa0hXWT3inZ2VaZwE5Emk4HQd4F8nAEMm6eUi
ahy781SZ0RNdcAcyEhXlG+J4pK54bQkqDVhgBiirCJ+/1YQhkzkbtT6StvVDRsbW
x/uHeIuz6esmCVh1jANHjyzd2z0rjhHLvHSMwOYnZ7SOmzRRE3yuJ1VBt+EGYHUU
V03WlPCryinQjMeBnqANGWDY/n416uNw3eFb6IlGOvTaWcN/+dxeMCg2ijBp7qIk
`protect END_PROTECTED
