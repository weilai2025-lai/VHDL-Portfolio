`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfAkLstGhX/kd6Tg0sSIdJzxN94kBD8Ig4cN+OViQdOu7toSYrzpVIZ1DdfObcUg
isLFwnDbK3yNLqZT5sIh9TtjPguLhheLSIcdVI4dA5pfGNx6UlZxjXFVc/b0XEdY
0ZvHWpzwUbEC9q6gHXmaHkTOh72ROgYn9nzLkmDUavexglw0WjYoJQIJANoHdHSF
WgbfDHQkCnarUMVrZN/bMKf9Mx5ZY/aIibpHb2VTjXmjWjyHz/jm5PC5mK/peyWd
K+2DWkh3YdIkVk8TUOti6XQW4wyYft8rR/U9OHzMDQhzSe5ETue1oKEMXYcifjre
Dg5oDDUNYVaTts+oSC7nIvhqyYVWQAsUaGbEGRuKoA2/WfQsKu3yS8RCAsB4Ijr/
WEawE0l3dAMaC90qkU/6aUHJBSM53Ya/kKhiaHKKZWvysWYLhTXyyLgF/gpgbnof
CjRaXsFxNlB6A4w+KE5pc/KeoAFLtOeReReygiDUP3trpUVtD+iutmPLaaVcECB4
29BuvGPmoVSm6y8S2k9gZQe5MtgTghFF+vXj6FDiL7dqdEottPznb6YcyGUVsZ+G
jvWs6FPCPgyMoYgLBAeumAYz/m4G9bBQjBrecnBpznBCH1Chb28x3EKvuuPEhaRc
5+5tGF9AQKcLm1oMRQ03JxXb+8UOkCRsOpYcR0zL/kAld7vX96BQoNfZwvruOqrK
27pE002rqoeqMjAslYweID00geAlfYNDzBfT/OjhbEyG27uK3NefqgycEvUGGYgG
XcLGNeJH9VX6PWV4aF9Zoi1JDcdTvFGn1oMlOhRh2DQrn8oyiz7bwnDfiY8oWuRy
SMX+FyyzlRwNp3GkDl+8Qu5J7mVvF7jKIwJz6+qTGButpT8DENIh6MRRIRy6L8gf
2TNfLBwR2fNxNLnu2hkLYOskidprWAYnFs0GiEU4t6MzSs0NPM6kf7kdvr+8swYA
rvnDJiwjlNEQIliL6XhaG4IZzZtBvqMNdUSZvspjcX13UsxUXOudvLPliNJxAVu9
j5SfpIYqnInSlPuHJlzJygqWBoVIcwjtJ6Z7UjiwaOlqx+E0kIGp1U8/HwtHwOkD
nC1StD/SCN36BmUvgwsgiM/4XfapAYtH2pnp01028SQqD5vvW+cKDD94rzhPuSTr
19SrpkfEdfX52H2+lmnX6A==
`protect END_PROTECTED
