`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7TvCs1y+AjUwl1nRt74pCyr5DRRLtl8UhbLz0eVkKiXA5t2VZBpTEk6jV7esQHX
smgA3GfZjTSm1f/besU4wKLZvnfV6RMJlWqO3P92i+oDNTuyRT/Qz/jHm440/uPt
rnA6ixkpECJwXAX0Pph0wne4biLAgu3V7dsL48FgD9AkrQ4a+0ID63ToY9m4kJuQ
MDNTBSuM0+5gC81yPd99aCkhOaIqzgppAaiX0AFvErL9p4TmzLmR5HmQpnnAlM/g
WEsjlh8GqI4eTIv8+0T9BoptfoshGU8u/S2+5UHcFWoqcOa2VDcFOFP5gUzb4601
TbU8hRaHOJu4KJxOX5xJVhdIC5TiiC06rrST+3RucY93DTHcNC9QfbIQrz31xBh7
YRjwTul+haFk07AqLWXlaz8P6p26Ah61/tuw8JMQQB1m7kpSJytOA5YulKI+o7Tp
0jD+a72mGNJV31/DaVKOYmQ4ILiKlqznN6FyruLERzBJR6+3A0y038bxjnLmeWix
Uvogdx2fof3gVQ4OurwmnTYy6dEnxFNgZIVlWrTNaN1WsTmhkikJl/Re1reb8Sbo
eswgOus/i+MnMCpq+VJxqZCY76DIovyCvoT7Ng/lnpFS8glVkis1UFhn0kUshk77
xXwP5nz8JRo94Oae2lNjAFJTmxeVfjnLho2iLzX1Q44FLOKbO41PmOl7kmS8firp
vz0qfv5ZEOfgypP/Y3kF2RKEU+NsEDwQ3R3iMHiqqSo/7y98zpEEyZCKbqX5+QxW
qa61SFn+4Pzc6wCu53VAgjEgWEbATXIShSRsWBUjUrYXe7a9qhQ3Z19pltwxsGft
Aff4MwbwuyWrs3yKWIBrgTqUcc7YUjgEg08gAuK8PeBFGU+HcGAYWBLf74mqv3Mn
E47eeHiLbg+aC2ueJYLH/na4byZFK7XI5ZxG2GQwXznxCf4wXAeAv8H+skTmQJtn
mhVkXn4QeVI6SkG7yR00KvbSVdpz6PjwHs9O0ZUpt7MC9Ziqq2o4yUb9rL3nlkE/
cxjyub35Ejjao4q8NbdYtru0dJq1hWGjBaMQo+ezBqQN7rp9kBbRFudgbsQbOAkQ
+d/BMxzRmrJ9Yt+Mq3t21YzrbX0kkRcEnGNhpAyM92pyxXR79Wz0DPgFJ5suFdZG
0v3gDUFHez3iLiTXEusOM4j/1VoFHwPR41DauZ9uZScy/2qNPSwQ9Yu5FY3IptWM
fgE7jfE1Re89UjjyxeeVMvsiX5FPv43KK1e/NBYOmLHBcwwWrGr43nm0N6FU5Rh4
Cfx+8SHR+pLNoQvCosDgX3Sm6y6hXMKIG9hQh7+gyc0+SSiawoQf0DsYkMVtasGf
8u5+rRL07r22Fef1MZ+EnCr0Qj8oVmWtN3dzcBd//PykKwDWvDelpa2TBLP3H5lD
P7GCKdbyVvyHxiHf2In/U02MXsvUMC49J2e4MLw5KqMGccADL1mef2Nj3BPPbe9q
L8DBL1LWPJigWKRzkV0kh8rUtjS2z5ReZTJcLRQS0k9DGXchVnq2PDTQoYXbbUK8
+C4/VevRN1s49cCQJOnJCk+lyEsFdeecUm+zAtN4RRHDH86PykFmsYH0kUUZoVOa
20kh27ooJjCX3Z/DEgPTemAKdoY5keC/41CVQrJg4JJYe3NyY4EjV14N3y1uA8IJ
Bzg4j6o7pOZm+nm1faSltuAakW2GGZk7ypx6L0G4U7/1wPbr7H/lemWYSZyKIKNE
+aCdoXBnTi2wV5toJDvVOr5TbYVszaIGn8Bs+ATBsRb3MG9Kgp11EfazY9Zl0AX4
MpD7MGUV9V4cEh24N3iv1lCQiE+xSwaEhpRGOjjvHYCUC2R7BwrqFeMR1UxIA2p3
pMvTs+DTbaQ8eXqW6QTTMshQ76fPYsC//Wi31M53t2RZzBaFLfpNgirOeYUwNCOQ
Vvf/CjFLDkWUSc8XtT2n740FXtKR04NOPhtwO2Xn6aJ9Y91skM1UGoLAXuLk3ERw
5wAJs4Y+6Au366B1iGbkNclw4Xk0fykT0aWoKZQNvMkB24c4fdzM5xzF8Wvu9QDm
y/npPh3fLvdA86P+bcjgtlfQU1f10WPtOtjRrNrn85iBUnpz9LeSffpN84u2Xh16
d2ADB+bqTo9gwMXNZQw69pXWEPyN22hFpmZsudDdnnxWKQLgKDGRY4m2MTdjU6d2
aTRVTx2o+I+dAJbC6ns0ldX7ZAwvBSbLqBCdHzmuzan5sLRR6TkNyFPPkq9Zf3T+
s1ccTGjcTrG/zg4p7ouGNrU4jWBzl1Sz+HQrjlfbOhaHhJw/5JKEgNlJCIon1wbF
G2Is0lycxOvVyHTG0HhM/ldtqHPGLp3NlfmXUDNkaU6V2fxFnmXRQdvDC03uXvFI
KHV/iOmw2y0AQMdWA36D6+EzdoQgtXcWYKdwOWWyPMQ2Z56er0hJX40TyWP5mxbe
8bB18Mm46GgjTe6iMP9OO9VJ2038V4BUB32NFwp46RwHh4+EnnZ4LkMPxnYm09qd
rGnZxqFP1UFVX9JOunfdAIfaM/p/qOPcR6BEwPn73ZM/RZvYMuWDC5Iu2Lyd6qNW
uSY4IpH95r74bv/lRnTKK9pNtsH5jH33KSjtKCF9DXZyt8ipgG4GqNlKhiB3iEu4
6AtgXFuwH+Iwwf3keMh5vxRrtT3FcduUUNp0TfSkCdo4XEpUqbT9JvZGhwQOzOpH
Ku6F+CdNusNxNuE7FRzm6S98bWSzEwqihylCD79V8MHpLLiBN+5eI/cjCRrDJSSc
4rLgfT9W4ZtPCbdINC78ZxC81o/lHh9EZ2OP6W42q/L84YuXen9a7Gc7N/sFVTCi
cfX8J2Te9r6Q4Ppdu0iayqHhnjHb4QhhNTgjldjkvx4n4fn0TqzFHr3qLSVyoSiL
cM/OBZPn2vocci5cuvpm6Zy9acNh6syeXEZcUFlc7huLjEQctvMnQ3uRFhMZL/1l
Q3Qb8t14aywXFpaEzkgGE1AGrrBqzCo2kXljoDvdoWjXtBSlGVmXMe1j6ByvOGn9
6WtO4Qg5x8V2jTmLF3CeOv19uR6tRHbg20239CibLy39MJI3Xxvgsjjwsbnu456m
Vl5fpVV8MDhhbpHmY6B2xPeRPB7TpjN/3RVv0ABFHPasmeDNhMNam/zwM1eIBywu
Z9Ku44t2CQKF1/RnSSRQvleKUOKiCq4mFYBI4qcGBZ8H0aQQD0A1GKxtdxPwsAuX
jkLoJtAZY0NTb1kCXnGaba3SXDpLXy0OFxeT3HunZe55pZuDftRFy4DCOzKdqzBY
5fWvd/FodZ2o8KD9sYk1++aoIyvZUErEX7vsIC0cu2q0jqPg5O9YhnMtRX/RJDW1
nXIZ3Y462rYs1hVDtM/Cwc/96T5bvz8YTczeJq30YpZKU/Yc3VEjfNPcAvkSOnGP
NRk9IZzveVNfJESmsR9fipSmnj/ZYzrqJQsOmIDGw9K3QNWAWQTftKOY03u6p+Xe
Tf7EmtFw7uyatYE0g1wRu6n3G6qmMg9qpDRTMRHuB+ThYauD/e91bxWRPWZdm5o5
rPquV/6pzIXH/JMLZeNtu0VDs52ofh8MlOwpaM1i68w5kDbjNVmsCVOC1+SrFTWv
a3rIZdLp7Dy+HH4JoQ6U9VDBP8aPGia2KqTBeZiCiuyB5egNQnJLBAk+C5VTVURV
e0leHL8uuVzKRU+5S2FY7eym6YnFXCiG3kb8o1xm96PZK/2aaJ1IZ9aJiYWNykTq
5Td9uJJ6XnorleVrZEPuLzZfRgq2CgOWkatjJcjnvG4pQVlpEVeKxJcaHWhLlGQ0
Ykjt6Fvjs65MJsnYpOCqx2ebYzG7wGArOCmhvwMHOWf4ym/p3R7j4EpYXnv4GM0c
H2t50DuWmQe/vE28Y0qQvk87ZNO8Vwz3mEkNJcEXwyQyuGWhFAO5dC9qXU+emnRm
0xuBw2CMyiv+lxu8rOALvgBRMnS5sGvfmQrD+yodHqYDlm+0GtpCiVPP1AoDAL5U
LpTkhN/5vakqt8hy/U6PWzlkxvpZOMJnOKhZDnuBq1pyhuf7nH9Y4v1yj0zAtvOW
+/q0v04KSE6/6uSyiTZojHtIF5981DqeTzCTlWFAlH0zx7Mz/pFQaUvLo/SFc6zz
e7IakdvBvydC8balenetdftB3WnoWJ3sqaA+ZDEG8SbpihFvZlwxuykX2L9d+Zbl
hv9vqYtmOTB93lWvbH4u6iNZ01skvUnOi/JkCXZm0xWha60+374Nz6jQFgrGHY17
z0H914lGJ32gcMOF2S507PVlnJBm3bP3UjMU9jzQWmDlTVqsHAwAa3XFkiIDvcDN
OrNsRqLy4vi8c1L5bkn6e6YINkIcDubQsUT1TbGERrNqilb2wOesViHx77Dhv2HW
8Ei5f3LEVJ8AIw7jweonR3RNBy0Bqlvy+Tg63uHO6kzU4UFEcNCn8peuoWIVCrfW
8B2j/RDtlGAoD7+cZKFzBCyXyAUrXTEq6lGIATtTruo=
`protect END_PROTECTED
