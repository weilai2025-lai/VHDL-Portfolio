`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKdhzhlaBmgb5BM4c6R+OwP6pmMIbN8KaE584t7zroiuvI0mqVDy4W6AFvPiWTbl
2HjlR5cdOmQQGWNsdiE1kfdh9u0kFkEXUcMDEjsMiXKyb6ahy/aI/vKXkqmG8YzF
CCVCW7n0vcbmfW5oo+gWCd6P0L382FiZ/uMcm4NapoB4j/NJQl3NMBTyTNLuUEML
+28z54/K4I3AFBckQrLQ/eRhNS/sw1FPkDskojobnIGpktx4IfvGjMYYv+pEiYbK
tXQS3A23zC9HW0Iyb/pqMRcmxA+pzWc+dnfRRyQ2aPZSvCe0TdntYfUcXfxlVe5T
yRtZDXPzWKwdFHNsnQ/qdvupv9SFJ+fZk7fPnasU+wmdAI7hYh/XKoXmmdArQmrD
f+Blp7YZdj9t7OZCq3tOAho7NfckRr/GIncIX8FysDC4U9L3Gt7zb/cJ8STNxKRn
oKwdOUQ3TbkOkhUklUsBGu0Hq8/rXdhMBnLnfh/UkTSkvCE85qboPSk0FIiUzEPu
K7KsFXt7fMAp+QBHxqGIwq2nd5hSDD1PBWTPnCmxrFK+F5w7lfcsxevYvZ/3ebX0
JlJjKwL4HL7oj96uIHeKA4wgOillmNs8BF+ElHW4FLg45jr+MnStoV/DpbILR16H
fgQslB6/060EnYOIQLHnU7ItixhUzaYt8dSRQlDEgC8jWQQXuw3RSLpfzwLqdyoV
kN9vqpr4XqNN/zw4vef+wodVn9EzhDEmKZF0o8d7ObTmytkscos78D4Tf0onmkLL
mhLClGjgkSN98OhQkncbjyJ4cD7Db9PCHncNhY51FJXU0KvxQ6Fw5vl/xUGtWMnX
cq1IEa0cJLRa3z2hIAFjhI9vODeOVZb1s/EPveK9h5292mTF35BJXHJMKbnC6PJ9
HEQrrOWtnKXxTGyKE2nGAKXsW9u+WXKDB6FtcmlHmP8nfGsCP+3aZoNiuWFoJEZw
TEGv5aNjuM8bQKoe1PwrQQUO6JSTL7v0+vVyurEYilPBipaITZW0pStcZfXOq5v0
6qpQDsw21tVg5G4x4lzQbIFOM8v2+dS1ZLFb1a0q54ci9hy8i88IavJr44AxRGXo
RVav1NthYS0yAlZTg88b6Kz0qfa9xbirKpIvesIMPpZkIPbOs7SuypSYYlQppfSn
L1654YaWa6nqRawrzPFQ8kB2ecWcHlsf0Gmjyibx5vegrhcIgvtA9o1v4VXOO2k4
xulOh7WxPrdy+BQoRpEfcL6qO9fYpr5wg6mTXxDZ4W0h13Gz8+XVZmu7I20f6C4z
HGhSQwyGFv0ak0Lj0h13+6vkf5WGefXyPEVnG8mUBncoESGM0ZQTStvfJIrHx8y3
Ok7agUmjQISTm+B68mNMrW2lYaGdMqd9h52iaczcw5Xg8eSdFDaavD63fp2nlPuJ
tuUqe3zLoXx9I1JtMuHkraLppieC1uqJ15ZRn9sMblzeurYzbDFq0Jop7ZU9aNeT
1h/mPZ9xXYPfeUKUWAX4TZ75Yov7bmi1bKRfOiV0SQLGwHDOCtWEOwVP0lgAw/li
47lBDyXlgfn8IUiK9XqGhF+rKhLpgojcXCv9gbLWFFmO4CGZkABkqEDTjyFk2SEL
h7P+o57gcq4LjofBAaDYMLMYwMxgOTOy5Sli7cfo2wXQwhndcgwQvepTzXcPj4fk
znSEGIihQY4yPjsF0Q7qJDME5+q6Iym8SF5wFh49tZe1MKMQiMAHibqTyY+nmhON
nys3CD+3ZeHaJGZba+oyL8hKn89lgCsZNFhvGmLvkDnZJf/+qHkllRtUjo8dJReL
koir09pMM+CFvlqNazZl7AzwUufYpNrDdIK/Okn2FEJUdIaYpH/yx+lW6TpUMqDV
jArg9Joi8J+PUiKIGlElo0OJ8jUTxsLZ+KI+fA+mERhJIEy9AFjhYQSrcr7p4fuX
6KzxbBzErbr/gP3lXi+JU7OMvBjgK+wqeBj9h1E5QxqkrhoyilzgGKN/ZKJk0mFY
/Pc4ODbs/XfZTdgp+1ftJV2k2YWNsI+Z+FcmtwpQTSFxuLhnmmrF6Q6uPjs8irYf
sO20k3iue3I2BgyzKTGkwZOd5PNaY+6IqnPEDh4nZTdhFLffTALzOj+t7FO9a0/u
c9MOBpBYYLI3MGE1K1BKBj8Sip8L2Na4sVnSXdjTCssbFikbJvVehzKAzNUTlaaK
vbJezuWZ3kuFneBMVLvvS9yjdrKO1O8J9dEKodJnyhB/TjnN7sp0nzyjhiUXORd0
O3WZuS9spx8eRo9BFMjtYlIBDHkcYTEq49Y7tyDqo4ic8IqiP1Xj74Q2w5eYfz6t
fZ1NN0/O3mKFReDTxaoRq0skAM0G7dFfVGkLbLQ7pq4XTw4q2es5Koy+OOIBa3Hb
cLZGaa3lLN3xoaV/cXnmKh9WiDi04ojXRjSi4QSoBiG+l7fwJz1ZKK6IhrzW/1Jj
yUhOiraZooPu3pCxyKrDDru+WXgLR+6PEBK5PqsmG9SepO23+B9wLzjUEOFNUtAg
aMQS5pUrQDjm0XJodzMY+CwzU6hnbqaZGHSz+lb9Jig5dq5J0rRb7hGLTTyfRC4e
aRAHoBiYwxPryyK59haJ/UCfPV0vGx1irmjZ50MPtlCf6Y5HSpG/2EaXFDBxtvX7
f/cUR55ZrjLzaM9mH/tEllbdaphv8NxQjXoCFNV4esJa4/kAmLOiJHTqze+/uZnT
DuhV+zCbFbwLYiRhAZs2uTg0Ig1gRvaGobEmnxr8G70ivF5EU+d3746m0XeTs9ww
pPRky+2x64ti7byPg1UWug8+A5a/9YDeRD/NTNRyNdpsFnk2VkDDuOObkPmJHXqw
aunlOkyZdLA7Cc6TJDTIkRud5mO1HC/44F0wxmwFz8PdGwrCKmtfgnKT9S0hhC/t
oC+C5lhKbGbGaKXp3AwaWO1dAOVUwaz3CRArFivLZYDdYGPYEYX2cKP6W4DWFnZx
0uJ311ZjUHU5qsC1qldXUvZo7FGT4P11+f00jm2mSlMGik4sNUnUzQ6s8d/w2Y1u
+Z1o5ZB9jg+PiiGBCDyNql0T/rOSiED9Ez8t6ZpYknJTBTTcrSvyoS+OQJyf+TfK
oQIv7u7uuLpFHsCTJGxs4e128QhrsBQOcFqKiwrmPinojmuKrQAepLVMmWiaFLcQ
8T4GmUwEMWP6IebHi5/AlTcjDrkAlEqBSEvsM4t0vpP7VeufoqtNiN1tSJ3Gxa/o
k7S1lTX6vuOeibZoCLEMHlHmg2HFnDCqZgBetfeHRtyHuf4IqDH2Nm+bH4OdBFQc
6lSXk1don/n21/29B0cIsSipG1dji5q6MhYP3+x977NhmO3HWNAVvbigZSgPynDp
p6L3/FyXE6lI3vD71e8YkFnxQgMc+MwIiy8XPN+y/8RtEAQXah8/WFqMqjPejnPm
qAiw2V+FVd/DrRMfiBaDgL6vWfNaidgDSd3ukRlm6vMUYHlBbZo5mXmbYtYWwaen
Bxi+KcIptS8FZ3J8Kmp28MT3IOeiyuzi9up5V7a61xMSg/T5nUD6eHhxrsZkKAFy
QhYq3eeoMHdIIsWm47LsicXMzaH5OT0Ry+nQ9Sod6AiqyOf90k5iP/s7kCgE7QVN
DwkKpHPzEIx3yO/LLJSwDHKeh9TPZCY0I53voRJHFp0wdln8b3KCJEoP+36h5mE4
YKzxPAyb4dgQcWjKDRUGdzQ/ElgyyiwqEpGiVG3uOzSyJ2g7CTYfJFj1nybqvN99
Tws+cbCwIwqH1C21lpZvmQ==
`protect END_PROTECTED
