`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j88WhilPaVjRfWTMlYRNP/ctZLTqfXLmfR3J4bxZ0PmeRNAFP0ICoJ67WIC2XCrf
a3aHKIZJyhc0KdGdb7oluCGAZvNovf4na522CVquyr0A3lJ32jLbT3str/myV6JN
utko3Fxew9aaBFg/jlqo7hFFsc4B++6cE+bBMkzYvXWN6640KBu5L8z1nfruLjOz
MBWx5k8RvjTRbdSY6PhUTuv6OTaZlMjSrvxf/mNOp2b9vpBWxnzaw24yufPQU4LU
QwyXqd3kklWBbrnK3PBTkTPXqRjyU23jXtLT/GG7XLkjeiNuVZh8p28krFUIXv2F
dV0KGvSrqnvE+jgnA2Kc/PLxe/G8cCxR0p9ChdWH7doslgJ3guVG8YZ5dGuVZk/r
9zyvUrnjBjNDiVKgYSbo+PasnTsisvS8nBWOWqPmEFNI0CB3jkWrySI3XotMTdf2
soOX3KWJQd50bOdh8YYKMyYcJjC0PZoFOr3nALsErmwMELct0iCkIp4Qek2xz/tt
N8MUQNUtyRY7S2Ubq106AkVUMx9UrJq5B6p0EwNVXPwWehFZBTMabeJ1BTZsBRT2
a8ehp2Or6aD8+F587i5rMPnmFNPcvnwZXjb1rIkvlunWEkS8m8i77dwXsZnaZeiF
6feg3jqQl3ZDVw61yzijPBdZplds2qThFd4ACzcM1J3RX3QGgcT+49gGQs9AfI4d
+S8sLvItxKT163JPofIhbArSjRXcNRNs2FiGBExSg7iGaDOtXU8VEXKXFj2TQUU1
IZCO/IY7delgrUcN8+s6HaluqasAipBxasHQtDkPeo+y/MB7QnC97ZRlo32dnClg
gANo76KQxCrB90HdETfnaYpQHnRDxpuqf1Zylr+yc/7mPqxxDDA7fOqX2Tg7iDf2
gjvKyYQ1Ul1vXWR6PGUi0Eba3fpXyvT9l2CdpVPojI++dQLxJAV7kKfZo4axXiyo
YzoRWznt8RXWZ6pLjh25wzhD+KSHPecR/eTGWBLeaMqCR8a554m4vW4GWQncm6Fv
BiHz5n08+aEVKznkI9EVfusxfNSCevI4XmyMtBpCZ2ZspRVNs3GliS3SHibghoP2
/iiKs6MMt3c1QVSUKmPaojDpcVFTu8aQMTtDsyDulh0LPUYebMvHMHZhby0/DYW4
mmNjt5Gm0z0LsAqzsF0j+8ufHZ949PWyu3qCMpT18X/M9TA72WaeDHq+KE5wOdmX
o+ZoQpyAt+NNaDPtawNicAqxDcJiVWlLAm4JFKRjZY/80Lvhrf0Samcq6t7HsDDp
IjH8DHdMRsV+BFSeKgz1p9o/r6V1Gtv0m1TmGxsh0zLJCxjREFiXi/ic48vE0ptO
AS29K9LbGWyA9LpCHW2w/Qvnov/Xrra3uZOGN7ZB9gl6EMQCSS1oTAtXNfl+ySoW
GRwya3TtEC61cJkaeF0ybYaHd4W3I4RbH/5ke4DmcJs3t3bTSQ+JCq2w+++feyfC
lHEyBUODMrV3nNSfTujZFrX/T4QWxtBIkDTe42s5ApLrJVe2Wukk161PU2XdVTnU
9q+EJJ7eB/DdjnJR4segxsXK1rEVzqxQBeKd9PdoG5WpQa1hGl8bSNI+A91xbrJs
zQEATnN7P5lNdOICpljD2/gWYTFSfer+6Z+ciInx81I9AqPrRKpOM22hNFF+iuWI
RnoZAAgcw8r0HUj03nGQaR0hTQLa4eh6UB6IdKhP7KQ9PkL97/eywXaemQXHm0vc
rSZN0RtyGReEGhuhAR7luBmP42g+qIQ6zm/PgFBO+85JNT8y3u3HSu7mkvX21BDp
VEdbqhg4oTLVfIociIofCGt7Yphbw4TAbGYfBo7HP/nOUwAjdai3PGvDT62GkJos
YNwuFFf4/kV7EFIjwGGgbRfzHDomdgDde4tzoyp4WOXhNV+oEcW77jRkkBVvokrZ
p73Px5ghPBO5P2i3TqPJ2bdq8F72kJXq+KXxCdmDJy5KCRZbELVYNx8Z9wfRXcus
J9bcH3sm7+t1bdn8KJEdPRRh0i9v1WcorNHXkDmdMaSyTCmRFYaAkx8T1/49/i0B
UhjIxFS/S0/+TnLnIgMWopLzWLbBCocTQey9aHGxNZ1xSP5I9sOnPUqCFsq/djTM
OMXVDcYq3xc/fkgz7Ep39IB398yDq4ENgwHI4gVfDLRoL6BsuJF5EW8zZ1uip0si
KlqS2DO7JucXHA4102sA7WOuL7ThTPvev0PHF2XlfpyGcfBtPcoJlV6crxf2pRtH
FK1g8tHN14m6ozYEmVPWJyHgFgX0tnRJuX6Ck/bFZB9AioMGFYAm0NZjCXlRhy3V
53QjUqFgrBcugLYkDg6RqTCePpRIw8q7Wv/xBIFPEUSc5bXyrPJnbWO/jtnYoWJF
eKdBEmlZdME6mFFNgGoh72OplbYDY6iiFzapYp3h/l2Je37wA8P28LtOe5M/PS7t
RyEgp9DnVb8WZmvk67IUFWg5Lcy/4D2mGH1TVE7gV1Fqg6xrALUuJiRVD6FFj50G
+diq6ZAyLTOepMOONhuUzbfH7pAcZqoDleCbIF32RFh5aDUKcNFev36uCgaHQirz
3GItIAartefmbTxQluOMRlX9xLdtduuTG5s1pffnj/18JNmFR76CQEuHipYaP4Je
7Leygj+fL8bm2CimQjIE7MqyHV+Mk0dF8OGGe9GIp7iAoIy4xbZPlOeH8o2XCNyh
rkEvRUFBYYs0qqCCt055Kr4z3c3bbC4zWa/twnFBxPSgUomApUyCmYpCIO47vwh8
uC6e8lxU0Jtr/m1cs4/MMBV+bUTyEoMRq8X1zf6hWf3t7JQmMzKoEXxpmFGN1Dc5
OeJwKt4tCuSes51YiHRjF7V+HX+3qZOR8bU5ndr/tDbSz7xO5wIzojhKUgUGXAna
/8ma2S/fXcdbc7KE/Y8XazZTGMHdnNo7EEFJpTqzmXSJ9DLJ+AtDotYE2/jbfFOt
5ePspV+DG0uZpZDb1K6Pub948xvI3fBPOuxTbeXCZUg7PCXDpzQKMvY421aBmaRh
TdIOkaOZGM4X91Dn4QIq9/DoSj2IFLiFTKbzZKNEOZk1PE4W+tmoLZ7KaDia6abc
pr99uFafoQznECSYFJ8kmLN+wz4FagJzZtx4jzdNMzNE0DLzQxmrPhi3nkzjNCZq
Kt7gagUF2T7VS3DOPK9mXXcApK+6CI3F8JF6zOn47pRewNVKuI/CtVsxrF/W30A5
gOoGJr6nDrnS8DBy4Xr13iLEDvfFoZJmMVYp1e3hrPvqnZWfxanmjgLAUT7o0oQc
3u3NTeN1/sSiLwdbZ2IH2DBrbZHS4UeuU2KzKikb7RCuBKF4ueG8l/JN8d4CuQN0
vcoj7RQnxunP83Xp5hyWC6GP+b6QONrdSopMR2fmwPm+QcPh5Xbu85PTbEI/qzIb
fnnYL0LaXNMhrDbqsYnrNbY5fJkaz6+Hqy50Kt/NRQEwCSg3CMOXppUnYhiBcdtz
kXqvWId8l8t3uurAMU9FKeBpLDp1dEYNG7RRQ/3+kysKo9Lipm4VlsrO83+T3IzI
05ibpGnF68O49AvFAzUaIpwkBa0C93hZI2T/aWbrZg9ZKXHi0ptgTzEtAjx5CpkJ
EvYdwsZRi6h6uuWeYzD3FrGbBTN5CbRTvHV+OCP7ZBFFY2UNDTdEZneMBQoB3OIw
FkjTUInk+RKVf0fJGEK8sFippM80YnEXOo7WxzWUSf/Dacem9QAE9PkClRnugMOk
aSzdFmaRRJ/le5tuthRW+rKk41uQpevvHnPdP6kCavLmMm/oehHjCZDqvk+TT61L
6TQmXBZWjn5lQBtq1pk4lZxRvTZADGlHFmbIa4mdb8993mT69pYKxuNaKvjBKpGG
dRECxne58WXysTAdW+MGf0hl0ubNIdinExZewvnG/sV8YnngkcZkpZzrz3CdM2ZL
MtF92SARSs+LADvJzsVeDGnvP7wJwDqkqK0jklClw0LZcgZXPEkVgLPqk2usSKPT
nTgn2qB6sZqm2MYeX+48xonrjQq26IKiSxvv0uV8Wn7fOWcVBkofVEpo5UAEPGDX
reoMTfgRcl//hkgU1OogM81anlouTbHvyHCNb4lNYU/1FMWg7fB3TlGqn7ZdL2+z
xPekf0yrt8nrKXsPwMPIjwWI74yPC490oteeoQmNNO/3e0nukvAdVPRQxfjvh/+o
YRBQBGIhikqYx6Vz0xMeVWo/KBU4LzXyITODfj5YdUZ3RD8xo0RXyV8rNM/uUJZP
7WDLXHuiqVvBxZwY/JQeXzKEdoAaKIwzp99FMCPgbj0T/Pn9q65pM/5m3vdo2OrM
4EHvZsWO/TNw86DsLmzGXuaIW3nT56fXhYJ6AVhswSKFPJ7W7TSH8xiRcpGFFK5L
I0ituxrQHQ07ff/YMN12B124a7Kbx+nmq0l1bP0RRJ5Zi/5cO1T3XbVv/CKllc5T
+OeF/wzPcOsKNIIvOOD9MRg0zZ0NDzw9C03JNQzwYjJvkzcly7LtyIlPCgHVJFMl
uLW+utlMy4oKeEd77QkJNV4Djqn8qxZkHgwrssie9srA5oSgoJjzqCoNZ5QJi37h
W00iuA6cksH2nJESKBuKHpxLnJS/6oEeFjh9nhezgLr7ON50uhMyfS/ibl0aVKIg
8If94cmp2gkFm4jlhY45cAcRUaL7MiVNNm9cY1IPAUjmUvt5fQJI5acLO/k91y2y
on89xaqCB+Hjym+ip63dYssM5EDZQ40VJ+GLrKNkIvFw5Hq4Xon9K1JfI81gfjTV
GLTrFVAADUjtkotuzNLMU6if7aENgTJwSBSQbJ2xtfBMaT/gjQWu5aZvUge/cmuG
bTaWHeBcPPIeqEDi49jZsH6zj6Lw+eEBSnimZeVOpaS5u0LyVzAufhbjNi4WTOEz
MZH2Cm26PgWUYJ5F+8HARZkkYBco0gWA+/aMcG4i5wl6q5heCyQLfFSSc9bbuKLk
j94kLZG2aPIT8vpeRK1y/AiEjw/HIrdF77q4TxmKSdGrfz6gD1yPtjaBsud7HuFC
mOwkDOJg1mHrHOsqsvfhfRDwuEUKUu5O571/tiGhSqXlcDgfUH5zxlysX+GF/qS0
SQjJkEnbhCPNOaTBUhUGFPoXsEUpuwO+sGoy/XKsN8aqHpMdPvmvuC6aW0zB+CB7
M5XvCwv+MFj9nLS0OlIlVXcgLp83vEGyYBxbr5YY3pE7KHh9Tel5HAwUI6VU5iPS
XjdqqGeGiRCAD3yAXwYjDRgBlaJ6oAbvvsjyd9nP9KYpUsvQAbSTfs20yshMAGMR
rUn3TnnAs2EGhAY1kNyeuiwrLc9Lfnl9P0SX7bsLNqpwUGkxmk5+VfI1GS7PZLI7
HoDpBzdYEoPpk0hjOwJvVRE+za8xD3zFeU+PnB9qU1MRjAmQv9569O01LzDBjjZc
1qWW0sVLaaNpO0DRf5PituNBdz6/q0Bq0AZeMzGRLLvhCydmZ+MjiATeIZdX6Z7F
144loxcMD31KAtRzvruM/EeRpsnRP17g1tBJbk/DjhnAlMa/PGLk1R85NNo2nWNh
UlGkwntbZGJsQpUbpmIkrmQeGoz5lSSxQ4jssUAsBCJaV/N+SW6AIdSdMIyfedey
vntOaxk3rhbrnVr9Qzzb0UHsjgLsDiiqnaDHE5UsiwpXHmqOQj/EoHN8xkE2l5zY
KAlbG/Ro7Gn+LmGeGX/P15A2DWYo4ZEPhLfMhmLMd/DTDpv2U5m56C8hDiFcMkYM
XjgKMkjcGECMVdABmXXGYC3EweNoiOIQWFqGPRu64ybTl1GTKh8enRTeWDOSE4Q5
jskfXKvJ0mvnSV2bpKzY3VhVULxDipBVjalS3JD+48aPsoA67y9LgHSJ+YcZUJE1
eCVLzNZPXIQwt+6MuHsgHvawSP9XF1p4GmHs6DUmEdJD+Z5IxPBs92Ol2+Jj42M8
jG3YE6UuABg+q1HIYjbiBto7bL1a0sa0vw2m3/BUtrD/JWW52RepmlMtGboxLbMx
9WNLkrLSMbr2OQk4cyh2pefzti9OE1jITL/KXgdL2A7C2m9/ldRDvOE+XhXANFhH
IgXE3yI+Vhstqanj8apyZrHYn3PWe6BIAsuLXMUAC/qYMJWHXrCBxn8Ra6ggaZRn
6Cfh/eQEp87h8j1i0yt14JsFyHQjn+OhoLbOTJ5zcqcg/JE/aQXNo9NxP5mByc/C
0FJz+RfM8CIwLbhvmbSjdwyI/iGbGKmwp6nL/GPKGCvO4mTz20pQvv/49QOY1P+F
zapKbNLH/gfj4HTuTltF2JgeFXvi8kPyTEWfwfMWKvkJ5I3Wq0abxEBbaZvn7fwy
RCvWCSRFkqinxNtWtFHysGBlLLkqFDGIhN/XGyTQvAUy9W+FZfGz3maPeRMbWMaU
WQ1POzNw1o/99/J2X0o4BmHtlHYZvdO6XKof6nHa/CsV9Atvd9DXcxiz4O1deRw/
tjBwYuZLj53hkxVumxqvwH30lYkLUzHYGlCCKehIEnS592rHllVl6JcI6DXHIAJB
FDlUASuRYiXv6xBgQ7Nk3s7cFg57Pgy12iZMw1aGUoTbd9UM988oQfoZd8WPX4op
aSg4aSqaWVW7/1K3pKvhdUzumwywnBGxNO/5fu3ZQcnLI2+ckjiM5P0RWrAaso73
f5XQJA9O/+5HUpALrAf3vZ7qItieoLid9sxnxpC0zi8m0q3K0cjpRgQw2wdovJzA
RwCmf5irDSOm5mva/533okzrxrfn25CXJh141fvBgUrz+hWWnwhRkGXSXP4hrnYs
25mgtCC6Mi7fai87+GDetz1vwHfJNpHULOX0PRZZ1OEsMr0K92xwvekRyOLCr9Zu
NtbPYIQ95HfkjJI1b8DOij4ZORtA8jYSUZ0htrVYmFHhvPlu455p76hCnAxeGSzK
FMnwdJRnvVQj2Nbm5zTp6rsY4iiafCjaXJ3XYc7aO6DjBStWP+uZ/kLE3Qg6tqp3
Dusevtrl2qqcg9OcL8fw+7ZyAYZeg3dA+7Lk8PpV0YU1rYs79eK643T8x3sEu7fH
1IK7d+jt9saDTwpJw82zqmK7G7o5S7HIXRkBwCSm2tErFXQ2teadQYwmDrWIK1C5
Px3GuqlzRNsz8j0kNGP2nxrX1YVUCodgVVU9C4ExRq5xjwNLmILCRGM3GgVUdmw9
BVqHwykcDrhBFuP6Ks0jtaY/DrIJVG2CJj/bLnAc8vHv75Te15sqWrUxjFlRYMQ3
Dwij9GR3kuOrUkksjEMbMb15oU0P9zYNz3dnkaaVMo1Wmyw6GDToUdXPL6cxbTL0
pOhW2VzppThyujLRMpOUQdQXr0mYjrLpNEXXzcc2VMcMlb1Rl7lWgGj0pHYEEybm
EHip8pmXjWHikCdXgtl+Cp9aAPa7JxoywBAxeO9oWLMObkVb+P32V9s8IYSQ/IT5
oDPV641e5qavNOmXywbvhF4KO2VP++D9WnW4QraUM4SIdXvdH89gBCqy5iKOJmWz
enQ45cExgbmIW8XnIBaetQMjYFl6OUsH8OS52PM5IveJepY2c5AoCFKmELTtdMeq
bMstLHuQvpKt9Rs//JpfvZQPdRCQa8/2hZwhZXU/FowIXgR/AjaO2abmFrb8E7VB
f4lKZRi4GjUEEXjRoYMGEm6jVgqQVznlTavfN2NjWKyKwoslp6nytef6yx0aRev7
PubQHZEkyHi++1oekZRZGS3FDI6I48yahcUEJACzXsgv7iIeaWBc5qqfZYA+X8nm
cL5Hh6jbBQv32XuM76CAcGsaHoeafXE6L7yORl09xiH6iUkvNYc9a2Bitf0G2Iqe
BZNbRT7G+oEpTuXTGaKdBAEtxPojl8nQcuKECh2hMQgGTEunTMEYJ/neC840Belc
TX7f6mgUeC0pc3VgMOLgaONylnSi9eCkeh6t10Xy/73Y0NHGO7tXpsGDgkmKJsGK
Bug4km4qmpn9+g2wQWG+Q5MQ5E+dGolcQ5rS3Yhf6lZamulpy+K6C9wgROU4UfOb
wgP3aft8JArA/uJVe6SSJvvTk9Kg92EJSdPUdHjKXHI4AnjG+Vk9r1C2jivl5s0R
Mlxx68MaHXOcNHNlfEv0mQ8L3MT62irx7CTF4M4z3hy/WqH53fXWX4z6B4slOy9h
bfexHLAq1F8oT+ynGYHvsq1VxtrvtTQRw2jW5ZrTatwYfFbEweKfb9v77aJAVQjM
53W4l2rFZmICw55tNylrh47YBZX9YLCAcNgrCSHBRvXNcBTd0UBJz3KHmyBS4pFI
EHD2iuw8NTmuJ/VnF/Ol/oWxPapOmNhKUaLfesm1HTRvURY45uhmnazI8sg6RK6o
92ubbjTqPNgXNuKUwdTjuJX3pawWugL2yEtHlOde9qCa3gBVKwm2tyMrAE8geWI8
VZimXXOPyTSwMqd4jiKsR27icpboJGDZe03CUXaYUYdRQDRtwD+JlUXHfuob6C7Q
Na/a7xIkCDsLwATUXrk9JcjAAFM/aYcI11A8t5rxSpldN+ObNUxLFlLpLv+ShCrO
9GwIvxCiWC1GHjZdP0qDboDXT4fRm4v3WYIJwbjYy8Ydwe7a6yYq/4GO2XxW5xmH
9IIBBRT7kx0747+SdEMnbJ3FBR03OZA9mg5uxX84/umJ0XJnn0JlRjhv1JmWfaLL
gWcVJaIoE7HgLHzN4YRAmiYGqENu8ym8gLJrs8fGe6ihWyE19uKF6l2AEvPZfQUn
kVhuEnCTNZ3ZMAtwbmQOGPt/WmJSyFDSl5VymRhoTEOu3c5IpxOCxi9+FXN8vX9b
AR1IAkA/fsfBn4l0aP8BHIq15oz9FlHF9v/p8hZci7UjG9pU7PHP/8r8kvXs4Tb8
kGwIeQutHJUcj8SuxPawAs9yzSaTRAi468ltqsuV96dJs4Tp0fs607TsdjGnXeqG
D2W/Iq4PXdvknoe0F5aWKDEAmTlT0Q8a1qbkUMdxfVasrWCYxleXXrdjkJFl3FzX
jFDksdUBiRVg566Yr3N1A091PEkpc8urABUdBl0SxxfuNoRr3Ebskin0gnk8i3N6
G6/cMUUCJGW8oGtij+wGXOtWwpb4xDUISPXP8dIWo6jbtBQJ/+K6dzLeqermGkaa
yrvgBFeRM0EGt3/dozZPhf9EFCRV85h6qYAQBmLcyPGRPBOxomHb6TCYbN9zipxp
G6fq6VpDtkaDBiPPeUUCrdBn9McGUTKASEkInt2dL4g0LhCQgOCAhRIsDyv7woZG
435C6t+JAeEbvYnyhldqWUNMmnjIqDFHNAaNxKXBVzjG5h3tuIkG2ztxxEFB5YhD
qMCQUR0eQEFC4P1URnRpQqMKglwx+O12td+dwIOJ+2frGXVUzPGmlb7rRt132xBO
OvieU0leGMzDWPwCRdf1iJijqkp9KHFenqRTxltTWWSbk/idDlIFYaM4XL8DWk/r
itOsm1oFI+eGz4wKAsw23lipBlwbuexmOkCrPZaGg+L13LL9RSYJkmwr7bQmAKtv
CNNU10ZHDt/4jcPizPFoU+CjDM6HkCFqMBHUMzCuhsnLdhe8xW4N2CmsGEot/vpR
w42vYhg8X0j0YUqRvmF2NrpTs2CdRgfDa5XQrJRSmtTjbWolXPXI4Gq8+vTFc56b
KbU8BOJloZtHhUHmRFPP+hs+mxVG9ZGvyJ6MRvLY0M7c/n1I4btsqRPSuTadV7zS
iZAppP7iGWFuJc1A807o8PbAFsJRDycF7EP5SobOBPALWBbIR200u2FoRgwxpwbw
OMUc19nchmHo8PsH71DzVrwolQ1hq75vDZYp98t2ycb5AwdlX0zv9/2Rz05FrDIW
ztMq3vP+u2wQ4br5SkRLIuM73FF+eXWOZk6ZPXoEBtX4eWWPn9lxfQWGq4KPIt2m
crDrxTwoB7n4BmaMt8tn7NBIDt1+u8lvL7h3SSPFbYok8E247ZYF3vENd8SLOwwJ
WUdHHGUsOKXKCA/8vKDF8tzndWApey2oAwOOogzvyxBbcHtcjKKnSjDW9hUgAkAw
Bt1HYrl/7EgQ/9zGycaUy9SU29VoqnfU6Fr25Sza7MW2ZNE/9/KVK5GBE8fsqtrH
n0MLdBEaZuqpU0McTdl94L23F0Ui4DePIsQhQ4/dvz6WtLjgQRaFZMldmFIoTR3J
1Ce4f5ajrbYyRTURU0iOWFgvF5hvbpAEWl1JsD+NhVbHIv/PkwGJMDzs2loAJruy
1qZtXGrBpWHgewKXCFJBvi+gBhjNvCoCZnIc1/OOUXgiqfCFxhFEske7EJA+5Q6c
4p8z/gZojERm5BcLKvBPKCInMLGCtqWPtwtptFnC6dcuuPVIPaqYwmOnjpYja22j
7wfTIagKoPPcI3QT8DamCJFnM0eIDOwHwjAfa8ZPEtgfvTKbsB5g5Xfex7th0nlo
LgGRFkifbwShylRK0+zCfH6QXTuIt5XylbH/LOxct9IthO3QonGv6aUHLaxNKu1/
G65Zl+wRALnHMx6FoCjutaQFjlT4UpzIaeoyVAtFww/JFRHhbIiQglM5CZ7PMCs0
+xpdaVNrUPMPuuuFWew8mPYUEa5ptErqVD4uBFPnq3OR/sxELh8yr+l6roLbqYiC
ewSw92Kdg9SCoTrqDyqF7a2k6KyxOtXbXnFxnYNqzfLRDVGju0Pq9y/wrCIAADtA
PqJatpt6caRSSkVM/qxQR2oiBOCMojDG3gtZd8X0hfcIGDdHd2/zwBpoqDEvQzN6
AcO6L8qLE/PBr+mtdTcWcVOuaTLlUOXeDqeIRHNm27FdLCSt4+OjD1Lp9Kaf3uuD
DzBZqnfozqfSzQfCBigDrnh5n3sOx1s6jUf5OnyNf8EHENjXQz6rmikYT3svWstg
G8BiC8Cv6abXtMXisIy7GnuJrG0e6yfzTK4Ul8tz9Bzk/pHwv02e7Jz7embOPdjY
UlIosHeywv3Tcvi8al6u4Ddr8sxN2HqC+6OA8UCeNbdjLFc8RKqwq95agSH7jjjg
hdUfqblBhNNhVLGNUQ/QV1lnFfGY1AfJFQgBkK9eVTvrglCBpuejH1JWBAACt8Vo
mjd6DbndXdb0Yt9sHo8ABlK+AscVe7PRNa1W9kVE2dGcTdLzxXxBnDEYZSBbTHaL
EF4P8pWU4IQ0GNW/0ytSwslpnDs5wtn8AKpMrEH9qCFToYlc/8wgXpJDXSkwX02a
vCJY6VN/cgJA/yl/yOie7bQnEvEVzKaCMNUEI+0dSuGc4sNo/HWScjzEDyO3PxTR
RhStyt3H4m1MaAnH9Tm5enQH2N/oofd443V40VRM9k2VKnfM2LoQy3q6VFifAhI/
aDYj4hCKjX9nwaAyxAzsk7Aq7HPdiJGDUwl7f0Djo5PFXaSi0XlfjO99HQXVayys
qaxc+BvhmCSXrLGASkHlJcYwdFI2n/uyNytGperfphgO/YGPjX3rGbGIiFjvK8Gh
Knen1vrqTZlu3ZVyNVw5SDD/OV1ggonaK4Yd3UU+8uhCUuSvqPbGG1zeoeOzoE1U
0CS2xjlCjKkrFOidNNV9QxfpZCGGMKfwD9H2Fj0lJ/3WE5ZrlB/zh575AxN0tM0b
EkPLOJ1C/QekEvE0U7nFwEWqSo/c/QD0D0y14HCrMv9+Yup7tyo21N5ybpyX7RKw
r+zp7ivPpD6oYGLWSKlKuh8Lor3Ug3kgSpNCmC9cTCbMVlF4gXA5fXbkprEESw/9
ajdbIBNw7RYNTKp7tnS7qHJ8IQXd0kKp5/dh1uarqYGsdKIfJKQLFIPl9+Tgkewx
CCKs44UTp+cYfiKFli2v5C2thRi1h2LhxhpbD2lKEdMoHeHBQWAb74ssLdzNcnBk
dTGy72AaK+bPay73mPGqwn6VP+LieAhJQrVfjdx1ktPd+mt3puq1lEY/KOPy3afL
3shjvwkj8QlxkS6kTiYB0qi5d/10aByLbvLcfez0BNpiH2fJqs+kGA/zx2E/sdAc
H/a4ed55YrdByBXcICsjxuFObbbx1bYOFQ5kUzczTrRhvQM2QDjLa8Qzd6URUJMf
T8UE2+8PIqySFqlenhLKr37KJpw2BFT3wAd6gSBWbLIge3WY9EUZAkSbjIviP28p
qAFyWZHF7Ok/pWaM7BIKwoe7KU6TOeamRiq2OHHLVIBzKeZ1KMlZX789iz3UsL4k
aqG8dpxWgt1mDMUPG4jVlAfiObxEkP7dubMK59ml1dj0raUZFARQHS2rYbK1lOA2
CJJShzfmNXdOdXYP3/aUSumpg7iXsr3RZwh2HxQpVyMJLwBOzeXXHHScEOkyr2sH
zjF1S9A1CfOO7j1VrSYOVdisl33L8YORFpCXGKQaPea0q+CkATdSwAHMTg4brWCe
jDkwjXUPKNsN0SzDNDxynrp3+HA6ULoXliG/SasXZb0k1+i6ZRbAn8+WY4V/DHAq
dlp72LsdXyKERglo1sHB4vmv4llHgSBMdzUtMCVXdfIysSJGFSFDaN5F0fOZYWWT
UDmNL6J1QtyLvJzCwP2SS2nS3nYwMX0gaeCQrZzD8mXwMprhkljDI/K1FGEQL8ev
nADN4vDBzpP1nZlbZ4dDxdgWmvN2mmhJfu24MuvlYIBpx4nBEUAET5WVELZGzJoS
U+YKf84FtNBK50MyRkoseZ+QrhkUppTANIH9k6mqb3RVPpJ8ijHmK7VWEJM20NQg
SpM4yu/2QUEIFFPzKOTAnNOMo2481n6BM5OS6R908tp8d7lxxYG+CMD7qLx6WPC0
DssesyO0PVhR6lwdUBqTcdBwq9JS1m+buLVjRJm6gvkz6cisUYfuBJwan8bOuD7j
1xnyODNmGIu3dYKOnZAZ97iV19kFl6DDqeKBqyN/Bf3rT6/tf9LLMVZXIHgW1eWs
tV35cj/OtnNfPjDgBKuKJDM4v2qWG8YobIAYEdMX2sk5hjYuvNB8Cs08eBojHSyF
25XP5XvCMWv+n7oiZWK9Lpykhpo4/tOrRPz2EbyR1IVQaj30VGJBKoaeMqa9H0TH
BD22X862Q9gb7tgvw2GSVI6foomoTfWQXbiTKa6Ds5AMljnAanXHpPoP9nq31Fab
KAAuZ65g3V2Kn2RyubyPIPjwVcELNEFbWHrDSP7Ne89CNYUUF8WbVbyO/FFj9sz+
fQC9XrnnFaXQkxQUC+6XYdpl/VpLMb1xDBbNlZFtRah+B8r7ATzujDMOvwLxtNVs
AVTs40mMrGn0imqwlOZh81QP1AtrDugktgFzWb/hCnwLzwGtOI+XCwrcNoY8+Gqf
ekrHuhus5+ZeDRNYrdUvjDDWob3SEf9LHKD014qVoQgnS25f7gQMA0PU2SRKrRWb
rGmFCmH2CZxiYLiZIuRJb5dAouAGMduDJXqyjxHD3VilVmTpdhwsF1vmkrEceLWX
UfJY+ty0RuX0bJSHBSuDU5m1IrvF+ik1dvtzNiYjMMvlmQgm80UKUCoaVGo0Cxy5
Gsb2sGfY4XFo7c7A8ACcYJctGqdJ2OWiVK37h/M0EIfzB48pktygdhMVCk+ZJ2+m
2B8LGXK8MF+NV1+A1jq9az+8a0PFT/4uS/gENOk6CqL7QtFBFLcZU6X7JrTcJgXA
BCPfnWMCkKUxP0Gd7kzsJctjLXImJFznjrg2VS13WUooDphQJoIcumyjKdygHnVN
3dQFpUv/B8yuDj//GfWxZc2sMikYKwGUt0t6jE5+kbI8ylOmsq94jKqp+Dww/umv
eRdnshlksGPS6PtgZvMoPMKkiJkIzlhL/XBbEj36TOxs7Wt7CnlwNSySlsuRcEgi
an/MYDLsnMkQe2j4T4c1IU28cq+8bnoxiV8RaK0c/AuCAzdECwhxf7H5jXiiaVV8
O6zWFZABc8xsTnCGuHoN77e07M1EY2GLYRujw924+GbQKAEVAo3DPYz8x5wqYbnk
tYexiUToHCSlSMiYF5d6qq4/wVmqK16Fv2logJkZuy3sjqPcFul16K/3rZxtJXPL
SM665Mxr3plkXJE6ziCsTbTdwmoudW4/PEuNMeghOYFHYE+LG38GEa5iLvP73zPU
wddTUwQP2N3/SAfpl68aiPj6WM+jo8Ppkkk8OP4lGrhM1jSX+U/aunVoTLwS3z98
z5UDKdHMSrPz9t4L2xSFmBZTAMXfw+FyfO3Gj5+YuKGplp5km3aP5Rlv3dUnTKnP
PuL4CN6EoJWB04p/m3WroNhSCYh9WY26txbV5iB9XBzjZI0khgM8sod7uyNp+tqt
glcaX3jpXmNbI5HAsvL0spDzZS5nlRSZfAeVT8H3bkow+Mj9b3rOB6JxEkYusU3d
SjVffdwBuuYMCk02iJWUUK5gBW3t9itM4jI23+lEiuBYzH3bPq5uozK/QbMgNast
UW0cwmTvNYXGUIgN9DWxXjK2JGgVp3NZUGLdem5b8nCqxoDKH2nXrLws24wU8q0s
Xq0BhcGCfn1AAX28DA0RjU/AHK3RUN2XK0jhfZPfsxKBiOL0gCGWeuXKeovnEwqw
hvrTyyp84YKfdCRPTYkNst/nvj1Dv6akcAPIUfTGtgorYd+RBQ0SR+2HbOI+YG22
UtxQQuC/RsaYzbMVnNigIPL/5+iBPvw1+deVZEjkMrZJF4XIsvt7pvb4dJbwyWK8
1BtsX+Jkch57zI4QTv4yLDVJtjbf+Y/8tWLZDcmVf0XUny5J0Chel1NiNY5s3j3x
RxhbPy0kjf7HJ549GmoBFA8GTujLN0zy2beCP+542nKkTrs5KjYp3WVbpqrf5RDw
pX5nTlU/nW7fgXnoKTBitCz910n6dfYkfvhVaVxni7OAPiI6uz10h+RQPDIlr2EK
j3z3WiJxLs4tJ/079HxtncmAMz0Pg1IreIdx35JRqBc+zbNQkGqxoxOmojXaKdHK
LmLQQLjps7SJExOE7m0O/QidRjbzJywVud4n4p0HcnoYGfiY2AjTWv/l+IbCbXF7
dYX/5vBtsBcEkKw8mkLOo6viJMpf75nAaZQ3se876B5lOK8cSlmHlYPurCbFuEzg
CRxOiYg1xn4rtvNAiBR1qDd0qZNdqnSh+5GqrGll+WCkXc5N3PMfSiFO51y+u9KK
dR0RKQWzhgJhAe+ayyXPnRu7AwbrLLA5WcjWGsLKLRgtokxzPldbYFXz5yIykYN0
OJPl+8KLc3vhks2MksmItP2uk3UnOkIq+XOCb0pMBRaLykROrIbAzg4xn6KvSuoX
Nu4jQsb5twUxkWPiqqwodvh9LbFxlMzkMyrLNrA7HzpzDeHQ2/8JldNyXp2YO3B8
hKNvSQtJlYIXCnvgMI42a7kF8lylwNLPU2eysyMEcVmXQCp4gyUsnvnr2cfqHmH3
F8mTyq9son5mq5EhGe+9fd1EydT7V1HtQWJ9xhDdPR79cqOatv+Hn/Q4mBcdcj+q
8ouQjfqPZXl7Snbilkw/O+yeRgESzkOJtYyO3YLTa57mF2x2uugTAtNZWzTZj5iJ
lr05MLSp4lcveyoebKPvYt3LXEveQ1TDDXeHKAIoz+6BM4AO6YHdqj6vXJpr2Y0w
TtgQiQCCDqzg6ZLXHsdH/bQq0Js/OdmGZzihYQQ/QUWyIuuyKJdqjd9SPBylU7ws
wTGv+bF4ofPAqroRjwDs7bUu9pIFgeOtHEgLuiCwdeKMZbj30+wZBQ5+a0rQDkNY
ZTMEroHXMS8h9TuFARk6RdWjB/mHZn5dw7filKyD7e5ZZ8gck1tSSJGIwAtEqm6L
ognUpskD0DS6iE7+oZPsSl+ZM8j6WWvyNNSJbL5MBXtq2JvB9Vl7WZwcHq6mVgiv
muAO609F0UqnK9cmAS9CREr9hlUeiF5S81Sv3hw96g2et6uBnWgiE7HKuzUQfG1P
qmAAKqAdxsSFgsmr3kTsKPuNOyrdXWUORw47e4rKuL0=
`protect END_PROTECTED
