`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZ3C5BcF+4l+yVLQk/Wg2f/Zuf8c3L49IU9dJ1EEUY360dMAI5ltUTgp+OHMYgSN
4tKj4Cielshkx6QfFVEbXJb1q1uFjLcYh4SjstsUue9s8qCRubOwHGkqH254ziwD
u+kUEe1SP42ZO713dzZ514KwNvc0/N+HW2Fbe2nn/vbQkQqHl0W0GDKQkdMLpj/J
KWfeJv5gvb2Wv3LY4y/Y6FWCqAp2mZdtugXH6hLIKL3cVEzpLTQChxaIA5ZbnfGV
w7WUl+xDohD3Goiv3dBtJCYxiq4VDBd05UvNdWoQgiNF0nxEJbj8gNtj7fUavs60
RBMfbI1laOPTTTuHKet2Y4UURgq/WodEwHVxpYjkkMxcensaYDA90tshR8Nj3Jje
/jySHZwIS6Nptj+Jy3FekRZK0oMbFEXvJvbbSW4QaNqgfhZZKtdeZGim/ut5QjaF
dTTeNW8otTpriYC43vzUuqT0KYTFhbRqsfdRHMYl9prCr8LibAq0QazdQJjNaZKB
neVnwMyV+WfW+ubTWGUMg1vk3b1hOSsMDtVNNVfMK/L+CrJttZWfyFoVTKsxG1MV
OZ9HLkArdd4uMvXxgQVlifzI5JiLqFoJDW/WPF2+14pMqLBWDt/+Yi57ZHzfLLoT
yiVgXJWa6HnJ/o530rP3Ga2SElO1VmXvupJG7rCNbnVNr54NOtAFWwfnRzeS7xZs
yM9DxakWGKU/KCklV1tlYjKAGw0kNYhXqJoAhpuxRaDBJz14QYoU97+GyUIo0Jtf
kxh89F60sYWk2FNjbgCoKyWZnL42DWbcsCmP4YbCDUC7yCrsyw5o3/KLkfgjDA/x
8nC7ArLcwhzEuxRN2poAT+dSg5ZcyGS6ChJzKBY10IC4j/2mdAq67PA+5HhzBU5u
AO1/wi2ffmg4M6zw0urupQ==
`protect END_PROTECTED
