`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8K8na+ACLSbT59z99NHnFGMH4NJM1eY8Jrulpb+w+2D6tVHaxd7ghFUtfVpAu7Bk
CL4Tvqb0NUatpT2NNDTLUo4n3ARGSNS7UN0pR4imDDbW/GEyYm7tHXT056ZPrBlZ
24KVmxNaWCTuoMxvXp8XDVKwN8GZX3A6gbRcuss8vTP9oBqWd+xDKb8f0qsRnCIp
qleutavnnwXq7lY9AL4JeazZ+su1ZyaHYqi33c+j4gnZmnGze1CTsdO8C0GtBlet
KHv6kFq8QnGThVWDGrx/GdsQZkaxeENxsoWTulI3fNmExUkaSbfQ2V6tJvR5vtbZ
XTVWGsA9x0khY+vvvQdWsMVje5mSB4N7+wBMgr+Om/ya6biF4knlE/ZgBR0e67iP
j8pFVBighBYVer2dhAjw9F2Yj8GDguuZilnQLYVFo9s8rIbwCx2R1BnMsZI1Dcvu
f4ZT91MBmk5sRzRjsdOnA4VdBjK0/J5leGTXuSBCz4UtNvPuOUvZrRXWM284JIub
wCffw0vnaK3wRgxLJWEsJKqY8cIHIWyCYhjwkHzNk5QcLt7JaZtxy2+NdxtTDz1W
sU8Y7KaQohkWmSIZ7bfC6VQvCsVUemZeobEAUDuaEo5Bjo5cP2rs0/2fkUeE86N2
/B02h9TtNGFCxLQtykk3p1d09gwR1oRxr/N3G/gjVpc7OE/TybXfHuMSkWdypcgF
d/SjPSkqlY53erSDwL2pWVQP7cnZzFBNvmIBHEJduD4V2aH+Ig/5BzqSuBEBzq1H
hL3sLoc9lOX5tLTXwQxB2A4Ne/2r1rC2DuR+jEXE/Y74sJcQHJxYYnOqqzWmgz5m
`protect END_PROTECTED
