`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S2T6Ge8/ve9Ld3EXkdUlY8Zkc4qvYiQV66rVNfgM3L3eTkqhI3WH/BsWt1RrcrQ6
pgwV7nqsvKVRJNNr2Q/2mdFWjrzSUHlkwEjzlumI4fUJylrXhKARsqZ8iR350+Ue
ccXTorebQAgxJEIFWuDbT6eqgS6D0KLPs2x2azoevkNrceuTAPGcfNegtwR486jX
LRDZYuTICOz14lIbZBxFeKARY8onsR4l7LYu+0/b3qcMAjy9JYlkOnTcfu/BKGiB
/zwcJrCGamquY8zlqr0Lo+hB9YD9wmAFHVMhZnUTU0lVA26OlGf0iBX+6K9tVnaN
/oKEDO723umo+drPEwYQe9ALl5TmDTePemB/xE9Leu9zcXwn/AMl+0XX01Q/mmkf
zmxbCFb4e+TvTdSUIa120KiEn3XkHDj6QDnPlPXmGcC4PJsty+7AsqRB5iYXRXcH
kX2xgv2NnMuBXJJlGExiEzvI1CeiefwO/sUnfSwF7oTj26iPbllFplmUKyo+9rUq
T32o8aoGRKwdyTpkB2M4fuOUyk/T8XaRyZWczMi7dLPXC969kmGQ/fhpcQlD0OEI
Wal7YLydjtD+BsntrUib0q5+L+3wWo+sEBMEn8y4dt8AaVC2/Lbp/kd+SnV0Ws6E
JJqxvKq8x3rfmUUudy33NxrWwvRbp4TGINavPtCZ4/XRQIJOORpUMtadxzKWDTnK
wOjB77QJzNJWvAmtVRNlLP9WFh/1Lb0hgZ97lCvtis5/41Dj3HAbflm7z+xQe42X
mBeNdiyBy6T8cw6mSZVKJPs+DoN4VOCLYYXIWckGFSFU/VKoD+ZESJGBWQ6n2rpj
2VJQgUFeKgliGP1oHQwOfag88S5QdaqOg2wrIW7qzA+Ez8+BFO5gyXrHsFzUZXaE
QZLY13YK1JG/QcbWEQgREgk386zLp0qezY/q/mlgZnzJxDH1Ez00V49gqggZ2aYm
nqZyeP69LBIe57Tw/0vVymbBcN58MqeMl8++8ggE321Hc234UGjuF4bferDPbwVH
kDeEL2F0kV/uasmX9gEaVkSYIuariNS5HcQq0EBJMa0XrLPRamBgX6/aA2gIMIeL
aGOw9xdcTLRKM59acNloLN/nLtmLpkRtWrdtQgqTProDL3C12GK92XdBFE1bU/bB
Bz5it5WCH/G2u0OB+uYpz5cOQmL2l4zBrd/0/eodIr18oMyuip1KKG6wzkTmDVrd
q28Ox8SPGX4uLN3VasJ9VzSiag+9QoLGGOGwWDxwvIdpDH3PJWinvVUTkpl7E8b2
xsrpzo9+3keAht2Or0TdmV1B5vjdt4eWTwgse9N2qVSpFUVfqSllAyXSn1kK/qJF
81LXRkCn1u18BcBhxOe5kyHhF/HCNe0uIh78vTOhvz1zTL75o+8zXnkr+u3sCmFw
2brmpcC38GCmYCXKw8E82MOfSZzhyIWWLhffmrUROQ2y9rlbF+H5xZ/AUzG+u3oN
slhJSxv/VZXQjPLyVOMGjPCHRjyD5IlWbUab0yoF8wVqEPkT9WTHs3j8NiqRsIfB
xu7bbaLn570yHYgGJfVwPGm56SgqXj5NTwQ79hJKSrD7HoGyLxDcGao8fKOh//ur
trb4gZCfJpwzAYKap7pyRIoIKWcaYuXbKlCBpMOOlm6b9K5u/zGbJXZm9wpxDgRQ
Yc5b5OKJPWBJT4UK5K4kfJI/CoBWCekECO6De0NIEj3BlXOmzO3jsco/poRN4DFG
cPP0ufbawKqPMhpmVuJoW7TxnMjQ28fVjetvOczRlqyaJsTcpDEptA5J6dwGezAI
KlzRER7nFZaQn2V3FoQqHU//nyAHJNT6Nrct6mKMVYJIJwZYjLxEUHP4KUvuE4um
iIrDTJ3Hd686ehjhMTfj0V7U/Z/Vq8iZPh9zqpY/Iwt4Vi5Ktra6oDF4Zc2lzzhs
y099B/t48gw7PHQb44D9dneti624bGI/ATW1JJiy8bWSiszwefSDA3hiC3H/3i6T
n1w6CWy2avAxO8bqJrL8yk3+7xaN6gc6z5agTocu6JmpYNp7oNBx7exSO/XTbxYr
4jtwoT6kVM3OplHIxe35cAo+p8cB8fOUOAORkK+y4ElFSPOKqGigpTWs1fi37VTz
ht1+bvi8QM+kqDoUeR0UAewJeFmUOXCuGH7FkT82FS/s/cg0zXsCXz04g2ge93B/
t7ltyzHKrqNTdXwkqp7g9oZbWcoanMdCcxE7Kb+9roJrPIKOw9eF0VcwFojGEr0h
1VNE4ymZ4kvGwSzKavbw5uTk1nzBKPPo8t6u1+9h1dLCORo8ajmIhslmYVLcJr9x
uUKX5rcc/byLmpq4rL51xIL8/Eozg9eI2Up3M5KaODyttaCYlKLEnQBl8drBaRej
n61QcYbybB648u3GDRGBG5RCDCj3D2LXfhAsc09Kt1bD+c0RgNn2tPIMWI1ypb3Z
cFulQcZI7xCkMJVxK1b2Czu273GBsoxtkVYaNyC/KpvO8m3T4EeYXDFpZ39SF4qJ
YdVm/I3Q6kijK7UCmJ4h22bVc5vY1LrVBxAZB+qFJU4swR5CXOkGHwaIghPrlU7y
/t5xMRp+PnSvwS4X9/NicT4KQXATlB6W0ueaTxbYlHfRzFqak2/x16YcrUEz9qnp
n3YEDDuAQKczJM6sXbRZvPp0XC/GUBxPJ4Y/xN7QzDivcGVLFbxb0u41a6KX/9Ao
zx1VJZs1uRbo1Ac5pGmHm4XY1/zjsx2dZwK5KrcqJrpY7gBUKnhOvDdL2CUrdorl
CqpCTgUqdGxhPxgKZsPB3oQTaSv1Zs2Q7jNwbn870jfmkztTuvKkfS2JVi512VPV
lRqfDIzGzXhtsnC5zhbiibppuLiZf/VrUiLan40xp4CPvfDQDBxDtrAbdMVLXrvp
BSVr8iS11lYq/O61v4XcnDsrcH9N5L00Ng3todbI/q1md0lMFtqHP9LqZZvzTqii
TE6O2nAPWyTxDn2fjqvw5P3R0KJbi7O6dA0Fekf1dX46JGafPJjJTo5mENXaxR/v
TlIalTOeGYAOR1CvPysKAJJHkgmqOQqAh6DRIO4TjYOJrQWj+tnnA+mv5bmgAlyA
j9nfvMSm7Mph0C1ftpqV+r9QG/uBnaKTZlx6yXGdHFTT9B5iPDZ8SBblmaY9fzOp
imGWI1unO2qYlVBEDCYU4BzOGN/AMthTK/bgjxXtdbvCI5xtWZnfemXTpmB1DA0t
l8Wc3lP3R9AjPcIvbcjfh/E7SdXWuG+hC+1F0h72u+zRiHL437xJxPmXX1E9zZQJ
hbG/78f8xOvZxyy6JHI/3XZmMucQTqmNOxi5E7JlzLADWtJ6vzY9rcQ6H1YSt3wO
biVHinGLZNqeiKQA4c+q0z4F96qgq6GRWcEiVB/T9HjNzkzGFCIXM37qy+iVuCWX
eh3TWLxnXNR38Oln/8bOJ0kwHanRzzd1i3+JdITFpwZKImRjotsO5KeIw/ATkUWg
7nwYLBCJT/fypfLINOnWrbyUsE+xxZ/2EkiGeJVYDhKsNdX4a2odh0OYxHAqVvpS
Uf5AzKWTwLgyXCVhx5e40xwg7c3TL7Kb3Ta3nqV+iz5gnMsav+6+hrZxjih5UjIF
fNogm4NfPsuriVVvjk5WM+2aydKEAyUTR8hJfc6puGPVFUjb71Rjnr+f89lxysBz
iIW6STEy9tJsFolXLNpx2kk0Cp7AuvY0nPTHAJ6ncc7TeipslquqUARLSn20fauR
+FIfzRnLtFwQNjXOOsHC8zjeFOesdVFcHw2wPywMUacKvjcaDcWOZPRUrc8PjjWq
0Z1k0yS3G2w7tzmUZwEx4s863VMbYv64LBC6nZ9K56bHWmClquHzW4K0YNzB6Oo8
QtMDZY145Fc+gIZWgxM6f28l+AtBR+k3Itq0LhuH+j9co3zXHcabFJbyp2s1HmRJ
69aAlLn4F1BNts9wPOYGSpYNZunk4hlV0BVbtteSndV1ezQ2B7PsUmpY6LOl+HDr
z9Zx5LVG/peaWVkie5L+xLoQYwXChWSwjdzZM7vEfpOfFLg6vtpBU2rKqpTF5NCK
nH+DyjlX1MIW0n1aEpKSmjYBEjazb4X+Xda4B/VGaE0fLjN4n2EvJ2tMj31XuCGW
M6aGuVwQMFfly/InkSaJ6VKVrkId8NqnmplZf4S/XatucG2d00UUhTZ6p0M7d1aN
wRUsZ/TZQ7kRdZ+lr6P0azv//pthxgqYjbWVGmyBTwPVz83RqnoQEKBu4TwsQoBK
IocLB43TXaBSkbPKOVeZf01AZ4ITLGIVgcqkIaa8KwIGTmQ495hl9PEw4wBot375
Fhq/b8/SBFK+Nohha6vAdCy0QiKFeaNbfy8rnKsDT6CZcswru09Gt38qLySv+SjT
kstbi4+CHigJv/mcZUZTuCIo+6Y78eoNAFjacXYw7py32MGcg84CrkZCkHQmJdhh
tcRI+gaXxo7nIJLh15lcKNzjvAOT2FGSa5WRpvD1Y0CvwcAFuMlO14eoIMLHnXwC
EzBJvkuVwLWYiG2QzSvsn8s/PkyP1kSaLnWcOVrPioDTFjFA3n219UA9ASvuZPtb
zBnbScCqHVv++M8BYwg+aHSrc4IpSoI82hll4Zg5TMimqr0V4eyg7+qX1Snw5uPP
FLAmO6/6Gul5nAZFnxKGcNg/701hfsSxs77r7IzjRWI31xVFgOiuj1IlotMVB7Ns
zXQPVF4NxUP5dmPxnn1Xw/mumHdsGOV8l6PuY5A2XlufHQq4MBil5wdzcTowsThv
kLZSaYmlcbY2FGkg1GsOXPaEr5EmMl2GWRuHTujjTsnlhTsjn0cIPvpXQRdsOT5e
EoEHy8A3r64R6LrLwhM8x6qwzQQKlZD4wggcGSDf6gNLMq52863kzHcTpswBuzHF
vWDmFj6/rJeb6GjepiegeFXJqpXUVFEHZUvzU+jI9t2TJb+RFsEaHV/UtiWsIJaN
KZSfpe4niwbQvGbIqUkR3Olxk6RVlwl+66aDySXgF44yx2o7FTgw1E6uPhjNI/8t
u1WMF/ZciUwxMRYUkJ/aNvyAOzF2/7cT/wtZa/0SyYJ8l6YSuPIE71HqJhI4J5qd
OYAiZb1bHUh+SuIxWUnpUoRAYEnKOOD1T9jOjv0D0sN4ligCIuXmU4korMgBJzQt
5/04utoyzCaj+j0FUFpQp28e/ESKSfFHREH+ufhRbbzuIwFhrGE+zOFzvns0TgT9
5/qHDU0ZfTqySykAAOqVfzGnoEoru9qYVvC0m4+FpDuJDhYo3jOVIGjz9tiJ/YvV
wqRJhlqypY0Cj7tPMGKy8y3ZvNnbSH1sUtPjmO9JwMVtXANIgT+CmlUavpBpoofD
PQlRFSm0rl2w2eJ5vZ8o4Z4fjF1KeAz1prGwM1fy2/Ys9sq0eyqtVAt1fXCi2Q4K
ztKxcPnpJe3V19EISLWaCaC4RVk4T/DpW+O0OrorEg4WM0k8LPconqUDh3uMopea
7VJinRAhCV+gE2zGw4U8AMhrGasxmR7A/LuB3cNNjpPw2dcEniD7VOvW8/YlGy+m
T8AersLfcWLswHDFcBXhDgrPtirYL0Kw7mPXuBzjgkVuvC982oleXKcmo1weSSMW
P4aJO2P2KCSLV6A5XZ5+hG/Z7H1pFLNpnF6aaTg9bcVRxiGDqQOnp6HAKmgrJjmf
YsWc7WyE/WPMD0CkVLrHHfkE1W8XAgvgKvuKBSIxxdEtAEhM5G2Aarg8IS2SRQHw
7INye848K0foM/V9qEfz4meJM+34vF8J7FChbOixpAlBGiY+Px+Mq/9+JUhtmnQn
Pmt0tnsc5kkr4HzaCnARGf78ikvhSd6+aF+qqcRiR5Q6iRaY5ocr9DJgUdMg064k
wNN5Xwftcm+gGZtzcQqSF/erBOOm11TqDAKkG3Laj2RHugX254f9VWP8V9+VYVHs
EmOB9F+4J+qVYkpJzdShaM3D61/9P7VcqV44UmpXB18pZhfdQdjlJ6pYzUz4Eawk
jNsj4Ck8J7MNW+dzU8a++wqLX8F9j9xcSbE6hW0NBkXg+loyA8Wb1SPkZg3aNnMC
0H0RjPspdME4RTwMq/MrTNBdOjdNlT16FF0OIuMDbgtgbxsUs4XGTPwRm9AU8qlc
3Cp+0V6SFOy2NBg06GZppfntFGBhUElGnIpxQMyNYar0NEG62bSbu/RId7QT9gdx
5APFZIr/bh4Yc74be1C9zfUzgWgUvIZxPAN0B8kJHPpuLaNCLXjwPCkPFEApyVG9
EdwW91G0sZJ8ZnDN9JGX8nSn4azJ8OHA9RenfSlzxHtOiauWe/MfACPBqtfZZc1Q
XPT8j74yKxj8sbuVKkR7woRuR7I6+2Kg2FELDz9ydVvtLopkvvSmPg15ythUbnfe
Rr/RJ5SSMUusU7CZuE/Fgpt3Ijyp8RNUdm/hmUO4eiN0GfBxG2mSJTv4nxdETKyV
h23JxBm9bCDNVkTztBOpThfJqlaoJ68N6MPs0qsnl0ih3fTuFdR/y1+U6E+EyGsS
kH93soel70sA0KF1wvfngFZxwWSsgh8d/g/nIASi12dQy6uK54os2AyNr6JQ/0r6
4IxukpoEWxJwuo7PyiFxiy8gS8tJAo4nQ5d7mcO+sNtnQs5iDrrIvNddvRtkPI1I
AUUb1zLf3EG2aVOzn1/OORUo0y4sopP/cbfNTBg8ezVBpi+++HiRzkdAcqCYlj61
Ni/mtMN5jkwpEHIhY6fUFiTCiDoBiFkegJ15x0CG9Yf1tc4cHfehFnWclfxhHpWp
bfsok/eOuA/5ApqlVVpL8ntPIiyJRvA9t3ypDKmJ5jjlZq4g+9bJbH6mTrArvBQk
nN55cLOtSgq0MWbR85wOkWOyvKgUOmZnNMZlJilykRb23i/vujqXga6x/2AeHpC+
rvVEBEa7gtZaQhAQBTBOB53D45uKR5AxHvDk2dEH9bM4kTHwFLQmt2IateIeRla/
Hc3rKB1xieDRZ9LCE8bOhtdUeDPjRyJcNPj/CIcxKHT8jMDMcxRuzrUvTpZBA3Ht
f0l8eZcpO1wLK4aNEawXxCAefbh+ZF0Xs+uX3Hn/DB5EtCywyknfRr3ycb0+oH3A
xl6JHQhBwE6/0eEFTTvhPkJV82U/wd2vRSMEEADsTkufJlPIb9KWIffw6W6eEczt
Fkl79OZOehKlxBLhSXZKSS1AuCNLPEvpuLleybZ7e005mumW01MHoX1ddvHaCmQt
4NzsjRlTvJRqHod9U+TkKZkCG9sci7sJBLNvUkT785VU06LqIeTnQWdkX+3/qogS
yy0C1WGghmEOkGf8A90mXuil50sbdBwwgcHX7QTUAtHYgu64kAhmJGYTYejDfr/2
O0MHMXu2J/U08UwjFMDwwNEq/hXyXmVyek6PkNPBFlsWtzVPelGeLVSpNP4/1sNQ
l1VV26IKDj0fpmbb6gYUHsxh+wa5doFV4X0OHRMzbGbySivxaIPJFWvH99EBG45h
NfGSCruxOQciP0ERCUvo9eUUl1168JbnneYYZUaijnXu80trW+WAP/LSJaoKUU/B
N6Mz7/z1uSNU7SenRTnqitS9daRLesmiGP+7YTD/VmsFyUc65U6MzrhdHyzhCSf9
Ps2KvRSwxKHUnVD7mF9ylJl0ZjVfVlgTfuM05+BEsmc7FZYHQnGJeWzuribZnH8e
PvBtgfX6fpaCOSGgYshQv4k2B+AU6+V13Bcvj3RxIRC8gpXNO2Yfm2DpT1uiisET
fFYzDT0AGO8XkAfAPMLlcRmbkzCXn00f3ZwuLmRu1FgdAmVwT7MFa8YsWCpgiLkF
Kc6SbFEEyKGIAyQJYt0+DIdauAe/XaYMnAMWAIDUUQpltk9N4+xJrZEWSGcT8cLa
8o3pfnIj02rgMSgdyZPwPU4MTj02e2HjjPfJ8vnmoMap78G1QHOM0mDoBdwWmYM6
W72gV6/R8yRr14ywWAZB3pKBbp+iZUzGfCDnDaP3GSDZYCCoUwaNpLuJk55OLUq4
YAGRrbVPmtSiaxAvZSNDp+xkfGCQD94Sydl38HTQxAx055XLgPYSwYUF6ip6cyYk
9GMcvHDy/4USkSTNnmlxDpRqvSzvGzlQxiQ9Rl19gQOAVrJlNoacrcEhNPX2JC/M
BaH4gO0J0xLFb/Sne5dQcWjllshwHb5QHo07gInuofx+QZETI9b0RYuGzzIFSotQ
ieindQc+wLhuKgI3ROeWmESQ/ljI6bWNHUlx0Wl55OTZ05IzIIvH8SeTDH884UPr
l7BLjcBcujsSe1LeHGTArp7QzjZX+Br5cVZhd2ZS07YwDmRRpxifK9m6B4YKhMT1
ENKJ9enrieVJwJctCF4VnVejaK5oj274oCjV/43pGQaT5zNe1AbKSYDAikv84qcg
D7f/YsuV6a8xdPu3FsIxENOZBTuqHYxtD1vjrAJ0/NFgUVsK8n8tahKyg/LpqntF
+N/A98qiLmBz3Hfz4MQNlAsbBRUFJoDGALkZXY8nmiGrUa29fv+XJI+UaEX8gNJj
JKeMqf0c55G6DGQlfG7Cyu0zIF2D/oGNFm39Di8n1oBCul173NOyTz5te9LNIUza
lLW9PxD795V0O648/eqYDpju/FR72qcIerLIHp5+FiUhzNYTLoAowbaR2lePv2T8
2Wc9UBpuU6HSxpNjrm0XRlFiL79TR4cEhVkgqDVtCHz+skqiyDDyTAdZ8PWWfG+7
gCkuf04yAsd3E+BIeMT/zac7vNJvmkpVu+VDDSb8/aT6MWVJH3TgK7oVcBZh/S6H
J681ZRaThmXjvD/dhRYuGh5gAf8WXkvZqT0GyZ2ZOwmmvFELVWs0iEmAD9jJ6ofe
321Pd8xy9UPp6o8E4KNoRt6o7ewdWKaU7avDNkZ420OFSW4mqFRQGTe9MzAcgVjA
IOCcaP2qAxA4cgG006Nax+PY0tosLqPQeMJCTHghgMdkBdSMzQ8i6yNcnlYCXqrZ
MiViP0Z0EFMth2vCEJY4q4n45i+hO45wf9okwYeEnVlOksoFYPdz7MeF0er80yuB
QbHY2MdF0cHVldRoVo2blP8r1LkwCOsmmf4mEVcumc0eS9eZQxBZXGJQIhF+zFGP
9xy4Muh97RB38XZvUz3YFfeOxPQp/uow5Bj/MYtPqaoUPly9RkH4lmbeGKoWRk4k
AQaZKspDGVkfqH5HKD54L3InCamj1CinDb8VPFhtoyeXEVEgX8Byppqn99oVIHAg
gUSWUnu5eYGNaPtchwdCsA2kU0Nd2RpNWvQMns4FBh3YAwdw6FjLQCaJpTd7mH8B
BSlMdgIYh0Rcs1ox0bZnb+/TR/ypyRQ/SzEx0CfCUdO54Du++JF0jAE/5L1e0t68
1rnx52kj2k4/r9qKPbJdosHUG0VisHr81iMPJjN5XBxYenjKvjwpVdX+HI45R4Os
TkgLiRG+OAVloi5Dxh/hXtYc6BOggKgNofRtVfHcKe/uWKwFTd1o7hem/gGVMPDh
+6K1cKIgE5Qio7wUSUZCl5/ABkJrINmoPyOZHkmI9i6qQs/g7oZHnR85ktfQwr2w
rxwjEvm/5+yAQZ1WjVa49bqzWrWWrhn8dsPjairpBlTYD2RnyfNPkLUUiCyXEh4y
umjDxswLBH5uv4CTZqOKDpRFltmosa1zOzzRmynv89KkvlsJM+Vckddxih3YV3yC
AGKcU5+QErRXl9lS/EwGHOzErlEkTcvqx5iwoILvsQTxl+Km9r11r28QwlfOKOpU
vFiwzD4USspg749BTi/XWkB9BGgs6CupxXiD+6qR8FtHNjw7ELfxz1ns3BmxnwFS
5IqXWTmluaW3D3+vmOBvGh00+jspmiJwKEp/TNz1kdZcdiuFy8WntYNWHHFZ7nN8
VyJ5e0O5lGbe57601/idfV2epCx1e/Jz7Xtz80BPmOcS+Bnuc7BSZt+7TXJrBZJj
Lie4oveQfhzCv4FZp3KwKI/sP+dXVJ6pz3Orh0al71MM99HDw6KFAWa2NEGvlNdU
T11hiZPhRys1MUCX8X/EYeyuHpy1UjgVwN5xCtXRD42R/C0HjskbNQ+/WIEi9VgP
SOzV87fpoEKxK2awC2Ly8qVp1dlHHVGtPl8nxGD+a1Obbdaw5hOPMFaKmhWcSsOp
mbQZjPh/g0WQdgQb8KOSVluGdIWNqaGMEnJatMHguds6Xp61SaqzXxYF0v0TFAjL
S+RC+qw3XmYoDiQx8vO0eFBlIMHuIx0cCAT8HVrL0+keI49YeDb0lTt16EbycMGH
XgEF/h6JVJXLxeQAXwAHV6mx4eaEP1D3aoKknJ0qLA2+S+jt73W1gJAyBw6doiww
qcFEUAjHa/93GMdR7ikf9DY86nRAw7XBn0Cm3yjMrhTKQVqU2qGvimYcUrRNjuuY
WtN3QoihWxnJkzGnf+mgV8xstDgtTQu58BhELNM3K4HK8uoyeG2Vv5uvYp528QML
I1Fk4zcIQ51zg2MrxO6fgZaII2Wei07inE9DoJ/A8MnulbRh/Ex88VyzkQ7Cp3P4
vgV7hus0VfimOtvIHQUV/OyEgNBDjP9uDbFl7GYdawBjXa/8Jm+3TdV4oTZvUmFN
uDppMUnugmC8caVk2SOahl3jhDxuwnVgn7KzzhEBGKPA0734TZwdGz2WvPTC5ZAq
K6C0T6aWX+VW/gBH6Sp3YWnSGj4bF3lGT5geZogC2K+TwilqakxyhAJRVB2rGKqI
smmVwq8DHwFNBUcSySK8mD38DUZmKCBafKnY2FaccH9dutjmtIKYpxbXvSV2UmFK
BZqdWn38DHn/sBuM7zC1ZN9rJeG9eILCBs+MsRLUU2cZZyowVjoHpK58V96xiv4z
K1MWvrxhdCseLbA2INXLICp3jdqRNHvH5TdpZDQFNgpgE+M0ic5jLJt8H6Mnqkqv
83BweaZ90uxB7h+U2t5BHFs/0uo1pk/3qzVQdoCA+39JTDmOtTIq8vqIAb0kHxaU
9Ixh96jbzPsSs2N5DRLsG+mKBYRRiGhzIUiOZ0AXd/8oMjCbwOsIgxhjB59n9/Q5
Fi99zWFaNqGYfk0oZHLzGb15Sl6wxnXioazhzePgD1zLJf18LGGg+uckQBly82jU
XWrIjjYMdozBiv5uhzHFaI6nmSb8gOzSXfGZXSKetnf5NtXjw9LaWudFXfkwvvF4
0hY1MYaEpdhAr4umLhHNygF3a+uNIFGDis75Oj6M69o+ZnBcqVJ17Sls0Ctcpt/7
onWY6TI6oURTVLEp1limqSBnsB6WxVuf5/wlVLD4Q5x/2JTE6ugMgbSjsQlv2v9N
GBv2SKHUMKRc+DHGhDFfflFAoVCumVpQTMJaf52ncvkgcWrOYW9XzH1KzIdAuFZD
YLLcYn5kUeQA4GgWkFQB6HdbOODqctuuJnPs/fLaYtbs0nSfzj/2ooCZr8YCbePQ
OmAhajX13ckyLNRwEEk/jkH+/atcRJ3GJcJfAJnB+uhJmjB0O5fYDsUtQnZZAvgG
UeK4cXtAghzzNTYTpTZEiNhG25hTf4JicE5si7XGeaFK+qTmt2e3VNZ3j869luB7
4e7LXLzvzRCqqgXBUG7wHqttdDDkr5zAK6I+IUGrTa75KanYBzZnpX4wcSeH/4SP
WFHEk9bQHV+jNyX9v0J7TxHzypOmGnJqV4QvO81MMLpgy7olT58v0yeHrLG2HEwr
tYibDiEHmHmKIVbzk5MtlSm8mQeeFjEwVnt6EgerZ74f2gJDSzODAmxEd0q7HQrO
VKInYGbIOunptTZvnCOy+k1xT4JQ1PMBwJiR19dFqvu7xPuhB9PcgB5B7SY40QSp
ZmmN0gVoyW4LpM8v+n9VFuVBUQEnMLfHNz2eG+nN+dzB0LwM2cc8JGOSvnjg9/yS
HbE8u1lZzYZn6NqhXWpa7kQqYtC1woXakJygxjSQV2Oz/zo3Tmw/TNn2ahZlsw1C
IUqKZKaYAzXIsvP4qpHufNcETuoI0cTYWd1HsozSrGuCdLcy52oDn1JVrNaxVsLd
itrBElBhkxLBuUqnf8h5cXOHKCo0oi8Zqy5Y8LV3cIcZgU3gwTmoFI7PAWM3fsG2
8TDy9nYGA1NGqXheRkEuyvUov6aNyZgPOa/Bw7/NjFp58O4wdhDYbp4W29Yo4J18
zRtfmOs4tPvDhFLxTulRhyZgGJU+tBQzK99TJ3R1i2cKQb3cLxzS+7aQVOmnb6Q8
H8e3L2E4R1kdnC6jUgZvcIDArJjcF9y+0Z3Q6WjQE+nlqLO90a0uEaqJAXrCjvym
uqISBUjJ8SpfbUMsYCDVW3k+/8xJFN5bASD3dxzgDvzCvxdwZwMLle/D5ZKZ7DUr
hETl1K0eEi3LfhrEp4t03OvjgOb/t8pe1PUpM4NR968eOtAYuqaw4XUKP4vIoA0Z
OiIco1i9OED5gYYV30aEG6yMHDP7VivkLWDrAynlAweBeMccaPI7kuy7qcYRVmFW
dLwbj3wa5Zk0ZvYTgj6yWTt5SX5w4mVP6euydTH47XhbxUSDxhKIg6leli0AXYR8
6H1+lFJ9kypNewbkXtQ0jyOWKjSZj19PW+skPbgpqM7yjvNVwxfBj1NNjhZ+ika1
OFGUfqodqPEOSmFyCdVEw79qV4IwrkIuq1lhJB8vD8pKbkqIdh4l1Fkyqxkio9wz
K2VpVMmHPJMwc7POGq4Ajl91YbnOd8G1cWYUukMPsHJarbRB32uPI/q4T3dowwGB
sURZxsETC7YaU6iNFFPBHl81Y2btzWuPYlcZB1nL0SkbP27nB0jxwUCzs4int98E
DXy02D+8fmV+xrMVz5pAU5CLwEL05oy6wTvcXMy0hPTpwP2LJX5HnUPbJXPSb7nU
UqiPW7IEKSeZ/RFvZSckL0IYMpKnqxaUjv0R8wRGGPgcog6TvxebQqHh8KDlPqgW
9pMnXcnZH9f/GB/oCnFxx8X5bdQFHi6Pmru1Bf5P6qaWlornwo7EmZTl5dv9JVTb
N5Tw/3k0L0gWgNJdp46E944f4hqmSfJPW6H1oU9j6VHFki/jhGH5Unhr2Q32eVgO
5PxZ08O2WizU8zxzqNOCNvWiwa5fmJUyEsaNVcxwd4piZbY1jIrKDH8zxQbM16hR
9fcqXgE9U7pdlIXraoMhsYw49qJQjLmUm8UCweITMM3u8VQcUW9xqv8sSQgT7Wu1
FsV6fjA/W0nEQD5Kq5jpk7d71CCdjq3dyM5cvZs8IVYLoWjKfGoPZptoXklvbgjq
+v/5WW7rRLV/fEu+FCvNIOLeAfieyGfjKkw0G+EF4SFlshSI5+r2Q2vFyKHR94zM
ld35N2xBdz0fmcCS4RgjzUdbBjg2Pw/BUAfwExcGzvdrOjNaonFohVlotDK9ZpNG
CfZK+P6JMTvjtH6coqjh97KpqwkAJJVI8vGmYspShaQFTiYYXGRj63pGzaPqoiuV
uiS7KpJ5mgjMiVwCrYkUpH/5MTJvHkYjYYkKScVOAG2Klym3Zvl0guZe8Up9QJ9N
eIQU9DSr56at3QrAYNAj/ZN+soEMIcCydohUI5bRM8skYnL/T6I06vXg+fDn6tXR
0BXLCbNtU3yB24lM1Ab9oFYdnp95hEQvd2sNp6J/4zj4alXLyF0Aswnfo342yE3T
uruv14Ynh9WkBaU4N7KgVNQd8FYk2msWjP2eIgMZuOi4rqf/MqzruDUFtRclEjph
dgY19hUHuype/XabZJsQn9ht8io6GuWiFQGme9+D7CvTZA9gD5MP/oFzkt/3rHNO
P2Z5lcFBXIFEGaxyl5W3WVqw5JBgMLohOozKlg6mpfe0k9qIlYqA0FZN1/hS5rg7
5mmvz+QDw04yS5xZCsv8KPeq6hZd4XluRB8aPjWK8n6vocqvu0fuHfovoDEXzUxQ
LwZcsq6K2fSG0G/4eFXETWmmzfKTReYnRyt3bqEc57CfHzQALAEWewWa69TqcjL5
VNe204pzXt5XP2Sp2tZKOmA0wW5NwHuF30EZqlYk5NFasq+17ISOh9MguUQgCVzc
FiSc/1+9JnNM9qglBikDeGVL5s3Q6muNVPvdkgIp6EI3uQowFQHP0VSVdAhs2AZ5
Nmvyt0oJhBjLqwH4xdLaGdaxs9Vlbrxwkc1SgLU8O5tcW4fKJFzsWUmdv63iCN51
Si/OEFfXRKQDDdDq60wPQKCS9drKWriOGYLpQ7ACc1glbJq/5T/HmqltHg6cnjHc
f9eU80vT24K/7rbrHhBUA797RuGdESwg+Jg+kG2+BKOmiuaEwev3ClbPBRO7NrH2
GWlto+BAR/Edns3XEJU+XC7YofYO2EZN1Qrc+EoQRj/FFaSORtTK/Bj2RqO8pMRu
GT5dswYkL59Ezco+WoLyei7OvF0Uukbs7HtAovTztas2kGbARA6GpxSJwe2Kvr0O
REREr4RfEr6OtQmZD3xGV7uUzeXEsBzuUUikhm7LY4TyRw9gmEI0FQKLtg9Hfk9I
mA50n75bWQ5yyrsLHmwBFUd5YyMEu8r0iCQ7+nmyLWwVTH2AJ9npoRrd3rPybDjA
fCGCd3BzDfJRQK2DbITDWMphJy0KB367jPWN0cr47O/LZkpGK9xJjbOTcHvgzyTV
vitIo0b92LNQzZ4r0W2yWc9tSC5zcp52hX34uSVzNUMn/a4gsaqhhLqAWTRzhVqd
VE5cnlTzlKoA+ROCgm66BojAhCiFyb6kBMPlpTho3AapV+6TcmGCggC+8J81POr9
mL+ockdoUhy37qxjUShttRCzSCm+yZkjPMzdQ12Jviv6HsDU+IByzYbUQmHCxAqW
9ucLo5xJI9MZ73st6u+n00WamDkXTtYFniRun4SVvQ27WEgWQ7B/PTzulr/Cn2Nn
aGjGb5X8rnQWiw/JZnzxTD64ZBfJ7SdTSM0uj0tHya+RP8r8DMA8WaxFmxDWAX8p
g2GmWgQrHsOqYWRJQM90c2cXEqCAi+8urxvh+fBSzVqVKLwMgVeVwfe10/dOGYF9
i+CuZKl5wjRei+LHwj4BUiOVZ7562UtDINHgfod2TWaZwERLDbuxfY5XXPz6HPD6
Fi8/obW5BUCsPyrdHNT8OUm4DR0aQ5ireh2e9CWkT+mzeHz4XdjPdR2oTwH0yMsN
p0QULK/cxQzlHfh/EA637BjxRGH8xjMAUqtvO0os/SMXSXwCmmMyVzqq1tIx85Xi
Z/6BALzQBiWX3xPh0Mh0bGuH54PhDZGFy+6N6DnKg+sPClK6Bzyjg06TMFJczkfe
yYyZ+OSBNQJrJxCc331WVYpa1dCXGw3uouHIlHIpr0Rm0DYf02i7jI7S8fV6Zrtq
JOs/ya1V9JxwAa2qUzXwiBAhSEDsLLP0p0oHCrj8rhElDNCy3DI/8KRnGAankK/E
PTzGa5TDsoe4ariy8R0J8jTSOvrV5GvD4AjhtXXWB6EJ9AS/6zMjaWsl0mfJC1F+
JVIIghDTV2tGgTrwjDbPUrmRwCd5PeIutlumZZmowNS21yTnMibDUCiuSgM5pG0c
GnrORaPsjlC1a36tL8eWILy//m6UB21tL/jCYnFUWO5hlGryzJ23dHrHYJorxu/4
ugmAUJGCBRRFIPvrfZNE5KAllrAbA48R7FBBxB/msGEn/IWvXtJ8aMEMWoUg8nO0
ADx+/PHTQrXfDs/9ZCl9FBJyE8cD4ib5K+GAxGZrlpMmYOZCbjBKNxeCJgvxzMtX
dHbe9oi01gkp8Wg2LSdBZinfySIhPg/SbTUtqW6Bc/sw8MIU00v10bOBGEiiHVqL
20ZQm+1Sx6l/9OPf2OZgMeywIOZRu/brH++WHn7Ch/Sewqxz4lLaKusgvdqbLT+M
FW2JkdEprdBwHKAbgJt5Bva9zA3/8358KpVUTmiGLYXLJ7ZCUm3alrvdtE6jHPvl
BnbxXvtFI7arOP37mDkn4GEb7sLLILiaydlvuOpvSMfKI1V5UuM74bpcLaM2GLfK
UHUcllgPdFbhzNRtoXDHo5r2A6henHuBvy3GYts0DLxDgewAypuANLvULBJndAnw
cMz127S7VNpuZqUe6Aqb883HkLYmeQpWRsq7QUI1F3j1fqtAwmOk1hvGb9X0T3s0
WC4sSTq2Oq+NZZKaHKUH2sBfk9hxTD/i0LWMz+aKCxn8aXL18MXq1l4CwPbln1gc
9KYvMmc7rocXP/dX0/yJ6AtNVfqNpTbHH9A3AXIa1l+U64ANNagcMEub8OWUgC6Q
WOFX51q07EiLC58gPBcIMCJewJvv3at07WfV13sMv/+9qhDtp8Cz29+o1piTCZK4
/tGY5inDzCzZW6QybWTcOiyVFv4YbhNcBJEwhXC0hrorDuxESD2/YmoLHEcIVdXr
JInTlKOccCVKcWNQTQIvqSDTvnF7pJdkyiCC9Z+jRUaczYxIJILMr9cskfeznUAH
LERbzxJnJk30be6CQYb59Wfou0nhrM7B9FUQcQinrxtRYI4boCKxXKjoraulUQGq
NQoBJkTmFLH1hozqqELFqWbSccI1z2TDYPw1Akv4evmTLfjVBVPfaB7TWEziMny+
ugJpJfODHHqsDuh+FE1O9GAuBg0hjuoA0taYipzuqLvBP+gfh9/mkjl2uzEybGP6
jpodvKBTY/MdGyqMRlDJ8lLEP8fXD1XsfmbrdX4+50wmE9GKMojlSDn8gAzM7nhM
luzfWfVuGHvf40J+jPvEeWmnr2VUycxLvNl1/FKKU05x0thshELXyQI1WWvmIrDg
lW+hUqVKAC3NlSKtqhV2RG4CDrOAzvz7hIjjuEhAzHD3YcDoXGROMXuhMS8Xy3BU
1Im2OhIcG4Yr30LRu6Q0K+Becec1lA9HKPFuIu2m1QdZRmt8wDrN/KYohv7VNEUr
pvCHmrSuOx4Cv0pUVtJCecK9VlkYLRsmkqlottGnOmk8WC+O4+ZMQfdXpG5mQoD4
2Vqr+tnFC37PDkwtA8zRIDkG813tRk4D6DYJjkWUz4HJsmPrIglaBgmDrKMDnLfF
HIuG7mLcfEcnmq0UGWZWUF7SROFcLpzHu6CRdwtq26tDlqNagU+aobb9AZu6k2DX
jLZ7S1UzGxnHp607l1T1Fw4Hf57FdoZjwqpaWWh0l9PK4sQYpc7fuxlrE5qQ7FFv
L10d5DBhY6wnSfepCY4UbpGsGy9W69QeN6QveYWsTyMmoOkzCg6b399gbLk2DCaX
vMEFawd9RpfsiBx0fhQ+qGpqXtjB6hgOVi8W/ezOUj8yPoTr9wDInOmUPq9yN3n1
zPMRpc9ySm8yx6mXYylmcyzgwbcj1xZfxQGn+lUuzXC6b2u62RJrRTG62ExQbBW8
KZ5+SfunYfaqwsGgRVVvl0wTikxTRnJbF0iNfeCzNgiEjtPx17YF+y294o+K4AUe
eh4SV75i7GI+46iSlVQi66HBWSj1eOuqB9iKD5H7wauRY2qmKQ4lzm5eHt2eddB5
BEVAcv6oSx0+3aPOa47D37YUS4+bApafWCXpP/wgYxgCbC0rwxxQTpcfCrQVFSpF
k5lhdrav3qaCkWMNo9BUwBouvnCP8W2TYfqEzWb8jETHVNUg9gYHLsv2ikIl0dNN
GNAsokB6dhCt+hWd4X+dDoqdi31fdkOAlCf/CjaFaFajpC7nkLGuShWCu7xYWhLY
csQd4QFRowVIlvQubDQSONQRoOb/jMuwj4ps02+Fb/tva2MZHxB5YxwQD7o8F/kL
bDSUrPjJ6c2tZz4zno7jdyzCEf7iewSPya/AniKywL1HH3zC3Hi5YvJBs1s0Vl9G
SjuZtH2KUEA95uoLtBSmNjAOYB/Od62E5F/z+S6j5ii/A4xC+6S9J4blAOSys3m3
2KaDOB8rPtXWYo4tVDIiwrTChlY9Aj9o3yDlZeTwUMFdaHmdnF3FmEPbCAhXlYey
4VZI01t/uivBdz+hHgI+D4wVyUWh7Sh17PJLo0MqGlb9pArx+QWZXPQ6CbYpJ6Z+
bzBPbGQdE1c2ZII4dTKlKR7WSPtx7sSB3u/Wrz1CImh3SICPbnAgdGJB6F9H6SST
RU53I/c1zIaZ/PTHT+xI6iSPulpqk36me5XGEoP2ocILIrcptZOznxVOMUKCnaxv
4b7bhCLpQQpafyECIw8SgyFrzk7/ZHq/ayVobtkp79RlokS6E5J8y3ZmhAwCo55z
QJA2mpHxjw9pBcXmTfxcZDbhn5/+DI78AtFeFJKEO+V5Uh/lPvXyFVP19kBrF50a
bM+D3DRZD03B1gPLW3JoMMh/V/Tv5SfwCu2lbiYuTou9NBiAjFDLiLtUr3aUFAVO
0S02fIQetybbMfFNDZzFyGJ3zpu5pY5rBfvUwF+B2bn/ZzfzMsmmHAyzCs+NmhFz
Hoz4SGaJOj4cKpQxAC7PVvBawXxSlYfjyjvYq2eDKC+Y4tNeTR9x78hiubeVda9K
p+jmK2h6lPe83lxuv/A12WeQ2kQp1Y9hTZvfh8xMmgZ5s7bdvwvwkqEOh21w9B8D
yv+Ur0Ed3CQBIJzjdmYDVAxbU5jqgAaKRG7Zg9ZwZBLr788ESL8rn9j7TjitWkdB
/uZPhF4eUkJA7rqBV+JgWhKv9Gok3DPo73u4RUzITYBV3NDDHfZJdi6sVj8V2Ot3
zstfdBQCj3aLeDSqBwnH3jO1X1UjR+lDJ69QG+8O4HPBbENfb9GGkcCNnveTyVQM
jrQf7qQOjY644tfbKmvkOQkAZqcGzy2duyddZn0bLvMH2Kn8rz+x/sRceOknE5eU
veWZ2EYbSUoK7xUYj/m6ImVuc4CzfcL05kFgCmwps4jB6PB8CiRWmFLUJfoDRCLA
u/PmcO4VPylPYq2KzDU8FYyFQtYosBh1WfBJIB57utWoPRMq8mcslRkZE0Hwb5Yd
7Iili4dGvQ7GeezspmuAzgKrhDDd3ilI7sJrSGe1od+iZBLo/mx3Aaf2td4DJj+6
dootZA3sglhOu67TDexxi+nCYfemuKG22RC0YCqcy4tmPFGB3sK/Y3qqbGHfp3pO
+ytCOFjfrqi0V+TTFQ1lF99b/lIqzhNZxfE1rGNNW2L98BlhYfS5vEmO7tDQzPVk
g7mo80AGQyJcT7rCxian5IZ0NbPhCD5rIxaBd0uOB68t+F0k4JUSvRtTk+l7T8LI
YwgMuwHDueFTQoYTlT1OLrrMDjWjvs6FIOKsufKhCShMarnX998ieFtQUoPdyPVQ
PIYLPwjaaUtFOC6qOq59fx8HU5tAOV0KV3d/9ReP42IMY5BAvFSsD8L9z0Tlnpyt
jBzm2KiBcCk7D68qmJGJJMqK2LJ/9OXMELkx+5+nTLFCwucjW5aHiEH+yYSkcFho
8TwGEGCUPw203SRAOK0hb5NQ4tQvJJJfI6Dl4DorxHzc0B02x6hX20aA9oHMR5id
06o1nsU14qrlb3D2lDR2KBICn5pHuM1L1TJkSXmyzo6FFkLSrmA5OQLxcH1XqnJS
AAH10gZ/8WV5Nq7nSsrzeejV14OlQ/ViPuTDc/rytC2K765A/SuCMwk7JuQ/fkqI
rV3BHRkFjbi+DXqI2w91EBCI39xn9srCcK6IPHrbDhNu5xC1Ig/9kRtPk1bq5640
0hiXg9XfG48mW+BQmCVNODisL/msVpB4cQb6tWQ6XOyqJXLJFcZceuzWbkcoxJkD
HUXyqYksZD9dMmMi5z9iR24Gjq1IkBNdwP424paLpPxreWjLHoNWpH3+KWLjP6xh
crnrftqk7kVJo35ihg0DxaMGHu/ilxzV9wI6ASmMCn5KurHCalt0rVRJgv3Z8vSK
QUIoPBzPM7vJrX113I89XrpHxOnZyVfvd/4U6NzjQh8hX1/HrSjnjb/r299CptLJ
fihlRraUGQAy9Q65uQJQlhGKDY15tnYTfxBVtneSaapWTm2suGrjjNn0TKvHrYRD
1GJny/2EPN++c+4mISMPyx3nmmTAoiLU3Mvl3UB+lNNIl9kougEgUb6Iw+tU0qd3
3FPP7GLen73zjMCh/U57PZxIjXLfDxAOzX5aPkgjlOP5sRwtSaQSQm6tIL8POUzG
RTVjG6YEH+yfNkEpzub0FGYnsRwF6NBTnH+iwab/aBkS1QsOsIIMvzxt+56So0j0
7ah7qNCkUyem85orq7KPwoerBNX47pANJYSrcUuG8bv3LlSRItanc12nEPW3ZYI1
M0dRH/plG2E2gMhZzv3+JKXxtr0k7ESh81uFNdq41ops7+H6pN8FqX9OxeuBjeM4
88qdMSn0wvxz9M6j6QfwQMOTGkDgDXJdZq78FD7qJ3Vn+Qhy+nSJ8wabkQeGVZZg
DGc0kZFx+CzoPkoZjUmZU6ofsDYeczq3Y5IX9WMEWkjSQCFkGdel0N2CxEs81LUS
esRe7A5ySTOhN+WpGelBaCo4Sh7McIjR7DbN7XcFy3IrTbYN5n9GlbvUyNNOFILu
67arMdGLMWea4RVeYfxhcpgX00l6TSO5ZpnTQdrmoF53T3SeU4Mm+PUbT+Sz1hw1
nnKayoChlArCuTD6FVDf4dHH8b8SQqVek38bhqvsI9BrFrcMWlPGwRN9sr8LlwXu
Y/xU5nzh/6Nqr/wmJraB6ntWrys7rSgGxvfqm9CJnx3FOtWokebArpN6LLAlGw8/
/+PmunaJvhUnPoY0CRkgRIzqq52X5CEb0k6sVR5voKleaMkTIVhLnPsZTHQr2jiW
mg34/4TgTTXatA6exhW3zBmfBQp5CXVRQqxuL17753EwpezMxlypGu5dZ3wuNt1d
KkN7IIUpSQwcm46mP8X1CZuk25J0/A9gtnzvKlH9mFTAoK+hAzTYdrmUffu68/gL
gE4ZwiExhp7kbVaGPfYCtdAAV0Ndz8bFyz2VbcNZHKc2zH/wsF6KrPRu49Vnaqml
oGg3uhY83tZ1LaA4qVn6TNdOnBKB7OrVVDRQ3EvUMOMe9guavQYhFbW6LjvOm7d/
I3SJsljsf6w/hpZhL0tAZsGQg5GRSTyP3C60SZ09JbcASf2l6EM4OuEYQq/I3oGs
QBU98XnVxU0PvYlWq4J5EolvMy/T43sKAQ+JMCWVV9NnZQujOtCwl7KXnWIlDmi4
s+9WE/x3yinvZSNqUzWPbREDZjg1uuhV4Fp84vcOuYIEqHr4NHgM7K36fn/16G7c
cbACDOTcdyYXWnB4ElPcCktNNpmS3lYa+0Hk9N1XVk3Njc4J9QXR1YjfL1mrLDr8
l9TPFlGJvS0LNRNEdauVOEC98bF+poT1cOxx+hV5i7Xb/87l3b3kj0fevWJTWXnz
ta3ZD20lAhq1v7YNauSq3ljPB24CrZYWIL25EM+NCxEeEaGqn6mjqS1w0SQR/NXD
82qUvto2OBymoDCK8xVn9lnEm0uNoRN64A9Gna+z0tyYceB3pnEhqxKlQWZeHU+Q
Tj54fIBggzi5n5fCi+ppiMN/PHa5Ziid1gLwm3WdM7BMXrJ/YZci9Ey0ICz+Uz1W
ucU9DNQ72aI6OEsL99kOS7h0AFG53sUde/gQ4dL243tTR+X2hHaYTokCFlJFaeH+
SZ0CEiGfcT8Y7SNLaK9xTFEBLq+xb/xjDQ+JhhMR9LOHlE/sSoPky0Ng3wf3ezEU
HHml96oAh5l+TEL6ZdZlYA9uUwwJUxtZx353v3yFMYVb2cLdRkTMY+TpNqog/0rr
pRfZVcHqyYRUGdSThxRPh070mCJrpmPv6yh7LdemTWxw77i9wCGe/sS+I//b4UXD
LpMeylFdmnqqCCIiieHneyQKsegIXxx/gJoHXG19gOef4bVG70VWEozcmsEDrzv0
6nPIvtm73tWO65YIeDCJRgjAx6McpLpGotKFpdvl7PC9Yp6DszAUHMIlKkFDxow9
tJJHps9vqwk1c4zIRFZFWexT3y73Vhpu4j5eZBPcR7Of+8mFK94sqkwg0qLij2Hh
wfRRulOvYW2JAP07neopA3KRdun1nHZXmS7s4e1LDmKW4V/4DilDL32w31UsQz/w
7aSG+wN8f1W0+wiUZ0uwUL9edGsOvlzOnBfU51JBZCgO7VnOxPGCRFpioc/tqT5d
ueTxW/XQdkln/X4FFcOrVNke3dgXQU2yH7ztiBXg40v93EnhLd8c+1hkHU1hTLxl
nf7OswJYzvKj+GpzD38d1EWgdcUAK9q0MXoEKHrmEhBp3rqlwsuqXre+I9bSzMyt
+8MJYP04e0VHWhvsdH9orxHbC3QtvoEtIPnw1srAIvNgqaZYJyb8EYnqSt/A5JUN
r8CEWEQ8mvCivDoeXVgCzob3PWRNxoz/zEliiaJ5rxYk5ARwW1bH+q+KpsZAFIYZ
VA/bw0pIATgA6GT41E7zXJyli2T0Ubi/cjAjocAN76ORIuekgTSugWKRTM8r4NQE
PW6LtRmTZGRwLhntZZ0jBTxrmYXSwEWMzi/7PLhnIHRMaJF0MJes/d+P2V2gC8UR
SXVnSzLNbyTNYMtvsCFg9KFVZSmTWsPJudL7rCjrBr6lvPVlJN8tqwvy7vym8Z++
4m2aRVPx+TRuriokM1LIK/EkLQbeSr93Ocffj3chZPp5R/QOkDy0EwYcuxg7/4M8
9DJm6u28b9Jmm9NEjM3cxkowT2ri3MjrCKYfgAgMNHjid3maYk4Tj5/gPDiIpJMp
6ZkpRMxy9ydaQtxr8x4o/3QzTle3KBULrDSMnBdMwFovh78KlvEIDUiOGPYXVPmD
SKtDvSeDzA1YKOsqFTjfOCF7isy4FadJKEyg7zbvAkO3wGdaZCZOWYOaj+4gh5G6
ppZKATShGurHa0GTZ9YZGj6lPr+dU/jqHU+XMbPAQVHR7zJP3uCC1GCWwacShTid
vDm9O40Bud7powE3VDTxiykVHuarxgKa510woFl1r27MjTwCmdk0O9GwBVn87Dmm
6QwnosV1SFUS8Gfy5mkzrFoPImWvtCY/4PDFqoKU28IVFmQoW1dWEfremwl84inb
PjhxQr8fuRceZHCHCeYIA/sgYIGnajwOy2K7F2A0y3VysoQlE+R52Momj81ms3YJ
1M83hZe1xUVsJSTu9cG9Fq0mzc5zn37gFJVDwQoBpzTBpV9E79yGhrJubb/0JOyq
RY9wUndoRfc4YSWepvEXsGglsKIeqeD4ZHlE55Ae4f+e6GaZrx2RdXsp1/dDpvs8
4qqGV9zk2hZCqoQULlUc96yT/EdyaAL6QuUdYylC8XyOQb7cNL4sjWoLQ3I8jJ2R
BVw+xKl6MR3iCLzZ7xXYZ76WsFUEHC4L1Y1iri3fL/Nfgo0+MmoizfAVuBm/uv0n
jIFdR0MA0dq/Rs5ZCJTr4hRug9vJCaajbOPUSYoiZF87r1akzWtxLzauhX9xYXPH
AqJfNMVRbk+6xF4B1SkE0ldWpK7F2O39fS6OBhVCk8k3RMA6SL5m8n+rJwcNeJV5
BsXlBhoPJCofLfqXHeLF57ue3IUXU9I7eVnaRUxvyYdAGrCCjmelQ7vxPcCNsCa9
Lo2KjV8d8qH4IsKbdYIb9lpLvsNAOVlZwl+tFBkCiIE4F/Ls1phJqlpp85k0mJlk
r7IyCF3j7LLemWQyfPsv6bwU0ZyXC7Fapb2WfmBXAg4MTewLTuDG3ZSc0e6J+Dk3
rFBjinkc3urSHui0Wl2LPDNTn4E71F5uy4o2XqWSYV0p4TxppdEOJO+wCfsc9Ljb
U79n6tR86cqI4ZxFaCUMcTadFE0w1+RS/5ipBW2BVvlmrSiTzD0951wIvUylP7d6
VZ8NtJYbrXmW4NdTwU5/cMRkU/otlNviyf3pO/DBHz7CjfFyNpHZ1gbLX3MbUFEz
d8pFRxllWhUm9Biy41RCbWHwZ0llISVBEjpMgFX/sLM276agnaPm/n3K4afNdVia
fkwKePeGWhaN2w5YOFOTYVwZABd0pbjCJTIPIWDhYttE283wuvt3fh7hPhObHAMJ
sNAHqphA1KKCAUS+c+DLCFX05WDf6F2kt2uEikuOzJovgsUuUJbjBPPhRoqvrnTl
Bk9ejhtWoANPihhmevvIaJhKpX2u+//87cw+DWIUOXf/v6wxg0EHGdO/7yP5sLAv
naozDUjCkkBuimLCIFIj/b7etyP7TSgbrKRJuZWpp+DSjQlFysB0NtnvVaiOs/R5
0MbtS0a9/15vx4//hg3mrw5injK+LQGdwvpHfjBTrsOztFD6qnxHj55vMTkns/AI
xiE3TfjSlXU1zuh7ymYx0bgHzEnhxjJwD+Fr8OHK76963BE7PpNyWA6AVwq9I0dL
Lcr7NTYf6pgKA0C2mJpY7LxfHjpuV8galbjd5/fmSag=
`protect END_PROTECTED
