`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8w579+O91KtEFt6mxifDsAAynVSwpQbOt+Q92ICePmluEnMbzfljmQt+SB4cqL0
cuRYmzrJ2ZnPihrQDl2S3lXQauYLZushEbOcBrvV++wlejDnqoChCrf35pil8zeQ
5lOGr2XJjij2MVidYanG/puCugfQYloLByAjiro+7Yhi4Zu/IgLEou6hZaG86tt3
9Phbf6kp2FqyfNHWN4TAIe3mLCPUnx3/Q1sfvO9AHPYIDSwPWCqpglSqvYg0HuWc
HGLJiKAaHAY2NpHkEX5tpVteDbhJ5ZUxxt7jBJiGpHiC8JWC8+zOuPYLwWrxFjhq
4n5pGGIzv8CRqj3t4FvFmxk+ddCSDpuvnv25Oiy6XfRLulnJUlgRnrUJmZg3mJx5
8WyxzRgpOff7T16SYrfmdTKMqBWvCEIxDEq6Cff7LgEktj42OEhSpLb1w4ChPl2d
aAijMVqVndpi6VQqGfhIuM8DOtB6N6BnFC7plGCXyePjjgynf1AdLYklZ/gd2GH9
WMAFSn1DepzHID4gC4GubpntRWCSLLT+L1MBQCeu8wGODTCfSdqZLwwHyiErSzy2
J2k4Zx26OxrbO5yKppQJnEMU82bVI34m7X+R6l7mLrARWKKXPKgEWdXrVYVAgUe6
xj2G0nhzKVb++BPmnEhgWCXb6F/cx9EitgG0Gn0qWTnLm2GndnRXe/c5xLvWlAra
AY4AYKbQP/QNlo8AEPaWZi4GUb3Tq1mgOT3vnNpzdaEIOIRozn4dKSyIp3PkkCN+
TuRHoKXfOYXi0kYtf6Q6d0MRi44BSalQpCjhpkUGfm+SyOk3ReDWLLa41iZzxISC
DNtgUvqsVfJN78lsWsnTirm2LjRqCvS8QaEU3bYNIsJU4XKMhPX9v/fBI3ANtQ5P
UiNO4LATv+X4Trlvrwn1qxcfucb3d2JAFec+Eom1rfoVl5jznaM6KsDpM4nzsDA1
VJPY0tz/NRBN1Rz8UmnjMswKDuGAV0mR444ZGltiBdYPoKcznq+Fjv5c300aRG6V
qijctxxd0uMNEqRgy7OAV07cHXYfxTt8iL/QDjDNKDfzvegGmTPDjEih7+kYx1dz
+0x7CxWxAFlMDfRk/18w+TUJY6MV5/7WEnxPEQD77MrISVQcCRiBPm+WwNO1KInZ
6BLrocpDW3MViRbtyTOWFMEpa3gYv9WmdvWYRw+kSZzntCNoffBv2GC06K6yUccv
itbgn/WmKvoN0yo4st+7nl7Lxv07wBREAcJnVp4HJVOPr/jLfbWHJC8OuF/4Nqx3
GNcNYEgdlJg2UJj9iXvgbfhcsmGpTgiHuhtBlGfbsWInxX3t0PHn6VBa7z9Q9GyU
lNZY6/q0EFw0dGFh+pLVlACOyYrGO50b4Ow/FAwrthUR6+BKgPckguKD1mxZxCwM
Uxi5e1BtjyHIdpLIBGlz+DBTQANQU2CR9uFBmtoed7mPAKNoxyOP2RcNVFY3a6Sl
SWg1sK0Wy7hjksuOuwDVx2Eb6dTOBOi8j89GGujbzrg/Zpa7ZDSrXlZ7W3fJ1Ska
pROX/rygRcflWmuTxSt57Es0BiZz7B4pXgXTd90UYsqvngcekf5SvIuwBUH+6D10
`protect END_PROTECTED
