`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLymqhCemTymOGXvvkeDh3jYMdS2TgbjOmJztY7U4O9q8hEKvOFDq6+0n1ZgXk+l
N2aUYGjPdR1w7vmyKwpPIqZDqmwCV20JQc+9A27QEMY9aEAvUu9W+0CdnBbm8nZB
gskzWWmL625yk2+C2Texy8jDzlyx4BT4/2Aw6AAZX6CrhJ/6xIgk/KE8og9zMl6F
AnRlDT/aUpEZv98ESNX7puSP8KwbW7i6uqt/tdnQc0bVfarZZ66zmQ8XmJFxG9Ue
2yV5ygvSz9rjHFcXaA7Gw2BnfmEjfdbEcvGadm4W18ayQfUMqrO6n7ivmzoPmOpH
qZyWJGg5uCso+gxJU2cXHEHIRcPeHiJRgUVtOncFl9Zso658sbLvGsCIxkVm4PkF
ACEZf5NwdshCvicLkJtp4nh8lXyL74gJ5Yi9HCkD7vicG8IB8mFmO94mljjSIxKT
BAH7JJUI72pL2ncy9tLXNc8TXVLjODVj5lGqYEVngEu3ycYk8zRL+MujxEFGZCFM
on742EkaBI/vNHElWdBbpBk7v5VyJtDfTOREuuPrJNIrL/k9zcQsVRUuOYSeYo/v
UzWYnd80MGuOof6RDH3m+4u0AxtRd4HbplGIuiJIIN5xaolSGLb+Sxa8Lx+BBGnS
G1el9j7Os9Z0z9fUSmStPKCVAF2sp97GuGpBT7rO/38oZ+jjASi/avS90DlvknAi
i63CIZwqN56lCt6tuRumZ79uPd0q5i0CnIxLveVu8QCE3BvVUlfFwLSJUt09mHpM
SCjZ0D7e049495CgUNR8SxUUqEfsHSlJ0vKzE5mZEcGHevmRFptqo/MKTlyCqgGM
wTeNOUwdVysWwGa4wTy/LziWa/KLV8lFV7tVK1qbBGvtafdP5iCin7R5RU2xG+gY
UKi2HwgMd7TtvX8hcA2YkRplZUa0Q8zg9+zOj8X6a1pS/7ERmE71WUe5VKJdh+9b
0zrIB3ip7+Ai61Fs4bfSb8PxURiKhOplRjtbzAxKMleve731c8ctDXubwYvcK1LY
0PGNCrXl7M/8ytIRsem1pG3E6kVjq++ljvfwqTTBgXAGJ5obsgL1PZoPezytiWFJ
c9ybyH2blYYwpLHy0wiW8yxTuqB3Q313B+Psz11o3QRIeVFwvbVgpndBJGlzfgW8
mpTNHlBtgeSuJKDGbYEtTUBqoFu0JDEtooQNEzTzJaZ/DtyFgC0bqiig9LJRIK76
jZeZWjbpph6QMQbTOwV3Z0jrUumnHep7GPZeiQhe8yErQjXtP0H2DOJEvFGFL7u5
79bH9c2qAOk5os8HMeuBNoadeDEbFtaKvSVfKzMbuEihtmCXRyNCqAq7EuDLeBlP
jIEY3ZSTgySLQTFpA2eZE8q3IyOjyVjvC0RamLOjsEIpL7YcOPTO/oUFrnFbHhSK
KmuEsQc8Ck6ebn58bmA24Q==
`protect END_PROTECTED
