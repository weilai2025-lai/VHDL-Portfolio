`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4KQXtKuONix0Ad6c8HOr8/osTBf/vmVAXn9ly7XjkN2K5aTft0mtjxlnuTQFgbl
/+T1wz7Gwm2MSUc2ZYuOf2QvKnnLaWJqMktrLMnn/nuBD4PZYse1zrVNpNT3W/iP
kSazZiW/hD33uH2bwTSUpIAJM9MrxhUTlSv00bYQhcsu/Y/dvQErIcbZ2KiF8/kW
HToZF8mJJ7kv8HxILiq4JFBPKEg6L/elej4MIxGoOPxLFKQqkHQbNAVqhCYP0Jyl
jNPQrgXQthE9k2xD7cAf+ytNEzIEg0xcdAG5JQmxQMN3Dme9xKgKdEOERfJXdOKU
RwBGdmbSwRjRU4Y2QxZIsG4RM0kE8pIeuSLXrggUTIqJxQEU1qysTHMYL+qkD/75
lVLhL1Cy/AR3hwjrrEeVb2XTq9ugWOinCJ8+PCagrVXFTU+hKhMmExVmzwfXS3xe
XPnbPn8WO4LQ2rBd4P6iAWHlpgZJqxTY3mRg+mqOIOQtIdKrwFRRkUYdM5fHthOB
`protect END_PROTECTED
