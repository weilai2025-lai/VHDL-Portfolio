`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwJCa1IEfewfnmT0aRBKNkhyiDc71/CGWWwQv5Rd5GZcBUhNZ0yLCWBIfPnq/2gD
+OXUZRquRMxJnxmi5m6LJfEOX4weJNkqSC0rc+YW5V7469UOhGK+2A+mUYRTrzp0
WBKGRM7hIdKLtGGVM59PnbEUwLN3Xm5wn0c6B+OsSVTW199hTPqoeyyaBjOrlHcx
1E7ADpJYRzPJApc0O/RH9JqGQ+XDOfZwSzyxPyxHQOpbuyBSTbGRTJSxwGYhJ0IH
l8W4oABjPbX4atkkUzul08LyTQV5q1NSt1SJCaz+AfN/FuozBOhCDeuu5Ig323mC
gIHWJQ/VpAdinYZ/I49s6rq8cfTtcpqdkPRYNzULCxEj2/4s26qbFPLFQsRCMSmR
Gqvmjaimj/qWuuqAH5oo5qNQZ5C7Nzgw9aEHlZ2Kx9QxoxlMbHk2NzAejgYgUGMt
YI0iOvNP/FJHJtLtazapNboGveSlu3ik8rH5C/iwrQNW3vLClNrKfXJfeXKbKV0A
GZqbJ5TGQYOEANhoorZ8dyLUIle4ETf0VatOlO1cRSkYnFdbG2DP+QEC/tY0IcqA
cOU4d8PrSRzOwRoJ9dY3E+SmxcQAIjit12IWPSAKvGu2ozjMVWXF3Qmhzsen3KYo
uELuL1EbTXuO4j6GH2FQmZU9o09vb53+ud622dlhg2kALe+AmTT7WEbmw1QHuVYt
n9SF2HZ2301lzVKWf+m5oNNynFDyfQWkddvKipSEJ2dATc5Wh7V+xaBybki/+vMD
/GBgARf3AqsFvVXvFQmNcG+JbjzV2v7DsTZkmQuY0EPBZ3uPG67Ce7I48LTBWY5l
FO578aypCU1s2ysTN85Ksv/06Py3/SwgbgVtTv4m0iy6erOMh9OcMiJAB2NRIrr5
GYTNq+XoCBXuIH2CAmyhKKd+R137DiP8zHJzi9bNshcZzVEEhxXjtF5nKb+ZB7Xj
qVVEKJY5S2bhIC0ujpjmM/eXgN+yXTfVNfV8tI3zOBRRR4v5qOzqrkHiln8CKA4X
0oDZrTeNPhzi1T3grfK+hrfGEQe+j3JFcR/P7mIAZgnotffhxf+GkfgIWDr1OyrZ
0tPcb66AGVVPvXY1IMQ8ZT0hG5AbcKW95ojQGi/mKgwOg1158ZKutOpfJ17pbHNr
BqXzw0H4HjI1Wwtm5ip96BV8bXOl9e0Sziy3hqH129pc3j92AMSDUxjTZS9MgR00
LYp5vwABeP8m/UfFx9k9X1Gb03Wjf0UIJ/NE5HAqnM5YCkNQQtTUXSySMBo6PUSD
4f+/CLuFhah8qd36uCrIZiPtrEVXQtYqqVQCQubUxLoZfRm6ItbZzbMZ4a18K9mC
LeovGVWP6qoojsNKGBhTyNrpGmmz78Q/cyaPeIfXrjUhbjp1KG9sfVs3+MzMXCGS
rP3MqOWFunyMOwybHrRolSJu/g24oNVuZsAZoUKl+pHX+1OWVa+eHZqa180b0U+9
5aioTDJHuMCYzX61AaQ0oZvwsrrc0iwhPvB4/tau5hDBuorAnKGlJ3vTLM5tjokK
+Ts6xLECDR0ddJ9n5L2bBdISdsDls9GtRC/mqnTO1oh5Txy6GlWG8Tk2xP+OU+Ln
MxYRy15jatPmKgKuSCucZlSodcHUU/ePZkte65MqXO2GeBn+hlTdIq9qhyH1iWDO
9QVV8wkXwZw/3Sf+pmrFoN/l4XVyQem92sHn/zDUW6McfoDZJAtr2MH8dBzHZtR9
BpRT/aaIjPmDn1JCgxtOeIqmAfuWqfpOF1rj3qjW4EU6ikiuWfo5j8yu0e4oW7VD
5knmoIvaLDYuLZswbQ1BJHMwkQxDu2PMYe0J+9Dcp4xMe144goiPqA7eSZqqRBkr
SxmTaByPseSK9yzQywBqa5QTn2LhVNhgVn7f2GjgnLqr+EHczC4dZekNpJykJQKC
927kLoJE0nYyd58NTlUAMAl7sgJwZuSTU8+UAc924sDMJGwhVFWrjn3OTXiNt+gy
Aw+z2JCVP2fOceNjoxendd8SytU92aWw4uF5nVb977oYEaMNGjk6F3j8yM+5b1GC
UMi8f9WCb3+v560E8wzXTathM0cGWGLW/luHUzJQBNy6Bn3M/qBA3EZWtasLMXST
WhdIfFWuaKy0IINJmBi3KtU1+n65N5l5Dk1pNgPFELormSwKnuw3K1OAS4Iewmka
kXU5j07lRK/QEI1tG/D1ZW2UoTSgV32yT46ps0CY3cdH4k1iLsl2apJQZOhkMPyi
Z5Fkeft4ZunjXE7b0s2n2UOVqdXklQEPWLmvdJ5oXhpMwQlw/js/4DA61W7kRSCu
TJ0cGNze+vFF73Wo+XI7cT2BrApIH6H45t9RqVQTUkxf5O4XDDEppMiQ2NITJw1l
wTUlK4gwN7hUiAUKImgpJhDJ9YsSu4JGQ7E3yRfk8ioCoq7YIXCYySCVTKCnp9Gc
MqSL6l/XcaWjqQJsSIDcIS+vneRtPyYAF49p0sbBWe6nFsvyuOQxrhswwnJBVmWG
E7qZOUfe299XCmvaqaYMHA==
`protect END_PROTECTED
