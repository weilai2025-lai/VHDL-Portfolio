`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rbduEV/Hb3gJHw8za5ChpvDBS0Da6IEAU2SUfDPnQUJHu39OlyTa6WG40of8E+pJ
oZM32zXnx1u+vip+GvUKMGmTWA/evOAjQxL903yTO/ThU3m3s5MPvcBVfRltXARK
WFWoEaWajbjW+Hhf7/0CMyellwBGYx4lfQ19gVW8qdT4OnVDp/p6M969tb+b8gE4
q+0ULGRPEZSIYj4QgwoiGDBGEG/9/aJg8NRNiSVU3LhHgEDhD5JkEayy0O1Q/R0F
pGk/UNakF/zw5sn0UFQUBPdk0Kq/GrNsiQPU6Az9eFrewTVhxznsqRKJQmzGr0B0
V8XAH4d+rBoxzMYvc6xOD+Smxrb0nU9HEMEIYRGr2+ZLdQ0+XpuEFRjIsEzpLRfE
vvpINAldmCokkyH8/v0I6xpKUCWwn4QetnDV/z8cuTSb+HCv72x4RYpfORH0bl8D
gba9pbMscMiv8SC+VLqSf5Z1Fmoifwmw5gtPbg/+UFkVa9w2Hi7iCtrQ4pG5M1I6
gthXFvY6+R9BbTTRaGUXJyF8JpK8uSFt/RJfPLtrscux2DtiduNIoqawWUFhCS4+
lY2S1dTYdQx/kktFw0DBAzjYk1nt0wd7VHIdS37UhZ01gypzVl5uuclgbfAy57hN
1Aexs3mDiTyxxQMDwlTMUdX2bfu20XN2lfCt/RO1qf4RN1gwRBVOCeYAUHtwBTjX
DcPFqNzSonFJxiuA7hv9/8/WxN52RQvEIstJWrPLi/DUZ8IRGTysM3EmIE+0msF3
edvxTzrdlcEyJO8PPxTqDelOrJEN2t/TBdErob3SpEkE/FW1kO6HlP1yw6BntYUp
5/gZpztoF/4IveqLC0jVzipwJaZN31Ehv21Z2nH0XIGmnvnQ+i3My8ROSrnKg2Yr
V4F5IaRcuV023RAAwYsCvrDyIGJ4ThTUs/DKabnlGJnW4XUzXSqWajQp6UHgl5KR
CRkAkCM7KQqL+8kKWEvHHuKiDr5AnINwDkY0+RuoSaAl860MYUHz6Cl65Wl3Epyk
sAEVJs8imnmbQWbW1f6xM8Wmqfxz/PImkOhJMm2nT0vxu4iRKuCZQk271rvnatwT
`protect END_PROTECTED
