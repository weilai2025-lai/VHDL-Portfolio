`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGS8Cgu70xE1vCM8AbWwzPgppR1fOs5LysVvW38wBIyt9tVZ7WaaJKCBRqxTYu07
Pe3m92SHziXvkIk299xRpFq+6UeZQjmIjkGM5J5oJNCSAsSY4H/hVwnTSrPPxhbn
N2VudoT18WnO3M8jYUzQVphqlY/c2Qmzm5WVd5XZ2hEESVqNmY2re9JcnKK+k5JN
X153KQVMMxY4AEn2c3eNz9WisERBf3Kqa3B3xsChjSNyc1H7wLa/A/bckFl3r1bN
lPH+cN/zwZhJL/ynRE+DMXipHNdqYbg4ro3RiNZbLICK/b0z0UJxJF+/mYE8jzFU
x+kt3FqtL0HxTUgLklIwhhg13Kr5uRsoi+k60q12f91B5RiFBvhdO4QzxOQM1wxD
4vAwiAh5KPZsPqOor+Xf7Q1kZSmPvhkKPlClH5qO42D+l8Sl9bZy3Wxp456Zjh4L
EdZj+gf1MzHFYYqw46WTwnw3FxTprGmXVplmVyHgs7Ft/2o+6LduYju7kpHVhqSD
Dqu+XQj9Pkub/4ciObqE7iftafx6ofbyO1DELqWPX1C2Yx1TTZMRNRGIEOJ4Lwd3
YTKHS1DLAjbCAZluREgEuuCOVF28ZuSYSaEBx7GE4gz8vhelmqFAOEpMs+8f7Z+c
XnzzmImT7sw5eTyXj+6kVWZCzjB4ZMZwP+q8jABK3uZhX+NFdP15r4oU5j3c+UkT
XvMZMRfkcH20ks6xnMbL4Eu54SGvFI/L/x0nsG4isGIooQkFlg1K6v8MEtkgoVt/
OXt22cpYyzlvVvZSF9exd7UkDmwuX1S35Ix+pIjHCbI/fokmYll2ywT/kBWVlawh
`protect END_PROTECTED
