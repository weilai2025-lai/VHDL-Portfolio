`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5o1qxRM6MZvfYpK0Hy/0AFWVtoxYIYOmC99NPRte7z+xzS914oaDdfmRzowOXS8
7gCdbm5UVNgZN2UqyITOk3T1hzXTkM+vuvEeQcTDKFRIZutE83SulkBydv5fqMX8
hDZJLg0PLEKM2wsi6+gIrFmy5zYcq8FOblFm2OwiWwr1V4EfeDzq66sMh+p9ocWy
QFbWP2JEHMllQTp/hqV2mctbKJKMWKoSJM5HNptlqxqQSrfBlH/h44t2bHPD0WWN
Svfa/dz4A0kXWudkRBm9pb00MqJ+53YDYc/Nxl4c21/m43Tg1d/zKMi/PaJRTKD0
dfqc5wOZTC5oRv9BxGbOA9HosfmkDZKNr1B+huefUB2vLfBnbbz1Fl3S/7fwUAFT
GR+OH0CFCk6NGA4QftE/3d6V9y3TrkwbxyC5x5eCSBV4cX7gZDzPRJHsT6Xp0wsu
Tq97oKb9cx2RNAwg6Bv9Lzj/ef+fbUHdjPu0bhvLxRvOc4uVJEvUi6AoYUdIkdOx
LKlzlnNjs8e10gculsNOqpklreqKgxigATGygKJxSMF1sjUaUzV1nWdQEibiZm99
Beg3c9FGJIB7Nkvc8j820ooOgdW/TUq7vl8i88rNgiO2A5V+jhO/imgcCnceGqYl
S/uKPZKdEiziv/J6Q4dFVt7w9TOMkOF+CIuBpxQqAWbYElDM2sicyNN8+Ly2XkzO
HbKFKmOVjKm5bEVckyKkU5vnOmwJ1eqL6+DA4UsyJdd7aTiVYGHYc7I3MKYOZUpS
S2/Mx+0mBfvuPYy8tqZbSSkm/ORzhNGLBZe0FM5g+Q6EeijZlJWaZA2Pw0vQbtL0
lqebPkQoo3tRh10oW9fLs9GcEW47teEpSsRdHhiKbIDiTtEMVwhgUlLTF10r/2c+
QmF25Ksqx5I3NxS9pz+J48fv9sdfu1mjPh9wBB8n+nU=
`protect END_PROTECTED
