`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2y7Y+xBUvijXTc/VDndxfLvnsQ4QTJrO1a122CriapsDBeoh77nIecvhvsGXi+xC
duV9ptm+nWe/jV28mR25P2B/wmY0q2HaJa3A3jak+4hG+VxQav1O5snxzlBHSdKY
2yp7A5XUZS/kPSnH4gieOvPmDkpAX1moMVzhzIkz3LzQEqosWqb10Ih+O3ZzXBXN
y/KTVJHUY8jwijJ9iU7L2aDzJIifV3ywBLvge3n4J8tGRn0xqKDbc1XsAjmFnyIT
BInol1szQPeyDYeqTDgUSParK5/8SKlSEdBaJOJR47EvDQeBZBO2+yo4k+0/u8eG
kTeTosyLt6g8TdP5sU64sM9MirvvqThIMlh1iDR0aA8OcEB1jevqTv82YPxGKrig
0tA7LVrWp1Vf+iST4sf0MwDLIhilJKwyOykaihDQqFjLw5SKmtihN8bTk/w5OXZn
4d3jiWntD2xPXY5R6gTI8daYzpQM8pFO9ec/HrqVVWi8fuYey0fZ4lbRe3v1WUs8
0k9+aeWjJhdx8JwgA2D46A==
`protect END_PROTECTED
