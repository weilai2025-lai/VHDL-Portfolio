`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c5hwKyIY6RtTl9YjKHOOF6cMgi6Lk3X5wH6aPjrA7vdaTjELSg+BfZqPa/9FpaFj
+AhOvLvKNpPRyl1pbi72gr4TtrLzBEGm8B1UwSmI/5BzQDlbxMx6tCaPt/9FKWh9
CElEZtj0sToMCUMkVA3Yblp5K5PTiZ0mNUSDlH3bWW+JOKXqFgPTFFVa239oTxzV
KxQDW9zTStDjia9TbDdtYPtzlxpJtAvTX3sldTVPdxe3EWgvyF6rrL8kDpWZTgmA
G2ATPqYfJva/7d7BmdjeqKty31HGnq1XrYHztm6t6OmyLodKWvr3ASeotLsN7Mrf
P4M3/XoFrQb8yNTf+aJgsNb3pIbbZiTwcFXEXB9N0pT0q49znKnmxEoVtwnxg4yb
RGYok4ZMhFGIVfZvaVIX0Er3MwIOODeSvDswZH8bilM9n1SJyGgDAZziMU4YSdVd
Rzr+5PPzh93eB9NSgEWZ8LxChAXujZJSS02A+NkJ9C5Z/KNwkbbsnmyyIVx2ze8O
N3+nDJIFCE6uiUX8w8Bt9f2Fn7V8YeXy/UI0/zfOmeuW9XkJ0loYEenJfrV5w0kb
HId7r7HVBMjWcQ9lOuV66aKVP1qde0zZHhzSslgURfpwPpwSAdEZfnoF3N01bh/9
dpwlSjhueVT3sE+S1noel7GIIHwiX1A1oowxA4/awXDLSgw5HrUcuEX8qaQb0wlO
ZSnXHngYaSt3yxIUiJR+G/wdzhYfp1GVSYYFfR2LA/pxPApSp/U2g+b8fFzm+cwg
Ck7woTZ+2AsURNc09uZpG//UxcN7OXgBztP1G3rijGi5li+DRH7DmCDQs2Xkm94N
NvfvCL1NDxsyU8ejkTpCBIHnlsLkPxaRqH6V12B+4FMyV206rjiAVZ1YtUtvtcrx
SFW4DhaznG5bOfbV+cdtxckBBwfwwEpuDW5RKSravK2NMs8wiREoQcp7rlLsUlZA
GEBKi4v1rLiq7VDLlaM9CbaIFrIJjCqS1sKBbLQGmcFxndZBBaNvRsPSJ7F24Zb/
DJgiI9BVQIhoAkjFK5nBEOTQJA3Ebe638Merx2Fudq6pjhyeEpg1Igm/2oz0llqt
AUj79pL8xycD/MfaiQTfXMeqnXa47Ha5FHr0v02p6MmKvlPg812bLlKrMOlaHuQh
+zoWJLW5hSx3teD84Gfg1N/SkUrrd78PKLdsyDyb+GiwcQBZI6WiRR8eBHXHGYT3
OqGRMcC3pGRTwUFdsOZ249OKRw9P+ESe3z8CRTk4RJGvWZWoD5V20/HoGpVyyphK
B4UjSmiMRtfMytoHhR/jRY3eFChmzIe/QCq1mgza/4Yrr3Fc72SR8JrNOxKNPJh8
oloAvpoARH+D0fRa9I8wtabmtEQryPYWrV66mIcBnsM9rqNZ29ftx7RTjGAD/iqQ
z7evO8hn9ipIY17BCuR1t1izDOfyo8Tf39XbI1rij5qRD0O4tKY4ZzxiGiiNmxOx
hCQav8HG0uUIBNTFXqKCn95htPX7GqjBvRg4mSUeunH/oBrJPRw+SeZPDSCnphvl
9t3qJMVFdHyK9sIBDqcUY0VOl7kS5cfQsjjh6s4+LQ9y4ZxHtIbhYu84kCj8wRUX
Zw3WANdWcY0tGgqB7gPXS136ys7Cva1nVWngJR9NBWibmfvki0fDL83hu3W2V9fs
Q/+yFM12nPzOcIDZ9hTlfsjPa8Knbp7DIl9bWtKYcuC2XWuuJDOiw8ezZ1KAVX5H
JNSJb4XNWvdnR4vD5a+CGGSb0+vF7ZVgVclTs0A7UTPESdlnQtwWRcvCUjF1y/dv
xFy0qeirvAGqripT5yD9dPj1U942xyrL9B/5+EPEGS7bqV3cZwI/yRuk9iRPKy4F
FDQvplG+irhd6jpJPxUZ/ZkTveMowV1zBZmKOtRRbg0P24ywZwbPH+3qaPYSSPH8
kNl+FUZ4iRna0CzwkicHBykBtjOtFKVLEPeDdy3uD3DKYcYUYn+TiQABM8J0E2HF
AkS83h+AmLiY6IptXJDkkF095Q5ES96fPCigVtoV5NgoYEBa0++6Ry80UdSjT0WZ
mAauBX+xbIG2UZndhYC6IVVo4Cjk+rfeaspgQVCjaHaC44NLSMKQdsHGGrhYb1i2
4l+FFz0+mTMePgyoz8VU75ohJa+GsXAMxMBi6LxINAUmj78HL1thTLYlcn6q2HJa
v8hwWdrBKXfC01Weijv1AA6J8Qczve7JBEmBvLgOLq+2NaISrVDCu/Dx62c9VfPP
jEJpeN6LrI/iQMnIZAESFMssFjqyxtpI6CCIwl4pkDuB9OFhorHZrX5d184flBpC
fQ63nyosGO7YaPDKyNl4HEOUzVBT9hPIbdTvzjJpbErQfiFaNNmDcgnPpHiVJ8Sg
eBiyuNfiLoCnK8rY9XDStMAMFwiaKlQ2Z/oA7TYEQE4vtWSK6Cl+aJIRkxoFBBBt
b/MxqXv0Yncp7L1C9myb1I3fc5SQTQMbcBCvgGDtHt/IE0RYze+RKgT0Su9WhpuF
+WV2EHYvjBm8EGdNt64hNIvX2QSmdqVMC/8WfAu3KXVeyJSbUdAW5yAHJYi4lADm
VJ46TuWwGiSd8ONnf68xfyXcCcaK8KY5HQL5r9heUVeHW7ym2mhX7xVbitjb6s2r
Ov4/ljl+VQKpRWr3nNm99qEDxjSP7BJ7jx+qi0rVwVhnt5mN0XOrThQjmb6vVKjB
z/fRwDYX+kyw2jNLvQUQw6hW3XcBGSj9FUkJW7J6wxNK+Bu8TvbGg74OTnS6ycqI
CuBRSV6ctpEn566+Pmh/mRYQZIBEykT08xuE7haCBQmjKbIyLCbjB8jaB+pc1zuz
kxo6GQTVhWEoyJbHmUPqRm43jtfLiHvzPBp6O1OgT8xFToQzSJBmCJGwXgChalya
gT2T3B628ISIobe+X3u+oE3pX/7PI5rTqBtmDu1Sfk8oRItj46Y00L/2qIbxjHPf
6Ra722uI3ZfF/WVhu46UYa7wy4eY9el1frElLr1D2IyDWpfKleIY9DPdphgaiMzX
PfCjDIqu88C62wunKHw3sxGQROFrBNAVYfUhFLatLRD5D1BBKUlVotu8E0IbUPAU
f/hvftwT76qx7DwI7X7mOB54D1f2bIdddUnBvhsqjiQhYrrXIs5uQx/NEkQIaaFh
PZcisqixpxe5mqhgT0cxE2cnhh+VYnhXa31Zfra8MeRbFmyCBiokpy7L8Dx714ya
kqxSO+WPTw37yeIhQHKST9I6HU9iv7TM1eNtlus2eWw9AgHFg3HyLxNkRTmZeE1f
WxeU54nW0NGlkKd0i7zQgzx3bR9VKC4kJl4t5uCWPN3Ce1LCAI+jKdXYDabovOKO
uPCxRArg7dTs5flGW5hlvols6OO0tUklGKTSjkDaDr0HdheOQhImbuII6+n3Zraa
IxmfIZ4upoFeVSX1UnXGCIQujtJ/OxUZe2woQo5vkQfRibhGqRN2Ym779Sag0Wa2
TuYbM90xS9ylwA35RWyWIaDt0Fo3qzb5dWQBW/N6hDWS/zx9ULsT8Dyu41SSkb46
wtYIRBEKTPx6vSLeowo8EtGaDAlxDjVg6ntc3heMI5eJ+wxK4FO7FRzPXBg5xbvj
GnxdwAKEgT+Dz7LdhgJoTujyhkGvX0WqXBt8ORHOPwxS03rv7dUBVPSg9dNRLWzn
Pl6yUMQsrJ8ZNHtCaxHxu1dVRsUQzcb4r/NiHR1fZVIMAfkoo7KFsJzccmfhK9eZ
btgSdYr4UyPvx6W3uwtDIrPYFW4oCpFaNvMTDFRqX1ZGEpuqpSt0lGSjLIGfZ1Dx
rxnLCo3TKfDxFeCwRdxmskaMiIo1KordgodosIfDf6+vV/taHyEXe1Q3LSicUH7h
Ea0naSjuuiDEpKHcvkYV4TNvbIub7em6DUXtmhKbbSBjK+P2eXqIpeDrvDoakmTL
WB3eUSCkkNHnvwmsFpTJ2ILY7x5wJE1F/154kv8lJm1tzxwU7OsREubgBR3dxFne
qmCsscOUuVS0z4pxN+1XXvOhEb0NjRDMK7NnCCT4g9zjFjsZkj0rYnXUz+G0y5KH
N/9nf4u1ZYT8SWMZDQFYO38fgjNwG8Vo+skqkxrz5e11imt+9n1AuT5ImGpmrg7M
XRa/fhS3S7yW4ae8MKXqIHDEdq8/cf6ccoVXfFF1VQNwmYRqL+VZXqQU2xJQqxkO
xngcUZQKTvFMQMxEYCGZuwHnhmIrJqncOrBUSJirGyPyd6N6gqMDCbOjEsQTUAg7
ddyud3sK9hRzVBWQuzNOOLXUJ8QSdkK5XAlaEj9e6jYJPbp8ds8XffMcgpwzhsLd
ieqGBGNs+vS2JKhwNkD/N5NbopJ+1l39+kIx0l6mDXAQBvNU37wl+phTFd3o580E
rkY8ex8jdO47pBSNF4fyy1jWqrYWrHTTGOH91eVJim2WDXKwZ9sC2TK2oo9Kb9MK
mJoXAOYPD/MB8KBEx54kcNHni4N1Km6q5ebU5wuaC/ZDet7Y/6RMV+ROF6U51OvQ
PEGxSwDww6fXdu4ZouNDFY/I3HVcclVqbr05IcZGn75jS48YSgbWoi1ph0EWCQoI
yR2CdE5vMUehHGGmHpMCuWWXLQwuthEdVXsM3EGN5H1xaW5Tl/UFEbn/zqoap5sf
MB0STbrQVbQ9+JVUHd9wCig5nrbmZP/ZWPkCK6qJMPgaQxxTuk1sa90XJNjKANI0
zFsGShmihUMdT6LVB/bg2yRu3ZoYEYzNGjYWNP08XKQLtNOgEYYmUbqYwDSEtzvr
p/HKCKcjIfilX/HGxJDtietcRFeph3jW1zkLLzQHkQt8jMQZNgAEf0xf524fYSfn
YQB8N/faL2018qwn5Ty710iJjBqJz//GojRWhOXKih39Qfhr1fja1OaW5vVuxAP7
xQyG5FET6/EdVeioKkVBdfC5JegPy1sCDVVlr/iLx717ywIKAWiMHfImhUVICtF8
Cn3uaQ+z/gFgJ8F8JPPYW2rqKbBzUJphytRTunock82bZBpKPko8fcx45lauuvXQ
PXKcWo9KkCCaSZefpebsFaMGd0mMbmEEZFwynXO0r/RW4yGf/c8uC50Yj+tmfMHb
6SbyC6No1d+b+Yf5JuZl/GfBhmXu8opraV9wESp7W8r6zlCCop9yDSggDqsN6G7r
FM0Yd1oJh1xyB4wXWGxYIrm3Q9nVf2vD2A/AsHt7yirmdpoHQ+qAeYHXfLeBTGaj
0LI6yLEaH79dzsMB1mlEDkmivcZ4ln9lmqs1t8cDP4hg4Fr+nA7WLhPCp8+rLK1w
L7+VlBbwB9RBylLQpRz1gSKoL3py/nFkSR6ecOrk04P39+q8eWutwSXdzxHb1sQC
ovn1qlZQXlNWI7V3XUuPisR0bMPRuCV+oGXEoaYS+WgvAnU5MuVJ5WNPdlz9j18h
yfx10mN5tDuVeUW+3l3TWupfKBi/1QLEKIRTL4F0kW2l9l5gozWW8cCTDheB59NL
+tKmw8aKJKnNKn8AiwoX2WSREnprMNW4kLe3BX/TnJTwDzC8YCU/YbnohQjud3kA
wGUAVJGvAX217+LXmtusu8+HNhouNRTeZ3MaSge2lMswMfLk3niY7+NsFsFWaI3v
XGi/sGBFDcyCAn1EplfmoGGxK+RZ7Ql+CFuJ/9GEVy3dLKChoOBu0Hag860CDRq3
MuLc4EzvNEVNQZLH4oS/veFVKXbC4uwnbVu5yka5OKMDGRJqm5glJ65V1nmRUtmh
Cm3IHa2ppAYec6+Bk61VBKcqewTQbZ+A8DHzPuinlhXDV+fRiffsdFnUOV5tgyLA
wC7G94XIRDfANh4B9ur+MsYcP5Qvll5hgnEFWDnCFT6MfK85Oz0rMTZhNYeMurhW
yQ04hvm98ZvC00RTXLdqqU81NzBLU2POLIT4K2UQL9WlpVnyz3YRZDo8XBHiyr6O
DU/D5urparbDMxO7oo2Kq3qkcR6pIaQRV24LWBgCGG6Y3KmP7y32tC4CcmKChpGO
KubGpfsF2E72RwfKEBs0rXM+06EvsgXCzteyFKMDUSXj3rqi5T8ICGcWqJYHbLJs
LowPbYu3T+oqd/YbBX+CXAw2b5/XDRNoHKsVilz1s50YY18z9nzX1ZvnEB5lGmi9
tyDvd5ra5HWrmfdufWYomT8yzNxnk2bLqiYmioKUJNxjgCHF3tWim9MTRb5REONg
T9B+s5zMxm7il/uj5xlnqcHTix7f//DXCq6UbeHgZHAFWcxjuasevBma5uU2/gf8
qAiBFN2WTzha/4RTcB7mg2LkdMcMCXMcSIyUMi1bDzkJ4qOy7Oj06lqOGJ3D5zpO
oGG2hEG8JxGE/xy3chCck4aa9ZnLIuodX+J2jEkqDKuCNcJ87P+JgDjjRQ+RjD1C
LQP7JasSUUvqM/JaVAC3LDdit9m2o5uM4h0efVK+ouII2qtdI+LWJj7oQBJcUVoh
9nDea5sX/HTjSW6/AoMCYWlox32tXbfvMfbQmOlH9b9O5qvmAJXDWT+1w6Ln0eVI
eKNTrYP+cpQTYetDpG6LINqt6Y8tWKpeKqZZBOEd7VawTUKaSS7Iz4GL5YZPFy9R
YczSQIM+t9xR9//9HRC3X7OpK8cQz0RC22hJ7x5J8JFy6wY4OTOduAjAR6myzcXw
R6Wgzb8U4gpzome7jM+hCZcn+jS5MQYMJMP8lS35T5jBvhVQnsnZgbqb5+84pDyO
0laOWGPhMq/42vvrn9SoVfIKWnqleehrUwaI1zVKSXZtyGcgUsHz8BVM8egPVICM
8KMhWATeIvfQ7l0Tuo6UywzNWFvKhDdkcTlf2mpAMzncXFqMjpABfygY8bgmMPKO
Ln1YDr8uKP+BISNPydrgYeNTA5GtdbNtf/InifLc9LGPX8unklVXb3Kl8HLpxgdK
+U8ciMEe1AiKcygZ7zp32EmbLs+sDduS1rXllFnLUwy3DQpRKFZLmCwMUwZ2scHE
m7Q7Ire/RLd18Vl7t8dzUG+D0TC7RZrVl5ktpY+nYfr3n/R/UnpWk021F19qpxSj
9OqSCgPSO4Mx9xLivkq9RaIDtAqBIOiEBlmWVa9U7x+/Gww4fLZBEPSbhS6qUksf
+Dg3mevrW9n8qAWk+mNNHqdxSQJ1EdLNRxhaGTVGyMQlP4bCRj8NsPSgxX8wsvc+
fEZSbiBmOmKIh8wj/a062PYrLZgsot8G1dys07JuXm445mqbR4/uujKZRZEGdjgn
wMswSS5+6J3WtRVIIJrZh19i+kP8Thg10TcCtGtMHkwn/GyaAsVy/+yv8vW2kul1
K1YoEbbmA9tHxmuUWXsYwCcYezShX5rzN3peoMyVU9odw08Y61lnlWbFFm777js0
PCF6rD5eb64hmWml4SzFJZw2VVcpt/dhfyn/8I+bkMZYN+yG/DQT9qLkjwW8/1am
XgAtUHq+5qQXbcHprErvEhA1416P9LL/iEJiJ5O+Ze9dJHf3WVSaWqVHUlhltTGs
MW/Qsdk/OTZgHzF0GnHYPFk8V/uxLMs95n+ieC10IRd1/PsnQEXDXx/VJc7gphcV
vg4VJVo7UwuK2YxLEifZ29QZb9KiZteYo29YgFyQGJiFYJYYrpYVKkTZNjV3G/pM
IjIn7Eu14EOhTZ9F+4XHa4bAKfWqPM6zm9MIU4PzE58f1L1DjQBRtDzJgjxFLSv0
bt3fXG/Dmy+wJkMuEgL4qxFEiuWY1mGOKpU+W/yvfNbpzcRovUbfbRYVK/zKwzmx
KRBGMrv/GAWbQhEPBiLaHjN2+YDpFoocL3BcDoVGKkYtw0WeI/trnXtOEefjdmbF
S+D9hi3PeiJgp6IlbeQIqVyfjPg0SzCKbFJiZNdt6lGYMm15/olnu+gC9tQTxVqE
FjlrS0Lxw1XaJ4nzVjSQ00hJeNIYjCEg2m0VVBgU8jS2G3csFJgUtI8oBmS7YzkY
aFmvnJGI1K/tf0PjMEKT7xSQ3NHjeQ1vA1wl9WDYKL41UPnkJGc1bOUY+gbDSk0y
QDxWFxa0kvXNJf7DcRzU4w1x54nt++NMPmi01+XDn8rU/Tgj7lI4pQmt2aAXYb2p
281mJ9SDywq+GrIHRAZgaEa1XLIZrL+hk0TUQA3FOlGXTKYNLHzT8otG5+olfrvD
4CEoDWbVHxhwD30csvW1oO0PGFFy5dePNLs7qweeBbTq4VxMNQ0e8rGiYyvdH1/d
CkfkQqitxUbRCHxgrvldWNQSV6xNilHr8eOQLxGKigpxu5KQsN2/+BSKDcHFFG5K
FdFQ7YdCZs6KuKD9M1ID6SpI9u3xrUAcloi1FUMGI6mmyDJuyGHZrJz/+141eV6H
ipcSIdvR5bLWUJSnwn7owbw8UToXKpsLV6noFjy4T8+cJI09+gZmrVwp37TvEr3d
+YMnJfoAPd9jDFB2Eixl4XlzmoGmq0JlInSkwftZrGMrx9QvzQttN43tgERDn9sW
DPWLG4Q/s3yOsocPvg9QmY2FbIKJDHTVfNivk0xyRbCOOvs0ShUq6h2GkZ3iizea
lD39npwa4CE/l4oAbxmQX/0mhq7A/ejbjpuf+yl518LCpZI11C4dWAlifZW/+5c+
dT3nRZkfGXuk2tgH0vcl2ca5RvNDCdiAoWG7I2esfB6n/Ze9NiJlzL0MMFs7KK5E
gN+TTigoSHxuQtGa+pZ/XbI+aBg9rglBFNDfc1JMo54Ht2KK0bGIoq8XYljFKq6+
5B7shQkXBxS+JTF9eyl5PiTI0EfV6IX2TIgJJvcokUiNNmJ7EIeAE/tCwTqqmMTl
c2d2zblHXgJuio+Gs281Z5nGt4Xb8lW5DpmU2iGdzVbpxgm1eVnn8yG4I5oWxvfb
Z+qFXFx4iq7/6hWdzkfeV5lkLh+7Wr2DFU01QCrjsAZEY59+/N50pJ4JAMBs4I2g
XmouLsaYiBDyV87qfXSKQEdM7uL28nNf7rSgYNh8JzbHol5IT0Aptc/484g2Vk5o
ljMqoVXq26mBpXM0Z7iTuDEfc/gL6Kqq9aHn4SK+ZAaQtckl2WQEdSOC9IgY6w2f
H4ZZsCnJZAhvrh+AyxBPxbq3ijfI0nhMKe0gZfv8tgCV02pJ18iU9IolpwWQjU8J
HEehLXZTMj9Z5vepXXNrEUCFSus4Haq6ZZJXkY6JtC1qK//0AQWJJhddv4e+ft0p
fKiC8a1FrNDG/0TflXSMc3JFXMkPreGm7dw8OwqSvlUkRH2GXkWapMLNAbfKW0BT
r8A3kfRMOIWu68oazmBY3Kt09NFAAwkRAzBMD6vvUT7C5HknirNqNn/gy2RWngiT
tL5vjSgS0RdhjqSfZDf6hytSJb79tr8sV7jIBU36yro8cR4s7T9U8uJIBEB9juRe
BOLZ8mCanAj+fD1l4s+0uOR11p/8M4N/4WoevxwEbLYd0L6UMtPA6hCKnfHxpdoO
25c70OLWRuZiLfawMQGE5jjukdESfqdK6uK1LctaSOeuamAb5DlAUYR5ZPbMktlc
fC+y4jsinupilvlHstppKMlE/UXSxpRhkO+NkEevmsonHChfdAArrAj3mHbA8VnV
l1XLBbXZx58lpZo9EURoK5r5DRkW7w1w7oVSq69sVoxM+cd66txrmBxrAfjL7R+k
GfN22VMwXXqd6LbskWrewK1xD/fm3zs1dYBznvvwY4p17ylPNKlhSPPokMcpQ7IN
SHm0TlLpV80yDaQSg37f+QYCuPcnSXwjd5oMvdkeAU8QJwgF5NL8nmBG4r5nq8uy
F/AuIleKfvGC9TNw9+VlpQe6ZXKJqnwK7b+9mmBxY0TpV2njYsZZvikjjnRDsG7v
BvYemkfnQ2P5dK6QK4QNm20fOhnXQQEULQCokMNh7mKAUE+fkCW8EDSDf5afELhI
pywjqdRKWUvv/g75KNd43frZhAO7BYsZgt6r8G9CSOKx0BE4SrrAJqcmY6EWjiNr
2kh6oUXuyb0cEDMxcmy/2DPRIIXdk5jYBkZMbH4hYAd8snRpdnL53kVwANWuAoJ9
ndnyzmcGjrAiOYFJUh/MF3AS6NAxSWz4CtsxxLWrRs04rBu5cjP6W3AmGRiE4wJz
XLKL1pmGr3IUoHzsiRnQVugcO7A0rJYqLrObm0rPTA1X1YTXTftiWpyVp7SlwJOw
2qpmc+fCDU2y3IKMhiP2kTvOITBNG/WNduRU281t0U8bH/uFeJiwh4/S4EmWhxwk
EdhSRmYYIJLSjIwcyD32MJe14lJ6zThBhBeEe45BvvgMJixcDOa1X8DywSHCYwNu
hGip45dEci+/cz2ty2vTBm2d/r3B51I89RWX/4qXQ1q3PHy2JBBh0yOd0vSAUSF0
cyx2OHmOvjtEJh11MlWtlDhEjrF8sNGrzP2aaS6QzWveFMUTnsVEobXnULtNuE1Y
mXcXhOdMwThMZHYBVJmIU7O9yLG/JgtkBHq9xbrKUYj6V8Z3TGN3hyGjmyfxaK/P
LMg2lvqF5IBpmU5F41AOmjJvRjCRNBf2vWyy/e4HFHj08+pX0uqVRNiuro2QUe8T
VXtcDZw7coCOfKTErhj/2MY0Xe6sMc3+VsAj6Pnv9v9J6XOXRD5SqpPxP2pJ8MkK
b7hgB0age/8BOi884mXjBBM6dLitNYr4oROPRG9pBytjTAeUG2nLGK2zd9YF8lY5
f980vjzqUZ8VhRrwcBaNcmvRalRACO3z+9tD7jG7Z56LGfjW90mmlDYIAOv8tv+Z
JbdZR2GFQdnqm7fL/D3GqwvGhXqGyv7RypRLeZCd2CdTqM2oofh3AZOvcppI6pCV
AcRhbiOz+2akOghdKFXbAnI3oLZZoG3bwwSBBGCUVW71Gychj/3Y1ruSEMVZmTbN
zuvxEjErRNgLjpPIX4m80TxkKDGUnAerFYTGXn8KeF8ZA6tVsAggsOYk5QOV7ap8
wj7SOb+2Zpq7jjHWXxvapG5KMzIrb4bMwQurxgOLDsMnPPHohTk6DP7qhRN+2wbU
NOaUKJveFBBMq6qxH+jablbZOWhUAe/0GIbWq4ZtxsQPzo75iOW5A/0LNzBbLUxn
KM5IQfQPG708NPKz/DHidzvWZLpPMC0M9evjeXetX/gH+LxbHfsLI7/3A78m7zD8
ugTsbI4+AGWnAIYbRFpqjPkGlODXZTZYclPnsykdRlKtwHJHHlCn/SG6xvRC0SS6
2BCW3RDZcecNOANOMskfaCLC10KhOzrjZGTelyx3mpdaF6Q5bCsmcfO9dEQCXd2B
QME2BfbXRFp5nhUis77N0wwyNVcI1jpjDrh6cQkAGwh+0ymT8JmYqVO1QBU/EO4a
FGWS781NRUQuqQ0EMwdkMOBVIVrVZEO4d9rKIy1eCGJBWhTaIghBiq7H3jO5ET5n
BBopr5CdbIwOp+mtXiXZ/i53itWFthwYw5NJ1wo2gnpoWf84ZhzNXZucAhtjKv/P
YUiO1uv+sF47RZOVv1tZVo8wQeu1BLq3Pzw48ETMt0piyF+kMhUZcZR/Zdzu8eh9
8gPemZ6tPu5Xs28DCY0Rtpu4PjflKUca/BQfCzIwwHPv2fahfQLqVQbbnpXnlz4l
Yx285ULvEBxjl2DrdDMVwfMAliBNcuU/up16zC+VG6ALMezSE2OZ2O8lG4h4Tjd3
mVzu7BdtILq23/ONyJRbjNbHRV3vt7NUA3zOMwBIAF4MKEmdw+q1298+fG4I66AN
l1U19nZbkRx3NFIHIfwaWEHHVP3RfaT0P6EzXQuFFrOrMCkEhrWKUo7+LygeyHHx
xuV8R7EtUVA8L8Et4wKcT6YxQywxwO1KUK/ufvZktAWjRCSJSogq6yJZTNM+Hvrf
jJ/cMq2jeAP1UvCwNwC3nYqp+Cxmezbxc7/0OQ4ChI+s6sM4X2kqjNS219THlLHo
g4e2upKdBAWvbHwtN1emh4iU6PWVRsbo8TTQcTSujm2jrc5pp3XvUaqlQ53WaevL
A+r/yBxnj96Ebmgy2E8B00kX7RELW7amrqHy/gWzSbMxGzuR/VYIK71lbEa9EHxn
p+e8RPptJQ/va8QQorZAQ3OibnhnrtR5Z0RLtgs2bQgTyp7T+ekHhUSaAv2yKIu3
EeWgnOVXYEo3h9m2dG6ytQnCrfPOIQ/epj5aiMqvxXwz3+H9NzMH6a6PSq4sAszG
phyB+N+2OnCQMWBETLBLJojezbSlUZrp5WaJu2JAetB3j8v642uNty30+4K9x+tl
sHoX3N+FpVf+2ICVB7WmuuDq7EJUn+U1T95E49qREZG/JUx60nS5JjoFYozi0lV4
EgqHHBttHgtVOHW9/9NBY7uvYrlqNXk9JHkj9qqFH6HAev+MuCJ22zy2s7O3fQGV
kaT+zpYb3qEwKZGOsMUYsy3oYLrtY5dOOTZpiLCf8s23bPEMbJXWgdDtz3y1d4pe
7NLTiUsbYB9b2UxkcuXF8/cIcAoKsxCjycrI28RbYuzUKwGo5M7fou6LX/qVNgCH
9wXpL+xiMh+VHbh0zZDLn3uxE7dTAFgYLT/R8ZUkzmmoMVj/WOg6VMg7OB3uzhQT
3NKA/58S6HdV4p5qK97DSsg8uRosX6NrsXoDcBbFBPwNq3iDqkOnzAu76crmwVQz
Ydzr27pHwxkbrFE2D3Jvz11KQQVDbVhJvQ8Q3t30ufmx8cEb0KUP9N9QmUf/gHHR
IXoJJda63yuykmjg8X7DmDQcs1llqc5GokE4AruCYMM8AvT5/WTPyJtPUG0zpJbS
iZqEiH0c9wsNvDZ2hYWA0twRBL69qNUHbI9iacw/keme4HcLmSoinvsvfLwxS0JS
WnDrU+0buDuuVtdOoVCNsqkpxrjhHqZvKRGytckO1xuNOyKGT2XPjRlydMzVzk8l
sQixFSpG0V0iDqdLbCqoPyaMMKOEOqnMNifjuItzU7VFD7cZLVxFUv2+apK6d6eV
1Vyjd5rm6uRMzkFChR6UrtCkimRMniQ4Ux3DMHOkL/ANxVjrD9VD0CQVQl3Sveq9
kvGsxGDTKxQKEY2W7ptZGDUvKrH0/ZPdvB2UU4PUc6ixiiGOplZz92RhgMciQi0F
7HtRMUYBOuI9S/36udYdFk3ISKiUJYG5rZ3w2qzYIjtG4NPyt9wfoibSujBg0CG+
NJg6KWIwmC9Qbiwx/sM2qzMk6IgHp2vef5LV7vto4JdcAfbjobviv+xBsF+Yq5A/
SovnYlv4cpslkZxYuDikRtHFB6PE6DFIPaJ8uo82jcHO6sAX+gbOuX+zZfcRReZy
Puqkt050KDjshgJzAKlu1GGl9bGubtxMDVOPnAor2SsmpmdydMoknxOLNz6Bs9gh
kC4ibTxsbucOug0erJIOA5E/q8VfXFCKvRY0L6rzZAPsMODtv90Yb35jOmUluEZm
4t0BCJhYZodyWe+bFAwOmInWB+uFwPY2Tvk2yVAhmTrl9yRJXX5opbh4kjJOGhcT
y4JwbSi/uND/hKQMDrLwKclSAQYi3cVGltJVpmrMXedgO10Te0e/Hft3fYw0wI6Y
npbwmz2cYE7asiMrz5kotl1cyalEBlOT8cZpzHPn1C+nA+yEuIj1Ydg9Eczh33xn
uv3Hhfv52VvwWdWzcITPNUIqUq/6VwVH//o7DkCJesOFMXJTOCkoT4ieXSswf7HD
qXsD7/ueYk6631SV9amBMTTVZ6EbT5LWQsoqYUDzCXx/zn+NmCy+zgHsbDe+AmSa
Salvq3Mu8EfssqDrsocnbNLrJDLAbJVkEbkibXBzlsFJEIgoYbA4ek12f+be8rN3
1B6G4S9p1Uj+9gyekx6UZBSdddfUVrRP2DLXDiErguqpghxBzAMAP1CiTzQmuXcz
dvOhctSsUmbiNz9El4AOhWGquy+hwFwonGIP2YBbaRtdSMpak1axJu1pOuu9EIxS
yC32JhK9XEU3nG0P7/K1iMyhaQIGjcFm9NmjVxLr+gbtdPWSQJjREbrwfp3WYICi
IOAefaMZLJB8+vwWbx/Nixzla5GrUtugHFzuj26uNsJ8aFCDPeRzi4V+Km3qbdTQ
ZZCPAbnLv2SHjRx/yNY/vs3MKY//YFTAoU58Sl0NvA+7cx33AfVEYUsB2+fYrpCC
n3LITTbM1+WnSHvBFYPhdzekDiAS9GsGzCOXy1RsYYDRg8/Op5UnQtm3l9HWXl6v
xeqhH3I8/67enj0shOwDYtxxz+yLhysr2QLCTTOv+MBp+XMZouRGTL+Og3rxfpUJ
Mfb4AJOahjIwyoHCzx4zzyMhMTUzf7V+Lw9AweRL/EeMDapnAnQVOk4RXBZFVYF5
+PMiK+GNNR8yhiYk25txfcLaRdNYecFwFHktE3nj9QsQO2kX7KwgXZXKuAN9xxOr
+5zic5YZtUCSlXEj2ew54wOSGdkH8+xGG4yLbFSATdUgnqIhTFp/PP+odDaaqO92
NoxmPx7gDYr6z44Xb51Kw+jkouk3TZS4u89uQWvH2oj8z52XR7ntV+e0BDxJMkI0
qHQRWzmYVOOFfqGR9Apj6ztZRRViy/1K/keMaDOW3RXcZ6j/Tf3/Jrloa6ZYtbRt
Ep29ezFM9/k3yZ3G7SolT0TE//rZ8VT9HGlGAaDJOsqW99votEb9hwd4nYjQ/z/E
SR7c9l7x81ketoUdFP6YNUFrSyFmd00XSTlpXPEzNNLUhHqqQ0SSh0XOmL2FR/nX
H3vZPIPBnUr9zX5wh7/zifINlvd164jcGn+biEFQk2D514o9VTeMSKaO7xhe3X1V
G0tP9YqizHhE5/MhXXg0MzDS2dPKYL2DoRPhcTSWrNJDCQcHM2RgnUqMtDsPqLou
ZFJzWGnRAvzS+SeauUfJ+77Y2KnZLIguMLkQrec9xUf2I6fzdTBM1wIc+9WYtKM4
vXz/YjtIwcKg85/1vsQnpBqj2tnEt6lkkKsnzEWqWv+B1X+qsvKr2rdpUbdHVtUo
zb/QMCAcoPK/mKXKmN7KVInx2ifcnPOV8jGjF6h2rE+CWfKWbAiRPAKKl3O6EPzq
VbIo62j8pbmm+FjGGhcNltjfNccFGES0BVyJWKOVmaI53ZgjleKn68MClZHUp7PM
+jm7cl6D2gHknhEauBPi39ENkcxyORC9jJMNX8VPh5kffPP4gjbI6jhxTc/VM1fr
gTSj+EHhx4xB812vfWmIhTndbdDvYJq6kLAZsjrka/bcsZOBovaiPH1kEooxbJvO
YAiEBP/sht0m3n5bJHSLKHLh7OPalObcHI0+KFJIn3FcQyulWKlHsjNm0fKWyfIM
LGMIzfpJ8MF0Fr3ltrHCFGK+rzfDbvvtOVHhk4Xxuje43gCS006I96R82G9+JnJl
qH/3hk3u+xOZN21mcVYbYPgUQSQmFBAnDNNXp8dC0bFEM/x0eBLRkLE8Dm6q46v0
+HHjN9TmtdJh8+jb3uOgcpqd82dzNP/z6co2IxwQ6RxpgauzI71QlqwdXP5vxMa8
1ajzOJ5qD4ltRgPgE+d8hadpw3HYh83p96AO+UFQg7KlPXRE3MEyTA9q5DLOTLXD
3etaeqnPbhCxQ8AhDH4jMhNKTwr7ET13Y8FE2jbtUL2ytAogOp3BqGeL4lfPF3h+
J57o0pKq0m8r97vak/xeqA9uu/kgPLoZO4BSreL33gIdUS7MYzD20MfhEGJ+KLhB
MxsotPhG1bkFkb5H9hYYOQGlXxsc8EC7mT/Q281MYQ/gjXSFVMODYYZaBK1Lu++F
cqPHnlNsVo4eoRxFmzZEg59/ztKcxmIfbUj4/YrT1a4Y9TVUhHqOeW2eRif5m0sJ
8HmwDLVoY8J/5mRlIl7v6rMiusJEiHGQYkVQpT+xl3Zgy9aN0O3qsNTznizY3I5L
+Yx04ldiKOThHzroEdqLaClLBaV7Hnm34/Lp8jnfMRjZHOAFFnP/EFzUWUrT3I5n
upq6FNZsJxtB6PaZP7HExV8d6MmrLu1bnpZWZkUfaQRnDwhOJxosepLm2F/nGr5K
M2f+Vbk/aCecHPKC4jvn8xXy7vGs9+dIAIOc7KbT2Z8jIfHMCq3aDxfCwa8h0aY7
ZI7wgPDVsda95hNjcW3cWz+n34dFiWqFGWEsKmKsI5vwu9eTx1oNJihZx/gIaGkJ
Z5O1MTftKGLXigKajUF46qf4Zc/qeCtrm94DHJNiAphwp4iXvwY2rj+xs70+r3A+
S2xpPjnmMZeOZFUB8TfLAWakvE/bhq5+79BiDXSgwcBzsOZ7Ih85UcBlBIqWzC9J
VNfZejFCllnVkIlMI8B0uUDucae3+70WRoW1hs5A6sPCt8X2V34dytD/lnS39NtR
6rQmh5772vE8WP9+S5lPr8UlIWl6xFXl5XICDknl9ULNsMRfZH2kgknS33IB3emh
UMXbqxt8t1vmTR++ptPWFa1mA9Efr5Gv1jsW0m1p5LpQB9MTnVIpTjjBqjiLic9m
zu3ZaktXwGO+0NbgQwbjoP5W43/Pp9OFTI81tqz0druMf90lDBwuKIiPj4L3RuNd
0TfhLIEeR0jQmUBh4yy9IhfM9iL4f4c6K22DakRI+/q8ptKFMooV2zyboFX3Xz29
dnEHMYA1eqbp0G9OdIBm6wCZ/gAK0wGZ2awMH3WPzcDfRJaTUJvXRN1UyQnoeEsl
5XXqTNu8dP5L3a2GXx17IszQT2aiX6hUmwfIkmZwUtCZhZrITGnolXdVAEaWzhwD
GY0VbOCxpxJb/RK7PzNFdqQJwo7//iOeWY3ph1ewEtV8r1oFpjZg7dXc4BvhX78f
EgrJM1QX1He54Btz/i5qkKJ/zbvxOUM63euA+1sscEj2cDDK98gqXG9fR+8/r6kb
oE0XsYISr//HAEGaZtn1JSLhnb5TO/m69LuGAz2WpWu3St/h3w7btehOSobPE3i7
+AmR/rY7EYsgT6uPCEk/KqRkmWCamgJCO/4ydB83I6LbKdSy+G7IVePjRCI43wAY
0X+i//d6lIYhAWyOMTg41m+41dAffMTotjJrWSEvsB/NNBLX+sD2DcbT+5khqUZK
fnUoLecnkhuYDUDQ+XdkcTb0A+ncLr0Zk+1HX3XQ/Rm+kF82MAkTJffWFIxfUFMu
R2umEdNE/y8yP+gn9yUD4LzeApswl5Etft5F4LjibI5n8FF3CaDb/92VjNGwU0nv
0k/E1/NBHHcfDSrdmS+XAfVsOZJhP7Mf7ZfGvd8/KxTKtAG7k4IIqvsCYrrnKYG4
eyZvgVd5yKp4GlQMnbxU2n/eolQ+k9GVootcOZyi4bYXUD3mvjjfiWXHMBkIxI1a
aG0I6ayTg/0jqw0TwwtZPka7pGw9R4Qwcdft9XIdgmoT5kqbMH8chDfhaCOC0gQ7
GnmyAZPem1CgNIT0nQey7iCuNoQKnO6GpqZJ9csV3yt+/FJwX1IkcMXU9GHY1+th
a1FCkjHKh9w2qIVnFskqU9Si4QxvHJOT8fx++KDF7e7YVSEkPSl1zJqm7+O+JZM+
vrwhKuegg4adSs3DC+F5NcEWMMB2w5JvMy/A8ytOWaNO6lOx06Kpg16konkOEoO4
+t/mdXmeC9PPl72xXaPpF6SFSy8+NccNTpVUnWcA7O9Ioi1QlOlTFQMIu6ISOy9S
Sfu3SyBB6rfnmhZnl6Xb58TX36KDUp3fvL+4xOMUZ495n3K1cwXAcmu8lRBcUP8b
KIV2jUpnUoDt+69AGNHKX7No/DVeJ1TEQul7/G+sME4hFp9bCgwWWz80U5gtRzsc
/xpDw1doWH5FBdLpX/imCUD3oyybJzcsGAQQwsXCAeasKP6hUXFvTjMK7I78SSBR
BgQmcN6B+e3+/NBnZbPQEtDTM8bn3XqM7NRPlY2PjIH1haw+/i6IKebsPdktZvE4
wLs/WfT84y+n3++F1A99tJB9wwrp6n0dqlhsQpfSRHQG0M7n0YG3OUTXvqxFfcd0
hg8fbDeGFWrZ/uV58nwZToRypMjt6cdKZumqMYGlFhzI3AVEhjsrhDEnXgBZ0uIq
9eMNW2cIKZ8vTbdGB3F5/vBtq9kbjo2vvK+htVMxTaD2q8hXJY5dDBrixWgSFYoD
z501DNEohTrN+s2mrG2JG5NxoA8PhsQ6YNeb8CvVnVqHpJsvZ5w0FV+O8dufrpV8
5uhExYSt70G2dRR2aOqCLWBQFjv3lwBKIriKTEtnUL+GWvX5P9RTZRSuWRQc9q1h
+Fjk3i5TjDFhEBhrJRvabl6svYQMQ1rxj3DChex4+cEMSwN8RMAgDyIDPqBO/NUt
wSdUxo8ejPaaAKipd3jvoR255xSD5XukFqWkhBPSTXHGDyeamRCfBO4A7axcZxS2
JP+7c+1j1Yjrs2UYKXhqzvqEY6Ljkjj86n5Tu46wTuAutwodUzjFQTXARBkWzAJR
LZFB/3r55cncIbfNTXHgxxo1+iiAHZJDRfPmwmMjhvZmfxN2W6j8pcn0oF+crwZp
D9MHC2TSK0+v9l/g5mH8eBMjU3+4twrzQjMHm78mikHsi/ZfExk/ZCajo7VevkDb
KaPSzYOT6LkUd9k96wNEzDlZqu2jQAHixBeO5pQwX8E+z6vtaWYZWAlJovo1A+yI
h1wMKcYaGxrYJZ3mKUehMLzd2swg5ySjSHq/NlUKc8nVRpJH/DtPzqQE/0v9cKAL
oU0XZWCzdWJidQ6ZekvP09GfumPkpbUg4XG+dapFD0Uq3g4ARP2N572nbQ7G3a0m
dGnoqEYV0lfiDCO51/pg5UefLY2uc3mUrFZhTyONF6hnZdJ2UM6ScTep7TTE29eO
OjWxGzaZ2J6Raw+tqQTqkvCT1fv9jsB7Y0cdkPn1Aktx306QmsdM5a2099rjgRb4
jbjh74RBaKDYQih6hzC3+D5/TKSO6f9ED6w+Ay+7bpqz0Rld0+/ICRDrgDIDD29q
h41j8xXgPpG9loIPdxtSXO+3yNI0jq+5hC/m4eLE3g3XtO95fUfBE4YwIqwIo8X3
KX7F6zoSxz9M2uO6cETRcO+bFeo6B9tKmTmpZYmrP21YAt0a9XYBJnCjuKtAvVtM
ClER1NeojddH793E4wexRF200umksHIKoWNtmr8DyNXKlenxYXAuQD0sDBze5oYm
CfDM4Wz4zzSmgm4yCOFRNXiWABwn3AeEBMI1LN9AnkJRO4fTkixz35GmHMC/7Bmf
+02DQ8flP0rKelqaFhODC6Babi6F00AgRD0iF9euoV6XwlcyEb3ANVPPDRdCBo7L
+tLdVxY9ZJgS44Ms+TkTLPADTqIIzGdxPfaJIlqN8ydJB9S34B+Qocmbn5TN8heG
1v9kGfqzXMvKc4qF09jcNTz267QhmMBz9ySV9mIE6HJ+0DpHLKLDBfC+kNhBabW+
22cPgJaJssCALd1nejPo1bLt6WKYo6OcfoPKK18AFsApBVfK2LJukVOmAs2sg81G
kYX5ECFLbUTCjPsBiXMp/sqW1fcyo3oud6NhdCwEoQmFGAhvTeny2x3o4X8gN72C
Ct2SqMzTOyR+W5qOPZJQuTQokJDfy7skPd+fDEqf9NzZAENBmz0x495ZRG/EEmNs
VCU++tGIOuw09eoKayWtmWQMmz8eaQggTBs4tpfFG+10lp6iFPEvIqF7ZsXnR+C5
98b/VYgnX/fHp+V1nVCALd5S24M7Ao+E/7KvXAtkzubswlPSkJ0tOn6e9k54c9/1
pAHfcGu/Uguus2ayMF0UISjgtAYLP4Qj0SyLib/DXx+BJ5FwDqcqhBCVlAqmg6oL
8vqjQ/IfANfVW5t8pN7+cgzbeQkdzVQNADi/XbO2pxQ+2KdWuyvljOiblmU4zKaB
OdwHbZsd+InSu8Ne0O9CKHQ2eVE3UpOgnoOi4Xau86P7IkDSYTp7bYKSnPOjPeO8
ft/5DR4XPkOd2+znJPbYIfYYbLDi3/OALmmKdha7EXGYTUw1glWEP37LZ18pfPx6
58jz4XrxddZMeXXt4aqrcARMhkCNgBE1ZV8jXBi3msJHujqds+y4sD953snYv5Za
fbdKYh0AxraYxw87unZVP03NW2MgWLp2+6X2eRqeBengjBdMnbUpPZZ3j/Rq8TID
eML/BJTRYUjQdPE6yyr5szOaeQnaZgbbIs4lh38xfoRpU6uwNHbYwhrI0HyV8pWX
swnNOZznrfCduN6FGgSxK0ESJgmBVauduUXQeqgEXL8duE6iDK57ckKcdC8FQr7G
gcD1rzHuiH0cyUS/9EE7gavS08gJxv0rlrdzIKl/hht67TZMRERmM9HC4QQ2R5P7
USV1XtqhUHOot3OorXsAa866N48/FO3Me1Qow5rAWB2gbQE8fFzSf/WOuqt+qSHM
ExS6l/RRSoOa0roOfq8hy2kT7+LldQaiqXFVJlzkBQzeNsv4uusiW6astJfB77HS
6KqK2boLH4ZAmv+lwpW+NvOzoToqwL9cPfiuirZ7Dr15wrik8U8I0g3DglyExsft
5QPRP0u70w6BTq7TUSLykgxo8AUeWxCZhj4vh7/MZX5jhMXLZiyHrPr+cEa9NlIt
qEuaio6BjuNCtvmfZGf8Ku/wSGh6gieYvtU58OwEwaKwRTenrA8XG/7WTpHI86S1
rN6Dg1Okuua857UeJYzRye/jiRKHdvdizODWa5wE0oK+vldBl+IU6y17ckr4YkkX
DPuwUaiJmE2cXjgdshXGy3J9vSrhc5mnlp8lRD0tDxkPFUWtuDczHmTu5SBZfUhN
JZ/HrjIh7d+rKxbQ7MnS3hucfhHdZe5j0lLyzYpsdZPLY5u9WIBiYYXDQoGSnd8P
DZQ3hE3pS+TbzEmK3VhW05mzYgRnlyH+/6JPWZH7UgbmwxubIopkW8isDobTAINl
Tl/AdjBhBpYwAZvHfK7l51fi0GS0PRwatjdCUjb0vDL3khDKbzZ6Vw5G8OnDUgS3
ZRsI8hqtMhyXSplVSo8PDP1azT3YBCvAQBcZqIcvJve+NNPrIES5Uh0fS2VOt81z
imyGBePG4WkbpWMUqirPWQgcBixnDpHa0gK3Yaw2eeCK02V4SlXjQXBF/L8bT6N/
Ur21veKeB3MfbRngoi8uLthmDqfxEXyyNppAZGvTNXiy0SPmLRKY51jS9Cwp5VgE
9dkDuHUjHqv3waWxEPKac6z45UrZ+kYd/JvAkaUjcQ4xPbRWxqu+v+JgCvPh+0bZ
AcnetQYhxqcHrLCWFNmRfEHHJeUGy0XBX1/JecXldT2mfVpLzUYGmon/vGJtLvB1
x89xdGgshJ9nxWfAq2o4qRcmUTskCAJFV6rDTIyvSRKbWHHaqEyU9BtzR/6ogLTo
iPLJyybB6gKTq8g3OMhYRm515n/La8IShewWTVzM2YPWcDiTTiWQUSFQM975V+8B
59ScU0Uw4LfLTZIcrc/F0w0BMDn5CiGjYuyxEFxqXqkoJ51n46Mjrxer2gv7LsUw
AOaItrcI5W6Q35QQULoN1iqARx9KGxoiHRWy7znZMRD6JDE4617doh9Q5VrEgKHN
SMQp1OwMLbMcUJX8r5taN/rQyZ+OVGeZx/4VDDZtbX8D30is/ahtCZWbM9Fv66pP
NiLbrQFR/9YfEL7VOdeFMNuukk3liHAsfyGBMt2+l3Y5v5VR95gzl4ed49ZN3JxP
i4oBU65H7VL6vEOtc8cYS06awrj+kdAui/0c2O4mfa1j+MRTJ1DhI53gD4ufAxMh
mBd66J3SCBVUJTt/4mQyiaGe6QeDx7KjEnMeSad9d/zeJQrRW+MSYQvdGcqgDUu6
SbPyz91NzzFG+5jzUjO6GB/IAZJ3jlJ4Re1z7cyxXzhSQmQ74NASJM6MZBcmVIjs
S2zEoa8AnE2psIoLBdx8AFqazCKeo7hRDbXoEz591NKX+KjD4eFqavWloBWJWCCY
JUvdirzX3nx7T6EZcf2CBDffZ5/WAVMuLToyEn8nHCDgKSERWhAl/nuWSF3W3g2u
4r8w1Bv07O3jAhBCkobmfA76pRPuFsfIKIFKxdSWZXK4HWjqQZSBUeFjNdu0TdR2
5HuIwsGbVj5eP8AulJ0JkwAQLwkH57XmZvicBQXN1TEl8ft59CJ6Y9mTV9wu2L6G
Py3atHCVZOyrw157bQXsY8FJ5UggOsUdzJMbmS3x9DHsO76/ILN0guJjGDdTM3Je
Ksa04xUCJ4zCKe8UFZx7g50zAS08D8ufFn564kRoOOCciIvgBSxPQbLrx4JQPIWN
RhMG9X+/7o4BTg8RABCGYklho2uOoL4MelwirwtWcpNW5AZT7IwU/e6yChTZSqJi
nYXB1eXBsEKwbhaDW7lkjqdgMDz6UInKPfU512XB5LdQ7chcVL1+drbpvfs4IG7n
90sW4H8f/9aapQ7wDO4Z+mcKf7D33yhCKMWuGDOe+FfGOd4eZZHpQII4mN87k6hb
QLcNGkIBAITF1NvZfLIWJ6ibMDd4iUqq34VOFmJMQYBHDbmn6fwBpS/+o00ZlCct
CjnHIuflrKVjvk4hTaLjSEpAadslUb2sWqddViHF5+aHRGix3A9sox2lIj0ZICMM
/RR+5fU9ARMtjHB8QhfZVBieVGof/Ij2xwgYyvZe2zrKVA2tqFBZhlg8WuR9wK4x
VX1M8est/Xl4T/z3Wh4OmuvDOIMv5XIsZYoKmyFcBvpo6H8UEqYzNO/hdC4UTQg6
NwNgX/RJODt0s8Imeb1xL8USeYbd+d4stPbz3v6n/JCWIe1REh75BLIAopZlJuNC
zTlY8KPnLFtoZ2qDcQzvVgIknkCTCrvqMFKgxB/emrQv6FAWBoznZ/DXPKzgLTFp
hFAlfOJAwGLbQ6s1vJZd+5RF3Z5JlITSLdREFuOUt6QNjYHJe5a7sgm2OFwEVQbo
eYJDh7PwntUWU9MR3QVbHtLDgYcz4cW/4EOnyerfBQ9nllU0QgRBqjxR/R5gJJQf
rbj7eXwVrmxziFzCYeMHHWbtXItLADSA2FyFScShAYqVk0Q5B2vxYzYQfiW/YBlc
r1yz66c95H4TVXPBn7NoKAVbj88S38t7uXEf7STp+Cma3Wotsk+3/fA6tVFY0yBV
C4anVrvc3x6wy8w+iIs9PzYQOi2h2eZ+kAhTJSRipSpyfk2JNVUD3h1fHE+B3DyV
BYIDfjVxOxhpYw8TsUiMTL35LQhreiPEe17gvuWdSCqLlbOExCtbSSYDm+RYN7TN
zVtabzMIyhzrP9qlsXbAofhvoTCDrluXi8Dx++X9ep0gay/D9jLcDew8eaIFlWWB
McV9mctpX7EA+St979bEZ8LRjxfhp3H+eLtNi97qq7bF4fs7rDq4H4wxmOJ6NT6U
BbaoNLRaMVggowmI8lDo0e9OTFYhuFy3pGYt1QTZXTKmbM7MBZKn2WYHNFx/bhM/
mvS6g3B13gtd66YxaaDb6UEhWsueySYUvEawvpi63QBDFeWA8Qb+NlozdHeJ+k5i
FfbaGL44jFSAfsX4KkKi11nybgOKiEastk/w2K9LARbZlxvzGLXIf3/KUgxu3mmR
qYi0vNiefSJB5LeaRU4ZI6EzZy9428PA6bu/PzkJUW+2y+AJYpnw1l8m+LQvJTAF
LbWPryd++ngjQxJ7/67yFIAloJB41+T/K09gkczdQf8SVTUrjNcT/B45YWchDHz1
Qx7VdDo0oVu6wStLmydv4i+AcU9AcnDK9wki860QnOG/tRfNOvMptwSZW4UQ6Ct9
8Mg10I1jsrD4iyqeHzyv0BWXfTLo4WLBeAa9ZW1dCCh6sIqM0kZwvvAe+TxDGGa6
BdmINYYcJsRgS637N1JrWShh9fIl9yJQLqHjmqpsSeLN26Okds1GbPH/CnyObsXd
Ns7JEvt+U1jF0NC7iBlBQBbiu296syxE3IopO8KewzcJkygHzy2dvcjmc1I8AYfy
TgeML5v/Y8KeFXveAQYU73nfI73ydn2/YgT4TKh0nCwucX5VCNwrYX0bn5LkaYIX
icQqB+0q2yZ4w5K2jY7PPsacqhaAle1EJCFCl+Z+3S6am9ywjB2zytU2YpjIERbU
Z7FjIB0kGMqEaYtYKoei+hGO8AsEdqhT23Q8zendrNkzQadad2ZHDO6VZ1eiJJP/
YDyG8/4OJucOfQpr33N10Y2PdeREOqMYOgpVhmHE5I8i+gDij37qhlD3Zoaz6MLc
ZDq3eT+BVHhWoHkQpQ6YTOf2nB3OsxryoPH+/XlGh4eTVojxC/jW/05XpBeg1k1U
oJdC1Xu3wKgIeTbQGz0y/bhkPiKmA5TASXEM86H9BTfKnyktr1Kko9tdZlNwqQUM
NDUwPxA3JnFRogbeSU9+gfimCcUOy86r2P33KUSNsG0WzNH6SmkiXkGD9+p6/EXT
GJWITOlvArKZA1xIkQNYgqjT5EOPJmqgHahXqQ7x9uOlGhPF89Q1E+HakGOJHSUn
s70aTG337O/YCp9y9bTbaAAvO6Nxa4D1vR7MGnamFmHcJ0XDhYaiMSaKskHW+U81
isjtXN5QjHy7xOXuKu3yZ3RUj0mDbhsOk8apx77USG+Z/mP6CC+20RcCpTjbwsba
3s77ekTHpxVoBrIog2K1KPF2EQUEEsQl1eaCUcCZkmQKKXMU5/sdI3n01jqTQhI/
m1lbM1hWMh6wjKFwlI6ZiotP5ZeXlIKSHXDZMKfYhVlOJXPeazu7SximqMULuBpr
yR++vH8ZB6LDDFt/9U9mK1BbPVur4plc3GI9sgr3nmO9p4hDu4LI6+ELm+PCzwZB
tVpnaN0qJsoSQV5+kP2kRVDhJV9khiU/nyzlSnC52A+gIHE8fK8MCPcKiJ2qNPNS
Qw24XALru84GAZ3wB+NOgWL7PoMGdBIRgKnDIuSvq7/Z7IuSx4CkphhTQTvKa+CZ
s4MM8p/7q2Gb/NbRtWKZqVOk2cF77aJ/9bZKQ18IFA483p2WGt4cjy6cQNB/l2SV
SPYhSTbuc5jHFRtHjzMh38jjw5UFoBO3ZVoPqjUKXE7GRk7Dpq+MCHkygDW6oIUP
Mo8PXI4qJhHgW9Q4b1Iruk5rk/DshyjR8niMys3fkTDnEdwWJS1ojOJU9cTUV0Pr
CjWC7AhG3R8E9zyX706EE5qFUNJ1iZNLA9lMttaok1Sl9rNJyrkWg5ZN8VRHbOzo
QdHTPXXnQeKNhGX2mC95p6ynvTmnmPuHzsxlLFT426PMXsBt0BE2L1ofrtckYYJj
7bVSe2fJ8HFQoaVLT9YLPISpw1D4HGVdiy0WDEqJD0oVlPtH+/G4aHAkn0/0s/2E
cUOVNKEGAQqXPTGzziTY+1X913Kk8206InyKNLSTDosa2Zutc0SJpUPSrD+3eAWw
5HCKBHdde/sV2OgIsT0SyMYBjmEXYX2nD51vT3Rf+2dkr9PJMHcJjrvVM9vfpKGS
sVEqbztOTgqCZ49myNPLZZEjNOtkym6nEm+e6OiL2AdUIfYMCoLHvVqjD849zfv3
F0MlH2y9tCa4FYA/yiaWOYsynHDUjD/GmtkVAIO0IprwXuHG45aj5dW/9qxPeEPC
u/VwdnHEcIZje3ruEEh7tMEMy2ClnsknZm9MZi0GRkitpv321oa+eJ0pA/7YISXQ
WRl92l+DVlMrHBMRsjwC2TW7cyhMAzJHSqLvhWkwrkqX0Y9TQejDfUnZf0tjxQEP
TLU8vSdWg0hkuAMzVeU9KPQoM94IAFz1QfTR3PCrP4VgOJqZIoDO3KLt4znWu4JW
M7K8qqda+sFxJvu4kUMfFxBFPFfuGvdo9/8Z1ygqovP9+d7SSaM42zZd91Ptb2yg
2GvxrofxZzIyvATpOqSye9jDkrYlJ2YdS+BqQmft9Vg5HQPmW3ahDn4qIFaO15Nh
OpNVj+Udni/9IfT86Zphs38jnb1xwW86Ppkmt/LVYAASiW1QUmrIRLqidpHcMtMY
zglpFzWQKSLxgovipXwE/z1STreArrh14Tm92btYWKYo+a2oDCDnqUMsHN8C5UT6
z3mRwqRtFz9GvYMkFnDDQ/eiI/+GlIFVqnZGBsK0/0jDABYxJcMHPzWUyxXwp5pS
cJd9xbR6Ua/ridxrnV6SWvj4KPZLHdGgl2MOLK5KkuCjTrxKMihU+TMBvwVfCHmR
c58OrRLdjkoqV0w5AS6JfT4DWBCDiRgd0Dr2tvSDBcKDfyyIJOG2Mi+ejxsH+66J
8qKdqOOEyFKXRO44rOsakLZjLjiXdrQFqPkUBTXGp+yoER+akvwmexYTiftSuK9L
EPk6Sj7dtsAPhDIXbMcTL1ZwVLjeQRPrepeXG79OnPPaRuGcKB/bb5vU7SsgHE4l
oOjQDdsODIm/Hjpv2P09QqMdQQsEy4V5+g7fH4a3K5ikI+TgTyTOkiJWv2OGyrcb
46vDCF/0AwwZQeQ+O3BRnB/Bw4VBw9dnHZAVO92WJvnWHOm5Hwjo8vTlRNRFI3K9
xFn2PzmCQDakf6Sh0v4OL4LHLAxu5dOA0fnvNiR0RKwi+6yA3IK9B97Rx+W2t6Rv
8e4uyqAY//mSR6LHTk2A89RtbgGymwc42sCCbuPECqElbLUe0NS6JjGTKcFlGimw
EBkZmW7yLjT8s+WOoHm/Atn1sVd/Q2FCzjKoUU8kaECl7bVvCWpCq1NxSp9kPfvO
CrVIfQbDmvVph1cIGNuk8z3NF4kPxWj4F2zkzpc1M+BJHyNAIMgjAhVXOSkYv7X6
eQBGybJkmgHAWhln5hNfPuVpuCvEMmluv/1hAj7O/g6dwjfekcPVfRpf1m89AVKl
nLuLCMIVcnj7XhsGKMEK6SVH4pKuJqMPNS6F5Sx+4ph2umROMiqJsBnKzoGafSyT
wOi9EEyiK4QJGwkLuBLMtxUO4swILSnD9tTruwetr1bjz9uKkgoXFTaZ8goald6S
y+nLg20RHh+eV/8iJjaXhGnhRHp2f7fvvvKWz09RLLH/YAidFnv62gHjNuhkhzhQ
Ypj11JUk3GroBCmUOFxQSWof6frX+tltERpvaHD5ZnvsVVVWrBt3IHpr06G4Qm04
EAv34szuq5sXGQvJPdH5yyp2MtcKXKIDdRzLhWr+VWYte16cs/yP693VDSuflUyX
n+FjOUj4eC5S/jM8Bv+AunbglyFU03gnXHcMjxIJc1uIYqfQqKhks2O//tCK589K
yamS2xe4sEW1DRfnwXAfcqrEg0rtOGqjhmQ7WRihkG4/2Co8FIulMsMfbqnfjmjP
USr2lWrw9fscVQRFSIZQkqr/ZVSpL2ApHyijBo+xXBYvF5KWqmxoHcjASPVkefsn
O4edQnJBW1I5bBS8deADNsVTOK84pL9tYxpMV23t88VDO6txblk6RpRE5tqCDVoB
IIhSBhng8MlItkOImXr2XIFF61CjGU/V8EfWxvTsBLD00y9p/5YGpPvf9gBY28iT
iSFkKa/0ZJilTps68m9nL252Sd1xC9sx2JYbxXRp07ajIw15ZlXGL9D8gEN16BE4
qyOo8d9/8CAccHFymjQInTDK4fo2ZP1RTUm42InR1gNeUrg+MuisvCkD0Mq3Wydc
pTWKvBLVScypNplzfj29eGBqLwKOEjBrS7i+yFvpdZsBoEJd8JxcOxJT1cxNphAB
fOttXL04NIRXSpB9JjQiD+dh3RxUxQ8ydlzlHNtKr22MQLh8eA++mWJOvsazzj2L
tS7OzvXY5l/I3VorXHdeJC25T0k/g3BOnkRKUQd6JPliKOMmSwCmvmvyHFh+ADwr
ztRyZI5kzn+UItXtzwOc2H6EnGfiO6iqJ7j7B09pC14fxhGDCuDK06Ik3VPeVqMN
IkVp+3Z9FooZ5yErt8RWBpJ/rS+f8TY8sC4RPtOITbBGD3+8ChAHRUKBDx6pbBB1
9GTfWehQo0pUWOs1PpYX2Zfo+AD3Kd9teP9n5UPK6u60O4Z73GSS6+M96nyaxNum
mmFWNBYnz/OMobk1m5goiS9nIJQyyoShg4Luw2ImDN44Fi+8sc+m3y6G3bxwVY8q
9MnOH6HSb5AMv+bIRIe2zPNlMIoC1DT87aFgXqREvzolzC4cAPjWUR5FumPWbUTF
0KNj2buf7vEjbNMwsF7VJ5ec9/Y1pmdJaedKtdc4omEyr+HT5L1zZPujD4nMN8SN
vaV0dQ7JdxJi1Heg8jNpbN3Uy4uFAEy29wkXIWyVF6Io/6tBbFtrW5gE3lvRwONb
dn6mLCO785UgFA04tCz+BY6X22240yxiFoe7BfN6Z1pbi1yq3+fj7wmokuZUD0sR
r5lZQ53BmP7Jp0essoPQRdA8wTkTBHWiAIkFEAo1eJ/SvfTEtAbi1mie7fW/Fh4x
o5bIf1Q2ajp8bmmOg6g/UVQ6CUgpi/68Uj45nPnIEpdKZqu214PDXPpCXk5EBzYe
qSop6h6qXj3vCqAisShL3Sq5BYXU6SLOH4eklCa5bUAcaq4WzVL/GkenBYLJnOcj
fU/ilVSSLddEDWF7R4MBl2B74dEtgwGTZr3jrHGO5Oo2vbzn2aRO+dNOYs/L3cH1
ITBSZbALPzDMWcm0pipIq4xDlGrK3JF+t3UVEx2Ej1dKxFh4jFC1W6hvvcAM/PKG
qRDeMZfBHXrOI8AzgWjiTJnKeJLnZVIl7AlYMcwFDjJ6ZT4NAHg5BEZQLUdDvBc6
okWhPiks47Q/9vcx0MUgaDgn6hzse+QwEK/hZYaR8bYaEdc31iNNrfz9Mx+GBl9T
7gS/80/54819/kqRNHuQ0VLI/FveRlVEkcfE1CSqb4M1XdJUYWVwV0hv/vjJx7f1
WpthKhLBu2FXkJOr5AUCmTfx6/3DLVTmcjfk61DtPZP7DsA4OSFxH3vnXkc0VlQh
WkRKU8IX3a/m5me+1Y1/elW8/tXDA0/iVb6BXC08Rq/NCliTySKqUC1ZMYnZuKOm
UniTToD8k2oI/LxyTLJhNk9ERxCtixoevKomwwuIMc6Nf3NBV0UNHgQWwBp8kgPp
CcIiM7n92FmfECpmX2Ee0eMZh05NoHVm+rqkboJzndwC5Cw1SLZPrNIaznx0FKIp
JdBqm4DzhZW+Uwfj1LVtLPb6qO+UWw4tUDWX1A7Bic+BvaqTGj9nQnxjwV9uK3RR
ujSZaCbOzA8Bu5269Wd3Zs58a/1kIGeyykvASqNOYrcNH/7TK8mF6a/RcOseIwyl
eg/Ocs/N9vATBlX124wxuBUW9JFU7Y/duvnunx1Y08W367u8CrUZE9SvIsk847t2
+Y2tCFYY3gyXNyJjV4poLBab++/o3kWy6JG5N7AfY6/0rUNsTiJW46LZXbiw7Gc9
FQA7dvwlKUtJZS1QgrOlU4HbqC7YntnCDA7u6hWmEHQcd1oPa78+o0mZ5X9ah0Xn
FStZmycQ7BCbJN0+Ksmbkfx7f+4I29kF5RQ2j8zPBNV1W1zW5mJeXHNpT0QZBJPD
ngPwp/cxoiCY6GtrvEvUZFG/5gfHNLRTWG6zT6CgcwwhLSzxSTsHYSHDKvLGD9sr
Z8K6dltez4jncnRocjuu9P61m9a1rZBfGnCXssBa28UmkkRxQ582GN1qxgvYpRNX
LnXOzogLHakwpw1/MQ4NHzF+ccnEvAfwKU8NIelmjRlqzppsG0UPJJDlmaxcDmX6
GWZcIoCmPZGEzjPR2D8IjLcyJ6o+5psNoVyNIEfmpgL4IQM2k07pIKoIJeFiIEJu
HnwJoOIbdZUhdEqW5QNWXGuHdXlxFOsUn4jE9Rco2xUvEMggHsp1frjH80iSsQ0s
rJKyv8DQ3JV9i8gPrW7bhZmgHuKPaegess5OtATi3bSG75Swp/LKegdPRQ9Y4Ncx
KtAr2aMPCJzt2AHMuJp2myVcAnUvh12GRhMvC1w0AjY7YhTJiqJ3bh32Rj25SV1J
DdMt/0e//xIJ3EHr/mMEdJAp1doWCT3geuXOV7eHvFDPzhT+XNreECDFThAgFu4G
bdpoOG6qnPAHGsIkYm2CBjBkqMZRm4ND8G8dJIuq+j4g87vNzlEObHWh+Bafg7KH
kVkN23NNPhVjYCEe+w8m93DUf2iOhqyI7uyRCpqBUJ3bY+DcPArkeVAb+3GfsEHm
KTjDUu3m/HsX9FS/hNNOzd/qgGeK5zL3uG3OwK8eLmIMjXPSlhWe76/o04nGH7U2
feIAt9MOff8GyNG7d+fAuiY/SVluVPcHO5n5Uu0wsH0TCi/8b6X2HnWDif3Gntiw
bAHd9pYJAiE1RXsMv9QeNlEMqSsOrPby/pD74t/AupJT/UL4ph43HfdBxkN7Mgtj
CKoaLuCWJM9d1e08NvIikaNFUBE/QiilHKDF1c9MVdUj64YYSh9IrrQhBCiC8TGo
YNUOkyxagUlAbeKiwLO6auDfvGTeC4a7Ulk4kYKkfY4QJIXyLQ8NhXFOFp+REDoR
N3nSOFo49JPEZk59Bg3JJwBfcbKbSbpsn6huGrUbQ0A6GUiZrsayz2Rp00RVq7lJ
NTnS5l6E5UI57F0V/pJl+yYFlWxoYCSiGokuJ0WS1HqlAfa7WlzK8tNRK0HX+LTa
TGB9u6qr4Kw9mDAY6EA2cStc5bXijz3/GAH5dbmhxmP028oBD26LKEpZnj3zdkXY
O9e6T/jeUFORB6XGHYcmLbUzRo0hREl3tTmdFwomsLdP3gUmWxjq7AITYmNBIhdF
jH4oLjYvHyzsydy2UZ5c65aqMy7O9Y8Kc9liMjDDMJZCA1l2lpfhGEdcbiMylhQS
ZW9fX5oYdjd76rbANUUTdeRr+rcgsL+Ebb5WQhwy1lsm6Hr93q0O3r4iUZJlyPe0
MqvXmYjr0YN0AeNVsc7rEOTJ4A861g+H2sTfbXbvUtGEcgMCqb2pm4K1G+RqmEUi
vCpcnsy9oshk7175Lhu+X8UPbUVtwOihBIOTtpje0ssw5B0X+oBkpQtj1JhlQTPh
QUqNJEPK3dxjhhauAyA221ipRpsbGl0p6U+ahN9RcjwlYznsYxOmG0IsvnAZVQBZ
Zud4eheOYsvqPvmDJBTGDvcsGrvV0+IHSXLfD4UmqWZrq818J61/Jg6Ultfv3epG
JglwmCyE41f0ypxPXPwsafAzAwbSyL8fRo2jagVoFum9k78K845lX0exEGDA88xA
zAeG4bE/UODXRlNWX6PV26iL4kQWWdr7/QGjy9DcTVJ76vUBu7a29Eyu1mgC7wfB
Myqw1CW4SZE0AP0UiL7OJ6jZooZcF8G31ZQjm3Wgk0cClHznNMGNb5Ux/evU7JsT
EpthZs0TNFFd7i1tC/PrdeZJp5d+tFW6smnc3x3TPyHUF11RcWRcuzhvklbVwfur
50by+rbV0TZjaK7mlY21BRB+EBcw+aClRJMP38k3djrsaiJDjOpX/NeirPPcYTmZ
FmbVvHvE4FFHGX3vcdNjDV80G1ri6CnET2mariQjN35WO+8wXyJW8MjObv4bLBQn
kRHPeCoQOEobvz+GRA8IA+izt0Ua/EErbyqSvcIoVQD2Ndy5u7G+rvdAhPZM4jUn
VTV8dfVOmRL+nmihA9JlKAiyH+/GJUqmo6lYX7E7iAoDRvlurdniI75c90+NnMEA
AnHjCgcyeoSbABZvZCbtroAWykFdke+k61UVPvKzIGJ00kXEBumbYH2kaDcw6WbM
xCqJlicS/NrFxwIVLNXEtajOV29TGvnEACC54FPuClCjVi15SQYPWBkLgzAjbTxl
5qO3l40HOMIAtpBivomFronRhG6q4b50EUs+xe2puAsrmdcivDkqoH8gdC94JcF9
vRLRkTeVLmgl4GTgGOjhdURio3kfLYEO7zNAd4NnqYlEW8mU6G5Fm9E0LQfve4C1
mgPFpEBuOQ7g5kIdk0zMMsWNtQ3GwplexTF9P+nmuif8JIR2i2CEbsqIJ4fsDuh7
5GL65eNaQTa3vQnFe2LDqYqyYRgYRjIrINmafNuJhaCnwzeo+NCELUlQV+3233+i
Op6BDp/GkkJw0JH/J8NbP19UhPxxVpVMn19CF79dNuiJuaGpDuTB+CvphHAjNmlF
2liftKi0s/WZUStq8WvJPJbnpTZNpP/xk2WWG/tIisDY60Wfp/eebMZLjYu+4YZ+
nI4yi7pu9+rHd557gC7bNMAHlwiOiRsRJ7UQ1AooNtHHM0ycNLtqlV2BuX2RlJ3E
/U8267RtZhsGQcbhkSWyKOTT+jbrvTw5IdCSt/49ePgrU8DjuotqBs6I2ntcmusL
lktv0xqsNT1bSFyZJfgYjtcjvyqRApyltV9hzKX6ew+S6uemzMMZbWgV8Jus0KIK
V/o05bvSs/1SwJZPaB7gMM4xwQFL/V3j07iB3iw+oGh+R5OQcHG0wBE2eNa9dQQU
Q0WRSpKXQY6eGn3ffR6lr0wmIeofGPxVCviNFU91PTj921y83EdvdEZt/HyOU6iL
jn/WiuV0jTJUe3qxF3cNJOIgFbK9FwuJdyN6jGgYvVd1q4Xw1M6jn94YRdAxpabB
jVZa9zNw76ayVnX538QBVEpfGs6n95Te7bwj3bMnqhC0i9buZLHWFIcw2WeEo5kb
rRncH930QPtmWuI1HyxcJ9KFWcdbe2HXSKM1vVvQbmJZmH9t5leeLqpRFaEG8l4H
MYsz4O7KlUA0rFSnu1qGmCAyAKyxMuXWrEPfk77cb2zmP4LzRb8RgB4+f9MAk6De
T8zDfmpDB1Ykg4zPhzI7fDk4p8p/h1245Fm66F3godxZlT0PMw4dkAlrMHDq/Rdx
NFsCis68hiUK87gF82MKpDZtygYqXBeCgwjgt2VpXw5f9hTO6yI8ZQzMVbyhTIdK
4Twyg7glqvMEs9xpOOaFBFa6iXUeC2bjrDFf63OUSZF34GCyoH3jSb5xwLeSi/27
OwSoTvQhdp94An8EMGgZsLOoV5MHasGVm6k2TS1gJkJ4bmjyzVNRg38LOYF8FptF
7EQ/jEbaCtwvQqXxDOjSH2uwWNEF/BerKXCPJNKkB8oXV/Z0xf+wsxWugF2le0Bm
ltBLkqVyXKUMGe20i38XvrW2pTuDJwltdq7LLTRWu1/HQa9TeHCiT1H1ACP1l3pg
YK3vWDyR09NYhlo+CCxD/efCZM3zupwWq15gPTlWu8JoaZjCyWceP6+RtF+iCf3z
Qbuw0rcf5KuFQWOCX+mv1xlApwqqPh1dobcLZ97xQuX9uxkAiisN4Oh3Y5slbuDV
mUgPYyftC0Bt8kaNYexxc/FWDTYo3nO1Wedx1Rb09O1Ow3yavCjivk9FLyfBq88/
lz9mal5ymNzdg5+K/yADPXsliEhmFfd7Pw9+Xx9vC+TOUG0C20HexYYkGSOBLtfa
s35CFAbgseQfhCqmel54bxmAFqqugKlNUAdnjGeJqa2ykRdFITdgOlWTn21Ez+c2
3NEe3Fj1tYrGwEGCPtgpTlKAd6AL7BUJoj8GAviuHkKpkcBGy64lWABpK7txs6eV
+bcfx4hkLGJu574FMOXnhAh4g7MWA45a0OMdB1wwpUMFcFwFi4sMAmB2Bbs8wu8D
smj1XBWTn0s/GQ74OxhF5J7/hswN1pwF5Im6jc+7nt9R34nqzfm3Qdp4tQqiG8sh
3tMpx5xeWDJG1ylDj8C5MJUmMlnf2ekBcoviGytbiTrL40yprGm4neEhZaWoBsJ8
n8uG79VJIsyigBJ/RibpxNZhnFd36hveEIp1q75nOvF2PexyaWHezr7gwNaupt7P
mta2Oy7LZlxFwsNW/JXVhryuGuBePXphe4QpgDekfYF4DroAMpYkDmNTuClu6DCF
uqt4pYUiTVQou+N4i7ykqq1SakQc0cgfU8FilmfYmGO8a/yYM2FWX6K6jUGc9vU5
C9LEc/95i8jePZDSWz9RAOZoWeEOsb+7WHsUAW+pJcRVuU1pr/fAuPH6WXMSCN10
Qt8myqGPYFHWt8HwQ5+gbYcKj7lWmqmDulsa2z63rHMZaaLchNDveULstr05oTT+
iAjNZYVlFUYIXklHaBf1Aq7ZbTNo814IfwowRQ7wcHhqePS7NGW9re2SLD51QQhm
VfxZp67+Mp9d3qDw9mgWqbhFn26GvC2VDfy5i5dbL6OiBaoLWJYD60Q/aW3JWhVt
XJvwWvUFQQml6CcBoXZQGXIdyL/gpt9zlLK2zksqZRMc7f+Wvjw/B8KYJ078oif3
yoRaRcqaHpa+OO5qApPt5CRbwz9xsbA3r5QlF1l+Us9ROoSEZSwD/zsY1UrIQPnz
KQl59K4bOkdAL35rpD8jvNmh4Kg15SemKWVVPWa4XpEKbsW0m3iL5WIbpkmGVRSh
8czVQ95nqy/lS7cRmnk7pllN6lGN039yB1RJzrbC6UhSXb6KZLjBoLF0cxFhUFSo
0RGHANy6k2kzXDr+V3pFa8K165lI+/i087pR0OMPELNoYJjj5aUorr7okgQnTkXC
NZWMQj1rQMZteGiO7zYsGtWQqzJ0w0fBo8PRr1rdM53uFue+SiziKh6Q2yHxQRXQ
rmvrYRqkaUc/LRgb9VGOwk/AEA/Etw/Uxb9fmu2hYHOzITxYvjL1YQkxfP33BS65
t8or6igZnTFvUvJ55De7FMYRWi1TFLYXv5xDNU/AyGoAjp1kkkCZ/Ue7q5y2o5nU
ZcliUB30YjegJy4cNWA6+7hEE4HaAoc8BVGnBAqn1S6YNagDHXPKPEkfcku/9Sou
caG9PwMjgFQ6Xa7ahcOZzUVuEItHjhOCmBUTqBtg3z1U7jqz6a2LMlP28fO33nX1
hXVVcJBAjuN1ZfUo54UB3BawYQiTjw1bid4DUmiROVJou8BrxWxVUa1gWxfFADhN
gXkqvqdkJAUnayKmeyiBkgnxRajkh/wcMUabZZMMMszahdYfpDJzrT7xPLoBcaTk
VwHpudoW631XUyXx9oTWx3pvzwoyfU/9aYDB8VaBEuqVWikxWIJiTgaM1WzPOvQn
mCu0+YiABpcS4zTo5Y5+QpR2ZpUA1kAtyZkSuvgJ001+fshSFOsTBzVk1gYIo0o8
dviMbIeFigUvmIiF7khSHTKx25fU4JTCkhXywbo6HTEO0vbkTAN4OZdMWkg6e8Uo
7sGleXPyOxKwXE1TM/jN3eBCONOLnqVPHL17rzc0HndKh9sEmNla0UFIhY1Km7d2
AgnZPYJpJ9vkWhtbHPL6ksFmiQRgs0CJipW1iIhCRMjPrfFj0bKfD9CeRqsNqlK6
oOconBDjrWOhNsEfsxzPS6TdkvVUgO29QYaAuz0rOgs1E10UkU8BNlroFQ8CtPOO
EKO+kSdur6IWRgpmkxZwP3EGno0NYujrdHmSkhelTqDQRaQ6uB1j0NkdqgQrVue7
FQ4BkoZ4yjG5jB2kvDoqvvHMmaOMNsZzy66/qgLdEUgFcmAG/LQB3FwfeySTPoGS
MNQf1MoNSJ0ojXIH0LdG0ihbQL3FiVABM8H2FyRYivTvnU4BSs5ifLorSrkL5t3I
w5pbGeb3M46yU60opjwX7G3vizwEGPZon1Nl6qJ1XUHsJAob/8daOiL2lGmrAm2M
IBRUKECXx4QHc6a4gDmtIjq593AqBQJPevWfXhXMn1YdUQ6Ggbc5wCPIp6kbdsgE
ft+yy2MFkr7c74l1j/ZGhXNuAeU6AM5x+FOZu1WTfcUaHQVfpdwiOnr2RRzmpm3F
TEd7WY76KDMkMPX05wwfTOR4IjWQ/QopMLnMij87S7vvXM8peMcHy858AvFI6ydy
/WYnxA/6vcilQobyLMp/CyUqjMPUC/GkcPL+yqYtDVw0Sp0qFvbijyIYDi0VYzrh
eYjLtMrdpKiYyJHbWMihUbdA0IyHDNtT64vxIZd92euaL7foRk3J2KC4xHblFQic
OOM4+RED2/OnlSLK1iCpkhF2xjXvI7ecD1EkwEhw/m/J9t22cFhaPERKCIQtIxsD
l4gdqQsvLltGdK/vKnMPl4S+S70MUtOs77Oc9FUx7IX2cv95GcvJmrM6ngPyzpbe
vxk4CnUuE+564pXU1ckIdF14MugpmvJNrfbCUNBXgg1uUo5we7QEObyQPUl+tu06
Z2m9oWcZpZnhdCzkJr1m1DtGOqXmzS8b2ioJ0zmctApY6OcC7L8BZWeFUvvAvhAn
78cM9j0TcTTK8cxvZfnM6kXBUsxDWo83k2MoGVz9KqDyHbssH1pvpvC4QthWFP1Z
TVljCLnPoNxiadZVtpM0ViSjJyEO/CW1DjXZUVI2P5nfMa+NUA5KL28JmYH1Jq1S
nZsihgv7c+t3y9FOnBjMLZhOblovdU5uzC6WAS/GSo0Oz0FRGUgW+yaVoUlzr9VB
r51W2zcKM1BcwqBTkrzHuocajfO28xq64hFD2JviTkXViKHBIqczdrpOvrEvkkcD
dLBvNp/tWSwETr2Mg424F8l80eRTHl2U62oVzJDkkd3zl2WILqXlBS5SW9aY1r7T
SaNxozuQYOq+RXyJYi7Gaq+kgtsDBpPM0Oj/NE4MFP03+X7rUcHGKG0M0aq8bihf
uN+yO+xamPFbt0KWDjOJkgd4Dnyd7cVMuOku91O23KOBbDLjl3K+6uCrNFt06coe
OiQgO5sU97alDah+/Uh/DYeQDE3M38GjL9EOpg9oYB8i+YcBO3f+I+hZKofkRozd
CY6BJcggbxT2f0TkBqj5LgAHOY3dc6ot2aadiP/3mOgPFXf2a4K749QkxUR7RAcW
vjttOfsiwTO5XwCCep9Jl3lHdwz/MFKxr4dIwVqbiFNz3iRUcZAwrwt72oUIyHel
ALLTVduO7q+0GuJ3o1zyGmqkC+yg96w8Flxvq6rdDemuYqrpLMcZ1GYQbL72z8Yp
uW9MNlD7Fr5Zuvfd+8f4jqTlsUSGFIcj4xYSxcIYb+WvWODSD9mouaojROdRNpGW
FoOuCEkEmo6YvUyf/zNc5FjWia1Hu5wijchcq8kb9131Z+Z3v8+CON9PfVwdtCGU
4IdabJWZE7Lqx1TKgFKYgSu9/h/EJ3H+anxnYWMzvNBIj6kQA2LsZn/NQTyrVTO4
aLbvlrPgOyK0WOWg8yDE2FUL/MsG5gUgh5XTjmpHcdpCr+YxoHyUXDduwgP6VJlG
zhE9pm9cw2hPDeAt6i152FNgQSDqyqV6JQ+UjJdYq9P56rB4MxD6NWFyrocVh1nx
WhoJX1Y4BSj7ZQupEuEtJ+Qg6PWXYD462A/iFj/Rfanx4qigRtNN0Q1FrdHYigUa
wAt4Nr5KfWnNn3lotYA3FbO6svnmHeeP7MWruEhbjK1Hs4w3a9pcp/HOAH/frITj
eD+F2bwAJALKnV9gnzzyhjWpBS4uWje1t9BfFwggd8QhQ3QDwpiWqAfgI3fPZm8Y
jYy5ImOrytQgKLQZNef8qihYDcpfho+yh/08hp+xotV9vwgHBCR7V/AWGYUa2rt8
5FcV7MOM1K6D9ggjVHs8lH1DVZV8NaF42ImUwH4tfsBwEuc+zcvkRH4MqxmyyxAs
k4Ncf+QmO3DoIR+IKWlfJGh6b1CQ0deidu1+veLBwo6BPVAjNQaZOn8SEde8jpjI
5/gJq8Em3zn37f+s8X9iZhCaD0VmgNH+6GZSNs/DSGkfiXMlT68u41qVIBTTntty
KheQRVzLtZJXanNLwC2xbG1o6qvzXoc6dQMGzmd9gr4WyKX6lOb/02kXGiOCz5eJ
bqvgsNADCv5CwoV5lDWaSWQjALxyxI7YPSuQNUGf/EtC7mISw+P3MjiNjd0awlD9
j4XKwIFclr28U4UDDAZnbbTzVLuEnFTn6rUneMlRO/ERsI13u/rIcM4OlibNlhKq
k+ofcVpEgxl9u6sLvy+NFNcb6KbnH7gMd7Jdy7o1OtkOQa0KXjX7ZkaQDQTsmaxs
LaQKyWoAo53RmLnqgQTAIbmi3uVxOAw8wxcbFVHTFuttNocvGloVs54lQz5uDahE
MtNT5OgTjbY8hCtNbgoZ6exeXZ0a+8U87Fojg9baxMhAr6NMzKXtuCg6AhLeRWD4
hxtS6Cycl9gvvp/Njz/vLY5WQyKK1U/li+GvHom88MuQMPAuw0ThXDY+44LrbuBT
jJTYJW0rqD1RKEM7pOmYA1v4Bd2n/bPOuCpz9hz3bimFHhsUvxmpSe4H+3rT4/Kt
gHOIC5S8M2hmO99Q+E03Lof3aWmNIuVHZUvBQpgBk2q5aBONVh1O867iKH1MWJp/
ibAR67cRR8HhHJCH9VGcSy2SaUGuGpNdKDOIiIKZykGRNOLmSsThnuFCn60gNyob
atx80xnRxefn+3WaeTGZiizx/n4PQgP1chk5DASV7M3E5eBexEX8/LgM2iEV9+L7
UUnDopbbz5YbEtQaO8XWt8m1xNZgvtzKahs6O/aCNxWfuIse9jJckBbVYgXMe74o
SYaPiWXEeQo2ZtFMU8DMYe8pwDKD6cZUwbKaUoZq82cknEDgV8nMcMuYsrSsIl4j
ux1j6YhndK6dsqX0UkPkqvfUEtasBrQ0Fp98goOd1qBeIK8O/vHVCQx52Hs84msk
ftEphdgBiq5ENLjhQA87m97BkQczMLWk2Wd+ue3iG7RUww4u9nN+JACWDRxWmlyB
0UVLz3XCJv2X48W3kPGZWW0jX+WIt6U7kts1fI3he912+uUxPkyvq8u+McdnmDuN
5ZHUjgouE4xx4WaTlXZQHaqrUEzWVih2uzMybkn/F7t1SS3DT/ckjSHXlD0Kb5bA
cKzVPOtunELpbrqhuwDzmJYx0f20D8JrP/PaX8HxkkKdzOQd4gyIoGivc1imw07y
nIQ5lEUNPkWQdlFVkR9T+NV3WNiKmxW2OMzBLq2gAPp3ERN0wWQVjbkNN+Uc1W+P
cxSPXBwe9okz7rIHqQN1SfThqB9+xVe9jxnegHjUshSkBl1eOXFCAV8N6/iu81LU
dR+Szmiazy/Jm38kC0VD4WsZbit9C9DZcMr/G3Tkbt07s5eb2dBDYVENG1oj0rSy
dH+W2jUjkL1JtY5vJEO4OsApdt0YMj7nkNMineHcv3S5c4nXNQDQW0kdbyAgZNpm
K+7sJm86YfURAhdUcX5agH1/uY8xr1ADDikZg7oTXyJgHOAIf2om8NL4grxuLfNB
l99fUE3pThWW9Qzuy2bhR1/fwLvDdyVowdxT2x33B6+CAbiQic3bHE8TE2tV5Ti4
vCHl3kZNs72peoQLdUxafobClfRK724wbvBXJ8+ZxJ7qkQ/l/b1XIAiN/d7Fn3n5
unRhjShmlrr/kNM3z8SZXDeu+ZiHWhNBIyAO7K+fGrZdhoSQg4hyLNi/HOYePUqO
U5nkTR8rnlUphc705YQDmKhQsIgbj6jrbUeg1OCW86tiADrrsd891+J1naCEnGzS
AAd0+30me44UHwl8RurKQlk/TURgPQ30u3MLjT0tI/oldByIAqe54U7WabqMkBsT
5ugRkpcbclOqPHgZFH5bk5H35iRTmuf2+t44yAW4vIqvhwSeqBiQwFbm3sbSTW7J
tHON/W0lw1jEZHnGhojzA+peMwq8P4UXsacJptuSVr18zkiDeLvr8exmUHUH0kXc
f0RNTD0vLFM5iX+z/w2PLwVLxA+WWCJz8fM78DFDBL4XaS7FtAXMHXLcA0leeS4M
6fz6XtQYK8aoK83SsG//hXRLOjJvnnZFP5brKIJsDbPe+HyKCuSWVdKw0G6glmEr
h7zHKN+rYhDDGuG/yjthYcAVAZxfw3CdzlcEpCmiaoczBrLZQm/7oSbOP8cS9D/N
7obBPVC0soj0Qj2uKkhSso1DfYgYzKGiqDud6qyD91duNlxv6q6x54dlhtIZNe9q
LcbitkALoYBc0vWz75dGNfQjID+aGnsYRQos9TW4JGfyJFJmotVrZyTclKa0wY0R
A17CTHBgoQXhsc7qeK24hqvZurcJhPy0I17rKNZkZMTJVpWj4XOfQn+goMV8aa01
xmkqdZzI1FQ7mLh1RtEQMFT0HeXMG7Nqu0JLHBii6qi0rcJN+ojBYnjegM7oRObz
nAn8JVoTaGoAEyy5uBHij51E3KSlYsZdCLFTEBJbcYrCrQFdV0JxtvyAyrAoBnRE
Zx+VjVIeXkZT1bhjKjabkuiA1lPdFw2hRiyPuJk3BtMWtDCeyu5PLxw8HNmXxYw+
QRUZqQ68d6rZUVgF+YZybp/X/pMP07x6lwyq2NkjZDXI6ZbxLfcntiitNCO51m6S
/f9kAD90w4Emrt5lTxu1BfpMLEWWAFv5zPBIT/+3GogohhSlWfOb/maUp3j61S5T
28JUTrxESq0W9vN/kzo+4Hd1yKjLVVI9dMpY1v3RgkQ1w+1wzSDQg75Qax6q1Lag
3rjgKOBuF+KJ6AiosNO5RHlbwM0kz9oZn/mKq9N5w9Nn6N7c6TWo4IxeQtrnrVmi
O8pP8QH5ABpbS3GC2d2eMM0G96Zy4hFagRpyVnpix0/aRKI6+Na5I+SQY7m41OAP
c3yYgtCtCeGPGkbxoVJsfqb9M8t9q6wQgzNPHclfmffitxA7UixCEovyPMLe1L3o
GqNIFO1Z3Vr3EbQ34vds6k92j61KmTNAfuCO6bAuO1UXQZ7WaCviWZ/JbeSTCwEB
s4uG2SFSihHsbM+R2tq//vgxcJdYjPfXU0VanBxua+AuOKhJa5+gY38efwff7oqN
5jeUIqvNI4j0zT9RJ0ILQeAxMopLIHCFk+p3MViWLYHKiZ+GzWjy8KJpLmRJBYG9
R5mAcjgB1UsnU5SRhT2OHKgoVp3rKpUJPOGWkISSB81oA/dIir0hrTfA2W8fV3N9
DMIXrQXX8Kxwv+OfYsnu2d7+bu8GgqoMcT8MJ/cS1SOYTJiEyTQg8wSJbHa2ibxp
YvvWuDTq/cZAZMNrB6EirAoMIdwl88BCGr7WEZNN2aeyirQeF4s87hFjpHldYNXW
HVHgRr2+UMDG33d69b3UoDPrku+c2RgdZGy01mjJTIh+VYeZfoUPm+LwK8F8nCdO
d8zHQEeTvPjhs6JhYUhQ9uLxBrJEcUqDpH3+uvF5T1L6K6NA+f/2OJtZS4psLxiq
2uFGhjP+0Cv5JDcVevYD8LpgfsorcJHr/VI8zhPxFQHxGjZqDn+Ketq7DfqixvgI
ve6J5YZMyckaIMEG+88W80jP4E9JKtg1rucJ3cdizTPyP8+h/somI3vkzm+LJGDP
uiwX5+tvIX5rpjbUaI2bOx2JgF2po5W+yYCX20KEyT6BstecJX1vVnRrIA83aR+6
zG0Zdk6ebDpPODdUDMBuxAE0s7Q5uyuW3+dk8yTSdYaE2a7k5WLXj1iXAb3azX+S
cSosTafcSxHTw2oed+Hj33FAybBrWbZXg+HnjQBtHcxJQYN3D7jtlPcpT6H9h2K1
T48y1h8x0j4JdFriP/Gna+lh+OfPiqvy/aNbgdj7ntGjykklMHwXp41ffshSwfcu
wEBoh61pTph9p7D6BMKZ98ctV4PpLLMsSXgoucnk80Qxpq0Q4btL+rm2s8U9fvO0
eBvRXE1lcO7ExP27jO2F8JaWJw4gnrG/pBJjmHc+eZtK0qdpHMSSrejD71p4wUJy
PIZgsCjDPIX5wnQp0NmUaeqtlAv9yJECmL2aJ93rBrjLlfc8HuX4E37yzGTewomp
LSrGYhjRUQr2uJBeIrthkTb+NNDmJLO9dXe8wMURt4gaR2HtPvZMdG85+t2WUQte
8nHsInFQjfj8S1U20pONjubdsznzDSKCRWW0rvRUm/wuX9gR7CvUezX19gYJS5rS
NGzuaJjsqFhkf5ipPHM3YWdktLgOE1rJ1IQEhUcmcd5VpnKVCX45W3+Fq2va04Yc
YqCzZapMhBsw4O1ZYuBNQ1CC0P77WVXG66SdnwEhoQ46yP/hfDzFal3HCEELUC8H
2HO6+TGM4X64B7HzBghdc7wumHfAT1PA8AIqBdZ1NLXa0y+j1XftLKKQ0RaOu2XZ
TraeZvq+MUL9gXGyD6Tf3jdhX8tLt4hPy/VIhK+Cn1pQ1/ohCZTGwd9izitmZq0j
QR2H7tMGbxe6qag/h0+y8gvbOakNdaOgYVttMv8uY/h0TqkKAI5AQU+iqjK0xxZJ
4lpc5bTvK83DyRKmPYlwAGBllpHzy3BpUZeBJrJ2OUA+7ZQj1BR1zCfNa0KbY01w
Z9k9kZ76ZJkM6utUiGFM3BpU7VcKQm7AfXDCrUtDsiCJhYQxaZiRKusUK/ryBoKi
DHU86NfTBBp17mbAA07EgpG9mgZDFIM4EpJDNCGUOcCIJ5ENZQpZ1JuD5XcCt5+I
gmkewyZRN3hgx1imiIELyC7U8Fvw0Qbyrrk8x2Z3yPf4tU0Y1KPYBINRtWTmquE5
7e4/d90Kd9pL7V0hhnOU7jrMsyqT/Tb9oiogpzJ20So9HIHEBSPH0WAfRFtFoseg
O2XMXK1LADGkjMooI0BBzAwKjtDGSdlMQTGzKUAhcYmVtUQnF9p6npdaPx8JB1v7
qFnVACSjdZqoa0UkWgIpwEZdV+dKi9MCsryNUZZUpmUs9KYToBqxI1gZwrdj18fl
dgaSRbYDr1Whd+gziOIyO9AfO3ILS3uaXirJwvDhzmjARNh/fpsafmeTnBVxRdvp
Kn8GBkYtcgbvsbNtDnvSWEZaw2j8FRWZcgs6DFZtEMFth30WnXRKfXStj0/qvxSQ
EwmGvBNYiPyr247KohTodvlJB4Frf3Zeb+enQCY0OynLRRTDOWeE6ZJuNI8N+JDb
XgEe5aASULCwo+++KIOHiCUrA/g/Vu4v3aksKIgOiLLLgw2i1TV14bpVuTmcjtnI
BhASm89o3tLiTZKknUPVFQIVwweoxVAmqQBH5Kn5Dz/IunrCcF3/Uvt6iY+5TZn1
xXXP1PUhrIfPxLJLamT3VmnhrWDMSvS3UPXVHaab5RGCHNVmxW/QbRk3VhrLE0n+
cEW84e3aIbN/fHS96X8dviK1QK+5Dp0/ur/OPTyWHWsa/2IkMdKEf2HvzidqshST
BTvm6yBwhBLTsCNXmpoLM3zxA1W6vJgWtCZFl5SVaaYtYhWFk4w/zU8DojRsGz97
OWws0O17bDgjb5C0C+kBeifvTpX6fK1UMrodFudkdf1fqblOpPv1Ft43GFIBr7Uw
Pp9bK1jVvqOa+bBCS0rPJcVW40dwW7hqYtcAaNmTR6/ybUJdInIfFcPIEXBedEdH
1o/oFdu31OPw7jDypJhd6xitYSV9uFmFv0hdCNm6aLD5bhZav9n/XA0JvKMBkzhO
s1YpbrvbIPcPQvr5XspylUXVuQ9M9clqbHPacntgoIb4JCfumaAqavjTAcqxx2jg
1FZ3VM/3AnUImr6yvILEXiWzxlxat1svzxpxaPYhrCmdlrrSpPesxRYRYpRN69h1
/zgcdO9IR8GxbEqttuTOkCa32lxNLatM36ivQcXpVXYQUXJSV6Pgm6TxFgSGthKV
fE0xytDmikW3q4nZK06AEVCtJ82qpa5gWWFVEvLBoP/1njsMQcLCxFM5T3YZWiEc
24IaASxHFyIanPE3VOvzHEscBwmPuWkWRH5IHs4m5u5+sTecd8pdp1lBKFsV0T3d
sZbKmW6JsJDp0wFkGWHzIDO0bc3Fpc9zJpzYPd1RzYfa6d36RCgHWjZY+0EbRb5D
BHtg9yQqfwQpWlBZisAmc2fH8/ly3EfvwBnP8bE0U3gpFmdvoVb8jDyHMRHAZlmK
h6lxBT5BuZpbTcfLDsFj6QAIG+Vi7WaS9oF5LpQuaCQW8hstJSRU1m5GH0n5KLUH
3az9TlH9kdHaiDlSdsgdMnzXmY/CmZVpLnOqvfPGFJXYv1Lck3kXCOzLK2CNAcDb
4ygtNZ+kmZTjBw4b7H8l2tAsF92j7l2xy6UcGDybAHlPWVTEwLS4F7bOhad35vC6
GSzAwbN4vSgi50D7yGVmMOUC4PRupcWL8cT+VKzlM1XcxsypJSicdaCLrGe1dFzr
m9w9beo8KLocyVOKtGBfci15CkvpcIXdYthxvr6NZa2zrhJ3P1zRHI7Kya2N9HnQ
nmjBvNl549M79tvMfPhAQWBeXGiKIbafQ3KAyjYi0GNT0X08p25GbZ4zmrb6W5vZ
s5Hq5Xak5uNxY4R2qD4wNHtVJdoerpSfAyIoJTuRf414/J4sKVF0iNsQuDE6QF8e
OrBScPx11PPzaHuNZixomidXj3O53MKgXKbMg3LwhyF8rL1jpcLJZ4otPdS9dzHp
LXrVYEsj3mqgzFnM3sUm2EtNO+FIxWklksJnTBeW6QBPOAdfU8+BXXbdiNkKDbv9
iTevCuGkCtsm5gyj00H6kA4mosMY1YCfKvAHvPmwsRf2dg7xumKj7MsQYRxIjdpQ
+BQ+HnaRyiw6Zx3lxQ6+H5aeq4mTWluiQ5G03maPNSvz7HbB0hOle+EjtzuTbqHT
n/3rVW4R634U5GuiX1C4XeqISQP8taDsY23wZU+jQHDcoxv80GWks1KLltyZj3fI
t+Dwe0OAJL7N3p88lLMmFM/8LmbvRihEdOudX2UKAme1kZ2Nea5jkc48naGIOWZk
jfmsp1GBO5nSGIdbSWgJvI7lDLrqYg7OqJwVsDoazY9v02RdJX1SaEtqaic5r8Bb
Q4XO42IwCoEaXb/dgClBaIiNbQONzarVBlizF9t5m0iqwH2YiVnab00el8tPr5vY
M47ZT/GfCmink71qQfrcn6oNIbZLb5XDV3hDKBX/oELs0O2GdJQ4v7UUBuapGLt1
m/AyLQX2WOLOuY90jVyjrWG88ZGGBvdYVd1mDrv9vOdfAelbHEcSeH/iChJ5a1ls
BD9UdiQTiAjrpzHjFQegM8WDYRrigHQMIe8qAYl58+xfCtH3OOrSGN5Qzpm3vAWK
sIlws7nkfq9uuKxlQadeim6bEVoPfeE0YPrwvU/sR+9TvfYb9+yeN615JudPi/+L
gowjW5bhXqOc2pG3g6ODVNi0Zd3u+51XzzsQe/HJmmyOjq8RJrNmVtFeHyFPTYPy
8wUGcmVVXxl4ab6WbQprJ8laCWkQUIjWcx3bJ/aw84RI7OYWn6H+s/NJisaSHkyi
EepYBqytiQie/bqslX+T2und3YtLKg8J6TG/h0e4kwirQD/oob2jQe/oHulGS8Ax
H/EN2QpuoJ4NgzxlVr63kQ2MBeAXkwMPma218gze1a57FefDO5wJBVJt4VkjEb0a
JR6wkLnUo0OkKtvCzgoUY3lBnDd1WT78vPzATWJK2/ina1YV4+B6jHrTsnobIAKj
k2lJdMs/FnDDY1yxt/sirtdMTR8WlteSW3JCoSppMrz9jJKWvOPD3vwHtvNvx9+Q
p219qbJyzCXG1uQnDyYhiLoVMhkGLNwG+tMXKa3NVAzwmOIyp8OLB3nQyv8fx+ho
wSdPx2e6vXkudr5Ox7R2XF3y6S0XhLG6STS4RxyClKfgYxfTMsoVAasYM35zo1W1
GuHTAUSWtpktK7brLOfPo0/zfCYXFntC+d/wFpsGnSV3sNryR7XO35dn2Kh03KH+
VfngA5kuzACLMaKrN70KxNcaKHGn21ZlBl3P9dOE6yS6e6UqlSfBjkgH1r9Fiydk
zprhkzExG6bs1lKfq4OeLzWEL9lY1Y50xSvr05ASXndg8TBcUwkTpAhQYUj2LQ47
d9GkBF8ZMkGBzYWYkzSzWueLoghXSUxb63yD1txgtWEdrJKNq1GJB13QRbUWh6DZ
3/GPRWsxbOlCZJA+21LYJ6aoqXuwI5vE5Yf3GmxnP90tmQMR5tk7WWFPLU7iTLEd
A4yzvdxAvSMuUTVlHbgFVKtTH8K6GLYtPoPx/otSxWIFV7+nV0cnf75qJDX2gS8f
pzhcVJgC2H9Z0L41o0nWQ3eje6wjD/G39vvpoQllzuSvfEXyV1952BSmovNKN30d
ifrdtl+NmczdxIOFMtm2qloTUlwVP9UjW1VO6eQkXmVIgB9/rs4RYY0Ca7rfT9K1
rEEeMms8L4i+bMADIR7QST4ptIOEVjjyx/p5SkPcIZSMRYj+gc+fDd9VxtptOpMD
njU4UIu7kiNvexUDF4y7UNrCabEjBUcLsMc9MxnS6QVvfJIpVSRTywvKt7BwSyub
FlT4ACnuY2TJj7EaNiHht/FLJGXFRaftglA1mszqqQos+Kxsnmm+oqVFnEwAxcVT
1GG8gaXuumO5rkS6HGbtmA0zYyyisbakAcB9NkSnyF+KRMccGWjkQtPQX10UvNmY
3why0mqVj2CiPbz10i8mnK5z/A+p6fHZN6QVyVklJ6msn7eEGZZtU3OdDb6xIfJn
jIfgzmrgRLd7aKl/a5gp6LCzKgX+bn78H4jKkMwxarXsyxJibWVZ2Tx2cKLYLQ8q
RSquDWxSKbNgiqLFozy081hcPhR6TpWhYLUrbrX+5n91spEl/kIxlxjvHU9JL7PF
hJUyZzs/6h+sJFy7xTvaOnnxEjUxiLokBo+JNp4yiZU0zIjcx1C0n2AKtdxajsop
m2BfG6mntD/FxQWRp/IAEyMY3bDkqS4ViV1xl4v7lFptJ2NEuPsMYVsUiuUO+wXm
ffBfNeUKqI3eLcDmSF0IUs9XwJ9nJfUYaIbKFKG6Hk+VJFQSm4SKKhb3h4rg0pbJ
08V3hz85GCG6rPmvr6aTVNzAceSySS+UwlePTDFaVxjyBfiQFj4s6RQ55jCC1cGx
18YwHgke6l7pAXOKzE9q+9nG0GgPogpEJB/Wt0cUCMWqRh37V0wnGryUUGrjprmv
ZhFxsrLpVow8IGjBu+55jiFAVB0ivc6oFtv1jEJJaO+i5YcAuKsrHAA6KHDNbpd+
FDDVRYmcOSbEg2rXXARfdbit5obUXWpan3DBTSVmBmkpRxMc0uIEg55DEG+OXL1w
q6gEOAIu6YcBfkWUwnH6JnVWAnKAl/9AU3lj0VPmev2OvMUpcQeDBZs5uUHf8DlJ
Xi9hGmSOCMJ6O+IRMMCgHIBhFtFz6ZerJMfz+tZFjEM=
`protect END_PROTECTED
