`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ffJVHLw88BCXBaDS0L1ywQxzgY8MRaamuhm05edpxsdAOfYJWfkhV2O5xIzNWSMx
ATBIc/F01vpbqpmRP44Nhx5dH0FmUEfxzZpjxnfb1K9kCjsCUZ1fyUAnEXwGBv4F
sJkl0TzbklpgTbkBu5uJreQsyHfrHpDRMVoZGpmhna4CI/z5Cbqb4+eTA6PIzXNc
pH2JYTp/RVZIKE9gMBZ0gaLKfiGw2+2j93U6sRLRUJtNa9uzNLqbQNA1HmqaD+ET
pJp1YqIOqFB/deVCVQYuutAuiD+lQZRpj/3pKb2utnOPga0nGPosNP/3CiM3EMnf
08qlStrcDL07HpXEkibfdcBLvs/taNt/KuodyKTd6JV1IGOGUxnT+XwS/FwFz45K
ukYeokBVSdWtU8c9+AVopf7I2LsqjieZJ+12M6MVYsB3XJ6D4bDxaTumgumucKHf
1oX83xw/4sAvyXtv30SuiULbhsFvJN2PSk4Qp08lPsbDaMS46xI/YnIxXr+1d804
bg+ea+0DilsklTccUKh6a3eQjSgd0kHGz5rg7VfKSvUGWwE/fDKDt5S9zTfl9rmT
hM7K4qlfLfZnIp/F4iC6ObM+qpxY2+kfPFnCSmNzo2KCyEmpyYCaPbB5WpxtXeGs
LnU0G02vcs9XYgGb0Ze5wvhixtaMZ6+dVpJIyvcv+TVISDxUOXDQ0jpQ7zbzzyE9
w3HX+9OPJ0YuVnl1ugHRL2DstT7Qn/c40VZnWWMQUjw=
`protect END_PROTECTED
