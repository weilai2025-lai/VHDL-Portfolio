`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CowwVwi1lIfQMWjWf65precMic73KSodDVz+FO0kSsvTb7c1bbznDFXWrFiv55+9
JlyuBseH5GH3PwYo7Zwi/4g2nk71nm2rdLRwPBT2UfpA3ugQbK8yKWDRrnGpQypJ
XthBdRcjw0vLZjc5copHkyqrn1gnnBKN9grfmWDyIsUCNolerZhh3vtEZR2pVW1d
RO5WzjYbNbUTHPfRFiH81NnEniKbdTX4LM6Scm47znCgD1J3JJxJq84e7RKtHLc2
wSVyMU+tAUAtyCL/T8PyaZjTUCtNrk5hqXxILeWH5nKfcXVNq6DJF7GGUyd/EMbW
jN5eU7Jvm0nouY2CGjMM13kjDp1MNbLZuExwgdcmL70lD6vkuDOg0/72eMZOMxam
Gpq67tQ4xpw+cwSet2K7FDQXSx9uNtePqB17esmEP3UHzi25lCPDxWa7bAT2Ks0L
AmMKJe/RGW00MN/VicOYYeiMjaYcJfmWAlv4LQw3frWOs4INFMA1zcHxypeYliO3
3c2Pf9PS8/h68g1ANPol/dt78raetQfreqHSIIEsYUGPzsY864J2cblQsxw1Ir3/
0ynJAf+FvSdlhMTIV9XNsdH5uhGcFP4MIhog1Vm1/ctVV4gmH5IL91b+I6FZ2LOf
7Vh2mgwp6/DJWGAeI5LgSWJs55+FvyArplqGpGlIiUrrXLb20lcl4H2AyHznBwDn
7lw+m6nhg9Ese0iOdxOQ0VkLjXyb65nvdoABxUnu4WrMH3cIRDsdB4p1R7ngp6AU
Wa61thEumi5D9Bh5lsCYRta9JV3Thg092mQA0+EG9QMEDI1SFxsHY4R/W+5lUFRd
zq34Jcp4Wc/T9ZWfsFBFy5eDc0IbGYWM+lt0GNVsktCu7zSpqJ61/iF3M0eMEzqO
`protect END_PROTECTED
