`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/4eREz8D0xbJ1EmfN1AAK5Zhc3WNWoOBgAFM70+QtFOQRifLqaPhS3sZD6Tsxwo
xbMnEAlcjD7W1oUj0+fnMr2TRInTXSv5msDJq7QcfhsdPxXZZlJ50Z7IYK9hcJ2t
9GmFSA56v/Vr/6+NvzJtGZDqmL4Gp0PSBiI4tGC4EqWpf4+pAQq7756KOngWiYZy
dHjLZbLrEyiHR/ApZvIFfc2xyxydzupEcphgsPbkKboBsxDwRt0AF3FocYqMBtuf
0mrG5AqfA20OnQbhWRypL3YIEY0oScMvzzxNpCNLK2xgVlUIcyhC7D6g51WPCkZr
6hL6LkwOe9bLoNR8Le5tJ/PgRcy4AF0k8ULRXdS1EraLDmv/tRbgsTDJ0LUjyL1U
`protect END_PROTECTED
