`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpQtjyd0VLu7Pq1RkkrUmULiqQokL/N5tHAbMp7jKNKLVCCtxhy4LNZQ6aGS6RfK
E7XhFxNA1jy9Gs3SgU8USy8YidTS8harcL4Bjx11uXko9diZswvx9e1f75FrgJBN
MpETmhXK83VF3aP0sm0YYEkbR82vja8GTGmlpQNQNN8yxgSuaaYDCObApCEcDvV9
lNfFRUxmcrzsZ8+ijZwvYGgXNUkYXhDu7KhU/ZIhNqneH4F9DM90lYoO0J6/WIwc
Q32soaJONNiPPcpcMrdEcqSrDYE4V/x1AhSNIFF3bfqLqnVSgWU1TTYW1+n7gtL8
jCbPhdB4APONqq/kJ9DlPa6Mk3ijtAqf+ZUTY2Wl3i1Xvb+wsd/cH+pFahf9w4c8
cAoUuFsQcscXReDPG9j30g==
`protect END_PROTECTED
