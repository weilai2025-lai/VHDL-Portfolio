`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/4p2RPiKbqj9LiJ0ECeKuMHo/lIMXTLZqS4VIH/YscseHcF/4anajBkSRzHNeV0
5fk/B0GzsO3Wf3vWuo5xmCJ0ztveK0mSA7h6sQIwn9Tgf8Ey99lkyugYyaSriwR7
jSNXa18fLFgrX8G4QQGTVKsML06TDtV+HW7W4Nx54PPdeV39MfpFqx7vqcNIctFg
D82EE2TpAvl42OKMmxLFhr1f+piuZRrdP5EbQbahoRktKIthOfhePERBtMAoHxZT
QdKd+jOj4FF50IpJILOxHdxas8D18A9NOn85+03LVWhs/HJGpKLYaI/sp1zhskiK
lTzXLpzR6MGqNaLg4td3su5oDYjVUeV/WSvmH5VGsgSngL8WivHO0QrFz+XkKknP
4QeFvj/LQM1mj/4m8WOumfsrm0Sgn6h3wJ11G30v14xtHZrU3Y6zsicqxkA7zJxF
CnTWrq30jyyaPE3RHL5Q7Hm2O1A6tMhq1b09nmTmS2qacYySaWjT7ZQ7E4UlMr8J
SpvJALn+EYYm40rOeEMv8sPPUfyqSWXTtdc7Jpu8rV1rPi1+U/2vSi86ePd9QIqu
+BflzGnRQ9MX+w5SsRCFBQFj64ct5wF00C72klyXUbuja0AHTdduFkq2Pkj+rBa8
COCSt0TnsVIfUQgwmMphP0w5YNjEGPI57RrXEJ9i9E9Za9kCHDBdbjOGDobxEjPS
oa4zEZEq1JCFMUUKKM7y16x6YvNHsdnXqyEG0lDPy5tydnJ8e8msDoLAAxDhpllD
KJRaiC+bd5NnMjkCyLTgZsqhzwHWiCZfk+SAOh+v1drpuOOazGe+se9No13Fccvj
T8hXGYu0OZaxIAbekQXj+TuxATWbpIZo56Mgoegcf6Twoiu2GGLHEZyqpfZlBibz
5XfpFueDmwpQ5YPvtI24g4dhPNqvzsFncBvPNmLBtqCq5rKNQUbolaCo8a+ei5pH
bVdCxIovIG3pMX1SpEktCcsvFybZblr4AqNhlo3PlFzp2hPSY1GarQjWMQA207mz
UKqM6c1kFJ1/NomvhojPAUQgLzAEThXG0PrAo+wdddOZI9aYESnlEQ1GSvGCU8S5
cx/jtLUfvD0K6qzzcgwfyabaBoe1DJpVKZX7mymhOOcU8qGqrldSscK28D1sTLQe
vOBqZeZW2thom7/jPCGsv/O6xut822dX+ABw5pHKRSlH+ZWcNSEF1ObeqCAMRcsV
WZ1At9jIo0j6DJ76DxgH+xK3Zf43r8uqSweNcOAPEZGm32oSyRkvFatrr4zQutVz
`protect END_PROTECTED
