`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vweWAtn/nK/YTJb3bpuO0MvJd6oj5s6Qj6a/zqK1DUdKQAqmVK2T8xqBDWEfDLFw
84i3sdHzhO9G6Ely8u2QjGQRsCizLVCxmnVFATLEAZ5qIrxtFLY94D7Azx2iJ56I
yXCCTYu74TVXVwJzFj7VVJdoFRCNcZQylxbFUZSHZr2X9sYEwP1Q+JXBYkMoxnwx
fPhwZK997EVsbLwqTGNUZ5YCjcnbk8JPnQPoPlrEP/jB3uLviykZcvY61WqkFBLK
U7YE70M80/XZLhzbwLU9kgiUe0IjznKWRC+Q9lVkswYSZj9xtz1MYui6QKQULk/f
J7/0Zp+DDRrrC6FtFmLh9zQuKKpZTwUPziTXw8yQUxgp+PI3xyLhz9Mi8DbglQt9
a88Msmo28yqzHFtFWm5RRhk2eBdRXHxtMOg/OJ+8FGI2+OQlmL3Cg5sERdQAZ3iB
/2+au1atpWKOLB1woM4Xuhh7aW8/ewexzE+eTXEYX88=
`protect END_PROTECTED
