`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+CS0xGpv/rXIAWn/+FvEnfKnGkQKAHl/r0kuxudsf0RYeh5KGHDnpXygUvX6hK7
weGgSrEHYAWz0NB4lf+/W8V57/MwBO8bd7bTknauJVe+ahWnnOezUcTh/xU5DyZ0
npc4sBjl08bKZdjujjKEQe4JyWL6L3DX8P7OL9BXx5ItffzWvTi9oIufEoOsGURM
+d+LMB5dip6fr+VraiKfvhy/eyLOhBsFrckMUc4Jub//Ru+m9z++NsHizANfMDRq
ojr5YImlML3UdWmBE8uVhu3OeWVjyrqF2QVQ4pGG4PapUP3mn36uepnwCkxVC4eU
QDFeGLMkib8h5mQNLSdjpUfCaW94Bl9vPxwcK5bgB6ZZnVzo+BykjL2FRD5hSrQW
3iSE4eEqecbH7dL0n2+z7awFCpun4LGaEjac8frHAnkoyf+iceiAW2tCq+qP/32t
vnujUHNgrkHQG7/l68J2xY9VgNImSyST9S2pYP/miLiw6Bf19OYzgmT/AlJdtUSb
oKIE2MDVdfEKV087VQ27E1hCxcRn9eMVR6aJHAuIOIDAK66h1IhjaGcNhbXENmXf
3eaGKGbEXA5tOfN5CrIk+h8GT0w4mns4FX9irUeGKOnFZQ1xq+S5ZqCj+zYgl9s9
f2zsJiHrtdwowc//C2juiX5TR+bpIQt4HWVuabE23UXzsmSu3ELjLmv7TxL0TK+k
5OT95UEqpS/E+9WEjmoi3cFZFNpTQnk1C8xueN9iIDfNRBMCzjQIIH1INhiuIeZj
Pln+xLAAfV/gu24xr3kJ0j3EIKeXOI185+fNDnMdRjOisINCejAiX443zvn2a7eW
syY4Y9hCHXVJ4A5eRB91S4jzwsFwz3xgTw9acmrGAzf2dxB9aMPmEWL8EOTwE22v
eCELtNgcDVWQCaEYp9AWbLtZkcHE9h3zBm8xSgnBeu55W9jrrmWcf2JQuCS3QoVz
xhGKGfhRzq3+9W2lluKjP+6maiysvnm7oExENL0RKJVVQr3QLhQkGpYGMqjXBkrd
VVbinJl6Agx0HULeGxT0Y0njDOkuyGfmS7e3GIxpATLydc+ooY0vsU3W9tS9x9/8
kY823AvykAaTcD8SBBPPqk/ZW0h/jF4ANGfHqo+BVgrkztE3Y21NxKBv78+6emu1
jkfPpYl84p4Gayi5sOOnARLmLB5NP8C4c/zhVp/2SkaxqAu8zU/xSOiVndM1h7ll
4+4takxUPiZjSPQWU2CGMh/UAakozwDfigG2sAf6JoPYpjklZ39h2ezwNqq0eZSf
F4cu5UGVACmTf84FkCrfoCBq7CWSMfOAAmrYAwcfPaxIY86RjAZmKYApN/x3kr2C
utGbUko/BTuPqAn3OQGY6wlRZhN8Qvpj4P2IHvh9Xbn0VxX/S1BmcpIVK+g0vE65
QfQlAFtVphbdvXecx/mL8fmkJLePXEGf/pT7FACknzETi0ruQgTzOI/Mfkr5D+vu
7ypsCERwNK1dpt/N4ePBBDUs/EQOujVjvbeoHz8t6NS+af1DTqaeyYOxOlRM2QwQ
8ioAd/5dRQJV8CozLdXo8NZn5vprD1nhxVJm+Of5DavLgBKhJjYLcny+uiK18bAR
037BK/HBEP+KciLHTzHFQUlVyexRqRV9QBpGCEzjTCKxocTo+5+8+lUtVx/+n1qK
+Xw6jwR68SoBjb8s8/H90Jt1WhMB/BrCFG5keBtcXHeeCWPBwamS3UiLgz1PS1Od
B3TEMMoKHr/EttyBhudTTPkf98nUGAy2AvvvnFxgv6DaFUXIr7C6ChDsvv7NkYE4
nnAJUdcDxelfnYRnMp4FJrDuFkBKlQXRP+FFmzS3sjFgOFsYU+FR4ZFqSw+83/kV
WOlMN2ibwEN7XFeauzFWmOGGkidiKnwjnv/hrrKK9BTgFTP+s5dwaKnC7FfU+HsO
M+rG29gYSpMdYINu4nnvm383TwFraxjNaeUE4+huanAz84srEbnFPc1wV342SSnu
laXjDvd6lKJ/Kwrot2HwbUuTX014PHALKRL7KYzxYVcWcSIH8Fc3CSwkpepPYyAQ
WK0bCbCNEbpYDpy7EmZxme7ObwwKTAdQ+qXb+jpLrZjG0Jtc+SAe4zaxk1vR2yLo
XMO0QhAYIUU6noj6oqldXmlBPhK8JesGVea39c5+HYRXG3VuXFJwh+Fkl70XR7qC
vqe07kC/jdKV3luMwoe7G9bTcTcgdvJwdGHZUpJ7L2MF4TMC7/KG+nw/nwRhbK+m
LnWaGVXdDgZzPulp9OmmMktOJ1DMvO8pJxarlQJ5kPdYoAOtqW2lX+7+FWF/YiKt
Ry5yHcdBo2eH0oseKI6NHvIcSXec2cypqP5SLgvzxrl5J7jjRpRKLoCF9H79myMY
4QgGN71jnNlNi4tkgPTRR8cHkgzjzqem7jdJYl7IpoWkIaT9y7fr2eevkygaFsO0
D512IiBh8Dok6gXeEh2Y6q8anAd5EnkP6qo68eMEMRT2j4kAtSqilj8D3csz4TkZ
OugciPuQQCjJORW+d0+hBYa6efb8i8gDo988jioicpFJ6DTd6YHjjXPwR4rTIuJH
BzKAeSR+u4XPutKsoFa+tonszoojJDVeMx+Ob0GXEsWe9FgvdymfHhAMimqjZfhy
hHnrg39fQMGduPmF6o14OChIjdJ0aumRAtxL8spo8Ah9/ejhkxUj+myB69FBZE14
SYoxdBTE/8PTJQFBSWhBsjODULm54NPf4gB50vKh/ih/n/ANxa2MbKw5N+kYRAGC
W2Ha9cD1aU8sETVzQFHpjn2L0zClQ9EIzdHvq990q81WN+mLbCY46t6cZPmaQF4j
AWmW9sN2+gRGqzhlQQLD3KzH3K6ADOmBLeZMfxms5vQ7hHjqhxWic0u87SHy8efO
OjHg4tjnFRmgIWHKzQIVYA==
`protect END_PROTECTED
