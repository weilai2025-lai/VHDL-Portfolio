`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oar5kGNIbNwIGvvFwZAgey7ngKs0YzL0sLdIpWYjBdbPOa5R31e3+9ZKG88Y7D77
N48XleZfI7AouJdFrA96qR0QDBQF8Qf00SdwIj8EjNtsB5irZC7HYyYgEoHVKMi6
wHaFLZXL3bDYUBVE3kEeqzA6OXgmWMXTmxqaO3sDhkIJ0tfWPxIFCqVy32Bo7lAN
QQHCdC/VqjcbzIOaXnWddqM9ROHpf1nWo71kVSduZFFTEw5R7TZoOz8P3bjI/Nkc
9NW6TZgWuXELUYXm5libM8oKLVn6VfWFY7Bs/r1qXaWqVbzOCQhiytlgtgQkQ3YV
O0re5ymY8sPRbgAHlMeIFOeuSfzNKnXBFIPGCFL1spyOZpNtFYd9K4DhTDy/fdLY
xHNns0FeCs2mz54DKJP1V3oypg26TxD+9SqQoj9gP/hS8PRu8o6AjtuwjUWCFWkb
CN95nxEVXa7mfpcg/PU8Toapgcj8s4okNC4Ksyvig8lO3ZBbV1f1Ze/QMzjJK7jq
ykICl4ihwlzHqt4wQvnLnWck8HaI2/2JnVCk+mcnDgQhY4tQLEq1ddL8g1LGyEr2
eOuqZr7lawB4lDQYxedhtpheCD9lqIv3e04xyt0XYfINh39ihNpj0iaB6X5lBnkm
K/GbQlAIPOM5LGsURwRPXwNndPf+4dfsGXb02FIuFyhChnyzM87GiTM2nemQITBX
BuEjfQpV8idPdGGwoSbrPfvRxS2eWD0zP/Y7NdUFs6N9dk/EvtYIuTK8Kk7gMzBq
IgWicjtPFJoGxByF8w/KfEz3HSPr5TQ4Q2A/tMvw/I4GjgkX4GF4zVoaPGLXkjMy
L+HdlSLZKaV4aXdkXFScYZ0cha5atKxU4XeWnWsfc2+IivIc5Bvlvi+KCkNUqjeM
5i/AO7uLBo1VLEOGbXaFgF/o7NERuX5v2WAdAr2V9oJ11lWCPnV6o7WqjbaHMM0O
0qs06olkVIt4gm4yRxT+Z5NDzGBEWKAB/Bw4PEO5Clqld323GgfD+GO3b5vlCUtl
0iu0g+QgqddJfXVBE30ri19xnDYQO4H2Tf+MnhxVoR7/elC3K3VMLxiivCEbCexG
zQyBKOxaoXxW2L0wNTrhNW5Av5ios5RzT5IxIS9iKZoAeHQsv4U2if6ReLNWIh3j
EmcWaYQjMXtZ0SlpNv9R2YFmXCSJLndKno8ROvs0Z8urvH2taQneSjO2jaWAPpiB
QtNAKC4X1XMPkMvOGJ9leUMGyxYI8owAB3EILRm6bckECvwQQk5NSw/nag0Lndvn
08THm7Jd1D7qRS0cAkogYmzGIhBNVN0sCbAIAS96sJYVqJK7nyn4Ab35Kqsc1d8D
FCjz1D5Axj+27488nvmHD0HUDH5dUmF8IsBWgpMUa8YK2BBeWbbGyA+Nc1vvPGzV
omrdwyK1u9WhMW7YB7Fx0QuYAMhyQzX5iay59MEG1byoyr2LcG5osoER3jGjEQzo
0tOMb0Ftrl9OVir06jDpsXPcaDwl+2kU8kv1cwlv/eL87L/uaI/PSkOGj6CJds8t
lik5V5DlPyBTQFMuT6IA8RKQui9vrvBAh7CnoWjGNvohRlDaiy18OaRDuFNh03T5
1nQ+RHdgIwhj2ivBuFj/Q/snJRHH/NqkohtSwo3qngE48hMQz8rzf6iX0Fv1gUKJ
jYxYDTB7QBk/qD92JqA4TFnDPS+SmNKmyKoq3yEywgl6OWHvelSOGbBvdbxTzQEt
G/s9IyO6kl71yAQ5Jk6NmvkRX71aFUvaBaBBqaCGJeWgtTszMt99yvFjh8NHwGSR
hPUheXpLRVDADO4LNtz8vquyLX814XZD9Q0UFzu7DyHeHYsShU0WT3ZZzX0LO7lJ
/g46Dbwphh7YpvITgMVRBwY8nyKa6bsP+EBZNZClWcZO0tSSS7o/BKTCFer4Y2xe
KLxqgWkcOzPN0gBapVUEtmO6KlRhmfD8a+5y58KtJ6kNrVyMz/PSLSthB7hgdyXq
fC/uQNLEr0YLHNvgtlD65w==
`protect END_PROTECTED
