`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Vsd6eQvqPEjgAJuYF97GqCtAHXfsPOVD8arEIBZN6+haLfnIrLt6lEyaTRtR1o3
l5RTSV9nSGAxiFlBNTmJG08FtVvma0laHA66GQxdaOQ7/2kiWfSGfTSvhNhyMpOZ
KEvbFUPG+Y0PoZS8ogkmxbb3j3mznM6PDDkdWrsXp6uHBGhbD+nxOubY0i7O3sPO
Ez6zE86fuRXYb5mr3/gJsQ==
`protect END_PROTECTED
