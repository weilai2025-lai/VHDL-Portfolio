`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBIuVWM3b3GhEwRXwcvEKz6AEa0pkPyg22moZOs3fghXoxoMxg5vTAMtiYFPLGNh
xuDqr3P7bzxJm5C39MZqAwnGjnOCLlEQ2pGxzXYBYUB8fZgnjQ+3cWk/4luy8ThT
0AbK4p+hAfhl+LfcnAO8JYKSzLkVvp+8TBUdsgpXSBt6/VcRZP6VX61khAvaxR5y
ILKVVLlvaKBCScs31/+Jc9vmAtRrK5XefBTyPJ66Hxaxg48FCJNikX1wpyMagpM6
BwSZKO+yJ3gHtDHmXFSKtzHwPzeQCxD2jIKbUeJ7K2Hk7fdHLvhCSKXr1PJBtdgr
GLDV+W9sTQdig2xmz6T7CU8/9sZi0uYGclMQp6ffLstk4GOyun1hz9qIsFVDxL8V
PjKw5W/SQgiCxSw0RaZzkQO3JYOLBRIcGzS4+DzW6Rf+kjkPOgMR5ZnLA+/8USIh
dMYAsBGO857wKn3c1c2FteWYRSM9C0kCW7CsLl6Xh6vT897M5mliLR9CBGhmUt3v
nbcjtMvxv4d9Sp5UfqIagW61jlomY2mH5UanIipWmHd2nMKkagIItph3OW651lD9
iH8/RKr5G9MYZkSKgO8g0QFA1Sv/5Ky8wcM6WDqUf6v6RG3hDQPby15mkQzCyVVP
KgdaAy7GbqDGZIG2zyS1n/x9m6SHhEyyvvkXFQ1LrHo51Buf4goKe02BKOw0Nr9c
o6Fnz9Taw/a4ffjo5/agl5Nroa+Pn163bJ0J3JOub8ia4S2Y0p297pFu9A6NleIw
vJITDkwIdJIEHufLA/VE502qiOniGVc1oC3mBrj2TKWG81UbRbrZutnCUYZOcNAs
1rTxsiofNrly7R91uGT5Jg==
`protect END_PROTECTED
