`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7VsALJyFalejg/w+pPp9po92l2RsSUECcTkJRjD5nBDZq7TUcwayJMWEXPkfKef
9uHrchC9OxdNROApRNaUWZxs8gOAFf/w9n2U59dcWNaPJo/RtVEIiSfLhu0LXiM/
gtBk/1HZuo01l0UIsCS2dj6ANh4+Rq1y1340fohixnY9iejyai27XpBjh1+I4zni
zmHiBX1qvOBkdq6ghHiJba0VXZ/7Ycf85pnK+D+/HcPqRRjZj8wNC44swZCe57zk
Ju5+bp9AmIPULN5hmlTTQnQowkzg36a7xk54ToXqbHu0tRM2zUvxb449Fgj5bl4/
0y+ohPfnaDgeH4sr6emY52+lXcML3fDFFcOWKxfIn0t+Rsngc5fHhH9RHFA5Vtz2
eONCJ9kNy+HJ8ZQ9GvGr0clDbSZOOBChQkWwkodUqlrcbaT/Tk2vSKieRIW82V4o
K1sEM5QnCkBlHW/ke1Jl1J+Kri1pqOUgLrbWufZJ8gsQ829kecs0dzvzv3CvszSp
CrHfkQQd6hH75kfspbu+ZDMKCBE+KuTe14Fp07xZBgspvaNkXHCIxL7ir8PMaRBx
Q6Z9OQqsMm6FGZVw0LH4395aj8DnGZda4VW6f5r22zSKSBFLBu65mFiaHJP8DfjO
rchlUrWlxGwvGQNdr/um7u2g47mQqGbOyhQcoRuySIz8ZjYRcE0FVcB60jCPXHHp
3wu/Y20+QPihMYgor5DUL4QdlxY9pKvHj07KEj5SefB/AnyYnqzGAU05uB2FnTpQ
LcmI7ILuLqGGCEfKU1b617FIyek3SLkJKcCwU7SKjkqkPdfzM3a58OR0mvPW4dHl
3HJ+N+NcJRuxTcpQBShgg/XAXeGuzjcHpVnFlWB9qhKNlqr/sOBWy5LBVkOOgPdo
T2F2HQCkuOPUiUaVQGy4GhufzK38hychvwAu/wsR212NGj7YxR+zQ4gUW50f1tbH
tetlH+Q35BEsAKNa5Pk3NDwpi80RwxdNBXeA43Vd0bU7CznC64zJKdCJ5uZ64qiV
uGE3ohlNjwyXLLo2EiReAcZhJGUlrobZ7Rrb0B7jrgWDvme/mAgpp3GS8XmUeBog
Isi9nxy149QbIcG15T/9kfTFaqFWWpzaP27B9oPJGa1fI8tVE+b13CkViHKTGa66
JvRbUGimp1ZFRLpcurzWNuLHcnK7PFIHa2HHYGc4XyFw0CopIKbazfm39Wf29dgQ
RdBpFd+NS8eU3Q8uuYGqQhEMnCXrOT5O2BK14Ron0zL4RT30QThKfUyOtYs6DglU
SAga12p6WU8cx7g9LG4pKJB/BT7JdY8bdaUfcP2VB9EU+KYtBxwSyLWFqCNwILLG
uRwjPdvkO/zLGrPH56yxVXdkenY1aGM02nCLXLX0f27iO4slsmA548L5mLVGRih/
8UkcJhOiM6g/YPlnFCRteTvplYb14LLvvsljqr6ZIyWuKAHYUXhrZBY8/blV3Wrm
`protect END_PROTECTED
