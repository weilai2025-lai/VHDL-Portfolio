`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1yGBUhvPr+Y/XjGThDSdvTl6uT57rKA0vipJYmHuvk23bXaiZQkTsg5i+pQSkTD
h62mb6021WXgzT5MrwXoqVzE3CUOwwnji6i6uXxMZpj3R+i1X2JiuyEUt/bqCrB6
zKQA08FUzbfHZNlJGBgf4E4OwL1ef3fTe4A7UQegxbUAyEL6F5JJ8xyvV+H4f9KL
6Q9VGq22s1RrAv9bxafG4fW1HMV/L3FkdqL5M5mo800aOJIBaWkrAOEX2Nqvdr3M
PXWyIyh6BlE16cV8BcpqqLmGcGzArXiY9HH3yTTwSV7iqeiXU+qsJDw5MaSiKS9a
x82GHyWGmpz1lMBs7sThQicSAYvYj+fMVZvN6BWfb3DXEJw7LU8QueQR0TL+HtDg
dnfNnc8l/38olCpu0MedqQkmO8OEGzDJjTrX0T55NsdNonkWJgoQCJKK9tY3HpRK
t0het6zyMavzx4/27uc3BcH80ZdEzPfjcV1wnaC2gTNApWFry4u5C73TbuAbnIbY
q+4bXKg2yPgVHN3diyCu45vEqDejRzpG4rLYcl52Mrvcfq0mNyvPELtp44g6qCPF
fhZDmz2bDqbMXZN+9igGg+y80Bc/i2ehXD4KjWYbb10RNaL/MrQF7gyXzy1/ROT/
qcgRApfiR/fnduNRaRl+WyyvbhZ6qdk5oYv9mDfTwHalLWSfwanD/Kh83j4WsI8J
uztLI1JkMY5D0Oev0/ze12YOUUyi47HUFe1qiBX14193N6f0J5PuLk1O56eCTTWV
35eutYj2VCU+Ab7BkFr+bQo/13I+5fVVsI0lcfM6IHWfO4brIxO2Kh4POo30OLiI
xaaV2CuXKW5IIVQaqdI+/jo1CN/1Yn9mkboaD4tlcfKMauX+g2lN1ok+scCSn1nX
16iXmH7lwwMhonvhMVoPB0NMRb+kjXp+0TFsvubGeyFsZDzYdmtcVQJUNi2emf7M
pnxUiLKP95UpjohsCv1/G4QIacV7IdNvkKHghMcjq/Jykj7eYHU4TUE+AXFAoT+P
Ywv9RCzKWDrykZBHm8xKA8yBoaUyFpfWzN9jjLzEHz1pWAQBHSJVtXm/pwFumkJ4
V2aF4NyWubx8CwFW6wmCkbY24P8qUcn5Yb4cwva5qg0apvAxiwXQlUlyDbANygVa
BTJs84Yc3PyETcCyW8L25PoaZh4njKklVvayYnmr5cD/HLFssMTJoODxklKaxBaf
AYE6dqpJ+Hi8UZ6HbzAyneQCqXWi3yhWuK2v48lGigIQImKcT48PSalnA+t9ESEz
qCkwg43SlG75ArLfbXYMjvKHGNOULIJ+Zagkh31O0O5iT0Li1IXLGcyh6EHWkBYY
fwKbZrPlDrL08nAJKQF69yBYzKZLUtN0YmJ4g8iOlMT1tq3QpMNHs01gcjhagKJc
XFm8jGvCmVe+YhLb9GYeYfKewHKehX3y/niZzeeN+nA=
`protect END_PROTECTED
