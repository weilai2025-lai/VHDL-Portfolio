`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tu2d7AC9YGsf+77p/9RKZ2OpOKm8ccfytRN7t0acrz0PhoRDi3M28XD2xykGnEkB
ZUCKKCVFA+vVY0HAEncbg0se2zlefRPg+/lKvq1M31IOhhT6qlA61VYUw0Q5ycuu
4I5bI4omO5l+wIVy+6fOQiuHYH8I2zQieS5Bm2l37ubSANW2nmdwF9JAolrNiNd0
hHXUWUp3xTTZkafT0wHgHtT/a/3QvtAs8a+eyyM5WxyQb7MNXXjEBv+30tYQQq1I
U6JaPDPSKHm5tbETIlwdtWZPQ7t0B+bQn7vcZO1aCvHvn8IATUhu0BqPy8x/zGkX
erf/EcpSGTKHxyjZEm4LtlUMlYIYgHAMblQRoLJu8gZN9YTDHqzvrQwiSdPCMzdT
3LYkdXfNt2Str8rCXtB5aDPDX44+JRkhcT+Y+YsatZNwsx4PZ0LYPUrFDq1zcGct
q5Zceefq1BkKGfZmlLrOvQOAmAvEmPwGDDa05T1eQvRfbrLWyp2/C/ZzzsAzP62u
X4xOrzZpTINZQXda2+ImX9v7v60bJ/VCxEUgy6l9iGCnsptIo9GLnRhtgzeqARyy
qB0ZfEK9khww11ugi5gS0lo2tZna/hrYIB0NwxVCESGdbmz+7goy8MJbo8xMaj8I
GGPzMgFI/8ST6UPLsZZVcry3f0Jn9h6h/rka+ZwG+NNfHX4T3b8ZVBWEukYSO/ok
5jRQKKN6Id0CrXCdcTIXCvvkxSWloPm8XpSAVz5rqYPU6PIGAokORULRXLAWKKRm
60/qXdEXk5dLYkY8IOuJ6owcZA8YDaMVASxLubcJVYFTwOsBoBG4O+8HkE4F47vs
abOOikYSKFgpSWlFYogUcwlCNJ718uiXRDRaMyKJsXLgdX599mqr1x+NawNFN5Sw
7ihVkdRi4umq8rmfo668vnuYinVMdP61MHkuGozBkMOl+OsNlzX2o9Un30uFDN9k
N0FY3eK6w0cQAyWC+qSJrxmSjmkMNP5CtZ08oUxkXz77WSwwIs31aVbbiMKVz/oB
B085x7tTXhe1Zl06NthO42saQiX/M5FwYhpwPUihLM5ggxnoNPkjlpwY2A+cK6sD
Sr86gnMB36O1FYzf0FsjX+JjIlFVTmOJcahTlrf+opV+sYA9WAQj0K2y2QO38kr0
ShVY4HAT/73HGEtU3LcdPJmQDpPjj3RUHr9oNQy0X+uvbxLAdD6Pd1RH8Tnv6xeo
EIjx52Cj0mEYYlrpyLBJEX/VxusJE9ff4srPgVKkf3S/skBv4QUoy+rrbz4ryxz4
uq7oiGEkyMjHur7M2xHhzqIZ/KEfkrhir9dyvqJZ1ZfKsvPnt1TGSp9J7nAdXnGo
V2kPB5WxWQn83p8Nn3Lnzd1XQkm1ev/CQj74WhfjC9oqPsld/Tel1sEHe0wka+DT
PDwTVTQUL6TX/3pXlcyCgUV7LB4XVabvmcFhxbAcFbegSCqKN5DBtLITeiGH1DQ6
Udc04FSc5xwIdpjaJzdWuWtm7PeBau/XevmaY5uso2QPd6n/yhKgKFTGH7e8q20M
SsnFnvzjee6vOh/3N/xfK88hY/s99hNbmEdufw/fIRewBi/DmRScHG8srzQuncIL
hyIjuFbJF0s/0OdYtdzo+37s8xS9dun1TComADoe7qmAhsJve0SIJMJpYTXAMObH
J3QG0xEztnLuEXa2PF4fPRk0u5Z+JE1YfLvFRDbw5LiL9OkSNZvDxgsqv+TcRg8w
xcRZeqNAMepR18PGnpfp2xL7QwWAK6y7pmYIRgy+qt4XJ7vnmgUDPV5+NkYXsOq0
lIqJ26C7GZWfH9gJGGXnGo4iKgwB+BVzqvjegC/nYVxmxrnyWBajpxIIHS5rcAKr
pbRWMtvYWfLgBez7cYSNwv3vhHuRqTh5GRyS5yfdKkzOT2O1XUM3/waTBpf+aqxS
opr4UJjHVfKyWjMwNDsiDLEweyNBphgASa+mBB096aM=
`protect END_PROTECTED
