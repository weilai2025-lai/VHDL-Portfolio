`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THrURmFsxRZZOHAoCPaasMK4mM0UG1zNaKSIdtZznRN29QhIo0A4jJICIGGesWuv
GVu0KoYEAuoztWITaf1W0CS2RjupF/1TPtxRqDnoHzXYs14zej4Gv7AktqIb2ghE
WSHHprheyp5F+QjteuzNXeXZd+ytkTXihoITqC4kE7Z+pYYyOZwjZ7ykkrIv9BJs
+aIY7LF7HDD7FLq9fb3NLybFka0rfapHNpU/tff9II+89G64FFB3YSjVNybWlNk1
7wou288+MIhNEtLSnZZItYjtL9iu7qy8JKW43+SBIqBVGLYxM4X6klps4Uy41m7/
sQuKmwpkptbePp2vEshwTIA3wpk8mTr6sMqZfKIkuluqiJHr80CcfIijXrO+fJP9
k3QMAeNCG4rO2QnMz9qE48sktTv+rNaKLPXPNAIY/FJJbuK7EBukKbVCjJc3YgWU
TnV30Rw68fPN81wdTTebLxX4oXBaEacLBs9K4ODQUn5DnJ/H7PrFd77Ul5W2nJuB
dUwgfxp4q0IKEDFDJI5FsEt5LgsH7iNV8fypTHB5KY4+n3W8kIl6AAcFnVHJ2f/u
1MOuPykFFNJwORqol3yImcq4b8wFHJA0QizCTCSb2QF3t7dS89gpcmnrZg0Y7VZU
xbVdJT5m2b/jfYHm3n+gsxfEf3m4a+Af3Ol5ASsNHT9+Cl6enUTZFTq2+4XMZWDF
K5IojbTL45Tfd1IN05C42POi54fww0rrxLinsNYq+L5/p3ZCWRbcVCXUdK9TxclL
VMvb6Z553/fSWrhsn1B/1RksiIG0xHJgmP2bHW7EKEfgOW3My9ntJB2ePO2K741A
BcocVxP1GwmrO7SMwL1PdqOHpqnbQL8x/xxcv3eDeboD93qzBiWYlAsIpR6wSvHO
6ciNuP4feMpheZ+3UGfBhJPFzDcm0BveNICLJL2OgiPDBdf62/7SzGqGE3+9O2DU
0OWxixCTQYhLa6EHaK9MaELa4FNOkXU3YANflW4/cl6gmlnYDvE8u8xVQEtbwqW4
c0p3F1zUDbc9By3Xw95dJrQyaY1g1OronZCOttM+LO+AB3j96WWUiAS/518AXUBC
7/V+W/8scSGyS1VFYsEvlViuoWy5s6/reBMf0TTZZf3KUzIAtf+R5j0ENZPU63/d
HwZ6NJtUXI6aFRmijjOpVYVOvRAZ26fcq8Uz3oE1g7gNzoiHbNOC0/z0AxTfyqez
Ooy3hS8euWAytEML79foi1mBI4U3EYvMHmqHO82A8DKPZMpytSVH0lMa7Deqdj34
jZIIfW/RZYWh9qd52SRXK3mI1c4y2Mbo5ArlGHXNF5jNX1Vf4ddtryIEtLZODuD+
MKddb7p7/KMU9a1f6scQVeayPRgbO9wS5hWxAcun1h10YGwRW/6qDO/aGQjovKkj
oGpfW+SK9jWwWsn+yzX03L8RKlRFO8LmtG0U14vkX/frVoV4P89C9a+/zmqLac0x
5Q7BuYl5Wlh1EhzYFdCnZhIN5NzhlzXGlbnKTNoR9/i1tYZr5/ZUqvlvDf2m3nwh
5lKrfFe6xmCTQ3Qbh7uLZ7Jae9l335qtSO52o1IOUWXm/D4BD8xhO7jK8PVKEE3j
8ZkcFqPegZoS0LJEr+5aOPbrnM2DxxRB/hnh/dyM3wLcmjLwsRaB150UYLwYOZFY
GNiY50qOw/bwRxZ/t0IJVpPGUdOqJtklRRrWI253q/PJ3oe0lClzd9eoCLXJBy4Q
D8Q12QdvB+vlzBKTaIdZhuvTjCqPp4NJINT9tW9pD1FHLCxQao2ZtW+fV/R6ogxi
hKmyHPqLxc6kkN3MYK6O8qBnMh2MxkgDtsv2PToM25DcH9UYZ7ZqqoPTVAOovmyF
4SBxACCQaU/akNQqdId7wkOSP1vC1V7WilbZbxy2QuLubTfhFGp75JCbrGWeGwJM
RqUaZuiG29NXRsqlrYYh6R4LJwHKbEvrHIMptaEJ4SLb8d9PWoLGIPy3LqXCcU7n
VjXjMozWk4Sxwrq5WaZn1VPG4VGd5iBieiAjkFDc41Cxx9gIyZ0zJBUR/hoaBWgL
VYlebgWIhynKZBBKVsu50YSEWf7trT5ASSOGF/dtXeLeA1VXFKOO+UasJuTBBpH1
N9JetXs7fEyw655UiOo2YDz3iJfNJMD/8PZi8bhCQgqHsCtyMc6eKPzr5ESXODTi
Igmw+X1YKqe8yHZEkLSeKGXnKU2Nrr+dm5mcJ4Y2dUfd3EeGvO4yxdKnqesQi8n6
v4tdLRP1GjbN2/U0tqktBjhL+kAOYz01sXDonLrlkAcQfqul+yB9UwBEC1UrSBDn
penIu7c7r3hjnit6uWgFTscqzj7N239DBmJiG34Tf4MO2wd+WBiKzqdxv3UH4361
ggjbhGXwpNk767j9HxJBM2GylU76b/E18PJiB7bWWnZZaX7JCXpuFvljE3swH6L1
cCK2bAFQeSs20G85/fX9gA8NOftDm4irHHJrTqCyuwdj277VwrpoNrkfDPvXHKKB
0qeIST/+dfq/BHtgot5kg37bHJRnSdySN8kaE3jIABaCdNgBW7uFN2O7a62XBlPN
9m/fCvLrDVTmtgN1tDPV3//ctv0db0Y8R5yOFq8m1M7v7PavAkiMzPfK9SMW08IV
vAGV8iDcGHXZj1TQ+na4bsqbi1E12vdp+c82OModPqGooU2F1xTQa049TcrNkPKF
kCO/7PQuSjEmYy2Bx/cghglwo+tqFKyYN7kAWQ2A5ptrKAhbL6lUtj9qlDzwZ5C7
AB+DiQoyEM74HKd2bQDYBgm7CwuQPPNriBx96qvRfV8zMV818XiBWDjOe+d+amgw
QHNsynIrDHLiI+TO3fgEzopIhS+kYP5ViwJABTD1Y8mK14NAFrAN+FKRkStDo2gF
BFD4IPh10eRK4BE+qvhy+ZGlcPfQqtQkjTYhQWK3ZZzom5qdl5JYAyC7oh/Zce5E
yt0Ujg/EODa3rEPrpi6an2LjK+WN34mMrPxg7IdNZBz6h8xP8zQupeqr3tpsLO4i
qCJwYVbeAP+p7I7a5cWjg1/F+xED0FFLGSHn95btDGnZ5KNOQMSnE02XNSHpJgts
b9nN2NHds+d6AZkV/yje36E7Qop4j4AZ+3XQu1YdZ3+lmh+sEi779ZIhkjuidNz5
CabQMG8uSUFecGdsKx+j4mTGzmhtFpcn+6f0z1Dm9orjJL5mXEPy8jvWz6f4MroU
qfG+TQ4pxvX6a9aeuvsUXxzBYoHqBdGEs9hJgw4SY6VUz2CpuSSp6voJY1T1344J
mOXwmrL5GCxeV/ciP0yEEyKvGRWOtufaL5+0hy+Bo+qPzNSgy8rok5UjP+2lvV0F
9ERAoGCIg6AiFFOb2M1uY8dr7MyDK9Qtzzs0DSlwHSudBicebTPjN1lc3tA7GARw
ZF0aMODezU39dM+B3X3XrTrZJHQD242dMYaEva9B7YXR54GO5fBVk0OpRXaIvcCo
ch0SawXIy/wgOPk4jBaWAe4F2j4iUJo4B+U7duou/EwqnH47ZrhrYWIM36G1ocSr
LVeSGs1h0dwLj2GulNT8hhwd3nIJws+GmlUxNnHJhfTo5DW3kWobSZOcOLE4BvwQ
6Yr2Gz7ZacJup7nzOzrL9++XcJnA1P9GPyrG86ioQHOM6LibGHQtQcPmL2SL74Qk
IUIKzBZOBQPzfMmNAFdQxFxVEQLPPvzT7C4ViG/hdoQcGd+m9OlMezqXkU65czmK
sl1nbLegBqSBrweNlIgJkweVM2vhhRkoT9nKn/2hRd9Wm4xj50apICa5ueQsLJm9
ESunDJNdNdUSfSweG9yJKumz6Mb+jQpsEeBtV67QXsgjLXsGwzri5Tko8tI2VwRj
F5f3LGryQ3DkbKLy7SxHKOQOyGZH+HNkwkWkwu5tLccgtUfYTXOhi1C9MpfW1Jd7
fF/A2QHydT/f4u63Joi0PnTx8WJMfVeTRZtC2ukNm/h059VsflJdWT5uJeU9cvWY
E0T5xJd6owgWuEqlQLP+1KsALtLXl4i3lca9BEUN1jwBX5Nn7/XdJdCXyXK8RNDy
rOzGy3yJel0iTM5ecdeRTilfTpqD/ox/UHjWGTvOKGIhw7c3lfQSQPIsoH7CQvQN
DMu7Rf6/DnqEojBrKQRDpRgiZ4tS/PO1lZGMONF5qLfMCRSGKdHXMjfY9ml/hqx/
FQJzWcp6vtdHPmB5UFtV40Hve7ACdXDr1n5c+1bnKbot7JA1bUzFhTEKqmELlN7U
jCPz7mgMN+nmBpPzvqojfXcs8MV5zXxFtfXeinQ45kSQtGe22tnX59rusykdsCIN
vss5BOB2MCAqvFu1B7LsJmquyGT18Ck1ELkJSKa8yhcbhMbGmSBZmJPDGqefIOB9
kI7ij4v/V+ISh1yAJDTqJqwSGt5mExJxvZaN1RfZaIB8ZIUOAUn220mQUtTI3KfX
H1P7WyrUhEmez0mMuXeDwzNd5CfdoK0SsG4mUAgMtRaxeLJfvlMxT6/s9bRbUjp8
4rxTkgOld5JPg7xX6mmk4ZlEzAH0kx84J+2NrMsYes+R3snJyYwMdP9Uneb7tMq+
jVDQXLo6tsfexpDKVxRDlF1Pa31Kf4PFaScHpfrlQP+6PfwgiuLZ2mO6t2VwoKpI
TqzmDdkRlEnWmxsofJbFuxXo+Mh3PcIrlDSh0+q0OKJ6IQYENQw6Pgs3tR+AGO/p
H7EHS5o21ghiXebo6PFna/HDFa/78qqVaIYVYksvMJAny7sEn+stxifKt7PhdzDb
yxAj/FubI/o/VosF2qqy53S2svFAo643pJv4XB2qOG1Ag10KMvhR/c2ZnhD87DIX
PchfIQa5MpWs/n620lVpvny8lkPOtHqXVUlMIEF8kfXi8lb4h5TYzP1kx0XaO8Jc
lFOj6nYmZLhp36w39qLEUSJNPol0vnGlH9XX6hr1dDeJ0Z47ppCm/Dll32rpBBl4
H8MwDp+ZufCXb2myZA7wDcP+mB49FHRFrgZUjq3Z262TWeq/egNDJaz6J7pcPVqP
bgiPs/ZfRbXhcn+s7BH4jo5Swc6ouaa+F5Ii4dHxkPPrk2Vks9VLkToO4c51JSW/
UFCPzmx0bqu8ictEoVGv3G+a9WuN20kOVrmQTTCBJTfiLbpbp7HpIn+cpOqkrGde
tRdJCSqS1+z8m+2o3VYbqCigCGTMD5xRI1JUt1hTchPbW6/UfIJK63aO22Z8w+8y
0EhRv9diZvzlJM4mnosMD0f6TARmgYIQdWLR9uhrV55frdvR3Zp7z3jTD8Q+SFhZ
OWMeHfUkjMyJ4jT54rVdqpDRikFgJm4j+J87axAeBbwJ36tlwprwyb8eUmYDolhW
euZdO/lrw1zm0feLQouXbkEa9OWJAVmEZYSP9Ac1sRFH3RCQPgC3B2eIguWJaEDs
kgr4Db41UYobqvMpavLnvYMpnndIKObI3SczyPNAATCG1hXuCnRdl5D1BEoc5VD7
ZtlZDDL0IRptrvUAqA8RW9DsTvdSf3oAY7V1tE1v6BFboJ6qy7F67261WD/zTx49
6xVxW9SH5/1UHNAaCeBhWFBkD7sK6UFdkJrFJVhooXZiTQ2bdfkh72gAKz7EFy53
JzwsqVdcfrzBXDIoYtc9xoRTXBI25Cem/xOEEeyPLatay9Ov2kcl7mfbioMtIQl1
xcG4wTFuDs7k1vUCo1CSTLBGphJWcQSuaqYjzB8qFj3lYbY3MoB38m8PmXcb67on
x8g84pwXhFpuIT0M8xSY3nZDFmTpq05hefLlfJDaXETtf/ocmB//Cafz5kmDeKgN
jdBLy+wOIzqcmj2Z+O0Zox1YKAJtc4ZYXZy2x9rHTZwvp5FkGBDod0RLjcuIU511
rLijq2ibwc3vkZNXypL04HawNHJEwwoa5BwtYN0ygqT3OD+n5nA3SoL4EzCU3+sU
taIcIBNlBr7hvC4vptPKo51I3iEAR/Or0Fm3f09KwizqysOshwd1VszeNZpUGXIJ
urmLKNDc1lmsD4ubcr5i4p+yZLeyHWlo5LwVF7fH08F53U0I9CSBRaiCUVN3EGo/
qkgcF2Z6MCT15cQiU3k7jI5Gek8YGh6zw6arOWgUFd+Br5Ani2Odj9hGKlo01kYW
CvPtBCS77Xui9eqgQ9P4z8oqrqxUkZx9elz+5jSGBNAun2owMoaCKpssxxFsRpu4
/7ahCC3WZMVCtESGapUh25jMmk3uPyok+BXzudWhRoQj4lg3bj1ForAP2HmAlNlN
Xpn9gG6HIXGGKDkC7rMuXxff8s2BCE/3uiMXlE/GPiZgxhFAX3N3SZJGq/zE9ai8
rf5vZhCrEs+ohOdvEEZhjaxeAi2F7kHwO8Se4R4doTKXAzz50UccqbPefT3ahbDh
927XKrKhP2Ia99zXkQLjMli5CMOJeBpNwyjKcB6BKGS493Dl9vG/PJJ26F+eKHnN
duEtyWs/nW3llZcZbGf+uCggvyxcvBNdsD4a6g0BquRzUqWsZKn5l8gcsmld3zRH
RgUqUbKqYrffx4kSZjNgHEXmDb4GO99qYBx6UaF4iGqJ5+S1wD2KiF9YUM4KsVwf
1t68rfIdxuD6pYTmHWuQQ5gxKxmUZ9SWgj19lF0QTdpAf1IupicdLgGxAvDmBfRw
d2Ulg3P1UMzWxS1qRhNKY9Nv1YIZS57yjQngYt8uU0wExnyn+bKqL4a7Xaz/dZ/Z
VNnRKn0t0DNfpvRfpeUl0sDA0MxJFeKfpDehEttoGoDs1AJypnJ+QSpHG+zfckNC
BJDzy+VrDDwDvDS5DFOIgVoIvop9cXveIy4rSVLAMb5V9wb/g691T4to9FjGUfyM
yju79HOt49PJK8MNxST+Jxpikqwy2+XisQwv0pP5TQUp+6styynGRjY5/fH7MvdX
flMZrAGVt2Cv4Ze20H7sKfJe/cRsTHDlgowNK21bHP0TJw2ZHNEDCqSEHqXZTHZ2
tAvhcpFWrlklQi2FH6B4ttg8NV+FIjeoPc2I+VGKavJmWSE6+1WaBP1Mod8yk/kM
vo7jaXC+r9CN24uVj5aEeCS4pqgR5evtwBe+5ZNpU8mAge6hZqfbsy7qFivVoYRa
hRRTablgppRtZOXUezEmqZoMmxSKbqfKTYMW0nWg90E2GxqrcfgIVYGhqBPnszCc
LMIrLDojDKeeaTHYXt1RO2GjuiM4p0HvhUUDAiZgFz/NILSvbqisUUNY4LYnUsaH
UGP0XKTNKLEwrstRySCBEvsA0LZdQ95WFadBGPwlx5lF8xFhYyE9m17Z9l8ytcZz
u+P/HysE40l0BPDT7T9RyfEAxUEADKmOld4KhZZv5V1fhbM4LxrPS3ylnxIfFK9W
ircQyXEDXMqUpuI7SFCvTFb6Z5aGjTnB0wAv4C9dSGzEMPkWHOJyk+Jsd0u+Jmmy
oBEr8QW3ZH8fTQx77lIOMYHzufYCCCH0q5uZV7rVs4eaw+YD8KR47g+uoGvgEpxf
C2O92yeD6TYNP6GDSeZMR2/dov3c/rHhAiAJUxHjKv6obnL0kOMSb+StN/ZQfvlW
Osa02BZ4CLKLQ9e2mPyrGiDZGLVGpYUCbof0OwsrhyV22iNgTQUKAIX+qSFL8XEv
YGKKbJo4S8e+7N96vn9m8rHTvMW3RzC1xPGXxKyzrDng/7TlLv1WcQdoT60Wu4k5
vcd+2F8FT36tdmGa44nxOdKmE5XrvV8zU03NCQPyDr6siYwG13eWceMtDbApUl0E
XccIsUtt1ZfCBABZtvrfchCEjILIZ5/YD0Fmdg9Ttxmtmz5n9eCFmb87iuuowtfU
eKxbE4f7FkXc3n86RAd+GNpjJue2WV65Ph9D+QWkh/a1dWJF+ZVSNKoB6B61fZCN
fgl5wV6ewzaNswTdF3KgYWeIzAmBlb4mlTE/8EioqMaKk/tIt9cN38VAHqRxzTxh
S2gnHfA3nWuNYLY/3cCDGvJ2q+L0U7C/tIRM2vNnTe4TTMa3b/PF2LUarzL8rUhz
OadQ1SZOVbpscyfV2O6w+bz4e+d4lPRGUJOr0LzefR+dy0JdNdz2lDxIs2EnzMNl
DC4aOPWjyjMJRGQvxt3e1rmkQeRR/LyaFHMo7otsLYX8vD5MbqaGxAmsK3pU77K3
x9y5crMZyrbJcmnawF8rsexROkLGxd7V7E5umA54DK/oJU7lzuSsJfLECGSNaYbS
C4Ce2pm3tTfvpTotgKYI47u7+cFjCQcPnhg0cJkJkKusEtOK20dUjD76egHsWWKn
Myrs1QNSyr+Q68a689qMLs2CeLDuz5pMbcm7mfTBO4GzUPFQr9zZBqtWEQgaews3
bJuNj8HwphQQBT6UL8eNDuZunTlf4lK/YZ5PdQMcqOQerM+t1fZ24JDNbgfggT/G
YykThwJazAYgccPlduIsHEnC1a+6npWfsDJk3n/EZs0ts0PK0WewupwYPqr7imGv
b3m3iuNc4wnms6o5Qr0mmy0CEfLOglUexzePtcZLC0XpqTz/k5boz6en3ujidhoG
HtAQ5YjyL078lgqFM0qyg2l7t5cRDNlT3Ri7vPnOPSvvgDh6cZOcThMObfBsRRLs
6HAj0uvmBxeXnpc6nn/Ub0SUgOY2/fM+1QwdhPd06bkDPU8kaa+KVulI7Ju7H0L5
1va5X8juNfxMfSdolDqCYz8trYUZ1r0fFIl0XkLon7yxX/+YF+BITVAWfZpi81N3
HTNKvki3fhWIS2IUR/EzlBfNpmpfXY12oqrsv15AtS0xVx62DQ3ZvMUnD2mlkjdZ
6DwwVthmzA6Uk4K5M3zoJ7B+bvK0QfiMkEa/wzIw2/r2xuJWTBzrPd2IAAvacBri
VwVb62QJDUbBcjfcGHVjl5fWt8Q0rVPeYksJBhl34uh5a3Ttw2IhDlARWNKT+503
2waRFutIhqH+qmgLaEbE6fO5u7/l0/IWnAU+jZE6mnSj2wkMLgCGDE8PJuYaUAk7
8NImZAa7es8DqejbQkagmBrzsAe6h/CzJ2m+O9LwSBX7LQAigwKEIK7CEpJeULw1
9XLiyQVTjs4lTorNVZUUqYXYkvv/KrxF0BBY6zV0v6gp1OpIFC3AmNy/jvPJd1Y+
NiryRiS2jWbXr6rB6eNLww==
`protect END_PROTECTED
