`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ak7bqCHWRPTaIVy1LgKnhtoeW5q/V/KRU9MR5IGozeiPb3Hoadf0E9uvX37CEDjS
HNhrJ0lbHqbjoebr2PpeDhDjs2E7KXcnCGlTf8hT6tLsikrmSwTWssYhMOdl4GFn
zMCR1q9ThHk6w+W0FqvbOcYEej2JAUrl5SMZikzIscRSGKpp6BdWG/B+fA2KrN1M
//+NEIWqVKLzmTeOojEPOHDLwwfYysnK+tlG1p0iZdC5Uic1n1fFljTkLBugN2Lm
+Hc9zzushwXfiBCRMjHxX+q8y7BfvOZ0FlVEUX9vMGsA8CFCJT45dprkQHjjON0v
SEZUQJPfGkIGvJkz1MCH2h2cpvQKrmxqe9FpNgy2ZYGU0rtw7W+iRrGBuVGSWgEN
rjna+dGQZ67xz1c2iES/xQzjDR+4sGj22da0BfYARfqMkLPMX8FHnl70KtVleXAr
07kM+vjeT+ngdeZe0yhBnMYu8tqxjgFIPmAi5f6o/CD/QwjowKjyD/TJ5+LbUdGq
TKqT8JCq5MSdaeScm8NWVL+4EtbKy2GTtnk6aW2pDZqYFCvI1atNoui5DQGXZmTq
tVwys/rEJXqVghnEPRpRx1ZZcq/qFQx1X7T21hHjVjUYyjgcOo1GLwKrRPEE9BvA
aIDj/gf87U6t3VUdvwLMB+1RPRh2CO2NTCmjS8/OM2DssNnIhC99Gu96IUZnd1wL
4HFD7iDwn7BLwc9u7wHkQrLH5xRxlAfYwhbolaU4nCUASqveP9hSPngDgStvZ3IK
jpJQZOpwfNx8PeE/Uz9H/YPDz2aPVND5LCFSYOxJEmG7Ry8mtfldiIqd+DPp6FLf
8XFlFNNhxxi63aMIq+O2oqO9hLQfl/A8a1EMy0pQQ4Aa8WVaVp8Wi9OosJP3sNDm
CF++gQTxGMhDnOA/IF9KK7nhLMpyTYhARVX5kCBVjgWkUoVLj/rpMJ/h4sqjk3cE
JtxASGZ4nA+jeN8jSrMjJ8s+VLcdnNheR7pXcYuQnpTaCpMmO3AW8hoiH8b0jS/9
ivIMIc0HyVNwgUNwDRDVC+zpCJ3yS7Q5r/7QZik/fKikAbk0adWrUAsSuv7cBItG
QXlRPAn3BvUWcQFrGHdjNISUtn5OiOtJyVQp2kK+JGsTXvVJrXu8B0JuFhzYkr2e
LZbsuvYQ08cMkQxdzU7rOIJ7aMgLCRV7JLhR0G2MDErCgup9ORmjpyT/yqpmzLTW
N/7Y8occxvZT4Q5j08ILkfA1jhiRVHz0NgFaQkqTTKUl8k5Ay5Nx4/8WEE/Y/EjV
wCtHIknpUAzvdTTwRJP1iuab6SHiiWsv2reKxR8BTj5dHLNJWzLjqDrGp/IlnCJX
8Bzdds0mJLed+9anVF8/cNVwEPSUwMwJWMqpNy8rHz2FVMklBeFKa5ZBGWuUQ+86
TU5YSFJQhznbld3UF6fA5anMF5Srb6UndrGa/mZkpDuRLABHvvU9Anky57BIgaIf
/R0eGd1wAU4cdpydHsj6zmy/Y8ommdZzNEJVWmMu9kHvmGkvrTLBIM6LkUOZ0cz2
OzBfZ1pC3GYM0zN9KiN7mxFGwhC86Yz2/Bl1n/cYoymlmrrN9oM9EqMXnm51o/ED
jxfwwy+pDdRKD39oK1jTNI00uuAdWjdlcUruC1Liiyo+P5nfxMD6QftTLDJLZFZb
RF8loXhqDGMoWoCxHylLXDNVXF4RZ/1G/iyb4JcUwo/90lliiLXXia73m/OWZ2bY
liUF6TZfy2T1rFQGLZGSkUYG1MAFx/QcXU/H2yixxUNcpbH6/Dghzlfu8+sbmhwB
63LuJuhWG3iCN+rZ0jnw6w91lmRy8uBkyfXl2C343bL6AthUHJkN9mb/Aa/NSxDI
Et6l3UMmkcQkCE6p3HXumhvuoFx4iDxgXfDAjNja1menWHRyHgs2Hc4ppNwy8c27
aalPcQ42mVGMTzg7YvkU4dPlLX8AGCpfIwAhFQWvy8NUyZo6+JOFLpRdXxeuqUZI
wPFmL+GiIRijZbvmoejpygK280hs6dyAIP8lvY4GIpcpPt27+NGbRkmYgWdf7rko
LkgieDf4ye0MnXt04aeNqkRL+PuKJ8Da2SVzXiqpByyi45AWnN0rz2pLmU4Vjc81
9GnyftDioMwIpRVSPovLeZ3vWW6wrFAv4BmCmfAnbZ4pfBqwQDT8GCEMOc2VmQvU
QbEysGeJm2mYj8VRnKvk6t7cA0yP66gBO1iERtWg3q3wU9/yv2jXpnZw3opjEZ50
LAR3xnx6LeIXFhfCCYWQZXRBEQ8PBpLmghVq3cpQvl0XJ0w/w/L0X0jbaz4VkL95
jqs6hBUVf7c8ZT2Zj9ruqZ9dESZ9lRRUOzfgYywGWgkTD2TND12VUzWiKn4pppDn
G/5LMzwOg8Cgpzc8SsQ40L5Tgl1aEN9E3htMqv4Pgvom3cgh23LP4HlvtqLyDYyg
vWpP23d8ubJi1gQmeW9XMp1Ghicg1vtSlP3MhFvAc0ocPgGh8qUz9X4vev1IIW2v
t13TTeQgz20LogF+4Q78ngIEzr/s3QTOlZbQVAnvKnbVvk5Bn4pMvczUNB2crhg6
yB8MredBs+l2XRMJwpiXYSWQE8vPyRJ0OGffzid8Ct/nw645/g8CCF6dXJpPIDdp
3mJexB4iXz2wRi5CscqN8/+d3zkUJjItjpTzfollRPKKizA/aL768d96Ubx32Uty
E6BcxS5bkXN71YO2Nj8hwbRRuR1cdYsZiKByMyqw5RcRZut+NjlA3yVp71DoV/iy
SgHddls9SkYKnbuxVnvXgyDIgkdm00bS1gOflggJBdWxe+eD2s6cwOdZnZ6XMgnI
2xV32CLWL2v2ZIg0LwFO5n4o8YHAp1EAb3VtaXzz6TJ6gVHUgDfj2lbY0yGgmYKp
edAm708dbZzNG9V2+VKFceQIfyLT1mEkE2Rm8GRiK2SbIBDxfsdaCiZP4+ieytKK
MEx8QmjvQ2tW4Zq14zyaao1FOWXvvI2wgMGfkFxPMBZxH31YQ+2e2DUZ0590r0Py
w+a2vNlcHAryBeZ+BUG5t9TVarfGQZW9hH+NoU1wMs8+SE2803eLNsjYt5P4bzPc
/u1w0aj+S3RsXP3Jp5/ZqqD9W0dNjLEbR+jZeow2LAfjUl7hUZkxF4P/Io6Ti7/a
zluN10pEr5SImtHx4X1r7KtvRH/fsm/oy4+F4m3+VT/mgAYuBGeV2E3AewSnRpmS
jzqpkecBuJRQacU65yMaiBFWMJ6yQF5p9d49xR+rKeW+HoPsOqPfKNX9RGDjK3Hs
PmbOA7SuZfpEwqokMjoav8SonqYWw8EK9D6osRluIUSjhTxbanujKTgA08KhC8eX
3N8zYHuw8OonTlxUPQFEqOsBFIlFsSN05DLbELKAq4Ljbup0WgAsqIQjy+LDclCJ
NPYC7Dtcx5jMvkjCN09gOFYPEsBrjiR3S6tuLKOEh9xZkFAq4ToYMofc3hlnWEbP
aYJMS/Vk3+nV209XvfDR7khQ1YF5RSGZCPTF/02qk2iPWAZp25MTGd73AdhJXMV9
BrLrKykVhI0BsioP1OUT/zW50N3zlKmSn3jTx6HTJcJk4E6v0Ijov2rBUiAy+y80
pz6zcY/3TWCUvurbKQFnL+OE/VuDxAELJUWfYdIKBqQCLHhkEFleqDjr5wc9O1B3
s3DPunhPM6tFKo/1MjfSJDdtMppKlFpEEcmm2BISiSYolKdS0MoNR4rbldL3zZ4L
tqBp8IXj5mCzaLoHdtA9cSA8j6MC7g8dMjpQ8h8EiWby00kc0hNxwgbmGYD+pypO
FRcoJ+JxBRv9oYwNMkFUbcN5FY6iCLgMpLGUkY6UixzyBePemyU9uS1sWEfDq0Iu
4yRUbcWOjjZAWCZXkRWLx+1kswy1coqIneFjw98N8LRAR8c2sUXSXDA++RGzuhTV
IuBNfmeqqy7dvuHtQ+f+Qb7jNBPmuX4qVvak07VXD1r7Ffzr9Ab4lMiNhgf5q3Pb
iJto2kJQXKewvjgDwLVBbIKS4Az9mCPDoRcbqGDdBqQKCztq4t2QL6eLnPls/GQ5
j2jCbApoF/jb9QKr1/t+ReKe0eZ1qA4iyiSNK2ns2Xn0VgOE+kzzHNO8UL7BjbV6
KMZMWVFGP28jNARQwThT163IG9VVlCQCEtai0Ylkw2dw2erJLwhKfqYhtnaN4qLO
jnVAlWeEOyFUU7uTvQ5BWUFBWc83xNcSc8VknU4C+M2RI7fgutSiX2pALqbgxpZL
i0o6JSHqVe1Xe6dZ8ZmKButCs+K66CFin7/ModL1YC9KIGt53BxVPHZ5BtzuSGGW
zuPVN/l5a3TxOOM6OFB0fHC8Hbkes67rhTQG72cIgr2NnYrBPUxZiLdymaZUSrok
mJTxVXJCvtVWY/2dXIfSL/D9U1rw+Q6+iDP424ER+oyA68OSCAQPleZs8FrGSzll
KMxSPXuxKZU+dL3cCKkrScFarNsNkSa6EnghusKorbt2HtEhilqFXWF9FMveWGVj
wnnfIvUwxYKA0BdP5RX0TvZ+GvdGkgoXPHPi98FLBnEF94WWANdvaDQ0mAI1aZMS
442QTmJmcSuYIo8/0dWQ3DNzsNIj6sbs/2wdwz56Ncpdw1vr3F6JOBBGoqijGykq
AHm0iOAFXr0vu+Dbj4WLvAg5F14+jcYl5hAxfJMph04MucpkIQBGe+2++uop+Mmw
Zk3cIYsRf/r549dwBkc2IX3O36DppLWmjQtFuXle9Ac6z3mcvrKEizAsUQFN1ADh
Me8grLZbFbNsyygLyZQGE959QRy/sN61TlVYj3X+H62wgMOeOP+dB0cmE1ba7zQU
nY/MhEPq7ciTSJj66ZtZOJmoC+WdGz4+LFR9EYr2QbRCjI5EuSnwoYCM0VWNOzX6
aS+Cq4hP/YSFnPF1Kw/hBnJdfAGXziErtJfWUza/S5iQliCdJxd392UuSGxm6AIs
YuhlRAyDd6aUjY+mvwN0bF5icQfxpYSXHeQn+CN36AA8X5gbnjGpYKslwPt0dLo7
+Pk3+Ldpzu/v6gs9E6aLmNGu+loHz/wlL+G8jfRO56YwxaQQqKWyYdWP10w9EGI6
gpZGtZgEr0YJBTh54ipYr+T0IK+IctJBW2th2/vg1OiRfkAhnmV7wpx/5qU/WI64
I5ffE+aj5PB/coW7lK8dRvHpjTi6CZ5uI6jWDOTgJr8P/yKVFfoin723ZC64Krn3
XEsSS/eJCs8yiUX8TfWFyWnQx+oxgXFAa9v2vL6f2HMmyaSfWKUMyx84PR0oJNP2
ohcdRHd98AarcyopppM2qkF80dq4hfbGmqK6YNdXVj4iK486/dtvw2I5SQPCGqBw
o881hfILGVAa9ZCjzVKxYcbyPAli24rnIkka/henaa39Yt4RHzDkHcAZqKF+d6Xz
AyOcTsiWrO1kiw5pLZpQT9Y+Sx6lCpPsiwuMPQNHn0xl9hy4EB7DiMbMGECIpsqp
3GXh00DPtooaQpPSTqtDZH2vyCPYCqaJibSRTgVg3aUCKjDHGyizuYOZK69SIOlT
XnrzJ7dNJqkXcg2vElsf4dOriSEuyMmM0A6R6O1q+76XXaHagQBlEExfc2IhMirR
iLqXYSBd8CnFAF1g2owyskMYlDvV9T3XMCzz6khmKHeMbYB7aMuxuOtLEL/WNLgR
kN9EAeiYUWu5A68QwKO9UH4PzVyKPHTpH/8vZc8HiuX/7DZp4jVEgDJ1F/v7nbIW
9lFHIQGV0dk5Im4OIx3KQEgco88zVrXshcCZICIj2T/U12FmDWwyR0LCxxgoEqTV
cRjaigwb2ASL55zHuWEM20daI04hOxSP6qUw0rU8PPDyArfrEIStBB7ym5+Ojcpb
nes6cbVJ+Nh7IU1pWvJR0ms5pLD1oZ66BZiIax4UU41emAXPXy07PPd/meB0Glq2
dVprhIdM1MwmcWgUPyTGmNJbZejce6BxTQB+IPwSRCuEsLJvv8Y1JrQWzLBDAkvY
pJmXGJqaF8MziByjQvri3ebi9OxwBA0s+GQUXNOlE7R1/H6fKn2dfSPXWslcZH/l
`protect END_PROTECTED
