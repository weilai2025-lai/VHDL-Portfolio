`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8US5Ev3rOA25Npm12vq7GbwKP1/znL1+WJQXATYHltUpZXVv/nnHleKlm/2ag83l
8vXeXOUrpYMj5jSPkx7dhZG567flRTUn8IcEvQGLVJWxZZvSCReK+TRc/Qt8RUHp
XD2JKi191PuGtw/Vq6JhBNXSYfMEJ/sYq6cMZSA564qhARndQyeefrXBk05E8YhX
X0rwTdAEnuwYOdrp+yFOR6hIpqpDV8vbFjWy3oWdhiXv80f2LXVuyWw5reNqn629
ongzWNL+SsoIYROeGUlGyoAVOl5op4tfhPJoxfZNSaerVWvycz87DokEeMWyNjND
NVAYLHs6lrRCsA5FL98+yMC2UqpVHjAMDrIiOWB6FWr59uwMyzzlWxe7k8+LX3QV
GAejcDwVn/+rx6mD4uBKuNjLY2zWAQZlxxLPnHdIyL12GgKVbuicU8RaXM+4Riu7
0Bg+8eqbwXQFRwzvVm8m5tgvJgbVt93OdvWmBffLy0B4eQPwxTjrP3wdxn8ohIj5
o+dbeAdj9/1OUUm1zWw66k4VK3w6SQpU0b78ljJr/oolMANzlATFrnBe08X6VCDX
kli/B6tbecShbvQr8MOKrNIAL8M/q48E5KX9tNdD/XN0j+GUP9lz30HHwCRDBJnM
IciCLs3GzBwqMP+ZRWGDt2NVxaGzPsEa/aMqk0vsAW06366rmWMi/RWKXzv9RbeF
KVKIkDBdtBLyXQxe0jgF01B9BQ6dMhFn2pagF9Pegt56ZtxxyplN9FKHc4UZLaTy
SAeX60tZeMMVNMOWxoBSf/WWspsYQM3f+l1s7ad2WKxjvW6gU06eYzNEWI9PpqUD
he2+Jzxnh80p89ilrCJVokXyJma14b3DTpOfy9LHqv8GUP5hiFrPdvU1riafPZMK
gFwcdzRYymPJ/76LMQCjdV3po9H6Gjo4JE4vFzuHK3NOiercC3aZfjCP0O5Kf+b0
Xf5X8CD+0dyjjx+3mWJ0aO5FN4GvZW2f7ew3Myghn+zpSTCI2yCI+hLmgOqeBd8+
9J5mK7ge+9GS/LhgviWIxkt5uHBkYbigseZLn0cfr8Tq1A4ibgOFTeaHkwIV1JsX
efTSwUInWuPHezc82wOgaNrbdhiSCIoC1IeYwPRYJ3XY5pnA+hJ2TaWT/IT3Ze6f
5DumXtagJRhufhxDmr7dGH/VyJqv5sTe4LomTuB8x2/HkCsrFPJ5SHWYM0tgBb3M
4L7TCGCrNuBDacO/JULpZPNBNej9DwYaFgN0O8NTj1OiRCcs2fwZBbdCrm9QGmW4
`protect END_PROTECTED
