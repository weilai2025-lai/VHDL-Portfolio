`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
svhkAepbhvDilkVety0rWy9YPxVhkzdDV65MROBcouuNLrbZwZXXqvhXIWA+wApE
HzzvR3Jxq52LJ79u8S70Mn+QqM+Sj2PvQt/86ldEY5bCH1jA8htHWCaljOPGfd6N
oXHhcroJCb3rWjjVyp8AemE4vU3EfCMQN/9Xgap0Gn+TPRsROtnmY/l0yOuxTpWl
S9FFZWcN6k6+yz96ORV8VOhnc0/36DwXSHWwQg0F+GONiUbZSHjqXv0HIYPySuN9
H6bVwaQLRDFitgIr5gvz1jVj42HjUbBAzvCXPSl4+kAaBKQmL8UwPr2wlx6CVMMd
ZT6A31ProKkizH9AqAgkgQQZwjhMSrTa1yaVrxs5JUt6Bpvo33IkMfezkXj+93wK
NjRGGzS21rLTwajYfGU3rJOQ9tscyIFdZAdbZ6iM85Zpmf2salV7BJgqlcqy9RpF
RiI9/AUd4Ci5thovu4Ab5xBZdpNItK6MWzmYlY2OXqCT6NJ+ZecGxOS1QEodxB55
eaIEql8c1107SLCGSRP8T6HLdmIOoD4RDTCU9lwq9Qk55KhCEZnNTWrhItv1o0lU
VP0LmpNVMPUm3UIzeQ0FhIkDUuKuRUcvA/BU5OQJfOXC2+qrJyU11yYXp1bPkLS5
rKYEeTHQfErEXSaIy3Q8FwK6GQRrXKVHE0EfwAO4p8MNwMiWCRa7xu1tnQQasX8N
HCCo2RhbBg20Ecl2pKcgcuDQBh9rSvdSGC7BBpMIskqM1RXAEA5VyCNjn43b25OZ
fWQzlDfvl/IvmFD7OTJrTZSWOGTVNqiQTYNJxIuUXplKEXskojlHPfsSk3wegU2s
iGKHzKCflF88y9Beyy0Bu3rHrfvT88klJoq2TY52WGaVMvkRTUBafKds70aqfUfd
OBlPPR4z2vTnyOgxMHfcdUB+U4Ny+iG6wD9ZXsby97dOLEXFYOKvoPnm0je3SQB7
ltbFvIjIcCqq+PqyGqwAoBiNmS1MRtyY/FDIrMeaubvRDpgHcNE8wVaNplciE+cB
bwfSXzp26v4SIdJwGEIudfYpvyOg7btz3uewQNA2OsYlS3+HzMoNeibg0dMQa77u
HNnpH/uasu7+FPHXSfrgyQ2LjKXIz9u/EeTLZPkHJz0rAXAX+tuNiMsnftB8ThXd
QMfTLyUagX6KX2WvdofO739haT37VkJjUz1+cCpl70PQC+et1bbGAYFkW2RsB3R3
wP/bjB3ZLrw7SIXj/Wy5Fyd410EPJAY4Hw5SY75b6sBJmb5dX0Ajnl+PeDBknlVN
zFszqDjl22Arw9eklMJpY95pfP9h8zMyBnZkyUj5CiYazAnC01Fz+fVSy1hvMAo0
kVvii4qYhS5k3p7Ks7i5Ywp0MQUMs8ozGGD+viZV+NLUov7weABbHrPebAEQeeIA
cgN2FPbClZeFMH4uxUtX+2P6lKwXT6MTnyptX5zhw5kK9BXSPJHyjaSiwBqgcJ5Q
DpzMMKXSn21CitJ9XVWcs39tPFBpq6NafyExdgzOvM4PKBEez9tM/GJQhJppiv/J
AZmIxVFtUon5PUd0GuoH7PgimhJYmhkCUmq+t2BbTvI9EGkm84L2CQTP02m1uX6T
0Dd2UbS3x5NuA4wXREqw+aQZwzzOPHwhwoauNkxfLGFx3pGoEKXyJjukAno+QTZB
vO9w1RLq8G4etu0MZhCdJZ5ruYCRtRC2YfBN7bb48DEKi284jFuWNBbLhlJ8d4+0
QvfV/tk09Sz3V75jLnOBD+7Vu9WzBN+Vk340IYAUdQfwJP/r2givZN0652zQWsfQ
c2vgTGAH+cPbYs9QZZln5bkvgNtPvUCzgcuhKQkNZRIRX7KYYZ/r013RHp7pWzZM
MHbrfRz2ybg+WeQUhFUGKaavm887os43pU2pH4jfSEips4uz+nIiPctBlPteJJAy
MQEBeQseB5LSlfW2YG7pBrFufonAeoHYLy0MJQiodI3G/Lq713GeziBb5qXs6wb0
G2IqvrpUsBsIXG+WWKtbm7lKxaXG68fYqc7fpev30mvpGzHwQzVn6jH2rAoCYFrg
aB0QcBqGJoWQ4APlTu/yE0tbMuUkR9002vHit7vI/+8ZjXcNY4gGODeseZOADNHa
DhhnshzaotddsdM8i+hHXH7QDCEpEZFftoamqYPVZNLdAaXVyMM68tUi9matT9kZ
HAosdh9QaPgyH2CgQtxWXg0yUEXqm01VTdvkgm7LSJgr5avUL3i/UbLwBEPeVbkZ
zwUrrasniKtuWwDhZDg7Ug9B+uIyzr5Ri25DM8P5At8WYIRuYyqEeUJmoZIFaNy+
ZVp6S4xtzNRScgW1ibH+/u81eeNJzVhtFUXok5hWPfJQxSJQarbB3YhR+i3Z+pss
2SIXq2AnM8reorofarD/3JXbisq6G/KCK6woZq1uYKuKj+XaWFcvl0+8dZCK4Mus
0qM94mMFX/Hm4GzLlGfjBxq37HjIgNro8w/egmozY101PUL5xaKrgPgUM12iG9qd
J/Qc6sf7bSJf4Fh8S3LqPAGKYrwIABmgovLJTQP1X0hlJmsLAv5oIGWhL1NlrHao
cQqpvJ+Jc8tLQV7YzhmygCqa2Ir0VLoOMbcKLS1AC8DEHFOUgRD9BSPPCrOTcn71
9bTDIKw3iESIdoLQmOWqhA5BJ1xTMwqDkmURVAdrCkDbSEHlOsIwxcNMxNahfd8/
w0dbUiMDZFuZTt/LuRMruijWotUS2QSAq9ChHK/1w+vqCRuQH0JN3aP9HRmwyhwW
/LQBa2HCDsArJtbR0MBVEae9x0RhgvKwEjMzX9Corz42PxrSpmj2+eSVvcrpeKHd
mLt4jVnnYrcob9MUt1+QA31//i212J/BO1frS4MSe29J72RUfVSc99LD4MEQOhAI
ecx9HbVClShNSJFmb/WsnHFnOlbVbLCRdHAt0Eq4HnD9P51ao+tHGhomBAzSm4Wy
ShMjd9QI8QYykJrBHsxmVMvFUOdvCOMPchiMbsCn4TxRgQZgmF3oHIw1GzVeGYvm
X4/YxIsNQiryad2KpeP0saAv7nUmFayuS3tSErjvSD1GZ1HFZHWTw+1K9w7lVJK2
JJnYNLbtqnxvbTCHLYPKE21grRD+Kj/d+MmmIbGFG914Z7H1HpzRC5h8LIpkjvmo
aoc13gp0IcbMC0H0IUFDwhdHcZyXcoIuDpUUxaaEY9qcA8dgsoftqYSPn+l847A7
hJrZCytLxAfQwOQz7sQsd3+dive5z5yuid3xXNh6V0kEwctDlFp79a1zx35wWFx7
7yA6UH/4lhiPzArFnH3OmQpihvkeH/3PpYJ9AurrJ8gQmxcDAW2S99e9CH7PvHVh
PBpSD6NO/LNDEbwhFjr9Pk/U3bgoW8yFOGBo31Tov7Bd4TAF/R4TVQLcTSsNWaCa
MaQMjla41HFfWaBm1iJSu81oBW4rndi9zzMqlKQX0vjMngV9KxyugzmEasID6k7G
LoEOUWdziKKV9D5kzAdODmsHPpvDl3gd6lOQjCgHCr0bPlyRg029WjmggDU0chgk
ilWplwdaM+DVwyzXxxgkbDRqW4nXrwzNnVFF4DL/axks827Uv/TVRATXkH3nY6Tb
jHZtzwbYC+NKKwIbmLmc1Q9ERBzgZAeIAM8efc8jgzP5YPjPiNmQjw+v5JJniOsY
T1QtvFUnjQ/IFOCMh7I3G3OskFOIxosUmsR5+FbORWxRXu1ISOYGzb6CJyL50jPD
26ile+QgmFyBk2JgByrPBFMJyYuTZkII4cpq8aHx2hCpzEgsUClIqznAJbRsBT9J
LeB8PA9ZiIo/YDeqeBZRPryjPXOETZyZFmguuyQhktMLeXnuZmiSfOmy2s0tA2zm
+hLktCBilhscZRbTKpXOHk7ysy4EnAPXcO9WJbpfzm84nF37OA4M2SpPVoqXlZIW
iJaPRlIblj0SWKa8GnPporaI28SNzQW2nZPHtI9aJhv6CbG+A26/6LvRRB9yscOz
M1/J2E8OHG+LVCcwVt8fnUmFojq3Jk76vBLEUbo1IPf5tEZTXkmQ0vDev7xjcUHX
kMinV4/NXejIKmtN4JDxSDXo8M6MZ3qjvWT0KhGqtA8me9V3/ldZeAjnIWjiW9Zg
pwZsedEEFRLCnOIe7Hi8AVP/oBrK/xM/b2VKnS50NQSktZ2rWwNV8KfYBxOGOWPp
WD6HMsndX1jpERQWOasEvsmAdshLtFfzJajeCPtbWB2Nwwsp4ulTJoUOct6K0QRX
rGH2KNVnO+qnLTp+H+bM+LvPXUl8ZPE8R3TRRgRvhY8MDo7FMcoCEjaFSGnG07jZ
JitXXdsrF2OwaB3DLBBBy4zIaVl+UIYrIk8u1UaDcVTDnxDchkdNOx7c23ZQOiLL
UsTAZWWsoYURwpqN/IXhSHdqGwCjn3f3w16ZO/2Z2+e3sjHEklFwumyNnyCGkWKI
u5QpEk2hvHWAnIIVXXTOf9lLSPBSCoOo1TEYhv0WS9RH6mFLX6gv+TcVYlssj+fT
/VWil+wKoUUOf/MITVRbSd4JX6V/pbs+Zh/VQe+v6IhnhhrW2BEMW9YV/CU/R5w3
KY0v6tgks/1MZkzEplsgBExqxZiknhHbOKdS85vXGFzBvjn+6UTlH1NRHwtxnPsc
Y5D2PoeOACtv9wawJTewgVCKn54vV8Zoy78N1qzbV9oA2w7iwVZ7hht9K9Nr6ALR
ifxIRChf8syVpFxhGaojHUehwT8xvFu93vLtwui8OMcWLpTpYNGrLhj5qe5I3OsN
Og2+qHtmK6vC/dXzQb3xYWZPuLoS+VMLABwkeTdTEHow68Xf2rVJW5EBOSW7WVCo
ruMLoCUpyQFzh2bDGheDdPiUK0HGf5VuydPJfa1ImLX92+2yt3hcawGTtYFutuNl
wWBGWkkvmje0p0TexDPzeo7uA/kLGO61ciH8My7OS3XVtOgkkGlvLd3pfADRNbi/
UfJmyj/4ao3IFsmAdRQ/4zDBumSRc/yWflC9mlMYBGy7y4NU2i+vPCsVbzOOMDMp
A0lZNAvf75mTAAy82ugg3HXXiywG6mV9tS+l5jFyOSNDjZOmbovl4faAdx0/CExS
L7IX4DdfuEO5+UCMv2hN55hoo5UpUqTiM9Dp+/Jt2zvqNPyTjOV1w+DrIFlJ9ro5
6fJ1Z6ibB2Q15ggTudGx6UyUbQXFyevZ6s3uUOBOSmIBZxvm7kH/bEuX6PcsJf6R
mR5bRHRILVhTfgX1oQBS8R9HCipB3ziM1Kg4j/j5Z1oUWsKETFd5IvH5+gNQ8GGC
Z9S9DQ7durGuWzsadgTFULdbJTNZfPS+L9A/LOrGCVhMwOhEYUMUsNFbzZwLU7Nr
iIs1ajcmbZ224rwIMJjHP/X9V1Fh60Vt+fEkXT/IxZhQhwWvzVipoeiXtVAo+ffd
vqdK8UWkYizApmx6Ku/Gvk+iPW+XnzCLKfRSEnC0+iQhuDZ7jAiWik0GUOH4Gv4m
OhvIUyF5TtuFRRwsC8K3HjQ8AjPYhQyc8yvJbQns5QtmhUS45DZeedi7jpW4hTv6
kLrANVDa2IHC48mxvs6jqd09Siyke1/evOEU7EK7bRbzZJqXLmPjT6Gkwsm/w5Cr
TU1jf8Z0gIE68cyVUD+A0App60LEHL8CU2HHKOLmBjRGoHjui4BqmZ45ODPOEUPk
MPFb1T3G+pAiBYjSxIyq/GBs+WjudEKeO/FpK0ShMUMmCbUiTvirYOC+XQzANprH
mN3Fo3oQYo38dvyIADmor89zONqQ0ucB/0b9KJkzAe+fHpkRtubRE1Uu7s7yVpDx
DAW5yOUGy+KMA/InFdLUPICuol5dtgRowiiZ55uucqRNBu9TkV/POBmOcvpy7SY9
Nwgd52/uL9LR0WJLTsrC5se8E9S3PZeVPUoJO+VLn4EaJu3qfLy2zZMKLkjQEF58
3OV1IzGN1gbTcAgiDnReuqcoE3d4u46kywVtX/eT/oDiGkbg5uXzLA32v0Xx5TOz
JxHL5Ab6xECULpOAGK5Ikpbw74HNO0C+BkWtoWH+BmWefUthelEL4r9gbuKk2lNk
F/z/M+qN1beWaR5Qw3TOM79xN/XNVGkEljn2ezkn4V+6pB4fkhd3W1e1Io2T2Vew
hh/4of0sGI4wDh6IA+HDD8EMpTfELVFVszpMVYnORPyMYyMkTA0COJ3Rbn/rY8zA
6rQT134XIDV1DlHKojxgYaEji4B/QvP0Xi+D5VinOvr/XjPfdvwn8jEKVhEqx+Ze
/90Jr+s7uM5GHDJkslsDdQyaDCqn5yNPO/d/BhX2g0DDaFgcbCfiIR/zBSfcFosI
/+h41+HvueZUr6E2J3L6YBO/JRAWMl/mJ79OjAEI0vhYiPI3ZnQad09//zLcgR9C
TeiHdAIwgXhnLgcR/vfi08Ln8UXu12hVo0+WMzk46Blhn7jlvjucZFR9/0s5J7JU
/MxwqcRCdbsVFE/l/mh6/B1XbAnhOVvM/YxgXHHidjWSrOGfMgivZHHFMcbjJ2Ao
MB90m79aI55/wlT1VkuitLUfh+Qc6SyWgsk3gOrrvxQFJv5+EfDn2JLowhTtaCBz
qvq7D/1TfHx91qUAXSOKQeKdNtgpQcqmjyqzWCE1FbR3fKHqjJ28Goa/mMcbdhJw
M+VrnwS/88SzRqPQACmAU9DNHcpSK3FulZc11tb390B88zS6IzbOGqSkxCQ46a5W
UP1aYMikOOHrnKzpsGPTnZLHNAaB3Nk9PlzXFq7S3hgjI8kplJ310TZkzTBSMhMj
iVFoXfnoLBV9OLuqnMgVdGIQ5gxN3dpSehWm5QTMck3CNe8zkSizsJcvzV7PJ2UA
YASrI5kvQ6YSr+cRSdtQBSQfTfdyVJTrWrc7DAK08wDcqL3YWdVxjtZhTB4Oj6lN
LB1s6Q1QZc5FOG5obawsj7r6ahzkoce9HavSns4UCvva65imxbVitrdKmfTDUc0X
Q25oyAUnjIv9NcMiKEaJxDlxtF1b++ED0zpzeW+S8rVsK/EQh2g4ATsvPsWJmNP/
XzQIwrtKgAQ/LXDOmzyBdjS98YS2RxLT13OFYGughhFrCzJ2SFdoyEH4MddT1XG4
I3wKvgrzaaU840B5BVs3h5CrAhsnaJCdQRSxF8Ew9N6GP4tD1NAfANlB2/mA/Hr5
e2AWPGD1s+HZT8vZERFtngKmrMmDtmYssOJP7S+EoPDcT829CRGM3tA1/kSi3nDM
0MB6mtFA5YOpAdWNAORyjarN17mbeat0lrlREIG0DhDc2Zqd6BRdk0CDqboAEF1M
x3FWfK7Xr4xL8raMKklMSzbJXdyFGFPxKg4lGTibkjrsZuR+JtV14UR2YAbb/pyv
oSj1T+jqZfWbyKKwen8vp9kPZ5U9xbtBsXDmgZK0/zHGjg2VqjywBA6j/PeO3roM
b4ZVsXyIvmt6leKFYfjrHhLw1QlhsDJ1fz6RxgZJakaZwfknnfbkCM8l+FzOhT4O
oe7YDCNxLIFSgvOu64tVu/pqWaC7Pu3CmDg2oe0rLskuiSYTY+6lUggUeN/f5WiM
VZeABtio4Gi9MlbsqGIa/Jh9T54yWNP9AppiTqQRCHwe9UVoc287YVaeMrmIxt/p
04aMSEfsstBqorM3esarWdCBcjrI3U78wJ733btXVFlYoXhEIEBqTYMwVK51GUHl
KF69SzEM93yLJShe9mB99VAV7cgKuduu9IwMIFQ9IlfPEKNhH8jYj76h3JpEE7LX
i0z7olro4NxWQIlkgG20buNXISZdHdo5+r1XpqCLPloui5H4P1pn/8xaTN7isIbY
lXCEU+C/W+/F8VYuvnaiQC4bzXlVvChyAhNsr31PLbyMjMRXMtPGJwax3nICyg0n
es9iigs4Fl/6fgKr9Skp9arDDR/wa8usVAhqndrL1vPb+IurQM2zIpBacfpksnQV
YWFwVS9udCUtzquUQjOQZbMBEqcmi722v8Y1WBeRlIYx6z1Mm+1vOBSq64iemBee
bGmmbd4TvSXR7sJCIYjBK0So4R8BA/QKouS/WYeS1laJi46E8i+H9eHtTqyfwV1u
caZ2QVYh2Rhph+0npw6Dy25eaBjnXco/XdreQhKtG/UDO2VnZaclq21FEk5RLdRJ
qGB8V4meNim1zbGjPnvur+xSLJpY4OhJge80LoUY1Vlfafq4aHZ42zs7cs9YNyUv
IVqwsLvoBKukuXgL1YVBN4dPq+Dt4sCL+Aikq6Grf+eejyzcMLu6DRDhz8dgVSE+
X4h9loDsLdIUil80ld7Odn8+8NZ4i7o5hmRRQ6yIfdG8muZiVm1GZ6UU0F0LxonX
dov6C5aN+tuqVFR9c/zzdKT5sX2ebqVmx3Wivsdv+ULEu/brjt0yJRfJPpEsGW8E
/HONryAbrDWcYuXfzLT8A2tbi1qW/aAiqj9a7J7WcsiRAOlxktxFn3dLbeD1+KBk
9Hc6pvtAGIEE/OjVTX9bnQ2kiR+UW/cP7ejCwPdx6/mtwHpwSKw+51qDyRmAR96Z
dr8WDGxkLrkI7HGav47ub9yX79X6lROnSXWxfU8gg9jAdTdbA+T69vIIS4LyX5oG
YJnc/8kInP1JDEzR8DDs1uZvPwpQil9A2OMqPWvxb5Gv51v+ZXU81dO+PkRotTeC
wu5oh0I5cmmYD179x08TqW54Sp2ud9m8+nHXHpd5DXrHc0MWiV1LoUPKMaMiH/Q+
S5yG/4wJ3AY5WALufOjI8DurJQYDyw5bCvvlklqCs7nWwCR09X5iF5yijdzmmtiU
FsFYypEzUegxxSrNtv5emI9HIF2rFHoR1aJ20fz7pXfaTA9eyLEdjq8DTZJJ/oox
Pg4n58k+ZbksITQnvApycJBrvaYI8ro9MFjjjJCnrsiRYkah6k+idzVYsgSFTeAw
RF4fwOcJVoGBRQuU68HSc/FdWcu2GbNinKdIcQBktUpcQSG3LavrPP13WJ5Uk4JL
AHkymfwW5CEYQT+ODf1Yeuf+SJgFy/fLUC3g/tPunEj3Z11nx9OT0eiDA8ShoAdO
6J5XcbaaRUzUHbMgwhfEUjTexOOjuPOMcW+qswYxT25h5pNYac233gjbGNyAVBBg
7ASyWQESxdCD6FbvHkq6XSOdy/0OiF+CSfbepkhcdw7U6bhqxLE4rrWV1b5mecq9
8ugM3ue31F22uNUdPK0Exyb415xfYYfQ3ZVQ46PbMMxBVR1S9WK2dr0rBQXcTKSG
BRj8T/JV1KAVVpT2DanB3VdM0Yr3hKyLIfVmyup39BPwRwcg2ZCCAsy3X5jGy6sb
FpS+pXZ7NGA0WsYV9HRc7qe5PBOQQ7lPXtfr2mqIOdqb0H/rD80O8dYL5+AFuMau
QS6taGVBJOrZWPOUxfICIvS/T67t5UH4XKLP6sAQiTKid550sRYMJxYYi9U73Rtz
0f3JiXrcS0/tdkDggRbHC694NmygjkiVOorH290QqEnSTON3Btr0oHwbv0n21sxG
e3NZ671HID7KdE2Da1WqIxzGMFJGJAht3mcsohJTtEqp4SsSus2l0vn/+Tk4UdkD
1/bAyYmuMRICUXejno2a2zQPnzdH4r/i2cZkFXIwNjGydx4MFlTPqiFdvWwFZ83I
KC4Yvsvs3hFm6FqvswVaYrBp1eXi/0XPu/yFoGLF3cP04FMsURp4+a/NYzjIb9/S
lwXvD+y1PFjos0Kmx/KmRXNT6P32BTjEko0tZraHnwS/HKITLB+VRaZP2BBIM3hn
o4coU6qDXLKgEQtXbYBoQ1zhnHa33j5kq0c8JYJs0LrfmvTZ8Y8Q2C/a2BgZI04s
1sg5IFa1vPIsOJVXI24x6RK6FR/bmBrRGEN9F5ymiXi10vKCe5P8KCPL8KmguEnE
7v+6ns1l0dZ+EvyDN6v5P9yrRvyYOSnW57B3cmESH54j3LWd5sO2Wap7U9iGGkfc
HF+tfX+2uYQnIDrR56GemBJh1i0hQDbbbSpTUGIZjyPuZp5hKA9ZOdtIBJqx2z7S
fgIbM1KLVCL8mxTuAys0jN3IQv1J/1+4TruJDwG6Up3yU2EcajaUaRWIq+zJKmyw
mh/kANkuJXeHWhGnnGlqbdrhNkQVKyvwJk11h6fhpGUZZwSP7i+3wFTG9IJYfG9t
T1Q3QHohVq2DIJpQWGKHqIfRLozFo+Cd8j4RPWVnc1UIFWlYOx3/N6d1q685ASsZ
iQp9FSHQXWg1TBfEUgnn4WnNvmS7K8lCxOopOVqm5pcp0yb//4e5KecVwUkfAiEi
YxEfgkQAwmigpRfILGUJP8vuGR0XfNXmLIw6FABIddw5lvA9lCQM+6BHYV9XN4cb
IEPiPsi4ga1VRINCSGNnq6XenjMKWp5r64EIdqTKOROzwMcxjYMAZeVBGcO+dRJ8
aCVPPS2ub0bIMaSzguCrtAmrmwJnVfGd7uNSjS/CJzAO9iNf8eE4/4r8eIQuLFrr
vDDXA6Ui8M5HkuN7plBpiGTyuSx2p03ghQJiuk6ALcSBYTUSrocOJMCKbYCPLUOs
B63LPKGPQETJy66q9Oytvz43sG8Lxsa6jQYqy8FD6kqxJImBo2slhGa6ONvPR+mG
yF/Wxa4lqtcTRnVkHw8Zc8JTc3zcfnViJYDs+p4veE+9YhBy6sprDLn2lWTV6Rpa
mErEDmeaC/TSzq5AKypKjlnsk3bfRrsOGkxer6E6qE9RAVMv+93RkpIDAnAPeG/v
4xqt1BMQd+7a+Q1DD37uXwLz6I8+65qLq9wmpVif0jWuufozj/SgNIHcPnx1O9ru
8tXQGTyRPcp3Iit+0/+GU1/LEHvD1kfj47ZgdKCDc2FNuUpwzLsj74dDxRjpqHW9
+stdtN5ATJgZTTLWK5eB7OsjyYGz0YZViT9f3H24AKVziOH6kvnAnafnAJaas2c8
OxIgybDovSoCTFA/JZBB+oQVQ4CIaXBQX09XXJtGKJIWNf20mBhEiuLi6ThOCBHn
Ie6UpTdRN4G7jbHM3u13mxnD1Qsmm+VuZkEhfbGf/n73znr11kz1LjuVqMnLIn04
yYA1oT7XWvLiIuvHFkrLXTUyV7Kuv5eWfQ7Me+PSFfypIeDlxo5pgAV5Mpwuf1Cw
0YmYlj2YBYE8JJkiWY5R/SjaPS+7om2zduSEprD6oe5A02tDrQ7EQHYWHANRpT5e
+o0Vp1txFhbHHa97Jm22jy+MyliOzzXebBuRsdsGL0vTaA5tOno4ZLA6mwqE67X0
IrQ6AwB+MdE2Edk+O/ynJvb3M/+iJi4aPytYQxe9wqLPthEnjx1OMQ+Yudqn7ey4
Vy+at6YarGEhV8H5PaNBViwaXfp7xyWC2Ur4e2vt4ZYx+2a+Gg6uVaeCMKNPT4MT
iveKS32GFm9znmKIUiHXzEkywe28dpC3Z+kF6ML65GrMHzF7kWcPF4DoLI/N9Uiw
80h7Cme+Uj+3zNADj5F/GEPZ6qoLac1ytAIDq6cpTII5ENfdzDHRl4HjsfNq3lz6
1UzJmC+CJ5SHHMkbG+/GXDy7fTGTIpWm+rvZOqMfLsumsv4ZqPDY6IMP5hV2512X
M0uFWXYaOEQSmZ2sOz23TUE9QCFdpXM9SI2gD3NGDbXcCHCwbyiIzPfN9U449XRW
uRnRaGSxtH+/SUUgJL6rhoY6jY6oA74JyYPatCAQTu2fJ2JVGNx8E65TA0VW/VQc
KgZRDRftkVpQpl4oQuovpXmDLx+GVUO59UR4rHRDZh9c4i1L19hqanxFc98MFdd2
bkKpt9B0NY6bHUM1A+l4+F4SzYjGQh0aJfcNYQ4Rj4wCTdc+wu9zH41lacJPyYtl
N/IeZDOgzHF4s7YIa3H1RwqZA+zTeXGoicgOU/ev8/VLnKSenD0zPvXYwvf2AMLO
lnQwRdSV3vgJtW3gkGXHn9nvREE8ZtjGAeqUw9nqgbAnCvO7hQcfnPIfyAPqxUBd
m4KWmMU+7z8Ur+SWPOHDK+7ztc3SD6HowSK5sCD9Bi0Ok78FIHjhiPzIt2K2sJDL
7bycXHAm0Ekgu8odndwRwpOha9z5qt48tTPsZenZHQsu9pK9OCQ3SyQZDYL3eRHx
ha7ypctb2TuS+rHf3ZjZUAV/yaaKIYCIO9FX5q9eoHJIU5EbfRpF0DqVCU6RRvAa
XWwfUICDiYJorhGGppCXT/chzhVjzJOUlG1c2sxoA7Evx9EIg68rkNIWR/FkeHet
eewffQD4V24g6Wfz0djgDmJ7AHwFU/p6zSJLEi1EQuGX0JeC6csbpWCWIXjhJUTt
rTAD6nNziAHurcLS2Zc7yPI8TntpF8vg63iigib9tUI69pc5qdqfrRDCYLpM1DFy
kSQPxcN1YW3GXcLcu3aMAYEpWwW7S1DsgLkYtq7hjCiD07LuGzX3uR7SqEj8TgIY
N8qdqcAJuzvbX+pYbRrfJq7X6y6IYIJz86RB5UStrIo3/mRRCKJho58fm1MWp09k
VLQ71H/KFX0KUHNrvku3FL7jIvfGW8/7cjEniKzad/uGaDb0d8iXxUphxTiCVJ2x
paZ/qIVy0spiN7NbgoRLw0IiZTzdpqyJW1QOMjKThG9R+CPN58UW3DLF6VwiuDz6
PyrE3D188pzdv0HdMu+D2r/qHm45U/wxfbauduRmBovK+m+GuqwWaPN4UHVPL+MN
togbOHvlJBzG0PyAKKOB+qT1l4i7XNYTaatEYxeBU4GGnRJ/kk0Bk4On1bhc4IUo
5oOdx44VdItSZRUwu/brc+rExHdhTR+NQYVziDurWbbnzWGAQL7s1jK6JXJnsFgh
VclgpRnIdUGnCH6IRaenZ1UkDBqEydMomNaJlbdLUrhbf5xwg3uYq/blIuEaknow
17vm6UEEdEoRLblzHSbyCaKnt3qsXYOFfVvT7s2iiE+qgf3ZQHzU3Tn9a/1d9IPD
vZSbsZEUMf3V13Fyz06M1kqg4Rpo3KTK1KDoowLgUw+EnhM6kRZpJCSETKcbGCOL
5XXBxb3oI1HgYuhrak6Qwd4lSV5XSKZ3qjXr6V4+9HijBYVNhhKlNvdWjQG+x849
2bgufEWzrehAUCYzElhvXu9TvYmqWzCPOwAslntpXVfH+t2sbs+VFqYu6Kne9HGd
xl0KuqCvjxxX+8DTDM6X6P3NkmSWivEwRSTTa1gZwLzBHIyRmgQtuJKGg9gMY84C
cLyp1VWEy3m7ypv46ZogOwJbfp1ImFXjuuWby+SbhClmGVzFiQrh8d3GPGgkgS03
wOto9LFLFCaD3m2nkoefZGbNxVlMc9Rl4rfIdbDTpssYiaMUvrnVqDC7pNYMAAxi
XafVSxb1IsGMdv25tGmvK05cBn/jHVaseVuBH/2OPTdjTkGGJlTaZLDvm0UZMFB2
qAVPsh/RJ1ztuhS5Hqb/5zq5zIRS6I4KoYUtIw2mVzl3+o+Jpg+D8u7CHi06Sqvt
axK+KMx94pwZ1k3vGmwz5h/sCrAVvLxi/eGb5uBvp8LkbxkmRfy+6PDZ97mjCSFR
PbxyICCtWQ6cgwTZcyLZU3YKGAWFnNodxoLNCke5hIIhHFe25kh9dz6JUDyVGw4k
m7jhTLKYPm2Cb0oOLUeVpvvp6sPKaMsdzU6Xqxsk0FgulKv8TizKeZ5PWm7H88Wy
YUSz2lwQs6LkvDss8oBogdQ+ftdpSrg3p1vUXvSdqp7BRu8DgbtsDqaOGrWHZ8Aw
3pzn8p4MIFpykKlM/lGksI5m9ugYg/y8cKv7rLbxVp3YzwTIAGEk/4Ypa/ZFcPJM
KoSOyBD8AbCKHO6hKd4YOtOyPVaod33U7I/YZWAhQqG9jOmbXWYd7d7maW6hkVHJ
keam1JTNfwsWUyJA+Zhoe51x/IEG2Rm/W/Wjmp6PKCe+h3satFSvGkhOCJMobek0
xeZ6alO74efkNWhAd5asmwuRlaA682XgH0LHk7dsJnYmQyzuFhSvyY/T5/C+PQl2
BuJBGaybxqIAaIZAlakHYvHSIEmsFYb4+Dz60UcbePQrgu+iNxumgU4oPfVedcu1
CGnl4LndlbQBSOyfOF0EDItP8TiYC7zWRMijKgALpJ0XvCBod3TJo04PdAF4iXMb
VJxoS9eQVLmdfNiQgEm7x/I5cCiqVO2noC+VOeS6Ja2IMIXmFQgcZdr4dbtXqVim
IQWkr1PJ+0KMX7uTApuSKAQUkHPV/TSDuPHFsOFwn9v4wIQB7N3pjNBQ7iB6lxld
RfgDG5e3SznUANGGIpvZ5W1fF3vgEZWx1FTm4IwQ9X4WfZGUxvFqjYBhKfR/ykpg
ya2dw4861YXy80IdmzV5JE5Wqipc6VEVMYtwuRiKCPsdhpGfP571AC427xWSpccH
6GJ768puUNxnCXDT6ZNIK45oppXM0FFzaKHV7gy7TriUGkQ+VmJN883XrHbPLCxQ
HU+BgIDqbPEyVW4L9c1kszRlEkIdtJxcfq3qIDD4Q5zlfUpBjdat6e5mGK2y1Iaq
RsttzUjl3d1cKk/b5YGLe8Fbs4NKbAARLnRA8DyHRNgM8yYiTzq3jy0bUWoIaLJs
CkpGsP+fqmU/t9MpmI2qpXSSYX2OyXpSy8Xlm0b/5gjoz/VIc6V010gbaA5P0gXM
fRQO7X1EuqHgXWFT6bvvaFb3mi0D6q1JIXbJuyOquSa8PiXsW3mdiD3wqXkcs6vN
3K7kw1VN3RA8rAmU4VAbYEqv68GALzLJPYGAjqcFiS2N7NUYpUIdT7faSIbCLNky
rq0bSUhh38FgLHTpCYL8gBsu0e2NQLC3TNSTsCSQEd9ufVrALmtovvBXU4oG0AkZ
zUhX6WQX7wUfUd1/JcqDpcnTEoudHXtGuzL/6XN3Vb0Np0ZE9dTVoo4VPuNgHYEv
i7T9jvn/bqYkG7/rvXGupNbN7xOf8CNUNG2TcuTvFD5YLnc8eCK9NqDQ9q70BjhI
iafqP0YE394oA5Toy32h/w==
`protect END_PROTECTED
