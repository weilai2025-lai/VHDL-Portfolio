`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGa+xVP2PfKI+cqlsUXm7/UMC3U20me+bupcwXiUuPmFTBp4zy5rlG3eCrfKyl3Q
wu/+7QRvSlmxM3uLjnjWqixO59qr0MdO55v9bT8ZNvO6FSeJPIPFjg98RXQW09XP
Icz/xQGx3qBIo/UnUm0FELz28jy/+wWHVY6Hp5Y4PpjAnmHaDNLO4FM2HGy/6j+T
TtmxixMzHvbUWgZ6REAJnaRB4ov5C4qix85PgWqRvXtgtyQOlKSWrBX2WvhxZDKy
THyaahe9UmQIgq/aVSCmfZt4HDW58uui+1Mtpg/HXD8B2rEUFj2NhjWWgj4aRNXJ
sX9S8qzSM/oS89I8PXZAiK2IhaYzjFMuPeG3sRkmKgi8HT82bIA5lTElYC+XYEMM
5juzQDLoymA2/rC+7qneBXejIK6heeK1rKkGT2VhqbPhYyOFaxxEIXZL4nF6TR0J
C4MtK3j7npDW67QE1ErzQqhJjTGnTkr2bahpDpMvVQSvTKQ7HPvgS69YXY/Lvpxs
vYRPYzDlbjimtCWUAUMZMDSeszI+uVybT8L8jDCxXHaeYJdwJzZdMW0qFosbhBYf
1gCurQ+GlY3pzZ1Fz3Ugoszcpi0m+XYD6xFfEebnO4FNP9PV7ZY8SgU9aTdZD2Oz
oeVaksY98Iawkb04FVaznRnENqVxRZBaCaIO/drXTh/gw+kxPzf4lg/jyGgkKVLF
NoLYa6zJ/2Efdmq0ipPwBRWZuCIl13Q9InNvH/ill6MEzw3hUz4QIJ/dhp+R9r+k
vsJiw4Esn/plffHZTt72jucBr0q76EbjaNUsKuMn+bf31AWk6uWRvsJ/Dloghu2Q
SXH1VRZ7MPNUf26ftYKzHM053QrSC0z3xK0UxSdIeK2a5mGR083JlAm8mIx6fFI0
pHPhXAOQ9nIIgaAkZn45VHTXjMWzHk0yB8hE/H+8oHieatwYfrHgnj5YCbiEqIk6
g/Ir5oHDuoAOpWVybkxLG8tYGgmX92AK+BRCZ04lELz5FPMlvNvK8uVYRX5z6MEO
rLxQpN0fZbLYlsxbE+SdoIi8g9UAUL9r8oPmtE4IoIFxvWgcqnljCRutKu468KVn
eK764zAOyF1eJtAFcCEkacr0iLccXBDTi4Qo4MV0cQh9Pam/SpoXt9YTcZW+l7f0
iYsoAAn/5dfKgSSZ6mvt5LaQmJYI4gHZJL0Wzh3jtczfTopt8vVi98ULFLDOnYAF
Qi9BCARg2QAXvPsZsXBhhPTB/lOyIJbcUEVMi1NbhUAbfIIlF4ySiCQaBptiCVAW
VjWkPnDwmei74tghym2L5VGVcNUgxT1hMPel9/3lUThUUVV4U1eXaJW7f/t3HG3h
yVg9JVrwlhdWI9jmeHZh/LHhZcSSpK/YZMgLVPITKXz8JbX1cFcCeRQf7z73o6/J
jo6jgAocWvg537vASwUtG3ONtpL2iHmS39rK2tGlUUGB3oYgDaFOwY28tC5qGTDb
zL8hZjO1lPgKuD7n9x79VNZe2w4k9AIUndV5T9cHtTXbAVCsKtkeekX2toAUe8FH
GR9Un+sW+eqXpx7z48CrrvzOBWgCqg1QLY2mvuDCMxt1hOVWzKccJOZwxU29JfkE
rrWMMscMM4GrXm/aJP+GzaxvnuqFKwNU9PCQZ+/YXQeqWYJfzE0sFonvqessaisM
S2WK7nYHM8qVxG3ABT+MWAp4DGYnYusMe4Juv+qLW3oxqVqoA6Deh/e7rmFHvVb+
J9+RSECLqsVHFWCKQQF9M162JuRPKA79aCy0a6uIqu+SQs3pQ4Op9VYtYml41dPV
GzWKByaIeGWuHu1p5YMzu007mKXsvXpcBm9phYFUoaQhJnmQZrqu6eF0MNeGC1YZ
GfRaKzfxi0Y0FvadKJTOgY0xB+6tQCQ2f9i0CyaivtOvq/kEsufC3NvRJTTpq9f1
pxyNtfUy83B7jl+frGUXRkNEMoUyEukES9wzUFqhTyFb00xkwVBc0ZUp0fInEtCY
QM6jeEyM3V9SWO7bNG6ETbDn6v3jGXvHeR2kNvtIS/J4QOtNomVwV9KyTr3Y0s6A
mheRaNDovekneJTBtyr7JJN8pWL5KLAQdqH8g5aC6uzsHmkQzOW20S8kncVxY7G1
ZcCPTEA9nNZ7LGS9nqMkm+XBsrjMNqJjW3zxCo9VWcN+zXLo5kJ2ak8I2abbkH1H
Nf8uXv97uyIhsKCQV7ORQ8JkhbYUn291QEfXpww+3gqskg/nJXOgwY+PXG3Mslwj
nL5wvKa2/pY/nXWLCajgThoCW1BEjc+LjNTqVQCFx6iobP5XVLad6Q+NPUfpCOh3
pGfvxtXhBXJDr6vgjHh62FH+Nh8E8t7TowX4rOQrChGgy3hRvQsSAvHEbyuPAVPp
3hijxZLxB6FEasV9kCs3f9MCMlPw6qduaHMZQHiJc/AFmBRoCFqL4y2JatKCQrFr
4kNeI0iIY59cNKQgLymQv/fIwEKFmbymlw/KY0cQBE/71JNDC0Zo8klL68iHXyga
lCuOKNx1oWh9WWCE4HGrG5lDmQGNrXArZpw8h7q9SupGPr4/Dw4bWAc6Nc3uu3Cs
YOEwgqVl7KvO6HKGRGz6kZFnEJ70XSLa/27rJzhi3sf4O+sd+hQGTct9GeMsSBcD
Qr77rXXJ33yOn+n5T7Ch3NUY9y6rS2J1FgoWPPKCKgeXax7KYA9OVqJC0HTbPjPd
v9aHx6FKESfDaPT/injLGLKjo2oFy2jn3uy/avlpig5I0RqQ5FyaHhvvuJdwoHQi
iN4FqWR/7cvFkgUKZolcRid5zphElef19wUSpOj5W6RYKA3qngfjo23Zk3aj3CwC
Be5ZkANl1PZMCEEcOtwa8VT6Ht+hTVUTTTHkKo+CmgnIJ5QHygaGDWJkCtxZ9Bjr
Jvh2xSBwD1jk7bD9ERLIPNpJyd9hQTtxzNdOp6PjkyNjUWgov6ZUHW1hgVEBTzg3
rQe57ubbfcu25AtAEGYjJox6a3dkPD7zXGcoDjeOQfKJh3Pftg/4w11n4q75fjgj
2VDzQVwvmezd9IB73uul86EuyET3dsmMH4NHWoNpj4njLTSITfaMTFSXDeWfZX/F
UeXMfSWCDHv1lAdJxLe30lqg5xDRhqyzKaBXkIsofQgL3BhdxrdpsKAvC46gt7Jo
M3rN3xd2mNbNHq271jG/9a2LXQM0mwmc3umA7ReHbGJLTh1yhL0RzB8F+nm+t7UK
Wgil1Pjhw0xqrDgH8YdsDBhg4uxGR6VzUlJunVV507wqV92oKR+SCEjUXvB9L5zM
TudB5l/RuAu5hXbrW8XrExAhXiVYF0kowBCRHUtEJlHn55OYnauMUPaIxgnqKPoI
bk6oewN8/XktMArhgBNpqQ8PutwK1x0hTKRbi6vsk/t1v2BQn2SnRartGQuFISit
uiNqPaUjD6SE44FTFWOwbxiHZFyNbFfVBdmXpQpE6YyTkbuIo+qRJUYBx71Oc69s
NoxDTH68d7wNoYno6nYKarAn6zMP/7xQuMnYDJpyniyvjLUkgO1ICXEb/EMcgr44
kymMWPiNCu9b3KJFbJ93w5IuZA/AE+7s18yfGB8rIT8vZb3WcNZK0IF9pvkDPWXf
n8mG4V8XjYds4Ns1FT56HWmvnKR0oET71uTJJcU8oc2TufXqu2XFIQeiKsP+Trlu
3kYIPPQkxXh5dQs/NtQGPnhwRBOy5MANhZmcrQJFSnmyItQp+hNVfaZVJj3DOmf4
fF4xKS8C7Qs0GaVZDiXu3wuQp5lT67PlQpLyx41wUBGD+OFD7fnq4GjNjPW0UouI
F4G2Waymj9L9cooQnxKbuTTjdBvtPs6IGe1zrNuIEVx5O+wjEk1FKmjA4C/Lz8z4
WeMw5KYVglf7N346TTevLBLSNqLmFo3gWQIkiHFwFORskXCQOGO4DkOR6dADOKja
ug6UrWohgXmIBe4vbdgluYgcm0DZjCUlDBMibHm30l1J+bTbsCmV/eeA4chrkLSs
Pk5ckSIHBXjapeLxyGNxkJScNkgmvPwNUSGrjLkBY1uxfJPHVnSH6kk/xtZMtTcS
KZ5d40f6B9wMQWwugFGhFFO+7pt1bwJsg7ugRguQ7MGf2US/DzbQWeb09vXpcwXI
QU9h/Ld/uZJCy4CUGJpcwBuUYJM/Yic7aZ1z9JB7IQN/3ivQb3M9Ghn51yPiZN3h
FgSBZeIj6KAIbqbESf+nU6pqmHivYUyAuSkMiqsAI4h0Wa/Wxj8Tm4uQCYzsKFJr
9cW4nN7v2gGlLqyGtD+0tmriY7qFcCxzeuXVzmRdvMm9/zYAuelOOUXPDwIsiGkl
BQeRlY599gGs9VRCliH/UFhfnW2QU7U5bBCBKBd9TnDaYLkAJAid/49dMTU7QkmV
V3MAaBXVpEK9OGwvzaTLEpg+9+pMqL1k2pT/7iOgw9X1Vbov8y38FKFvhqEEJiUh
zMrBVzVLOLnU4P0AI2CyEUCUAxvKkkelZq8By9vFwuBiNLmVlub0Y7GQUAEYkXq3
8F7WKHsAFKSYvkLBVbYSgBQBIyJprf63Yla+kmTkUrMbhbgdLhGKZBS611P1Q4cb
JQIdjpqryy0KKOIiqY7ajhIDh6ulCEgy+lyEwAUhh1oFCPjAM8A/ZFwyz1Pp2fMh
uxw9eiv+d5uCDT+shjeI11Hh2hAS8tiq8p4ybhg9sGNSdxapXuTrS3ekEOpSA2m/
GB+nYNvoxA8fT2w7mcUJrW93GQ/mni93eAqOHXePeyQzsA3hOU5WOcAFRcSFwGCc
LAGSViFAdw0T9wpKmC2G5yZ8/+OzgLWUTUq18aKkPJ+N5HAvQ32GoJhahTLCgjSZ
sQTG8FtM0c75zsGrEMX15LcbfPQBORnfGMH/a47spsOw/xD3hQC4cbuE248I5LHo
DYRQb5LfCDShAc9cGnLrQFKtalbSYyQPvN3uowfAcD4i0wMRnH096l3RvrjbtiKX
xOfSRxE3teMhL/s4iLibrV82vR1tJER1ROqHTe5su4Fo1YNc3SgK78tQD0w/kbBu
CebLjB77v3oIV0FJ1FVpsL1+Ht8J9wpMeo3UKDXZf4y/XLjxwbYHZAtMSVY4YucE
PiIRfP/RZQ+qWwJxerhCjtWWhZOR8H5wpK+XjuuFu+0njUrW/bSUZ4EpbsojuIfk
/BOkWxpEr0CSeREo6ffUI6GvIqpbUsjfE30dEAl7mKZWj1CA29Ix1eGpKZ0HMP7e
7gOWJ6LaHdP8aMACzpV2E+t6AWh5zOGlkWLpe0gBgXbYYoIoUweA5sycRNEo/PK3
mSjB9Vj9mBFSDfWfB4O+nahX9wR2RDIEwySzUF0YhvMhyq+iSDiSMk/MeoXtGeu9
ljh2HsXu+skDT2mwP1nN13BV96WOgT56Zl8HQNmyR2BzcanBL7cG5pfdseY+4TH1
8sDmQWtzMf6vLIW3UMex7Vwh5gSubFJnGjrCdn8ioYgvZZkMJlkgO8InPvWxATkN
joq6AwjYCyscyhjbid+m0K3acgoFACJcaCZK3wjzhmnt4gfLDx9/V6lvGHKOtj/Q
VKFEJOU3M0kssWu/H10wp3f142MoXLCuCnZK1jgpE7/vLuOP9w4G6h6G4QjRTQaE
7t23cKUm6vw4Twt+6Z9tYLi+1TpHERzD3Pf0avJK2bVo7Zc03Rs6VuIn6pFjZDHm
JsuvyNdQ6wPtoO4pV/faz/NpyvAWQ+NxTFVeHxJTeIPxkA57COrpYGmqHe0d0W8C
pCVw5x1LKl9QRkvsAoieLWYA4WJ36WG1MbhhEpSQeHYfRBSzqVXwYnUReNuGzbQ4
fpHwD5Wr88Pr8khx4IuF4CPy1/CQbg6yrdgBc/ECBCbjLj6R7R/D2DthiJXKPBhd
QW3HTp0lQYeC+PrKcwe28DT8J4szLfrc4Yae+aMeDYwzGZbquKlFDkep6RTw0RZI
YZmCCfUrKchkn3a4aITB2TunGbdg9Tq8QTQ/CQONcQpHFUbqz2sLCl0TbI5fUtV3
lmMr+Tpo0HR9IVTKiiKoej4eYCHzJLNM2KSt6oUrrZ9fyObbofc3CKRA+J/C2flm
18ryUVzNUrISsI/HymtqdzSlhXBKPAQrU3dEePq4QYfS2HepNtOP9AhssqRZ8C0O
n5xVYjgD93PhW15neZ1djnA3RMvDy0hFUw0OZnjjFUWg1EcFHjkCmPBP6hWtOz1C
nzlHaI+rN2ZMzZAa4E2N4xVNJK6+wLwOdmnZP1WfaSAE+OqobgoBg1uZr+uZlWiX
hrmytz7CKZW22bCaGvaZpvCkqxmCnW6u63B9boRqZyOuBA6pSIkduaKL37JeyH3k
H5fGq1v4ddkp26qKoq9yFTZOXlQlDclNcDU3JmJox94cI9C6iwKapqOKoF2DQ7h8
3ER/Q9pZnOh7lP58Jg85dDycYm40G//RHXn48m3U8wMyiAV8x7uYK9pQUG+ylvY3
Xs/bZZHhlURi/YEpDTWOT4KHyrsPiYf3sZjxPm8gLM+4S+6xXxTGCUOETCDoQjop
Ihl1bA9yKOZ9EATajM+6qEsXVxeEz3ZXF3UVlOSLKSymXPUjvvFRU7BfCGxJNv41
3c66Sc/BxlYo1NnNrcEQPd/irBMS2Nb+6Bj88wtPq+1UFiBt3JE6/SeLLQ+ynsxc
ZWun/cbnurk6erunHsdvoLDbcDBsOmU8Sk+4BudwDc3BlQXPKvzPWXYZF7wdZqGY
d4CwAD0reQ+0nCbMhXY67bmZU7Mhga8zQg15Gh/HSY5fIh9t8DWagz5WvMnU+TSQ
T+H0b0+kPNZF6J/1Q2LEsxIt6Qu5ufhw3XiXhgr+VIGLRRPiiDRQyCsISfP6CFzJ
btUc30XvjcT6fvETz9kIhsESfdXHqw9HIWttrjTzGBN/MqNfIfQsetHOONiz9rDU
J+tbctZQVkIO19oYKSL9iVbJ/4CthK95LhwOpk1NfNGDDqyPo9s6lxf5gKc2G5Xl
8pPZ+C7r6f0WbcM94z/SQ5mlsOxjNmE06MeZh6YaawrNm7kmUmvmVhk+mev0jFK4
nbyrRlo4br9WqgtK8ozVfy4ZrM0D7Tgfjh7YdymAgNncQcYe8J4lmvB1OollvNRH
jf9GPiGJlPvRuhByO+3QdZumnqM+scOx5iCx4WRm95OTxs9yWEMp4z0fIVaui0Y0
/ucU+ljbOlmUHzngZko677kZfC3hFNdeM8JGosOPAlbFY2Jw9KCHIKPwcc3SvMt4
kiHO2ccpXROLnpXa+FinokguDRVTISAHvBgd1vN05bwig1qduTMDfoXMBqrP9i25
xAyTP7l/NFIw81Dbf9YKOf0eUGsxUsQZ9ba28KENldfCXa7F9Ip3/U5tHLOeRHfa
VUTAqkmAlmvY/AWbzvUyfqnXAW3Tv2XJRDKCcfpcqHb/j1IIpzg+jWPCizzR6PPO
cLBt94DBzlXA41nT0ZZ3QP7jljsY1v5CriYv8dOySK+nMAzTKhFpRk1s4Jo4OCvV
lppLSdXSN6ci+9p5lhRCxWqx2CxRDBx4TEYUzR5eLKnKhcX1O6oE0hqKs6gv2hCa
zKja+cfJTgZEJTC8vp+WkW6gsNYw6G0sp6N9cf1CMZNGfLZrhxAg0ephJP4dTR6i
7eqi71++f4vsSmJ5Dp8rLAzmrvE+S5khkvAba4M5SiSP7dhD03XegzUq7WztWzV4
yMI1tGo0KrIKm/tsbDh1h4g4xmy9bil1HlQP56u4fhcdwzc7dL0F2gEihFOeaclQ
gmpQaefQotxmUsb3gPz+f95KGJCdxFr45fMFCCONCMkG4ks/650g5WEuS+jrtVWR
xJv1v1+LYjSe68H9oJihfiPD2fbVCWX8SiXDdQxkRtqQwsnt2YGdF8fzNEBwy61/
uzMDanltlU2DbgNlTooaREgClQhm1bj0RKD7I0wjzH4l4ZA5VsLFlh1Sip5LMCj3
fI4Y4jP95gQByo1RZ7TBk/AxACYzNPB3h84X1kR/+rXw4HzkU2V2Kl+m6y3Kz127
itGJfCjB5uVv8jSzb3GIKpwJcf1rEEDE6p6BWqzQUTG+E7T4SVMv6Hp1AiJlPEuN
UtTJCBY2EC/9pXAemrAThvByopXuicitS98+jnsxmbadHyUr8q1THHVsHRZJlfq5
65o2EPPIZs44skxK5u7fbex9RKfbENUzAnqL9UMFUrBDgQdoh8or64zpOjPsjH/r
DVTmqpG4fRXGqFjzfLTj9RVnMbJVU92Xp/16uawWvfZBqhRqCDrjaXOLxYBzyP0o
r9Dr2mDNxd4DPFTM4MHyYjV1qWevzEZCOAnYOGyct331oIHohv2FsIsNsXCeADHb
5ZeAb2TSuSMScFdaV/dTRbquymhiAz1GI60JQYy/TkeNTLxj2y3at3P0WnxKZR9x
7VKndeNJb0RthpciF0akaeAdzJPd4TVn6VEtTZA5LXb6JdZ6iVGLvbZ/UvFcw9Gh
Sof+1W4b94XwzPUD+7/Ju140+G+PUxnWJVclI03M0jJhqjEdeS4eRYeveC/ISqke
ASar0vrCunjMbkceJ7nhiPAX8pHl9QlILdNnd0vxh2+O6Bgr/iJzBam0vV6xUC+X
HeprmkdUmXz1WuZCIkccDWFDFJwj0eF/ueuvBzkwa02GDIVEH7mVc/yaRIGqCFBD
v828rED4mQHShkivL6f4sDiGexCEb6SigxkV3gtOa5qemHy2rNl4xsnAXfn6J2lP
PO3476QhOI/AmZdPzI5GpMWv+OSCxCPJqn+7Dw0QaD5zqM5y6tl99rpEJVc7+Ffx
uSA6XBpr3dQtpKBfyTakKjyw08/2olx4tgIXbKGP/xduOpkwr/OwCJrHXRRTBymb
tco15bA8nd9Enm5YRR47OgkxrV3UpJJlHDf2GwKMAYXVrYci6FgP7Z6tajREUIFw
vOnTnYw7LuOxAatkCHpPAGR8/B3PDz3vy1G4eILb3Du4Y29+BK3qswBuSknp1xc8
P6b/S61SMtqoz7rahQkYLL098X5k3QGEmITtAukGYUN9YJ6guphCtA3YlJc9DeEV
fFoVTYfOwdLvZI6ajCqQEWO51Tz0BQaCvruWzY4cziF9ABU2G/654by3zcn+aq5S
Zq8/HV+hkK/fhqUVNmaaqJXo35qXpRN1mAVXx6YHkxgNlxNwuRdZtxbYWqfwfX+S
be4ibLmqP2NGwWQVMPXosR3mC2XF29oiCWa5N2XwtTdTOVph+66SuMxHHSMCoQtX
4v6gC9/2tPYan82/2Lfep/Ya2vqaITAOxnaAJEuQwPJtHfp+Sjr1vYz1fRsHBkfE
EOV66pnHWlVMcwjxhkYIqajQe1oWSNuK0nqvPfZrpPDJVFHk275SDpK5ZeZoRViX
5ZG1LFnBgnfvl89VRABOxjOxYQll6unKdfSEfP1iT+p4sumZiBkL8WkGg1pbCVwq
srLvowFwMe01RelFNk9t1+4pi3vzX0yNdqge+JIEqf52IVpIYnL1LC29n1/JVZqc
OC90IGeDSYvvg8MUlRM/GgsGk5rFvc4ZtmKxv1bNkvZeL/9zksn4xtrGPacgdFgq
iMX/FG34FwqSpO/+vZlh5y74h3C3kgA5f7poh16Xt0fcmfFojwxT9B87jiKfhdse
3gG2g7s4qCC8LkLNvTWGY5iNETDVAE7YMaw2iv5rNyzUJeb6M2BHo+3auC6x4+dE
o0OmRV0OQ5sRQ/ldBks2cRg0QxeZeL2QOQUst1OtHCZAf8HEFb9+wqfo0Z6Qq2Xs
ER7LkrqAnIzBL05V86wLlZdkTRqMxofnJ9DusMdsDoPMeQGDUfdJQy1x+NFZzMyl
vS+vy02ZUbfBBJW9pOEtubmYqoOJ1xMmbY6i79FR82lCIfd9yy4Qw9AXSUCazVI8
HzVhP+w+EDPY6UdzTvwhv6uBAQGaAtUqopqpdRTurM/BS1D/WHVM8aVIxZoMTo21
wgorUW13Oq0kv9gPokr2EsGg9DhQUAexNVI48W5LB+OGn1aIBvbTkHaYtp5cSBBE
u16Ynx6Li/DVWzThdhNwLcE9OI8NGYiYQY76AxxDpv8YQTA832vdeP5adoXLfM7V
4ebPKH5IUBAAE4kF7w6Z9ijxf+5CmJbojpdnQG5SYli8q+1VO/8IyMMWY4jcjy3R
eSKvlCpFifC5MXOr3THUvcwekL7/0nLULv+k2saGWFaPYf2O2jFydDOeb3qvIgXs
bD4i6J2H8E/QTHQwfiI+il2tEiOfH6bIalEFBqn/pswJR25f6AMTykQyk6H0r/s5
jWSDQhcoHG1QIpOoAukRKPNjFNo7KUknmXPGayKAlYW1RQUkPhfmi12qoU47QtFX
Wz2aki05VcZwb+Txsl1LehnH1WO1Wji32XTsH4yjU9hcX/TXCwV/ocP17x914JBc
0w63lDhuAr8x5uJmqpocXpszjZQ5EV58rXBRiOEVH23rSgq+prKI/8wKG9iFJ5Eq
Ccp8/oTTCORjdoRCJhxmx8oOE7pLEeAW812js/7U2WS0+ynElmQrQujcRh26Mdb6
waKyVYdwsf53+SFQ/m7FPGA02Kgznf2DgkDNbXi16xvFwwlrrCMV3v4SBVW6i5Hg
M6ZAz+yyE0FkBU/p4wriCcl3BODZjjleMR1Hi9JkIH7LRtczbrKr93yT15aHNZdz
CnZEZt5AtzL3dof6Z8S8cSkoDna5hkBwoyt7rFqK6Jqfj5f2Y9PjweNUyA0exR15
FRvyYGX/NvtbyyPHX0AJlqnLZi/1+R008e/v9E5b0FfJyiB2AmBFVPWf9FXxcN5H
Y+RTGd1/UjsmS2ZT7/30pQ==
`protect END_PROTECTED
