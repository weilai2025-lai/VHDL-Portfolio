`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SY2pUcUSoZcAQMrhHR8/2DkywN+N+oEUqp+9HdxHsDqWruX8a+dGqBGvsizIA098
uZGQjFbXCiYIL2acVQ9c5e6m0XehJ5ZtinCwe7ErwINwJFBClAVOhlS/tvspwDVX
HoQZxy0p0YMas9ib5aH4CkgvlpgH8QVKGpBK5ErlVP2UFSTEW2Dl8LFAeUqyBPQ0
UHAcwfcxyOKusvBPZYtNF8vcCUqzEE+kDZJJUOZD6sySeuDpOEfm8tHBrNw4BXmF
cgwURMhv1esHRAFNJ77EyCuh6veNlM9gzfAqkBN5t1/YbWMhI50RmltaY1TLDlL7
7X/7v+pQ55Ik7naSHE1l9TaBaMepROs5WfpR4JFK+DSa3uEsxdh0a06LSGc5SVF0
y58D8aTw0muwG+usgHuQbqF5LhWhJIEQEs0yS/sVr+zY0FBHL3q/f9pfNbq/Lo7M
Ur3tACyRjb+czD1AIDIDd4L85P/kh0W9tNEDxr2r+oRqw2aMIzS5k4mKxF8XCe7N
wGnORalBTXP68zxBCyFSnBfhgIoxK8ShJUAWzmbZzex6KelI9cJeRhnu55+PNjQY
`protect END_PROTECTED
