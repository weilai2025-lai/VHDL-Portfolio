`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9qsqgoCg/I1cf7Ww+D2G3R2/+xmz1lXVBrMI0/h2wVp58emlB+yQNmIGLsrBAXu
Ngj+oVdZHfJBZ0xve0XRXBi1s0j/iuiXZYrNaEScBOYxmDFyJ2Zc7AqL/J69fZe2
nUSMah66uo2UrSDa4ty0s3mcPbOXv4zzVRtt30KgCUbYYwNfSWHMBHsx9d0EnaUA
PDZvEiu5jG63r9LgyE4pDbN/4dcFAQM+8OQ3JYamkIOyygLgBZLVLU+phndI0LPd
eihCqLU2bzYLRBLcHIvuLFNnTg8+FDWve28LUEp3/7VnkxSAYzUo0jlM08FqVz/O
4RtvKu1rYBU0wmbLPlqJVdMfPSByb+y9l4dpCZr7tci/SDbaFoHVXfRNYnLlZHOC
wAEwczdWA3FkgNjTYbaSvXOS+CgCMEcxTbODJckJ27gWZEyP6wQshPQJqv565FPS
1nGUiVlqBK5tRVGRIsdX0ztIHqBpcilAQJYFR9cHlBkcBAEd73HU+pXhjlwmmaq8
a2tw2qJEkJqJ/D0/VvP7ZoJW3hWmASZxq1xJ8Im2nS6nbDj2mIYsyMxbn4luD9Cy
Fqv30Oca3dt0pEhejLoqqWa2wut+bHveZeGSPWN7h8kHcO64u6QAXJzc04EWF6p3
XK8b5uSQpIrv38zLJmJVMv2ojvWgXWhp2FzYunb46H5DltXJzEIUY7OMztiaH7q1
mfphz+nyff8Oh3tCIEEf8stTX8TCZ24JleuONYkuewraHZzN2Ck5HQXSGSc8/CCk
I8efwuhMzzhQZ7ZSkh9rG0beXpqMAzcraqBRSaOeqvx2F/AuetrlQ4vgdNlnNprR
dD22lFCHCMVOXtKefirE4RqFm4TCKq8IA5WDzTnBVtgkBHpLFkdhyIR4iH3e6SE+
p/OuitWLlvBH0KHQLpvjddMX+T2y6hCjbuJMc+3Q7V+MI8+i3eJIK9JiWhLVfFYW
qSBZBYx7fnc65odmLFg3MEqwQMDApsqNB0QxeoX0QQcI93bJNi4XfplAk9PmKs0q
bb+7dmg4+Qi8TSiC4iK1IeGFEbp1CnjE9Ofxb0xnaxvoicdaM+3hVmaUNBEZ3+DS
a+P8Oi/+zWukkA24k6LJm/zIcCP6mj2RBQR7tgq21y8gDqKc+g8As8QXcSGemtd1
Jb/M15uu0W0cmhlzAQq1euIvf7y+6Fd5y97Tf7UYkKd8A7FehcVHoyiyt82A9ftN
VO0npKR56yShbLemxpHSah521JYUH/dBpT1z8NdW8KwjMx3BlIZrXuyzrZLWKlC6
goMBqXaAhLsAj1ljWsXPqBF9W5S3iE10zIqtZAq41/b8Fy6FfPlB1qVZ+KPOYwQm
Za+38NGx8o50zVRoXeadCxG269AoAula087RJciFYQfINTDxfjLy5EW84QtJncnN
T6Pc1pdGE3iylZcxLXC32W/9SWK2s1/OPt78CjDWcLrNGMghNgWGVYVDf3hjiJ3Y
`protect END_PROTECTED
