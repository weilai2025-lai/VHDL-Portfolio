`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNgKXhqUi/H4HJyeH9SLdAXgNfXmRMUkY2Y7b+VZ0WNt3aRpPib02CjF3APscTlB
YDCn2UUazbpdXRhZnq0H/qf0WTgkQsIhET395XlAhDN+41gqgtc1B1yJfLyTo+J3
VPPh5Se03xyKlDXL1zgJMhTkYRifqBIBGB3EhIA9meN/khl+s1FkV4BcBETe8RNm
rBl+LULUICSLLakl1+IZf19WvkaLYRaIweIWNmx2OutzoLNpzJA/L7OGgQT9N6TX
R4BUNuhaTM86nFlyyxQovxmK+wogePCVjxeTJ909IqzxFLDdbxzZZNUctP2buyZ7
Kbysunx7w8QOM8416bD8lzY4qL/hSSz4DVNX4GluLw/BTiR6SlZxdUGiatvReeQ0
PXZVqdCqOQNM7TNaTIgOK2Zkman4UuM5mfQZc2BO/x8OU2oQx/r9kenG6hLSUYOV
MieX+Tg3Bp5KvWeXFR9VTYfCB3DAQp6RKwh4J3lspD+8h/VC64a3xBl42+BX+a80
sr7lulQFw/Dzvk39d/Eqxok/nWY/Y49XMv0GTYWKUqHT/WLpbYeYfyn0fl8R8KwT
0PUdtV5lL2Ppb5U4/oiDuy/l/5gG5neXKTbI3m9y7vPl+F6mk937evqRQAiWfGSP
4uR/GRpcRFzjiatalmEqakWkHNVi6vaB/4IMvi44/blYp3NZQJaZ/Z4AqzlD69dX
q8wOVZ03V03ifo/zXvy5c9JZFtiLZnTz7MaK3xJfNtp7M3rQw7jyjqSpPbx3P/yY
ExxtzPvrlbTQonk4MFis8ORUwCG/Q15krReLLSxLozncttieFi77CSQuqd8aUiaw
X4mGlM+zZWxWrTXCsv802nhV6YTexNSczURsu2An/ED5rAfDftoXiQ2ZPOcXuH30
+CkSh6/6tgiq3BTunqLKiC638zbAemZPZMBf0V1K6A18fReiaU0FrxZlhdHlRhiN
qlSj7HRqV0j/rEiECkPK9TfpVX47Qwa3YaiPFd8ihOsVhgBBtb2N8F8awzs17YoS
7ZnR0ff0cFNePb6Cwg7tYOdeM402UEhvmXxur686CyBHtkpkFzAgh05+AW2bEHxM
s9DEa4ruAuAgn2HqX14tvQ0mr71CnWSjAqRkrLsdbEZe9L+FQi+23X+oxfL13j+O
F1WYyLe2hlx1C0VbA4Maw15+gjL+oQ6wvzDWNvPzawRK+DxT746eGzekUXTI9rCF
09DDnxX9oGj4A2CFpMKqotg4OlGFIDacI9MytyJjsQoJK5GAuojWGmuHAzKO+GFL
D6R2Xnc6DWX/y7bEoI+CibTc0QDcGGT7hGxhXohQVjRepj7wc00UiwOvRG0tJ5Vz
MdP9g2hO2MLq8CBgKmDjZjwAVsU4vz+hFSJoQoZ/VjW8mhyFVaVjH+Zu8XaWQ1KW
nfCliM7tdWuItq3qT1aN7isGpdwj5A9mnkUlvlckYX7XJDVA2OfapgGqjdYRxeTS
FrKcfHJ74SMdZ5hIR1dRDxiDIicoQvSyW2kcuUmfjrlbJutRM55k7qGXMPIjgX8y
+WE2fYlU9yf18MAPZwwVdg==
`protect END_PROTECTED
