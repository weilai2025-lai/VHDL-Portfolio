`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mXfV5XGharfewJYoXdq12d3SzCNOfBJm7oSria5+jvbQGoqzKOgUBACVl8KHesD/
KD24FCSaeQykPMOqEEeC/hEK31v3HSqY11hDE2RMjR45r9S3QdekOdUuYQPNKjWH
eCFPm1ugRAslK4OIDWEFTIFkl06v0MEVfwRD+Li/htwQfcumkZNIQl7gAxVsQkUT
SIVRDpDJVUMAYRJMrZbA7KPOPhHP5WHcO1EUOXijI3pod2QEWcZj+VytjABHXDZf
if+TEqQTpXCi99mZzO4CMmwa9wpJSk/rYcwYy8EjfoRFxy9lZKIUJAnIz8+2zCMd
EPwOlJ3bp+9XBCqA2NUylfnUol5Bf5BiXuiVjU/JwsvRDVs4akVEyiTp3huvopBt
T9iXyTp/QHJ1d2JhvicrczSjM/Z6hirE0gzbssurXjEdXc1MOEKLY233edSRqgLz
+cXd2uq5eY3JQTpiWNar3hQSXu7leFz0aoOcZcvlbJoSsocme5QB6lCgD49sy8J3
H38le5ulEBQ3C65Fv7dseuEIaJDHuYaUI/CI2f/6+YYVivlq3UnJDWEfxBV980j3
y0gCJS/1VU5+F9b5qnDzP+/0qDfNAqgdsTSaP9WjwoWtFFiFxzZL15o7c2DB1TyJ
ZkEfKIfybDpe6zVSVH6e1Rdkii8C3CexRJB9Rh8LL4MbmlNLJROH7IUhKx+WzKKV
L8M1fVEABeRbyz77LXxFIeyS7+Jj1Qs/zvp3Q5PLz2BjWp1LcCzw7R6hz7OVhm6O
Th78/kDre5EAlUd6K9Tmhmj/5hbxfNVP5j7+CYiAUj2ZjGBVAU/Ric41H8jVmBPE
OPHMPn5GX4QsmEDb5XS6CzxEmG45jX0y0QwRGI/3LbTlbwo/TZCgrn5tO2EULdPh
PZ/wuvBqBGZM58zwpc05MRwd3zYLPr4LfYNYHIJscjmp16xntNgy13Ucn5WF04pH
hvPLRP5/hCbNaN1htUI2ItsVi3RdzZ9A1WggCeGp498y8gke4b8xCIrttFZy6mC/
y7bmRHmUjA+31K9/nosgYPCN2Xtx/IG8TmETrn3L1j9eOIR7jJAFbQBdaAvNG+Ip
ltg1wHUzFYmhUMkJy8MZBNHRSy6v5gnT5+dW7E/lc/IARUSqehRhrtIrkWMRbcly
84vO67YDu7+srReB6uonxacmw1SeDZowYkAcNsb73Q9oa0bMScCCG+sMfTFx5Cph
EKj18Lv/+zkyb11+JmVRbnuT2sNAUOjImRT/hbDU+Ao73TI2aBoVa/vfv0pVp9OL
GEzRoktJzbwdvOM59coQkSy00+9vh4C/zL4UMWJOZ8Pko/bZ07S7SWOv1m4a1E+P
A/z051rnd9RLj29hBu9eOziKI1pGfqjIoM5ignULPaaaB6nqOdS/6lKMZ53sEwT0
GOqV3T1QD4pv2Iu/vGQ17HSTUUmHjr6I/w5XJlmTfCGzfYt4/uyrx9+SmUoXJe6J
gncYQp4GzLB2mNCxuGBeKDNeLw8FNeI1l3okB5mKUGhJAs9Fjdh1cokkS3EJkqAa
z+PLm1fn0IQzwNBwfCgvTkXj5cUgLRXZ4sdveHzNXuw9DPG0QMTSFtVSWA8Wdopc
3x/5GPiZC0vmuN/AHOfRnienVOm/uYFfrcX2jrYaoB4USDe3AFZTCj6Xa3xXg4c1
2u6wiWm3yPpiV1nBy9zSWSEX8AWl53/JJL/mVfoUPbk+WOhCfYsZAnpuGt7INYAH
PbzPp8JiCuO5C2DmF6CPXadyIPLCJEB5+XmoWAHUzzdDJaYvYchdJD98dh6C87jQ
g6quODhv8ZK/CnibqZ6HQPvuG4b4YdEmHY1VEPEZ+Klq1YVAAlkNQMsNj2G7qFuj
qCValWR4hlGUAWFceLPXg110fJVleQ9Vkzw2P8FqzOMmg1G78XWFrdybDNkNVYOt
r1ZzBgwrvjXm29WVwrY6KDfiOo1NgFdbSiMG9zI16bhryf8GFOdu7WdG2CgFKPYv
04BSa3naBcUu3mQOa2W10VTcbxc+tnceJezeBZJD9mrCcw23LU/ZHsrdQvVxV2X/
Lb6ptKNHetXSoH5S6TSvm9qFE79aqg4nHgqzkwQG/0H1VPLQDYPP36grhuabZc+5
SU9HWqVv4JlD/tg4UCVVcm1Z+y6KCa3ikdlfxlw6Iq2izPKIbmDQI50GPIlUrrPq
EUAsZN1q9h7iux7EHITjXfJMzJX0pkxqnPqmYKYog798E3bhqLnz3CzZ4Pkbulyc
0rGXAimRqgCWe5wd+uvZD8MTMzzWrcHtCvErHDbkI8OTPjxcZsvEpFh777BK3mD4
zQhySAckqZLtyIO9zJUF6/qtPnwsGgf8tV6y1oHd1aTQPha4A5CUduGS+lgoyaM8
pz2pTFf8vrdZuJV72JzGrtRpsd44HTUpsoHUq/bBkA6Grf+Hbyc3B7ZsdQZmh9mh
YEMk1deqb11w7uGNG4kklonh6n2PkH828tkFxvVTnJUy19h6d62Y6Ge2Le7oIXOp
yQPblTgflNN2hqZnWlqdJ4M7w1KhTdBaYxQNNBIBj9Bs0gWYyOobpdNon0L8g1rm
2dqANphcfhFDOTSLtEsN44B1LH9i+kCNxXMHEgUWCsdwun61Vf6D+QEKNoPkg7aH
Y1ybbx4gBnU9JwTWOuLTK2ysGbfQ6YagUDOZcAL/zVgCbAsxDfOG6ydiAXr3VPm1
G+kXGm5yl1V3b6D+Rpht8UEASzlH0HY3lFIqvlF+ULtVfcNd1Gt4PE0RJtGvmRS4
d2mZy6CZ79bDm9BvGqF14elmHKKOLCdRkPpYmuUgAEzKMm/lDTNP92kiWqfK+dyf
e/ODVfmXovlD9FoskffAYZyiifG3XZdmsqmOACDm1J3EIRQemsuyUQ7adOqs31y0
hJ07WxbX0dQQko3EgSLOR/0OQ5xHXzIS6nY88p0zu8OX/aSgpGCWYyiRWV3ptUDL
q70TTBsg7A/lD3BJwxeKtPsaDxqwPJPxZCagoCNLEXpfSt/l2iGIjxHnwOk/W5Qb
EbgMiIEvIhyvPZwyWTYoe9EGvlXlZiOJwdopvzOFCbZbJxlXM7hjFZR4sqaVccNX
o8ZLBoja7qd4AIG3APsjI6xTIZa/PiYh3teg4jy4Sn6eA0FOkd6hHdKQ4oiRpNC2
dSeflgE/bnj5gclDMzgsdKDvbq7hyo9MFM+nBHOhSrz7lfY4cv8ahDTwCFOj7+3e
jUxDHoeWa/zN5GcHPA8Bwn+CNrnOg5HZppNRN+C0QwzzXTwnshBBCgpF0ktF67tU
lrcCNUCvGRmAe67kgKkzboFOIvL7kM7ipq0rQzXQVVDURqKS1xPIFjzZh5VtxUXl
8b2JRR1KCTJKtKYMhqgrIq+MRs4l38IEwOtgfdomKoycdfBb3EwWr7OfwxMaP8b4
RWkgOS3Hirmjn7xN/cKAr51ajoo8whOQt3UCnf9AF/2JElskVKkbgEiTGC41FjkV
CBPBMtEFBrfoT6zMrGmWhYc53ardMI7zd/Df2SWMTDECyl4XC5BULggB8mLOczXn
OCmnLku3K6kTIFUp5fOep9kfKNtDCvz/RIzcMzcwZiRHFtfKIk4dn2yfNP4DRD7e
8MSkqEG5GSJMJpIY4dqJpLVG0zyScJq7LbT3ec8lrCOcJP2WnY5qUDhnf8TZWVmr
vcc49UYPyhehCBzo00eRCx/LNH7eBD4mHaCQEQzm9Zh0E9eB/STtwyyZ/KWyY7hO
ak9sHbJvDEuqLqIMhp/o5lhG87IBO2wT0BNvLlDX1ru4VFu2t7BI3IsJj6aJTHRj
Db1nD+bX4zaoTm6kKvEgm9/2J5eTC/79LH/knRhawfI3m2lPduh814TEVdYWxMU4
68Sp2Yxse0km2DsJ24qTeH0QvPUfwbdsXxy2ImgaoleMTIuJuXvY+ZsFedM4oumX
KzxRixNiZEXMFhrTf6UpBFogkTF64oqvziFLwW9oUM1KgL6WRXXj61MXVbTD7T/F
HN5JXfYbutVlGnDnTYgwIwRnn1Rr/j72Xd0m8ejV2leQPJ6tknnxEzoWWDuL3Zav
rkDLi+QOWlvu7jpLgdVlGxqUqkT5dOU37COOoKVD9/yKdVuVUuKlzY8TJWK98TvY
fGnFR/O6/dYkwZ64Zo5ifkJWbz1e8ra31xO5Dsu6Em9K1ZMGu/ri5Y3DHXGe56SX
h6dIMKdZsVerRZPk9ZBI8fM4eGj6nH8Jp+lw0QcqF/Sfo7QFu4/efrh7iWFRRo0a
s0pUT85vrU3GZ2NNFA28uggsoY/Pe6NCrfFC53byDKQx0m8fhVus1dgePGUcX2lq
f/Izb9DUVvkEuDGu+MxwUc4TchFT6EZkmlpLD4Jv8PZAItQph6EEQ0HSJhegrsim
tWfsE8Ur3WmIh2STqOy+fuFZheIsDAvLLSkIDvOAfpVBh8Hxv3tIFcg+sqMNpBb6
OKVdE+2Q1g9Lfy2ySWoELD2atZOmexPaDDqZMcJrtuBv3LB4HjHlHgW+OZRv4m1x
zrrT2C7Hqx5fhmSifG+gSKY6mZo2nH5X0aF20WJsJAj5VFpSJfZOjYKtlHMx4xUt
hJBkqunU5J1cjY+q3hE06r/zoNOR6Ncc3qqpaoWuVZNV6k46jR6JcvzD4ORISPRk
FPm/XboHxGmcgJL9JvQr6bIwCshcUTJ36j0TjkcjxV7GJmIU3EkX/pt3tvLuZ/I1
1cTsjoM3zt/GUbsWk7yFxVCE5qfYuj6we01N0+yO2KjzfgHBIxIDVgqxSgunCVKB
tN9OxPV2FqgxK5aadYDAgCAwo/ralvhS/J7jgTP9Tpqxq7bzJilSSE9TTkQH6GZY
HMmn9sdrzMif5TL98hnAYMschJ/krCk487FxZQLfXkNS6vAxwx4kmAifRqXUbnla
Magv4Fi2d3v0IAyCL0XZvfi83zWL9d5LnUlrvrjTeZJCrWcHBOI3k1WbEEvVKaZ3
ziAtXLHSWd/i/BW89tm9XASYDASjH46TidvY0BPqoihQogtpC7Kdoi/R5LKjNs+O
tSC1JxDEDTWy8yhs0EqrR9Bj3p6qnGy9nAbd6Jvi8emTwJweVo/OFw+A5prHSFbH
nUPSHKI2XBqEQ9kwX9K2AM6wc9bQa0hzBSa0gVxq1sExBF/OSetD2j42yiKA8vH0
mB8zwLcyYdFh67WNt30Q28WJrsrDaaziypq+nTGFQNeuZ1ArgZeve4auzxEkfTvx
4BSlrSElS9rmNF02m5tiGk+tlstlsCUHNqcE/w3RO074LGHHf1Y3w80HxgNo/3rf
tfKFUEiMVFrVO7HP1ilmCJThyB+aNLl6F4kwhh3yUNG8emicwt0ad/RQVrmpswZ9
v+x+pWStb2839XWRkJfnIqypNM3d7uS5ZaZDsRLazhucsEb5hun5L+SXlMyYx3JN
CnP/CzYyLRJFWhLjP+GL/CjI8x0UZqH6BJdGT5tYUP4ze1x0/Nxj+w1yC80D9Fkf
5t55fXYHnDw7XdaKIYji5yrYEJ6OD87LrZ1QCeY0AVJsZ7BL6I5m2L+gq4iAfTSi
O53FzK8tl1ZpZacTk42UAwuDwqUsWjCYz3fYbB5A+lretBARKRYvOjFgHOaN0nAx
hBH40DQOQrPHx2ZCJBjk4Dqh9IN0gjk9GVxHo6CKY6kZ0JWppMFvzZxbnXuCgNbo
Ynr2/gR9mGvIlVIPSlmJHJb+7APgOdooKmu8XpSgJOnG25ilu6udNDwY88FGNGh6
jcnOmVzWX8e/bJpB0fMYfHMC8jSmoUI/nxiBgxTL1ijcz949/wb5kgtejkYIdrQ+
Q+cxsHK/fAhhPpzjhux7md9Q5air84Jll9OSmH4jkHQGKLd4LD9EFg1WZGWXF56c
eMaOqU3KZ6cpVQULNOcxhXXcQ6zxL9YuUECa000MgVQl/oi4URnLXf4G2q8wLLAZ
gwU4QdmJnAif7Sm1KlT7ojATqwQKznIsaqPF7J7w0tnOQH+EF2GmscOjY3gayVKL
A9E11eJcQPh0mniMQWJWebSSIwII88PxBcL36zi0u1NTi/onrRgkSf9rkt3avjcG
QRdUrFrMNRrPBh9hvGQJt1kHzxryulZMA1e4POaFcn0q8T7uXEjFyinOH3Coh8SL
o0duzkyXAAgJALVlEIGx1BUaTglnlY83kmW2FWQOD/GOvZhzBcGA00OJHokay3Fw
kQEzeItVQQogqTpXUYFvLSx+B3ahJ+RWlYd293lVJWZwNH1kpO5FgIhVb9IBF9mT
dSaIM8FUWSVSxGd2txEqCQG1lPjcK4pHb1+HrjGTckOwAWqj9s7ORPqisJon+849
WAGqYniPkVwnaFr2Kt1X+aAunxao+Gyrv20/p5JPKa8Q0wQ0embxBveu893KvdAd
/3mLa1MEGP47YoxKpccHLVVRIPlowGavi9fqV5GLVehVGDunAM8oAJx4d8dgh6y9
jxzaGBx6zR7JFLVCwmUho+8BYat1MDdARr0lIGYem8J02S8giLnhXOOh57oErlNY
h/GmeXISnU5/6MGW0tXohLtjFFRGiNrMaJDk/gW6K04OepHoyPHtIMQ5OHlPDSSH
sa1A5M5HsUs3Tn4O8gwkQjoJ6D62hpCEwDu7Q2WWExBCaPAwX04qRxd6Ii+8Hp05
wODunytv8cz37XRQPJi6kIDiG9VBXI7Tftn5wxG+EsNXBegyFz5yglkdWWsR6Cwv
UehVoeiIlSn1wSlTZjHh2XQ1dmfHFEnQhJQO4XIN/Z7C61HKgW1e6NQDUHZ89aa4
omdAEa/HGNsC5k3woaLQl0PmZyFv+CLgW14CWeQKMik1Vlns9oDjquEo0SyrQ2ti
5lU5rcxLKW7yGf06pjfSGtYQVQVc1tV1NZA5csTOZwrvszgWCpcYhG0wVVR32z7s
gyvsdRPkuQT5e6MluzvPwUklyBW27t0Cn/Xk5v6hFbaXGRRRmR5txCXtHXcZQl86
Mjrn3qaA02YE0drc5Va4yH8wgxDkzGEwrwcvEH4kFZ1fi/hw5OtQCu8EtPgfnzAY
gY/9UDAu7DjAjqWzA8Im3Rx3Y2W2wv1Al0vP/2MRmpVx5iieCtMNWIowpiYK4vAw
G3pc5oGKRHFjSeuAT6gEgLzciQmfPuyIKEOLv1CCGZjdv1EeZUMIIU8F63for01/
TKRyT4fHFjPfzhSLh8XgB2ICS6Kl1k0uzrPoQPKv75URedxk/sghdI1plNLVY8Pg
CJBEf7cDPaScFSKA3O3yF8c0LZa+vk672mAKDHVfXZQV1AOmWWx1YvkoEKEHfi+e
fnTFnq4IXdnEOBOzmVr1ezZ87aLbs+qR5W5CTb5VHfcMlOF76DzXxsSiSynECqEh
4GVXL4VidC6uYL+b3z73/QFE600ybfNpdEXmG/m+hmPrCwl245ozeGUwfPfFxKbj
m1JcrQ1BwcEZ9OkgCB46Z7AQ40q6fzs6qnTU6/lKR2StX3NwEANF7BzyMSKoGuJq
qpMCI7PrOnA+GFU8Flm9lyCBuAUCSWnnnZ7LctxnAUiU4zedyUtJKbBcj+oN6L0S
e+jtWsp9EawPq+UErPsU6cT44nzG5XhI3M5gj2va8HNUVcFYtwlVrjJd1dd1Hq4J
lG0yWIaQ51KsHZ5tnZR2rjU00KviBYDCimBVVGnIcyzKj9WI97sLSev7sqO7vBrW
NL2SfgIk+YN0bkambsa3Cb7QFux2jqDAlXZLb18JjwkluqCnLzQ3D7zxg9Uexvdo
8o5X/a3tYqiQ8Ksa4lFZP+fQiuL3gMGpxJ/XqhNc56SRIYGknGzt/J99PK1syf1X
WLkpJ+U+aFE6q4kEt4JWcLc+lEvY7tTNPzo+Kp6m/9xZtXtQEdf5RrrYl3y2Xxbe
0sjvaXOAgM9zHpqRgDdQq8ccyuuEDbmXkP6NHUhYSLn7B1Q6PGArGiYFnCYxT1sJ
MamCAguMEXAhWBt68m/ucTSPSiBbbtwDmlv0j+HSrcm2qsbfmbrlxp7tzxE+2HuZ
eqd1AaWTtSQjh35V4QDA5rh+Mi+3Ikm3pC7+RdZ5ABtxW9qHE66VN9VHEPTEMofM
AO1TPV39x0lskKVvgohuXvDqtG8q/ApToxO3L6awxP3MxoBOiVR9vGSW7l87eX9+
okOGJ1byQa07CYaT5eznkhbkxV4KDPr6Ihg7Fr3x/+h0DACc1VHhpygADHQGFNjO
oV2QPwC7TMaDjYPyYVKhuQA1etOfdEiJRHdceIRprPhUlZglIXCP0xHTmzINjHCs
n1Cdb+0EfdB5fUJ79B3RXoulgX6jtMN+YW/DBTIP+as2yad2MNGNKXSkhYJuS/XH
2rCDrXMn8F3WZxAn2tCHJdRgnAPoU3hruSb3KqHPonLCMuQIcA/YxW6NsE6IrUS3
jqv8aw0O2QXjxU7W6p0dmhFUzYZaTqcXJ979ZtYn/fH5NWKjc1jHnw+FRnXpjdfD
vhmgd9VIQ80Dg0yUlzYageurUc0N5ZEKDaHlDfRHxGFDlkR2OGmw1hxjLs9iivNQ
1hMoi2yebe4IirnGCLnhCXm8eRD8scxRrc4Z5TgBoOhEWqJ0+znw2tHwxs2YXYUJ
X00W41bwnBaXg6NgBrG+hfJjEMBlg2h4UPDIS9a0L3FjYB7FQfqdQ6xy0sh1z4FB
A608iqpNXuIyZD8qZeScLZftSmedyH08Q2NmoamedLDcDn6B+LmVvBUDIzQEknRR
Zdb+fkw+Fvk0A+uGXY6gvM4UgrEnW0NOJcMJ2MxM0zs/zkJ5ZDdpJFD+Xtcyj/u2
CeQYwxtCBRdmBIbmLysGkRoj4IQbgsitW1kAtjksmktZ8lw6mzFNzNuFoHR0q0y6
TKr/50dUizYm9DwgoSaQ6Bp55SUlzRdGZc02SUIgpSWTXFU9Xqd0P8fmEeKS7tUq
bBvYDSkpMDNqWcWAPoUlP0fjJiy2nNrUAFS6+GC622Vzx0o4XufnOhmsqXnX/sw4
uwSrvQRqBw8jjy5yxUITfCTp3+goWHccuBEOQ/fvrFOvg+N8+CRuaigGu1G9ujG3
tbUxbBy+AI1cJ8CVNco5fIg20dQW/A0qiAMkuPLzOeqra6YBXo+ESeQcWIg1QFXe
SYTR/NIxWQuJ+3EZ6S32m2nyhAN4FHLbKkUTnblXJWpTR+wouJ1oK4+uOx8w7N/o
gdMnQjK2tACt5EnF/I1helV8ANugpagW9woaOEpELIdHy7nN48nQPJ503OT0C0WE
rpB4jEQFD99dW6tCq0GszgSiQ+6xL2Du4xJzgOetz3mwJjwVO2yX0YbGa114tUAd
mjEM6CAcDCzZq+QyJrSpqV26Dtr8HZCclXaa6UIU7iz35AD9CPtg3l3jXPBjsN4X
9ccHLlT8VwNw+TPkyEvFaV/c0B4L5m0kESoYNJBzxKzAPgGZ1lt2Efh8qiCl6bbP
OuYGADJB+w1svVNbSTXzsQrmv81sXHEnpEHPkjEEHm8P2QbnURSZWAOGEvMjVgJn
gzyeIJbtqb+d5ioP+70V4j4BtOQYP9Eth5p1aQOljXXe6AZLOEHeaiqy+XBJP4T8
P+Z+NdLT6wkUnMuHmFQEmeB3Pq/QHtdS6sfH62ds0Bznf+fr5UmbkIOrfI0P+9Wp
iT0TkghPuSXsFiT//pTxMGJAkIOuw6UkCepByRRGN9uTwejhGCs/dtFMIrCjQ8T4
1vuNaA/BdO6+cf/Gxpzb+jNSkHDesAqiltFc+zZTvMIUQONjxzvOe4Ix1mfhVF27
AF0039fot6np9+0J5TKe+Ld1IDbCR7BfWeHFEZdXV/G7xA/RVEtCBrgdMltz3NzX
SRgFrz2lWZXAwbRN49lIz1h9JQFWp5+g+0HwoRPCfBjDHUTxTK/YpKJjm2nDr+07
55xUk1OldWB0JxfOIKmzLmQ+paxThYbv7F7oalNJEsqigS+TWxL8ySIithH+sho/
fpGCH7367x8wezXzVNA/NLBPNGn7AuTeIM8xBugUng2D+qZ1K3YkGKYOBjczGHdT
nKXBkRUkEzIovoBELima5rGqJm28t6L6IZO7teaCs0UtUCrmTBOKfAOImFivuuFb
MfJGC9mwM3lESDhLao/bb59T7YrNyFgTYhK1ZbgT68wmx4onQswfUbmQAN2CNvVE
In43KVDBlZR0eycPCuaGAFS8Vg4mFEVxRIYRx8dGIDsSNcujSCnEkYVr7YkQHuT9
toNSzwvyGR0OxQ9TqCUqGL9cFL8G+p5n9NAIi2GVDxP/AcTau4eyhe3p9BywaSj5
VnShq1+xumBSzynPAiqSU8I6xb8DXDD4m3w9UGqHPsEEwaH5qUlcXPRxeyioLFqd
xlpUSo+XZ1cQBVLyOl+yFJ5Wr4wT5BipoHOBZupX2e4j+troH9MHE4SMp6M7duWD
uPnO49pWPKrKoeNNGoc1d2rtraehTcJGB8v7tFAHiZPPO/V/CQaQKBvbcFB1XwdL
IfBzCJJA7XiG5GZthWG761/cypc795CN3ONCW1FP3R/QoL6JGGRa4/I2C0elS56B
b/MY2gRt1KGilaslM9zkKdRMstrc0uMXaiGRL0DXO+wbTly7k/8EfjxSkn/Py8eb
UupeL3jNeiNozyFMeIx5lvx3cpFoSImhxffpOg0LXe1oeJ7v6VH5z3uOq7SwkcqF
UgSRI5fBucMTFDpnEhIMIeaRwegMLHaNIx0OJ0tgHQIrwwiS7juaaBE2Fd+3xMvZ
YhdEpLrbYuMX26PnCWxxrrzWyN5/gslEOrHL/F0Mgkh2dAx+NMZnuhW3HvwT26PH
tSRsrplDnjbsQh4MLY3C+u/5lhEizMoPbsKOa0FPUZYId/m7v3ME7/Gi5OZaWMz0
8G++Aev1RClHZLtD3m/O7Xsz5PRJcSgS1X451BDiq6TW0CL4NcHe/iV11SvtryWw
kAqgIfrwGnNNeEVFMpgKtlfCa4egaqu82Zr+8U1lefs6+9cjp4PG37z48gy3vgme
l2xp8p1pI0rLJ5FiWr5knRyGMxn1G2Re75rNY8x0d1ERjTx5XKYmAY2RI7CRptrh
jjQrF1QquUvIVQYTy8C8+dOFf37yBEtqwy0TM8AxUTLJVJ73moMNCy+ekYvaI1V1
DBdmiTx6HUXtjWMbppzmg9VCwAXyK8BIvOhheJ/YM2wI3mQ2E/1QO0/dlqVihY4T
K49/lOB2VzmgCgwLfvRueEpKGApO/sBwA+TnYeC4+8nFidsQnaJHro3EXbiSlg42
bqH8f9M3CS63xVwx2jSbj5MBfFn8haH5dl2QVZRuMRo8kN5e0CdprFRx2jCAjYsg
rGDTlhuwzsBJTtQ633fV2m684BIU+14xlkj9qliVP1Rt+WIt4jTDAL+F3pLnxV1K
DVVc8Sm7807K9BP4UsBIQ3mN7QhxyFEKaeOrat8DOJbzPUeD0jNHeo+pz0NHmJLZ
gVZuxtY7NqGhstzg7iJCPcC7PtZDwUZmaGmt1fP/lFqTBqdnU4I1TDRvpC0jNYVF
tXiWEAejXEK/AJ1n7yx4XgiSgEFoEcVwoN5ZrAQPQNCgGWngxbB2DmUDMjOkK7j7
zC/sV1pgFx1i1R5+CK8eCeb4pGI6EA/vCpxrTawPsr1qLDeoqTuzl285DOe2YwI/
qUmaD+rxM0FNCN7jUq8xskmz6/Iu6n3MTZWnPjtKQDA0lVHl/C3hKGCw1NyC1cXn
jJCX+1uCpSwZ+BvCaDDjFwOTYgU76BEvPmm3kt5TMYryRnpZPtsFWV31d+SHo9PS
q/QBAZGQ2pcI9Xfu2CqJDMzUSW4Ac2OAmH2Ywmi2Wk2Rsvh1YoYG6P+Yqfok5c2Y
lcSSKwy+mgeV2valX8G5SGl2qlWG/d95G9lITSfLPCOXNZdJ8/DDrbQZIfuGaP4C
QXhcXcpjWVY/3JoTHqLsHK/gUgi2YNGjPcFEVsX+75QniitEqCH/YwqIANM+/2Z7
EUnRU5h5lOYPpitRMADHOf8C6NRH2thLcZ5W7tL80W/nW1IxgU6HU6TPBmM+M8VF
eWX2ViTqdW2qXajRvOZJJwt4vD+egglGtNvBI+0cCBBDTA6MUL7VoIJrOkUG4nsu
d1gE5CQAeI42eLx4RFdADOTa+/oTedhtKm6/YLy0oz7SnlZDrzoYczQRMN7ucJZu
NjXECH+lXYwlqLFCqPdbXKe0ZEFPhfYxTO3a+vvoYMKG7kk4bHnQH+IST02x936Y
0j+B++htH7KecZidg10pfP4IcyvxGF/xJyAVgpKpeX2Jf7z1QaGvnHdKs/PDauhs
zP9OndsyPLyLlFy8TldwFRpPvXpmDheiM/Fhx0DyJgkISBVzxW0fY5vMTbY66DYA
b4dRJhr95O2x9xz0SeCZSB6oZ5kzqFL9a2sQnn1NW7j54Y9bTqi4qY+mMT4XFzDO
kj8m7KM3Bjzc5pBz3/6QCeBB94ySOF8CSqLNtlbiCw6Ah1hOfOk5lUtBE69WrO01
gkubnl77VA8IBc83sljSJaUUYCrtmfNzNLAk5QcFnPCpt8PCz6i+da2Gbpb6Sljc
pcnFwGW6oOfq+0hNMleF78TkZoIosN6YVekzzTaTDcvFXN5AHclLx6uL6eNGAmz1
vM0aToQz9XaIfD4K25NzQeCnbdhuD8apr5RF9Gbh7HVC0l3hsspN/EpeV0AtXP8P
IYwxVjpQ4Diiaag0+zDJ6kPvXrOl2TtEFnHT24g7uRilTerQFQ48PpbYBISOlwlh
yn0pubMZtQbRe4GHCTiAcblNZGsG2XwpefgaDN/uoUA7uABiacSqw6I2ijLybXdV
GUH19GqJCmN9+rn7ZbyoSYtEiFiLJAurkF5u4aKbg6WhOoP0ooF7IcFLV80lxbGw
lN0rNYcEl1kMLDgHeuFIG5HOtKwIhm0YLO8oYVkN1r/+1EjqOZ2M4uYjc6gn8iRW
xml3t3XKVH1KsThJJhKYk12c9skWrifu2uXXTxUrDNd5PqpaXcxSD0j2agWzQh6N
ifjTisvZokG+/aTtlUbcGokL96/u3m0sz6hS57q5/Irp7ePhw4D6JfhCcAQsbSuy
J5UCEf5iqi8KoKltsI62cKsyEd/32ld6ohETdk2dmeU/BPqh3/a/4Iej4QYBBUxp
EdRwtYz7qQx6x6R6+wsMVyQfXVNejoN4oHuBoHjz8tkjsZqcGf2ymfOdfadiJDuA
VDjKKbLd7c4Nwmd709FLALK/X9yk09pV5UJfr9eLugMsm5ScJI0i2sIbZ5RqoovP
xHgp+Dj5lsvL/lwiRuvifBZtOhElsCVeytNmFyHf7iFrfMggcrHmXZXO63886Vde
Q6M+op1ngarucziE/2x2YzI+Uj9LGIR30shluSjiKcKsp4NVfbeEXCbWwE2KJdnx
gdzl4hJ72OuRB2Sl2sMFqpgtrJ9EPi1JiIO/Gcyx+5mV+Rg7jQ5USYVsVP04lCee
AHxgOeGvELjk1O6hGVsapJwmJXMyGPSJd3p+S/Wo4mi8FIjbHuKxh74I6cMF1Stn
IAA0j4g6vVSRa65E8+8ET2ZYdFX+Hngl0UxFBFCJRVzrtxHs0Hl8iqCdevVU6jXz
3/mkG7RNXYCdbmMe1BnlwY7yU/n2M/EAiwaOBwp/hQa07luO9iqpFPUcnXjHnh61
s4fsoRZrqjmEXpg4xwbWf3IPJ3ddPUixDtfvqv8oIlXitG7Hi4wBgbGt6Mi2A331
3T8W5NY38HDq/nkIOjWEQPLFtY/vHZUBTV4Ujzd1vxlrj/BVAKUWMpXMDiZaRZVe
JLKAKVcEYx2mjZF6ivAWxyRvV7Jyui8O3LxinSIoatBuPDyXR26ZIVUVSusMpuqj
DycS/tYyVj0DXiQ/fVYq7RyQqfjG2CmdGS+09bmdNiS1VIQRoB1Wg1cLfF1LzPHX
pfFVfpFrzwheE1+jiMBStDW97P8Qj1hvuJh8qj9gId9iJNq71phe3CAvTdsw/+XD
wgCK+nZSJsT58wOTa0B6AbtCilJrJRdwLRw/dAP75qWmMNPNCR78nTEXeXxPiG8E
d8lsMH5albCkyBAI+hfO/7ntxUWwlPaFimI1fcSVMj3P62Dk1SZviuHMGCcwnnZH
2MLQLU+fxiI3pC44RavAkDknGSXTuILXuOM9Vf91iMWDyqKEf2eBQh5ukkb9na7O
C5K6ymuYtM3ciA0cInLziicVAY4hJGG3TRtsTavMnhZN/Tlnw/jcYR6cNrkPfNN+
gsWhqYqH3gkZC4fNTw9vQYUnV6A7KNqi4sQmxUaNZ2qqnvu5zgjxnNNIjeVpGX27
6RrnoKEbY7L8C9xI20N8CYX02eczDSQFMMVy25emjTg3MguczHLu9clJ/aVlYC5J
ywl0DRsdr2k0E6WfpveYc+brPXCNHU0h8KTe8S9JN8d8K/cA8oNyzG3jD6H+YjHt
Vt4D9qBWN+pIf4wHUYMgP8VkL7zlFMlKokZu+NGYlFqXrHp68GIK8SBgTNBd4mp2
lPaZeQBVJCC8Uviq4bAHwlvv60t3oaw6FZy4EzvoVIaspnDTYS6R0BqkMrtgxWUx
+l2uZ6wzYiRKiftghjaybAMHHuHomS0/Vj6UiaP6tcO3Z6rd2pPcI3Wlcq+iuNzw
aUK0fQU6wt4PKIhGONvKGkpeRfBEZhXNL4YS0uYzRAylgzQLJiYRxJ11mAbjsYyK
X2sR5zzXZp4cedozIFizD70iGLQql5IsSsQ3Xbt2/Y7aRjNKRX4P6wXmUsTYDb73
JZK7xNjvg5ScaQxFer7MkgfW1l98xKUa99sjgqsl/XjK1rIpoHu596Z9ouxo8aQO
vsZsG0jPXnp+nvZHFePfTtRLeHZQsNS1eMQoV+83WBagxycmpHOh7N/FL+ljETwY
GCeBlrEY+ABkirKyRuRjHx3xjzSB1lNVLHlTXq6A1SBUc6bfXNngGRDTNyKDXKEq
VR9ZneoOTSqbQrudPFHaBzUDdVgQBQ4Zdu1qwKOHMv/R2tHkkI8T82sjeFUyUBh1
DvEKF7cgbyOA3lMV5rjEXAsLoDRMWu6lSnyUSKShQ36rQ0ETsTxhStoWyNlqejdH
Vxarp5+0szvxU7nsqANH/GAAO0+w7FF8oyZ8AYEUcbygCPcte5gIT6d2Q+Qpk5ae
r3Lggxai54SFBcMHrCH/n7IzFgmYlF2GJgcbCjZsaE3i7WC2vAzdAlyK2jVbriDt
XI+E7PIluEn/OlT9aZBesuG95pSpTC56TiTR3dNWmhL6BD4Lcs0bOBbSqmpipGKH
OOJ+5GueNyhBAkzHALP4LPEDrEIlTueDnJRTe2s418666RPJOFmdrhIUSmVujq2p
tjwge3wkXA9GebkO/X5q/HzvdQDTVPrWs0eWSxD2yqelrEWEBC7q95Ak84rwf9Me
3fEOvhtZJmhs8l6TCcMmaWFUxqbRh1D5PCmIq4Aj3+Ew66lXCZZaAhv3H88OGn/B
FyiBV3toZP9ecWsG4MPBbft1SonIPOFfWna2JTmtsQI3/lNQ6DkEHr4bAd9bVMOK
zhZhN0Pqtly3BWxnF/KZBIGDPTKQ/CzICfuwQPkbe1G+gSs0wnJXxxSutJaNIHho
0bAMgZkDMN+jNNivVaDiKXanA/lEyvy0q2wl6TIy+MOoPE6tsss/pDK14CaNi4to
hZDLsBmhhKpyiExInRyguFyK+2giCdMGlOc7A9nPlxocde8s6rkH9U9W+dWP81OD
NaUTesqyBV7uVslRWwmlat1v/fEnDGKtpGbVAdAnFUN0IJDyXdOigr8oH4dtl6eH
zfgQXiAuMnsgcaqW3qAiiNoSw8lKjwlvjpYQ/pDdartkGWyratSZ0eT6e5R4HgND
3PEvzr3hIeKTeOaex4Ogi7S9p3SPzIdfELHkHU63q8qZIaXpoifWb5SQIiODdg8Z
MouFrF0ZjH05VeiTedvpiQHraqT7wKYIgJEGsrxn0PsMevDPyC6Er6xkiBxNUzdk
eTzGKNtdnsGHqdko1kwVqM01PH/lRrkwiv4TKMllqzgT5UWohCdNQmLn9gdW5yw8
U2+QHTPaQcD1GII9Bgo4uVNjHXE8zE6AQ/zEzp9QP8DkCFLuhrHFF0QSKike6XAQ
elDn7a6Oh2Y7Oy+0SveIeWzMujoRaoj5iW+K1+a/FRlPAUGu+oZ2SGE8sn83hdNZ
WJT6kWKKQBnEqGoz2qSIL4ystxMNj2ORHb90vsWLyBmG3r8QNHxfegJ7LsRyELeu
eBvBWOZj/mVhTJ6KGr9BpaFJpwTBU8Tje4Atb9j1Fjr8O+vx8FiOzwyDMfotLDKF
t4ja2xf59zMuNmiFHpiJ3lcp53VfZ0rVlBL+/U1V+HragWY4iabUtIGQjPmNgNyY
akfVol3l1SnotWNkhzuo1y8q4tvvq1J5nRUSbBjndQx+vCYGndZZvIh5LIuFIaaB
nXKUYhvQV/is1zHpz/1e6sSfF2zsR5rotHne9y3ifKCxZNokn1JxHbG7VraJ5xVN
AQNRSiKBDdoUh2fq5DBmVK3frqKB/zFvpvKdzLLDw52Ten9PyvLRZQBrgkoegnk/
uG0YeF8xCE+x71oGh4+oGWvsOfcRPn2zDg+MJ1ShxcaVv8uvDs6DsIiNbCN811j1
DzXSNqBW3xiTR5GDrWc4KOWcZZ4s3uqxeJKXMcm+mm+E/ZwXxNC3iSC9FoE8QMFp
O8AToX9lcbqiGJqszGIORYAEAeMIhuupHBKB0aYR8hBvEwmhMZTlVkX17qCPd2ZW
oTp6Gzx9UNTadRgNvhvl1xf/OqptRGmKSZOxPX9nl04YKPizJ5kSZU3JM0J8eGQX
/nhmZSdZtgpwnO32HQ9V9Mtsu4fsz5UP2agADPSPmUNiW0Z0CGMbqiTp9Hac9ajR
+LDmhAcu6L8VdWl9Fph35LE91siNbVWDoPnWvdaD4URegvP0b6arjH7+pCd4FWZy
QtNWIy/dAgeNiO6rHP+rKYdEkFMO3DCzrH41sq/unpxjIUSBd/MW51v90EjzmRIQ
U8d9KKc248b479txvbYqAJFBY8Vb/HHZMukeyivSs72fzfkthcR/m182akZIQxQ6
i2FpuJnxJWPVeoDjeHJAmVISu/H5NLQFilwzfDH+d8alhP6IYx8yb8SAPBgukSWf
kBGMPn5k/CZJsyEpK/Bsu4GrwwaksK8uIdDX92+TiDf9R/9U/RWIydhr4vKMfYtI
SWKxn6xFqXCHybPB/y5BjpZwDtAIBUX1MCv91TJLy+GFAuSgZnEou1y3G+/Qks0d
9kpcmV1Yw0bGJV7QqLUv7dHH76ZnzasHUONyTLqyhLbPtjpNn1y2gCupDIXF/bII
H9eqygWNa3yZ393FezsClmX1MLJV5X8IjJHmwaQn0G+2EIyRqzHbv7+z2YXSUtnk
SNvqvdE/4JyuFKdpmADgfS5h5BMUTcQRezO64MmKfdii9K9wR5JyakmSNHxhffyH
wqKC3PrNkcFcIrwocgpFPTGoDOGslsDVU6xgPTz5aFdtqY4JhLom/ewm+Nh2BKXq
ZEVVYXkT9hAw/Y1DOjQBOt0Dag2ufKXTO/jbjJaXyDr4IripevTqYGpYoKkeOkdk
5WDSQohXXQg5l42enrAE+8GyfVIVIBYETw7MkJRvBsu0/JEgjY2TpGCWesh4tuzR
JrscWAukzHlncAbZXQF++fbpfFOUKPQg8lFO9RlrixFG0ehEriqSW5+r9a6GNtsg
XGn6M8WxB2PLaOufcZkDRVgPnyvlylfp3uUOB9TAmu70wtw9rP3GV0fmiAARXsiy
NumhtBfzvFPEq/DlYlwjHs2cslycXK1cucCUi/arBZnwHHIZGj8U5TBHyUYq6Wbr
1mA1KpMUgwWDSjH4o/Q+Ildg+T4Ro61wg4RZ16RH9GARcX/Wx75tWJLv1ihMC/Q5
WK43ATr0JXumSspOR5C7uwT7hwJrffX5ASdMgftAlmS4rBk/f0y7JN9B4iX3kaNT
t41d9m7sVEN6DMtGDRAgeI1dAiem6IC+LM0lGegYmz8mc049a82rftJk44u8qBvl
oMj6vUocOD58lGxXk7TBvqdD0Qku3ELf8l1DDLUtrDcQU22o5NoYOzk5hjVZKhiQ
33U8uQavuJ+liH6hJYsDfCju0Z8sdPU114rc8bYo7WZhsUoUmB2nKZO00WI3FOaB
gLrzKcsp0Es8izbfrCN8wfSUxZ8NBuBmtQ5WwOwxQe1N1XbPb5/4b5Z5zZbkZghg
UE1f/BMtqvqD5JlaWVLG+D3NuYhxjpqnKu/mgInk6wQqyFklillXGYdHeJdU0+yH
0ZnuFJ065ZLB87ok1Xi1Jh8eY+gkpjowKht5nh7+DlsD9XaGuVS6T4InHfupk9fX
6vNWYXyKaSEWdACp6y5Q0wb90HPFUopniqi9DuMYoQcYcvxxubzxsnwLm6nfK/cw
8L/Y3HDkK4CZ0Ez3C0i7gIoVjIYR+WCCmFOzZeG57kWUSKHSIU4zXQFNJYGisGrK
NESahCDCzbYD22IuJGD8whizG2LdOQ/kVYKBsYkzDDqUY55Es0qd1zJHauSOVwth
qM3HvbwG7h54ypiFLCMsA97YQgYPpurXc2QEUTs+cMYbi6lr/IMYIHED2v3nZHAk
d84KssDoNR3UwaJXs5bOcDpTokHKs8KctwAoaUdOr6DM5NbeKzHRET+T/ik6pV1c
EQ3DkLaURV4EW+OyDbq6Fsebuk1tSFJ+ku6r53SA60mJyrdLnL9GSGgYyg/7yeOL
2ms+cuhPAniFCpaYXYoR3IP042Dm0+4Yrn156rEFWp7exR2Y8PEMy2S6Bf/HfJry
ao7tpBOHcKF7nEOM5q+4p/xAcE7w8kmYsXQce4htu03Iee6xyg0hhqx52ltXxNOZ
bjb7nXvIdoqbbCcBt3mSs0MsiDzpFsvqzol9OkNSmMU9j2vGe+biW/VR5SKpZXDE
gFHMvNCIaRytDbFq+rexGj5Xau5sMUxzcCRzEyy3JAZj6Xo53GOmwr6ktDOmkG3/
wNtq7cb6l3y9ojcGwPvBpwQc0iwidpnha5JOHbsRhw9s8Q7TxpZKJcHuEOxUIWJD
aAKOd2jQxe/LcGmKxhZHsgfGsrmQEMFBC44YoX/6kMfhnZNJCpErjcg3ovGhJQmf
74T3p3t0mY4HAGoO+rG91n0R9F1jnnYyYvi4TvFYlGuJTgow270W4mTubJ9RJc9v
3yYW5F5gNGvufSn4U/zGghupT80Bn3A72ppxfgTxF2zHq63FWYpyeIwYKvU9rvrh
Q/XNpBYf1I34RoPLQnMNycruLFsDBD92o8UMuFddJW1l8wOsFFfKdyfGfcSKpi4t
B9U5P+B9MT0S30mvs7hPx68qGmtFGt10pzZoc1yKusbHoC7F3xVruNmVK4S0QR0j
nCFO64T4IXJjZSq6/dG3WWk63C7wtgvLmUUu4hdsB9tB0nyPWaH0cS/UCpYdKZbI
kLDnkxGnLzEsLnPUqF1HJCkJhJHxsuHKjWDf1YTcVLLCE/8xmm7ZoPMkwTrQP3Zk
znOMT2bLt8gGnJvyvLGTUhSjmsxdr5kzWnZxdpFNKQzEbJEQCfPo7juiv95E1BnV
nC6RNkt77p1M/F0joZjL3B2+McmMm16mEe3CxrprS02+9XyGs4dugW/TZZlnOKVe
9mq6DPo14ezjiFULzdSeiFD/pcyx0rFylX71zf6acCNNjJgGqCZguOyjlKBjbyhV
o+vMMTgUkMMh+vB5R/xIYMtuJ9VuWpbH2MUDtER3lX59/7L4iTtj6McNeKW3ypHb
T2i9U9o6vqCivT+sAUvZquvrX8cXnfL+jjDnSpdU5KevdtqNd2S2Xl3FzgiBwwTQ
p7tptjV3lA/duOo4nYwmYgz8zglr3CMmJcIV4Sg2hJ4p+8Q+gPqUp28kNzBYaXeH
DC95Baq7nhmO3m0I6Djv3tuRkWXF0DrLhG8hh60yww1A54L+ZR3niJETxPBJS9Nv
AGv9Ys7tlSz6LBaZXEt7lmXaen2H6KpywU52E99tdu5y3Hn1/dl5s44Bq1HEYIbX
oWf7WAZaCDYchZUQtwQXp+OTbjiAC5HYLiWfP+3uQ4f4JQB87JFNcVDCJIT/GyJt
ZnXDU5EhgkwlcaYwoRI7b1VGljYGvhssctSYlLLjCxav8Fg+ANND2E8lmAub8hMa
TzkndXlxH/gb4SbnJ2TfwSs5jbMUx6YK5SKFIbN4R3jiEoXBmekTt/kax+mqZjwa
XcvvTYq3q5VyZfUvKfNhCij3YM8r2jdHZyZ3EPRlt4FMIbE3QnZyqehYbB+U4mWZ
5LCn4yNDtUkLgAHJpLj/xhj+snWKrSIDMQ7xaD1CiyWu58EU3bSLaDluPAttVVHC
i/9AKwerU2lM1/H9ynkFu4K2xauKF6Y4rWDTQuHAIGXS34CPzO0+nVbtIQt794QT
KQsxrPdbVukhmWQIPP56KT/D+v5VO6KgHGmaezQ8em13Fjah4XNMKyE2n5SNNXIK
zTEQk8njdEjrcDtA/akNBzJMulbG3QjQ8bsPJ7916bLB+dzqducD76mhGM1QP3u1
viaKrzOjcVRK5lN6bCAN/aKTtmMBGUnbzRgIbV+DZO2bR9KUCJ2rh84bgvqsDjIR
if5VDJIDcky8y2FAe0adWj9UT6H2uT05rrWTohLL2Y3u36s+CveuI90JN4EvKJTp
Z3EOHyCS3837GDFPbRZ7QWoR0HbOBgqThVd+13ifjga5reNdOaUF79uMRu5AEKss
F0Znpkzhhabune2BlXWq6gN4BWfS8BRhD0Ww54QKLxAW52ZMWgkQU5CdflC5NqRL
zeb4RxOiV4X1YnCVGfJUEuRVCdIGUYSPQHALu5ySPtiAleFvVLjy/qHsd4VYVKPm
ru2nmMszip2mv/XgavsGdt/2J7gugdNXOUfZKb9mah6v8W2DIvbLmCizhFsI/J4k
VeuMapqW02J46a2Ugmao1ynKSDKlIV/3hUgkgWe81XFrPhM698QKB2hL7R2I+jeH
nJbxr2OcG/mEAiFe7IKxi1AcPqopsEtqhs3+XfAd0T6Sxm/60CPnFwF4+Il+Ipms
HZJ24V1dqYYNnDpTARICfjUAqB2eZmqg2T4YSiqclFHhGVYTsHFHmjhQuG8zcbTD
iBsrdmOnEw8lSGK3v3ms36a4ALaCoNkFxsCTKBA+qgE/4TjDdY5Z8uI5oFhaYxDQ
UcYj1HEJh2EXIEzKuKod6HVxwlGQNXHvc9h5qc7wjOkVMoGlxp31IIzLaYT8yDxt
dJwAm9xpoQihoSNR9nw2BobFDQrWV0SioGi4fSFbtPWK3dZBKwHyUYr2Pw5NcwCH
X980egVKXGE/UoYbkcRaUdz9i9C3k83wllnnh3x5Lh0RbQJ/9QCu88AzH8CIQQPi
QROfFoQqYy9hsdQEXxGsg3Qhz5KdxDCo17051UGOxXHAHQGMZ9j6Fr+YqzfhBG7Q
aNyTiP/Y0HtTaYoHbDt2nMk8//uE9zXYhrPS6xIdTkKWTzb13GFs/oBzrUr/5yq8
SLvR+sLRvq90XJJwynIU4iqUGNE3hEaRTo345htAKcpY+IAJvwK1pKQMhqOH14bN
H/ZGQp7bkbIxP0pfAN3CWVAvsZ6hD6dwtldpPa2awtDbuMrmZksmfmGCLlS6KcSA
ZFsOuvxGwVrv68u7p/2aX2n6Oqe2ZnpSkfSejWB6uU0rUe7VBmgcD/2zEfh9+VUM
esUHoC9pU5RkVRVblLOgKbRwcdGQpCRrPEgSEd8G5y+D4d0+405FaxDvOX+3ABP1
xiZyRctUwWtZIM2Xf+r5AaZieTsSa1JBIRWTZ5JeFVC98puDNLYtEVy5fdQppS5H
bit+jn77+sva/MDMMuAPmguU82JvO4mtqxpVpMVYcwybkSdPQsXZ70mjuDP1F9Op
w+Z48nhWit1QT1rMS3oos2GwoheI0qP/oN6RLhCbMOl2CS4GHN49Ff9vqMgpXMMv
i/pUNJFTRD737iaI3/zMDuRNkX9eJjyTb7Nr1hv/aUfTE4n3FxMpP0cgelts9687
5ldDm57GO9Xyqq6UuQErnBvWFkhyiiO5JKM5FAqlLMBFnLwKWZDOmqhtKNNJxcLC
r3a6qgByiT15WQ0P8VVVuAirvfMr5kRXxabPVKgFbMpDDpyuHxo8A7RmQ4/BPP/5
sk3yr7RYlVJ+c8XSkqf4LEoi1IsVXcl0l+zloQ2PUqQzP2jMX35p0K0Tf1xaYhXY
vavIcvLOFokOE8Z4z/O0l0XxbpaXjw6sGVhPAFw0Q1mlVpV6KY8Gg+IvMwyOpnK4
SJ6TOgbhKsiZmAjk1T+0vmSCnsLevMTm484vg53eNxpY0qQ/YooknBOPJ2BA3fw7
6hRNMP90l7Rr/ezW3SMyQ8qRxwixNgcAcd9kMkfYFiAiBehtBqceT5rn1N/mNoud
38WYxE1Dcd4OY9JjzBgNydD6GOmwgGKdQMZ/FZh8ws2hpKuXoXHKrWK4sNkCAe1X
Nxw+Qze3eQxlt/B07whvps/n+IreeF+tfJH4qOXSJ4/jrARDkpBs1xdvCu4+rlxe
bb+rzOq5Mcp0wtqifirqqP5Dm2ZsbeoPBwi9ET7es7VjmCKlPTDDF8ZjY0+Xz3HI
oEMN9GSoGguxN513cIocqmcZ6nlXCRMzcBsomHwcr4fKFh8KJWwfkKSUjh6GtJV8
ZPS/WgcFaCXdlXiIFj8HpiqXtnmwh8IstjvAT0ZuX+SuNVkzUSoCwjfXiwtg2o0v
hzk/PXrafC1CBzhZIPuIWzO/g39dO5sPfxPTZgY6n54287sJ7lz2o34d9rznxLZg
X0DxXdk8Grd1BfdFN9dfUoBdfgFcDhHi9UD4boWLcCda26GozQ9ss55Mfse5jqCK
otElLzbbGwws/1kYK9wtMe41dVasOTYyYdI/c6HmCedDLHqSl6R7uXmlrP5rtuKL
KGiHYwgJKiqbxt3HkXEjoNjdSjlqnpg2rrNLlVuBbbOnLFEKtEhS+Faps+s9MEaD
m9FLMOXETSYOWfYgIL9DfwHyba8cvdWJ4QvPO7nio9EY5ACcAsVTC86GwcG9/2wZ
jfVNhFyJCBE00ed8pDlFnwcjTdeMI/42/tJ56ifkU79kgIGZ84gdnDwGyTRchzfw
v2cNkuTkkzcLSKx/FReu03P3PBybUoiNbsQd29fYWnQkoaHmQVVniNK2ivlPuttN
Lu1tYO72XSZXhKxBGraoIEJ9ifcp+nPH14ITgxN9Ofozs0Sirv2yhBF/CMSXs5KB
65dGa3xrewfDc6y6J5iSGoURQC8xbE6CmGhiR/6Iy6nULaGeHYjABGUj+NQNt08F
AClqLuAiKTSigjFC63bZ+kpqyPpxAemDn4YU4MDdZgcuwzrkfYQp7Fg9HZtPVcY8
uttQ8d6aPKrSngi44ubQCvlBi3HNatX+Lh0jtZU39U1WSjgeJEPbOM3Ff1wI4Yl2
HKCRCnxZPelOc4zDoncJ8sJ7DIWkAbFq+fEtC/7PDC3I7FFHdgG2sUyoEqD1g6ed
gBcCL9cm/YDAppxhNnQO8NcYRrNF76kJqCvi8j9gt+3Nq0Gtp4mFZ0URXdiGvHP6
NbA94B6jecaj07joPC8Cn5b4KF9tLmarb4H81gXUzCdwCYv4YV/YIQjnMtJKwoiQ
plRfPeIzbq3FyaFX+0A5HpKG8j3kJlVU4fovTpFBLR/jYLLtoUwUHjz7/1hFid8q
63BDsL2J6456vdfF3Deo+UqyMfdyH7ltBPrsbGKkIDzqPo14l1PbYtisn/B9aWVY
zySINs+Vq3CaKw7no5V7XTw27iT5iVtMmKeFkw/I9n9tBEv+TZuCghwm2J3yJWZX
+v8lr3ZHFwregtv7s5fJ3QBgaE6gow6fN1j54PcGBP5UsPw0/ch4V8vL2H/Pp3e1
IyketeCosFRAynLjDPsxV+vnIRSlkJwbsJ7/QAiaF9whn6kC8wEzEy897UUW8ZoR
XKijxvedo4Mmer/3HeiOrAoV16D/rTXLsr1GCIxtM9QmJAP6mfywZMXsozculxs/
0qhfDLYN5PGfmfgymGnm4oK6qERhRff8ZjoKpJVSD2cmiAh9T66axZ6zU2xT4erX
JxIxPge2K06z+Nv+iwlOuZwrOMCmY+jFPyBd1tDmpSfbS3jXwzuPuBEX22obXdws
Qq0Wfj8LCKJk7AB/oUSZCCV7RE1zlzh6BN07LXyqrxKNLq3PiZHRe6CsrGrjhZrd
kgsVAdyw/aXx+afTqkM9YFoiuyHaOAWIkLKdipYTDQmZ+WCu7xlV3jAQvPkM+ODa
OZwrIZ/DupMUi2l3n3CCEASonYM8Nd0fToLwn0XsFiOWdTNXjqkF+KumjY+wlgNz
xpmld8h8ZrpNOdZ7aikWyu7rGIuMyXs5uAAsm8iIx/adA/H0SKOQXmuqTg0AQvni
XwvOFisT8o07j+S2wCNsiHG90/IMXPEvEZVlUPB3n7Bxt589BdqHqMN16ERyX5GX
Q8/u5OHx8Yf8e1nFd7Rx6y+0Ha+G2S3sUx560NSQHxzuO9fvKiff1ADK5e2QkXV/
g+dD9tau/GBX0ZVi4IcVSgcqXv8DXNRDEF08uqSeGCLEXSlfU5NEpxfA0DIoyyJC
vz+Aqe/2p0Ffz0f8Z57tA7fXxcyMXBjohm2hlWOkn6LPg6RufSYsNBOI3Mq+cnFe
hZylrxSPWSbYEj15+w1gxUc+03cUE0ZacpRXx+WheJfaNYJfHNZ/HTNWADjB3kmL
moLlUew+lS6SoRHHWfpOf8DpwkId9uD3CRpcDYhC7waLCjaSt2ZPnR1Q6qzCbF+X
mgbPiBtkubi6bYk4R520og0lKklAwp15sq/C+plE9KIButwrzNF3jv0TC6bTmyC7
DuNE439GHBrSvcII5e960AWlfc8yWjy94MlhroTXwe67P3p5y9XnJ8GABiwJwHPO
2IgcBiqxKyjpvQl23f8EiYm3+jCOK2F2m5gDcN807MVAORd2fTgfi1d233AcYs2H
oG/2ShasiMKMlJiKSvyl2WvcLnxN9seSAojTDD3lIDWEARtf5ko6egCNeRMOTYaw
yw5kTASt5TktejT0g0VHliLeI1FDx0LmnjnYS5cfUEE5a1G/61QHpapipdt0oMJG
aNKGKnIwBy0TJGMr1sg5N7Af3JR5NL9gA7Zl7bHi1RNDesYe7K2/CO2YC6mU++w7
JuXaRWSVwrqetfM2fGxX5/2c0BRpI6jPJpo1MP3l2QK/pR0apEs3JjDRKzYJrrrt
LXMbzz5bfZcGvdJ7hVemdHUOHMovXW7ZCk0HJXQMU9ULQvlAzcT3j8bLJcuQ3wrO
ChU8gdPESgJA3J/72bZDx9SubuGcweu7d9dz4g5tlsMDRLPBuGNYq0JiWQKkapHO
A/CAlxE3ndLHrrK2uDfyswIPWj0rIveTahBNR/rjUKyZpzgbd4RTqgMIa8Yzqtdz
50Vn4uYTe1RKZlXKsCxs0zgs3RfrzHiEPthGeGW3XF3b8oADUHVb4IzufIpBRk0D
m1X0BKwfsTqh65hQCHXwaGEriIlJ6YrWeGvrkHJ0y9fXSoR7b3QuAeOWBPSV0Sz4
JLMXczGe3gyAhFGIXS3rKPOyV1+ULn3t8U6RV8imrfNVXDup+gMUWj1MJMp8vkNP
ct0hkSiSEYe2wOYUE5AgBviOxTSMQLPAv0GN2gosbNZheR8XGFPAs9iQAHm0t8B5
uzCXCW6xX5ZOwTrq3U7BRZehxzwKa14w/2yZ/nq9mtTYbchEFY0E7wBpPZAlyBGQ
f70lNj6DRBqcJVhcD8UbncOWbCjajLs6/CdBActp2MgQgE2c2HseYmQA9BwcIQDK
4JI3IxtH1l5cNKsZSFnacY/QAFbidD0jOf/lrtPOsSxW2zw3ZVg2xV2fKHJe6w+i
clQcytlK151VynHdd/JsdPQLb7UQF72S+ceHMPCcQaIxRYSHngLaCAtXfhjpuCBF
LQ5o0lo+ZSSAQakgpGLrX9uuwO/EOSdvGhZMD6ZIs66312MhmlI1n7DDWRzV7XGM
10Tc49fJsHzILDXN8v96zdqWW6afK35KAYSUTC3xMsyO0BKiwybeTGUPKf4TQTs6
CxrdZUhOV1ZKXyBcDCes0i31tR6x76NPJhiokd5TUizVnptP6Sj9bORcVQ6TgwL7
bOdz4kMQBhZQdJ+DmhVclGjHLM3S3KR6ikBRShmoDLQ7rgCvMrPs/+yAbzIeO6zX
aPOTyo48Ictp1zfBRQfGSiwk7Pvh9f+o/sdSjYhOKPYADtketki06HQLN5QCHkG/
E7cI67Car6G8rS8KIsxPjW9Jzj4na60YMbXgqIKiDdZ0GNXMoX870E+Z/b8Q2ZgA
1ie2L4dD9v1DMoh636XCZaX21E38wYwRwI+fuZZnRNLheup3OBwFoepD3/fiYUAi
KZOlbYH4wkquDRAMeC3cX+taDmG5bJ2YutL/b55eWIn+kXFrrrOYAt16fSULqDlC
hZ3nqu4ptrE4hx08819QBBouXU/qTGxe/K9At3i5tqZQXMl7mLae7Zm+j3RJaIua
mbPN67EVJdEeF5bHO8tN412aIrIatQgq8AEfZjVatRQyLhNsJJBWeMwM3jHae6lT
fmrkBdklcU+SMkm7v9QocJ4gV4yWIHPNpCL7PwekNJCjwuVRLHFWNY0OZu1GxPlN
o8ec3G9+k9/OsLasujAzPT95SyzFw8FnJ1r0HFvMMq2+wihs6hPGaoaahFbwjAsK
jkIgmykHIA8n8eVLmy4tGb8CbvXlkjMWX3QkyrXnqdIuU04dXHz154Hj862OXy5K
yyJNLwq+p3pJN2Mv+SZCRm0Mv1icPWdcbZC6hABwfXVsHdBjfKvvjttdOLJ3DKSg
Ua/uAcWBsZKHN54RVxurMGHK8tWfvld4X7qjrcTitoM5Z+Ab8eEbc0iHvYK1Wuk9
FnUasRmwy3H2sWInK+AvRb9NRzENEExQdF+ve7h5uNaIA87B+Ybr3afo4bn/F6Wy
d+HYEmXokMPsBJdM3MyQ7blqSV/ulGVPx6fZIt51n31T6el1ykIUwgZ4RC4BGuBj
wzhrrVQ5Y62X0ISAx7lyr9CMn0H7989tvSDgTigJ2NHy6dOiiVRuCpN4dDCEl+JW
UmUmwMqV2fTdZSi1OhJEEHiuuru26fnyyL8aamek7DRnw/jbPN7F99/MMCi08hSe
AtX2nLomKYc68ZKk8DNfHEw3wmj4QFWQZjKEUV22/3jTV7l50HVDLfWNi8k4byBG
9ZH7Fk0X9SJvICWp+3U0CrmyivT6MRxmmSmuV7rpo3+fA4y8WAitZcy7kJnErCTq
uhnmZlJHVs9KEDzHdkT526oKSlHRyrj5kwI1CxaWE41jffALsO/MJfQ37WEeYJ0+
xolXdzNRsJpkK+stAbdFdqepd4KqEifudbGSh8Ut0mtD1dsrl7KnMMXL11NL8dX9
ieYztzwPxS3uw9TZDbNG22rXDHar4DqhEoGJOIsbKAyGg5L08U9clHX9ZNKHwU8V
0bEfyQlYqrliX6dSXrSwjYNmkpjSkLD4mEcVp0r8NxDXAVeboeJXHqcdCeIVg5Ot
OEHc/ufyjnhWVEscjoYVzJ49xHeKROeWHVgZZv46eHRqx56OozVGSk8bEejfQm+z
Ke6vERpMkojYdzyt/jwVmS4A1zRp7EhfqQDLNV+73PHi/mDTtGUiXL6E6LKC56UG
n4wTLiw0UT5FJ1dJ+Mqj6IREiEPCIDHlLotHD9od8hCAL9y7nr54gu8b0ZDUKQvj
ZjixsX8Qdz9EFiz3eP6yMJKyWN22X/EeIiJkzIkcpO6tW1wcdZww4hBSytiwVPqv
e80ROpnh/yN/ITu1rSDpuwDEM1UBXRmPuC7yrA2/SB7qRxcbUUyQECc5K6OvWEoZ
3WHVuWH4IKXXBXmVCH9axQvvJW6WPQDeZw6fhxXvPl2fIvxZ5UQQZ0o40jlONfMO
nQvKeWE0e7EtxRSnswyPNk1uTMtbfqNUKqJzfmiHd25U8FaEg5b/EuXD+quwpeYY
BrXwc/jggg77oIBBEqW4POWv1BYzdmNl9meK7Op4UGddx3gWN7e40Q3RBb2yWXFy
yIxQjah+3mnmjm0Yyq9W0T8GjG891OrNTH3Css+vX8stHIZIosGo1JmJtX3CMDFK
Niej1ubM/aS8ma/+Xa6XIU9sIGqqZmjRHCT7ERI3wsWSRIapCwOejF3HgAMaSLmB
J///oYItw33ugwMkN6f8zF2Pjsr2vx+LadqhMszt5LTF4qdjtQbNVqVPgqLeMwQn
YGwowAB/N1CLL0JETURaWAUvlkLytddvX3waDsElcz956nrrWdEQxuWknU1l6XBB
/3VZJ5XUR7x7Jf1F5dY0ADp0ybUuNB36S+I+gUJJFal3GmJPAP9l6lKSdpbp49bG
cuMbBTCVHJKTNMzpFyRumU2iTR5lsGM68kprYSyjfKVRBzo4dsfFoUXUWGG46Hb0
DYZSJtvk6c3YCMtTxls4eypOAYjmRpABxoPUUjQOLL62ZOmN90BKeiUkh9IIu/uP
kqQovYnTaXBUg6rUop719KVrM+qco6d9gGZgGaH+fD1bN6FHYcSsVIFC3J52AZlM
Voc83sLfDV6gyVTAF5R0D8W5M65XU01ba+pxcnNmKzWVWBUe04wmH+UA/AsPFHZu
NWYJzYoKfs4ZbYhb3yaxj/ZkGNT3PHyy/9AP1XSKPnb8GRc31phM464igASx9vyu
L6qyE/DoxNUugrjO3sOBprnkFHyjndFVqes7+McBfp/QRyxDxEaGwlNMz6biAp2R
20Fc4a+R4aWyN6q3pUa9vjXHXknRuGbQKP5VZQEG6Sja28o9YniJ8SOBp2Eq0E2l
ZJmbKzLBI196VkRpQ2yqvI/nakZ3lTNFLGi3MlfCPJ+7QeqeCKTTNHubGWmzIp/i
wNKWb4wupaowVH8J7a0NhXg2x70o4wa2ZqIzobN0qbWVcyjDfjXX27RV+KX3iiG8
z+KcOjBgl0eXrNpv7OhxGVbJGRhuFVNLYqFyLqi3CrKw13SMAX5EKXIRAXwYZGuq
abiFhaQXFdgUspRiUKr425sRRYhfDss8aXZu3Rh3FEz4Gfr8SA7zVqopr0kMJPOn
JcJg0C2IZLmOQWO9yBcoIG5dUDzrAO6nvqppvpyZa27Zc4/ITK8F0cvqd0vMMCrH
VK+FjlFF78KV1gmkiG/rfR0mjQDieINqvN20wa5AK4Rg+CM/Lq/gDnU20AoP2UTq
y7mZIyPjXMhbZ6jEdogARACb/HU6xEcARPgamkG+/H/CaPh8AUvdPQxTMnAW+lMJ
xhxHU5m6SPSB15c4XLDvxcQaUhVbfgBoxtDOCl/yY6IyK53nWZB/0qmpj51TNDmz
U4wvmVVBah9eD9vwA7Gs6FxL4n21OBYWK7d8ifCJ00ey4b5AMhPwujdKwFY6dQhh
a4nE2mEC713qa73lzxpBlBoX6RlXUPFTrnodjZtBl/AGuJ4JXqRVLVpp4Q7sPBei
uAQCgcD80/A4zBQTzQKeugKV/Jfu+/BxK60EDm73Z0ZGzCDfxMR8/a/VWBmzBCKv
tXHKrdkNkRWDJve4OwICMJrE/yj/EEBBoBJEpRQUYji0Ux9iRWVacOVOkzgz4cJ8
QW8b2DnmH18u8H7H5li2KrKqH6JaQTXIzWg6QHxixIwgZe7pdDjqMV+BUofjKqWv
KIOKRfme5oyZpkcOX4Drh+s68Gwd6JPKfqJoo7d8wLL3N134YTj5pHiPz7Gs4ld+
ySnxpTCjCsqyIBAiklNy+9HA4fCJxPZVTxNz9Rz8Vi+FNSbPg+JA/EMLySxh+gyg
BHa23OBZ91w2DpE4NcnOmUuCJnvAKoEoS+Z2jvSN5z57HhHjIsVyB1xl3ntg9niO
0ZjWhYN4/t+amtKPzXcYFWEydoXl3vCEeY0Rr5eAkoHP3/U7u++/kR4vMHa4i4YK
WqHTxKnpMq3Oxk73Awq05/M65ghXFg0cI1P2HQUd0lBvG31AShZSKVtEQCOqJClc
/3cYoW0Ryj3yO2sZxGyZtFvyMtAWkm54ggVYWXWqYTAAQSCL6ROcPwFgTYrdnurs
1B/vvUoUXiIUyPMQNwiOk8udl941fU30wtrJ0DMsbdvH9GwkgIYZx/f5adU0q4Oe
hh7HTo0EoFDQdq714YkkaKpylGqqEgZDpNYKQ2zXzTLs40r6CR8hnJKez8CNtjvX
nKDBEENBFJCEXRccAHZURAFyKf34QFmb2mYWQCdvtkTZhfqFdd9wiLEZy4kjD9Vj
3eqVs56Xv2PQCQKXJCtO5LMqAldt1+U2dTMuBN4RrhEY+07RNKnPhOhgN6y4omfH
OU0zxl/7GZ1BhWBBo//ALszuHnCvPgwXW5kK0LZ8wdRDAQ6PwWLfI8oLQFVlM6pg
mzNHs0j0Amv7B6IloROS3H9j9mgqQxBMijxsVqrTSRYYM2KjPE02L2xlaTy1rWmY
t0509hRdPsKJc+KQYQ/gSEIoj6ARfXFahi9/bKyhweKl6QjTA8viD9c1dgWeTQvW
V5z1wyvwiXV2eKflXp0dim0Xc1mf+J2PvJ5w/Dm65yAu4nIJXa+rDuNQ3O1AQP1x
IBcCvR7TvYGie+uzISwbLM2N1QOUueJ0fmrhQ/93B53BiMb1Ka9ma89vKeuNCEdz
AWzXqvL9sJTU550Ok2PJcPNeIixzrLV/RhimjBzGkQwt/DampuAuxHvGePdSM5LB
WzXeQjYxNMQ5yobwVkn8F3okFBl/PrIh88pj74k4bzQFzs25aUtlqYGXyLlQw4YX
wLowY1fTdztb2N7g8R8e2M+ihOSkfzL/S3Un/gdjCaFTl+Oja8+ay0C3Sc/AtZm+
EG6bF5nJ4HCw+kmaenO0he/iHbOuyUKhN+2zF0sBrk5GDfVQWl9Wt9wnscFFsrR+
0xBuTeiisJ8271IrxBLBl+YX+BKjNnZhYhw3uwfiTxWfMYTjjL/6AT771bI0FOTM
gVegadMtBZuLm0awnYHCqVN3HYGnA+rMX4+1zqGzC2gLMPDaJNeYUD4ZRDlGg8yC
wPz/VHFzqoM3GV33XgAOjZU/mCjzIYBykk0CTD9HlgZvb7DSugG4xcuIW3c3zVAF
+CPxUCQr2RoPLmuaS/IGcX+OxzlRQanC2vK6bnYYNIk9HE9fufW8vkxaI0HMfri0
z190yFce9zTyXxuscLXu421CHPNuANzBTaCFUX/z3yMb6PwdrP+LPyCxfWKYMBMv
7XTs6liAATeo50Hw9dHN1uysh5N8nUccHMC0feQKTRBk4NFvc8p7cKE+TESY04df
uA8xJ+bhwdoKpXvChwPzqdREsTdKMyElsudpnpPVMnHVEhSHRGqurTWYL6GKmXty
8vrvNJ6AUf5iizD6oHTTG6fHehQX48eXoRgUciYL2HcsceNZxBbsIrmOaCh/U6Rf
2rDp0UtSnegI2kdi0dHSQ1C4A1huLiWpjTVr5tLoWTvvglR6G3288Zmzn4B36XwA
l0FJF5gFj02+ZDFWCO1ECWDHL5L6FxHl3YmNUhOgVVJYuPV0o8G415WwJc6IBhWM
23OWEsltHuafnessGy/Rhq2zdWbXKX69UB4/BAeiJ4vdTOs3Qs9iSxlHvdPNGUda
KPYQ29awCHbK9lnd1U3fq0Rk4JOvKOBsSb3mNI2ISf0rhQIAOuUaR3zlOZFkXzih
emR2xREk2BV+zQA3OURSf5eKkCOeH0Z6Okaox3uH5kW36HFeR4cfy/+eOYJWrFtX
5jznMEU/yU+F8XHsh33fmA0lv6/x/JtfM7j2j54aFAcXUHxOT+jUOrb2FdK39hGC
FMawTwdv5NfR/oLIOP3cPM3F3EPpyIVbWB+wguxmMROkrUGdkfuH3ukQt62Z+sEt
/j8R9FYJcLzr53tcfNEUTFd4psKjOKaO4vxMlozAO1O9w6gjx2z0Zl5QdSMaZa7n
31WMwjRpKvENwV2A91HFJ9N6EFHgPYD8fsCwrKJDtk4KqwOciY5s1TaruJCVv170
/htPxI05iinR6j5w1b4BzBl9NCeeYMCLlRHwxco4+za3NKmzz8DkjXfgPVdNBvy0
EC6NI6QS8KAe3mxdLKeM0F0JBPGyZmEA/aiTIv8ZMJ+7vJRExciVgSOWhA5Dkh+B
68iOn4yu8VdpyHl3Sh5IrTM8bhtC5GOYDHvrNZTtoSqTgZl1P+caxssItan+Assb
gGbtA0/q7xu9CV5I0rr5X7AmWNYbEsPvQu5A2o/o7fjU/ItyN8dCzLpzHOASMT3v
8duMEyPtCngOoHuAfoKIllIZ0zBVbsY8ml4fGAK+fMbXPQV2u9Wkcxy+Zjd7L8c1
pHMzBpvfcFpsW8HDMKFkU+xAKYFV0ZjnSChbZVn6LAz9oKbLAyusPauFSMKNY6zI
ZsWyHzlLuKOYA7FfGU6ejr/J1RHQCmnfYddumaMyO+o47bL77jq/ZM32LlGHKn0o
08fFRoOOuJVGZKtSLe5k91qNjnGuDVh9NoZwIZVIYDMX9UirApJYIFKR+LkS8TtW
hs8A0F3+udzohcd09teJDwPmaMrT/H3GB37BCb/0Be1wzaWcsP0YQowy17QVqA9D
TBolIu/yqkvqR2WR9vzYyeXjdqB28DPW32kQuIyVECDZh1Yxw41cIA7gls2obn4a
WLxKOXElwCVLcYQLspuMUvX8NulooE3upTOJVzeHwqy1tL45Y/HHq/emY91e1RQl
qpn3zR2oj+1qAZ0cDj8AyTcy7Q1q1l3hJNuQXNWUgzyS9g3unl4KVxQjqCAy3LDI
yB+zHl/boFxRnO7TD1FPValfY8dXjbbTW3XCyPvrR/iMe2hTCRvkIbP56otaAvu6
GOwrvihI/BsQfi1xwEl9rr7Yxzib8dp2G4OQ82mZfoZbBSCW3+jCWKwcD6NaNld0
I3zylFdOMTTiaTKXgTHCVn4ZU0P1So6VXGyo0tcvFxzz3rUe2tPhz5w9eij7Zepw
VO6Bs5EqR8Wo50rDsQtzQViFtVtZHrTtFYRDaEkAKRAHsjTPKj/RHBXZVYG9IwvD
U/JvttCxEcYEkwy6IapvI48VOMCwvJSukI4GLhRIY0NyK0B5DkoRzyFX/FlmeIlM
T7Dt5K+DHKjEDe+zJJIhL63yqkete9PaL2r8cGqKk92FkQeoXkrrEoKDt81JJlVA
4fIbMx/H7QXWiulZ40WkvPaGgzmcUVCXxp+Ax6lBtnovGL6UR4I7lH5+V7nFpKl6
B7LB1NcMEhDKCxKCoHEA42FE0OJfx2g7UW0IVexAutEocqEqi+YatY46LxJvZEpX
pB/KRhwYZIyzBMxjD47PhnHm7g20PYBzjG/ftVD0qbcs0RNI+NX7EHxYnWKCkIKn
9MWe2VT8YmMf2sWMwEzCNosXetrfibyuJKHfRXlAMBcnLwviEJan+6q7Fy9LA2Sf
J+RtAvfdf8xdjm5136uCGXwlgfAa57YT1bIwC2ictpifn88pJwkTIJahzpG3KFlB
v3x4XBcUlrv/K55LdLbbqjiKSx+jTX1xQR0MaA7YVd457M5xhIxOW5KagpkYYnzK
Hbw7ba4gi9FwZm8L9nFaI13byp5iqPSklUXCFY98+XgZB5JNImNGmRsDRqTJ7HUV
hkQtupeG4IekNZGM7BtnftrVCeS12tR2n0zI3+ZuxN5YUftM+JnS1rUkko9HQLg9
btBrsKJePPx4Zsnt+BN51VwGEVMijgRU/eDDDfOonqQTtZsuUHqO0mYlPzRaaz/K
IjOesi2lzKwaE176aBjmMb4qxi2saOsVTKvdR59erdnAcTnIN8Y/m49bgTpT/PEW
TSEB9Cf6wNTGTwnRfDt1bRoh1xTMwfS/O59/t/PZK+SpuiUrX/irSfraN68sig5X
P64cL1Ni9ySbOYL7IiSdfnhqTD5XvRxidDQ0BPCkbGELNGDRw4JUSX97nSlf3SBG
1su+yn17mlW5QamXjfDJxS1yhYb7hXTgWp68LndLKX5ZdTSP1Tz1LWJARU+RYUJr
V7AIARvE/KNXpm4P4BqaxH8m0fE1JumbZ1RYf7eQl9A2SUwP+At7ewEo5zFuy3Yi
Y4KBQSPBAiXHmixdhyfPX3NB/e60tpFxpHEgCxz2j7UTk3XK9M7fqQSN32exyFCt
adTOPXMaK2ouizyJEjjey20LbJlWo/DWagg8d4e0T/eiiQ6vJM/njhBB5NC2MXSE
0bMApB7WbhEs8i2qxtrn7nNqCLgvAVSxSz1Uc2f+gmrfPWEROUvt8MRaRNXWOzAE
JRbfoVx4Xw8MUlCma5Cb61cTVWuVJ5dlpYFt5hQnR3d99wjQfnWKbcxlAuCV9HXq
hf0P94L1JDmoCkX2cUxrIJGTRGjjeJ9BEJ/thpgp39QOUNjvFGaVv9MeXPUfv8bq
pxzYCVmriIt4KviiuoQZebA8mg/g7VL0RpU2AWjF60A6XJ2C78mDjJ4Lk4IRcpJf
28laYGyjWgzxpGPlFyjs++qMLHA/wFvcbn4fN5WZuD0hIsYBrtx1FavWPeW8q4Vk
KawjcSjN/TeOIKPrSJRCtY/FMr+czzajumbY+M9aK8nLZMgdISHkyKrd9kK2o2PM
DhoxCEgRLvPZp8hJE2OnMm3QNjSv/Uxogqxj84W5kWOfzHklzrv3komMsy6gWIIQ
Mr8PRwnQHXjMFz5Qw6VNrf41KUbiiZHcIipOxkZidZx/h0FXDEe6catdhsQt86wT
/zoMoCsHJoqmHTCHV09EmYf7FvuqL2ivVYYvOfWlmgJHDmohkYsYpIxxJciTdcaG
tGTIqHz2mRDxiveM5bhIVPT1ln70uSbwuuC+bwIHnzioxrnFk8umyQvlWAtSGs2P
imLKmbKdsGJ4WEn120sNf6Sc5uazKypKjqyN/ah5OlMbkYXSpiewq5nz6UZMTv4u
0ktWF1KYBoGHMSosRwp1Mqj4MOxdAmFAdcUxBbRMGPAuJYyZYQ0Iu+EijPmX63v0
H+857z4qGdcX+NCQmY7NVRqW6MTjhzR5QEFQQBz5G7UF17Gqlwvu6feCuLvqCc+c
imZYiHrt1zHvKt1DmrlEsqQVVRYm8EfLiLN0DxVvHLCAmtYqHEmjrUbdV4ECFKao
dKKk1DSBJ9plkFMwQ6UNSKb7yfznvy24sTJ4+ykRq38g/opecUuInXlZx0YKZ4Hb
s2vTY5J7zoFQLVtOaKAAz1f02PLOrjH/BHB+8KixV+3LcFJQEM52TIf9Kw6U5J93
0sY/Ad0AW5pCTTdofknZyf1rJOsXNCgPVISCs32ARZIwnUt5tciMaSYixPs6hC0J
31LU7g9ZSV9OW9Dh6kxGay26eFRkngJtERIjVEXL9OjSE0bPFT3rLM6516NMtVcb
zxtu+YzGIbhHVJkrPzkcuplsLtfL4xfnN+/rEtfhjQzngD4IYbekJs+xBhe0ZJyz
5M7LARl8nb4TqbzLiLpMEVEj4TPRKg/u4xOL0cQJlqgu9Y3oz5Lc2xDCAYujL6cr
7nuzsCsBYSrjfE+hg4HiIAhX1haJo4XFBwY7b6bCqyBs+SX2Pf6k0OllxHuH+5PD
KpZFO7w2BNVASbwdDF91Qkdd1C9aw+dVNsw7/QEj3rrbeQnd2kgzSB7XAyBDPRAK
Jw9OQU9kRNM+/s2/O4MOmMGFKE7I0PhFfyjyybxHAbwDUcI+M1f6IAsbeeZmWquE
pTnJe71fhPdn1zB49AVdeOJLM/ojOFj21NiHdR8zOT8kXU5BponRa9mLSFnVqe5W
cJaTX5fCdJx4KxpPt+uymi+GWWXtQgUE/6kP3bcZrnKYVAunT4PeogoRT4Z+IbXi
2k4VNcM+E7pOGV8b7ZIlG6p20k3kxf1pHLVBOtVsw9OZlIL6tJXWbMLedkCDqpVq
VkdPBScL8qvZ2dFP7WKGoAS+sjfe39/tjdcKR6fvU/C6wd1Fctgq9hy/qdqk77z9
h3N1hDfWFRjihYeWYYr7xPqlZpBgsVXOEcwKlsG9D6C5A0PlH2RXmSJw79Baq5RO
MNjCXKxNxz8lwX4OBO67G1FdKqb9dae+YaHo2tt6vhrDoIZXHfeMqgLC5mdbE04+
i0LfEKyce3ZjurO59pAAv1aybfd3d+zgViuen9jyr4i08L8OTT8APlch1xsHgBUW
A0gSuR1034XQc+FHoPxG+QDubHw/VcudWLnQkCm+u+mTxt3x/C9pVjPWrJc90WDt
OpZ4IpE0F8lVeUCIYymlflFcO6MDa7u1W/Er4ak2BbguE4myzXzLSWqUwZrstBsr
Bhwq9HO86P+QuAllrAkH6pKm6gNkQnjyjNbn8Srjcjgy+xNu9s5u+c+ZBNIAn76p
0HWhmCaELfOzM36hkMZq4W650pCvTEtWBVN1YEZx+a9AQy0/doK3VJ9VXEhhcl3G
7qh6trDJPQQi7K23kdZlsE4f22I7mEOkqJVXOPEJ1OwbzneylNw+uvjzMovS50Z5
heuWv3BGTUg4gl3iLM2SC57PbuE9eI8rpU22DnZe0lH+G2GFRDHTmCVARUAHsKdS
9A4doEpa5TMICSQa9ANwI+iNn+s0ISB2QOZpDPxFtv6ImDCrQuzEDN0WFG4hQa5h
09u/kpP6Ht4ua6hogfPysHwStyd23tVMe0t4NnRCjrDrEeR0wjs5tYuMP5HdRBvm
fYjlDMajn4UVytb+BMOpoOR7raQJj0U9YbB8uMNQ0+eHIpFd5Lw7pH3e6g450LNv
VfWhcHJd5hbn5L03ipE30W06jKRfBAydRoz9UFnQgsmERagLceeK3GBDLuaDo6bE
GDfy2rkSU4obtZAeSUmSn+5jLhYqrqRu8iTILeFGbTPcuqABDsqSyjfnA15pisbQ
okDdA6MUJm19VBd7Dw9rgcet5SOYVGq4d054j+9tRtNyjvD4zdMzF2oYGb4HE9un
N6GqtYC0XROAQB6sl9jBzkLnqk8LmYKMCU78DX+dACpIrkxiuvbxJQBSdVRzeRWw
pHhID/LdRaphAkGPk82FQMnc0X8KzjMXFPsq/ZP6fTJXZkvWeNZRcTSCfSIOEnWl
khvbMc0GbWsR8UCQrOH7lEeaPv2Hipj+HWo6OFgNScWpkf19Yw4tmtlhtUT39B4C
FvHX7EaQ4noHlqIoCH0JInnL/MPxD29eZGsKQ1of6CS5NNntgs4Xw+pTwmrx1IUq
Y3r22HXQqvj2mbzeT11ANyqv/8/e6g7hJtXT51riQs7sesYTQB2PN5z1lFaxGBlB
ZqSaEHqRRx4dT1i67HICg1ilgeU/Qf1ZF0/jSYEf6ufKZ1CKI2lQQAS2ith33lB4
VGHwVT8f2buTZ8KK65tAeMh3u1Lc0yOtxy9IEI/6rmyfsaq3UH4auTRUyqTuDhcG
8KoBaNvyrdhyNiZfE3xcFswGO79VQ55BRSlDr3qhzl3rGCFuXidOG0VdKqq7xfHC
v7iK/MZS8t9jpUvq8GULuuDa5ggO6Qpfrzpd6EpTvhCmF5cysInRxFsRJyfrnQge
F33/erhC2Z3IgjdpJgePU1rT4tzW+N13ApEwyWwldsWFb9q01zqdC4+EnBkHkZ2L
UQG+xWffqn1o+3DbvTbWtUf6BwQXAiDpY0kvqU4qGz9rN9Bx/cw4FW8HzoMvsOgm
ISocAyS0f4L2yAqUJY4kRbIoPZ5V5ROMIUB3bHq7UIC+V+naa2DVTwVj9gYLlpf1
i/HgMebOm9hCEZjq/9/SpoUEfMf4P5cx/QNABaAEUEP2gMT77fl95FwZ6ISQx3HQ
XB484tix2v5XIoRlQOFqMwgK/JJDdg+L7tKOQ47BsTFTU58F4gEPtipU1IRcNAKS
NL/c5OG0fgORS24gwmSHfCnyQCvl4zQbWiQKwDEtGXbiglUqnsdE6+ZzQ9xieNp4
PBPyTZD4Bvvx1qEnbHQLWrIg5cUdzhLeegY6Y9az5LpsMEj61WRzydG7oXylhhqj
9Qu3UjPfDPckhuj0NcJUtRpCADbw4TJDe1h/eoc3YI5icQSwpa/CCla5lrRO5cGt
w/xcBaiMVRpFQ4hkGfBlSy+M/daR52nikxUb9C+ZGvaMDVagRJBiXQ4puW7azkIV
utH2fq8KujRK1vSiVzlDm7EWaao6Bv2zWiM7hRhUWVjcijKsvCioZDo8H6BUMG7U
aeXVmxO2dZVoDet9LY6OKYRIdcw3O1oYOc+Jlt99u9E43gazEI219Qpu6Z3SV0Xd
BLUVU0o5lLgJCaP//J3K8Qd6A2DF0xnovH/dWgYrJ7VMAcQMmBctnO0G78U+JxfW
fdH/wWcVRlEgW8FENa3gJNyCotU3hUxa37IiN6qZZtTl46eGpZ8VNNL8E9BGo3nh
amGd86gpSbOeSQ70s7Ojg0kxPFu+EahLnF8ODJlSg6toVdATVHcbiNqpcIweIpb7
NuI48IvQcDTDR2x+IQv/sTxhlkzdDR09UxwIzCV1NvJ2H9uZeip7AUkCyW8OXq1n
zm4GNg4CeTH394DtAudVXlNXsUTjrnr5Gh4AEYpoYHxbV+JYU2LEkPcArgdMoCj/
gUGYdB4dhnOGawKgIJE94WQBpXp7W/Y3rMukUz0Fzx9EYoG8A4GG+Nh495XFKA0D
EDD3us6zCzCsLsfm/0yJQcUfCiXNlb7iwgTZqaBVrwdyyYrTbKJoZZoxQNYSFzKq
Fpm+Kd7VACetv/MztXgjz3v/ozKVahnlVqIU/0X/ddMiie5sDRSEkZGValumo9Fo
zm3UmjEdExVdVObeX6yeZfwHOk9T5UIlxfjUJ6un3g8HWWMZkC0EDVhB6ToECxPD
FnBpagqjv6loOyWQRo8x4VWXDBNwN3KqvUCK0xw+nlrKxKYTnzS0jrXK+Kz3CyXe
3mf41858I9206LIDgd7OlaQ5NIRM/sco2H+TEV/RPymq5K8eGHIXSvM7wubyCcim
Q5c0PtX2AliTF25MaXwoiwCjvX8McftAvtD9mwdmbIvsEvZaKVaVvZGXBHFX7y+W
Rg4rSQv/Ir9XKwGTW/29oJA5MY0K5YLq+43Wxt4/vbzuZcVltt/KVZ6eTrVJqk52
rGfELuzcaGK047rlAaQWoJT6uQ6vVDFFreFkKNH6p5CRggLirQl2t0MuE50cp0zr
nWxT86hNEc0cnAIuh79CeNDBwqkV8xQs2Krk2UGuFh08uPhspnB+Pr1FQh0gjIyW
zmongFrBrg+PQPA8/VPG1509Kh7Kke8Pffmueudh2OC7JL5OvnPWaHEN4G7CgZ4I
b8pETO1bKbWwo3DZ1aC5SR18e3NxSCBmHX7ow0nmyA17EyqKVroznlQf5LgNnyVC
wnPZY3n1d2XP32xkwmRQiSH+E0kAF6QTnL+XZgMEvm6cNMGbJH+2+pDST3OkdtZ/
BJK5p7P9ldNMc67pPQmq3b8NhCfxyF9dk1eZCPXH7HV5rphjk9WwHg+Rvwvfd+rQ
2+NPL2zsAii13TFWjNqdMhM2Wpu0TkSNuOiz15HiZdiqLhg8WGewUVdQD89lOzFQ
pZZWz/Pg6714FNphapyiQZ97lDjUlS4Ez/SrH5H9geHAovrvAZCRjPLJZys3J4zN
jDpdvV9WLBuwo/SzP57+EGX/uyhaVP6Zf5bJV537qUyGMRgK/h4PbqDX0IR6eXOD
yCDy3ui0X2xJ7MbmDkG9lEojQlmwVSi6Qhly8rBcGRMWCRfj7J3ua69a7x+oCIoW
10Au375jw95deT/6c0Cr1eaA+N7AIQ2J92BsJ/hpqMocYXw4ZGT2PGVZSciTkKk0
swpT06i/AWjlia7MHkOg8PzEcIv1P6EgAiHDnMGPMOrtWpathtG5364y4bAjT2fy
WwBH9remtXl4XupdnsC9kFWpjSLAwCErAs++KkZKnTU+rC79+f8HTKlFgkHi4QaV
/N08dR4qz8qmKAAvk9r3Vn5WrwhURKoZheKfsM/N6F2DRCv8DAwtOxI0oseHPgeI
Ik0H9i8lcI2Zc/SaQjsQPORmxYlHJj0NnQ57qvPyXkMRBtLBqzVAnIb50izMQzfg
d6bYmxbTNpY/ymxwPKq1kh54+m7c8loeySP4QjMybHrIO/sx/0JmirV6Vq8v5Adv
xbiFMo0CiA7lDTvqksq3SAmEAnxiFM/XTGpfWFK92foU3lRB+hAH2jiQrX0Zp3gZ
oRZ09zAkfD1qfM9xMesKVxD7TOF0h1DUk93ca4aeRweItdd4giNe4XRLTUnnFm7R
V9roXtj6pBJ1IMnw9ApCVfFnXG8DhHAK7HVwfw6ISGHS3dPqhFAWLVdZQshBP86b
mDqlXJvU6fyGfLb1018V5h9BAf9e4ut+HHfF1hmsCQWH+s5CHsoDpNFDnDkPuo5S
PVjOhnQBAgBPIVM/9yCWxg6Qtt4F/NXXJ2o+pwgnUHkNFC2J6QMuTQQsLo1iCtHG
wpBsiHMt7iKPwq0BnjPUnDsR/jcOJ+t2dLdIPqOLqLnVZLNKbEDyLwGWHAmWoPuV
tkItyKv8V2tK/QuwyN9aWdKb/RGjzNpQO9Hec45nF8BAIKwkR9MeAHyZUrIbjcVL
hTQh1+vVcp5DI6kPbNTwZ3z4cB6rEUUbqDQfS+uDKF70TqxM8gkMpEY3V3Q7UNeI
qEwnc4RVsYsh6rnqMswRAPDBYCUVuxqALiR8Uc7pv/iuPRzsaG+npxPLN9MsoieK
RLO9tEufKFO8g7qxOI+ms7Ro1X7+R6oquXtwhd1fReUm/L50cTmiubbtCt4hRlne
IePtluCywT9GQ76w7L559GQAuYW328ylnvVYRBA5RMiPflQ4B/j71wuNrBoRIn4H
yiils5svngxB7viDBOJYdS14bxcJmF+LSYyNyKqFEBhwb/sDCmMSXNxbLF7f4U2w
55zMKiNkSWyh7nvk1DnVOScAH8r0FhTXaqvGZ+Avs9YrbNS99CwlOzbirVTZdThc
jtOY7JWevXvMyPtvenQx87wVbE+Aw59yRRAr73i7JWt0xrBfirA3IdJTBvm/KYJx
jxY/OmjwZa+Bd6JJRtLZvZTG++AJe/LAfhlfHA5QiGQzOHEroZ84bkyAxY4+RdFc
oACiIWdjQqYKvElzfIBz0Oh7TQ0C7D4Hp1oZPa7wRC3Dc5Jf9DMQ5dZVPvAlQUVl
py3S0Uhz6nWpaMcJTmS8y71MlDUMjhNUWesL3cy66XjTTWXhfIqhAcna1Dwbln25
IZauPTX60tsVZCO3XfoeqVmOrwEw39nNRh5sygmV87IJySENmLHRL5dS/ddUDBIz
MzLRJFYihtKABgPr+x5mFSVsVqkb35TrVpxjt59NqjDp5r0iFGTMzvWYHUArpq/T
vJ6B+1XMaML4NchPMZmSWkgJSzTgCktrtJzW4Y0CgF2FWu6+qlSf+HA7XsbYlhbG
8sYI18BycS6ODGZqIKJ6jvFiq9TPeD4OCBaDUmrYFJwTFIIg7ARRGQQnni/7yY+K
DteTsQ5KO+whUSIVFl0QnOrt46b8DsBI+Kg5QNzCjxCyjdf5E2eS81YNlzJulYGb
/fE13ERkL3awEn0hFwaJhWUYq5XIysk4mTgbyg1QvnpX7UnfLNjvKL5P0LhQnT7F
t0dntflH6/b5vFAVeBZJ9Zae/xVtI2ZhV5q5Ep3zugnerk4Vvl1jqWpT4A9U31Dl
l33Ynmf2SFJCsk3Uld5QmgTWnWbvUACGaphf6/5iAikFLhwpG0RSh9hLIIbM5GNv
FY64lyMGdrjGh2TW8EqSepditKjCdhOdnwCsevCgc5U64CqDFE3rUsTjExlLoSNW
xJ5sHevAXc8wpkYnvwNhQa7jGIZyYRM6N9uWwFo/krYjI+qzGOOY4mG1Z4ODaxeO
DrakRNIGLDW5NFCnjqkQl8S17RET/W5hy1QJ5Dbj4uL1rc/NSuzMDR3E9iRxkGrW
qMnrbtkLUW9EaNNVKf5Gz2fASpSJwSfnxjW59omOKa/tDl8jTMN0zetsXrP9/t8S
NoVAiuGPTIpxUItyhOZty/CF/DLy2sTAkFZ7rQ5ntimXQimDiUjG1knZZe9vYHFG
U4RBCm1ClUSsPxVxeL0GI16i6r1X0Dac40OLTuiL0K3ZUBbo/fuanu0cSsGYdhWD
Dh9aPbbmouSwGzk3j3JP2IBmNEVXqWf+H2SS0WI0taBv5I6Y3Fzr3cdbhPpVs2k0
behfZHT3d4uRE2H7n5qX/xZdp1veIiOPPL6DN35WP2x+ok+cxGTLYSqyBvUQygHp
OTvJs8ezmNY9hT7P5AwWzei2irCt/exywRKcWaQIOfklnINCmqHJJAHQo+RpZlJZ
QSufjIc33mx4LSFpPOF9Bem3Mnft0ckXwL7qEuHdwmemPqjgvyzTnfjmjkv0WfN3
tJynCG0ZnIHTNP98LwFrUJd91+d3ZrRWofsHm/qTajYBCNKwqxpFRXo9c2APqniw
gSOxaSoUZ4yJVE9h55cBNs1f7RnCZmasqLTyDcIt1GigEVDYRnOlXMlDv9yneTjg
Nktirq65hjMBdVaoKb1SzlezVnUYEjjkhza4S4n41aIJWMTcn6Qxm3b+8EOsySwO
pJpWl03GMsxqx48ZI7p7hwGKQ+8rsdGqbYo+Mfelrfcqc2OsgWrirDCH1JUVjwRC
3VZquaUIhg5vLBLkutvLnIRIsuY6cuXaRg4HJEDgnyiEE5q4/GDYKK9WbFxxQnW0
4cMWm1xtGFwjpV2fE5jSaLlnTzRlfkKB7zl3KTjLSMAhTSHhVFpLXL/30rxIPO23
0B3mH5IY0DORv2+/TrQD2qnwsDWvWDxvjpPZaF3JKYGmLXMIJ2rwpuxDETlCB7TF
xLsI1M5TA82+ZeIL8cAzdsxulfc8IQ2buBpKCnblxwHHViuMF9OVTNKO11r+R8yu
fg1ps4Sp6S117AWWZUviAQMLDoeT0gF0QgHbHUW8ZjRu/RTEqfaZnACUH4lpjNTQ
EcgL6kPTR0ZgPyzXOMbPlsutOt5JGPptx/yt9gPbZ0557NJHIly3jF7s0LYpi3b+
3BZQD3/EF+uN/k3dSFlZxvi/nnOJjIRzXrpNZPURYqYPGoIuyErzNrPuCO5PyQwE
5ZaIWb0QjkBnxzsVVu8KGoF6eDix5m9Q6ArOO0Kk0Yzqqmm1fDR+Nlfjk6/cGcNg
UXGRoWl6kR4D6PoH+ZiU+9sqSOZV88T9q8JmHKiCawV4LYa5tk2Ob/jhiZuh6dJm
oyE+lREmpE97we5q8RmVw8FPBz+kM9jeT1xrfqBY33ihNfgz6uo6YokGmpaJ5Jbt
OYYeQVsCNXQ7NxxSGeKjGF1IOA6e40651s2NTVcFCOyCf+lcoQaNutKxa5iDfMCr
DNw/O8gr1PKsiKyfQ1yRnWQysLsMz5W0dCqtbg1tsPyi/iCIA45uWULmsE50AACw
74dnD9JHEJMHfsW1s1Gd/oCTDAFSM4ecAf/RTMiMsXzGIs6t0jpvP/n/MsSXh49U
2c1B/y7gZmjzgonctzv4CtD3mPQ1i/wV3ZT+s02XNCjkZodCfpoktrhf38gg6VMr
RzmKeH7NkJCOTe3me5RXsbt+S9pKSW+xpDfoUb+a6B1tj8HevnS92VJ+DLZQ8sXU
VcWKi3GAtYINlTvP76imhjn5XPZdUfWeyPi+O/z5SBWiQ/lY48zq/yNuVS4ZCve/
2Q3bLGpvFMjJvKt8HM0LBewHrrNORAuDIYH+zo1xVdR1vCWkVKmMOcKB1yRu2Jfn
vI/cqwEqWi6/AsimBx29d1CoXSlmbO4EGRrcpzATn9xdW/JIEP69++w9dfTgfXE6
ze264A1WDh2FoSd7AahMLl41pa+bUvPF02Nk6nifKup4LFq+Qv09mX0xoGBbHyXF
VPfaH4jy+q7P+tzpcAlFK3HfrbV1MzqLvsx8M7WmriUlyRZ805hBvMG1v7wqsde7
uvel77Vk3AL0ewr4LYKvd9CA6xxEZ5oiOUSRpvVS1/ysDNTQ7Nt+YKkc8pUcCNRB
DQgkRDq90g1cN2miB2VYIv79X6bjV6v/fmXg2B5bdr/fIetLkDFGofr0wvHnb5fP
Ib/nPiZUDswqhHu73yUYUNEkS8wI7YwtdZeYb5kaiOWWLzh3L3853v1zi7Y6sYWo
PdhfaoTaAm2QPrc8x4ij1dpB6hXlr4J/gzeZRCGcsGdCfXs9lSnRh/xJ4tGo8Hz3
PBqPl9Wtfxk7OJS9KZ5P+gSaxUe4vwZy3+tD5wfjp0mpTEgxQ9LvVfLA9JANK5sK
3Hh0/lL+Wtv0YtopzrriaMR83wtVhesPVdZRED8uXSaWmf0ffQnejjTE9ZHEOcjP
B0NdUK6c9k2CXgeiF6VJvyslb852KwRf3kripv9KzapLLE5TApjNBKROU0KY6c5n
oTN/iYqo5eD3T5CWqQHB0Yog4f35iWXm1lUkiV3qPDQVOhGe627u+g4KO/Gm/vHR
ltRVdtBvt8IyxERVyB5cnLK0FHYFFoSW92bFN1+XMud7TypgTw7eQ0+AenzL8EPP
z3yEaFB7pF6xS3+SwoA+Ya1OPDSjeIHilfC6Nnq4zibclhxHVjNjm7qOODyE3Q1a
0vnBClbie5Y1Lgw6IbVQUSzIsIzi687rTfHUcKKvgwX4aPHgvlTMYrMZnElJk1JU
9hm5QOMfun93shrCBNu5NnukuvaRcltbdx+MzuFRFfE6lHZ4r4g2t49vlGQjamb3
25+MjI/Qh/DbhBt7YSYoUigzrHoIyGCdIf9GJ/P1WmRWJBfZ2eKsuUqFhAnifZmM
gSGrrh5w7UDt0ICedTH/3Ftuy/gJ4lEsYBusTObX89o+NUGwtVvsIVjOOpsku+p2
GkC5NUrnqT99sTlWmhlE7y2jvGIq8gT6WnZ6eJZ93/ygvKfbUcjst2O2fn9Fmb6L
iS3jrwN0rlHcUqy6mh4txKHrEetnYTcpNq/TADXB4JecmrEXDtjVUH7MoCpeN+i7
i9W6OdeY+ySo6LWorncjVTiqhf88vevCkWlqezBrzuZ3QsYVtfes2U03Im4VSq9v
+Rc+VmmRd0C0hXBaOIB2eB6YnBI0vhcQul8c2QcVgw3nJbUivy+AZNI1jjOQCk6E
2ISvayLL6MFxs6ry9z+JtRYZaCEdLNZF/fyCYrDnnuhju2l4np7rjSVaiypK9/lt
YKk5JBjy9nGs6Ny6ml9g887thvrkW3rIFB48RLyRdzs2UYyuYZiQ1j4xqDfXvuql
si61elQUYcTJoKrrtyy5MXpi1yeSrs0qOabCSg3PhWZuvWg16liL7Nm1PGN65lun
uoK3DuV5WxGOGHON7JNuuzcSv15XvSD2UsqM7VSz7fps+6oPfObuOL/F6EWC4MUv
JGd7c7azVSeGfhY6Svxz6psm5Tf08T/8vVnTE0goc/X0NpIYxoj1rC8f33WnHpe7
wUUoLvA0b30vKYl+KFKZOvT3EK/tfCQjWrU54eYo/esfUTTz+zEqm4hl1Ww/Sq4u
0n90PQDV4y4fPEuCI9zeacQ9477Azzbhqa4rKG+DQUpUr22D68IpQx2aSXOHC8gE
++K/t+PcjynhYrB7BnF0lUCATtMxGSCg/aUzJirUOa2wqwv9DWf38b/Sb6xfNTlP
zAiCW+KCcR0J10/WHkfv1Vwgz6vA7zbBu74xdeQ1cwqYXyBKt8zgrfYDOpW0n+/p
ILiCEeyjBEvwhRzAEnhuDkuhHKR2Q3ek4NS4AN/v6ilvBI+iQwkcwoBZgcovscIB
MDPd6Z4SIsLNoMd5UzyzTy0MdE2sdYkCtTviCfOj9G3byVFEodpSCg4I4AIp4HC5
B6dwBQPF3hF/rfF5JrYgjvCdbIxSVF10Rg/iOxvboPaCYY5aeDrhxcdupxvrWjVy
y1qfzP3nfRfItpazlsdW8WGmtdC47uk6kO7J6apswjipMPPG8eVpsz8AbA2fT2ci
ThoDL7ZWCz0SZ17kVEtrVByneFfQf9BOEjrT0SxcuuGizBGAsTzwpngNzNoWm7eT
PcT285KVaMXaJ1ULApA17w+Qo0F7yi8NHlVESt4Ix62GxxhEGXDJvGe8kMo4IExR
+ycBOiT03HHw/OymkhVwUu11y4S/m2F559ut5Wmp9TqJBuLSbF3r4U15Jd5Ks4Pi
3ohMfaF8s7rlj0S3XD0qNWeygMEVNeV0FLkD+Qv7gdo6zwKK0hBqYewyYsrMdRcV
iMmgApOJfasFqpOWLl/6m7adJt5LVCeZSA3C6b9+GU0ne7ES02bE4kjavc1CH/ua
ZH2UNZdGr+z9vKz5GrwlsxtZ8BqoOhXzqXmzK5rBtjdBN64XKndo+3PBP+RPaGKC
GlAHz4TJSrZgOrfYjOm1MNLBwG2YpaQaGikysC6HgItnRv7R+jmj+pqMCYAJ4xlU
cJeqOPP8fzlDqXSC6SHm9H85sLtbV2gX49o031U5XjAHilGkaHIf+Ggj1aXCS7hW
eatN5P/z3Q6v6cH1nKOR/lHX7SbtS6Bwl1g5EN63MtUuPkQOPWkRwshoJtUTgenL
P1cevVWcQevE/xhb0jfc+HEGVY/n3PuwFlil0wRGwKff4CCKFPYmHovQ2Ajw6//y
yP47o3SLd0a4rpj4cmLKcQVfxJTdH8SvL2aykLJimjc0qDSnqj8M7CDJMXllQn64
IZdG8otLv1HTQBOgKwCnPeM67w7RZoNoun3qeA3lDbQhnTUJ0kRnzKyhSwhNwUwh
HX4fqNtY3wcs3fmtSwSTsWh3D+3QBhGUQYb3fjuLP+AiiUzf/nfzzE2R2eKg6EjH
vREpucOE9L18NQ+hnideQMzc49WgMvPdBkIuP6Yobrw=
`protect END_PROTECTED
