`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
enM5PF70c+Rhc7SnrQymXRU60scBTmdXuKOy0fObGYzwDoR77uNOR+rmoqZdQmqp
1jEOw2mwGp76jBftoufUnuxivS5FK7xDOfpzVQ17iaKux618aNnXPD87Dci1gUow
kr1n1GBAhbg00NqaWhIoPGV8+pt/+47t2m0jaCcpDO8aOm7twiLy7qjm/2BAZ7Am
kUFbL4lp1B2Zos3O3iiMrdaBOE7alftUirpWFPGF16fxuCiJts1L9I5rqzavNilL
dxzXsQ5ch5mQ1zOqS1NttvI5EtePMV21InBefws6OsLAfiI779gXKkJ1sQgzjvsv
wvSMHB5q0S3SVuX28pqZ1I7J1Q8hemrGTbKP1Oqc3ts/7aJ3Tw5RDu1nhVCAACZ4
9Amx2Jqk+CidInY5pnPyYd+Utz9hBhUzfQ6fGL7Svyy20/Z+F5wjbvOtF7IWnWYE
Zsb7xF6SgDNGq8ty9bBsxF1zYv+EHTsJ0iB7eVjMWFlwlI8hWLH34rWf5hnnYs2r
rg4cCFFIDl3prU1X7a2uMExP22W4PhsW6/DYGa32z71sz8lcj28pdvxgWmL6Q7To
MBuMeB3+BjZ8rGidNzK/SNTYvUBsYw1Wgjf/S9aBXL27J2QwKQqsiEsrFgvwqSsc
1Hs5rawAn5BoxO4JtI5Kbi544LZdcG61lbdPuESKQkwvTOi8dyVuS59sl25Yyud8
ypAvHU/ym63+aWDA4wZPyQKRnfF5n8ueThZw07fA+FSCsjfScGiEQEY6kys/bOko
IT/8bCRhYubiD4Qxk1tWU2zrPKzWFtRg13+SvzdsDYWTRL+AlJVPIE50y9A4mXkl
+wUUaA5P8eERXsD5j4ZWcK+TJMtuOoY+I4rJd3dDhuXXc4BexccaYsbQn/nW7m6l
Nun7S38ZRBZs4CSgHFECdTZISYOKTCac/XFNhaIXbJV25EXAJhwHQ0ikqmBoKxi+
Cc55Z5wwcxy9nBpQrqHzybyNgX/TNV/T0ggE4OgXmvdBjj/3T/OzaYWtGrErb29V
d9e5Z3x1NxuRc6KfFW6cwMKpWXYPFQettTJFnE/r+Ab4GCtX7Lyx6C0jTjiv51gL
XQ3FXl0gM5Ysl7/zBN0TBfa+PVR4+ThA3djFHJxKqKCedgBglTtyBBNnxKQvUw80
G+PuyefDMfkyIUQsTqi4l03agSCYL+vRzwHxHDHbDimTBHvV8oJWNWffCDFdfHhK
xTnHhTt+COrp3fZBPMw0rCumGJiy8ax+MCOdJEQXc9CNB/EfoGD3K+CS8A2X/PrY
7avh8UmTjdgV1bnIMJHncPL5lzxYn3Tak+ae9TJrgo8PmBUQBtJoqQoEjzwEErgl
dAg8G5b9tkj1wJ3DYiKZLiD8oOZtWOSHGbFzA7b0MHlvtHs5OHUGXKkbGN9FBSKB
gbDHOcWmn018ZT2161kIhYDcmIYNf6gz6tFEUrd8FhlH15fomlwQN1vdIvxc0eBO
fJX7YMxVJVlDbQqj9cT2w7MjoNcqcYVtInBMrfrIKBr8zztb4s8crMNJwci4S3co
bOdgz+DxVswmYyPk/yqElb8tMTclYfuW1b3YHBIpvI0IO2nIyCbl7HS4rzyQkXjk
YcI4dM6ufHiMEg2De4UYSmeAiM2qFqUs5Rzj4Iq1gtE=
`protect END_PROTECTED
