`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n92IAXGTsKoQ0tzhiIYzPOpYJi/wf5X/n58jwjsO9m0OVlwPy9lKK9kbJqYryoe5
r6b5DOG0GuPboAafK27DhXon0pqHcOVpeLVsxUc5UpchVsILrYq58T3cYBgNHk5E
/b70/RHDKA/yQURrROFQ0XA4hdp/2l7QbDcDjpcd2U8=
`protect END_PROTECTED
