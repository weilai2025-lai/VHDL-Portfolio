`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oUcgi3w2Ss7Tmi5HSqOyyNB3WsyThMa2q9RXmYn8LMzDn1b5LVx9UVaVfjZJhJDA
EBDoR4bwxQzyfpMLgyvVnEA648RF0gJsC3yes1FvClpwaIOG2amp2X8KREfXJED3
Xi8ncKRs27gB98Tuk5cWzV/lsz1hzsYukZ5mE7WyIA+8buuQRMywbCM8aeUfyTg0
OuoNGkoVp8lMWFEU7BQEkAYoxNF9wWwkjWoQkHrXN221i+Yn8OnFi9hJvIBGVXrQ
BgomHO6wHioP6hONmm/bP14bz/73h/JbF0AQehbuVQWprCibkXv70ouRmoYpx+B/
p/rUaHXPlo+1AXSjBoTMwg6olFlv9o37EZOoe5HdoVWEeSA6D4MHLkp9TanekQe/
xDxBTL+Ef1n+wP6a37347rs03g4WVJmqOt4p1/Vw12LyFWRB0lvcTpPae0mblmpW
gp+ON74BsTiEJUcKz4Fzi8r5cfNZEQMPa5Coh4tw8192AVO733pRaln06G0dbB4P
1lFDpjNSymPgOeIYZ2Df3qcDmxeBECUAeMU7u9H9RLkIE/wFzkUsV5kbNgo0rGOd
mB/jOtiRSLVpQjGH/fx94ftammaRru4asFbIFCy9nBXFFhQH7xLkipLjmL7igCuj
YqRis0D/eBCju9SXVXscxnjqSzsD3ncCZIz2Eqg4v+QP9zR6VJRlrTiQSyrBbvLZ
1S01dFOl/H7yyw7xi44WQHeQ41SiKHwmIj/1lSUALiPTiibDA1WoZajQbI0Xr2Ek
YlJ7f6KSVgV535zYf3ttszZppMZ2WlWeA8tXd/DYKZFfud/TWDbNmqVgff1hM9Uj
D6+28j1vhxEiJovx90z/2RiBoa4eXAAydhi2oALvqZNxM2bsFdZcp0tDIWSq7Mtd
4liabrDKIeHeyiLn4ZshzawJr/cobqgVGTzv95OYYhEnB+FH4BN9JWIK1KDeIM2k
ymCeCRQTen665EGCWDNpD1lEWiO9FfLXRnGtiO4fP016JB3aUtDaPH20m6eSCl5D
sArj0AH+aaeAYUaJqHzC2SLBjhSwkLLjWyXV267ZkHgwJcNuwYULZp754f8g46ac
JJRcGGEcsToBzDGq4jm07JUVwGiL89PV5fQuPWyX/MojNw8y91lHFbFQcD8DbcOd
YuqJN75ymSiFNbaKcnhm6tjQ+fE9uini6xRSDdSRzFKyhx3LeHvKi3dufjfvBhHX
1xPosWT9Vtc/y2GjpiQtj1CKSYTPkOG4StOvK7UKgFiNXGEUTQUmclSz1doAfD3m
1V1TpOnqxcKv1CaXY1dE1eEidwoevQlh/sFL0R1zUex7mnhn1vSjK04J6+GOJcUA
53f/9zqVRyIbDFmzUM3w/fDSYTzoFY4ir2mpmbBhqnCoEY4wgXuZZGs91NAMFI9D
WXc8QstQH37QqXu+h52gEqrHKP4iLFCotUq1j0aPn9IOHDp58iD4p5sp1fpKUWUE
1SYHyu6z0Lb9mBZGWL4JB+nrAIfr+z//Ite/jN6Ly2pklleRg6EfqrErxbuxcGlo
APcBkl0/jWeHYKD6ADDOlhYKibzFkvhChTfk6EQoFQId66qin0Oh1HCGAGv1mAVq
HmMwIZ2x4OfyqDZJpfivnQkC43utzrQQmJUBpJIvl8+6Wpatl736MYuZR13nWo/W
p9UetHXU3/eGcqy/PBQSYbvdL7hWDx4enxg88SJlqoJ18lcLkHmaZHzQs0bhg5iK
Se2/8EVN/TdSoSFeATo5nVUF9VAR1ebJF7CSeInpn7Ckkf49rKA46vYm69Kv3rYI
W8YCrwKJo/zHQ4sFEGowWbahrRhqaLl1N32ZwXOTtX3Sd755eI9lihP5pMvt/hR0
EF9t+FY0GOiDvdCFk4zGSH5gqblwzDW1wpU5dpVvfZ+m2W7aNsNuyfKuBfvNi8OL
TnWGB4I5vr//KYdztQm4pgog3ZZLsOOYr67Idb2nPOUZySwhI6Q9HkCIpPNXdVIl
4zSoxP3xmuoBFdiI1DXb6X3hZdg5sL7v9wfZbVDvlW/3W2fC0raNA+RVJtgM40v/
IkMbwyVy5i3/aO6GyvyJ7CkOQuUHdvNMDxgQmwENJ0+je8GCoRBt0CtUOCmaiJZM
qKAJhN39+b7wO3IOO2oNR4CUtatgF+oou+ZSC++MxN7Y7aKv/Mj8ykWVrH8tRXou
rhYVS1mcwdFX/vNRJ7CFuhbUh6KN+bscQdrrKVrH/uXL0+tu0AmIh/hrQ3S9dcKX
5u4cfkvz0C5Z3eFxRAFAUBuXZbrqIH1R27l7jhALSb6MorqbR0UwyIv0xO5KkEJt
53xB9+QegNJm2mb49tBGNk+CNsE+mykYWxAP7EXNci9UqgXEfHJtFK3d31p89ja/
tuGaV72FEkqejIkWE4+6oCWKASB2TE1SZnyTKr/yWtfv8zO7iETw3NmR0mSUmOZg
kJDagmxSesZc6P8Bl7VYUqN/E2PuHPydBHRMmhB9opBVc+vLqFCMU9MaVifxJbMp
WTR5enK4Ghl/G+Qn/munw7Ngx1isJrkk8Y/h01/9Mc93jU47PMQCMiJf/a2Oyx9m
iW97AmzRui68Nh2YmfPCYosgWeSDNRUuxZuWd2zWUKeMIv1J6Y3CI+nJWvdck55f
98I9B3egBy+jjXvEMHkclw==
`protect END_PROTECTED
