`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdKfvZP8E6huZdivcmv3E5AA1isaP24oRvHdd8NKazn1Yk0boqhiLdLhBBvYJ0JR
ygt25zio0W1x60UwVD8YKqBeDPMDSMv/z+hmOtSGDTnN5Bi2PozgeKpMmdBxC19m
lucBEZNFYqYURP9Q15pQg5kYzGspI1TN3/IQcTC7GGV0gkBQ/bSXSUs/pGtM0TCH
jOS0HoM0hW3kWMpt16Y1Xm4g0b3Qk4YxCxSB/5076jeVA4cqg223J7ZcOiXopEio
7qCtdQ8N0KC7O+GY4NmqU6/8iUK3XoG1zghmcEBaP9YCzhmFyn1gvb22piMs8sNy
ezH49tvIwZhDLcQWqx+cCZ5dj6ief3dCd5VkTrX79oXoV0b2bC7Cmkm43P4DmAS4
9+j9ewy/O2v3KrvE0xnMrOVmATrHz88rbZPuSSVx9PUEtyE5Znh3piYP0/qg1aJM
k4pneKph6M9OeL3K1sp79/iuE/OJ3rso5AlMwE+rGmwYB0ipGDU3bM5nnjZJtE6K
0wODx9V6mpx9ZjXDI5NLqusqKtPwB4kUxiDAMyKzQcjey9E+1bn8+o3gV7m2LHyO
9niV9XNkQnnVlV/WgcqRnZTNP4YpIfZ2mWoLdQzMH3NXmYQEqnEiT+vRtGF5ZOYx
WrZXD3UOasHnZeMqZouNJPch7sBmYo2EjFucBff1G8/VxCO8GB9/YjbpSvDVOFKI
4hV/KJiGVWZzEgjxfYmOLc/KS49eFhIJcHaTqEXh2uCjrByaV0ketQ/19KiTebtF
CCcjaHrGKAto09KJII5c59KB3EHKE2f0ldqssIYLCQ1NSnIOWZVSJ0JTwFl7wfCf
5IupVBdDgvfWs+BcrvlEUionmA+vIxogV9r2gyVQhFY3jCfpai/Yv05+2LVZVkkG
`protect END_PROTECTED
