`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtjG6nvvMlgHB7GCZ6XcTIa0n8NuD3m7JG/hVdQYDXOyPQfYHHMkK7tSNO9dZhSs
VSn4nr/MxGJJJKKqchCVUME7RortsEAifbl9dY6PP+r2OEEmOpEEBE/UEM2Z8KH2
nAHC3VXyJcLW+S8XoYmw8kpGaN9ds5GfzaaLQuIdF31uQKmtUYXZxanXGv6DBKpK
JDGlLxaWOQvxWa+v9cBPfkVforSBehBBBhj572pKfGf0mIco6rghpkbpoV0wbLg1
YfEB3mEia5aHAEl/yd/msSlv3HV1jFifVboVVoxZ5iLA58ZtWiep6Xa5nILTRSB3
PNBQ46zdYVmLCmXiRk7tQbvpqeJpGAfI4SMQ/v5dii04R8iChOJFJEahUImfCACQ
HFees7N5cI9QPIhh4sd0vfoAkod8DmZQzKxT+AWXZSDE3qrFe+YHfP7tOlHly+H9
At67ba3kH0M5cEb0eCvv2pnSotVSScSmdaSzJFR4VQzWK1kfDnwryrueo2LI/7DH
sWyJ6LtQAuvRWkFw7P0DHVWsV+m1dkfCS6VjBfqgrhiCekN5hBLJwiohE+pRshb9
lhAiWQGQ6gYe8jdjsRhN2IVjDafhknvTzBM1QUx1CfUhUgL94LKP3S+eCFVpY8aa
tO6zUmHULLdBbVwkpRF0OiC8yr7od546xX/f1mPYeu0pGvxj/+UvhMTNM3TcyjWB
SsulHPuC1ZMK2euVAVN/hkwIbBO0F+9vyA7osZGPqOivVNPG16/eYyoKP3nupV8v
0KSlW6ZKi3y+NmTorpb5d5MjssYBCFrojV8L8QRNKtEk87/EEJgCG0IZsGua/A9A
vOhRzx241rjpYOs16Y3aomUWmaLB0ew9Et1HOitLY23SBpLHro6JHe2Ns7PKdAcc
1pglT4H5wLl52/e4DrHLtuBzmmqV/mZ+ms3HqoLgUKidm4smsost2m2SEkH94K6H
1MZq+x4hzj5UoTXuhCJ3TJ2uKzahz7GVk4QMvfeJCm7FCFuLPltQ4bdcUGvDxYbH
qNcL7WchDZtACTPhrHlbo9b0wdjS873eqIkJ4R6ZmzmInCbr6qqAcljhpYr5lola
tTgMo3bpEf0moQr6McRRAhi8KssENSLrcry4bh50DZdPK2iWwJ3qC1kZNQOJf0Ug
oi0GhJX1jsNISjCGksFzXio6duv/h2rNJeN7bcQVV20qRhiAJF+iQ8+/cTq6Q/A3
1FHS6NJjHgXfiHI2YWax2QbKYqN+DslCdCEc07x9n8fhn+N9cZ5YRu/Jtg+7Yjmc
riuYH5AIg6tzRBjJhRimaic5kV5Q+HTFWwtrGsuMdZ43rShvA4cGEk9No0BQmjzK
RgVhq145TjZ9miFAzLp7JQM1t3Y0y90CKDz2Imuf8Gjiil7kE0UZYDFUflN0C/FI
1hKU7UJ+zpwtb0LUjNKNsULdI911VTkTn1ND6ese5apKkRu4h6rqk2EdghM/eAVX
az+Z3SyOuBPsRqCkCNgS9Zs/cDTuqFMfYmtH/Kig1dszeF11DxdhxzdLw0qrjYlo
Jb2OtYfWj2FUDzeuiwoF10T9PVHs22MkssgWQ84d3StMeCpxhJYqiLoGl0xK++GY
28lr3s9MOvC7+Fr+t5nxac5pcoMon0o9ajwVUQhtVWwRjEwRP+mbKRWvCzpJ6ro8
gxGROCyy2xcd/Z7lwurhBDlRebcBOzxAxUXWgDpOYx8Jw4X6F/OdUUS70PwBOwtZ
MCF9S2DqxFoQ+Y/5ROKT4qoQz8mA/dAU9yKsdbYjbELTPns2jvt/jX3mFzFCpaUQ
mLBcL7mL/NrC8RYvVw5T8zdK4G+zaDf2Y0pHkmmWoY4neSMBYZG+PtVrL5p7yqWs
iFSrBKD3TrkAyY/f1EFDa03xzG2cTczLzu/DSCn/UZAqkV1qD/+xafAroS2EhiKH
Ww+7YyGUzCzxPDKUZzD5UoZFNJCp5r1kvG786L9RFHW30bd1E9/lPLyl65svaUQR
UaxW5n0MuXMzDIIdZs0T0U5ZE85pKfmaz8sypszu4i/Mg66DcFf1f8E1bmDWY82g
cZLF0V5lisStwi9cuWkV5mv25ar7AQadkviX5glk1vOAfy3ZHJREJ3F/iCkp2oOd
MPTAEwXLge6ijv+0hm3XbqGIAHRh/gGbbIL/Y5XnVANpshay+4oMJzhRhVBRraD7
LM6mM4Tyqqyi7Vt+wsR9H1KD7H/homAxFTJ3CKjuRFGJ8aenXTC0DL4zq7l4vsdQ
Tv/cPC2po5vyaAcgPkIF/K+TABZrOjUImBlIWexrBbaM3JAws67X4bKEBUVG5MXc
LlQ7tTl80xvjK+5mg4Tko6zaO3kHwfbrEKyag0RKrYFgIG9ir/Lx+lsS9ZCg3r1O
oyiwLG/5hnRk/817WGWt6cCC9ya6Sy7LRxnqeqJRuPhU3cpmNIMDEtYCDLxF6tNY
BJcY1c37ZvgZTC+13iQaarxF3FmJUImDltxQdb7yNC8MT2jJT6E3jiWcyr7iXsvk
Ll03fQYnR5oWSHF3kz+DXOU0vUP2msW68liGtMnTBcgk8tqqPOZDOhJYFyvlNPUP
vNeBKnSyK0H7HvAqXKPCke22tAQ3avVId00sJEwsevwPMh0oXxO1iblPAnEaUttQ
BcQamI1U40Lzh8FiSWF5MDmWGBxqR3HjPhyq4XbqDmdiy744Ku766YnCe4FOMcNv
nMpZlo8Vs/7cx4/wlR4nmT0UwBtB0Tosgbx00QGTponfaIrZEtxX8sAelOKTlMb5
F9u9zMH+L4aMjwwGzf3nEvMm+42X/gDULreWlZxbkbp+tNvFji2HWmQzmH2sDu6c
qPPzQ89AOFHAVqXfP5Pj8RsNEFXyysZZ1mLXMzb5GcUPH093XfZ8EbgOrAhFUQZg
VPOL4nvkfJ2N6LScbTwCPUxCJzHYYwx1lFV2OeI5UOfc5bbtIAhVJu3/itfYOQBs
BXprBToDK5n/TfM9r4hGUvErhC8qvs5lzmcZtEtAlDO2Nsvh6wn7+GhrkAPrdavI
cK0/vP3WZ4D44xPe1rMBWT5/kUqB6w8qqeWsfB4r4VQ/s8DDfqLnu/xxsYYKLx4q
mL/QrXA7YqYu2D5WuEzxHWFjMWNxSzO6Bt647j5t7hMZbipH7G8V9f/kTUmm5v7c
ZTCtToALYs/4W7ejF5dFeY+Xpb7Fi2FcTorSmdy0EapDADzfgKk68DTto1vFm11+
E1fNuWIZ6oXotCbUYgJd+FybmHzNZWVg58oCE0aSszICOVW+T+i8lcG6wga+Xf08
/KUeiAcHG0ftq4egq2UYqq05QJCBx+/9CDyuZyXXA6pg1qVzheTbKfsysXImd4JW
/EXQxyNfm28kzUItKMNR2+joPfxwfEGH5KeDwCwJXs/E94UMCO7EZ5G9A55FIEei
3xZuhL3mUYE3P+F72pohmK2ZYOHJsSvdE8zMXM6Y6TmPW8VXkRvY/PoSUyKzBFBI
oJaydQMh038kPjwCL1nzNq8LnPX/Yf29xrIuKIKGKUSbByUCG8jlJfZ1uvFD9XQ5
i9L3i+xUjnbc3+3uCiPf/kP/GkuRGhQ5gJcdlp5HADaLdIPK2Hm7xDgPmiXWoHbA
U+g9N1+V0x94VWIPRQOY+Zj/1c8d7u9btHIOqfPD/3H24LLnJCT4eJY063f9ShVL
A9Bl2g7kVfai2d31rnY+R0ehbn7wFDx/QtajTs1gdhgHxt9ZjohM5DNy74r/rIEi
u5nGiKynbC4DXJA/5O8GLZpv5+OEIK3MYLjfgdcHw8waQhCswsgBGdFcifIrKNqC
0dkJ9BtECCPFU8gUo8KIrhkJ7pjQUyIw+8cMxnbi2OgErv7XZ4H2fngxB9YBYUV5
4PvJtVEmnGZtDPqBT4U4mRodosAT95HMFO0L1gAm/6fOvwFOCE1V0FQxblqPfKih
gRKVi4fVMFfKETCQabDY2GEjTbhSnoMHOZVo9u4VcLvAnU/QuDSEEVP/2Wd0QGW7
ZNvLWhisI4lyDsGct+iopQHeEsp5Ho2Zrw1Qp/cJuzxqjDORtewSmADViTaK0/U5
BBv956IrF/Kq7qTeKPxJJLX5qBPlAfN6qIkerHxbCKX+wRAwYmisHr/4sGweryVj
TkIETG1rYsMrMg39/boDBWQ3pnWf6IZrrvvfLn2Cw9y140fEZiJxLLOPGC/Kcznk
22qgQWz2MPfNV6LWZa4WCYkdOnJi/GkucOdcJOIT6Z8mspnHc4TZot4FIZzjf/3z
coqUtdybp5B105b4kul2QuarTzMiyE7jdsrLA5M3L1M6goUn78sunHwWEnCSzK8q
sjhSEkwezdzUy1EBEgrsqf+o9CvVx5/6Rw6BwOmCWnhGLpKGiGlhHRHT6bHUM0JG
QBCTdfDp2FXX3IcNCvfXH5ZFXdGtYu+ckXzmROMQmP/gIbEVDLE0YIgt6wqezgDH
ONu8PxTw5uyq+JV62fDUFlQqHKzqXYcpzAmLIWG5pZVRfHKcHyPMTyj64d07fz3o
Jbbf1Lm4lgZKbr5v4aWGOK7TXE5xKoZhMWa9ptJuU/SiFGAQ5eZZjZK3P1IPXoDx
z1NyRMnI456an7cRLZR9108Ikvju0mtQS6WCithzy0d3GY/sgZu/c91EFVPtazgj
co1tcFdfK+8v6b5F0vh0t3z3vU/aeZ0ssDfx3mVr1PE6J16EbevyvTY+ekIm8WJs
zYj2/6g8TMDA11hY+xZ3Lwg9ZhUrs54Em0igvf70gI/+otf+L6ojCay5Y35ro2wU
wvZ2Qer7wBhnC8ZPG9FcH+yuI0pPUnWW0KD+kx2PeMACyuiiR6+SnP12pVYa2ZUl
pshGHhkkFqT89YKC92eIiVAIpEBCc/bnEK+b1EMGOW0awQLiTYKBbjFWnuIldrGG
tTD7at0scV9zgh1RP9sAQ09zIk53SzUj27KfVOQjL9TnPIq/qVf3im4LGci95+1C
QpBA15kTOn9NLfeKZrPRTaON0+HPyz+WF9Lh8jGfJSJnz/b2yU5BlQHOFPRzau5g
g+GPsxt6V5F6NSoYJzwm3VIo1OgYKd22zre0MWLe7QOkxzEcnGSy44ZoRtqnYsU7
sTLVz0m+L4xKlYyGxldzlCgfIFZjeSuSeimdGxcSW9D9blkzbFK5ISBMm2X1VIb1
o2aDdfPQzVMorlxl/o5kFbsdye9kQnz615XSLvNOeIXbRR7O9UnMhZWVB8ASAcNv
P6VFcaJMTSbdymOaoUsqRnllXWxWIi0F/9TO5wKdMa6s4CC2oVlgKXd5m+LsWI9o
16i+KTDxEIgdX15KACLNknwMB4DNXPLMm7QCH4WUE8fmy/5CW0/niQTm1F2bFmNd
9Vh2VEbCNdWhrLYTFin9BYr7qAncj1d+TiCuNme+lbH/dsDDRzbL3mRuZlD3xNHn
nKUfyMTC6Xc28/hu6emlEnLibXT4lfz7yHafgHZMAgAwQ3aPvebegQMnDStoPb13
BkIRJ9r82sxoqEILb6tm+B7H2Q3zUZcV6m2Ihy+b0urMK2gN8ODmWfA8jtfyec7S
olROp8FPmksy08j7CmYlGu0/k/Tuc7ycYkSgZEBT4guIAHO9/Pd1uzR8tllWuSUx
RI3kSBt9MF/2eD3n+w1zH9X16ChdBVF2naLvUlg5dfd6scVDXlV9Yqbgq37f7N2+
oKPtmeUpKcNyix+Wum6l8ooUkvPnyXi8LUcsxbTh78d9A+UyLQTE119xPUJNOrqz
GJpwEIm9aPB73DCfe4tGivj3kXJah4DTPBZzGT7RRAoT0hToeGyq2f2mbe7oNDgl
jW9A594sIwM3AdMttPs5tQJkLHZvN+dny8A3eVvBtJ+zFVo2u0NQdqbvBf+sHTy/
g3BJYCx9ZaEH5Ger14Ur5dFdExqyIaw9g5YaQiFkBezW9HdWbT6U2Tv/6AnQpbWZ
od2YQzWoog9JJj2HGSR0ino4YipIdtXi7W4YMUbrcCSAli1dBdjEzdSusp2Ezg4K
WnqRSvj6z2FqNqDMzYgDEcqLPawjjm4RGTsVqA8dMK/yaccxbQZhCkZzVONfRGTE
bCvke2s3H9GckdNLEPzMHv9wW9rmylKmwJE0eeggwdqxNawsWbvImHW4BJpeU8Ug
T5zvYHfEKdBTHI6R/T8taTrF6ewLwGRzMMsU2lUTkzI01HhuCcSf+8m53LZ3pBUM
ZAMVsRWjnIRT2LYnt8MHCw==
`protect END_PROTECTED
