`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2HoSlb4OKWgYPlK1cFjOOa9+Q2Rf7+BG6SKabsnSSDZNVv/4MehZ2Ka3ylHQRSzG
b58oqXbV9jvMYCjy98joKhb6a7m+6K3u7LpYd6QZe82lkZn8rko6tHGQDdZor8aX
fB43J/plk2w/P0EY0MeSD3Dzd3eWz26MzZNMCRYyaZHcpU/NBiXHSRLI6fC0iAKL
t37Op021aDHUM0vVCi45tV+a6ijAw35te2dptQb4BC96nxsZ9ufg2ZUMLnXmHRb0
hLuVYCx7s8fd4mJNTgVZeSP8M0ilE8jlCTBz/rLc369A/z/2P3npnFSHRAVZqJWT
eoMnmKPZvilwbmEJH0HrHPRTcZMN9MQ3UHVgvy/6wvVnOWS19po5cvdthR81RS3l
mRowW0pQPIxFKR0a1PZRO1KTK59M4QCqPR/tBh8qKoJYErY2iOk96M5f9ymOGanF
onzVARod2+fvXj2e+tPycqbKBaDkPRMezOkfZqYVe71KazcfOh530dkaDgidM24c
+ERPe1g5xt81mVR+JMylHuAgtJx6/q5KkctNuk0kv2yNQxAkBaydH+RRumigpPZ+
FymgA9CuXo7WgXk7d79pf8TRw743xjd+CDjVTCKSqv4GFM3X7LhCLS8vL0RYvK7k
asvbhGbDeJ7CT423hB6quzonEKN9py5XaTAgVCxklPZFO/9W81JLiXHVq0jfkIJy
zc/YXsdD/bcOy5kiekdhQIFMhSsiDAX62zlnK7pIzQEvkMXn1dWLDJbnHV/gead3
b5p0KifdXvXZKQ7xihykJp/rM+CaMnVLHrqtntkEwN7OfvsnWagbNbdNfPjqU34M
m+VNyZPr9JaOKBj/tFXF4XLbyQCDQatCRU2PtS38rxPJ+pamc0M6l5vqkDzPew10
q5R83jB4G/CzCkWlFHmDU2/xUhr07jimtzZwqxaE35kGQwH9qxhhTiO3H70y0gYO
vr/BANpQZ8IhJhs7Z9UBbNJ+ZpBI3VSS3tM5cODdxa+mGAZBxtp1MlybCg/dBg6E
ZJXqyeMyCUI4SDBW2wjPW4Z3sseV5OUyyKH4b/YXl8kIX356hsgUM4/YyRJPPfbk
`protect END_PROTECTED
