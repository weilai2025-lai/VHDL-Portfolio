`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TF3rsVhyMaca0CXJIquGn77OPI5xyc2b/MmH/un3EGEuHFvpAV+uSPCrz52tqJc
crNhgYxliIfKWDC6Nqm9KdPv7smbb/n6hvApYbeyIAVZud5bmtap0gyFHR5lVUE6
bVmR06pzV+t2ehrY0hnEn5QsmECMi/nHQOJfD73nFOiNrMvINktpkJSV8FezQuNX
ZV4ykP6w6FeW0WJpWrwVCYg25TTB/2Ll9VZ10j437X6o8ktvU3HwWEmnei7zuDCd
zvF0YF2kJL5Zq2/gaTteo+VcGrH6G/xhX4kGkcjI5uKHoNWv1v0LWsBR2QR2JpgB
X/DucRmITd5/CBNbOvz5UxQlBIwSMAuBIZLkjc0FUpWzYUwTQbQjx/tGke89HmlT
XasG//UOKiLZ8RZUS23BjapjubdMnMoPFh8QObe1dteEy41dsA1dZ8v0zmJ38hB3
lKnzF0WNb09iQnDN74ldVY6Lm7Mniyxkmp4BEYXe5CQKhkeHwqdVsIivcCYbO/CX
lCDO5ui/f/1QNmbkMY6j00UN2ybu+p3jKTqyrG0zn7hZWj9uUmbjA9es+vJuoSoA
1cJ3qKn/NEm3C9QcXXQ/pxZ69L5bD8lprpti8VWqiXphjF24JSWuLIxAiHvvqKRz
eP9Zc66a9KRqgUoxn7JCDs7jAOJI28r+8YIgfxQXsb2oe+iqGp/H8u+2WRDRYeF3
RFdh/gCM9vcA9KRw1qME8egM+wZDZt/kTh6tQkv7BcvjdM/JPnKcFtQN80tsPPp8
mrGADO4ZE9RvUW3+YJeW5WjIjSruqSh6GP5lOQ8nHunDYAPX1nVCHj45Qe6Ty761
GkoLM7xpHK7M0zFKFxzeYnZUpRwXsnM18A8DzhXF3tE0FEmBKqO7DiY4l0NYNH+K
7f1Vx5c/vhrR5j0bHdAf9GLUKJJT4oeYQoWBfNnp4LyRDQONN/xqwlUKr1qZacE6
xMgqONd0OChZyTL1Gmnm0nCMqPyA++XkiesG8L8GMMCNA8pIr7m0xknZiwsoysCn
0Ik6dMldLAscGkmML7NAWvpMeNsLbUHTz0q6WMoMbAL/I3pQY87tceOhZyzfsm7Q
R717eX9HDTIOYcOJugk3W+CtcdN42HOf9ylfuCOWE0QwTco5CS/PjKeR/JPZqVpb
62Xge8viWDNJaGDf1D2k6abl44nf//ooVOgJHV6N4YThEEAQTZZU+guHOQEYyawx
4KfpYlp4+cLabYg0eFJFQrEq8+Gv51TzzLW1EIeIlGAeIuiiPpFzji79bt/JRLgE
JpMzK8Nz/pe9EP9FEBWawKkRQRvUR9nhS3tQ1zDaMI2Ei9UivoNHpEqBRyM+868S
MIg1ex8uyUE9vBS9m3JTVSK35ns97KtRq669GtRxhNIecZjTghik1YeQLa76BQX/
zSiMw9cUWhK9y5XFY/QPRE5j2Hx+iNrbnH+lN+93Fn7Om9O4ehW15jHXS05TgtH1
OU1MB6FY+p2CBhoWdE/8+tVGIftLK7pD9aGJ/J+faTplegwzsSqoxBz29pnqEJmB
M280OdPHIOvfm9tLtL2rdKbGUtMd2KWUEqQdWQJ5TAOWFUrw5r5p5UZhuRLXF6da
1xQu+1IO7w5wVAXVgutujUexDkFfE+GG5i1ZM+IS+MqIpW4VvUQpLGhLW12f0IcU
ZRmKOX1zXC1wtDtwAMhdS7l5NBvEuphLWoljyjGtLRWQAoKZPoqEMvspB3eUNFKE
Qt/y0+pwsB8pGgVNQU5wQ/PwPNriRZLYpOaMofpb7rg3eBiR/TWEW6ZB6HXt4GVa
`protect END_PROTECTED
