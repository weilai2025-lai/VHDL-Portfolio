library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity multiplier_unit is
	generic(width: integer:=4);
	port(a :in std_logic_vector(width-1 downto 0);
		  b :in std_logic;
		  uout :out std_logic_vector(width-1 downto 0));
end entity multiplier_unit;

architecture behavioral of multiplier_unit is
begin
	generate_uout: 
	for i in 0 to (width-1) generate
		uout(i) <= b and a(i);
	end generate;
end architecture behavioral;