`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0q44R9gnGLt24Ga5X2rnevux9p6rytl8aeVBGgIkLhLF6i9SQD/r6a/UtCM/oVEV
J4I/1UA++0yyYE0Q287ybzdEkxah9Ipx3jwElJCPpM1K7vF4qzNpF8hgq4wiVSPt
mDhA/wvWiAcCxXu3livw181eTzY+DBB2AXAISXLW/uS+qzirJ+pgax4dJirO5LUn
x5a8dMeV2C2FitzFxmIaL0gvC7uEEymvrfbWBkzKQfAzbzwVd0v9/YRJCo+ZVe8k
uLIM633OSAiIVFx/YSBpaIs5M8CLPEP6V+Qld1XmNLoLi5Z2FIq5eW+cMXRdEfYf
VnpNUs7AZasZpqSzlvBqyz0dYsZAEpMfmwN+xIZh+eOubJasQQ4u9xk10JYiFCbN
L/vl5Kerv4/Kx15jgzdgHV8sp6ZJDgLzBjCi7Pj4UHfzp5JgEm8kDxnKhDb6XU8s
z9rNMP8eNp33HBU5dQXrxvQFv7Z2yQWPd3uyfW3ynlaJ/U+lQfl6e4KV00yefgMm
LEhuxbkl/CAXKTG/h2Qm8sWtW74yBgT3yi2BeIgfs1weYwYjt+GNPFwvv6/yIM2A
BBL1Q4A1glFkV4+JXLLS99eKL7eTnF76npc3lr3opoCMqaFshWZPIAdSy97EOg+Z
g5xkXsxEKQJlJHwLoJiGcjPll1Of9zTbDcDm5c6XZC/iR5UXBrjfRlmgTc5+4U+o
y7/l0T54Ly2wPLPcqi63yc51y0JcsrNEp3cXcweF5jJylyiyeLux2XpZ8c1HpJ1q
Bl7wpbkiy1ZX8cr5tbFPLBIyME50kSeJdPaxJBsRDxglb2QsXKf3c8fC3atGOzOK
pSzNgdOMSuYsVPOJM0QdziRJTV6zsneiAruNP3aItQp+fY2YHbYS1UynZyBlmPxH
R295w8AzBMpc1ud3WJt8moMrOQZrHGXLDRz1KK9sTYfJWfU/G+h2sM+MIgqqGUBE
ZyGikQlTpkg7kwjs5bq5gYB1/enmynLYiWl2zpVh/SRVgVe3xtOxZ9u0IXX3JSJi
pY8f59P9sB+YfU36JbC+FLuTLVRBM9IRLzo2+KsAPB2tZ5HArvOnZAHi1n2RwWm0
M1p7w1U7w+UXnl3SEhJbdEbWfX+aKjLJagZhHvxHP6B+WLPGuXrchf2ps9UrwaDz
R40ZWqTIIa0Vp2FtvP74FwGFEMrlnM2k4lxZu3qrWhPnY+LhdT1dMS6IhU7n6TAf
Z6DxCLMPzl3URNdwBVRUwPGutL054vsvT3kdXwnmyofRxmNvSTj1MFDBaAHF6AWP
CBQwDEEq07Wf05WmxGmOAuOw7XOXczQ67GTYsYVqU4Ttv99Fo/q21bQuTuIJ7sqq
9L6Sg2R8Fh3/EFqKLh4cOwVl759q1Y5XQcRNDzVcSaV6wE/CshC4RvZOkDwcKlo9
S0IA6p2ENUoLh5hznVqaHooA01Oy6Z2sMMWQljdhvloIBq+mcx1FRtRg7jzJhY/E
JFRUTfaAUl3nuTEen257iZ2dfZk1d3VorbL2f7lXoGkKRJfIa0lmih+v4JJgi8bs
QRKFvRoAomvn2gkCtn8v4tAOIKFn3rbamyfmtXZ8nA+68SQvqTNZPYgDQreXEt1k
hPOQEOpute/wI4KOqoSq2DLoV+frBVuWbM2u6bGB5p3McJ0KP++sDpY4XV9umofz
A2qcoIBWuGqSarBhQYlI2/o6r9XcI9VeSQSbQjZkHGvQqHfh5+S2uHs7pcrX6ZlO
Hq/ZvewE9DagSBfAazJkNhcxVVsLIinlLFRsz57lQL9yZCePZYWwl68t1/ooKB9Z
7bCXx5kgrbjb85KTn0GbeBAkytdubm8crR1F1Jj4i+gsc/4tj8+hC/Hes7OiHhsL
wPwP1drtR0dp2EWBqVrJcbTH7H8TM47nwsDntT0U7gGOkCmTo9bez1Q8770H13p5
H73ZWGHwFTOaZ0cvbskSVRfoSAZvB5LXmE7gK7RorgBGpb1PM0pFdz9KMfYKzIeC
fPQkLOyq8zwCutMuK4aG1jDvSnYOj7BvzcYq6QHAsYeDkOwjPjVBrdvrsDnXcUne
RTPbrf81bfaf08O8CVyb6YQJuyw9vrGSpLhT0i+uMoU5RL20uXkB6cE4KSCeNGU0
6lYlZdcjtEk5+lBXySmdGneIEG3B7/nji1czbgD0Nc8ByngG/q/aZ7tAQSnYujAh
rFyYSS6PUxUA/uyAPTgTuKBui6vUXlP0q7jJgQZXZ/kk6V9Fbqxks/N8gLrYjthK
T4bLHBQBUx0LOKgU8OkpzMu3mTQweZl+/dvKy48aeY0ZoPkxcYlrseij9iDi7BWO
tuEbzLm65AHG6qMFXC2YV/iNVJJ9PHeh85hIFLyO1yEY6ujLgePg/cK5z0BEq+nr
DjlFRz5KLTh0jwbmHgsvp9u538z2iQhaC9elsCwa0kJBlwFoqkcXxCQl/NXYbNPN
cK0h2ajUviUmuq1/HHkZk64zE0QftnmZnyqqb3qOkCaSrduMM2djqsdyEU5NmD0q
IFARkQ2ELH+myVVM4dRvslVgdAj0q5/AIeYLPpolC9wtp8kDFuvWKxVmyzCRsBBN
Q6cRM4isTWndKNq5NdOHL0ftIBbCEmLPp6k0h+BPp2tZHpkpufei6v7s+brGw4L4
Fv7XJ3I3FrarajNSwTyT1ndUnPk1lFAlsKnEHb151qug4IzW2/t/jJO9tqxzXfqJ
bDhq069IG5iwXQ3dOk2KJQ==
`protect END_PROTECTED
