`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5H5yYSqhFkKU6g1Utk8o+RUT2tmG8RVLMAdOTPc4jx7FV0YwTRR81qq3BgcJFJuO
CG/16AnyqhtqYNf3Gem0Tljjg/n7cVVPargb1feQ2HwAu8rv2HUh8aT9GRpxuisD
eS4o8HB69jqIamUEm/RNGMLh+ouOLTS6JaHDJ7O4r2QWtEiTggJbuPgQZMhjec59
CDkloWzU76TuEyEh7Zel6QF6dYVB/gkctbXkpnov0aH+OcKMnmH/hBqWfII+WmkN
91gTOE85FUM4zWHWKztguA==
`protect END_PROTECTED
