`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umnZVN9e/IQ6DpIAYYoRCIwBhOPwBQ4eDZfhIU8d0JJB6tbyvlwNodAu/TOFp6z6
fRqukkJ07uqQxpLTEqKgIJMvpEAdVfh+bHvn6yTAGR/Qqq7Siykp9x8h6JIHvUk4
NpuJ6SYpzAN/GOPMIk6y/DfPHjKxgCkM3Qyk/tm26HlcyCZJjjX5Ol0QScfJ3GWu
VvytGN0jhtIQqf5Qf0aQhshX6uct2d8I1Nozt0am4pQ4mCguDkDBgH6Ddkb1L0tN
bJI0IUYzAFvBi1ie2SeT/8g7FB6B8Ux7obd7yhjmt2WO/Xef8OtuRoX7K96crNaB
qJDFzWICFLLk+OXrw6P78Zutk6RCV//eCz6IeNxk10MQvUHB6XnarPYs0isUxf27
rzkZyFhYiNQzNsd2Z0rKHYeXlXic2e6Pmm89seJbgk+kYxWCN1/TyyCE788hamGJ
/WnDH630d6Gtd86/49g1Q8LkZ3FYphLg+3G9KWpbjzlh9TAlUR4cbfh6RoaafMor
QeahajC3KHeEIYkHmF286vPzXOAeS87ZaJ3yGyMOIbN0E+98Aq+EOaXXmFza9fFo
nx3ng5v6BTTE+QJvPTC8jO/3DD9sLfEkTG95yBZXZA5ovGBb1eur3iHzEYmVDHwA
ffQ+4ly5xOSu/laWAFKjQlvSJfSd9mUZHsri8cHKPF5iZSDBXiQDyKVZfmJveE6h
hYbRt2PjSvS3O8vxVPBkyT+25MXNiecHTalCWt/Pl34M7uF6Q8WdfT2M3CuN4VTm
iHYYcX0a5IpGprkA3BOEaLLI0vkh0W2KiZiTzN3NSR53lwRd5Kzt0ECXLbUwb0+B
sT2C4g4Pt5wboVaMMnHqRyLHTzkPJr+QTP6yovLjgwyOpZl+6GWWBnQ7j/4FdwFt
Jt/wrwzU2a9+wvyUOw71KdbMsy6V9KWVEe/oRtgr43rtz/puVZBuXTe4mlIH+UQz
u0Qd22rAULq/KX1Db1FLI8D+6VPEYq60unlEdmr5CUOeq77CrysVykFgikSpV552
TaccnY15+DBnqTwiZqHsp/jnwGg17Q4Toxx2E3+XnJDOP16AeGatFfYWElF/yIhW
OjPGenM22oNR8TaKdplt7xV3IlMYuKDmHPSUEaHYNqQpPiuS2KTMmEtSfQtFERI3
P4r1Ogz0oyGBrl88+uzYQxNFYeW5HHYvwLmigbrO7QKVKlUO5fqNgUHMMTehb38Z
jxkw3p1RfQRwp8TwUhbGNEE4WQDUUJgKCkmWjmVmwmIsPiR7/xDHMrfddV9M809Q
3LFLBOYuyE55+tEXUggCdF0YFlIk6YnUz5ES6/H3zEdbeYzbVW4SNeVJ34WWbHT1
XMBBP1da6rmw3chP+JOPrkLqcuMaNh+QZV52tmq8sAURlhefwsGRznTfwDhhpRJO
6gShRzOqlEvqJZIKOOeoRRiFoLIm3l831ZGyxsvrSkWHi43QmXnpVzZQo6EXeOeD
LE0PvJRAK1q/qTipyrpZQp6uSRhl5+bMlKi78tGrG2R56v5nFU2k5APV750bZlJ6
e5DU+KjSTlt1qOCmCEFfcMK702f3QK1zX2zp7xUjqllh7mnwQxNeBYugqge0uPy5
YHGLyQssvMYA8rwNmbswX5M/HK5Cpn+f0py8gV8H2r8YAhYZtvmlqMJQ7W+Axo5c
vR3THIpt5yQ1kZS5fdxeeTwlehao5Vutcvob+B4Rgg44lNBuFLzSjzU6pkGxFMQw
/JOekdflbWoxVxUzQct1Bd5BjS+WTIhC/abBk3uyc+bsK5K3z9+qNIq/eeygoI/a
amf+TDgZPTfF5Eg31vP/ofVS3ZSHMaawbDYtm0tm0UBY3DWF3qp3k9hiEw+3SXa1
RXkA8+HOUhlGuoj8f7GYR8PWsvIPoR29KFyH0Y84ngqAGlxzqZqNp0MyChhIe0+q
/GKPcJJcMaSwbROrhFTL1XzsGjqp74w5RHSa5ItRx+JAosPMa0hg8jfmfnCteZk7
YaXEF9gk5glnfXhrgl2whNlOym6lP5cnXD9XG4NO1NxKE897M/gW6Z59rftuXEOH
Hu34AQABHxJWx4A6ymG5PQE402janTXvH9EEHrJodjRTebUILmLGoymGTcqadk1v
5wdw14UaDVKgagT7rHgRspPJlxCM30ww/QIJ7NhRkHnMRn4mFXn0Vczt03//p8ak
7LEnhgfsyIs+f5UTKOCjJq8GVPNlpx4H7XGwTgEhu6ZXgkyu8Mx8e+cPDxMsk9ru
r7aazsUFgnpUq5mPoMvntTCO4K0G7uVpebpaElJ35vk1T8qtuJjQlHXcsqowj03n
NNwPTKnB+goLWaJPJ6jfdKMx6KzAQh8DkpGRnCDFSp5SfKpuMUYxr+46DdZUkQFN
vgTU0672mfZ/87A6vjjOoXPBgu7LPaJ2RCMSg7lcxkvJfhcBdNfx20f0xV1ErVuc
cHEy9J0TwtRX8sIwuWRazfTDqpb2sNdqjaXgGBuBt6PD1HChHu3mLCIjE67rENOo
dudd8y62/P3WlLM3T4L8fvC50s9zoeJUHOEWc/kLonHDGmzeY2e4WMiZjNUddKUz
amllmvmf5sOfx55kuVtdwma8KyriclWoqZnMLhGixfYkH6KThunvFmNeh0Hd8bAo
posW1nEZsm7LCX0hjP3E7nH3KqF3ysWg/SR7HFO7x64voOID0LykDWZ8u+BI2uPr
dzzsHFqBviqVPXdvpvyuSvFTlGT0u8lfAVfnSJ3Jht6unZpkZMlP6CqZHjZm9UAS
ABxlTW0b7guLDOSxudX6QRdw/MF6Y7J1UiKrBPPr9pT0M1Nk+o0SDJswSYWXCS08
PU6dLVWwZQrH2EOtfmpN8gRKU82lE69OdC0yqcZiQpaWJzFnqOa4IpRhFd4lZA0+
/oPN9DSglV0c2AjioApfKU6NVKIj1ycHi6x8XH4WwPFrGOUjRfcnxYIi/7k5x/qF
1+agKdZzpsIxBxF9Auf9jXInHOLhLEvwjPzL5Y7t3rlGyavTlpLxuNxzqCp0gaLz
kWVqsR5N3wsAQeVligmr5dyLBLJVPCbrw2/40MT9iOAfZaoVTTR+QxJuA+qNjU0p
vOwu1TNt6DCZjISpeJxJIxpDN43PVE8Ms1vqaXn0DrH7/wGIV/NK3LPjlbUPT/CZ
N13k/gOVJnhIDoEBzISeQVOVz4UNsiKk+uZABzxjaFwvrP2f3gNC36RJjSz1Bod6
2GmfsbBRV4HRFRwwgBscXEUVfEbZMNtmAOL4gclvNWx6JiK3S1NMpEF6XVA9ga6i
8pkNhO7dnjNFZhLP6giAprR0fQ2HXJttcGswOJGyAj1IFMY+hXbqhqLSJj+8CRUA
056dzG+XTgA9xaOI8hXagXyYLv9sXYbnUaJDV374hoCa2tSEVeXrPgB22TbaTPO+
L/XbQSYVgvQ3Emtkn5kWOdKGGGpVrDb4VAVgxrBE/FHT3MhDMcFM8PKScl7UN0aR
I6uyrSL2CJOw/WSNMhLvP8IN647aeU+L5DlGzJ6DDBjF6kJXKDJLdQDp22w6IUJH
xCMQPQOTr/TKP5hmRpWUY+U7h+PRjxVPYFz7YnCpFMtPl6Ef6loQILI+Jkmr5WNS
iVMtTHTCa0AkY0IBGxK4DMlX5ZzA0RjggclTEZ0A0U8xFcI3FhydunR1R8a/4sLx
/Ic6M3sFhZuHF5oOuHxGZwr2VQA7/VHpwUMPpZF/3VREVigf/tgM4+V83XAlHF8K
ZH5ASuCft7c8ZHUWqcmYAhrjD5ks6LfGIagtDDr3AaXoGcORffPWGTboZo7tAkzx
M7mXRinDf8XqJkIjyW0eEDbHtPfB7k9dOdWtMy0us0ozbc13nHIjHqB7gfD0YPql
7hk462WlxQspzzoQZX0wD0V5iv8kR7rcfXOF3SYX7ObvqYxG7OfJtsRsB2ll1BXJ
5sIiBvjOIlHzvH+89NomPhL4OadT+G18Bks1frDKN6BXDAzZv14zu/KiIoFRvNiF
ouZFctc03UA8yX9l6rH/KU+I54cVQzuKWanaX+bzVsl5bRrnc4afEpq49MlmgFHV
pB2Anx+gGAIBV40V7qJSryMmkVOpNtB5u8PQw+GbnZtbMGRqfv7YO0/tASwXnhr/
wpOyvO17m9f7Eog04PORqhwv3WuLRfsAmZjTrc5Wm2BLF3Rb3+heRa5B9UHwHCZE
oCC6zMAAmc5R+to7qqNan8nzyN6minJ6CI9NAw84+4gJNSF8zyhTAOkhNv3gNor7
4+8xNB4otzD7l0P+2UoMYFHCSJezAOvXqmvI3z1c1h8Oe1nXc/UXlwCWaQbnqUWI
hj+KE107GRzr3Bgr6kkx2o9+H2tkOIagnrGF0FQ6lHcnnhj6vXED30gobekdppY2
/uSp6YUKtKuUG764pusTk+AlL3ThfPv/ObAnI2I0am6jn4VQDbll1UNgeCeUNsxt
1qGM7hxdI9WUo3KSGnNrBZqtTAWSdKdMiIDkl3hM1HkgNoFnCXYfF755OrkluAC5
5s7MbauH5rO/ehWvT5PjbGVc2G2Ub/LE+REAJT4wZSdqxUQC53yRXSZMJlyLuc7L
d0BNVk/c4GqwF0qeXFW59U592i8tb3iB2ASSom/Rp5px4npmzt4RQeoKDygV5Zaj
+OYfGya/6RDEY2RJgZwSVG/oMa3ISU+pqLBslvDb11a29QekBXkyrnBIk2vBFeP1
wvHlXnRyNH4NRKNvZXypRzBqXsNRGqYQmGm9LgGZsoBrjKEnYwy/ccOqjUL1QV68
L0SXGdkjcSyTjhftJcZyitLYdN3L4ieors2aesrV+cDIgPt8Q58gVmoTOtr/kJIC
Hq/yEI1rsFflsfawrzc8dWrQfSyAPy25O+KFE2qsAffH7uU2PlWL48cdLmVTksEi
o7qGyqB/JaRm4CB1kblmtVTCy5OSwsvwP+D76X1oDgX4I1XrI+W5psdnPiCPBcuc
4V9Ij5ghGU68gGSySiWI3k3l+O3ekYS1sGCMqH0weg2fZD2O2adK1z+4T6gZsysd
1tPwGz3fuEaXfaEWiZBz3PNc7cvPwSNAL3bKXAuDI2xNjamNe9tNItic6hgwOWkb
uJ9gJU7HsovTQSQkg6aaelKPwhWPVtiNgezgf+agQqPlTn0mQJTq4Qi3RqqncVk6
3mcTDw7i/XqQPU9LOiVo3TKPUQEAAaQJBPSW9RSVIe+tpSO9+hNPacvR+FhvhBE1
AF4ewXamta4wI/l3Jzb51ZrXYazGsUJRr9GRCYtGHb2F/+Snmk+Njx0wJlmJi6/y
Dq9xdQPhuzHy24LAXA7ienllGFM4cr//ZCjhIyXhDkHEsJ9Io1u/khx6PxqsZL+X
8l7FXws/SciCtAuNBjEbOCEgYYa/6vbv1EEpuDtJvCsKZS8cYmpNlR3KqptfClPm
5IBLUWTa3dc95DLbMKM9egaoFY9eNsUaquITWt7E8+GoUj2hAYvegTelQEwHh/3C
GQN0ydtgFqztOkeA6dxCrUFh03UBcNUERx/BUaQ80M5bQdzy6ExwR0WKt7iyWN36
W44O9E8M+eTn/FkFHgEBYJk/dA4JPMAkOJvfMvQXhN1tAaFJLUFMMDU+Qg7TGlQE
lx+JoMSB1D1Lx6h+o79MFmBqp5j8N9lZ/uB5MvmlJEwUBXRgxbPGxgXrDnciQOhK
6nk2KZDBeQLU2nYpOZjTPVuzVmcXWtX3qCN5Sh1mgdxO+2bKRrKtT4P1GBpX9uJb
cAZaHllJl2ATlU7N7kWFScYzEEB9I0nMbp3HwTWUzWQA+7JcCYO8nAW1AVEStulp
ZGUJvTcx3S1BKO187Jp0j3YK+6B0eO4AFNGjXrsD7dqeYcVvcPMQOBmnMWC6oozl
hHAamCO1+/4x1TjHmzjF4PqFh1Gw4TLLcyJygOHkj04ixWXHt4no9itT5dnDivKB
ctx9vrXTJDv0kg/JXhmV0yCChxu7ySLBFKqD7Zw3fxQz6K212Yp7lzwv0/Vt5snZ
LnAcv5OATCnC/JM7+/aX3d3Zg08qZNtG6oJhShSL1PXp0I3pH6wNM2Cz2yfZOuyL
ui1nIDfTAVPaJPCwka+SU8/DFE7hatL11a61cLLbp0UW999AyIdrRSeVh1ztA0bm
5rUjiCjeApApoGsaDDgGkMi7o+K2IJEoDMSVU2dH+iFfIoPkjCwvDKyfC0R461FD
EiWuXBtLiJyqAiE5YKjTB1oL3wynckZlniVyjBmMV2RM1pESCoMZFIbw6eNU2mtA
nSye7RXkJyxigdtCE+ZNccuSPxfNbS9lIA5tKsEEjuHn5adhPxahGQPNOISIjdCm
SHcNtvOYirOlXdZixXt8oGMipS4OS/uPsuwPEDAgQJ6T5lW+c8kj0yl4T7i92mPE
/RbgKc/wpjXAuUPfxr/0ks/PNF20dGmRIunMaNeHSUqgtejXgaz1U8TvVoxgKVw/
9TZqvkB6eKbi0usx0KE/ECEgPcGbH81Sri8mWjRqxvdywO2YBPFGp/+rQN+RiIqD
+AU0Wwah490TZub1iV2BRZXVdBumL//WuEbkK6TP4PffIstdivThXd4fx0eCAr0M
E/FBuE4af5bw3nRKw/CxCHNAtZ4JLAMeZjOPxkyaX+7pK+I5/2jWXKOjwhJ0zzOR
XmgCwe6mLW7rsinV9qxtG6fRDMJSg34qKfXF5dnXEN/hD9x3fPwaTJNptWN2ObSE
OOgSqeA0gcPp3030GrlNm59Xab6+7/yboEgmCRDUe4GUil9OjzKW1DpQwcZKoZWt
jK7+IoEQLV7QgR6E9yMwDF6HS4WNR8Hq8ARARPdiOBHwX8WPY9yChEnB3IBA7bBo
KRAgxevJh6xzsYuFSI2H1iPnKYyui/3w9f35tPLqYGF1/zEKAIz7xeYFbRH3njtZ
g1cGVbbw1mdV4jYIuFaHL2YMV2ZdtLVn/24SCRNMVhy58sEZqKydoJyolCXTR+tl
OGYbh9y18TcTdLvmTNbMBo8ckhJ+Hg8niPkL/X1p5SXvEvzpX2+JuoR3aNK1T2Rn
gYxBtM17Z1on10pSRoFuC3UxLdVQBW4RykrL9zDs40unCDkKP/MHGm8ceZHtyD9V
2upILkOlRpNEY8+DYkUThKcjShHd6GgJHjnQj1ouZrvPkdWXE+svVimNgotTeZ54
cWFDbHCrqg416azR6Pt6upINdtvL1kYvOZksdjhWGPdVYmeyBnZOlMbpnz4GfFFQ
Ju2kLx79s7Sg+JXrofo54IJZ5fxoJCCHIDIgQb2No3lD4GiphjHr3o9QOpfsWqOb
n3/IERfRFuR3sStrXo01ci8gI84C+3tFAO/0i6Cz8pH8pqx9KsHNRobSj+xL+VG2
I0RRJx7B9dmJi2wT4gSvzFLWBhWaD6xjkpMfVict2uCy0xyp4R+j6Tx6uzym4mzm
dNo6U50Cub6Ol389yanX5BKhba9P8BQ9q71WErKQWrAkbGSLA92SpagGFeRmILSG
K9t38lOgizOVVCQV0wBgx9n8mW//GfE+zM8gbCrGvOiuf9c+mwthi4w3bfx90u2S
MPmnxLr301h2iAYPgDCk16tBAdR0pRvPojzDGDmAyTsmtQx9DRAwcas1L1YtVXeM
Ya0CUfMR8+sZNkqyOnZPX/jX0EcefkQZwbr1Dyh163mQP4cVozpLS8DtH0spH8DR
pm4DZBV7soYV4C24Csi/ZMRQzD+16SV2C5ZoqG74sm6grpKLtzycCb0x3DDQ6bYr
BdNcCO17fWM5KHG5kxUEx1yIGbRnQ3R+hIA/jaqKXlP3pGK4/UNdg+jl5YPNxG96
G1qzscd/tsYUYih9UkCfJqFI1cMDDxi9MHOsZTXEVqKzcpH7EbMSpLuDGG7Qr3fk
Oiyr+RdZtLOBy/pCdCbrI7kmQ1aWHuynD3+X0lTj0SQFAXghI/iWCwy3EuYnxKhg
gmfMuGOL4JvN+VIFAWwp5wGIf5u84cnE+Sjtecv5Vrk83hpN743tiPPy+dnxWK8x
C7MLBbnnNeVS6lKG/Lr1/dJBc3FVf8p945TPGCDxumIc83XqFWnvnGYGTt7FNVf7
cTQp0CwumGwSmfw8s5dl6dmunrYow/ps6Pj8QEU5JSBqi8me0sea7saihhFmX4xj
mGug028xfKg6KLMjcZ+NBSECL4+jFhE96AOGMn+2w+aFWz6T2vVUslrkJfowXdHA
UIdf66PDBrk0wEayQHxfil2s0xeSll9NiltDpESS6IgCzhXKNRzgLcmSvw46TaM0
EJKi5jBV32tWL1bR321VV2ns0HNO9AHq9cEfEqoO2RWOAq9lZLBn345bEr6UEPAf
wGAII9HjU4bsw0XKVGydRLNyalsoac2RrHC0axsXI0QQw9q1YbnGM7dpAe39h25W
5YAlWifU2RR7EI67ZodOYc2eOSrqBvlvnt/VmRNk+1ZLQjMyjJRWYsTW3N/7+81g
pOX/Da+QJjT2uGXIdHWvFj/allGoCnKxa414mJlxm+U5WoihcWk0PXJudeP+wmpo
nW7QvyvbhKFZAki2Q4yAIEER4on/wcMvEcMUsMmNc37x9wKPK05J+a2NqtQYju+G
6S1tlhTCWc2ua0NrvQYplonAR/l6RdleWOgQQmi3tj23OIHAeSAShgf4kxWo7FF5
SmdHRTElt4H/Vc+sa5PK58XIPUkxKksqa0ZI9nzYTJxTOKdL6YrjRf7J1Fihkykg
j2KtyRfL6Rw2Y2JFkGrpapNGm/tnyiU1CbGn2RMzqfhQjEa5ok3PeFaBt4Z88wrP
dfc7P71rWGXupy6VpodG2m/ADY54W0jz2UG9cwiADDFak1uys8Jm2tUW0TYpruQQ
dgzBG5dfC7Q5wWF9uTOcZcUSNG13/dd/MPweiZRCW7AVp+wx6s/cZ4ICnz2ztFJw
FCYUruj4dbvoyQj5qhsDJRTAfzr1Gh74ScJ0H+8UjdyI4tlDmWF6ox3ePmDG6I4Q
lq7NGG4kKOCSnCIezUPYbD69owk/rRGtRWXnYgJcDubg/YvOONmKD2CHiJzUDI22
4AGrIHwzStcoaYX4wCZsGZ2uWks3uWdq1hGJUiHe2QXUVAwpNGyGgCYlQuPRoJyP
aWLNOWlZyTic48wX6DqsnGH/w7G58AOYCheTJXbVP7CTS5W41xg1FzIQXMwGzlm0
eiK+dVu90L53rmiswuaHIM5Kw+6eOPVwi3kYEy9xOdrj8pLLM8eR5u5kIRJeCvRE
JIVfeuz6o8GD5naYEbsNFTvS94EZFrWufWTjcx2XxwbfRixLDvXa2JNltcsSMnpz
7HahrVmWfgoQCVQuEygqMBCJDgzPAEREGE5LCXDLt2meZNSrcQNJ/r3y/TCcZhfe
BPF6NE+b1Ms0SH0g3yqKLQSLegDAWWetf112gIe2AqTeABP7R5EGQpHamKBXg3jg
EroQr1glzKf6Yy0PCZcldVop8SsAtLqmGl1FFswMHvsxb7doYV0PRh23Pqpncqwp
2yZYBLEr+minDf+KsD8rU8GkEUuq7g/mkJMfSXCGAgE7KS8hoFx4nL/spDV2Gi74
zxwQh+xkgwBqcrbxr8PedULqoa7XZbrk7deK5GIrIdMT5g1TafrrO1qK9Y/NsDyN
C8nrXgxbQl2mYM7Pd50TVn+NONsvV3L277mVIP1E7VtAXDbrizZGpR7y/osQOrCd
u4dsUckVTDcak0YG7DKbu47aU9uldcrfju7noiYG0fpbxqZHrshc55PXs9BJ+ziT
Z6cjlFI8vPDXjAfVV8ubU1sNFuJ91DxIecicq/AbNid6BrgooyyORmCI7vH40STW
nFdA8SKEd69gJYFHBPfrsrSIseUqK0zkgrnJqkv509OYkdgbDV8ZWHpbC7BDOG2f
91gP98CTX6po0z9hDyabGR8U31TqQ7F80Cy3wDSIDnOmK7Qn8jCjWrMbvzfz7DgO
y8fwbqQVlGG/Q3ywoRphTcCdVvZ/X7kD99XXoOLzLvHPC9z1GIDgjKGRPUqq/WR7
y0TitVCtIdNcvjF9wgJZw6sJcRQ4ui5ayfuPhPGbnp388KrItWzRdWlV7WwUEVgR
2s82j/JV1Nz+bPoZ/F8kXF81lYYx3qPJ8FTNRt3sZBXUhPgRH17OGWSWbT975Txx
5l5INWfEu5SOMQzyg2agrsqDubikFFeY/b3nCgg41GmCzjzW3qBJ3SyvrdyrR9T+
ZeCPcPl2KVN/SwjrJLYoibeZwO3Y/M1U/lHlgw+8MTkYmlk7BFOlDb9cSLGWjO9E
92yDSrQhE6XvPC8lSZEDQzVv1Owj4n2CSJzpftJKFs0SwAB8kMwuhbR9iTCOQ/5g
dZL0vkeBC7e7dqLTnTDtZc2kPL7u2Vh6J0WkXCcRoCGtPJcAuG+XUDC9q7+t0LYH
e7nTYddgtGHbDkDpDI6aEt9p16GH0sUqrAY2C/QMTIZZiJbtXtHupvbxfMrDv6EY
xpP6lOQttDgAJSlvigIjZDI3tnnOSIeKS498Qz0uqiA1aPX+BjmOJnkuallQUyOW
+0quHFoxP8A3WfUErHSCyEfUXjO07OLXOARfg6z86F8LVknmOJA35YXjLzgqduFG
KtzGB8N22W1GDn+LyDnZWdz3qZJAIuvB7AapNkovOJY/8w9DhK0SY7NoN04ytYwr
ZyNQZTBV3BEE6Izun+ZbxUQjcUPgw2tQJnwk0X571oetU5HdBM7+Lk3UA3AzGEfd
liq3KavO1kvKki9I3Q2xSAPLi7vTva8t3klFDYKc03qiKc5dkRR+G3lUrbwAlXQ7
bNN8p2LNYQ0BQWcP7zQLpoGnW4Ss4rjq3+RYf04A2NjEvGQmOI0P1hKgNU+7Cd1t
cPatl+XCB72jwN2DAHoCV+q8K1FIxC1HeC/7GXJzmoI6bB7mOZsh190p5b1NTHF9
Fy8VkOBX10G3O5rw4b/KSlmj0x9/HNyDlDyYCtEmh4YrhZ1zAb3q2L1T6JZB5AmC
V0eRcvznQD1FPzqcQ+SrrhplhEpmy3oSj+GksAw0D+5TwRcriJMgdRowQPhcHOou
bmA2YjXPnuFkEiEZBpQBNJ/kFc5RoK3MXLKHb9KMCdrgU55t8JT2AxqJjoMqzSdF
VFvWhhEi1s4U9YtDICwo/gzIZtcy3MpaqGbV9JiQs3WmxUClm9YjRmS8vA3S4HQg
jFwBMzdnW16FFC6CBIAsRpchHz+zpqlvrVMMRuvpFLIA/bU3vdzvafH0DIXBC7/S
7CKh04zdgMwdEuuu6n7lR86g1fCxtowFlITHSGJmHM9ILdRHeIfTtbUS2Y0QZiVi
n3qpsHA6/A57qZynbXigHevMcP4wY+5nev7WCb2jfWEtzjUwOE4DSjoirW5wp+/b
nmGkQnztZz/cIW5pp86qkeJsdcr2rNELZ5JIINRGAdjlY0xMrdxUhhHauPXsUlNU
CJ+c+xIEH3SLtKgVadGQ/4M6FvR3Txuy7rbX4eyo+beFvnC/OjA5xCiao3ZyahjX
FKafZ6wOLc5h1qcKE4r5l8L2iFLfIfnHqBrDMdp+ExCySGcr8xRmDpGjjI6vL9cX
TfdpVqw9MIz+H9kbEoaGPezQBPJdC+ZiY+ry8W5dp4bifMRmSC1euweKR3zjvLv+
QOHX/nohpeQtHayKTXNL5PXXt1ILYz/C+Uejxt7jS07PelpVsz6NBYOoakVwgmci
mad1yc5iJNxUWtQ8DncIr2Z7Il0vn8fbnBJjEIQflGKdGyqnM0T9UGHbJGrL/Z1W
FMi9O6cWBGE452UsNsXAcernagF5BONbmzMT4I92EXH0awi1fQjWM4ljokQnDEWB
Ef5KH0XpAWm6xaOJQetDClb5OpwMR0PFcxHbJ8qWjbT2kwM+k9NJI0lK0U2bPcwl
kESYX/jRsGBZPPGn3Myo/5mRPcg5htE7gehJ8AM9nh9cTeZswbHNyUXzqREpg5Y5
Z9aa9GOR5md0wxg0I9Z3M/1XW3knXfmD/X3l3B0xxF9bvcgw7xPSK9BYbP8kdRCT
z9fzQ2KZMtYjCsHvSD8uGKXX/n9pMQUMN53PSh69eNDy5OqBm2jfOypizegt1hzh
LQxaPeSlfom5xbhcWkIgHhQPMKgtYwPhycWVm1XqV72MZlda/WSoT+vmKVDIi134
r3G+6Mrp7fGfj6V7mWzWx85kQ54AHjN0z62vdKMGJKiRBuOkRJIaUXWjruIFFTus
qS1vMt6jfbZ5hEf68xH4kyoIr70PVdC3FHQjn9UVYSNccQqDTWkYrH/BBuWY/WE4
LWvGg9h2gqs0DMqFhZGHIbbs073Pj1JPypsHTiltffvl/ZJyf2HowzOeWycGVkOr
ENPR98VlQc2cun0YX3VNprwZaekHwIISFpCsuTJxCAWBBwXaqlmVDn/Qx8EWoY5H
JCGZk1E5W3vOeN+H3dE8EC6YLCkzs6NpGRdpotqLbtHeZsQxerhPiMmqkvSRvGAe
PK8rdCZioP+fR/nLINIBs4NQmPdoJ/o9t61nYwOUwIJshJWfvc4abSvlDHnSfr6H
WmzmCQ6w0LiabXhasJ2d1iGrcFW6acOpL32IaioF6s0asqEpzblz/D9Zw+gY58a0
iJolfLY+gX6NKIoceZ5YL1BUCkAV9ZI8TU8ulqlZ7nP2KyMAX/Ke+2uOSK92Mhl9
5zp00NXsPnpA0OCRckx4ORe4KSj5DlBMySYUytD6h5AYR44cSl47SsBK0YNCcHU/
tOz2bwuW6Zg1ZOgdLuxOkWP5kZGaAbWojHi53IwKDviZVQ3HmcmF1jLkjUrym/w8
5tsmES08hpRV38xXdQZng0KOsQ1N7F63ogbohJK6F0r4MlEcT/gBKYtlGxPYTFZX
hbua2pkBI9SvY0g4TLtkSEQoyi3JrG2PuYKgOBuhydfWNXx43g96dWEd6GZ0Bgiw
00cz5oz4S6WsFB4pj0vLw00Favsr5Ldw+y6SH2W7n40O9lGgUn4OEpB3L5orlNc/
kXqSJyduC3nyC748W4owuQq9Zosy463A0akB/hLGuFXWF2T3IZJpRmAFx1Mvk2NM
JxhSWqntf3y9pH+tHfSFcHTXgZ8lsdXwQDD3ufClOLD00TiLp0HzKYqBDEYpdndy
7/UypfjV3amL0MkLAhnyZG/tBgIgJBsvunTkS/MU8RxbhjKSG3w6FM8W6ikd9Q+u
YwACu6Jfk8047FLzNOWeJpLYZZuI460Wummu4NWZUEaegqCSuNyytFgdi3W92gwv
WYfSbQOJvNOTPtd3oyQdYS9kmRMkUTzY6BUSoSd1KVM5hePWu7m7j1vLjjDzV/rf
8DifLCwCxUpIRRaLbRqJaGM5QJJI+zKaH5KuPvPwIBRalQvf62vi1uh5B/acGBv1
QoqKTD/uKZ1W3hzRPjWJgQbBBnPrsPhVB6wL0n6i96JqOqALoeW5tmhxfzECS1j1
Pgl7hp0OtSJhIrV1Z8aLnjh4PiSFiMVW01LMmA39UucsoGe/8esZi2yDi70sxfyC
JXnk0nMw9GCcNKuy4U5QyiLSFVZFU4mJdYOD1/opPPOiQl+dttdkL+xjfSiIbucu
roZmsmMXhGEfCF3yFWWs/4U0wEVLN8tClKkbAxCBUnJSxLu9aBvG4eYdy33GClUA
dxylrtK1XOi47FYWLfMlQgZL6+pW/CnQJjMlqkvIkCB3TiXbgI9qitfAhYteCe6E
JZs4zcjPIepHSZvwv3PeKouvRYT7FV8TZOtjsxOYJ+3NeKn1TBgWp3pBJ4VAEBck
e6eqYkhIcFJkANJyPxveNn2rM4/72rqFCd3gyU8O9aFbbmtUljhdBeAaE4PWZ2Ff
kkNidPDO1fA60dZnbmgqDa2sQTyZBLHomnA5J1xYvx5+20fHBD0xnmKtQCztAmRw
Pt/uugchZYHOgCLT5Xr+8WKWspDndKHpvN3qvnBlRcMopmcscRtXCOIVm/KH7P+E
Vz8VMIFF69nm9bGZzPg9ECuPdYqY4iKeo6FO2+40/VHrADGv9qR2q1KBIi2+e2gA
ecRvU1LE+4ksXAPkiY7I8FYyXQH1j7MnXvdLXpdT+ZQdBc6Axtmywng2fZ2F275g
wu2QrPCjKz5QV9de3gE9sOXQUSrbdn/kTXCdRJWG2+fGd4THCH1BvWoCe38gliel
qm/JIudrVs6E55DV1v8rI4QdW+x7Gk+z4hTdP9gooJnSixKclB4JMbz1cBD/ioyh
88PBDjoTsLWegc2xkbVzJG2zHMO/JgAfPFl5DR5WM+AZbSlJ3r0k8qjjh2Ngdg6o
jasgrHBMhh7d/qgb8pD85JzapVxnS8bRVQsusV2mITI5hxgl3SCazf45xVY99On4
UrpUbF3iDXUIyKmFFGIj5w7SZUtpz2bhhWVulGiksYZD7IDfLzkVqO/0dVF+0hLg
S1XQejSapKAh7Y2AgPaYYUzGE5DBs5v4V4cpkoxADLSmwi7atPO5XMI0hU3RZGIA
8/Cx8TkqYwUcCSkKUsy6Z4kEInLQQRtyti61SFAuvv75CU5V8y6KeA4aaI2wlMlM
yXP3e5XCnkBrjWNI7JbNaIWWy+5OmWPzOlbrII+RVifp5s2mnd7DjuE39r2HTZqn
lJgR5Q3l+FMvc16hjRkw3TTEUkg/l1y5lMvdE18jqgGFV9SeFh5SubXrJqV35rgh
gQUC40VBB/D2aOwXe5fXuVj86/PVjvTqmzU/knAafQPW5Y/qk0ZcP6H4ZNmXASrM
4Xveb+Cazuc4z+B6pCLqpWmloBnbQBIsmAV0dbqP6btDPGWFNxcYiCOz6qzjs5Zu
AppiVhdzumS8VV0b7GmSBlHvZpV7DVUWsSFLQXQX178y0/wTRcjB4j7aiJSSg8U1
Yp4ljBUxH/Yk2Ug2G2pRxHr+I+zdLtonN8U15OTxGgqpr4A+BORWHOBFlkn1Sx7e
/sFBuniBsPIIm4g2LbmjoKxEdc/N1kxrLF2E6aj7v3C2tG0us/E0BvGAFv8V0eE+
9FV4Yo/y0M7f76dD5cUqOzHKJeqkJZEQEWfEsbsUbwiALX5Yt77BRbjhQj19KL9b
Q84dhZypKVAd5+1kqsjyqynAI6LYLHC7Oi971BEOXfCOAFhX4T0CcGRP5vmWUCWI
uuZH8zhfXQ/tvj30oZRObAQA2CNpPKygaGrgdNZg44fDwGt37lujOiFo9ubeHpUt
6wwml9z8VsIvJWj9mnRVMfDuDHI4J30wccsYbnc96MbT4mOLze72bsCA8p9RwHpQ
Yoh/+tCE4+Fwbvpp+OYg7i1CmU4ltUTr6hynRhEXHeMwucM0JViNfpFF/Y5F+uqt
TER/Rq8AZSXDm2DZ5cRwVXrxCUUCWjm/zwbIOP+uLcPPy9wa2v+WLTR113RIENya
hxgJ7SReMPSwUAj9hdtL2Z+UQFzsVkTSqje27OhAIGxSfHGMuyxzTEsifWtl893Q
q6C+IYSWG9qEBbtzlUtyCYfZuHF8X8GgK9xSwHy5LBVaajwoCeojBob6tXVq3Zx0
KYJ/DeuETElbu8F+eNqDqt85SU2cQwzeKlSvjjrgD/abbX/58aAZ7+rKEAWK/Bnh
58cTzwMH4ijq/Y3ZZmMsFOgL2iJ3R422JWfEmzSBmqoB3A85qFXWv93Efi+hB3tN
kVr58nSuEWgCo2OFOWraxCVJRMET+dVIL+zzPwwU7dNK2ZkwPZbbEcBCDOnSzYbv
QB/T0m8nqZHSjX9kmHteAALCMcZl6kAtprc4980tAf0YGinzwZ6PY9swySd8iqRv
WNjeGJsMBN3KU+SnkoEY+wtrgRwaPUACkcrB4xa2yTms21eChXpLxrp86aRSLa3w
RVGB021+abZAEH8SpUjNzojkbqUefFMmYRWEig07yKGcFBPezAArITck9OIBKnQq
1r5yioz0ZBxws+u+vovw2dC5Gajr6uwCotXOulAdEU98oTeAduI3jLenwLN2aYey
egc2BWTpXhBDlpl6y7nHDHy4L+W2/PqATMogDM8VfMPYqxeUBk00FA9+Y4xRW2Ro
HrAqjMXaCndu4Q2S56xlUQq/MkuQxVM4AFCbFtGRMCSYhhhIGtdQQNkxOpB4ruLy
l81RtKY3QNreRDjY5QYS6DLQ+FrnEriY/VcJWyaSW+1ZOtEa77S3ObUeFv2JHMjX
gvf/JrWKbVNTEKQBhBini8VksH4VyJSYQ0e4oxf7u0fRdHHEY/vR9a8OZ32sn4ao
1ybHQfpyWS7Eks/LbxQirbq96wrsLJL53w91uL2J6r6VUBBFX6TjcNDZow32wCBn
B3IknlyW0bYgey8Zdt0ftnWseoG5xY7wog3Mv1yTtmpoUEWL8Ywv+CaHnshNfnno
CmdMZCffCHWrqgscP5Ksk+TmtaZU0I+LWP3QA58E5WFINSXlSZAqVjlG0gI6m/5F
PacP90rnb1X6NlITjz78KWN07yoFGUQR1+ky5g41BH5qdbSt7NdPr2EvrD8TEnbp
VPeEmRZ/1eT4Sr4xnvbc0htLzlmV/+7TsTn7xoaaIomyQm1vtYsmyBiEgIUF/NX2
igFET6uV4pP8RFNe6t6E/9Ywz5x9nEfShhAXQxpas0QRk/Bms0NEa5u348mlSoyQ
Vj7Q7ZTqTig6ekeg4LnoN8zC2S2ugfa17OqrFQuQqksIevB5sA5U4A2MEzEymMis
gW6pHAHCNO7DpuQA0P1ImVFsbkiTK0grkG1FwJlLM3FgHMXwiaVpekbLi2DKhL2U
lf006+DYLsXEAhdIA84oKVamlC5n8/QHkAS0bmrSJ0HPQXBaT3lyZ0IFEL1dHDD7
+t9AYTS44Zr26r0EVvYZ1itpF2B7kj67V6s2vlGaJW14YkC8RWid5e0+aRkPgTsP
KuRSWeoyk0uUN+rT6wH3Dpi3guUNx1yI91dlj0SYXtncT0yb3bYstX9OCQGqg9OK
GbEGE7fDC9uyXLlFFzVEGdS0Z5i6t1twV5BlatUSLnROw1/JCpPE5ryuYT21hLQ7
qathGduftkjyA1kRneQQpEttT9BH/bL0hAL20tbTWpuBhgkduMudhOBpjVlwxomz
C/KcmMToELKPP1kPBQ1SN3cPRw7nBcPeIhSkrYlvFfvKycLaBltwTzWIrug6HHwE
R6lkQ9vcxveJpliUciBKIkyTgbUJRoVcxigJgn5SXwRjxbk9bWvx74q4uNqp00Qy
qFbNYl8YWPgYyjBiCZik9fzXvYH9PZ4pJ13f2bZ8ebjvcFN6CW2xGHjXFG4ud26H
Pwa0d0LCqbikdB7XHb6Nl5IkBlQflcOZyvfuZEG56IWazoKUxr+7A3DcGwI6di7k
x7m4FirESxJ27AThvEo9I6yU/Mc+u5f1OrOEaFXaSDGgiMkZT3nqj/rOQDXxVY70
eaoQ+0ZtU6/e3qVfs1Yni9NJa3/cMwsxAoc8vcfQzenFX9nkzi5j7dZZFWL4ronz
jcey9jtwHtPm+2zLcHxs07w3cgQJGoz/wIviu9WUOJyqnQEIvlYScQIxyBS14tc5
uZAzBAJmrRLeIA9N5HXprBEIJvHjlpT3/BE/CdocbfNtDmII+JJbDvwztXbA/se7
LaY5h/OysGWrebiuPdjFdwaWGcTpLbVmeQ6wtTPcmtfy+XfgOULLUsPiR29jg1Qm
jVGbaaavoK8j1lUyYYHmn4wE0hxOsI8Fegzlvi3k88hTKX3FZeHlp7TJ1Xpa0Y0O
hF2lHA8bd5U/TgG8+/9cXO7WyhOxol6qFKPcdjzt/U9pCKaMRip9r+lxcK38Nb0v
ycu2+/n+XLwmWzQMBeCpTtZdkSkit2Bg2siNoXfxwBuW1qyzRanpErsDiub94ny4
C9ms7l2AaqzJNn1Q3WSKJQ+gZ4RiAHngxgejSGuoeqIzhFEeddu4+2ge+YcPFgHR
7N8WmDal0bM66BaJj6rp8FYtUp61pJP9E/O06LNO4yZ8u/9u084Se+lFzrXfGudL
e11XY3Bn1vfxl8CITWfQktLgs1qIAz3oyLR4poIKPEUYb4kofzQzn2VesLejqJt6
iQ8TsQO6iNweV6iSA+v2btkLMQHi1P7XVxFeHk7z6vHe9hGTUPfbA2xnj7y8UMXq
ArNMnFPLCSkNNVlQSxqpanjRFeSIl1g+6ygeHTh1FJfEvtwrv2yZI3aEYBxqBHlR
CBmKSvuHrr0aCvclReE+MmOJE5KVr0HU7p3oUjFvA6HyJ3KjP9h/lQlZXgfRg8Qu
TDO5cgqzWB9nfQ6tmxOH/XBCHM6B8UaDbR1juc6nRmg60AbbOx4dRSmDB8B/yxak
usNSAPByrJyzC0qiRlZ38RQcTnInNJCFXKpJ5l8sqCfwuQkf91CGaieMkgcT0P41
w/RqrdD2i+lfg+6RrzevZxLkzrUposFVN41kVZyQOvtMDgWC/vxJelugmWSFBi+i
xBHB5fM3HK8aM/1WsqdPRlb8zfbPNIjgJOaOyMvR+CdxRI7yUf+NFeZQELYVIhB+
Lhoif9gn+OHxJpw/j6HRv1czRGDU+eidvvISxXt8VZZdDl8U/bz1fa0ADU7x1gPV
kwmr9u9cJYd9IEbY4D9xl8TE7K2S6rLha4gAvi8Nx2moGEIhsvVSKxytCud6/ty1
2zJi4/0bIAQ11GeG8x5ldlkyhKwQ3LBxV0nPTlbzoFNgqLTbgahsdcskuaT4vA55
hJ454ZJH9e/oM8kIuBbt9JcOylQUa81jwi6Z+B0G7HIwwhm1xulwgrYlAdevmjN1
akFAJLY0klSjQBqZFyqYsbMRvRB/8QbijHjXDQItQxs73zRmcDwvqcEZnPnSvJ0t
rNeDtvSV172+gga2EwI9sxfVwfIJPoRyriXOh5M60kgOcFqeOWwHlFaR4UVeM3SD
MDOwg/VAbWUzVqCiCzr1CyN053UxeIFCzpWjFU7lTgSrkiI0VWmRg2bO4+nesYxz
+RBwEGToCto8HRzZSv8eX8ygYxFl/nTv6KugBffX/vVH0cMHY7VlRfh3DfbuYHBM
y+4gEBEIoScjX9wv/D4Mhu/akiOFR0+G6J8N+EgrV31B1mhlajaxaDF4jQ9a4hUP
iTgcOiZnH8OMVo9SaEy7+rOnBguMhd7PWdYSGZsEetcuMGuCPcXlZTRwIJhKAvOn
y5qHu75GQmfHpSbTn/Hp2YstpRBszacohEJzfvd5JGVXxwMvLuWouFpaLsJUWUGY
ZxWAp64ufDIkM8gi4QtAJFKvhd/oXq03mQoMZURmAQ2+zOKdk4SLa9i59AhDuF4r
SRt33YWLb+/5fUd90X5720laUXIXrc0pzrDu6vyD4xgrIF7QGF0IZBQNATFshsOX
eok2Zys3yxzrzK3ecAw2nDLpzho4PrZ4Kk7gTzZvRLGEo4MVb/DNFh32AFgdVnDc
oALct9GHVCXvFVxwm/ngtbWs7BkmxSTLLjceTmew2EuCCP4uocEwQRI9AnkLabGt
RNjmptsXe1wsBdXrPaM9Xaaou2wk+ftHmY2qbAgxFnRFtJuH88j1BdCFj4b5AA4i
yFY1O4IEvoZEpOHB2TRqq23+UEyRK/ykion1EK22PJF/JrsFXWL3drDNVoZo1wTI
l++31zS3rdiWfNMKJCmngyKc2gbW22zwXcKWJ1r+7n+XuumGVNnNOnZKDXxgwmrE
pPaCYLDOBjW0ohJnRqoNgUerSe8B6Nqymy51n8zYhsfS7i66lUkzgXxa7Z2L+p2b
6jemJbUtgiqPFclaBCbC6VAXVe9d3OPMYrQ0MJWOXGYRbULKXqPuGau1O2nupkhK
0rGK7HDl34O9BfSPTTUry2CtFzdFOOhbR/RiwgjS+3AWgbD/N9UaumbQBxWxQ3BA
vDV2+F5ziqn9BJGFjpniKmIIVRDoCKy67Nd6/J/M4nOON32G4XKH0quk08ztzv/C
fqHd+DU66GlbD9NvVWZdTFoRl5iKS88SZ7AIEOORTUmcnY79OTCsIQ3Z8LbWKtSI
xgqytQayE/lrz7dvmum2JMYXnQhSM/djRTWV5bVtRpB1ulaTWONFXKKHztsfecoS
PtlkUNq7ubKftavQnWdVNX2G9TQy2dd3m0F3sa3ZdaTcWqPVdps5X97mnZug0rvc
g2wJHpUOsjkUt3iQfkUfH/EqC9kmolzaeo2+XrnHz0EJI95TnCrLhAEeWVffxjNv
csyclxkkJu6OSPyeGwjAb5hqfhQLq+/igwfvh0YIsREjdlcMed0D5x4O2vDu7Jii
kVIIoKFbI0IvR9mD1uSEFE7AuCi1LjHGcn3LWpwguDK16h41NM3qW+joYQ8g4a1B
jxBRfGjBnQRdNl9tbTWFBL0U8qT+ptgcR22hL5IU1/Oc92/lRzD4mflQ5XIUKoBp
QrI4ZhnpUjmxjfYDhEIETkfPgZKagQA4PjGp+WtJCGIDD5DYo29sd2fAIHEG012o
YgMtUKjOiMbSfkpAF9oGjXZfc0vL3jrhGvH+K//McISIiY4TR9Z4FPvl2W2pSkZA
k2ufqYx76tqU8OvddjFjPQsRlXH882aPlXwWutxxN1Wd5zdzdNuGFAk3zdPj25Ai
7iglgeupzkgAU4S0/6rJJtSibCc5CdUoqrHQUvQoiwTU90CAntlfwSqYwyRjK879
PBXDe4CtQp2xZqOwxV8Ow0oPHdeGsjYZa4ogVDV95amxPSLDp7t8vqjdqd3JnU9s
9bfP1/U8qqEPN6rhVnQw+3imPRlTHblh1k0VA/aWV5o0fP7Sj7FotYg1muMnRnYs
JVImZrXguPQwGRb5FLyXdFc51HWPnsJezg0bcFmuGb6XRXeUwuzAnNEmgO1iBk3E
OLHA1v+55ld71opCG8c5ofS/6T+90pXfMQWV0QZygUJjzMnZ0l1aEMc65WTdWfY8
XgSPQvELUKko2dPNMkuBymXkdX7weaKcPiv46+mQsPsPmzLK5ynsmnco2R7+vPKZ
yi29d4ahdUQQRBRZHKeNKZCiKXSIooMKbb/VxM293wjOvgVkzn3UMWxeJ40B72iz
3hBownY9tqbfnYcOxkkmszEL+46a2SFQLLCO1eFkv0M7X02FF2k/US0P/iDTjA31
OONzatVY9C4p+IfRTGlVRZSAyusrYdfVpkwPu+RWjGjjStdqXue5sDBCkVd9ugm8
cosn1E7/tTP2O121YLwcmit3ipEj0xXwptAoaUBjQ7c1IjIEOKv2fqSXRiJ2ij3C
GJJ/0bQlDHdU237xVGGkY3DQEXPMP9Imy7xn5mNr0dXdgtgxTeE5eeo6NY+sUk6r
Y37JNXjafWcdQ8yqfa3SVCMPgj91GrKo2yfOpQOWW8YppMPV9RRgphIABtMK9+Ef
aFR8rtBY8ghkoYgC5xMunmpTcxxzr20f8hFrEVDQP/aMkHDAgwM3QAxJv4aa7lWt
tr4oxqeGiWumc9d6pKDHJa1gqdshXUds6XpmFB0mVEZFRuWy6OnsO6a0ZVQnCCDx
vHIExxC5X1duvsTdraJL9ChGr9+Y7eyEKisiDkRE4XdMOsQ0AMlmB8ovNbD2tggt
qZfFMnxKTJMH9b6iDaLLLb5I1rkX0QULEGILMP0fFEwVaAOCQlhY/xAyb5pd/9sl
w2z4LcC4y7AFnh4L7xICKhQkLMRrjuZJOnnj2QIR33TbRqPa+7oSq62Y/nU6Fsy5
4/7Pnztk2c63RRYRXI5YuSjuGbNyj8g3giXpt1VMCk/f+VFYjJ2BxZgR2Ty3Ya1X
XRaLaG1Uq+i+BqfU2vXE2zBaoxct6XkE6wgdxwRwz0dGCP5OGGzNA0XMaHkyLgkB
dRxa9fyfERv+ZQSFQpVCU/Xk/fMvGBiEtWAtZs4pTXdhlHgyWftlatz5BOJ7pmhB
sfbbTK+Ul/Yvn8t9hwqSAarI/YbsFJjbU7aB5Ljvu4Uizk0PvV/tV9rA8TG4K+hN
mTbIUtzPIoh3yCGBeMjJDRD2I1LsmYoDg8ifaoFaubuofrvfV0vnPKwZElSFEeWU
PlzKq2WnRYyEJhXyQs2nenPkAH2apzhQKtXRh0uqw1BfG+aixleE3fjxrXsjOIWi
8w1U9dBDJyPOH6stZCOk7ntlvPEEBcWMaVICbPAJ+73HukLZEfIq8nf1WNDGKzts
qqAGN2LEbdg4cVqKtk7b3s6VMi8WsWat+K7v1R+4dtfZgekNefU69nTdaF0PvQFG
7pWomgsTFm7zE+lgLVtz+2KfPsGc0Q8EZLrdzlN/U0S8PDxSaKT/GsCbKGCORkOb
GwnJGuICk+8Sdt/8XuGPJs9H+1kKml3GKQ3HU/YjNWPm7ACTRUxOcT93d4bOt+GX
4FNHvYHUExpUSqDZgB/hLX20WYj/SicMYvf+k91cgYtqMSBBhmJ7fXl52CB6tvem
IZ8P0lntv31dOekbhGKMhhRn89CEQt+wklwpZMvmavBD3R6AmubJNXDNAC+5lmkX
ZdgpWpCG2sOwEbOyFjzqBxEO/LQESDl9uPU0bTQqMhDM4AjvJweQ386YAiHeTsPG
hsJE62jMP1hHqcARO1lNpw9pWGNQQy3AzyTU8l/j4fN70oyEE1IU5UTyvl1RxwLu
az9FWzDLBw/pvoy3LyfUgeu4BS0Ksp0lVxkcD55zZr0vkqm78mVgvLuD7XCVDWDU
fbj+7Ga2PunJjvELE/zOOx+i0Tgc7I4LAo9f3O702UszNYUJqcc0/WvKW2liLMrT
i1U5vMoE4z5TxCptC8E/LmDJjKHHeQZ4fmD0QBE7o8AXCz/1HtqqB6VvMmF2c8am
wrPTZC060rHw5FDLOXqnQuSm740FTvD6tdlEzMDc2AMP/j2nCqQkzi/vxR4MJsDs
lpSfmge7TQvDgqYyiJpmjIBAr43ac3fdiXE+6tdgyLb2SjsDjctiRq8d9gAvbn73
Qq3/sjb8pdyEgkeGu+P0PuU7fOqexAGBkuMSmEQ/zHG0PJ9d3SHcJkoordCAGoS4
x6M0hKA75qRzenttquAXAcYxjTNOzU9iUF6a8Zi3ty3TAGUJg+Gp0FzMz6l/iBOS
BAEMAolIrMeffwqv03dDd5xemndr2E+4q7isu4FyIDzts4ernZDpjNAPIVuXKKit
MtCVx2SdSaUdORqwHMswrG0+KWeS8i1hn4CJXJxyNYjvPPLRhwyjW9sJC1NLIImo
EWC2WNR+OheSF+6q5boJ+q9BrqMEBc/zrrHQDz1p2lmj7lxg3/k6J0rf1t5d0hF/
sqTMkU7YhBuRd6aTegZNtZ9x/mI737Nu0Ed7Ht8hnDzxjn+rUJoFPHbk28EhfbT0
ckbMud6KwEZN6BFseeLiDi0C+Qb5hR38n/d1Huuoe/o7B0ifq691yYRMbG9tU93z
GnUE4thAJBWpLEhpOaqPTA3HqjBvMyYZGyRahTl+lYAP3EB0idmf+Nh+kU9dpaWM
14KB9jKa2qKGGZ3jh7BK7SqdZxisz7s5P1uwhEccn7ozHSLPoiyjAY/nQuw7IYFM
y1b4UYAr5eLOXUE83nzx/WAp8baDfOmVIgkApN5h/I7Gcu+hK/v81T6LH0xr3wMH
Nn3u/spV5wzaNTH+1UxEkzDdOupTUvR0YLaxBuNJibc+V79m28yqzFSkB1oqG8TJ
lcqW8vEIg19lxRMp35jDiuQdkfC/LHDcSUBd4nPCBbPxydNKN1uzkzakVaELb0bS
JwOZrtWYg/YFlnilcmBm/AXPoYydyzZk54Mj1AwNJwTculgYgwbAeL4XeXm53KD7
kAESXdCaP3tG9jpWlHC0igb3f9jaU0HAQpyIyxqfhysDrGk6oPLFA5o6+n89IkGU
5mUYGKejrOtg3Kgwf949Xu1uYY4h78IYfooyJ5QiLU5aDJY46ZFiuQcTSi+UvzTb
lpNTgHcCUX0givDVa/3IA8ngbnuT19+zWJlUtAdlbpZG09XKJWDYfr3+VwT1dYus
SpzegKxFFstIpDqlrV7efeZFbC+I71QWnCip+kQ+zoSCZlBeWQyczd6K2MCrBezd
8y8uaxbdSDbvaivdW8zXfiwS/Pc9eN/LxVaHoN9cpYbH3uYujm5dSVt8HcbDQ5m6
M1Jh0nAQYhS7mOeD/tjYdPc0lIA63PLwQGoxW4gShlvCau2cvLSyZ/y7ChJz8lXD
78z9IIIWOlYtIGKYOZUEMFdhAzVVqLWfAC1W2mPX41dZGXlnRX14ZhXayHp3MNrQ
EWNaKquaQ5G4rUxhRvphbNXxzjhpwRYt2KLSVL13rKTDdZykNwM1c3nH2Bc4MExZ
oeChDIf2Es97eP7XQYrJkc6aYXC4zPDbnVrNW1MQJt41K3eRLM889+rfvHoGb0Ol
X8WGaoKrBqO45IGDFjl2NGDpUooeujw0iX9XCw0X3VPyTdZqTMKhzgA7rQufpklI
tPGEdKVuKUO0hk/BIvU3/oigieuddEVJvYMRbifKjq08PMNjHf9tAesgYa+FecPr
Zq7GbrCqWZ98fVi9U4gafvARGMbc7pYspi18ZhDeRszBx2QImYdt7ucJmdY2cE21
A/UoKPmnOpHz0cQ8w1eqz68GVr44mM6IKnlEHPSffZ1CNqjCRcH/6aMLObNTctD1
nqiUNfF7K9jkgcdAJRX8cv0MdbFObikMDyBxjwZn4N5OYLqYpjCgfp72pGINowHW
sNjrZpjMEdoaQhKDytM2fZ4m1NaHRM3MXAogW5CA1kyInKG6LAtmaSl1vIHSa6AU
Aoo7Mz0PEF+5WnMmtkKhsIztfF3FbwDj1gQsHfPoVypdphJ46JP5HTQ5wckbwVlU
tmKjOs6ZfqmPCA5fHbjsuArd5W4UR0N1bXq7Q2FDuf0=
`protect END_PROTECTED
