`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
soGActVIlCkK1MxiQSwZthHrFrJyRjA6z7QQuNJUd/O/XorHBI4z8z1yExjhWNM9
qGxljdr7B9cl0vViAR82NEjPasWt8t1LdYrld11H7H0FKIiF+RqopSLXA9vA6xMx
SG0zPGZECGs7gy/GBBcBQ0XiLJkVaHJGHVdFqLpN/0bVCJ6M66KWNE9rcphE2H5o
GtD5rxx/ZezE9vmDUCHuRqE4JN9LOfx3051wvu/MN0vtiYjoh0sUzdvmpxRGjW99
EzMOnM2Awp4nE2Jr8uXi7jjyimZj842w59DDZ7LeQ+UEkPy9lmrFXcyGvTrjwWWp
FQG5MhCvtXr8Q4qhWRHPjHT7zac37+0ZuWzij3hw6NZulwiO5dBuxSjAa+PbZYrC
cjeHrstdzYlLEidbxM+W2dW2vsxeNVEkL91BA91RmcSZwdjXpwvPkxjBiJc8llDX
ltI9JzbC563GRWfYrZRVJdkk27ESZ3XUd8wa6+7RHnEAIyrQKoZAucYcR/PZK2tJ
KHTKiiHT9GbCSfgRlyU60o0c2IOBiAjkPuYYbO5YIDCHCE587tVISXzbAZ3NJJtT
GM7lIrlAm2gLALGljQtwkk2TgD/bQ6v7UcO4wJA0pMQc3aB5pmdzw6bMQSfxHFsp
uEHfcIDlEwVxslwUwOyxMvIJg07uNBFGXK8R+2BjQs7rkHC/FlbeyHMwdRFq590R
+9X5wlmZeJcpzDysc95yObo28DIkBo5pnQ67qs7XzoVshnRGrU8j2hOTAvHPQ5Hj
1RaTis0rQMU0Clm89bFpM6WgjJV6Nm7cZyTCF7fOWok4Yl3B2FiX0gZeSLHqKrHr
Ft96G6gcmN8/cnEwmx6E4Bbp3WMoMw0HTW29RGvWQuUUP6KJxrt1XR8Bo84pMyfY
rL36ivk3edZr7n6USXB4xYj/6jbBC0daSq8b6ky/CyjNYwgX9t3Ll8MEqTCfQu0z
BX/1fHvS3nQQBx7KVPZpKKwKIq4w5DKY27aVeuyFqOpv/I+MA+wvNV5sdpCyJycC
8vdRFKqDir82qXAEjKOEZ0KpMwcwscM8lRAEgBMZFS7B1xXELR+A4AASpIiohap4
XzFf4xuvYxovLunEwS8SChxr3P1dlJVclJjxtez3NmGmIbtWExB5Z7ibqAAiEGZa
Txsc40R/gTf8sgfRkELKHyydztxIULPZrNU2c1snJuTWShMRFUWa2k92uggr/UsQ
ZWCHAQmVUvpUhGmRoLCIJAhd0PmMwKPWD9Q0XM2gRFt4IWeQ3crQV+1IXDyQfwKp
a1uRR4uljeOszZMLah4hB59aOXne22NWk+Vcj6EywEsm483pOeE6uJVVLe2wHI9c
i3ehND5+fmV2jNVNdJ2LrSz4BYLqp5oFqv2Bkw0enZOKLLpIQpRcRSBpuH7QcMgb
zWsYHZBhYrsZ9fKtYsQCyfGhNWiutuOznZ7aCQXXFXmjYj+SJw0hC64KSXdP1jLh
6e0F+izpzPuzeDHvSFvIVgpiXJkeVebglTUyObwn7wUhUHMqrs8iYNx4U3cYQjsY
KbrzmwhREHNzLZlcT/FgQ1oltvkVHSBEjXxbBFo2AcSNCEdAyjYpHXARHWToIJtT
d/v2oyz+xNOFxPYrCh8FMebX/LCynebX8uWJDO3LtbzsHn66yRVj7nqC9O3MIXoV
c5Mm3fGyt/6CP8Wbm2syFFtBLghgPf5Kp/6fjwL2kFaKeS9iknrVtcmJ8+53b+WA
OkJ609vgNlvdy8K38SmAL87BmY1tw4L8ntj1UU7FBpXoBP2FAq07owmF9kbMZ0QZ
H1K96aqqLLKx4LscHDxvkWDlbiN0oAsQ7Rq6nOgLRzsDyyW7kpWJCWW0fApi8dZo
YQ71rtSX8yJokh5+GAKynrUKULWHuAAccmmM2JRK14SwN56WfjLSfqVnnX49nKAa
IXLlcr+XycvuCfY0Wfr4RCps3A8XiNdJxWPTm8NqHvATvZcqv+W6OoUt3QolXFAA
NWpAU0UpAVd4z3VVagE5RegvLXWacObEtksOSvSqgrn1Pt2JJoDZ++WTzqDFT/l8
UnX3XEW3CFLJINt3+CTz8UaYHQOZP7S9fpvbJK/S2vTT9KAyuucmzPQeV4WWlGxU
tWQFhup5ozAcSOLxRdGqBnlTMhMob+UHdjOzNhhM3Wrp9bhlec/YykM678LcdNjb
Te54b9lOR2wr8xliXNmo8gd69M57xKfZZzuF0ms8GRJw/8ixl5uEk3JmpvLfM/s0
fb0s1SoGoXaT3QRvUpDiwNej3Ua3dfZ9yzEaNlgAoAh+IboteOXAPRKCbIGBDcAC
ly5TKjjEju1RfHYhg9J9ta1E4A5Yg1kMFJVNm4/cvt2C/HPcD7uLGl8QYbDz4Y/y
PENsPQ4nj0j2r2NVshxHEox9up+aQxVLMhayh+BPalo6yEGlDN3kqgmHAVNukeqC
oxsgKn4PHQYZrKMj1XKx5snpxrvfNEiwK2vptaXNJz/3+1mLWGo0DNIZakB9tEI4
OxK5z2Jh1FK/Jf318agxBQXuBvD0a0DdkAULDu5f2iO/YXOgQDC81KIQEtO9Lehi
8zqhXkBf7kQGYianu5BXQ8zCYEs4X6jQqc47GnD5AkI5bbUIndcZrV3sPFmr9N8N
LubI6+jVuHPsDMoAyOr7ZVP/jvo7SO2bMYfS8wPrLw+eMSRInWem3lGhlX2zdnBE
5qzl010peTsHyfZiN7nEs1Yd5mN1/FfapzkktYSh2qLtiDUb0PQEd5z6yPLHBb6U
WmajmG2MPMamR3FixTeCyU6R7ue/JHmg4xE6riScY4rdnY5QI0TwN2UpszORdGb/
+M/zGTkQgFZCwRxxE1ZTBk8Q0mif3vQuNvBhpCBiGqxTPBi7TfFSk9g6R1cWegEe
xTQto0kregGkFE4m6Dp5jE8iPgWcaUd47VrEVMtLzzv9WbvSIWBbNo57YA6JVfM8
5FYUWEEfvZVZHOqxT4kj6KWlPQkC3BRvJs4eQ0Aenaf/B7tGTvNLZES3IyHMXIto
ueZV7d4XuETNwP5+eMAYcj8NsHLkC/gv2sEIURpNXNF13/EwshxeW6ZcMNq+Kdbc
MjeaR5bA0upWKG0x5xB30aqQE62Q+mdqdiQcvhbBQHMBmmS2nA+WjYio27mwtcLp
kzwCM4b5MYsbSYTYgDB4bwb6J9cUQiy8J6EhQyLPH1tjzJUu3vdn7aQWWHptbPAb
8/o3ami6cZRhsJYVHnPcyJVQOxfBM1TMff3SsLXxJg7KFGhfcX9pOtVXP8FsArR0
Ibk0KSxJY3UrLvSDlUJlIGVFDCP2f1sgKHvowEavcgaxNafNtPXrmIEiyQtSGrqf
VKjOrXW6zJWfzglv43Ben3JAirDXAb/pyCDTUsW1rhxB1tircyjMa1C8SgT6Zp5G
F+ZwCmac5L/iZqpfHyQHqpEzIyNzsJUYvMY2cj+ggxNrKc6a4H7F9Qb5+pKD38x9
/U8gGpySdgocLAMGNM8JtWHcF01IxxmPe3wrJHCGK4DRLXq9kBjQtjyIxpv+UNxz
8/FUHLZq9NAotjjHCYr8olB7yuhaFEVXuO0+fiYPpz/y3Xs8jsD9LEM9gRPGrlU7
dcq2nrkDqLAI0fJ+DoekvYEcJr8SP9WeZVt3PkO+l0fpQZEWJIiRnPepQfCbLKVs
XIWxJXI1Sx8ZYV7XKSbpH1ED/4LxBvXoEXlnjT49phszqdryuyBY2rJOJ3E2reQM
mVJUJ7RBACS++DlGSuBex9/ENQYzoqiNldr1n+bFbQVf3tKBg0EOo2wms1Y7TMOQ
Jynk/rxoYblETN5SXg6Nsn+RPc4ZbI+yomp83v01MoRlyshYKwHTF9Mv1U4622mG
sULju+Zi23QmtYwKMCEsn+nDGPylrooWp6Lc2DXEK+KZ5cw5578tSEEO9LLAFMkF
0db7g9l8XwwETWroHQ1hsc7hH3CCg9wmZacl3EDPgPlxq4u3JXNzq7/C57zzmPSR
wgn/3tG3QuGGHEp50Gq0cmp1ZfMaUoaKzW4/BKHQTh6G2fdR+Y+fu86zpPOsIIlF
O5GFnzRPHweIecWVVVALomuBJEukcz/U5qxEBTBLp0+grW1Z0bQXiqMh7/r7smql
jCLxnvz/1yTWpFT+9ttc70gYJnsQSLfFXGyUqPsnGIiaaVPDeIFFg+zIvYFQW7ZZ
qmn8zL5lwXpPhHd33q2B2PKbFN4Zh8vhbtAYn/4/nHEvn88Aa/Qq2HfBNlf+dAfG
CsXshFQTxxb94to5Ats2nttebDa9rTyyA8eduUhCJQ78wyXuiXbDl83iKeBMS++d
vZk1J61w4R5wKcqOVAaPK5J5fs8c1x/o2hzBA8k9nlmtpZbAypk8e+Rcw0JBD3zm
5hdkbgAiqUGVP46hsccR07kU0sjlIrnyWCjwHJZmvnjw4zIS+iDCQkiWTCCNIjvf
GTpAzndUgctfBweJxgES9M5kmDRcy0PPSX0lcV16DdbQj33+2BR8v2w1RGOIweJ9
`protect END_PROTECTED
