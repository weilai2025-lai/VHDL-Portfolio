`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZaQxI3SyOnnYHXec7i8KE/mp3D/ehbB+fBXx/TBZZLhQQm3nhXFqGZdlARUKSbZ/
it0P0y5HVzgHBFc9YW/9evQAYDaVDNBZdT6UTmy9zFM4D4nfC2oKiS0zxkcXmQ8Y
zUfo+zsBjhqEhjjuguzNt0tout9nSYmOrld7APq2KuvoOlBmhj7iZYqH0kI0kwR8
Zqp91oPf8La0sEwAfqutkjzvqHgVcrKvoizr/bZwX288bGfst8mS3ZzxmZHmvWIx
J4D0o/daPQmnOn6GsfoFB0/GelKUJEWERvQEZqOlRFbq/1wVvq3I7cykB8IXRWTq
yRvRPiJFB26HindRNPvx2pawqDVIzka0FeP1SUsBz8V2LO/2LhSm645YpBaNlPLx
+2VrR1y0coF5uZCJfTt0Yucg6Y9Dei6H0BFHFNO9zrANue6juPupKXKG+Zm3e+ZA
rqvjLWVbr5o/kUN18pOjtBbpN8o91Yxhns2b2ecIxyzU2CCWNRyzLX93adAnygJy
9oGx+mMXS/zK3SzZq6wlpaBK9JbwhJlCmmGeCXezssrI9PHYNCtXUPcIYS7tH8v0
9pocyMnWObBItCZtIxjhCp+/9L8/oe4y0DTcoJNeIlTYRX1jsXsoGJLUA88hg4/8
jU+m6dWnKXZUg2k4F+008mBcq0laWMAttU0bxH/9eMaBCmO1TDGWQKtgRcPr2mqK
F+SZtAi4LCJ6BgkhED/+hk8dLRPWFEaVhCg9mFCpVfFOCFktzPrH9Dr4DnBwchyV
GQP0mVfyYVxgllg8HyjYoIeeGSCf6LpgiR8zSOs/TQOFmS3F2MxByqXyxXvVcgOl
PDprEPLPoJABubPrMSb7jiRQK/WcC89HGU0gEsuqzFaU3hWmHnVK6+HkmBD7HDsB
u7GlftWbdJ5hAt0p6Q45qTDsWVnpz6nDiCzcLllidalAPL/ltaTsw6C1lsEvjR0S
cmPGhpB5s3D5BVHRtoTJpdro7N821xuj8y62c6sl2v/KtBc1N9L6TVHMIm2VizXH
xGO09LZy/+pb2vdbiSy1zxtlZfKvYk4DgivlmZUlki6Z51d1aePoxLLvxLJk/G1v
rnJh1Rcay/NSCOXHKIYgCHfofcr0sJBJ229pHPmbkwV7esHh9fEHbVMSh4qsc+5U
CQI7EsUc9NgWFPIXpm10OJzzICyXQ0VF/aIG0u335vF9XfLyEA0F/6e33yJbdzz2
+YAmvL0hyJQOoUyC/bl51A+rQTCBVd/DwFpbsWZrrIY5ylbFrH3XVbDpmy7AsNoP
4NAkm47bD9vQm1xVRvplhi+VUPtVKF8/9lO/c7Ek6KOEs0TC5dAypSF8KV4yGhZM
uGkcQdnELlepl7xBNoaHq6UxPoxNdzKUO8XruNx0/+6ReKbMA4YyFNLyIlTzIDcz
rB1Eu2eJ6WMmF8gFXCzzz11nrKX8SjSpH0utZQStTWsZwYPSk1ZiXPSkW0PU664T
/iLuAdn6s4JS4cU+sOOwBIfmhNzwfCVf/sQ/MsH9zm9NHwo7G66SrmpfylLZvTfs
JrUL1LSJWCAWoHFkYs+L3t9iREZw1LKhTPCq6G4FR3msoOfq4smPhb7PNiLIjW6S
6LcRWFV6VuSgCD96Qi2cLSIT74Cg23bxsnqJZnk3V4QpTnRVdFmio04k7Q0t5Q+L
mG86KgCRYTScrWxDnkTzAGhkt17FxDWts3ltea9iWBWeYyCkqCf2QM6E9NbTnu/C
CRVTdKXWWiqTNqgbAKCZbhWycXUnQRPQU7e0T/6UCAorOkiY1ynw0pU2AvWSx1wJ
woh3zOYBf3e2fswZ2htbkV0lpH4JyNldApH2W0DUcop21p3D07qlO1G+NPubo73q
RogcdmX9xyiI5U2BsczauS6BODrijwDOZ08T1rLDvWwmXhKF/gVdtlLSHBppMXRt
6DStP6SOdSRpc0RKxiFiYng3L1waRDn+1+w+c/bpWRvE9YaBnP00BLAVWhFcOFie
cit6lmEBDIlErswSSrI3gWu1Y99ybuwx4mUmSI+5bJmONbHdUwPD7v6j7cq0wlzT
wPulqL8+yuKDGg6dQ1SWRD1mGc4HFnLD/yszbDUcJmb+smaaafT1y1X/81oKQJAh
0Sry49jpJ5J6A62DLS8tUczTbY1Dl9usb/JMS+bXNK0EAcwmWXhp35ozYavwHhD5
oZ9Lo9RvQNSljV871+fpq/KT2iFzIfsD8/DBVAwphBWgdnYxreaOB9luGqjr54jx
yO3KtKEkiJjgqhHMGqsWj+ejbaQqqkEJu2anwllUZsaZrMr0rc99VAWjUlNw74Fl
pZtCPfgR/liGEL/qMtFYImJ0Owl5NzSk1fX5Dc8ETqTNVTmuhQf/Tk1Cl5WQ+nNQ
st+gHM6+RiVHgIwSkGKvlXyIaeuptLQag7FxleeAkVWBKW1DoBBj6BUEphk9m//a
ZY5PSqyWHDwhMlyqbVQn/rFhEMgT5d4DV6KU4NO9qHqirveUXTNVsx6SzAMMf1et
RVImZm0H6Oyx6OJGMg6Ma0rpIJ2QF/yYUpU0Pw9D05ILn8jOU/v66hl6Wynma5TE
e0xX+ZKz+1jHx9QpasZbKmigEj4iwTvLDq+3EFjNcV1/QsxtpuntbJUd5rJkqLXB
K4raiwwmsg88QwuTR1LAjPrIxe2FdPcc/n9YMmvC9WfHz5lQSYu92PJnVDcw+iyt
+ObYPOXG7iBjHzro/OFaoyDu9qFV1sefioB7/8Ix21ZtvPE04r7ogqlr8ti5IMxj
kDtJKQMJEBTTM4vzN3lyMtMW9GFjEvfBHgfZ4Amj89QyNBW2lL7lrJJlbZdkjHTl
1h6ajojW/tUmb49CU0Hfpf1PwM9vdCL4YzExZ8uKLmidzh013IvxIKF8SffZQAKP
t/XzfU2CZDecTKrcKXvbvAoAMXfpjDBHYjiMTBVEH7A+u7ZmPmASuz6JL64HAdOk
J68laI/IvPicw2URRrzjsk5ujvjHFgxc6apUs3vnF+MmT9pt5YBMAEP6rSaFwrfq
WjEF65Zj8duR3Pt2JfpYStavkmq993t5o5dyS43QKqxL8DofDP2mmOygohEPiwY4
iXrPguvq+chSj3ODedAJTedre8zFdiwqci3N2/hgYHZ92G/0CoUfoXwjusrT4B5I
GMYw1xh3/jhEaYuCamL2pfwN3u+UwSZlzoI6Xn0xOb2pzZRGLAoEbiCjnz6eCezn
oMulP+Ed8VyLVcQRq7H3FfUv8ECupNqRzkFAzaaB9f5b2oX25SxKUOotUsIqZVkH
cekZ1/qHDVZ6rx3sgRWQtS3Gh+/hTB8UyJ4iPEHL6L9tQvOHhqZF57wXV7hRjxZ4
8EOoHYyGTGHfeC+TXWBuIqOwXYlxVPMdW3P8M+YdFSUoQ+EGULsNHL8HR20vOUs3
P3EJx1DLTJCq/9z9KcgaUvjn+ocJOdNImGoepCuD+y215U3R4XHHTOj+b7Tqzte8
o1ORM78vgXijJTdkJ3V6ryJ7GcJF4mVtgnFkYfUqEvAb7tqJjVvLkxVj/iJIe/z9
oS92HYhSMMxUM7EpqcxfgPN9PhnrOFAxcVI9hRylNS1CFv3ADhkNumL+dYe98cWr
1/zdIFyrorAd1HBAepEiS8+6bQ8ZeSTbGlVJwqrxa3y71fR+Lq9nzcmxGZudJdGM
6IowYAgBeOluPj22bSxdAawn3DHYkSq14w2OzDiIljVDyejMChY+9d9dKwI/ID2A
gkDXT/NMeSiJ8LEW9PDhMub2XGMI8uuVOcNSyzs6pOt4TmWlC5hvW2W48IyBCuyv
J3OU+Hf0nFGMcfrnR1mXI/5qla22cUweHeefFRZYi315uV/KlHXv7GdHHfi+khev
KEa/YJPCd2fEdsbHXgLB0l/RTkpOB5DZhdOUSiJeK8Jrcb51vCFahrLsD2AR5zpd
vuilkhlIRqbhVqR0lw8f1I8mYrxOW2rUsTkAh53ASclJHHWRVdR6m2wH+1W5nfcK
dCYdT93wUdFUkwM4RVEsNNQRaCVMrgc0AxxDb3k9WiHr5W19vv6zopJDD+5Z99lM
WkEjNuudkmU2ZRE/kHebXp5RVwPksogPoJ5UKk1C3BeFMib35NbArw3z2rt2c1E+
HeKZjhg9mRIbgrgvVOfxsndpJb6qWP4yphlWaJJCw1VBQoG6xzRGZSHl5lXtPzM9
Ig0jrdblz7YmKxYxBD1HQJGVmdLm79stV3xwI+ESjqGEsDi/2na60RFg1M9e8MEk
QJQPnWY/jywFo8B7lNpik8SlZzZ9YF5GH8/VfniiJkIymtUENo3AOvzt6FNbFE1r
ljYVyJs14xbPiiE+ZVqNMEEKseyYMxu26tAjMdCni7JSfu86bwUFib+Yvtw70kew
d24I2uQioDFUZAELc2Bf+4kk1p4r3zNQeV7Kq+1vZWAjThCFJwoj4Ilj7FA8D8wM
5f/vNyJ9UP865j5XmUlzYe4ratyNFn9BcEOGFBYitdb9z5S5x3NbahFtg5dFuCiq
98nyRP83GXyH9jPuIMwCchDrsfmnYeCX/gdNJ5LVu5sc0aSHB6SkugjbcWIUXgD0
6kENtw9s/3sXEgZ5b5yVzD8Qs9wivMinAlF66PlPtY/IRp18a4lMdcI0d8EGTwgo
StydPMRMlCXoLYGJJqsiasv/GFeXEoNpiX5GH3BYDm12ppfW671Yh59a2oh0jBox
LWliji60BcvePp1h2rJHcDL0KWPhdCim5nP3pyEC+gmzmx9m8DUeQwXcO9gEdX+3
XnYLD9v3SUxH+UTwalmOludICqMN2JCEHLGVICwki/eZRuv1HJaxflBY4HmH6tUh
CLYW0VceBH9BMTSUiZMbD0GjT4IDaHt8HpraDTyR7XCqXA7A9yOO36SODfdpqkX8
lZzv8xF+kPXGPScxdjnMgIMAPEDzCHzjI4zsOsZkRvT8xpz3KAW10eaqD6m+QQMo
K1wUu6aFNGWocCPsEJ/u8TQTdMunnyRDjN1FC8jxvMkJKxgxEkCGzLnA/POQD0gs
BT+gv1qKl9jFXb8nLO4ugz/l1ROgURQwO8/PBw/U6lSYru0REDTtHLMa9RlzBw3X
J6YjyytmWuwXhvO2EbHK4mHIY4It+5Bq69PScgy4sQJfbMQdekF8uzVFOtP256nr
nTge/UyYZFOEmBpHTqhL7hjRPicpx9Xyp8BvQp+YrPoGlAzNNR/aAoBhN03eFrZS
GmQ+uXurYFqZ8k+anV6Y2FazIgwCXFNv5NnbCYa2+iYtkBm9EV4pdzF793thvmN0
akmK7nKokLxPqWrZnxHdpWJAXQyHNmdbd7NA5GkYwEqeYFU/GOQMWGIIG5y6pV0m
LPYWtB3e+17BWdUetF/MF6UBXYJFU3VycoXwzNgUXwCQ0IjfP522+qDjGg8VuPrv
5clYJdmPxjIxudXS6PaEXJ6nBgI/dx6KtIZ9XhACTaq8mmdx3lKAEia0w1iOrWm2
++ndkQqcIWOfqHqMR4Olfn4AKYDBmqCzYkL3nzZeG/bX3Gerrxb52ifEhJIw99F3
LYhBGdsXzsEeR1djq4YwbZ3EAVuDQluMIH7pmCW/k+43ChYJuYLDEOj+2VoSqg3N
I8hVVaRXysWsxsFnpdtP+IDJBRDSfFA/H8GnbNPSjtttlXAeHJenEr4CQdAe0dnH
Sr9csy9/K/wxvWerhExEE+HZTAfDGaOQNWUPIv7yuwSg5ztmSg4QswkpZ36vuIeR
UqCGRP1f7hCORrSYRbs3fqhnqIok3arcO2LdLG671FouG2vWBvHbbrKh29sQPvGp
KEjFN7KoxzTtE65BctV9eoPczsZL066RPIMdNlW10ZBUAABjLh3ZiZo79cJVixio
tqWOvXdleq5hBu6zz0XumvmxqabRBqTMCjS/s2GyaZttlphuq0gomIclvVPYXi0i
3PT8R2Y+44LBOFtNAXIfsNW+mOmGwo9ecxLHKpAIpd6kNGlBlPdxvLoapBxqkDWH
CG93udqUduQv8denq0Qe6rM1wfsCPT9Mq1x/2aRKSodf0ump44QkCUiJijUljt/h
MkElSNq64fue5/jUag/NdFQfnQ89awK5Sx8VSF1ARwOL5E+Xbz+Sv+/cjbBDhzMT
AkwuYaCGlIe7pD6BuV1eoMzn8VV6evXvKqZHswnvfphLEE34Um/A2Oq5Cf2+zMb2
gdFi26LNE85eO7LRCoLEM/aGmg1tkvvBbjwcWMqmOzIypuLt+Z8fv6lEUVballQb
2I35JkH9lJ5LAqOD57KnUc0tong8WaSPjxM691fzNkesZ3r0Nmiz3TJL6wl4pqx1
XrFj5s92Mi3UJsdAcR3lsyHDJVFd+BF1N98nxuGFN/ERnD6jhj/+wXY40q5WkPKC
D26N7JtB5vbTBfLn4FJZhKpLTImx03ffoXtJ6gsUHlK/8SKsIupvNpESvHVu31bZ
rOgouXqdGyzdW1sWiVF39FGi9QNCds6KVZEcUPu9WE6E41pDTeIAcLOQBI/nh+aJ
rqNhJ1zk8NlGQaxW5AVf+r9Py4Tpze12UYOBMY6roO0xd3X0LmYqTfyFym0BNbbm
scpNqUTV6Jgf1IjpSh4LhoVdPBhws2aI2d2SUKWUDecCtT8yFm3CzWTT876PTNcD
envm6aa699jGss9PeGIQvk/FVfz18oPk663Vke8V3mE7TT8E86QWNBoJxUvG6wbC
46vDIqZbk1UD09v+nSTdoHsjS1PIZpGs/fQRAodrTaIl+s86zvYewdsYOtwS1cEE
5m5AyRl6ynPS5YwUK/S5psZGoVpSW5aeeXBsas6B1zxf2ZLRO4pY2hHoJk3L11j1
hjJnAe2ScnzDxUjrH7jiJpyJ71AqSIadvTcLz8xnMG7TnWTYM6i6i3olL4S/xxsK
Msb7eP+tmeOw4LWM6rsubQhAp6nNtcDmCtgGJ7KLAJCGF3mQwmmAr/fA2L5RDDGs
UbZLTQWjHQN5EDZXxJR9PvONE5xNZENMuz5qEMAlPr4Lr36MQjWIqJ0CDHFBVv2J
+3Xoclv4S0eiggvcWgBA/ZU/S1OTdMIR+41zQhRDHKSM288/Vc0/ekGRG6HZpeAl
zHF0OBupNVeb+dh2y0MC3iL0ge/veduhkVc0vIMb4FKnqXi2WCt07AMaABVG3mYw
0kHeMWIm+gnKZOCbCbs/sKxI+rOn8NWBO25FyWojvmMF7WDDmJPajIfA/thpheFz
Rf1JWQ+orRI5/jJ1eS1KjT2ywLqXOwyIniNhzNIV4mO13m8fybrAha0lk/CYHFEG
o9DGrf3Fnn3oqVool6ROhRQhsq2my51CSQpJUR4oCrHMDAvMETFtovs+izrWXYn6
Y0Pf8mdM97MkGqKL1d2O+VD3n7JhzJP9nISJHrQPpWI3eAxoqKyLIytpjsobqNit
D5b9IqT9V/BO9H1iFsmIt6zfDeA7mm/7OOxRuG2FvcRFAfqwQOqRrHGhfPrlI/zS
nUOj+UuTShiRjOLUUF+0nhg9LwW1CDy6qxdx9HSMkdPNdydWgqUBulgaROZwEjft
Ybgxt2H9sPfyctBNMszFMqfCSTy5ssb4xqqnHYRgwLzEVkbpAVLZ2WaAS1KVnHHI
75SrbmkL7UmrPhZ+wx/vNA8lDj9gpWLqaG2eCCvhjeOf9FDISzMNVQ/UvvqH2cRo
rLWdFohL5P1Jzc4BefeQ8ESuysNjx02YPx7ScSo4L9etdvggPJn8hjipp0c3rJLA
KOwTTS8zFJ0oFVBaXiihGMKEQwobVG6W8uWuIEdEd4UnkexuvG7QcPF8bT5Ljldi
5dPs7bEitxgePLzsSFL6nuqCqlgQQRLzQP0nwsS5DgvZd+8Tw58fERQU7wWdQyjy
FycLYLKkFIbYQU633kzmDzZ4srFJUcm6frt4FXtbDJ5tbyT2Qzc1JvmXXCqSsvws
0MH0e1ztWCQsrxucvjPsJC/iB00lkchA2Dl5xhzkxA2PracXxxy9ETaTYeE6d6wQ
LqRbbjYiEs24mrRPEKcQVeH43zYq3BG4ucpFRtckS6MBCqkU3aMT252h4HFaTNEM
UVFrGEvJ+me0erGS2Q7DMgHtB+XoNz4HbqCYz73EoIRDQ9MLnoKnWWK698ElntrC
Fezmy9Le/JufJ0ywodcGURdcydw2/WK9jQQraVW8qE7s0uFlDNVWvOY2YaA46lHd
L4paAciCDLEaHQqeXRpuYAsqjapbCNvyJE/GUoucYUdCUa30A4lrV+1A3MPY9Dfu
lf8VLQQ+qRGaQhoPHAKO4VpivSy4G/5QU7PZvB4qAom6s9YuO4WHXQUKb6wOeQmF
qV9u1Wp+4r4GRB64nJ2gbmhm3eM8QHOM5g65WtZAL62NNanRYRZjtgL7uN8oDMGH
m02kOerS330fXQBPKM49Z3Jlg7Y299mSyLZbKFuM6gEeTuAo/QbDN9UoSszFfInB
gQ5ug2N3T5AMcDLqjH5Z0oHHqMRAkl1QaM95S2zDsAiAnVl28+kwVWIf2CGz8oVG
KfM313RlLaZy4o8cb2ibpECVEMrnGIHLWAwkroUV07UY9EI+maaruGy3/3C4/pV6
AqYB42qEUCPOkL4MLzaj8TFuzqv3vJGKAI6HSHTTgZfpotun2RkWTw/E7TPNMn2X
cnbvUMcJDDjiGn0X2lAMRw1qmWUWiwX3x/fqD87d7U96bHqFafFrNTVDeiuuC0ba
GY7pjkkSWc7VnuMQ4FPB9u4jVgIB8wZNrX9o8i8ls37WQpPKYXXvI4qnKQIjJuVp
2vbJia7ZVlogWUaqFE2rPsFjaZ5RUrqo/FTjwhkg3dPyNUVDXicDHgqDLdLKkM4R
kVZZoVm+DspVbLqM9UQsC8A51ggFWgqkRVokCpiubCEEEEGzUT5ShfZkbpGCH+Rz
kGTBzmRsmgwQCW2yTuiI55V+waBbAxe4zpSEI/hRHvzwyHxmggUKBFFjuFFXeVfC
VFxuba2XDKkSTI/jOWFrCmLvkc5rK/I7oHfVeXRhxSeWIiV8q79MK84aymQXESxr
qlfXjdc1K8gJbQDlIqNHWl8Ba/BNroyZtuz5cYGo8ldw00L1eK2VAQyPS4f3/v38
YPfcg+H3Qa0op7D9T37CtHHvhyceusWg4TidNVOsbIlkT6pGKV3aqKjjiULOM4oB
Z6DleLJNo5efDL8S4TE/OqWpp+7PutJaU2gGdPgrn7XhSea4jqKIG4vqCxe5W7VE
3s0dd5G4/rHLWbMfayUQ0p4JFspxjVNuC7Czq6O3Qv4vLwXZMEwqyqRlfth2HP6r
pOsY6ooM593JOhp/5aa6d8N5g18TDCbbsm1j2s7Y3kYIEDqmdaXDQDn6CtqVF51h
okTKvHqPUsaYju7y6CVI6YNcl9oCYJztz5b1Zw+E2Yi1laMuTa+ep9ouE5Ebhx62
FXWzo5tRqxXZznY4EbrA/FB3koRhnIAnTyfNB+fDgSTBKJEfTfRfgDt0xPz/R9Sr
yaZ1Q3IkWh1TvRBfXcXq33fG3XpN3xuehBob+k0GInOlFakr/kCo2hEbDpLU5ysm
+27eP5a4mbbe6iLoPRVHQhzruzbtAJDyeEwQv8CoaFXqzfW2td4y193SRmOfSX6S
fjloQkQKnxIV7emzMjIaw8n+U9KYXhWiOp0ZxzBHo7mltA7+LMMPWPbkZIKIRma3
Xw+Vys+6N3jlOm7LhK3XnbClFTMJpcF0obustcA14GvNltmeddUv/jwEH0SVxfFW
2Ww4r+TpQlho8qAySA+5WfyDbEsCj7BNmZNfaU7dJfpnFBMrwuebNqBP4AGBBga4
DNUIwItjCQ1lat3e4EBuVDuDwCksinS8KeZsd71iM87xIrmvdRlFq0mHKU6bGbGZ
hWAGS/8H0A/cNBDUpDTc0i5EH/peJ7c1tpN2KlI6UkaJDmI/grpo1bfXB+I20NSz
qx/+xRShhT/P1wvqfhHLMyUpdmDI2kKBV3ZpR1jkgkjfQHdUkWo9HWCfKOICt4nf
b2Jip6J4cnamY7F/y4NghRQwSALDhjaQxMxOOweo8fORqO33Ik5loINiR/uk9auf
DManc9gI+ISy8FdCD8b6I80TwYc/N37N1u5X6W3ykCXpZM3CRGQwbpVOzKui+trz
fFEy6XlSTttAMUajD/498/3Qpcr9IdAnSg03y5ZAB4cqk4B1dkTo5qMoBsOZiIJK
b3BLQXk5Iau7VevKmsIASnUPLnJg7Y7tR5+7cH4wEZqx15wUsU2h3OQipNqgXpaj
U5ptQHrITzDkm7++xhSVcyS+mGxTYliQSFK+xobh8uwkeKQjTVJZzqJbVUhj9p1x
H6QRfvun/sFhrN48zH87MCphzqrdtNnoRDOhs+LbHT1dcc9E2gJyDXX3HLp01HLn
QpjbbdUPHjdIfvGtaccFGqyfPE8wJcRRrndFPDtxiQOeADYVuMxd1GtdRgZyUYF5
g3PA8+VErmUYRZDkKErbOwdcbPDm2e3zc722NkBewnoNw9yYACcSa9taPUgG1Hp1
GwZ9YT/DySynEurjqF1desCqTlLPXl05ZjBPsYwNAhmcMHJ/Of5rfd2dt7mdZoBR
+IOqh4DuPHMRQiXN4xf34o+GlpWIljZbsoIFSRC3BmDYnRbt6HbK+TzJu7JMCECj
d5QuYfodq0AwPgqBrpfQVITu5JEc1ANDGEJBFaKjwYv/lcMHSTBXfUtaLu7SgAGw
BufsnwzEEwmDmt0OWngLfY20tZ+aPmTVHvB7iNBAEQj2ni1CWF9TjUOpltglRTot
EYzYUDxw9rOE+B/yBdzAB1AUC86rZ6EbS8RNnifIbZbfWftRlHQcWUEAvb4mY5Fy
/EkqI19F8w9X6NwRxhPf9fM8p4UHmXNhRJGEvZ/+KSte8MRMe4IZJOH5TYzYt3zu
C9LEgkI5Bq4GBdpVvElJxQEZ9Z9ZCjJUBoVD7GpOo0yucJgdp9dkyogLVqG59KeH
Mru0Pd4yYMYKu+wHAXCMYaoYQu7amJ2Vde467jX0YdsgcSzJpOfGA5Gz52vtd4up
DHPjyWl6aQ1M9qjuMpYf1zqtfrqHz9uJahevo89GA4QAibF5XrpLlr1YtanXgV5I
qOczIrU9WMrOH7WAI8asbxNPrma/Ujn7YQZLCUhdNdC7Hi8t1DdpRwlZbB4+N8+S
sYgmHd0oSjLE95ZAa0NmZCdcNqfTxO3d/9IE7Q/T7fLSEKAatvoYIy7vvv4d9/K0
VcnhP0n6zttaCDI+jmeyHd/DgRU+yH8+DD2QYEzu8wEtmzWnGgFpmFGnAOlVsRvS
aRqNji35S9Z7K9btUnc7Yz01/X9YrJ6aEY96/YrTYYF/I0+CYYWsvRih5Gkb+QpH
edxXhm5jdJZ0OntewaDX9jluDbeegI9TO7imRYngvTHvOumHbPeO432Z4EqOWZUn
I5/g/Japzru8yXrlq9ab9ELJHLYwCovAe5HXvexdcOFiak4WDuafqXf95I+jNsUR
hMJ+cjm2RcONtV1CkBbUb7dLmCVwYhrIjw9SvRVUG8gr6JLG8BxjiUFyGxQNSIzP
5mQ0k47Vc0AMZ/yIX+KXGTezrw59yDLpBD5QCull35f1C7f6oj1s1hKWFLzJrhgA
cMWgkahpKat1dA8IHFqOh0pRi5dZiizcS2buYHvmlyBRu41n0rbTVYskxPWH2tpq
wYsO+inRvgupuDpwAyMEI8RH5IHIKG84onApLEeAAQTc4Q8yakxZm6r1onShL4+f
gGIRLxy1G9DzNzyaqzvT4VQ3flt1m6LWabKztpaa9iV5UWIvUunCNzrpL6Zd0yet
kRZQTLVnY67IDzHFWAcRLCtXyC2c+cP4TDL/uHp+05XitvCEgKXI4d5FSpKNcMhE
GKSJHonAfHxyb2CPASwlX/v2A1ZDJ8mhLt095ffAGxuoyaYcvMwj3O1zLwamSRdl
e85wVGzNkoeH0wg6/brpPd6k1QWISeI8hKSQv+zRKnCNJQfSbc7v9vR8K/7qjBtT
mkA0H3QAKLFWATldC2FszRmW2peNYTcTvzhF9AIfJ1b87QC0TNw1vSm5JZHFK1Ce
Z6a0lC0bY4aQEAjt7wTKl3eTaYzYYRlRhAzG/JSFIX4WtfH69+2E1l78HJ7VxAfJ
VfUtk8F7co7m7OCHX86SgSAMF/ueEoh+bL6g+MtgYpA2nFq8zCeNe5ZTwyitH09B
fe/oaCHrpH+XWTAP4W63DIi/AV0m+pdwrnZXUJCQuUT+G0m4UVHD3xjpsmOUkce8
4Mc33QKydApHqvgBjwwWXGAM3MX2fRuHQjRIX0hPKIh7l0/GOKVBO5rYScNBQa6X
YAGlTCRBGqeRj7+mouxO27spDa3Dw6Y4D5e9KPVeGrzupEojTYEx3ph0tx9GlPva
D4vSTn9ey59vpaYyYGxStcTMNrXfoYy49P8xOkUgcMJGl02WBs46jv4di8rVa66e
QRhhVmAIZiteYmwsudUEjeNtS7wgzx35PLzgTHPpZJ51pocBzSQ2KcjgC15B5hR1
Gew6jqiqknoQwy9EIQ5Zz9KUCub5b+nzEXwhGhDDR1C4S/zFXUG6WP/cK4M9VFbd
SMTZ4o/GXm0+RfLMmqn30hwYy4RDdIXAATGY8Zw9KJjQLbzqN4B/J/jhkWenbIGz
J0JTF1nrw6F09bdkfqCwgVu/OHR5113LbByxiRw8nLKtC/3On+U8iylZV753mZGW
izhB9w7aQO7lVkcP9Vi4l1HIX0cvNW5VOPjrEecOiK25H/cLg4wJHbkfggifIPq+
QC8BfZe3zA4zEsIZ2cbDG/Q9hnVYZaV/a23v9UP8Lo9t/1u6SOnJfwK2jGiF/dU7
RwKe30j7QQGDILelQmKmk6nsNUOX58rSKk476HY4+A+p5/NnpQG/XpJnsu0VlrxJ
EO/OA0l1H7PfYFE7OUgcJ3qFTvy7qxU7h/1KLmLcZFAz90JrgBc5If8vp1K+RQin
lkf0wLuYYokbr5xkDs3nxIXJofN9G/X5fwZ0DdTXcjla0RuESAQCI8XBu8T5Ldl1
ZTk+132GqrBj88kQeSFZoU5NIIPVh4/6UFBjM6U6A91jDfHeHkLdmB2y31yTdpdX
8irMOV1f0Zi25CHa8nWrM54xYlkN5H8e7j7GIl3FE2+d0Hbw7cScX4JcgmryIkvF
PgQLoUwrFBOcUFijHFoQN9k8l2a40Fq3FxTNuuCZoFtNPc/t7ibnJ3+0+A7R4Nu8
1ajwLJZji2RWlJz1qtPPXT1JbWGGsJ/CFfMzx4Gr3DT6lduQchqMss8p40IDJ+Nq
3ELeTXAmZ8UB2xVylO+JAQ+Co3go9AytnqCrm6uCUm63OVT4B17+P/CJJKtMHoYm
`protect END_PROTECTED
