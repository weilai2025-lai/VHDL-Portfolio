`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
no3/0F0k9hUEQaku6feL0f0/lMRXH8qzIrVKBeoWEtsH1RMjwQdxfMJcpZa/uTtb
HcdgNIIUOJmSeutqqVBFOM0HjD/kfqo0N0nDFVYl182qjpL3XGLVgf2g0zwqao0J
m1f2YB4ugq13jCQgJ2J2oE+S/EqaVdb+TkMVvnA9WUEo3kCT5l9LydAGeqMWe7lf
YNuUxpYzEgq8nPP+f6MK1PC8PigAvBDYr1gt0atCjwrejwhqRnVom6QQMVj/iqcW
Zzg/t92X0geKWz8caIBe1mHsrJ44OpQW3Oak32727ky0raPNpsPGnIVfGCyJB4QI
vaKKFgPtyV9cNJLar2W6bhJR0JosFx8RwmptJ8RcfcGvOT6eZy3Kb6pD9U1HxI0z
//8lguvpkgotBSi+Z9K0fEjgDz/eBfTRf7/UCcTLHr58Y3nk3PGsDKD1876kfkoj
vC0t4qhCQmk/QEfXSzUqFGFCmi6/QvvhWk0mme78DaWk8BLi+jPwLE+D21WzIB5E
m8MxxWraAjSgKiUbMpG1r0xV6UBxaLmfLmWewQKBCwprF6KFflRkwU+Yry6Kv9Aj
UkAPmHrvV2qkhanLQuD15cDZQOcyKkVQwsVqurc5koTSVapiwYYKfkmLLfMGm2yJ
DmDniobDtmRfejCHelajI6IEnHpiie2/QmYJTeXvriG9ueGqXkyug8tdvMVFCVIJ
QJqgomhoPhypg8JLweZ6k/DWwc3ApsSlp/n7x7xR3Hy4b+H08lzot4PQA5F4Ml3D
0axIZatP/3XFBVO2ym6Go6I1UzRAlcwCDyTyT/5iaJidJLZxI0ptQhJs6lv3vNOO
vKv5LnVHJhl9iu5DsMSHOjC+QNdhfM/YaA0Vu/+8j9Y5qjj9ZMSf68LVt15DoTPF
bkp0gy3Q/ayiUdxTya+2NO2ZKKA02y65XpAAO+HXDtG87c9ehy0mALRXlg02bDKg
YXt2yopyGjedAvpurCqWCAYR4Gx9sghkUBBjLd3KlKv5KlODA1r9EcAagBfKZtFA
0Kk2FTH2aaPzMyorObhHUuJTD+wtYQW6HzLGWP5LBraz7gORngWKnhXFesvYzcOl
zeQoD+ZpYJpIGUPmm8xhwmmVwWDt4jLIbDf3Fk7x8dfSmCjTZ+dU/WGx96M/0uxl
/BNMqrYmHViAntsW3kyg9uVhbt7FRsIUIDaJMrISr12Okr0E+EmrTLSeTLJLBKs8
TTc7hVj2e0Wau/vCFVCSkcWJPU6alC7Bt04vwU4bhitd/JAsbTxx6954wlygJMK2
/US5llSWrSkL3rdYUT8xChQHViO+y2NDJmKf6vYC6JhtN7j+izGToFZHRLCiILxc
qSGJE1pD+60aZ+wKIftBoou1u2Udoe153O11MiTlkVXlTFTAJioVukeyLx2T4Jp3
SlF9gbuADCzPftE6fEVBJnUALtnOQ/c+X4AQWsYGccFxoFpid/P7w/WwOg8FdVod
8NbmR7Br7UpJDsFiDzN1XnJIVCAHp5u56WPY7qL4RjkxLUEs7fYwroayH2Exv9YW
aiODlLjducP4c8YxwqRA38vc4CJEBVrMEyznoh49xtUCT5DVd3sTuQYRUZgxVLKg
R+Jk/zwBLaRM9V+7ABqcvV/GJWHoBkOowH1FJ+x87sbIRa58tVqShKT2NPzj1ob3
NKd9QBX3Pp/nEk1kQtg9J130RX44xUw32gbF0HV/nG6/jmi5MjeNXZLgVkDIfy6m
6BIy1r6ATHBFBih66xb8EJO5lLr3ECMuJlKTgJOg5RZbFF9vr8vheOJwTk0rImr1
xHO2WHw1JEJEGgRDSLVeNzDPod2I3eVttffzHKnxcKT8KoUaZB8QbqvvLRFq84Iv
E70a8joTQZHechj+Yt/cw1sKuxljyuLXbQ9IbwYhd17zWOo3JpqS2znhE5MOrQ5J
8ONVma5z8I0GgykdxWohoT+p+M47T7CooMl5gHW0RPc4OjiGMAhkFaMq3Thg7vyk
QZIekiVhoCi3UwfwfGTUmV2HQC9xmZw3B6ZHL8RSAp49gFNPmpZt4mDWy2QUxal1
u5GAdXAhwtwiDq4o43BQi2VFwJCtPNZEkKAj/kLP0GYsyZLdYGZHAHTyr6r1HLR8
k0w0RTd9rrZIaleasSdyM8++AmyuQ5CejgNF8CNMI4bcFRcb2BxRfx5DmLEzQiX/
bcojjYc+pWd70wRC0VhQaji9OAnLPz16pe9LiFA7MgJareLzL/CPZ7qi5L7LjSwU
ZMljeH4IXCyFvpufP9QcBLoQmfeMTn9+WXBMxiDqCzlLF/M+FuBKpRg44uUoKgn3
ufem+KI83xZ4KSrcYmQ+syLFqrPWSOvvCV3dlo3GgWRDCg0QBojOYA3i6vwKJjtP
p+oE6KuIQw2+bAZCR28jPawhlqUyn59xC6HYPkYbe8z1IhCFbTQSacBoSGfJMmo9
1JxkzRHIi7jOSmnI9H8x+XD1OGRmHka3aVbnbBqfDVVC09gAsvlnLdsY5YgYQXcd
VXhMFzFVeew8C4YvOCwGOQ==
`protect END_PROTECTED
