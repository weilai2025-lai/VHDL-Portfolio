`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yEirYoNnt8JuAFpR1nRf4A9+aZZvSvEDkiRJsCqcOO6faTMrnpxuJg+rWuKnyo6
WkkO2dZRu/wMsI99fAczGHNUSPLSzcn3rsDzovfGymUlcSoegxx6YZpaau7H49oM
afMCbcNx7qI0tgIE4v2aKgmNm4UH/VAvXN+mqnWhV0w2Xa07FLNXYVZD38PmNPq8
M4g59aNo2WMhNEoSaWy1hpGWIINm7csB98sWRw/CsVEhMAw1OXuhMy2BuM/MSysW
Ug0yev3zdnhzXTXaXinLV9voAA/qFyNB6XdyJIBro/LrusWpFdbufYFtAmKhtoKK
hWWPRSTxB/MriUsMjk4/QRVUyJVSUV8RE7gFyCZxI5X7ZTAjgtSn0mlA/Ri+4QPz
QHEZDRNO5OlaYmSp7l++RmS6mfe8MB+QCz5znbBIRNHfXfA8sC5uGHADK9upy8DP
UWcByTrpWh9fzHyGwz+IBE9PNZIxcKkvAeAVYxuM9H+jqPQHPXo8nVNqs4Q233bE
4qYtyRqi0lKyxw6RraoHa4UB7iY5AVVaNhSR6zcxsxI=
`protect END_PROTECTED
