`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ifac2aQ8UBUyhEpEIJ1vVawEglnruKkORxY2+sIlliwsI8U+D8ZGhOfmB0dPDqGF
VCwOkSP2KnlG+ffIcrPKzx5Orispg5yDjx9lpdZ5qEHQjxlXsg8uafI4AhCnozYt
NpJXOumE/SAUn0YP2FppasRfDKidig+jxaBS86Cjx6XtO97LpddOhkYxfCoNHHSC
RW+kBpTIBc2AoyVxNzxuo2VU48thLk5O4w0btOD/pjcbCXLgUplx/LnMAm5GOhup
Kx/U0Llrni+TRXgfM4nEBLbu/lI70N6TLUHx0UpYbUgMfyG7mvD8SUjv3QN1I0dm
wEZB8tc2WV8581XlJeRjLc2+Yp4B+f2t1md/hiNoxD5l7u/5MHU7umi2AS2wzZlE
bPbstTd8NtLaTKS/1jiBiSO7YuY9pEc2tp6SdJ3QT1Eg6TmNb3Vu608L9huKxboR
Z9Ir+RZ9zoxT7K/4ongDnswBZAlKFIlAMQl5CadxLVGUXWSlDWE6KKPfbcxYcVm6
D6jAHOToTh8F/zgElQueqh4VjdZpmvGkxlLoQ7L5N6cmJT6vS3z5QWrPMHD83FvV
PS6TSLusJFIr/uaL3SnOaLt1eOcQ31N8Wuvm0Ve1N/dEPHGcKJ460xkDAqEFBz+/
jKJBsXhbYC34NiBVS2czu4ZP52vRjHDhptqptj7EmxJL92BKN69WB17xMec2Kt25
Ge8ZOm8esyXaoMep1SRuFQ7rqYSxuS3kdrRlHQ5tjelRgOQS0J5EbXCVYCpq6UGe
dycUGUum/GlBpgeCkXrN08qe9Tbh22Zhf2UoLU8wxrB11qHMdLAL8jzHygQEiMAB
5Rv9hu27K3G85qVw8c7aLrTOOgf4+lwI8FfpGm4280A3m6yt5pmFu0wdp/SC4v6f
OFuNGpooGnN1n60qBm874AR1JawghCEIKPaMuIYH4yJJZCl+dTswKhVHIvTbf7ik
bb6zYCwOg3f4La/oEZL12SpgAXFcXTNxBGAQIKS7X8qHfZS+TNdFsdPe4GZp6ts0
T141z8p90jHg4fp1Js0C4UnWZFtS1JBcZ9OCid7f7ZT+/dIsAnMnvfiUJAp23PO3
XB094V4laZLDsEeCS/JfNssKndXzJe7qofXWk6GFox9jamyNAVGzba8UumPx0Jw5
qmNIaj2dq3BepcCygiJmiWco4z4V6wTV4q1Wbl/K9Z3LMCE0QUrgJalcCz4Vrz2Y
vr3mZfsnjedv18d2aJPxH+n3BPYDD4GndmsZ1nLagapsXCwExIVVbhYdjdeOc3s4
DiuCdvuDthVDn8FhZdvO8Q7C5NavsxpjDl7K4GSdtYwt7wdX8SXdH4lSl5livhqV
E++LRuKX3ZBw0hmqfrLvBS0l6X09+aBc5hfEl1AwwxjPvyD9+rE7Ex0BuTz8+/sZ
dko6+uKmAnlVPDIjx2WwtpsCenWptVRRTwOoQBSoc/iCf897HbbtKcfCoUq+yiTS
lpcHgyO8qX3SSvs5fCG7eJFFOks8ZflV2kNoefj+8os0kUiGR40ciW9w8JpHleYI
WxMqH6ykjjHrzB9xrEBsc1IeCTcg7+sKa3Bc1cs24qQ=
`protect END_PROTECTED
