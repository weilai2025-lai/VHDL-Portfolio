`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TqOdIxQa2DUhwSmWWqQaLgmtdryTe0Pkmiie6iBBXNOXMGkkxZi4EPZXUypvpRWE
0nbX+/QYm8JuvTNMEKGov4DiVXY82l6v7V+iWwhMCRY9jHrK8UMOi3wlIjfkwBLm
jOODAmIdQR3Bk3wIT4IPjYzWchUDub88WXNRaf2b7uvJXQjoN7AmOLMhaf5By8XS
XN7w+USaL1gQXrhnXLC0V5FRzyo8X63rlr+XHJN0tfgH8gRc9u+RVlBvnFsGRSf/
6Wj3jmQ768BhXfgX5q68LvgAVrdt2JrkxKZjAGmgTifp5jgaZACQRvB8BsgOTe1u
ToRsYrebRgooh/jqkF8q/Lx2cgpUEYLwLRK50PXwl980yJQJQr5AH7cknhYSHelx
/Y6pMz9tvWFUK/VTDQy7ulja8ScGKzc9HGIfcD7Y7sHbPZSYT3BsnmL14Bsdc66M
C7lXdVKnpWz3D3/draKdOoRp+HyqQiSKksOT7p7l/ElSXsySMNKEgff7ePSi4JeA
mf9iah7AgL1fTR5/276Hn9/cjmZfhcYPdjKd+5R3086nPgVIU96ZYpvqEBCthaTL
OuJv+AbaSKPunP43Ra+ct/hEbJKwUEgjhQC9vn8uJS2CLR5uwCUFQoYcgHNuqOAM
sW5kQpicdJQdhtwj+8zvU7h9fvFVqTRGyZQCyEEmEqE666mr1+Bvx8vGLp9UQx2t
1AH+wRu3iJdsGHC80yziJv8bGX3ITE7kXRFINUnyQLqEkJw4IMk8nFmgiQBXcfqD
ARlyR2zhefXez6xv6O6uvBixINT7ZBYpNK6leEITVgRgsfIVliPJovHsMVLlD7+I
`protect END_PROTECTED
