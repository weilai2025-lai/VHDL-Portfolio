library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity mac_int8_pipeline1 is
	generic(acc_width : integer:=32;
			  sat_en : boolean:=true );
	port(clk, rst_n, en, clr :in std_logic;
		  a, b :in std_logic_vector(7 downto 0);
		  acc_in :in std_logic_vector(acc_width-1 downto 0);
		  acc_out :out std_logic_vector(acc_width-1 downto 0));
end entity mac_int8_pipeline1;

architecture rtl_pipe of mac_int8_pipeline1 is
	signal mult16 :signed(15 downto 0);
	signal mult_ext :signed(acc_width-1 downto 0);
	signal sum :signed(acc_width-1 downto 0);
	signal wide_sum :signed(acc_width downto 0);
	signal acc_in_r :signed(acc_width-1 downto 0);
	signal acc_out_s :signed(acc_width-1 downto 0);
	signal en_r :std_logic;
	
	
	function sat(x :signed(acc_width-1 downto 0); wide_x :signed(acc_width downto 0))
	return signed is
	variable y :signed(acc_width-1 downto 0);
	begin
	if not sat_en then
	return x;
	else
		if wide_x(acc_width) /= wide_x(acc_width-1) then
			if wide_x(acc_width) = '0' then
			y := (acc_width-1 => '0', others => '1');
			else
			y := (acc_width-1 => '1', others => '0');		
			end if;
			return y;
		else
		return x;
		end if;
	end if;
	end function;
	
begin
--stage 0 only do multiply and add_in
process(clk, rst_n)
begin
	if rst_n = '0' then
	mult16 <= (others => '0');
	acc_in_r <= (others => '0');
	en_r <= '0';
	else
		if rising_edge(clk) then
			if clr = '1' then
			mult16 <= (others => '0');
			acc_in_r <= (others => '0');
			en_r <= '0';
			else
				if en = '1' then
				mult16 <= signed(a) * signed(b);
				acc_in_r <= signed(acc_in);
				en_r <= '1';
				else
				en_r <= '0';
				end if;
			end if;
		end if;
	end if;
end process;

mult_ext <= resize(mult16, acc_width);
sum <= acc_in_r + mult_ext;
wide_sum <= resize(acc_in_r, acc_width+1) + resize(mult16, acc_width+1);

 process(clk, rst_n)
 variable next_acc : signed(acc_width-1 downto 0);
  begin
    if rst_n = '0' then
      acc_out_s <= (others => '0');
    elsif rising_edge(clk) then
      if clr = '1' then
        acc_out_s <= (others => '0');
      elsif en_r = '1' then
        next_acc := sat(sum, wide_sum);
        acc_out_s <= next_acc;
      else
        acc_out_s <= acc_out_s; -- 保持
      end if;
    end if;
  end process;
	acc_out <= std_logic_vector(acc_out_s);
end architecture rtl_pipe;