`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPMaGC0iPID1v8XNB7eFRr2bdFGFPmfu1b4SWQH9aLlWykBImK/a5uFzAyl5/4JN
lOvRP4DU/3SoiOYRymkhadxyc6ZjgAfrL4OAxEB3wV5atcB8+nVFrynrtE4oi2zj
iKvw8Wj3JWsrbuIIc9kzmOeiox8+IaCsyR2FtLwvatd9WYLNymvN6vQAHUP8f5so
Kcb+3bKYoYu++xt+O5Er8CiBwUTrtFpdon9oA14ekTbGrGbmR9+5VbzrkQjOxQuk
OFNhZaQRcCfeSNTcrKtLOtYklOHatUcJxgXVXXfZdm4qQNAtqGrJBtkPtWyHX/1C
geZPwrFdB+ig6mpTClKfEfkvFFlzxYdNyCxLCNFDdJ+FomXupRmZjfAjLHS/5LE5
Q1CFkjPxrel6tj1BIoIRJyjpf6hn2ZmlUUBFcbq4ON94MS69wmk/kTXjBFetL3iy
1T9lwXTrUAY3VvV3Sf9GU+Us/rEC+MmBqpZ8r19QOwxOKaF2MY2MVh9NonG0PPGp
v+iqYXsEvmDKYHAZABf5Xlya05q+0N+zrJgGhEooGr0rKOaEIBSPMPscwHWVnpQp
H4VQel/vZ0dQnc49I3JLQ+wOGQ0GSE9DCtS8BWTz+ePGcvFOsGUEDq+SuP/wyF4/
kHF9a/cRWsAkryioLr2C5vM+F0Af9WTXpf1n58QuAT2TSG4e1RIq3+pgsphse+AH
AbcnUHLkl7Wre29ZrF9DWm/aFUzdK7uJQUhXRVvQmj2jxeqoK9gNpO+HeT40O3zW
VPHKpxJygUGDA0K5HDwXC91pLIN+cHdUwHiDkOt08HKHwqqupEBw41gSe2cldw43
ifiXMqYP2s72gxcFQ5uxQZk+oCeyM9sySTb9fSRHctN/sZuSK73xyOAgtjd1nKsE
e9VYysKc4akXExfFNSJD3wFjzGMccb3avUPYC4LP0u7vbheaSsHwuXxYatJDF1hH
aNpTwOFEoLk9on9wjCJ1kN4p4wvqYbQCRAv4NPbbv5O+N7sfBOfpH4ltGQdBUgzV
3Ew/YoeC1+gBDM/+zCBiJXN1UbCnuOD4bM7WA4uclLWzrgcLcHCh9+U2H5BzUWlU
GctxSayFJf2G1CQA08MNd2m+QHXIAK9//HyMlBUjZyQBZJ95SuPf3npso+RNUaCH
H58wj1WDXFhII2PETTUCoYJtPpgEQuE6iyFgP5HsH9j11ZW9VE9kSwzTT5oykf6V
/sx2Za9JIOuaFWkcx++IsijS2y2B3nsaSvobiSE1KTqTbAXph5yRvkDA3QMYnByV
bB5IL7F7rVPKWVMQLdFvo/vFunUCIVOwHWibuvpP8xABWeZgXN1YerHYI36SXAWq
WwLdunVavAOVyUPQRP9FbUz0E7PisWb649Y2UJVJapnPfFk13ji2FYwTLrVDCaZg
rCwjeOvzpDR4heJ3pcMAZj0ov57+LgQ1rDYCh/t61bI9hrgVAE6gbwaWup8+AcTU
L4k+pAIKRX4mSFeGVRO9X8EGRdcMo615CZq8unt6j694VK4iU0jWE8Gdn3pSgY/n
B9snAmEGC/XcETQiIbdZU9ny4/8jkoqbMrr5kKD6MjRwkDWsJgU6rLgghJfx8UBy
tp0jlCqwWun6+rL+ixiBvbqxhjKXpOvIU2YkcP8p97bkB89oRX/MX6bA82AZvxiE
8Out5AP8TGH57BW8ydSvCOCI1HqlfcYGFb188xOiodpIEcYJNXD42s+P62P7HcYi
GUal0UnE7IoXrq+LCbTZgd4rfXB+HrpbxjELZC+Lo3Yh/E5Uee85QBOYl8BXyy3A
/kFSBdJ7N6DY0ZI15iAviYVsvWz4Yhmr8rCXew/QKy2tHdzZWy+07mQNZolzFGJY
CsrohjjoBImpTbmscIzs+DOL+4VhwHytC/v/sAjjKVg42h0dUvKuoC3mFZlBHayh
ZgUFDIDJRq4Sbdq0sw2/i/auwUMasPuAS0DChKMUbIenHnHF7iLWFHCUt8wMoPSe
JDqJLyrYlJnoz9cwxOH82ZkVBMRTEi0iMaRpUprvSmJH+ygEh/FLqK5Mi7snB1jT
nmA5IhtJsd/dzVEKMN74swm3xyJVz1SuYFsRx2IyQyx510dHvu91BAL3/E3DPyT6
jCtQkXMTPMy3sBos+JvTEBOsYQg15BKSwBhcNW0uAm8Kol6BpVOE/rA6Re1D0vWi
f5tIZli/Jbb2OvkGqPrNaHGPXU5yvrsYjTVAj4jU4rBJ0OZWxzuHyrZoRwZj6N+w
Vfc3ZKGXOWkbaANccWDJtux4NNjKoTLuQfAr1LpNRDd8kAGS/uZ1x0gC/Xyki/2x
y8IWxOtn4KFc8oA2zP0k0Ah+iVTH30FuT30L1q3Q1IFPsyZCMv/1u9kKrLC/I78j
0ylsa4C/dRb9nN6eoVm93oBcCAOyTgFlNUqIAkK2LiTnwIKBrxIw/9MQHtxG6MA0
I1DMovvP120lDNWwJQpZMo+gKgAzKIwh7C0EZGBPFXED7nVLg05r2Z10ldyvW8Xa
o8A39S3C7jq3tyXdWEF2rlkItFRclvfvYvkm8+r1Pb+xTBi4ZusAEUgnMf8iL3rf
BeYgUffamMAZv7TggTmotBp6ul8o9Y2+HLob0PnkgL30Aep6Tjt+7GE2wd1O41CH
P9VAuMMEgPrcyRBNZlLPYA+HNw9aEBBqkSJcnq7SJV9stYwSdy+2gGynqsC8ienq
IktOK5NkhmxGJCNg/pirq0dsUy9GJ/kcuvc6LoBJzn7X5bRVMZAsJ9mMX5tGNlCe
qNJg57qXOuqvmVe56TjNtj/xIOdmhoSKEoMS3h+iMN5iXx9DgINP0OyyX7KSlANP
tFbUaA5ShZBzn9aIshyp9ELuesIA2/UqG3pLOC0MsI7rdjFzYMEa1/g4lLVbk6iy
os1hWkinE3AOboHjh3EJNWHJsmoppRooxS1+Xce7jx/T8+5uruKUjFvq2rkrlbFO
C9sTfjz4WUQiPsPcmyw6Yk7nubEVTAXDkQpjrlLgcwOHIrWmfxxVX14jx5MCnDke
B8DShzl9zaoHc34D34U1el2Jh9R3TMlyxZKSWKYEDNQROgsDJDEvpHHbmlkOixJo
YVYxEYKJ5Xu1i0mU6dDXlxnw+DsUldMig+hIM+//6IAkSrM8qY+gjxJveSLy3Kb0
BA+uYBBlnEkB+dUVbbGbIV8NcvG6uuoRb9SCl1yjJmJqdHyi9lLUvlpeGy02pmEU
DA1WiLw+6uRWyonK3rHgP4cwdwObsXxX497INsMi/h/JJb6q9zOAkv2Bvyk58KGh
bXgIyJWC5XEmfaYG7itjz76OOsdbM9t4Kir5xHT/vAYw7ebS46Fz6fnEp/5vRn6n
1LJnvEN4sspbFqG2KGv5a0shJPEYOrapQweqzei0BzK/Ome56MblqOH/s+8p5I3p
LJm1wMMU5xh0z8H5mkMzif32obIfDv2UCh8P+P6wc5s6piFMkhZwiR1ll9gviL3j
+OXrRw4s9bsn9bEtmGo+UyzyoVV373AM1D6OJxRJ/vCFTySW9gzM956KduhQ0ZZN
RccCA2LibGGgdKvV5spZfRQn60pVVP2s0XFUs8wm8uIbs+4/OOzGAgy0prN+vTX1
3pyaW48+98X+8VXk2HhOskx9T6Ud6NZ1uDbqwTC53KmPtLf3nBfwWvygKr69Bs2g
HHEaGXCa3H5iSF1M1Nz+mrTgPyAgy8uDTHcEk/pG0C83AcaB53xSPuuJ+tE6mz5/
7mne9wgHDIYWvuCufIOa6ah4fX+CtaYVu0U59P41dUbLX2FlX71beO9nrTqr6wLZ
NTjIon/IkXq/X/dn2Sa8h+1eaadC0rEQzpwzfobiUJBR1qlTtM0hgdwqG+mQfR9v
JeI2DPM9q2dpK9pMBFu508lwzP+9S4oRDFqyJijq6hyAA5I/NVxjNp34Wb3WRbeA
PsFa6buuQTofwcSFRmfNLEHSP8jtUA9QDfm80jyn9OrwDbeBepGtCIgSBLLl0oZ/
Kwp9zWTTEKrsP6BLkElFNq4XE1ar5AnZ2tbKj+GqRSjSkD2J5VpPeOT6cFu16cT6
1bgRZQSOfqyYhhgkpWrNHwEzWf395oD8ETD1jy4YnRtFJOblrzXyjdZHakgpbwNs
KSeGEHSMMY5C0YzomldgdhLflQPrljqr+SOm0x63frSbP8xEWc1bayYZ9EMv9eYZ
/XVMiXmfVVBvUpl5xOlQqcfNrfnOdTn0h01ZCoxC8383mDbCyaos3w4x42suqD77
E3+1r2/P4u7+RdImmrL02/JeOcmBauehZ7pydNp/OrYNWfqNXSUdeXcM4/YUW/ZB
ZF2fCD+4V5juDT8DRr4biNWAm0LlzKm22/FalgoDfs+nMa5qxCrAiwRhxZgkUipT
MYQ3dnVPgv2anEIlBugRGUi3E57FrGsU+aFuliBwiyGY/yNCzfgjChQ0qsIsfrUe
o/9k/UFMrIsF8TCQiTgQRvYvEnyqImahLfKrcaIVyVx9a+03CAGUfPHLoGRFRB1Z
a3pNiyR4pHc8i3p6pB7QUMRfoUuzg+YlPeL5XRst/5oyVnOflFvpuIT5Hvya4VQn
xw2Zulno0xdwrrLbB74ms8wFBOUVqlKIKkJFdMaFdSyRSMlJnQZKkWDwlxhJZVCc
Sp/HG1qoo/Dj84o47ktxqBxdRXRHD5ofEoMwLSfTRrZq01i7x56HgpzFcVPKvpKy
9XoxTfpwWX4lT8ScSJ9KLLTepvH0dCS7Wp71YoSecJ70FRvluLZU16dMmMew7FEY
RPb3bVia++PCT0Ue0g3Q+UEVe+AMSle1k3Xwnfg0xx4Tld61v3gy0FltugEGczXo
rHQ7RwyWbbB3q0PDIjGZN27S9rP8QfJ2apLGJtro1n+1NwBIIoUKulchHt2NX917
Unk/JfC4DOSyJrmKScJAUUEhFLlwlUP4ZVsucJXfZzNlSrQ+RVjaBmD6n43+jbyp
gnDVOpHlQElmSNScq47PRqH6Gdc5YDuTfkZUb6WYKCnzU7l3OX70xUQSEEd8Ky4Y
NwfGVwMc/DXFVtvn26uhw2JZ0wfsBo4AlRQSP+iAI7bGeb38n/GYJDpmWYv+plYr
oFnO72H7grDTGR2P351ZRTIpcH0g6Xr6khOsHtTQGANMbUy+qSWdEfblkyfil1NO
lYRSvthFIkRHnJfZCRvw5qUNKKAVzI7BtTeSMKqeK73K+RfBytVTkow9VMdVHtQX
62eZmkpQ8UozAXCWr6uwIj4h97iFCMfK9IbxszIWzWSQ4PNNOlrANAjXSYeb+gWN
GOacswA65i+fRkp9CV25TNC3BRUS9bLtrSZ4wl3zG1CW/6Hv4iltBvi4VSr5EeIy
Jjg9jrrjvUARmmWcSvgx3x7E/D3jWpWrZKZTZdQGZ9PrEcc/NSmRLgG/SbnMNY95
yurgsNjKEhEMg7LHg0F7FfE9YVHz+UwR4txf7BRCWZYZJ+OYnTeDTFJVjBlBhqfl
WJDWJprpGa0z7wGD3rDmj0+igWq1VvY1TojojmEWu1Nl10S6NaRZ0mGd8tz26REa
0+GFLJ2Qlxr+r4FlhZr6vQoNOXLpLa+DZL9Jc+WVpDykZbX1ogdB8bPGCtde/qN2
jZjodKlg4PJYVYN3XNos5+y82S1Hu4b2oBR0ZoX9BtsG3+ymzx5ogPNynRF3T+cn
wCG1/33ajRas+cLS0eAgYVzFTQcITA2MA9wblaXNems348iA9cYsWY9gJgrMDm0/
VHBeGTAIPgknBANaqJF3ORVHjp9ZkRXRG1grAT9LqhHxDhtmMdRlgdSMOaZ77cNO
SCpnIKJ5Wk6/NgvDoDbcM+pFzr5/pOthtRB9Hh4QD5RyjZDCx7+fxieEmBNgSvQ7
gP2Kd1G5isrl0PNNebof3f63vZzSOYUBLStwmX7YG/9dcSFmITM7lrOlZjJbU8qR
oU360y+XEzHtlhJRYW46kAMTZqrwzqi66TZjYCttw+8v3OlbPCVm1NEdzmGzicd6
NKp3UIGVFCGsDpWyhMTtEr9hfvayjzahS18vdbK8kzr7sGvkrM5vqzI5jSKW7BOk
DmSVpeLGXVNcwWGHCn4kMesr7DceoQSooTINsH5qDznfYYJ1RlpBKLYbXObL8yNJ
rdvb6eiMCoewONw71hzrdj4aPDAKtMHWh3GaIzbNGmdN+fAASAgBHQMKlcdq/umR
D9yInrSnDjoFfHat0fiDAsQyVBCKapeoNoXWw5lgcx6bO7tB8gSgv3X5LsASHLhy
3ewjr62YrZjcO39cu6I+SniTN2OblvTKEoNYLONvrSmzNsiglZGVmZucjtXRv4Io
m1/zeawZo2TODHhL42HbHJQaEQ1imo3u13VCBykLFK7cgdO3CcVddOxLiA+bV5Fy
OORp6QDoSQWdrUITUmpgw/BmwoJSUReTyAYh5o34TRBcOlJwCVZdL5VcV0XUawRB
jL3sVKRaZI2Bf4CZWUBxT/gV0XgBecZS0RhZwAQfNXmVx35Xj3uQfKiFqmNnjR7t
MnxSsFzpFkd95DfqIZdvBet0ghef6hoTF3Li5RRuoNmMCQawzfHV8EBjKi1RdJGp
bZe+0Rc4Gixao+MKi2olcJcCpuO2wkFvFPF87RA0THHyM76JdsSKYA13FR/11N0a
dgfh5mlZ1s0JyCYHMIvLT0ZkJgafuBmljI0i345YQJ+yBj2jpb38wxO3SmBOkcEP
tax/LyVGy644a6CwzBvLbcugXp2iQ2igewtTGaJFTF9rrRVCneC5UsLyXrGC9ee5
y9NFKmVerAeF4iF64qMG4lk64ugdqqQq55fCyQklDNk40dTx18vVp+SBhLKD3bO3
OsJjYq3HjkXKwdFhEHRIBzHqcd+5aXUCtE2cQYwrys+DQSS8Zf0NlStTYeBxsMx5
VJJCuBIGk/F41llU4xrlQOL11VbiWXsmZXWMWZwEif38z+WFsa0NbQ7uSqqQBCG6
01VLNfSgTqJgAuDy8DpxqcZYCDAEH8XPamWYkgxbZlBnQ4Q16jzoyMY38C6NQPv4
ldc4xlzY/OmPxaIBfs6I4o50ycVD0NYOgYCCUt7EbMWEgjN853frGstFyZojEMP2
xL7FWYOe6cnFkTcGIUslMF85++hx+IRqyLUcKK0++LW5WhXPcOQU7wjgelTYihZh
Iacql14Uy7N4nS9K2Fflnyvz5fiKRycyJEMopfhVZ21nB3TYoSYcm4mwR/Yj1XKZ
Ic3akGm78MCv+rHnICdUd/IKSfq8PgWNnbkEjGiR1WSx6sixzr14XPKzNDGvK3EM
dRvzigbUHGSNeBPuMN2UYo1DY+smvE/vQFf3hxRKQlT3rjcFdeY6ZxIzXItcwpsp
dFSIT9zKuLQucdPmqPjIRmtUtFWQ3c9pNYAwOq/MpGssOVtp52IKmF7wtrA3OBO7
LB1jyIWM4au+WNAA3vLxjszQGeWHKkkKkMAB4XyGJM6vjnpb1j9oD1xyzgsaYXC0
HmfXo5FgRl94iHTU4lwQjD77AnPHO0J3Ft55MCktWmmGLAI3yJb9nmPstWFzjLhY
L7Mo7shGhURyR474bNWRw9TY6u7J39JaRvRyyK+goJUOa6TGynsfoFlEp2UYbGT1
KdwPEEkomhg+lkAFjkks8GBXXgp8tjBoLa5ABcQ/ReLeAyJn+YTQTdnDFkHcXVai
CWfUIau5dyf5HuX6ZcvMNQuZAAXe6zPVykeI8d0KElu/yj4GJQV8QrfElE7xY/uA
msPwkaN0rWkz6WKe2k2dh5o0gBDIhBRv12W1elzHFRwA8npeFi/QRYrknLC2PNk6
up2xZ+YYYE7XT1eWkNX2gYUx06qo7FvKdLK2VeNRMoPH+68wTghaX7qt39PTCAU5
xRsCr2jAh3E2NPwdgWxUE1up/VZdkKzagQDGjdXPX9YAkeVosVE/4VbGDmoPnBdL
nzC5QxBHpmE4DeMxQtDnfUqsFM5ImnbQJn76dH+zlNV/RPxCisfAYsOq+ueyt3Tg
nkiXowmq9l4b9k3WmPxHLhuPocAwiEoP2zsNwE+RVQQzDynZ0kUxgq5TS617ZQXk
ndK5+oxfYqE+BB3k5Yr7DlG9Y7nVo3Gk0OkyrpMUeFLVGcIGY+CvQMBSEWUhUoRE
0e9NT1w9i6zuSnOJcYqCuIMLaxQjqHhU2raP3ybCawecJkv8LTsTx9fG85vpjmIe
beLCovvGgpRiQnXljK4buN2YtEoalgSJUKmisOVbYkFHhHw4BT4r4EgtIoaWxZpd
1Bu+JhhQiG/fwCacDWsKsvOMdeKWu00i6qmiAM+Kh+g1400iy965XF4EHXR8dOXM
aQbMdtAP6hnmZgjRugIrcYwEqDQMYySie5vZFOhoUrZJYTfE1HmkZYzibR2VaUip
pVv6ZIVZLFd79a0YZqoyZpSd919kwMijA/yQSjE5ZZAfZFQPfNIaLr7C6EPErGpb
Tfq2oHIbOUIrSlPegzX6KD+QsPDfPU4t27di/nUZ1bJ4UJnyBveIF/DIWfV/mL1/
es1aIzNo4+dt8AviCFDUADbYk7URj5evRn7gIGVm0pBiGifHu0lg2f2fN5cS+gW4
DEaz+PjV40jHGAh6OByG0vpMgnIBxI/zbLkenxYKBhH1YyVS/PGHFBRbCKVmz+Av
Eoc5q1pMZ+4pYDzhXLoigP+XFcIruS5mv72SVzxtEzCs1Rg4pcwn2fe61M4DLLg9
sDFgT6hacUsExC3PWpIdhh8sQ8TclyVjPKT4PwYn5P2YeYQU16z7ntxsjZha+DEG
HTOToxeUTTYiyT0zfs681l6HS0gAohCZj+oVFjKbM9JD++6mUCS1Ll/+B0Ob0wyQ
TgGg2Y3lVBS0/z8HpRMmARKVMZ9lR8lCHSjVBhmauv79DqL2A9MdZqRe7xaoNiMq
enMeuXrF853lkuySjqU4rL6UCMAs5/VKL05evZ8rzwHA05VVwsTSGCcGj3xGcx4o
zed9dEq1pvi4bztBmQa9LBtVBimgUD346apMb/ClELjdPvNHQ8pU7hIxvEKl8WaB
8CNMynyLO9rVq1DUemeSb/gLlQJqEtF4x9fE/gJB6966ztLmscv7AVJHBCnuT2w3
1VqHUAZFi8yaQkK5ZtTY/6ppbHXyFRQQ1vmRuYDVBh27N4oQfUCE5uPG/8Xs0kQ9
rOYuvPgnlP1CDpbXDGl0AaD3achUAhOTsBrjKd8inAtohjm599TFLLQD4WbuQCp9
GAPZsdtgaXcEuTjj8wqR+3iM/S63MJtsa/haz5ROwdyUQLrJf42a7tUt6LHDvQYd
TIA9kXhpMzz8VILB1r0mg3P3YydhOdiFi0/Rs7TSEdgYHEAFuv4x0ykDgmv8LHTV
0s3IG1+T8Pcp8qbuLj/84qhK3IIi+tGE+PiVX/Dt7cZFjgjeVKABWJ1bHmXlP0GS
jBW4VJzLUcVvED3gaaNJGkP/jxpgNZt8rIad+5tOCRJKmHIJlMWCIX/tyrd8g+O9
C62PyHTYJiQEv3DFo+QLxANb/Vk6C0DprG2QB8shWUNmAXwKl+4mOJy2QF7dFYa/
c3PVqVQSg9prbmHumMhiOxVol6YUe6hk1i7CucAV3oYHRqEx5foaaJtEXb0m4yD9
D6zEZCGIQD87643mi06lttyIGdiM4CsvrLKvH+umqAN2YktSkGxMVm25uWcQd1EK
d652kEpiVKPbIueV1fglNM6t7BchLWGwnrVLdEYhAbfEqLtTyVVzg9JLbpBVsPke
rIzgYpuW2mYN7RvFissDzxJ+w2WrDawlKG1K1kTMD0tLBdBdbrQajm7ndvDdJMUJ
/1Ocae7RSy5qxFibZEP1V3VfnTKrJxZ+Bsp65+xN/LjiUHnWZ3CEbVyW2PGW+LRt
/JCncTG1XPBPPKkyUL7aypin/p7zQkqwRzupRL7ZFBmYj3Co0PPwWitJ+naMHiPO
+YgQ/BKBjwGTdWUM7Vahj5J4/23J/ijqOM8EwWwZHOEhABledSbFQ/yPCRkyd/f/
AXw8Uh0dmEQuvpez+AYlVga7BzP+UWyK1Uutv8TM5lAqlBKNkYO/PXty3WhVBAqB
uMbdUon/3saQmXmQBQIx5mzz8EpG+RruG6mJsLKOjxpGecvD7flzD4WfY2to/9o/
bWwxc3JYP1zPiHB1xW7UzNm4L2leh4qfYDFTfOnDwLnOaQji/kyahozz/MFPqKVr
OIyofkMtGw5H/ybecift2RMi2OzoQl1Br4Pxmkr1k0cccAdEEi8FzCYtirM7vD2w
pvTbcFsDRg0Znuc3KKICOwwhkBUfeKWYvk6vgMvuPFZD+sSiUDNM/WcurWb+Japt
DwsowndkPcMex6Ss4tTPslsT+VtQtM2+HqBFCD0Q+Us7iuIvCdSmUu9AkuEje8dE
/MDX2Cj+obj1qsqXcUoV7NZhdIQpi8nYeKg18TJaj/IgQhPX5gOwVyOGHyQWbLyR
Rzt7RKc5p6I2rdoqgU8M0M81Uxnaz+4rNjuTzyojOTPoyP4n8mQUQx3GN5zmW4N8
QFSwuSvA76xjZvXu+uFdT4z5T+pk0WUrBlh3RShaPp+5DUCpOCD2rQeUEDlvl5zb
ywie8eAar211xs283xfkwrIZx4v070Par5TmLT4v8PUNo0oJG84lLla70LPYxsG/
M9W+RPr/yRIg7859fOtMtQTsZZgpvLUh3tn012uh48TKJqd9e+xlkge619reATNC
xfMjHaaoA+L+qrBR018a6+KUpqZOPBPlM/+suiyRwETXw4xcRoAEjvlYGFr5Q/+L
Vb5EN4v7+ZdX5ExCyD5NeHzwZQuxZjOG27GwKr7th3FQdpXOJe5nq7M1UUClr/zQ
Kghxq3N9SnaKXS8/6GngcNl6OsYPj61PyY2fJSv2bsXUjU226V3y6+2B+lbzz6Dz
O5Yh8fWAUAHzjLiQM2hlQ6I2yVyjqzsknIwN8ylY2XqpQblD3O4byqhTmoD8lkSW
fAQqaDAmIju9mkO31wjqRfSsqN3GSxtKFGTRyjFZy23ooQxtBGvMMpYdZRiTTb6r
XosenxY7TGYM9uqfM+IChalLYVt34PP29xk+RrMAISPW3JfQmSOJPq7zyLLd9lAd
5mfQn5ajBGw8nsfly/S+ytT2gdaGRioILqe5SPk/ee5/Djah2yRFPT0nApxibiaZ
raVAWUfvZFtkPNsb9mv8b6oyDc4AE/0M6Y7AGehPE64XlkquJ8F9wmSGYzD2WZaj
sOxM2TKniPp58tg2vNxDjZICgroLog3zxfBL95c1hH6LHZqo+J7hirVI4KpL2qQk
oUuXgWw0h3y7CmSZQxM40buDRCDzeYuydSIjz2UczDn4v7o4o0V373vKlB57zhC9
Cx3O32g0oEymRnD6IyoBp8cXGmo86YgY0ZRamZiBM47CIKCIKL4Lyprizt1EuKsh
k+UXPVseNjE32kVLVwf6Hc96A4QDHqbTRV8mK6pVlignW+CZKcjdPJjWjF1Is0M3
6aSZ+K46kW6e29tUWlgNjpwRXrnnb9fhABjcO2WqnD/JesjpPry5OYK3+vU0dU1/
PjH0UVErqIaP5YjdM3AcAfaNpkosBs9bRoD3SeW4LlBDeI+SEU1Ik2sJcACwYC++
m7DDxuAzsKyyKRXLeTd/GSZ5E7OAc2k2zm7Ey1BwcBp7Ndm58n+9m+3QMEGIM3f8
ae20j+v7FVsvR22vUNMKREYkOaJSEsVrgmr+z4Qm3iFqSlkPTEg5sPsXmkRxQ1Bu
xFVIKte1ytKNSDSvoNwkIuWsnA+ed06dlZx4wMFejzyl7hRnXDF06nLGNsH4+4Dr
0RSxSiOve0c0vkRz5Oe7OaOXuihnMaVMsSHWEpQqeGZVp+WOYYwRQvdY17Bts2zq
q9p2KfaQ18RJnRCnI0yvn1iMPYjiSNbZKOSVhTaXwpQrd6CO6mSZVwayCWP/oPdH
WBwy1wGsefLOXYffh65Le9J9XxqqVwVl88hn8k6st7SSghMc7c6OAyxRiGk7adiZ
e+mkMp+CAbAGlzSvq5Jbpkh4GA4XssqAKEdceIRNLsWEsUhoFZvOsq93LZtv0CbC
VxsmcnpB1WHu65N1pP6Yu99yiYk0yTw+BUOQDpceL8GO6xHofcN6bujjmtqACgWF
NlOWyst612i7sNNmGlgXl8e1TMB8gsXJF6KsxDRQxHr0dt/c6+ThZTzC568kbPKo
Wyk13tk19JSrtqgSrPg3fn/JzeVZnW8x3+iEu/cLSyyKv7drA34TXSRY+XPo4C1g
oaTiOvSuqyv430s3cRxuPWcRgf/wrZUBA/Ua6NRKV/gpsrSAiI4Bo5J8PPpi8o2+
EvJ+HOMRytLSTaCFIh8wJf3Z9vQaRP0nOcZx7/K+9lRO0pYfTnntHmcbIytCjt0n
SfoCyADzLETIgERHSWDbLm3ujcv/1nDRAkfV7eiAwXY/a9/b/d/3iuVDrGHmCFhC
bAKCyLTtKB4l0KOu/wjtd6Zy6zxhU5NsZqhsLV4Rzq2axqrG2iWp+yEezVJFnBYq
7twzIJOMmLFS9i1ZpM2kmqaUnCLVqTVUALDNab/cj7drAC1EmhqgdlYDMwkh5iG7
2ky86SWfA5x1Cl2CH6fUUwBOkqa1WjhKAAsvvV+vhZ+D+VTss+3pvHg1nRFqLjxk
0kVCOlcPhFfGqnzbNI3IQFTBXoMCgtSWhoOp8qTcZU+QzS80aJY1/cTdpVWVEvUu
21b2DMpoxFlQso49DbSR3mwkOpgheBwN4x+B6xgEyxasHY7qXHTHwan2hFR0sr9q
Xz1hJvL2UeleMrJjtdcvCvdMCVQ9STdewtcpH5nPTFYcWhajGVpMcH93f1dzw4Nq
8NkuCKGZKQi/NNL4mNxmv82zYXPIeencfNuQWGwLWoB3pBXvDKS7h+Nr/RdAqAnZ
XYHNGT07JRgcEvlv+GA4HUa4fJC3+ZN+8lIvGZt2uEzL0E0hDXn3XQ5iBOuchU9N
EHAD+m7r54KnlN7V/BK0LiwVF+d7RHvmLaR1pZln207jCdCmowwBQo4KyQSuCDPB
lTrhM/PbNZ7jnbXXMhhziGANai4p/zr7NiKl/PCX0Vgal91W02VISNmGm1X3YlxS
JPy+9qcOizrNGMcGmpCQZaf1ujTblw8xYutWUL9AEe4nPARyZ0lBv1OH9ObZ/y/9
CAa2+b2i2ZqdZs2ELEaW430B2Qq/QsTNI3x60JxBOQAMezS81c/ZAGpjovCUd6sl
g4k0OFjbKP4bMNt/fb5a8mRX8BQAd7sxGCM9h7NQO3U8s0V6qYneWI1zQFxZr2/i
u2Tmxpe6RmfOk65+ek23gOqverdAjsHAs4naIS8FRN57FuGsv96NOTcAnaWRSsrm
ULMw0S8H+rKSv/intfiYo66s4RO4jtWsiz9UNGlkYqI=
`protect END_PROTECTED
