`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1wT+qhrjStf8tmpu5kjKvCyKZvygO1Afq0eQH+tVmsMCOSbIziBqngT65J9Me3WU
dgUfo595+Ca7YKFR+VzVH/O5GqbZdD/XxTffBd+1YN5Ci8PJSQhkbBY9+d3KD30U
Q8vIWpZhwzoY6wv1EY5+eWF0Tcy4jR5erofZf7NvtUqk+xtde/Y+d2e7zxUqzqaX
dc7e4UR8sCrX4KzzOXZ6e+S8pMtPxW+ZBptj94WmYnqWymLcJqEDcbRPRRpA4UIA
JZ+I7oLC6U/+UghwFFgCK87ZCLOtI0gUF5Aw5KUFbFf28vUU6iUpf9VxZxldGsAp
WqtOOIJ5Z/zexJI20q4rY2KiMPRhkViH3ZEUR50cwyeu6XmEiKsZx+tesa4AXfir
kwuY++XZBbsEkoDboTqWXyGEu6ZkKl4Y8hgWziP9DnvhOSGEowsCIDF1jgcrZBk0
/vFrV0TRlD4HpwH/BBLTo+P4bQKfYJul00nQ/IAlN1F6O7gqsmhy7Xo2TN2fNP2+
bLnggJS296d3+iziVueW7RuLvhp0xStqocDDjnwT9iQiuR9uJhoqSWZoLYGfOkMX
V9YVL5LVVybSQbRFHiMK5Twy/RB54WCQMXxqkJiGVpyUgqVCTjE/ByBQxq08EZ4d
7RwTpEd6PhYYfiKUZMvxP9wGhrrho8uReKI+bPrtolLM2mscXeDNsfNAx8+Vwkm+
NBGAN+T1Qyi6649RaKnDk/rA7gg/c0G8lOX4uSmHG1QcQwxr6hutFcDfjjyDZweD
R7+DrG+Rtiwdz+WJra2DVsz7z+Bc3GDE4/U+6rf76DDesZQJSkMP0vauIq+aXN6L
9RUylH1byMOcbtmElu4lXZjjwDPS7UBluof7+nDlfC5pSlk2LbMaAhShT+JtDJfy
xMXDLQ2XwNKlBr2FfNKWVlSN6/9tTp1DEk4nIm3AmQ7Y7VSciezn51rkaGoa897M
7kwianwXKsJVa8DO9F1vSuJoaUleGlBx7eooYicMIezuKNbzHUZnMv0ELSsiOA8X
76nQ0PSOLOAa9KUm3bOz0Rs81lehoCBLos5WkPjUxhICZBL3dYPx3MSbXAFsr7cu
`protect END_PROTECTED
