`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6G8CyNDMxZuA97vV7p1xJLKgUrbAD6COJAjnKU3+1atALAS7KSGy7NxdTGUqHFnd
kfQA1zTAz05askjx4cOBLA5GR9FXhfiLtwBq82n2N9ltDTvL5/tH09dvaWlMEqe1
wmn8pUzk6IYlgwvrnXYqILTDtoxZ0SUhR5xuMdneoEShg/wTpZoSuR/4qnc/4R4k
DsPXeZBuOP3CWB/yuDFGxbR991oyROZrNL4pf1xlFXzshdxsJz0Dj8RpiLfQ3Ixo
gaWHIC0O38XcrvxskmMNo0C6XtH3t8ca4wyPHoVTSHb8HVU8z4wB0AjlJVVxs2Xt
sEvOI7qEFnDuahqNpTaA9uXrmTy9bo77eHZnq9iTVXczuWHlt8uvPXQBxBgMt3UV
9cP8NPjg9YLyEPdAkiF86X7Y1/Nxfp2sIfvUSTcau7yFxrtJa7OF3d/s9mh46pqD
MQliDlTajzdeu8/O0H032JM+a39VU6kAn8Qs1TrasOJwGxkcwlIPjkJbB4kOoiCC
0tYdcRMa3qWFHz9hWX6Ot7i2z9ScjKNHRcnZg2lTT6srfhX4jZK8duTZxgWU2jRQ
L3jFGdCnRh75FZhzxztBW8iSBeBIaT47HDrPjZCrUwqJWkxCUL8DM+dGgWV4vD2Z
hzRcNmWHUGDLqXJM+pGNPZ5nEjXrE5vT+Ob6Sdvkw9jfVHVz6UXu5stmM71sUL1d
r1YehnwlJnVTmy90+XF3PNhUEYgUhknezCBvXH9KopTDbB5iYuctFXfMY6WQr0hF
wuXHqncgVlAJx3X19MVZOadFSHZlj5NGoPXao/sxG9nmdT/mDkDhfOqaPynXNhds
oPpv01JbOs1nJm/LNhmyr56wGmZQN3rQwJr/HZ1bwUgP2Om3+x5VU8FhBJPtLars
BBqQg2DsSesCF2Qp78Mov13F+x1fMnsoe8656c4+eNxyTJ76MtUpSGJenP4f0D+/
jSv46lnoXJamm0cC4FeGOtHhqpC9mSLBjbQnHTIi0eccJGC4UwXa+cbjZpWDPAtg
lWxPxJAVFEFY3qGnROzMTPOEqWUz6vUFj07YxRP4XhLQ/b9XiYQZwd3cYjtYJVcr
eaqsmsEAd0d3m+b46z6Tu7nPaEkP+wOQi8sTjj+UszyZIqWsR2cn4E8c2o4CDECv
Y05MA7uVX56U1sfSVLP0ImY6LE2qTkidNaK9pGV7m5mWsq5Aw10hu2WF0c3sZS4p
K7P5X4R+FbuFeTwhoJTKxL6X4SXHw5vP191v96dAsE0qfkXx56WyQ7iYXF89A+y0
i4ncDOZ+ws5CFqG5ncWbXbbbheMLsrv08gMq+7P4nfJHk3w/PIGxrJczlNF48Nhp
QKRl6D74sbSht3ZrOVGjdcGa4HDeGxvv9nHEeR4VWyHIK3nGgirOtSQdrRZiTIq1
957UMWJpHvKQqpwv8eGDUuhkiQQUfh4BNb2euXbmSVctiJnf5FNMS2YHth2sx2dj
JG0PrxSMwdmoHeuILeESuCUVxqvkNc4S2hFhEaPk3zWwCNTsAOyb9r3Ix848R66t
7GF64mNQC7E5SlyCqnMCwIGscjBYlaK7GRxzxSh8JiztExcRv2TSFIPoGvyqGbaz
URynu1xYPWxj9WSqPlLsYxGBL1DMpaau3oHH1M3r7O+4NIFXrBCMEKszEzdX1fqJ
3bl2tLXnMZsDLQeaOhfE0iPH/Nuk7ICMRchXzcpKCFxKJqZY5XheN9Rl5LVlKU5Q
b0YeHaX3BE/8YR3bIi7dky4gu69ECrZ/vJroTjtnsRFJH4UaduDlGMVgCmf6GtbU
gOUixnamUWNzwfQupVI3fWd+OhZSQF6DDsEzzmtV86u56jwmcdXs/44oZGwduTyK
QLpCwnOKt7/aQvajPvyq5Q+V1w6y4vUlv5HiJEviWDvQgvF6w8BOAqlhqav21jfB
bAZCR5R0P2aaRG2JKeIApxFdumm18+f3hmR3b6TrWy5xfQ7HSdlWhzua6Nv5apM5
2sqeqnctQ4/vEF9INQWDA4QvjjhR8r8770L+4OCtIimh3nMmcRqbaJEjkFYeHcu6
jCvAhaKeV9Bn6H7whWV3BrT3MlqQMuTvbfKgT9kfF46k4SmrpkzuSuXd49w+rob4
FEs+pLS7huOMoqLuQLz8lXSi/vCr4IoIzJDM79Czcu5uF07h3pqmFjolL4Rx8Sm8
/bmChSX6cQePuhQjKBaMs3yfIr82cuO4UDV5uYEuX2J/fyDxncLD4mt0FHKjuE8L
4USmZe1jV3dYg6+Va9N7YdreIwBov3MsJLthC2uY217T69VgRnTzQDL/3dONwpq3
2xxGI0joZpn753Lj3f2vL/dkoAdq9JbK2Y0fDBFzP2njRudNGRuI9BXWp5yfzYJV
ddA2vBRWQIJ7H3zSvR41eFy4J0UJ7/T4DhT7V1EmRKaLZx/mmo7Wg5Vr9JXgAun0
UqS3o9N595R/xzlCq2BcZzOqJ3mb9xPFYpG8GAgrsTCGQCrz/bnkLDgQUbUEYKQQ
fcI+ph8dL/lxZWD3riPOmbuMmAdR0Kej+kSSq8mdWewXb+XOSi6f8DUdqc0krdUS
cnwChAQEGyFlghsK12w0kFLvZTrndtZ0fSZjx3Pakn2H79TfsPmZKGxyhbSAZaTD
3npCZInrs27yi6CEke58wDxZ2Kn0Lf400mfrHh6HdJ3Yy1WhAu8jtcxTFhsBIGkA
26saGVfVS1HFBMmmVfzFGbKCaLL0xP5e2OzRDzzD9gy3xZn+a0HgeFS9nWn5amTO
6s0GPw1syKToN+WraH24fyhyUwsdTT7q6lp9TpnF3goWFqJAbvFRI6VoeHl0JFsx
DPFU1P+ZVHCGZmoUXMxZ+Oihv074Jef2Vw9zgLKFPgzkvHg9FWcVFpd/RBR17LhH
61FOGsw54ZDt8/6cAEwcYjjdfEORfad8dZ3kkjt/1VZI2L/0LKVTrzGSXqtrHqEz
BZn4DriyRQ5zDrOuQQVP7qJLGEbbmGDx/4aiZDpOqsJI3cT2kCFB1RnckA+TWwAD
5PM3x78gy9nMzwGh+4/+fQmWJUL8l6njzMz84teKuG7YGkRGiOaSg+OVXndjBEO4
cYHG6BO1k+ZWfeHJZECrIlQJD2/wbpDNmpVnI+OE56v6q5CxtGNRjrGRYQefZwNe
WpYLTZarWaTaByLhXDOFvXsmn4CMo8abMhXGoefyv+RTQJYh8vVcbMd5Edj20tO4
5+tbTreI9n3Oy5BAQb1CeFOjiT0iZAjqAaHUTAcIDPP0Y9KNGBmvjVKYQW31LqxW
KB5LPwdgQRqgJofievb24DwGpE5m0LHiUwTDDNMwDNZjqct6F4zolWgP4JY5YDS0
AXlvCeTd8jwY1dU0Uh48mQECgfc6ofhTUzKydkbN+UHoSWZYQfzsda41xCFgTnow
sRsE4JHNCghahe22RHJAA7JClD6WzC8fOUZUkW/9+gtYopLfNQ3wZJlIOh8Pwyeg
9ePBBNdAx2reAO0RRYwZhCJAsM4ts0h8rt4UtR9Ka89pozlB9mspQrMptrGMuzKE
F8bpFZgbjQKh8E42IweePFxL0O1pUA7Zn0X47hewL2fK/OainFetbmnMEx+gI8pA
dXD1r4CVG/JDaoCKfJz+wfE8lXMi4u29OGegOHVsp3hNQr/Xf4Drk+cgMgYtSiJe
zGfrPGCDgI5+tWNNPIQcv0AZyZWuvlLIJDF63OQFRAAOSmm2yP4ICJ5WWtuXIrb1
`protect END_PROTECTED
