`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FtUz1DFQj/vnYqg/8PRMpfzNc3BCsT8OUyNrQrioDiLT+oieytidpmpDJcqpR40t
JadkUxPR+1RJpFikw3OnRHviqDrqw5CiCXf0TUqIr5Ee0tt/m6F1cjmXSYL3/wrx
D3WRBO/wm37uOeYkPaFSpgR3pzh0QlEYgMCfp9a56FfXp/Mq3HMcJSbPkfmvfzQ6
kcVFngq++rI9ohldmiLLgC/1HI9uyPZOgFgLBtpzR8jJd2lYZuEVvI9HAX4alLt1
AzlwLXq6XqedS3blmljkLftMqwFgjhXuiKx4hKQsLz4SOO+ZE0xJwEeoW2nXAF7g
0FeHBokLCQLzQARz4tT2XaXRz3bfSRnxVDe3YKJBAStTTjhT+dfg76rxbi6HAq4x
rzuTri64Wz5XyeYBV9d+McAGvpq4nqOLfRWDbO/0lyZTogU8UKbVPsV/o9afbqF0
3NmateTvhEJtJqYNUf1vRabbHrYojYrdbst0dNWCvjf7tpmiEeHfe82x+dRbfWyC
OnVSYWqKng2pMDnmSQRYmQYlOEvKBTa2L9tjPKiMXxuKiiBywnxjuxKVHRGlA/iP
bPEuMuoqfjfcg8yIyf5r4+7+yA9YQXC5aDssGxhIB6oxNMOd2WgUwvBSSry4ErAi
pJvtZLF0fdhIFxGkaNC5o8A2RBhU6Dl0wJFBK9qaOEPgRw9oNzfS6B4U0lKSQCo0
FwMMpubw05D1K0ou4IUh2BtD9jr0s02sLANPVW0+HV0TuB1MCcPsDuLXONb2FC2G
JEKdRiETXpnR0vn7qBrRDXvReu9EntNSeafVVKugemFO5wFNanQes6zPOXid9xjb
wcEQL9rBl4Y4GqXgcXML5gn0mbxLttHfXACFyd5oFM1kHJAI1ldY/29wnQjOXYep
d/mnv+eseGmBlzIGLZqk1UiGeDawyiCWU5EwjSYxpQTho6AiEFD2sEiazio1l+Kt
551ejH537V6ETthopJ0OOisDxuLcNijtqWcznTnGO3dCVYtoFeSUjEhiNbkHLzp8
zFLHC40QK52U4RQZUKVtISNnGFP1I6ZaxUp9SJ/idQkhmR+dJPXJc+yL/QWhcrLV
qVUyBpZi4oYymR/Ai3hVqHSSMAyiv0r04hXjEfgZbzYedZ2VA/KZsC9QuXUMDyuW
LL16AZIqNmfZD9tL4P1/CXqiJfXMwFHL8rCnVWTtEK1eGytygDot73/HphiEcoVX
5E0JID7atO56M0e3t0s5hNbzZP4jqWZa4fC2dGuC26XQecOWChwpyFwaeEAJoqFF
IvVXxr3rLbI1XJ+81G0a5tMk+U50/l4f4C8puu2pfXUVUvSHIsiVbP3VRH7aZSZP
MAzWrLXDVtkpRMszO+GB7EXKMJLULFsUmr90eDHQs+XEQdaCxowMHxoUmGr2+H99
tst7D8ljUrvQht/nN6Fvq1RMHH+O+kkBFwYJH8RODB+cV6qRir49M0YNGjpwe00g
cnINIvtUn7qgEqGCsXHtykL8w9VkhWKQMJWIvpDVXCvTyTeKDdixH9D04Yb5TqJ7
qQ90FGXdCAUCsNuLf83ToEgaXeNxpJPOU9ATO0DdcOmlxG53xR+wHz7snHALnO8K
tUKrCov0hqosYz9SRl30Hd8fo0WbN180wlPiJ9Mv193G8H0OLBfqCychhHbKKuOL
58hxoFCbKAgHhlsPCfHi2T89qy2pWgPzfYNmlZ/5WcDZbeyaLRsB9tHmyWY7EAAD
e1z5BvWkrKhZb4SCOSy9ad0PTIIFcllqWwe8YG3grSykTaAA2jc751FK4lLopUwY
mVjadAHf02zIz1kw1yrm3ZkFtFLzKzopVlvb3C1NHBIMx8osoU8xkz994uhZfd0N
48K6N0oa1q3WWtu3I5GRoua8m/6H/xJzX2AO4y8T28LnRgNX33pKIoEjYbcB0Rpo
c04vFqE268pSW41IK+WhUkXOEEUXF1TH9r1DwFbS4C4A7tx3nsuih3BJs1YQmU35
D222vVBUTrHz6mnWa0QDVIwLPwUGGfA7SaRZK5Jim+psAdYzb8ISbPSeqYz01Hfc
f9Yh9Ot/LBowwQ/8Lp3bn/7HRHnMUPxRM3apuUMfVU7kncHKgcM0YBjgQxTyBUIq
Ht2uIA228WPM9xwnB4SGBOFXqCsAlpTWsWbgXuj65AMAjmw3Z5bh5fpk0+tjLCUX
V+4i94kjNSIdv21QN2e4MDrjY/GxAlao5TH9VxjA9zbGBrAOYzYwjH7yi4G11iUG
8yVVG5NFUiV9L8Wij5bzm9DPt0/Lw9HpWQrqWi3kIzE+AeDKUqofcaFrzo1WuVyu
dNCQUdVVsmX5PjSfILACxB7SyGWLqXUfs8YauDx7j0qvayqAnurTEu0fSpYE5gbE
svGp34jI0v4x/YjSffJc1XnHWXDhmSArzH87R4THkcmjxI4ae0RB8EsDey01Vde3
9LIEK1E7XAWqY2ZDwJ7z8PLiGIAiF6rnhzSqwOBV0A2q/PAwOKMLRuWbvaoVJ8fo
fPvk37gfl9DU4Hiogcb6EN6ScURebRNXrcCkpsgcpK8QpsmotqxStGmWfYPXl2E/
14GoxufeOZxKTFltz5xG9ELVPIMcCUgYjWg/VFCX1adcbKgDOAnQpvP2rDU0Aj1K
+AlIcBwAw6RjKrsqaUg14WP/y/J9JoOrzrWaDjeC7+5rJ9OKulYsZ6z/EG+Pqoeg
AzWhL9Qio+BBokXYoYmpP3vbnj2M/VZdz/qy8xbiGfZuwnfJ4wtOExjj9STPdpuo
c/s3IFSRou1dSECfIvG9YOGAsPPAYlIinCWiL1eAtcrJyPg0Vjq4I38xonONfVn8
gcD/Wo72ZjcYVcAQ9DH31J8naV4AfirIBV3mmPoZohAaTAzJv6rO+rD5id+LqwgA
Du5Ax1WWB5aLMEIbxSowjRkMI1SzgHKV7dIQHS0AjcZuQ/iOr5inG7SKaa1U2Fgj
BKxSZeOF87vs8tysitMqwiTv1sL1WTBeUIHxh5/c7zZxrTzx5Y0bvds67lq+7jfQ
381/bhaDb77XWiRlEaB6gQ8q4FCkV3lgqm7jHIhKiD/Z97MyJF+33oyOA47cFrD1
5jmqNJh+NJP/sOINYSNgbq3Ze2436j96t8Ib6BTQNl8KvJ6LYVXrqBEsWeRjFU/M
vBy5l0k7dEaEB3Gg9SaQ7bQqPZJ5tJd+gXcHslECi1DHs9eGSlBOfE8f1874okXR
HnxEUFwhdmDfQYnyR1pob/QLISH3O84vTx0QDAc1saaQ9MnD3+/70Iw1tJ8lebU+
ZkiAymtwvzfh413Ls26gRr3yUhX41pb9gZCU9uIarELgQXgkKbBQDmQb7ToxINpH
54frpAanZ8p09sOdPVn2Z8XaUXto2T4XfnUYVvjwvw3b4cUDfbYZOKGeZo1XREsR
DDBwXLfFIdmNUfiQxFuqADgukLOW12zitt9ZvMs53nTV/FYA34U1MagS5vSSddCS
PslC6ZCVela7Q3Ad1p6r5GNQd74NtNxZDo6MMFwtDHN29twTaTkVQqPfw3C6R8Un
/y3yn0dfNr2smhWZfsZzqg9yBcW8yf429SRp4QPBy8F9gXOBPrnijr9mTgeSP+Ol
HdsOe798Gi8LRyACiM3NzgA5t0H3TH30S84aI8u/Q2gscMC4zl2wsBOFxO6UHE77
ip1MIPTCc1UWHJYF8ywJv0X2AP92lTl1PB2fJsQhKRi2U9TVskEZaK6CqjLS3Wna
XBCAeW25Bkmb4WauiELF8LwnmSGCGs/IioBIIy6itiwFWWcfc9o9QxthVUpi6mUo
5wK14eGJKQCjUaVmv+GrQNgJnzBbe1aA8RwvhQPNoB/bpDeRt/9er4EvhFg2Bi5s
2Juvo7aWFUiJnvCRGPm0JyrH8dyzNyr/G9rPo2OFRFz7V1y+N8dKtYVkPxH0Tlge
Sjmb+hZOok/TSgLjyZp6nHpZ0Z/oMhjzpeAOu89wmn+Ws37NaOehUHgm+eigJPSp
NdZCzwHTf4vUgBW1F/woxAK9H0RzIZHSbXxyPOZ63htTrJ/kQ36bojN4kHrjocLF
lRoPKFH3f8TVlVBWMiZCSwDdc6fG91c0p5M/K4+d7zi+H/7LjEX37GbAWOx0n1c8
FRi8mZ3WoC4EUSPjVjf+CwyzayCE/SJzUvDud4SbVomp0Gqtdgk73DWSyfJlUH+y
S8sq7qWRsWsN0iteoCGEnToauqMiFrS57aAd/ZKEAX6l+7EBb3dSijyFtaBPQZxh
q81eNQndiuwHrhAOw7EmxVgmYLJNS1AJ88E6XEW6oIZ7HYee+64yfNsgK3auEU81
XoHbTIvPZ/WZauTAT6xtfd5B4L3hjV+3H+SF4846u5K0M9o+Tv2Dt7DEDG1xsIqz
jIlyYSuURahlyutx/faw54joxEwHsqokTHrBjx9AnxqYpye3p/pXwl/HIukVNwXc
/Dz072DpTAbD5vOMjVE9hClc6C9M4qGKxHUdvKmFfPmrS4cZ7HDegGCDBfgf4QSi
XdvHoivkplP0AjOT+Z6dOvJ6pa/ReHS4JzDR3L/MC6MwGgNQvysX9BaQcvc7n1rH
uHPIJ+kmiQ3DackvfoD3pDTcZNBYtc6p0RUDO6X0zBCnbnhZvqtpgngAmgocDmNm
kiPNxwgquiE+dFb62CBUKYn7jfauvpusQX4q0uKvQ6kFNAtTGlfNo3joeRwsIKom
6hmilIeHIqfcDArXiPcaqxO0sKphCXC14y38riKoXxn4Wnp+ZNFRGhZjpw8QIoG2
UvFlGTZQ5/2G6YGOiWw5RWAtBFxBTGSGvrlTd7h5Oj02q/84AioW38SzHgOmxkz7
ik9AumE9RFvPcP3JTj9PIM3NkHOQhGNGJFmnIVZ3BHFbs7heV/joZGrsR/XJHBwD
t00yewgK2goU+mNgSQPQqV+CJDRrl/H43cmMZ0ZSXjWdhtdo/K1Tb8wtCuRC4LKS
I6xYw2bN99a2e6wJMfbn4wrE/lcU2xW3xAy8XPujJ4wEv2t8qNZE8/Vfsx4m5J6b
vTUst461Id3PtrDd9uSlyNC+37jyreEj/nhdfH9gWMTgpcn5LWWEM3UASgt+l9nn
CCryrpG3vPoUgZizF24oHQ==
`protect END_PROTECTED
