`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgJnRXss4Hh00yb5QTFljrHO/J2SB3e6D10cQeM0y0Vt9MH1i5TjC68UO3vN02Q6
7n7pRrRvayf/C2rYsCayVWIP6Q0iXZNQkvdSCsm1N9KqiX+8Ju4P9Pc2OESJHe5N
yHNNpWWY00xGTVKpqJt8LIJ9FFmnkVTX18KJbHOiPmZXXpNA6Iu+zH7IjeiE0XTL
W67/yVbnsLLkgW2nicVt8eI1Wa8S4CX830UGyOShlbxzFS1v7z7pOVbxCk8lMC2U
Ky73NNNF3eeTUlF+cz0I/Yim9QWKRjAoOcq7q/bQFKk3+W+hg/pY65vzVFnlmbNy
C0Dp5Fy+MEGPk22TJWFZ97I5XK1uXISh4rAQ2zlKLMGQheFM2DhVfiBUWMGQvXAK
oUF1zEMlBfCbHxDt7wpmPFgPJO0D0wnWXWnwCtkY1KS0rFyJQPvn8EpTydgFR3jd
H7RA93yWIBIZGal20Byqkby+g33nn/HOAzMBwqPxkHezz1sCnXCbJ3yvydmu+5PJ
wGdJptsI5Ozxekr21+7PQspILVFtcMaJtFjirNfhfXQM5pa6W8XlPhoihw5DS/N1
ui5SvcLKiYOYjEfKCRa3dpPKQhhOWcSIYkwNe+xuq7SgvBXzz36aQvuew+I4Qa4Q
B818df5KoF3pnMAl9DaVRjFLq/jZ/b+pUH/27e924EN1Us7svcYEnQg5HTxaYsIv
7aLwZqXm0rPVDoKlPiIqwsbWvSLqudG58jPYf7wcDmgIV3h6RoGlPEInvfLmqOW0
GRPRIkLbVa9k7D/lnbNH0qEkawhD289jxoTwso2rVwPGz9wk71/gZPS7xPSlFMjx
LWbb2NXZb8NjysDX11NxSQFfYr6wOcnhaS1HyfLCYVgIXpczmacBU/fQxsgdlG9V
QAXzmeaiS9gk/VOF4UUeUwnm520DKm6+Prmf62XeA67nXWA+jEB9+DnkKPfw1du6
DgmVjxHZRu0ofBkQeMXZhnW2YhcvO1W2/TnKVHhJGiedbW4hzSwE9XTGr8zWLCZm
QHVgtKpEJ02+EpYddCfNgRYZAHolBK10JCQhCwWv3PLWiYZMzVYeptvKtYYH5Q9t
uWDCnVrhQjirsLMuIHG7/8Pe4EZ4YV1HNJ/A8+Hm9LsOf8e0DP974ST9yza69JmB
QVePfYRfJoq6CJyg3szxCNT6mazga3NBm+MhiqemQTk5mKBDNOVg2KDTIaZRPlWW
cisjJbJHjE/qZ0eMdVz+R5dU/4CTZamTb3SxIy9lF2CBfvOgcB8uzVvBVa++pet2
t6gJKIixTkCkaHTEBf+GNrPRROr9XzXOTTZDpIGEUFOfdfyfohHevRDMqpC+ywoG
8EbkIbIz14hWEHJ3Fm+FoXoE4NWHhMoVtwbURpsReBTEqqqRMwu7t5Xk/4J7Y0tX
18AdOqGNkQBVe/Tq+biOc7SQFDE3y+1jNkAYjmQkvhthA6imcTrjaYZLuvse8f2F
pAADkcGK+mJtY3nz7Kjc+slO+esO/JrA9jRLzaViqSK0Jrf+irRtlYusrTDJfn+j
otiQlJBBiGD1nxwSwpBVsT6Yp4K25w9CVQzsg4Ie82DXmDQFhO45QHAQd/DL0Huh
qs09Elxqom9Vs7Tl9XHDeWymVoobygVbU9fOCKlCH+FO2m4kzspzWnJjDofHMLSS
lJNA7bmNzcU+QgX5XYOjz6qjYsLcxl0VEjsmZvlDGIoeB0DaaB8aFkINqh75rTpD
Kz1JnLhXZcQJqc2lUv7GGS6/G9hjqyszyHVX2tvaFGdnc3zPf7WYvzyNFsCBdxIr
Mgdy1/SiJDFS5IPCbI9YtRLITTXY7xWxrdopdPytqbptgWi0rL85XyGfuyU7NQGd
oSjVTQNAblYDM9UneVrSncg53kjewFWN9PL/5yKCVmkrjP0y9gBmclEsrCmpuJxA
PZNW3SNkKqzEirY524GFZunj8CnWdYVgS9EEXKaRre1iHfBiv1KlBesI07jMyLOC
DKxhVFxuZF2wgftxIdkA/lnPGT4NSp3SX7UpIy3aS1LOBX/kTyffeyrMK1cB3Owa
65CPk6xkqavDFBnqiegBHA6g1WLjMhDXh3UNDt0OI9iLarm4W3Ffa25ah8vl6p/o
tOtdMHjRi0rdr06irf0JBMyrwIHqaiopbuGPdtC/zr6hlRy3h1RcFmaYbHZgubIV
5gbpJtRP0UwCstDM2iE7Bgnp36dtq5kfAmwPcpfDDQZhWPk/Bium6MwU0wOrkInQ
JGLQgwPg9SC690SVA0dAFUhA1xhaGu/YDsU3lDjYsoPslFKcRNDzE5+8bmzrDkhK
WK4vLLMAYh97bNVOiAq7j4NX9428VCJ/5OeZ8wtJ6E3gkODjf74ff31hmljhvbin
YA6g9Y4GZE36hlwjiVai9Ezde5DsMgMbDvCuCMoWrWtJyRzoO3ErqAz66n1bTDYL
m1nFtD4JM/lzyYh0n7NeVJGhrEy/w2nw4iRDPlyZkbG4w8WnEeiXyY5gnXrLqjIS
s0uRI3SeVKM06tLTbErJ3qf+nwJEoMK59qzzL6SG8P0h1X5w/HYV2Jv/ABcFSAe8
3wVQwc1hD8LaDdX09eJN3LWHMKoPA4VozuY2v7Ktpc4jVIVo9qGSDy425LtiGf9k
f9FAFndzytKyAC50MzqkN5CnIIjF5CYbjYZWA2qdOvp3Ch+tFuwbTdHP8Oupu9dJ
TREVdkOcOypmbcu7fZpHomgaNG65kNuSbPbjNcqDeswg2WIBHbggx44kLpNGTWs0
nqg9ZRN5YUSPigf3yOC6vUeyXKXvJrNv+XOgtwXd+jEShT6NKWqF2qu/JeM0o7Q/
hn+H2iQuMONEJga26MqVQAcrGBY5svUV/aeiEseOmdzmY8rP3lBaOo39Ori45x6D
IoRbdpvUcTibJfYJCcMXjXspOc94nfH0dkZXEjSY9rufMS86mxDdxCONpe/qgrCW
qw9qvzmITU8FvL981IQxoryoJKzew0gB/TZMcPOot3WygnYb7g1cS71vawEZXqHE
2ilmuzVOZI+TV+yYIeQ1DJOVUlOxh8LnOG8XWfJehnd+BQhgKBLtib8h3alFnOHE
aHjgj+e8kh9IS6i/QN2h9e9FXkHcRPAaTPym7FxKdFcUFbRvg4nNCcPtl1rZ0BXv
V+v+tX8yFV96Bp4FC9tUnxtCUPR2g8Y+BQQc42o8tAa4Ek+S7M/oA/dunytHusw4
UAKpoq3OMQx3eAGkOj6wWtiB+Hp1gi17tspQoslVRWUvm/KuJKrxCBn3D6fTk3jV
NztxpC91x+xmyUInxtVRv9DMs+trqLLRDtKZfP8O0u8KPmyvxT6EKMaDrugu5Yzo
h9bYsLRHGXsav4yHf/jAp4uZhPgv1TadzQOarpDLNSTkAb2kCiDnJNOZwcXuKqhZ
qMB/weDWM9FM1w+0sAq/pRKoDCLLRgr83odHqjxNlmtAtSsD4BP0fTsV0h9vIGYS
ptWT/Z20hPSjwXcy3V1m7oxTPUfifEZhyXsbAhrd3DoQ/ebPqIlBh5IMh1a6pj2J
3N/NboO6OPzD2Q8c7s0vMlwKsR+zBCUzGCuToeOkqTxRh9kK1IscEMZQdr20l8Dz
IuZJFjo5iqxudIhqlBgkvFTklftR+inzoWqFfQUDJayhoaOSrdMXqj/W6Ztht45r
Cn3u3/Ik/o0+oTQiJK1HoI/elABeTsOQ18UCdI/v+8qfADFYAB9/DLwp6su1mn1c
Xq6LpEsZ2qj5Art8LbDph5NAhbygNvBGl75gOTFugdTMxF25b887Tnqqs3+yzzj4
xx3lQY5XJ5ILBK0JvWuZ4Tx0+V9fOkIVebt09oAa/taCAuYnlUCEsnj+bSZVAcLq
/2E7o09XoYdF1nUsKfFoIh5Lo0BZmaYCj54rJUAbShz1U8GJNWTKH1BEyR49Lg4d
FCFL8GTeuq+qGi7Q3TedsQsUsUbqS8agZab9ZUkDSaj80ehcvr+HKha62poFRSzI
qwIq7gIhxcAfxOgUt5FH0BrKXja2PkepgYV00p6tCkSIlr5472mQxN1x8zX4rgtn
k5+BkVU45Wt1V6Tp0lN2Xh9gULQEra3mYx0oGFCtL1BRSkYJmarMCFLk0zlPH61m
Si9694xITHHu5JqKCMoNykyNSuMfiaVUEOugqtwNw6EL/WcwQjg7hwI/uU2Ihg/Q
RWodxBREM9BLtzPpraPTmcG1/h1yR5Exo/7nVAdD+cwN0OVO51gAttzUKQdWIl4y
eQ0d0Ds7RTxRIbCuTv+ehrJCyrQEKNoh8cNxhBR+XWjPbCcKHZQFD4p6P8WH5HI0
TBQwgbn3qO5IDs5jYm3uhCeRajzDN/QF7CDSQGlHoH3BGd7kuqkGlObEnOiAS8F6
P8SUr0W4+ZgxtT9LyhYpUmrUw+cW+geeIvOXa8si4pJp3ZDsljmNlV9oDpWQsWZB
3HuKq+h/UvOr2QeofwEA4zzC6g4cVmOvyI5n0GLBwAtfxXj5WORo8KfSaU3ReV/h
r9sbI/vDG814dY2NwnnBFvuKmlKzRN0IZNqdktERHxqp3Q+iHd4FHFprOdjCvizq
JXQ4sCjbMfciogwZYw321A+JeJJqxEp6lkwd/r+4rYfvHk4HK2kEbbTa4DOGFeJm
xiCIv7tDOTTc49GBBl5EFEvpmVkClyaU+yZajouhJslThMO0jyTIymdW6O/pR7/T
xepxqdHDiXzsFIGTGn7v4Dn2J5/xDxyZNYMS7F7+v7rB0fxo1t+IMJYeqyCManTX
6lVl4vVNY8pjXkOXJrBamVUtGYwSjU2r+gBZ/VD4RDWXHA6D+XDIGyD7cT0MhLh4
scqHd07sqZKNPWdigBYgJ1frqmiPjDAnPFfVos87jkUBGWPRBEG1lvKuJQvgY49k
U20uJKG0mhB/E0piSsj8gCL3/GcNEvd71mpgG3gLWHXR1XcRK8/5Bv1slqIUc1TA
1ykmMQ5ljtusMUlqm7qVPl1NCVREus0cBw1KUZ7Pmp2VaWZW+62TH0xaj1X4gIq0
bosHbUSvmOGmoJ6TrptQAibuAQTpiQdIjWQPp1jcSrgGZ3ZVwx10GCSUKlG3X52z
1UayGw0+jviV+4Qx5jc2/e3vtnjlmpNscJOe22+omiU0wFtPMHZinAXIBkpBXK70
E1Ll/N5fA9gGuS8f/SF1OlC/8+QL1emj/CoaE6ZtuTfQKPnIYuvDzpIaQGDZQuE0
3/eOO8VyorATte5EdBQi55vlQJBJmPpu/zPcNZfri96M46aZ7dJOpH4y1btEQcJ0
MgamKncMh34fkrj3O5OyyhdMsvXjGlX/e/LVAHaTYkEkjnFIpMRuiVB+xwBNCXrh
sMlbcbxGltLvlbLrvQ8glxe3jk393/7r/QqrVWUno2GFbi04RHEUOxPvaMT8AOLG
st0L1kvun8yGl36nyUCvmmfFnv2YK4tONW7uUBVgGUn2vGTTjmAey7CxlYl7Drwk
2KLKw7xY5jv5nf+rgbp3j/QhEViinVb2Id3l2toVwGBn4+RIZhLwEKOjxi3LKiXM
lw2N9wVKKrfZclimXSH56Jd2BpmJNbRE3ug8b5jGU+BpGvctSkM1hVfH8wpNdfUP
40QUMxm2wo3K0boxeKnBxy8HcLss8wjiAcZQzEsJBhxeCs9o2PrAMTP3cLOfYBYD
H5mKcqXuuzN7A3ZBaiMshmL+NrYbwUG05U4ta0B4d0JIeJz7d8XVeVZxBJ+/hlaR
yHvO/OrkyuoBpUJWwe4WU6X4ZXGEv49uxFKDmDjG46UihrDLBgy9GZ/k4+gxhlsZ
TIWnM9jpFHq1g5EAM6minexI56ywvZKTi+z8x8+pT0kHhr6Eub2OLlCkM3pIUBw1
1Xos0DCOCzrPtQ7gDRv7dgYsCAT41XmAXGCgxp6IbaWKA8GH2Y/kI/s0rhheNmOH
4iW7JNqD5ZPZ0gdTrnTPP/KqkFqE6xnYyCbK86csNkDucZ1a9MGz3Om8wycTaWNM
2NcXOIh5fc/DvTJmIg5+WpzrkFYD8jbnBFIxB1y4Tbbkymvwobtr1aTrj3CeeIic
kj/r8zpaUhPEBI/TbcrH/PCCAjxbgtPWwL4/r0UtCAxWFfTPxw5/FU8XaflQnjpH
l03tKsSL9MnpR3LfYZx9ymwfbUEfIxVWe+au6KqvJBY9d4+Fv7GqCAKU93Vz4Pz2
BTZdg+hpArXe8fkeDg+E+oiD2z+1bXU3JjSj8OHpOrIYBMKuSgRJoYt3GzwpTcff
6Q/XV0y80z3gjVoT7rwo3b9F8ZtUURX6G5jMbzp2hTkfVEclmafKOSZHpFwO3KgA
Vaqx5+Y4e1VLHcjK5W7U6nbXL7zL1cfXdYkE4Q61/vFG3hx4goeD4YyuVRuQ4FuI
bGxQtGydTNSih2PvQWZQZfEan/ug7uUmmqusSGdk36l9fshmlk3aEeNhlbcdmX1e
wnE06sShXwORrHwXwUqbBrEscbthZfIbgXFdERT01ESjgUzQzY5sKfg89XajmCoj
rXKE52aDrCPeKeJfOVAp+8wcaOwOO/XUQO4HbXOKCBvVHMzD4S2jJc1EVGXj5ZJs
JMD3faFxa7BSVy9F6Kt1oYrFQz5+OwkDDUwcbGDapjuH2dPU1tvxZ6yS106MNL1y
wB88uL6QifZGIKPpP6CEnREwjXEsBeIYn8k0xhNMsMVG0FWXWUQQxrJ1Qn+c//QL
nZ3QOQ3Nv8Ibm4ewnovb1CnaEZnM9/JR4zhB4vBVelR3/67lYu6z02pGHPK/9xRo
Kqf/aGvVArCmpsLWUTYZqao5Fm4o5BBrINHGFKZiTRQaQCpJK+z2Bp0OwZ0xnHcR
PBQ4O2JQg0e4siEZmFYDmU9LErZiWeA1blk+3rmUn5Z2RBxNU6EkQ2to5ZsIlNOH
GFRCKh3AFE5IpcwpC9dj8IjBxkTx5VAVR9EdGRAXojexc0gKlNVtRUsg0JK147Ev
7W6ZAo9gSkNUrf9zWT+3yNrmZdM9mZrn1ooH6SNrVabSSJuD7TODR6WyWR75RdJw
aedtufqTfke+Rho6Af+27HllNqOfUiNNxRooxeEhmD1PnL4IYuhy/jrRd5gMYh1F
hf65nzv4HdXOePraDyRnLKgKafYUrNXV3vjN13wtzS1zE0MQbDveIDrxj4dtQSm2
vt4td8ai0S2eqRDHNvh9GUfJKtPyCAOYqwvH7RN9r7P+0gWvF6vziWMJJbriNQlE
scB/f+BK76SeZT03GHgjpsBX0miyIrORHPoVfD7JpRBFl3KaSus0vH0hv7PLabBE
UbybHDVtKq2/n3spBSj1jjntjhxAV3iWUpVldX+ZQ2udKi17+q98xWUETZRmSW3w
l8r252RFxIE660SvUE6/aSk2p36PojkmXIy1EjCvfJev8GNMNi6/SDLKRPtVfxYD
QzXJDsaD8Lh9jFBPz1UEMUxGvv7acVnmFch0G4zXhhVVvgDjTeHKH5cd0dHmTGj2
IztUU2fHouxb52qrhMFqCFXPJKAyqas3nE8sAJYbM8q28fIZf22O62ZbTGKRTEbw
dOi7GdwCJzcagdGTZuy23bjLNyeuucOSZ7zHDJXX2u+2kLYujH7enPXgj8p0ECpC
wOcfS3m++8EYkNASDnUVTDSK665ewhckco4++6QL0narfASg8qJ3fWgjp9PLsKEF
k3dObhqBd4koR7QAyWfnDBbwRw4lH1bp4mYH6/JX2hY13F/IoPb6uiLUw4+mbTHv
7Pt7VLuSiMY1k9Mw6GB7IZjJC3wGhi9jYO/yaQMPgdX8uYQy+M5hlIvNuNJyyLsk
0gPkVgMR3XIJBKCfMGGI4uZLlk2hDXJqjA8RB+VdRo4EnMrIaWBzxsblLDA1L2Vu
7TxSbRbUFFO8IoIA957WC/R7i5B+yhVVcKfnlJy+rFRD6EFs4CE4gJRFOSoMvaoO
7E0x74eg4AkeD7T+2PV0bIp6DaDana88CkzSNc0ubyB6VmiK2I/ytdyrnwYPB2A8
s1dxLHK2OrxJXX2i5Rox4pfiovO1NK9WoQqhbZ71bvD2RoiZYmV5z8Mo9Ozu4TyC
ZP0RIsGQ1FaElLjY7yDl54uSTyvTMZjQV6ixYnDtTrtMtISOaal86ej5crMaFja2
hEt7x+ZMrZg9xzYj64/UGexaDwEIy4bbDTl2y5JI+VyQiQozHEGlUyFwSQFuYYUr
UcHvTDV8YQ+WoNbn917a8CU+/Bs6FgobVINMB306deu/so5aAtBNbZ65U3hB1UIU
QuLG3RgXap94/V40uQuV0d2qNvqkvufaL6JOod1zIW3p3+RXz6m3RlcUozaaWB/z
hWjFwIfZq5hS/qBe0I+PMG7n42r9cH08Qvh/bSP599tQzky2cM49R16ceS0OOh60
CSgPhuRSaXXcH73DI5Nc91msu1WuqYSdK2Mjf9vPjQcimWmO+Bzv/Ly55sXA0xak
eRcUcXeA9UCCGWeosIGLV+NIAiLarhfMqWxpP/W0KYnZyHE1hMJGjalQgcPluQsv
/b4Cvn7ca/XEvrK2dWT5p13CQJLkZgqeyzLG65qJw6jCpVBhqjHOJwWUjhTuPTwr
fCa2+hJfY7Qu6yfiYm87vmdAyQBM9u3+JyT2HyIfBSdNzI8j//OL5+FD5QzF9F0o
2sdVuaR0ATudxYlNMxU5mFoAtKpfeFk7se7AC6QJJIPbfAsXNIT6FyeLEmerzZ6q
2nLCoI1e6wx/dvr2L9Nc5nHJisW9QkpjJQrRDX3cpMRJCSd5k1i2He6tNfbwCl5z
yCcGVcla3x4gYHctzV5qW+8FqIjd9zjAVxYIiGe1orkRBzbrYRyJgyybSNaud/y7
31mwrNJCGeGlXCfp6mj30kwuihN7zQilzVIvgIqR3K4fEYZKxWelP6t4EvEJSE6k
NSDTFJBBF0z3Zwz6IMHSIWFtCtWWVQRPGQUkCK9Rbn6MO1MCIrt6geJzv3Ze1eYz
gZqDRdot88mZAY5C5tZSI7JMwK/iBBAA6j77YJoxtsQHnd2q4elYF7SsMVd0hRyy
9JjMuzbNRimgNsW0G/GtcE5B6xOj8Sf1kmC3nGW/kVA1Bk30iolqnTMBKDD7NLWa
nO+3Tc42CkhePmuSE3pPhCs3ROj11j+Q/UzT4UxiuWUk6Y+8u9ahrXGu4AbdzRIS
/Fv/KY1niNpa5Df2Rx6+r2ScbJ2hXMBQiVdt4PN7jEd7nfhxxn7V+N4YtIo2e/nl
aSNrJgeomrCQ9XKcIK/9KySmJNNG4WhjFmejYfiHfKbwToN78VU0xAH6I0ct56zl
n8syV2yllQVAudqSalLz6s6hZWMXa8sAxa/YmwGA3hVAr6SmvvCi48j1fiGbS3Cp
V6YVpJBADEccM5LibO1RwMNKwj4KwVeZFdGNFRNiwZtBW0niWns8m8qVPu3KhVBl
G706yd4it8KCMp32jLEDo3x6xDprlt2n8v71CzACIRAvYe/t0g0rPDgDX78hhA1k
lG8frXlRl7KpZQIUgZr/AEMtF1CmhS2WaTfG7TLBPrBJGS5NKMUuGs5qaMil3XTq
lnRqdjXmqu96HYDZv74rTUmvCYX65/EO5OlWGF+WkERD1lFq6tzfbA3SNMUF6fHU
hv18Rs9UqeDbTFm658aXCm0rArZKRQ9biVTI24skNVbZl4zkrjxlIvnX9zv3vdSS
W1sphOY8E/nJJgpNa3GBhFfRaarSBKS+RngYmssfxiviKHlEmUllXgzgGHZCScBr
Rdqv083cgP80NzmqxFAnYxTwK8thZgqZwzCzp4si/zp375Mi6lEzjH8jGRXJ/Ci4
hQxB06P/jJwmjPYepW3CKu5uLP8aNV9HsL8SaIOR/litujwbfoXk5D9lBSc73l4s
RjStzu/Dq2r39iGFMVJTgJqx4Wi5s+C2DAZ9LRTEYb30YZPLT3jxVx2S8WTAgW8S
77fbztlruLLguVGWs1ExN6pm2PyXfdrSHxHVPT7X3dTF35B/axFnnk7m838YnUnI
TwHGs8azSxEbBPUk9ldeHKzQxp3H7khcn5uaduuO0X2gRnF5QjP/CIn9P2voOfUi
8tXYOHfoIsKVT7RUpEayR2Am6fH3961r+euERjA0kzF6jWpMBGhIRmvubMfBJocs
q8gAxAOULzy8GudL1dkiMTwQU1CiJ8EWGlipVUKb+5wFjk8VPOXR5hr1eg4LvRDH
vEsJWXr90/cJWEfaOz8dsrVaDK52j/pptUau3JMIoOWuQiYhQyaPR11+els96xhl
B5o7fmNbGZxFwb1YBK6Wnx6Fy2+Xcm9t+oil3bSJukozG1/DvmuyWVxIn0d8iA09
5c+JeHT2pgDxncv5PVvbcRBRRlMAMvpfbvvUJFnh8uM+/XqJbhROiG6RRIOTjhPD
QTlUFuqPB/NeKHOOiOHvS64d3TDN+CviMCLy3FlSByZKGw50jnzblX72JTQXq+c3
rpbutrd8Fvz//auCEDN6hquECarbbLvPm0LKoryhea5aMQfH8qZ7bniX/d/k9gnL
7qtok9L1B4r5vVQO7BjjWxYwCQU0ODrIFHvakiYQ5IjJckCTKkbGfV/JetXYgHKf
VOGgD2NecSjm4fTSL/+oktd2FPScwD1gcDKxHOIsKl9wm7mIfEkNvCcqo3sx3gWt
GNYWHxyQcoh8y7G0IfI5V7481CqqakJ+KSa7W3p7vl2R5cpW1Np2wT7JsR7g43rb
wWpbc3/3J86WRvX79JZxBXu/H++1wrYGEPbkMdBeaweoBlemGd7J4qQp1Z3Qp6lc
Nf+95UXIZZlBb/WztWjrU0hfatv6hxjMHNmOBlgWN4Jl4tt98Us69nRglxsu81HD
qcQaVeSCXIzxy4QupwBSH57PDlbuvdI9vbPVjShRbzbEzg20y5s6hMnuSlwT4CPf
DJXX/GhTcEWlxCVeM9ySdMTb4Ic1+lf7DQLeC3J5AGvtZaTq6vt7jAL6ZZF/Nby4
73NQYKNbvwR82YT7hCM875KB1Vv93hsAGR9JO0vXTaZ5KYV/iZlxo9Naa3xe+ehT
b2dIbZVR3oPlMjdcIT02Z9q9QfuqpZq5I7NGEH+66Jd4TYrVdvedWa/wh7GFhG/Z
38NMDg1wM7Ksb5vxdnUwWDz6VcppEz2fdc0afEncaHgQAxcsrxkyUiuf2XLcI55f
UBuowsJOfAd6BvC07fPqa6hMjBks/uvR87q0crknenhR236rkiUYN1avS5J0vgaR
Xdb0SN2AjezR5peZEySa99TOUnm3zehxkJ5b5cSmoTMKVYe+jfKXbcTlUGylJ3zx
bTST4JnzmvRlMWX3QBcZB/obwf03JecuIlGCFJFQ3lVSWheg1xGoQG18GbkATT3t
USrskwU2lfWPTL2gztltKu7tl1FQrUB97eEs/HyIBQcD2SLQJ1N729pqxkcjH319
4/PQ7SriZKP681v0IXH+BLBJ3rZjJYQf8aM4M6NwNDkUTTfECKMLMl26wwuoXdFx
DDx6vxSSJZStsC9bOlG0cjuUrXWWkTzJGxlAOtmU6UwGSX7YBePA5jWVF/axdEFf
SrkAeGgol+CXFxt1P08TEbxYx8yYvWmNwIAMxaanlXDhskXT8WALCGfvhAsIWk1m
Uyp/2Nd/P4VEAn9OENcgSRlUeesfrkx1JCGFxk64Dth6KFNLqNe036OQSVrcTvCZ
oF8vdNEWEnV1F9MOG/tdN/I803GVG56ht1AG7z33/QZJ03QeGs+lmHEhKwzTFVme
alz6mIl3jH1aY6lEkEjLydytfAf7zTqIpFRDVueqp9QQXToQV52qu2sDM76wqUrV
mPFApyCJYOQp8vQl7K14YG2ZMvsNhmBqskJOHvMF+mBdD1f/oMplVpenSuHZl3g/
pZ+g2Y+GyzhUGpAgxq+hr8tK5VL0DMIiasYgydmObCcZRicICncvz5nnoemnkC6q
93+WoHu02bmMXO5h6HmaGDCcXNhhEmrQUnbiHqLKSTyJekkCaTz1oRTMIPCQiCx9
8YTIvMiEPulw/st5E3hnW8A8rmO5Eqx04GBVSL5mEclcoREJiNHEXBkM0TmfScLp
CQ2bzTOxZ8ODkVF34l2oivh+eyaNR4mnrxWrzj+d/7lAh7yLwHFgOgDrAiHUvZsz
wqY2SKAXn3+AOJZ63EfNVPbIlyvwd/ccmgHxzsc+sVhDE8QE4DF8WPdrclIKTid+
ugmQWvDAxyn6FjkmX8PxAmS+V9BvokPPLrivGSTSHdDgS2pTkEK3X1aLy4VsMOoT
I/uUMF8pQszFil0VMS2MzwA09zI7qpLLp+hpkOtHUIiz1Sn7VM1LqASnVpHewBEC
YQri8RU4E08wLu1m2VUrIZ2wiCR0GgOAtJkmpVfLLzEKJ1hzenI7DJuglpOtQRF9
CxBlKI8oVaDf+TnDVzdqxZrQsXQwrZx7+lIz/HNld0gas6iOWWA2JK0d5QcZIlgk
4y88O9NlpoLiR0jTFv23uXHwTxzOJ59KuNtdJqdIeK7CDX2Kc4jCH+PZgaSMWEZ/
PXj5F8HrdnsnOOBNRhq08IY3zFACg9SMBxmC97B4W+xaZLT99tvi3q4Q/NcmG0JP
/rtunbKxKb0Ulk9zc9RkB62Y1ZbmiU8cz/JVtv+ZJmFYB7RRGtB8gjKjUfr1Og97
0QpFwAMPF7IUz5frD0ZaPh1v3bZShEFVT1mDNS0JIlkwwsyD7YwjB3frxy6A+yGj
slNRJDRYQgWMfTkWsinlsqLstdos3gUlGfgiIs1gqjBqxJyzW8hnePJVjEMLHbbt
yudAWtfEcEFmxwN+8YqdnmmeU7p9985tauVuE9k8crxEogSK95BjJGQVR9Wjv20Y
JT6TatKfdpHJKTWbccGDWThqKoHBIdZ0gGzIJWMOMIbV3sXGhfcj9DlJnzZV8jBs
pmmUtLIq59LKffbV603LuOrWg/gOmugFePj4uUhcf8EaFmbONaoCEyqCmsVT/S9W
ZnALaYvQrnRea7lSXkmGVE8OkYhzhSF+BZ/n8CT88dnSiTzjkUjVd5BPwVn5efHg
68RwMFHAo/0iumdhs88oOMm5SYkmExHRGOflFMPSk8xD3md+t3G7zmxDFBJwXR5i
ObFuHBeK04671KxmHN3JjU8kQlvdPPY3PI3qZXLZObbz6TGiM+IMK9gOl+UwuMgM
3YFz4Gm/UaVVRbONP5eZ9Slc4yejI1dvMLcgPOQ/hNYEWzAjXnxGu4yr5JSWb/Ul
MS6XySiXEIi6TPMKIa87mKpykYmhqesy6E+2thXNUXqHO9oI8kVuutDwFDzpUdJO
EcImEsZMqeHNdihga43uEKmZDNj4LZruSmE/rXGyEEKak/uEstdBbv+WqMmqlGe+
ttoyzemIsE0CTbAnVp8TEFSH0CoKWVgZ171sRdAuKRIadTkULb/ywZ9HQ7Jvdxcu
D4pvuIpGxozXF961rCK+W/OJa1akrjIBuWmNuxKD8zgGAb5ufDVBX5F4HTbT4xPQ
IDOb8MhYAiIh9xao6esH1SUBh3pONWlV4QNRL62eucxS1u43xquC46e42lZ8o45o
2n/hVtxCsZQ70ho7BBSeVJPyjgOAxr4G12t6gjVhZGnJvX87cTNWWOe8pwwRRf4o
qTJzA4PO/9zETPzJxIxxYUBh/iCXdj0WQJ7qjl/AXDYNS8oCXLhMhtAhD1bvmJvD
dUi5RJcWAjKFKVqA23H7sT9G+duqjTwmMfBHXKSs35fsto4E9nkzV47vYU8UFehi
RloT0fDqDVQaQjOwzYFnY4K5lv2SvczVmoPZfW3Itf94DnhtImxr9ocBuqFYhviE
NJP6wDkwHMv6qgZ7psg+zdsVgSLU8vtQgt8sZ6J5wZZrgPnb0yP1t7oPZjFyCf0/
kjeWLOEHJe+2Z3sxBev7GkbgqyW+cWW3HYOzLKCVqzMOKZ55VuSTaIJJPe1vXKNe
5Hc+aq7UpNvUPBkSBg8XnCb0QTfRB3kTolNOnjtV30S2jwqLc15r14uEmcIdnZxJ
AvNeaxYBilaOymVz/flQVECIY+sU6a5XHt0+YFuwvoJuS40ojo3gMHJf6f+E/hyV
+C3+AL6GQ607ayjuW5dAKc56Jez9WCknCg7WkqBOV4fnNUvcTRz/vfQtA+rtHvjG
yfYbiKJKUrPXOpNxGUJb2NWXiaUVel+Ay7ZOjB7goFFb7Jx9k4gLsrYdCCyxk2Dc
YbxHfKRYNH6bWmT5XXTTjzEUbODLk2krCyLUL4kFtKbDETld51SECUc9pb8Vdkov
x+SVinbp9L8aC3XAQX6zmY60REWq1KcocsjNvwxoN+7NNhALherOw0RKLV52Ewjv
h1S8FiFzUwbTDwP4pWXWinQFsH4BE8j8zKS9Y7sQAlt64Qwe1J6oTxt/F5gRTFaB
k7t5nyl9Rq9cT1OVVJykPyQN9UJntjCFgS34HqV9L609qXihnwNWHLaEuTGUHUnB
K/3zfsQUV3sYtg+qZ4uf725eUBxF6+J1G2RZulbkQpKnySu4gKnJhDrLyC2rC8ZV
+6pi1l3cSb1qfEOh62Xkm064WMST0623nL/lQZsKdJsBnEPoci7ajl3PpA8ekFbC
azV59oVjyFrv03o6ZB4ObhUUNKpF43HCUuoognidtxC1NFYQjyKadqbIH1gryIpe
i4sPU180/lQY7T+TelZyo/zXfzteaTsWEVHhx7Onj/oOM5Ap2bsJA6Koq+r4+DCn
S4dM0b//HamUpZPpzJ4T4N77/kOuYagaGgV4CBzc/29WYzQfIqgS3EcB6JnFRL1x
XkEfFCcwrA6/n91JRxujI1HM3KFMKqiYIDpyVokC2eN65/yuWBRLiRcUr1zczNxQ
JBNaIneWKyAwkHbKP9fhXENuJpQNbuJqfBrjiYFl8aL8T87mEjukGjqvkBapvPyH
V6CGMFmO3A/Z+JJykzcsuvImyyWJR/UkNCdVFvqw1zJyd/ymzH/R7KFScFttpac4
dQFZxzoMCgqbCavGmD5zjewMNBhY2dfba3S51q7FdJmJoqRa9Uu8+1tEIOL+psL7
MuPSClR9A7Gf3iMuHftCn5JgFnViA6C9ha5fP0wyJludHL4fC9b4XuqmP5O0OZeX
523nj4pOWCFJ42TiUODk5rcKYy59gtcGk2ckHek557RCA20S4Lnb4pkcE8D139sB
XJpHBfhVgOumzK+P6T506hN6S4SogMbEguJFysAgrvXPHoGmDXag90bjHDRvKugO
xnQTvdBKLdVYmhqkREePxdcT7QZuWjga0oCXZtIt0DDzKjo4cx4VSwceXz0jdjNS
VhRx8wOfElh7p1KDzxmUWoXreLN1cBGlopYaamUb5f+aU9x0s7Vl0Mb95nhrLmyk
XiE2WqS8Ya6Dv99Uh5xqlsYW7SSl1nxpx/PtVO6iupnL7qoE6RoDqmXQIpwGT2dg
h3CeSLQcZvaA4HPKK1drbzQMXuN3kMZ52c/1tIO2QP/vavoNyq12wtZydaSIZ37e
9ktT3/LJjGgZ7lm9fAPYKLvAy4Gq+O/H8v2O7HEwwOqul8bQlKJSGLNnaFYoXJC3
5FbkuDx1YDLAxuburW+dNZhH9YokslQZe/tKSm5txClGQtrMgur7UB0G5bAbys3a
oXRKWD/+crztOiB5aSz+woZeuyXOLPFNn3JqgsIdnj/kX47uKwySt3Gx5DupYKRn
4AbxvD8590UBcfXSec8trQNIdrwJi9ueRjR9/EF8RA6qmUILU5T8bWtfYwAfgi6t
V+JSOTU2oQSbLBbdnnK5TEgaRx6yPvdnNumxWcGwj/118DNjfxGS1+Wa6Jb8LJxC
rPefLnGbLCQkQC07o3EzeC3PEJ99oOb1F+j4d7PqHAVky7O+9deAkhnWv0kwwINn
8Evb3Al0vNWKn0cvo1h0uSnsZyVeEtZkrM7ITyHSLG7hLEiZPgm1NvI3z/klI+7t
dEb/zm1oQyPn+WbpfedSswvh3iZ2E83AGEk3ck0U1wEoQTInxzJRasvKQw+VOMAx
9Yrga1gcHmsmHtRbg1x0Aew67zNRt19Ya/qfoeVTL2RPum7Aq1BW0sBK1DdVD5Rc
Jdk/RRQU4wxzm8tIGDnlLoJnCo7nUFasTUW9nMYO+UXBdN/dy47ig52CLonjh5+x
ex5kUn3tNxNYPthUVxDwjez4m3O88q8069pifsBAa5gkfSzKquAuQi5snPDo24Ql
xHHK7GQbctB/f/TVU9RgFK6y2DeVGsYlM5hSStwjZooo8xf/z7xGAMOaDlAp0PbM
bYFeA8X9GIHG+bAwhK7jprVsnDNpMrQPYQfNQ2wtedHfVixtbn+pKLuw3CMNYYdw
M3JD1GE/Gau+G6FCQAQHuJBfuT1nc5c8Z9wuVE7UKWBjmU/I7eIqz1vapLM8NzuI
+rxhNBAdO0FF+wAZS9FDSHe25N6Qiu5ZCFWSJEPxewEnaqNXtKap3PQ9Ve62L3kc
ddJliXnTdxGehrg/O0sFiLPa/23JnB5PTLid10sz8gpBYI9tN1FxllnD4YaK2VTB
E+M9siYuAyn7lwqI502WWiWot+qNa3jDK14iVOqhenB+WPd1Oq01tsyYIVpqST5Z
zl3jLK8Mts6O4NXfYCvbXoLjmBzKRMY19y4zPE9o4O+YGDAQyTfnGLvGkZq1FUWf
uHknA+TAv663oAxNMeyyNp/nv2Bzk0cs6yvFLfFQC7CZE0BJRvILIyYPMjXk/GsY
x7zFcgj4ktk4gj2HEr9HtLDksf7JIFX2U9kH3S7BZF0JVzqWTSbrRp9pnzC6MeG/
ajiH/1xj5WWLKpIKjPHH2S3DLqeF1HFmmqBVjV6SbaPc9+Em7v1rL1K2X57dKaT2
nTcUcFww4d5W48Us49ykX0W0IeSsXq/oD15DD6T5liDNM6jhW3Tc1wLvphYd9ZRi
FsLIwSIc4xW7DZVpq3xupXlQAAxyrPBawsghIL/uUEiqn32j5WCGdk1n130D+/Yg
Sq4f+wNYSVwMJw+19VmWIrGxilQ2WRZxWd6QCLy0/DbnUx7lY4sRFBSES2uOh+/4
PDm/mtCn3jTRsCPGua9Tak+lWAO1uGmCVbSVwHO2NQe2xWDJYHDG5WCU+IYS/xEQ
Vrty37keJcgBw547AWT6lI/vGDERiSG3dm7C+OBEwXbJgkeXLKQYR1T4bEKPfGnO
aurP0LL0fRoLHGPedZT/3ubIOD1EKzFxmj4mxIrmtLJLWb3kBq9zkkNPooy7kobY
wiaMLIp6cvix33xs0H1dAlHh/04jZw6LtDBEznHQytPElnNw1kkV1TfRWFkNd2wI
lJFCr7w9SJfAzS5ba2JPWi9vgGycVCLygnfpQnapqnc9OA9EFnL0mxROmGgKishU
lUFlhUaCpxbWyYh8D53PnHODxtwuftfs83iVdgoevhxN1WNiLgbU/SeqAJWqFyUO
Hl0kXfN6YqQ41e3UJK5MFLNeYZYCtSh10vRot+ObrO/ufcsAtFrVX0iy5PDli4bo
mTahAVovrtyW2P5U52hQgkJZIjbW1OkW97KSYyFRkzi3dAq8HwLLrKqXIw74BjBD
KW7U9CURCiilkWEdZcy3Lx1oMc7r3by6/iLouWsetlQ/c7W2IHgkYBe5H3dehuAu
kZItD8/NG90vF7HRnD5beXp51IM/DM/hO1CKGAlqHadZBZH4J4tgxJASSFBtduzX
WtatLJFJyACDA7PjhAwq97fZwBCEJFvTamU1TQnlcBLzMe30YYPnVviiFcJsXhnG
syWuwvVzDOhO396ZRM7Nj3bm2ZAfbGocu1hUqHcnweQONIff5ailD7d8gViJb+qy
x0BIcdcSilXxY4OZ9PV6cgjiTeI0tjLAjJgVDz02tnKwOOFe/APsg6huEP6RzHNh
RJZugr5smLPpi7fpWBQLslp7TuxUTLINZADuuT4kH05d2SmrN06v3yb3IIYfjHQD
CJhLoYBcxmsol6pBP8FaGuT94NUMG+g8PBi2w+RGnLGk57/bFryxB4wkM/FaDZx9
ghYVUt4dhxLSn25yca0G/qXkMCi4Hlv6wFXyhknX9C6ZsPeuaAFfM8p3UnzdYei1
AR4W14cZAQy58tUXS2UzV6Z7FC7K2Cxtv/OjVVq5u0xRSsBHw+4Sedtd7Z70fe82
lbV69YzhuPtv3pJEne/AORkpuOcc0zHtTXA5zNiVGUR1Np8VLUGhad2geso5iwUX
mzVjERWVRFr4gdGzhRMYzOdn0o3Q3og2hdAJCeViqk/QfbKk4+op/6QNvgEBfKd5
x5pwRrnHXpLtOfEBJDykpjwWfue2eAFGlgkPfaMZIV43Iz5fOzv2RwwmhP4wK1bu
nMJ3JhKxvruqcNkcEcKSvL+WaSHaW5UWD13DKIccVN518EjWgFVa7ae+jGx5aiG5
3Mb+tHdpeSTdiPGYMoSvi8O0JbAm2/s8TN2xE5jcxiynV6e5R+90f5oPza8/MZp+
FmMKmQ/MqmPUHy63nAy2qI9Ig7ne/Sva9zK9MxkxuPcOnjdnmzLlgvW0Lx+VWOWP
7sRKjzBGl2kAdaBOTfRlhgEuwWH/By5TgOWrFS9yAc71c4Wv6YUzHNvmqLpImSgp
mgBk43888TAiZKfMFX838PIAeTN+P4a1MBNynplCDCx1aJtGFjo1bO5itq7+y9Mg
pRCGu4i+zdWrLRRuYmgepyLfXHn5ftQXTViampqKlJ2VAWuGz1JU2l7t/9RpyK0C
IEULaB1LugimBkfljyPOp7006GMXySr9UJOaz9uRy+452X/UqEknv75uoP9as4gg
t4yT6+dgsxU99KXoYOkN41Mv4Tn/VsljlFQthTzJj2w1fDjbPqnPH2PIeTEsBHqx
6m2F6faU12Ib2JgsbMl428EPyPxti1t49EH+Q8olRuPWZk/1nrtHoIY8ub3BSeoH
JS4w8G6/hyycKetVdVVMrjE3tZ8GnscT/ySfjdV1VJVodIjx495Gg1Xx5jg6XJeG
rQ2B1z+GBp7aJ6V2I2OhAkvRAY3XXI5Ho2zGRUoqrQNVJWnJPpNV89/bUcd79zwS
V7Jv1GjJKnw6fImmUwWkgAySvIal4lSfEKM6YGvvaOOG+/UWTqq3+9XxXu0msa9W
mbNXduYR5h3Xgty4jpDWFjHX8AJc/a1xS+m8nLwPBdnLI1Gd34EKbqu78cgmPJVW
F/g+mm7Hp+x9V+WEJE2Jtx8RRNUdnVS4f7xIJfqVZ56wRX9dvq0wwzavJXPNsrC3
+ZlszDZ0gfXIeu6tuYafxGasToelt2ypz5uEpTKTviK3aEPPV+/YWg3SJ6twQxs3
4UOzDuThoADcN9YnCsb55nvHbU1Tkz5F9eJyfqzlrb3P1/TTFelnrspJo7LeTR+C
VdjCrfEHTfXc2E96WyzT6DisyemiZiSwlV+iWxtnKq1nYfehQ8pAGU5blc134u3n
SH3TBBCX8RYNrStK1F5RG0TeNLCxNV8gtbSo3IFQfJ2ytlEoYkoD5SNHZP4AN+4M
eSt8Y82GWozJ1aLfVUmnETp42McieuuuvPVRDsp3Xaks1wtgKXMsLPh4tkS+RSDt
eOvCo/mcEn4BxwF4c+vcYYBp4xy+bt6kdSVZfZLD5OQebA6PXVIq6jcfuoqgIbI7
erUeryLPKlINPkb6h+JucTRNfxR+S4dvVJ/T2oxMu1r6xkfC1IOY/lHcSnLkkxkC
0MfuMeHpUyqi28f3BPX9HLjT9wg+inuJsz5nPuB04qBIBtarEbB81zfrVzlcRt6Z
cCn3xWYnG1jmCri+XgK9EEpnyV8iRnbrvWbOx7pc6WpLAXeAG9MmIR6ZoKtcKkHm
WUC2kIaI+y66TIgx9bqWtAoNazuq5nGEPt8aMP+W8Hd5JA6WV72gcV1ISjnIpJlW
SeI1WF67nlxRaflJvYq/W9QWTaDth4Of40So3JXFvZVssCCRSlQ0RsqCI60GIxZ2
vfaDgR5RCXrVdCU2lNST9WmoTbZFNLqECw0z8QFTfsriitTKsH2MXC7XcVvysHVy
ih29fB0CBXK2xXLzhHKi9OEF/4o9/cFqFKnjpodRFn1Lkb55SpMMgnW1NypcxJiA
OKVZWIvMSZNl7AHoFqEM1c9hPzbxOzvU/FNuaqoFFKIlWhfJ6ADOrzSPQpLsEOhg
soPLwaDuaPpFmKO9pPN2x865gRV9GIk5i4XTzsT6Ye92AU4e6pbsX0ghaTniTVJf
G9U1qcqKwce2g8rGe84vkMnCeBZd9UU9cmDUwVuBvGmkZ8mCCh0zEGiI8vSClUtT
8BtSFz6Uh/YgMUsgVSlewyInsWRb7mlLeZfVL7o63NT05J06Np7gINTfCRlFtfHD
S0SQXObL6FNzNzgB7MNzL8OKG+Nz3TsqE058g7oR1IFKPM2kURJVoPTnAPifdOXD
gFTX2Vh0mP1sURAl7FQu4dlHz52n2r4rM14W4dYxay6KnAxU2a0JS7RPIOA01MPS
PRHxW6gY1ynO4m+KtWH156fn1ezxJ1t4dCvJzmuDvcJcqvtYXBUdEVnXowmLAJYL
MoCJAwoJ+j9JeLbgdAAmDaldIANM1Th2yGRs5QLnnm0GKEc3QEYUs/KZlXdq0eZr
8Q5+Z3IKo4PqCpe4hLlfQMnBEntpPK4+TRb3BD2jLqyQsy4rhpMCFpJ1wq6zy7xE
Hxlfd5J+AOkDYrd3cad0wip5MrSxuqbBMwem6ncBlNEi7wv5Cu3ZbScWpYHad1b2
VmkltNiXmZ6J4k9v51raBMJztp+dJuJQenkY979S2Ly31fEkCXwmquQdkMLX7qLf
rzOKTZ+waLeU/Weho/jgkSrGHlktXEgq+S+eiqs3pajtYr/DYRWHp+l+rRnQ5Tai
gQ+wz8cCtGYuEMIsvn6jgKQwn98zk9iixtcqMvTi7Dsg6nlNn3/wv0TM8Ych+2Bf
pdEyxxKNQx1oxHgV9tFymj2lG5AEPOVUVFwJC8NG95dk+wT+5Xizi+upCM3EZQtI
InerAmPP+5Hn/RyIAw/1exnQE+exoRqGVg5IGc1Lmb8/zjKq1z+ZGk2uDbXktTZp
DGGwvMZI1JBWjw7JWxpnbAGvyw5OfkObf2nHN9w8LEleGoSVh6EJhiQpj7p8hKWu
mGkJw+Roe9hbkwQ1hi1MejxVvWjrVRnRzXhom7CzWkSz4IUJqA074LBvN0n2dJoe
emFPT7KGXj2EXLpgKTz5OiSZ8Nu/VfcC7qgZnWFcuoL1GnjtBDVNtSv61o/NxKCU
glt6gPNtRhB+h7MCs8FycB3XuI8gEwhOm8GimPs1nEBnEpKDyy+M5lo9TQkXDU/4
1gCb0kAt68Mj171CGlwGoFZ7UZAy/gnlTWWQQG/4ET4LZ3Mpgt0bZzY2VCuOdcqy
HGIeemqCC7nVwCk9EGGOFAyr4bFW7NNRm4nIQiL0ZTNsmQKvPqoSoegd9ItfdG4U
8yx/YjX4G0a7H7UM2FMahG0fMvOm8N08F6eT4T0AYiZxOgUT8+6X1bj2Sof9/H0a
7tLCzrU1vQSULtYcC+a1N/MhQul+KmNtLN14f16YN+4H81+ShR6Argo0FeZ8RaDi
d3Ju0DHfjjlj8gHG3CSw5JSv2+OdX8FD08u0EnaMcA6+K/7ImHa4iPHqONgIlsOr
VWie8t3zHA2A5xC36WBjjxOOoH0FSaRFCKAR4rzG/m39qpB3o2vo/l9eFbma3eU1
D2pPyqeX9dW5KEyJxG9HMHl0yU2jL5JXWnoG/qQsbedVL+n9xoxkiIIJJdVD32nw
LlECalPkEt1w9Mo40DWPgkhJ5Z8Jo6ZGFzUif5bzYGBOhz8rOhenml/eCGHbgHyo
N8a5iV38RQWzarxxQecrQwqh5+S0h63I8J0NoW/sjoYesnbB6T/lX7aFzSsoEZ3j
IIZ0Ebh42aiybZsUt2/jfYxCWk5Wys/phcXpJtQJ6yENyQPqXVUD9yWzFAxv8jfF
OY2hOl4xyy4UyzJyqNIi9uSUjvhwUH85oMohly95kdqs5R4T4QzkcOytlSBundCm
UBid/y/FWH39CU7WlrbzFEfz19clw6kMtroEOZveBobfcJT1tDNtUlUBPRDUdQdr
D9GLN1R7PgwVRllwUrx8XWYt3rbwqZJLTArvZQiHZbTjBuu3+X79wktMKbqaXdaJ
4dt1o7blHjtQc5jaN2Qzf2h7akdd+lkLjc8H58HFgHmgIQPmcbXyPZdWgOImRhwX
TczWrmvKmnbINxEuMOnUjwh9DR5UU/yqper8NvVDtgd/lg+872RUr3mxlTOa/WSS
8+G1scqDWeldgYFQg2/V4O8BDzzL3xoHKahbuQP3Ttd9eHx2vlJquFTCaxGtI8ci
76qM5Z4Jo1JNnz+XVSnTBcB28LQe4iDlkzAidkf2CB0h1WKw6yG0beB7GSEt12AS
lkgwvbGvpbzihuolENwpaEFPjZ1FUV4rrl/SVn89/tCpGYU5eeIqBAqk9LGVAwKc
K12qEDzu+x5Nc4US1DdZDeZKFVONHqYX3xho71GG7nZXSNWV3cLbN60FvSXvG5UH
34I61ejXOVFejacAUjWJCSadm0emAbVhnPocZHQlhh48pROh9SHKzWg3hRUEq9RT
Mii/Tcnrg/7rt4vN6/6R5tdRaunExal+e7LIO8FFS1oJ1iF7fynM5YX3s8CU/ZgC
Pt4roYFxGiOO+lfbjPRgPrVatih+aklNNGvPvFRd3QxDbtnQwyg6QbTTR1fjX/hi
v+5AiRv90dFpuBbzARy5ekcqGG+N/YCVb+t39WRmEn+a5HxfJzgEp9h2MZPBCQeP
INjcG+cowJToJyeMmv5NWzg/513a++I061YLxvLbMF+1ifjdhxPpEKfOMuHFXhU8
uUPdJALJTvG0woZg7f32hnseaKOkX+rpKYk4zbN37YH3FLtDtmwBdCVsDSq+Viet
cBxJvYSqcOE6k6CEzM5IjEByyW6X8nJXdTbw2VsavzZHnl1hJ32pukmW3hP3Zhvs
7bRXo4+k69770kjQo/iC0Dd7nAPdyG9F+pjRkhkW5uXPldGuM9uUK/EqDTJ/ayKI
n2LXAkgv/esWnP52jkpC4D6Z7eOyFmuujM+5jVATIeSP5oY4s+0k77j6yMtPB08J
HUOxg6obgKV8e+udiZsTmjSqFcbC2RzEFnWDg3O9RkQUZ7qGA4cQUgv+tXWQ7UC7
hch+C0nuJ4m3x6JQRZICePP1nBwvy21BJYoJV6QEvCK8qIIalBipmf/btarH2aj7
yZFdL/uKMwRfqv1hPAUcuzKXEfYYUUiF9C8h8v8DEmLKp5pbmhegIj+4uGWD+1Yq
WEAefWuH/k/Twje/UmE/ebY1SnbB3AB4n/9denUnQuBCeHt3/yKECk1uy+1DoNfS
onKypmaBi0oyV6gwds7uD76P3Z+lSOikojuvKt4TEn72/Hzt60+23ABPhyC8h0ej
N46ZOXY70uPaJkMSBa6Z8fqecnbY3voylfDbmHlnQLVOnGCJhWZ0Gax1X42JjxLi
rUCQFrV6Q2eMXa/EI/ptXWcERKmwiNb7tixYjWO3hUljC1jxYmOWg1eg2tSEtVvj
yXAT1W7++IW9HoOSsNcu9guEkOihVVJghF5+N7MyQGex0XGDvnTeyprqXW5A5OAA
HjhXWZQAvIoGLHjuxzsbKosmuelpmgr7oWgaUws0QK4HGSHIKIs1DQWhhXnCxwrC
C4FHW9qN7qQtw5rgNM3tcrWwHq2kqKsYP8XggrGFwSbZi/y8DxjKjwRGaslaaXmW
2QniJ1jw7J6tQWK6RhWyZVIxA4PW2IvB6McAXdsQ6mRuoJNIhXn4smuo2MBhX/1Y
HD/ew3h3+hDW1Tzhgj5+zbhCKVPD79IrlRDwV1idZPyaooG2V0dZGWLsdHfVhjZO
PrWWyHjUsIH0SUIu3PDOS8AeF2R0cc/n6+84Gs1ojYmkXmMHl2YR4+Hl+aKN19Bu
7/uwmKYEk0773Ec3dwemZWCuJ2RKkLpVrwvR4KA/vvi9s0aqy7WBTRGQuihKlfJh
DZfuoha2u2MmMX28KEunltXxQJjNRsB9jLLI4T1WGcD69FIyIJFVsfuPOky1GmBz
vttmtnXefCBH2FsgGi2oNcEByhThmkSsCtDk0LK+/7JEHH0wnX3yfuhTDIzW/Awg
5deoy+PQMa5dv5tv+ySW0fSmGKnImhZxjVxGcz4DGBh6+6qpIKdnRfhkXlLFgrYG
8n6lviNUzRs7ql9rmDTCW2mN9vcQpn6Pqoh1ck1Tuk3na2c7tx0tXlkiMmyv2SzL
bTlpOA/3s6QjNmjGiKrsd8AuCp7EgntQp8Z1ASkY2p69uBrA3ZwdvV6PdvFQEJgk
7Uy9uoiXW3zHYtjp4WC+wKTA/f2Jd+e/0SHwZMX+jcmG2gYNxfpootp+GcqJ7Z7w
9YoALgjcmWoClu020LfXHm+AXw2X7SVY/RpfQ/05ljtF/n89ByB4eLyjF0tpveaU
EPdTkKdKWBD8RShI7h0rq7aq6txS54tOoHjpoelvSrTApX11QcehJwiyCXh8/ip0
JVc6C4N0dm26SPjXtq2gqy5J1WRQu1DxQ0lcNbe3iR5fiHSFpzFAs8tL/GINk5lC
NV3EsO6dRLs9v3L1cbkeEew032uFFtVuGWh843HqUQnVrV328a7WUFqIleyR8pGJ
Oxo4KVHzmOassFuvYzU1K2GQEoLdnzaeDJpT5xxk3YoIfwb8CAI2d2kHwZaV9/Jb
ISNI9tSEPdPph0QyAsaFVhlytzr9kYA4aClNCerlw2h782yzdNXdxRVhCiOcHdsN
YscbNAVowF8HNkXLP9odJjz0wm8VefDQ7RPJYa1UugOIal0GhcDCw/oBPkBIYTEN
3Nt//k+9zxngIVgdhs5SowoJIhbdW2Am+qSgaWytHO2HGcbx0xPVAC6NEfGqTrDE
s4HjUqfXIWaJuPtJrm13TeBkL/KgfQLkcRAQerpy7UPwVclbTOxTxFt16TKupSzu
E+q/cog+kJJZmC39Brm2H+jykvifzUUaoIhxY2Ki97cflrlsYGxEQb7w8apc3yo/
mJUz6XOM7sOXRHuA3YJCC5tWz+2Vxka+3A2zaLSyl2DjiOVQN0R+B448dkfifp+u
QmcFUYhTHfQD0Oqqho7oCVA+K9hlA62Bwf4fBEkMqv0FKPfEgpPMc4gfHUVukWZF
BekSZ++yUs2VzJmESfk9Ln9L2rK70xAJ4gH2ozma9+ues7t/yTWfiGM7G1kgGqlO
Zl+6+D3tJiLolEx88QGCONQxHhPGzcrz0FrHCD/9/rmASsMJgPVDgmsC1Fl8vZeo
pQpKI2dVq+Z+J44ZfouwLz1duNu3E3/poyg6QaVMa3cJf6wY0qnCYRBp9jscVHAG
7w9zySG97QZ4LH7/VeBssXakt95ovuJZiwIoBZOUx1Sri898KGikLHCpklirWlpy
7OYA4wfJ2PtPX7tj5A672Y552eXMkyhm5k5WwBeR0RTmZu56j/Ut2onHQmKtXxuY
vmWzqXUHFfc1g84/NjIvpGgtrd9PO2KAGEcaozh1a24ggRUYOpb6b/VVODzZrrY2
6+UZwNsXkSbJZTUSNHRSHZGiV+RohNHWARSN/SFVAchc6nZZaBzIrqLBbwpcz6vP
uuhsPP71Qn2SVgqcGtnln5PmS5mDl9VDsij/v184+5NJca2EuPBCf4URNMwXor0B
F0hjif7piIVVWhBEWFEBi10pbHPVqJuXAX5NjubgOMHCUoT5WRI4IIMYXl/ASknn
uZJS79NDbw9jxRYH/ks9/wkdgqDNTA1lon9sSFUBUp3srF66IQfhxLOvx5z79g2v
52u9hEB2dW+G9Y2g21RHYeHLMQYIBSsroH18FfiFJ3gjs7yoGmiaUQ774XkJl5eL
omFZOr7x62WsEf077XJUtndg8D2S82u0yPnZewU5+4u+bgtaUqdLUlMDYVgyLSh1
4mrHK8oeO48zUN+67vWFunZvg/jLLakce/rMZ7d5CbWjjDImFATbzEhdLMcwEj2L
z91YfG09ED9NU/mU7JzCqnM4nZwMxQL6ONMZi8L6Pj8XPVtS4O5Bhh5o9OsVgy/U
YkncGs/c8hmXYKC/enPvLx5q5Tm1qwe1pa6UPIm7/HUAxN56/CRCL0aoK+dthvyP
2w2ONKI4386m0O3I37iUciGNu5SE4c6TdAqJdhMeqaBOwn826wvHHQLWpw4ErWlW
f0LpxIbEbPI5QxoduosSvnfZGD2Z4wyhGoJoe+mNQSXyjgeyqHDDUmIUYcxgoMZL
HVxoW1b0Ls1zQgFGbABvA8SDcax30EkFJoxB8vlU8XyzqLDjhT5jzZhpTTX4h/Vu
bSWPT2PjmzwrARM+lCH0dDMAkvf8tqaytVyuRZnEJFiI/10sq9XNX5sf+LoTGFwx
UInsdwh8CjBJBNch+nXFCblV1NXtCFjnLqTZvA4BCbEbFcOiZ2V8ElxwjcaUNy8S
xFJ4w81LPoSuqx64gpO1XqCcE0FemwMx36NdEXBTKY6rJ8OyYTltSE9d7LloxaR7
gIATqPkLkWHGOTxA+GvmgJ8Q/ItIhOE4Ec4Ek1RQI6S34md4WRi9Th2poAoSS31h
BA9ddife12nEQZFu+8g94mSiBbYFjHMNlPeHwy6Et06CKz+eRVRNRDAS/NN50nza
ZHQvr5z+s27+ypFOIttyNgK0/z6meDCNg7gYdUv9KngFGpLQUcYl4Xl6ktmtJDXJ
fe6QXQTSp2X4mlyIrFczW8UOzhZLU8IRn52JZftgrhkzV8eGpS9PtEHnF8INkoIS
pNWBSu9L4RG4pPzh93iwyCUuyyYxvAlf61og/I+GImq5QsSxY8C+Y8B3MO9TK9mG
J84fKthEt2YUy5MFU1UPO/kzkFfypDllb+2UZKfDdxuhM2tlXtOi0BPiigfPBXll
gzluiOV7vRcspJVXkF2YRoyPaoaD5VKyt+hDEAqrfJz/jQ2ScO/Bb4MnySg18vgF
POYLXRbh1OOaUfXic4Ud4rDS8uGSOBDLiFydbxmtbzS9q4ne1w1v7BF7s87fHlvT
Wp9TLxKalZLUsgjdNJnZIwy59UC5TuDRRer2Z1y4xPn7mW2Wltmbiy04XUyzqAQs
0FfG6lvIz8vJPHBo0AOrcmtIQ3QtQmv3bXrEYnQTajoPhPUwcmJuQnS28K7LlYze
/KW9KXMU/rzqWwT6gI+PDGmFhXdpVPMoO4BYNF/e397baj+Yr20d1LcHSIJ7yM5Y
/8n5tpb5RVer4I45sQ/OPe4tSDhSZPJ75EJcBzlsNao6UJoNSugFr7xPD/sjZFe6
imJFpwlNlG8RB4d/nTGSXXmfBcTUZfJl8zRIZCR8REpVn8Md/VDCJbc2fOc6P5D+
fQf9H3dnWSb0O4ROUXHKcvFSAMbbApK77SLa7Nn6wm67BKXk1I383IF4EjFJWvun
ClhPjLPvxsqmZPRYLKmoc2AwYi+wZ4ubmpbsOzeRSr+j/Tt5GyoItz5pu7z9EE/p
/aT4Fq02TraalGUn6RaJuIJX5XAGLZEe5sBgIFj37sqTdoig5K44LojnvBKOQwcz
HtOJS6SBv+EMFmJRwxFNolpZgDiPWfxaKbZfLo4rM8StoZkyB0KkDgb7imLdjBRh
p7wvAj44DtAI2fNs+6K2FomUvB9HBuu6nPlJkIsgqNQbfcTPe0zN35jdhQCgS26M
UnUHpohPX5FrqKSexCj9ob0+PEx9FrtYIZhT/EbPjbHzxD5tr1JVJEg5B2yMkDNk
29M4A8r6H3HH6bcg6r/eO7JTDxKQ9JGWKQI91AbwUn3ATMQGb6qH7qOL11+VDlbT
6ChQxiIfq+S9TNigyxlWJgsFquVjafFB45V1nL51t7BDtZTmnbWlqtygiXd6RPmN
13OQfy7qMv6wx9XKjQXNYOyAnHKy8n4avYug4QnuP30NlVVX7rsArCq35pDsv1F1
Yi1tRIfJmumCWCDrDtfZTgmJAGqXoVucBMdI7CHlqs8yAODNq7LObHjtWgWtRQEJ
Aw9zC56l5L2OImvtum/VUWpsBZXlqQt5FZS5L1LEqAyOr1exoR6DRe2Ayf9PSHQK
65iEkoSy40A2c7nT+YQGH70XYFGJ1k47AvsLFzud/C2Rypkx6jxuxDn/sxyZDBuW
G1H2ioj/QySnT7oQCdPiIQ4XlwgjgRaDKcpKzFaZUd//bBFGLzP7/+oTMnQ9FMop
7mKZYs81HeiD5appMMVFczcRDwV1yywYLIWtOR/4jqORWrR1OrYUgvHzlzvV2r4a
7TyxMrUuz33qampGjGYLqTsu4BUtLZzivyaLdUDPSCfuuDQl1VvxORyv/oMBrY2D
fi9fboLlZforITiUonKxqInGWQyVJagt0FedqGu96nJC4xDqoi1qP2wMFHfhcl+q
cqIQioZHTmcktMPg5pC7gbl8+9btoHaVpiVNW1fqvuiWQIYAdhfB1O6a5TluHjSa
WdKMdN40f8VQkIwhwedPLWU4rNcy7bTEdz6g6heyCgJCqGKor6LLqijWcyE9HXIE
o2vmfOPOAgtaaycGQhmZewYd1igV5KhDy2aqsQHlrj+txJ72UIdqx9LNPv4tGIn4
hmNOBet9HblQ7lwSP1m1jcUGA94LZ5iKN1qX/fWn2a2E1qhaIkR54IBP5NhgztPN
jD6Y1vAS8YsGgYh+bUB2vWaP7YdqN4gU0q1fjH/d3qyfUDxnzhuxSLbYzLXHU5FH
NYEey0iKRpvRJZXkOuB8TOBTfuYEWYcvG7YCYSA203zB5AP1+c4c5+lm36wMiJxc
Wx6zW64pcxZmEXc4Wn+6knLmQkB3pFmElQ9n/qTz/kMsGnAnlfOyiSCictPeYZCR
nsCVX/OVoafMZ3u3cLc+Jcg3MX1s53dz5Fb4lIJt2FVQVUtkuJQGaTtM4KtftgBE
OmvTIwnx2YsvR4z35Fbe5u/VKoIn3hIefHjH7LyHvwqDvF3BL6ZJAG6n2NnUluGo
IxQhRd9bKoazHd7uabzdiRmvJ2fq+jf4d06RyY7PSiokLxDG4NDbo4zmfSxTlUcb
JljYxN3nu/+B9clyPGzA9O4WKZKn8rVHDKB9A55+s1UOavZLYzXRzGgYJ7De51hu
YY5sf5HUd3MSB3EsrrZ+FtOxB1QDfwEwudxfQZ+Eico0Z7oIqp4bwcYOdVPRSqLH
gUOtQzCLX+Zlgg1Li4wuGdIepXKY1o5oKxMCIKzOzKTJG+neifWbKGIQFl189CPC
tlrKl+7iCQbYIdcYoysQp+/YEhgRRbyCqCm59bZGoeMEcNvL58QUW6reQqKCngfy
A7QeRMrMxWMLnp0TO1o60b94+1VNG29EUenbVLL9FvZuHFWTAYfYsag0uv5951cq
Dd1SMp0t2Rh30xjahnrG7HxGPGSyQtmxryggYd6kSPYfhhjr2A7TJEIFQXNdTyBL
v9se332v21848XN/tJdKTEx3BZZnX1U9glLka/7gwA7UYoxxIoiUCEDi8ZgpSQcS
gZsDTpoYeCN+GD9wf19FKV0o9lH9YZLcuxF+2r3/dOGW/0VF8hNUsqEbE5nrZGxa
UoE+Br0Z9JiwR/gkMDstDIcJXVosPrhzxXPl0gEwBMXLW4VjA4vcNKJ2nkII/7pa
wJM1Z87RizV85swqIVEFE+VR2hkPgtVbvNwm8qEaXpKfFJ1ODKJKHIkTkl2iJ2SE
UaUxmoJFrP2d090yW+i4sBVVtuiD8Id3CErtDxa9xlM3wy4SmYyJzUf2LrK3yPvP
sDQAlIsxSWutlX3TLKY2SkO5cYCFFywIr9znF9T3a5vtQjAIc38FHpOBUuBvR8T5
5PMC3nNlsW5EI0Ob8iOL5z/eSptFIy7XfXDuyQJxndtXRxClP6DGEqtWoURAT0vf
8KPqnmMOXQsjG5frhZ81ox+ndct1NKsZ+/jv0l+R4xXFNFfTeC41VRyHXau4SjY7
BeAglBU0jQ8GcXneL6TnsnyHDNrhokZgd+qyKKObANSGfsGz+Pdy0AR228BVjFIH
4e3NwtqB6WBc/8G+uZT54KNngcMnGEfSm42RwvXSsF3ckW+hPqD6zgrXPP5/l663
0FHYSXFQDq+NQew1POGCDxJozJ2ZDNOxvSTf+1PZzCgbSnT4ZVCdrmWmAm+mVhni
aT90BhDYRGhw34rPNKPqbx3S4P2lIUMGgltV2yg6haQjqCKwWb3yY/7cXRB54e6O
LPstXcnEanoO7nnNtELxBaUZsS3iZ6IUcTeWU19Lz/XmFNBZ75J14gmsBQjTboND
EBKiCPOUj3UtJy82Ql49QU44qjuDPm8qiitztsQonAFVXnkTrtxpwZQu5nkVb1zE
mXN84qDmpc1yn9ujEU/sz+kUVVNZg2EqTZeyRqov9VvAClZO/1O41MhvnM+mD6T3
woklXcu2O8qM7dB98f0L3+HTAKrCMJ1eThycYKRSSKEgAOg959dp1k7aUD+n4agP
c1zjmxyDnBAWKag9aHtMYIm5O/KyyRO8UcEIkyowCIJ6KMh6cPu7vMRgFsvW/ntA
Xk5Hi/BDjxFgU4QTJFaH6jpOs1z3h8oInaqL7e/a8OHdlhqvtBpA2TAGzT4P3g2F
cIJs1HPvSZ4jz8j5Tvr1syiSPH0tqdFeypNqECmshZejHd0MlsQEveCP7OqVqZlQ
iEfV7IQSfut574XLwCvscD+ezqcZtSDE0DOU337OSCKBZXpf488sOIIVydNzCMQ+
a29gghThBXdIj0nvOwAdg2JhvJTxEtjkPZfNyL+8DItHG9FwOSqLUFUx63OrMdGd
1yICr7rX0pmJ5nAcNpuGqKAQze5WGD+Ii0w4FDoZIH0iD2besIDaKwoEEI3N4vPe
rBYybG3mzpm1x49SJ0E44UF51k3QCwRPxQ+HjasXPF8La5LkCCFys1JxGeeNe1Ug
J0FPvRwYPu2rbDwVZThR/bK1rz5kIUplcj+Mgb8VvFbK/vAe7J14q3fpkpOajF7O
bXck+Fjs7vWjqLOqSB34MFznmcx4Ii/Md0UxOyTr6s0nPjXgg2KLKoyBMgJGhVUi
aIf/pkrFXZQqvsCbzVNlwL41D2+5CRtaXQ656UdNaJirVrdiaqQfm5puWuAvRxg2
JVmCZuThCYI8QMaImZPXvcgQz1LAnJAxMg2cBEdeIBq0Vzdvk8TWaF+yKrPKtQB7
KP9lhNs8zTvq0iBjPXChdISCnEpK/siKMLBrtIJlZ44PX4C0xYxSw1wS8KquHJNC
kvG4VqXysD5kqPFZ8ynO1UQXqtYiMr4E69yw7JtjjXLV+KPk/nQvaMkWP+QYSA2m
qnQVRS7HCug5w872vp2RRbP08+p6tohFK3DvYhLv0rkHxEBjLgsFTyRGOsjb8d2v
VKNCYcief9Y+y31OQzqzcgJtO/BzTbtYdD9pJ/gC3K6sbQkjPkBa8XIKhJLFRnFe
S0OMUovZjPgaXY7oiWxcarjta6ZcRb64qtK2Zc29Q6imj3H/CTX4paVTkgyNctg1
tuo0GqaSR1zjM1wdkYgKxMYziynXBwZ2g6QCK0u7Tgi+Pbl7BPKFhnHedWh4lZqh
PUmC52o6Pl4hbGGU8ho5BD/YMaNiqDv00wHsPNqIlnvKkhqoVh8BdnoFgeusYHeu
SUVyvIIGgz9eLDqtOeuBFiMOyYYB4vtn//x/j+rwIrPKwa0IVHOKHPOFui0HGVoI
HYgv842EBsflRBgw90QolssOlhJ/RwfzVQ/xdsNlFHpH+9gldG81MSGw9nA5jOZl
s290k0kTGGXvxzQV9LoNSzSW01R1BMdQHBDSxnFErz9vtKTjGu+5dHWYx+8P0riG
uWX0sY+RgUZ8ed6hzYVw+2KKkjSID63j0+WDdNiUV6zf3vzXmBiUPPeWi2Xl6MX8
q6RCv4fmb75ugx3m6srbzz3qRAJLQeWJg4QtzkzB4wy8hjT2Q1Bi4DUoCxcSYRHF
ZcT36cx491H44qWVMMXwIzG014olR31+nRQWtnzVrLxjOA8IQ96fWXo5XNIM/VTG
fitXMhvgQBSYOyDI12QLu8ROp+F+fXdEJ0EFoACxOGuKDe9r2URW4X2/aIIrDPek
GPW+JYMaqmv+Z98vIzQ7fFgeaoCOqxv5qcBshFHMqDl+lb3Uton1/iqXd4OuVNzE
bLNE0z//Kj6EXUQw0lK/C4/wwSWKWt8jUo6QL33PlfgOHNQMwt6L0Y3yI/S9fEvL
pN+fnQ/EB6UprkwmKTrb+zSmo4WAw92UVrwaVBVL8COORO6cRRHC5+xq06np+u9F
8O1PmSPgdgf4BNrYzBr10UlC5dQRcX/ECg371vqfeUMqmhNhDztte9h+8/ObIrFd
km9EcN+cPF//Fixl1HboDDV2rvZO6cZsYjJzCTKKXxOqts/zwun+Z70fUtpSM06D
cL7uZYg1QRNWTLBK3BRyiKZx3lE3bYi6Ou9SppIToMHraAAUO7HHhCl8TIQM56VD
kEMz29mn9DQTAtwOx8tISC0paqyCp69qjc4tVngTa6gWQV27UhR0oxTS0PtqDKGx
v6HRPmJkaYUDlTJw7Slr/jIKiiQ6zD9IDWPlv6hn0vcNZDAjPKZx31JMBIkgg5vz
9XdFMnGVvJmtGQ1zNIU8+/IATly0m70eNvMvx2hzxnX6uCLrriNjYCcDEXJVfK2o
1fSMLnPK44QW0W2GZC5+IfTrCU9JjdF+u28vM8aYtfbiseoETfWd619K1REVknOu
/bfpxovOl/HKAjudLrkmwCL46i6Y0OBZY71wogeixP55E1BArN7AwVPek0Zs3O4C
IWKgf7VpRgoWogdFk0TP72fYgGHU7e72JLP3HIpj0y5cRA1DnGdPscYQyZjgAynb
0zoI5sGW3/zSvrYfrq3CiDI/qGB9BwqI1v6KKvpiNiT381q/zKluGrh3zPPFS9tX
h019KT2WNAm1TDXYtzZWOwYPHkyhXu+1EcYGswgzwFfjm8ellpYP0dDYeXqjQMdE
1Oe8gZjoO2sY224IkS0EWILtswwS6c3WuwXPCVGVYiXMTPyStJGGde7paEN7FYyx
mxTfkIXm7jrEWnN2go/OWfXorQO0McQx+zaBI8oolzmLUei3JWq1MruQbLwaMocE
244bnFCEXUYtrJFgLmd8FqRckdXH/hzot598922s3Hgj05OfqCF2I3xhErWjVUOs
39zJTl+rexlE5WqiWM5mkyF9OR2e/JgPAL5cDl58FHePKs4fkVZdLFmrcnV+Sgaw
ZTcQ3BBpmXEH4RJhFT5CD3bsnMv6yJO+2YqRuPePAYE7MAdjzLdDeiDEoyU/mcbk
iPnYQ6pADnaKA16zHQvWCrxsJbDCKP/jmXKyVPbWgIDWAwoKTxxJMXqUzDCMOANO
R9WFaCidKmxqYO0nkoWuGzDQvojnDZR7KordEeUa9pFwWKfYEryewqVR6r/3Z92G
WoDn6RFPGs3pc0OtzwoS0oLK0uMwXotFY4CDcugbbw3tFNyksiN/bX5flkLdZJIu
J4UmF3ns/guwf7hxWM2wFQnQWlC+oRNyWeGJaq825afoqAHruDXQY8Ny0EKTa36D
aMr7ZUh5GEF9jibiUgKrd7Pt58swy1RJMmmy90ZRufhoXR9uvbucqDfeNhGbwR8z
FQdcHGVvXXhO1rXBIYxqrPWQAkX6ZGXXT1F8Wq+E+T1H9D8c9Pv8bM7XB+sxtofr
sY+AQESlEohmNqa5VJDLxTGm73q9VSZFl30V7okPr822Y/sTAnbkXVwb9ZHkmxtJ
Bs8o9mTbZlhlBkuGIB6Qe6aICfr3NpX+E29EpryabTGCivzQKeUSoW54roE1efDZ
T14tXret77fBaisRBwmVLKxYUwL13SA8zCnq4jOgLC/1CR9YXizziH8xydYeoZE6
dpMnjG3xC/BSPf+LuYFj45rqATs/kd3BxAQ7vJ90D47yqoeJa10l2ft1Ifi8roP0
e8bD7y4Oh9+XxxTFPbUvzRaHFiv69/HB3OXGCIH3X384hbNpSetzSe3svLVfKL06
2X6mb3i2V+MCYjpgfz3dqIMl4VQ/0UHm99u9tPfWwzZgcKpTuuu0/063HRWD5QIv
5Ihf2bZ03Fgh46LB2tVAXz7zS8PigaOEFe9ZllKKS8k4zg+w02dy6fF3qVyj7pQ9
I7Cz7wt4SeUMhRybjhMA+N3o4DpnAabzrTKDZ6CwHZDqnhadv2hljqM2W3AIbc7X
XNGJL3xsg2Ha6oxCp2tdimcIcFkJ5hqJokTbUmqZb2Vbf7JMwTYpceMqwI3I0qp8
Jj2tgQTczYXyC0lmH0H9Z7M6kg7OJ9YLgngn3Czt7u42ots81He4qCu+QMx68iZJ
coBFg7ZFkyHzO8l82BQhIrEQHjOVBqq0mZjZEQZ3tXaa/r5LLd90KLdvWtKJ9705
ZX7YgCzy90DjF2iy3iL/hgYc52XoPIG3sZWVwnJGUZ8BNwVJjbGphs5GhNisit/7
LeZbO/0QzPe+K9McBgl7AZCr6evTrsFNzeaowgU3qeEN8dBRFBPV7g23cgcix0Ud
Cfjje/MCn0NCpgWcHRk3aFO2j/GSB5LTYxRQrgvjgKCFgcAEZsZntu5z/DsYCnTP
Dh9TE3JNQFyI/ICb8qmq4uSzS8Lz+OXvi4tteAqmCPXVJtio0IA+vKTY8igVkTZ7
VFcF42452FvWt9dpDj8OACvP9ujOooNtuLjDd6Wq7cjhJCMuAfzvGybo1W1nolCk
My5XvCEsfroaMs9v9U44UVWEk3I2M05LGieCM/TukSUwGUb7j9ggmQxBFDBG8fN8
0i1BEWbNZJWfqGI3BOT7VXhGM/G6MUG1BU2WPioq2Aj2Jn4q1o46B/WH2R2gZMKD
8Y9V5Bq4Xx9AFwva99hDWchjIsOCvtDg/IGY6pQR8bTx29Q1cI4tuNMhKb/jNd4k
eW5grCEvyMHRvm7XzDSLJeEG792J7obLyr3heHUbN/Yq1n6TeDYbKUPY7LGgkiaq
wtmOsLdjhCk/tb32Zn2AG7QG0V2Hk2EfJcyP/3DCSGBdnCICe2i0ZVopBbwNaeN5
y0sCWC9VkAos+1yTU6b+I24hmSwrJpqwk3unr2tZhSMUoiVakUVKnhhIVxyr9iqi
GuFUxeGZ1n8Q/84q8EwBou4bRFdP4F6D+FA3dvHzqd+seKI1uchJfGUZzR+LpnJk
xBEFrB+B0cNGykMUDDPQfvHgkWB/pwtX1wHewIxC8G2yXSqxiVNF3Bj9EIhltJJc
C4x6k1zueAdUoXPchQjOoLMaOIIqg/j8GRJbOVSDHTuARJ19/2hv/dweG/m2e8Hy
c6Oy4K7fVa3cb6KPIQhrM+Doe04xQUw6HhX22gPybT2yEkYP6ido/Dsde23XVQ2P
voEy9uSu4uoS7H72DtfBPGrkI846dMtZAp2p5gRSv7K1+mhVSAJXDoH0+dU4HW0Z
Ue4ZAH+pUNKp5QcY0rmHOOBBUcjXrk7rHe6W4nWNeYKM6IYgsuhvJscr0/3MgCYI
Dem0yVb59At3j+N5zL0lUEUkZGffaVoMsMsPP36juHrIWEcKwehQSzWSef9H/QP5
tM98D5UYRMIL7Ex8qQskLG9g5S/Lue/FNyZNZoD6FDeKiWhoEC1moRPbvBLaBaPA
VqIh/2PNMD+9f6CPjKAGzelzP0jjBP5o3mUJ/0trqRYWk0TXnCiRwUFm5BLI9QZQ
9F6PauulL2wCJpjYgOmW7hsqURKziwmbSFm9ESmtPpooSwpSjLRZEB1Cqde+OWRa
fvP72cRvDO3f9+e9RM7LKsgMEbD/HzOpBTN5DqpH7OaNieh6RJATSB1GD2DI0aYL
YmAGT7lzzCvgwIqoXW4t92+Gwo5vuY9Bhc5bCrqm0AALKfWKjq5wP30Om44Y0RKJ
4VJY5+NxOdQ68rugtVYeV9DWJiHIl4SvXBouG2J9CdBdGy1b5IyFiGR4fXJrDm3d
Jif6hQHgcQl0mUwpvx8z8grg1HmuvJTpM+HaCaia/oIqkqbSMHe93SakFy5PZ2oc
2e/yWwL+pMz4N/2dIMAiqkkIMCYLeh0wXMO8YXsS1694GlhFUFoCd2IdgKIKu5T6
5miig8uARnHu2ePorYBjKUas0WZeZdVoafFCxe2A6Buf6c5omnp0k6cvmZ/7Wwjg
O9ij654kS4pUhq0Ni68Af6rhSC/5DzlgJleamxXnzpk9eT7gqsJHJ9hSQhzohRu0
SaJJtqMAupjVE+4H/aQlork+fI3RVmewkifbJQFigLh1DUt46IRnwIuNpemWNz8s
F98gb3V/DvDZYCkl7unjMjLW98lfq7+1GEws3mgNx3tIqxF8LSn7K8D54IFQ1jiF
HSF8uv8fsblaM6TCXQ9uC/GCuJBfHzZSurmORBrP2VIG8JbjEAaBiY/D62lsa10n
djMQGSdWxyJS5A80bWf1WCtj6GPKhotMS8i8hvk/Z637LJd/xqkQ1EQF6kowu0Hy
XeJ/6h3hXdeVwpO4BHyNhuLM676sutfPglOtXvelwcQ3LKvY/2UzmkWXnjQ+1Yxy
OGgIabnsESr6uYjjkw27Giy1bYaS/6m0KuXcovpQIdVDCUc2kTySglVdqYB0lCIL
h00P4jjiPWhakOWwAgZ6c0RZ3JcKoHK+c/8hEbKo75TMuRm8sz/ApjVDPUNj9rAY
ncR1OQz1sxBQWMlh2KnswwrEi58cSiXqGYIh1TnDCvOcSmSBolwy4VfD6X8Z+5cM
NbszsnGKg/KVGWD0Wl/9Msjtdr6K2lt15bB6ZPS60HSEkGlJ3gcVKAYdmKoFFnGg
C8io/ZDCXz10TrTjJKuBFyGE+TNbb4eilg93nDiX0s6aTB1rVT9Xpr8p0C4McgKE
p+qQv0KqyecyfioRfXG2qbVA4KwQGh97Pp9CoERRYXsPMQgBF6aVe/LQEotKoew+
kItw9Bm5nvfPLFANxHv/D2wghVaoioStA5cCoXoqu7y3eATdez3ZTL2y/0uM1GCe
PUsLTBEUqT6EkNCmTrzpXWmm1Gg3pgp2vvitQTc6eHT5xrs5TrnyAlrv+yWWgVXR
jwu1dWS8gdmuvNRoGEm+mb1OyFy4XzTyOOEPuiCunsIOzSPr1noieMM0Ao14uVc5
ALhRySog1eLzbMZf3xbL+Hwyg1ZpPwdWfqtN5m5Dej2BOHid81ERlW93u7XOVQop
vIC6kuLEL2P4HVEMZA36Kl60lWdKYSjjkTU6pJyr57Wcdii2fYS7nvyDZHljtxdG
Oxa22wcBTdUxJLKVXvQDMu1pq2En4Q0uRgPwPpGgYLdqQc80iqMETQ08LRXbF7Yw
MD9V4OQAHr/lGn3muluoP+DvRSY3AWJ+K8yZT/sbASA56HPUR5++x3sxxNhLhQ1W
7qMg3Uz8rnQ/sWluTe3YgFlql5fMU4Dp9ab5VO6kuL7Bs8WeTSgksCa++AoIR/Zp
OZs/6qBybeFz9FMPht5fElUuctzMa44fPRx8fPlyTruQdGIaGtXi+Qg+brYEh0qo
yZd2iDf0hhJ/s5/pHneiMHKjjGvFG2wkfbv+aw96IrBlfZuzUIClMeu2uFzEuwAd
GlsNrtD6oeO5Dlb4uDvhYdrhK+AGO9MU3daXBfRihRV8he4BtnoQcB2u8AVyn/x/
RC60m1944ilBLgZdGbMW2Pn5mpZ8BU9e+mk1Hs1zkhKe94T34sk0o+9SMWChQryE
Dp20TrKIwErBMe9g2xXTMHx08cVaODYdG0+8rEFVJlV3Y3Kguo46jy3rkFwGCWWr
3caujjL1MKVbHyTA8YfbSphyWDuN+YnHoNzjD8PMCYxtLVreM8yC3R4beieZOi/p
WbzfqDuWhbG0DJAG3z+aOHKjorqwN97RWlvk+TTr66QDRW52nC9ejqh6kHo8OnlZ
Afwo8WO/dHZDQ3RifMphrg5ARBEKaVzkcVbgqLFEtZ6wvBR5YxZZdAsPn0Mq1IMr
PbB1yw6t4bHHxMCbnPQHHXY1o4mRjd21GiCO3lmXy+gl04aVLQPwbIHz+wNZnpO6
6l++qLMQr4GjKOTf6aYl/ZWI/Gg8FMKRtkKoo7kx9EmEPyIAuMFLV8l0lfHHFqek
PAoN3+RmPErVokgGekBKOCITV3ka1Vaa7Z7cZ0t8jdMDsb/KMWMXkv7FxSYwVva3
x642SFk1UAeNVuUwxiTFeFRrL3GHDq1HZRsUAOfvMR/EBPlBt0+Sa8ZKBG+3zahF
Og9FJv7m+0r9Odx0L+3NFVDlDyjfHgDm9T1kM+5+ccrkU7c20j/p2Q150onm9skv
SrOhz7UvuCTyyQyomhxPBxYHye8zcFoMIU9ByjnUS9pCUf0DJSfUMYLyE4Qszknw
xxILvzvt7IEL6qxECcLYTUzuzMqaTp/vU8+4eWGvUrzjWh6mFXXcurZosq3G2nKB
wjjwbdW8gQzLgabDbHtbpODzgQiz9TX9gn/VX+zOzvb+6TwVTv+asIfU4Jc9tGGa
djNd7aaKljrhQyvkmmftzGTEvK16CymRd+9Ly2y/kVp5v9+kgC41rDu7VeTo9zTK
FrV+HA+S2/ViXUe/mzQ7qAkVvz8NAGbXPonZGVWFJThF/zQ6DJJsnkf6+eSP700M
jIB3JDBD99QrYiks83H1BC6Si7tq4yPDfAPboknoRx2qPWxq9onjemgQyZypM+Ez
ASO/ZBRKBoIJQCao9ZLAvPI5waVA9QIGsGn/qTN1aJIeZg/rNW795bjXRr3aCDu0
nMlqhsiTaASkgiqQuGhbPCf/p8qXCXPXliihSZSeT69jRDibxjdtuy/AARxZ12Kd
qhS5E7gI7iujPJw/aCvY14gdNhDjyE9B/qhPG4Db7IRn0JNkxCa1tlqdiZUnck+y
O6SvVEtWOPVKIRqhY/0HZnZEMf9yX7JJxmEkAgx/+603T2tGHVq5NR+uIOxdf1vG
YRjzMZLesIOV/zsf9w1gHmHLY/5GUOqwcfPKpQ1q+XvL67sM0nKMDLHSlusP7M0M
pYddwhd7VCzdBj5EaotkV3RtpGcAy+3XUbYIja/GW+EFxfMtTW/AlkXk0lKjpHM9
9TsDAoOvnM4G1PWrSSUAKC3JtxF54X8VpnnFgJyckiH1523UgiygTpRyxR+q0Ygl
9gXt6QnQVgaRleFq6oKc1sbdx+dT1gokjLs9cFp+RDsp8BlwuF+kJZlsGeZNr+nP
yexpvXS5AAPJTkfk5Q2iROsGJKQqja/KJZNZSFPbS2zX6Y7oJKbz1B3OWId92EZM
zD5c2pKcS5v+fUULv/YH7a071EQpUMPqa723qLqbvVjZqMrTHz/LDcWFoV5sqK4j
2ioRNf6qKWgqQ3WfOhbmo69ln+Bl27+PpY05vubahxAyxuRNVN7vla4XSnbvpQSB
wu70SkcE+aDHpelb9sRCyV8Fcm6Mx/cotnTj/Jq5m1jWCG8Al3zGn4uFY00gXyiz
c1W78Rnd/oRM/lbkAfDGRssxUI2BQYOBQ4adZNQ/1Dawog/rFJVfteBeZP9XGLi1
W9DMqeHwYC6nk8N8t7SaxnKhJH5/ySPe4tYZewr61UJs5S4kYzjQBogy1jX2u7Fg
YBiE5rY1rtbZ3O1a4Kv2d7FlMZ2ITVnWcGOJakTrZGMv0V9eEJGvUXsjBID1qtEa
Rnap3MGirJlB1gZJiEM1gqmNhvb959V7k4+3KXE97lmQpi3LKBxi/DlmxSUGudL1
YSx2vYlD9hb3T2BXsXDwSbJt96eGtlredqQDLaBunKsBK3TgRcF276SGg/UEMA2i
x1PMM88nAVmsJH/Zkl34EltjBvf+G7zA5Vx5fULmq28ULI6JW5BE9xnL4/9yISGa
BmQKAwX6LHIy0iemMUh83GRM6nV3n/Aw3FzxijmFLCzkTGXQwL1VFc8NSZNZaADg
4g3WkdZGHrMLVZ6YfL9qfi6YMKqy9xazVyIRwwKeEiAnyxi1pumCoVpOgAcswbCU
s5onwFKkPPdGk279RoOkHFD3Bq85k7wvvqhX5vPgpI4BcYRTHYylguV8Ldm0z4yP
NFX3oY51liz+pMppNd8yhmlel2E6YovcQK9I2ot1U6eIsuxQWfbniJfZ6vIcj6bF
Fu9JyDig4iaaVPyKfr+3uMZ9NjgGy4abmZv234X/EaTClvgTCKiXAMH5stppb3HM
Wj9TsnuRuQbV1fLnvVmMtctzYl2PVCmq9D6+SiYFAHo5PEcUffz0+zhT3lUDriid
aE5532t3tO8PBu6oQy7BfhQzE2uLC+Hdef84TTQHYbUs4tOiDZWg4Ak+x/kT5sGI
RupdzrJ4M1YZdOMV8pH0l/TfEy8hwdxFmS1dah8ISRDXhcJhHpherjDSfdPA+qkY
YG+06VL2pQeA6HwZyAr+dze0GvS1YfM7pcZgfTFUn6BbATdQQ2sEXG5oYcmx/+eO
R+JHimejJV5j2v7vAtUUo+E7aViup1tL5EryD4w0hDeIrKDOJQ0a/zxR115FQATr
GQIsEFgHpsbl771CmuIU8clxlTmezMj7FLPcY8jQhzTfzXe7AC912/Qa62fPFDK6
S5Rlz5DfPjfq/2mHVPOGCAbb/YfirmhYRWaQ9BcyiWutVivHe8E2IjN12x6xmeT/
L3oS3fWy/N7qnpDs3thiMgPMmVKRCvgOQ8TfRLHbYvKxY5gQ4iWkCpaAxqT8DUy4
57UEoZcPCZS3TmxymYS3buG834mYj0JIvyf+ehDlaPQkf9Y3BkHXSt8SwwgB2kMJ
J9RmQTxMDCsQCssFa07GhcFE03k6WNjYYYOQ7AhR9mgeIgjxbZTPxR4AUaFw6w4U
wF1ipMqKnWeMK1Cy0iPHywJatVzV18OkZENOqRXmwoyh0HHOGecUgEI5c/6neaKa
fkVzZzx7jkGg/6onaZvVkEktFKfBzugoZtKDHi+P6XiCA2e0TBrFu83ONFTePj8j
qFNDSJSMgEqRQQY5Yt1fQEIZGMZQsI/88LC+RAkvrFi0Pv2dbG3N3zUETox/dFHU
en/nhS6+fAG2CEVpvmBPYW2QlmnD6VxUXsiZMiLUqzJRaxvXv81J9weus5MVYsWj
cv3Np76iQ/ybnEe4TuhxGxajA32vojZc91m+Wey5iN8YUO8rgQDrCau7WxOufzLR
lH3lSgK8UTrJMyKsakMJYQB+X7uz7HcddtU8GB4ZiyHer3diM1Ag1gkbFZGWjc0R
EQEFO3xoPPpumknXDE9WKmYsI02EGcJJ9DE2s0bD9jJy5Ej9x1A4vtEg4s2juP14
hHYkAZTuIV96NNOhYTOIBbVHrY6QUAvUgv7324dLhUR602Bkxe7PwGa4rlg5Q/Ay
4BNOUisfhiSpbhcb2RwMiT+6Z+NHqheAVA2Lz3hB+6VgJ3NFIVRQY1cH37EitrR0
QgNtMHZyuo4fBo1c/SeSL3Z4zZQvzJsGoYJaikbPTE83iEA2U67RE7RPH//DoKgF
55lz2UoEG3zQXtYbODGJq5H/Ti1Cw+6/9ZiAdGyRMFV0tYdEBB234E/1LqZxhfqt
e8HlcOpw4ztvX8f2xheetlHLaJqp3aX8FregqdOmE7N52G5KJIIAF2pEddWoW1ho
ZyUhTWGXIsA+T2zwv6UegZUJwy37a/1hDZF2vtmwdS3C1Hpqm1R3HuhPAeo83wiz
e//4hWiz9SDUcAgoUrfHMrfjAgYM1SKDdnZEG3y1MagxCZdecwCayv+VC7WCnrtR
j5uYi5ym1YkWrv+ICY3t48DIivNsHFTDdGpq19XYgn5iLvKLf7SS/pCJ5oC9AOa3
/rlwfDXAtWD7NUAUorHo5YOhpqvhTz/OewJaFBg1S47F0a/jiLCBtcas8OxGcAGq
IQW7DbvBXxsNEW04gc81G0rx+HALH7NiX5EKlY2kvxbETc3ugUNMO0dbEvQB8Y2X
2me/sRVb15y2XTiD/FsZGb/kjvJpBLPjjbtb7g1BP6a8hashcT/90reXM97u36Gn
nGHTSHDXzEnnVXjMmTHET+s5lr5LbPppNVF3gxIG1XKBN+mQ1ygM66rY904mDHqb
Ac/SaDfrtJ+dFvkqoRytDJctxjTNk8GSVOPWpaHJJD7rLWi7Z/dOJ0YGzbm8txBN
OvIySQMXT9s1/oDlWZqhRfATTiSnEb3DXJz5IMfxfm7xXszVD62mkXjdT5k62QH1
FSJkkrIwEAhF00leEQCu3APNhSe5Eyt2mRoR2cqGo2tlEK0QoQdaxTGrVuqp9R8A
B17v0AiTsyojifD2krI0HD1MwjGHnX426MAwDxAZheWjA282NmbsIjuwAotMPjOU
kYlEc7SUAkvY8oktjr4FGrbGZN7MDUtDzaqTT6ZVWbaebEBiENdyAjA05DhCXF3/
CGuPJQl1WIQZAUQslo3mZtFJ9wmIry5zaCYimoiUOhpr/DBABI7zVxM9aaNuGZY7
iczJfQ0KsuApcriravenfQwmJKojqJUCs2S+w3r/jom5xkPSlCuWMdMmeB4YJdNu
Ze8zNnTidabUZgyIfmcvyoYptsw4NoBsHklP27RurEV79suI+a0u3QVnXSGO+DMo
/jcDhbzCOfHF/GMFXJWNoxbhYD24dZovM8nGpw2W/me/sxadr55rQlLPINBr845U
zYxNXSfxQy4KuDelDyUhlYmwYXXhiHfwDRwvIboRSTk49BWk7rPCPoeCBVZLunBb
CUBtaEBAXa/GRthDaM9vP0KjQztzPfuMjB/X76FD2UZdmu8+XBxMLtCcIwuSdVFv
DsfPpDR6Og6srEIgh3FRZX6ZIfayywv1UdjiBukOna196Xl5UqpoyZ+5oiBfyeTv
Pqw2YBUZTQ7+Q5DVXgRDNEQ98UhnrBapNu5o4X9ITF/NeIMzZM+XxJDOmrKYczXg
LmMx/EjVxy6K2GYDs16rNfs5MsrWgl+DNXwMYi9Zxc8NKIPLkqQHw6uCMBh7jkAC
0dJF/2/lHex+nQpBjxkLhftz0nHtZ/QkBmm8W76/WeVVmzvwK6IjRbIp9Ub+efw2
YGihpMA4xmX9Rk/gp0BFVoGa9SPWt7Q8r4HihmDES2NiWyeXUKWnfeXJe4Ok1asV
3qUZvyeZkmtLS9SwfYhVDtNVLs6aQQbBm/DzVlmwlV8wl4bsF4DyWcTn1C+1Xl1U
VokGaY8Ohn2ATYlTZMSi89yEyvJ8SfkXM1YK0RtP+XJhuPJ5kTUMm3AEemGfkaL4
Gm3mTAmwjv/iT0iIIRUCM1jRz1ONsMx7PnGDyPW8YnviSOZ5IJUtSk5UjugwiKsw
GHuUbKKKgVocDtrjIyn8WlM0CC4OtorQvrk36x5VsiOA6mHVzrYZuCeHPe+Xhpqi
odz1MJSB00NoyF9f7YtyXqLsWQndp0Cg7A3xHzx+2//EXeVy6sJqMStDOyuuDrgP
l2Kep1iBHGK4iApD8TCcdaFH7P3muqrtquqSrQU4ZY8cBJelyzRLq1Np23ZvN65v
Eyo23i2hnG4QTzsG77YktwpR0wItijvEgTzRpdbsXLSaRTn09zxkzgYxW3X/v5QV
Z+Vt20xfP9NLC19185aiWJiQsxNpCGHfAZQuMLnKoXiCEUbL9DgkG+NpypdQNTFs
EwMSU9Y3cozFLuQ1HZHG5v216VKpRH3JyeooFDH3qABy95RNJobWUkD7+YaNCdK8
MUMY7CDR4BsU4dmxBZQHC0/KT+tELQF76rVYvjBfUkLlSnhKwXOHd9wCIqJuwOl5
VzEmvBcGLFHGSMdn4SUl9sP4s5RCRgpqUHonjW9ODkNTdBFD3+xcIrDx/Btivec0
NQHaufBisaumv4+w8zFGx9pbFqYMI3R2fyvZEsMPDiXsDusuvpQ8YH2WSphiGP4N
GDdKPjXDTI8ZvVeZOSpMcMxdgMbeVkPAGmyf9xLfc04F6dQWF+WCJVeRRcqUbVYf
368pe85P9gLc300YLVFrBdmdTXFFil+o+itn2SDMqCPBJIWuasn9YhDEg1DOrgOC
Dq4Xih+RjLBwlv28mM8w6RYEIwbrV8+Lt/Fz1inao3AiHGThn8UTun3gDbdEKDbL
G1VuXIlhwekO9meBH5wIcijF8AKWSxu9gX/JFBh63q8AQ/oKobFHb704skfyPkW7
O4bHFk5wf60TPMCQTfPVN6BOUbKbbQKvY1p0IdPnlr0dLAG5p7oeNqSn4QZlgucO
CH4SxLNeVFJ0DAmbo2mnwpRXxW7QgRsbc9BCnwQ/HTKlOamcs5/unbFr6Xuh5Wpn
80PfOsn0+ptdfp6N8RvsiUjtwhc5BjZpWTpqid+IAOMnGE5yCK5AtOT9bDffMqko
xbmjUqt5dRjjMJf25ECZIEbFB4gBODNXGKmdoOHrJX75clagTFrwk9JD8EHhaGC9
JHK5Q5ETTOfI4PbRkX5LcNIuwWhAWibd14TAkKgCdUcb4MpZCNkOrI0gDO2UcM0+
BU5yKS7yuRVhLPkkPnzC5yrRuUETib1AVMi8yBqDYMejP1pt/SPRd8/mtJNuC31F
h5+xGciMUeAjFGFaVKjCctBXYcPVzCK8qLAyOiNVhXaZUdnVMcZ4Yu2h0PUuplva
eX+r51McCZ6Reyl3qNAto7OoJXwhw14BzttxQWUA4A1mQPr1MKNt1HUw6YZJclAd
9B/jPD0CU7NhR7d0fKpT3sk6IIdFdzbVlRavigULXwkEV3YhEmxhdL+gzvzs7q9Q
N4v1lQMrlEdcCqS43IaZUUR11Qs3ML2l39k8+GZmTTpJPc2KVC3lB9JrmjoVs28i
W8xfNeiKsa1s6SV3xvfMZz55dOwZKLVPLLlo3TFSgtPcN5I2/Cb13vGxtYcA+KEG
So4iXZv/EADPWgHtTDgZt6bHKExGN1J7FCkCumVtkxU88kuUYTPYxYLa3c4IlpIh
Y0+2wj2vY2q0RrF0MGxEcR+awDx4/5IDMpr4DaJGMdsqlQ0HCVoxm7CDdBq9tkzi
LYn7+aalZE3aCcQVkQyBlHgz5H08ZaM4/zwNSErqBZkeMG+LtuHTkhbm5ylICWiG
KSO2v9meQ5/hrDaOqRN7bsPJ/Hcomp0JTp2slSAWaon7SMmiZ/2azCwNk6t7pk+1
KH97PdM5WfYhbUhld5W2rrrimtnVNCcFo2ZgXkxfZb7srIQAhoiZTmgmwez2hy99
vJKoAOZ/b5EYtoM/KBjD2ygGRd5d8AtwIXTfzu1kYc/cGKWa+J2T2q9gteh+npbj
eVkZTX+O/vUqHArI+tgMSCzLFpDL0s1TDlbXHXIrnQGG0vkJhGXkSailNDziyce6
frt7zEH/cd6YvzckL1TL6R9evaX6O4Eh372cr/gIgoQ98U8VL24TaL/MbBwZNYXw
xi4pBiD0x8Fl82Y+BECuXVmDQhIJ4YFGPYMDXlptg9AwyxuW0iIsXpWv95fBf2gX
/OHGxtPq0GWGpBMvp6vPrOz8VH9rd8Wr6ZI+CgqOxxTWhZAORai+bEgZ1j9f477J
IhYcKiSqs/QgGtxJtITjGXgZHN0qJmsDodXnZTUfd155GgfZifMGQ8XLtujHpTkm
mIYRsFx58d4olZHfARxlv5cBseBcFIl5dG6ha2dIky9HbWAfmc7Nl+p7IKl/9hxN
tqhVYN53Bh+WI1xexNfxkSj36UGEQLzVAa2a13QtERThBojDdYaT0goG727mCv6b
gpy2Eo7Muyc7YQmGc6t7ojt0UXwuatVHTUOQJmEZbUnUa18bUcW7B3YFyywU8Mag
EP3iqSY2/C6zIggCd2a2hGOJHFxIjXtRY0AwuW1X+cOCjwu282C6Wmzt79b+yS9k
//cGq5YtxD1LZf3yi72TEmnw74mIr+LiSYAylBNJRJh/RkjhPB6y5gKUlUCYZMjc
K/J7PDG2QPpggSbew18tfJ5PT0HXXEpeCsd5HVTitItHwIFcoiOwe8ZP2YZrzgk3
MVEvOc7X4vi1Yac7dqBLG96HdZBOyqTM1gSHaB0NyK0HV3/QU1wx3beyqDAgIpBV
JdZWWU2dDKMkNwSoySll//ZnT2AclaQH/5kMENVOEeLuC1mJZIO2ASCBKoJOCwfx
eDAp8k5YR+D4C0uJ5A5z8E6I8MErjHTnN6mKITSymF8advqsAUtFJ2BATNezIAaX
0HAVLAnOZLG1K64QDhqFpTMvRaY0VdvECdbUubqPd86MgOecgEZjEJyIY9h9TXCe
NAb2wO/q74XGyIaHy4Ba39nHw6u72r+N1UFr7Z0MLvztllq8FLzbXO8bvq15daab
0FF+RqJlnvHM3Xqy2BRkcUN1RS2HG2zXGOAnes8LzAWicnieya12GqZeo6GXQh7W
1yweAb+6oyBT+fuR1COg5oavrHS0iGtILL2zvHFAXJimULuz7AG9/4MRuYfzydat
jus1YL7VBU09tQ9YeXZXgpWJsv3oE+7EbOAiipSi8jGAynGlLQ8zL4ln78UPRuCI
xUaiZGTywdxUjrrGYQfmsK+mlyDQn4h1z3+gAcCtjXAZFloUWFwdrS1v0d9zXR6n
S2yU/nNOMRk0i8VbGrbVyyGhCQczo27zIoyspb+x8xeylP9Wn19vdooABgYUIa47
557OcK2gpcHOdVg7vRUSlsk6VaQi5Cf3edbvFQ80LtMvtEjXr+yVjwOXxu6JzzD8
XmlpDNjv8mocsJWtO37wFY90jiGB4rm2GdcoAEhN5iFlVQ8eOnDi6bs8dB4djj3t
rTwRuUOm0t853mfdbQFbUuJAnNYaM3UCevzQCKbX/rsBDZkrzzhdlWER3eSR8UIN
dcLnPgKL3fXtV5o7cipGru969eCXzenR6wvhpN9OsMDfpiJrtC1TuUjp1GrEHEOA
Y4wAiuIcrLSsB5w7mjC8yhaCNQrynmKtoeC1l5BzdCThnGfmOvC2SHpzQi/BgEwi
rpKQtTMX7JArO7gnvIBrPkoPazOJV+I7eEgpCLPhGadwthBbkex0uoEkDl9aOo5U
5tmGsM/60wKGkL6qZeOsuMMb/fe7s9/DG2V5iGhqPjYxLi2pWwrBlUqE78aGB9g0
OK08HSZTam63jU3jbR4cMpmKcfPhw4re0BJUvyVFDZhdKCAPGQtXrjWzC3NiL4mf
NSbD76yRMIhWiVkUbMQmdJWyHseMqiu/KRhqeORIFHcJnUI7k6SdrbqiG5YbdtTR
tOvmV8EeRx7I2dmKSAXSmNub9DV2qaXyhs5awy+19LRbMEpG0W4QjemyJi7mmUSC
LbHCuAhzoU6786419L/xaXSBFkXyl0X4FvaViflZNOpE4MiWfW0wtRurbFp4VXv6
au0gkPs1a9ZeqYyl864KHty732x1Mdgtg7y8kaGJI7t8Iolip4WLAjh4LqUn3L+Q
Rqx4qBC5PGvdAfY3TrD0467CzT3f0+EDRoRkXYgq+5ghH3htgxw6aATW3EtXeBI3
Ej3QUASStn5STbJ1ajDRiJEf4eL6QTsuPfFU0AAjxuk6Q6XrM9u1pvgbSoramVVG
ofYMqH5lsZTS5ZCg5a3uJjAduJaAt23AVnjEClgoyEhyo9R+tKiWE8d9FYkIniSi
IbcS03jFT6VzFInCttxX+FX6Pa5+LZkA5z4kqaz5PxG3OGaDNSMo/ZLOdyts7U5I
/1kigIW6eINxMZWBPZGNS54rY0AW57+6guHaGtKUoX3CzkebR6GLW4/KOPyB4+aa
2MAgbdW4fFTsRhcXNPIuIhUhgQ8cWSy3ICdV7C4PmTrLkqQUUC9OKwlHn3mZ2BdF
OPpUMen9ZG5sKUSKoDMeY2ZvNDZavALOyT9DIixqQsTGDekWMvOd/jNPFVJNbX5l
XTqUEruGCsQyVjOnnjfQkLIdXLzfSH4B89MOKfSMeRzSWZJn+k5cGSe53YVRiwqB
SmcZDVGKAoDoo0ti1z/tJQG3QynE4a0lHJ9n4ys0EVobMCWjA5zj0Jd3K2+MVBTB
k9pEyNULWnReNzSQOh5Obes/aqZ9BuI7WrVEybYKld5ubBNC+aKJOna7SSMYAtHF
eJI4O5mU+mZZfuXgxGmUAwX+W3C66VY8PcqQq/093jf1NtqnFcPLqfHMxsXP2s8I
OTqaJPLSGsq3WdZ8DK8SpZxKshmiqU/V0wqkGRQbqDfVgGbgkpjsA6iOFVu6tYFJ
SX5YNTr6UqyIDLnjI9n1RJPUSdIaAtHaJsL5APJu+tkTJqxjiUDqKoyLzzbCi2kg
XWxGkg77ymBtspywzDetgxyH/y+thmEzE3805hEDR4FxWIfViLbVO3lzFOMsLwWU
gXKAnAkJ5cdVVYpdTBZnMevqggN27HcurA7KI5PbFYNZc3g3Ao80JygCYPuSk5cF
u0puudHghYOMKM7sGQJD1s7mZ75uBLDDj+0m4C4o5Ee7yZapZL9eFPblLyzswy+H
kALqcXKoAqd253uXKfbHUr5KmBt4/P6x5Sz7s7mdtKTH0en6cX6VuL7FkNCQxxT7
Qgu/lu5fb0fw3+XwOXyEiax6Lho6jTEONL8vqB5AFlm3T4iylK5Cdka8IGjpiz4X
uW9y/0s2yd5PsMwmuU7O4K+x4Ff7krq7VmRu4H9sv2uI5bqFIftBmefoRFCmNjo1
kSPH+Vc5BvfPtuFxfhHe10C4/ElnN22n4Lc9WLrT/H8ihNUuc2X5Anb/e4mwshfo
NouHsqeNWuD6SwW9qql6RODV32VGrWE/U3BBDd5kfyDgXKTfMhrxWvkUgrGaKvZ6
tXHqwXDg5MuC7XfZ3A3tsfNZQfUjwPMPVl5s9cekjpMrnrxOkPWsX2V/GlwwZcES
xqZFApS/MxYlg3F8axMSb39A1XkspoCIkiTFhfFfC98061lZ5A+IEAoYXlSHqNk2
RIj9vM9hpP5WY6+297Ovr0W7IIpTjWZalT+oAJs+lUTtHSTz61Ey/vybaU0hnrTT
JQQnTybn+TcwRIwqdHaYfuWMbQB4B+7xv7hEgihB7fGPXJSZV58lXehaK8sbklE6
bij8pA+ArKLh+N3F48Hw7CtQmmVO3n22g1XVaE4Wrnp59QTVyOJaSohIbETHtVBS
baUAK5qHOemunrVigwwccYiHTLxIL+/LAzD6OyP9pnYUj4Pg+axls0zy7v08Xy0o
kWoQosFZnpv0MEj3h1tg9924wjwXZ4WVryZAlHn2nNxRZOSqWhj/dJCQBiza6pOZ
TOuqeYLzbQk69WkMfJAAYDydo/OVHNsOi8/e86gGusVqoySgnvLBd1LU6Wr8RqjJ
mrB7UkWiXwloXhdxBxF9H4mWKKV54zqfVn2ZbOZD7lBA8QuMlhWRzWbFzBlCwPPS
8TrUZWQomXXFNYsZ+t+Iy1pvSw11BaPp5wy/c9EFHvtJi6+YvZnY8TzCQwXhNNYk
0kKBGb8M4y12JSak8PNJd6qRS2yMCpS0jsindtgE310ORyjXF4Fmk6bFdv1o5wJv
9mma8e0LWTkODOtqpMBoVlzeyI27jU/0CUKSgTvGAoVRNYWyKDxtei/Sinagwsoc
8rkf/mDk1QT7b0EyyAhjtjhhaE8kOcQb/UmhdIFtfMcNvHu3rPkEosSOBZ0z/FY9
E0C8l1KB81zMRsWRMz5+JHbXs/va56Fg/HbRdm9pFMW3bzlwZjFUUr3479LrKFRN
MULfNJOcxaio2igJc9XA4VA2l5bMQU6dwESF7NPrhqfx9J1eohoFaoc2hUKI/lOr
n5IFfL04rVpQGfa5oUguy6BPYqvx6TSwYSp7pXjvsQ5OpZPEj6jBsF75LliHftxM
6Fp9y8g3TV5QbuP/EZcFjljWFarn0SisuUhdOHCh3Bq/zFpg8HCMB4FlmPiJWZt+
cLtkto2o2UuzjPaSU0iQUiYeT7PtMWYnaEqYiVFebEnfE61S4XeHDOTjf0ps5lMl
+DwsK3IIfCyJKhMouEQrMbKZETLsSOVl0cdhZlEZ7HEf5C56oHsZRMoiTzo8Olpq
R+8GyIraEcziVTMRvwxnwttUm7r+6XpUrQ65wdi7uy3ueGAvTnhdQ8euZgvlFPLP
aeYnTPgOG+gQx4iRvVK3tOVKpwLatF68qUApPiUsjKUyxlwECTBp+CClpJM/5V9J
9caA8ZxzXcnvXFNW9GXk1xunoFoWezWV+/q0rCtp2LCdOx2+ogrO3D2SoHOlQw3r
Kh4u4dlGqDxR6PwD4BedzpC2mjHN4QKQFORYmOQW0D/CZPtyDwdNS+I5Z4+g+b9N
mX+zO38k15JqMDeVc7x1W6647S2dfmB+KEOtffamfxBuo6GGR344CJ9eMxBYMari
uvLQcq8PGkl68ko8zIoAmiDEGaJxERsnVg1oBWY38b0JrQysbySikR+YONk6l3fD
QU0gO5H0WK/YogKT2IKBtz2DUi25YATyySooY3x4ahkJg+9Y3bg+mdlQacf7t9XJ
KnXI+Hxrxb4wFFLHtJV0rW42n2zoNH3n6REhPKjRZIcA8cQKhC91FzkDjfk8Tkg8
UT/fvwQNtgi6MKUZCo9A7X5eL2RTFS0i33zxMdgxNPOMN9d5lB1W+GGzE//MRZSI
YSsQHrVAVbHhE7lxphNcvk4sjRVcmRScvaMgFtmkywwZwDFmh2J349N+6uAVWNwC
XIsUEJrj6ZmBSUz/qT9P1dgg3hWmrdfsdhQLvTAZsJkB5/34UU6gIEjCRA1W+XET
Z6d6nURSR7amH2rDlhcpAokrliPLMRxLAcA0Kr4Ji1Bw1NYSICqNsbDKTbW43eYQ
A2d/mIOoJs9R79CVZAIBluRJvclKNzodAftBkSYaKnhly4UAV5pspNFlvHi09z6d
`protect END_PROTECTED
