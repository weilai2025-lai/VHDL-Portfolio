`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xB/SluWtKKs0aYIFxq7l+mU+hLga4cWfOe7gAEIEWdS8QgmHLTojP2at7pXjEX69
oIcDg104mdt7Ww/v69ejcPzyvCRq5l1P62GGgVaFx10MsFNvJx+eGjWxeRRPPPvC
EIY63UKY62SMNwTjly0lLotjnwf9+C4hE8HzAZk0BH8eNao+p9fo6dlkr68ge/TX
72ug9cS465nNf1EHx7CXWK64lQPFp3JQ2nhSl1iADBblRny+D3kOQqcokFpvvIBN
8YhMbgSlzHju4cWdAlL0EE2oKkHzJHdfqUx7uDn59rL7n7cpDmA6cBcjNgNP73p5
im4Sw71mOsQ1JWGn9IYrGzn3+QhwyxBsWBLq2qeZHeOa6GpgPO8rDUitsMdZwwNY
8Odmph12oYAM22bqM8Skk3iLmcqWxe+nlgBv27kB8qlw3RXhVlyOZ8K+Fqjtv3zY
TSg87URLOMBA7oeZIRL9WczE6kslRdQBSxj8IR2VGyqLSXvZ+LXGTEgaTVH9oyTY
ikV/xPaXawuQVLPr1BoXqZ2/pD1f2MzY4+t/IvN9HuxhrqkcgBb4W7mhmUimgSMZ
wXYSLeBVM56RiGnD88DKSKEUJjsiJMYiRUdakytW6KZ9piwq959LkOKT1YsqqFKR
6Ezk0sBDzrB+8WouZpNI2gDprI4noC34LyBQpVrE03jLf5gQKNBZTrxBzfUYssfi
Er/3482qJIw5JcSm4Ma68+/60PxGfPyiIrD0covtiRWgv/ffcU3YSr55Ngn0ssHC
fx2bl+xN0UUHUTGcO+nJn2Vxqls473Ck+j1XIG4e5FQqOM5xwFIty/BjkcUI7PPT
`protect END_PROTECTED
