`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8VtuxzuogIRYZfhzI5AfN8ykW3qamhNU1tqAyJdIqzXhQmhiQ8c8exPP2vYH3Tz
OAD7wmwDKYZOdSquelI6AVbEelhgTZq+XxymVXT1aefwzXBXl4RdIeNOkUnc3w5g
CUx52u4ECOMGyAgMBar0ka+G7Yc5YScAvUIq88cHonsbcPRf1FYMfHd990ZC6kpb
bo4NXW9vdZepBCrxobT7GvuPRy7OWExJF5QcmVwnvpgihIonAXAGlkWFk5YCyRK1
8goUnPWEgCVTlp3XMPPa828em+0l63W6RkU517Fwuj22FmRtgkKQ7Z4tf64XscW4
vfGiBCxWayCtAqNiF+ZsjFe+qCAcEqCsSGDdrOc2w04=
`protect END_PROTECTED
