`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7u3Fa5UR76DPso7iv7aEp4F1AfoZ0BSYcJZONit4ovqiU8MGB/JRgnt7MvWINOny
IpWsHOAg1eDq4d7WgPaDThkoxuQpLlNeHWgKtBC1HEv+V/Qt/rs65MgbfZaK4gGY
PA+damV4y7GfTV0zYfUP/qZ1Nm0ojosAtEilqObRJoo/ju6wBlmMFiIh+dt9zr0o
PHV3yzOeJ5jGZnA+o0gb9qvwZX1UIVW0DGUgy4UyRHXOFAlH9ut6iwJ9QpTQm7yP
LQscOmAAN96dRtlrw6nlq3xxIqH4N/HTHxucIrDG8sXw/YFeDItgqXwJHvou5KEP
8MjSGzSTx04DD7zYu6qkt3a4R4wDGV4yAPBv84hLYqSUk1eoHNpimeQ53O8SsrIK
m4yvpNkBI3lyb1vhqe6wLHfy63rXysfPrVxZ+juLX/0EOI0LD2cAA9mZWWwpWj1q
4fcHY8MXH3L6Hqdi5ItPs6F1IWBiV/ejURl99vSI3fyZAt2Zjct9WWj5LvyfTFRS
CLsBDncNZ4vpq/UGY133IQHwyHSIMOxozNoizKrX2rvlUPKI2jlUhcUmRTJOj35X
1iRdRPEiRUBoo8M2rZFg3YGGxVFKOcWGxA+CdLKNskdQKu3NSt9Dpr54L+8GWy5g
D1sv602WWX2aK/Or0cRYJZUSXTa7YXds67DM53CW/OxZ/uKvFvSCHbShusyAUXH4
IAu5lu8cLidKMvKlLOGUrlEtY3nmq1HW2y9asFkaIvW7YUl8CndmWrPjmHnpT6Bz
qVjZLCZLFNuZW7LikpNQ5KGxvDkz+gTRnsGTSkMMa9MrMFOsC/bh2FH/NMjBLulT
SSYcI38LUkUGy1IR25jDB8K8lm0W7GyxpB/J7we1/MzMwJ9zfdsV/fyOT+Fntho6
n/AJVMo4hVto9x+SUHbBU3JcZ1vUf3xkx4pIVR0R9tLBSx0gMDjDjbAVx5GZ5G2V
z5my6B8zGJ8bGHWXvWy/QSkRPmWzUMyGgfuf+g8RQ+kFbDENlU/w/Fy+G11IQtsD
AqpO/yOVdM1x4x7dGezgaAHYcd68vsm7ygp1cUmnkZopgjCcmpuGhJxvIboxuC/d
vfSWlVoA42oGYqUHGBivpjmE9Iixt5xU7gdVjBqF+8nDKWekfTof90XhRdl+rVy9
RYaNnfce7RCj73Fe63/VpGla0sF4GquK5/fVjJdKdrMCuqWVXrZdPHbABMJxxGri
j+iu7UBSJAtJeL/V3wtR+lZrYOU/+ny+No0fyQUAOxiYTKslPVHDqsMVAbw7pKX1
JDi+PBd4Nar2CPiKN4/XFRiRC0URsxZQH4idaSo8rveKt01qqVrK+xKWx78snYud
C+25Psq1WteRTpaqg3O6hfjMwmJ/kqdvouBbFCX57tak3RI585i6WYB51QC4IQsR
+VEORGw23Utc4V+9g1RYRHyfwJifLGVTT8a32T3isQZvAEWxPLxCt05aZvamqLgk
YiteTD9cAemOSMAH1jMQ9QuyrMoPW3mT0vfjt1xh2mYOWHXcvEshkOKjhul0oQZT
uxVe6cvep5eLAOFmIFDL0yquJ382mZS1UWGBBST2TbbFY0TyhKPOaw+COa6Wk3Ml
Xvl6nWbYfKeyTXJufF1fOdl6x3RGTClEx0jYRr7FE9JJBhJzsW+wCeB0IcQC1LD3
plmklp21+GqmgjYz5YKqeGN9O0VVIHQOWSmOkkFb1LQGhsL1Sxsne4eYQaCmc3AU
0cPatueXAAYXEbXGVLRcxwpPVLglacd/4zTpj9171NGk5q5q1Qw9umJ+j1J8nytm
awGGOahlH/cgYprMysXNnEuCbUvNeOA7+fALP9tnKgVhXl86X9i09WerVMxJvlcr
UDNPhAqhNX5YIAMDQcBCjxqoDQf8AWH0Gq4ydODJMoIspxJ+tWylkU5QxaPxQVvW
mjgJz3oenj4h11iVs4vxPmDmALN5XqKyGVIyXqSFYjobrxaWlilIlu6TAWSnLLp8
I3vYVOA0frf9K2QkMkEFeyaG9BHGDMk4+YL9eLhIaR+z00La3a0hW/2LjXsEPIBJ
/NbritjpjjqQfQ72w51Kq4O9JFdXCdV1CCSY2qW4JN+clXILcgRKJvgMfdr5Gp+x
cWgAa93biP6Rbxfr91INVKIlUDOz1wNEUHM1yjwIH8fiPXBuYUL34PcZhVTT086g
/d6HMgRELA4+r+RyBksNJSXbSwv1GD0RhMD4B4GAgkCjFuEI7Epz+fApnzQde4WG
uNkKQSgZrMzqQQyWrZ/Cu4GClEcXGWODEOsiTvccoHNE+fB8WHM120uYyDxyb0OC
I9OnH5i6nqxLRFJ9whjqs2DJ7WXBikzDQhfbOr1If+w7d5nEbvD90qpUP5MR9cSK
FOFCPWImnnm80wXwhAE73tQXKAg3wYTdKMJkY3zqKDxOxnEArBTY/u15BZ7IqnnY
GiXrGI7up/H0XRc95IQimm/cactLNc0Lc/nVc6bRicygZmGTEVuYgzRxba32rMvW
TwAnVvxkkd+8hkJYLgOCDxdgFUUJLopPZfQlYlproGBJLwrPxmq/XJ8hDw9oR5Z6
lCPMpzBPeWi3h20NRW7brY9ARyES/iPZn4fJAYRwXxhG9194Hv98O3JVuWrH2Sp3
IVdIxaG0ro2O0xfiw6ZO+g90zCi3xjCjYRwcUIxNh/LzIEHm6Fo6sSRZneTHWEvV
z04kIDuIxkAIKm6r3jzPdHLEsFX/TtFvVi+QPBM9Tm0q1FIictGw8XCf3kyAIG6D
57YXZl1YZu97BMV+ja09/Dq/nHcm2khdBHQIjGharkcnHosoS0IYLwwUt3du/kCy
WGgrlOWCGs9dFuxmzcnFmhgqgJo22Zg4NReFM1oyblE9JWOeNuvVusuKGO9GPwnw
Q4UyxAibGy+sR8zk+G3/2qdU/qhsa+Xxu0uFbIJgfXXU1Z+S1Ua54ZW+nu5KD3LD
wWo8bgV3LmFn57eMnK+cQE9d1HQnejSQsYweQydaNXS+7H1z1gI6nGSD4D+h+eTd
seDFUZ4O52JiESEBpBId5u5Uklwce53r9n7IIheehN92kfthBeMTTmZnY0xZtTp+
0AtjDii/J3bBx/nvANlQ4j80rV9/1gTpQa84tsy3yBpXQRPU6yn+rwUANZzvcPi/
yyqAh6ViMjWyS81o8YjJfmjDOKE7gay0HL/pvhAWYXKHuEEn6dtuAxJhEzKBAeJp
x8E5BehQI7syLZDe+aDr0d4kqXSY3OCr0gdQSBvt1i82leuw87xpXZnC1Pqbv/3V
oZWHB2OzqYSTOia8o1j7zhgYkR29PNTPD01Q5gtO1L1T2xjf5gweP+DNiUe5NanL
Jkg5NzyVsCAWHroJ3Tt1B+4F5PrGjj162wcjMu2aU25zDKVcVv6v3RCDowUgX1Md
OATJgsXqXzNsh/y20bSlDmvlwe20gKAWkYye083FnFap8gVJhrSZMb0ejGACakiV
+Sx42ey4NOkPyqR9RANheMItBNSkfniiE1i8djVVkcRIzZZ4Gtg55YvfpQgy26bL
d2rzN4T+pgOExA3cDnECL6/1jHZCwhYye5FWtSkjtyGptcFQGNSyF5lnY7AP+jsK
/jOV7xQvKGlFnc9ZcvUeb+ZmTGTC2ZuYctnXFIyzfuugUbfor693Z0XCqUzRk3/k
LUjEsjWm/dEdP3m05arfedChQ88IiqxmWLwTnJYTxYk=
`protect END_PROTECTED
