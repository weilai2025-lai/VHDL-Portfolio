`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I3Ro32zA3ont6R8oI7QPsYuzCyxpSqGnDGouF5qy6EaF4jM9HYkCZ1y+LUuwx8Ch
zgG59AKgO8Okq8dff4Hk6gAPrVRhuOEVPZwJuf9kZvovVq1h3gx6kLhuLn8XunX4
n/JQmKjljimepOElzmjt9owgaWa0C4KXMSvt0HLf6zmS9UlHZLOUTVv2Rxo+EhiQ
Zfuhi/3rx0AkpaH8RS1vvLtdoUOKdJiMyDdaLTBd427ybtxZuKJhuvnibHhKqtUv
58OaWi/Hp7Otle2lEO/tf6NHalKUuaYxwfcr14n3WfQYb15jrj3s1XTY6RTPqLLw
RVQkJeYasD6fpTzgEyWRS95eZVuz8OXhOfe2QDlxNsSj4FCPwBrApDD5ZdeK9SAL
91hE8DLErpKlS3zWFM3GmW6lj8ALdtfeEyC9v2dfqjZ01xaVrDCKsW1bxNq3KrhO
RmTOvxNGbSD6LeGiDdf0g/UqYk0C9K5loWFxhMzLE450zsWlYmf/4Tem0Xxz2mwr
QBKJRYx5GiFS3qWeHset3xOOLLIPomIpp4z8CFYrzgyqyV81Gaq8I+4GWPYacQUl
uGGNNT+hhZF6LOAw0LUqu+0RsCVhwxgXtT/K+7Y9HbFQFT2YNxVEdmrkR+AtUZai
sU2OrkPADl2/0TGc+TEPoNj1X/w5gCKqghGecF/wviSyBUFXhsCyxKm1130fBFrt
DHS9OcxDlmiZ8TFepy8EX0Qm7M7BS8vAOIcFtEYUvw0rNCwJFLINs+mM+/EYhNMV
RsNvnr2NUYG+Qq5oduTncyIK8Wu0OSTY6mzmStwAnvtZsVX7YFv3B1V2BjvvViL+
`protect END_PROTECTED
