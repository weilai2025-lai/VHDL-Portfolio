`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SoQae3j5QIQCc78ezk7GPDtn5qKNOJDkJx8xd+9Y9ddaURZo3wpRqjP+eSa33PAA
84SfentwEL/mBXdNDSzYjLLVbajWowOL/maXUTzYwMmR5FCsIcMqMOHAaSxKdF/8
wTcWLkORvHI3IIKWkF98sHfelG7MAclF0ct1+13IL29C7uVztzYh0Dzv815ttrVo
/bbQBFY8h0aPSHFT547drwE6s58OpDmT+4EeOZ6qXpuRJtLKRKBYd6nGdNcbHJwj
IMXRhj+G15oAjGoi8LjKAR94frHzyzmC/USj5IV7VnUP8W8jJLaQOHWreIQSE5Uh
CaDDsbrFwxWDqUUi2AvyBCVA28++47acZd6HWj0V9ysZSYIGjCk/lSNo/YwHaN+f
f8hIWzUymrBNSoxq4rqAhQ==
`protect END_PROTECTED
