`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nIPrIiHfUytHbBh4LjTiPmTanKTZ+J1Vc77QK96OAepnzRZGOCFdGrcJxmP5gTLv
2afmaZDzxgwvsjuDqFY5vMlTINGpU9Gw9i5MPSHWHSKO+rzPiEMejoajwVTq4DzB
9zHSFZQkyofJyQNc7oyEL9WvHV3hTMozt9XDMvZN84jyMJxc+hKvC72IgROA44vp
AfwSRaK0quF/Kz9k90h0UJmSofig6Qg4agOIlVnriO+g9G9Kj+lxuAl++XbLDxiR
vmz4+cRUlqw283fbxllNxwchNZNDPfWuOSV8G9gQABYnAivvPEMbAB8NyBrg7/Qy
QehKSm5M2X9OYuljSAIsc/4gfHyrNkVvgSRv+09L5wKOiSfJmPbBwNFwqyq7xpyH
SlGi4GE5A1olHrxaPVNy6H0tfGpMMPSx3pSdtNJyubp5YJQ8SY8r3C2OcJtJmySy
JZSRWQ6EbBL4fDCyy/l7pU9JmirimQ+VmEuuYkWxgVMIYz15KO7EX0ER2T/VAiG7
D07Otlw/l6tuJLnaQETI6birYNTonJiYpjsgauUXMQWxET8MJ5SxlZHKB6dW9+Fk
MY+g+Q/XltA52v33Ycv4kFEacW0EnjlQMBBloaqROBM0HIj2WYUQ5IpaWLzXbnVg
ca6oGeg5cY5aP5mR+UnLbjAt5/PRS+Ln9l3yE/5L2zoA35XW8HnU+gKmzZIxro0e
JHjnNNdN9OiRJuH48iLhhePexlNiXHkLTYsP+vCcyVAto4YUSSiVW5C8O0Ebp8dh
isr0bxm7irMJJJuqlry+2JrLHoJk882Ue/EtaHt//JMTwT0tKeo/fWDq2ZYluJrx
H51eFgcohWMNqMz3iZvFzX+PvuAhia6mXYTAmwVYrvYuQivxp8p3joS/X9GbSNqp
uhrRIEUvC4MrHrSVE/2+F4yDVOEDIdnHC/AOr6fVxwNqy/Q0U35gUfChkxqjEoj6
5VDCU8aoyxg2gtSnO6fNCq6JQiM6Ja58CPQ+AT0N0PzfnA/IKbYLbzAm95+TamJo
OiuI7v5UXD+jaFUW6pwVHf/gzqmGC7b0Qcd39FZ6qd4ROGG9+21iPspHsgjZV64i
zyCPgsPJJUS8/n7KKx/XnaCvLDkZPGL6IAs4fZCgTggtjcTQI9G9e5eRpAQ6TOP7
U3lMmuDRkSEsMWCEYwnY1RJbChS3sMHNYDM5VIrpjUzXrA1+5LgpleZbv3cv7WUy
VJjrOsaG/xdHdy3pGMrJmwaUERLbV9Utylxo8EeAr5KGJb1dii95bwzafZP0+lwe
n6wPNFqcDalAI6J23lEFB3Mf8AG0xUcXoMJflsXtT/La8E9DLV4Fr9wkTOA5GJj/
4GAJiq9GzV17p90UcHaIxsBObkmPFnKjQwjSWx6HDEk1S73+dbDWsuA5baVMmjlr
U5S5GPkimO7A70O8fGJCF18dJMqfzfRG/l1898po9m3gNm8SNQokGC2rWRGH1sbT
yRwcwgbMwg9jhnVkfBrnte4CRE1PBqQRpLpcKru+lRUfM7hOysKWIc9TsCeo651H
R2SdP1q2BkRvAdet8N0AFkLdGit36KvZUitj2pgiL+KhWbLfKAAtBT8xIpSyqzpF
DAGjKyD9lDf5T1EiBFI5SvtRxk6oEX6NGhIBw+pNL701scxzE6uNLtC+NADy8XcM
18WWGhdCnJrqBKP8Hyq3QeGBAke5cD9kt65V//0NXIAbRtrYrRfHQlL+bhM3hXQo
7osxA8VP0hfppexhfU6gc93Cbg78TKXbBYdfKFWPwSA/U6R0ZAwX8eAsfCKVVoVU
q+LBVglCfFoCpJCEfjO5Bbx+Tx4MBn+XcuBBBKpm7TJA2UR3U6fhAdvuI1GPCGmx
Z1FeiXA4c3AqcEDtYokEuY7R8erlPyDSMu5r5wXfZWzZkEGqS+5gn2oU7NxIJWZS
U4kCSswwmdtsOxelJGQEQ3PZveWoXfeGttXKE4g7nUvf+7LkhPWU/VpvMnii0bwZ
h0PVtAfVWybT7U0MvlLUXFhLrG6SceHNRCkLxNXB3nWzOL4Vjl03ckNLwj7pnOsu
Ik+LttEkQG2U4Vwpa1OBG05S6tKAHdRHbETwEK7h3K/qOBIQM/S8WNW/xV6WNpLH
lcTGNuOqshLFcvlvmr302XrXHh2CRYLWtq6atC2zj8OmqxQDEx4XwxnmTngd+5jS
6uzJp5kdQ4oBuTY4mds5Fdr+WOip/nD5GK61w3EwftbGsXjJh6sKfSSno+SfG6b8
S1KjtrCpNHN0nFHS3HPEn4Uyt97HXx8PXZ8Cf9n68dCZ69jpe4EkARpAHFd1xhKx
gQLVlaKszOIUT85HaqBXpur9JrEMyzDB7qQhlPCt+LD0/oPywm3q0lTwdboMnHPM
8XEZSjOGN4LkK/0DpN0AlhmwL7LWtFH4LN2EBDSi61G3qsSASLxtSVti2af7lmxK
TDEuxD1ypnRi/HNGSEWZvtYYhEgpFFceM09NQ7VT/PW6Azq8aTIE6PjVZY+uTfn7
qumbDuQrZDrEOSKvooP2djjRPMvO+sNtE3/DwhWaJHU=
`protect END_PROTECTED
