`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FLzP8dmnbN709jQuVDVMYkPFAQfXRcoWfY5cW6j3Ik2GdhqNdwRacz3MjVUNYdJq
XwQLUHB4afgX8HMFDXfmx000ErdvUdSJzpEMtCtycBj9plkS7vg067h3p6FZ7uXf
E07hEk4T4IcH8YDbEa+s9UzdaIYCQ2kFSNdk+9oHptpTy2Y1qkBXBSYX80+eMNFa
iQG0fQyD83NLpIp7SKpJJqAPa9IEONpoqs9ZClLpfZZUHGil0NQe7ZcNMkJvtYGw
syfg8amYHvdgcWiTqEM3NqpWXuK6ce8aCr4Xu28k3vUYM+mqYAl7V8AmTj6aKZWa
26njbiB8ForRcDtMNUn0cwypw3O3ZV3P3x44C7QEsEW+G8b/1+ws2FJ0D7nvc0YH
GGa+QVyeD7f9jT8497wGmEvRZJvH+wPgD/CWqkToMoPpc8u61bCvW4X+Gnvm2JNv
3fUig1XalJB6U8m1CYS1111r0EbftTKV0fEV3NGdikf6nHOVSlg7C3YLz8BUopm9
PiH3RAmE/RBhOB8woOu7KXC/Uyljy1C5I1XbWpmR8s2rfHc7Znb7HxNx8mq0mfpp
RzXxlARDuu7hlElN/3lZg0V3SeGoYcd5HvEIoqZpLNjVJRS+C4BxNHZcD/SQKy18
IcJLqmXQKM8rC5ChsYLXKGw/UyAA/k4v4uDEYou8WJCMIGIUdSZf50cjlx94z86C
UnNhplfvzUr9zL/hlMC+tM8SOY8656XCTDuhxsFW/8RT6lpOch2nftKbQOOfSLMG
aLV243Fn+lxSwDzIUkHddEqSeXbUUM6bLSSOcQW+CXBV/b1c/M2/jX68uzKt3Lra
BCK8Et3kSeGIayj3qsFRFCFy6kkv+V8qZYgPTrWmkbGnpuvb2SOs3Wg8i0YslWy+
SG0zOL3Rs9VR826htffwxUX+415gYL//KB8h0OR2H/CY3XV41mq/DM9eAQ0gyZTz
`protect END_PROTECTED
