`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLhiQa7F9tyO9VT1NY8btJJOsp14RuDdzMbO283ZZRKaw6zt2sgPo/QftjOoGJuF
R8+bNaBTH9p2kY5/c22To7xsqTQU/Ai4xOioqKzi13JK/URicdVj1aCaDJ/wgjmS
ml4+RQ4jaqf1cYlhd7o/fYYjaDTzpPlvvtxfEnHRb8inDHdyIQ5l2Grx2eVah5rF
GIIlwxaaLfmjDWUgn+Yl1hef+NAM6Mb3eExrF65L0BhqNsTcmiwA3yczmdcScgrS
Wpr9fSiW2dFzzVkIOnEC/PRwyjiy+uFBtKIMczsHpCSfinKvZA2DSAHJZnZky7Hx
hOaCxqf0PnSLvkq9OvamHvQs9+7aC/tqyK9ygkj4NjyDQLdEeEXwIjFoGRB7uM4i
UmatVgKIsooo7u/GqDdCINbf/VAwFS/pEDD4K+NXB//FGVARFC4CtodSJ4A/Zuha
t1iMEgFrpgNLGK98wOM25jOJ0Y6Je11HLvPnfIe0RXy+T5Vc9QgF6IRHD0liLbtp
pDIs7M9hXSJkvNwf0KhagfD0YwyNSanc99XsPlxBeA3qD+MDKqPRyr4mV6Z5FOZr
KHJTZ21zw+9EmJ5uJceFEZcYXRIKNP0onxFyhXBt3a7dXkYtJLAxusP8RVVz6Duk
dRjB92EsY44bGmbo7n8pT/GSI1xv+AhLTWZoIDT9bRiaDbs+6b8vLYo98ck6lVTY
AtYnC0PysNBz1ORzn85/PNXbPQ/gKt09PJ+sX/LtTWe/0+67vyGNnU0ooh2I6SnL
yz4RIIHJAPtpBFPkxUihSGwlvixjgXb6WfeMCIwjsTTJDOdGsnjQJJoPX+WQAAjM
dH4MEYTJymxYSFPUb98ZHFMQlVCbVqcPft8Q0yfsUbJWv8gP6Di1cORJtX/eSueX
kR+cCjdgUMPGJLnwPd2DXRMB2FvwynGX9WzJUSvA7mHzbkdGkufGID5+Nwvt5KRd
PxNso9VN9UCKTfoB+1QdtapmaqkgLEtkzwISKfxKsDUimuXvLjjRKpt7QvE27Z/t
`protect END_PROTECTED
