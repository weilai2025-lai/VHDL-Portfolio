`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AhjF8G1cJUt3eLxby8djBigip1Dw14gCgvyZFYrGfhefHS6WjUicHMG6KhhEvt6D
pGYLI+L58uENaxRx/cbGePeUy3PLzIMsJ0CQ4Irgtu/RqkfJc/vrTbrvWSYkJEly
A52PGDFCA8YzN7Ff9ffbNxH5Y2piv/qwzS4G3TAn7DzccytgIepSMyJSaYjbCXda
49VkUcxl/SEoMhvM2+R/mEZHV9J8Z52x4jDuMsH25/PbnikZN7Vf+rMGdBlLf+oB
5JwPrggcTEdQKW7ZiuPaM8Pu2e3rd/6bdCEDilC6qkYtD+bZF4nV+Dku/q7cSTWH
vEH3wnCqZdOTfREw3VeSoocrUJVq+r7iN+hRb79hM1LbJuAm/WGYYKGKchMTB/Py
dVOhunm8T+AB7FWzOC6GFdVcNHyqEM7zIuM76D3rxhMQ+Lo9KQpnqAAK9ic1oOBR
HulWpUeao4FK7ekjyT5JhA==
`protect END_PROTECTED
