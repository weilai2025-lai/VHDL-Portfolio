`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4tukXQt8Msc5voJyd+I7SJe3kJi1Zf/G41RhGBZG98/IXKidQ0k7aM4xN9LMSIM
bCgtcUNDF0ZDdfdgUi0Pc2qIcMb6TZdrehQkpEHqv7FygnCLt+Oxcj43qidrdUp6
UD7bybXi2dqk9cPhCjCULMXwQUUu6vk1j1YE+/SG9gU5gLC/yEYKtxqhetjM7EvF
J+ZGfzwGqond65ZLKk6MmIh42q0rEXf3K4OTYKgbISJ7yhLskYMnKU8TBg+CwKtY
vfQOi4rXAIsLsV7Nf+/J5THceEmp2epcinlp2yjitYJvYpCGZ07fD7zzhGt0DtTU
0P7NvXOIHutOtgKe9sWgVrIPWfRwNoPkFf7Enc7Ao3h8Vfrfx2ZGNbrnv74bmZzs
Qwnp8b4rRhtZ7seC8Eg1UQORh+cIx3WqgK3rF5pk2FIubh52tz0wHujyHjhFQkqO
CnYMSsdxqI13FVzMzurevKE10AMahdkkUOUbjjJV8XrZPoUS8AFXq0edt8UbBJnb
IMlv2n7EGnJLDtumBRMH8Hljkt7pkZLB7fGTRiV/+nuSuBhWjc9Rpvz054cYTcdz
5qaH8wFdLy4EN+F3cm+9MAnJWemLOPyt54DiwGfwl52MbA2XyFusXOcE+V+Y5TD8
wsM5rpR8pYpfhbPEFLQRUZTsCL/0yYkp+N7O2sDu4Kp1nvl/sTZM4HcvBMV74/iB
diDhLwcq8t9WrHanKKy9cNQiSliydjNQU+hUCHDRqU8Oi90LG2bbDRmo2BZSBULD
OlSXvjs3H+HX2IF+YEssuLMtufpIzjf9HlF437VcmTU9hgbTsR5G2ydPR1qiowBJ
/fIwjRPArTcFPbWdkPWHwg==
`protect END_PROTECTED
