`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzzLyao1tiZ/Z75vvqICRpuOmJXMMWnY5SeCpjbg5cUdCHG2d7UVifVohuqKacHf
mG6DDAqZDkX9lMseYG4xN6VJQAT8D4/pxu98+/gsor0+meige9MKlx7GMT1vqNEl
fkgleHt2AUZ3KMyDyzxE/n92wa5iYoB2jV8ipJMQ0tpleHadIXvZC3QBq8MLexsg
sigVi5orKuZ/zbl48hv14KqEgCDL7lpOVL29J618OFlba9wP8q+VECG1lMrr2Mlw
4HDAJahJeF9NL71s6dp5n/xKnTLH7r4acRreI+V3/JGdDC2bNH+XTM8HzRtigSW1
snGh/nioeZCDBCJgIm5py6NpAH98lq6guYiXe/9iTA31Iyc5B9byjuPYLNFAUTLx
NlJZ8kwJYhDQfGZW7zdrA6qXbOOKH3dk9kqExCz6rq1OSLm5i7SSVpZh4usnAzhC
VALyoxmNrU9QxKrRWfn1lXIF9yaHbFsamInBjPqz/na6zimucpiZsapq+76ZeLmQ
eiOEBOrv1dvaX4+AY8Y47NgK/HbYYYLs9Dy8ScL8RQa0DT6UL95HqnfuxwoRzyt0
2p7P9Y8MaUO70NxbRuoLbppIpwFS0y/FW5QMf0oj/xp4vHkXIdZtqauzKWdedc0R
qbfQpI3zKox0YceqS/h3Uxf/+GQovkbg0u1vs6UhteUkXwkqEk/n5gYjWRFgGZlL
V1dozognECjYl7PDOuiw6cwzGcYCTts+OvrCrv1SU8zaOvNO7eSwOG8fnoGA3rQu
CE2PahESWVmXIZR62cMmlexXWqLbPwFnK8Ilu4DerwIQrSHeNz6qv63sJtD9UBSp
YZ7CHniyVoHBQSDOK9OfxPfHdKz516I+mD5tRsnbH1scWVa8jE2NwBUSRvdj0faq
lxv1EnZuAXcz4dxLZ7laTc6B8FPIQK4INAZeFWOTa+15yjVnJRbvt2ZYy0cGfF+i
jSfrsLudw6hvboMVm12GmaX1As2dyTAm33G50kyrbqCCrHh1/p9XPHNqp3OOarrj
+VSYvd3vcCW2RN1vsU+nyVjKIuemBeQI31rUYb+LKnOf5At9EZXnkDI0n/Ih5MN3
IzLj8wFvAJPygt03ZxJIHiiAutmL1zRqsrHljuNJ6s7xCw5bD5PGxgyQ7KPLSJQN
0znK99C8/3mU0HTbPzPojqEoXijI3qBm7CmCDR31RedDlqnqiy17Sn59n8IuRhDe
XtGcnYHIVnfZ05ltGmb7MQ==
`protect END_PROTECTED
