`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UF9UHWT1zPByypz3kh+R/lWWBvRoe5sKZO/+OY5OWn+X3laedMEMrIvn7hxMGCS7
MpzBFuHyQ7mAwoXXdBIrUjSZoVqkokwzrnpxdmMZLL70QSbzpwIHUQ/Mbi3YTBQ0
wvV52eW2ZcLl7o+DXrJ/xErmCMHA+dlbCrV9/Lwvf86pEbqN/BPdZ8Sa/rlMue/Y
mgS7QVxscM5iq4sLpJ+8UclZp78lKNmE/+fSNkQ7/jzavEA+dBQSpKT0g2rRIpuk
Rv2M7ML1L+rx2qTRuMWcXRxDnNX+zEiJhAfmoJqLFS/lUeW3+b4TQIvWFue01uzr
D7IhRbQeQ7k55SS6nxvjuAenQv+jf6GYtRmsdDgc+O4R0jHpJ8ekK7z2/YnoynmF
8TtmE+87Ujuth6ItUX4qPLiVLg+SPoPtGbBcVuPELe+vW9XADJ3R2S6+KyCWiY4T
z795OsxBOVXH8AR687HMHXYvU22PdQ8v8GtsexlBrQnFVujamQ3YycYuIxFcpP2e
16M30OUF85U5/lWvMmfRsu5tngQ+fykNi0dt6l+LxaJkcnvL/0oxtLtcE0LTuofT
dkIZu6URkg7ka6qFbkKD/9KFqXOjaxSnd9CilRUOo4RarndwJlXMemT0BOSUWPkE
i6XlnXK3XdsvAnAVTDi2Cw5s3UlElNOHT6xTp1q21OcN2xK/v2PS9KCMYEbo//HW
x9C7IQNPQibp8uaWnEAKE7trHMSl0oo4EDp72oYteGhA0sZ4FICb2ICVSFEk31oZ
JQBJbt7RNarNerJTrt9MBmKBFx15aYujOHrFzWsawiOzB/xXu09JbOhXLBX4i6v0
GtuQCy/zlpkppM3LfZoLeDlQA5AGvnUfR3NGM5IeVx6AhBdp1/MVZz9zSIfzqOhF
JLOP7cFfnrxvKv7vDopdnByXRGgUcGTdx0qLT52kRXqvBYRebzH0vDsSuFnO7lGq
4uQ0KgQCW/I5sSbBM73wGOU1nCjgxKByZhYnEf8SsYf8caJ1gMQIMzGzV7UEpuYb
ffQnNvq90H2Y1JNAbeEtavTtJQ7GFNQGFU+zUnD9jpyctSHE8dlt3KnjATsJ2vAy
DmghVPz5S6zqW8kT7LYPQZDVFs/uX7xPG4IFh6NDycMo0UvKt0l748m4hMpt02Uu
kydItO67SHhP8MFjP8ApzNsRBtbbRM5ngdOf/efdkVzQLHjyKFDncsCpX9cAkZ0a
nQIGqC++uB4uob2gltWzun6/K/O1KPVVFCagJfGqETXIgtsuGtcW1szRCn3LKuPR
As8L7jOUDF41DkdM8d8X2njbLtla3ntOWSl/1uFxEXxY0cgRyjFmYI024C7BxFL7
i4sWWC7eIr74ciS3JzGnDmjECkBktfE8IqAqNYfpAhh568hQyHAEExyrpGwyOMtp
ssStZMcrbfQHFS0TmvyQ/Gjt7iwTzAeYq8PDtfc7gzcCuQo9CGLIJYBLKW9hpHnt
BXFwQeCCPGfA0ByoLw/22eLZNt0NFrGheDECUj5NFGYZ6w83hrJH+ndX16HU0JUY
9oDFcQ9hPfw0ghhPBb8vV1ovtioDOJC0oW9yMXe8JXHyDcJNSNQD4c7UNZ3uZXZl
us7v5P3NnlzSCavF2wCvDtFmRXcqpFdvlc1piiDyHHTUsiljP5HkZ/e8LvrBVVvJ
59BeTQ6vVpubsWuYt1ba+vcuuHOwVrngYX5LbunttV9ndj5Z81tEcyR3yw5ofBgE
jHO9c/w/i3HlWV3bA4p0RPoOlLJ1As/StPmbpslLJSlDEQrX7NqA1lrAjGkdz/fX
NsZ/8eRtMmCii4YPJ/5eDQE+hcahWSB37TopGAtQrNfFrygu3mAFli3kHWX6LBCr
R5lH5j0TT3adSn7Aa8ii0PX13PdoGfe05D8V7NehRoO66snSJ7067nkWvhakTJ8y
VAAMpOm04Tq7vHymKBTMSh8NdK6RSO51AQwWdSUhAssHULTXFLfBbIZLKj5jLwCF
ueIIgGdYBurXSqR/LK2H3DrcfeXSRYY1+zxtHca1PPPgMtYuwPrdOJZtujzd04zf
ytvHOHVADxY9y/O0ym3Ivg+Wf1XwLjrwydLPSIG43D08OSANsSqPGZS9yXLBC0wi
iM7wr/WhUt1FrAeZ47CIRsj9sgISsHGcSUbQUtrtZ27F4OK3yyJs2hM23tDxie13
8V++6ocC+WiJcgU52wEt0DqfPxzyatWQHK510pTRVzg4xH+BACtY84UzYKRP4f2C
6SHTCNAhD9g4oHDDRznwHuqQUaRPoRXdjQpnKoRdwddjyqQE4dHCMQhoHz8qM9HX
oGSZ2nRwgFSN11xHnn1gBynnf5NzxJWrWsiUST4rb87DIrfMLNvJ0wG8qrt6DPgE
4TnaiHVUmgiSp5L4z9fvSVo+gAK1ae4bB9H1ZDr/uNgv2RYkWaFUXBTvSjHsUKoE
PPJcD6f8C80HX4H3/Flg4+uW2Z6pX6nXbB9zOEcQlaq68LRL/DH+qRnOmc2l68eZ
lx6UPlKVmX1NisW1SjKlymARooMx6h5j16+KWUUVR4vii3AgF1KUCjsJQ7aN6/Xs
wmTj1Dg8CJiqEb5bseR37oJDPMnNd7CaAlCTh0YP+xi38ajD0ozIiasDUGL9tPSG
kgHQ7Hcx42T0vtJLHUsPhuGFBPAXQqMpvO0HD8ghxPUotsxSEJychseoCnw/FwWV
tuz6V/94Hx3ffPz2cXcd341eeaxseV87Wqzs5nEM1th6eV5mEj6nbGAk9xOTliAk
Pyp8WmieNE8i4eylAHEWPnzcAjVl4Kh4+/COHjGEjiesynBrvZ+waJPDHlXJW8hj
31Q0o8wl5ig1l8S/jteUtb1UdkSb9WHrsjPyA5mGMKKAtxcVAMIbHn82l7Mc74VB
JO4SIz0fa2ZTP7P3ODHB3CRM2OfG7en/RFjbYg8qfDHxhr/NREdjtEc3w7+TTE4k
hrG25YuxtpmTc2AQ1SLO+l3QILCETVryWF7qPTTtGan/vFN6NJZR5WyoIO+dPvbA
UrSjiCTd/heXSe1KC/wG8uwKLSuIyAs0mn5BgyUvX2LvkfLpoQrneneK8aMaWLsX
idhdoXrqRrmudlQya8xnwzU4uU8Ayz0y9Y8FuYqS4hZRM1/76DNPv7MSDpV1KFJ0
gnSMFNjl2EkZxivuoWK/H0jnavy/85AIXrPH70dPKXeb/+thgBzlUrD0CZhbr4ba
PqahPh+aDAaU9IKhloEPxO2yAthbPmtXI0dwblenlW4qU1hxwqV1yDiDLexm/jBe
yYtjhNBdRz102RtoiOoRIEx9ik0wzo1mKiRbfjrxhGNijiyGwHHnEuZsw82RLiXI
tB7Iy/s/m0AilU71KnvUMdHG/sO90TY17dpWZqtvvu0QBg9Ba6mF6KwLORRcb/1Z
SnIZOOtm3EJrUmrCsHxz3XemBS498OLLwsZcrBnY/KsRwz58rSWJdZ58hZZdYzCd
E+rucnuQxbBn0PtmsCEXjqGHAhW4/C72CpbO0gQ/e78S5R82/9J5Fh1AvozdG/cK
HhKa4ChMtyS9eLufqzzzB3Di0C2JDxE8a4lB7Rl4trp0OYCrc0BZ5qp/BOfymISj
VZtBBfhKdSxaZ6Y+VmGw+D/w1as9Ytn/ZGLR52gB5j7nf2Jf4vu5OgXCJQvVN8Ze
1D3wbaXGvCZZo2qymdaQ6SE7iJ0DVua8J1EVK81VdyaCOgTwixpdETS8g7Rrt9VB
++uVvm7mpWDoEJRQ/lCsedOlXVsR1iL2O0uL0E3vOwrno8KuzvTT5i76KmqA8Ofl
Vnbvz34ZtJqT1t/QPzkuGnRt6uGkmHO1jJV4wgWX0p9zb5clDI/9mWDTsoTcyIK3
p7RBcxrFrqiPOEhGa9GP87yqVv1KFTLsbIdhWSRYpSaE+Ld8EaHxA7iUBaysWNRT
/2in9MuW4GJhh1sPR0MT3t9unvrkEWOczMH8BStTeqTifG6WFMw8Y5q8fPMcrPsX
NyYsKtvKOarIttKOML23x4s6jq0mkL20BeDI1MUbLqZDDHzVjeoBajh2pcnusnYQ
ZHN9oKijs0SHd+eeTbN6krAJowuUo2L0vOkNF6X6koFoy5hpctLALVuLgvJN+a/t
aUmKEuYo6ZmHWX1eBovdAm9CnPw1peAsSWjrE/O/65n9Or214Epz6r+KKUrPh8z+
V3SN1zoQ9RFj2xo7xD+0PMqK4SxMZwZmPU8tuRWqPphwWoE8eDLaeo7kg1rQ6GCN
l10IxDV6XmNZl3ibmnnaNnon3KVPENP6fm9Pjyeg3QFZ2O5GvC0o/aISIcgxx6Ji
4c2VxXTDX0k5J0Os+He/B9viII4gzAguhdozDfgCpRbHL6JbLFCeSBpqA+1VvmmH
9Bmp5SNpTIT9/Yz2d0A7KHcdPdwq9o/GCMktCXDw0sPY0Oh8kqDlcPqf0wSTIDIj
99GBFY8ejoVLnyJoCgrv9bBp0iMLgKsfWADL5Grxrswh7fGIRKX2HKLcOYIG9UqB
pjGP1jczgcczzcJSpdr1B5mg7yxwI4Gh5AHnubjDH7kYcKf5m5lSd6SdDgPeGQld
ZQha4Hbq9d75gTxgA27ahFRo6an1fYjJv9FEWoN0Kz+viFT/cWUUHAZ1JH+9IVXh
8kF6gIeSdqeRo5ByS9LWFoC8npN/W3bWP5gIK93OUaeV43N4K/Mg+Rh5wDKZ47Np
C9nY563xNIkeN3a9S+EGRR6Japy8Ozh3Qe+uvC8Iq+ySycCtEkNKaFwo0xAdFS3G
iCjnKSaUd39McvB6KdEWPgqYKEn0BY91MZX3xPXdCAwXB8S8SDJiiMZu+jer4n8u
afHixIsxsvsnz5rW39Wa3nh153s1AgWc+0jpPQXgVH9B98KdMJblHNIfrnkHVduz
K5VoEi0DDDxS/qZkb5FoRQE6aLE+pOyaEoG6IocRLevUi3WsFa/mhFhm9nlHd5/u
UKOmoLSYI0UFrKmF0+ZsaiaedcVScgh259QKW2zotMuDrf/1cCjEf45VA2ASId7+
zbdV+az9s/e2qFko92yqq4AL7LntlT1tehN83KsUgzUlhxsf0xTTiAMhLSCp7uoi
3YPge5Hn/k1btI450wZolMqLw94aeNcXfs5Cuk+DPQQSrooWPsCGiAZfGuxCvZPY
kYjDEd9CRZ3QYg/59EmP6foYMwyAkqwx36qs8xTxWs9cLV3axZ4sVeL/sAy/y4ch
7gtLAkpBzby6GwiEr80goyhYnVVYosyQvWYyn7dcIS3kbH/9mnf1bCs2nEYac+jS
8DQOp4XGkCu5TSP93Ki6yTnJ/9WH5wMxD3wktSPmDXbdDgQlRbfYrZjOkkJUkfdh
iJ7DyDjXHKhDNvpXOA4Pg9QHVtJ4Gcj9b5WUK78MEJ2Fu6g+6kIb3NiihOQd3mQd
5MEo3qrekWeh7fnE4rKY04z7a0G/EP0NM8tblOIYEbcrTnzp4P9lVppGpNQzTTp/
qwVz2qCB6iW6c2Mkh6AnhHtHXxdbXujPkUk0pIunZJ+sklVSb1MV3euiogin9raj
pWmmxR/DpFn14JoydToxljr2Afj5k11x0R74mw/rYE+jeA46j5S46Oaas9NW5Lfr
g4sQS/WzNhK2hfAEhp24wfUfTC/iNOfG82qr9Rm7QafC/9gggi/Pwz29rkuzJAk+
ljZ1lHZQaLSn35sM2OHdOIfGJv8uv3yUFocbsBmCOxB2bYNeOkI5C5DK80Ju2Jt3
9ZKvHj2oMFJtkVY2Ht+AR2bPOD7u4n1P/yd/yl7RDSIhy5TBl9nMa6vnuE1UECge
T/QjPxAaitlb/S0y7X9H1lxFKQK3UKLNL/fnqDwAgU5FM/s3926XAsAxVACAZQnh
1Og4hRhg4rI+KSygn988v0TAxWs3X88VTX5Cak+ikP+opOyWWWbSqwFIJy76mMGP
vs9b/vmZMa+ytahZNBHbeBJZrBKbzW9IjttVN6Dv766wCHNpbwWLLqduO/vZiDcZ
bNLp7mX7giDsIIa1INMvrK0CIufJInZ+La+yzxhoLF0XJu4xIR00Fcizs/7k1hiY
qoUSghW3Q+o5AUZe7KiQXZARZgi2c6BOQ2vmjqYVYxFl6uC6db92RK3jcNzXrOxC
cFwz3rKuy0dwgcVrjgwbKSSY1OU1md423sH1AYdZDXf3DYzJ/0dykLhXOThLSbZe
+5hxbt9RAWDs4/xgcKfUbh6cG6iy2LgAjdadwF9uqCXLnyiKy3ZvID3VhJrXalaO
E4KEcVarnWlXDlTZE/gCl8Gd7EBG0yHbkdyXURLoiZ7BpWYW93QsuV2lkDizPFSx
KqOuMTpI2oFy7S/RUzMn2zwe7aJ9GrwECgYzMz1a9kdQV3Uz0tMrv7lm1uOak/fC
ag+DXhrgkhp+rimZvHk7ElOm9NUKCfRzK6gSg/EydYNHnIj+eBdTYzscyUfdB3Zl
YiDE4pbgNPuwEkY9cKEj9SmGHV3SNq+D6lGokJGbkLaUx5OmY2EXjuN0WqXD6L5+
IaiEcmy4A3gqevpmjYD/cFTHqCg1j6bB6HvdhGyAzkgB33qdgEn+qEcVNNgxY/n0
kJWjN+InXoNmPNU0BDdZhC6oLtJuYWyBGMoNQwqOO5UrLv0NbX3jQUHSexLUXPwh
g7YtW1E3o/vq/DVuYDJ1kayfhyLd4T/jvm9+I8BJWXZBP1g99y7w4sbZ7HxOI/Z4
q8mPXxf5+FGrIiJ7Bt0eNzUv9z+46T8tS9ABe3SlFYbZQJgU/hJOXfp0se7I8yME
LigQeLM8GfpJFiDujt6RmQb9pVUtSkPx3fo5CsnGmeEwS1gU6OJPVHamr8wsok27
j1INkDsWnsLNVZ2z9d7hJEURQdmWrK2THpRvZJqE5ib3APaEvECZontNyjwWMJKH
SfCAFZnxwpASmDJMH5Uc9GjnVBfqKbaltkWRCG0XJQ+xyRtU9CRVMkiEMjedfo0u
u1raq1WwW50LfKOHKyNLA7FTwm3Vu3JSxH+KJWRwSB8FcDEvo+JZ4WLiQMSs3nln
qMONmlFBGBiS327Oul4coWDGicrLgGF+MBghlsJoGz5dutvkkD2bqh7grQ78N2SJ
U++M2dtAGPhHS0ZCGV5L0Rks2ICdgSlpix5QLRBl39Dmopfm0cL1J2LI6gILwMG4
Eq4wdtSLyXJFGTmoLPQ8cnOJXxVrRzLRVdZGw2/o1UGDRxae+uMMw6LeoTibPwOL
+6IMgSFTLYAyhjWIw8l5u1yeR36YpZ3LKKltCm92J3Mv/iub6B/ZggrZxcNJ4HfJ
o5pcRVk94uwet5XSY8BpWHsDn69P7FkJJNugQ0PRp9lI+xryCjTmwMNaLlCABBRq
yQG0lXp/Cy7X5KilAV5ikLBZHtv2VVCofbjiTfHBp3HDX2GZVBa5PdxOeB0HvIfH
j3bIn6AdSCxoCnQaL5PY8c5xS6y+KrtMyX0m+HC/gi7mqVU7ckStVUUN1A8OrXQv
blNsV3yk/3eHJCJvo/XW7TJtDhsNJUGfpyk39wLL4HHW4C+mFA504Lbs/X8QssYW
jLu2n4l92q39bSfb3xevo56Tm+8vq7Sy8NM3thpLZ0M+sdjVKqdrN2Lb+mVN4UUc
Tk97FX4OfRjXJwQRx35kVtBWsHUtzjIXA4n0RCzV7uYcdcHjPh2hHyr1yD152VQX
AbkAD6w9moqxAqAm3Ye4E4X2cFtzyhWuSTIYzQ6fwD1g2JNqRO0iDYCwdlq78gHl
Qqjd0LNUP1uzdYj3s51069GNv+xY5QfiF7UwCd+NdXxkDhnRVZEFodiX8r8namGs
xPGTIScHxkmnkJTImmjNVWvFnOMEiWqQ08/9V7koHO5LuC/6JU7txAROy8f2Fvkt
8Ff8j5jI3QYrki7X7iPV2UZvH5k4V2f/8lD5Mt28mdDrRqSBPX044PJxbsuxag/i
n2VTMDRz1GtUPG+dATo8iLsmrEacyrsVnTQbzXJ2JFgUtnlzzFa98z41wsmLHkSS
fJ5AwLngd3YPTjKmoyGqnkaqjAIgiGUDUkFNX6v1fg5TiwSuG0san90xiWBRKlu/
JU9ZIpcA18wYhoCT6NX6xNtP1Deip/NgiuvHO26O8WkiL1ztAM8HuVObZSWfTJsP
PHFp4t96fClonwaf75SPiOuxQCS4E6DZiHnsBDwIK1D2jtFsE79ldw2eZOa/FS2Z
tb8p2H0w70Jti974yMMNdJ3oLXHaSdzgUKtKjoZrW+rXEe/ytzvMpI6KDFL2lBI0
JpdceuiJODj923kIETCH+Tv7LTwmi74TRT8ovrtGByEyDln4qsyFolqTh1uZ3TkT
Byuot8NRGqdeJcUSqMzXtNkfE4UNR7nkOpsICagKcpSMfqfBqPcLBUBaWE+DTbs4
vQxeMFhGYaE/UJdbCv5M9iZWtp9GYIIZahXoA0Uy1mKBEFWj6hh9CEKrJJojJmFv
I0NJff/I3f7mJXCSS1sH/f6DQrygFt4dLgGbqXT2KMKNEVFsnE62TH7OsoRyvWkR
Sjm03UyNEwgoYkSWT2VsYYg+E5FE+RA8KRLa0Glg4UFdOmNWzc/6yyGofVPVrYJp
7TDuB2mGhHvBJcLOn55mvWP3vKqr+w6VX1O3EaCrB+D8NQoan8G1SdILpNCmVTY/
JN8sBWVyGdlOQZlVhOsLmdr2eYL/7Oe0XEXxpA08gCEfwGEOX90Z/xNlSXPotENp
AxdlfwI9IPt8fZ+DWliKDATMZLrWqZr1uWYR4+f4mL8Ee2dgd5C5fjby1KKfRc+S
UQzwjHcV0tDlLC7EWZuoPHE5MzJ7kZtZcHEO5ghviGIp96RfcTzqox6Oj8KgXq25
MHoy57kD17E6A3e1gMLi3qd5n0OZeEkLx22/lWphBeCy3CPH1m0lWAVmIA3lv+BD
/siFADkiCIMaz1FvJMzbZ+gkqb3L5J8MMMFLdBSIf3KUcZbB1Mz5RTH90QwZynOq
aqKnp5v2+JjsNh9uk9HrBQmmUxIbK6cpIkgb27AEVJmraUl1+VTpxPfGITI6wY/s
IcT7rz63N4Je8q7svpoEvGRk8vESZQHlvQ9yLhOVAtTW776GFOQS9Oms1GQOwJ2j
lqzEyzN5lYLWKJFMIbGX91KzSaW7YvIEp4MFp+7XFgaDy1MWzsqY1FlOQR0Dhdrk
F7Z408q+Z5I1YjI9cq9J0x0gEY+VvMq2Y9N4RT1JR+Gm6XOS9s3ofHOW48iwCNBA
Wo/MY5cRsijJVTPAM9xLviBgfRsxSFpZ18mix+EabUDO5St4zhJn8jSHw2O20fZD
ZLZBQuIdIBHDGZuj5sBrbj3Ss7f587Ths7ABHjiBa+bTgqQHyH2LoJxvjuJ+XF7P
+at2qUDZdeUby3fZDTZwg66gNAsQF9Kysz0bqs00wwEQ9cjJyZIFldC/sAZRSmhx
u60wGPKzsxf59h0FDCELYhwwkWe0dk1cpUPPHJFXJ0+olpqIEE4rrjIgjNPWNZOc
gvdPCUApRnG2GAKNSJ6kpk8I8uPDKCQAPsGujnQkf8iLM8cK0cVmLKNB9FgJ74WC
zQxd13GTgGHQtjiNXGUE3gFeeJ1Zrh2p4j2SLjsfNxIFWGA1VlMYP4kObLwbqf2Q
rp+4P2BlJWRAWklkBUdbajtxrdi9JWGsqwGCwrngn8t3ZUa8ec1eTaxZjo+1J9uf
u2NG6EXFShg+U75g5QXeEqN/z11bD76t1GFZOl1HIMwx0pf5tPUwK8q4lp5EQV0D
HXVLzoAbeNRUaepbqhVLcjVw8LGbDdAzzLHsavNk67oPV4bJzTYgLvvo++Vc+KGU
86Hk94vAEYRMee7syS3p45bkEPqhCzkPi7iyRMXai4Y7/gtpRE9eogM3B8Uih2sq
D9SF0tRnxqUEl+F31QvD1HUyMMnJaNDcWDxoOyeAaYmblVGtLl49E/tiFPLlTVMs
lwLH83zFCgESFqEpC+VtvCxVTInli9lbkHmjpzmboY8NWweQL8pPeGCDZWddEhiT
HE4Ai1A6iO/LBcnrddRF2/OTFRANHasFEIg0wtU6dsKQw9AxFoju9JPxi6f1wmjO
oU1AhXl89lomK+IFzHS6AD00QiGM75IvgrPuLWOm18nS5pr6efo6uqep2TWdkGDR
zul2RQAgI+iajJ7VgyYRHB70qJho3cy5SG3qhM49L0Nq+e140fYoOw/zYnia/pF0
z8q/PEKzfP18ZDDgRowuWcwfPXq2lZrNzXl8JPiPiygGoekLAoAAZzlk0KGJ0AiZ
IJcrZYaoKoMJfOM6vDUHAvv0oa7+bBXaQJ2attnxQrhIRYuGheFw3Vd/4cZTQzU9
NoOBxhWXSnSdzvAvt7lhr3xshWfaCH/IAeX/Fi1JfFCDn15RKYtLqqKKVFTFC4ya
ROLIYhy/TJLKtuXDO70LLkgUm4EjklXEP7sgY6IBRhqJnjK/FzAjzimgr9Hw6b9h
Jz7r4FNgMC2V8TrJwZgqFpnheSFiCyzE86iUq6Ve9Vq/fbE2KpqVXsI2VzUf73vx
8l+plQXrBxIYUjwabhpmHs5T5Am8zy029UtpUmurFAXPb/qtdyVoGFBSwEegrbaj
EZDIvq0nuhqPwXUdBVx3VsN69350xHLhrcEALU5FajkklTTdas1lhwJyyuZNkJxI
fVtnc1Z2awv4Ev+uDp/PO+z50Lk//TcZJ5TmhaHcoa+KXsaJdhJ8j/VgApiTcXUu
zQjcyC9gDnKgdoFHlyOGbb7XPivqypPVFKiZPUNNaQ00kKnnJ1PP8Ofpe4oLkhmz
iWUW6jtmzXc3S3s1YmmaWe9wcNKvzLxldb0V0oB68ZaeSOtV8b6pl1SF6aPxn/Xc
tKOvBD4K3gLdazUQwGTttk9fZbpznFsmKMyDk1WYSGv1jsCr5gnyu0qE7JuTeP23
8FJIYO719TNl24ZaJonGMKQnkMEkifLWfwK1yuA5/Dy+9Xu6aHreodUfHPAAm6cF
UBK1/SSvYj+z9xLGPwXJtOJTHU7Fx1IrcKE0zwBhdiEt/f9pSxGUwRUa0dk/iPDE
TcVkkyyIkEoMNhCZim7DN0mtU7oKz2bZvCoz89cV3geAy0q+ICGzo6w/cYhi1sNr
Lq5ispjqSdaL25+YCuEBpVfgUzM6BjKK0VoAVdSYmGI/+dM2fYEMIUhDMj75N/wu
/CynZuVQXvjYUjOuvTOeT3c2StshgR10Nya5LivlJdii+P4FEeh3XWaXl4BfEPtX
2H+2uF1dciehwj/NXwQYmg2OvMxoW8QBtJUm/uJEbCSwwUCpWluIw6znbSNx2W1/
Wy1Uw2GeZLSOn5r5ERjG5nHYliq4oMwsHMwqcSl40B1nJMtbZ5hUmqYjVitjWeKu
ZaP+KGP4wf48nJQVD1FqbhKqUAxX1PPoaMRw5a5jZcabo6M9cVA/nCY6n7amZ+Km
kypQQSAlUhkVBNcw7cyhjP4FWrhJGdfgCif5gq1xck/3HpnlowL5aSCHUzpkFzOg
TYEkxV35usW0vK4uE+wjWWWnRL6wIUPYqwfGR3GuDDP/xRyuKbcQ10JgRWfdIrXo
TL3JvNIWKd63wz5mtb1VsvZ5D+0VryxDQMOH9Otai+9QhzSnaEzwdODMgrfnRxqM
v1WXJR4V7ecera8icbNU2IVu/pMUYzohHtbJFMa/Yk7E8bZEovTOk50PWAUu0Pdm
jaSXPKg3JANRgJeh7GBq+CIetiEFJolhjUQsXiZKR0ap0zVzcc+aJCfLwYkB6gnH
PbltkUzkd5pNPK40iclvNULB5W4GAGLaTO/E9MS+vt2kaxO/Mpk9sP0WrjIT/odU
Vg8JYUuEjQAgWm3BNUuKI0aPkkd3aJ0gVLme8B5Usv9RsKy6MwOT9PHFLp+wCbW/
c9xqFzweE0odSVTJsco8RHD60q+lqF1wEXLImd4jbCUA9XeeHTLnDxUyN1GAZuqH
zmHGwVKG6l8fHRR+D1389osGhQ4eqlahEKBtKKkgP7Ue14tdaWQ/Z6dNXrCdQXxg
Fj5Bfw/RCbj9GqM1elG4LZZR6jiLpkmT5aCEG00g7PzOOzCCWIv7Sib3VU2R9+5k
5kjsitNC+LwYeu7/q83tYbHQw8WnTvRb4hXGLiljffVFtIa+PCIm0uhzHrfMMBZa
m9uJncAQ955TJ3FX4COLIBm0vPsnSYULHBbmIzDZjHXJbfXOLI4Npz5RPRmhg8b1
Yz8i2mTbLJ4JR2W9iXiD0XLXlT+iIGWB+SrAne80fU/QJMQjO+suVXAcIu0S2Z3n
yMt294Pnl1+j1kwwFP58LlvLWGPuxoRep/wO3cQcgn6rFniKU6dvwHCbuaS1yVaq
ZQjtOC3i4Ft+6HYd7xF9+R6WOmRfNmPeCBdJqDfN8P6OnfCjuuVX8pyxuJeaJh0t
6CC3onmtE8Co74yGFNLP/eWvwSdg7Sqice5ycuUhGHQBUtQcH2v+8gpYKrAH9Djl
aEMG8X0ByiVYio67pey9Y1oYIZ70ex3DaowWu4WAgry3jIWbGCcG5n7Yi3FNvgoH
6Ou4iBDbWM7Xt2iidmhsoE7aVFwLO0TbETiM5ypZFf+9aiBlTwGNJDoxrfLH21Ea
L6KqrO/TvJtj22VX+wN3jyiB8bPL0AXzrwZZN9N9oHMPSCe0Tu/DVccAUTrw+mPJ
VVzXMHpKQY5V84c0w8x0OBWtlN55FskhqUcps5cKfI3TRSBGqkZThyV9VQV2/DZ5
O/DtkSXPvyiLWQzRQm6V/V8iy2xYU5Wxfl5Ty2hvj4LU/M9LD0ry6wJncwDXsaX1
vDFdVgEWQv1i5W/VFj6I69sW3ynd3pwgD8/ErvsMcR7BIf7WEiw3j/9yiqNYoMIm
q5dmr3D4gMlcnOCy4QRcEHq97GPFuNx3DVCLDGx3cJ5BiZ5F152+vqyLT1o8c3NZ
+1m3Lbf1NRVqwt/53sfeWlDCp+2+18OvvSZNsrhBlyLbHzLpPEaH7J9Muv5GfbQ0
k9XwFWBW7A4BeDkbvqzXMfev9AulOlIHjliLVneQbH4yJguQYshTRMwKJ8hnOckB
14zpACNpDE4y/2x4EMTCDEKXOIZ4FM4ITfry6Eb23j+cwZz1COgJvl4dgBQTHXwG
zBOIXRkztnioqFCoRz24Svn4icjN2nFvADfa8po7QXfEX/yw+vQm8cyN/azY0YeQ
rqsM/ZIy5bZORdjVjIzyJxmUPmSAG5q4tQDr1JVdWfhLZhsMvm55B8/1Y+JC9zEQ
rU/YJwobkFnMT3u8NKrK4FLzpehYHfNCGWqblFMECSnWr9Wpyy7DtD3TPdVJcGQT
7Ei8jZ3HWFFIPK3yQD9XSinxGtAyOiGBhkgw4yz/oPjN30wgBZCjtpP//V0u5F48
+Tau6+gc1JIL8KW5ZxSY5BdJgVVW7164ys8YVOpvuvH8lRTHrV3EnyVjOrY3YinO
8XTZ9z/SPf8yyqpnST0tTtt8VNJSNx4rTDq/GpaEZ+sZ6Ov+w+6+WIp4RNDt8dEr
UC7cX5CE1ee+cc5lmbLfTdpTdQ898dGa5qgHMUo8DFL7YtrvlfPe5zlMdWwCVHWD
5MMdt8Hm9bg6g68GRePqKCaivvrVEwl5OL0whr5q0bMQHbX6MQGrwiH+eXw6lPQl
QlkSRahAVpolLpPCulXaYR7BlU+TD3A+OxxpXmA4aFr/gOmBDP8I7Lk5e8OKfHC8
uVDeiVyPkgbf0OccFX/UsRMnm2EpsFFjiyD7gk0ZSD9Ls7oZayHbw1PTpJK2y06v
JUwrd/SuyO1eOoFu+L6WkrzDh2bwaDxVHWRf8qWI88b/xiga/6NvUMsExQpeqrNG
3BKrSUYUclgM9Zo5LJ/eCCW+T6QmtGXEC/qI8N+ufFmUNabXKAheD/SxmvP94fFd
AyfFWvPqr8cTsLalF92DGKAZsm/zn2983Z6V+e8/VLGwhraQrE73eZdZTzmpzzhE
xuB+cxiba43Tg+0f5i6BYGGNmg/3AZ6D+Y5Tr/L1fSVO8pRQz53fQ2CqJRBfqSuJ
GtENozosQr1m3mxb4hlbquPkPq58SvfhfA77bQeIVoJ67fCgJVnqJRl9bhYy5DWy
A/rNX8biOhEBzGnHn5YJK/OjY2UEXohgto63q1WvdvrmtTVG7tervNkPTf/TcG7d
2eAq9YEDL4mU8Mgbj6auzMC+8hzhKWeHdwIoQM4ymtp961qZcIXGD/Ik578JPpx6
g+w7BdwSt9uMUEiRX/mMFbpL8rLsBpszHwtVulxPP9Jt500DgG7CsxZ4BnjHO1ik
oudu3ZiTcLCwUOJ4IiPSbThXS9H2JEAecDigfU2LT+1jZb8gyYPOw85S+qxTWHIN
2mepvqFaozf/8BbvRmm84PEKyOZqnsJRGBx81Gkavs80q/PE1c/ZvQnmhnoF1LXu
FNnsXSQroMMkPsLRr4BUPLQJjg4HixLxdikD2McltbGpnr3HtOFjC+JUg3I5wYyv
tV7FGpiY/LKw+RZUI3Tg5jtIsJY8OnnWgzPnm/UfIPwNsywZHtwkua6RejOO5d/R
u3VlaP2upcEK7Mlt/yjWyfMoyPvFLEax7x4xYlJbZzEsnsmPHAbIJZLrIZDA/769
pohmkw9QTrZJ3qHPX5hxQCDGHPv4j0bdjZQJUyLVjPY0/nyMW3GcRElmsSCMqIJM
eYdxHKcp2V3OmYUvYjPrA6IY35dkp6TzPdGZDBwrb13rFkPSrwuro7rj6E0HWPYZ
qIIBdImV0sqxtNheprHEC+GMN+hVrVRv+qTrdmGjlIZXhuVBNjOPRocxkOxbd4I9
IIewYTcLi1pem6nbaXxR8KO9L9WcOFj1HSe4O7eHxgR+61IBr4Igvlx3w6TKUfIH
HzcK93fFyvSNREWQYMQw1GPihkP6x4+0mzq0r6cEeia5tZ42YxkHwF4iidwsmiRA
y5XkPxvDpxG/RC5GhT3c6w==
`protect END_PROTECTED
