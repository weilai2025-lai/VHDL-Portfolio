`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60UhqzC1AHjbhIe15zrMUOvH2V9dj6YaAwWxRev1uEwBYQRvkeHeKtfkqJ47EW/Q
ycVgqMQZ1qnZi0C74QoAL8NdBdZyp8AkD9Glhn/iHQ6i5B5FUXn3bQsckDJT4cJr
PWcWFsUn4IPG/WVakEmDMSorvdxvUIZh5Gb9Hvtx+2FIuctbqxc1hpvCYcSy0B5l
+WqDSwAcCQOQSY2lvuWwaZc1VQf3+0y9f0eLlFPE7CgW+g3fDucuEjoqc1rpsinP
DxfM8DGLsVGrnyyfsFugDbXcwQm4XFrstDCrRzvzdKSLA47cIW2gBZPo4e9rPPGz
E9UznDZIICzREzoN6Qvx6sz8tC8BZn0JmKy+4GknIU3UdrIDCneEKeHdgB0zTzs0
oK7cuJ68q3UWqnML/uoz9teEYIxHQCG8UA6kGntvdiKxm/KfkVZp/21aJNkUQ6aV
1kn4jW886gW9CHP6TDvYLaEzjzxBk4osLuSCMIBvxi+R136yI0Vd9kHBIxbrOPvP
J1kKxUCTwBdb2VMFvIvkitdkq+5JJvVDXUGjc7q37/WFLsFweDYj8tpHpF1kjmlY
B7LH1EZgQZmduZ+RlAuR/SBZR87sA4Www8mb1Kf5byZqrHDI92UwzBmzI2u92Jsm
slijaWUGbG9mr+vBzgDaBF7nGryzJIZWLe/uBIrA0LlIoMzBTChsWDVwuO/WzvwC
MsjI1YPeNaQySf+HNu9V8qihl2ZsM+EINwdp115nnjT6umgIECuGOCvxqrBdo7sq
ha7SyStNjR3PUVLXgP2yCn1PorKHBbcMSDVCHHCj1QWxrRPSddFMF9gdrQblI90R
22zOYpDvJYn/mkVB4zBePpxgk82NMPpc/BhmsQZuhEqXmDBGGwVSjS3Pjkg+X1YX
BqpsJ2O9YPzuqR5iZzeA4rHWIuUOCGntIsKdY2l/MeZtOc/13EAZr/k6gM7OyEPI
cdOXc313o7v4OxNuBkjng1Kd+t2nSEMlfl33Cuu1xQHOY+BM7Tvbudiof+CHzcLK
uK/CIBcmMTEvBe4HUYANv5rduMcUHwniv3GNcHIA2m//Jt3QRNtV+CwZQOvcQoEQ
TSad8dAir7v3PWsvyEfAgGu86BUXE9aMhSwzpTXqgNlLYwtcM0gX1+GD33FObZNz
7ok2nA1r/tsW+pDoqQp8I/uqdorbzEruVq6CWVJc5ThunKVEqVMVu2S/LsMOYRDM
vCWY64py3A0Nkc6vnIs9A8J95ESOP/TNxUSg3NfV6i9kC+sshnEDFVkJw+pqTNT9
5dBLBkniXjRSlZJrHzxrbBc/9grevRPMv+3g6J8bjH0M4ZjbcNPQlTtihsopQ2wO
aKxpW4YO41VJbCFXU46ZRX54pnW38pbVTXMACiDGI5883Q4p7D4A5yZyPP98mQgb
Da8/UDOPJKnDASLbzlNegftJNpimokPwSHrlhwOmpnOVF5nrNeq/4YgpijfCwVmG
lubrtWkSFiPMm7XpIt6SCEdiNAVjGbx/PqH6RdxWfSnX3NlGjpDohyw443hGzhds
LIDsFYY9tvFf9DQLM8v2hHu+I2QlhtLZJMeGKXx9p2/roWDoaYEQ9Q4zP+eB55c2
CG9IiClYh7729u7msF1lRey3mEXfja5CU9YAxxi3mlYmABTKNtFHypXNzFizx7x7
HHqyL4ViwjBvjWthDlzRWLQz++Cz6KupO4iNXUCWCOs012rf8yOXXP7lxxcN+2dm
FIs4fULUjNTU6PgH9l8LLpQTdaJfN+JcvjDGNzLL5FshrgjGTNxUD7qLshNhayIR
0qd3ITuSRQ8rYazGxNUunSRMc45xHwEVb/lB42S3vk0aoJ+9zDdZRaUk3wgs/Mh9
1O7cumW2Gn9N1QeNX1ibj8D5r6KrgQnBLiAjVBM87BCZ4CIvXCUYDWRwsE/7DlPu
5NoVroGgaREyJh/hv6+zV2qj+N+AStmf+QmH+32eAvA0u9JYllJUqRwKIAD/MENh
G62UF2sPyAsZiDg1dC7j1uUAzURZ0/FGWJzWdzTvB1wOPQAMVneECsnZjKCmtT0C
xjv6YPhJM+00flahwsBoIfxUdsCJWgLdk/GzcszbFoPUMTU6xYip05gVtvQlas3S
2pL8dLs0dIWvpTncVVDo/KR+083XJB9yXVOndUWD145f+ydCQP6M7RxhzZY/qNhl
JGKrK+jlSmfVsy0CT6p9/Z5u87Ed6sOzdHbfcSG+4F2AAFI7BRciw7HVmbXq4NWP
J6JWV2NEiOCEutQNbS4ztUm6aRzeDkWrOZfUnrwI4yCldg249vB9XzzQXoZBFt9f
5saRiLexO4b6m7hzmWS+K5ZcoDzjEjmlEvec4AO10yjHySb1giIMlh7U4B1VmIv4
bTlEMCjMu5jjPz3XWqosGjNKf1eO5JPjsikhiBHKZ7DjAn2hfpPrtZeEn9IYRaqT
REvKsGjMOmTZVsJXGyWrfTFCjN7X1mwuBBBF5yqOEroEEx1LY/CnkezIk2ubQbbX
tnGflTYNL/OjA8K6TcSunAP/Cwf2LY7qWjQbaluNmRARN0ipHcZe/V/sAF2BdrKl
3fmT8c0Oj6oPBEA3POtrLsX+qSor89koqtZirMNSTdR9+XN0Fz8BGNgQRAWXgiQJ
zKG4qMigVSd7ejW672aNWatxoqM+aWYauT0NMx69/GUNT6BoGioUsLDw3yZFBJv+
OTGYPfyLhKvnGrAE8S/0y8dJkUgCL1eIVseADKk/rfwBHnPFm/5KM36j9nQ0kgYW
bGQ0LpC367qFzTdCjeQCezUOnFdIWpoo/AP0nBa3jsoxkQA0mJoBKuNM7aRQPp+H
+8HVLmA1FAyt53yqI3yHizux3WfR94R/ojxWawrE2juXDxsVzYPdHjSSkQcbExog
plQaMRFTKPsvoWbAVDLK5lfbvoIBdlkTpCupQAUQW383FO+P/iyJb8h1OWzIvXZ2
w1vJK89Up3Gn1mPkhepyZ9fgqTDkB2Bdfbc/LAOJk/+ovkOK1w92/zttYVyKFlI4
yvbfBTr1xaMs1m/AIB2sy2yWDfETEU3NvkRU3EbzamJ6HckqX3g8uY/hFOfKWDyX
cLNbcU9gRvcRg2CbP4SdrYg4/n1YdF3uk4hpVg+yh8zbaD7nIn2lhyNsICe2KpKS
CkAfrmbsRcsPtVQnTtcHZPCwShe/vwomD0laus8vxsQ53nKCkqsczWwpOpuY/9aM
+t8Wpl6XZQM2JJQun/x/sRso+MkWi2S8h4yJVaPg3jvO79chBODtKo69UvLKlipd
BNx50FjfYSQgwJp1ARlx4njLSf3mYrU4TgN7sfIPyj8ivnbpMDOMvaaoeZHAIIRN
wg5H16iYsj63PzKKmNhHj/Mwd11/mwl3EMrG3L5Nj+WXyjQ5ujceghJdahAM5ZfP
hJ/cmAlTj5qeVBzqWLX5Uc6pFgK9AWQD0gLYW4E0q2HgbYst4HdGG3ADSk5Sov2W
8ES6AR6maBC9twhYCE6LtDZzB1KqTxQowp6oIqZt+uQcl+j7DmO26iQnBPGU7dnI
ii00sGkymQXXSPzF4MCLZeCnsmj+q/doX/TBdOrN5sjO5PN8Y+HTzPCOR25A1jG+
lon9eYkWIXaIAuYe5aTCrj57sJaLClT1DfmWlADNnKsBAEqZoz9Ch/tzMjppXOcI
nU/ZdvNcXXUCNNGLyop1pYOuVq/u4zBk5LE7+4c9snRQzjZ7dNolATzB9bdJAvPz
88GVIiBXKs94tXXuzhWc57YdFrGgzx5VA+dZuAh0+a124m97ZAGPcbtAHqDHkat6
VBsw20Ynq5LGeeoHvJYu4Qv3pcOBqm3TlGBfZYzA/7w/cgu2EkfAgvEEPGgmq+Ej
Uyn+utiljss2doCSwTGUBEDqQZSkEq+o0tDeTUfVWStZVLE8N4g98Mbk1/YToqcD
cwGxrb6YRCwfRcx4liw9OmkjpfhuLShJX7UVqvQXujX36H2dat71Qdtcmb+gNNhI
Yc0uQfOJyHGZrvMLXpeGO2KQOvESmAw8AP+E/HUMeKiLiZX+6jayeSbnw9UhmgeZ
cCR2g8nAJg9F5c7/UjxufMHqwHqw/ONW9pDe5CMDGxsOyvx4R/G8Vnii2nVa5W4+
bjIo1cYn1BM2QB7vRguj742GGC8GREGNy5CpYR9eTj4IpAKWT1Zv7J/wqE4GCIvi
PkZe9BEC6Qax5lxPJMowoiyPc2+Oymm2/OwjOmqPOgIelCmU6GhKmSlO8JYqPBPs
TQxePTCTRs4itQC8e/iX56bLLFaoMbJ8/et+I8xeMlciJgZ1EmRlCIPuQC3ROK/J
sLnwT8MHm/nnGW0mdx2mcUY5tVWl3mDAugd9Uk/kYmF/da59l0AvRtOSnvsQuo8U
TkLq4EvMtdXnsH7CPqHacqp7GGLL3J1KLhgOJLXGfiXSTA5yUIZ8jrRPqjEbFAC5
dyvgco0K/ayFZo12rckW9ASRivgw8K27/G19/I/IMvbJj/PxGx7VC4AdJ83BKEOg
oESnLs+shv0GWzz//lDwuUoEVg7gDwMsV8h4dH+kiaoLEXemNpIxJeyi5+BNzubP
XoPR9rGoiaUIpcdaq0RjnunJcP+8oklxLJgDf4BM0sKiEncjgFCp5x77H4hyITet
udblNvfn6zyy+nTk51dIvyGUoCahX1QFzITNZlf2HS6F9om4BFycq+0TTFxM0Nhk
rKSXEXLiUSqW/OOpZViuw1/gH4qz/+Hlmxo3IPqrwWiQF0u2S0Q9bGyvRPS/w8Je
fwrmZ4ct6O6+2tbDuxbUkFoRvJRN1+Lj8z3LkPp1L9wSO3ljBG0zZSbKGAbWxrwr
RuYO6TggvZuad25TZEEUiZlGS503FVKWCbX2QHknjT6hmvIp/3XVyueQxan74EOC
F6W/yaxJ97UTp8VxO1tuAuG67dw07IjbqrdrCEaxKdBREmALJWIL9aPdKS2wi1Oc
uN4aZspedsW5karT2XdSAWbWjckT7V+B+7wmDUOLo1CEfVDY+GgxZs2THlQK3pva
xqfZdQw+zYbHZmoXSc5EzbLSU6C7mhFG+YLSJLeS7f2RiHto7MelVUKaofoEvhn2
4pWgq8M9jIIqyh62GIhWGjBjlYwluKXOfv92rt/lShgEgKxOzdBfpcaLdqFUl5BF
OlHdYgfFc0riWh1TTGl7qtvlqG8hVXtcYsGXxCGmEbOrwjICBkgCUBeFK/5YqG+P
FfoIjSkE1Cu49KEHMTZTJ/SgHOFLUdrDXitJgmbmMj7ms0KCRveK13CTnrEb1VUn
e3qM/SKOXWLpW93k5dY/MKpFiPmVVhmAxalaI9fjIJDrtNxPGN3i/FnaylbGwe+S
3/27IljG/wzmW4HG+puoFx1pXUkFZoQaGkTA2/ayZwQerNc15KZIY7OZ6FCbRo7z
xSSVwrwcbpZ6irjLMgkGCRnqfCs3CCpiT3OErRiqM1B4F/j33/CkFDDLOGx9RGs5
v3/tIew80OalRysPa58zkVRLio81fUQpK5rUl1YxLeRDJuRpSDOTgJXg5O6Ju8Z9
y0K2je2eIRB+tWRXNT6LVyDIN8iTF+lfgDP87ieFX9Pgav/hTxr9aW86TmPc9PPJ
wz8ef+yrWHFmDcjltgGqXUoAvPv2q1xwCQPf3ocjZ/wcvTP9yYgtSKBmmDgH99BA
BW8ES51Ujb3FHIP1DYYWWc+AMIxpHoWEodHgMzjA6PqsmVN/0UQmmAgH0V2KRdLG
JixXKTlI0TsMsK9gegM5ekx6R6ZGZdWO1augqSTydX5R2rjxizLl+QQBA2yiXrR2
8kzTBIbIITybY8rVcD4QXeG+zK0MkE+Iwqc5KDEkaNYUDEzcqvTx/wJrpI9fP7Fl
FWV7I8929bIlr9aLVUX6aEyurzf+TkDFVqGg6yc2Rk7eBEOlGkbhqDZ3bEb+aYJr
Fsj1dr06i3RAomVk4cBu6phePw4tTZmRsaye61/5PA8AfE4e0Uak/gJj5iHJ279+
dmh1tf86Qt3kWynnd2enQy031SiXkz/Emr4KHuKWjA97kxlBXO5juWImpHmBsCQK
WzxOzlLOHdE3HKur29JJ/DGy87QoKNGKVChunwzhModjoBL5XOk0zA38dEc4v6Hf
qk2pvfffT6TEP0Z6j5vAK0KhLwPR6lozDo2QK1pOZJVHAbuZAGWVTb7c7D/ybE4L
jivGmpWg/IWyQMysRs8DeTA1UMzL5UVCOxVUrMs2B+SEIKefaAsoditxr2cNmm1n
rItr/T5Jr/evgr1EJHUL4pVyP9WSmawst+QLMVPXIPhRBaobrp4ryk4THb8m2bGB
f2aKUQbclkl4jIDxtL5Yt1q2an4N0z9c1z77AVOoRb3vbY9gPo7o8vV71Wuk6ujz
QJU+/7553sXWlf7sddzN30/0c/Qtd9mkmx5d7Hz2AVZKc/Ui0VXqsD+kbxAnr9A0
Z5OTqkgtbigbLakdQbk0TAHo/IHPoTcoRUTaT9Dcoylfgk0UsY8CO+z55ix32v4Z
nHylTgLOt2n1kUP+sGiAqp+UQtPoQUSVVE/xPSDLFCR4Sm7N3h8/ZlldBZLR5KYl
jtQ9GLcf4gotj9ZRoIUWmFqLRE+mUmKOcs9Ukiy4NKU3oI1ccxaySTVrAnfCX5Gg
0hrFniNKZGhkDYs6fEHMKPwNA3pvGKIr4kpCKfujZsWVpQ+nJjF/vwsViu25VRgX
`protect END_PROTECTED
