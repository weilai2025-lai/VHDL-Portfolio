`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pI4j0bmz+RoA/eugFIubySPUmddA0a17+C9Rcwp7HsgI0HBsI3kNzPrdwaaIlMqt
w3RjLnq6WKV94PhWeZv3G0FzF+wMWkLcAsvbcAEDDDhDbaf+d4DBDCFOl1b7PZDx
NGscco3sIWXMfX2wXQs9qBQYu/mBgw6pK/V3to4smOMJZRLQQDse2e62WHbXkHbp
KreBl0JxEmMIdmRXNsYxsRDkhxSlvYYGvywHjunEMBJIoMGHcSN17Vb1zOoCM9Vv
fhip1dOczmFFlCCUGBonzAfwJc1MZF94zUjOpHD78wOwrJnfjtkIKzVu4IQFb7tT
LIW0aoRaJfU4PeocOPV+q0PizdkMIsZn+ldtnvZbB3MYpRku2vsS9XBaIPVFCJS2
E2OER3Z2OP0pe3BVuzHhoA5Clu0S3rGYhsWImcjj3GqTm4n2y/EJu+TPQ0vgcbfk
SkyxbFeXPUE1ckzyVf8TkOaXjAWJ+P71CGfmNXpFFXxxcZzCDkxwbH8RT6o51rOM
73GwsBh/ZA0cSEX8DH2LwYqyPXRMW0NX4220W3FF8jKQ6CdQ7vP6eUg3ifuNpxwo
LrogBVZb3AYSNdwNHFG6/iHGQazubw25VOmKVSDOETU4YHaYxoKI1gkE+pCIUGQW
nOpSRczp90nTjUtRGvZsx+8OmNIoOjDzEK7OebQ+TUJZD05JDkI5Mfc1R3P3+Qo5
19N8JR63HYWvWAuWkqOZgJuqI0uN7YKVcvT07eTatlN5xmHf9MoHPOEcKXwLSlcg
AFplOpwrH2R/rz2m7318E6pX4ZGLAbHzzR7jWU1/7SXvfM+aVYGR6EJ0d4i4TFQc
jIw6mmHaWqFAdvTGlAtSeMq9ucp9slEAl1LgOmUcxrc2cA+qabzgIlURaia1pNrr
0tDL9kc2lWn+Bkr2OzqpFRZJ4Nksv/C6CVM3i96+iQjPaFB2NUOxEG+KkJMlDdJ+
bGOpgIjbAPHciAfZ3R5g6XatSDFhysLL4Q6JXx7h5uh0Ahw/XZ5eDkM7W3r5VuyE
rThzlmG1Ur963doks0+37L+E+sDxjg25lLb1Lmug3PiQ31CZwbYcfXtNcuWXRjmO
qR09JzUOeoRuyZY73DQ/JhZbFg85YHe8zKMEPhkxVnM+2NSzDmts1IJEPs888puS
Yn/IXlukGnMwwaM+pL/elcO2VeFdtLW8mZcQf5rRvQXoD1huWdUTuxRMjHCXvplC
KQ+k7PrHsZfPsvbKXdO94QTEJXR92BNF46PVpHocFdRBDNCkRLAHfC14XlwKw2QW
CjZEQmPmM/46D00KB9gRWxDxJPH/5ex9ZoJBKepZH0+NAxFNgaz69c/kcaFbbnDP
m4nqPrkiCG9p85DNp296Ujeujr74l0uHqQD4tRUy5qayWI7CYa/coD88oLJ2zV62
XK4cw/BaMdmBx7aQnXMWD7XhKNKZOi4AZQUxub608VCzQEcjTUD3L7KroArIGhX6
j4Cdafn765fS22CjDXHMZZuWA/TrBEuxIAWnDS586RtP+WESHdtzLXTNXRpd09pe
vUuEwgNVq9Rih18sG5GIekquhQWNB2KRLbvDxwej8ib0deZJjcQcGCJWiXwacfKB
42LSKQQ032cFe8tJRfc2jH2UGTrbBU/lGens9o1N6t1CDv3QjjaqLeTxwIYeFoug
ZHHo8skI6VkGfT8VkRThNO2MjBQzLlcCXajhSxlFlztRvwFNEY1Zf4gcLneSE9zO
Jfx+uCmpvA2HsFRKELKAN6U4fVsSWG0NxkdtdAwhMiz9K5asFMrWiCoJkRrS4y8r
NQErxGW3knetmE0NQCM8SKwSPZadzUyM019K3FUAHmBHOYR/UybXLJf4HWWsJVoG
ilGwj5zm5o+mesbZLcwkZEr1o0T/JfVQeQze4EHr7nWwxkVQtF4rSQdz41Vd4onI
544czPqLJpgcWo7q1skf086h9u7kBOi+WSIA7XMMcPEM3IOjD05qkKfmRLdiVrkL
xomAPYIjvdL1nWPisBmAImtfLLy/SWBAgIirEdGU8/hTeSYgvRNU4h+IV9Ryt9YZ
mu1DpTsuOcATxTd+01ZkcnyxTi7/q5SdXKD+hW+1cZgyRRo71Q/RVSpB38hHjbix
tBT3+itr11Yu0pXtR6OMBLadEdryPlhzrppnijLn7qXtIrvlwC0ghVdyCA8LdC61
hMOz2Y2eiPAJlKlkoEKbB5aEZURB1xHdXXaBn8DZ2NwRpqQxfPl+AlFvxdY8vv6h
qCqQKzpqyc/aemw+hFRkomgBLHI/HP+rgx6h++M5aQWIhvdIGwgcj1bM1/0BJ88a
hs9Hi2JcbVYh7KkrNizf/kX8eOfuKwDEzb/ykCQevYDN/jkHzhvZ5bru5vBVxvqG
gq4lNm3qmyFB9x5JrlkTM7lW4xIU1fPS3D1SfkF8lj9b6REaVHZEIz6bxzw8dWlG
K4Zw2Fp5w7iX+TdrIJLPalotq1catXykiNFbmbe27B6+NyvBWa9OGvq3bdZLSV8L
S2xh+6J15rZusnZpDmXW1nf2GGA0/eruHSM+Y6+heOBGka5VSNaqB9cB3sKAuqkn
qtHhijiefmmVSalFrWS9Ny2/9md4+UIr1fO6up7V3ow1rXzC+D/VXB9HmtezGQ/3
H1O6Cq+4LOxdGx0zo1m/SigUyFNCDnJr2+uVxRIYdrGPSWetT+Gh2+X+5SOYh6Eb
EcAkmokDfqDyq3e/N0m488Ht27I7oxlCNKe7YkC6cpaJ6PDDDdRqZE9t5IDtnSI+
RP9w4Prl8zGGoUGyX6Wu2kKLOfuxNvDlUNyM5pSoP8M7wh26AajDIyKsQ2zoUNmy
D+TnHt4mXyk5mhDIKW2qqwQrUnUwiOWQqxnlk9jR0XoNuGxq4U0Kglx7KUa9cisj
gEC4V3QicztRltXfNVWE9j1lbXT79zzgkG/n5uvkVLsbmmwEYqGyOvaE27+K9pC5
J8ez8ZRUdHjfrI3sKUN4zOuP3Iq547BcEkXF72vK5ct4ZyKA9mtmCkFE5UjCeLk0
NFTZ7P4zyOHdu3TchbpQd3qthsMWzoarXmiUYJWnInrzdRO0RXRXPgtSTRuwpDpA
rv7LkiJuJmkoyPFsnyQM1JhzHV3h343TPnJbLLAciT+Y9+36tD+rIcl0pt8wlgIP
2CKOwAQnMvL03eHeIcLiMsxT0by0riYhXHqiv+JfJ0+CHhMFXgzyj49alFNW7Ohi
xXU3PHR+yrdKfwVPmLX/ynUhIRcEJT6UbaMPOm/TTeobif/yQuFsIrZ8h7FrwLB7
1sUmIO0jImperGSH//n5rUbxbhBA0sKKpNxVspL5Ts9PZHq193acTCDF10MRzgUX
V5IzBYB1a2Yj9FB3D4KgOYrzO4zI7tmpkekL1ecnceFOCARay8NWe/1ovwoE+Dhe
vcdHqgGI2Zj7tBuIqh4zoWSWLY7/xGsj/QRK3US5+7WMlOgr3etmE08QzbQMc5B2
X5s8jUWMy7IJlEfWHdm2GOGBOIgI0Bv3qD3XDf7U4ycBItIOtRYqQjgOHX0b6CUZ
hVf52AYUf8+3/msjQv9JOn0D33qqz0OF8Bj4mmZNfkDWzv3JxE2ugHyYO97syRzU
pOQOYM7F+FcXlLcR3x4hPQwiwILWeLf1GOiQbqh8BM2inXSxu7Yn7YaN/LptlbFu
nlxK94lkawKK3hkRFsbpNE5n78zFlxZcs2EYk7D5DHQfZkXhgicIkAlBgn8x4aG3
MgunGvIEnCoR3Tx1J3QQCVODbumcPZUSuri85SaEVwMBKt6wAdSbJ+CNVAB9A+TI
A7yO27GPsKtuakNx7Lt7Ozooen5PRN+W2PFaxZZt+bGnAtPZ6S+riQNm0PZW28Bu
iYhlKaehPZU0dTFooh00ltBrYCvgHgeCqvrfBMlzYDQaFdrgTwF2hlQSRym21X+u
KHs4+zaYgzGRr6+ECwTFb7JET6Frdw24xvB2ioqeZt6Dhhwqh10OKGbr1Xva5VpM
SuwupiwmLpcrfcAkdyTj5XoPPM+pEoa3v9XyGXrAlN2UxvrxtsrP1zS6pw/FN/1y
DdpR5Au7NOCUPmjWuEVKLzMWT0TyBTQS0jHkmJLB1MDrfIxR7UgQAFZhZIEkDug0
zDybmsDk71BgzXMNLTsC8znlUnVxZ+YtymN0HMA1QCI3l/u/5gTwH4W4SW4lztZC
AA891xx1i/FIG3DrxfNfJvCjgT1cqy5SRouyVT0Av4uYwHABP1HZCWqJjTy7zFUK
8KAOBAkAfEqOtGC78pa7dfgW9fSjhMZ/FFInaDHRsU5MK80EzTBhW0UK6rpi0Fie
XlF0ovrHHX9qRDPrBjeEY0p+q8OA4B/fAi6Xv+q6l4ktYy5O8UTJyPQjD7/v6Y/P
JSW7F56u0DtBZB8+5i+8K1EqtpaLlE6XcQh/PMzH8XBrPOCBrogM7glM7ysqDKQw
FkCbstkwE/Lcnc24yRSVv118brGvJbKFbntDPyiD2m9GRBUjQPxi2Ua+u2dGtvLh
VllLwqWxKcYr00GHrce3BSSYjTd6PiyaqBYjUR1EZTGykZYlpYsHJAS+UekuGm+3
15Kcj5ePKyRxTwtZTs5QlwjucjrsELoj/Lj8UKvRCMLqUO21tx3NSPHx5WuXeHEy
Eq/Kl6hEivY1ZfWuoiUss+Upmeh1QGHiw509WRfaZMws0zgvATcwmz7I9RueXP1G
iNBuFjQOT4FpH51Rh2/SwueIMwaH12CvbKvJ6up1sLeH7OljlI5OkB1mNCYK8JEy
DmMNia0WWLeTkmi2cGFp0LyQvl4A6Nm+lwA81uOBZJFHUhDG/bsVwGF60WFWs87n
OS6MKIc/27DgsxcPxzOY8ZnFa7N/QMuiubxicSfhQkHRbspaJGMttVzzhHADXrxe
VkKyXdH0DeW/mVRVizX0li4JIXqz6r0jWvWbFrJr7sv0EyhV1N3Vfc+JTusLYd0e
ZnLdflx+Oqnd3oSCwE3c5nr5P7k5XXa/ot4nkLEfyzJzvWW3vaCWW4jewDgPXahq
TkyMoqA1uFQMwg262JGnSEVnk2h8+Po3YnrfPhxZU8Tcm0WcO2K2+W1G7PMPmexy
mwXVTZGIpXc7/LbkOsw38amVgkrdnNzyuMh0dI9jeso1OzJ0X4ZknsPQUwUhvhRP
GLH46mrtiv4Jn1ItCwY+u0fLfCLJ0UQBZ+m76nTCQxDlCxUJaYgsRgJTgrTEOOod
CR6kd0q2bUSD90YWhz6dyQ3fAqQOPM7WsjZKBj4GWqrZYHEfYx10f3eo3lH5wK/J
uM1RaHBh2w1O4cI//hpEEVrGsgVRZWMICFxibsYMn2eWuhWJfcONHyFK6O9NSQrk
W+TYWzvi2qMPO0JZsJpx/035LQg2i6p2ecdKuMqziduoihVLiN3nqitvG3l2Yzfi
SCAed0X9PZDAa4L+wmaypSN+4TAdFQ0ot20LVr3KV0pLGJGvobAyjfZsGmwxIjoN
iS68iCHbow8SZfl7H+GBhrcHCT7IsMxR1bM37HBXmv9j163DhmIv3hTzQXUU5gaG
/WXBOuPyEkPpvTvko/g05ee669EkLlKSkb4+fvfaENXNG9VF2JkpSeSQblI/ZlT0
vzvZcvQB2Ym22NHXVtroJBjCnd8KsMV38XuanL7K9jahn+0SukhluoZQ86juW2ET
xV5dHM8UXUs/8ssF5RodurOiNpgV2LLMmizVAOejHCNAR8cGFBx6idCRXt0ylDQy
CqnTYrz3cdit2p/7segSMismyfL2Har2Z6psp9Yip5bQ09tvh5DfuQkner21W099
YiK7gz8AFIVh/WrP2XBg64kaRnUu9mMr2nojHq9rixd+SZiI0doAC3wzapICwH9Q
EEDBBbBDB/T0O6F1cOEffMbmBW7hRI6Z1NqQNqTUcPgUAR4cgfmixrjMPyKsLqNT
3D7kxUeStKSH04hEA5fj5PkDZLwcaYEOq05Qo9H842yC1tN2yIluazg3YNHqpjPD
rVppx5ffuDs76oBd8SsuuzJ739jN4OCCTvKItBKe+ooqoL5RFlYwIoCd0/ufcnBk
sV463NkzwOkk346WTONw7FoUg0LkaXq0gl8KFj9WHlWX3O4tkMV7bqRPvIZj9V8G
ogsJ70ixmINHYFBhpk1yVOkxk+MLMuMdXdP9UQqPyISZqwjhZgIGbZwvjDxFe9JD
r+QguMVWVLMGnwC6hkWOORR0TyPQgRG5DgveZM9Cn7EVkkXs7Qw/k4kFFDiAi6ff
5tuWUXB6zEj311hwXcaqtGsj9IBCx7ajef8bwlhxevq5gCX7kpE2DoHZzz1/Egvf
cs+nGPn1MjpaUst6uRjW+XStCPOShk93nr8crxgiimBGOnZtLAnfZjwLz9mK75ES
siBIAzf33GGXfVjw8Oahg+Tahsr79ifkPk5sffi66p3DGyJsHohRp8UwZbAlEM/o
GWymWYK8a7hdix0H0SJZOcn/Gx0HXKJIwicY47i9+nL1KLTDYW0+YCRwHVMS7Tsz
THkhTQhLdt8GH1kE+47pwBKVNb2dBprLKH2u38vyU2DUjQIYwytwNPMb6/q5vfQL
rzoGVFMykxXewvwBUNv2EwawHRK2N7vcXKFpUDjACks40rGqcZ8s6fD0X+tRjmtV
vVaMjzGrbzFYol0nK6nrt4FgByvuzldEY3aGv2KnxjyexBSDDpErFxe/1N6fTBZ2
ftxUaMe3LG5XVLuLN6GnaFh6lJEW45uFLk7plFMZDZ+5z9aWTDyEiOZfqwDLYrvd
k/CfiC7cVLf5Jciovr5hiMiQSn4ACqyiTi7ZnYpN+/JIteiQP7ymuYlaHbShtmim
JnrmN4hl19KF5c+IYSobAAdbHNwu+QBrYJnJS7FDvvlR9S3KZq1+w6jn0HoNSF7V
hyAjlsY9vSzOIfSJQKV71plJ/vPGgDmbxLPQZo8diTji8Gq9yIO2kNtD8uJ5Z0yC
e8uOzs44QDTZ2VQIjv9Vm8MQE2i4UcRTwiVvNaUqbKOKhSzx4Tvi07CL8A7ZlZFn
lbZsYyugydLMbZfzClFhOVpbOCnDMNLhs32qC4Bbng/XkL3BjKbmkV2jWImaLUAp
x0wsmE+04EaHhx6uPGesCZpwqJXRZcjZ7l9FjJqxsocFfOFcERPMokuRJp47jH+q
ijd2gSjkTIvpoOK3yBJo457U2Iec1atTFb8Xtb/loQ5VhVdIWT7RcCmAuptiCnTZ
VH393gVfl0u7lxI9DY+NtGH1sz+N0nXussAn8xX5IMXiA2sihJO2tOWqNd8Cvk2J
yC9377RA3YDDSYzncWVguIlSDfXJmmK9JPAkN4rvTQSIlzS1fTmYy4NRS9yYUL85
FVSmaln/zbUFqGRc7O92SG5gLUn4RvZSU9JDdBvk46dlltSZV0X19VJKpxifB04n
pulsVJXi2XSEvk8v8CvwgpW8WOpKUuIpk7DiQwYz93S1Ust+Z+kzZ/X1milJFBuk
7F5RyNa7lTx5f3QiMnbwJu4bodNF9EWdPckD+D4IqpFo90BtlY4wZVlZxI2GoilN
P7D15U4hRCvzRzSrEORCbVL+OZlcp7Q6Awnb1YyMqAGkUXAeZ/9e4rO6pEcdFCOI
qCD5ToZOyukaSCRh77l4oW7mfmVRFsh4lE6LdyJYjCDdM3b+JwNXGdLESVWA2XZ2
y4ppVD/ZQWsEdl77ynXoPh6kPxzXGrr4DEklar4ISvEqzCvXC8LvIfmER7YXm2wl
JC2WL2LuKDP0Kk4vCJ+dW3cvxj+/s8NxHy5Itrs1DTlBLAwROgV5TD9aOErJzVIy
hb4b6Zcw+lbm8BS8YM9vHGxjqnI0pUEo6rlGUOzQDrA9O3yCrOMHSXINidAinFvf
wmJoSVcd87fZ6+/Deuxx/dB86OJtgfZO4fPdLqMuRXO5hIBpsnAq0DuD2lNFxl7P
CD/6bEPBJfbLfpm7Ae9zoZaLdsDAldAzm+Jb9pnFaHVGbp3z9ryMG63vDR+Yh8Z0
10C5ysyInQ3QHK1s9jy6rqT8URZV+aTntSUPEMs2Tw3pG5mod2Zz+/Q2sG3iasyj
0V95M2oBt/RkCxNQ64PdIJoLHhry9KIjrpSc7frZszYtm3s/GWsKRe4bgWFjvQ53
98EOoDPHgqBnHwu33tDXMxiW6WygchwhiDBAONTJ8oyq/zlWAPfxVRllyjPIedpm
rvb8FzyCpitLXU1896dbtd5Iqf676tBnmDZqEoYsVpPy2Df58IoKtt2Q5nnAh4D1
taEoQom0/TLhzA1qqgE/T8LhmSgysC4cg4Jc1J/fhD9EU8uHUPQdk6c3yq1WPS7T
K6Rft2viSjpQwMReLtz5lhK2y9RWt10g5LrIjYJ2S89o3Q7uSBm1tm6TQ/c5DQvO
0MdxoR28xjwGa5L3K870mJu2CHoEt6r0b2rHyyvbh7DZVM7YhTpKTPSCGg8tx2/Y
uphE6IfYCXuWh0/kF4vZmbyehGCS0TNmPvdG6c1jKQvTVRY3bXtl918ikCm0TZi6
5cQ3qCtFOt1k05eHGK8Pdgy1k/jLGzMhK7UL7XohW1cLt9ZqJ87FWkVZ8ybgi+Qs
rj4bu64rcdMMPVwNU+9djN7YU/q4GuT5ofa6VqdYkwfpyw4pmbzbaTgShmj9+Zfp
g10nt0nEvkcmfWUetpMY1DtAbClShZERka/fAW6QHu4DmtX1NWd/TYtlu+8p/t/6
YTvkrYOPpSDYPkvkN5GRbTEUlt2ORXjFTtlW6XMoM9+PPaYCASVcgfKSkAsanj+G
GzEJZRvboetrOhKxn6ROZlGr4iVW7obduZ9znr4LZ3jJbEUTe1xFAc2VDq2Kyych
tEtEZEpSZeBRVh9bMK7ezcAGocKi2qfdlyJX9xn2wecLKUGQ5p9pek/JRtTi6wcQ
TFhRiHe35/gXa3wpXSV+8KyZ/6X+hY24bQCK1YVjIEv/NL3bgAukXjT4Anyom6RR
X4N7lTrJLoaWmsaBnoXauPScMadoT4/KPKCRRBauQ283m/vpk+DbVwTwrHfI3xfu
O87JfZEWIZ0CfsUkwRTXFMrM/iBz0AdKc3ZWTlg2QSD9mQc/koLrnq1VY4hjrZAE
rpR8zZvxPwM4DpjGJXTTytZwfjdOuBn+jDUSSzRyvg2sbVK7PzaRV/Cnr78AK2IW
ciqrLCUlM6oBBreAqFnVQesealPvLYRhGkuZcSQt2CmAIGC/QqnbQSOYolk3ZwVU
q/Xh6iGNMLWVQsvVsbBunwvKH67rYCb8mbySpRzpfcaXDpwcVyb1Hcu402Q8OhhJ
xc7iAgMrBPnGFAwiSCWlJnQ/gDGgL6lgiT05gAew0cNhDGaJV3ftsXhJWvYFVAou
JLv+hVKds+KwtvvaGZFWrAKy9GFz93grbHfyt49tmmbUrYHjPdkdHNKD5bqOymRS
tDnwfdO1gX1jKX3pyKMqnWQFrXNPK82bZbCILzlpodMoCvloHTFgFWSE7WrAhIJ9
0BPc6byq75w2LZz4XNa02TEJ1xKnWObFkRvTM7+obBTwsiJAJ3wmKpOfTGTT5GCd
HIRtjlAjrr6q93v7tYWUDBn377Rn/iwtemW6iHuY9mpfP6KIoHyIQNB9Y5ifrqvg
Vr557SqJbmXWSHBaYD5uZjfiZDP1MPuOywZRIYbiv2EQCeDRRlgVjtEE6J2CZKGa
FU3rDyq6q9x6ai9VerObbFIpcV7O34f2gpVeoJgl7LGaXWyJOpqEb+Np+blfOZxg
uU+ngNWaMZQLikBenM2LHd1sUZoPPwd8dVOEdW1g8bjLyziJuDJhEV71oSkyzUcf
0dTSEr95+VHmnLCX0gZKLWrBsdk6uazMZxBZa280DLe4QPGdaHUB6ov32rQFUPzz
Rh+zwvKt5qffx+PLIMSv6CalhjfXuj5q7dc5pxMUO0bdJrKhtoMjhbOz8dKZezIp
D+r/wmD8kxBpOmS3iw+wByVtMIZUUyLVwpBbp5XT9Nu4BwZEQTvl+hVIdjmpto9p
QadepUwAwSH+AhzJJfKIUOzhHWCGzIy681qqoEd0kBQQwCV34GVUbwsKyeVJXZ29
XWNb+17k/rCWhFFEbF32zPF0gTSGx0Cu8+SvNknRVQfx+j0/HP0Aei+2SW/dAaaG
rKXMcgJdnIkZzFMZRpc1QOk2WwQ7Gm7RzshSqemX2zzk8dxX9rgajiYO0F9LNQze
MCgsIHRTSLwKzF6JCUT5ohxI11HfTAFWq61ZtAgYxNM/fZglHO6uaNW2gkXfzHV1
TEyiRNlzD2Zsr9l3s7z46oZLTA9qAzB31PG2IyO7VvZKA1HGCP6uFPCO++dg+QdQ
RHQ4j157eYiGqBPO7UyVR9ktAI9uyAuSU8IHudG7B5AlmUSaoDHYbJJxUuSeIPEP
qf9dcksJvE94ph4LZFciuER8az9oGGKMnJlTsEa5WvjH5wT3gek+d0YZ2MUCJxVr
JJt/tpMT5HjP9Wpm8vgcgsWYU9FTMAdAl+RVK7t7teGlRVMlbkBMVKiPiDQoHAUl
C1GcpN/LbJy/bo12Xq89mkq+lStKyKA2CzwclvPQdLN/7RYrOSDdsMgdXwc+3gr1
Mowvv50AWWOiC4RF5bYQD761XUbaFYvGA/Kg1mNGq0nVfjcGWhblmgovWRaZ3r2C
zzKpsVFbtToMk3dNkGI5dr/9+M6FnXLCFM+cU3W5bFXMXVRpLp1mRFSPwaIxuPwb
ZXhkulJ18KpzwccEslPu/oX/LVENO2Y+JbflMe1rYFdLRf8G3s8ZuaPltD8V12Rt
3mV+xTe8eP5kj4b9mCBCMatDvY3AWABJqDcOCq2fc3ydUvQ5UXGPDXI6XUbHbeeD
QnGx4scsYovc6WnBdapNS2JcYNMjrVIyInAXZKCMKBacfobExOaIJLqBF0AmsDux
1/ukQj7o4i98to55CAUrZ5Un+Kmq+nmxCevkHbiaOL4ebON4ymBxHQz0w1frmFvW
u0e76eI8EAHGp1n+FqktEuZB7vCEigx11d6ajMwztRgWVOqZoJxMEbsyY7CCvRPW
ugiTGV7v8ilWF2LtpmS7eijNyOMx8hvb9tsqg7KSC6RNybzzFjMTQVAfBnlPaLo7
NYdf7j+HXM27nwVAdOf3reqJ80nvwHGbC5S0HPIHSfwPrFNuM7LwQetnp9cAd/fu
9xNMwjBk8j/gFI8RsI9vCMSu0w6Lh/XJ0/2di0WUqW8FSyQ/+b6voGncgfqjVg2s
bVSXg7kjUdk4a2NeD19sPxBP9SSAjWMzJK06aucELGMeD6JwduXwhQaUrH9iEJ5G
rbM+gb1vBoppzrygUckJvMqC8ibyxSDRTtsCsij6OZ1GUHAKFsBZvw3EC86tumHc
ZzTfx7IamX7j7tnnhPVYEz/oyGyj2NjzBnS/qUJHfhoFPPIkYx19B52S55Hw6Pka
adxb3azOZBLGV7KCQIledGovCvfdFa/ljeaGEFyksyUTVvUosN4uaw48EISopVVU
zT9YtVGLcPaVmeCmNugZ/xx92Wbem4cPr4ZQpPTjrj8UV+IqK0hH45++43Ht8MGq
+NmmZy9aNCbZZGzov259JrOXf+smb4DnDWUPXbgd5Il7AztGOJlMumzwCEvVoI8F
qogvNbT0SvbDLT58lO5tCLN6vx5oIMnJ/v2uJsYYigrkJIz36BpFlVCoArZOP75r
HoJXAg1ucfYbv18x2rqIX7ChLkl97srV+Dd5C/ozz8N0VUluFOcIOHOjYHj78Qog
NjMQY+APU+msXbEmgSgGPfJ+OD9nJGpd6oWnt/lbtx+91mWeHeW4WU1fAaWYZfE1
WpAu6SbGMUYQwgeW99M60Vw3laS1g6yeJ1oUQBpOWuKRS0uIG4iNbPej3qsuGXV9
5X7NV3LvDNE3NS1MScjNcHFLvcCc7WRz4K1kfTeORJ1So/dl6iYXsfQNBa1OK/Q+
Uda04Sk6PgREeHlgpP6hBt4/Pmv+25tZpw8mo9qefOTa2p35MWeWfy+3icBYJnLD
VHKSW/98g3uI3NKMTR7z4U+QhqyCaPzWWAbm4StmoBNgC1NHVIvyrGDLiZhA0Lt9
8erCysm0aoQTIxXX3rTBEE4WJiJgvf5rZfa9PB4P0oAUwsYzYmp0+EgoRYBNRSJ7
D4ttp+tiY9WK5fviwCt5Ia7Fe5ZhHouPd3myhR1+6pMSjh4WZfYLcWC9sqROyCAW
5aSHbgD3JAneITp0xiEbZRfDbg5Oanwfp7q/CvExPGe3vA4PuJmNzTZzI7iaqU2s
a4haCTPdfH+B1WlQQIvbk4G14pr7TFKl5oyHk1xrjAR9GDcvCBHoGPyFD3MgkJEy
eglt9sN+w3C/yPmI3pcR8hExm8YhqvfQbvDMwZtHkq68YMfuy4lcHDeFh3Xo7AgI
GU5930pHqFozpAh8zHD9vMPCPqlx+2y69j/5jBdlbZ/3KmqUFTl2K1A3wyZJ9xLO
4a3yLRslLnasD20GYVkeGUYQpdhOqb1lLUa7p+/Q9CMh0aVnsiJ+3ELEHpM+WyXd
9aD1JLpD4IZVHOmuyLQKXBK9+xvVfic3eG0nIfMOh2CZgehss6tvBDUdwIq/4PNi
uJPxz8/8m/u4746PPF0smBs/uB146RibIdZTYF9+n2kEeHFhHK6L+iuDH5hjBDyI
E51+JoJCKScJ/JCIzA5oDH8LzCMR+InT6z8EvvlL8jKVI+6/YuUlKZsnkQ7zAvqN
7FU/iqXyVUduVmTNEX2kSFn+++kteeoxGYeHWkfqHhe7dZxWIGndM4g5veD43e2V
DzMtDjOkYcqZm7b1RaqkBKS+BcZhpudqw0V5OFxGR2wF888YZvqLr9uviqpqDVTe
7PIMcqffGI5A0W/umC1ArWTa9ldNW9UpbgKLqzsr+1u2R6v46ro5Q3S2F5g2hJ5R
h2e2ClLTZzYkGzRz/txkSSJDV6ViKoBXJA3G6D/jo1fiEpocETcwYT+KqBrhtqfm
+hjTvSQGMxrhasppfTM9Rt5u99Ym3D7m1WEPtMjaHy30azHRk3s+Ck4wFLaCw8Tl
RGy7yKwdnmsS4RqCpjH7UK9wQc2QWWf22/PnGVWojVf51MSEqsn0iOBeoVGW+SkJ
FiiLze+RuBcDdPRAUNpm38Q/LxNtgi+LCkr1sywldRu/so+cQSERU0BB0Qp27zrh
I9Qa9YlobEYiMFmKoeYLYue1d9f1UVj5yTgkcDBBqAmBmCyA8ZbRIVJmKh+f1uWk
3Ivgw0aeNdnmrrQ9MqUI2ZVBG2XroXGVvoApMjrsOXjuUUFhQXBnPFiVz65RoSOQ
`protect END_PROTECTED
