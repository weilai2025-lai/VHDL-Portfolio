`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfcfzexM0gtFHIX2Q4jN02wuFdagCQHjTcF2vzIiFjLadQHAUDEsvQGMC478Tm8Z
VR/+yR+zfHOnyqtS6/JyN08Ay4Qh1hEaWrfi2gGrPGbLn0vx1O9YDZPacCfBr2Th
6IPRCCCyVXlURoxeCW/UYcfyZJq9JoEtVNUwn2v9eSlrprWjVWvehorwHGbUpcKG
NHmmhQQj88DrUeuvoO9xvHmtCxivdrHFFOPjC7YLsLI2CJ8TSlJyXk1LToejUeUU
L4mBhC4bUj3xnE3i436MJt5EwHJtvVuDUNYjzj8eB9etMTCTZ1etfZpMp+4u1Qlu
DuBJviXy9x/wqjIvuC8Ww29V2R6Xv5FPi6SdBH4PhhAcIzJUqARsAEZM5wxGbETr
UrMTwSm5pcLekgQpu/JhSLY6HZjocJ+2hmAF2TSSof+IZBqJS7EEfUTj8/sFZ1xK
WyYpzqWSgFHugOLQBHsXxVfAZrN8wfutPYZi+X1zd11DrqYon2SuyVikaHHuchtj
cUeNXIDwlBFqhMRaYC4CSMy4XJXEE3rL265pcyXCBPSj1SmtWreWu7P65DdPYJyy
1g1tAfrv7d8qUzRgd92NNTB/jDcHok28wYcsFR5vHwMTVwyUispuVoCEUsaUwVnp
qmXuyJrxE9ThpCTgZ/QQX/KT8ZGBBm+vRrPJgESKqOVru+LdP2nz4ryFlEVBB07p
n0/NSRg4CadElQ5fZy2QGOHkB4CUqKCu+U14e3igoE9uWejtWHmRZDZPWR/DJfwp
N/JODfoQh6I2vh/7srWoOl65AxLgDM6M4bgb5ZOWv4WFjTqljk/Y7DrogEH2SC/t
ibL3SW830OculzTyoxuBIJjIDZvbIS9xPDvtaRrbY4nNdJx8W7uo0EQmPgnmVViK
pB46rZ3XWIv78bOFgZ9gJRV75pi2WXA9ApHIBgy1K8xtwwmLpCcqnT2Y786pSQWW
TkUVmGqiKsu4sbx2vP/k2Vqk4dinqwAlbT10NFGx0fBSFl21VIX4fGEypziptEyQ
5Ekkgnid4gIXQlnE5Z5e1szjnLchfm/EoOoa1hBx4HQbEtvh4k8mMqLKibmv92Uo
XtIfngpdWzB29lyxfD8QdNHowI5/+yvURWWofnHnTi/FZCK3IxNVRXwjSonEQoQ4
ZdooIl4YB6a5NMDBWHZXI5MJ9zscZrizVfXVfv5sQv5MukRaGMqNaQllZywBYWG3
4QopvC4l0ecle0itbyl6yy95BsAktc5/LswG6BKzK5m/pqEBUVIvvtaNOcV9fvcN
fZWSZeRZxVXm4uCJhykBaVrShDRsopMQOnDksJeyICGzW0cWQE7qH70kN1aNG1WX
lfB3RjZu6aQo7mbMHGJzQ/P0/42Io5yePHFu5lK5cwHV3uylX03S8ZlqnejYexee
eIlF0G/ekKWcmqvMjPzPUgvhzXI28SxfR06dl3Ci1efN1l3WW9rY+qmae/0W0plU
cN7ERFoGIHoqO4G5gVfbQEqWK2TSv32O0pp2ZHLI5pj/4V7F4QHNIvpTYj1pxRxz
Gdclwyr4yr6/nfPMW85HE08IYfrjjNJS1/As1l6xyJb2Em9DbYDl5pjgHNFahn2l
3JBhoUcUjYySnO43Os+M/mQenpC8kuqLXlcDM5qz4N773C2bQ48tKZckyE2K/IPE
cVyO6aHfDQ1wyTy2oehb4hBgNZGr5+frZc5Sn1H7VwdvqJ7/2j6iwhrLHC44/DlN
XwnVcWPwRLgUW2o8dF4pNlwADa120w+bhF4vuYifNZZ7GHDaT0MNyXvpwPF7VQf1
5b3G/hg1GmQyKC8vVSJFky8Kh3WEpFePJmigivKyXcOf5omlNs0M4X6v7+p8dy/P
qmHIK4dmIQcHrL0C26ksCXZuz0cCTXVE6vSjujnBw6Ma0FvNsUMsAwkqsclwoDyQ
V8Bl89iIAVWiiofLOhchHbQnH/L7kwp51+KS/txurIJ6A0qu+kc0kP+h7xSQ3Wgo
dAHVoTTR4pDeYCJqrWNhIo4JtZx0nMW96A5AL/D9xFlOVyhw1qmvt2gTJODQE2hV
nZ1OzYVkDnnxmZazsCD3CHqHqVVHFdk6EUVUN0Ee7nuWDd4i288pNpjTmbV0h/TX
baQFjlvO5Sg57yqmssP4GOAv9RQCUgHVZ/D8Z4GmHYdXwO9leA2vPPDO8ErMhTdW
cGAe68kL0105tNvrZzLZwtwt9NnSDVduO73hGTgYRa60PInbJPFFfVXb6i+oWwcN
U7GPSk0RcSbzcWTIuNYXvZMh+uK6Xh00ohpSB6obc9cI4KP7No9NhY5VB4nRKfdx
2VSIkVCIdj79NzlSWg5ska4WqFZ3kdh3DL4zkmsRR4MoH8qqrXagNNEo910CRjh/
s89QnkYWEDiPcDHr1BAh0Mj2syGs/rNf3GpQSQhasRMaF8nnapAzG3WKB7kpwkyo
S6r57lJcr9eNRMQeUvN1xWVbAac5ZJbXuz4ZikePUv5LFoePcdk+yjp6RXjQwcbJ
y+T8LK0zjf4XHiGI+Uz0EwQVXE26skqiI9H78FnYd2nyyNVW8wGlZ0dpxbi/btNe
qb4b4iNYWkDaOFk/FMgTHlrxEULWENqSYowVAYqYFlkUP6wdT/UJoym7RYgvXy9x
h/wSkPy8jQfaDZSyd89cxBmbzGcEqGMliJx/Apzk3vl7PKUWb8znLsEL1n0L/lj2
/IlONd9kAxG4nX5CoaAQadZ+ke719Yxr/zdU2etmgcBICIIA35wK1BsLWEpmscfn
LuyXXMpfEuXkxYSajf32IwGjvk5V8HOscuyrDHcrb7gXSAHUeR1LGoaz44QKGXpa
fYHStvmprFx00qx+h98TWLqSPKDramGdMEwkpcBgaMEtGio+caAdXdgC1P6+hIeq
k+2uTuK/rb5kycKJktvCgoaeiSZdhmTU6epVtetsJ/1Smy3oNJgIYzl7cnHT5lea
EkLlii2l4hoNqL5k/cCEaZSxVYFbILxuyAub63C3wPpKWPyKwzVvBbl6/ea6BZHP
CfG68p8DDrUtH+fV8CgdmJkNoIQ/hOKW3Wp/U6IOKKJ6YsI9tLSinUcCWHM3NL7h
74SLsdpphHU16Cc2rxfHlCDqKb+KhV0EXw+ckTHSL1ZZ40HfJBW2bDZaLWsLbgvw
0AOy1u+0tsn594YVnrO7a9bWZ6NVimBJc/CLLmO0AFmrdUlZONT/oaSA4LcTuLhw
zADs2E7wezC4cLOfP1oYb8nDg3flrzv+EGJiHo0lAxSFf3KJL9Hn2N+Elg9ihyiI
fgaCECwLXt3eYyDHf1rGlFh4S32id4E2KeHJkYGivbrdD/tUU9xIL1vOCfILy10L
ol+B9id16Jr2KcqzPa+gvJ56m8/Vd9CEL+Sw3K6lDGm/1+F4HfxLlX4tv+HwdB41
zZC+V6ez3eT2DYguGp7mxASTAK+nadipgsIFrVbLaK9cYZBD1zPgOKpnRsD+9oEG
JLwTU6IlXD1EoEbrnqAtAVJD+uSMvbpdj1VPHpzNu3s=
`protect END_PROTECTED
