`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkWzb1Ov81XPa1uQXqkjy0hFxf/inUyHNFs2I8CCx1CZhnLF5ZWOHx0pR4OPQg9R
NF0eH3n2oz82z9cKhcrlwXM9hXu6+ScRqJm/fZO8G95W6yJZCStB7bOcJ0oPA396
P/lmrAZueMMTrHpv2paidmBEs7Ed3eYjGJsogseyHfLlLwYv3toib9u7KZqzCSr8
gfBG2C7e68WtheHhjvfFkPm1gcbzCEm05q+ahmLxLGpxcNxb5WvX1hR/dW++yxe/
auMNYXS9wm6jRw6rCHEamedKbPh1WqOajCTZmD9Hxq7YD//vdeRD+vHGDvQFxMbw
WbPp254jO0rR8D5ftzPUdrxKBxAv0s45k8w6L3phCKMau20MvyP63rHKvxkZnF4o
B5htQm7zzjTA224cob8DTPMZFr77wnDNo4NQ83xXi5/Ml/L95RoyEOCJlnGbzkMq
RHwD7V10bxUNhf2A8+UrBR5HUEWvg5lUkTVYpKiaq/fZWGAdm0n/vekgn+knT8M8
Rezamf53aWEpk6GlJrkUaj0Gc3HIwTJKQ2IpAixgrI3Wc2z5u5jtDcyzCkPNkvLP
y4ZvGoFOKYzzDstRO5e12m1U4oxLkU5Yu2FEp5QS0ZgtaEWq7Ji4LppLNVzm4JC4
prfiWolIJfcFEXWXF+niiyxS0MegDyeyWDd+CBrz4io9Y+3CkuF5Jrhngf+YpmVO
U/PukRkPpU+TpiEV2t4hTG3Vtx7b5icw+wxUYiGetX5UZF5WmNvIQhJOO/ZYwVmd
MJfSPbYAkbjAWEusmttzkZgcon/g3e8QeBsfAPjiVcWkL3fLrInyMQdlwsJ08D1k
LvrRwj7b3byaq2nUl8ha5FMx6OsZPPt3aflSM93Rk9qYgEvkTylD3T0w2isyhoBM
BB4i+kEm6Ir8BeDogMAmtT8GTRTFCEXsp9ybh+1pWQEFQFQxZNrUTQj9Q5gcUiR1
wQj8zzYi0jbG9HT2bJBjzeFJIbEzUkU4aTIMsmJ9rZwMT59q/+Xr4AzqCGHX6x1f
VfHZvUe8Xb5bzDgZf4VpnA+CkdCFmB/JFIbxYK1ryQjr84k1hhdmUrFqngfU3I6L
IulsUTb7xU12Tfecrlhx4czXHfNhfJIaYnJG69hqHkk=
`protect END_PROTECTED
