`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wnCWvxqV6RPfc6eaq408Ir5yUGILuzluZHWpfBeL/TzKO4vMszjJo0cB/kF6Tt5U
ngnC9uC4ReY5xFRngquiLLNbc3Sf/3cuauhXW9d1z/aOn6DdLgc7rVRS1sWmEeZ2
4br3IGHa5omjjm3iKlXrht32MzSavS+zj8VESYgTpPLcNFUkpTQoLON+dvvZIo/j
v/D9Uro7O8AHE1i+H2DTmcS7ltVIRiIPA924QcUb+LDOa19AbS6FKh5gnTGfD0RX
WEPrnv2n04tEnr46Y0C2UrvDlDf+dG0Fwyf64A6CugNCflyzsx9u/8lS6czoVLAb
rFkxgVyz0sUcyAQIDJ053BBCgsSAUqYWEXgB3/9XvLejYsKgzFTu1pLgcyBRR5Hu
lfU0p5Vu7vhEpD09DI9GR0tzdoDfnCpX+XrroQy57r2l+eB/MijeKxrCcbxrTq0s
qdkO/pEIcsuEryAny6362YEYgThUKf+E4CfCAaBIDO7tfaKenib/SCbs96FxhwaJ
nTlTNyS70F68lDCcBWmHKsbScsxxlB3oz4mn7cAIbrM/V2Nb2p9t8hbRnHI6Xn1q
q35ZB+1FTbn8CJKI0iasVXYLdqpjF2m96zzrUxIyzAxg7RQWoJRk4DD1tlImoEXf
uJKeDoxwSujWAToCQhJyEo4sqEtBSSfghqgKlkWs7mkrQ8FaOGaM2kviK08Q6rnA
RWESvy5jrcxgSHlqNFB4NVMJZZfF0clnXNzj5Ln7uavnucZlP9IxqFwXkIKRYJai
dl2caBTfM3lzrE4D1Ij2WJIHk2OMQfF566OhTVNHN1OyKJn1aUwlTWuo5uzhxoqq
fgxbtOf/unsffkB7IgFgbcuCTyeY3nwFaoCfW/Y+zE8voW/YNTyRCqI1t1UcE5xm
1/hiQRB0pJEZbcyd+7zJsZIDxcWsF0c5aglMzPkTqMQv8xyPPowUKfbWPKEsx0n1
RaRDM+yDHr0YkZThPk83d94iMMiaQz2Dt/VcMdWkrqFnNA7GiPtdQ8PLBbkRbmrg
6PCrlf6J62PQpsvDXYVj5Hu2tAcMr4KxgKSGFd//ZVWEJvpu58hwQoDrOLrd4ss2
SsNOIqxnzqUMX8O/bGATLsZvxF83jRZ068TEEAjly+oeAEGDgX6Qhft4f0BtBIaE
sTYFNKBTQgRNjBLrLFNCengaMN3rb7J1AP68e9skVl4Lwzx35hZUwW9rgoE6tYYB
CDAEAxuaeET6ZD5X/B3RNPAoyDXimWoMSLPvAwSUca8JQGHMDYvCzHW/5EaX9FA8
fiRJ095yjb31JKt9q8Pd7I4rjfXU4vl6zwyYmOFmZmWZ4/tiBETDbCs4m2dGPWIH
epiJlEvL1Om/AE90+kkOb8oXbieHBCivrdPMisX9JWH25AJvknHhZ7JXnq2W8cMi
Qg0CE9uS+MpQ47jC0l4tmF0sAcLABMP/5WWQo35AvL6SWyDATMoLu1OO7Irj0OVT
cVLKHyB8pqUNpnisD4lbygBdhCRddt//hj3Uzi1Ge4fzZOqamvu7WKMQih0gBl0s
ciMyVUvZOGnBh/qnjsyl3SIZiKWx5yqYq4/Jmne4wCWfeG5E4ZYnCoJ5WbR0RANP
5SfxJ27txtoffn9BmEzOARuqV1g41jJXY+GK4KCCEW1AATblxoduOLnrJBlPKRz4
4Ce4VjI/Typbdrv4/r0BpNbWa8hwgZ29dNytAudwxl9jmJ+VAFtBXQMonKfNxyES
K7ZmXCr6DymWuTKPWX4pr6F4OuYwSch9Eu887ThWWXEqXj1494QjJLoGg4b6KV78
hqPiVNIvJ4fNBgQ1K85it1he76Vr4kcamHtqpvTfIoBWTnnjIFbCw+k+VaLXmpuq
8egOhazglb+HEe5fhgyxC9RZSrgzFSvmISw6kvN8zAOTj11eBqPusnTEeG2SiPIH
vK1VhdBVDpdp4J00P90FtJ2JeoFAGMMH2dRuM7LqVs6Ncw2RKotuK7ZJ0Ri7y40i
g3e4wSmIQP5Em7J8M+YHM7yMJJVzoe+yV+fJwen4Y1GsaQgVZ/cR68DriuNmQ4yl
oK04LVTms41RQXcbr9VxsFLDdzvBe/BA7Fkf10S26nmJ8BefbyRxKBobT+n7L2iK
vsQbYKS16VYtTODnkpID+f6vrlpTcSc1ERIS+l8k18w07xYKajJL9NV80TYElrRP
l3a7OA5pS5HjBz7lcREc5FrsN6wxinFQpembv6tV0P8Z3+rO30XP173dH30D1/UM
+v8woe+0c/2Od3t4l2R0NhEO3YSldFq6N0Z/yFKUg7suKpC5Izu4N+kS3qIrWhlx
Hn4w2fV1r+4iaVRIrt6ABw9T1Z+V6WjqMOEaXFu3LTlO1okWs0TwhZEz3jIGI7Nn
lbHi9T6jALG0h6ppKNzYvUUvId0crc2xKMxu/8sx1qjEHRDrokrh/DJXBWaXJcUB
K8ibbWucz0CZk98FvytU7hNwdwZZPFFCUo9P4hhatItmAKXWF8biGlPfw26ZIbK+
HORdqt63mPBWREkm1PNfFp6ubSkJCK9TyOiUoCuqlqLM+W/hw21Z1r/gt/E9/NHg
oNJWnLoA3JVcaFwyA08iU63zVLka1DQxHwCit2sxQGng35sMUQgUxfpkVOBh3FKC
gt/zM3veNovO7JXeS43BuAsueCGHqi7cTyzTreffeamXCgXCj6CRXbSCJSNJMyMj
e9C5n22Unt0lFLG/NEM6AxAJaqsJg03Z1hwOusFVpZi75uHb2SFVLyqznFO+JDW5
ZQKmLX0ZQh7IP7LjoFVPtzuUzPeDr0WLLGz7REFZEmp81KUpDHaQ9AQ41Az21QCo
jNFMNqjUWhXfVjmmTKjSe8/wzYiukHc352AcmH1cHbitJ7TZ4iiItmRH6/5mH9WJ
kGEy6cyx2hYr9LdGW/uvCUvidwOoJAEFKKRi0n0UWQEsKa/bzFuyCj2myLLcEe1f
WBQ/4grvQs4O11JdRfNpfhr2OuZ59l6cMAclhpzA8/0Df+Xleb5FwTn4AisosCZJ
dQgfDh+aTNrdONcLc2XsLru7Z2tKvZqiD9jxv18Cmx99uQfBCIaaXZAxAXdLezcl
/aqq2RWUueQKmvPpSTAgBMuf9Sa6dk4u53cvAAVQCAPM0fW0AJ/o8cs3V9AaQtXA
Gu2JeURCAQkYxt2XfCgtHQ44rcx1vG9s5f3C7JLemDVENnvap0NEz72hHznxGRPC
sQ4y/0IHmEsPRLo+WegCCtsfu2lCZvwm1XjbPONnm9r3r7GRwZiYcoliN/IROYEO
sBvZOc9i47cZVrgthzggHQgwn8uOX0LD0gKSpphG1wU5yPzvpOfAY2f8ARBlcur1
wljsFQZUCVVSkgRC/y7jtS3olTVjDAvDGQ+/gyJ9NpWX2Rxik9KkYd6UP8bPyfZI
v5+EmF4ZueafkXetL+Lu/IoL5y/VMGZT1P/4TGdmOEr2KWIlT2FKAbsz+r0QwxbE
IXmq2s+kAZMzv8JZZlbq4I5TlSUTsXjMmgBunTvtCkBnGXc/eBjrlaoNxu2A4uR9
tTwO0MfMPjLstVfYn6+6z02sn6KWQ2PPmdP/O2DmjcFCnb3N/k/hIBBFmFJuXOIv
Ltfw8OMMcTSaj0dryNCnuV/xi7KJ5UjcMYlMwETL8HQxwFbuV/IM+HQBQIeRbS/f
xnLtl1zem3Okm8bIyLJz75hxkb4pvR6ZpzIVjoEzfV6t0ZmErC5wTwPzmvbAHZ2U
1UpcecmvpJrZGc5ufY8/OBRLkJJsj0PBO0KW7elsPNX02ogKYIr2jwNtvj7jyf5z
8cW8OPj/xLZ+2BJNtvLTwcVUt5DI+CJX+sz8dmLSlQxWUhBR4xiGbLUe0Ld85qsr
TDW1DAr6gOFyZZjKRVaXVfFVhg1hWx6yRf+bc7ZxY9pGHoZv5QrppmLG4v5Ff8Xy
W6kvrkx1AydXPON3f5rxH8YVLaF7IB2ClKF17a9pc9QpuTsoKp478wxOyyHU+iF2
woiXiYXIG7uSOEvNnvo1a2FYhLQteJkcfV0/9TkK9XpARo/0kJqyXvr26tTVTb5u
c0DvVEhpyXBSaPL1LJgRd1JIx8WMicoQVEEdMP091czqx/eccspwfBhnjvFKmFT5
3xUSWfoB7WrY+co3+B1+cZ5bBCtQZ1fwfCsGnKt+KUX++oaPpgF1ICdLyA+na630
2pPf3ts1q/9+Ky5lXPqerO5JLIKf5HQy2qFN6B9DTA8VATGRAPjUJ+Qj6XbSt7bs
BC/xwVM2iuVUSysMyMS6oVCRSdKaJ4Yk9nfddfo3GbtMtfEG2OKmaBkQ7kCCYQBI
mDHpZrkuQLMTc6+OGBXoldYF/OMvYJOynaNYtgm6GT+LTnoY7hv/jhdUj0RdoncM
5nuv4QW+jLzNAcTyox8urRpnookxxaQiNIVplEZJ9+2Zuedic7yLfIqrwGzWE0Nh
aDEKTevAwTADeARqlMcMPIl5WfT2vdPCqb/4/kWnkeLf6hUIpKqpxf9MTk5UIBsY
D/gG9swjFLh+YkyutmxuIKmzWz2OQyUhTCEJDrz1TdfMTeY7D9C5NhYavqJiV//9
6avurz8kQSur0mI6CJTFAWCBEpu7ZiYGQ1vtNMM3H2dPdC9LN0nS/2XN524k4qNU
Uk6zQkXSqx6pVdjXDsuu9Eitc5z6TlBEp9UPqf/bBTBnelIMWIJO5WHfdQND+tAD
FZDD0MqtZ/bi6K8/zUeV/T6pugZ8YVT6brdGeyvxJhgV+wU/wPqerWOoq3DwzZ0S
q8HRvJ/mIZ6PRn4+cztiyPhQB6J8b1iIsh1COZRAf11MkKLWM//4FSSqmuIXHSSV
So2MqLkvaltFUhj15Rm175mNPVXnncKSwbpGXwzZR8AX+j7cLhXnHg2jN7E+1Agl
pAMX9f2o8JbOM1hs8iMM3HpKquv0gyFx17IkhyjHMPkhVdGrM6HKL4GkM/eMLwUO
0jxHxcuqaXgP6sfITPeJb6vW5fzU/IIt2bTz3kH3EeY5aIS4gV7OmLpLwcDDm0ov
DPNhR/BQoklUYKW/f6XyGUrNoUUFRsjBgtQKtex8nw6C2SR8rmBqqygY3TlzpjSc
EnB4AQCKqYjgSZHZE5o1s0EfxEYIce1+eC5UYd/uj04gKxJKvvJ5LHdyagJuoZGx
kf5MiEn4B135Cb6sI3a8nZECRHcW41Oe6224ajpt+CqroWtw969CTo2AksjsR8n7
vhTqobe78gB+NG9c7GORR/AfXsh5dQbZOtqjzwZ4WfsYOrwrMHboHTJtRfYqw+7a
HZXVtnoTyiYSL2SjOS0d21Yao7j6+DzEH1SkKvcV+3svIwUj1OO9sPf5RQSymYNO
VvnZgYgHfMrWYJ5GfKv0PgJP6jOrjoYf9x/1m/GUgYH59n04c2P6ZUqp/kDKPPbL
GCfriJHeEl+jdaaq8fYw8xB+E+1PjtdM3DjN0xd4/VZxvltAXUpyUL/LmcGZXpsK
P5+PdlFMzbilKMJgH72rOatdSOjeZSmzw8WXaOpRQe2J26tlSKELZ9MTGhGAepIJ
XvJw2p15hWV03l+NDL7A8NPdl5YM8TLR6ARJ7NBapBsM+ksIOKjha+79aunWEIjG
oEVzWAeMF1NBrhTrndqF9VaQpUZDjcM5Qj2OrBqZVyBWwZ7kMzUBzYM8s5NQC05v
XcADBOWVPtE4Xz0VrpMsBfZEsPF+FvOiDpx75blqrb//D2UikNY6zdA5+7yXndYV
7uTB9vbrzKBAadAod8ddFBMJAzQOEJmdY1X3+vwzkfyrWuFRAlv7e/9JdV04Z9Fp
dy9TnLL3j7KcJ7cJYDFGK2avB+hY63YOcgmT0be5vKDFCUoc0kMwck1uW+FOOZtV
h2X1E5PL/ljEhoCgAvP5LpWhRNL94TSNv2EGO9Jx76KORSpJU/QhouSjMr3KWKV9
sYGn4fXTHthFQXvSAafcZTZ4Ll6SN0jNh63xY4m/ebkWpWvkz7O9EqHCegENl564
1bAlS4aIDU0pc96vcU4YGqAN+j6hTvgTbVQUMLyTtIBquDlVS3QSYUqncmgObkma
SvUf1MS1K+q75dwBpYkHoja5cv/obvHEiH/l+hQ/JYCiKLWkft82zOoBGTBMtZeT
`protect END_PROTECTED
