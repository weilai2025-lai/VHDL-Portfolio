`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZIYc9rJ/KQVcvPfO42i3JLH/0fEZEnRfmVeHkivRR/AquB0GIHKG61Rh75J1IyT
aMqo5te+hNO+yWd++i5NDf8J43tAJ/5hDSLHgMxM0lOmja5Rj/DXLrz1nMFlWiqn
89Ifl/hckTmSda+Ps3xvv2mmKO+pt0P/TnsFGqUwVcH5OOp9oDFB9JDwZazSZUiK
gzH7hrsl7/12st2tt+z/6V8bemqmMHSINRwo4jA8mYv+SbAuFAHPZBbtvz8gTDvG
4s9h8zPooxNc+Sh2xhteqSXyMTl9VeiGvxVWm9oEZb6HfjqA6uElZR2+w6GEmQ9T
yW3wY8F32d0kuFTNYUq9+ELfES+4kcQysUx7zyxeF2S9GoiBRs5oKktWZ3P6WX1n
29xd67DeK6yPPTFobkB+k17PJwUWNIr0JcYjjJ12v5DlEsKo8zhmL7TipKgvb/Cs
BGZeVHGHDCcFXQWPbJgvmshkT/iIH0LBucvV/95veiA9VdOkUEC3PZk07duUdnPK
Qd9pqOIXMnHKS1BD3VmmNcUuqTarHmN5m5ZnY08YQHmx8B86Aj5JtAQYrQ6iFf3x
VY2FQq0CqzHvj/bTXmUqIkuI5LXBuoieB3BxcSCp4F5o8U8o/wMppjpsn8CKmT/n
ou0NuhYeQp2Qnbkwal2TmSvI5J11idUVSzSpVWIBX51B+SOjdcH6HSPbAmuWyjC7
abfA9ZBcifyu6kicp8Ba/RKvVgmIA+cM6XNKccTyEqf0CSeGFJzRF+akzV51GYL/
LU/GSHRXbV4EGnSwGo2E+mSrrgmRdGZSdVZtQC4qB4DVf/L0zRmttr3LC91It8jM
KNyeCG1BJxRIyVTC1iD9aMJFT2P2upmlrkCcVN+JNbv7oxtWvsUOx/sQMyNpMTXa
`protect END_PROTECTED
