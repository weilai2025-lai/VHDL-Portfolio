`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uw9utKzJVKNlpfYh/EtYnlPfPsaCXaLnaEAC0E4u/ayYDxbSl5QdOaGlWpb5ynt0
b+0QjHkRkQ7JT2TJJWnMFA31PrtDk2P8BdvPc5aTRwbncFf3POPU+SpIyBIEEcNQ
3GOb5XUwYFK1G5/k8m7jdp2iRFnSVg9sknlgXT8RUjvc9x+B8NJy8LTsV96UhvWW
6UoZQVvdmqRcn7T6txcd47CZwpaDgBOZ3BI86mmDddPtutg4eH64Bwx9UhsAa+qn
cAOFMtgKZmvk0yrkTkOOupFQ4KApJf+OtIRCCYR/DXoLXQNt7PHAbmSgzp0CI/Nd
gqyskb9rymI5d0AaoJHrt0nyWd2r4biqGFfDRirmUyum0MYGxvTYuWv1iVJnLUJ2
fRIWLKwd0SLVFJIWtHr2goCyZdEJZFfYX9KUBpVzOxg+io0wgSZy6F0eJ2tHGEtG
3c+aLrm79oIFUV+O/ymyypmoMaVvla1Du+dNMyyc1PHScgZFfBQR36V9bV2uBxtK
is7C17GQPGaXxSNYoEF5YIsxW1ehgCBMJLTiiRDy+m8Z2Wcf3yXZGgt93SSnzDBJ
3L1gGgsnt0MOxl02bCIruokfkIDPD13qiZkUCVWEVee0r8aJExIX3cZpnHW9XdYz
8+ZuNUsq0U5G4IpvXd8swAtxM51XLMG4kK9rNkHlXIW0VIOjOLadONfursvgNg4F
fHHfcw0rDDQCY2oUUNTEhdlBrAhOfgVD3ncxvgp1kVZDk85qYPt4PC7HrsPvhu7q
qDaQ/D4uZwi/aVBmUVVS2Vrj8Uf6ZH57+MXkTeXU/wwKoVa+mU8xE67em0n01Qxq
TRGQ0lIuGJqiJTYO1sDVWqiqEXvqQ81kild/jzpAXux3cssc/cMbeOVRPOon18ar
O62efVUrMFsuK9/uUrFGz7KAuvXGroGgNR/TppTOngjrDQlpCsgrL8aIjlEMcZyT
OOJJfNWOZpHgHt75UIcaGvTbr5Yv2wUWiW3zNcncLXxpM7IzW9bbcIaWN3KJUeyS
lND7Rfu6xLEhGn/LJ8HPqvLk0m8P0wU5TcvN88OFFvDRQZprtt05vq1hf+Xfsde8
qQ0MjiT1j816cISK5bfAlMi+adyBNtvpEg5jr542UB0OQUEut8kEHhMH58goTS5Q
EcmhpMO18lCHUMdt+43Pte1uha1u6rqu7+hC8nqjaLBUOtQRYxIcem7w7vF3X24o
J3LWBSOTBq63TxcnpsOcdFbg/wgf5MH2F2znpJzYs0FaFFuETe59uJlRAdlc1Ldo
wHIADyt5hZ7oOZWv8x+iJl4fgulahdCTwAGS3yiaOpRnpliNNi2VVsHKwhQXZB/c
xhPU6MupVNur/V08DCUOF4U0WtesMFY3JyXIU02GpSVS05yEQeh55PjSG3kOtrTd
Uy+HEGqMs2T360dEk4LaZa4PfLdD5YTpyMDehE1zkwgFhpbkGHrzh4utZWN273PV
ACm383SDSkcnxsC/yNbIXGsjCOYSQfTnOEba+DC9TeyNQt52Axgju0QLPKdCFqPg
kxQIAgtv6FU+iVeVbgSeexqxun7z88kJt4vvYb1dHhIXBq6tOHlGHC6CPeJszI/J
LB7XB+wQciLoUsQMcDy4T6hfyBDNFCS7KDVCyowsRSo9C9I8u+SSOyPK1m5SI9ps
3Wbm6Gd0wONNIVZ9vM7eh4iAdFiEwSCuZwLWtNUGrNthdei1po0+nXgnWZhRdJt6
Cg+sNCha1SGYBfVGq8FNsFTevTh19/MA5Oi8BJ9vot4K6pNMoGgKrBOKAlLf6MEa
b2SeJHxcFGI7135VhfXzfLyvXhay27xHxNicXqAHO0qcGA0X2R6A8spPbNgEVvYM
Enrb1o3A1mXtJbeKIKetEHmo1Ex9XS0ozOS1WiinNtypTTZHb7Q9t8tyHgtWwDJE
mNHBwdZY1s7W5PjtIXXg5s9bJQAfTWaVEisiSsK1Q4gXtgcjtfPySzoU06EI5c8z
AxcbwLO+4Nwn9wDq644qMowDohTxAiTkzw9jx4md2KdoQ9m2y5AGknJ9Yya8yHCr
FFjUlWRj7kLdZeG7zlrBLgLB49U7gcXTNdA1v/Jnk52DAnAnWxL083zqxM24p4Xa
MFnXMLGDw89lwOGDAEXGpISkDbPPA1m98eLbYD51dNMdRZGV0hELqASBU2bvUVDz
zTV6+oYF9Wde8tLN+I8aUZXjA0+0IQT83y/w1BE6tv5VstoTQGqN7NSB27ftuAgD
cSzDz6LG85slhDwVOMue555cyCLqSLOgfCaQI/SyyySb2od7+sEfNlOAG1h9b8BG
CgAEVavPi0exkMqobLRN1nIznila/XUL0/eS1FTXzGpCOnNFTOh+sRdb6OWpYAKQ
P71bE0BRBO/iJZvD+VS8rY+pFF3POtSOceld8qzYRZfYmPiQGO5nCIZet9RRJi5n
Pe41tClcfmfGcUgQxBDEnyBCgGDZWmmaPy2qHj0uFlGGZ6pTNfq+iUxD8ZnF8cMG
S/bWsoup05D6GwEb6LkIqWfMIZAh9RfxcHvqgVvZ82dHRVh0UW+XnkMeeNyYdSOa
uuwI9+26+UvzVZPVs5iC3L9i47NnZX6FmY0JuIb1BrZbhbB+VbPcb1dppyJmkzza
r15wC94Be1JAO7uxBYi8krEgNNm628Aimhh5pAfCGnP+o7heDBsuM8StsE24XAc1
aY9Thfy22xCICqHUM6FqsfQvyD9J8Va6CQ1uZErooiLVcjzK/55fTrBkAuI+5u3O
EUzVi2Yt5qTA/CEEa/YkeOmuTITiuG468WUUvzHsyzcmzo/AOt+1OseXtNhnu5qj
9VPRy7oAKQNRcV8AOtl+/LP268bZyHkOaAfnBPF9ZmPUyoudAbGnou/s9xK8eGVc
bs4TmxypPGXNyiCnyAXxC0hCxfQt0Llx52bLlCTkFzoANHWyJCYgLAIgrd3K/3dQ
eJSrwxOpGxMB8Hxn3wZGyqIs4zhlNQzLmfafkkX0/HwCKjpEKc7e9OAyRExOVvDw
7gwbN+TBsX2tdrXYRgV7F0rkfSARS/JxnJ5/m8ak7EqxdYFsJq7+WP/UWn689MTv
JFGO+w4qyHIIEf027WxbWPxgWbBPhvsL5IODuYyVL2OMHqllXZaRUD827ACT8G2s
glROxAVLEdXB6jtGr2XrXzCHcCqziH61oBG3XS2ubMPg9ub4mH3pMa5HTEXNvKqo
hNMSb2W6GOh//lhZ4BXNyFKxl57sI2ju9QcXENc+QnV3rK7qheB8PKXP/J5BcnjR
XIdtH4ECm8RCSayKDY2GOzt9BL7V+mSRCTsNaXVVI9FpvWgspW7MweKxGyJfEw5s
OBVNnfj8RsXT61ESo63mRlaUOFEsaCClcYKU26vd2zjmeNmkWURRmGRzx1VQvJ/2
xACiLoIyfZIOCFvr35LZTpH4agwM+1KTPHmNWvhgU3EbRfTkmfFhHftAfK+0CE4T
RT+OIYYYmC/zqscYewFkHOe839rrTeQ6Uy6/bNDwEad97IhesbevWoVfq3aBVToB
tgGud+CzxPsoqyD32fQjqnYCExzX7K/J903KVePpSCxQf/idk1HNxY+lK+RqrjAz
rGf2tKVID/qNuzK7EtTJWwHy5TEQuG6mwTZTtkxTZNZuKBw2eFgjvuCOd3WDNEVv
07uRD2XEkfdoPSWTIGXUlJC7mbe8rXIXRDSQzhgN8uOjzlj+AlZtXLsyut7jPGzZ
pkZu45kagFErHx3Um51IvgzQ/57EtX1a8ajWwJTaXQL397/s2UcU4fGze0ANxPhM
IAe73589ocdROnTR4dMBqXisoy3wx8IdTsnFWcTZQ/ZE+JIOAItcf9szZiaadBlZ
ILNrhLDn9ADC0wwjXsnc0KGoXXFahe3sMCJ+16j1coJD8ao8zfQVj5wjO89U6ji1
Ijc5km7ae4dykCGrEzF5n89sVacGk15tVdMk4Ru+RPwAWvQB+UL/G5itQHFOEUyM
np7brPwZxD7BYdyLsQ8HSZE5jLa87fnbk0tR0d5xjSoAOmGu8Wl6cuxiGEwFG90U
j7kq2O5hfpVnC2CU1uyz0CRVtJzQcaQdCS0eZn0+Y46m/wj7USxCFC5E6z7leMUt
kqkGT9+TF2Pyi3jIGEjlWdKplfxWv/wN43W5PrfeJ+YILkj/HY7/sHVoUJt4PqN1
Y3NEW4yNwttA7XqZFBkhD8RJaSSB2nF0y2yKco7+5neJIwpwyGyU7nChWs0Nabde
THb8EtBfg3uO3/1bHsnZHRSwZxXRLSm2tKHPf4z9EYg9StxTRSQZXumDN9lV3sY3
uIYyv1qnsSOoWV+kXkrtegec45/uxtWNXnGAmqtgQgyJLwZFFNvjf2t5c19IPChj
uKctLSCpYk5RQEOhBhhQ/sM7rKybVqUt3SkdfHcYKC8Kk7gOgTC9j5L1sEK8lW6o
VqRikkYkDD238FkqF8yH22KJYy4jxfjEeafETGHwgrrQaX6UJ8iSLUkTW1m1LuM3
yL5TnR/ha4o0HMn6fFQHGJ2gOZWTQF/F3Wq2EwgqBNpmIX0vLHjtgdIXRLwcZoRK
Nez71ToUoijIz5cTDGCGsblw8GoFhhFn+rw+8fN7RnV3e5zISov8XWBnwyFaGG1D
NGIXnF2vIOCIOL/3jr/jybHwxgtP7Y5xtrM0TyVDYWN9bdJmRr2RnmShuWnjrgW+
Gf7Ze7T/j1LTpiPVjHcm9RvUdoagSnzzZJ4jyeDcwiYxJTo/7XCFjwjGjH0PjXTD
5RkIQmQPo8eXPqk30VEx3RvV54JMJlgEp9zAik0KwuZ14v26ImNFCSGTInFD3E8O
AEY1fmMVVJ+5sTutgbD+c3j9i0qLRFLXoo5iN+wgUQQ+m4DJXln+RVPzoGdWPCIe
MhRQa3Gm/II8LTs5GC2HvH5KkpjgIPAIlxSY1v82vgvv5vBJXvftSPcDiOqgJPzS
TY8UGAZ0Bz3GzJrIsJ6bd6sVPVScl+ABOSvSI+fD/LyK/TONdcl1eENq45PL7dMQ
lpOTTUNfQaDDLeIBcMpbefsF1t9a3OyENBZT/hUyTUPrO/lIfAuad38lliB/n/kB
m0jlF8Zx81iLgC5oipiczUp5KrkeD0FOZfPWsoHH8PvI48nTOCjTZQeKoBFzjCN3
jTlQ3xBQbrpYllcOhUH979Rb07Jba3nbxiQb/qVWBFxKWmr+QQgQ1cwMrbfMKpMw
tJ0u4MoNp7weJgUjiyrXDOoHDXSW8u2sg6XbbPhm1pzwUSVHM62kiu4RLyerj89n
oMPsvuRQm9KLwnmcM4ZC7ABnphGTkQXeutfuSqTmphhF0OqrQhdxFf7/N4d4flMO
Jc+3CmWuRqpB5RTefcYVUi5j8XY/P6Va5TGKEpX61d2mIVpGc01RlENZKYF1mX1a
SW8VUdi9VQXCI1W2WSDFRKvQcrrf5W9lCzx2eEureYiPvCLBEACFzbYD/xAa6sgG
b73qeGsx9x4Xwa7xq6+0Ccm1+NTpPOvD2vd2sQSWZHYa8o2Up3xRnuJ+lLUoxNx1
ZzCnZ8iQooZph64Hbz94O2cRkLWclIbN1A1V+bQOSWCqWF/cElsLYQ32UrTMUvqd
3e1P0M9BYhjGa4PiKDNILdNXLbQ7ckIv/4LXQbZrcYwfdqomc6wUbPUc3mQL7CrZ
Y2PX3tpydEUB5xnQLbe9fQ==
`protect END_PROTECTED
