`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x08cZV8EWAejfKqnSaBiEQRxws3JXxWRwkPcym9aiyCXOBMwgG6v86KWl9a2fg8f
9qnsSLcQyjNxaxGq2rCMbNJevJTIIjrSC+0/wY8+jR22DX73dut1T8Nb0kvdx1fs
eVqOiqQLJtgupJx8crex4Tx8z7zQ/UjaXnWSlPw2/ROBmbt/SLIaEs6NS8lOvc90
ZwXvb87WmvqcSSPHvooIEEDZkcjskjWFlTappRBUMQa+zprwbEY8YkoPyekc8FgB
0t7uUPaC4J1rwC9u2UioP94hkhjF8t7uEzwCp6XTMx7aVXyI6keh3M7+3rVd/OJv
P0vdJQoBcapOYUpe6ZVNX2CdXzdTCLXwnzvJaFB1n2rmosITtISnmS3oJRW2izJ4
FvUIvzxlzrw5srM7BFpJM4zW4T9kI+jhP8NCZgve0sSfvRU1ITQankpKp2s0/sGX
Ij/xybUsEalqqRuBU9OBlh6dTEqPw1bCLU+MKbaM8U6WBUSXiVDoD0/jnR/ewqJ6
xy+A9jU2yxkHyGFSUGX6eD6kHDoL/nyiojqB47oCZCkeRHpcCxYFQD0cNmkpyqms
tfg0eZxYgagvGn/MLzxRv7Y95KkBOWIie8uiaLfgkpPKkRajfl4vFLWxaL+uBVfN
iF+dVF+DRsa9F3QB/2cJH8GxO2u3NuTZi3W6geZQl9CBqWsBMdMqXRe67t9D8Yr6
cLYFfFREIY7KkWkvD789W33p4klBJd0tm7G5PQQq8H0J/cTHnUf6+AvQvWh4xRhb
EVX6kwJRj1dNf1GuB2LWGt7dhIE3Y+pcdRhzhqxncX0khGbGSozuCxMDEfDc7qp+
W60+AzMbn6wYuJmJYjTGQL5cNnsC2e+6jcqbuMhr+0M=
`protect END_PROTECTED
