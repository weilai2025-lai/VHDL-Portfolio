`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TRKAJYjFkL4Q/cm/LWm+pr7ABGu8pEwwor8KUDXJBJFdWTkI7G7yEWv6Mize4ELT
EINSC5bJTEfOI1yCF5E40B3JPy9HjoKg7WQwHW+d4VAi1bbqzGtloXqvv1xiMmNm
eTnKscYoOV029rCuwAyVSgFLRifl8AdWRi+YxbZeWRpP+N+XbUcKSb6skyb6renv
lAWJzP1RS7SJnAg+eqt4/9HCK9hXbIr6Wz9zlLTyh8Vq4Wdp215cL03tHa7JC+Hn
USTODb3os8l7QwVEzbQ+mUyD0UDnaNcsF3a7ZweMzWtQjk3Q7nfQVBEqjuto18Kb
oALjZjRnNxGSuV1iKXxYUMPSPufEcT99IT3wqIeeO/FvcRMN3tLGPNh6QIe37zWJ
dFg0Kmli1Zzkt8yLG20mT5Sa/pyEnDm52Y6FAa8a4xiTNog6IQX2SGhvnDewAvqm
477tI9PIrLXAwUDNSs8t1isrMNeFxC/jaiuk6vxAL4SZCVNt5a5m9DYcbH613eBo
/M0E9DNQWHf9mFX80xT6mKxkqMOF35OU4tJOBoFYrgIUxPCA9bsQq9ND8Bt7LJMB
QdO1lEEg4/wj/exsm1W6duRZv6oB4oh4RKMmPFaULE5vclzJEdwqAMHKR7YqI2m6
JtJtQ0KKoza7+s1KwDmWOAqH6HAgYxcadYP6JCtRTp7/PjdwC1XHZZXPQrWAzU3B
Dq6wVbDNs9/RfZlc4okNLnpJfoz5vaJG74PCJVviozJ+WlLxXkBFpMiXLAzzQ6gb
ZhBr6HKBVxHPS+jOMet7axGSjGl4qR6m25MIOj6ih+tY90efouMNuHOla4K50nhA
WrpHTiTz1+dezpgKnmQ1TFnJqvZvka4A/EjSUFzY/oXphuqVAoloLrv6U1YNWQ+E
YRoXrS7gxRN4yjRdxWcqyGkP2vRXQBkF/ij0Y/9f97gD+Yj3ui+zEKRZIlRIIEHC
a9/EuFfeem4rAuL2pDwncoaH/RKFznAZq488T8rYX3hWWX863Ek9WfPjT7Nt/eZJ
ox0JhzO0hfH3vAWySxaoTXHjciIMYVz2l2+hUR87n/vQ4t0LWWFya7r6+hcCrNIK
+sb52e56bNXnTu3+DvpbyOQNkxfNDjZNOuArGUJoX6IihrIDEULVmUxX4uCrd/qO
D4PKQwbEtwaEqjkJvfDjUA==
`protect END_PROTECTED
