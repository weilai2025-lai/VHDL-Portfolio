`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hl8mgeU45EO4CmKJIhbCNczuBkjzRuYAy7Ofp8AfQ+sZisw2ZgK8ZP4gR9Zs5vp2
D2h4Tqf9c0QojBfAXEBC3p/KzY9ZgHGJaQH41YFlJRkY/AyFxAWOr38gLxDq7tKN
0Cqq1jHlQdezoD0oHza1yuD8uJQQgIcrwZfvMQggau7456fSfzdCjoytZQ38E+1o
YohNYUdBx2ZAfhm2kzDVvZN1GTi/wPAxj3jARCADzWRU7Eg4TRJ6csIq+05mNs+b
4c7W0B/fGAojLhLJHBEIuU6iQx7SePfCKImySvUQy6rMDlLpQvXLYenB0osR7gc5
NoyQ/9+QO23Cxuskp77r7T7mQ8tDR826cX4oiRaD0u6y7XZesmSXRedTVG/YKf+a
JITXZb9oqSrk6OsSgypJ+XLGuNsMDfKvj+c+xVQEft7CdFnWflZ4R5bGA2q0u171
KIFxEFtmdBUdwPC+BFJX/OxOxT6EnReMQiZymTpBn2+EiJQT6c1KAMbh7yQFNU3N
cVmZrWxxsc8HV1qrKi8txlLWJ6McmG+T9NocDgMxLKZiYvb8Qbn6QLNuYTXhgqxR
3OBCsev3VSoifBDqJgYnpy7h+xb1UCOES7xEbHiVaUJLRE6UAx/CudF2sCB/8de+
V0NZKCQ7CELgLoOP5TSIiw6l7tf4yW+OQ+0eT8dJZfp4VL6AEL/bOCgW9C/WkaIC
5PgIRdynnA9dlOqzHsiirXIANQ95343zXv6YYyJ/lkvMM/r/lmgtcxwVJ16dSawg
saI/TSmgYx38JceXBFZ5DNkTO4CQ+Dj/gr845esXjXy36bOyw8kpT93no5f/R1+p
kRZlyQRAZiy9ZC4U4i5UYxEnt6tjtX/TUg7JHaWQPBUpIC9FT+gYLIP0FZ9Vn1VI
5IFB1phBRs745Tr7hhH2s398J4fn8IZscN+M89Eg0sP03oeCsDfi7d99OvFcDhvD
REPKvgVTNnRiqzb7QK9l/7mRaGRrQMFP2uebCBM01xWMK2/I0fXl9TOEfZG2WAP0
ycpkUcaM3WHIloQ1zqbFICTxllMaOEk5NSIWkJOmdAkzL+wLwm1Oew8D+r34NwCs
CbmJ7M/XYERGltVAZtzbSDk1+GJocGjldtuES6hAa95ZnUcunwNYdWSYnHjmThw9
/duYkuvPTi9XzrJxndY2wXuknhDXckDI40hDA/Yi0uGG0osXAW5jzmhxP0Y0t53o
hTJP2PSvsH/oVg1b4D5mbYyFxIt5lxmpFbRS1tLYBCD1XwN5MEdSEaRS7Qi4Lc2C
`protect END_PROTECTED
