`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ko4dlsL9k1BC9sTPKZksFocLD1JjuLtLoED7bxoihu5Ab8osECjlkELvQyA12rtQ
vX89VkXxjSrnreVpkegAkhgT8xM08n4QSqL0c3kaIDwp9isMd+D4YJJdJYjsMKGN
rtmMPRPL4zaF4AatiuXzkHuBtqEPI98k/3euVLPi5gsAR3zM1ZBW8jX/TzwLvGrG
d95o+11HtmqmVUFBzDdyQlbmTag4rJTKs9CzUuXQm7Y86BARfS+EVHpYF+3xxrO4
unEALXG02icMyarxh+8IVvDHqjjtYV1byaLrQZQm2r0BRugkfe3rkpdqGDKGA2+d
tAd8nUHJXOuskP1TFQAQKr+EyOIkT6Lx5m7EU6W1UnMrGRqEFgaA/LlHSUcBCUSs
dY0NXNnHPGK7JF7ZaiyWQnsdJwOFWhY3aENZAbPlRasDv6LcCLs9nX0bikuXvkH8
e1mX6gyVUkLzyOSISUFGjLzccuFSwThwl8h6ufBrD404MweHJfUOKAevPSbbHrJ8
O3aZEYUeGJm/7qeKhr/axn7QuFE7jwU4vKyCSL4ZGcDQz08HisW/AyMRjW1WoyvT
+eSQs2V0vB6eu28EfPVZTfpaQKO9Pmb4XaYFeK/V7XqiHeANoUpUl7bdhNoqQqOT
4FnJW8C2rFdtXxkaru1wEMCIpDrEyFLGw6NJ1Rj1eWl9gb5PDj1d8DBiGUhW7iK6
Z25a1MxVGe+0iGkLlT6M1fqDpNc4VBEt094cMeQCuGR57nkygRi3nClxP/2wMGI2
JqjVIj4Z/bzGuD6MT7ubWRR1dqx57ET1rFGNTYKRrKEHTnARnz0+4+sig42VfTk0
2OuV79Vi1zD7/9iBhWv0r6nQ6kjixRODQZv+my8GLdEPn+PU7t6Z+sg2zzkLviEw
big9yIxqwzYI2mVwVxd1DslNrgHb+UneiEPyaUNq07PeKrV2Xb1IaCavVZ8Fz/Hc
UQZe1nRQMAMyai2wvYybNeZXJZ3NxKkw0qp306W9O69X1RsvQDVDG4uRRgaN3opI
DyeOPi2Y0HVd4etI4DsAb5NDoBzNEPh4KbXvRaQ+jQr0V3O2FBk8dhs7S0ozDuED
V6sk/jIS67RE/zbjuWNJv6u9FoGC8iriPXb2YIu35pMC7/gtyG5TLF8zrjMM4eqx
e1/1fkogHLfNvbJe+Tp8FQxVQXsP0vE4fhgHEnas+TaQZM1BhwbbJFT5cRqPDYjz
kHmRi1LCZ7QtmmhC83tNZkC3O8TzRNHgE6wcNNpzgBn/gKesDnTZ7nY2isb6ydQ1
+HwrPIXmuM3U+o33YDpPJzYKOTE3KdLT0EA8klQz7xME63P0gotLy1gE0JEyB1Iu
JJz107FtnDuCV7ROTPI+jlPhEzyX7+7TkFAQUjicKZ+bRWK/YfVTTxeoWMXzTZGE
JCJL2cGBZEAPOUytICZMLCjFAsmX+2I8r0YsQS0GAD7gbLxyxIN0H75V1XDBFwjY
4uaJqr68L29eFIvMtu619M1aE9dGe0k1M+8KcH4R7AdmeAxuZYWC3lG3N0c0pjIo
/0sgjek+wZWARVDmhHD7iY8u7eyJr2T+8637wZzjZ4G7PKqGZr3Zi1sDXJtQ5dWi
CD6VqVNzGeUc+26fIqbyCHgFHe29PAkJwNpnCPx2Zgp0VDcuNQAeADgd48WRWBHv
p8ioI2kK0vsW67ZKF27Qxqn6C1vtcVekBotZshQYyDVq4W7h7R2POe4Pmrpux30C
M+5TpwvvzpLeUu7vu7A99l7d3FRIFZY8vAwxVuBjfOYc5ryrhPIb82MuDzXp6Ve8
k3Xnx8fOPbN+9WVnPfXiNyUcudWaM6tQIwXVm4b1LQF7EkzNuoBLQgquMWw9RWPZ
g8L2t93TeCCDYZwOO8zKmHCftRGzpqSVdevfEYGFLDsDT1XP43ODBRtFQbdsc0UM
RIvD1e84FIYKbUnRvELZ4KgO3Y8nWkSVpaz+xlv1Sz3z/ox+lCRa+8rM3GYVmO6V
/f77vnI76UoCIW0xAED7yQ0oDwLESShzqtOLXc1CzlnRsXtMnr3yx/pc7wluwsLy
S22Xarh1LJdjMDdHjuSZF7JjH9w9Q9FMj/fvc04umugLtdeDj23d+gcHxmB6lopZ
cT8tLWmgW5X685ON+pRklKzrlZDn2f0d6cZwWSFn1N4bRxaBnx3/3/b2eUQ8S2KH
3BKfHunnrwhH+S4h7eNaRkmNxriEGFzm/zZqw2RSK7Mes1fXNgMVF0RLc+Z+mgSa
XU1cWlmDY5KYAALbGJ8tdirU2pSP9LLhss4QOYz1XLbEy0OmTbGTWvxJuK6nPCfY
8qYliBJZpcZIUlhHDgHapCN0mAVYylrNQ70guPomyaDums58xj2wWqZpIuNLlWa4
qIMc4w1peArzlWqSL7RLWpg5UG08rTkhtGjxogoTiryWuWQBv0GIO5OrVVvobrPc
XzhZ8UoKOm55anUN7Jzaa+AbHDGu/TUP8f3bnYmJr9AjbJx3YiusPPtClPtC9d3r
SZUBp4x4UJnlsi48zOFwuvEK1q6tnn32BPId70M6xkx+vrH7WlyZrtz6sZsUkG0p
ovorhY6OWtIBC40GCKLjuqvbBF26NUgAUTVGnY947BXvaYGU8Oc4/pUumy7rnClW
7qRzV6L66+rsVJkJ2nw+zx1JWHuqb6TA3bwMhh9Ku7W3N5J0bS3W41i9AeHOmcKi
U3rPMqaAwkvzGDpu5ZZrd5k2L3govJkIIQH0K/egVKvYJjihqrFuwstHsHjM6UgZ
KM1WSc6Er5cs47uSqz/cHi4bV5POwl+Hk0zmm3EsZYkqr6lS0HsbKY8Xsnco7PWG
iOUD0z8IjAPKCV/lTghmI2k1DRZNl+pzVQfISqfB3g68qCiqTVuOOluXXlJRsW4y
uv8oronZvU29ddqMMCglBIHf4ubKGgLvOHCEOa8T/DkhWLDeQ22QmcZ4UYtrPzso
LRQuoRIePKYiCPNo7J9ts/f5vGAHUYUSgIuaGsKZyB9DXnErU6d7AHSYjbEB0Cll
AxX4Oz+y8VsWE/ZVvqScIctmn3kJS4O6tMFwdq2VR39rvPmiFrbp8eljGTFCIj+b
4fvhWbS3xy9Ot7p6L5BUVfa40sSSrMN4rMoqFYWWz1s8vY5Ak6lp9iC3TtbBBS/p
D4SynT/19YpYxbDiCyQDp7xDAHV1tb3+YY85X6bwQNgUikpMSBLax+xN7JvpQPaN
yNQAe03eMsX8t6qocjQllR5PRGc7KX5ZvlLyj+G9UkVCQDBFbjQRVuQLHb6Qd9XT
RUiDZ/Akh++BbiAk8B56AGZamlKSmNvRWLjjq4W5b/5ycl/dKmy9ZPUKMeHIcqU1
ueUJOocvMXTaZKUOBZsxAVdJmsC/Ur7OmNQO6NFF5WSFvKX2rnzqi2Mzlljcoucu
HkTzzHRbh4RgSpV73gh0fOburiJWIKnECK8L0Uj5P4Oc5ZSK2lfPzN1WiTSSqiUr
u1I/Za2pbBTi/hemYWE+C/UZlGVQhF8mYRNfJTgF+Ojs530i9Geq5mxzrcTx1Zg/
Yn0yXX1qurwNWfdvdQ0ZSzv9DlFPUrsRippu7pSqpjADIAtcqrxRr1/EyecbcHK+
w0NpSNaFpX+Ow3tOWF/oPV3UwVU0lBZSYGV4eFe3mksv2Tb8AxK2c0B4URIQokgd
Uv2vfFtBygHe9K0FZrcByOqiCN1UwuIXmXLxxibM1KqN/LbyCwrtRY+k9MXVoust
KA5g1kAgKxXBgk0MS/WgqA==
`protect END_PROTECTED
