`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+x/DG/e/37senMHs7kZXc8fVye68Rs0PSnmWhGhyyiKrMC75Qzm//K1F+eXEGF/V
u7MQr+Y7rQNm2ap+Z2S5FVMOURBf95RBcmNSFB0tXbSzzJIHBvdRmZWo3VwUUJBs
mG15kpJK/I/gmOwMIXcOQJ1ybdGYvoQZ2x+FqmaBpljJXwa6k3vCfTS3+rpLTCE+
z8XcVdGpNW/0HVCn6aB/FRvlx0coj3a9GsQCUWD++tPwnlKgkNc0gByDUUUEgkEx
0k/1g76VOf2VhUR6RZZTlS6kmjkL8hku7qKvV+SId5g/DZd67FdzlYVeyhajq0oo
4a+wnmFcz9SBCS5QYswwWK/Wad/31Qu/YUgieUnkK0vBY28k8etWi30Z3T34Qb/8
Qtc0IZPqGTfD7YScJBBYFhjadbgkCnrW4PUslLE03brIEwmmu2u+vp9zNfdwReHb
Cwx+cEBcYdvv83rxU0dXolQYzHHRJeawvXB7Lj4vZ5/DhhKhwDNyAZ+RdEcJm6Kg
HYQCpPL6dfh7IFcXt45ZZMbd3Xbb3B0/GRFdIivvVRlCWXWjQVfETjlldRAgbxCc
o63S9hHu9+UfgDXZdlgjbamdQig4wzhJ35h5K60eeXzNUOjYEQk3umkqAM9IPrpb
yp60N/DUbFjy6fcsOolQ6YEZLTiDmwdkY0TmyEf/EMUyU4di2kCgayy35Jp2tTgR
hbRHeqcH52pj0Wqlm6GCDXTQ0a5+4jmOBSrM48XmRh8nxkX4T8dechLlTN+/CMQ3
Ma3qk3JCuIlLZNwpUC44YGrxpgLTeZ8Oe5oN4ySMo7uqi4WdYGbH7YGDfHiKbGcs
HGkOxPWgkpqc84T4xzhHi7kgVA5+jExi//28adlN8tbPjLVHMCPdLcLpMBQbgRir
fXhYp68qpN4F0Gya/PsH/akcWIBVpZEGp9c/tbgy90oVsNcI1JZCvDzlbny5uZ51
KxU2Zpx8e0VnPZa/LFUCP1Ln/xjG1ZpuRv8R5F4yqoPioTSw5dsBSiuEdiaz8atV
QI45nRERtxSvbu75JyVIBJwT7HJKLBumJtAsh/hXNA4uOOw68nOtE1X6p1wKNbcl
UWCkHNLIrEl5jzEWQNq653vJGxcj2CQBWC0tjfyPjuT+tX9ctebtY62z5eXoQatv
l8hdsMWR5GhqalTmTxya7CWYGK/J5CBILsMRvA2zvhaaI3ikAdmBkYwO+aM2PaH7
zoerZK3FNyYkEE6Rh7wUn8Hcp4Kc8x14a6pJq3ImTDYTzMk66/kuOwO9Yf4b5aGj
oUswjejToKi0Vw46cL7JuH3+SlTJl4Y0spogzlToTsDtIX6tEXpidqLvve82Wg0X
itDQgLK9G+1gfAbrZwZGA/ZTMGzOFFNmwTzn9cIXnS2ctnRkG9p81tWcvE32qWhm
WpbxzagtZ0ULLnUWdC72Z82QN1z6X6iogixTCjKSU2r+wHZmMYf3xVmFImo0tLzo
P8ALktiS/Ooj0HwJCdQD50XTMe30TM4N0+oTVw3rK6Gn54YKd5/ajw4MAQS2KBxF
tUGohIsoH9RRkFa20pGlrReJSvIr3oNdIYTt7RraFNDSUd/VI89pkMihhKEgWhBy
4HAqmJyirrINQnoCGbevVA5tOFBTmz7jdF9dLrf1nU1Zp8nNYZGW6ZGCY2yOMYWD
64gYw7ubsnfmFOcEDfOe0mJe2wgNKsQncJW7mPEjL0w/FYpo2djuexa4MAABOFWn
6mftZLoh4E7hWQibZCqPqT2Oi14D/7KooA7hiAD1kfPWzGaiMgtjYNIlb1M9jKkE
I7rxkKpiHaPvZfyR0q9kCZxzQg5NbbB3VUVW6/NG7Zj0CvMdKnqcpqXLAjdlvh46
dtAEdgoJA1neWFdfz5/hTPKGIC6Rfs9+7P8nffQcMv5YoF+HTgl7ZBQb3Niqp5lA
uqBMWJ8I0orc9t7bBelTR/3h8uJqciFdiL5Ntt8IG3RYHiOFfsbtXlDdLr5XIDie
vH2vnBTKNOo4HZtQjqMbDouIGwZrOSCwtI8KwZpu1+EQXm39EOTGrdhme60Kx5hy
wfTRyTu07W/2fXDfyFEvz8cyiWAzB5mnykkTODtG33E/3oG6wM36afeXrRrX1R1W
/dZLUbmU4tMUIfwn55G54cArlYTMlC75ikWA1EACvVTUigCP0WMsusWelB4bY00W
fSe9QLFlZPHNbv58HN3EK3vg4pMxuxfIcRddpeWZbQpkolsikYXKDf2zRi42J4v5
sVdhE8GZ4BzKx7IoKSOsbcxN5de0o6mdQXTQxfy6APbJEn5E/RCzkqxhFD+uavC6
rA4/GGYvzF+68kclcJe4zmjt1rXSqxNMSjvzI1JYwSzjKPr5i8KlRjTliaalgHyM
kcPeFWjlqlRtxNbMKneWJRLZO3vV3GQa800rSPB9amelccjaVI69Gcfg65uTyrX/
bNRq5DAmaayr4g3Jds2jTGbUPIemOILFJUEvVCBek7dPrQqF8yT88voVE07fQ1pu
rNm4YWsv7E1mgfptZW41qTJcGNI2q9AdYs1qJCNl4XfjMJV7qoa8n54v0WRv1l0Z
aE431duYHiuoxO64o4hy9s4d8pyUosOQ9BSBEO8uBBKrNZ/GZyFDJC0U4iP4iVbF
7HP8js4ObRBmgBdBTOQ37vkCuLmN0xMUDefb6HbCwLUuHeEYLwBIWPha9eE5jdjS
bV5ooEEHZkvMadoCL25jbPReY2yUKCEFE4ZF0HPPSL2nhbk0DNZ95Iz9Zc/WkFDC
uyLqesiw3CV7wOpUCnir+Q7RC/jWmWYXeCJ31KTw5JwQMktmIZTQcPJ07EqRRenN
qldBbHyg1iQqJfpW/1np7BVMrnRHtlsq7ehUV54ODjpqtcR5QRKizs6Eo+OY4L6+
mTrroOMaT2fnPhH3E4ISeh8j2phIoSunX2hpIpeAqDCiXAg6E3hTnKDydYz45Xh2
AuCgfLHQvE6KVJUXn4kjqH0V+EXJuTBvjhghPwxwNHxmpGof4mZeuLxr6JLEQlOj
wwXlzM6QFvCvdxcbD/4QbJzEebyFPZI9YBwzjqEfDVSidCujDK7ow+OYbR2mrSIg
p0Rm0YCnUy/WjOcQeXeviOR4pFQdagX6M0A+1FbwTagdaeuVSU6UV1FHIVb8OkRA
ZaQWLx++Fe9nYLJP4AIvy8IUA+iL6KorMRF3BtwiEvokZLZd2LY6QA152F4ZNZqN
uq0TMnP/xWPKoZyazdKbbOcNBdP1m3CqQ+KBp0rVuEco6nDf92G+GCGzc9auvBdF
Xz+lxfKCtJNwNyQqAIBdQoGC6KOf/DZicpOEMlytfZ4/151SlkC+9xP1gZvr+QXX
vTvmUc5LfAWgYApI3prLf5dEFkobjrEUowiw8oTvB2+ToyT3Ikxktkefy+NcpOyf
W/ERb2ECfJRpRUNIcrfrJIJ1BMGzzCPTB0MSwSIXlX4Y5BPjhZk35XO41mflX8fh
BpHwoX/70tn0X5uvHUNNZ7QYSgwOXEFNgen9HcZ1jpZPsWkKpoi+qkrM8meV0Dhw
sqU2Q5N0phKdtWvzivZE89uRiXAXKj5CN/8WtbZ17/nJrtaD1oF0odWOgQ0yKdCU
9t8d01GtGwnISCmboatGZ0Mg2PyQunR9yfzoAM2VwqHQH7wq7hKhyeI0eWvKi8I5
pYmKbtp683zEGFEyBNBu0UIZb8xnecZx/DSvvRDBPbQe0TyQ5neC4BvLQsl5nYiO
0sLUSc0eXlnIugseHoI6+jMthbAW3tZYMJgB3BYvhKJ10c1aKRVfibmlQrJrkVXY
KH4NR47/5wW+s6yQwM/hs7Fg0n5bXcdO68ujUGtTkq0wXmHfspUL7MOc8RjpaLTw
ZXKsZff1BgZg6pQM7YJuHH8TSAa/zlr1AvKAV84lbB2h2ZqtW2Tdtsl0rypj/eDO
NfSdnHfZ03Vuy4Q7btpD834cszO9fp56B1F6O2yiiUJrlVc7R7tBUyTJXT6DSG/9
6GyEpl6sEkFa31hr/dbP/I1yIk5puWQAiZ1uH7L/5wdsefLfh8DjYc4UyZBTDqey
sPQA7lKDkNJwHe3BiUxCqN7sK/vif2BexuUvex+TQFalQcgZ05jbRU+PNZFApZtw
eLswZdBo3WagnbKXQ3H/n7zbbtukidFBX1O8xaUjmbgKfxKlr2VuOYTppvH9TH95
Om8qflW5cfe7TW7o9+dHihnGzXFQtGJhBbPcRfJZmAFz3Qg1p5DHHBmArpiOVhIT
V88PszV/maoWYLvfRVXtqkQS5oKFl8tJbFd4AHlzlkkek6Va37ZVAuxQx7ZhGxPi
xAsaIpEaGhEkikxXgKiQPC8Urlmm7GBpN7CVr8yKoGZB0XJIeUUrnfm1TkN1vdu+
8A3+GwA+hQzrfyZcJC85YCYj4OYRVKfHDSHdv+gTDZcqy4oDXxBpR34VuURPtavX
PZ/PWChXzMSO6wpKv2KmFh5V/44wYtf60kzcmWeV6VzLdlrQu3ZA3Z/qvUdy8wYo
LlKwO7dxQTggP6tbj+rP44GtAiBUnu8KlLMPK/vqB17YDyHloZhnuZyt43F8FETm
cDR0k6GenlXw16sqkXF0Nolg03PGJ3j1Ae1jJj9Q90+6Q9UvDzSNPUn/Vclgv9U9
tN+wIeHTBo/HmHhx3XpJZiZd+TbH71zzSypgP4GFNJVnqMKzDKvlpdXtobf5gl8b
T0ECQjXf5SkPgWCEhrLfd7dxkMcCZxmNv3J7tuwrRTgtYJ8CYMS/lH5Eb1Dnd3zz
39FH2aFMHlugMs2+TSv87frQWhuJM0rBUUCzlWZCF/NAMSiQb3glKXCHLtGctOuv
RUJtsnMGlkuzDNQlOBMja5T32eKEC6UhHM7RO4DxHrmJpfgxtdUB8tDwdcdYcuev
3vaKHUWGfYIiDHUcEs+56fkFWdIOMvy/4bT7/yYo5aQY9BPVXawtAlcpbg00AKLv
7KjsdN0GAhSn09Z8Vm81eNQG+xL9cJ3cNWcAUgA1cvONDTQtvBAfWt8DenEw9pQQ
bOJkrFoLU+o2coEuc+t6ZGd/yHIN0gv9NtWLbJwZEFb2qz3Pz5Pahpl4OBxHKEfH
9otydCvtwFp4p5isAYHTkzMdGxDZNpboeJSm5IlTsge7OHaVvs2+mLiWAFB57KeL
Df7vdxpOR9qDnmrcGWqzvv39Q++WFhr2iv0bpWeSg90aWkxj2BbFAkxFfWo+0JMv
aWmOox3Xd0M5mCQuiOeW2EVZ74cye1oXDuPozQ08hylsQLymDw2KHNBhCtt+wop5
MM94gy31H+m3B0uHFkAuaSO+97k0MJqjSXNd7m0ysKAq3H+5VDvcPLFFQq+6WpXH
kGcNFlpXrwgNG8vVuTYQVxGtztbRTIpy+DFHhSB7pijDFx2TiqohUcDjlvDuISSF
SGNvYblIkH2r/OJ9O9w6jlvL4YcJdUQ+OA6bMB9G5PZmtN9fiKpNvP4Tm1CHJYyF
u+EpfxQT7hw6zWFFDhi2YfXUudCyedsalWQpAsJTrhNHoHqU4mvJ+me9Y6EhBKYk
g30S2dvCa66juaEG3OUbUB2erlmfX+id1K+OejSmhtFIWOfKYwXRAtTue1fHNSso
4T7Nsge6pOezXIuDYKBnhb+OwiTAcSRv4VdcN7UdpvNuXq4PdgsZUw3l2gbK/szI
iesFKXMa6vIHR1fQt/Ibv+6EAQUlqfBaOvzBc8cP3lmZiOJSruXxt9VXylLCKNPq
70/DQ7EPysyWMVkRfJ5s5X9C3JWw2WzT/4YVocPqOQ/xTgLtF3IVTUaXux1orLJ8
/vnYFjMdvq7/JltHQiMk/9Z0rjb3y7NH5k1jfG4uvKwH0W/XN6fzX8CpTS5uQvDx
tkwc2+5hhdITZaca24mUaDWro0i9x8pGD4JiDVQ7b7P4aMpy0TXr3amo9LccApw9
8Lo2FfRdVbkY4Lww4ZedxYaOtqqY7x+x2D1gb2hTi0NNA2tfSHOVSe0nn/hKNk5W
yHIw74c9NtQorcIlMwA595Lr2g/3VYeKXR5vmUHf2zQVQRiJrw0GBB9487mWr/YT
tqLAU48IdqB6V6Zhh/FSzN/Z7AaSbr9yr/TEnO+8vpY640aqjzQRlurKpLPOeg2c
046A7FMdy7SwAmpeHGcOFz46UVFfcRyVxrrGvuBzxa+xRsiqsuW8snDMlOvUlxfC
HPMlz8O+GhKBGeDuXnTx2g3HVeJcfUsDbdIXsSXefhYGrjBW5EiOFCCvGbOAEUBT
TLlvjagj9fK0gfu9H0PhSZcaZcs3VlHG7b+D6V+SjgxsPcURaE8rzk3s6KJYLXc/
rDF0lj3kBMt1xhN9fs+iP4D8m7OpHK+uHN8T1DDdhXRG7qaNNsAXtsaiNswx+OYX
qZHkl1n9w3shPKCjxYoEodaXa4Owp4NV3yFNxeS0org1/MOZUDknkD1HgH4OeCLg
JuyWqYwejDAV/ZuGms1iTTeGERVpBf6gKvLPZELg4cezxQG7gLH9p5cFfF7Uj6NU
sWxPdCz9kPvW0y86RbeNR60KkrRX/YpUgxJZR8ncNolDPYJL8xVfnq/4ZWUQMRZD
pNoiFPhSiz6T18OJwWkdYroV7PVFPs/dst2AMllgPFr5jF3KBX4vAdu2P3qC+e6m
SI5lI+daWk8QsmVTXtfUBYUabZp8QBld6+xyy8miWVygEyXn9UviarkSnReT1MX+
OvAmJC61ihzLRmSKOIx7l7ho3dEj3SDhGI/Uk8I8IiJZjTpDOfe/jwRMYak1Kvl9
JV8kerMUvJhhYxP/n+habXRbMUGn/BS6OAIIPPovcWcPvojqGDrkyrX9c/2Zte6t
tA7xmEsbmVTSOYuPZZEqGBkU3WDv0eebLs8TdT5DRpgb3krzwCn9mEkd9+QWE/l8
pPBrO9ueCIRo2GQq9Dq98mpWYD2h0TcPQH1EnsoN4WewECrhvhKgEl6c6HriEZ+e
0LE5txXDSB5PQE/HlqBFYPq947WhMtxR/OXTQUYN8TRW15KR3qqIJ+GeSWuLo25m
HQdCSPjiRYN4YWOnHTR6MVjm2acHmf04SzlMz1yyzcLqLBdhP3pjhWYGS5/YSITU
4aD+PilqNzxZ8uOLdg9y7iZS+grw3GYGq1NAd2H+NyKqlcSe5X33VF08AL57fYYI
wBhYLCIqKyzQZ3V1YwrqQAG5JQcC1yP00VeVUNUM6fRvqPzcTvWD91MEbTMfTjkH
ArZkp8xkm1fCKjc2KfVSbmzpgDpnbT/f+i0qML79QO5t3t+gr2M9mXoH4XQG8ht+
Tid0845iS5YDXWGQhxy2EB1Gg0L8lrAyxs4fwer+lmfszfyKgiu/WQ7XwNkppkhR
+EASMoWSyIrBrKzzzUPh1zll9B8W1YYl1ljNC1ckrwpttXk7Lv7BiTcJwU1BvW4b
+1DxZ3f3SJz0Hy+AXKjnGxilOD2nW+E1z46qoBX1QrsDKHqpm32sgUERXNGAy7RT
p5jjewhQllp1kvDhVhZdeOsFH4Ib4MzkRHekBRABnorIR8+yZxVrGO0ikf9VbDOt
zEQf+50rDGT7f9PGytRGCYGNKIzvjEoEdn/S23jdR0OD0Dbr+nOz4LxB2D6bIOyG
IDU8eUsIOEBQ1E+sZPDq6FQ8F9sw27YJiM+WblztNI1YRkoNtZPSqWh/4XBQmiDf
uEo27qoX/sQU0f4LJgCLigjbzlKkitcDq1o9BzKwr7gqb9vGgoEjyK5qEIY56qp0
4+cNnHVVkeNUKr4Zw3iX4+s+tFr9dGRQCLMHpd8TIxHNBhDcVRnmPw6E1MSHzJTS
04URA/6MTWdrXj6BKulP1eSZLpOQFCcQj3HotzoSGTgEJkVtFWziw7o0BOBHZs1o
JeXuZUs7vrfBnNvQvw1avw5mZfqcjdVMsjorddOKL/5fbx7aZkVR94CZESkUFL7W
irOAInoXFleNkwvxbAvJtuQ+BOsu3R3ChO8W8VOR9HHOJJsO61bIfpBp7KuHP7tT
nEMOr3zEMRIsTqLS+qQdY/hSufDDugvlpI/1ZcZBzVAO5MGRY9/LIgFHUd96Bjas
9tRI6Loa9rVt2m0KZzxqM+whsygeIqFxyqW40Zq2DlnXQ5Rx19n7CreSV8cMGq5y
DKg3Pzw1/INiqi3ItrXgvz/6xoWOG3dtg2XUTjs+H2LY/dbLyaYZ2cz2JEAIUfQa
nmuWg8dLTo915YsdyhWDfPz26WQkJ+yMcRiimv9V262ayf2CrPKmB4OhLGsJJfwT
rmaWVoZAWi5bnVmpMDLqN70kdHzu3w9mvJC1oRYnasX+3af7ulfZpIO/ugmZaskD
1E5GHT1AM1fyZb+nA2EsA+Wc3jKxmDPLOkZL8FfxzIdHegiSaPZx3Qg6MOxZrqj1
XlMHVWrmoi6trUQmmtm3J2BTHPhgrtK748kOa3R3ca0XNIbe3s9uUcU96aS8Xhj1
ot7x2qIQX0gzRG4K+NZjSTSaIhvNXVaWIGLxl4JxWPHB4Ji5aP8cqN14Gs7Hl8f/
pz/cjX+1GYzUDE8NKwy+3ZRSgzHtjmXx942Y12yUprjiOjl5sRD35UqAh+MJABTr
NvdgzKQe5SkTyWIYuMGeRxmL6UOBQzHh6x8J7BepQqi/d42YXjtt5ZELLfgDxiFu
9qOqr5y5n9F2tiKdwJriP0oGBARDv61ZJDFnX8Z1nNJnHdmbYKblOWYRe3eh5Mby
b/DFlL5RndEqR5cYaOs5s74hkpIrRqN1YZvcGDJeLzHgK36Qdz9Wcx8qtd/RTQoF
W6zGLIjIKRAe3ASpNjh8crrK301U/iMCQ5qMCmtKvDsyMwQxFXzlgdda+usYf1Tc
Wcz1Egqclpvmm6Y2CLjG0wWWgP/1mNbHIeleusT0a8Bnp7RA5Ibd0ZNDSO9ZpLZm
v51Io7aHh0WkaghU9BB0cEuki7ngb+Hg9QmImpVvaZRiN69nY2ycV6fEWlhsFwYC
84cB2XOluAO0DZsPc4JmwMlrnjG4uwq1zHjpav7/nQwAsn1XXDnOF1HHmL7TfkcU
QrSdCZTm4xPOMntLh3E4Hii92IZAeKhe2XrJCmfu7TnDwr2IuxRNu+/UgpJnyOhE
WPUCmdNRYS8ZM+QMpp5fKf8ceG8wwRq/SlpiwlpgBzQ6v6YdFO/VeGXPjMuzX8Bv
tqFYNGtPTpFzE6JgNFvmDJoBUS2LBdxm66O+AD0In/BmWU/6sA120Jhmp2ylYKME
wFjyHmaZzXq4tyb35gU8uA1WtKN2VWlMW+hCBr1my1vCl/3jYf1RFgoJJxGLvtme
IyUHXRt55N58PNUiiO1TZsYciZpFRh8DsQd4TqArEWtPvh+duxGPh14PVhi+cJYX
QexDHvDHV/uThkQ8yNZ/Gh6Amo22ymTT3MY38m8Zf4OeUN9ysjZrLjrNMciKhN89
nY5vCjvpVsmeXAKYhjJGXmLOBbQ/1g+FK4GCV7JLYt6eUfbpmCqZY8urjtzC+yPo
/6mvidSDOEITqWPkBuOqnCc/1I/TrEE+lvRLRB9EyZWixsZEGjAQx9/MwMIuDVNB
vfIhH7lpNJmgLHKGmBskevNlYyp1QsM7dx0b6bDRsKe09dQHfSdBMhZehbSt7135
YlkB5retxVmuB5JQlxPtg5YKuqf/J8gEzDe/X49+WNVoGPiBj6Bj/JymJSC+FJQD
uL+59pDVCokfvvMOs6mQ9hyczVDQEAam2kQ1sT7qNagVu0m8yWTU1cplYIiRcK14
J2xIerITTYN7P4Gl6WJcLaCVuIXJjZKRhrEsVoZyXsZzzFwZZtRwG3X/M+qxMJSw
3Vc8V9MevqX9dF2AWcxfvqDLfcILkm7WkyBZbKGEfpR3v9K3RCeEl/5dPrfIpGKu
wqRroN2Fpise80VkdzkPsWV27ZkOzFO/Dp+GHKDz51Z5ma/Ky9TQfKuozRKAZeLt
nv1Cy7LWZFcHooI8tmOUVWtywi9/O9VKAGQNvlh5kxWRCnqv8j5rcEJxldnkc7Fg
T2/AFbExfdwXa2SSZdNZ8eUMeWjA1jUffcUVbk6YBE9/VrWZvpGQ+Ay2L+jcF7fR
9WwIlKjiS4Fu7IPUhU+y8GpJu1rXrjMuQ333Kh9YNLtbPc+s4PgZPHLm9PWH8uOd
57BYKoUXBrcXMi4t/maKcvSJ8DfKIz7L0XzD1hmzZuBcV8J50uyLj4ppp8l7WgFn
BIjlwo54kIaad4kmRW4bzqWu+0skc7XCzDw5oLehIxTnmKq7do+4/g/0RuoOlFKM
QfSmLASOW4JnI7rrYQZwrtILZy8yF1L6rE04zNi1Nji3jMQqgOTp4If8bWBzsBmx
c/oiJFjRSpixOUd+G1ulC/JsSp0HCXHvAlcKeKf85CCAm1cAbbcP+3EFm9cwuFmm
/wNdpk62tRE0gnXFmlF46vXxDQUSGwlwyQYMBq/lEPPoe2PyJKEUrnwDwEKtYbRP
3s2sb2UFKoCVxWp8hOlwA73+iGGuh40hHduy07ZGArDVW3F1SFc3be/4P5sdW0IK
iihB1KbV9Y2b6cPWuytzrchIbJbKtF6XqUsxDMi1AfLukZl6Edvk7SjAYHwc7VEy
lRfYqa8n1Dgk7pZipWsbBfcjNDnVlakjU/INBVtRGv3JMgcixyrdUVHhixUYer/K
UPAlPiCGIiytshzmXYN9NmrfUA8S2TTG3252ZCOOy/Pyvsl69MuBXttY+EgeYaXF
vQtOJEmAWRSQHZ+tfQ9mzeYI7PLmJcYpX8qyfevD/+wk1yHTyFfdmlNaguACg9pf
ZpIBgyAsxesZmJ7tiMxJ3cdA0jEyP3ZpSNWgpIeYlIEH9dhlckBl5l4UE3y0SkO5
ZYVLd63KIMpLqw26oBZ5ifqJ/iwm9i+qwnf9IZA3fwwCkpY4M3/NZu8pwyuJlr6s
n/VsGIdt6mXOnvA/OVO72UkC0tZx8knfjjwjtg2FWaozaBz7msU/cZtHYEoZ2ldV
RABrDCZP8X6hHpc7+WxkgdY8phyZQH6/6EHAtQqtpiBuXBb9WrR+83cgTOFjZl8s
hLnEUw5xWl3aRjj8SqPhgqLKaTZ493+jKYVvTMOSwG4AsWlaTY5njIcpQjDADy7f
CUxkJQg91yXFri8lO/LhoEJAFJC9LawVSXpgj/qmJao0RXj8+ZIvmxc5d92rTdDD
c+h6G7E1CBfJGrzuuq8ehsYbwm8v3eReP2d6ljbtMOU6nzNW00cx8yJqib5rw126
Kw2bAs4Wr91RV0O0kdEDl4Qx9R5NOuqeeb44BOcRJgrrmGGi+a946GIitbiJsHey
bVD7vP2TWrQ1qSSwZsLvk4+t+MLHnPWWasyEPZHJfrZlmG8NO28hBam7Vc48W9Cw
Qeq5QiJvxP1dGCtiFc3XqHOndYydWCsvZa1ub2sZGF4wdqMZpjV37A1OLjDEz+zX
aLF5L1yFgfz/B5w+AWE9tOp4pgIHI4rIpb0L+2h9wZIHYrIo9AWXwmi0jF1mGAMy
jv7CrbIyQ/dSrp/4Ng2YRCIq5XOF5dAufNyCFxaT2b4ZWKx1AJo8/c7/etEMblpu
Fp8yUkehZB6vIXyflyKhEeH9lfOu0Jf2xWDGkgE6M7UXxDugcfCnfPESAJtcDBT8
0asKfZ2cGDhvb5FlhUw0Rv/kPgiGJXl3ntDbNC3ueEA8M55qJTSP4AifU+ZTEI1I
WmxpKJNn0ooexKBTVpQJY7ml/LCamKTRspSyHVV2VqWHWBF+6hqmBR9oHSEazzPG
JIWAFh05p+wlVWe6yZR16L+8hRj803jpaH7hvEDcnpaYnxTmHapxJlP1MVPHPxwV
pFAkIA+ojwgmvCqL4aBW41BFFScXen/k79JWBhIFG6hBjEPQHyeMVTvSBN38Wpjb
ojawPWP36Odkd9drPWZ9G6pCZBvn+felMNpWVLOM+VxfxOyH/ob+JjKVMsoxzxfv
1P5qcOZyNmfY3lwuaHr4aa/W97GBik8P7uPlpeufD0XGikGdj9veow6sbzaClVup
a/h9p8wCk0iwr2PLedvbuyzhqzI4Zoov5VG8l2/KehKV4+smnPuT2oKRWTi5l8iM
/uAVN4f2Q7uVqK/+2YMFuOggV4q9jUhyaUjaG5qilFKNc9AzUq3WhdmOZ+5YTUjz
r+HqRIx6XkEJbGUe/wLfZj2/0uoTBSi8kBspm/adpgfmg7XXBITCXv0wsfc7uayR
9zJe5wPXEZriAFgh+drIVolhADfvEvOMGfwVHaGK7M/2PlhSPTolwtAtXh2Uj5r/
OiFGthjRF+W0sOKzPid0mmS1q21mK1sf9JWCGpvHu2/2LlEuWXYCSgbpPeELxcc2
R9rGD20XhSDV0224WodkZjilHMdAvZ0ZmCFC5GCjKMZ2aBk83Yf4foOhA7AewPcU
CNKUKyx7zI0VdditZSZ+JgyHYVegJu3dD2rEgp3RfBa3n9rJ5E2T28qJF1O/wycX
kmkZ77WWoxMSYv8sP4sn5S7M4ukdAcfumEpKm8HJ72oN5KMFGP1uOQk21Q9ikHKU
R8zed+Q0IUQXt1ptuYM1UdIiRRZmx0LMn3VW29Y/Citza5GZhuaDvGLX3uNsC0DN
R2JP2zzi/N6m36iUu9rdFs0GKNBbm6jYShDJKbN4JGdFgf8r9PbLDkR1oR7wfz33
iZ/M5vJGZoN3dho7g4bKH7jlWMXlXJOdSq+GALMfcvQuLZ5aJ/jNiEUH0pyrBPyN
2xilKl/FydR01X2Fk4vsiXQVptRBJ0dqJ8G1zBLfivMacMfuzyhZ9Y7wMEX6t1FP
cjpavo/DPW0nA/8k74ZA5v9PH8bDqfYk5VpX8Ns8ybVlXUtWF9Ptjz3hFx9A1GAY
Vwc0wPHORmxns6iFwpvDjeFd/aCv2yOVfbyRpzqDn+Cb4TEUkyGVxqIfriKNcUQF
i5UXyGDe2aECAiuesX1PIlDWebUTg4tTc/Le6NsoT+bjh/aA6zfbxx1cHXX8YYH0
eDAMfdKZ/YgIVJutvM1B5/IZ+r7oxs+5zJelf2EO8NyDi1o9NM55mR6AwYD7DOx/
jVaE2PkEIDwjqALFoLjglC0Uw+Qm4VN+sG8NX5wzdNOMVDOmalXwvn4ozD0MWxay
JtSOSBIEEIsv0WBt+vc1UUjS8WnENellY19Y96DgMfyj+g8dMifDUKr7qtFeKCKo
tm/Ct+8E+fVf/2BFEKnMG06SxRzRz1Hv1d7EmXPBuRPsyRlq6T4NZfX+THWlBLdE
mrPO3rBmvXPblY2jkbyQrenU8wW5ncnxuE6thhiNEqwVAHZy7mTxm3YQrG6QIXIm
kr6mXqHCJLt4ZgdICQXfTVb2HIoAmbmEsO7GNiWlG7us7zXhkWVSb9ij85P6sw1r
64xIOpsmK9naiiYfRP3Ht6hr9UoJqU8W9fSAMHctzizFuUX82gDeVrDqYwH/hUu+
7bm1+lGxfUR0DUqVgDeL0w==
`protect END_PROTECTED
