`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYdcV/4JEOPvzQmd7AX7lT4HAq8L2YPfAhI3zYLuqPcPFkFktBcB3Vgrqa46hzpG
3OsSnbzdpXpg8b1DZTZ9GtTCOiXNDdqBcJ1NirgXnDZVrU6EWMngi+mDRVq1+WMv
YIfSgjlcxSaa8CeTBVgLsY6Lt4cDa+8bwFkRdYqyMk1DCFY0+KWdKlRFpBhJXKHw
vxN3/HD4V98MwATPzF3f6QQRbUjvNQrDpDK9+n2bzEc9EjNGtnzFCz7D5EoCFvOJ
54JICrStQ20PqV5+58nIhvOCqnjyFY/b5Hn/F7JZDyMsp05RRQ5NaDaX9HU2Aj6S
YNgNZXxNpq2VdfqAKKqYcQIP/o4ZZ3Et0P/9HZC0KD41pSSXpp0NDmDDZ1J6c58n
0EaHnPtghXlYIgY//qRkp2hmA6U1Av3A/wcmk/mUNP1FrFpdiO+gJRMDPRv1VxeX
GHS+i3Ac52Nr1dZxV3klYGNGjA0jXPrmAfQDrmkE0ikq0xLNx2abCqwnBZ04JJyi
M3uqBA6M2ZOD8a4TzElzXxcC1ff9AACsRbmhuR+BSTjmhLvPA4Iht0+EaoPdFap3
itV923Xpgt/LZh6ipm5xWkisiqJpvalyVOyx1iE1usmlo47wTOq6qERt9oz5/mYH
nAonhj6nhkfQDEamYw3+Vfv4q98P6GPMstlJdX5XkZH8Ri0SwUaYC9j0cnG+JCj/
zFEDYmq8NSgYSYN0CBcype8d2Su4Iha6/pCGoTiTw30=
`protect END_PROTECTED
