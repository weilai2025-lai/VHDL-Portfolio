`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G70pXMRrsE3jm1rgn6lhEmRqqHMeK3QFRF8hAyQYyR+vg4JSc8sOsYpa2e66RysJ
fHgihKP7Hbfn+zwKRwOha3lT+/mEwdyEtDVYA/h3577IpSc3VTkiA60F+zLXVxCQ
1JmWWFLAkS46EB5p20XQjV32XABgqyFHUO3W4v+XnXwjDmJSOC1FLrp9CmZOiHHH
gr6O+w+hpb/ckbnkMj7yv7n+Ii+L7RZbEBVxn3oDC5Gtm8i7YFzpiqRwy9BmTvKk
dKRyAUNhcSyp0ar+t10LynJMhXlGXFHMqoA+BvTAME3lnb3tlKFyDTfET368rszq
xa9epf6K0EVIlt+bA8qRy0PoDXDNX2qFWwFg4Tf4sJ+9mCW2+/4xjUk7hXHFKj4p
X0aKpi30va6CeaKX4SImd+8uOOjsko+UJJ9nJsV0Raezfon9s0fBF8GcaYxYFwj3
wBisrVAGMT9D9J1TL7lddsehKpDpAH/kWs2Y+u5hVd6EEo9mjLRCtfqIXSknnE+r
YYap5iMlDJuewpNbuPOEVtXYJYus7uQ9DFO1jHLd6b0=
`protect END_PROTECTED
