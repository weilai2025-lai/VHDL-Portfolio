`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qCqtfnqqe6lpMwZx75BbofareueDK48J81qWBOg5/Fpd3dVZEM1SCAh6pP+QXPr
l9CCms0Pxn4KfHYx2U0yXg4Rzu9Q558c3bpbmjIX6TZkTp/4J8PwTBF1DGQXCY2p
oC3HxB8l+O/4PK2qazTL5I8Li1XyvtKFs7fZcAH0s42gFO8Ll5htC4Fn6WaYxnxd
d9HDXM7GFqu/B3H8h0+m/EsQxtnhhHRJo2oaQyNt4Zm0bqy22df0GfL8tgsMFO5M
f2hRdQYpvcyP+VolNO7kSHYlQLB0jHpl+VXzvvfaZ+zuGvs8sm6zkUsd3h6Al7Jj
NaVpK18ENh8IOtJf7RSdjgUL9QjMN+LJr7FnH7/vwRUcYExdDQ/aKR2dm0l5F0b2
lJF3QGCvDRp9APglmfhfUQhBoEyttoTyC+CctVMcJRGAmrjznYsjnxUYhtkWzcdd
fJPYRUuXYHU08ZyiKnHstb6GJ1m5N5n+SPOdijnI5eOF4U9lH0ybrFr6Jb2ta+Gj
1+DWdFd9JdTYwXVSqLAqWJdlJ5gp9tOIgoaIlSxWkeDpBgcUj5UZYkwwdWCiTTpo
WtWzZZd4sJKs1DqwRCGz2he9igpIoknsNQEQlzGDqqufy8liF74n0HYPU77VjooT
`protect END_PROTECTED
