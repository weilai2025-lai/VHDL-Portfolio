`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMqXQojAtQjano+KHSoccVHo+LawKUIiUcFV3wiUEDnUEOEsdLVaSj5j6ZY/hzJm
1eZbVynIIuAPyflJqgWN9eY+0wrOyV0svmvVa7xTdSBeRvfYRrFcoKDmkeM87pms
pKGSM6dO3wogRvK3vP8bFFZ5smkQutbCetZ38BQiumRlqs4zSrXKA/prnzUBIe6U
3CP8yWVDWbEsvP3tektypBkFB8tO2G+u8eJRUFx4WHlyw7g1a7BqxQTuDK9pFOgR
SiTzlnaf5EhgWEXw6Oh18eg8P+ayH2hSSbJnHU9Um5RSkWxp7ckdku2o3/Wtrm7C
NSRBrtLPLTMgTlgK4zmtDQ==
`protect END_PROTECTED
