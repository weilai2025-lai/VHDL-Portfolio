`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVV1U8RUCta6xxPK/cKaFFLUNUatEYCunSr1QXUr+YXlNO04uyd9swjC7Mn0Ui/3
3yFNzNaTRfJuyCJSSCIcMU2VqSBBE0a+FXqSZbXkkzsHVr0SlDMP6o5SkVHkaaQ9
eW+8lJuq1Y5AYkd7N03zy5VvurH129p+yQReKFGbUyGhHhcIp+ixJg03DBSeeqXg
92u9JAgSbzJK4Wbde8+gA6cIdc8j9QhJ6fd+/XLE1HYIABxx/Z9cGzmlVECg4roN
vQ6k3DwjVR40dClTe4jjq4xJSVKe66amGcRI72jiIWXfsZJbzaUliTCfjEFRPbdq
/Y+21kC7v1rE0MSZrtT9XbggjJsOSJweQmw18/2hegbHZtpZRFKYIxoPQEg9U1D6
uDB+biQEAYjMfWPcsgpXtV+2z/rt6putM3+vmTY7DNHspd3SSQkOPSEXMjIAVIh2
VdCROm6Nwtv9hNf02YpFY+pJiDcjCtwpbTQ5tTbN+ooO/6NoNg4NTLmz8rcGo0yV
WDiyzHKoOns75yrvcXgPeL2/9s5I5HouCL0UMV782KD6NLz/4uYhkokg9Jb7MY7T
SNoeDWydH/g799gk3RyonA==
`protect END_PROTECTED
