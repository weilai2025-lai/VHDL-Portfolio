`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqwDyQg2n32PC4aeA66ZUb0BOo6hKzZ0jrij/sjW9PyqL0f0ThbkUyy7a7IOSKzH
gr3LG+KKetHccPjAnl8ATmMgGCfrxm1dnRw1EdEtzdSzFHztJ3K1QJIOKz2jiXIE
CwouGxhu14q/48eynJ49WrQfHokGmaYdmEc+tuDlCVjV8Zx1ryTHKMIsKwi9ABDi
Q0R0Ja4m4YLaibCgeqW6xFE0i/K2jwJWZcGCYyg0gEpOuzPYbNA54UpxGbipsvAd
FvN3Yw92YlCAUHGrmPTabXE2KdvO8vD2s5M3fyG8+ZgOzYl0hqeCw/pIbo+zRBtl
k8LzUGvTeN6zoMozw+3w8gDloBUtn0Zlh3RpUp798DASnTRM/ZK7BnFX07/LPgZR
zOFJ96pyhYAFRRhoKUujCxECaEaQQwWS1W1lfkNexMEZOt7cUeUPxiCJEOLeSMlU
dMYVDzcds7cjlk58575WD0DEM7D3f01aUIGzCT/trZ5R+TbgYrF9ZFiN+6oe1Tma
q+Hc+vw9CpBcb/l+51ZiIQG4948kZ9ff86Gj79Y3G1KD9qD7qsYy++0dGWSQxho8
6vuPncHk8QmIMoAvTuZkR61B1vYqvB/ho5+nXX1TvTceIuT89Nw2pdZUY24AgbFZ
H4q71b1upG8ys+ltKBLOQq1jVKJ34XmxlDg4wyvYvgBDOZ6q3wa+NmHTzHJVg+2L
zwO3Yk2twOk+OAYzyqfOBvrNarINu6KqKG7veyex/xYpIKcG8l5yuz5N0XRLOJ0a
ilxzbib57wIy79vXD0vxG+UzvEeMiq9o5vx4nTVy3XBIzkPnnwyBDdKbP5SNPstR
nzPNuKx8gQqnb7EG5H3iogwk3dAwmj4sztkA3oyEnANNyU2Sty+iVGZnye2TBRJ1
EmceVbKAswQ+/56BKTsniCBbHkF6gIvi4csNY60eQbk72GOJ630o1QIyq8xaf5pg
VsDO6PbgAhv/yFYFRUPZzxnvK8JdXw1yGvAcM8jSLNnBdc+wmTH31l0T0FWkr3hh
h1rkOW8KjaAK9/+rmYeDqEda6ib281axuLd/CIOCWccCzKTcqNQ0EMGnU7WpWJBx
pOWPuTDfzvqgMbLzg19fxLyhQrhqCCoe54uCcbSToRS4TM47C0MEtjluPOn7DdBO
z0WIHZPeOd5AdWBWVTfvaz5lfyOG9pX5HZjZDfInTwuzdcpMbhzmK45hHY8yuzYQ
U7FPyNUk28ouhyIWofbJftzl0bbsaMgnVqw3ZtEnP90HcjJzOSgyomVEkm4+BLUq
yVfRNvjC/rGZOjUUWSryUqnj/rRNzuy53t1UHvZ49tCLPJ92VSvprxRKL1XWQZI5
gk1qSFjT22Hpa91vttXKw9FvZkJDcjGU/6Yfr+VODPwUuUcC84ysnCInJcuBt/iC
BiDcjJZTADRbHsKpozo91gEHIZr9cyZn3dXNh5LKzMIBt4IRGZRS9nkle5MngijE
8RGu2PzN5TSFMuhw/CGTZWuaCsJJEfFHTfVMxqHP0KqlD5P3A6TPye3Vw20zuzmE
7O+2fSqzcogsag5EoAHdNwJuJnezutXJnSopv2+pwv0LqRRxI0qTslNgtVsp4E3R
XxhruEPu99eKkNm2hjyWx2Z6haQvL1EOQk+NxWCLLkKE+ehvr/LOFAEHuigGWEvb
r5LUJhp/WkqRTrUZPkSC8VmYtDk5GcgLeYJ9IJ09Kf0/QIntWzo9kgCKuTk2l6JT
8K8zPQeuz0R9bbUCm/vDaS5P4TWxP3ktiYdEar9HiYcYmAnp2HOWFAqdbFkrr8pv
OQKhK2vJEtHmwnSwQsVmvFcGbTL3JMH1K+iOhdCmRpdX3fLTBmXnenPUr6PdbBI0
YfPtR8r5AS5VrLUVKBo/nwfTDQerTTG8BxSTGieaQ4Qfsl6LrnudPg9fYP6kq4OY
I7G+KOALYs63plBw/JbnPeUZqG+bJaTBbQjhnYcIZjWyTiDPPKXo7w3kwxMYxg+e
8Qy+91pHAebbI7hecHKtJ2oysUlJ1Pk5lafzKX703vJHoLpBty/2SGmEXLlgS0n3
y1WeSoa3TGv2/5uIRZ9SA+r6i0xdpi5dM5mQzczJlCYjYfO9AFppZJ4nOVHk2oJE
y3U5V+ICuNns0+AKiZ4i/DhMNKqAquiWWlf7pu9LS1xypXM08M+J7QApzNy7I2ZY
CNtYC89+GvAX1vaEil2opL+b1ZNJxWzNJbMeCCwi5Tm7DQTBd3vAP2XVg3f0q9IA
bnBfpPaYJ6hwZD2OGUYkiv0uKBlQfPc28VTE6zBLOK87XrCIu5koHI+CWmN3Y9Ya
jEUSe7+XbIV1GwGt/BorGOwbPK7zZce4ucDdFbSklK3MHKE/S6E85dRkJghIGzEl
kjR4mcprDsPcnbrrWXE8VleyVa3wymCHKoOuYUZa0vnBseGB+lb81NRpx2bqcUV5
BrI0FVLQJhv/ME2E9pQir/Ux+0bngs2oTu4j2SqkjLbP8IlqnzasPxzOD1qyG+Dc
I1nx/7uQZgZHdt3qxXbfdA==
`protect END_PROTECTED
