`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4T/lM01z6wn9bqUP3KTVR83ufA1VYykdVafb9e6qGOioljdh6sBjUzellTzjdg8B
uySDJqMIEmxEYV/YgJleQmmw0qJOv5UGEmFpbLagmk/xi/AEy9aYWS284BQ/g6BK
TnnqggrJXbvdeR2VvBwk6QJLsxI73CHhXqWZ9pKupWwd0druugRJobVh7QI3b53Z
JP2Ocn1JWZCVS1nOsHzLl5Fkzl+JR83qPZKn5/AT5CRh/erjiZr5CsNRB1FXhDt4
5LIjibs2KpUlAu/op4tnFS037BYoZPirFatjSIQt5S2J2qq0uhFB19mCcHptm2i/
fxZ9IHLXDZ3KLRfwIPiSLk75449DuuNOw+jTNIL5MhYx/jlYYkTHxj1uq1i240qJ
yAMBOJnvJDwkg1DLphK7y3Plv2Au694wTvoixlyZAG9ct6fF+9UI0Oyujh2y5Yv/
b2QyPmEoKsMLjlWYTA1T4HzAMS4MOTRGgPXb6q7V84wq9dPbVDNsxaUsmMLSqjkS
CxCgUKq7pI5eSoX4OppgLha9+qH/2S0jXjhBU5Byn4hTfLm6BnY4Kg/oBt64NgBN
3qEsLvpMFJhQ8oJseGq+LZFYHtJTGy7pAnnw9LID/5NJukBSStqls07ecRHQBOFF
o5mnxLsm0NLbv4HsOVnS7Q==
`protect END_PROTECTED
