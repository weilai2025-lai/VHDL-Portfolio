`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdrcPLMw2NAx4ptEryfeK5XRqg1SA5Tsecrp8SGM/NBhgElRXL/D0k0ffzxEIEHy
sRhz6mIOY+NifrCNHu0p5tZ1f2Y0gASBqE6OuTU3h4j5HDhS+vJ+Yt6dHxwZPfGK
ITWLzftmw2GV0rrKF4tAuMlnNcSyTwGKiLPFQtJNZ7ibZj/UHTRLREplM0Cp3jS1
mvCkS8fyz0a8YE0cv98KKTkd9grbYNShxqis9jnOE8AC4jpXupMyAcXFZtHRQsFI
+K7C7KRlPWE7wVweoC4Pdm7yigxXYtwL17vYbePHypmNcimwyO8Ux8T+qCzfAr2+
ICKn4dzmvbuF0pb83GjRhraOf/kSXxjRdaqXuhMr0z8zz6u/Lc6vO+etQVL6TUdJ
43LrkoUIUpiXirBPFN4cfKjnaClgcaaESe7syKpLQSpCPrKBjEVVQ1/CD2oP932q
xHZKdKZOC+D1poao+con1rBFJLf0oOPQeEOJPJ66eDD7UAkjXz9SWUIegA/uN6h7
JmEENtiHXKrhzVtpJPQF5sMZXzG3ZUQofJoFMjbMneOqqt5ZwkJUqqiWY1NB1TyY
GRpKADkPK+vAqw87vdAGPLgQOzvXWYyvWNLP72hKZ5AUe2uSYVDhBMWKYodBAcMD
Ho7+xuif1Utb/Lxsfy6ou85qiLphZn/pBEuNHaHHxDncgGiVKWFW2TYMl09afqHu
D+Z8ayF7kDYoyo4h5kFX46odfW1RQJzlErhE6PsyIMf4rupTwKhqlwviLkQI1X30
2OBxJi4ow0kHukTGbAMv554HSQPQD1vQ3v9xCB+8D4bLQbJLzE7Pxc+78TI1mh05
Az2LOaAVOuZp203eHXaZ7gFLNFaEGBiqETps2SROkhd09NTn7uPaAUmng1TEYola
dO7YaaR7TK0MQyz3HLv7E1443bdET+tce4LR1jkzaH8=
`protect END_PROTECTED
