`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBYY3kp4r9Z5GhIG5nMBmiM6JlIxeYV8LPq8RceKUIqucScYVayWGPpgHBAz8iMa
94mVeh/4YsDE7VSUsOgI6Am5psJ7491ylHsPEUV92AxBmGfCMERDUQz312Y+fhTH
x8eq+otTyxiUd/6pupvNWAjsxSNaeoyUkd2tvEOd6LpS3BVjpdFP7iKQxBjnujNi
AN+aH6oDRQpnlCyrt5vqmNKwrHj8mBOLuznQ9BXsbZi81fMwuWJLrkV01W7h3yDB
FZ6jPxtsVvBBwapY0Axno1WmJ7TrwvEntZvbAvmK5vebqPwfnI1EE+V4RtBbSh2d
y8JH5wZM9XecfVp9PXiPpsEmrbfr/VmJYc0f8Q1EFkAY9SBiwL/WI8zBpd+Q2d8C
8PCSCQEl3SwFvYDRH8NwGpuRV4kUbzaxF52Gm3/b0JAeIQrK4xrXeSg2YD8G9PgO
3B0yKyLSu5mE0ONX3afgMkcFR4K3Q0dz3hf7FdTcmybQeSTPe5RB1+8gTvLOZs98
H95CEO70iVXpipCN46d5j8Z9W6+lDuNND1p3fC6bsbFZ3Qng0RzZjktiqltxSD5Y
Kx9m7qxapMRx1WuEWoWXJmSgSsRM19Rl15Xgxqo/yTxj/JjNm0LYCPYHjLNmoO3s
3VE+Y95Dx5gFOdZnyvaD+e3OB/TJ/ykV0htK0Ov/nnPmIChsqQKbGSWpF1UHp1hw
dePOSHR4lxAiyW7rbA84EGQHCBtBmCdj3frqwnesL5iEyg2+PzsjfgoknXniK0TK
Q755IHJeNGfPckCgl8NCdgY7kNxhwhpi2Ab1RekBF/B4aHmR5+FY6hvrdFiMyyGV
MyXSlpv/ymqROxFrsxNYc0vTJU+aLf4jtbpUZnsY+wc=
`protect END_PROTECTED
