`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpq13P9oYydceAfl3hWTbNmUhN7ftXINGiZKW8g3QC2K2dsccjG/5I/ilI/NNQn5
SHK3t9w6rJTuj+ppFg0+xMCDI5TracKQ7SHGMEHDhvXSiKXES3FsiD6q3X8QL0dz
nLg3vTpDry9Gg4bULbiIy+GHqIdmGq45hS8dGwCqiVkhe49d+pq0DVhXrHreuIAQ
5cu4wKhouvfgzQBDwbPod21GXSDi+QgjeN9ipCm1Lsx9OCDHdHTLKxwn36QJzVkC
Zw1MX8C7jHgjyykRfOT/gykmjTsQqIrKINZQL9TCkpy2tYw2DhsVQKMYKKXsk/M+
cAiQ6tBoKC1jntQaDeVrftlPu+TqjKr8Wnvp3m3Y2Dg=
`protect END_PROTECTED
