`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tNoHS6067AcjPtdfssT96WxS/J2AoX+ymgw1kZAdefqecDNwEOu6yfjTu4bG7jp
D9xsDW2MfFeSA674+nAbJPZTczWdg6nGRMKmuNN1tuLZskbRUEuDEKOmtMF1vwmv
njXFOF1EiYetpAi6TaQhlFuy5ca9stTu39uUgb8BYX7oD+s2ocEq4GASZrfD8TsU
xqDCPZtWfTfsBWx0ndAx/z/Hl6hPHVSsjVtoJK04f1vA4K5jeT8tYz/8coKSB66E
Z5zEq5mHK8lcHFdN9xQMglJSJHpmdhoEQIwGvqOlHLdV9M98kRJaZ5U0vB3nXI9m
bnQOFsVvA7o5CEexAJCuwoPp/Qq7MG/p6FG1PeC4TBI=
`protect END_PROTECTED
