`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17Tx204bh7Z6I3OuIXmtFfxO6qkt68hwMzxX8o9aJBXecIIL+BWBiyQCb8dAx9tk
tQKklm6GAzZntlndqMz9GXlBBQuFiEFPD5AtTruyZdYeFSLKQ4LHyAWvLopvOQFV
piCfRJeoYRIco+azbDEVucQkmgNfQ8KIQjpPRJ8sJxwSezHipx9y2M0K2zY8rGKF
c7d3Wpi4XpPqPVmaVXmuWa3ED+ygxoLSoJvprYOfi7F50hXo3/uAqdY47X1RJmCE
pFKHDJ986rKSze4kzsoRabolISyl1QEhqP1l4+k2Lg1P7O0LFQxENChhHMc/a//8
+3wqz2BRHga+Ocglm251HbCPB/K8dfGhkG/+svRZNuuEmoVRodFgAkSZwfnaUq2o
Q/To0ZUx58/KY/iU2U9pBQuToNZmI0iqs6j2ojGooRPmZiRIoYx1RJNciRqisc08
vBnUNCWt6dWYoIMvlp2AJYTE0NQopH1RHKpsq+Fy33oQmoH3oF6muJEVi9FHUvyJ
MEbk5bklyMI4GQfqQ/CeNQ9kw3fPQMNxlxTvJ+thMCGRIAh32BSx4CQk5CoqxdZ3
ElFaj5YkuDEwsPmyS/R1aylnxnGtbvfToDbr6XbtbQKV33dex2h0yK1Tx5rzVTPL
y/hwdxArEJM3M7S89E8cFtdUe6T2uo+mvUE/GO94RT8xiXTViT7NN49UZ4UrMvaK
2LWGvVwBVKWhVFPE6f9a6Hb6ee5dtiG7Y60VPvlqANCbSLJ8F8cBf+w0qCOPURFe
/7BTxdH6f7xRGiXjrbQq1fWqZPoiLHXJIH3wvlumBrfRI7H1G9wIwl42lHpB6Pr2
IqqJBVAdURbAH4dez7eYjIT8UgWAeWDutDlrRfZJvUHHPOZZibuGsG66YXujHuyI
uLMvzS5+OvKIUsJk++H0716VAMaB94Gr+tHriJGnwoo=
`protect END_PROTECTED
