`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vj0HHmstDpDwoNcPiJ/BHp4N9trhUOIrvr7knLbcDUJlJstOoxdbqzqgrPqzlIr0
rplFj1ZPIs9FZN2ztUzbIi0ywtJyEG8j6X0+2vTUcW3OhiWzWS+1ii3Pc1XAuYHL
xO3dhquadmbZn+rv5GynN8tbrtrKERGw/ScQJyBIczJ5CdYD8CrJQbai8qz8DHdD
SguPZ1GH/6KkxGfkAyQVNiYpDtszQ6BBNhF3475R2YJ3ZWdkR6qw1vBvhd/6a08/
QZtpLWytCRRCk/Lq1vnQPuWscYms2muKV77A4OdR6EL/P9SVCVl388NunAlpKAH5
CUM8pdQ7jjFHNd/08OS9POO0OaO+n+8OtgoF6yOo4mD9ojSjQWsXt579H+WW+Hg5
lmW+T3OjhKETnGzFCVn4E6O033jbXDNfVk3NxLPEHcQ2miETZRajQGKlxNxkRO7s
fkSWDvkzEoTR3/768LwbCxT4PtMr2t3ACN2bBzUBaUrL97A6/y9C4ZuBdTA5VHbU
lIu20/JvA/akd6OlcaTQ48IvTJdRXwSU8plqMnWHg0IXezCRbUMeisuHAo1zbwlV
nu2E+E3SbloSyQ9vr8JfSnDtVIUi1AXQH8CbEPlynuupKQxVX/ei5XGawNYDt0FZ
hffV0nxwv6uumlUTIrPJK8qlAtRc7nH06sGQj+Zcz0jQn9jcTJABQ7xdrOJJp8cd
ImmikVgS27HdFUdwDtvr+pK647/Q9HJPLfw4JnJMeKPYtpUjh2Me7qV3sQ/G4jLh
Hp92rJZRnYzSuNIEuq4VoPxCDDjvANuW2nzIQpkFrbvLFWSR33s71/Rmw9CjN7QZ
+jMI0C+dtlvJIyV+PdckjSJqxKbGLiUwncdw5P7qj8hSRMYyDlsA70N7GB+Y1Sd2
RAlALr7UArX4uzOpWv1R/L3Fp+aP9bnboUVDtbRiPebMNcupRgiUCCMvoNxnumxD
JLK9qilq4PgfmMFQ+VqkorGWBqaJQCzDE/3sDrJCe1JPuDx4zGEcXKyrbheG7vPO
1KVYUPs4uFjxuVwvAaXDZwepmkw3BoQnl+G6RBaPDP9FRacJHdButFv64ywRO5FY
A2vHU9ysvyFvpUhT60qMtg==
`protect END_PROTECTED
