`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sk6c8vE2QPQij25KNTSSSB/LH0WCogbXZ6Vyjd13Dh6t163mOsX2ydx+pJnUjzV4
Yvu4oPe7VeyITR5MkGLG//I/4a0vGylsufXP7WD8JjXUbqttzbVkF5Yq6u2USKYg
8g0f2sEYmAvilzcz6xTKOQPv02/dQc4rgIEbuOhYecqYbnGfsjkD5up++mPmTR20
PIMemimcqpM0qP5TgqRgpSfU7kQjfYV2xEn1LNZnjtg6GArEbc2h1g4kkH3gIczj
0Fl5kNLSiehP2i2u2V/McohkIh+XgWP8dS2JBCXDF5J06WkHZf0Mw+zruQ5OYmFk
QfHUApUPe7s3QtVOK69ZLbgnhQUf7N+mgvd5f05YE7yadkpRXRE49RxhiO9ZZyaD
rlmD9ri2R93FQ4ZWAHtgcmJKFfOtL2Zw4ajK2G9HzW4JDrHL/CvQJS6/EcHk8gDY
puX/9qHd0UvPVcCwBnbOzKlN6oUcXg2Xk3yuz8GTq54SYhfU3Aul1vju+qHnteMt
gBaUsER/Cf9pgj0NRcghjKFeCUOaB1uhpPp1reIuyi3QxyRKStaZJulG32iK7WrE
0FrrCZm7goApBibl9gf5E+8VM5DHoVjJEkEeCce0TXobd5pZ0xEJO2y88uaguhzu
Q8KA/cufzmBhKUk98RtldmbOz+uPWTvn+JvYGJmYYCLvQz7PIMCnCBHvxO7vFnNH
DD9c1QZSzNKwBMWLPavjGxoDMgF25oGCct9BhU8wE5o+jI3DP5c2oxyXjxQ6X1U/
JaSBE2AHJjXfNMFIhjvG4nQ5kVwtWJu9GQ6db9kLqYY0aeGSugAOz3MsuQn5f/gC
2uX2AiashSbQ8TVYRPp6HK2UOnq+ITs9NgJBMQcN0evbh66yRqW+ZJByWWjBbrZW
+Z85KrtiGvhfdpXVwqkQN3MxGpz5TedzRg2WnkAJbAE0k6mnitCC+BjXCsi7bf3u
jLF5Xpl5KJcF2lc1AYqxLaBD1e7xrwh9RqBm6fAsnE7dR1fYGeajqXNV/2Sc6aQM
NLIzpUmCQ0RKif0gIoeHHeUfBPZrxJ9F5YqXxiFm9OOt9VqT+XBuatOS6r61eFsC
AW9iDMvqF5ZyaAn5q+W2ejbdLHUamsj+MJNcpQXVqt5uibgCZVGUChOWx1fw09Zk
EZGfidDpoGOkWY9Ar0bVQ94SnpaRhAV/HLWWb8c/P0V0bYmRoIAJLJXC7GRUHArX
gXU7tEqJ46ce9St8Ko8nEaCiutk+fBVg7jo7mqsP92KF7Q12cYTEIvjYLMCvBgFD
0xHqyFNW790s4kjAjaJx1qX/tMc3N/UuBGwH53KpXOFF99hgAQP2gS5Xh5P7exvI
l8Z238xLX3m4NHfLbnJqWKdviT18tafuafl7/ZidqyRHn21vIXOlhNgAGGlVtqlY
4kb+cZsUG+oH6WLt/FixPxj/kFjwjFd4szbLoyjrVFMYgTdr2bHR1xKsYxxbVmwb
y98lak3YWjVmobFdjg6BFLCFE1LU7hyyOM1B+MC7XtT9qORiF8tKbISx9xsrb3bP
Pjau3BMURj6ITKsB5hJH9q2UN/U6hcoEH8CgmjKrTY++QyzPk1GE5AWvafEia2XW
1MXGEG7awUiyq8/DUSExJMDxKQnW+VfIbsWz5Tks9LbH2aQbLd/tvs2BOOTPUV0D
yaSlAvXuUHejSOM2lFwTZ3/5M6CMGchkg3jLEAHGfyxY4weWL5pusROKeXoBzGC9
Xjj7f9qDxL7k6SxR8dyqs8DJukbk9+CeOkgVGPrwMQS/CR956xV2AE4/RlQbBiNB
k6G4WgOmYl0wL9Mrdsn7ajg6uvLjw/PkS3aZvWtlG+08Q+jLcRvTSfZKwH4b1kIQ
d9Pyz/kZXXdqOZamvaJolkLH/pQCBepXs1aDtPkzVcdOV/E9/XueYtv2+/vJM67A
NEiej+xp5Egha9zdn1EGlXqnPPL3iEXZMWEzIEs8WYhZxBsWyRB/kC3c62Efb8ev
TqLJK31Eb6I8cLPrYYYP/CImYNC5fnkmbLGrWyJnuLGtj/nzENDvR4ODwWVAlnhu
0IRprp6+93WcxxGvSp9xNJTb8qH1DgpVyzb1gsJ6b8yl2KdjVrySMBBOdSFS1SgB
xsMXDso+6O5NlSFsA4pWSpHs9QwRAKWcS7lp17S/dPJlsiSPD7K/osZdy9eA5emQ
rsQsPEVtIsek/PoG1/LEjCMLPIaO5Ggc4QC7WGd3oHO6PzB9G/Gd63IBOOHawRoZ
I2hH08YTJZEUVbCt1UBPBvK9l/nEx3XtN0iYPZcrVeiCAp5LbRgCrqhZmIkaQ9/r
olMzPimrrsj8CueduDzH4JcpXLZLh9k0pDNrTwFBycNxtP9HrJaT+iYNLWVYFNTw
Rybck4DTgAGJLQAth6b0omtKGXuJv7nFGeiEMmdE1DzqTQKvqzx6eRAuv4xO+g87
dG7zkxsynX0z7Y8daS4Dde1kMMWsCAOISyxZ2tL97c4njxcUKoSK8yDwlkidsogc
qCpq3vn9WN0egdpTwQ1GRwdKUMKBiivjs2aNW1e7CNhi3EqrKanbInplG1MS06jZ
Ogq1PTmS8yP8VC+Uj15JAArdJVGBkY4MfEH1muR283x12N2b8q1MvxtRZie9taoP
tFoq91ZP5ENfKRs4ZrFlaT+Pyi0jFgbwJQCOfEMDX8KNXrk9dP1VPI9RUH34TEyX
cUyaNG/pl/bVD4TWM21PtjvPT65L+DcMtm0fZELqTHTb73L/hquoipLzqKTY8O+S
Jr2Rp/XhToeqtFZ2ThT4LhM0aHH4jn9vpSDY+xYaQVLegOd8ymBEGIdijp2mc2p5
qyE8cjmNQ0p5Vc2seDkMyInX7vADbX1sNu6uWpkc1L6JJroXZlWZ0z8qvMayUJmo
s/SGaRboEtl97a2k1im6yFksjuiGkNx+efz+PgAbSYDxEMTPd3VTqoN4cqfp2Eur
QlC0a35QO0jNb0HEkzH1S2aAt4UYXdM//ZYHz90aQxuVZ8PWsyiqSXxgnnjfMVdS
g62cpO44L+ELSXWnhctzLhyJK2LkZSwmEHRKN0LB1H0kcJ0FqnLxlVrDlvj5z5L8
TyuQXDIN+OvVpiOIF57B42vZQeN2s3lV/u5X/Gbhrolo2jDk/wklQj9VQ8MQAiEb
c8vbjxEgFcO/LYusfRN+sAPzpBdAQgr/OvLCOhLUhkdlBvuZO8tEkCEXYlwVFqJY
DgDuZWyGWaz6eWVg/yxKcJJv7HWXln3IkkmKThuU1cj9GtST7KE8Nl0eUDSVlrc/
9WlhkBLJgzhL6BGu2DkJSUA5fW1YRGycj9Sr6fn78xnhs/CXdJfMkKAC3eozNxFD
KeBy7w0V2kHQ0A7++YNbqex8U/iOuvHSFHqyHp/hBLAPwJSVpQAhm1FlICeVoAnf
hXIfExz3EjOLM8eRIQPYv2hWFV4bQOlaJlNYoId1TwKj8iB+Sv8nFCvxteZ86v4z
B+FxIQJ8fv59w7geFi52ix1Fl7ozybVqmYiXOh42c9d8MYdUTPz3o8vwtWb9mLn+
nzNW71p2EbvWAHFLgAQ1UP/CgppTF4gdfRJXyuDZHkHlRCtm0rTCSwS7xZ3hNCUK
USNQvSehlgOXxZOubHKWWCPpZTgKzC5p4YpxTBAYecPRLXMgy/GDKMlxjxnXjq03
Qw+2iKdUaMn6iwirtV/a14fIlnm3NXuJwn7xk/S38JzPU1NhlaMEDAPd/CBw6zg9
r5N8pbkqneSGGfokvH2YpULWAjvYOTUScl6TfkhPxqdCU34CizOzbHbYKXDLAi2n
PSMPXSzH1YvChdhwZ4cfhtfWQri2uGoM/c5GT1kn+56ymMBVHasXmoJZQwdk0hcv
+cB5UwzwHfYwcM0knzG9bG0cNaP/BwbTcUadoui/8NtLQGl9bUOcD0/Ps0arJRDf
N9V1l8t8B5dYvl0jEL24C/OmtPswBxNhvShIEk/+rwBchqiazsbzgojmD9gMnnFy
hwyFbK0MDbsF2Y99wo2/0dLFkJMkodhEyJou92Y/bn0nhBXZJBuOyZvCiPn+0a02
kKHJsHh18PvaZWNByx25TZNvBK8nVlbCDFb5nv8rtpvqxrZSARVoyXxg/LoHcMJg
l+skgY4u902p1qjuQDyE9GVrHYkZJ1m9YAkZFk8s2bwUHgHrMg1OCBCgo+Y9AZCH
zU4mbhzzl6lHsDLDpConXkcS8xyK2kKezVcv1D8lAaklVtArw6mqkUNDb1lNU6eB
sTi0TrSTC7aS9zVv5d29c4SZSUI3MiumrZTH/gVsaAK+VhuhqssX/0FNSOUYnkEb
qR/ovbol7A0+19uW/m8aXyfNFF4OPlHU+ygv9E3Jc4sEnkISQJhJb2T/P0mLMUZv
d+l6Ph8RgULCxM+xqSdk+JEhkyiCZOunsEj/G70S2ISQz+8H/IfrnoQF6goXzHS9
qk7p02EFt7/ReaERkdiHVYjVsLupGndcSsaSDxl2kAL5eNzTENrqq3U3uTZCxVSh
36nKhKkz65wEiZ4b5cxLv8Vgtj9OWUfaB7nQob35ueJwSJXwHTHoUGu1co3Fp/pr
h6Uru52pneQYt5LI7bMD+NatJDkE024hn21aCXTY9Ii6+qJfhg51CL1BfQ8zfUYK
jY2HFXwjjrF5svzTa/N+JCAJZY4O/ndfB79ulWGXll9KbPwCWRj04rt9aDlnha3N
FQu/fckuhaKRatEYK2Ew6UZleVluNrF5XT+mwE8fHldA0i14NpX4ArN/GW1Zee5j
jcTkbSK9HFRSVYu4P6rrQJ85RbxTGQ348nYwHuh1SevMIm6qMFsASB2d4KyYu2Zq
VW0/1OPxzqzsIzHlKTDgfH7FXdi5/2YDxC+8HKzYbotN8kXDJ6LaSVgUXvrVkrCB
Iy32Zm4t1NnyG5FotNdRNKPQEcQrxL95m9Su1VoAcRakeqExYxPFH4M8x+j8uSRk
Y2nb3GcdZLvbtAtgrGYi7uL7DEM06GEbrgSOeSswd3XdxSaYw600XSBGpfKeXnpz
lOjDreJGAK+fwSRfpc2QYJJBgBUG+WkMn3L8xOpt5yrHe+dWCkpAxUQ9y/VzeL9Q
yJLFaPS5QF/O89Va5oiZyvBV8WrMTuQn4iR93plpPHFYL/gXN0Qv72jqPgWrgJo4
FBu9i9G4tN/CNaUDGeesL4mYFHcS0aHbKOW47Z9R37U7Fzuj4OSpqYoTB5UZeJJ2
KFjq2fMWNztxCV9q7uXa2Sbub5IMb15s0b3nlK/g0azGhwPgwNUHOcKi8jUa9Kxw
gs/8NJBDFG7dxVJcwvsqQKyRhFVe3vcHP0fOzI63jZxHvShDCwFuLQ1XM2YpQ876
kLRM6r47qYVTahXT4YNm44EAWZReSbOU+lGG1iuxT290qIbSr+XmVndFiyJc63Np
VOuDuoU0UdqKuTW3Bxlg0r7cTzFo0pdLpfHg+7WnFeLRj/MUowAzVPC3Uxa4V+8B
xSYlfdyMTFxhCMjDRl7PAx7Y6iTynk9M2zMd2bUj26WwlhE1dxhIqmzcuK52a0AK
eI9LARx/GWQqsrmglo/Uy0zm2+M9Ojugj1RYCW3vy7XU0ikANo6bGemD4124uwd3
rPpUN8VCgPKLFSCMRUOgWRtxU7lrfehiSgysVhux5dTh60ylmA3YXsDrOtCiMxRt
+9Zm0F5uCfEsTxqnsnoUhyk9nE6iA2bVx0VU3ScUG0V9yRL5TINAE/5rSq0IYfwX
t4JegucSJ8q8Me3JDQsGNKl/WfSVwu6K8YsTS1WkX8tG150+0tBnOadp1QApJaYk
neiL3hsUsTWD+Y5E4fHUDv24zFtfhEJKB2FMwGSxECqgWnKpyeqUhNZROM4xqBWk
9tTbZ8HUzHBSn9uhqfJO5MiRCUr5gtdG+qs54ZbNIl0SdFQus0VsH+yNG8L4au0j
TU21K+r4fj5KPRIm6yK1syHyVbvX+Aa9ZFNF2Mwi3RmHG4eYniZZfV5VbI6dUXJw
D3ge4S2XxgFOTuP+EOdj/JN7rzmKBq1d/HUN7hn3c/45uaW5uOSh1hg3QU/xm+VU
aB6GbJW4f6z3ujCmZdNQZaUDNqN5AHDp/lspZR7xioV1JAEj9zI6QvVTYAndBSjX
`protect END_PROTECTED
