`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fHz8InyDlbGD7urV9Hai8zcRbxQ6cBjo3Rn0/jW/p8zPTgbDAiCkVnRAEl2nsGF
HvCQLqT1CucZHpc73no18mGuhuVp7PL6G5u23qNO18Q02li3ON0pbiBYo9xrEzpK
U0Vcet+lmdcnw3W0fASpQByM7cpId2/TIUEfT2AiJg0pgTKiJk2WmlH9dQJvbyDF
WXKk5pzdZIzXuBOfVCruTqbjbkLCgDTGFP0ROeOEHZO4XnD3g2oekZ54Vzo9jUoe
WOJ0kxqevQAul8LC/GinJhIAZ4f15tXuraWtifs0+uaIwP5lO9tM7wSH4bTrX2v/
KTFKft2v3lwTheDc5Nqqqsrk/ksZ6scfFHkwwADmoQEqEoYbwcBwEInfcn2uLILo
/frsfAgmti8lpjlmyCDdu4PQ9BAebuRVDV1otfive5XVkfzbivnVaGw2Onh/fQf2
B5/RIqsojAk4t3ekd9t9d3qSvKBPckRcAcXoQBf4+IQr3W94Kk0aq9GU827g0vY5
GuHr5EsqtJzdhz4U5bDRxWvmn3Bq1QNbblfjmLJeynKrzjQHcSTXi16vF01uSlWZ
yn7qiZS/EB3HR90qPbnecgMBpdXDDgw/gOTszPnSxUPwnK/GxFDxoEuT4lPmdCIU
OsrMf5XFkVRIMtuyrfZKcbjBb973VbMNrBU99ATefU4cqQg9rCF9uPrb3c+kRMyb
GhV4sd6fedxQGeRPSGYM2G1dIT1UZdaZHPzYMqhEHOZu3L3cBtpj0a5zxq/X1jHt
Q9nRAH4BNiRsgckvrGZCLSkj0HjgJP4D/ob380tV1cHcVEfZRg7HqyqzoM95kXQ4
KUNHzi/SLtzsFYfYHe7y/kcGQxFj/EeNbVfscBfUvjAbWz9EF8WfdPcfgGyuUjsv
iPADbaggr6yr0KuDThnVORkbPU/omuBpzwr4HdWBanEGQ7yprnZ+u1KIkJ1JjGnT
aI1eE/SPPq3p7ynBAKgVm8FYZi65xIYwrhaOwkSvhGYhTkheTaCmxE5LytfdasGw
/1WsQ2G1yCMowZfF9my+oue0tpqMBjpgBKOdPiBzxIN4qHOoGwPb0zgKyJhIPl+R
ALANokb5zRiVyO4FD34vOXBdqVyBHz3VaAX9HBBvNNcWubWObs4wSlgIH4LNTDlg
xbiWn87f399mQwbctoHB/6D+NKKoHDcl5LLzHhBDko3A0u3vdcfWJv1jvL6IlJ69
CXYsYsj7zDbCqcyoRQMTCbIK3mPVTY/PL6HgzyF68JpciyzA/2ao70XX35lBXu0q
/htTU1igZv2B1gWAuzRhlmQvQXfrckhnvjh/FxlU2RGaZ5sRA9IM9i7r/ZsvXf+N
I0QPHLFFmAepZH4Il1sG2W1QzxIUO6su6KD+L5yfzyfQxmkCRzVvTnWEkEWqZ1Qr
okDLzNnGxH0dX1Dbif2Cq1PM+7ZA5U8esXnAblxUFHDrqsN8dmthr6q29gPGK751
F4zEp9c/CldfsUiC1JLQ+sCzPv3jT4rJehTrfyGOGOGqE687K2RN0T42DswZ4kLG
69LUpwuq4kcA26gF2v+C094skniXMKbU8oun5NR9EBhPIkneO5vrc0d3ApD72lBi
YKcOc3MefaCVahdfYE3mGJ7TZfaYE456oF+bW8Gv5dgAFQlz32SdgLI1+l/cTLvh
f/vL5sRBXO0TcXExtPflK1XbBBb4Vm8lqVboT7B+7uY0fvf5DGXjJUzmGU7G2gPl
ZU+3FQMaRqKpjWo/flKMeTE41lEJNQiSKNxDewF0if7TFAE1+DKG5Z9WcJJ8QuF7
IIdCL+p9c838X3JVh1bMhOinhE0I5OfPGO5SzZDQmX30hhRx9zPb6bP+/9wJeYXr
LG+T2jsgXorBFk39iifpN9eiQTv1mAiTlgZpo/HPEiLhQQVTaGr6knBqS0IJO9pr
zYONdAAtqPth1lSEuqGzD+oH4OaukPynl9kim9CgPCa0SEOK+0wwZl/CWg9cThIP
JcueT9OfQ8YPv9MuPEdD+8SZ1DeV2MPc/w2D+UyvMeMC/+MNn7ou/w6BWWviQMUx
/5GJb10E0g79WTshoif3/9NXvEom2otv7bm+mBwfMusNWmaZNVfqD9slQBGqUeOs
uKC81ZCqpkwF9xouRa8Tx+jEsYwv9EIT7PfdYR77C7bi+Et6Rgnt5qx03daqzzGj
fQNLLJcoOaGsbdPQIDrfLicLDVj6c1cnxow53C2L4+5kjfZ3Pp/7cp5dzuh3HTka
yhK9n1tjg+3SF5lMezsDj6vb8Hg6jgeCkq4HvNDhARdgA1fLTwIuLradWEkckW8g
Utp1I4Q5T7azOr5o50Fk60cisBbTM0H/yXvWWcqUDKRlwpOACxz9c13+dIVjhPeo
9VB19ZDvOqMdrIryB1TUPqtNT+RspIDNSz+/TuEIj/BP0J5M5sOG1zbQwZOWwbcc
usi4xrWo9qC4vl4LLrf6eh1IczZ88zz2/Wh0kUs59yuvjhTuEmxjPdhPoBJCIRd5
m+A965w4qBCzi11whjNCZ/SCz4kXkWfZBcLYNHM5wjFttR9lYF5jEA0rmBsZvrVi
DnDiJ5Xyy1Ekyhm/vb0vnMKL7X+AlQAkZ96jUY2TixArKNn+Bh9AHpMPvyvLXpmI
FFCrzk4o8g+yAuFvGQDmC46lb+XCj3HvJkImy0rE+C/7RMJ/CWBDNOxTpkMdtnzp
AhfkhSfsf5hP7cjYz0AeFz2byIuwXt+9i+8CsKEF3A9pR7T5zhCArobCDiCJ7qME
TDus2+7BT9REQKT+2X3NZKCuigQZZI5HOgqFFGstmfGMveYUeJyfNWKHtFbgMxhU
ARgWBjMNOLQ6ab4hTPc7DQZP6Y96kLokN4ILhQLO0vbRYNVoj81m9KDD5I/YOsI4
NVbNKFt3F65zrnYp47hTsGsjG+TwO7nYfVD7lTLJJMcM0hZ6j95Owc8EqjUlZgd7
CrBHrxAm730b4rgBGJQaMkXh0MYseKgFal/5X+F5NI1FbwZlkGr2NoCuHj+RGypd
zmYF0kwUZrSXz6YVr7EsfoVoVhAhglkSQeRz/nkKOgQ08LYyyM04B1DGso8FZ+p1
F0oQyIsv1qcEpC95JRfsBAhqJGeq4sb0IlNeVfqxDPnrHxgifjFWkxQnVgEApJCg
2gMpklZS85ADVW0fMCXSgtXa3/kuy+ZnfN4cjwXxTMAJkiVAhBVjK3yhUjytTqG0
edpsP9p4nPjVUgiCPZoGwzYoevmWEynkgSKyQVkI+YbZ4Bbz7ixJj4qjBYrmYGXH
EmvVe8ZCXzd2fsEeKgXHhxLz9j2h8nzcZf6QkfZwio7xcsXxrzeynoA7fvwprzH4
D337edX87rB2y1fDM26QdtZiljQ9lr2mIVQ87eg9a3UJrKgR6IwNQRjVR+sxa7h/
TMM2cUP84ivQDt6CC3busDQoeedmFtEGOsh3l06ABYZhHMpfQ3Ed001OvvVm1FcM
u+X5XvKHn4u04e5vkRQjHVN/N5Y8JKW1SxuGeOlJzo9KhNOdr4+t7O6SYaE9H6HS
bCF5jvEei2lIn6hRAIR8jRApP+rJ6skq3icKAk8B1w4IvMiF7qE+B8Jp1GWd65br
iTmSH5FUxrEsVXNPB4I+ujcj0VN9CG3bHqn4MRTaB7VvQMlpkQXxQSpkNej0rpuR
H1Hdn6bWwp828UJ67KtpCEY+MQkJC8akuwztNoKg1oV7Ux6iJvGCa4MdplYWVoca
aSWU2OZ/0Xo1nDOAarJLi1k+jZvY/N8MNZGo/h2j5k9O3aUWRqkTS6u9z9+mGOKW
d3ufKdP+u+BfbOkr/HPnnDgCbPlDmYQbApy2TE8Dkdd7nxWC59uiTcqIwII5QwuF
n21yr5EWLQMrMs5mlI0RgrLLSe9MH1oFmTlYpcxDW6tTkqqCtydX8B+pomRaOmIm
CvlIKXbtg0dbAh0dWj5CbuwVBhOhqphi9+drDUAfJTN/sPXj52fSwMRlem7oVDBs
FnfGTXX46Qo8i+LY+8yDg90b2c0RLpB1BgmxXHsDvJQABRZWSMrpoq5erjMOPGPI
PeQ9n7siwkLpt/huz9/RqU85tbYZsNAA71IryOjRGt7dN6/P/hve/QJSuTAjv+n/
7MSLPzwlewB3DMwQd3TN8YV4b1kREH0vF74+KuM53dGG0mQmh10zwSoGlRe+tTu1
IGg9A2MsaDQH9bbUgBa3oIgGoNyRAgcmPpKAuvFDQ+iXrBrhHnXUxIuTdiAs7XQT
Waty98z+hlXULLG537PmH7h1OTNNJ/blFfU9o29dW1CPeayxXqPl6qBGk7Xs6tEg
oNWRIorX+J0TPbyDtQm3jhTLn+Kgo9K0LmVMdzw3zzT4cOgFQdYjw8GRjzVDdazf
QV3iYHqTIBu6n6mAORdFk2lWrnixWvcJ5D/5N6VMaz8=
`protect END_PROTECTED
