`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBEq1j/F1x1hNoGg9OQjg4XFGT0fq4BAW6qOMpFmpNdk50U7u41flCcINX1xt+6+
id0JabYujd9At/JRbsS656XnnLHtM9jqYX2UJ8bCLev/dh/NoKP2g9GbN9Mu+VTk
7Z10AoQqjitjmDhBtdTZEbqxmyu8VmJ1wk4SraBMjsrnN7UiQQb6Rmr/K1/yiMwF
U505aIXAJDW2Hole2KO1ZO44yDxQQ0jdRxLx42yyVZuHFACnJB56jhIzgjIiwuIz
Oj7eNoz+JS1X2ft2n0G+L/LpUwhfVF+FZJMbWDCkPK4u1o6dnCM+6zAvX3j4CU4S
CT//VXsgPVFnNYhfBgOm+T6ZNbI6T3G7IOtG9sU8l3XA6dWIwGJlc3+9k0M7dP9h
casY+SuMvFgSKF1ZMozEDF2rqCAgTMH8Gwb9h1sIYZrBnb1hjskT8PuPKOJjRIMR
//PczSFGQQA0qyLP4Q/aErx2lN8lfPx/S4CgsjIBtYgJWGKfW8HhtK71RF60tSb4
WNmbjOJeSF+XltHprsRH+koDCpiRcT5UyDCMgIXZK8dlbKsCNudxRMpMxJvIaF/o
rYBq7OOsgyKtR9etqKtepee2ufZtcBZXPNx79SN52EOwNi4w11APZWqIwlXO2QBH
J5rD6VhGYWzoJZi7OtVwl2IaT89VrPxalkKY0NuSOrjz6mWUrWZQ69R/H4qbrI4C
uiYSJTS0kGPQ+G0eszIs+cgzNjkZPzzy86brN3zVJ/wzC1RjIaERkxtenj2LKMXu
TBt+i1asULborc4gj+Lh4WtOlXJoUUutukMwK2NChVVgjZRefoHtiYtTIKGyFzMX
rCmHTrm92zwzbQTYgBkk1umXts45GWmvbaxhUurBqeB8YhtqrPjFxguhNvyaK8Jj
DSuaUjRVEdBJPr21fpUX4lquViZ9kmjX1PKzsjvcdgEwnGYCdV4TxB5lrtOzvrXc
d/t9wkywiwVlyiHHN111qk/x6ffD2OKlF8ImvT4tVHm/WW892h1rp5TG1ayXdq7u
lJF7IRIIdrLtnEa2nbX/GWnP81dWinwy7yot/yBDtnGSz66gTeDQ5jEYxPPXd7Nr
ZiO1wBTNckXvipbo4Bd6WLTOzayfNHfD2eSLu/zHeBlRLRwouC+JsdWJsYge0ZLW
R1v98W+m7u8TlGvl30g0v2UKCUvAQGJ2jowlywb/Nyp5eOYZxK0hFR8bWujcoy7F
po+x4+ERjAiO0TSv49ReXFz9uDq9T+OsjlgzL/C68j0M0tn5olJkJIixPq+klyvC
9FkVJz+BOOXbkcErR2qkWTfOXPx1k+AM3Kf1ScqoPOK5HV2Qw/MFmusHDEHeADhh
CnHu76ZPQBqP6MPGfKAH6i04HV1Tuzi+livZxjLuZLwMtSeviQK0m2o3FP7MvtwF
H/PiEhJs0Hqtb3cdkC+7jxzZz5KCsMkmOQOWp9jzSqOUwBizTsC7aIUXAR9cLqM2
PkMGByWsT8hB/4ndKtrzWNd+hGNSDS7SFSxvbhoG5EkNiW81usinZwFcvpeXdt/2
zS3WsIuHyQBn/3RHi/iPJM5g0Wv95A452EHie5Nw2jglOZkhaLfxIldncdUNLwJD
3LhyIgOH9xOOop8EN2b/njUmoTnjSJKfXnGqQKUZ75Evuhiiz35Cag1PShPjfO8a
h9EHD51gFhzqSb2/uNeFcPyZqqp5NYhugYZxSTSHfI3imsxomRjhvAEMKym0AKPp
b2dKwts2E8LTjvuusm87jZl0lM5SbfSFFn1L/iAkt2c7F1YKRL2wM6O+BZ4tGl4y
/y7nUgI3YdHkvvRjxN/5zfwTWuUQdkSwTLvfrv4IYUIEsEgNrKDof4a+dKsQYW4N
8k1lW70f1WwRNM9jz1SjNhPGCTF7OTxw3snbBgobYaoFwcG6u/IoALkD2gkTffui
YVQzetuhFyP4i+XJDRx+tFLQizXDF/JCkjBfWHvoV/TNnVpoHVokW+PuVynrTZ+A
JjrP6tjQavniWm9oRJbqHW647xdlsvwetNs+XkYfLjgg/gzFQzNqWmcZVhgpubaM
eKpzKtaYkILsDJ4XVanSZ6XFHYQofLicA0RE/u1eTJ6WzLFf3YxJNYRDyHCWoDW6
QpnYl3L0+T59JpcOx3YX4OEb4sgpIEnTN9CvmpL4OrOBRGR2TC707aympBUYSNMP
P3O6YMduif1ckEqNESOFa53BdavdwH+kt3SQORqdsszoVruvto1iKKtKWwDLbXfR
p5AZ8N7X71GZ+Cjn+s6HfkCeaAs5afP/3LTaYgHW5usIISDebBe8GHDORXRDdtMf
Oh2o5irGiDi1oIB0w7wgmsOppPuIMAgM5edqYE8Qvb465CLj3+MlgCvhPX2nGdsW
kTYaMHccBgq8fStrF4nYTIxRJnmedxCOJUF2G5TVtz0IkWXVNzRvr4z+JaOopLRN
v4zL/RcCCBQGvbbD7KsnPkt6Vel5wK9H7V7M+JgdplvafW6Ana7YmnU7UNfrSm75
nRwMgAG5L9/eStbUL+fHxiL+GYxQ87ynQ5keYBWcnKGCq7JDjbVYntH4AW5JnPur
In4xWOVFQIxU0z/e3qwA5TVGNHoMrS2mHz23GUBQF8zVQ7pwr0z9ZcIEzxnBqTvD
F/AsNdKA5dKATc900T9dnGOSocmw2lXL9a1VyKfQTAhD7nA7OpdwrdnG4jinJYm6
lQUxxdpqqv2BK1oFTy4ohjui0dvXlfdNbklMyJO34GeNaqFlqA+lPLwVyMYr+pcX
JefsSWoXs5vRRrkb8znVmYiKAV70LrUNig79SXIlSbrNWENhV98FefbQggJCO3jN
PLUEGUgbPQXl90AxPcYQF2tPDmpky7EYuJMKlRr/iB+Rh6GJwLHcHcFXIoFyHEgD
4TyAkimGE7zvoGWg2larG4LMlxKFfZi2drO3hg9wy5bTIckcIjozKpAp+CYgxicp
ctWbENRrJfI8dSYJX+ioEmQZ/UDcVq+I0EyZyd5uDRaQc2v6jo/03Vg2QjRJEDd3
zMu07W0nHQ5suhd67trU95+d/ScXfmaJB03rkQPx0VZlMqwblEx1BDL1gv9T179t
Em4inXyJC3NIPuZRIiLFJh7abDG9z3nNRslef5lFGKQBZzY4gFPhGmsPujs5unvn
rNQxclMw5mDC8icvQf36LdXG96eFc77KbRw2Jx4HEy2bK3CSh0Go70n4+uZ/Qdm/
74q7YPLl+PRObjX8PgGToPpxnA945G+EVlBrRa/aFUCddqh7O7RRe0uiepJjkOAB
wKbwojSyMOC1Wu+vOa5cMLzjuwf73KbLEt5N8krKW5qNI96+VRt9wr9orI72NbeW
MhM6wJFoA8GCY7o5UurRPs6VsbEOIwC1MxaTKLEb03eqBSzH/dGIdZ4FIzxEnpvL
eYXTvTTtrswFfyqaSkZF4TQAZeyNbOX+D2lwbDhzQrW/WRQUVGf/j17uOdCGWHri
+k54Yj3/IIVXZ8ZnZgryRmB1mrMOsSp4YHw5L5QmJaZ6asw09oGGvEC8F/vWO5PB
UiSxWJNTTVMtZeszb3skRd3dlquYinlvDHSp/UR7hX7jRfY1Zwd4I1E2N3EXhyxt
9Ct70PiUS5IAWGR/iy/XPZQ00O2Q5R4q4d561O+IebE85RWYCFP+AEp08CFIzXRs
sI23BBXAc+589u3D0UxJ0dD8sskLpeL6GtsI46jUqp8ZFbSmQuzapoAgW48gPbRT
bIbqZS31TQL3+w+LTEguXPSGeZFJOcsTMfPH1UEiJ8nlcoVhN4NGtYNZ/Tu+9YOe
2XPk3jqcBZKdgEVJq0XUwZDnWE/R0aVekbHyXbPW4kBmF/p3XpaRzH7jpWtMg8G3
9WCuq9wg39i22/y+c09bSv9bGBPx3lPDIYOeRTr0YyPCc7ucK4srIjQP8zXVM4gm
KaVhTcp3Ci0BjNZmMqsL5E+7lL56KPSIBTJFY1VBGR5Vt4yPzNMyWPoKWBjAO0Om
7wQ0SI4FdKiqje/ZK/6pGbCVE5xroNlYBh/r+ontQFBrCFrw+kQv7RoE5aeShFaG
WwLuPxoB47A9j/3nJXc5ZwEgx5n+objUqYDvWI4CvmPh1iLxvBEUwisJ6G+VxBOx
E/c0f2DobXfdNsigNB/VzxjXjAOBKRulosj94+5KBD6JMBYLsWzDPWgvwB+054/S
mnoTrw5TvpnxEui16LLjnE4EZ03KGmA2v9gij2GzjhDHkAjVBkjKbSB4+LeC31Np
aEs/WpuQbCvFA/My/oz3l2d/06gaXoJ/AXI9OAVb5e2ejDrqGlpLE+eedrKyv4qo
EryyF7JGA2NhBZHbdZ2DJPlfY7DIcoBt7uhmyB03Uh1ekwv6EC63Ym+X9WN17Q48
arm1iw/gWBdh0q4O+b9oOlRvrv5w408iKzfIYHbIrgKEWehtXWhQJz4YHWnHIKEK
qjXWW40NJX7fPNdK09RVoDEIbdHqa8eoS61B3tEaIm940x2HQXIVK8BfUCDypdRq
TNsfYP/8t6Gi/E0HtjBzyN3sl4MOJsEhlXjklTD1K4YDnfrcNh4CSKYD46G9ji7I
8xFPZmPYMqf2YpE2T/IR0SqCbWpw8Aymmiw6x4n65bd9U0WO6weTLrqJJzOCKiZP
fdEi51AwvPgsrNFVRossGGF1l+OaluJMjDlwjz6i7eKU1fV/lX9ua1jy0shgr2xh
BHOi1NNsGscy/fLvLjGzXwiZ3SZPTNtBIp+tNWXWG6zRRDNFQ/D/ST1Ef8cUzSos
m0RASA5sdSuFXfFY36FBsjUbxCb99WgS+bxcog9j/zfx8TIexxV2mohvuERtPgHd
ok9WDTQpKYQqumw+1XsWztjPkiAreJcXyKtAE5WyWcmgsQFlv1zXa1ze0o6Ngifc
2WM16iYx6FOlu52j34yOT+BU55KNW+pJuWifXZ0qrOwZH2jymEbN7ol1VitaSMJr
k1BqZQomWa594qUboq3SAU0dYoxRlmPo1QqPLO9QUO4fJOIJvZPBv2rfTkIAATQ+
bkVki17AatpUxWWaaZ1oy9bgc+bH11KVypq8Q+8XAkKHDwUzEDrwZNWYwj0hvYo1
OGbG6+EZkqz4ObZrcQYbcQd0gQ2gsFIl0VHtKESDmg+g3Cg24TkAZ1YUKzTdRCwq
4rtiIcd8tNghc3TZO1s47+M5EVhz5ddpUesrH6NQ640HDzJlKgQAk8BG8oLqPMG5
wr8VQNMCtv7Dz/xbKTgt0588i5Vx1JVriEsTQzG2iurhYrKByzuBtL0OYGOms4o8
XUpJFW5AG8Qvm2adG/JuItKMir9bP1Sgy0q1cXv2nqFOH0kBfpNDcp6EBpb2A3hM
npOAU9mSjBrBRitfhpwOxIrf1P5wFP5FIco6RscTDsLqeIpCthBwYktjNqRS1a9D
xrsZH33EIAl4nGToobMC+psjBhqnMNbQ3ZUXPvhp8nA2vGZmbHVQBzYrI4Wmdjdz
/k7MfJ61kTl7PoLbbnQ4KVrdADsfspEyEznoP3NUsVOL5vjWPcSo+VqcEKJbG6Nh
qPwXOc5tsCVCzPdtVG7zERzjuSiVtcOAIxY+p+chmNKz80f0pmX9yVMl+HyipbdZ
By28I+rNBl2lUG/WJjto12OiBt3vf8mb2aZP4dRM/GQeJcL7GA8PQvPURaIIZ4Gn
6ckWlsPkTQBfqNzHlL5hF/PTAXTAu/5QJiQ9GdGFuX6prZy4A6/WksHawyPY+Qh+
s0lcD75ztH89hK/B1bjtosbKWCNUZFyHxbsukxZ6g5inlRE/Zkt8JY480B9uC/Cv
z41F0vjd/gZq26LnVPq037DioVqEXavbcVOcenC58Ui/i6iHe1F3HMxXy/y29x7P
sAdiciyvy8iCf6WZrMndaMFyybRtKUPzmwAKQC5AngYS3Iqm5RH3kFNa7L/JPj5w
8k6z7g7ccLFPQvGNhcSKhNKJ5us0OfEos7/w2gZG/7ukv/AEgSKsNI+OrfanuWIX
T/2hIS3Dhop/YCB75Geku49KGkARgHmgbRsdYyJfqzsoXFupVdroH0RDZevqvlID
feruotUiehZ4gTX8e9EgzPoSZmOhag2WJVyPqA9ukLF6pbmqbEkEVqpAUkFheltX
UBbxbhXa//RY/NUTRCEHM84Oan2uc8pgUZGo7+HkbMjwTsW8bQpuaIXbWnoizTme
e4t8ACuuTNYx3qAjmgJPyA==
`protect END_PROTECTED
