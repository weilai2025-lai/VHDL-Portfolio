`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6BWflx0nVBdANB3NjkdTeTeQ+qRYG6DL+9DfOwJtQZyvOFO0+aWMMIkBjZRmQXC
gnImeW56uPYxa8sXpLAmCzYNox8WbEjGB39+pgNfcwH0j6y6qnInRiMtt+0zW5An
jD+CAE3/uT+9/t1kYO+vvskaW5XfIXNPyRw+3Hn0XBSJrrvTf0wEDniau41pijZH
rbfbAQ/WvEbZ/lXdCL9+3sB04VLn0Bx8ChoiwEQQTGZqDnFElMmFqyuQzwA7Mpl3
gUrvkZOXZKeakdvzK2FwIsxGdr+PHfgZsIyH6BffQc+jUFuJHlXdNm1Tyy8CW67Z
SWvLqXra9QMjzzHAM9AX5agAw4oWrWMZmjY6zaj+9IrPEG1diSbC5dxPRPuaAqm7
fow7Pd9Ed3fzWzaZCaB9QpY5Hl0lyClBs1k4jKcDTQAyVIdFaLWgvFZgLDvTygIE
phUkhLhoDNx90pLRFyyxkHy0PV3XzyCVg0PhrZIDze+mK7kRiRCvG0a6wrv16jpH
KXZ7KoGaElkuuLuce7zwu0EoM8rNJwr1+D/pXCHlIq4mO4mgoQ5JD137IptL8DpE
tESaYvi1aylNzar55EuM1cAzBjA3gRTTK8sJRDY2Lnm5w7Cp3byRMveNLA3ul3Hl
4XlADHggVXcNjJVmHRyWfar0wbzpQ7A0tBaG7SDmqmy8BhfnIsjpf3Wx5KgJ3Llh
mlZuicF7IKWbZEaLkXQchXjmoSfjrZx40gjN6LGZOPbS5GBn7Jg7jdjUa/ZRGgEv
C/EYYjCyG5B6oJoBmry3GwbItKCQPta7TH6ZD3vWrTjg9pObHPnO4E2pGrOnyq74
5GRsDSiXVkMf4F7wZ/wujyPpJiFdpkNq7atfsEOWhnZjisHY5QVy1YDVKnQ01OnM
X6t1JrRmHjbRDk2Fc3B3B4aNqbCNC0FFgUye06in1torc7hUKwmFjSFU5Zw9EPs8
AEfkU1HEvpXNkWrMftTbzBSpP1AaGyd5dnp4Ebl7jwEvUbBgTUmOl+W4rzpqFHDZ
joaA8/CmE+maDJfIBvUg4bd2kJBdwl+lY9f2hn251WPLPc1qxd3iw2x64hvxMWIW
QDIBCne+O8cJgCFwVwgxVo+8iQhvTPt7yfq5EBFP7tea62gw+dsGf27mNB7mGKIJ
5o2CSIClIZquZz893rg3117y4Wld6uVoNl3sbiw8liFy1TaxARVHzkcnNcfpma8j
qhzSEeJM9R7Ig54Ie55Ss7sQtY2+OL281akIHF88CoaPx9V3l7gzCL3q1Oon7D8C
I3K/Kp0r4dW5wHyH7OAZdP1pJIEqxjND6TO5lPce2EvRTtJ3p5v7OmMA5bCwaeGw
y2D26tk3oZKy9T+VTkAsTSN85hWbKIl47+uFveNmv3txXQgeYSGb2yccsDu1EarW
/2c+LQMUW4vpL8nidzRks2y/UOszPvwamWETECWeASTGhmc1/VLzu/Cl3Ti41zQq
2JRX99TQd/p41zV2ZmnqFcFVaRQyRwZJNaFdavHiun+Fwx/zpDhA0qoFjblbCFtW
InA4SOwCTciJPOsIOKdybqOPMpmv7S0Llhjf8SVDiBf6CBXs9Nyu0W/kMQyCalZk
U79xoe0YXWJnoHI91q2HAKLazigr3EuuIceKj4hhZ6E=
`protect END_PROTECTED
