`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0RAKL2VPhGtv4Gpf6Sd1uTaC97aU3cB0qXRlI7CHG/zUm7nUHMz6QmbBENCx1qU
qEdB7CsSsliPka056WNS1dDnb/SI3EkMyrDX3DZ87QOfa7mX0K1Owls/hDM7FlEy
m8I+0fyjeLOhfToGsqyCwmH5heAQBtLvLY2K20ISCb4e9jD2qonyNOvi5XhcyOHT
JBT6DP6EI8NxpiYXnCXivLVkecx480X8sByBx57BFPwFaYBeFjKYyOG3izUenbPR
6Ef9IjmDcsDwzmWiQRBkqjVyvWNiYXD5V7/4KJZu3u9hDa2MeheGcXqBzXef2M6v
VMj3J5bklBMqnTwrt3Fea5GvXnm7pwccJ6hglnyPBczi5hFHJc3WIjAWLT82AzZI
FW8H3Y0EC027RlAHXEfb4t0f/AC1BvYLGsvEVyy266uc9ZP2s2jIskYg6U6CBpbB
zTC9o+QsEgRCBJyGMFvHLuW8o2q7LSuA0WGLXEHu6XZiosrIzYFBgFTTrXVWBQsP
3WtIGDt5BsSzytUaAaixK1w2gZ+YLY/ulQuNa/VFJyUIIrgQESJm1NtdC9DglKdz
qt83MonHCfUbD0y4isYDkxaX3TC2HjF1iAZskbr7wmAtW1MJwa7OsFpIlPZ2jgYU
FTPYkclLb46U7yRpGZi6sCSmBCP95ZCi9iyWv/GpQKTy1Gk3hx5JtAnPjP72+Jk1
e7QqIvArO2Binlh3TtxH7dOQSQRmWfklGKon1nzqKOE9C0RaIE7l5FqxxydrcJk4
e84cgrkeliBhPAMmLy/fnroVAzluQadwe4NGsGOTb5aNvG068+SuOxf1zG8MkPlb
6ccThY3H7Pag+1J4Ww3hXeKJ1D+4FDYz9YKhKLtSl94CHL4PBbkefAVwjJ46VfwE
xh/h7pmSl07RsuO2WbtVIAmZhZVg061XisnM4QZ7cKubcZzuzuKuUwxMzCbguR2E
AbzOJP/540/9pb+y2oIhvWFBqG9CBdpkj9q6sjS+bKJFKWhrh8ru2A0Iutmaa3g8
n1bEnp1Eb0oAPVr8AR51llH7rV4zaFcsYP8SNKmVoYdl2GiL4/7jZDTwO2jNH5Ep
3xFcqKys9v9cwv0z5M8R5K6K3o4AsHF8ygY06fhLIZRX1Pj7aZlUUvjulFyXs0Fb
6xwaHhvzijxLUYo2LC3SDIDWqCJxqBqIzcB4OkLBT1zYrN2gHHtYcd9HHPYyN3Ea
hd9fkiHysNJDSR8ewjPc+XFDORkbREq92Hk76Z1FaQTapbCchlmSXt5YpIrebOZJ
v+xzjD4rQimVIg8YWjOlyoYXs1ZxxO8ZQKaR24PMs3cWmk1cIAHMFnXCFY2irvIy
yNtxeHdZ7MQ38wNdyD9YtLcKA8GeWpXGH3AvXKnDVRCRvQ5Pebi4gTvDuLW9l2Yo
ekXvQC/ODsc+wKASon/r0c2N+C3AbfIpmfJJk/R1QcZcnsDzpt+WFfUIF3CeE8Gl
Qno1uasmvGv79JTcCg+/8FEqn6OtnQhS/SHOBufAW2qn14HcXzJVdzPIj8RjuUYM
fMJDYqu0wkx2l/kTO+Z0b73DwyvjXSQBJw2/P8++rgMLtgUgy05a3ss1Z5g5HPqr
bOjLRhcjKpkYCBYLA+UdZNsr2m+kekeuuYxH1f5ebry26nxyykZwpSfiPwUsS0Va
0s/Y3V6l1yPOB184V+eMBbUuc6c+V8PUHZ909zeBWdzCMO41ncWFHnVi4749QB4t
m1xpLaZo9/qHudOU243ctdM5vDXg/qY90nAiVnzVnlzkdmDWqi0ttSl0OgUYHN4z
hfB79oC8KZNXV+QrnX82KPih6Q8TZRFc9ynlC8lY501MQ4HMHGH6x9qVwjJPInQy
5Slk/UJk8ZPRCH0En+r2tWFJGVRHRrlYpzbz1ScqV636OnZIQZJuIH2GcJPM7qJD
Y6yttkiHPpNY1zQtCrUQTStLRencsAmLbNDgmosdzR4UxcyycxJFmpMKWSzsNUt1
Ff8pY+GSXvx1Hwp3SNFnd8WleCyRuaIxmaS8Xj3gfwhwcffGhlqPtGwm1s9vl4Yp
fTgg/1H7JAaaOqd9xU1E8hoRekGj+Q8YmevS6mJEMXqHomOCP11DjoFNU6XlZVz9
3wxmS4EkvtwDxKJcpwcLthVxBus/dLJBQY8/1zxs/t7vOqskER/JOs6PT/ryOSJn
2Els4z/K6fyrTYszJKM39JpcxwKaqUF5uA7Bm4sQUeBKWI2VSw0rMug0y8xNoy+b
CAMMwiYJqp+G5KVpw6Chy0l0+Bl1cZ7dCyaIONv7vFt46liVU76s7+2EXB3EQlJ5
HkQpoWyALsMLcYZRtBDm8+EWbmLL5XWWBSxaj/lX/jGrHGAFaWEiFyDzaK9d8Wsc
hLBFXFpksQ8jBm0PSEHVSj5jrZmjdc1JwNjJ9vLep4U8bOaH0P0EGb7Edv/rATZg
0J4+eWmlFMRNAe5Oy0wwKdaknGlsLGe/Ua7zIYfj6QAHqg7yZaSRQuud9b4IlQAn
HBQF9f1FKf05I1DJrtUAbIfF1y6NdG41OAWw99u4Rq4r0GEBIGCk2/+Bog9KYdUQ
K60Qc0yWO+pJhYUAeO7WR8uJZGvvOj/b3DbVokLDiF9ElO5NX0lu+fcyrAnVRe1j
wziXUR3Y6IBC5Li9VfQJXOjjsjr/T1GH4k4uQtzYi1WxOcPAAHoWnzoJE3qkI/QD
VhFVKW77qmgf/RMST2l2LONYR6yOhxQG8pwb23Ty3nP008b0WCpv8wRmYSR1+t3r
HxEz57QUwWuodzuKAGXazV6Rx+cfBXtpZw4/hWsWbedHFeRn3QsqT9pwAn70cs5i
XDcyphvyIprsvKQxiUwOruDw0L/2DrADPHILDB1/yNl9wAgM5+OgBRa6X6WGKFId
2/czP9uymtZM95XgspDM2w5uVZ8mGKff+ur1YwlBvbnzd7K/3fARmStLKEpDlrIe
w68rgzckdIFPC0n8bVwvX6pnxgdODZ32wq3izysMQI/zN4puZXNAhTIH9qGuYspJ
9u8FbhJjLTukS9GyqtRdEgy4p5ZWCj8up4Z1PoZqsyooTfreoDTl8gZWUS8P+bg8
eyYxEpMTysVFjoy+iqd9fwwKm/Pu1040P18lvi+51/WCFz++56bkOQjQihb0jXf2
YXadqUNihRpGY8lzJtKFvmdXghR7LQPyulpYtyMjGwgLIjSe6p4GQM7dxO/AfREA
VOd+m3blAvjjC5J4RywYZP1xDSl2+3W7s3eppJYVwzwQF/+67RLL66Loo4DCq5uG
xa1efa4xc5Z5z+bcKdTy2KYrOHlFXQ+AGcf399Z+Sl9B6BGdh6HbhFsxSjH5M0RG
S5fb3JfHU98UxTy95pftuNXNHSKYrC+si5pwuU/vKDyj0hi2i7S94uAyWHsZHhUv
XUGaNGdoFZkRF30jozSnQjbKEhl3ihc1GVvc/1GhV+ifkmKS6OotfJc6HUl/1dYZ
ZA01b7sMYvdgrLmafjVX7TjQmUPQbFDmLBdrUZwH2N8cLlMKfLDTVv0big0R/OSg
M2xBg0d8gglmbbyXbXtikFG3l0rHd/jnLryQ4vwNty6GEort2Cz1nE9s8zq8/jYe
mHO9cp/ErVq9SLyNAIYlzmTH4jgQ0T28/R6vQ88Q97v5Ikg9blR5fR6CUfjAWNQE
Ei9Fhm4embYpZ5fZlSPbmozYZRIOMFpFh3kNH0ooGt3fDSD5cQ72HCj1Q5BPT99b
wRIUdxBt+1vcT0SaMjL6JcwjEw3KJZpMOCkWeh9PzkwyLNrADUm/x3a0DTHG9Fxy
6aardMDGBv6XL5Lgy8KqIfstbLXXSGHZBIdlKrr3LToSzuOmkHPD4x/AaP2+LkqF
U+Mlicu5Nq2LZcb8VjAuKyMtnsJ1FBIXacRs6A4Hvce1YZZuwrGf95iARubSsubD
uANqcbqkZ4/wcpj+HE4tI4EA8VX1g/SS41O42s5IeARzoRZa8kfx1iMnYJdYp66W
WMwRV3806CAB1rAfOK7kybeqcP8YbRFV6DzHxFdOGM6+XF9lCAeqWZPFh+USvvRn
bjDj5Fw+tyNldBO9wI3PnC3aPdOCABzOkzLrFbFMs9Cn7O/29WGvDRBg5BfmL4r6
Dqe50gAnzEGZlZ7c1EhMgHIAzS4gR0oudrI12+tsdQ41rdmi+X2x7vNYsethRzD4
9fB8Jmk9/1lOi0R//4DeM4bjvQf69PKKpgCxIzv5VgoIT0dlYJiEefomiA6QQeSQ
+Y5d7R/SCiXlRscNlVATYK4Cw6nqfN4WCaMLs2xt9vjDofNeg1T87U7rCV5tCpaA
wIRwRmRnN9rUrFYQ53YwK66epg+Ub8BE6r7ZSXwLo6CbPYe+l6LJpSwLVdSsbfxP
dwslm3P+nd1Mdhg5/s5z0KN/b4D1IVO+SUatE+m9VAiBGfnPivhjHT0EEbl9lTMy
CAjBmTo9+Klsbqn6+6Kqfaf+An2ZlPSUzq848UlHuURICedFHVnXOAMEVrKl4S4F
uGgd4S5R5S0wGvjhFu4zpRj2sRlTsa8FpAjKfEZGkVD1/+yDXMnN+LSTCnMHDQTC
/tNzq0uo/XKm71sVEJwF5wglI8htwyAl7UV+rUQegF7qfQr14gU1/T5+l12RlGwQ
aedd4Rwo92Zhokntd9f6k6JmOwmVUB2a88WVrdLRBuZu1XAe8jhEoFKYoehE8V/y
EKg86BTgvaoFPZVE6Lbesq1TjKHSkBI/IUpBBSBj/hoehq+9wNgzv0eHTL3YLdFN
llx6kSZQzBWHQ2GAQ8h3bPEc/DAIPk0WdNZkrcSVdA/OwGqgbBL13FqVeLZOSDIU
dOgVPAukPgh2y+gsjqm6e5OTgpv5PclmSsFjuu/q+NHgZ6aU197zwgL8KhB+OP0R
hTf1eOsb5n9a8RMepCafvxJ/k4nq4GGxkC10f/RHPAFDSdKFsDvqzBbBpo5V352G
ySuslK8DmkZBzt7duGn7Y7az4W2eNjwzvREvweLrcMjFsenDwxnubgyOL1P2NJCd
d3ryAFxbiYHS9+h0GtbLD2F7OxWUPc2WsGzZDr9C8KyWfKXhvxgNQcpRQ2wv0P0v
CzavjywJsCMCTVRyUxXDXox5ZQ+4+kO6s8zsIbxE6CM6NGsNNde9A7aRdR2HpXge
C0COD8RMCXWy/b5J2lCP3UZazgQYziyoOHpFdTQp6T8DvT3mN6lqFctfI56KYz0z
m96Cvu8VQ9NOLWSP05p9xsvT/F88uyhzsl5n/diTUnT+lUDBFkdPAPUrTF7jpqlV
4b5I5jC23KVrNJnB1xjbyb9nU6wVsfsPomIHQQfquscE1NI3wGftiqz00oAAXr3A
Us+Y7s5z35IugdpdVkCrpw1kMOSrc+8U4M+eDSju8NBXQgKUvYGXbrUlgGs7hC5Z
30/787L3lYL/BUgqKFJpc1tRJd0aIeNljP+1mZQN9OGQy9SEdtvKhEiiO7Jpnt63
xLkoXrLxuOryxkKLUmZRJGv7iw1dTdGdMMqzJzzYB++8FttYi2rOC2YSx25M4Wie
A7tzYpQI4suj2Ie75XpIbsYVo+yZG/GeYGv/3ahuVW9WlqQGWWS+27W3h6qMV+wq
qrjMs/0ckrx33oCSeIFKBEVbou1DDvtp9/ZyPgu2owg6DahTngPC8Ks2ortnVRFH
tSI6dp2OR26EBEF8SDSa5kTPtYqU71pWZHweGC/N8biZ3YuNDGcdeTELVvxVquXl
P7Q6TTy28UcFtL0N+vyRXGR6Gsi0IRD9TcjkQ5YxplyZ4+sHAzzc+geybMs4YZG3
FMrO90HIdg6lp1cffyzq5uTW29lgXSHUMzkjRuiwa0JkQyHKMa2aH13BEiHfOeib
6OVs6ulxlk73w9LMEwyzVuW4KBW6MuDBExGN7eyl17HTSmmB9TUZXMBn3wXS7rii
FVnK/Q1AP1o4gj/wmGcukb4anrnaQXKotAKErncNIdgGn9KYR0sf1b2cSn3dFVZU
pkMCuDvhzNy33xbNzSk3Jax9mKAJ8C8lMxMScuPhGBuNNVLJ+I+ai85sK+bczyZB
LujRaUck+/1LSAPoHspEA/6PS/ei4I2rntQKBKp51Cgkw+UGQSLEyuR92fsxwAqd
u/BBTES/8GDx7PmONKivyoyFmZUrOy/Cb++3ARQZwsv3fWRSKiEE4bUHcTaXFB15
0IbGa9mTDLB2vQkbZBafj33Tu9x6yLFLwphacyqWUwcYVogKgmgmIY8bIg0FqzT/
LLgOVUcbC48J7hS0p5cCgw3gVsLWFSEBo7TQCRIZsACl6ho7oH7FM/1W7hJznuev
BqGBuq3NT2RiZdBuN8Lpj3CcWC9PKZTV2SSTVRjmimNCyvf/V4agUbz9E7gpSjXB
qs26hf2Ctr3f2e98/8TXtaPCe5yVBFk50Bh7pBavobPwZb5Ir/3rGuKRQaizyL5X
bKWfZYhJRicQR+SPJnnp7WuXsEDIbwvmiVsTzPMlx01EdOOdujKX6ILXbHYw33fB
rot/Np7DlNY81zYWaB9Qr6kTrFWrwOJX9HRVXn1gfmCCXXMTdwvvmEgP/H3sl1rJ
leQkQWhu9wx/vNkpfHJAmluHRZc6wMPN9wscT0kU1Q0Uuh2tcB/vyzP5xTM7LCKI
PdY5o4gxLGFVjWT8sOJxPnGIDNHE86u4aZg6HOTS5279ngmY9AgI+hdx7TMqsWxu
tcsH2mnV/9Ow0WU/3bVVtRCTIIXEPK2dKuPU5FgiHfjJZyf06PcDle9jqRxeNVoG
EOar3YpIRkj8kSn9Om63UJLaRbkZPYsM0BkKkt3qrfi8h40hJeRL1lMPjYyHbtnz
ofDdVq7cVLjjD3YgFjU/nKnkS65g/EaCXXwsckQZJRpDf+4w9F+83FhT8I/Sh2ve
soIt8aUop4BfBFfMMMqnEcbFA0CQ5NzFYrxYsltVD03WIkwZ2s25dAtdEjjZtQ1S
wc+DoWHWOP+UhLx2YHYTK+hv8YBzHuGOUpSVQg/csqKwFHuCB2ts85j4qjSOU2C1
xKqGNWJWL81jhOWyulGz2ReHWpIFZplsJwgW83ipf+NDJf4xE7RmzibQB283xuCw
NU15qzJ5GeHv+DF6oDt+VCHvDMC8G6eWpaKEOF6gQAM/Hg6K10+8HMt0xUFO5tOb
sQudovYQDVkLRMFoxxyuyoIRMPgmdKIUphL5FA2iRFjrdQ8Be4Oc2joicx8VapsL
d4uXIDR5NFejVflbyTMracafapqXAVR1LgBlUMiQ35hzdIbyXtpkFjPhprzv6oWG
22VsJqUzrjpmEcoQVRloKp0SPdOKY2cXVthvg53BPyS4AvcFz9g+P+NOlVpCn9eE
WizOTwmdOCRXNCBaPmuR5Ybg9iQp1NPTX++FY4NvC1C9lNiUxhFqgxras0sP2a3B
QS4iFwfzCJXzHu+WpdmxvL/BQYhjdrWSJw6v577t4bTQAttweZlNB6qVVGZDCy93
nHoXSgw9CrNu3nPfTjm9VH3vN9f2U3tCORY+9SVIYP0xk1d/rtiytqwooqkRF/TB
njxaeR+qVr3/pjb+a4crjqDLqAOmGJSdnzXCthhlTTdhZ+jHSW3mRL/XLbKMtyff
ODJQ7VprCO6H9vYxYL7DnJzgXxw6+i0C5UBvvlWg9/vEl0ak+fexcLKtu+f3MpGw
dQH522lxEbnhZ8YNuCT+FftRL7vNeEs/Rb4/7ajAVP7NDrqLFmiavp0HT9pCFAF0
TrpuV7lwV16rVx3URYVXiOsq5Z0FAfiGUhy9quIf71RHdRudi5wxDpH2LShc1w9G
mPQPOlIJYhWFvbIraprT0h15c5s45Imd2TMyIRH5QEnrbEqaQu7Wk2g+QC53ZE1w
kcO7TtbWZ3sD1L58tgZIdUgjvkKAmK2akoeOVE+485x50K/OsIy9WJfvuwsyN/lK
GFYh6q4hLz++p6o4r26I+E1dRAkDpEBxPU2S/N/7uKRymNyXAZY6cJiklhUpaUzS
U8WZz2Cc5SlsRCpmJ+IOy5bM1eHGB25I0m4ZeVMkFmvEtnw5luuUKSIk/hJsJztL
VUjXtujPR6RD7ZsfAHHBFPKjceo0ERhUDZqoEZKpiO2sIc9tRB2L8tukZUnrV7PO
MmZzxbb+BDL/ygs50SG5tqohvzZb8n+SsT82JEtQG3pqXbOIG7uUYcOU2imBOohf
pp8A8ruKc9BWrdTnE4+DpSaA1PVL3FX+wtIW9jt7UhYc0WUR23+xeVUw4cL7kq+A
h8KVpAM5DAAqc85uKfDHivTo/SA8YIyrf6lXRyiliAXrfoPP1/9JPyjsYR4Ewj6T
2RDlzGhaigf1pnnrGXPAbp9ryvTJIaaFuu2lXB2ofwiiVqZasDQnKEccIz4RwAlL
aTu7Y9gY/j6g6f0jUUseNNmH9MuDZ55NQ+k7ynS8g7pHeYUL55p0qX8oOQBtNG7+
HQNp333EdEMMDpyqZ1ZIJq5Ts2Iomrh/LqS72IoaViP729pU3MUku+eXAE21hIVu
ccQiJx+e1lyKlEzxcz36qxWyHMJGG196hjLcTvqZ7eSdIq4+KYH4zqv2v0GrSFH8
GLbAwGuXulv0hAv1Un80ZA6ZgFXRBhMcjoPchmHpbmeWwzlxstM9LEOMEKtM2muz
mbOOnHbYv/dYPvq6j2dJSeGGwLykb0iDXGzXphopzgI3oFAoBJMgzO6I7q6vYrII
xnRSG/W8Y+AX0Pv42fY8EAm9px9cz5Z8SLsiBQorXz7DBQaMFXKQ8SEuBRB9dOxw
kvoleIO/DcQhfOS4hQa9Sl+OJX1fyJ5b6DE7A2m2IuMBMbHx/HH8LKM68mLk+BpJ
bYRN/7korAQIANXBqB2Eo/qnhYZtmZcjr5QlijDX0SvphBp81/CoH6mS2nrHJGjz
6xEqVwaaS3fdC7HiH0JDdvrr86ouFGXdKjhqiFw0UbC22cgmoveXZnKqPYjC/Wsm
q/69NNnnv9uFEFYPnBDbA/X4TMQWVedGU0GO5i8hlSyFPX0RJBzieDlRP1kulMJ+
II2Mmv3PqWvyudY2jcNEtYX3SZl+5UZ7gK6p88LEutOk3UszN8poNUQBYNKUo2T5
6i17NfpRphcEvHBPA9AK8wQA+2EuDOhN3Z0K7S6Z9LG5uiRycTOd6SKrcwUPrh38
r85cVAWbH1QtMS73fX1F3UvZmGYNrXilHAIDGspRfop2pxJoiJ4W83UwKp0nrB1O
XXk0LOK9KLgOgZMNU5IOYht98MvP5G2AjVUTQNBGcjwyf4R9vQzB8m3X0WaNhRpT
8SOxExcs7CTdDhUUDk8tcm2IZccYgc3m/G9Rf0o6qt1n8h/ik1cu2Q/nqLl7yFNY
ST97d9AcgbIt4cAdY8dzQBF7miB6QW/B42plgmZl6SmN9d8xclTS5Ir4QpHJDbHk
sy3PPtSUhMrP+gUGckJrwz0KlpgWk20xZ5RXOod6j7R6DnZaAMvoThDaCBE83aM3
jsR4OP2hn8DvdTlM13zX0r1eNBu0DpuWnpfCrMYFdgXjPbG7dZ3z7GxA1czy6XpQ
XyWrZiaj6NcAMmacrM1eeTk8q5TvBiuEGKMpSpfDuPi729EikTOpJbAtMEpUWdMC
TJslqLCi9D+l4HDhc0l56WnUmJcRwf/jLmjh97TO7XZpM7ngmzzjpUvgWQUh0K9R
h5KcV90aTJ0McJ3PCP8TgxpxeKJmmwNf1TwU5ljZw4WH/FgdSb2+plA8Wz2GTvrI
MQr70QwLamyiMjQQPXk/tQuYmL2KgoMV/w4Wrc4lFtkb6KXkT6n5VKrYwrNH9auw
9MwWD2SIQJcFX9AXvxrXVFFIxr6idqP2gOhsy8RU4FFubzzzhu8F8WkiZ6o/mubw
s92c2MnJAimiE6LUbTatWZadVZy9V3dnwtVEzs2VVREqUQC9AjskSLRSiYEjNa8n
x0P7DQMcJNXEQsusgKSZB/2YuSuRoYHVQOl0eS5AUGDENJn6mIQKyGgP2tW5pBYz
8wxKVU/XtPYr8hDAKSRK/oudp10aAUtpPmAYcfZM7wvVJzGpAJbHB4Sd7ACT4yr9
EhnfZJHye85r0sGb9YHXPHaeXlVKLX0GYblgnhdS47ORdNmXqoQXRmyI60qPdmF1
yc0TeLyovb07YFe2CAQpZ1WSwlR3B1XKf8tlrVWZu6wPKKeM4+QFGdkSM3wnoAdu
0KmEMnnmryhoY5Yu1fdIadwATN5fets16a1h4MkMuw30wM/LrkTD/Uns3VKO/ttk
dZhZdDjurk4rg9amNjM+Ce5Y40dmFwSBZxWt1HkzirpfmuVRLys8K7mVUOloErQo
RldEsR3/fETmsoB9/21CVdMjK1XtITEOTysLsApd319/YSjdJflaztDc+Nx7Dd+d
MmU7mntnnjwqagloraJKVjpYegAPr7JyXsKTpRoRWGPYPla61Tt9B4YvKqh+V8pJ
Z5gkeCc+eYfnI37+JGGmlII/QRv8wUE4kMl+DArtXx+F+HleTav6oxbGeePZmdQp
AlOeomdHU5oKg12w1B9gXC9Lu1lqII8JNL6fm9G2TZ9UMm2OaphA5MvJUUpTlHwc
0CrA7D28FWFHm1ZKmxL/uJ1KsPqyVzD/ABXsKzuwzQ8zzpWa7Y945k4N+niVqUpw
tOYo/wZtbX7VZcw1bbJZbZBBqkWDs0UUecw4S3FkoF5QJn2ilKBvRCCOR2HfBexh
EmeRJTrgN2yWPsyLIBvcXatlGY35tNkzl/jomYcaHUTjB1vbvceec6ZbSZN4cAVU
QjAqDDQ38BFpfwaTwa2ZQ+M3JyowkrGAP8L1ZHpoIRIAlXCVWqmbUDje+RYc1r6A
qKEGGMREvAroSO3ijiAH98fQScYDkyV3gOc3BUUubCvzHXfJVHcVywZUQ4SmSB6P
6c3XcWI/3fFHvxrioiCTyx0xTQbC9qGBb7igozAp1JzFx9BIwvL7x3KcmtAqLNzR
FF6lXTKHTxalKggrvXODo4UxVQSaxMJkj6cVb9zuYNBxCHwptIZ3eK+gmZT1YjY8
BgMQWZXH5VlACXP/S+Wptv1kzCzQeL3BvoIKHUbaNJ03KNpKrTWVgiRtsrcBytWI
8d3LgipW9UOKEefWg5HFHGxFZUZPKqxmBXcGQysXArXgyQXNH0qnTESWWYOVZw+x
bB81GJnogai3NW88o5jy9yRfiohRnj6fWgz4U569i2i2sZbpsdRzZD0BsAjvSnuj
87OBE4V+ET+qbAgQLz7NTwRUyc9ErUQcMdz2Uts9/tcVJ/dFDaWvkO2BGgdZrKtk
RfCFSbCpckJJCH+VpDUnCTZGzQ6j+Oa7q5WCgBXVmwDJxFr8mvWrCh9xHDB0il/L
rJzhHNRSuurM8VAst5VtuHtlgm+W46xq6ky+7y1+DZUN+W41rY8g7T3Y/gEkFHXz
Hiese4KtU0l92JfnG1SEHMmonFiyZbXzw3EDeqkYAify0BMoQ0gNZ9C2MS53/74j
AFIhyMwfGBUkP44unsae3zGTF4Ltap58MBI02FPtaZegtNNJSKlJ1BMSjDm4wcyw
6idVzt4Dy5uznk+8I4H3+t+aD3OTp63HtrTSLob/yKP6HDXyMRyaDBmFo0Ahej/i
xBLDNZc/pVKGivNgM+QWJ8l1y91nWHD3kZSKcueQQNxhy8PCJz2GVfEbKFjqrJb5
VQ1hNdejNf5vAcQ3/9jGuKxpnwQTcmqGXz7y+fSKcCoKfbgYNv5pMi9h/AOe6Gyq
6jQf7XPKWDjwwsy1VLJZPTD5qfl6lf/MKpKLjY/Nk5WXzDBOPOlTQRjMJ6VhBxp1
q8OETTEAU8zYLM6nEQfOjOWqu8muCG+YlwROvfREnkOS8po2PSMcK3WPEE4V8q30
FaPnIQGIxDc44INDFYtiwM7K3dIOJNRBYmaxnCyBV1wwgc/2F4DonBNcmg8IpU3R
xYbJ/JLwAgi4FDsjeVv+2+Qr0zAIEivoag3CoV8c2BL/gw4lgp9z9r2yn/HKuLHc
VT6VUHgAM/42EkXT4PLJjspl3VWp/Zc7jlxsGBsBIg/g3nxcdWY0MGHTLwSXenuZ
UuxlOMuKY3LkZDO7BqFNOQRIa87SOSnqNNrymn5Ibr1YTCEsWwD2EzauCUXF5KD1
8VC6F/mL8ykjI/ZL8GGFGo1tkPVYZVFUfBcUqvOkQ8t016oVWEYVe14k+qg/fl50
JplXLPAiLRqU4yMOjHy0SHNoxsSMM+H+KgjcYVqSgSxGnJVjEwsWrOoeK7R3uejy
ZPdLbcYjQNCtz2z0yLMZTA/y1kiZzbzxoODLj48P4Wr3MQUKUqRXGl0TS1ymMM9Y
3TXt7bEQNaxwvxaYqAr6KUnqlw3K0lbDbOf4dY2/4UHoUnDwv0VXlLgCSP2iTp4v
Spiuf2AwYecuF97zIGF5Err++N69TLPCTgeugZm2oiHzrvsIbXUReGbhLh3/8015
K8ARfY7jAI3P37z2R7H+ehBCoIYUPhJQAzvJFLyo58f5M6bBAwSI3cBbcz7ZT91e
KlGTbZmmevNIrbwBAHP20OFkgcg3KjguEYlwnBOY7xeERu8Mcp/uF1xplhFzsk88
wn9So4WwqSWzE65u1FpDlPe9pV3XqPep6cXijquBhzzuclKjnJ8wuq2kvwLumOTO
4qWePunOv31lFJQ2Sy+1bDUtIz33ERcFeM08Rf4P5c/QdYsAZgok9a1Iw2s8yHH0
7XppANaS+BKypbJqlxNP2uk0FyFMT75GdhyprQEoyPgKI3gh4BXlHbEUDEKlW45j
zdj4uuyUfGHkADgj5aQa6Co0kjUSrXH3P/MENkI69TEn1/IBC2t2o7zAfCo5T+oA
BJMKcnAvaABN9vtsjhgJr2SrySlc+8ntdJJszxibrXDtbcnG8Xojv3n1xxtL2Yhp
Hy0via3PPtb7+urV1HsDDS+05YQkfPWOAlh/2HuLxkRaj8yorcjZtsdHLqavPJz4
cadPoii5svB+ObI3gCBtkBhoUbJptEcJaVUAMIA7GrGh81/fxoh4gC4IvZ3IYT50
XRAVO07uB2DfkRctADnKvTQ9b5x3wG+eFRBJtcKGNK/uAzC3mWWdCTamR9+jgfyB
WVsOI4a8smCJX9PnnGoFLyiCUB1GnJHNJ+0VdK7H9FYSixarY38dhlOX+5Qx1jhq
7fr5RCAYkuG2yK0W8b2u2KGoxztVyEXNoJauxw6/WkvDRPoniP4a88gRDymIecEB
ARYttH3E4huFrrhHA5UCiKH07fSvjyafOgp8pu4QsBQRFcdB8bWccmk/pubmIv0U
67F8hY2zOSe6TD8QBT99tbobTLodcjTBJ6vTi+BY/UbZ84CQqw/pUIF36M2uhdhg
Adew3JcE7xdo0F9nCZX8F2sGqLT9ZJemQYxoJMOzs8E6Fy/NZTxVPlGg21OiX0oe
hqjAZnt2X7zgL9wHkhLF39H+PXcpkPWuy9LO88IFMdpfnMasnYfxxOcX2FHGrfl8
Iw+dFAfwU6QWhSA6ymNmCHJIvLznKCcnqQNJO+dSprdLdfvTJ5SkklWP72kxQH3Z
VphYH7QbXvdgQZRyOabutCbMlRPLeTXr/7vrOKuVH6cEyAOg3mRG86sbKH19sH5u
92FFcKc8GoHRxCMvrDiYJXz+b6h3vtMod48/GPoUW82CBtIJgLLOwBOQ1CuTvkru
JtOROeyrX/OQ+raaq/ZepViUG6HHE+8RCc5eBX4BxJ9KVz6fDU5wyRzxJlpFNiM+
V05dhvd4fARQvs2CROdsPBmJ++dPJtrFUwgXW0cfJrxKeNMpLGPIsWsKgWsPiGTy
FL2sHDBoVTegkqdcJbdz0EokvvHBKQJmn/4LatfVnDwC4JCjyrUmV6yUsNLnPBC6
RmT/l4HjTKHBYjHIxOUM4hiyFEs0IlT1udLEkOn5XPB9F+KuQRkRz+6sXmHv549o
9a53zYQxalxaCxbugWIBsmCbF3t7S7L3qemtHpHGLzcxAjiVGRfr4h72JvRRzk3/
ZFgQ9xw00QVW7Y7LyNkLWflA0hWgu9K2Jj2WstuNFi0baBiAPzZ2J1yGOyjP58AM
n3/Nz3FB0JBg9ykIFc/afulUaVZQrSsTNYc/DtLFUlZ6wmp4/paZ5EKwkFDB+p6A
0Yqos+aXwSCkjeodL+SxmX1WEZ0MSDxdFpupJ0RNujVzQVyclfb6EeSBMZeJLFUk
Xhl88G+HxfgSAxyn+EbxO9cvqz6ranaKCvwwTO3GLm0BDp/zLcmfYI++o8PkI0Bd
zb64j5ZudirG66LifG/ZbxBW6LW49r6QGCm1CvqMkog9qUL1G37ANEIog9tL/4Yk
uHqvfCVUDT7PRupoO8g56ZaP2IBOBMFiGVhkLB4LT7NGjH52wo/Nv6e7m37Iuk+/
`protect END_PROTECTED
