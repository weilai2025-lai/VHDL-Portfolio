`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPvRncuQFzPRL2Yo418YjXeB9ex2+gUJyPVDZxf9Mh+IoUb1bz6Kv+7mgbWgdIcH
7dz/ESrqs4KtivgdbhmlaKU+PxbjSuDmQ6D58FjZyfgrEyBOTebgkUYBMyD92c8O
N/8lcaJRCsoZSJFCi0rNUxU0Z5VrxX/GOufa3gSJAaGon8SHKnwDM6hPDYSR2rav
7v55JuzgxKFVhhQ5Uf+TWawzk+w9mP0FFf3XedhNMy8XwWAnv1ay5lRm/X07UW+2
ds95/qlFhBgFHIIsG9FgjUr81c+2PJv5XCj/IaxAZJynpkXWv+Ye69s/1vHU4KO8
3MoqHHVvx4C0IKWKzhjLDvRMZTeJh87tdnVsmhwurkD+6nkIfvmrGwzYDiIN8EgL
Z3d3vQRVVtYbDx1r/mD1+F2bggFWmPp0hdiY3gpRscay5Y9BuRb0WwescfCDtUIQ
7sRJgO33GC0W2RYPevigvtP/EpVM/FwMkgFcNQT9/1sOCDeAOrP1kHz1ZSupOVKz
IWkLixR/rLa98iwtf2fp1Azglbd03qQzz/dPa1g40RgS6gyVHpDCgerTIR6BtmAk
sG7E6B0vhcOuhw5tkgo2RLKnEzfgBd4wok+F9lBUzRMwUKJYET5jvr/Fdx1QkOFs
GS1TDF1AhqRoMi8amu5/u94HYcrXOCdaV5uS2GqMNMc7Z1zg+YIWFoKaeP1PEc5z
quxP3axIw7fyWC2T7znuL8gDGB7x7tGjDiSMEPQpTLDQrf4CdhoR04WMwGjzSiRU
GtftDUqYoZysssJ3mY+rR4WchQEL4skMio6VwKGCF9DappIOaH4iu0gYZEaOYO6l
E8aB+VJfSGVinpsXOgLe40o70Vbx3TLFqgxPV6p+CvvX7o13QWbUs/ZIPoTAJDJ+
miywVUFWKuDxWQ1NeMmeEH36TCtqQY3CCH1ryR/zi0Hlf5vMEuwnHvcV97uwp8aX
yGbCLDW465PMFJ5nFU13OpKqKpgs4ygjCyr3jxsKG+XJkjM3/y5M1Yw0Dw9li4pV
kCxLINXT9Ky2LCXHMPwcjZuiSco7MPDjD8XlORbbayz112Zsjsf0lYYvjPvvuioN
X+hfVDhlUn81QYjlXr/xDh3TDAbGyZcrcdgWu43EVsbe00yGYJo7mYZ8wpl4T53X
Sgf0ExtGgxUqCl3Qm8tGncsA+vXfH7JK1ZHRMh2pruZfLnA7jCPKqRsNyiHhDJKf
DzNQAUBnxGxzPXMZovo/TYWZPB892moqhNjEmHc/9u8aqwKjGTejfUhgAfrN49hR
kPxR1LRyYRD/rPGiBotzSXv0SmpxTHlxSY8X2ysaaRfH0nPEvlw6bzbgDXnddM/8
wcMhZcKdM5Sgkebpf5LsUWB8vC8mUNhrGwlLhCTs3wrJ3CEcOBlfifRiSvI7dcI6
ll1eGkcvs/0nIVb3LwaurC5CiA2B8m/K9utDX2A5P0CHMRarRtdlpec11POr3pCF
t6xMydozb12z84A/GCqKMibr/yORbEUeeyZz3Pq4oeF7L/ZkLH3aFQTjao+T1zpl
6V2vdXJu3sgcJb0/UaCTlTZrZy11jPDWxKff0GWra6oW6fe9x0PUAxrGcQomKmX1
OClwQoisWHD4/rboQAJKZOC4Zrx+XSORCLlMgJAsRhWwuTWLPXwbKBMBYFJqOejS
QguERT202zdrrVeNtBKcUDGXfKg53o4qK6azvki7dBzYQw98V9KSylFdakAXymJe
YSozgOK9XyVlwix4LXCpO3MHQoWZ6OF+7ycAPRl77NbMjQ9sX1W6c5tQy5vq0oh0
XheEE4t+4L9sAxH8+QI2L/chvtD9E+Y0BfvFAgvG+p/YCXeZcI5qQadULQ2QN92I
l4jkgmfj0gV3j+jZ1cZ0PhkCBTmXZqZU/BIWod/0VzgmtbcbcImJhTGQ5WwwFJbC
CGdSFJYK2iBIQf00yJn+5JoQ/XzuCD1iYGzkXFavcXkQkYEYLvkjevW0Ux7VohvB
IYDKkD85SWGRqKXjxfZJu+LZRE6O88sSAN66Jmi5DDWP4P+nV46CmDIwTrBKgCul
yF4mT9KCASfFIeYvzbViAuMPImgVzSd4vpIlZlsjGheWQAS4GY+6vhYZTZIDNAiU
AwCDNVCg9MrsBDs/qeSUaHsPQlthxotpGoZvpzxCNuO70vPaJe4iLyr7W9SZLFwV
saCUuBtTE9syya59DjTJmrE6DQty9wOmQ7ZWGTnIsYkN9TyZJe++EuNQdsGJQhGt
RmUUoXfbF/033gfsjsfg8gcWzYfYowppJfrE3RSEssCUR71DvYANiK8VXhhE5TYk
zDNgE6vbTC77CDmu2jGMElt2DAJaTAt8B/spWomaVTuUr7vyHx+UDR/egh3MboUv
EGwooGq1LlAilCm3w5u7h5uTk80OEDfp+a0XIFSo589EhuFrjln6di60V5rwjVlu
8rjGqWbRFqxGqmri3WALIlNa3Fv87GfmCpL5sZjVDs7ieJNtcYpd25ajuqDRPVse
T7GJg2zOSwHbrypTBAKq3icwwV7uZ9QS5zQ+oczXph047lqOX0KpSk55mykLOibJ
JHhvsdc5opuMHvC122AGZUMDpi6ocp8pwY5aXMJn1ufufvksMXP6Ek47np3kaMQi
ffqfM3YiX9cx1XUe+clNXZnrHiYcLCkru5phM0rhkyXbiifbjaJPuHQoOJB+ULh5
e7zUw9/xMqG7AGH58pLW7VoDLEwZnS0xGRTrK15CTbaQ6d9AMMhzwID5itMrbrMk
oPYLnS/gFra7xAFCZqYKwgqFyHqk65DshwGjbEOJiodBm9mDRAoY3NUlb/HQ4XXO
PELFGQlKxxTJlUqcCKisoE1cGuHq8KmFsTJ2n/GSTvDAfolPu+d5n4r1rdaghfD4
Ug7Lk4de5t1z2nM7n2YkPbL9k8GQHLx1WehF6PaCX/+Ife6WjZzJZvdlL4HXVDhh
Xj6DJ7FPtDSGEWeBbYREe98ZmXbyPhLaCXTiiAoO+C0jggXlpRx9aUij4OPjoHfX
+K00kx82zLHQcDQlvdeJ39XzCDr+h0JbrEsh4YDWgNNwQIp5UMs7nORsD4zV8gYA
fNknetymvHdLYWD+IDANHGVYnWA50DUOzBN2w7+dHhIt6x8AQgBoFnYBwA6jMCqz
Ulndw30E4qXRioo7LOe8+NsVlU/dVLWmFMdW0UnwTwlZanoxUZ6ZzbqmhxJ2SXsC
iWGuvmZpx/mZ6OOMolAdTZsot1/aFOz3wUMmOsj7BrciQbhg2zhKab+wCrCBZQ3Q
7kGkeCYiPf1vsNI8MnH/uFth5RFRLfoWjocsmCegueqsGnrdB3JMtjuH4dinCCtY
F9EKo7RqmySB7czAe0EJFJWZBtu1G4naCpHFkK4SaB8E3A+HsNTfVFawAfaj2U4Z
aBa6bBL4k0VfMHUdvr+i4lFYjmeHs2JPXIFdBDY+Q+1qAfMz4hF5CtSc0uuRaWDy
v9q5c7KovlhF54DKCJKsIG6wOSpt3mXTBXRisRmM6Mndm9VhtGeZqhLyXxHe3tok
oke2rFsfZResjWYCwq49u54QAueL4MA97A/hL0CLhv+9wtoE4rMO6m7A+ASU4ZdM
0gMbyoS8kbXIfk1KiT+ZQaMc2vGTm3sETC6wL27wPB2tasiSaswjLN1j0i7G5pdG
cLQYO6xvQdIzdci8x+4F2YqBft9OpQzNPl5BqexLGIynuTgGFJpv+MnJPH/nyMlJ
+tHIjln4IZho2/4DH7gg4aq7IcXVctqCLMJ6OJSsGhlxs1QpqXP5u/hN7parL8KR
tbuvJQL1KRItNuwBDeWdML1/4g8AYDxrHiHSVN5HirKT+5SrkL/yZ7WrvQqzy2Lm
wE5qstUTxOKr9Xr4XMwlEA==
`protect END_PROTECTED
