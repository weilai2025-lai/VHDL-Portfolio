`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0kpqpwygMfgsAka6P1H1kzzdvB+b6XFWM3ZFbBHBc2e+XII7FbpuFp0QcrLCK1A
su4Az0WoiWlrpLzvoSrv+9zoKSGGIA/QiT6ezh8+He0GZjnYaDm+mAB60UhvBAL4
1SGSUOC0raV4PN4xuUSwdCgPVGkNzKXDu7ghVuokO4gqOb0f09+3KBQnZQfzwDNw
PmDBPlcypw+sHsYoJThRzg79MyqXSJPLkmYv0ZjY5Y55pvhdxw3A3VmkXXvTOTfV
W1Yd0JE+HzpDg+XWFlAyaCjTBuomPAmgvDxaAATmKkQcaN8aoj71z5Hw1eWZmAiB
jak6JJ58ZpGDn7sfYF5/qMwLJ1DzedEd/0IPVeioBEmG8bZOZbFu1R5wzASWRGX5
96Lh3WvXPmDFs8dCKWjHQsobFPjElYIbOOVHG41C91/VW0AUHtKGzMVxgDka9pni
m1Q4qafs/baoU2ILxE4LgkjUE/F0SIhxG2uetCUy2XXr26IUv1oKyPwXNxfSVD73
Wr1T8/NP6vLjkip7zjj6cqWzhr7x1cJc3mi4APdQKaKEy1w2XKTDJhWbZswPXKXm
hsXPpYHqFljnFUlHgM4/6yfWp6PovsuCCBwVGhbJFcJM+yjcwOwxHIQAOMffMVE5
aaI+pKvP7Qi+VJ4x59KWiraE/mLOESgF9d3iHGR6nL6bCm9jfNYKGI0Gvsy6i1pH
B2EVb9xJy7TJW5Fllh1ZJi/0Yss6wzwDAluD+u9hT0eg4Hv0oq5TOjoRpx19zshe
OPFCDlb8EBkieCc/0wBE+h2YmcF8oX/w6ZbZZrYIyP4R0sedSC8AjGt1stvxVPbK
uKwuMkNkiaDPT1BUJnUywvCqLrPPbJQ6JyVsX3hbl2rrRvlPUW3buTqE8KjjH30r
BgkALB4I+ipL/bdtD1RSbPykqUEgKG10/93oop8CRD/cwUA8PiqcaAykmfBj3F7N
RfMeEPXzvCaSm5wXqD3mvSn2csKwyAoHlRqhzYra3CUnyzEGSsZ9Qn2CqdS0/WFX
gII7HYoz3TllUfbhpBKvI2lr+1YmD4RvpXhy85Yqcazmzh0LfWlnoriQEtkmK6q6
IMDgVPniFJl+g4GlzoCy4qSDd46pU7kcSIyjaAavNDlUshkWH1Mc6/QJjQwBI8jI
nWiLri5r2tlikBd5kQt+VzQXtRB0sMxVY7DJlotLVUIjN7rh72zUXB0Q7VfEFySt
74Y03sw6NYDsUOjI6/oHwxbr4eh4MqwqRoSzgSVxBu2oVA6mtPyoKFg2oKy5Ry7+
JZkFY02UFzDkuSqrGPpuuaz5hz8lzcJvF7bchijfFX4zEUpxYvk08irNb+5hk77i
N4KERm3QPp1AqmIGI/S+N1s9ZHrObQ1gk0yj6vP4XdkCjCnzsXyudsBOaTPE3iUC
9MyKN2KBb65fXdmIx6ulg5bwombLN+JYkO9AcXTzdkx7wV2nJcswkHRy2LMaN3Cy
50D4ob2KhhFAjnNMFk/nSmfpY6er5tX57RJaYJXY5/2pdRqlhvNghJHzOVTNwwN2
t5BYopdNwHaYZIDnNb4qn43osrxI+uj1DVK8u2J9B2zHqkLFQguUmXkslK7sl5Wi
`protect END_PROTECTED
