`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mQVEA4rw8oxlmUt4mtRRTUbSITSvmN21qQJ7790/2xXFZQiZZtHaRmMlPH0vh78w
LJ0jusgc/oLdZ5vZbzKLF2VmweP1OI3EO4GNqFBnS7ij41+Rba5a+/NB4nLl6I+c
6FCOhsqamLqYg2fv82/ZdBEA6tjEjHXMygGB6sEkYucDmJubTBS5Gtg//ka0M+qO
BXGlbFZbFZGSMpez9zsYocVq5iHZ0kxUr6JXx6idSBpJSTEpXd3S8SUWry3DwP8s
8m8y4hqoRAG9Khrib3CUI2KX4hDDLjKEvF5EHA/5xpgQmIld7BXDx3ZgPQ8gRYfA
lTrt9D/dvpx8hPsCtBGf92via57N5SQ/EJMud4eLB2k+683gBcvUCSGmmIxMabk6
nAo6ZygSLRuRKI+cy6ezhDp80+FTMug3542Rq3+8+GItcweAGb5Kr57CMqScLKD0
ckLhQ7w3UQw9TK/iCcHXaur/rBC15w1JQlj6OrodEhE+VDJFnFEbyqVlUv++CfGt
WpeFZNSUXPZHkM+23HhONSdlwhOq+8u1+h88PLmIWOK4b/Umstxq602Dvr/8Yn0o
fYcXU6lycBEagwnAay9hD6RjhWlb242m0tEUgq5BiSeJe04Jk4qhPWoWNzpEJka+
Qs1ujwGRmpFwaCgBLWSEHd1bkqqW/bhxiHRhZaq8a8Mvd0p0/X497Jw6e9RF86f7
/60zhL3jabusQP3aYY5tQA/zgDs0pSdA8zvd8ndcYvwnh/kmi+r9QCacbGf5L3+X
luDvA7/jYz6+1QuVve80lKnWlF1+egqEzhSj+4Vv4V6jxAcI5YWELGi6DfN8jZ6P
S/ebGAlbXq9baLg1VqwcanU3UT9G1rJQm0kUkJeLwl1TPB8z/bBc7mm0rjIKYG+O
NObgDv5yAR1DiiyFRumTbavJzp7WBAvE52N/kbOv2AVlFQ3AI5ziIQA3/lrjweky
4pHrBm1tIdmLS68bJih+0Yjg5GX3GekfRjF3Qm0DPr0DvR0SOxGwBmvIzo9zugfT
KpmxZFaPFuHOOgoGZYvic/p6sP1odPUnjSLj1ZP27vu/a9kPgk9nX4RiOcowoS3r
gshRuf3J1T8MQgSvtK+4rfpgFJHo/SvDWkO+mXmz9f6uE8NNrnJBPyhbDBmheXf5
mSWfD5+nK2HBggNpBRC2WCX+/Q+NPjUVcZ6/Rml40UwLPZ1XqMKKMAVkFgslQ3jX
UNVK2zNYYQylN9E00OCOTkwmcvVJ5y+EPLGWFrJZYNrpMb61e2HbeJc7vAWZPTRz
NI3vNEWM8Zv4rQyzM571sVF4cG3V4B/oLRu45C3mZDf7EVm4ikhhb2KSLitffq4u
3f2sUmkQqNOLe6/+51PcfLJpP9U0JMsWbfhcOAnkCuRrGvMSGN46EeGiKVIyQiy8
fykuslg0TXknXo7uqcw5B1SHjrsmTT+c4nNG/+sWuJl5INTevA/XU2yuNyYRx04b
R2qoxW5cCOep+21ssTXNMfxszpBWJ0bgMDV0oCUL/LfTxJKSF4/IIZPnXIPZOux7
Gz7fWRGOoYpLLZoflkIMGqGHP2wj/USxJ//1Vws1igFjikT5z0FMAq68RGf6HSlb
My3hwc5zoXPvvBHA50ATue/jQ0YjzSGiXxQ/jnX6S3FXQLN4w1veguKIcW0Kgy8w
vHNmFpYHXI00TJ9sJACKfU+x4BNHZDRNKjv+JiunqjH0eCaKjxt568O3R/bo7Crn
7WL9NDqYuQRySv7FoPAJRs56G7/4+h8UiCqngzBceqPQlSgYkvKdl4okTMG7Yp1g
qE4tofR1KTJbn9nXylgu0Ti5duG3PFAO7x8htvJY4naYCrd6yZ8Fc+JHwqoQrvg7
vvZnKItcz2BwjSTIBFgwI67ikeNH7KaHAAFZzl7Om70LRKf9jknKINH8yHkhCcyc
kpmfIDWwlF+2Tq0e4hsuctBuvfbQeIhZQ7Js3laT+EfCUpA5B/hG+e6WumX0KpKZ
0qQ+cTi6S6IrDK2WCRRR1ZVFSk0UfhlS2vzbQSziO+FnktzTlHH3vPmLCszU02AC
4noM9kejSx9HVLNB0ff2QuFSOPx+YUVpNzkZktzyitKBmp4PtfTLVj6MFTzGtIBn
F27WamWOaibr4cMltYxq+9Tg6HCfKjU/c4SYQCurwC3BtCs73mN0z1vrjSFF1P5F
mtzxVFWY6YSCFHSYqL9Yjwor563drsiaf9vp/dSg8H7qTzM80Esod06zY9wAcXZB
H6qOU5YiiKN+fDlityx+wWDKyG9+VnkeV35SrNsWqcpgeamMZqQ0yRNn2xxpKkQ8
hmUWQ2pi7MlbPN9Uf7doe5JfbjxtGRN0fLQQUC9vRet0O0E5UKVqqnqTTL/OO9Nc
47oDYRXjzpYIi35EeP05U5PzC3PRlQ5BQ+n3c6gKw0gyJm7anXzRTrxMbP9Caquz
nhrU6inndcXY7yUg9R1uXYc69NTZnY9H13HswihaL1U9+Q1m5aE9CMkuZqn2xI56
6VxDgiZcSd16CZazrRBJ+nonjVdmVlZCFndmNu1/W/vHgMvHb32uB+BCIc3v7xnt
IIgRK17TMJ1ZQYF49ze/vkPyfIe8PqpKkBec7XQtyrVx6RkenhpK2KirQoPjxpWs
cpn90KoSxbEY9GTD+v1wsmHmmu/nLWXfySXO6iEI1u2VvlaxCmCoiIEOkcw4zzBy
G5WxJsILzQA6zlSM0UTQY9JcufdX1BjOVsgFMy/0o1lXpqoU8lKPp2G+yJR9QQCJ
cB/yWPpOkBk98kbO4NkuBjlM5P01WAj7M/i+MrIkJD2w9CpC5Z7sFoj5D7kKwpSr
s0M+H5CscRUvZdTL+3B1WMQxjShhvjV9klKRBgDHSlsnqjNxq3ly9+eCJBuergI4
Yp1rFNOSWkpOg25gQsO3Jsy2ufNjmLAwG/8PneKUpQsHYg8SeXh9JNPyhdu9Mm71
1TJjOa8L4819hS5lx2RW6kcxgFd7tbM41ONGx4HgxlLgV3qWSUE1J1oxR31j6DcW
trvJN5NO9VctL/zfxFrMri5zHmAUD3DnExgzoavE8QHAwkNTS/tqnnqXba03ltNj
YNBWAcMVVfsKMLjxn8aL8ylaN1kFaTp1l2L+3yT0vZPN2YC9xHFrIvS1Ng/NhKzP
Ya7GF+jXoMY5x3zZrzkV7Eg7OuQOopjzHCugZHtWYBc7a0pLAez8DommB0WmVwbc
BP1xMKJLNAPis1MW8F7NlxwUtIv/c9TBUb8KwF57fyynaliF2aaBw6nYooYCVQH7
EfZgXGEHOv6Pz2cNkOdvQfFkUx6M2V4hEaxOj+QKHGmx9EPsoPL9ovqa/nsOe8Te
wB2IDoXg7Sf6yi/ncZn0eNXYGkcpsLc7r736yd1uRBq3Bcrhvr84lCMNehXSyhGm
dhNPRDjqjyp+hQ0wK0fpm1/Lcd8Szl4eWCvMSzKBpARPXbLGOT53OTlSOlfoN3lh
T6yVURW+A5uGo4EEgGZSquvKzZGMJyA7RR7rcuhPGhOophOGMsLgpg3hMN61TwHj
o9JfWXiA4SLhkt0BmBTRryCJvpCvsdcqsGPh4iHlDwIFR/sixcJ/eQtdNfPwIGLZ
7IFZhHbGNlfsqMCO2TxoVWyVs7JMFtWhfxubs+zQS0A0d52SZKMRtAtLWzejZjNl
dOjMRUNK6f1YaaBIx1iQjpP7VJvKEIPlGnREBwN8xsfqS4VSK6A6se+IE7WzfVqq
vAI0IyziUzhJ8rDN5szPXbNbunoaPP7OO15wx0e4aYFF+TNhEWo19PINIrnyIPuD
mojZqiDexMhPHu0VtvcbCV0nTraFlAD1AALqGkedALzdl6oAnxu2w+TlZBI5Vrii
+CAXbFHQP1Qrd++BoSA917lJ/sOcTNWkIbstUToFIgUyd5+3QA5bwz6JQWO1+Dat
tM6kDzlgb9YHWEmGU3/otnivHeBU+oUWvVKPTFX0rmX02x1G6HeWo1PwkD/d6Wy2
qzAla50ahGD+iNT9zgwlQmHT2DShT6z+bl/tdaPvtD6PWA+vijpLTyYSmemJxiDT
SIs0i7d6enSmmzsPGL5wMOwZD5y2kYwxwGfnwdEe/w6HLMjex3TzqSZzBc1YcC3g
EiSTWv/ur4oC+c4kQwJx2hM1ux5TZ8R/X3FFSFF1dgmzZ7eTNJc3EKTRVaxzR80o
9zV4Q6u4Xl3wnj9/2dS1k6J3o/BlVdCvQJsYZv5HkTUGRtOOUG6cFEkbh3AmzziK
347/HwaUnyD0a3mRcbUYv7ZXZDWNb3zR9kwdHYFbjtQqFsYuKdZZEhP44OgYl3Mn
bUmY5RH3sOKnypMUPgdfUFPF2O+aWIig3QMA784XQZ9ZCLf3F1lWw72yt8UnBe7z
Yar2v7QIOGX2ibbqroRt+3tlPkGlizITEe5Q/gIiPgjX8RVheQXt+iVIJM1q5odD
RV7IzbDhb2Mx6s0ffSK6SdfIDyywyXXNZIW3+07g/P6BordTRrppw0NaJCofphOb
WQzPUof+wlKwwH6tRBfUOW32ATWqi19U7Aaapdw+UKBebrPpOBcaa6JyLd2UPaa6
Zg0+5g3gPRrz6zpbEeey3pm7d9XsKjx56roA378MGAqC8X9zrLXppwjXuBr6qqGS
G2yGGAJO8+tpk7aWrnVtXmv6+Mw1YLLjXoTJd6pjRGUGItoqLTG2iz+ukZYCftT+
MjYYSu2k2MYdZ9Jh8RRlffrVG54I7M/LgCIw/UB0bAAVEPG45gVLPkcx7/h0MZmi
8iRsmOA6O95KJhB3M+k3p52HAzGqlgZuXOy+HfKRXxvWBIs1+Xu4G7mU+3QzUHmg
Plxr1TLG69XGXl6SSAfxs8QIMm8EWbFzkHwuNOlIh4dHIwXjmgL8haZPzD2qhX0S
T5FkXQ48mkVOJ6hoSbmx4TBBYNqM/8E8goT5lN1g5FqUsD8vbQu4SylfE+nRDfc1
Abb2QB/u3b4X1wiFFTIqKb6nZNmMkQ8Qv9N5BQjJQbicGQNU6K9OmGufmPCk6+Mh
Nx2GtxbvnyGhpafI9uHS3RyrPlitmINpIB1TAOFkKHXrqa53q2H78TCFzNGLExbu
RBsR4gSdZlHnhSD5G0NIczsMB3qBR1xPxrEq6N6f9Hz5sYU32jZmLTW+SA9NlgYk
U2/+t+xSuoZPQTB7JzNr6zifzatz4gIA5fEjM7FLZM0m3MVkguAy9/bGCjszVzxo
8CYlP04hU2JPXIRMyqonJGwLf9pC4IRWFK7LOkmOa47wGQW4+IXdZTl0fbof5Bq3
OXhL2k9FujdD9LqIwXIdRlzLa4z5iNsM8t8b71bRTWLz0ktd4R0n/5o0hgHdt+pr
eCA5gX4WUMLRfkSxRZsFuvNZ4U9o2P+Zx3s31EQws0YR66o9cJfrGDL93FGuhlVI
sicgqbZUM8rtfAx25moQ6UCbf4UiZocrpui2Z+v2NM6vAl5Ga4kEVQolW22ELcRq
eGsM4fv+HTBGLU7COAxaq3Xz9dHC4TWDiMCkEmcS6VbccMNV6YmWE4Jqlsb7N1jA
ntPPZ/mcNFBy5f3F99DAk8wXFOAWkY/SqiFvU9aKYvA7Dmj8aPWT/BMGX+vHiryu
T3dHY3wU97FKfki9F8408gH80ZvqkWxdcla8JH2TNu3gjzsYmdqAZoH0RNEJiBnt
n8n63kf9iwRnCnofY/P3YHRs0OnkSfpTlQ1ud9S5W1uAftBIQmjfV1Qnf6TDBdsJ
uM6v3UmCO55cVekEiA1/2qZdOzaTjxsYyw/Q+7I3YqtHXxc8VxLEDHnsnFEgo44z
j1IPmrIIHWIfcIGWFIdYtrXN11T38t6EL2oSIwyzvQYeyVP1CuOqEUD1i/JKZur+
hBzJypY56ah7f1c8LlhAm0Dr6kP8yquFfOgjpWzlSNHKZOnpKaRh40SAZksj7nRI
RT7iskDLeyCt80DaDJm2AJbn90ya/6m9gCRjFFbFGOV2ILoPpwr1nkzzHtGgkPXk
ttr6OwPteEQCcxGexgA6nokxr0bBvE4IlmysUOsVO4DyaXQEBRSGMC+7vPjtdkA+
IeVMj31s7AH/PyYNtygC48CgExb1NYjShq5T3xCEuysxQNeqtdL64hazwJ/Z6xdC
4D4fOj4WufUAqPAKOKTPJb+nQCrCPf9LZH+9TMyni/s1df3A1R8uqXt31Z47YQKV
DEj2hj9lUA1O8ISyO7rZs0oCYqMe3zBnuM4UCoTMWpICqWJndQZYc8GDCLXeLC0D
9dfuT2Q+E/8FOk78yynH8nYIdFYMyma2A5BA+GFxES3gsbUrLdYHGA83fDW+wL57
p1zlirKl0SBvkQs0JqvbpW5rg1GLnNfWFazsolIT3ghitJRFXx8jKPSD2Mj1ydf5
peBNX/x0nuSMR8uIio0htMkW/FqyMo0kP4M/MgJOjrwQgdX2maqpQPi0AJmwhVwG
1XZfA5olYVEr86DAFvB8drT0B3ffGoJLcSJsl39T2ph1HTZS7uzGWUKHWyHO7UOf
S8Ow9+p3MFHFBNFOmG7M2ftM1WDjpjUQAMmJAI867U60TKl1v+LIN1FZNhVJrDHD
bjBpUX/l39fWPfx6FNd9abif92iInlxj6w2WdXQc7WkxJvOMJoQ6qzvCR9KIFQT9
8tsPhdS4vlqArpTUNm1g2dYqM9Wu4zcH5l38Fbd9nIlEL64AR+eItvDaCNaeFXYz
QmKa5nZeyUkQskWjv+dfAurD13pvxrYqQfMQVwR0YXfji2De2OqpQINKBIfsX8Ap
CT6keovuFG3UjVwEnPlPsqfj7kzsXnCfGSlyb/8wQ28SkDayzgrk4w4ku9R0K75G
G75ilz2ots4+tzFIPT2tzpqJW8wdrharHvhUN0qZoXUul10uTXj658T5DFLOU93V
ljTgAlENQ5pfZDK6V4m6t4OC3G5OfjW0Pv68mBRfQfSyZzRalMy4r9JN/nkSq2sN
hmF/8llfbr3E7FH+/XFrC9Bzrk2iA3YW/Vl2b+7BUtGNoahEpqM43t6UfBYlHUlZ
+2n95VrQooMvXmvYwjnqpGtYK1W+MS4NdJg1DpsaXYKWs5gzAC8SUS901AoOVsK1
NF5yr8mli5BJPG2HcpkMOrIMJsB38G/xMOnw8vRVKf3TvaJLA0dOBTGh9N1JzJRZ
cOh9qNfrjR1ud5AsUUOEL3TAt/8L28JpWWVhkKLLZOfB9J1q/hj5gcMgE0An6RSD
BSDfYC7a4Jtr7dB1GpPtijeHL9kOe1iuNnt7BfAR+kj51I9DtHJfBXwkipdtNw5n
HIjVb/TuUy6QOVZR3hVKnum/MYpbL9Rd5oW8zA/7DNmYrSPgPJdXBvGODWjiPV4S
VoDeKs8Yj0+qDu5HS4grNBlp6Re92YTkkxtSg9om2D2TQLYgC47jQ12PBiTh1RPQ
DOKieFg1o6uJk/nDVpmrFB379qsDi4JvRAZiZxjWZDMaaexQCkkoZfWrN5zufr3s
IoU97ch3/tzKvGy48VJy0Swykm+Rfj9NdmSgFQNBg0FXoH1IPdrurZbmsdpTr/tF
gKsFnIdqo173H7DuqhjJu8HfNZHxYecemck4lAnR5C5BqoGo9N5RnKHHbThq46w3
sE73J6ruwbiTIGCGvZIOiqCAgqYxV5zgbRGCb4s9Sw0ct7rVNRB9+VdbEiGM00XZ
62hS8GhcDgYKRfJVCjtWqPtDlmrpaxa6CWqrjbAzVDmC/eXAaA2o9rb7DBd5Zy9s
dPn2tVayrAvPxitDzLZNs9KHggaypTqzx08m88DOBehIV35pVV71Rq91Fw2+P7Kc
AxPlHiGpagYtV5apEKtj8L1Ce+zcP3Hl5olXUJymTrTDHBgZ15c1407gfluEN5TV
+UXcBfr7OClQ4WFMenIlFziYcHrH8uT2X7Ws+eQJs2D/oo1I3m1+URlA47MR9XjT
ksZ/vf49nL2gbHTRt6/eAPpq41u/ZLBF6I/iJdk39xcWUEesqU/uVQcJS7zmaaTM
n/Qhr/VtQVR/EW01GAfV1VZFFGF9a9nrMbJMIhY8oLcYZSDMK3VGLiQ+IQOBQoL+
uZK7q1HwlAKxV8ideMnfUjM7OJiMF2fTWcl3havK1YuPsBXNGTsdhrKCG673LJPT
h4K5PK04Lq6wGB42PWE1FeKKPKJfShJA0qwqaUpOy6K1MMj+ObKbdihKOz3wnQsT
lUs0BYcFj/F7yrEMgT7bL/G/LCBTxcub9ko/anMq6bSV6B2K0z5MhCL14aN9er/U
MD9PZh7E6ssxFSvk11MFiEOs1UoLmZPg1izoLmU1hVlOgPYQAaF8VNnQmwDeLyfJ
Eg1gVgyb8QJ1teW1T6iHqbDX06HeqFA41Bi4RY4/MhKKRAOyE3zBs2bpdS/izSmB
EYTIz30FannHRVrVstNFEAuYBcAL49BIce3j3RJWcOXqPstD2dqMDdAFZcY18x/u
Impi6nDJ0vrmW+xDBxDgKgaWgrket5AbCNkWKZz3k9b4O1usOcaPSm1F8Cp8vNwN
h6Rg3Lq30hOqMrqZDFSstDtLbm1+jgJJi2GAT+fn7v43k1scnwmr8co0fFSXhvGm
wII6xvhInvxJ5fYPtBZVB2J8plIMbLeYPpYnrk2zLIXto9fq7gZD5TCDuQJ7u7Ww
KVgOg6N9cMn4HQL+b2wvrQ==
`protect END_PROTECTED
