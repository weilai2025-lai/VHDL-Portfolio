`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X93wWInKwLYsW6Z8oolctoDMUoqKE/ZYNzUqMsfCGaXdxCHSlBytjNWUooTEyIiM
q/qm2lgY7RgSd93PlmIjL45SkCcQa2k1qw/3PHXxo2iatDD96pVF9IzidUZru5iG
h0WbWXLYJSVpgA2RH2IS7OyuE2a7w0gJ9S2Hhh19XmyZjEczqo1tANK/62LLmDy+
9dhwLqM6y/LV066LWz/guGQ+XSotM5DGo07kc0HHoeFyxKoL7F92hlWSqBB8wxK5
1IdbYDeEqeGT5SjhpqKw34udPr+VTdOsHu+qCWDjXOwVhju8i36Fsu/2f2G123dG
SXfiO85eN9DwkavvorpbPzFK1hqhfTx2/NRFwzjjdUWPUb5+LvdkMasVR0J5myBs
paL9vtvV/uhQhYGcZ+Id/Vj7A97+kEdeCCGAUIZ2Wd9VnSud4Az4YFxmbCHyPgE7
/Lfl6Br4+E6HJ507QlVwzoQEdFpRiKiOmD18k5lXjIPy/L4+qA2dayhZ/Pbu2Z3T
+YCqfOWPVay8CaVkklK0ApJTtHZoRDWxkkO6ar53ZvQtH0NLtZB2eb5wKDKIsi0z
z3yUSKcT46GXj+sM1TNRO35wK1byXKgS3ZxhY7yyCvTIhUKR/ttiojhw8MEAEa2y
tdWwDw4IplZGzTcNkw88wnXdsmlDLtpJxzUkkCJGw64rIdhhsN+xe+bksyaemf4U
1SlpNmT5o6TFjDr+rkbTtQtrnadtGczduB6kYrIATrihjZpOfym/hvDXoS6OhHif
qyGVPA3RU9jinw//dh6QGMNmOOSElEwffI3mkreiV7sFTadnC2MuJAUewDFDrS5s
aODUN5g/vLlk+YZGG6fx/jYuyrGvY70I5kJM35IyjeNZrg+ubO4hhKlCABR1hh2j
UOlNyj33YvCICo85TcDHirS0w49AWC0V9N4XDeIfUEZeL/FZN/ABlKCmORflQkTk
IZT60W8zEf6qWV3c4KFt4sDt7OStT+jklTXcUyyUfbN/P4g10opdkheZQes9fC4p
RqFe1L8XFkW5+LSZqCKfWzFXh26Re1ysQnNlnKpD3Or4usTan6MzSPNAiLdhd/MS
weVprBtcD3OIHiSgVQ9+cV8ZAcNX05Hcd13mr3P5AaUsbXqux+LphJi51bCdNMHD
m/ndAD0qSbTQa/+HWNDf3BZXkcYnbSpXQkr187A3PUfs1sP65d4ofeiOiXqib0sE
MzB8P9S3iDC3T30gASOQkzGJ64jDG8KCq3ENZgsirq1j+G8vDbzWiw5x6yA8Pmdg
BbIplBW6FAdTcEqoKj0EArIZT2azhdn+oMCE3btzrWbN4Ny3HGv2WGXxtyXLdwfU
CTy7YFDzVqcc6gH4JqhSZmIKvoSd+xPGsws6DRV0KiCdsB2s/cGVE/tKiwJUQGyV
6jqM9HIurJ+YEOq+zLH+dTd2ZSV7VUnEFt48cgHLAeh/cGCnIbVDPrvNPSl0x16G
NBFhhxjf/2L0mtPtMeFBodEK4MHzbD1Sxqt1Q4/b8DlyWiMjA9ex5xbBCXbhKJSw
qWBRmD097bcJ5e2AqknVZk1Skybo/gSjl2yxwwz50PyOOe//Klpuvjw+jVncPFvV
Uf9vi7LCrYHjTSADaefcDa2oCZs8LNAq2gbiymKHw8EVa2GrpNokg1aROI1DRrGZ
RdZnnMewKAsqpssqeCHDVhibKR7eYF3Vgedg4tnQguaP70r4qa/TdHTcdPOq4pha
NlvuJFR/2bILY3xAlsCpK5Xt0incxBX6ou6QgHlq5R542xkAPOXGIdaXtKkzT/uI
rMJyMD49smCpHLJjMx0WbOxRo3JRnKg7dSX18w8GJtPut9scw0ApMskbTo7JGsD4
ZkG8kbUScUcfsWBp6PInE4Aqc6hOfTngCfbJIgBzXnIrIqvwbPtyIleA2o1IiOyk
K4We0c/aKjcFZp7W8b5vVvAJ480NcOQMFn1yz+CEBlnvV0HJy2XlP+O6fCPvqQy9
VV0GpOdozuL5AvThDvXEreoKZaBVJM8okQ+zLp4N8g7rJjMpmst0LAZsRonmUZlx
363CzWYCSQPSCCkZah1sDcFmG+0ncJWhrj1WS4T83j5bJnzfMuiVc9zL/lGzCZ7f
nE2l1Iq6joU6F1sjG9b7izCofeB17myrDQxo/N8oRilJrUfqTJetdjN6eY9bSVq4
e8nhKmuKACxcNWf54Vae3naeADYkvdtQ80AERMGy6PvJtDC5uSuN/WoZf/U+jSEq
zhtQiEH4gSmtwXHk4O3c4KnAJIj6CCsCxbvHi7Z7KekcMA0KZ72yEua+4EURoLQf
YxQRnlXp0ode5NIoPPsUdq/iRhdmkg7yaBvbcNy1ejdKpXyijZFqS4vyFWTW1+/u
OwphoUn1QhcIQ4JfergEhyM7xsfO3OhudhItEwjvo5FQfQJWLGxFHjNv0N3wi4XV
dZVrru2DIyKbHT/CDMN0s03Jl3gGlNS8CSAEjwfZb5HL71PWdY9BsViOeFVD2L81
4MzTY1atVXAwP9ygGClsSmOxBvY9t6HB+A9eq98DxQesIwJwU9Uj3WIaj0TNAAv5
+S88D0gA2Z14ONx7KFXDq5H1lytFbjMHf8jmABWUG2BwPUxvm9C8fTaISFl0jZMo
8hmMMHZAcUGQw4olNzbu9W8mEOw4oBguwZJzFgg5CYdbrTufSFExmunEXHTCNrBa
r7WdEwnXZznT/c7BGaMQCmiOH+q9IGFi2ZUWLmqjkMaogOi1yNefADwq0IKFiy67
CV1y2+//aTnohRQlaholPdSWhmNiUfzoWxw2t6+VMx+KDgN8/yBXnpmj2IdeMfoH
6eQn5m67gHRFPggvs6TT/ZJcjcql4Szv/Jc0xDqXhdUH9XagkMXcYutFQGlb8/F/
1HkwQiGx2R2NWhKg5k1Pmj4hwArLoZOXleUexU99f6qU1pqulz9Rq8a4LeXuc344
rc/iCNBaxNuinqFBHCKmHfP5ATkqLefCEr0opMeh4orYeg1DgVuQjZsDhqyfq6Qk
KsmSVLMR5o9OuBifod+ctd6TmG0VApL+lcbDD55GvIVIQYbMuDi0ZM3GmDNshFXm
/gBJacgDmlBslWj9DhPs6p8PVhVmH00eq+J+D+KSfsvibrmK7yYWW1+kLFww/XBu
HnhkoWjsOtm0zipSqAloGWAuk1nVXlUC/u20LYzo7g/ljM9jcoJ0Pxp5Bjk2NXIz
S2dFl202I1lOzLsvJg+xa8wVaAfMBD1lwIy7ftVuH947NIyPTDHTDGVTaAZq3TRU
MIPL4J8MDv/KkZZAtMbyZzeQZgSo7xtdZTfRvnYyvtsO7Kh9q2owZvnpVilReS5I
O68Qbq3tyYQjohauHQJH1jhjVdiAms4UbARuXAMOJiI1xoSkS3vaNRH39kdLqx0H
YDkX7MWkNMDw6lme9+0cMczflDN0p35zE+SAzJDPs+FO8bHq77LcFQyGADQAj1QY
J/PY3h+vjdt/X2TUNk2Z3gTYAvE0GnN0LvM6bcBP5HmqeSYGtz+Yka9tgi5yq6oQ
4QViqR5M3Ga1uwNcbM4SCNwAB5V0M++uySjxvjMdKg92h9DpSAYwpnat7tiL7iES
ma+Sy8uLXG+n7bmHXBQtwzhOA8MJXLKHbrTR4RveqiUlPGor8ogF/imMQsBnNk7x
bJocBwkHnW+C6emYmyX/3Q==
`protect END_PROTECTED
