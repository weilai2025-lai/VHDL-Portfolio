`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJXmuQ8Btii4Cc2f23VDUQTE9QPPhX0OYUGrQltvZw9jLnH5y3k+sJ5wFz6/6Ky/
T67CRU4rqX1zBym1LbbP9Vo8DObHQqdd57VZD1O5FxR/AHVGdrwkwDWDcdRexEsh
0q8aTn2xbdTJFKw/hVlrxhZ0FEQu8OIDkqSU4l08kOjLeYy7tAAzKFjlZT/qn6hx
HrK+sexCxlCs6pbidHsj/B7B9AD1lb+MDox/POhIQD2HP/x7KmuYf32WQU0SWtNG
ug91Hm4iYgbr/7HuzPFmN5vuWnI/F4PgFMoTb5XN1qTL0oNDXbZ/NUys8yzf+nxG
IaryXuQe+Wz2RDsayTwsErIo4zaJwtNiRU1zhSFpa1klctWoupaALiCOrNUF6CPd
YNgynVkJdrYHzB7MK2isuX7O4ZEqRxvqT6RjLoBX0gXJ9VprPmNWhd3Vx67LMLyr
xSLM2Jo2sHl5sE8a/boeNIO/CeVcQWkCl+/YCmDZbHfw9ecrL+8gUaOc538vOBdY
W14ReEkJqdCXVrOxebyqdpiG8/GhCEBwwyvrHQOq1bRWrlZbVuxo/hyGtfSr2LIl
kpXrQuLivR/85EfcLy9bP6+AXH58REgMuZ163nOHkhXcDChWnnvT3+g3S7arfKGR
HFuRUITBywx/J4Q8S4wj0sabNE7twqwLkjrelyjxWep85AK/M9hYDLtzQBlW7xIO
RzNYkkzmL/O6v8Oq+4ouqGGAM9r+2fLv1iD30XVC9+ILUYVVzqBcvL5v+XUX2d0g
Fsq4MKOJZzwo1TVSOLT7ptDDFTMB6lhdjA6W8WZWTBfpcPGn4DcyMKuX3y0DRDkf
O5RxJuBdoaRhE2FhERSYAaYyl/XUDgelQcJNRLSo60VLHRmHiHodiRwZoxg+0b+E
3rIIErSJo+Vp/elNwOD2OGaMjGBi/ZRAPRfkJOTQjxCF/4wf8idZNQijFFJOouXs
WlMrpHIk8kZdNJETpBUtprcaZw27qdxlbe9il/w9OXqFTCaQuDjAuelSNB3DIycH
dfjsxYaAXRPApf9opkjYh2i87H0W8GnANZIhZL0NfpNgNd504gSEvhNKd5UN2Z/v
N/HZhfQq49QeKyEHwuXoCJcXVXQR+6ZL2Rr7UGmGxcshXhwhzUk1P5PLLlA2XEPC
NooFKNs26o+bqmRZNBS4ACkULm71qKEl2HrsctnC7K1qbTTTYkEBLNwFbW0zltTi
Fo2fRVifMZHDEla3maTG49piWS/PmwYlUYtZiP1hVZkbRJltdd8BnQXmFEpR98vh
j6TudL4U9lsFRyoOarWEMnm/o2fDRZAQhRe33zypJ6xlaxV7GxEM/nTMfvL5Apsy
bl70bwDBv7KQAUcrz95z8I3MEXwFlyNmKA6/vb5PHjt0NncaCFy0wZo5ffsdNfT9
tXGg02gPLdrdT1Jm6U7ZqfvuemRJrQ7Wrh9zm7ngWUvZJsWBdWhSMl9k3fHYgFaE
u6RhO3emiydGfuNeSt2966Gvx7idyltOdEIgmSbYvMaUu8yNMoXiT3xReTkO9GO6
XHsDCr4uXgw14cAWuublzc68JK5eLEjRXK/mbwWON7asNvlCBiOCO3BoGfY0kGcD
b7+hq5muD8sVP327NFX3NTe8l4cuPDh0FotcsUMaYS3izCR5qc4qPqVsfQ8v+o1U
NddRH8zClLfBxC1jxQxobjzBspXU/CYhYbtAk+On0NgDKMpMMfkqr3PYB4MYI6nc
dAJ/EOPYhKAm+inpEl4OXzxeFjBsD1kWmhjjzWLGqoitb+Fhas6Svfo2+Pi+WXWx
g8KyEM6YAiJ7LyHEIv2ciPJ0jRngQBBRrfpci7nn1uj71QhMmQL5nsNySJ4EnQGI
nntmv8m8sQM1A4zV5meV9gaFLY3Qr4mfLj5V34XdPAK84gBeKrISDcS0tuTQkRHM
vk0CMg6GzFN3dvqbY15BLovden4W99V0zVKKMHZ8Vc+9gy1CTDRsm2tNA0zyDez/
W+Y2BPufOAadqCbGTW8qpIh2vGIJgMVK+XXKM1bgovNB6NHMVFlVk1TFqeQXZGZt
4xZGyRyJUcPLqClH8QIOFr4Wov9Khens2FLk/97M602Y/Y+nwW2cPELXYuM3AsvE
a1ndKlHeqCVhmR7/FSJbJ6+At7hCtiXQHMtE2WWknBPWTiy1/n1HuKtKXyyiRQuQ
fI8D9WXHN/pYoxrUT2tah9tgc2QKp0CgbZ3hdOoBIR/mwnAomLSxeWUfbpEhmBNJ
yX5BnjisuzCxrQG6Wu7Ma7p1+QxQGInwvDFFhheQB9vELD52S6AgHP35yEhXeAGg
iT7jP4YDmbDQVI7rL0hU3b1auLO3q9GuyqcQuHeNxq7RpPyqbmPdEAmM38hdZWaD
f1oblPJVksomHoeNJP0uZ4C/0DoNcnduto6chXJNkIvE5BcPUn5rDAhC3sbpBdgR
8kVMu6ftRCmBS5ngYQFbnRNcoxiV47XUVHgESKSXAONaYQjInunK8Rr3Brp2WbFh
EAyBLKBfNiC8z6KD+3NtSa+kvpKkeuMZPJrXJBaXMWeLTxCGZAZvdZWEdBPkyAVq
r+WUxyuidCkwJM6zp9BDeb5SwN67YrftybsLEZT7uYBf73uvZGkVOTiuRCOMw6Px
2hoeLg+ROxl7qBmsHI4uCURylPyC8DNSGIYHnpB1HplS+B7TbOBa/BdmSg4KU89a
lmd4SwjwQl4katoPPjhC0LRsdFeCalzORLPaogzP8KBTBL3vDI1P0beEY3rpKcV5
sJef3kkWjQu5SzEAc4d/JalyZ4s7HiV4f723sVtUd18EzbZgCzKl8DiD7SzW73LR
84Yd8a85P1kpMuE/NK9Y2qdOE+of38lzr/5dZAU3Ikw/JBiCvBYDqfzf+tRH32kQ
fRVf59ShLM4sPVnrShnpDaADqIsvdSDMMPmW3cNkgcqOZ8bPib4D0tq7gmULLk2U
iBr+YYB++XDoVjZ1fJYAkp8MTj6FiZTlOhdVFFJGPSe3DeZbmuw9jETdxbheqFkP
ecUdUJaSDsnt1vmodELHOTDRlpv5/0+RxcA1Xacx0pqlMHoJbL8fn2fCCd41SMRw
12lz6qnpXFkJ9ZpQnMW7FP55izN53IDDNLfZF3ksFoU52g4X0mb7Yp+qLWp3uBGO
O0SugJyzqspEdPEK4Dhb3GcHo6WaFyF2KSztboDSOwPr709lCYTnYe4R8ODI/Wzk
bSvYyu2Brhw3yJJWrAXbxhB4a3dLGuem55UMbZAEab2+nbOIwEGe6iwbWxw3jr6G
8tMAPgUhx9WYhZYYgYaW/43aDbwo2DG9ZnVC4BAvpkpwRARsvHhKcBotOKGNgy0A
5CXaUGKqJoB++Qwf97IW1qTcONq793ac64ZpKkn/QiHYEXGbLBKGZ6s2WZqPcqmv
a38CHg+bvOXAEOV/HXmPikdP/CitbYA+56/7PYFedRxUDOh6017NB/AUmjrVsrtH
qzICaHpaJcMFq4jG34AbHPKuq+52bBPc6gKJBehW7H1MWFu4Fq/LK8nXSlcXqTsF
hV8Srb+shXK4fjYXMhuExBaup91OOLYXx6UNHqod1oHYhKnIYZp55n91+WQp2sXB
VJnypb0xS+tURiAlgAS+kNDHN4vpUbaKpd5f6ddwm7+BgrGaNnf4MfgB0ZRW2Ai9
EYPEq2EclZYEfUbwj0IRdSUoKBkqi97k8jLXKRFb2XsM02OC2Qgy7jYKv+zWEO1l
d7Waqsabm6gBZ1D84Wn+msrLYg4FM9nMR32LKqm9c/SAFp/EhcFHGJVPVwtGc6yR
eBQTUhFBC7UilKa/pHSrSY8ZIrlGST9pw0loX85Y+lrN51Tv3m1+AlxBEO3dKVaZ
cH1jUZFxV1telyH6wun/pmi1QbC9QDvSlw23H1NaBAKjxMdygdyg+p55Y4fjcW6x
O2B0fVg5P/L15uXK/opcbnN6DuUZtUUtUghd4c6azT+dDEygPwf+Ymj+b8ujGHip
7utRLZUNnZBB1S2PfN83tich3B9GE2Q99aSDLIK3NdB99K4rpeMU/HsoGAZTKAww
/mf07qpB5MTKyo5YT0uSKx4kHxpPDE1fnMHOKibp7copgvKI4Eo/5MRs78JCAemb
ZZOZCHLBZzM+Q2arnPgCGuqP6DJloovslbqNljotj3KHo5MG8SfGs6ArxeyY3aRH
dBFCCLpin8k7yAMFebT5jhokI0BNySK5UM4pgsQMoBtfepy5EjXDgDNWNRGrzUps
CbABFVI7Zkl0wFq5y+76mWcPOEBvLYB9s7C/J7sOMjFP8vI81abbfPngyuIdioXG
D6kOFFTau1q+5HFyeIjf68xIibCGrkBCyWlvjbMs7HW6PwuP2gxFDHk1IJZKhrEX
Po6OpPtZ8Oc0QPSan1/v0XL6Eq7X/SV8vSU5/0S4wvk=
`protect END_PROTECTED
