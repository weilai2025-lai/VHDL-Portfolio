`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sElT/qKU0NOE05pv9c/cQn7lucqH7fd1zRqkwYHPx+BI8cXzAtQLGVCDqGKM7ozS
BaGkC76MLxg3/yjBR8gFiEA9lqxqiKqUHggoEkN3ryTnpeYlZThOP2o3gT6SbpJG
5AEFtcmDcEXBYLVKn6XBehGRiqLpRp5ymD6e3zA2ndoCDR6tyGGVN93VDrUoyd+e
6P8AF5+e5qLDQOfXvzVSDiz8ktvy/wKEPxpHUru2f88uc/WJiVdM1GSuYYt6Ht5B
nMAJY7g6DLLIKgbOPQhCGIZ8pOZaf02X8OB8tXjkxC1H5HRn2r9PyL8nlnCokq1a
ASrltiFY60DvMUScZQ+oHxhXuDF5qlHqGBKP2U3s0PoK4oUx3Avpp8thBph8A1AI
aYWmn+zGvbkx1TMo+gtmnA2i8VHuPbOmWPh88W77R3RP8HKIFaJiVSjEtExaRodr
IqcdHuSFm0t0w5PJ17GSY1nZIfyv9nsgTWjJfNFlmcCIaDZluDEHb2upogeBk19h
v8R7MRsfv5ckbjvBF/m5wAUDJi65q/TcmbPlA8GJobSqrMhmjtACO4RPIgUbuHIK
SQRrv49TR/IXlxiD05PAeoxljxWrUNc7SBp7NHfvtWPQ6Bu9KpBW+WFSoPau2lXn
SVO00I9h/eS0eUmUvTNHQBnn1KBn7jYvusjfiZTGZmL7is1H9zw9mxIu1snDiS4I
8ha305zrxOyynHV+vQCnG0ZppGLLbdL0gy8gtyNp9pqma9dt53ZO5JBwS6iyLRSH
yg84lljU7bhWTWL2tyqYvIu7YZBhu33VYlZaddl323ZeSxM8JRIl7d3eWYEz40oH
kuGTzEA0IZKg77CRlmG3YhTcXskCtBCk1+lTPuTux4NHFVz0tvVuwcvrNOnDznqD
n3rfOqEQJgbvYWvfXo5zXPistpLMTFHBG7xXuyyr9h2BRSW9qknbMU8CLLa58Yoc
1erbkFMXED5eO/5/poKADGtS+6o/V3lLkQQzuBcAmkc50yXIpAAwfqhWilalNfxp
fXztfncR0olIWZRclc/n0tFT1Cigb0EQpLoZa+oI897O7j6O0ZTiD1qwTMQ6OjYi
zYVjnnRAmNceNloe5DoYFSfCbyVza3WMlLMIIWYEjowkQrD+lX1z7LWCdgOq3MLS
nSAS3LFTBYPihPUvt9wLGejlz+UGkKs342b0hsosx+1WbsHzTadq9MHOk9CbMa2i
4S2WpGLfUAzyRNTuf36PMghAPuRN9JmIrYMns4d7urdmT8vTCx17VBJU9X/TVrDZ
SRiiSUen8qScAmWY3pZnyrGHxWVieINdq3dZcRw/sIjO9+IRCG2ArgeEzXJ0eHpx
s8gTazQ05glHQ3GukcTAhO2HJQphWtNRtgBZ2hsRhc64E5oHaggQGgGbB65xdJeJ
nSbCVELdbZXBdynDtvmMnBiKIzLpLUfWVF+raJwHHvjtnGJ134NDeQrlM0RK6hcY
`protect END_PROTECTED
