`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdJlcminCFrxc2EhVyRfoPQbETNIAMc7rNWf29nTL0+F/GP8p3oyaUFFgfureUYL
fnjMl1i73kuKoufAY8BGzezabDe4SC7poatwHjv8xmavNpYIzveaHTglloPD2qVQ
dPDv0nET+LELXB5daPSkrF5igCZ893JlIMSkUnG4IzLT3LYZP2Xo0nbx8ah0UI0X
bRrDF80QetrGBw+Q6DtMykcBf3cG6OhPvYzjceXmsPAPE3U1gd7kWxUBOmKhLFkg
rKm8HOlHMsoAAs43sc+8HvVc9FTXtTOJ4UZ+yZAu3FuO4qe9rRBT3ew4U+ESaRDo
HJcri8p2eblmMDUNCc4DRUXzpJiQWjNungTnplSPNfTM8MRmxbj/lkv9sfpjRSux
Ea99eBZxvyb1TQFxz0WUfOw20pZ/zF/ZGaLp7922dhafUUV1P8nTB0ofBSxj8Do2
4cNSDEHF9nbM4c1ESqEhVwLRHIvogJ8cWqCXv6KJfVWYBWHDX8CipNOWD+VthMZ3
u6EwbiagzeKYX1VRn+Xfyo/X8zZvNWr+MEOf5mG7ZJ/jjXMUfiITACBmu2442gz7
1spNhLOwg/tFvP3BLUsIdudEJFwvEMEOSEjuo6OojKR7UvkSroEM2/PF5en/RZ4F
F/d/H0hF3V7NMy5Y3jHtkabs2uYgFCBgBT4vNh6puKZI3omthjOMawN64sIrBikd
LG4eB9s6kCucrL0mqDOi96+lbAPsZ0WzmmctT+ukZyKO1Igw8Wlq4JBjr6aFmo2s
yGe0/AMP+digRwJT4cyrSQSQ3uQ00b+Q3wMNEobrGaFDFPTk3cw8Tb4Lbgl5fmzg
6iMDo7mGWpeuW8vY6MtqjTwZs0CfztiOgJlhxM9qegk=
`protect END_PROTECTED
