`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vp0Y8DLRXfXf0kCYHxsw8G/YlpHtEOfcnjUuWnag3cvbYGCJ7PGoOpxGYYO78EU+
9X8DrwRlDCjTsrLwNA02FqyfVS6nBoUKXoLqWlZWUAfHy93xNrLx57DwiZ6dXOHm
Y9kSHvgYoa756G1nqmtVa9MhLKGz4BfW4CPCQcUdSzO4p6G9RL20K2IJMt3Th5Xa
c/Tq4p2LxNG/TvAAvhp7tGQYM4vqTgU+DiiPxqofC8tUdArh+JNN3Pnc4ymexjtI
9e9Q1Qy0AFm7oS6WMKWXczzXpkKWPjXQMXWFrQMjS+a50ihMHYIyiQk1X6EK/Gna
Kd0PFC8zdfLHTixEEKG1dVnGJ83r6LrWMxVp06Y3krq5WUwR9HKRPQyTRoQO8mEu
5n8Q1NhL2mO4Z/fMn/+aUFOgHIWL4NSaMiKkvzZibJ7Na/KgKgA3Caj00TF6W/2s
O8PZAw/6NP1ros4CXhmGRIO1ybSJoovgmIvr0992c0DNH0Rb4Qg+HhV8iMgw3VW6
o6Edep6tbf7ZJNlFtTfli+GO/99SFmhipUgq1KKDFbhryG4b37g1ux28q4QCVs1e
Obe7psUiSzzhJHvGrG5ZBSSze2rlm5dO2kGYcP3AlpkecarV8/nsjtiPqHaGTeH6
xP4u3lckvT+ZEVDd7Xp3wvMXV9dUCU3+E1N6+vfNmmen8HT1rr+rg5IX0vQDVJR3
zNuNB8Pac1jGsO3AecgtCJg3EAAJzdG/szNM8OZtlGb6P8EeNvW/JMdOZ/i7ULFV
+KrR2Z3zKMIfX0hbd7HRlOoZWrGfyyi75JtwO/fr5Y38mKh2jUCmFCQbAoyPzabg
mPKcolyaURjnIZDiZ+q0bMBBwSsv2f4MSleiPbqABHdsg0EO3GxTemn3RFSSdR6w
vjzZwW/8Fca1askcGtHiOwFaUTSvszuE5zRn0ckZHklRuzLXjjnquBB239DO0dvc
PqQlTJfUOH/vn7CtuaRMF/IFKNX72g6vmmZ8+o1hUWJbSOQa5c6laVhp2DTmijnh
8Z08qF+OCeV1eb/FdGjEsfozeybGHoHdn7OR0Ty67Lqqemoi2hfY/iO9Q/OP/h1j
qzn6A9L39gvzXYRLrvQTy1cnAQsAmsQn3tmNVn6nNR+9bDTU+8/2dYzIOF/G8e+x
tgdlOn9LbfcI7rJ6Zn1BwBYSNpiLpAEdKBCJhrcP5wZDdvnEE+zNLXDBOw5KNfVv
/VJBtlOR0ENxGeUKzTFk9qqnYGrk6ZTyTG26FAjOszCPgSEScHIOG3EDT97gO27L
Ivt4KRc/HzKQgkEPrOiOvuvf4/ismrGI71eJ+bR/wJ3uhh5OY/kbEkpmbrHIOSDg
WuzM/gWIaFVAylcNLnisOiHXk89cXajHaInk2jrbPwRx/Ig/1rmgQv4mEdd1cLvG
IlUJ5W39yqYL5gJ+3nvewj8x/Id2xxghSIfh2ZfS/XqVzoCUMvM98ShjO6RdQ9eE
CYbWTDuqR7s5M3u9XPzUPvPAvJXgKvIctdZLAjS5PZ9IWkRfGUPR7NNAiJBNTUIE
1QOLZRxwBljax/AWOjBFcZTWaz1W9LshHeBiVDHE4N5118hCnxgD4huO+ayek1ZW
HdHkSp1XWnL1gPlYpy/jW0lwMbSgSG57NHBsfo8SBecEsUrc9W5/oLokxBkfEvkI
4xAxBKOzvXllVJl3lZVx+qLsGgDUJatAWUstxro4vjff0UhqoYXoni7NoZFzmR1v
Ex0o1YIYSx4PvjZAfbHOdgx+K9/qFwhmTBMFZUkvS1rXSx5rZXAiI9ADH/fWfdzs
FCrZKWGPO4DRxbknaDZZ2+I1rjhVBXQnriVWTa19jzLCipH56/hzXU9Z/UIn6v+9
Xzuskmj+E3YrimyYAzGSmM1j2fYX4hC86hYowdbffnR+w4vKIF6JHIQcnHq9/pIV
`protect END_PROTECTED
