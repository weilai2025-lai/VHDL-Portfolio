`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDi2TFMaHC1tlNagDqJyLdUdZR+juFWWhrlZX4KIfyhJGM/6x1wTOeG4VxgQgTyu
UN/75gHmy4v7GhO4uBBkKo7xdxrl2v3/eOZfPrYyuzCzPU1XqaDg8MiF30Q9ZNQ2
OZWb7wpr++HKqjwrJBIRT6m2mLFrRsB2YSpD/o3Jc+xyb/QdoGGoFOacqJHw0uUO
P6ldJTlas9IfpAsnIoV18ait+lXIvMF4oH0Ksf4EGFo6BFiDA0LfJqDnxFHLFHEj
N6KIE8GVUKZN1srckapj30hhQKMXUAGt9vFInQrTyopBytr5JRz1cbALTIA+Ckk+
FBcfXLdLpeusNGmWCMDUe/dbCOjT5IcVH7W5V+VdfsQwyflD+KCpMZ+aYaaSB8vP
6vf6f7oZkJLONhGtQO7mn9zhB2Rq58AUgm3jpPSAhf2sZAaDKwS0aAUL4rXPd8un
xlhk8VXbVZN1doEwqA+bU/ss928hzEKPyEejJWx5FzvYwUFIXYeWbDzn4y2yfjSD
rA3dcR7T2BwZHsGmAKDjTeu7pcS7KIECriAHh7hu61BMIeGmCWsFgmLVDWtKac3+
NKFEpT5dHLtjW9m9Navd8HbGlE7/hmo4us+FMY6HNPI0bLZN4YAOxCr0giBEE1yP
MuuPdfz1R/hOz7p+zooxmDHQCHsKCM8pwZcfFFcJk4iehf7BfERREVj9VYwZVGvf
VNNYF/0WQMXj63Xuv+0GeWu4W7guboKfvkBwkUc0cuyZDXvDrfCki/AbWCSnReDm
xbFVch7TkXoBwRf5eHZjFupjZl+8i4d4YeM2uRmortOdJgoaasKaWHR+2OBvaCnI
uwu/65eq3lAiDKwDm3DnvwkMpzZiUSw3LXYClqDnLtBHDWeyz1OFpl+4zAQZD6Nr
LYEtB+GstSxB80jF1xrHcIJINtdiKJWkfDGgivmmVQpBYo2ZDLz+afXkXgV7KjrM
auJljeW/Ge8ipmhVhuCLunQh9PGMIUFhPv8doik4MwmenssGlcDLpV4TVSmY/Ohq
Nikovhua+8vPHqcEo3ofzVZEPA7HGTrJbzOMXcuAzKqqf16o/CHL8kq+EBCMAWgR
CrJunqPe9G/eRfaskScH1HxjMRwSvInJrDZf5cTI/53gnTZcXQfW3yr8Jna+ws/W
BOTiTQXLVRU10qzhZytG+QCpYl8O+yi5hAZYiGP6hapYauOwcND9ia6toDr0acu+
rWBDdh+Cm4UoNfnBYZaBX4TzK56t/pIIlug4IZC3i9tb9ZWfcawY6ekfQWLvyQhF
kHNNHEIUVeihM8l6KS2m1eu9qOR4unBzYGicvpH5281bQoUqeZE6Zq4FrbFaxPfw
3u2/1bRjt25Jkz1mwtGAkigrHOn4Zg6qe2DnujX1kArs1pMuFEyosVgwRJQJVCCg
DxndDQkAenfjNStfr8Bu9ARtkWxhA4sUTZPxYZfwmk7hdCtd/viPPAz5Tw7pNrjm
lEPeBYK4S2/qcZXzgciiFPac+KqGBRY6hb4b5q2IrE0hJXRCuTZ8UJF4aBicaSDu
Gm6te7WUsvMKcKcCgW8o+LQIvOK4kNv4BhxRWY4BSL9o0V+S+ebJvPyyafN7poFg
Ac85eTlN6Hg/zEXyLlz+WIjQ8rvoX9QOAAPua6Gph/0BqhYvBeNcGvmDW1+kCM96
UXFOpPuuL9koChlQ5kSFs9JfmsHlRVwLZhGFCm4N0sCusAniZjBPO3XbkLM94m3l
VZNmjDDuqJxUk64jPzPBwBCICdskm8ZfPnyuHNw/Q58ZgJztUDo57SBveOq5p+zt
B+67rtn0LxB1MpjU2G7Omcpw/hxThiN6E1fgy/FsZDsisH/TKAw+/WDiuX+VzHTe
DYgIpdt8lzkOW5fIdr2VfqjkAX+6CGpA0z9Do1yW5ThYY0/ooMbWAg6+uL0S6JKr
gFOWtRZ4HJmAZKG61Dxax+2V7euSCTLre++gAVMVO9Ip3rgfrBMiNno8WdcFIhrs
v4JZL/4t25iCA3xCzWeq1UJH9Q4kxXaYe9eqlzWn3lvt6d2swwvOcCZN/XikFIpY
WKQdaTag1V6gGlYy7yxFQYUEPUoTnP+uI71D0tSSKfCjXZoEw4b3LiDPE7i6uwpa
Mlu4I7gR7Un929UZ7yACIxFqBTwk0BnZID4NG1Oea4g29RjS1ntVnlbHT1RB7BQw
4IvNye7K5CXNNpKxOoypfL6VRBW2RYjsBj0mU3hXqfWetN6UzBlZB/yUgUVeVRuk
wbcUOtW5CeHgnO6p57U2Jo7xgd7Y2RfqHlGzwYCcBKHp2alHNDTtAgUd6zmgyX6b
4x+ex2vhXByOEyY07bQoYnbQcYoyFqhXwHmaHRaXq6mk6VjYOHvWbewFlkbpjkyL
5oV5sRPVFBz9E1LTxtiE+NYzCSkIxyQslu+5OjMu4AAu4Pfm4D6mFKzBup0ugKNg
NZnUhErg4U7g6i8QHAK03jfaaYwAufGQ3IheSOD6UGrZ5NfkVi80EQW5kc3DAxVt
5pxicDX+TorvwEkAzY2QrnO9/1YDcKY4D6w/U0QxUF+mZ+VThyfDe6k7Nk7pqkPz
mCKQOfQj8UH9Z+JBf9H587krqYRB0B+8JROFxmGsio0s2xfD2QoUQwjkDnzjWTkw
laUwQw46q8ExiIvTrvc0JjhBLVjs+UWZ76dZcN9L1b35W9jYVr2dwM3UDAERUUQJ
Shc/yTAPLlHSw8pRUmWRwo3XOSJ6ZAcpmKWiPQ9KMiibfv8t4Sp1jEuHLU7JmB6p
940HpBt6+/F5GlCwla46jFJmkKPcc5f/uhHK5H7XUbw5VJBI/wZ1XDOsPLKntzaa
/BJCGbMLS+k2XByFJ/6aRwxmu4u6q6Cpu8XVgHYP4GXG59+zDgeOVeUuTqq7vZmv
cIapOg1sr8SKedb1MFvyjS+UtSForE3k7z4bTrV+gZ2MvBv3JlIErYsJsPZjd3Iv
G5qOOmWT8suboNYaHmUlpRu1jF+Fc9M4OVRXjGws4sgfnTEBhnvpEReb1cN21a0q
ubUKZUeZkhwY0pILs4ue1VgobE5y6UaY6bBVy4xT5GXy1pTiucdvPsRTI4Cw3Ngd
GtrLbnooLbVPsCywHChdF0fYfXX1MxcW+9yKNuyHxz8QbRu2f1gilqdCLV+3j6yW
S1ESdhkBeri8mxEnH65VjYSA2003Z5KBjylKji479ckGRdDzR3zC4Q52nt4yyW0n
Mj+TLj/4qnGkA8BbOHozfz6K30rSbLoe5fW38PmsHm47pBPvyidXKCAkbhwhGxhu
KLCjYmJ8cXe4dGFXIz7NpLWthaM+vxzGpA+JA8mXMw8ziB3Jfn9na2zesCc8q85f
WXF3Tsv4WwLliz0Eg11zUSXsbqNHCao3AGyrbWXqsZUcCzL17Z+H00y0FlPRS5E8
2Y+BMUo2UZDb/TzufhyX6BEVtbyT+pXY85CPcHxOoK1n6BZx6MTyPG+9dbTF7yHf
LseZBeyjxkD6Au2m0qVjkGJKZk+mGpxaf+P9WpTeUHU8dInju0L6smABUdR+CDkV
7zgDW25ANJihsZrSvdkfwWT9VT9HiDiCLfPjq8nNIt15PB5inJdrtdxy1CYnocU9
O6Ce5MnAKu2feoLNJSRTyPV7cgewFv6mLRXyG/slx25DV75vpHRVE/bst5+VXjW9
vJlLluE+zjF7ooNK73eFGOSy4ONq9Gq1LPCNPKalPIwWsy+2x/8N4RitvW8eiiW3
wflEbP9n6rBqgKIdUAXHOMI7JQ43ipcDLxQbF6402XAvc95gjTuz6t8G3XAN/TQ7
8/O6LXD2ht3BU3shDx76XbvQkyci25m5Gk1oo9OGgvv11FZsW9lYCBNLkRhIeTuE
iVe1+IVJIFyGJwCswXHPeQPzfidL2CPOaNzZG8VLSjBOPojqi43KZFIN01Yp2MXv
b9XA6mziu4FZpMTxnlJYq02ChfApGsUPnR5Jl6/pFW6C3MAimW4T8jYYGm0IaS8b
5dS5JPCb36oXBFjo79CCbOPO0Pnx04OAh++o4i+CaLUl2ASHFdDNjsjVrvGJaVjq
KmyC3Kt5euOIsjHfYdJCeJERdECRgJJwRAHzQZU3vXNbZd0dl8v9G8QLyZiOcXb6
WJHoc5ZNWuRl9uuCT3PtBfudj4L4NlVN6U2ZdNSceU6/SgSl8fIGlodiPQw3Iqpf
DuM5xwpBpwscvvCIR6D5l8Lk6M8gQ4eaLOrXn3brbf/MplN5RQsvkRLssWDU42v4
mj4PwZkN4lOjx+ny0Ao9kJhkFC4AbBr4SGzDaw/eCFtQ2/fEqyL1EmmFfZ5OpRzo
xHeYUk0Xb9gQVh00Zw9NkyDJsv/jiufbv2vkhxa63LrXabSt67NkloscElQMlbg1
FoDIffbqGFc6BkxzL+E48FujD0iOiP0eFfDi/B/G1GuKEGNtS4Wol+sVXmKbQnPw
5bCUp09XyN0xfeif82AFj8zcFxh8Pp4mGoydHFvBvqYfF8zUMMozgwtAyQfkTFVD
kp72veeLvymz3jZ+qRlZ9z8NVHN5c5MSVa5uP6LztLWa05ZadH8GRI+m4iEQXyYJ
LQVGCsofm2Anp/HeDVGx269mwm/euKu80FoTCCeed7iKmIfEZkEwcOpspD70cDcf
TyIk11ZzN1x0OY0wXkLFhghq4EXRfELDJu72FXIBrZcFPbwc8xKnX9uhYDHxb1Lv
SfZCKppEm1ZCZDjF461TEwPEWFbr4cH5GtuTp1WJOjE0nVVMuaRnD+bIkbO2dbNE
0nxifsDiUIKk1+/h3ZG85hW0ccHvSgPzXhgDAS1mZFKirNEK3fk4y0ATi1PSDM0J
OWOgKKD7b5d8EiG+9TstbccQtdJadYqaSRvuMRxREmtc//4IT+Zkj8D7lNO4cpoa
MMTmxqfI7+LS0UA8jMrcKNS0VvQUAOMMlCiwK+qGyZMBx8yAzZl7Hub4MYj6Em+W
hohN2tghzmTHwdwghkGxkQ+tsXQggmKCAkfPo6AWLKXk61ifLId4QYX3WipdUQZV
6QeezSfcO9oqT1tAv4MyMdiBUxiaLvXEZoMun462q1kokaD4L2UD+KKsg5vmTTMh
KM2bnbrttG6nBHJrAUtx6+pNNjMNOZbiW3RLdJEv816QOMEswV2jW6Qao5HNtfJ1
wbg4iIMOmN1ph854/Y+wg0tGVyiL8r8mg/c9HkzQ7O+o1JsQXivtpJfV8h1ByeZ8
xSQ44P+wT3XfoAIYg5GcwuSuXuf2FO/3ZbuovhsN9a1iVGu47HJs5Razctp+thL8
6xuBqeWc+LfCwA+Cg/lfsxF9AaRl9V06+kTP3vqCmLZLWF8vCHaTQLX2hbQn5b/B
J5jCmF8twO4zbvyEr5mErpiIXJYu1WSXyUIEjW7Cp3NH343pIWqkA+wMF41hBnMF
pdSwerUGuq6azyVzbCCZ6VKpaCsi45M2B+lqZxgii5Fj84hSo1KGLo+WPja091uq
aFzXZLhHWoa97lFcjy29Lo8x9ZuvF45L6scdRGDPd3alaxEx+oWZNELc4KSIZgfU
0fOQLDITHF0boQw+zN6q2rG/nVsCs6eoxumIPxsohMTM/bLVxcrKAIDA1yk7DfVX
ZUm3sXoX8xeLwivioegR5ltojxN31TR5+3N9ONdgqX9q8UGACxtH0Hq4JIJIzE5w
ah6ntaoI/MaW9kpK8OKxc3U0HxDH/ZfxU+SgFRqsV8FwWLkG5JrVrhJRxO7g/RRz
IWX3oe0uVeEyw+0p8OAgjk2w96IzoIu/YWec4Ou/z7OcKa2Rhrk2GqSvu9h64tlW
04kHQSa+tCpdfDepxHoKPizfnifyRTKU0zMTEmY2ykZ7761LZ4El2o0Dpk9pGjf0
Zy1hAAsMAj7Nl9VZtH5HhkKSFFrarE9C2nxVNljtEzMjnVa/HomEZH/ovc7GuEAa
g9Y5CLAzTsjEUiCEiWFbDK0rQ46GA8JfENtcplFIMSVO7/UK2IJzz0BNYlvbaNXC
+MZk2IeGDEy4g5+2xOgbN3v3N3zcCQhs+YavzRN/l2lI39mQPiO26WhxYsajsIJy
5PAg4Rb1DCeMhznN5UrNnHgE0dtVwWED8F/fYGoOrDmCijCJN53mahOaMVS+Q5wv
I/gaCvf//wWGn4KVIfegf0/ti3RJaucyJtTKFvItZjNp6r37/Ei0S/sC/XYgPQ3A
ISUBdyN1QN6HGACfs/Yei53wqzxqR9jnFYvovtetZicbiiDunwLqbUfY0QlhDynH
4e/gdNqycw1DDc/d22afF4m9j7gkYE0Z+rF1TK6QWAVY2VIuljnAPUx4C6x1tz4c
24/ws3dbpqiSMjtImeNhb1MCtmeXEf4ADV4tly9FWpv93+Uh3GLpqRJs6tv6lvt2
8b7peU3RnIfkupg09MXm0Bezt7mjX0RL9c8cjuVinBnWDhpx7GbISEu4P6yJaFbf
kX/umniEY591YljIJLiO7fautEmX92L/QGeUnRBtq29JYDrVu/EVJgHYotsuRCWm
y8mWwY1tB1A86mNfrJms4K9jsdG3pIPVQt3ii1O4+qwDcKMitGPGMq/XSA2ZCI4a
twZRaZ9K3lYWUW/IDrT0WtmVgLaVWw3jx1l0VGwjCuzA5AIsEq7sYWmY5C8WARRQ
RitbZPmwyOk9U+H4BBAoXDl+tBZPb6way/8joB7TMEmjDBtEURcR1n0sQk1yy2yD
DzoP/lVC1D78IhNsa5fKqmGb4LjyZ3t4+yih6KoCuputdmZmVJkvB+8JoctiOX+g
Bxy55uDcUZkmzs/6mpwlCmLqIYLK+YDADgQRvigMXj7IFHx9T1gGe1huMLTchXuT
/s3afuXh9+pLZmCZRtpLWziDupJWQ0siS3IMyE9eG7yRuTJ3MFDCyw+jrypV6ZFw
N7j6ux+L0t46u7C+hcwcHYK59yodR0Y8jVa1b0xERC2HR4LkreunjP/se30Rl0JV
MqifHaf4eMDTpWm6fz8HlXqrPGFBtvSPJkfzWyyazpOGWiyRn0ZWaZN1P6Gu1rs5
lISDYGG/2nwkNn7IeXN/eh+kxzj7QFVXnfKVupd9jTSQBVhocHO5V4en9nCFP7H1
PUvI6BN3MaMpk2M9yzWIWHiD1PoJtla+4IuBJOYARfkOUEvo1nqI2VuRpeVaB/1q
PJUKdzcuuvXxbbWra/cRohvzf58aGqcUdX/+j3aCntiFnwwhD9oO0Ag/YfcoPJUj
M59g1bCgeUDgDUS39dyLUPEggtRhL3V+ZOeqxubaqqjzJOI6fJj1JSZfBcn1f9Fi
eXM6VtzppAvHgq03i/oWZD7GcEmDQd36uXIIh1U1nB27mil0U1bDrdZTP0Nr9J3B
Hc3ZrhCQuD7AtE/1bybAzWC/mR/Wkt84TgB5RjBWS5Aib41re0T8nkgSAhFoEgFO
b2eNBDPFMF2I5LwEkwZgo5jzBLV6uRlPOsy+Oljph0+/aJWxuC/C6+rFPm2LZY6/
vHe/+/drFPTZX2v63DRmRAZfQev+vcwfMpZcO6JGGPuyZmdTmzp0K9ZrOL86of9a
xsH/AmNU6XMutYbGHnw3VFffjJapmkS9fF3ba0X1PBU9BPxyOuuG4De1HWOULgen
lmvXMw/9+S0Tob/pu0KSwiQmEJg5tyBFWbbgXbxWMNICqP2w0XkAI/qWxmee9Fuc
b9M6qvUjmq6izGCYaCY9v1/Zz4cUQLdnNqDgZri+SR6rI+TX2Ss0EiqXoTRgFN5t
zFeIwmOHQd/0kYJkvcG8YSy7UFNKfkX/W9aQb49k3Maj0La3nS3AvVqewVdzeWba
d3Re1DKSzNXg+xgv9dP6KLSQoku1qZMp4ew38N6VE/dpkL4AV8qKQx2QDzm5QyrG
jbMVmf8g9EELnjofvLGila9IPUHdrxZyu+ET1oaE6pPOuTHRZREZyiOR7m9lZTin
VicWtwwU1ZEtxIQzNqhIoKExQpnT8qSYDiS9HKiMbTic6SUODCp8Ul+2NSN3lnki
FWz42F1p5UHLFlVaDGDQbvvnv7yjGmXuWYoK+Fx6YMAnS1p1w+JR8lzJhc14eMjd
O1TUE8ClynECdO9Cx4MCs732ILq9ZjKa3Fy3ClRwrhfFh7Tg7qAoGbSeb/w5y7Kk
WFT5cgqZn2o/9IitwkQehBA0uKNuFznyIomJnFfMHN0H7JDcesblYtZzxacEyPqb
1sBM0h4TbiO9SMYLs9Z04N6ltq4KMnZaJz2pctS2R2rc1VVmEbPpYyH6VfpU3Pcq
dhSz7ChaZ9RrLGkP+yZ9HlI3mVcqiYFkbRugVXTiKCXaIHWuQuTLCDZmmECpxIKR
1lKh+Yge1s1XNuOLKUl6mxZ851vx/+sAVnxrEF4wtl9GCe0JiFHtmKl5t+Nxup/k
ruHLE+ctsv5UZ21u9rM0Z7mgEtxmgwR22uFDvmtsZHrZUPtoMxpNYffYmXF0AICY
E2ef96ACoOiyCWEZQ0e/UBpMK8uXbreHt39SR8LH9AM1RwX1ixBwoZx04Z/6hPnu
aaKWF16vUMUHAR0MNWWnovQqU1KLGpekb7myr6XMHQZ0B1mBgeCrCFKVU0YfXIh5
Dg+d07jWzVhaAoPI1DPC77D8OZbnvqQC0EjWnH/lWaDDgj4uY/5nsg1f0WXco0Bz
sQ0NMDXyK/RgDzY4pJ1Y1jqeHjsCqlO7PoLNLyl89wiGjlaTMW/wbJOtxtH6lmIX
FGZ8ydj2imh6fwvWk5kgzQJtoSwI42XGGDN/+k/BLkiHT/A2RyCeabW/1jvaBDwf
XRewbW7PZJOc7CmQgQ+uguSLYiI862HXhdzzMGsEUCrsXSCa5ZdRqWn/OmC0Tz4j
upFZImhUCt9dCgnRaa8ZSLRnzOqoS4jO4j6hnhHuHjWLE/py0RaNkt+defYDXWfU
PknIoVsu1UYEEBrvdl9xONGs4UWS5/TyjQp8QKPs13srzKDgZ/ItCSCIsTaS2ZjK
cjcGSCAMleZT32mQRZmM+q5N6hYFOkQZdyrOj1l9UfCYbIbv7czvMw7eUQqyAPEk
hSpAJB6OYNrZozQJS5ZyJSufMjS3wETDX1MryNQdzNLr0VUpdfTTPp1A9ixAXj6h
cnah76/YIjYO2S94J3wrlW+uF6w82G0Ag22Stv/K4+YrFlyfaXzP1YUly8Wk6eMf
dEb4qkf4JblYH9PuStkWyiopCFpGq5VlJE93/i9vUfOem12TNEtIWUgZgBIj1JOv
CyqY2IVN6iseQtKVmICSE1qQGhGmLYHIXateyBfTEqI4xMahs3Nwx8Buk4YNXKCv
j2QeB3nP29+dPGSTf8pdwFLJGgkRi04FE6g82hKfrygg6exFfvTewPqBZOXhKfow
bw9CRNFHOcyWyIvj9sugZI05kLvYcciLnHlxDGftsJopZtMMVKENRDi758Dmb6C5
dyCw4R+P0IyVripWgnBVJI0qH2AkrAa2sC75d07xA6NUIlS8S4KIoNn7Czihw32Z
bir0xI1xPN7zH/Lq1p3Insj0F3/TzLEmdTmJVFp4jVBxDlPCWhMDaR9cOaRJY1A1
wVe9z04FE1fUQ/envCf97eqTh7ivxDHlQkp+jIBOP8gNykYalagXQrxl/y9YoRpI
NqdhSm1y7xZwWQgI3/ZjmqgX3bvrwhsybg5L2TIwpoCgVT9kLpuTir7gXNKT33ef
XY+8p22kaOrhBurHPgGfXBKmFeR337p3qBDbVRQRNqNcw/WSv+SQHWAv3goIy0jf
SyhHGLxkj/KiWpyGHctJFrs8eKXrKpJfGe/QyDbsE9kFxmpgMOTl4dtduYpN4fzk
HBpJgjmJPXubgKPHvPFT8Yq+ezRgtzNMyG/6LtgcWWkOE1oAhBedidOzCbf3Da5U
MtreFAZgeqLo37okCp3FeJmNDXyeJgRx1dq34AxY3fS4GTcEUxZQnK0vn1EMPxNK
cXtjntUnm+I5krek8MIF2HKy5uf4cY7LjAWMlFDKVOZLcpl/t4YJQ0a4wJj77/c5
Yc5U7321NbrAvxC/gXqm/158bcbLI1LblE8RDlY6eyLuhil3ZY53fpNclq8NMRe4
dCchvqhsqDk1oCFomX7zSUj2DiL0vcCbzBpdjdK5yI2+/uzV7t9EA8u6hU1sbt/C
JPkaTH24P7I4WRQG6vrdrSHcnjNk74/YtNUnu1O9XdK2OHnUUS9+ENwFVqlLvHor
6bL1l9Z+fb18AG4a3NAnAd2DI2yg20gwhDMw8VDk6pm6HbfD6NL1DPPHdW82qLPs
ie9dcPMbDdonNpn+L5OoM4p/hgk/wiTDi7aq4icYwj4mYFBcrUkIB49sJOA1gNdh
s9r0/MJMSG9Y8PeTC7B9QtVrxKjiq7+qwaySHPrH42C8fW+SzqQsAERv1k36qbf9
4yyrEGOXOGzEMg6mRA/wuixYLtzeX22rB2dVSFj2TcbpyzkH5vTFMcRD1rZF4pzT
1Xm8BjAJXk5SEXSgChGYbgrDod+u0r4aD87psnoW/lcDCcxBNcJk8qVRDM5JuoqF
iwx2YXKM2DxCRLph2xH7Pe/V7BOsUX2/nBa4FVV0nXBUSfpmQPB0r4hvmAPgLNgo
t3UJ7u51ZNNu2tnsrnVPV8p2SvLlZuUwO3rNVQxZWyFjJjnNDW957PVoHc2xGEWE
EclWDLF95rkeqrWcYJapE3EOUafIybsmd3RvndMXHReBhdc3HHfMMscdXRkHhiWi
USPcnM4dkg6Voau1ivjPvAXZXVz9hgCZMPAtZDW5xWuNm8/PPyn+/pc+Kt6KHeZG
QjBaAmubDmzYsQ/ROWfti6lwqJy9ZzN8oc/36T+ctngFgMidr/PejSc0zveTdV2W
Qr/Ke9W6Ma68X4RSP+M98XChdAh7f3223t2sqVNMLBNA2jLIG3Uc2ZIxtkUAWiS0
5CUaI02aDCXkccP+iofLxCiWvLsXnc6kNJzQCaZIBZu3eOoSATZHVFeasHX9oTBo
09R9RO9uF6pVGa78x5S18JQ9n83EoPgM3cddPtSbyhJC1V5mZPGQSgkThxByIgn3
fWT+s4Q1LlhozCwjydwpEK+3yFfEw2zDpvukKgz+y8mjsNPYYy/GRYcWy8aEplCv
uUjfkLELEpzxaaeUGnGtOJeS0uXPUW+YkhsgwULpWpt1FzOluul2XSh6ERB+2UKP
2kJkqAwnIpXfZqWNix7dOpIfv9FZfZNjKWQM3foICIIi4zJKk2ffZtpjxEGMlXeC
zdM65ViCRfNrB2qg9uBLgr5TwUVy1lUOwzCmnIxR1LhN1GAjLe4cX2ZFMY/IrAN0
v8Rp24BMjEFVoh6F0KpEfMy7JjkqBp4y6YpegYg/fr8Z3Y+pB45d2sycdH/ouaoM
YPOMvPkEC+c3/NSCw9B58lh/l9IODRgXjUbiGRkEbiPeu7NKE40OVMKkDShX3ws0
uSwvvYk5NIXI8Yf55MWczjmbQLx097XWeeMVuUfIxJYQQyqiDA+zI3c+Hv25wS1y
+PFUKFmXHj8xzjPIxZwMMYn5qxQq2Djh2e4WVVdylEvnRlp3VoN5YvVzeasnAZUR
K5r+Csr86nfJmuTZVHikrK9d1cq9KXYCK75DsCZ4LJ2iJXtZ10R1eZ0HS6dL8TAv
ntol5uKxUTZgVVUKuudmUf0zClO7LiPLhS5bRBadMGhOr3HYYad0XCkcn6eV2A4M
IKlUH9ZrmKh4+7MStWOVRw50t16WddN8NmLaM/1pqeFDQpDaGcVG9mYxT3dnDiiZ
In4vyFzBZU+sg9iUs/onNfMhrHtVVAU6P+l01udg0WdB0QlcT4/Mn1tULTcyJWjh
J9H3/LineLvuJ2x44OhYzT/8T2iyiBaNuqRg5wD5xJg1DGIw+/uIeuK1Bgsj1+tB
4LbnG34F9HJHz/gdKZnhRpXuPQQOV/9QIkt70pzhtGA8241Y0HwU86g9yU3F5Lm5
TpP1NOu7f8PxDQrfrOxFHZwIvvGU+153gKAahZ9ZG8t/57R2jk29XztFsKi3bN2R
3uGfoeCLmDshrEzPZpxyXKsDdqyadqS3IoTALsaktIwaHMaS8yovdbxhw7E3KinV
ZgMjG7jBwdIvl7sKaAWMWCKVsv3vQHCHCCi/BJo7oPh71J1vs9QU9fVnbebcPVJv
fvNWj8f5dS3v2zbD1kywdF7rHQSaQMibGE3xQ9xhCWWXdscyhXnVGzD+9jFGLcuw
cWF4blLMAi7YIbTSRcGO2iNUcW1Iobgbvbdmfe9s7ev03ho5YX8o3a/5zz1Sv5tT
+I/nz6W9geBlZNBQd6EkSYRq3aNay4RYcb2cX0FGFbQGAfuwvuK7wKd0admzSzIu
fNivy8Um1q6Jf+OcfkU9DbUfYuGGVLXOHHLxF50gHQ+ZxTxRzW4VOCfyny1fROz9
N5Nlu9o+Wgs8fvZZmKyKO8ynB5JA4uQQR5Yu9dfgI9e035yIlPZ9HwMHDGnt64bs
w0fgqYlLjogJQ4I7G6sL15M0dOP/UNvR67luqdd9Xle91nQhODRF1nDiMVYqqik+
y92KFncgXqf1ggeK+Bx1g6bGSko+xZ1Pr5RtGd6cF00qxpDgJXtxL/BDTMFS7RsV
oX1O83P4z5ak99SWXCoPuLddhEX00YNW9RBunZT+y1vGN9oKkbvtg3cLGwV223Ai
xkD+GHcA0zSkqdZwudz2FudD1JA+nCKBsxWYI4idFPKPcniiamFIQCKV0e/81E/Q
HKOLO6QnZznzs1rVPztzQnRrT5iUIpC4MiiWOxOQfw0MG8qWetRVgDmOTwhwPShd
oCDCSepD6avVgafBs1VdO+LPCOrWycGwI25NirvEUku6txVVghOGIAvTKSCqd/w7
p98IZpl2+mecDdY9wcdvcgdHhPys5OufxYrypCUBS8hYg+2A90FMF3o9xHYbnX8N
WLU2goIpsrItbWd2gt7V5pmw/t60fAD1E6xH/aCFKdqXUHQkWSZKG/aVhNKcxsQl
JVvQCR1suS8b6cjynl48E3o2d9WpRkYQhWAeuPGtR1acEOXPJDUbFrY50/O+YZRW
5ImdPC30cAKCVAGYI1PiW68iA7w8ul4d6XJuS9rszDv8nN6WOaQJVS7SziiFKj23
BsEEEznfLV7rw4GG+wXVXYDqw8GbWFXJ9/X2yJ1HGWccAcADRpAtMIs+3q1wQ+qh
n223wUUb6Wa433JEDRGpHG6U2B+hol+WjK82fauWn+HSNdz1dpClxZnZldOpif9A
OHCUitIgiykTmwmyLFO1KFBiF0Q1kmOUT4vat7/odj49hv9laEXduLm4eZWSJxh3
TY1v+L6qtJldXcTrsEGeMjryIZ39XsAtwYLiPv/pIL8BkIh+fTR8tAK9UUtLUTnG
EtzkFKdCZs6ibAmoN1h1Vgegoy3nRIzvhwfDZ1qsrk49T0U47uZwJLlAA0JGlSg+
ea5RncvwhRiOdy3c9TMWs/kLCiTDgeHu9nLePqbCNMD12x9ODWt8I2gbIXPtDGkr
bgshLUXPKXjYtzyE9qE25N6uVpcXIacbtRlAkKSi5Fwn3FLcf/gWJmIJ1XQeuQTO
U9a2rVW4vHhAS6IGYm+kEiEoOK6VZk9VJ1fMfKxQP10zaJUyyr15LaGEQwCckwYE
iHE1eIv4ESNdB5FfsEBhcPE3Zmf8HzWf9zeiPYm7ajWTkAlowm2IN0hel9WxwsRq
0sVLQIo2EnM6/SwgPacJDjidDgvi2rFZNhOuZdg3Xxv7rC7xVtNVhWJX6IEECNvL
aMli9mU6nruHsq1zptEViiJnOgwM/M3ZvEZFVZd8yPv4EStETsdRQrkE1aqP0b5x
GjZtLOGq4Wvw4A+rvTN/074MwVzSZcMosOOvi+xVEUfFk3taKrYF2uyAXT2CaCD7
92hUvtMueLg4EhyJebB9BRca57BqedABAj18LwYjQ9thZGw7Wd0NDwWxpTrgmDSi
az4SmL+SYwbpcSdxG4n2ehc74TjbpSJtgodc1W8NMnblKfm0r8o5hPb/1Hk6EUPS
6TOOPYNsuySpStulmCT07V++/c+vjIUQEbdcLw4tvwe1pJ0Rj+oEsowY91OEmS/j
eU1zePlwuUnE8df4uBkJ0+6VCEgEdj+9+3HR5h0BP9d+zgkzWjB4jyRNAixoWWtn
hbA6mpGKKQlJf42QZLuJUxSHN6mWmBrrbnKMMWyOcVejmM8Psv/Pd5x6bUnWXBOP
EO7RjHySVlIUjf0CTeYGPQ9MqVYbTPLbdCQPYNIxUobKCj91mSKLS/2yuxgEB9eX
tLWkBrAYBYIy2hT53LuwLZpJKoijhKSYebrZ1PGf6855gtptSACfcBCOMqkWYxYp
A1BkKZ7WsMACeU8Uf9sBXGwt//t0tBuFG1yZdRA/Q8VsjDiQNIXz+iZXC4Fc6bZD
qHztwjjwo0F850RZMYTpJMWqag2Oe91HXZZQL9w8w2FZ3jyCntW20WnqMM2rcc6T
l8NMwOM07+0kAq/t8L+OllmgkQtqlN2DbqOyHJal9y/YH/FkEI7ezxO3BlqiQlU2
gIiQjXdj+3uFYO84ZzuFvGti7s0v+1GDXQmAfSImU6zk7+3yfz68DyyUmJH15RVx
wAb5DGCeg+2LvRKMRL/jjpY5e0muM8g2mfu6MyWe/WLpdiRUmSpjt2LUWuxXPyAA
iDzBMMoDvytJp9JaxgLSGQo84WzxFzQ5pIXM278QdPPkxKP2iBTVPSLdyE/LdBa8
gPTvvPTaMsOHaqXhdxlfKHc7ZRx71BOJH5Mibv2+Mk2Yk/mFEIk7uSGweFmmlvWn
KJtFoU0tKGV5DEX387y5xYiU0zdZZ+AaBjaJpc2y6THeL7zcR53lICYeCOJnpG0g
7sYAZMk8eUvvZ4gWkO0Njn6fqkL68z2tVvZw6fTNwbdCYxz2MOA5LDcg8yhsIbI+
HcGsMBWq3ysEsj/1PZ3LIwRuxDX9WaJrfIWorKNTfgSofymI5xAp5IDkU1bTPvtG
LKq2GPLsfLXRytTLuYONlbQk0aLcu2X6GzVVuHvabsjETHKsmhADdDIexK95gL8S
bUgT5YZTxCqpNCkpiikzTH91WctiAx8DKV32YfBhHxixzOPp78jag0tnpjhZhQYR
3xtMuzMEuuzCyiXDRy7qXlDCWQyorKMq30wyswyJEhh7FGdtaOY2retjSLoyOzb2
CpK/MNI65v6bQDLZvdup8BEEtbKrKpOAI+B18AZFmKd2OgSuKwItTqxo5z5jUPO4
YpoP7WlDvaonLKyPjdJiW/l5trEWSW9/OwAjd1OPc1XMyfe5DCltf9M7Pw0CQ1ML
lyEcuBuEWaT3BsPeFdRq75BPeU7RNE2xqUZm9RL1Lne8of6aj239mlKE1+7YN7gK
x/NshmtKFB55BEgxVQdZxWlMlIf3nhslXpNUzkRUsdHr8zaY6QvdgRWJt5J2Erkd
lODE9XwXAZzRZXJ8MSNv69I30UPCm0GVtu3tI3OuKBzysnhrYNpb9csdB4fx+ksm
6WTztIFd/ds+O1gK2vaJD1imSVCnZdAW+E4YdwXh7oCNYCp98YHlJ5VHUmKhs53o
SRW/Ui0teIW4TQMpp+ra+0pLNTtzYG/X5QnrcGAGa5KXv7I9fdaDOHaNXTvb3mOG
kL+PYUQRi3Ruv21TbbyqmU5aGhAGIGn5P9TDrFRySruQ3yP4mHdOYwy+vajRCqi6
+NEXn5vQ8y3o+q8Gznu5Pvq6vjyEkMpLV5G8X1Xunk8m+NZWOOHkhuXePegdJYAG
3p8BwY7nvTUgV7G+UdCpH1Q9sPT4arsh+S1r0Wdu41X4Bci/Yz8WfPKFtV6GFMWN
RY/Z9sNuKAfCn2kq21/6O4ftLWsjfCOfuKcVdPRf1o5ausNyEhMfZTXJaUiRnAaD
Zim7tB1QiKO4UKzyZGsZirEbUpSzj3zaHUrlfwrDNVp5f0dRfrtIavFItG+JCM5A
B2i0yStiyJx45YJOukji1s4t4UDrVQ+X2glaKIs8Sf4DCxQDRVCejfAyryKAeQaH
GockQ0b7LeQeYNXkT4YwSWM5H7R3DoumypLzTssrS0Jz6nuzwxb3UK5Wn6ng6qdE
tGgbct0l9qdAjp7T3qav9YHnIAMCEX84IqK9+Dye6VMJH3iFc9R0oXiIxXxV4v/N
nf/Uum0mjnXdkyrYkMMZ8BBNJCVr9F1lbDztto6NV2Fi31kQIGuI45fsjSxzQgVc
zMFC8XGD9eF3GK4u2iN1kYpftWh/pT6O1wFWsQ8nbxYZACgAf6yUHDb2xsaqRELr
sHMz7JsYBMHG7BuAfEL3XVWp3+Y3S4kQV5BJTbyJAR+yY4inUWOcSgChnHvtHEBl
cfJrue/ZSoARzb2FCXBl/ibnUo0dvrZ7q5zDiHuVaRkRVRMriuOydR4+HteUHYk7
xSWWJm0SEJo+oXiYB2Cc1e883gI7ctUCJEglLYVN3Wk+SoGcIcfSHmXyxHinhbfs
LJIlK5s2aYnPIsmbQVQ8aA9ZKt1ZCzmTHu7TMGYZ79HVF6xiIbMnsiompLEmIV5E
GUp1wTPzZNOYGWmJzYGFlciDNB/vKFxWiPQwqWhEiOmFouPUDZxXXbhdJOhB6U2K
B1s2Kf+beeW6QYkPFpBCtm5tjkwF3jAVuL14RbvpOrMmI+bo4b1OcZznzaVVNCXp
Eesn7G0WMeuDJlqBAHJkNIIBmiOGIcplGttzZ6h9zrMCnCicJOmuZhWsvkGvW3Xx
vBCBRy8qB5HomlOP7vQXWByO6e6eHZUpRBSZj0H+j7PknY3dvlqMvAWUdp3y+jHY
nGFOOYjjtwW8kmENubpXpo2j8B5d/6iQdB7COPmiI2RXLu9EbgKuMi69ORgq5WiZ
THd6ilihf9p7hmvJgeen92FYSUD/iXenDWyOHEmg9ZPg8ULjZBCVM2LYW0Qb9G0p
IO2CoFvckdYKcXh/VtigBDDXyBXdkWNRYPCYpoggHosNFw2ZmRlcaZrbtNxaB3Ty
6Y1EPtF5yrItlkVEDFksgO7p6k/7/7hnbqlItG9cQj4sBiVRr/XZgu9jcJ4X0psr
8ladqN7SDht6Hvd0BwoM20b3mR8mFYeB9kI5gemvOew4clhjWCE4wd9644H+A8yP
K3OJIgv/Rfp8+UIgwRWuvIoANwEq38t3r33SghqE6qI2XMpvU3AG4Vvh/2hLckwP
aXyN88T+ORLavoiOS7Pq1I+oAfwKdojO4nTqx8pT2PYVqD+IzRbkRuYFHFAWp4zE
jN2iq699yfgXSPtODcuLIMv44BshUE57NLeUBEWVgrM65rVU7VGCwKTSJOWR5pTF
OH3UX7AFBXdkYrDt5Pn8fEKD988THve/FuFrKOwD1b4kKkF/ElabNnwMDtNq7L6R
nK5xGSRG/7Np4QgYQHcny4dqjIEtxteSG9mCSQDtBlmPv3K6C4TEekKZrnffMBPr
TCd2u0jteYb94/dpMWdoDFBz3Ospbbrsoav4zuNu88sJ0Vfxyi32ZWJUE4bSWQZ7
Of4g+E+CcHwFpYHSwbScJgc2VJeUOCdGtROq1QZLVTyeACNeN9FT6dwE9Ri8fOEm
7t7VBXBV6DB4PT6hyFFMCBGU0G2rRhVroqfe7l4kvGKNjOFxtS0Q8O6KVoORtkaA
PHWUQLA9gfBvwVY1H1A/vqiyIdddEcc5Ay5qWZraZvusSCo0mhIJ0I2f2r8aLLVK
cCRB0nd4ULu6VNL+ZTBncjm1gx3+mbJwDJyKSzaMf47LQfHsNsxAdGs+Zj24Mcd6
KOyky7+hmEH9HN6NgDokPQsprP1eecYESt9BgJcM/ylqo3HdqytoHD8qkNJ+rzYf
6b3viSKTKtpJb5fdOH1hwWtZU3jWYppO4H7VQeJ4WwCvCHlSrqFkdqSXaWhhQYxt
qM45setje9/7h1TE/heDuyuCd9WHuGIAJETyJuIyjD+re0fwEZglISy3Q8uLXbmr
BCRLDlpZ0gJi1x4ZHId6YVbBb+DC2j6o/wlFSFai6/S19WaELYY7hOZl+5jx+LI0
uWCWnDTMRPkqAD8Q/aq4Wp65l4tnVaDbBd49+8tLKbtGBku9o54nNo+QiiVim5mc
9C+/qRsj+6KXP/4qGi8q4B2EQoYil/OlkVs9lyIdgCbJ3r82dB6Wr23GXqu5zlXU
POcdYwncZBygVbc42Pej5kTUjwwEp0gXwCp38L52aHPBMasO2F/SUMF9mkZ5heLs
OjKK4FRZUJ56WsazEy+UdmR2XPCDweejBer6z2Eq+Y14PrNWMHvBsHyWK8SSqT2R
chi1A6c68kE3oDbc5NNigMb/wd/KlExIgZK+44iYtzizRI2hupnnkYwEINwUeTlS
g43wYwqpWJDuC89lFxSekybqvgaiXLIDYmlnDsCx/ih3ef7wdb9mrTfXLefDHh8+
JGTGiYzMA1PTGVcXOAQqt0wY4abP4Edl8jVsjHJXmTH7fqM7fvdiDZcCF7BFVKH/
ylayra90mcsb95yT1SUd0iNwzb1KfyWOpd5JdP1Ka6cFgDq6DO5cxcM6CkugbzDi
wIR7jO5p7HxrJ1tCqmBylKWvD0JhXphlVn/gUXtXHVRg7ppCfsSJAIO4hxzOb5dd
03HeRqTnnMe9WNrU9J1DiY4uwj5t1/Btpii83ZU8Nw7UbS7Hs59UkSbdxpumZDp4
KdIM6vq+l+5bx3N4k6LAoFq2+Nagi1/UPGJAiXhM2otJvShp9igE9+Hpjfj0BbUw
IpZzpNGmGPoRRT3mk32//T7rp7WpHfyaNZP7J/u3WXaIIU9mCw0DHjXBMBotrWtR
PkqAoktWdGpW/e/YRx6Qv1KIpsdYeoQ1Viw3NHKSeuGESjOjHds4GqR8xBxanVhg
s2XC/DrJqxwquCZfTTtdDvrc4kzrtxb0KVP4TyoXq1bqneQ3i5eJK/0KbVejLgUZ
3YGUcWkKE9fV+ZnrQMW+0hqa8CGIVIblSRCcICDkVPqDSNNrkTJCgHs/qXaTc+6u
QP/ffnD57jH47NIUy3rAuLTlfv1JoPpIZRhzaasiiUcZpmgdLGgo/kE/+w3adg+K
sN1iNxX+WPfZv/4KXZbdvkTzHDQuqiBs1UVm5CzY1DrFOaIaebbY2qIJ5OhSTRqC
kjlAfaYTY9oFwhzI3KnXhYZQRIoaI2nmepGL23720IrDxuezLTPmxBs8V/+cPk3W
170XoUjHxw6xtYlIbDsedHQYKIcPxe+85QvfyzubWmUJPEs7TjPM42NHokJr90fc
9vAzvAfyS9EVsZzLmj2K2iO5sKQWD0p/6SIiUBEue2AH03kJN5EguTkckTxpZpMv
k8/ZPrVTy3uD7TAUXnFB0BSmHRos8khMtPDEzyZg+RBnKNHHyYOoNk/pXW3RRZRZ
5PMLSA1Z9RWupf/lEwjISs8Q4eZrnoIoQ4ok/8H5ksZ+C5TBcZWA52o06NAC3Pd8
NNTu7KxlOjj6fCXrz7H0u6CwCIPJhwRM2B12CaUwPTfoT5zDhoJcQRf2EQKb9y3y
KM1oo39f1Lv3bzk4Af/WUUkPU6OwLYLQVxjaj2R8s1J4rIr10O/Yp70JqHg6UPYW
96+M6i4akDsLlF7B3TapvydWw9+ie4LA337pOUtZWkl+g0WXKMErJW2xqyHb4m0W
CBNqRpbaz3jP2Ex28T0hgUiiLFnviPpRf0U+3ueYqmE6L0eGeiEZch808mMrJgnS
0btlg6pghTnH0QlKD9D/yS4uwAhbq6pKHzBkxL+pfR/EgHpWL8X3g6BiYgrPO3hd
XxIp96HH4KvgUaR2ULpEUVfbwNrzi+nrSXlvwaOTh5dyARp/gQ1GE2GZOf1HHK5T
UqwsFTdskaT/SJcIvw5kv8qTJz1hMYQi+zt9jixefbAi3WNxDjKVPjiuyt7vznxY
W4fqahsFXWOJAg+aBkY+//ujhXjNRw1PvsWSz+yyWl+jPe2Ts72jdg+pVTxr5Je3
We+CZ/ZxqYzTnhI66t0qRdssAQgdo7qLTxZl4iJ7ph/CtAEb25oBazVg/rHjqcGn
irjAn1Ztfa4rWiSxUJBEVcvnhSHua/huO08KFtvAalnAq8aH2WF14yAuNqVvsZcv
EUBcSzbP1LbhiUeO9f1oQvI/buSSf6bJcKfpplMouUOtHcjk3m4f/HNMvlaFPZcp
XrmWDv1JkCIduPEIKCponU4BLEiixBXNmEjVRjVZjhONy1rffhrjI/HqoJDw7yoL
dG3Dq181Q36k4WIqPpXbnbKi4d6zMbNi7hz2Jwz6e9TSTuMIjYX+7cXgoGW3exLr
D8eBRTErbD8/n4qD9p//CQoHcDD+YPAokCtoqe66k6YbRWIXFhexvPgW/vT69LCt
uqHP8RLIqQ6viIZCNhhYe+dPCPGBGOFmVwR3lbl7j4S9dWQS+d4qCxIaX/gjKtcv
sqFMPyYODL23+zp971doAC8u8GkVmWbXEL2yQx+ml6EgAgP0Fa5HJ1fNvW5AoKWh
/mNx6O8MGMM2aFm8zWvLkkrQj2zufq+htxSm4xCsVW4lOSeVC4LYl5ECSm+TBjkx
upRErdlWdnS2MpZWNRmEbD0JS3KqlA7/VkA3svljzRdyTloRsRszbJEU2SP3fwdQ
sYnfs/Tgei1wOg6DsVLILg9bNtHYlFcMzb/WIvbnXhHjg1sl3Sg5fspF+OQIXunt
WoWZlDbjcXGGm/z5KZJ7MIr1zKLrsgiZKc+GWuFKOrPKjGdP/3Fu+G6iAmD2HDV8
trOfKDBIfACxMxKanl5P84tFMsVwXwqxr4z7GzuFtBKrsIHSKAVz7P0gCa1Men0M
DmjpSs0fQprr3OHBiksxZUDOlxfhUfNkETDR08JUMlkXwCu2bqTsK9i9wxEJCKmz
N/8HafRhTbuhYLWZ1hlLC0cgNq4KH/hq9+qUddfR/+m62H449v4GvlUKE43lOBdW
a/h1nZL4Kk7A0wPjqPVeL7RHj61wHlB2lt/MMdWlxhUvmH/Sqra4I7t9EbEtc7Ug
sHb0kraCa99lD4okbfgt8w45vb1u6CmcDQgCBxRd1QrxDgRZheXzstNQcHDKIkGw
El07rUREWU/tL5vZ3CjAcRRcRV8TVUPLLBmkLIbVGg+3MkZ5OFeQMQso8WoE/0JT
VggQpY+ChAPc9fUpsjVVa5QHxkA+RVSYhpC9gakWKpQkX/GIbK3sTW/heoV1v/m2
BFeVeuvqXPkNLiuMsO7yjeskYTCKdui8/OjtuO529Jk70/H/QUx17IkcDg9lp63G
rSoFIJMaKkKqAkr5MjCK/HUwYUBIqTLmHeulcmUwqB+aIvosRmYmcqqr+SjxGr55
V9Cm6IvoKwgj0UhoWgLeWoEfEVLQUpcLzC06aBI8KfBxUANOIBgJ5KqTw5OHlqYr
0oTHHaTCCzPODiYB+GbiKF976C2qMJra+vaEsSpvQYd5+Qqh9WwYYTDMsgHaHsbX
PHooOPa4tu4NcRMOZNQhkqOFY+SMlB8/k3JQjGlW+NhpKTS9uBimNbTKoSqc2CLL
D9yVL9VHriuHJhm3BWghs8lSZP0+ODgauHjpXJISolQPTxoYOykkRfg4yB8LAEOM
eQt1kVTSxazhvlx696tiAw32Pq/g6mnnPzhVD+G8Xq906bG6Ak+ofOvdFL/N2ej3
Od+K0cNDAf/XwCST6C1EHvtyqhsq4eKq2YWsXeeJielan8uK84mR0cHRaHhClBdG
vy8w+DfGjtPQxZx5ZOApeUCXgySCZt0kZd/38tNLeM0iAkPLSfu+9H7d76QjO92t
R1cdpbPf61VDw5ZkPHDDshIzciPDWIDS0AFTREmGr4aXbFcvn9GGvIi5R6pEAY1D
+z3fuDjWpLkOKwGeBSHOVKC6qtpbzmDz1hOyckUcZer0CeojOYln82L7SjaUBr15
F2AtmgpMVlt6tzZ9W0uaCmWb0tyee2WRFa7vMl98kTFKAd73WBr0fbdQE6P3nw+o
v6CgWewlmimoLg5vb+8xQzhOWk/bOJBA4dj4RI2JePgWoId75o8MD8hzpmiXVU+2
O1MNHpTmJotcgt8aJ81yzeX0GEe8kGYfenmpInHvLN80QR1j0UuQGyoLavWHjv6H
WiNgJPBRRYZFTT0BSv+EcUwiYU//1NgWl8t0H5O0n+rcOyvQCrgqh6COzhVl5MlC
9S9b0X+/jQeyM+qDXpsXiAuwebPm9UrA61Bwm+VM1Ql2cLrx9X950cVs94oKK2F1
ibJGbHsRQSg0IIusZZI22XaFNK80AtaDXim6BfPxPeNJVzqSDC9reSjhc8fyPXeP
p3YpgrAKPUlFW3Wd8aAf1ImXWsOP/P/6Og3mlQYvfkrjtEJ6QHBGbYNH+p/runv7
76c/LMhgy/dloUmcL7y9+P2aK4qQe8aSDkEDcQDNZ+hUA1cTUhpb0orR4O0Xp9/k
tnOpjTtx/RCUtlf1FUQpEXn6MBji/iO5rDgCtp806i38nbZZ4zIa8Ro9mZpxluGq
yZbWOxd+IDb1yfa495XZGdROUKuds2Mnxb9SoATsiWm/jr0i8aoIaqhkZrrFmMFn
HxkZXebOMH8eGZ9ixtLznTXabFnwsF9ZhTYfzitmvYWwungdtox6gFScyT0kzRrA
g4wLbSuyjdCY7qjZIx6tDDfswMkQk5tMWd6OVPmYHZCth7vsfEtgJ9Dp3+52LtM0
RHeG6eG4JrbSsSBP9eKyXYDw7/51zNnk3ZEcoXQy5ZyE7fwjKZn9zzHKImBSjsz+
ZEzx3pbfsd1ZQNi6XZZUs3FpjOyydG6HyaFIIeHVZjm+Nhy9xwRQHMvKkQounyBc
xs2LOwX7pNQzFFA9EWMDfPEj0J2O0yGRPaqfjW6F7+qHWIrJbhkZpvpTaziwDq9f
ENH+4V5zGtgdYgJu9MmiC+YMMSRjYr+IU7q3vdgvAPLXZjWiHlVzzY9soVRkRqq+
xqEfXLOS6miYatKwnSBcG++dpxOPKbyGGQlDRbUQtpqdwe8XhICBwxrEklaTmJtD
fys6yrZgGpudM7Emy+drmZmxliKP6nTlA+1wk7ukQGfm4n+NEbFNSEjO3w7uY9EC
67UYYVoGchQ27svQ5HRx9VFftfXpCN9+Gi5BXmZQ288678fY2XY1mmXnzTUGlidL
pA+PkvIaMPU5JVETXWDGAumJNYoycn/BVXecSTbz/MupnuE1sOXLodd+MbAn8s2R
TxTYpmsu7ED9i9Pb0btI+O66JximjUKfRmjNQfhzVySmJv56Skgn0FGUKTnpvGy2
ogwDkd3Sx0eo+RhlgdFeTQ3Sq+SUZYnebPWhXpeeayuBY3oqGviegKFJa6nIb7b1
4AlnmuffWyfB+lpZrERAOMdCvIMcGwPqXGw+2cLbVB1I4qiKDW7LLRBfRd90Uk/B
fq+wRGCd51MdF/fOC+ZAc1LddK1t1WW1rjlmD1wmuk6fV8pNZewokxUwYv+vNCNn
lGVM4sHDItSdt6FF3XFzXVxiqcRCMVKD227KG3TeP35tyeO9iz8EP85Pl+8JNVoS
PxrW75UdpgNcNylX6kEDw3KkYvjxs0luzLAS9p96LbRvCKKxc4T67pJ5ui7xpvJd
+HzNVsjD/nezNDG1cB9pYu07EaXUEOspnOhLuvSl5KGh4HbJ56PoJNFLu3sHiyEZ
jGINRxvYH8TuEY79HRj7HcXuQ5cS9B8JE64Wl2WVQwumPNsyqDKknZUNtkHpjj5M
q2i4Eq99FOuwINjYff55O+SmAXeFwN3CJS9nqXUbdZd10FZWxj1WdxNkSmc21RB0
sbrVbwz78N53UZiHjtwHMVy3BRaIJnldXLEf9GuVi0i+T/UNqLPBZOY8rfKQRMQN
GfFzw5tkd421NeU+H9Zm3vIkrDS8HB6BKvzQeVeREyvG/GvF8VslrnWq20FtNcrn
UExXlKvd0d054wq5bKzyRr4BNg2pau9i5onyg4mh81qHQ25Qki8eUD9KRfNt7fCG
I1jmQ5FjhzfG7+3VpMOBSldShQMgg5PLJfz3hhZsGnf8vKiXRQIJbyR/+EpnWpGJ
cMz1/AHi8vgD7tf2pwNwBYijDcwpLSxlNDT38J70WMaqzQyhJHJ4eV7nP6SxVpNu
LwknBatUTNcrTq7G3GF3jkBY/PgZNvwP/V6iXpTxnwri15mLqTIe7AbMNWy3YotZ
vqvv0ydATGr0Fo116p4XIArOYF13OwbKYv5mJjEL+1X15xmNMhnv7D6TJvxI6Vkr
2EhnX2a/h6g8msiaQi7Hitbsat200D+xZvjtTnLNse5G2IGmRKVslVA5rR44fEvq
xhMUcgv3fkuYIteI35epEsnEZShlnEiyZDR/3pB2tI+zhssJB02Mhxp2F21wcO84
5RwLlIXT/0Kc/AHZLzhPenLw8QBG5M0URIa4RxEQrpnGIQkIorsA1Sm0CaojU8Cn
efrDqnFGSXKbfI4mt0zqwAFzJYtvwSjQ1PuuuMNT3RTdrPQGu6QY+0ntnTiGbzWm
j5GdSaCFKBQFYSwILi8qPhftqRu5HKmW+Ve4SWXsSCJ/4MIPadnqi2U0WYyyq+CF
wuRAPvqxgS5is5BFl7jeWNscOPEs8y/d8yWTdrMqY8Z+knZHfczEgdmBkAMrZNB7
HJvJsSGyd+6I2CqWRNOYNRqrn4bewURigmKgO47l64yaS41lc13o93twI45DS/tt
FBhCkT82HMwCLX5ibM9yrHtRaFUyv0WnaiitERSByCxdXjw7Rl8w4+r0Y4Wdjvww
1GjDQwg0Xd7oi1nBfSbgT08U7PrQc2ZXotukf2JIHeFEeVjpBsaj7pjt0NPmxJzP
byk3H/R49gewGk5ipkb1985AQzSGjgf5aCNawpEuVvX+GHKdzYuMtxOXsLWWN6+x
8eT+PeoUHsWbEUEmHeuNxzmrsd5bphtz3b+PDp/7CXQeI/pPe5s8dMqJ1sOYeaXv
jt22qmARN8Qk7hXHu9ogj8GL8oYFx4Li2mmwtXFiF29MlorrJM0jr88jXFTJl/XW
R6GtFAWWBY85I4iIejtzB2myVGb4v7ICgtrq6Ql/VxA+4NIKN8DImQLvNjIqE4Ti
6BU/Da+QdMyyZel2kQJjmHPFFaTWCV7ZZf8rZkQeyWd9SRhqGfZSdOUbqoeb2X0h
9ujNuqkgHYLuqG2+DbWP5b5X2Q1qv7jhdScyAp1Euw0OZAJE6DuEoZiysMoCmL5Y
ttBi6ilXDS6FpEZfHbrGUq7X4xiq1HcE58oViIbqrK2GUmV1PPSnENmg7Pf2zRDL
LmcsxmbEpLQsI/ibUC1wjJTSkz/dd8BKSBInnwDjXPzhYM3dtTcFEDyE03ioZA1C
JZ8ATmGQS02nVx04fB2/IKPvvZyeP+to/HuVGIv/+AJqkC0fVcdg9TuwyBOlYfPA
8InRUrPCDgJufABddTa6nG8M8hw9mtHJ8uyPQi+BR4zqG2Ip08d8+PPU73LAg29x
IDy0o+9QfPaDRPlKtqjn/POvvUV13D1834J7HEfrJ7WRwjTsTu8ON9YALFRA8+xb
hyBTbdhEvrONNd9Z8f6n9iyhsbvfakW9pTZx4NylOQtlMiR+dRf3jEwrC7JziAmj
wr6iw2tf8Qy0Zc7MU2XRG8vejX05ILD1ETdWfZd7c0LSb6aUxUArTi4+EXLfOmVO
rARbkSDfFF0dZ3Cxjy3Mt/wrxK+EKAvDej5NWOQLU1BZG8PhXCNoMN9aV3Fprifh
VXX331GyGjZ9bihQ1u+yQiF8Kpx9b0I9suxURQsMmpD0dm5ff5NCdJ83i0o62LdI
Atcc5Iikdge764JWW+ckldYz+5emVI/mP4jf5sauiV+lHOb95ON1w/i672P+2G9j
PPlhYJql6V9qbgn78NkoXrvCp7SrK5nMlrDBq99wgBv4aM+AcRXgcfnpC0t2SYjq
RayHU+mf4TRNidQ3dRrQIG/QQM8onWj6xqX2PJfKNGspype4ofU4RoTAX2dpn1W+
+bZmXX4eDre2ADQJfE7q8+2XdavyxqBE7FGwYhYhr+uVvyataPfg2cYx1bD/3f/h
x1m8SidaHUPqYtAs8P/Y/zLD57mc4XlQB8D2XaQ5gl/lbqvPDydhXHnroupDvAa8
K7z8IKDvI1hWpZONCUCVU9RRKxbaCdCwq9vr99/Q041VD3XHvQHNrMGaNU1OIh7l
WqBAjvb8xoRKkCemHgkVAqbUj44rYyZ6QuTSNfvOUgWuGc1hmq1nW4zD5Ak+NwCj
OFQdVU3rgBRWFKOs+Uhkk+Ygr9E2czu0NbuS41/ITb/75d+QYTyCCq0iqWGuwmC/
y/3Mt43qWpOx2c9+xF4A9D2YoAqJVbOsEUml8IED/G8Ho5++DMufc+0HrHENH2nL
uQca7GxqSneqJ05VR3V4jrFndNoRD81vosUnF8n7au7U4Vf84X7ZsnulDqzkDg1i
8t8vl+1BaVRp2awkZaFikndFeezrog/tdaWXKvLGqydET3qqG84kINphiv7GtPE1
aj3YOgY99lK3x2WbFmHGrRnAGMZhvFpPoiq3+4gYFunWQFFyOwBaoUqLNysFZ1qf
/WwmEPnkv5nZjoNxnBN4n/DMCymgdyNQquR2ss6vnWa7yhIX/I9/RZe9X6hb2uHV
VmXTN8BQvIm0jzzZaGzoB2+w66gu1CDu8tm2sa8kXLD9R3UqVNhPx68n0q3lMeHX
4QyHif/LDtnon4BsLo3kpQkbRrZz0JlTgLXvMqUfjg+imJmDahcQ152Yh6Q0fNn1
Fw1DYwuY7HWil0ewQ0gfJnDZhZzLc20P98iplgKrqwMplUPE9YLaIfCSTYs9Fxl7
ZfTfIDgl5i2eOA5mA/wwFkvuhUVqD1QGvcWulUlsYq0lNkUY6WqfYVDmQUePrTVE
K94WbbD+9Ek6lMoZ7F2A00biGlKwghFDRspaAAwt1UlJqES+IGUrRzkfOE8qz/VD
cx2FkCWjqYj7DbpB2WCIpyaxenZF87JHuGvCxdjcdQOhPNyZUqIR2BVYrKF5OU8v
vtEey/enMOD24fwXKDdwdGh96pQvoVN8+adkZVToSdd3XVlC0LchV8k+bCFlZkUV
WEZYZwbvKqyiPD5hZA3YeUgcFD3gXraL5JR3MEpIkmW+U6MH7sabkECCdt1Ckyno
udG+5XLORLEQwqO0kCj65YUB1ts7dMog+PCXfo/2eIdQrGjdZWrXd0Z5XsIaxK79
QiJAMwNl96TbAO4s3Xh73uXZo7ALls14JxTVlP4ib+nYh8xxPi63eTFzjFzWvcQS
DjW+q/aJ9NPjYjeEMAB0cD4K/VqpZtX1Pxy6QlhloZQTuO/HFp6mE6fFk4g9ggLE
eVjRt21cr2TUHA4TI7Cu2L/SVfg2b8IUSm5w9yWZPDL/rRqAZ6UJKupi7sUI1gP7
k2IVzcm/PTUZmyn60n8hntUE3gD5LSUv9KUfKqX6WkjIAdoqBSc1I/u2SujSY5OC
Q23NfteAXh71ApAjUM3vedwJgNc1estDrA5Tr1i5BaKN8mGAomm8q3J2IpqcHFE3
vquzG0WsUaXYiD9Y34nYQNXPR0l1suDAKdz3SKGLzOUZWMLKVcnpRriQqQiBr3aU
JQE6F5FcEW1krgucnMicOu3iy0/3XMfnFLUpikuvloMV/RhO4pBvlb2i1KICfWYz
jHwSWmofbtMNesn5Mvv1Ag9Zc49U+Kud2WDwGztMg9of78hKCHq6WAlJ2vEBSfwn
lw4iqxUR/jpmonm6OlcPsMMX4vMpC+QjwTcmv8KCCjg0+nti4tEUAjsAsQPAdEQA
bCDSrJYfgJ/Hp/YNGTUMU0cRghk+eDItmENODPcv7YaEaJW50y/9XoB2jKNPxRnH
3Y5ew75B2xQ0fNFMAJYqsYvjOhM+yobqxjGh9Vrn08+um9sz1sYj3He6BjMASyAS
zt4DnHB1LthViB5D1Wiw190r9tG3KKa3VNKwAb85xz6Je07DrrLGcC+64zQncuHT
4Ezma+9BBcBnUDZVrLYTOC6D24Fo1Xq1vl8xizN2CVbtwYJXs+ZUsBz8dqViRMko
rqtOH5rhfI/dXhgzZwI1lPOuUsSwNfO4527T0GcryzOEt4Nt+Tw96L+KopJHrdcZ
Jmii3EEXz5I5FNMd3tgYo0sv7sF8/ZBDsvJsfn32man8pXrkBG0ktSk/xqfEyz/R
HM9i95m5JIbGItxDvnkeAkSP8wzlL4Kdb8DZ4RyS0khAlMAMaRZC+TF91RR28VX4
VibOv2ibFjiriz5H5Z7xgIVhozOwEyNQ/SdR3riteyUxwiedABVIuKmPtXrZzfD5
FKbNo9b20vD/YjS8o9TWhiKdS+ZvGjUN3+FdqbfohiVh7DzTBusyTClZ/gTc0SZQ
NP8tt4bZhfrVNj5D6rfOGIskZfsJwBtExbLK/i8cMvppkCg8fU8DPjwG+L9Y3PEQ
LBecK9ClE8ondHxf39tBlNhPiRtSE4cwY2OSQRJqeJFagkOSEXERO+ADS9gQGOjh
Y/9g6Gapq4k94SUeaR1ODcwwDTnJ35b2vcA2390VYyC2jzOS5d0p/P+GKO0JDwbT
DENMIFk/lyHxvHmnC3TPXfFDL7feizndpZjSZWOHmq1ao3j0+0NSU3oFCkOQ7v25
DbjYMzt4XCXWj3ywMmoNDZyV8+q6fQ9F4kz2zXVYd7h3yeClAURnedQlZIOmH3n7
GF63LS4egFNxkY3jy7xFhN+hC8irkEoGIAaKOoOo3McsV+SRKFyAcvARenicuNxd
zqE53Cc0Ggc2qqxrxpudJdJxAGk+NZIC+5OHUJ7IvwJWROVhtNli07XRwvexydIw
tkTF31PjuvIY+Xh7+LgULGRODr2SYvZadGeF3aHBhC703fVztZ3MrZ38jX//0jGj
KBlsGW1o+VppuOLFmMwtBVtZOf1wdMsyeoxvacUjFJCbdKMShG+kcrbKsRazQ9pU
l8p0rfIZ2YDqXyrsbjJsiNJjJ5jWqlJjKwz/+3YmF2J1YOtXfB6Erj9c124X63iM
2FyxwxUR82OiW3lP7bxodj/cUx2FN1wZGPbfIAFqQFOQ99NypISIOnN7BQp9fekG
MJe4c5hMtU1Lr7ND0x1fInieDrLhwyknuCYc1JPgL12kMu7JUwWBOft0ZJjMygIU
T77mezzWBr4reJEolrJScuC+fQM4xLmAKZGAhDo2qW5zkdkZhsIxhEHD37uooLdm
Epde+AcPek1Qe8xCd35K1iXl5Y+m6v6niWMAy6+kvaevirbB6yAkztD/xYZVYymG
ctYBFR8ddtYtrtjWa/GhU6GKLQAMWoIY9isgP+wBX18MW7o+PqeMQN7Ag3jUTw4s
Vw64xFUfGE2BcvZnBBZbQmFc48WqLTq6xdAfUW+G8qLifqniuoWzBDcnfvgL01A7
EYDOVUYZezKQAApc/Jz9r6kvgWlnZ5o793+T/Cv2lAPWuk4JfixDP5ZzYOCXogaI
zfIRnsKQjBh2Ejt/SSCzZZhkld+d1iia8JDEPBvfIlXSdAGZ9TSA7ZGL5bDsMCWz
pBkuBGRURq28DgfHc4Z1xDZNKRvWdpaPbTNTX21MeQLjEwggssQ/mwRUYNpU+UGZ
lZcNXdYWbJ4H3NSz1T6G6tmkTzASB+v6+QIKdCL/1WdcOpaZSY9iVljQviRapPvP
249q3wq5TLxMW2j4hrmJo/ChGrxD5vesa0jN5PU+kVXfK3yy/Fg0E54yuKpMwXAw
yFO/kRodmSGrESnfVyrsoki5VgT8mIM0P9JwfAwrJzdPhZoJYlbCP9ZWvEd+q/PQ
hmYBd1wNFAX1G0L8L5JvXpl8ll4CBGuWAd4iGwRLcv/ZnbNmjoIQaEebvQJHVEnB
+yEC8mSRtedeFfzJBHqeyZEo7yvLJOryLuqEMuNADufDTrwdZEl7MIbBQEUCkjYq
0HoGqeI87TPkQ3hO10EufK4TpYRpf5DONkqR6sEDKD729LWytMMtSrVl4vKR+6ov
G5OcM/EHiIRariPMqhq0nbiFu7kso5roS6FSQ4+Lw6upCCyDKrVm1FTqKIu2KZiZ
94GNaTboEu0yKagAXVXK5ldQo7PVML+6pkQQ5w7pVdM7pr79ycm4b+m5Qs5seP3y
Zw7d9qnC0cO2DUhD8z8u8RtmcY/4qwfi/hWrEYzYqUQOMnu/PrYBVJsK4UwrBlCb
DAZ37zdVHR/77WwIqfbgCBc11wNYoKj4s8Thj08jUQki4kmhC8JG8idM4TK0+Hri
EhyoC11XZophG+nRkUkfSLd4VXeezru6aNVxS+1F4dbOOVvIvow+WRwM+TSt6Q8I
PAh7xTSJGJKORE/fYVjDVGCQDmVEA5TrdUjQS7HnSvE7aA/QJzxGusW0sFXj16rz
JRgVzGk8tUtq/lVllsPDIjZiSRhkBth48CGLQfBNnLBkUmWSB/AeEd5Za0nzIty9
qZcvmzMzjgUWGXJWy3mQL+srZNcKX4Mpn++HQ+hoW2dIo5zO3xAHTW2Dg6QsiGyF
w41LX5HWgP8JRGenPDY/h90JjYqJ5QkCG8Siph2jdrc0rud9F6DQiACEICNd2Xsi
qMXKUjPfrM9iE+GzOEuYuLDi5dPROPQc8vPaCOauvQ48WuKsMsMiHdINSqKq1+Gs
HzhR8Uz9wwY2jtGP7SHwC81TeXDHPT0A6dG9jESoS9MdEHKDEFOmO5626hiSRRfk
DxBpd9cvJHB8cn5fnrQyCGEjXetMunczlcEKSYFI11wSVO0SLxurSYd9Ps0z3ZGy
hLzWxpbVAz8JvwWglba796oXY+z8kqsvN+qM6neVA8NucOgGD1IGjTL0KC6QW5jC
hNjC2DleI0eR/HO32kaTulAmMmjpQPZ3rmDsJl6kcub9xZYpY54OHZ0WTtj5JQA/
3ivc5smpVfUQIbpXdoSKJ5/XigPh25yWRJn6FCEvOluSctEUYwtReFolQVGo6a/j
7O8Rme1gAD4lm1bTkHiAkmTWNFhtdqdp8NBbtjmg1UX9qiigg6Hx3ytOK+85xBlW
asD5ayBJ5kn44mcyKAd+gYqP8dMVVGNips0HqAa8j0QNxgVi4chUEAlKw/a0YRYY
TlpZVpXufy8EaS6ZIr2xlFM3nwGjeuG0YON4IPZ64xWUakSHvmeizcyNvMByWHwI
eB2H06VeOWPBhRueeEISa4rCintyM8pCzZlOeoDebuqrSLCJUQXtaqQW5PlqLunH
1/lzfOisNgBCZbQltNB+5jPUWnPiNfGJ51ucTcaM/CadsmlX8t/zaCXVP26qthRE
B4fU8Cf+gQdGPPKPZ2qwUN7Uak4nV8H1peZaeHt12ISO5vfOaHAUtw1DSkKzyofV
Xeis3VkxNbwGX73wX0o4J9QVHNrfes6N1IUFQJNLrX9UJnct1xrot7l3thP0m7t/
kALC5xDz+piz+URXS+n5fawuNGTQxFrFSfLV9/NXAiZKjlSMBqsbk/5sUvupKaK4
+QFdDmt7Byjeeo6ICeEtHLsqMJ68/ANp9Mb+3bMZuMQfNET+teN3zN02HLPM5fCx
BVq7Fy+MwDoaEKRDLb+x25qanBCV7Ieo0STtsAz3i4n45wkoGdNT0Mkig64jUjA1
nyJczJrKbN010xkYmkpxN4McsjhcE9e8iVqy1KJ3wPxFE27qT9TN/XdSbqRv2XzG
7IoBCMmXNNfAbn9nLr/6HrjESQesjJxo8unAoT4xl1XpqtzKBQhMNHJ/aMbLFiT+
S7tPwSRWXm34aOeEKrvgFf4HJ4TO0Daq1iGrkbPX13zf9lKiMwK/dvRc9VqpgtCC
CnLCEBGN5w0dmFTuGnXDXMBgKqL6PxI0Imb4BpaPvimOgotPZpay/xUxObEht1SK
T54p8qO9EwTsFZZGjTYmQc2ltSTmjMuaHl30YC9ya7bjoPA5E5Y7xNnH5VMwCV3X
FC1bemnSyL3SR1/pOGss6/ImWJsBXpVeaVnufreFuucG9UCpHr9uESKFrM6IRjKS
a64qmzeml44L4M/Yx71le62vFehwgbDqjKHSM5SalkWjamoxES4EdybCYSJKvHUj
b5oCj3UExbWsHHPFOwpA3yLlCN/D/ec85bgu3+ugj8060B2yWvXAXIFRgRF3nOXi
gqp2dsTI1tJV2tfU2V9zDjpe8gy7CoXpjjiGJAVeypJRamvxHM+IKN4QzR79/ZQZ
dYeGvFkAqtAMfXmtEUIl5ZTrPKhndy/yXWC+mF5MBHfiRJ3PNEImScEougghF81o
TCfRirg3MbmlkA8QX6SbT6CZrW31injWQSfHEetQjBfLD5wHHO+eaKNLT8kM7jMI
5u9aYOKeUFobDwyFBKexBydsvfsl6ElPZOLZzkkLjPmGEBtVl/NDJ14Ko5wBQA1p
HdGmWxXLi4fSQs/eu9+hvh6b+DMQg3GVWgz4MegAjFOC0BiKaoqtCGvzt1lcFmkd
7G3BqKzNijz5ye7G+mILCmwjXOccDA9E7oeweUXWQI5QWhkmJ34igmaqfl6VXLWn
gUjGn2qMU8X5c+Q1Yu/hTUL/jF1u3qtNVf4b9Xy65i78bcV0gKuFEMR5OG3HHSkw
0C3bkNElulXMUPwfURj7lIZOHd/txxhKGDAsfE+wXPSVo4ExZ3k93vYffGMHjV7Y
G4qTW20xof1rh0Fuc/Rqt+1pXaYioumY/BhXauprn5WgDfiFCeLN2xx7kcqeD2Z+
9KTodswvQgz8L/a10fM/0OnH1139+sWtmOPkyzXCbsd767zKutMX4t6Qw3GNGIJP
puWYsVHsBcvrEu4HKdFWYd4bBE4M8djYTYG76NjnAPyeyJ0FznMxbvEoUze+tYFs
SjYFv43aSAxCCpXTWuGp3zLRaNfPJNnG5m0P0RwmP+RxtXUnN4n35VjJrCaXkGO3
ddZG1f/o/LQ0zFAWMB3Aw8ohEZkhEglH0KHcOsJY3Nhw7c5MsRNYl1WIayA2Ui+z
VFnuft9kPBLPGuJN4YyvluZYo2FVWXlqrNNpZbPXnPvaAGTUyHXYZ7rf9Y3BfBq1
p8L9AWSn9W8/wgLrnRRBr1V/JpHDwfKVDPOySNg5It3sD6bLtDXsXaDeV6SkMbSK
aBbAbHInL2LIPwttRjMFUnABnALksMIdAHmkGlb9Y6QELVOojvweWaw/kNNb99Qn
GBNtZB+ODX8sB8xhb/dMvolkHwdtNKIqm9JFIT2G9cxhYhWGvh0W6NNZmFFvAjmA
z6f/3T5KKKS+w6aA0iJGVHhrOgDQggmt9yDPWQbhfto76rYFdq8aCozc3aqoOW57
gJ7uCUfl6Y5dQ3yUWpxTQus27c+ID8Q8Anyw2mkKed81AxGX7K3wVpZ0TRbXAbw8
CQcCs2zBtOVVHnsXlEuhNlpWcrqd1U35Jbk9RbVIB9FGr1mSeAxm0rAt1irvRc8I
rLKIiXVCy46ssQceiGolHooqKliczhi1bXA/LxsnFFwuHdqX5A3ZcUGkep2T8pMu
NafZqn83u4SrCEupcwY07Pn/O0KrluoqgdAcpC3Ckz/ys50udRFSS+fqWqAbB21H
HH95tDrDpvPGsJ2qLqnVJDmW14ylf8EpMeyr37I/gplVOzGRp8/t9DTS8dlCYHdp
e6jUHJkJQ3SgqM+VJMJeXJ3P7j3481gFti8E6bMR09kA3YPz0V8C1nShHSGmLt/V
ltZzk7oJzjLhihq9NmEYoc+PjpzKM842As+8O6yLGm0czYyqKydAk1dq0XpvDkqc
74+0Zw1JQahePl2BB7MBEjju+2Yy0t+1HMhh1RSH0mk7lQUwFBtyQc++5QtxxTQ9
fxes+5LCcUBNsjYyWVtbQ3pdU72i3HQhUsWcNAQR9LuAv/vgMR4KoQiIk1gjkkU7
9cqvW4Tcz9GhX38LZ7dYJ5unKffxWL/MAxRY66EjWnAknqACBBJixLqaUQAni7Nj
pbGeTn2jEBIT1IF34il6s4Hxa3lu+3o7CrxUl3K+tTqZuwfaZnKtSi4eBvudpqdb
utXE/9BC3CA40E8m1yYFsogg53FhiRnnS2BV9UuvZ4q7EV1J3P/hoHKLCPK5MXGA
lNe5NgskAIYlkJbP7znQTCJR/p+O8beD4IUooTW0SkJXo3ehgSV3nsNUjpkpEciQ
Ej07Vppyg2CwVdUzujZ9SHx3uaPCJVgVJKt7baMMTmDq+qu87Olh4xMqe0TDqNH/
QdNuABd7UZAc5ZtoKBsfuuFZc7rbCk/02sQoBmAh9eTukqAf2J0oKh/46Tsewv9l
OgqZ9ssu8bYGr0fYSqeFgHxRJW1EVtLglE5xD6E8V9uspcTY++cirQ8AHXFeYV4Y
1kjbqUHhkfy6OL0HYbIaROJZSQvP9sGtnEcPXU9aanUJHSq7Bkj7MI6ShXjP6WvS
yHcDZdHAa5R4SYHV2NDJJzL2espPYNUGVCDtBjp3Xzi67kQNElK6X7WgYM7z0dil
RTZkaaBwBgXO9VzBrf3FjtAVCHoljIndTQYNZbKcjeBby/Lf4U3z5mcPeFOacK0a
c12T13pPsuhg3WtOcjgM9weZj/iFQxrhn58mNawtppw+88Wq/PQpNIn+fuK0rKqu
V0ZQc2Gi2WXPupW8Vm1CL/1TsVgoTSeP+7kb/KNaHxTOPVfhyPBq9jiReXietl00
VlyPVlz6MUzSAxx4qXH4n7l4+ga1FhK9sKM46aOv7R3WhFIEZt7g02qO4L5Mzko4
t4rHHW+CDUo34YKhi1sV3egHQkrzR8lMasRXQC4M8g4v7YOD2w21RuOZvbjdr1RT
QJRSx5JC67rr8v1R4trzTp5LMnw2mFsKaKsnpf9UJ4pvL/JP8zvEVklH32Ym3pf9
GJqzzaZ72KXsWskmwVG+U3Lqy9TY5u37pK55vY6UVnheb2LggghiKiwWSfrMhXkC
rcBnMrQBmAlLpcXPAla4q+TeRa58F0hccUEmYmMkMdxXUFWLbN5oDU3WYSjxIyh1
5WWNtHB1RnBCPw5qC0Y4TkZueXWQDbn1JWnHMRsL+LrtuicQaGa9uLvNOi7GyTpU
q2mSksR2K1FRB+fLYWxavqAhA4pLD2HUnNvRZM9eS9pcA9IPqzMdwBQ8scmVnZz2
SK/Q3jxaOQLMLdPWSlHHsA3Q7FYX3V01XYSX9MGgXuh2kCmESbCZHUW01Vo+dF5m
cuFOPfxfbi/VacA/9Oe9JWykyxFx0aVLMGET4v5BfJ2/iDbEreSuWL9Ynz5/Ns8H
Rz8G+eHAyAF/BRy6PxVH6iGhNG+dNUGgnbQbu7P6XZnS55azKKkMxUAp5hLQx9M6
ySs2QhCwWPjQIO7BcK4+2H8St9WChOQsWUxlsqyxo5lXad5dp/QNegzCqdHOjnf5
KyZV+/y1s8o/Ka91YMiE75jiGCa2xICn8kF6at9qe/5ywaW0uTplTx8orvIkAlFK
j4AZ2j1r0s9clL22l17Bf7vqtl8ks8G+eC4ItbP4wNv0Q1VQE5YsH/ExOtrR8x12
IKAO+7C21nd1lZ/evdSL8LIxXZK5m2vjqJGQSJENYeMljZ6UugiF7Qld4y+fAgBA
lvn5iQf1DptS818d1nNOQwug1iKF6b+w0AXnhjJavCQI6wodYBCZDn3otW8DDl0W
19xFI4SvjUV80+8Xd/1t0NyytLQRcOEcfnBQgx79K4A/Xfjvkmufr2ZLqYT/P45/
9+mI57Os4BUUcaCikLVpG79FQe5uX5d3z6zGY3GNgGUlkGfO4Lzk2to0pGnuomV5
JnKIdo5m8/3HwxgK5Xj5VCAjf3NQkZYlKzUfJw5DHPEs8AkR9G1pNKmMNyD1fJhp
Q4Z4SzQF8ppVcYebzSa9uiSdJtV0sUhpAN9dk8u9fJqfxQ+z2EQaV2MT09SODiG7
54ISfVNIGSY4yOydN0q3af8PrGxLvrdjRha6uGf35HjLvvNHpUp+QDsZWQpe3diA
dy7bOMQqTUuyhfF1BGrXp1lFWEDY3k03maAVRJByYo2KlBCI4qKZgizbigrT7KI7
qwksCezcbZ1fWvfoDKIVsnmRzTQCdYOe5BOsyGX9XdKIpANDb8mE6qkbu7X5Pa3H
/mts1eGUjS8Kz9nf0ygjGAk6AXEUPa8VlyAg5kAmCZ+rIDi2DMURqv9oJv8zKEir
ytKxLiT0QzD4PAAFqnj7KSKHf9Zk+yIpGPhVU76efajLxLOiiPH93LthMiiNRR9s
wiD4Y1EWAreW5OistxgBQDORpzhpzcWyj1zlBEklFUiDSyzv0jHz6ZKhjPz4Cx9E
5h6tYJrZ4YCAjSKLmqw9mDC1J0mhf9CSumqLfs+KPQCjtTtOpAloJCpOClBXUhr8
3h+xz3xeJadeWarGXBRcOLSFpiqH+AvzZ0v3a9jH8/oCEBxpgSKAHOlIsqBP7fv+
iM4NtKRd+FGM1GHMlMlnq2FXnfInDCv/bWAZeEyhWzkwQ0/cYO2Pji0K+Hnuww0e
CjHtZWKYaIWjw3er/wO3Seit9ow5GxO87M5MLZOdKzMPn3q8CtZvD78K5SsAuM/y
NirLNS0PT4HsIgZFbtsCvxTOvOH3NYYECmxbFaM7UOWlk71TZSmXV6dC/LTYjUeS
jkQk0srotfmz9qYHMFqcZMTbYS18UXhrvle9T9pL162xSQ9gCKBsmuPe4D7SzGcC
W1hgcHalDxn/oZj9ghEp/EWIGj4huiJ2rpi2EPswz90gZOQm5EPEtb2+nUoYekJP
k3wroVdo+LWfJSS2W2Uom4YZ+mr2i6/Ik3Y0KhYl31YWOaIEzjmC4kNvXLhAoSpd
Ddf6zElY5MH3T5sMJPHIDeyfFPyfL/1j2C1HjC2Lqn3VcYfvjsrJqwHu3ORJD6M5
rmR6W9j5p5j8KQf+dXvsATd41+oljN83GkyESBrMu4DxUF0kfhcnSPqDSl82Wkp4
am9TXPmCamE5NJa4wLez+wocp0Hduwxe82JUIWPa19bzmG+OG9QGPylU6XRXQHl8
pFcxTAuEEwu1W+CNbuEz7OZ2KeN5tcVj1+RumyMu5mbGGHh7ntn1CgsohT+XLsNV
IDRogbKjtU0pRd+IFfNkc6KxOdUev7ScXvS7oE+/oPPxnrF0MmeqObtT7JIJT28P
P2mtqsaeSA23wNyCG/KsPjWJkt7+yAzRz7HV/GVN4GGqdT1qewqjepsoQKGM/jbi
BN3ATry/pGWkUesJRBObzeWAl6LQH+oAhZ9qBZI8tRPEIFQ2dpOp3wlLTNfGdCYq
zxAZuE5A/WqmOeIZvQ6e+NgC3SwMOd1SGLisnCA0tHVQrS6dx/9iq5tMRZ9j3f/1
UX/O1wPscNSojPWnw72uyB60yJRR/Mpn0gHEFWSn0i/JrCy8pedhnmQFzt4DxxqX
Z074eHgfRryAE9aGKLJ10p73uMMyia9NEGAJHssR9/CynA2DV47YUEBdUWph26G5
+1ecNFO+vvfMOr3O4o60aoA3koQ97haH9YYqUxGe+TESBN2jn7pCaG/vE9DPPZ2K
5+yAMU9CCsDK+Ydyk8VrmmrtOji7WMXWjgyplsu5aK5TMTJpuTL7CR0HAT2ee6dy
rR9Qn1iQAc27kQupE7J9TWwknGsLyu0K6AUmR0qMN1yivmCpVB2iyMA4vVNknpna
R7HFpNqR5dKqvF7zKYHuDE9pMiKohegUJpV1wVyouG56EePopIh+M0uOyWVlsYl+
PRg4w3xUrBR9DrQ6BMSqnYuwp+iY9nxNeQ8KDC2rEGJt1jIHC261FnCLGKPOCVul
EHgW3EUBqKu//ksvXDLJlz+bQwtkJsA6SS4vsrYnfYfyuUjWbG0ht4MGg5iEvQij
fAmHtf7NUQZ0qXPjQ+zNDDu2S5+jMp1EDsHXD2xeGzwCAyJDcCa3mqe7EdvKikvj
6TLgN6a2tZLEXjP2Yho7z8z2oaOLutwWZmF4vcavc6amSQWDLb9k719/+h51Xc37
R5TJOGOwZdkwnbzlMOtmR+dfIL9TtYpZu4ZoiKPZVZjlli7q510zZNQjvyWrWG/q
m9aNJ/Yej4AxtICyiSjQdo2U6GYlDMttQoX+yRWSalMXYcWWgVDG7P9/O2GzC2jm
j+s06XusTJDkg0QvSZOQA6ue3ezj3IzxDjdt+4t/YX2cL+RcuQhAmBtjxZE81iVO
CVljWt9zT/v/P6N/sfmA61xbLyRK73Z0ArcwEblgPwVwW5QMG+Hfs1hxZ3FoOQ4G
aSTMPFwPQoB/pXPskoUNvtGV3tqStOh3/UdheAPBgNViaOBXO22p5ZniTs6gjjwr
YwLPE/up02YgNNbvtT+RZhY2nyezsXFNBg18QoVmhYcrPkk1E/T8pegh+Vc1m91z
Cq7YM6AMPXNhUPzeYfUdub954A9oif5CYByt7Vo6BQI5OUpHWTZlRZ/A15pjB5wi
ojAJw1FlP2DINxiJxbqz62J0lBCBUSEoBUZao7ZhqbaPUEm4OBBPUxD84vo4hEWE
oOvvR6xxSmTmM+4dl41B0Lvdt6yYm1noXhrwRSK1sckuEevZuYku7IVXu+sI2QMJ
xUZTq2TaezQ4FFihzCZq9av16gSdPqnKGy52ccrKlJhqADOf1OVDZh3s17/lz3Jg
yuNIwUaSrbdHI2YRRRx3BZW36daeQfmi57jnxV/laENVZTH5MF7h/yOX+ooQVp1/
PGcdZgJapGc33gjZbe0dm3MO8tb85zMS4xhMNrRzZjinvCJYT6lnvJkPFWZgq41f
KdvjX2HTBEB1veqr6YucSB8NvgEtm0j6MaBIKRXNtykQITBdjTbBTrMJe8CDfMMs
3eAp72Ry3PfChYLj+ZGeSWbP60Tfs9UVXFNL59lmChfFddX2jpwsbdj5MTznzxtJ
IJKbQTJJz9mxb85BdlWuOdQMx+78vxBKK5wBr2dC8UCXpm5egmkRHjhgJ3BESaBl
G3YjvoS4YtOp/Av3hfm7/VnFzKtWomeM0Jv3ghGV/uvTtsha1OZA1BZjeOZmaEQo
JrXfPwnJ0gPSdDX4pujA98qxE0U90iMysjnN+7d8yO/Ul8S4ejnYJmDEJxtYzzTh
2p1UXBVvfaZFIm2dDzqM3Ysyu5YHnoy1jhA220sl2R0Z67ax9M1/F+fDjnAYa6ZT
CLTIVBtpXaOd1U8fALBUnnFTexdKJjuW9sFay+3upz7IFLM3xzBt7+pHV5+5Twsz
2IBudOzEguHuRqqUDoWCdmS7uYuMY3fsxUMFm9iuqqwj5t8jP+fyfxIx8PqV+tt4
imomVtLyNCbMWcl7+/JFTJmBYzWf6asw0vHf1vWgcaYN/mIhmT4ra+8tQftLZnkc
7H1ySzScMmTV+0I1+sMDYRoK3fcDkbT0vUTWCRPCBOEk/xdyNWFoLyxPD0TyOGYY
qdyRKy8p36Qsk4Xj10TuTeTvelSO4dIS4ISkbgDIaE9C+qxd3wvzfJthUEU+PP7S
ByHdX5ihcMRKePdAn70s3ooDLhxFNxm4sd/yrYKYt+ZmzkifIN7hM7Ui/Cz9NlBn
ZqbDFYJOsNVqKlyrFRyqbUziK5smNA0ZSCRjzDFh1H9znuxLi6FbuElGKhEcqJYH
b70y6y3clqr7w1oSlpyjUYjxstJ48G90yZ1u0fLzVBc2jYJaps2He57Y66/cMXI4
GXWp4tOi2iZ/eevVkOPQmhxtzhD3EHq+0+fJmP5E+IYPtk/T84a5fmsnNNriqsgr
XIyjz1cehj1BFBvRjC9dKkZbOY0LQbxuhvu+gfYAMe0yNJNu/ML6nIG0rVn5vuh8
bqkzoHn5v8Tz4gNi3ZGnvmXxJ0bvd/AXXjURZrQt52P/I/VogN1gExg5OSyXN7JE
9W3evBOn4+SwPYZDyoQuXDUO3Dj1JrH1623ZuSMKfPPxPYfw8ScTMJALs6Cskmq9
5qe1KFecYvRAJqnc66rIut3cOuUGikPXOLfkVTAXpZRK/oohsRcASVJmzt8Y/+NI
3Cv07+bu3I5L7vLFAA9W/UhHyV5Tmd+V/qBs5aZXl59bnL2gJqRCweDbMDf02MtR
X4sK0z0zVzNAH6BXBWLIVOaQto0ZRqD9RNenDNX1y8BUnKHpclat6PshrQ/VpJXP
t/AonuEXPmrLIZOZbUnYVmfp3NHXZpYF5yA5YACZPf2ZZsRQUYOvdekeXOaYO1uX
R0VKXVxfTgvLnOAwwBmyypZqMQwqsHZibzb8Ea6iBj73Mlaif0ZkOiYtSKsMCp8A
RURqSPjyHQTayTo3YybfDPpXx6MftTI9eVglt2V4g81wUQvdLriaMribQ6G3zihl
LMjmzv29KWGTkR1q5P0usjVT2mczHOkR/8izBtZ/Duh9ezjv014yFrvpJPOed7Z1
FAWQsxQ8AXsQgZQpiB5KvHYZCSRHFoipW6EOjNlSo8I/OzQPdaZ/8Jkg59KkxT6R
6lbDyYxp2E54BcFLPjbTQm9k2RRhkzeVACpKwVMCTn/sq/LPg1OiSCSLko8zx7jr
B84/GvkxPUB5lrRAm4CqtT1Vg3Fo9s++UkyQSLNcXhAA9/o5FmkgezT8t5n/uiNb
ikEZ6eB2rgROCvksGxMx4DSFiZttWr6Y93RYQDVQ/eDJLyBPbOCSvYw87DdH4S6d
7BGfB+8nwR6EeDbr6tbpvhagPozRnCQ/vNEa7D5P8Uc17uLdD/jM8L8O5mD+igoZ
Uzk5ck4sTW3WUvi5zoOtIsBMpdnNBh+kJcY+xQ9yBuIrpMnqe6saGxvGeeUnL+yd
F6g1rlN8HqN/EenWX4/ebF8rS6xRj35DYM5bFVKTD9ctuqhRZzgEuCNl9rNbnLXR
jdSC1iZueSQKpR1cGIstpRm3N4h+3ZJRe8h2tP5a0zDApJ++Rl1WBnH13Pl84FlQ
hXilhvUeG9gA+O3JRteTkFhl/vmT6LnnTy9Gxp32Z1FGfeACIwKGhQov4Di6r7//
gT4JSFwjarZ7auZWVLUX/slVfyQqZ5wjI+2wRgmtKcez0dnFk78dIAtQaceobeAi
3WTPU/dUJs+euVpOi8BACws1735rSREL0diH9pyFfl0Ja/o7Yww4GZMSNtVJmvR2
qaEksVs1Ta+SF3IOlttJpfN8T2l6b+GXKe1axEQtpxqBr+c/ubIazrETKdErtcnJ
urjffIpbrs/1ZM9M+lPQYmACHZTOos5DnabAEQvBh2GXI8axkPePm1taH+FYnljX
TYqizzBoO9eI5kUmk5Hd6+yDkUeHazmBv856D08jSVg6I1byFITqQ/4vICW2Olyb
LOc3RR/ymTXdWCJkJpxjRjKCdax5kOpACVYGyTpLyFipud/i0ZCuuEVLm2iBqfOk
Eygkz5TuB8CRrK8uxBUbnLXF/3nQInECjzzNxgdp/2AhQ64ogUS9XQmULiwhiDkL
utSidxc1vTKlcw04TWw+v7Hk11toqFVd1NGUqQPmFjI1VZcQ8f+QE9FIYn916Cjw
UVLdAJDFdOlp92FgGdzo3X0tX8/o4YqMOEW3TrjIn9lwAR5RalpGOfe3HscJGYyR
DMY1zqy3BOWuSsaoOci9tY2+qoWa43cbvy+NBNB8/b3OMlH6rEDrD/DRoWnxlIA1
fNXYVsePvT9wKi4dVV/JY8Qddp55wx7QSI4JMYaMukXOqUCMbbHYwvY8bf5/cwaU
BHsU5cRUGWx0KR4KU/c5Ul2n18hVohRDcaAyq6gWeafFsTMXtPgrpFkVThIutaAF
BoWbzZEY/We1jhHoctRX8ZxzfaLJKwcBXxx3l7jddfLErjurD+liSweDuSof3ItB
/XQpBhkxi3RaqPHOwRIB/nVagpCUpPN6huqVCDSGjiRtFpt6PRV0V1k/ImjFSjsl
nuyEp6xkDcsyqndqt0vlRY0jXGik+N/HLEosOtnBuh5LtOsVLBVoalcyGYT5ZBDv
XZE7sSvpNEi7dPhgbaNX0VYH+5yCywlLEIUUKfJrDLDrYRSh62VLmXc7VZyKJjDr
K60tfpKid7R3hvrNNR1OlyggNwoviM+xLwxNi0q/X6xseF0CODNib588e5T7kcSX
CSHdTO5CNlV0CA+Wf0sT/+WFvOd8r2IzO5FWiDHC6pokDZdegxq4obERdkPVYX5I
wjUoCaJbIJ0eOtjI0WpvtbBbmtm5nj5mqMKPXm5YyiyWH8d4osWwVnNhbieUsBqq
lgk6vvk9blsZMxWV0zkZVF/yA0mlG0S0KAvawe/XskkULh0SAnDVT+45tQbhvfya
rnsOCxYkFw0cRrroMFl1VAL4Diad/fC0q38Q0uVpDM1UVWQ9Wpxkj1chQLitLz+d
/ujUbc2o+ay/FMobWkfodxaG/APvTp2zkA4V0XgFwRZFMbrxPVZZV6HlwrnOmRf9
peZaTpqU3wRg10YnXGV+frFUWGKUh9coOHF32LqjtVqykwXrJu1/4dEmLMXKn60i
aaLIWEkuDvZKWyuZ6jyYKxpqdohlaUW0ax0jl92LBRZn6sQM819PkcMafzJlWHHe
wIONiIyyWr7+fgj8FEI8Xg6n7hzANro6X+xJw5Y2HnNN20xeBztFV0nbBsueD3dU
vUdkYBWTs0YYmB3MlabM/7aYMPP1XSuDrTN1lh7G5yPesSi60cyekPEado/zf8M0
b2ORhJ1fa88vZGyxJP3Ioxmk4xHu8spefvkdhj+1PNY3CpBCsuTYrmA1FVlRk4cG
AdjSdoo7rGprtgJmnmQHRBwF2WO66S+S150w07t0gLhFnsoahK3hcUUoS1Q1MYBO
1U5hYjDwd/Yk8t+qkIASl3vHjThHuPG9PtAb3EmsGrMPw2VHBWoMz63bOr14F83X
YBNMQk/e8uoT4LJaJYEiTOgwXlyH8DGN36MFiTBlhECoqRcxuPsbC6MhXWUo4f21
emTS4IGwGArVsMZ+lY6zjLB9tdYqOCRn0ifUPvLe2XcDuw0eHRWbXGePO7pvsC2P
9UVaYX7KsOapDRr45VcouwU/5CundR6l5/bSbkU2OGgXcbY4xY65lbYNUD7hc6dc
NuyXgfGCULBwQGcf0HW5crG+XeRALkzGCEfmgLgOzBlWCxGhApYJagjA0cdSdTde
+95IadQlW+dJyT0HA5obj+31k6WBFTbkcOum+OMktYXT3y/zW6OETYvxz/75w05Q
/J1+KhlwzlV3jFCV2GEaXkMnZeysD6nQIdK8SI+n0ukW1F/SqFRvHfsI3gXs12T8
E7SD5sSJeG1Z5l0PoW5C5BvBcmOZfQzVQz0oHTWIwBrVpydRHbcLmuiR2PatDHRi
T/DluMqwwKCkr4cZEqQzF+pWUQrN0004LRU7IVZw/4ua/50t7QNrys8/5/uCuQ4j
DEYnBjCs3pnNfRgmNK13pA059+x3iUb1iaWnIbMXT+7ieShQ17n1CZHq44yxpXmP
bIAjUNOksMvZPMfaeNo91LLRf2jLD3o8NOjdXyoWKiZUogK5Fv8Tsxv9LkZ8GGzw
4+dtsDpLbuJPzU+q34IUOHb9EQBvNI6SZvvbHAAMacG3SpS9roILPTLtTCddU4ck
ikFFW49UrRhZNgWe1Dy1z18CacvBrxHFdpHKhFF0QXdwT1yw1nQnsNW7b1LwdzXY
I+4PZrZ0zApZ/faEYpALC0sLXjS7lVwoFyRJRGfduSvb+n/q8AasuYn3w1+h5Qhd
c8uSlhAxSCPDFbuCLZeb/r4OMn+eF3Kl04gdH8c4N0sNtfO+nyhA4n1fL1UNmX79
5CrfvSLKH65fncQ7DtjUq8zNz2V/yqE/TjBBNCqhdJ+bg9kHsTFqsjbEITZqidST
cjLBmrpb3Kh2mp62r6y8IudO4sgNJSyCGtu8R7NG1OW+qohyKcGBGOpIJQkdhWI2
Jy6DUXsKWIr7PBIP4fBfp66yDe+qFONHRjog5Dil4s7pU59r1puUhVZfIu7n0Mpz
iZ1J4aZy4T5rIzSAcvbwpksVxsgz11HaVtNvK97xFJmJaWUeppROO9US8CzgLMLO
WL3iMarXnty5DCcinDTDrnCULzTGQAwXyl3zbVwmdVGM3VSZY1eR45vu/+Cj80Hp
UgYSozHndiCZz4USWkzuDd8zVL3HOgrlf68+Dzahji4l1jrVkPieuyNXoEDK2M/m
I5GUyNAou64b0+3pvFl5bzGGud7wnNlBGUmdx3btq7oNa8oHmTfydKBJm2epGdgb
TcRK7GBDDIIEyDGrXySFKZ0zR84k8q7tM34hc681X5dntGnUsJsHy7FIPTkt4trr
MrFrxhj4zgC5mqv4Bk8yE2828Nw+mDK48H7s/oJsZ3KFrERccm8V/dpb0t1e7jjW
kWR+7seNTmLv9i/AGfEapKOKlnvT/oqJsEI0Lj4nEATwo1A/Xr9tChyxFVzJhCp3
6b+WN6TjvUMVA30Yz2oZ6MTbeJxo6onvfEDq6zHV50L2jgb1tcQxTTVmPZdAf0qI
9xtu9nsPQEEZNqz0Ik+TND3HLXibFqwJz/Myf02gAajZTu1ylz/FXddwkmE988Dt
QK2TQwauQsyX3u2fJpUbO/o9vRKoE6dc1QsssPeD6TaB9rNDjwhbG/holBZ4LPT+
LBjZS5jQM70j6y9Cp40YoHKJY3smph/8IWxGJL3wzRmrt1XF3Eol542MFniSMUwk
IL4JXJj7SOXwdTJ+G8ygfQae8kaPTB+B5weJFHPRhdwsvuzHlmPulwUjuw+hQjrt
04BYYKYU/nIL91lptbZGzGMUHJ85aOIxA5whcfz/mdKmPJLaothKmEWNIDjUmHLu
hKIGVIAK8YjoYRShGZZ2kn7Yik39TCTF3Svt8t47Hf2FGqu7/QlW3ddtiWenm642
/xwrHGFuuWpYKAu5Shbz6KajYsjHvTjKhPD1C0DcWTNjlIHQKjioTR48hbYYEpAX
XpdFw3wOgqfZnkv0lW+tF7KhHWinI9cS/Fk+rIhmSha7rL1I3OZ4jp2HiZficAxN
PRj1XVZrXb1lvNFSdW9bBixN+LWOeXL/MQfrs19nDMTJKlqQIHx9iJDED4qzGfxa
Gfx1gQDOPIfuI5GAXpuLvMPXTiV8tX4WII+wZPKPfDTEcUWoXYupiAjjiCG75oVW
lXkxHreNoX1Apdo8A6MUqnwyNq6FM+e8yZm3tmq7r+NBsmFkTSeJ1LddrvjIRZVq
p4Ow9Uq5j/YExS/TkbhmVNLsVXc2YgCvwTpYxyTKECKjgPOgp0hmqJs0huZdM6oC
QEwVp5VngwkfeB4qePkJdX0PvQQWZX/fGs8VLdJYaKgS/NJGl40OTNITfqmM3cBY
VIXtE5U72hTMe8ab1ghi3njpv4jck0WqBS+HxGRtEevXnYv4dY01H7Lw/ufVfR9+
OtiQg2WryE46sxHHwLCNWvyHZHaneD+VBDi6KPtD+P4/dAs2XOPbl7TOva9xabb4
2UmKQuuE9IWKrA4WYfEYDHxYRn0V+bhGYN1ETBV/C/dOj6UBphOYKwcnaJNwFhFb
SPaEw8WQZVfezaT9wylzMihSgYGkk8A1SD/ZyOrTvC9lWAzuWWxwGeE9eg7je67N
QGhglnccSL24BPxXTIJ1Re6xNB95F2v3jvPF51rfJ5lSyOj9YtMdue4DCSZWRgZ0
mHvUaKB6tN+1sloQECZzuCLsdpGdofuFGtrOa8tSstN2UBBlTVAAB1sB27eZWefv
KtB1NE34BGX1l/EJnz9U3C+YRUa1VXdJAFfOlujYgioKNGFOqCisMYK+OBA9RkJH
eFD6voVbHq9F2e0oxR6U9DyfeVWPyNTS3F6iBJleAdGA7KXMtZMIMbAJzpA5wznJ
xO4K7CrnhlGEn1dWSK0oU0jSVmmqz3RtMPRu3lBMTvLoAyuy5cv0LtdspZv9a5Vh
sdkXHr9yLCeHIudIoPRmID9DqFYf5YOPRZqn8PRxumZ9Zq6G6CCwaAIVfKC+UxCS
em1Ig/KUU5l9j5+9daxLx0unKUBItqiFnKgitQCeSF6F+qbcsvbKa7bYVAAvOQHN
pR2TVJYr1yp7siNS6X8KZgu5O4VY8OW7boy0cBBf54Bd1sKFH6xc67WBBOW+iJea
+eFhx9jGQjyd5utT4iXLdPgNa1U+Y0vN2DiZ4ilXgJgPOcxivUIXW9XASZPJNI4w
DKCCyZOlB2SIzM3DaJDaryjF7QhR6vC3ORfW1L188Y6sFaNY3s8Aysgpl/RVnN7n
9tRBE1K3ikq+8b/lNcCWk16g3B9ZqgHcavw76LHgOgUUc7I/Q/reG4Gr/8DEBhJT
s+qk+ENc++xW+ju6lS7731+AleM5nstXpoOjbfCma8PhPDLveP/SA27jfPbo3frH
DMb9cDnLLWTTK78SPD7axXq2JdFuYQjG41NbIEO0V/kVVmklycu40vzz3VN1N9zI
YBeBxaWmMlqbS/SSInm/pGKbfmaYOcyYNXpKKQWNNZiZdKRVxmcuODUWT3ih19/o
DwvMO8FGmB1R1RayPn0GioHrfNAyuYk/hI/uGgfl2SsoZc/ih6tfyvFkzJU8JwVn
KI4ty0TpWpcuvkfMJb4EMHxvoIInPKxot55ytpmugz0U3ODY3h71S+oPRmPDlky9
P5NcYC0Jv3SCzlXC/GoN0Uxgg7F/xmACnrpwKAIJ4306d+et+tpsv9I0elm00VYM
j/mgQLmL1hfck5MiHvo4VREBxTg4EjMCm4X7HusZlXQEezsAJEjcP3cS+OAl1rCs
T9KdL19IRNBbyTtiEKw2Vrk1Cq7CS7II/FFAhGJId4vrue5VLu3NHrHjdIyu3Mle
bBinReaikQxe0Y6ngdAHf11BdPWuJBLNG2r/MLXSqWcqdseu26Vf3k7oJtA+NScQ
xndejOvwllxDvlk18ciXp4IJG8cq9WO4VcQPws6yNELeAWlJYT8zlUbA7ZkgzVyZ
yhzOfwgtrTnr7WRUp2GhFMGe4YMQfgzmhmeJyKP8E3wXZOiuAaknQooaox2NyWV7
pxfKiCe4vPC8e1I2AT8IGgyCTxjDxZGa6SOeVAXvEW0LH+WGOxfPB1tcCwD/1x9W
Z14oc+6pcosCodsMUAkZs3gRaqwareaMxER0SVKjl4q3rZGw+MXEdmfka3z073se
OyU/qZ3XTezVo5i3ADxyr+F+6xG+upEbgjjVpoYbPC5+gbAw/P95dipyJlx/wRFu
IQAreJ932UNU9o6NRaOuCvvDNpeKvKK9JZQFtUgooO1bnwDJ5pIpkftybiz/bGzP
7aI94yp41a9jnbOlhbylzmlOWF+ocAiKZu52AeIQSW2g6G9y/c9FofOXWJnLniag
djh8oaFQgYhfO4NtgGoWwpmS0js8ijGwHtGY9EtDM9/TGy/0RXmhRWsEk7TXKjOP
n4zzy6eSxvTxVaDv/hutnTzaYJEsyuBlRYc5l71CKqwQ/ybZNFMkPGIKZtocCt4i
Xe6i3oH8wflD0BGFZ6I156k+9XpeJRwve5UAmg7p5n3qE9+7pFvpOmSV1r4HP3Mo
hXY+/tdqoqYVFKa6n5NWrxkWdP4ak56e9M/dYTGdk08yz3VzIrgTigiqaYxQEJQp
iuuOgBg4hJXUmSNCJ1rvaxgM3H7DeFMXaPS8/csxrt7W1P5NeCc3lgx5SXaJKv6X
KK68F4OmflbSehmB3Gx9bwA9ejJ5+zkR0B5o9LP2x6D9SyS75UT6mjbbUbevQ4o3
+uCPIEyAfRHf1ZHUX6KY4DPX/li8ybOly/qBGkOzUwyboBUWCx4oOZcw9cBAi1RP
mnKapyJMr+OBPsnPya2XN/i9z1e9JBCPTe10tT88TsxReeX6OsiOoiOAW0+oEUtr
VcZIuGzb7P2l7V5gMsXShZFPCadgFtlPD+Y2yxa+dluRIsqzEAUjWD0EC/BwElEz
lQFGZTBWX33vTB1N9KZvxM5q7cZS4DNSZnLdJ15q3gung3ghpCRLW+KT5vkADM8z
CAkSLHY8xOfhBvhEETfm1lLCPFZVdz1k+BBM/wySDSJwg9uXLjUx/21QW84Mlo6e
XXI5jsnynYE6ta+cOsdpfVSdupgH0/eoyH1A21QOA4u+T6jMvTYBmSIKXOY0192E
QDEu7iWyA6hxbVvaqt0HsR53VMffysDgiSAgZBJaNzOZCblWQP/VhXhlYGbf3nD8
CZjqflcqPXUsyxoUltKOMMzAli26vv80t8bOkJ/c7anlrlEvvTFHx2NArlUSZCs7
aZlPwYuOw6PNqpw3tRFJqjENPZ1/KRTuij3ow1lhrtOAWF8AZAVcg8patF1FgHA9
8bmtt39M07EZAkZLVZE8A6ADk02jkrL1vHR7nm6a7h+p7m8fBWBAvzo+5YQ78PeB
jp+SIff65VMOoU/ykDZ00f0ig687JhNgrUCX8O7acJJNO9cXRbzD/o11P6kK3DfO
pv1NEaH7Mxpjn81TklNoC+Q1sEDWrMx0WIHgTszSRUN9Fn4oXV5A8XfGiz9O3Y20
zTmHhNEeVW8emBHCVD4W5W8egPVtUcMnp4Nb03fN726MMhR/yOVIgN7elN8fWNGJ
ZP46irAVJdllpZslUSRmCngpnTIyxg7otV+K5GTki8/inh1iVeDy1hm79qT53h2i
7uxsJSim4ox6jdfXBCkUt6eIbGuz5qEdzjxnkQi7rIhWQ/vTrK7wbhpKgDtRFyGX
mkZ7+J0ylJzsRptVJKccVeCHS5zKyhDTgNDQSkQGHrsHW/dEbDZE/tBXuS4unTug
NSlgapyhLguJ+1lSWWWO/J4FJA35WAN+EkqAwxcizslZpvoC0M9TEMq78qAOn/jl
wAtZhQbuSReflc8MosFt1jqVdlpxp+edDCpyAJ7G3uOCR9LFUJ3MK7crVSiF1/7o
GcFyf/ITWAGXqRa3mHHHxsIketZR/kHBCFQXNkcb1iZRaChFd+xB2oVOLACdXqPx
HtuveMcxYgNnv1Rz7kkk3zOKsVCBqE5qO9h9V6oWbbgAl1VrGNGpPzEOJuh5YQCN
m4FejAgsiFrpdwxhXvWEbRXztNY0aTEkaFxUhetuW0IQARWyS9SB7d/t+Jz2WdTP
RV/DN+6V7WM3OaDMAhtXxmtLkpX6gEQNQ2x3WbxTcAZIHF7BV72Tb6s76CME5+WR
6pj49oIxZD+SsYLzOsOs/Iw5XIfjXSCKULk4rsh9rh58Nr3TWOuAv5MC+aA6JfRl
mYvn9Ntudxx1XzQaU5057CfkOCqMRL6wcrGiXi65Tkfcag57gPP0sXnzasWVF2Qg
NQg3tPB6HTx0wxzFvZMF/VG0JHwmF0BF1KECdfrA/1JG1LdR4Db8o8RbT3z/cPXj
ozFpNZEjRyjxUmeEGuV4evVJNYHPGEtYlRNOlhH5ep/hd+LZHhi0ObbgiT0EZqlC
O57hUF/UCKHYE8+7fKdzblf/fNWjSqjqPrp7tS6Avm5gDdqm7UI27LrTYfuKr2Dm
Odx7GL+4o05asReFknICFYk+LRuG4mz/Gy8e/V/QJkITsKIjGSXE3jFb3L6bumQX
R9UL01RW8PqiUeniextw45bZO4TDHKYAuspiOFi4/7W3TTdO9Ly0R1+gDRE6QOin
5HntNBiU69hPEEt7C9EZe1GObfbGGOcPAe6mRayIxDq1StrmoCrLt6QgNamAI9cu
k8vNNMqUXLjD79ZrKgsw/IJAdMvWW24ckvMC9b2UJYirxeYF41ToaxWyoGpb3PIJ
FxEkpte4knshsbtAtXQtmFIhnbS3KyboscTfS9VKfa1IYMlBYYezUy3/6yj2O/3h
ehdi6NEvETfy/BCRevCV14LMAiE0IaOwfFn7oWoOOuf0tJVR+jCf8Yxa9xi4iR6Z
95jOD3hOtQ5iFHO+CtEtR9Djar2SA5NfGuXDai9WZAX8gzZ/j6tlIprxfJ4R1gyL
tiCvV0uog7X3vVUafzZveUgPDq42jD1t60iLTEoXJOIOilVh3pHIDAWnKRu9KN3p
2hahACzQ9OYYuZZXMnrNTSnVZnOnsTmP7HyzzGUlM7zxfNsK/4crxVZvhCcCJmHC
focrx2hUblu36GAQF8n2uhe7Q1V3dSZOLpCzjLThnDXZBoOJ3TgjhOzi554eN9Fs
iwoqjZAsc1RwuJwQyFui9VquUDn0YFWJ/fIn16Ab5W5fTMFlquyX9y/ingBlB6XY
Urs5l0qO1PYafgth5BrwIVo4+/fRkHGhR3etAzYdY8vmx6biYvgbKTPIe6gZlHKs
HRSmx6Dla3ecEbauxhPgW4zHRFDTHQD4egB0heK9sanx50kJWd992FGXzFgbCDPa
OXwSEma4zS8eANtFxR2mNtsFPf9XBxgu545v2/RYrQFXSKyDPaF4fUwI4abRcacN
RtUvFHEf5tIGyq2RrWFnPuEf4HkKbuOMK5nXt7hwoed/m0Qc7DMi2Jufhaq1MTTK
PFEXu9PHfPmm52fZRQFAOOjM5mEM9Eb61AdsyR4Ky7c0YTVLSRJ87EHDRzvnobSz
Inh5/4c/OeFv+rvO7Pu7LzYFvWaheXROCcHaoS5neE4NOqPudvdYOmnDFrcKLl2R
9OTuNiAouNSVNJ2Wh+sMcnkuB/Gakx38mmHxXBULqt61opVoDCDrkjen4g4QJsnA
Cx1wcPRExOLnZeGTnpgHsw9favwBON1qqNA0lkNrNSak96uHrjbVio+FSmlc78bi
kKanX7lCwQAajjzenwvTQepxxfpuquvmym8gVY0E7yNgHHRTnnbGQJz7TYBjUD4Y
oT3Vq2DyP/apqVcm6SWmVUNIHwf3dykfyx/tB+5FyJLMIJaSiBm1pY7d73Esj+WD
YZg29SEKLawP03VFNFbKT2IDj9r5Nk70zlVQ/UsxoXsAZuK+hiZnc6+c5U29HqDx
hW/OcSShf80Q9MdvXhxVAnSY3C6E8eTYcGOi3qQd/jSLCKCLGiEC8hJ4WIHQA7oa
eSEVFE4+vUZPjyUbb6EfFPQM1oC2W5Yko7wy/wnR5dowjnpdNwnd8mR+C+DUWvji
ktOsKp2JfiGphjuaDHu+0oTh2b0FnwvknRxi+zwzhIx0BT6TwacJjVy0kS4JDTe8
H/8B5jeBokT6cj/lqwExGHXqZZT7oXWzklL6pXCHnn7h0PELWG4vtmOXJ2U7zkYH
Vms0Pfz8Hp2DrapsDxOkrMHpSTWvKwk+VxTOy4kkwmUl5sSA3123tAJqNdtjliA0
Ls4JUw1qfmpGkCNWmmglHxBk0YlrNgCL5x6PQj8uHQTDW0BzZ5BZORSNWdve8uC7
qzwtBm6v3DCsluy6bCupVAwmLQOAYLwmlWqQFuiUyzbVi6G2O2AOeGplzIqCfAqB
IJ/eAqK/XMyfEgEpLTUssZ/BaANt3kYMEMfEpvJtr6MeJn7Ahy8z0kkryALZ1mQk
czrfyeBOYfMi23pBLbT41sgr6OxKnffNzmpgM9KiVD6JUPxmMSHGyAg9KKzk0dU4
GkucliNkLzwW/3JW1QHrWbS4K2f2II8fPcYjfLf+bNZjVv3pYsHnZ+R6AFNWnxTX
0sJY/C56QMKP/j6tcbSShTMezOb0LBkdl9z31fui3TfkoGnfpNQ6LkZuT/5QWfc9
DesqNuEFrgTjlFhAO8LQa/XCK5as6KSiu0FRCMPNNeyaoSdW6PyKJnHXtlGTTp4H
fy/w3iQPbsb0rJ/Mf8405x1jyMTMMgbNFqxW93ujCssYk/6PmVTwQkxrTZeIuvA9
yW++Llir/hjqbpmeG1cp4FhY+iGt3xzi4zMdQLRPAlNZiZ0Y+jcoyBPgUeKl+wdS
WNM52EUJK9QoX+m+l1E9ybncgFjM4NJHZSKMdfb7IMIA0j1m5wJvm1pTK7oY7c6r
uhenW8Xbkkihp5OaYrhXTCeP+DzkD1+kbooPwWSYNqsiedb2seElSxc6TUFv8Lgf
qF7qpAIMIr4ZOamv41G+1WKL6g1yvHPE6zLNAUwPTAI9gpLmsCH3T9Ki0ubzirrJ
cSziiUBSvVFrdnsxTcsAfcVCCFvyS4TR/kYXah2mlaknUdpGCDmR8NlP1JScfjdu
iPI6FclpWBoetqABUxBD3zl6PzDyFVhjAvjKTP5zvD+/cweV/ma2v0fxt8SMRPm5
YZ4RkKz6GIGQokElGnrnyKe5KkFuIMIGZFrp8jA+s0Duo5ZzMFFP2daNYk0duMih
k1A91DU20bg8oJIK8qWeiYevgzYbGwWxKARPj+0ObdnxQTmFdBLguKpqTpcp31+9
b4TsoPI+yuYBcBRrBRRXE+zeUynyn7vT74R137zoyFPx9AapBS66qTNA9z7HHLKp
dcEkgmi/Whd37faRNCz9ixWsfTXgNx2+ybrDn/1LEuFjc1L5MpXYygLxQhxat9Na
IobZzYhLA5L50KyuASihsIpiaJqyLdTQ2y2P0BKE0FLJ5gbXQtvCMo62Q9PyyoT4
+yiZXGsyGIsLCRSSFycZ3i/j8HYSlmj9KcfrS9A80Pj9z6cUgg1yBW3YQvQ47eVw
O0iX284wrkURvIuf1JQKABZDUGVggJBGncjH3jcNp2yKVJs0dsx37lRv1pw7fd6+
iGWlFlpb3q7SmhOH/8/UVr8lKOSO9EhjZFRtL82u+D1l2gRgl3egda773o+t6wdx
BcfdvFR2xn6Z7rTI+Ao3tgN7SGeDSIat1UZ8VN/vKc5pFnGDo4+y8lCJAd8LUwW6
Qj2S6rlBHC0DCxWIO3T53TDm7OzVrEuO5ceyVIzBaPXYUuIHethJTg4WhqMd6oo/
DBHHhP2WlJ0EYUaYuoI0tvdVlTVLYKTOJeDXXuZzdHMC/p3Xdlw97GsGTPFH1Qyh
Vmu0UEhxkiP7olusrETdJS5LH7DEBFJ2stiVZzxYDS5SfHOCIw0m3dqJDoT+zsKo
bWvngpQ78HZw+sNLEUL9vFWBmN4r4Vwj27eEwt075kHV8JjYi9dTesT4c03VjaTo
pa1n9GIg7MNj0Cl0iMHzCgTmFjVbpjCyKncLCjbslzCqqRZhk4Ox99dT2CdtBxUO
Nm/HdhfpJZ59z8NJWz5Nja9JPnnIy9ArlRoZ1kRvETTg7weKqqXobn7m5jJG0/96
8uHjLnU9RsvoChhRZ/gbzZ00+8FbfbmgRASZaE+cQ892xjFC1RdFoe7vK55kkA2a
SkQ3sg4CqRL7QMLURimi1uvtchG79T/xEcbdzxiTpMZqxIjBKbo4LHM0iDe4geZV
tYbXI8xIFVlN+mvk2oeo8nAA4zQWXVT+IFYuwomw0Gw21KLBxC2AbvvwEGx3GouY
vjN51KEkCQL4S29JCYUnbSPIuXGiO852lCQaenpcL9HlfNQGx49Uyof+yKpYkoat
DCZk3X2LWMgNDxTOYnGYjvKsxuCGCiGjhsIudHdygaZoUZVgc/2zO9fbbxaYz6vU
K4/lGitzxXzR5F/8rK+/l6pW2tIZKKVkPHcG0umI3EBn5LYFVYWti84M4V4UgyXg
alaccZtW3md4DkKvQYZPyKiCDh2i8Ti9ejW4Mk4rP7Nw0iOI7kRL9VdiZTDPTE5L
FwkuyD5g5Ls4NmdSIHXEGmnzy3aO0mATB+lbvjb2Jpm0E3HjmHrjRSztXCUG1dFC
Zavu7LiWVbZNIJuQC2+K5vpUuOY3oyB+4FrlM4mhYAeZBRCLY2qjUKNFFytatHbV
pEsh8kmfoBx6M6ju9j2AQmI8GWmV2NdJ3QXm1CjadrJsR3JKUqU3PubxuQNV0ikV
kZ59Cenm1Lz64zTxSB5gHIPv01qNGIww1g6digWB0yamlPKPTjnVnQpKhHJhx0PZ
UGHq9RleaBd0O2OPnEU7ftVwDDie2494EdCvdqu7ikRcEQ1t9ripV0WhBh0Sb+P+
u9d++NN8OoAGJS4HrqO+MFLeUC+L1jDE2YCJNjryUFql0BzxUITBaCoONY1SbpMd
TJGHI6eCcxwOTni28KE5beiwA2Z7waDWtv29NTREvGbsNXakHX5gMY+5BR+w6njZ
/pHj35BIwWvQrhgKWqQ5yqvDXaQWAU3nH7lW/Lq8161x1bYqegHwMPCglzjmA47l
4sgOuUiRRv1KCjoMyn0cgkiYYXmMsyFYLBoS789T2ESZ/LqFfUhelcnVZUx+3e7Y
YLhEZ8PLYdZEdeeXmfKFqsklnbkUJD9yNE8mqGkW1zX67hYVVzRbQ++l5Y6N3yPJ
dvo7lM6Wf8eWKBxzDxlKlVd8q7SQs43sMDG16MsL7GgV0DdK3ZDQ6Vrvf0az7Yaz
R9dxKvEPRzIrBJc47a0PJLpwTgtYuHD8zqtf4BhTyyOvtOe1GNf3SRNOnARNtsaQ
6D+yj8xIaZJU3HYjnGNyp4KbEqNz6Tsf8GXB7vBR9lsM7VGW8zTk1XxMa2XCypRq
7HlRvy2ZTkSYet8i1F4xW0ygpQS8zFibziwE0QK+X4IaD9z6FMkdIzXvbBnJY4Xx
3dZCTbIIcDFY7AayXSIxsrS9dFMyTPzE3HGZg1gaY0Xs+gMISTc5iCMbOnx3jJB9
0kIZc6hbdIR8r60qSXG+IEbgxlX5b5ncqQytYhY0TKxZdj32FUeq+bPsNsCXXObp
es4JjfJFS3CD5YeELZVN4sBXLyTmenOsFduEfhE6EQU2gxpi0dR7l10U0KSPf3nr
4XKSABqDVqFwbAsrhGS0usFzlNj2Q4FcdON2pY5FuTnYANo4w5Jt+AuapqsKeVrW
xKFfZ0IepkjTkXbpAmArxWgpuKFvYRTcA0zwGVEgxXTBTqOdo7kXZl7dx1JwMXV2
NQPIL2EIuo0vOBSNpK2Xnvt72ZrY3hHQXXcJuGSfOipw/vRoektoy66dz5cBst3N
6ePURoMw1LxJTU77bBprH3U8NmHyou4bbGO1gKOpbsg9h4uUK82OHbio30E8sXrK
fqJloJbhtkQ9fjIyzCqE2e6SFSYIB9AY8DFuwxQcNnEZZkemEyzXGvCJcsYAR9IP
e8klplweqWKKsI1hqmERb8oqH0tWunLmrwJH12tp/gLub1Z53efe7sFDR5+ozrXi
r22Ql/xQ4vccKCzEQwYutZlod9MrDsG2BCM2Jo9J6piHhUqTeWxQMZ21TqFbTd4k
9KfnxvXJafqu+GFD78fXjC1aCQMlHsTibfcvYS6v3/IaJfxLeUwlQD2gCA+gSN6i
7RMshThQCVspF0r4mN2TvNewgt5a4N63mtHoJwrjZQbkoWZY6Kypcz/WeaJu6aae
4RY+vAKGd4hVddY4evXLNjY8na9B1EkqHHXF3rzCegwEo2RwzEaxkMAKcJyCEX9F
7YzygTB2Y8iedlITkL31FbVdS/SVQAr5Bi8WNV1fXB2fuR8wCVq33jsjMy6fPe4w
Nek8k9wuyT4g5FMWNzDYh8qnlQaQazfCJyjM0qnY0GBV1PVJ05Kc4CnGztOAFtTQ
H3V1pjrJBpqg2MRkilMyUbEjlv8teJkZ0tqMPx2SD8UVONKLil9dvsLjmN62p4i5
u7PYbFyjEKUZlHYd0dTxroCa6TUVlFmerKtZR9BrZ3ULRoj5asMNwEEHNO1AUEwY
n/3Yw6FerdxXJL5wnoE51HRIr8V6iNgJJwy/3g6uWCFtlpsNbvZUWgCnFkxc18si
aNkFpVgk0WRix9v1AaB54Ygr8Et08FyxnVKZxd6SApe2CPVQiNXRfOgshmDShUlI
zH9uiEfQLEZtjGLBqf3ZheQLtSNfi77IoBeq5tCt38AnI8/5uC3xfyScS1dpx7GY
QRYdeD64/zwbTB9iVDtNsqkiXD0n7PWoJxkowMckcrYaDAv/OzIBVc0LcyKddUqN
A0Sspk3HNYWjBSqSsucSwXLNK7vgc251GBf90YmU98g39UrHWouVNzRFlWfyxj0I
yHDHot1/6zGS33mlIE4xr93zqGC0eezokV09tp3UGT/uVYMqLxrIs8NEAaW81Kuh
TL3f4D3XnKONIiQC2FDVehHMSoEuEB590kt8Om7Z3U5byKfFGZsVJ9L5zZ8jVbBq
stTBt/I+sERuyl9/9QKF6firhaazZBsCrbfDNI/Xik/8wVufJV9cNqETvu8JfHfe
uTlQVrklBwd91r/yNlZksMpw0fQLzvAb6zhfmhC8/M/hveV/pcrkh6CZ7ySBVzxo
XVIiHJlt+Z4nTrYYCC9sSLi/F2KaVka/t7x7XKF6jIz7YuyXvYl5fzMHx6fPTlJQ
nXDh2t4k0FBY3+unOk7FRaSR8z4wHawRAQUQhPdkXisU6+Bag67e0vvl6Z73j2GY
iRipk8yFHB+EFGK914U1PUUTLCh4rOjRAPVDAHd3OpL2AJ9u7IjCPPiY9Y4C5gjY
R9Ti6kq+xH4cq2OxJj3220kN5N9KsSON4hIiprmB3gTXCBq+WEjs9Xf9XLYSyHbV
fEJYwxXGkTjYI2WOcIQKtBrNvOHLjPy/5Otvtc+YspZb7GO6mood66pw8c37iFtT
Dr+vP2kuKWoJdzyASecG+MIXLEmEQlolhKMNVbDFqgbgsyvIEloia5gJKZ5nZZfW
f/I/0krkMKqlKhaN6GabVMaOUSlLOcdjk3LfnZjO6zEJZQcBb57Eo1bnOGUtQAPl
6bHvOr0ToeEPx+R70dFIzzq8V1WP6KHUs2uYQJHsHi1SKUpHIPA564KDMDgpsBFj
RQIogu1ZlY2t1ythxNndhhFTAFi/P1OQNyzAxj1+fWdKRoO5ahzxihrTXHY2GPV1
WYhpbBGcmyIqfJXB33wyBGPfSF6mZX0mJoAROf6rrEPkA/eq9G7o+e1go5O5TN4c
NuWkRmKWnQqwuToF58QiRkgK84/lEHiwftgI4pf8eJLcb+wR0pFYIkqAM1efRv70
r19icNB+WajO9GvNsa2FEmwgtThsfhZKJACLkgBLrAz01XEv5CRCyNZwxCHgbAfi
Gy1csKj8qUuKJc2An6pJWn+KxSiGzf6vOjBf3CCCf6OUYEj5DLxBKeklRvV2Uq2K
imHcLv+ko2pB8VB5BE+iKgL7pFo4ncT1YtvAXzSfhm6KCwFv/rC87AxB4zCw9wOi
WN6gvP/jgMHkbo1pslyQFz0hRWmYDOKfg32UmCxchJ8Ihj2K98x9wQTxL4G4Rxl2
IXL2JHM0UD30kPUswDSCtViay5YsjhqPW4WLDfI04HDUbATI7WaGAmBn7M5VzriA
7ezuyR0Vy3KPKcr7G8OF9zTOzdv2xy3Gm1vSwlE+mmW80Oa98enahla9Zerf7lTT
53Bppt2GvmtQgVW2QTd8F9/W+F4dPzRZwDFNb7fziagoUYGD3j3DOhST01StSJd0
BRsM84OAPQR3/gBjQqrP6+hC5D5FMe0PmEjl/u5zPtv0Obo52rar+15zjpsG80Hg
dUTvj0Z6GyBrOzIYTd9DxXeDa3aZj5bdZzuuharaNfZof7gZTRsDfgyVezQvnorC
KYi44m7zA00YtaujRDI1TC4qEYjUwfhwrglxgpNQ6w27xy6x2noPUIUvLPRJ3s5x
bSaaKM/I7cX3Bx+1/mnEx51aq/FHGMRAKY6oFnjvIrMctrAIUMpdDZ6ouNixs6qs
pZ4DPxFsw4d4JZHnyd1FjIGaOYQdT3KEHNuCqRfY0HNwi2rYhLIvkQSHex00eHTS
mFTvLtZg4XRjZ+34EVby6PPV2QghmSqjboSWcoNbCP1thliumjvXzLVgdWty2/Dc
xOgJr9kx9ZM8Xg12L1JFZ5G8HV5rZlTTWAPUyk21ZdHqGZ2e85Le2GpTkqns4Ahf
qLl/H2b19Bcyep97FI4Wht+b33QNaG9lMbSynPszEPxxKpjuyjNNk2Qk//w/99d0
39p/W0Fwv2O3JeVsjCQYgpwj5cPXEznHeMeKoaJqttCTDB4OxIFPfzjUe9MZS0+a
AN7uP0dQ197f3mDEJV2aDQGZFA+7TXnREVpqC/h/BROgiqc8ipjZCxpjtVYPcdp+
RCEqW360B9Hv8jXk6vmiK8z+3kY6xTic9M0FyiLmFg5DLTQaB7NQLVMnMGy0zgy5
WclQ8woWEZSa54WngeqxMQwJ0sIWz0rIFWoCFI55JqGpYWN610XlT19vGdn0LTPz
GXuH0oKCmbrr8J8LSDNaHSdgenIdIdXSLfghZtfBVChzhMTjfsWfaXzexNqkSmWp
INTbn8iMuXbbwREXuqvUQfANx2ovTABI4XRuuijexyac/SuPvONkTzxE1cyOEFSN
efwlIvlSPb4TWO+CrB3feb6w7UMKHQ9IuPFC2kyj8LiKce42pU92Jsu60/pEaWeI
rf1fm+JwDq757OIpbmLl7qfwNFmxkc0s3ztSukPFA2uev7i7XpQ14gOBn316Nb5O
1xhCSKRQD8zODSJYFhr8hC5IAItOObtxefwsPVtzoItl3nAI3QCgh2t8glAjK2Ci
gdGPk8bji2O9AHrwTfulaKvVk3oF7ELJv1cAcE7yj0hogxn0oPaeaxsRAvgdY048
Je6HxEUcsuF9+nFvnzMAXfOAeT3AsbE0suR3rBsho1DxMQDmNGxLipGjbNbbstCx
ptYqp+A6jxte45bjzAoEnFc7c4TedRWlAOrfRiMnxlz9w932lOC+dcC6TtXgvxxL
ST93ZlxV+kQ3XA4wr38utbmdbnN1CogbHeXVipFD7TJHXI9id+W0AUoMWDWuFwOs
2d8H6P2UVjyRq+K7nRqUfkpg8aO421faceljzr1JZ5rNhHJ3OD6zmTBOXGvR85n3
jG2CGRSTDJN1igsKVg/3yRcmkINxrU1D3ELhRaXMMbPt11LMxvysbUXmI9wpQ6ll
DRtZkncu6D+yl0HAo5AepOVQMjE4chKzn9ZhOhDHqNyRz5A/tYF0SSaEDBmQRp+T
9n8JjvTDYfF5oU8YcpPg2JOhV3YKiQcIsS5S7XzAvg83Wb8iJnxUWXtHvZN2eoE+
J6N94TJZ0yKb3kUNSXQevf/yGEwVdqpgI3u0390JKsf7hMHf+deZGh+z/v5NwMlW
E3KElQXIRDIO1BOi2rTEUs1LbbWhDXphsxsDxuuKzdyADiaaxFMcn+x7HaR6/VJ6
pSreQe14Vleh6kV1ueVIoTlPhWC31faAVCP4hSVrQXatM8XyWWstH4pA5AIMExtY
j0rcxE/BQROx+B43u2pQDPxCasNi4AKqv+Q48g4k7Dj3Hp9Z5U29t93lymVc6uat
JOMDtf1057vWz3FY7/G4ZFpVo0YmQGuqyq4hTAQ3WJJkU/5EOVvPDfIb/xx1pnC6
AqI6ti623MeqlcAHv8IYEUQwVqEzKf5ZjhQfPn7L3YutZcd8oi+nC4G/kfUwhWGQ
oG2Ip3Kh3ZLxfzGqCZhx71JialLPgPZNq5h7f5NO1jVPBZOgqlDDt+OpSYFOwuU0
fPPQ42QL/Obq7WFTEYeqyKOgQm/ROH8OwoNRjtAfTxlqzjQF8CMHSr+T4M79O4Nm
yeRdpZm3xIsBwopZ11jYML8baEioZ/Rq2fTy6Nfh+iQaD0pAHY3X7aYL3fysVNSL
ZVr70O8QoEbTSLHUxVbfrGKAmvmTRmPC6xoJMz99yZjeQunR9mEpafc7IWrBVEiT
aLys6yVuUknrMJtrZg6rQhsgUILOWXaZcn2ngLNIo8XyU9IlE0IfkuBH9xhwZXoM
rioObuLqtLRA6QkMQv78XqW0nYlk6pRWZB9u2HTBP5I9n1+MDkMJnNTgH3Yd2knf
c6WDLKh+QcmffMmmN2Dgbo/nFr7llR8aKFJjscCckFbL+Sc5AsNJJBzjFykRKeB6
2ag7ibP3K6LE78lMrHCbUx7hU1ydJsbAddVkBSzVLgf+U05LIrZFkEkv8s/Nu2Ru
lssdbFNBT56pRsWR8q/3jtoub/QMyeK7VowF4jvuwmSGj+NS+jwJvPQVEdsxC4RT
EENi0UQfJhdu2Aq4cFfwJcD0QbUtwL3fxqDEkHCfJXcHfyKqt6v5H3brTXMyO4qW
NsXiSgU7VdNH0z47a8BdBPqYvUAixiM7fpDNw8Wv5/vNa+0d+9koxmgHgWTNvjtP
twTxRJIG1PeKsC9d2jow364xeqBLnMXsBBUPNnt38hXB8q9/ItGj+CvZOOFg1RkV
s2OZ5hdy3Dy00dQKrVmN4Q6Kcsku6GJWrvDr78ncBHQ5hJaqK4/aJHbfD6XJdGJq
UL3f7KN8ePFM0Joo76xTW2NhanzOHJkzYS706Q30bo8uBUOMSAeSMrhyShR8hpn5
JUfLojkYXy7a6eqoIH16df3p2uRan0WG9ZO9eSSLsaSLe/QfNtg7KF25BEy8ZrIb
g0LO4++R4AKvTCK57QEM+iRocQ/ONyOWWyK5O1cFRAqOuXJB7ZfJpn7d0i6ov3jD
iTEFTgd6NFvGdcjVyIEYlqCikzoEXNXHuHqcOkixrDDNOs4PH3AXg8TyVEwDH6u2
f84vX31I9QNRUcZIxTwmLsor9lM4ooT6grkSS1Ca9MyktSONO8waWO2qkw2zHTMr
TgDe5cm/4TeZpNNgoU66ZEyL7LJxLbjAftsLJw99w6g1YUWVi8L5AypxGpBN5T4B
1vPKilia+bzNST8MRiFNQy7O1E5Gs2fUrHOPQ5oLb28JMq3FlVVxx74AhqnADLEN
4PNSBa9wIlNJiLbCuhZC2U+AWJGI99S81gAZid4LA+Iyxh2ptNd9145EwFUXtidQ
ps6iiJO1LWY9/QCCETh7MGm+kGs8sRDrBrR3SpaVoteSRIKpyU4Oi7RbDFUTuM8f
p3054Nf7RH/ptkBNftD6khcaXGaN/K8s5fDJoMwufRIRiHyHk7iQASMTN5pas235
g6P9cp88B/doXBWkiMhj16FFEb0I2o29YWAqxv3PMUZPzz+njexYnyyVQnZfBX3o
vfTO6kOSbAvReECK9vtcLFbur6xUf9anjOJ9zxnfsQ8wd20QGVcbOqIvmpHkcXI0
SEPI3KkydfyiTNUp2lxfn0xM+L7yo/irTY5sq11kiCAst9pd30Ft+/U8MD/ga3+v
P9kS3K0cnNC+lrVwQcr1GKbbcAksXsP/IM/5Ijnlr0D/AG4RyPuYFoyxNXT7b9YR
V8zlhtNEeEyY8bfdidQ/nndPL3rPekwL5GpFIy7UJkVQDs/HEETGpbBAjf3PCIa0
9CTK0ZMgQgIjAOZVu1nrvUK4RtyVAQcwEYnUE3Df/TifOpc3YPkjT6+RhBk18ADV
PYhQt2hVO/oQiF4iWtkxuG8/3VHRJE/EXeSUL13VW4tO7PGsCZR1+044B+cHvwvE
QiaKyT4qaKPUjW06OuLNTZ1ezXZFZgl12vn9eUiFH0SPETj3mcxd8N35bWbg0FVf
Rfg2dVkhjxFhtit0tj5cnkqL73Ea0G+ynAVj62OgT/8xR07XbjBT93QIi+m1m8gw
RqNK1ExADUpOeEdQU2HWOIpYhZc1Tf3debf2P2ORMIOU74s82eT1YCfwL60fgiMF
ofrD6FUDWd7aAt3D5ALo3lANSWW12j45tV8st/WeT2L0FksxbpIfHCi17y6cAF77
oHSOqQiGvBezWRkVOin2zG9ep6JRjkai46U1bNZZtA1e2REb3OsPKNvSQfwLrGjz
Ezw5JLFTy1zBm+XJj+fkuwQyne6oXrudC8u3kTwCIAqNaLERq83Bz1o7hOXITEPO
WO5l6/5yX39EhLNntQrTCZ1+mlMdn+2rUagqnxLn4abwG+yeJKGDC5Bkw1GD7ORZ
jRkoCYOtDLPFF45Ovjb4HDpyg4DpnfkYY1p6m6S2imem6DMwhlVB67XAnOMTy4G9
i2PvkX8Azx7q/wqKb4zkW87arIaIzkKOkkrfwCuFzJ0aYlAAi5RorqC2ChYAuxjN
VEOF9sClrLW7DeVVfmDo5EsGpyVWTdXsTvlt7bGLIHC66A1sHyFqn2wexLTWpKVT
m8elkQ73zX8++cCBulQBTQl0VpabSg8oWxoiOlZXdzatJdRjqGSvlwm+4XEYXm7g
Td/G2VWU/Q2NdYbwLs9P3O10z5TpvBUoews8g4kJVxTsDTupzkOM7+qkvVqrqOoG
uhtxmhmCp9xaLVvniSzJiWCKgKJj+PVuegl3eP7BXJiCNaSvaca30PSqvjIyYgxi
g7qleyh8jG2zH4UzoCKs2OZ4Nv2Qeml815SYEvYncflK/r0aWNqDpBOU63i+XlrX
EioI6MctZp3tNurUlGsGDpLsHz+kay3rNVf0K0mHCT/gdSES3xRRn0HIQJVrKlDk
WnuvNKXTAYW3YOED51PFFkiv76TM6+bBaUiTt7DL02ca+3riZ4pzKnvM/l+VNlKV
NQFn/JJOogDZ22uCBpfpcI76l4mFXiZrHu8B/YovslM2uJY8oWdC9uts0U5YDhB+
Op9t9ZB01PD1nFtinyCk8m7X9I79oS5sxmTwz5nuYqeXWReOSgnHhyKs8/e8mVV/
OHN+3si24KX/YL+kt3rSKGB4pM202wUsrAX6ub+lSdtP8VpEZ5GsaZ11layo6iA7
t1YELcyDcStLW/dkYsT1gifA1qljCHdQcs33rywx+wUrfVyLg5Kp6P2xFPGsDodN
kzFx4xloKihjpcBGVznsvuxbslxBx26sSHwiuDDqggWP6b1T4V6uch1kG09mFcGt
dfHsT8BvXH+cPo1SyhQdknI/DpJWiA134zSPXxHmUw6DnYATGfDpWjDRxSEpPI+d
TT0qs6fkF/zqpkScVsNPqAZgAZUXV6+bz5Z2OT343kVkidhHV++DhhyABmQW3grg
MZxY0fJp8yhFRvz+I4jWUoJLs46ZklCsL94vQ5pqB8m3wrflylyyETPfkBKjDyC3
r2iTnrAnDlZ8R2+hqwWUrTYUvfbpJkZPAZ3iAgx40UiSrRGZC8le9G+YzhaHgkQF
afs5/ATMWxS22OWrRKegUF2HAv7stB2bhvOGs0xVBzHWZzPK5y7dmJGJYpKybgXv
YvvdS11kRTx90Df31kVVi4whyB0CaJmNdCEQgymX+AX/F1thZcnE7a/Em9Hir3uU
dn4a9AvSSKNyNzIPZKYFWSDKuUNrfabZL7gKerQlaIL4ITizsBwwaZuU6icNzJlA
+68lbt5M4JqK9rBZvaVZ1jnYarmAPvVR9ZYcqiThKhKfmlHwUOHbG5QDxR0rv8xg
of+sH4+oj7z7iGK5TFf/5J0FSVZedtRQkm99QO0iLa7rx3x28mPE+wkGs8a73DI4
08ybRJK+APU+2g6Dps5KrUhaCzYi/57JkbnUU0wCtQKRqQ54atAGglnzRqvpGeNc
06JrTHyUydTALKK2TWxVM3YO8MlVZHOzHrXTcO1iGgAqNNebAp5Ii5edIu67Qi73
zz87xloepk1EfFKbKHkuGn/9UOrwcnN7KlDlCfZFmGNWHWW3xC2rsOG6+u+tEu4Y
F6ZsUDBcJdsjN2+l+zgLNvacFrvQ1SLooAwlVEYJIWWWFIoiECGB47HOZ03V106l
bPd7/+nuXSwdXaZEyWGWuHgcVr/fgbMC5OwjfOIvfT7RFkKaG+dTIvuQn2bAIFFM
SDf0bbLaJKRekmbegvraljKK2G9NDZEskfZrHMrHm76PGENg4sbnLydlaBRyna6A
lPtKsJoP56foUfh5IMQhg31Ywwq9bA+C/UQKvy68g7BivLfU/OBKHU6ztslLxwsI
i/D291gmZlLkwzTYN7eRJ/CHb2EBlkyfJVTq/PCXlsoOs5s7D1SPk0U5Nk3NM7Lp
kQtPPrl7CrLTQYiu9adeYG4shjSzvVMCG4hr1UEKcJXe0JX2fdiWknvCn7RoETnt
Rjw+809cxohUKWuuhLKc2uU6KmbNPlIZCbIXKuIZnAmjSfB3ziop2Lvl0JFVJIQL
koCFL73Sr+kZvnNwSo4q70uWgIDaCxambagOq5JYkYVothhxMCP7E6obutGdaCTT
ORhr/FYn3MYQRNHWiTMJAW1LZK8m9WD0aXUI5+RNg+Roy5YKkXE0oIyp1IJJ/Uvj
LUej0+RE9eXRJEzIgVxvwpUNDmsLHXwlrkb0Q5/a24fuPNsyMur0Ppbgwq49xRkm
SDNFOi+fRklYD1Iu+XsZ/t+wmpqg0yCE7Xz6V47L4EPhHhz4f5dWpeqCos6uCGi5
iSmtpstdKkLfJbo0uT1pX1gBMo8zzrrr0TI6LVlrzx73u57ObTmcM2tLQvyHSTZ5
Z/21dYR+eIOzTpL/eGkllUk6+rswH/x/Qm7iJdQLjfVpx0FvURd0HI7OWXT3cVwN
pBKyJbbfNRqtPe8Up8WKqbPgAsqje3EzKT6OClSMb/OJ6gdFBn0sXcR2CycZ2Eb4
vmQz1kSXC5vONKyNDGwA8y38n4VgA2yHo6XEUI4eBIBOgA/WqmK/Bl7KfQ+I1DC5
N4hD7xTu7JUkH9dL2WHT5NLKP6ySPKTAbKI1ZIc/AvOw1ut7/HG30fj1yS8SksrH
mowjHrdWkbWcgqKomgC8aHcOT3iUj5PmrtaqYQOkJ5foiMLbCjLhA1WPgwJ7EiGr
hI47Osg88HBnAV4vWhmGGxV3FCgEj9W1J0ZIpZG9j9ROF9bBzBl/WYcdVIcFBdWa
raAnlbMy3kb/PKZr4nTyFVWs0S/s/5sylL1TIvVp5n7Lt2PMcJjS48A5cxfRId+u
Z4drgoGhdjDFUjJ0FwP682axEEq6mM+fu+Mf3/xGenM9H6ql3jk+HARn7QDy+tjL
EYV4DXoM7pCci1OZLKBJuK9qmKpgTnlQxI1xIf6nzMANRdyCk+G9l/6uAW6i9oOY
Un+DQzHuL+n6WTIKwmiQwbe/l1cOkOUTpHCj7WvTYsAR4/4GfdyuSCtAsQ/UEsX8
8PoKTq6bpPxfsBGehjxogEsMjL7VW68FlXYHJqMv29X/YmzIF/wyBBfGVysZvak3
YgriDP5wUt+C6n7fYmQaq5F/xn9+UTjph1vBYACfpIvbX5MNnoFX27H9VSX2qU1B
PJP33x0fFYNXgxbRBVEMz0YuBZTzp7PEUtUY4WCH3oMrYnKiJiIDbaZLpcS02vQT
Uf1yxgyL1O/MgJPfOc5D7Zx3bOZyHEJyfnrSUp5wSBNmifP06GEbnVgOWoloiWw3
gTht2WGtP+quvWYI3WNRfoWDIlTVn/6tvVy85Wib0DWAJmcg5S1vQ3be5XUdHj49
XetwAWZvgSC43EAoj+9eZhEDP2T5VIMTa9xqCibyLkuyTXu5xKI6Wqa7svakN798
kDX0G+EduoUI/0UeYH7ZgUheHA1bByn4dNzl5HD8lclgcwz+xdfB5wT3ypiXyKxN
cdHU9iaIvCR13RV4nT/mHesd4wGMvwONBQbQF51njy27/cvN60A10T0fwoUO2tl+
ZJi+olRpQ1/bJADDxMCfCCEJR/+xdiiyY8EnQuRgVfTcS7AGyUS1g8isQIRX9CI1
vzLasEhqTniyJLgJUPvdALNqX7F/VvMGpqazMVQ79Pr/afeePX/eY0f5YSD+doXS
fP43imCak5iYo3TJBMgxwt5G9ORQrmCt/SRgZ2bp/ma1IUE20Tf0lElo4syBtPY0
NewkrlpejgiAJMLU4zvYEtYVWlTs0xFSiIPU6wuqshJnmWoNHq6XBnAq65ID0QRT
Tq2lRq1t5CU1BhTDKjfBGAMln2j3iRGcrB7oH3cIZXnBS+M91gUXpuTU25qA3xtM
M9g0lC0g38q+nmhrgpdoqp413TI3vpjrENsU5ydGMv/u30ax91tIVH4QzmNTzo8v
xVO9m31iCUveOmAox0rL2wpUBzukg2ZJW2zJJMJ+QyKqM73liRHsD3zc+WMBQJW+
CD47jTwnSk/kUedT/uM22SfO8jTuZUq+EGQKu+92qjJbPYlwbR8MU0rGSAoOlZKV
wEUnC7Q97U49dCZrvoHYKZkzA3PHqOfndOKFBTPxbD1osw/cBJ3fWoo2NKmeXpxQ
jrXrI84CqzlapCsnqwlRZ5ZqbtC8q/Rytu5X+LIru97hFzKHft7Hgw5GSirRX4jJ
rWBktLBmEwcCCAyfp1A2vz1fgAWvws7BS4FrM7HvwL+5rShlxf0nqZtbjPEnkWbn
ENwzlHhnXWiUvc8A/YVMueKKAulSCVU3rJaT08UhGNjDo5B+m3DMxNH71lTknQIp
bIK304+EK/GXzXQt8MSxM0KMbe2fKGDtPKyUn3dBdDioZ7N/1bNGaIi+PIZsX9eS
8SrQ35Xykbi4tgVPd2EfiVxJIo9/JqIlgpYm0ImzctTPcMErFbVNS8DjXdC/DT8B
8NbVeU7SSkRLpuREDpGbM7hb0u2dQbQMfJRrTEwAWNH9qeszBsDIExnqRnTjf2n4
FXbJIW4L9yCBNKGN8Y4TRJUAUcIFveJRATKRRKnBrzcooBvXz9Llyaw/RlN8fYPX
WaD/opeWyybQYSrcDNp1LSxxmXs5l1KKmXWZj/MwJBgdAGnc+89SYsAafYjUw3Wc
MovkeRrrah/rRrzGP4Yk9Xk4HzzFJM9hbrESANOrNPDvTKhzoDK1DEpSrfP37qti
5dc1+Dv9rE+RqOj4UCS6YMTaLoVfmlH3CRiPLlVPTuXyv8ll3G3o6Dz5tf88ffnb
Jb7COcFG8fMO9WzKy5yFoKUCakPKCSoqrISc58kvnhMyCZbIPT0gVOJAlmtD3Pjn
QGHxZUy5ddlAfMmAIYWpalozLsHO0WNO6XVSoDxaHOeogteYvx6hovXZcS61oBIo
SCvbWUkd5ndWgRaJ5K9+FoqQ2GPnq7EmhQPIgjuTJhhZ3Hlc8j3mHpN/D8lyv7bS
YnrTg6BtBUwaBPRfPQphEOcjJkfN2MqH828uNMzFZbxxW2hSN1StHNxJqp1s8JRf
GxW+ogUUDCS/usI0HsHM1o92o9LO9sV4//NNz/d0aMkWYF1I1o9NXu+/lZT2NV0Y
W8SQqYyaMOSaILn6iFrEV0XEUf+/hAA4cNP1e+/1BExecmN/cAwwQs1qt7yJjB9s
Qn+9VwQ/soTl/SSVckZlz0FNsw1LGGojabLfm+qN+fuEMylhhur0TtpOg+j6NjLc
YdJks5kHz6IhPJWbJuFuN7KzmmfYM1MlYiVzVQFAtb7fNaVyFs5FG6eH6E8vq7U3
lEra7qxw/fs+Wtw5Rs2enPJMbrLplHCrlAyNj9O0UuJ5JpCPCW0/IO2F0ydrTLK9
d5Wxi5exopexFE6dA9hq3TK3lytpaCcrQr3VfJAVdxA2rAW6Cj/zpg6l/PzRCeDP
SqtmIeCzgqtUmuhs4Dx3GR0fo07k8p66jH1aawSiDow+czq9tmdbHeSLJdgGrTKw
VnTFfVWzNGEdzZvjbyjyJQwMANN3hqn67/s0G1/ZyAZH11GFFdAwFJxSED9WBJF4
o3bnurTPlFnsBA1tow5A3qEHmv+j22hz5+cAZHW+Ju2ddbMJXncKrAVwhnJ4qmuM
9YPKIVFtMeBbO3vVNjN8SBFnSPFi9tWBIYlUe3TrzEJ3xqfeTGXB8IRmGhmwIb9d
4CNluonXwEpUbvswM99aT0CZXmgfl24lcQzcL5Tu3Q/gtSWQMtABK206iDdw/GKA
uzcPnXNTu9E2PqKZ1LPnTXLGbwgPMLrpBuBZaZJpUXsNMsKjnw2i6oGHa0AszeeH
b6zUQ7t+K5RAX7QZfrX+okgRczXMo8zEDVXx+ZYjF7vrAwhOQ1/WcfhtX7lSvEMt
3EeKAojEnA8px8lGyLxSRPXjEIKo8TqkvonnUbRaNMd8Cgino2eor6CBu+wyfLN/
cYCt6+jBvmuV8t7ndaT7XOxtNXOrwbB2aiPIcWqyPr3T/EBpHkxyaqsljmTGYq8Y
2LWiMWA/vsvZ3qZiG4dkR2Lgoj6i2cka/Xq9fBn5bfI/9rX/l+HWevWMxJRHdqLH
Rlyt1DTIIssq/sPSSzRnbZbXVp2n97U3j/6EqOSox6B4fcwk2xSp6zTy8QP71ZAY
XsIJHyB58UWMBaf17C+ftd1kLQF7YDO6zxoVddbYPUCBy7KoTep0R28avU/EVQfV
DHIhmmXin7fEKs5BX1Xejgh5lIb2EE7JMxHOvenkeHFC2Uxt4ZnCzMroCAFXPtmV
eFCyjSeWnKciJG3JNG4xywX36fTRErN/O/jr0c+kGmvllYhn/he4p6fmg/pDyHEu
0XWC/xATna2vSPTaN+CLumjKaRn6FzUPOzmuaXhvHZHSyNwIAG/eoJ5E9VcHbfh+
rFW5Ke5+G6L9gTFKnpESKZ0AbOggPIabMrdHTf8YIsd96PXTQ4psTVilvdJHgrZL
TO4Y94Lg/Uq6hl/Vo5qwg0aIKlQSoG06Rrs35n32xtpah+MCtU3KOwyNPzJSI1y2
rkDSWjbuSVmWjaeNIgJ1wd/1ti5UdrxxlrORtBvBHkXGekvBB3cpMpkBvqrlqAR8
GtLuCRCTMFnRtT7IOPlM8K8YzU5eiWVEr3g9CVvJLLWnss3+Bhr5Xyfnq7o3I6tj
awYUdSGYX8/zOv0hrsYwCl2uFiwr9AozJFKfPlA+NMa2TSwaZzbqiQNuvK3FXEgR
oWkYTlgTB7ndO/uV7+sIFPcIE+Yp96U6ywN6UXg6n9blW7NXpAiOs0JjnZcJwpuY
iRFv8h9dgPni6stIFNYy3Kk+FePDjbrblglYO9oc+IqCGDS8M5jqouTa2WdZSBPI
Dgjwq+a4blmWcqc4x6XNpJxiFMD4mgEB7dORu0UTBoMIGGuDtdeTJtrjq2E/nnEr
47dt7Hods3Lqw/4geipmG+bHbz0lh7UuzWHRoltQJkF4Fbw0k4K0FSrRf0Xv6yfZ
yAHTOBaWKQRmkOdiN68SUOEMXhBXwCoF9n6YgLAyNz74+vYf0Q9ztCUoVUautvo3
AzlfTPTkFXe7CorNnTBxopiTn+mu8ePQ2RQ5vZ8h2RxbZ0d4wcs9PKMzf+xcl8mj
Ocpkbcb0fnN9RBIIljEJwhCsnI/TN+LkTOoX3Y3t8uQqSARUzNhe9KFEXOcGCreL
n3qhqT+U+Tq8yexnCBJA+SUbs3d6uPcIIIO5uTPm/4wIvOtqdC4U6T0SVd4BaFnN
pahSBLM6syhfs7IC8P13NN0ZxlaeIUNQ3EJhpmekqyVvwIuqJJO3aNWsuy1kA29h
Rj1stvORAq3mYTZtIJAul20cVyPBtzZgK6+pFXWmc/27e+W0R3SRQ1ps6HozW3qe
CtXpu0X/7TezCuIVmMUFgY2oG5NckvUtNMgcXZT1en4SkaWo3Q2cUpxCgE/v1CRI
iz9rYesfi4b3D5UTGe694Nd1ENKy9/O7yo+SyieIrZgwJdxP/P0zykv/BqmoGxHE
RDEwGDXfbYjU1PZ56PIVLhibbUhjdIVfirOS5ecuQeyonmW2c3E4hzqAPpcY5eIO
B8fi7GaCrVrP6KyVG8xffExYHf0dJUeccUPVVUXPRzP3gyVBxc/wS4qXFCGw6IS1
WaXuwK4qM3g5SuTuUN7SKcexrarY14SH/cvbqv30HU8TvmSOeaHD8HlOL4VBuk5J
KbWhzg7fieO1FUjxldlm77C1GO2IxxB9FJr+fV0OKfyYKKIoqZQObsyq6a8cnSK1
LFk2dGqfKqaNV/4s4rdo/KeT6qfq8cYj894dNh6EGEW/b4WtV5q3H01l5cN4r18X
rtzDk5vwKKUERW0dC52/c6VcbONYGONhDriTF2PmQRWV0BrHX2YKYBdvQ1edlgHU
IOP/sLwpxjlkq6sRwqn2YmIinQ/HgqmtTzKiWWv3sWRqJiNA1phll5N4ycgXwR3D
Op+j3d30vppTJajt4zmDU3BPIMglUJTD+Ne8mhxFxzAdPGha045U/aMswk9gkpkf
W+IPySTH6u1CXjscsMTXBSasL375r6PtzYz7scFZ1p1x5bD4MTqyZRpwyUC5dBrL
MIsbf9Js94DpY0Z+b92SGiyME+tPde2YaWRBPMhiUKH2BQwnHxcagM5SUVbRBwHO
tEf+v1pY5ZONKsmQXoc2FVHpM40z4gJvx9MwSwbhlKDgO6NKP7W3FlyAvu8ERnXv
e4MGLFpXACXemZsojPkg8FWK2fVM/j+AdpWzvEL/ROQ7m5oXgcDzCpurvu95kj+N
a0q7PrQpeHoMcayOoxBU8f9uEieO6YSHHgTh4VPgMOtuPy2+q4Ry+Oi32r+/amg0
lGnlAtV5xwNCOK9Bmy9AHltDaMa1mEkFVVPBhs6dXlzfzCWqH3cw+sV1KJEF9Kdw
NGZTdZ68WaYzSPm+2VpqHefBs8UJ9RrytEaN2xHJPGt6Rw1x/S1ZZw1efowwP4TQ
x/zv8kR14T5uwvU9vx7ifjzlRUCtTxed1TZQx2VLfYA89CY+p924U1P4Wk6zggXs
6Xc4TyssBLR2DJ//AGi7NWZlrhHHJx/OZvAFvoJ3qE6iiU9PZ1Do0Ekgt3QaGgee
A0qNLscoFm/ja5c4lprG9KKmjCNR1qN4R/ca/sJ8PKZRDQZBZYc7T1aBIaQ8uae9
CtR8SSHIBUUkz15OzU3AudyeW2Sd3X3zUrlfisCUxcR9kn/K2hGbbbz+lVVAYAn/
BtreIAFdx3/j3A6fBHhWA3q5VCkmW3Or/Qdi+LkwI+kdr1dKos8NAdedVR75efZe
BDzUyeIX4lapcOac1XTcynjRj5bZGCy1ZebH/2QbgysB9sgcd+iES6SyrJL3Dhji
Sv1Yd9Z8oYATHu9cWkPhfEzUvwnL3Bv6ua/838hacZ9jG9GMF/Lptfg6+7OY9xRB
jYHM7nKQhiGq++UJJ1gfmqGcpSQ6NRDfHRRhNxzaC6wPiOPww05grOo//Z7mPT+Z
3WniNge++dTgcGVGZUg2+FBK0tevQyeh5SU1UyBCUXtBXuvD3arqg5n8ExFkt24N
hMPd64xgOLNRTLqyNWAoGxa8CRQo2KBDYZVQSGJBDdV2ZinykGiXeSu+Um8EQQkR
LerL98smX+agwzNGNO3tR5v7oSFuWMBiCyXpdZPtN6Ob8nymXlbJ/90q61tJlaBZ
vUP2VB1J8TkdOV/IOvFgHBMonHSydAX/LYygIt4t5iD4VC5rQ0n5CnNzMbsGlckl
0suiBiO3wApRE7DdjwTLvxVW8BV1FpAeizu6oHy5ve0z8kj61/pcO/MXGzyqpqXu
Xo3ZYWrYRE896G5to3RUOBWlstYqlpzgnzut8H51AFriEOfqI3egGW7OdzWkCgXs
1Asxl6jjex4jmyKZmkrlDsA6iUe7MvOre+j+q5QjrNdLQ/CpDLY8b6NLZOG0mgna
+lGXElBqJyhIszCXWfIhB59dxn30Xuj/yik2afMTmyxAG+0uwreIPU/MQXisofL0
LjoWSAO6AFgmSA5cDw6eh5Kd248fa6PXqoI8y6iLE20NUFr43D6vKQNQToKswnmV
xaCDqOL9Zc8GWgHu1ZatvC1fIAaoYxZRZZY1Y83+BZ78s3rd5BBqwCjJ/9tYz+LF
XDyKm2p0bX2ri1/MbCiV7EUBbKnoj9vsaLDI0Mv1kDxvL4AqfIw9zVwzFX+RYbGd
6lf+fQBDkNMnHlhMAevNzdoqA5gBgiG5NYBW35NWNtnenPbrHLTaDA0swgeb1uE+
8+CwIAfxpVnusE+4niWBJtVAcaqcRo2FnayKGUyYjRsC9ajX+87C18Rq/GNKaTM9
MJd+huC/KX8S4U2dTbPKIlY8QtrlIAXqkzqRJmpiSUG9UTOLquUvB14SQvp7LVIH
Y5hK90R5i9Tss3ZRNXpF5TfSI5WHGO8yHQD+FoIBwbee4cLRFvxaIDOHA+P2UtwL
UFmSym03hOIq1ejWgrfEaoGn+9Z/DM9P9O/baV+a7xRHxbNamZxeg/eVWk3gYnHb
d7Y31/FHMs0S4ycJAJDdcCbF+TeIcYFLG+JFTAnOh2pst3Pte/hAXGut1G05y8XX
0q2jjnDw0rOJC/gLo6TlcVbrhjI6ZmXmwLn67/T/R4o2lU2ktOqViLg4HCR2f5BU
Be3o1xlEVvYP3ksgPjHViHPhogIE5MXQ1+piHj5TNf1obAJjnDtsd0rEW9e/HI9w
nKCphED1/zVnpkuIFO48BbbyAofIMUqjx8VF4RA0MX02uh/zfVobCZbNLI/bC/l5
B+/zZYjLIcRBWu9B4R63jZjXhdz4TFI0JpEJrW/zSu6W88z4qoH+RvtYxrjkVoar
plnzqb+7u95uGcclaVtaQYBbw7j2AoH5rMTJHOo/+JkLaCfXs0Hfbs2EKcvV7jNw
Z8Q618sLetlKVGIj2VFJDyiR6MuhplritsbaMIkIQfSMbpEnPRKX9HQlqSf7XbeS
WO8ZBSnrabqdM7sJlHNxO1IUw4ljO7cgzTK3X3Azj/SU4hGm7C5zb/a+ZbY3J35c
2Ubl8mvCj2SwGQK0+lHYgpoeHPIIjZRK1Bq/hddnfcTJDRsZn7nwAl+T/mCjVfFz
npkL2csdbKVib6mN7Go34SQrzo492X/0QZt/vLA9tC1A6+HcSE72A19PEBws905S
RJMj9BDFZ8aq6btABYT6u6Qngf/fyN/2zTK3+L+LzpYbz6plAYp8dHQ1QxhGkpxH
GGKJ42XMLZ2EEBw5GlZtGsumIJkpiZ1LU63LPM5O2WQs5E2cWDF92Lce7TMaFvk4
PSBgKI2wRhzhgG1eevpasXCTfXE5EFHgIo2S+WUpo6vHgxN6T2jxDrXD043iZtl7
wgFepcpQ4of1UX21fff7dfizUmLNVKebnBcWDQIE2HciHC11KkZFnQlWReZxpXSw
7ouZ7WzaEol+JUFhu6Wpx/T2M8WSFWQsJd27xRjSU5M2A7vU3+uIsS6F0kmOqnLc
aJKF3o/QX4EIyHBCvIadovigRxBOCeQKV+ChePWSC4TtKYr2YCmWVZ5muhcFlNpt
L5YQTFOtedbP0AIAlPIgBOoR/pJpRClIVHzeULTCW3J4py5Pdqc7cg2eOWuqZpdJ
/KP/ziQvQ0dgnaUfjPXYbyccC2G22km7wLjCFOOOY61dO6k8gqxH6A9TTViKcNNP
/7BFmbvd2eYxH7zoRkkzshGW13SfDG3LJoI+kBLRoy+LMzumcto7LI7uei6X2MX6
/beXVehfqDb9zpK4syR5IMqQwX7MZLo1fZoSHZsTCocIlYmtnYq8eohfSvFp1m9U
KLgMjjgf7El+8OlXZJPlhrZNyWVc5xXn6GDx8SBBSVFps2cV+MhJSmnSQttjZF2e
0SkdeQvpAdCDLjF2oVDQOyIv5NAFeZIkK3vq5KqzXawFHwitMmYcjekYFhK0L+iP
p1mgBxvjDT4dG0x4FFWsDPQXSvEehcKpbfiv5V69hwsGAQJxBUPN4jKMkRzoqJ/1
uv44PouecHm8mxgcgacg+T9dBqdqDirCLRCvvC3ikgyheX65PxQ9s1/ZjaSEDNJs
mTK8Cp3zafDUo/9X/xxOGnLTh//oxDZjudh2T1hx8nlpzP6Z23ZZuoExWhsIeRWt
cxTlLS8dZWjdzdzvdx4KT6EDUtb9Ye8QmtPRXARhoDqizTsFH390I0e+cUQ27p/4
EUp/RYJAKDM+T8ha/DUJpAUY/patvz4cusk74kI+B5Ud317E2KJZuQ9/P84rsUHS
4/gCzZLlTHkBGEzkcb4KHhW1yvymcO+pBs4+Mh9v3p5KI9/vzy54VGqShw/nSEiH
ebgfV+NHW1K+kX2LOafyE7t6rQVAC2Opzz6TkDCUNOZIGMwg/A3EmI1/UdFPUUoL
ZMMeknKBv2GJ0We2RgfysB61grymta3r2s83t3ZTtkxDXlQY7yaAroV8UD2DU1G6
i78mT+kkk5EAADd+Md+c0c/OtpVNqg1Ox0lm//c5KMXSW7oadjlzEiWx45T/zEaw
g0lyO3zRymeocJrPUniRwe+SbSWovkq6NN3B+wL5CXsRPKqZKQd+BZLRf5O1lPfD
nnJV8Dd8sSoBUEHuz3kcResndukbuh9/5tV38LigswwhueZSmJ4L4KULGRJ+0xic
WQU3cU3tPHYWmDUVuBGcyIcCo4k2o5yigJVrReDxyMhzvtCAPDjjsCLbrWFU/Caw
NSpDFzJOiA5YQa0j7wUAgNzjx8/nV3TME+86mjKtfquW9SONlzJyaUfT3m+1BvNN
xPGQ8oW0Sxo8NVwhFHps+Xvr86LTTC5GchmkEUJxi2wZzsKL7YyVWilY9pLzXHj1
5uOrt9CxyYJXmh5GReXp6XrlBcr+Ihv5gd0Kz7xof5IDQyOM3e3gcvrDdSa4Wyyg
f9rdDqCUOjRRZnzx5FYnJLBvFes/3hFW+aF6DTpJLOgVzeGkZGPieqHHZkEWYS7b
jKoEf++/uEx41C7VVnwj0DgZO54KKqz3+vdWOFBZUYZ9lj0KrWZp5mEqOleeBs9w
TXhysfvNQi9/3QJVBzWRgNoum41i8wEh3R0hMAMRft5TktgtuSOwCzLa3bKRp+ci
T+Kq8523F2U9ZBxtcMwvTn68hXLcmh3zDHI/+ydrOjMTBw6w88DbOAV3pzJtFq9a
0gYdq3CHTjLjH22MFqe35DSBYdGgl9aNUnPjkAxMv1pkKmkOGIBexAhPDouZZW5B
bWlBXo11I+1moR91H34FFJP2pdDmopHIS4il4KBm+mAoAFH+H9jM2bWTAhqOX5M5
QckPjhfkZaDXOa0wazW9+GCcfbsOGJHM9E+pmevOFADxEnZEubV8ygdYnmQFtFDM
r5eIrLdjDQX+kgvzuG5ofzvfXJWeLb5cHJkP6orsg3BpYPz03kArjYg3u6x7nKWm
TnMY+t4EelS6F2k/U3fBHMC2iXJI5PqiGOQGwOPi+dYF6JKOCwwgpXFXXjySZxGt
N4E0YnEv+di9YqB4gEwlWV/I3Yv3o6PywHEA80v3CbcOnNLgHWERmw+/7/yeK1NI
Yx19WWP6hsswoASRT/S749GJkalSnXV8zfov9ro9yqD9IYCg/PRngBznPl0dPNi2
W1g+Vw7AuR0zIBqlPPk1byyXGd5lRQy+7LG0pDiJuSQPCpkvTpfcK3PtTtww/1Rd
HTdyvTvjIzdn/zJi8Cco8xqBF9V0hjVAAYLUBeFi60SUkhHfefZhZ363S1auIy5p
bo26ia3xTP/h4Armq1jDe64MT0pMwswkHemz7N2m5kz6ylaNgn8+oSosv9TGIVLS
x/fSQMnKNeQkA/xxh4GxKluNcyxq+Bg/wHFu72wXEUBR1oxOpAGOCuMVaqFg0jxe
hF3qtwDij2AhoVI+ScgkDiGkGQQ684cD/Yx/IIdBRDDh0e6vsKUd2sw3zjmPCNM1
69WGUcDAQUoMwMl34SVQgroCMd4iGY3k04KYHWayPKcA2sMJUUoTezpkZHBuFLj+
RcYzPx7DfEZd3XYy/WKqir7jYCvxWTS0aAHZlZgZ6eIb14S2XtzJPgx5pQ4T/f7q
pFV0rZymZdQypDxBjqnUroawmlhnRbmJq7670TE4MpTPfolxGDFv8ibk7Adj64aR
JY33YUb+bu50o/yh69DyVbXBh/BCEo9beqYlpswzHzd/zafQM57E1K/D2XsblMdN
mFMQUv1iShBQtt9CHzIGDPGKdprqTO/6VFCGuGffvSobJxdKjXfp9qAxOHvdW2p8
mIbd+xDAZttLfxu0aUxfWvOho7EeU0XrvV3hblMXGFiJrlNpsuSQtF53oVV2wAsh
Rd5hyFywkikznXnqw+zjvBUUNtG6iYVpFnI7w5g2EVlhFPC0FkUAYw4Zn9xmHHuu
bnCj+pnwRyYmaIpwNiCaMrmcEsI3Hl2f5oiaO7AnZnCcSF4iwy8MdJilghLU2nCQ
i0bIPhg0saWK/E8ZVc2N4E8xD8oTQLAP1Odj86pSFRVPh6zZxajjJGP1eG1anZzh
/o3kDo7k3Zkd1OHWQ2PNlvzPGrinV05TImje4bC7DbajO/IFwLpfBUvw1A+vGY0u
jye5qWPmNhyWwSyzFbNi9LWq3LwjEzJUGuu1jEO88hmy06PmWFhwu56gP7v2tdjK
85wd4/hl2+hT9WnjAPW4ehST3DLJlQrMhBvU15PEeuSOAtO/+1NsqJx3DLa1DB9w
0SKQU54eKb84gqtxvtwaKqQt7U+s4HJdzrb0xGtzzsSjVKnysRSbNJgl7+nTWZ3P
OsEhI1i4DHOXMyK9KtL9PWtFJQlO8RIK+LrKwxeSf3g1xFi4IW6JZZ8QbOPKC8Fi
MQQ6jijlAMNRYQburuVK/xj2Q6ZbEZmghZQpViIIwHakTcmIj1Dgyu3lJ/3nspcQ
PXGQ3MVRxlvEBNwUdvjWCXjcKLkPJqTJJhFEZy1sK1Iiq+WPce1WJ/fpPYwvTQtM
NCpPy/EpuVIrrKZLoTVj6H8duK3X8o25pqER+krDcvNmQO9S7Z802pkeTpeUZ9YE
Qdn9TM9WlRJCKODrWZJV3Qcsv4QFIQXkVYWa19pCnp+LJHnw/qqBzbAtM86lPuXj
kN7hC6ghjzwbP+e82qDbo2yG1DOymHXIM9zhSKely/vunf88U15SJU8oPqsSuy/U
XG9zFXJAFU2EairPutvOS5ZkdvEZw9CDpYHcbqP69IiPIeGFPP8f+ewLZQoE6SYy
+i64BODCHMJQb45jEo3PchxaUor5JPnKmjXyFI5DOuMdYWqntct07i0qthr91Ana
FQTUkxkZE8XVNlanSdh92Nd2eTfb80/jyHa93VCAUoZYLxVV5frkolEiTt/BLq5A
lhl57gV0ZmZRt0KrpWliZWtTCti2y9AC0zXsM6XFjS6uMTmdjlQ8V96CmNWXHNW5
SyGXLk0L0yJKWCQfI0lulquZey6c1WGyDMqXcx2CUbCDz5YelfUq+9Wh12LWQlUP
+NlWLjb4agCAlA7PZUocXtws5QkDvzAQD3JxLnjBKM3qut2NC/xBDoknCbQmBkDh
IqDWis64wDRteFdkGjsp7O911mLjXlW+OYXNt8aJMtDXUkw/WCK9t4CWsWZ+nX6S
BI3JyzyU0FaDBlBxV9Ju+OMC6QWStvUtiHFMlk++wg6ox3zkWMoUP0JkL7KHjJhu
0fvdUyPxWKrFGsREBxl3ibQLzz86/ObQk/GDap7Bn49T0SHZozli3WByKEiBFiwz
yD0frOuCnFKqUHAiWGIlGw9PkbwWaTU3G0Pu3CJ99SsYQaDGnvShUNrIT1DTV9sN
DQq5GJ/A2MZzksg3JEPM4xSpw2lj5QrNmUTcUcA/hBxz2Ydf3Uw9cJsMgMk+ZSBq
36uP6186UdDAC9WW+/t6zItcmI1k04Q7r/AOy3ZJ+16Nupp7KLRKcWPbqTa4WFJF
8DXOeOytrF6zgyN2tz7AIIq8kNr97ucuXIQu5rayrWZKrJbhvooY6mj2DW0YJB1Z
wlz5iQ52PuSHsSRsrwe3CjzL31iJLztSP63mpauu9bLpof4lDEd403HhoJy/4/tM
QqONllqiejgP9ffPGE5tb6yDl0n1MHXv90H1HqQUM1QOfTk7zuKLPOmJOhZqm+xi
ogJwK01YGjhfykevFUpjaWSKJ/HdesYSAOV2ceJyFB8SPWAzHfK4VMA7nHkGbsdm
nOvw8KvB6E+OXARAPO/O8ZI2gpo+ev/XEh2GxI+5g3s48Ub2EVUWAQOUgSY3fhQO
9tzbzh094km0giN+HZ4gx4fkSb0XesYlOzBkRXSoxAodo3SqpcLAUBOgVrzh3aT4
VoUbkdVDgr6wb3hdWUCwR2ifeV1+IAl9i4BKCdQTu9OpeyI+8xnxIV7aPlf/gm3F
I8UVQhhnfYY35bq0hz/jZFkC/Otxqgf8y2oyCpx/dl/oNiORra5mSw6YpIyqhqin
SYedZnR7fmUtjLBbOnoMFaJ4voynYXxUEjXqHeUHE0bz45dn0f4/62XMeh4XML3V
EG59R0S8HMmyTtTD3Znd4qIniV9lNs2vedJuj7/WjgpVpRAEP1rhP86H7SDXPqbd
vgx/kWcud40rItnPVZenQaQUXabG5Sf0+PwwJjdreBlcQCae6rBJmOQ/KIW7/5zV
gLuMMamec7eix/7tqeeJ8i9Skztacllei+Nt3WcDg8PYa1jDovFYKh6oHCEvXzRC
qIlB1M8ppfUbHMVcqocTYxsikypV4KU5bdtxbEvPr60T2LlHuEz/U0/bUg7g5vUn
m2BC6bBRiJnwnabevHoicHMmD728s+p3tWFfZ+sybSAepz5jMYfhkXTPG4SdZT4b
gRzqhJj8glcviWyr5Ls+iAtL2B4WabI1d9TACHoZMbS1DwRSxezEsG2UVeYMafD2
Eo+W6Fb7Jr4BWKVQVkn4+OBub4TtNnHWvvSZnDVnMC5CVGH4bh0/v4mJ8H0Pkz+p
J2VXB9iko3t/fnquuCk2VJBEKDo5XGsb0q9LUW/WM0k5+tMrBbANYLqtPuklksUq
1uFHHrX1n2q1oKgJ+luaV3lHW39KTk46UH0vpo6eH6occaw7/ZVSN9uHYD6h01BN
ktUCohKiS5c6v4yJzer2VTNpqKaErr5sQgqIq43j5P2Enmkak0ETdB3pz9RrEQxX
Rj0TECkAvK9KbzhoS4fifdWZrNdDtHy8B4/aLVfdlmiM2VqwA2SC5ifPydUlOcaC
fmPIeAjQj+rZNuyiiraVMSkbcpju5F+WhAZkofK+WZS3ARxJx0aryeW9x6govjOc
TrlPyrUmH0x8H1NSI/PkjYii1o7q/zDdgvDsyIzMK48ZF4FbjKVyeuq9XXnqicN/
jdkCnOd5VCKEvJM66r9gTcwUZnKzsz0cPAhZV6LesTw/2r65v85lPDzwLYu/69sk
abdX3aCt//7NEOPK4S49Qp4ggUUHg6ZFlBiJm0oMTHMUNfkzc0kn5xQe4vMVg2n/
QI2JrA9H0IZnt3TKd+HqBbgddYKPH6iDmvvBgTNBSpeXLRWTH95PCCuHJtNmGwIe
fvWRvSUE1BxtoQQnXFXU6io1Ki15d7iHwR2/L5618v1ttMTPBFpn16wOCH1K1wvN
wErXNIfx8VedJkSVduCfmyfaUF+PN1S+t8zW38IRYPiPLBB6VIqXgMLyPLq7mTYT
yclJMPZr7ihOuNPHoZEWPHbKMRA+7YoGtUQiqhjOYvgqq9RTp8GttAHe3AGsR53P
zWC2kPEmjtn4Iy2kNgxPr1PNcqJaa7rZh1e7tJUlmMJyyKOhHlROWNpDgfCccl/A
P/m5/sEf4F8aJ2TQsaCRL2uMmySTiCeP78qdGhJTlTSc2GlmGL5JEF15OunSoZPR
dFQ8CEw3KgjDOrOUgYUmoCdpS/sB7aKCjy8TbWXmzHRjM5XdgDJNpbdum9whlhqf
SVtMMuej1MrU4JVoiABWjD7xUUpA3ZKqB+lNtdxPO/cLoddAhsTM/LGdX4slHg68
bpziZYXEx/sBp+g5Io4h9lbSp8Z86h6JvbMFn1TirJDskQSBxYsEvyHdtPi7pK58
zBXJzPp/CEP88xrphjN2b//kItqmv1NnFVC78r0Io4ZK8tQ9kim1gtehahl59QN+
rqY9+tqVASnHXGkJgV5zxPEK4Ef/PkMPbXl4+b+pk71D+aD2EbuPQbBxq6IAxHmL
IvXlhtd0DtyduK3S3kus9c0nqgv6+id8PtpXa2UQP9bbSDzrBBDn+Xi2zD7Lb677
HKUY8jeWMv0879GR2pRKXX2AIHfkDjnVVf2/tZ2ZNxlnc6Db5iOShsNwgLILx2Cl
pDSgzdxJQnH+xSbJ9en29OQvZfPd5ge69bH7v4gtUIaPFyh4GPyKmZbWnuXnZWeF
MEio0VZjJsFKDeH+U3pk9APM8MEvJiqFpleNiIqI9VxFeHjixZo2df0a3qQ+jjxp
/nv4iPOpeAr1UlaTeT/PbtEjP+6kVvEVvn90HVW/BAMItxmD/lFaoHF0WSjKF3ME
Ws66tBNe3cQwi04BcGLoZKZXJTr7CN2zy47T4m5wtrc4ufe87KNZNqge1PtkY+Zv
AS8qENfwsDY/yY1jbsEZIT8KbVhcjmZPPAYNwiB6pr6Pz3pGjDbP/bSteZyyBLot
tKixpsvFNykKPUieGm3Q6dz8a7WDU0FTkvi5idUsQnaNI08iMwc3JlYpSgfbUT9G
vqUp9xbrrQOwT8Adeu0jJL1IoZdThZvbcz4u/96Oa2y6H+hnMhIS/fqZyFK1ZJh8
iuWkpN4Hh8d8u5yrwEjqkdAYDqT+6g1Va0wwkH1mZuqO4XDLTJXxFJXbhqRiG5zY
9M19moh6RiCXPqrDEFL1lpUkpG9kF9casiyAFDssxlG7CrTVF+xPwrO1zwPjeFH8
XH8/117pbh+b+nEG06AMdydVWD4ahVYBlTaA31r9oFfpi2OXqjjyIPOZsPvjb7VR
e/RUobSsGTbxA9RwnXTPZUv01FWXWWRcRGotTt1vIM72HzpfzMZWgKCdRKMdmlR4
cPfjhe/pCwA4bp2vXCzfM8BFWrV8wEqz+7nFiycIEVlHwkOW0XHrmWzYEUyDv3ct
ggAfSxIqdN0YeHhWULCx7SFIOyFWU5OB3D2kkurxizFdwKUpJflyrzLOjPBjULbN
kiyftv/fiiPXFDNhroQeHe6WbIAz0f8tcsZNLOW1gpx8BGOzBpvXXIIR+9sihxDz
e9ml2Lkvj9iFB+dxbt5se71hySc23mkVaUb8vBI66Zcmkx1ASCC+5GySnPsQaoY6
q0xqqMjdSqvFbzhYJe57uIeebsd1wWzSsbMS8vVpjmVnMBT/3bCEQ7cxXMjwr3q0
45NXp5HVuFQ9UIqliI3Gh3UwSNwZvDrp19strkDzeeT2KYbJpIq2cPxvZcj+g00R
bq7Fxt+pE0ePoYAitDIjhwpzVrgfzG8c8HaAWAoNQ5rNGUxabnS/IhZ51hXrh7eH
ehhyg2H2Ne/8iFPu4Wpx1bJqWDvaKJieXAd8SFXMd783rOx4n05ZOqV/24kOxudB
85WTdgtLPlr3l2H9QMORnVhzHH1tKxSRxMDXblDqo25/ATQoXDDLkYea7pGnm6J9
ZdFVYQ12KQug7wGx8Z/4oZgDZSlwQMyPQZ2JdwzpDptZjmDbpVUlVHQlTIyvEHP1
INpq+Sj9oRzkfxJtLIWgj59R6yP6VQGlJyz387tW6PIwAYYWncVFrdI2c37uLUzn
EvtlRzTvpgVzgrq15JeCXzNwIM0/ArUHvsVZXRmJcJmykiNU5ajEhS5zHSHmkyvu
sCTBwDOIDuDHMJ5FdcRFcltMeS0StpAswH8F9kHEDV76l2aYv4scjM38ZI+tAywl
Fg/G8JDl/roY68dQN39HgRabajjwm2uOhnpNafPsU5O9w5evn+fCr4lfCzOQprt4
IPP3IQvohbNRmbBZrH4lDEtvnSRiwY455JbBD+tBILd0ZrjyHi8J0ZAJpiGLpFhS
+diWwt3ipfjn0+smaLZkd7lrpOobAzd7zwTVzWhqJp+VmdCT1T9sQEYLIlUbeGyC
snZjj5KX7BaiHFTTibr0h/7+5M2ux+Z6UUZYOR100NYbbyzZQs2qElzn2nZBqlOw
rMSR7qB5P5jgnsm5iB1LR6BbvPrwVhP98Hivdm20sqh/kw3YNpMYs09smTHDPzrD
3X71aSM/ocwJNQYx/0HjgyWTJAhre1KOt4AoJ66CRuW6grPR6tL/Ice1Kj7TvtjM
gnciGzyQS69JpE6sl4mrSr89zFjZ+DaKSFynG1eWlSYe3KGL5WBCm5Mf74ZCMwvS
t8B47Z6EbhSi92DYVQayumV7Jcpuuf57EwVgUWGW3EYxLW4PdkM6r3jXAOhAa/dP
/R7tZzfQxM9pTX4ctX6Dnp7hsdbXjg05/YyNLDgtzeL2oAWBJxTpoDM68zpxWatV
gOHiSQuk4lXqhqoFYEEhoPK7jAE5Z+jM9Z6GqgSn3QtqWWBBHAJb14B3vUX/B3SK
yNzfSKE33f59Q/2DuT2fFqe0m8Gq4fE00lW8E9YO6nxwy4rlT7YXFh3XUvBi5YWO
PIVeV5fs3yepgjwlg8i+lNuY6ZMqqBZo+34rkX/gqy8osZX7m+C+H5Te1gsmVSKh
7mj2ILteIRq10CW/JxbZuWIZaDDsHqoM3gJuWWMcomN34nxpczbOXtBZc2kv8hqI
zBeu1HZExtqIHletsK6lsCAxnt5jY5TxGOiUCf87kg2OGrDXWpmC/S0YvIBSGLwy
ioGrLHuD42M6du1Rn3TJnY2WxmXK01shqIFM9wl2GGdAAospl8TbOrPHRlmXgrKr
/ucAAxa3hfgk0yxkOUgjAGxoHxdkXC4n1ChjASTVSALz/tspBMH1cuwdG1hh9+f5
HrdGCC+HCriTLVv5Kn9goDQl//X1dpmCOk3pWlp/jsuhdDdTn//wMFxcgcaYRbHU
CNGBCD9vIq8c9I6tiA2UbGij9Gi9YVLa3bLG1/3d7r998w9hlQwW71fC7e3OwrXU
6sNHFxYl526MxNgtPaTRbDcySUS6RL2DJZNn0aQ4+DO6aQ9nU/GCB/U/0X+8GQ9l
e7KN4zINR/LQBlERO8i6QZSYHdqDCJZ+0ixKEbPzY2cbUo7x7Ky9tXs5w+jy+Osn
x/20dkv8iVcCpSTcQR+xmyQlxLONVv0HyUvOERmdiJ49v2WX58R50f3b1xhL+xe8
DFVSBXG63s/crDOThoc9rjxaYJZP/xA4feFX5iZkG6EN+RgHG3+vmCjIHjaxCcRc
wetJricbvmkOMr1D/K65yhsndGspiFQJBx3zIX8PfUh28NQ56HSCD6fGTj/iuF1t
TNpOXg1gxENhHbXvBkY9ehs40+rFAB9ISz7mqabjEz80KHR5sofYNPcCtlsp/EGL
yhw+LgpV2Wr8SQn5hwUR4VeFVzoAo6FyZP6ewO6yiw64ojpDMqPB/fZdc+I+VkIK
HDmcGkZB1UUrRujhm/54RseO76m1TCfmsFwkj3AklczvtLnshqqFIhKSx8j1XTLp
6g/OxZow3o9lzk4zNFa35HWds2Ct5/BxfrI50nn3IBpt2r5MBFLsIN0vz/wrI07t
HeZXIQr6t0iaUjVtATi+zU3lIGB464cAsiJxXXsIZUc3Ru4OAlYOFdaVUKqOCWRY
TU5WIpfUIttg+WkSHwSsDeuxdMqJvfFjkF2ZVCGj0DRh5QAkGSzE7M+wBVoKhaJy
5kOJ25JvFhakp6F5ACwn2zstZjEH8sN6L51J38BC9DKVrd0mAEH3QfL6ylL5/Vlu
E21iz3V/EpF5A45B392nGV9iZ1sKBtlv3niC0jSAo2y+p/wdom/ura5RA7VE3IvV
YuHIRZoKNdyWxljlKShKTqv9kmaU4L7DZutjXEH2UMq3GvAasoks5dydT8a+MnLB
PraVJc/BeLyDrDhF1wZqPQUNO3D17Iqo1tUvQWNrz0ONogwsXV5rrjUwrxW6fh5h
IyFnsmxA39S6Y+K3tJkrfJNOR28dt/tXRLtmZ2C3KO0K10g2Syq8ajg9EPSKvrZF
g71yUrY4wCLLouseCL0Su7O8DHhYjpy8P2E3dAXXjuzhaGXi8AQfUCkfR1nz7rlc
Tf2tsJMx5CjnxnGo6Tn0wqBZR6ES/2GgAImPhIKVdZB3TGDCT7ChVF/evC1NiQgL
pHnS8euBQSXMwH2Yb/wuIw/bjm9kB5sMUP76+YNdGDqc7RI69jSs4MfBmtPQZfE8
yaBEkJ0b0OCDRm4dB/H2IoOU8+I3nqULHS6figgHYJrX2yj6e3ztn20lUxzTbdQq
K/PY4EL2Mh6Cy9KDiyogwBgCRNDXs9B+aEU8WiS46qs6MHRwCksnYzaCj38Omw1P
W9AqMRPQRwKler9D6OQP5wDJL8CJS319Y3CcVj1f/hIjmDfET39MvoblteKigGIX
ZvC+cF1Sie67QyI6f/ZLrpfYrUpgnPhfc4zEMMR20rH+7kDkg34WzoTe9wQzuvkd
LbO1vHd/ewiiqUojS9mV1HameCGCZGvdF2pBOuHQmIksj+AUOrQcHNGkLKXml4RE
5LbAgZHRsjanJ1Ben+CTX9gNtNyC9ObzkqC8+CN7nfpTJOmdomuJ3KV2WGXgOKHK
a75hvIiHJQ7+dLD2cHysdT4r0jEkiL4dlKwI+3GWv/4Pw4rQx65o+IQ6BEUubWwf
bipXtGGUO8ERtX5SWoXDIyVurw7pTdicC7DYdeSxpHLM6akueJ9KnjF4lDsAJhsT
21cRzlwebYsIWsq/KjSlHuCtmWUrNtfDONMxh0I0ZVNMOJAcLr9O1rMScNcMUTdB
xLxnZji49NcuQOu9Rbdviy8zX1gFrCZm7OunfTiL336vNrM1HOypioeAX1NynQUO
JEIvUKrjfOxyLrk0ul0YnfzIPQJ9ySIxMACfKSbErtrgtKeocLlnAlCDmJWOdbfN
ckChKEvKL/DqU9w7eAC7odKUZ8DVZhkT2RkTw00cJvqetF9TngDw5RjP4ci0MVrq
1oxPAO9CTSVunZ+vSM7woEmnU9C/7dF/ZzqPcapikpV8+cGrPif+6AN8ifpg6Mek
3iKwayKiwaDIFjY8gVw39icn3iERQ16OwSuaQs0lW7rXyv8R7CIbhMUo0xrvqyZ5
JUmrwvD/oQi/fFYxaCcLRrBloKvTn0PzGhSG6Cf5NQHsBYB8xniL8fjidXMy+Neh
ywXPfBOjQEh+MW6VnbBATn8JoCQAcci6WVpjydaeB5NOq4gC3iR3TL36hwA1kjGH
Fo8CDQxCX6iztsrYXxRLnnnetuEqM6yLEs2jfIPG/EOH9UGKQ2IdSjwAqUayooRz
rmV+CyQKSS7uZoUBO4eY6ZhP2isARUTt7+8fCDJr+LpdKBTbVItPw6qptk9zsj+N
f7jVrQPFPmZUGRqxT8CSGDRUFN5IDo4gP57G68HoFFZuk0DHaWNfVcJBarXd1gUC
rxfSkHx/WI0cDek4Yq+XFX+yPLfdKPrljo1gH7D8YOedwMW3Gd21dxF/1/CNdRxD
jdJx3pFjXbfWcs7oWfP9pVyIkNaiAf4c1Ipf3Y4S2hrWfz/70up68dY2vLwtT5v8
uZaVnP4XW+FkDLtpTFxc5AEvQK5obf5yQYdy+nyCLqa5UnC/TbKot/IXJw41wTFj
oBbaoacP99tNSRaASio9+Hy1ZkQCS4ZU1NE5MH+M4zupwpN/p7Zxt+PS6wm7gOFq
g85RR2jL11ZvQQ9DEi84lkpzR2zOdsdji/7Ogw7lsdA9M2goC4mZWHM1rgzHg5E7
UuOeM4zEq8Ipk2iMdcKcVK0g04n/wXkrNPbhBU4VepK1L0DSw3LJZCS/lXIRsksv
sevO3f8WzBYq1VrlzJnFOZizaz93uXUzsxhsiYDVf017J1YLIG8CGd/hmTDo4+ek
qO0O8hREb1HdtrY3KWC9VBvOCOXsaRwOXiWWZjUrT7o1u1DeA1rLnlSh6VbkkIhO
jZaNIiFHZhZF+LIQaxyMx5Fu5HKextk3991+fuCw5AqEGVP8+A9dzgHmSDipxlnX
vNriiG7jFXHgxW+ZYmPrUH3RHE1+7JvKjJoQbpxyRLFK71ccyO+NzHD4fsbwq8J5
/zdOu+GWzXir4fvSvbiWgNBQyjYPkkPG7/8B0v5gG96ndOf5ybsh+uY5OrlYHBvl
3IE7i7xDaGsOTH1q+yRSftWYGzGFKCyKM+OViz5ApqgCMVfYqYjelgy7gFjyMt9o
J6IgZuTGqftzSkDaibhrpAaFcz8jEN7Xsy0GvDIFfatEydZApkmWf0D+pFslffIB
15wRPqh6c432CtVnWIyCNNbYnI2Tvx6ybGNEnJbfQdr8w8aKnaL3rhRM8bo87LDp
/HeJ+GngjbZbbYXfTUbRoxzbLcrucKeioN4RpSJe86AfuF97rUskeMAVlxCa8AAv
2dmFpigDhfkLb4vjuYeIydCov1t8PdCzF9gC/NTVexHP4cL9cu6IYUDFtdLf/IzJ
GgiYPcjWWtJNkcDEfoRh1rLXMnDgXymO6XIqRbkU2EGGgF49u85SnSrpYtYYPqkI
4T73rh5GyggXaYeaG3VW4LyQwawqldATgFJms2ou3QjTcMD+cKoN+4RCkFBt+lVC
dRVN8F9qNan9198hvBVnInv8XjRh61pElJlxXbCiyf5VIJ29jzn0M0U/bKBQqvY1
gmAoP30SV6bQeXFnzF+DCzZlWE6JlWyzX2KgQG3X4/OKlnAbq6pIjaKdn14Kgn3n
n+V652ynxMW5nHS+MOxw1+VxenLDF63rJ5L8gofz7i+ihC9hJxJ3MdvXViXYXzmQ
upH0ScJqgJRWziwWgjiKabTRTHVEz0B4Y7Lap7DBgfB9Eq6HC23JOtTnxerAalXy
awAth1QxpxsLeAeNwRuIWf1gYk+SY7lq7WKVcdZ7/yuZ0V86DEUvZ90nvsts7mJz
mg+jgUz0dm6sGbSVB/3FQQjwaYEQp7tb1jivx1/AXhwxoHFP+oE6vHYu7hxX05el
eX0NCdPM+Z1oLH4ONkOjzVta/0PZEwtRlT/5DGPIjRrqxRyJWoAk1zlI9V/S41gK
WXlfEc8WwcjDVDvRQErIUcLuU4yBumis9/rDCCEzF7b3h3QkwDjf/FG/YWZUFmON
azJ6qgIABBuiRjS2v86ABxRn4Bc452uCpvIEwh+i3XVRRcHbeP902QV88W8h2VIp
M5BrXU4kCaHPOQ8vqcMrLM/DyuwXNFyiEwfkx+ZCBMq0Z2hukf7Ha9e/WtzfNlyp
mX/o/EEeeacpos2F42Jvmsn34fr0cB59ANeHUF3nBNicGNl6jOA3vbkpWOrdg8iR
f0ekHBZU0v/r2VfuKOTPYA1zjluUoXptcYTTymYx9ktN+liazZ8icr6LgweYm+DR
1ZD9gwPxmjOo/khSWwn2rb9MjQacHePY0jtkUKjNxLcmaZ1+U5ocLQKoaQZm+uHQ
di+pCqDGScuyG8cwuPOMVSGksDD5zUFIOOUw/dASTB0uYc8CSN6+ZqdmzuRkc02/
HYDz4kLHjm+SsEk+SiHonEd1Nxjl3aFkqQwvvUqK+QKIeUQXIVAjnbb5go++lDQQ
VeY0l2riI2Aqs5jMdtlFdbexnifmIMyGVx0NI6dl8hwTzbZCJJwUdmRHUvibVIxb
ArB140LoslopMHDCq8S1Rh4k57gQKocErCe3w8JIIKPfH45LQoPyuYsmkzOlKZ7f
4uChx5lJik3xyB8iNVJWycKIx2YVSaffp0R4q2v4CwR1+ncY0l0NpZImg3XDhlrV
iYdiOtwjx+DYWWeCNom7/Q/uvjW78VofS4VNlOY5bOLEp2mDSs2+QivBoogxSAAC
mUpWzF5RsS4SMEdOTe31t0y7jWw3kHstAbDW5DOjp1Q0zZd4HkF71MHs6PGG+Z8i
qFX4EMEMg9ty+TJ6NS4qMIBslLfSqv7qSX9JYyk8+tI4WPaH8mi8byK6RNlwdXwE
ZLOF6y7QM/gnrJeP+khGAJvnL+O+vlgy90IskfyLoMKhVU2IfKPz0yLoqaVR7ADw
1e9tMbOb9XLPQVbJbfF/izCHjj8LhguiC/Psfi1gw55trUFUx1z6/8s3juDy7nab
DYxtwx/OpsdvvHNIQeijOwL8O7NGf1rHmus1Wg/KtMEMil3hpMT7Cw/I564LOJ7P
AkUQAKb72ScH/2ofx4gUxu4ZT14RDJ39ITWP4ve/XAQq4oQfFKHFiu7991HBc6YF
2W0uF3fP5NCegNlNKwdAceuBGdiRqYQW9kQi9F2Z+UtCnMrcTnFs9VcJ+YTIkRp4
zhZjSTdEBjrTZyLwtdFDe+w0rNQcPIcnPfzmaHHRFQlPEUqmD9y4pINgubByGPed
O+61yS2DEXN45n0otM+ThWNhqtdwRrw0wB9cBESml3/3panVcZHCnpdLoYKPssZw
sWFRCk0UTrHLSl52hNgrho1Ud5uUtUWIrwyIn6L0ws1W8jcZPPxMW3DOVPr2XFvN
GU98kcVyTg5B2izyV6YvVIigqgcT1SBZ/eK5q7i7EhM95rLBrpwS+aCnt0KE4qzI
arKefDNeeygVHGvtKrcAFWk0UA2K2pRYH9rZAD4pp3caGwQOP3p0XTJsbbC+lWPX
163cnyZbaog1ekqVut0CY3u9Ycy2b5bsXLJ8BglcJdTH3UdKzRPiXWAls7CHHBJM
oMUkxpwta6/M8Niufzvr6UriC1aYWePqOSLpiMloouB8IWW1fyllGUyMZXfIlb27
GHaaeA5lUbnD72TxBPgXYx4tQ5hPZSBenv9u74dRRNH0REPb3fW1iik3IiKcJMjK
YlR2ps1Sxa91F080b1QevdfvThMiEOCL7h2bGyYxG4rEqmxmp/eas4TOZP5hR0kJ
FM1BDn0sA1ijwU3C7azwAQxII7ijJC3QLH+kMJwIZSFm2WAkTESFawQpYJa2kEiP
mBftuK/h8uHsRItdSiajFhrKlFnvSrb/umrp5KrOi0L+eph//AoiAla1MIMM8vQg
QWfUWct+O1UzrizjUGv0jTSmR/wg44+1HGUqd5D3H/HXlsQy18lqpJSqR85CICc+
UeuHkuxBw0kW52LscigtrhDTk/AIVdaA0E7vYeDXF6Jp5P1cJ+PsmPWh5/I1zgl5
XF5+cx3GJV8Z5g0scAiEW0wil4wzVqwRKHbxL7PPy/56uqe3Mbb9mTsyxiXoHEM4
proKouwPi+U4QzezWffRE51b94EizFA/p3QXMu6TeuXI4Hb9ahKgySIvw02Pk/3e
TxNH59lYGOyG32/VHBxePPil7sGPWBMj3itj0B69uNyfXPjuqHpiJQMPdjbmwZIt
P5mtEogopDJdpZqdyBXl/9xJWeyMP8MIhQ2kcm25NLRqJzWd9toWcce2EnU6gipu
ayr2ueN6A1F94jnTlhhMfBul7eN8xViJNNdZDVOfjeFtB9BEmZlc7l0A8Nqf4tBU
sUbRSM2wiY2/q4oqqN+x27E+pPPXP+Afh7MNXRzAwldj8ojAwg6JiW5HA1IUm7Cy
6Qvbot3jvI4fT2VJulA2bE+WXnik9M33d1+S8HO9blgJUHOGBL8whAvVGdTxHxLi
4gqJaBa1enaynNNwfEqdNPUeyfPjir/W3Ffjm7sQsWdQFtLwb62rYNPxnD8/QkZC
WROzDPQET5Xk0bhFhMyggkSU9fKNR75b2KqQ+2gJyS7J0cfe0SSkXU1tBEOxwWwj
WOpgcEqQKn9dPNqGPpPVPyDh0o+M7vMqPwbP/xx0vFJq07fuZddTIkDpA3MFj9te
sLEpfHel2fdElqwTww/ENRFz3bxD5lm2gQ8xdARjeyjYquzZwSvsf+VNDaTRJxqQ
QTPf6lniuuiddJPzyqcurxgiVD6aqyNRtwWL4JB4KgIad5CWNvHR81jgdWe+7Mjo
YE2MBAcwZLbXy45hu5UWzEiUG4cM2GTtQMFdY+37jRKatg3TmFXk3QrJKc1sDNSE
uw0PrZLULo0lXP4J4fohf38CKRJHLjVa8dG2wtdgt+9i8Qefe6VrRCO0dfuqqyyI
stzIH7hWdzcAEfnod+geWYgwYNsCvpnnAC9yVGt4C7vC8n74J1k11fRA3o/M+Vhv
HemTbWafdBA48vv1BDIXA8d3/Vi0XQCY3PPj6FhuZhaRHA4MWC1B3BZvjtu+cGdj
RUVMaoayiGWCJ03iSg8EI9agTEypn0SSm+UZEAEgMkSiTXIZ+O4bbV97ojhtrlku
NS9iQanhXpBGASRhopAWR0uO7PneDghJZvfhDPSOILaSFBYqi9heDuXKb5tB+n8n
ovC+PyOuBvAXpmXxXTr+pJhoCur5f/ic05xOgla5OfaqEgTnP9zolL7vvxPLtGRF
uFI/IgL8U4bd/rq03NaLpFCfnypYs/2haD6kE84JaN83jCXXYyWVYSKYcViV0c9G
g5EXpw5tPHRLY2IjN3ZReX51PHVzpViOHWU+jxmCADC5qe2XxkVux4QRD/ElM2+J
g/AUq7wo/MBPDnHfhD43asrrECXEfQqwuBvtuXixiFCfK6ppoqfPWM6K1efT80Qt
WUltKB9UqzeCJanmcp5RM/jJHLbuuMtmuMc5n3+dPIb9cyhvMgSkgt3rG783lo1x
Nfewp/9rZHC7ct112bdvUuZxgLloF1qSNsztzxBhp1KGhXDVa7xe+sjoP1X2INKD
wyE8MNri/nWIwWptQiyKA5mc0hN19ounxJWoGS0yufKnsa2HyxNWDC1TfBsPhscu
5xtPPNaTPgB6cQH1TLbpAZaM/tjyt+YfydCgh0wrF5FjpO610/zkvsZ7XQShmS3N
k12+8FAWX4kCBLTR3cTLlkw+bNJal/8rkIKZ0Nm09xkjgEwx6dCOC2tLAjU5XqM1
/JyMt87sSFsCR/orLJzMnDzjnhLQwHWv+FHjFQumn/+R9aIsFVbb0b/kUwV31aml
9s6ibzG2/dhDgKrwyoKIPUBtUlhF+YwFpxKEwvz0oxpI5xe2wGuvkWgBMHNO2Q1z
pZHFFAHJcPE3iwhGZCcPWr7+DTRbMD0e7zSuc71VSZFQmy2Gqhls5HUYN1n+/O69
WZa/GsnFOsR5mjqvbA8DOFwJEGciOmpmzwUDcCI/oV+/AgPMvZZXtPrbrTllls+J
7ZovJfwD7YOGqGhlbtaYSALe98lrtFmum5qUSEJHfVkeGX97Je233rZRb+hb7u86
quyDXydYcwmUBs3skgHObmdSPgeti+AW/N79raZn2FFBqVqDt5opsJmcE2IykQ3q
OdQtoLkvibmgVRMW+x88u2SaA6hQT6GsfPfI9bhaubEg2oPGv4okAuiNHrweZi+O
kQbUePnHk+nH8y2TlQ0bP4C0oHMi0B8/k3d5YPLim3+iAFhZsgUlxPSfuwRasdg4
WMzImFGDfgkEfvrlIFAvB5JyTMhtEy0CKrZL86haCZJaT1O/bk6Ko3F4AbtVXsH3
uJo5Z6apsw0DQOCuWZfi12w8zMYmKCPRToCnkimoDm9Bj8fRL4bp6Z4Bnit9vrnn
S83v1Cdn6mSnFfgjxW704Ke/rQnFDGgPovUleoSd7ybMF+J3Wd+sX29LMxx82vIW
mC8XJ9tI/JjuVCRVF5EAWI1S+cHgsecYMP6l7B6A2+RPNnkZQNUtqRXmXwrAGdUB
+U34IFI+nyVcG96m7sE3KGnGtKp7kwU7GZ+BcBE1c0OnrpNL+8IzR1BYcRWRAgLW
EYs8QQ/+YMqwyjHnICP6eoFGSDL7ZOz4x8z2ElKf8bVsHIu22tAP6cT/Wy9ZKjwT
cIVm7iqSAD4Zf2OyD0jvHtpv3Ca4lAP2BvItWMnU2LwvR9izw/rsxf2aCPMVeqa1
c8qwRkoriNFvSpiR0jx+dJSr+xu1zDcjrt4JFrt9wgxniU3HMBpQAZkdvkVYq9vy
aO51ko0WMquXLvV9AuY6KKtA2vzqEe5UZg7nvmI3JeIvZ9Q3cApC/stRfl7XV0kU
OpLjYcggkWAYc3t3KektWpqUG/8A/VJRYGoIPSukgTQ/8b/TowqTXyqpR8ZCsO+N
qQC3L2X9/vmgfl2vtlZIdiaw6tvHBAg0jV1hqcYI2WDlvaGH7lTbM0r0WqC/eajm
Xp1pRNUSj/9w0WQfZjB2XE+c8kq5weRO9DpSRDG6Q/viwNIVqZ83P0E825xJpGYc
1LsdiTj4HObqcoYPspnw87TA8FjCLBvc3XbM3RLQ+KbrIB3N7TV2TtL9szzXmiW5
kzFVETXa256C8jogL7FIQE8w8B1qrjN6eKeSIL7QIJO906YGCVECZEfNdvwp8Pj9
hqtsKg7a/11JUFkMptAZrGpmZXKVYEAFs69cIo3FvA3O59odLnJ5tGDNJ7z5LVeG
puA1TIgzwV47JNK1CjtW6tP2M0T9J/iTiJFrlGxNkj9kQk7EqL6gvrUdaGaO/fC+
e5CIeMQyrId/T+D1Fv55oUdMbYnNTH3ijTWpsBMEnUJu7xmOW0MTfWFZ0Mg69HsU
OJC6j9O+4pLVReOr+CKS2P8UUfaOUUbxkPO8/S3BeVadWL4dpQSD7tkaNp57jitd
OAF62WZcHvITI/RjcOTz+OdOa1PqRCkBJmwFz063BI/C6T4JA6IAyrDersTx+XEp
92TbXViOvZssdx9kqmLe3FMc2wW0L+5n/4oIrG5ZD5bRFC2rvywd0Salb9E44kzy
o/X6nMGnbS8ChgBFIpc34M5zMs2XS6fcAdJfdfyEymsWWvq9olYmPI+NVJ+rZgWM
9D9SVeY3CkCeK2Mkl726mW51T8PfCgYVYF0sgt8LBhSXwFrEbX2uvgKYn/cuNYP2
khwm7/ZHioNl7VXgL9k3s2a1eKEh4QTGgEMRwgJAtNTp/wOO6DReZsDnnjtzPfRb
w8M9d+hV77XF9QLW/JtSonClJwoMwmFwcAQv6lAXtX25W6TOtGA5FJPNZWx/Q3jT
JGPlUio9T7lwCbM+/BnOicmYwhhXybLoUPwvxO3IXO/jiHtcH7Rt0XQQaGospPP/
3PKHvsiv8XWqRv8U6lIJ379tucrZ37ranxLfeFngY4osiX4qE+bKhXKx9X3Q5mP4
EkR4TyBKbxw6o/vNkR/znKLQshLZkRocrDW9I1elKNS34f7KDZ1ymBSxMpQWIv55
SPs5L71U6Lry74ZRoE7wehzfAYIwx+3CaRGcRnVdGxSiX2Kk5Nk4FL38ExKQ6llF
ElHp2ICygbwtUXeNqFbdYDJAlqVR9pW1WFVCHpCn8qkfHZYAKClM/on2pRnYWrkU
v4dHT1nmp9SsUhuTBRAq2Bt3EXUx+JKjph42k4lBm8FYwVCuxIjGZEsSb2cFAVYA
v3V88MWxoeET0lGmjiBj68ypn0Il5bOwqtS+2ZV/vVsOoQwekLkWRrS1wNE0nmX8
z94tlqqYEJOON1UPf9Qnxf9bpoW+wJisqT6aviNHyMRpYns3DCquZPkaILraFK29
gBlD+glcmmsZ4treUgQiY0/nUtfosvXqzl876OEjHobPSCJuDXuN/BhpHHkJ3c9h
CntXmrc9oLVwqF1E9JXNHvIcwYai36060NphDj0SgGMvQgBEY7S105zEA8GolPIu
f16OzP2oYjtyyd9bzY1oouuh1ePVvI3H6hX1UVJj7D5o5LKeRyqSwy1/kx/XPGd9
Kp1WW3HBeHyGtEXGQCOMLFLN7I2VLCJ+6e4Gw+vCwfdlZi4QHrwx2zAfuk4CCYdv
8mnukxiHPiN/t/LWUKilhnzYlDtW5ppIbqW9vNlYRpMQywI6FrHwjOmMM2188Z9U
KGL9/OZ0KtmPvKDvbrn009VqvOVXxydNuNDHq8+MShcVq4N8Yeg8c16baGT/OXJ/
PzlUOHTfdy0mvkV+miXXAyH3exxdpNzu+/yzgxYDOIFpfLbXHYef5M5fgLBm7xAX
sF+jlZnnAf/vcqBYOtU7qSwz3aml4Ns5m7RCYvR56e/B6xDx6lzYKivxFNPjJSY3
+IJvvLCDM/GAoHYhCKD8pOqD/Baq+ChMiFU/19Sc1v8eWP+ZsPtttTGaRux7Kj8D
HumWAitdT8lguXL0/6L8YRgfbgjxI6sSVB7qhiW7BL+PWNV+DHfszHClqeSM514m
r3T2QWKh9D4h9P2ROeIPIjKfuT2RVHMOCtE19ebYJqEJwa3nDsasHuSNqYOQxiH6
xo4j9YNJse8XNR8UyG5HwHFvEVJ06s094ssUo7JYetAgvUKbhyYhyeKZG30Y3Tie
/YHIuIk8XARK352oANWGHkL3aPUx4Br6r9pKfjhgAmTbfmAkg3i9Kb/7EJoNJJ35
l8NHCu52muGcCpav8djJT0RStdp+WTlTMw1scOJs51GVhkz8SFuMtBu5rH2Tz97E
d5djobw2t+zHVP5qu9TsHj0+K7UQ6ykQAAaCkIpk6Z95vO9z3VEFastRUg2cSI59
p9QUQCcFhkqBUoI4mG1+2qI8LeFCeqL777MayuFsCW5IXi1axvJZBOs1YjM2D/Zs
GBAa4tTdKVRA2/UGqZQkqRxoiq5VG6cyA1C1Jdb31HCIc0KPFiTrTKwgdL9gUimk
mvEkEWL1IGtNzaxdYiQ35xlG2tmwZqhU7JOw9UpZHNVu3EhUME+Dhda3RzgeHBFV
yuXfzhG7xwAa9uoR/g77ajLVkV29SXJPToHyqzUWgWn33vtH549E+RPcm/iELSP/
X3++FvykvEfRp2RL0XcG3SdfVq6YOlyGzFeHXtEeML00C9f6TQ/xhPlnl0ywqpw0
xPMhc+p3Yp2sUQ+64VO5xHlxiljswhbFuGk2FBGHi0/xZsn9EYbaADfamTTB0uDj
UdLQPnaELlzkNyDhLwXIupBFOAf2BJt+DZFQdvHnC0YpIA9rtG4pk9N0QH9Wy/1h
/Nqy6S4rHUL8SzvgmoaC3wngh6A/11JJCgwo6fCNCd474XLuz6H0ebvkO8TjYYSu
8lIXSfCXE/Y3EiTcOjZrSKH6UrvTQRoYwFG82CgDCAEHcw4ZCcmWrYL+EBuvIFMK
YczLOioF3UyvotrdGtA/+UGMz8m2QWCxRqnJnQBsr4M45Aln4TOg7bdiAb9dAHbR
o0J83kByAWRY2mVW3eE8qUVy4IQd3C18EYQOwAWO63JyBcAesr5XjLf7wiS0BqK4
zV6bv+ffvOCVPVewERVxk/cOCH69L8odmtTxPvPFjSE//xFt3q9y77fUnMkWfTX2
kKfv9qUrccKghrzcq2or6n5+4vpZKODH+rtSZroPY6yeV59QMmPGiHZ6L0BfmKfT
6bpTspMP+qZlQuVjYI93+CqCKROnlnDrOseaeAVdD0GIMI4VYDN/NqYwShBv0rTF
TF8NUh0V3kslj6uNHcYVmIFWCjuMTRO7r6Cuinr1q6j/yrD08V9ghF+pevlU0AFC
CDO4v7I0hVqEDirKjmfdTIRspyEwd/17XA09uG7MvyDR/o+DPtHoo6h5pdgGt3Ua
`protect END_PROTECTED
