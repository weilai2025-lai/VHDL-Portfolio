`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2ZtnUJDIU24b5sgVNbG4lSiFmhCbtVIvOxbzgjBWtjfN/ikPDNiC8y5PCt/UA/V
+JRY6XzBZ6IQMO5AChyU5jbjQljPyPHwxUMBkHlvFse9V5LX6IkMVjhakKi+FaOI
g7cRVfc7yCGLxn7GRTPI73dWZ2jvjRZvdrvJDWitqUeDttJewMIxnEzpShCVAZTK
uFlMpVx6eZhxfTa+KjNHcgOzYZV5fujeXc1Wt4lW/+XqsBR89t67P41mWNxKRIOx
wvo2dmpJbsrOF4t8FuTEwt8VnugGhinXHxC6m32JI8S/d2JnIcgZA9tE9Ehij6FL
z2uC58AhMv61QwDN8O75sUsrsLTCN6By/b998K1ssgoNYN2oeFdfFYbehji1Nt2L
4afFSo6ISI07IjE/iUhPhw5+i5bLbRA4gpolug1fTKqt1hNlY9p4feqv4CIJ38cv
Fd7dMr30q3uVmO0SEqren0fbyNPfkAOBuTvWVR1GIUl9sgJCAqCz42tFVVeFFSVc
TvSpxxqqsED63l2LCjtIliKZijma6uYgL0fDITrw/o61tGu3Wzl7oaA1kE1p2/yj
e9uRnyjKRw0o8drK+NwS+i6oZwPNyKYB+SLjkBPDXxDXP/ddUC5cqW5xinA+AnWu
LMUfaj2SF5t+QTd/lv81XFtMpA/l9JWtnwqxlGrZmsHf57nTxw2JXBgO44KMmbSr
sVeEJqLVPlsLzXK2q7NqP1oNsppnp5fL6U4ZwjpR1tqv6sBBRfdfPSnn46dkLG9a
QGLGy+CorzCLZ0x5GTIzAEcgRIAN0UMv0FX1EA13+jUUsBFoHVyggBrD5TktO1Oj
cRS0Eu1koRTVfsJPyjZKc+KdQOkTCGiqLDxpq4rwuBHXwQZmNxsd8pzlWp0mHxzL
kPCsmqTUxYviZtVwBkSRjfqKqnKljgpokW7jJv9ySW054rhLhvjbYdK46biKWJvr
+HtEa9dKPP7sHR7Zo66vqENOd7C2sPfsf3yr/0Jvdd8bnsv8547zgYtTkmJ/FmDs
jgWM7pQ2qOeIs4h2C7Afq6yC/Fp+nVv0jBMjEfVerqV6vO1ZvmiBS3qjrYDxQ7yG
YCwLuFRpHw4QlFwG84hMS9nJTttqzQmqTQvfyja9ISf6E2HRP6dW1qPjym+zfODV
3PUgBMKA1WQ3F2lsVCtqaezU9/+/od0Tmtb4cjllOKLeRamgKpUEbsLp+zxW0ZVu
RVlZWlzlGI+DVE1QVrjIUa2CcDVKewEoYIREC8LsaLsrEPpltncpvSg+p3J5LlFl
gQsCMrLzDthC+kJItqwpy9G7uwwAwYe8m+ZOrJME3w+1OdjIJ1gLwb/K64S1wPt2
+eiOOdsH6t+WgFUdsgw2sjgd4PiND5uC2zb4JN0ZL1RGgYTSbhqL6q8kBm3bmxaV
05Tx9Qv/CTavk9xYrgXpdQs/5lqiIQ8T+pvrbYkeevM=
`protect END_PROTECTED
