`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axplQ0Y6tB6uigR67juUVz/6APhDVTKSQL/0Eis/Xo1cA95Cic/un72ubECA9idF
dBfzOtwwbwshJWy1pE0Rt1FMihuR+wcNWbiB4OaA3y0JwtdQ6PsfJwJ/9TPHXNva
oAxhcPL3wyZ3tTn+KzIsM7WJYgjugmLcihVhwovJ0mMLOBLEnM/jugqAobcNouDc
MH8M4sXEhqNyDNdAtrh2wFpaB2XtdzhBnfIXDZB6MLes0t3DUghco8HO2hnnbjuR
9O4QDA6C9nAl6Fa9P7qQR5ilE5RZgSt5yD8gHH/hyMGjLX52odjHF7GfFAUAAGic
MZqkSuqPDgVK18+D/RDsDx+MJBNQM8zIkFyTqGC/myI1bcuWSY+yWTxmL9FVFnKa
81zbOnfnOo8YUzfnVtL5iT1LN/6w5ty+3HG2BG6dRpXaC9KN75m8xhZqrqLc/AuK
23PnLrwJm77QJHHXIEkXcWf5JnonwLUp6dvwocpZXLA=
`protect END_PROTECTED
