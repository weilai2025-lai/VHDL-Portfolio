`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZgvTSRiryHoeFbcLwjejGaa5lHdbpdzB2OH27zGmAc0mKzAykji5VXoOQyypMo2
wve4VoG9RlmZxCsSvrgPewaj65GonczAzd9coJbf8/fjexK6e+Zckg8kG966YdgO
kFGAyFvGGXdtFJBteBgaXZnKFnaMwViOVGv+r1nvBKoxEC3hxBTQLBedFfsMX4ms
RB0wmU4TbN6zP4iAnkf53gEeZPoa2q4D9jgl4r9vNMs1GN7QsWqpkQJCtk7BWdKJ
bqHctZ/k6bE0Cap0bF6K+xMtaXcXKwRBZjAuzleoNX8KI7oCshrwvV9OoIH8y5G5
sGMbNMhJ1BwFkxKfSJkHfpFSPK7YzKUsxINHBGqczZj79LC1q2Jnu1F4gTlrTtCP
h7KfCPrLEIYFtQ6u9M/QPqHvpNVguTNGcBSrl+5ynFzy9d6WUtd9Vn395xl3umlM
n/etw2em0VB06kOqZiQ5Q6Ky9LmAmvvI/aDXsxIe5kL2nBk9eahUMOPD5q8u7hw4
JJMaUp4yX+cosGb9KDXBBvTs+zvo/31b37TaX6KSby1otWfHB0/XMSVSsIzQoDe8
L+T8Aorin5OfsFW/EolRBvyFtaZF9INhq3uiwnWQF0oyWqAKwoK9PS1BWcP9wap5
gnAjlyBe1BfqEbe1HQp3E/deWRQWvL/CREWIaMDzHuHSnycvIDRNYCxXUWofmBLa
Ds7+tF69OJKj0BkVjVUPRfKRvkRzFv872sbePART5+5KCG0pxatxwfJ79kY+sLre
4+VGATXf0EA/aff+ahqhBwgSMNrJy55AKQdeOxjYQrpjHC87Z+pEPIoM44ykzq/V
vhmFgljZ8rBZSkzL0NZXgHFCotSQCbS8OLB6+Cl+S3710RwquEhUeReY4SxrrXww
uu+7vjvlwBgZJ6cK3eGXsteYiTDZzx+2QHcTzlZWdPzD5Lo1CNt4S81+uWLxQ+e8
2ESDBtzo5HeK1IyjYv5cOQspao1ESKD4d6S28CpH2LqC/b9iTTEYAX1V1K4dTPEx
9QKqrfzkSRf85nqSY+qRgGdPnVXRAxo6K0kE0Ar/dlO5DzyU67bxpjjKwPypM77T
y53o0UVkDu0nCVdCGDqxHe7pkuAgJUkJPcnAzmshYphvHgBx8/QljkHkElSVMse0
KzNeVRIOgQcRwOP9bGzMGZPNdpc4TB5XYaN1mUFabivFNNx5uGJVd1CQu3PeIlPK
9xmgqKRCLLaSL8odcqnHPzsdnkOx4Se1T/ElZYEf4v8WUwPFe8fJ5vsG1uWv4xjv
kL8Lwg1/kAEk2IqS4fMCq0gzfKZ1VwkKPKfrN52TumKaAyMXKGihw9rkjNnQknbB
hmbseeQt/Xd9HhiVprh74kXzec1Kk+UOGdOrI2mXN6TQ9iIp3fVz3Gega+gwYDYx
G9+VA/Nui2mV8bWaQhcBAPPd8Qu1Yqyx7qyWeS4VcpCRqviBkDNqhqyOKswkvYWi
`protect END_PROTECTED
