`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yi9uveQTWHO5CIIT9CQ3YKxIn8lQt4cpi+dGb+QBq7iIpN9XlQB3CZl0ithsflOy
7AYLMJiwSevoVSZ7DBCTR4XAAEP1WkehFx7RIdX98L3tt7X6rwR1SJP59WAKdOmw
QZ9tFZt4wBQlAxpxb9i2qgDV+V/ISEAlEcD0wf6qMg7eBJHhfyWOZ6Iw6WuEUSKM
mZk/ppe+ag7Tmez0OIeNvjTqM8KQJywEbj8L5mVAQ9T9z7C1sHNqkruTNNucdGnS
Y8dR0fvBG9AhhMZ7e3+ee1EmS5pP4yegJHK3C10/fCWnOZtTbyf+pY5xf9m9liJK
CB0BIF58mJinaGqDakoISEIrCEd9A2CNsV3MYiuMV4hMakUivfWm+z39WLi651oe
R54yRyMpM7j+TeolP/MXaKfpGbyrnr5cZ7vUwj/8FYwmgsmXlSlVIbQLnSQ+19cM
DWVpAZxt13HGDFMKp2nj1CCJzUt7M9nW05hJ6xtoSTB3qbn8bKnhicEMykXwSaCl
oY3QJnPmsIh/BEAhALzFXTpEgXXJWh+GYvvQr7kI7wWWGjuS54yrf4B1ZSfhuBhC
sEL+O8W6IQ6T+f3gttryHlA4sn7aX7mF5GujwH7iFPufnABCnNjwsnuZkuby7MIL
M3ZYINwffFSBn0LRs1Qj0Qh/ft4HhRWRv8Enznz7WNQ2YCWj2djuAzFrPSfZJI7y
gU9oaq8uen939THBhVdty3gezgV7az0sQWEzY3B8kVPqn08ETJ+s5rXp676KzbV8
frNy87w03eH2qfNxgrDVhAOZ4OspBI+LG2tA5C0yLW9viVMovLQ4/xt1HobweDm6
gcrlJE4/o93grEeqSOj4hKby5tJLu5lbq2v6Ji3/fG0WGq4XiuqTLgH2DKddWPNg
w0Mu8cm1p7zLwMIX8nOnuRihEDK3hPTpWyUEnDH3LMU4tMg5X97/9Swz+74+ppsQ
tlzCSlwN7wpjIT1nB44TDKacP5WEt0Bk/XyghB7mpcjKsYGZB+GKJdY6tlpzEcd/
PLZcEKBo1W2rMxFn5bv3jf7iYseLhX7YfQqlm1aI7JeCETQPaWPbOIF+SRiYqAQn
IJRQ7TGF6NzKXRiZfEBmQidoZaGrs/z583viD2hTyMDlMx6cSSNhNxQKvtVQr8eQ
BSGGdbSVCAMJ55nnAMStFi0z3FeIb+NLaq7v63R+yuQD+wQK+AZ84g60kCE4gLfe
TrWUd0bZ6DyB3nMyHqG67dN5yCzcuhF4hqI6QPgapV1Uu71TZkBaSY2NYAtjmH5o
xHm/czLAopJKYhDou8swilvs5q/dRsDztzqcyoQUzLQ81CCw8fqh3RRxqM8ondXp
3CZzffjUIH4/mLFzMYhNvxyMyQEXp/Cr53fu6uveJvMZ5sjbeY8gDHG43VWLwR4i
D7MDZusa3Em42QA8l5zrS7unPScHcsEtfzZDsIgyqwJE+NgCwDCGcec69MpaODje
`protect END_PROTECTED
