`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
om173DwT15glTdNtqU+fsOX7qvYXqrHe1Kxq+XQfsY/Oxi0LzLrhX8rweo7DgId6
PY26wWN2Q38+U7nE/0rBuDTlH92xZFVLZ+tDaQWwVHT2PassmAY8PClVrR9bdLhO
e2v3XKuHa4+WkTEu/fa93qskjSp88j7HgG+bJwdmDbv22nFhGd/rl00nt5wYEU0Y
DtZ2fV+C5P6DaUoS8s2nwgUoCN/tp/NiWfcycVkMfttEpZ8Ld/al1lH7GTcOH98Q
my0ZVz46vSFSKrgrHd+VJ9VvIJTImEDFN0wVB8Ix5VOQ39OQmOtpFl0rguqqpwPR
UbMNGDFV9Is8eF2nZGESdeHyttzcHpeZ+lqCXxtVV8I2aTGYCtvmNY3F5TCqm+Ms
dM87Dp8ijBQyQ1yGYlskulb9BdsclAv96QLPXm/19sqxvfiz2BIxYzfzXGNu2Qsm
drzDkw9drXZBHyQPUGdRmC4uLVe3r31KnOp8UzoRZQIqGJhMYWzbK94GwA6hAA1F
qB/47Ug+DebBaR73Skg/dlI6rMp+3uEwwj5Lfa9afUTrknrWm9fu2vN7JmpDUn+b
EERqHfMiEHGHY44yciRYtg396l1SQ0/6XanuejfLyCawsDYXc8jIHwlC2/Ub5CNz
Q3iKCIwEROsTuU66wzRtLbTfBg6GcZK0iHtVgdxujiv/UiskhE1Y2syyuFITBTfI
h+hGGWFIHdColJHWZeJ+A3wDXNbcNKzaIO/mjteVYXriQ6PfaLA61vsh1tiNgVEh
DVFWU2XtFVDUmLsrG7HSkGnBW0N0NEwD/73qmlDdWyjUNmTLuG0eflbcGI+PO1bC
OwrBovD30DLuK9gLaBY0DUKBuyIsXEQGod15coj2PgG4eConWdBTsdBXx9y4N/Wr
sNUZPob2+qFaR4J6UmQWfnsp6MCn7xLFCAIE3B7VgSscKx1epqqNNB5CTZVpmztg
QoX4mdDB0Pdml3jApME3xB4kOSqs8gZjt8YIMXXAaoM/NFsjMwF9TH3yQxJjTorj
ouUPMCke8qX90nR1p7wUNdtLA6ogL10AOjV44js9/IS0/KhS26Hep6ehdVMOTRCO
AZfcDaETpI72RSxEQ1P3unbbtSAkpjnOi0oBpHm+wZVBi6kjVCPfyJ8MdCNRKiYa
pFaJM5cpEFvOP0juTt42g4/KD/GulBLxtpzLpAiSAmqkJDQcJGVCb9r9Ee16fBR1
YLITeCg9/OfDzG6paGcC7JOrD9iDUqoP9OFBOSaGyEBDGasubWLo9nbFhg0jyOkp
nFGIsQpnoIdHF0xvdfXMFyzBcFUjIzhF4Y+g4igSkp5Otnn2rXxYm0JfADe9lhaU
MLwDMu5PSQBSQhkW3CBc0XRNOXPDA/106nR/ZZVmrZ7hqOBJj8ryTrEvKgufWJNk
oGPvSppgRes5Dme97cSt9z0E+4Rf9q/WzKgwfb1S8faYHr3OGRWU0M8CgaAI0KUL
Zs22gmRPIwj8kWbc5eewzUOT6HjYPxuEXNchuU8O5XH7JWK6nnzROdPAg0rga56S
FIo8q8NbjlaZMLjW+uucfujgHzNMvqNe8Cix8GP2c0OxDMc00sNo65OTHXs/5/sa
7EDwZBqd3r6dhfGXRyvdHnvO6CZ7M0rpL1fgZaKQffP+cCw/EvIkMsuyCotsKBqh
2+5rX+CiRMd7aagKTXLF5iQrSf7Sq4AFXVNkHQ9nJ1rrmIxLzs1KD27Vj4mE14Qi
uvT7ImFGuFGDkwxTwfPsNxzw3UOkHyRtEmqHHFlH6GqjIp9bQWj5hup2uxzysdly
XWTW132Sud136eyf6uOZb28Ou66Du6cnTGZ/2+vuVIo5E/i3gxF20CwmKGOj9eIA
QLjgg0Kd+S5KSXMNgr58/lhpiZt1oU0yc6GUpf9ChvvvBcmAc6YoPMrrpU1UV/W3
Nu5EPR5gHpu2xvd2wRXRkJxgdPimaw8c4BjMjCOJXBv19aXR7giuYoMnxc+Spa2x
AG56Si6tiT5HHq3Zkh4iMnfr/6sGHzKrhzUj+Q4HV6e9A2RN1u1FRtT80vJ8R/oG
zM+3U6xfl3iOVRvRmhUR879yflNjHnBy8rkX0JmBECrKA64BUZXw7bJye0XLK7MK
w2ZMLsHk5AkuInZtoOj4pvzU5UzmHKbjTHkc97GfFrdoTaQeFMwe5TXXA57skbSj
4p6RloizVGMlEB2XiP16DCEJL5YJXHXVYE6BK7iMQG/JeahDujhqMmYCX1J5F4Rs
krNBNudJ5F/61F20tns/Ze+oW7xsLOSGGbZE6CSPAnWH+YnIwuYxfheX8kCHsdJE
6KlxZVEruSmw+wIgORSI2W/CzhBv/7I4JfpsEhw2/LDqKeMCBRfqCapFxVBB+/Qa
sC5kyHtcANJVIwAQwd3sHzPL/LbmJXYe9qmXrEmZrwGYKu6jKRYIlQU3UtBPBedp
sNAQh2iVWpUr5P3MIRndgHEQTH1RcbNvPPG21huwsPD588TtOzbiksZ3SCb8FqMI
OKyB9uKUm+rFvLpFFle/SmiBYDbIGlZIwZul0wQZiHOygyFr7ZT8VZIl8qCZaQ2f
y5YnP1CQ5cbldqmvXsQOB8uFCXaVFAiP/U5NepczHdoHAV4UnYbTcfEPdyBPnvTX
MJkRK0hNcUdzteLRWP48m6vSmkOUo+F2U3eQpHwwEF+esAwQuj8v40PfxCJVtQtd
8JQ5/0JDHXupVf8ROUpIP17fwDQLxmp38ES0vzSHEpskGa7t7QKH5kyUdCojRZKD
8ALe1wnQa5PmAvC11j7C+AS2BdFHWFSKGXVQvScu587mhfA4gEDsDL3sNWRAHS53
0CrSI6mkpp7irHUmpofReB2VwKJm2DHS8hXqcWFTAUewyR7qNgcQ6RJOcLm9Wo6w
sKX/wzT3J4s8zAZeguy2vTS57fzEvdYrthzWb3OY5fenDsk0KdfXjLPoTnCQdfYk
2H2kRLWTWezssJo+GAsSe4nRgXBU533BSYdYBfZpYbO3KC/vBUpei6Yo/xBK8p67
QvcdbaqVtqx5X+f12KW4eSv6YUwcCQjSX1dnCV6UkY4BA8i0gZTYFA7ZVUIlwdgG
RyveJ0hIKLYn6F6ILB8elfWZE4AOm/4KC9bEkgzUt92aK1hwSS0u7J7ffi0924U3
WY5vDRbnCjSsx7vPjCEZ/OcfM6gdr2ngiu+CQBgyFScWszvcDEUuzrsYbtRsj/ud
q52GVpDQ73HHXlBezq6Vuv4kmWB8OUNi51xREHNJMam0EWCoOuGy2/FoJWf5IpPm
mIdBH5Eadi51CWed3jlGf9DIBTNdJGPxDHUfng2vlxQm5xcCgFbYbSt+3mmKTAvT
OU5XgYEvJG4w22jHqWVY0m5573zc1xc6eHwdH089snecFUuuE7wWndQ+7M30oSej
o556FQm9ZacgmFsAxW5P+zzV2YPY2xoFGy3YYBU2gCTphOZ92gGZn0TEEtYPI15c
aJ3VbYY1ft3AduA0nN8jWPEtHSS63MLPBbvrEVRh5YGYXBwL10dCkAx/Tojk1yBU
fXHqh/nnWP4YqoK0T3eOieQmIb5I9mGCCmFmNCeNhsXW8MMIhVX/g3lOoaCbfMyD
jaPgW2GiRKeFhF60dsG1+kKTBHz21zYeq6TVd7r3/jFu8cgbXGaTxAV8EYimI+NI
wQj2faszm7khJDhIOsCMoGYItRxAZxLmIk3KQxa/JHhKdoyK0xdCHXyzfjYi0g59
60ehh7f/pNa/O1TbvteJ72kW1clWNgExKcxsx7tgO6qHVObgZoXI13NU2b+dbWSW
88h7bYwkkQ9mXEL1KeZ9TVlTADZeMbjNxW40VsnVf9ETGDyG0EjCBpFvhtzIe+v6
HLXv7QOPntbQm4rk0MSlegvKFRgm3TXu+qIC8BFTuD6t0eTN4aVlbKTg9ivJLM+D
xwtrTYLeNcYgEhbXts+r63if7O612SuRuEvirrltw3pk2KXF77u3mOxNW3gEeevE
yYcNQC0lKmqvtnkLuqfxdRB7A7pR6p0K1BVCpSvTdmXBCh4xST8aDqiCMm/HT+/1
+c6gk6ncd5Q4UwWO69FOY/R/LobVvSzpMc66MDDPv3uNTg0/zlFy3KKO9KplPunG
7DnDW7W1mJNhtGBMwYXWdKjPl/treYKu7Fju1xbydqZlSLdTL+IhyYevP02iH+xK
+RLIREKKYJqz8fyDT9YFOzOMuQMNwKGR/5fxO8zWHfQfSo4FGdHCKqIg547hENSa
Q4c1Hu2OHjVMdfpGTG3n1lRE8PMCgWW0MKGDPWwKvg+2NHt+UB6iWkqNb/ajeGIV
QousXUN+9yDo3JJB/f54B7SWFvgrp8YEB+Oh2nNkNHKv//IzLRImSvCCHuKAGSl6
t5LZyCfdWIQUU42a0x3iMrXUr1hhFF2Nwhut4ivq3cJ8WC2LcZtoMjeqFx11T1ew
qakSPwBClq8TwBvnKkihpRaq27PENOcXu5a7kpJC3YGYGTk2CfIH+Rb55SX4EVLZ
qrR+h7DpJVgyJk+5UJD5uGwd3tHecfDmOi9Uu+837GzuHhxl8Zz2IY39Lxi3jugn
sHYwUBvR+ZS2s0EL2F8/4vc36ZvQuaiLzVj4dq6AarHRkyIogqa1Y/Qt8QQofIL3
gIyCm6OAjHRtwJQuaKW14WCiiLtBozgmf3RVGJehCaW8mc3o/a1wVhe0QHPVmGPs
y69RZXe2dxHepTO2vyXwiHb4e2cYkOzNYkwbrZCN2+dHnPi3qrbB/MIWGkzmU7OK
C6+KhmCQbbFSx+63z8q47gCm6Cs3ZaZ267XFUboLkxFs3j6u5zrNi+TWi3neA3cj
k4PodMzEIj6i/uKwTwWMehOqgJrL5tgVeO1wZ8MFmjuYmX/8aCasRanSItJhDlw2
VgtM+XFbxt6CVpXbu+TwHC3JwrVCOvVov3zHt3WiNPk6d3r2dES2XvSP0ALG3pma
sfhW1LxdwuxZr+ZFPaNFvmGlcGb+L1N1uYwJatsc1kp763Pk1H3Bj+bwSI8Dn47o
GDKdMWOIRFK1K+KJM+wyfiCqHg3FnDD9dh6+nxe0WzreqVW6KoxI20/EpFDHqGV2
83g5iyrZLvCpUDpL26H7+TBwwkSX+zVMaIX38TpxgIVeehTomvXUJ1fnNS6NBGDE
99IK9nKIEtUBpfGGkyfoUNPujAIRrX+YLAu9sw2hag7LiJtvwV0m87KQOXbluHE/
ufBZW2s81qns9iPq6a1pqvuMHBk6hEKOSqsieFff7PxwJjTQ2tCm9Lmxl7vuy9CN
1PECsjkEW385/eN0F5oTD/Zn35M9oLrOb8RIAYk0B/YHgkmxoFwIIf71k0/CbRnq
LiyIrOZj+QgToemr+G/O2SA270+Co1kd7uSB5ADeLIabaIyo4htcbsZOKNUA84iw
zrEvzp00g2ku+xXcSB1pEPcW/2gwBjF9j1M6DbbH0ETQqgn09aIbFhBe/EgjdiMT
GR/SSRu1t73D4lOKCIe2MdLNNn/rKezJSBep2vJoxZWIk92s+iIyuLWi7zDUp7Fv
LTyF1312rzrbhnIdIV8bVlGhPWIJqy+7islfVNqCMAQTPPNz0WzNaL2fD2gXWST0
D8XGkw8E1tTlIxSiacqBC1EuNT8ThkyxvtGif+XhzjAouCy26ajHgTEIL451f8OK
IVf0NDLkftXMrgDE37Chan3fonv8nvxL9NQyb6ZO/YrRkOOioa3lmbtsyDvdaKn4
6M2mRJUscpZiQG/MiO6YPxzFacxU683ZNoCS6j/LMbqfQPQobneQYChyf0cm7pW1
zrhTEENUyzQ22was4UJUFz9caNgoYkA7gR+xiI7bsRG2NRHiRSKSFUzR+ra0onaL
CmLUhajd9d8UrmLI783KvTnFUFhUPjY2PhR1/Hec4Xyu7yIHkzfJO6XR5aFq4QJj
QRk0CNtb61jXSHaMT9RU4XGyWRWpEBUkY8EuG0Acd3AHJTDaJ/n9AYyZDEK71+dO
qYUOc9ZPdUVaYUhT184tU87R1QU95sLIj0Q11o8hJDgoK/V+pAQDvuhm+/9qk1ar
mR7txtj7HAes/GwFxixy1s2NKI0us0FvtU4HXZKQfGwWve2qTHQ5RrbDcHAlOJaO
5IxncbbJsWj9KYLXPcjfQe+iITwWSCreVCQ52VBB5YjoS8XzCrA7awS9SGTYv0wL
txNPCGxykAtQEItszAWYUgmM9s6J8N3GOfKS7xFYJwB8phaFsvfPaBVr9VPLa9qg
IIk535a0pMGKb3izHmPRqAnR/+iW742MxOF+k3yw47PUpvdwwZGvJSiigc68q7BR
ivJ2gVFcA9DgXWWYUQUFJOS60anzwAYPJa9ChBjd05uOyoNs2Q2zX1g6G2C9JN4j
UfTmv4xKbeREBbGS/LAHR2MbKeuSOCROmcKQ/TRf9JowS/U/ogwDd/vg1Z342F/u
pO1tNn72cmxCkg0vL9lNsqiozBX0luKbEu7Rz7mGYcjsfzHGU5rgkckEf6aoytUa
1FZUbsxLl3v96eQiCMwTMTA3PE0HUYhVpY23Vx4OOazNLhQRNWLm9BK60MAbvQ1z
UqG51jq8IOo0BXmJtzjuxN3/BDeFFUFeDictKhGEiwFZ29DBHRi9B0L/zHkVboTj
y99vTVEWxRzfXQTpTIPoSnnUxGOeX8pfkylmx0YVI9S5LHjww1P4C1MCzpmAd3B4
xbX8FM4NxdnJxRUsT9ByV3mWyjv59iga3Q6ZXkPHyKFMg2IMfk25gQXid+Yg7qZi
vEZqswiZUV6GcgNkJbJtFZUfSwgKyul2cgwG/kH+479TB0RO6a3TJFzJDdNchMpG
2ilDhQpQUnW44taaFwR+RV7C7mzSphx9zLhO8+DmZteBYn9bXEN9eYxr0nBpsXh2
RDvyoSlNaRViip0h/Bc2YkiRco+Ofap3GmJlt84wEfDQZ33joDxS3zRT89NEksJn
fmIL5glwO+FUP/nemLMa1dpuYlR10b2R576a5kKJurjY5c6ZCt+5ccQOnwhYKJBN
BtxrCMFS9nBo0aKnLjRxFdA9b89TUcfCSwbJ6EFjxhfI/CpAgetesMSgl6lGauvm
WUXo7l0qVr57DCoV2bMhSU1YSzlpSux3WaW/3+GqNREjS/k476Y1wdiS6ZISLw21
Umic4dDWmyeHDsTvoK87F5HmcxoQ//BMNVQTTpDIPu/wke5DZxW8RocviyZ1u5uQ
aRicJi9tTqMFtA8FNj6Iq/y53gW/Lb45DQ+C8t3UxdIbGrwLMBj3QqsxFVT1T+Ko
E4PZsFeut+QyOa1ssuSgFn+a7vMAsVnMLRVOJqO3p6ELR1SoQbyGXcPLa+FzfuWv
aE8KWML11nvIOFN5WLwdR2VERNYLQzI8dL3p04M5n3EExLIQh1rzWw+AMYPG2P3P
XRKEGVD4R+y2RJG50b5CbmFGlpEcRBV+LO4Ld49aOsIgwo2iBGk6LI6P4vcB1DTC
x4r8A/WMstvwjW/+7iKKARFqZrdCB8+Z27Hp6VaLqpCmq/4M7mAxpxr06aPEaf/A
/bQglxK+cXtomuRklCXo/Ck5cQjhgQstMyXs9VT0BXkT6IqYxzbL/HCncrfjnw4P
0vRNpNyAwu1fUZCvfCMnvnryFSrJcAKadBZZ6KIBq8xlrxMfKb6EhGzHzIyy0TTH
0TpA0HLfWxKLA54brd9xTrVj3m7yRrk4qCaxGbI4LgP8vVgq7IuKwZqEjJPxocnS
qLHmJ0AsM8oPRzGu41/G/XaOck/XRBNDdw1HA8rR5c+5JQUgphK89NayPOOviNMb
gqcVoeBRdDe8506oMfMZoroNBobBMi2vBUCDPy/NB1qqg0YjneL84ZyXLG5HEi7q
htYbiSA1yQTIr0T1ZbbKSvPUSSWqQOMMvR5CGPyNkedLTDnAwwbrs7wH+w1t6wdX
OBuNZxsNrAd7Kgg31DVoNq9vQ5ZmGjJKtXhAjZU4pauqv/fzoC7rTBdfDi72uVGr
vJemW+2VBTdlv+1f5bs+M8Weahz83CQZEoUfeybWdzzp+IzNZliALpSJ8CEqnvFd
1mbgAVIeyz5wOj6FxuWhHuU1UTyoIieF3yKHQ0pxzYYCH6Kcapuqmibie2WN89L4
ThsGJkbO2mrB2CQYX0BHQVLEIWLAcgKoqJ4TChRGDR5LtAhLpZufu23nxcUIIiNB
OkunyI7R3cu2hFHLrshWE7hgzt7Vz444A8XK0CCznGRDk7vg+ypR3dJ5Hb+aY9i5
uief2SBIykKkoNBGjdHAudDcJdpVJMYt+iae2v3aMJykPn7Yx7DnzIaWnGNsOfaJ
sszpp6NgB5OeAz/iKcP9zmSIxI3f/85huG6zFNiyXPJRTOofMaP5wfq7P1SWGq9j
YTaab3oKdc1Jbi8YQnCL/kwwHhfQIOOIILwzuL3dMooJNBiLfJvBD8y63pOQ8teN
UwLDYWC6E/eI6qralC0WGb+5Xsxb9VkNC2X9yzsWZGFYeJbtj693LMREvyg9JGXB
ZzK6yej9lD0wy93irT07i9F1LkOIE6nOzEbVRSYtUGd6RkO+K4NydsKbkbBvzVv9
iH7EdvhtCUIHs1z5kBWmAP4NfOsDVfjwFdk2zFRFoG73fBQBUZ89xha9AAi+QLsi
lYaq4p3+H2/e/7tjNQCnFOuHBWn0Q3+v/oGHwW5vwON4gpoq+bbPnyK8OZvgJckQ
pU3zLM5IZBkzTIqM/hXUPTS6kx0gt+5I6f6T2bGAe0jxsqZWAsDtMJXP7OQkCZFU
Kit8woGE3ksqzQcxM+IKufthj6YtbXxwoh05Opyltx57711ghKbik1H0rGrKCByW
3e9DxTlT6/H6izqIwWA4GddAL3p9kZAhk70ZlgSuBLrjprds49iUem1ap7frK2Co
S718YZRjWY2hicwmoDBAX1OQ80VQWE7R/jAy/3oPlg0TH2UezKBUgK+HP32gtMAs
U1wW5PqYE86Besg0WK0wLMCuES9cGUe4+Z0yfOrtPP8WBdxBzU1doEeG/sFc/Sed
mAHHSlQOPUN4eOQVIlJTdCR9TYVoySUu7osQ/Mlce1c08xHQ085KPFSi27z9svqv
NWfS0Zlb3SC1nLXuc+IjGf29ptdIAknGDS7GtlW0n61IHOUb8CHTIkKqGDThoOGP
/7ZU1x48fOR1xELQpECKFHXgtZzGbYu2LPSzbLKWWY07sb/iFZJu9+WwGADEy22O
0fMoGGsV/ghviw0qZ2cs5mTtKFcc8y83vV1jPZuhLcpCj9ABpLU88HglplrnPgKt
OFynuZX3mwO4+M9iugecdou8kxvnHo/j1cdVCVPJxGLU/+wPrMLB5WQ+YXgNTKdP
2J8qR+NdYvwaGPGFf4wcoCiGccdE8RupA6EiFloU5242D47V9ooGpxDIh2vOYBWO
XQHOAIZ8Rxiz0OXVT3RB9ZJ9DMOpydcdi2oDrkOXPttO2iNwqxuYPaqU5dGmJzp5
O0A87jklSRx4ondwlYrGxL/A8HEL/r7fV3TCgzuGcXOoNlWvT+pPPJqnAYddAf9c
h4Xlt8FdOjt/zSKDEVC/249wn6/InXspTsjwHaw7UpCuco01YhYcIOVfNmA1WBaT
pTYZDcYo/FKT1g7h5kPaaGG6oHiG42qk3ORW3pAuBLhQtP5JUb9aTiNJjOu/xl3l
edWyDfXRtt2u9qNj48Ta8LE94LuZHrBzXcJMmBEEsMT7FEKEI9wcbLzz18eweYWt
rzajelaAIQpmdV4mFX2IN0S9/65DKSK5QxrVzI/WkumzhsdxPGS3aMMjsN8j2nM1
EC5IkoJrMT2T8TtCGVcyS3y0B7iOIv+Hzp/S1FyDZEPn5fE7pYFvv8nqMyzUZgV2
QI4XIISh1f0JUlOVSh0hidQRvTlWAyb5VjK5ZxIXNenkm/ud5S7TZWdWex6jCIJo
xZiFmQAR/QQGTQfEF7mOSGYJjIxA2yFS86fFiwh1kRe0uG8ZR70mo7D4cFM3s4EZ
2Xy9WPi4ZIeE633Qe7i4SzPJ4/xVMpZGrHvxs4wmJpegQj2d064SFCB9Wl4kYwv7
iL8PLaedXQaM7Opa4spWQXUGRmqcgJj1bbb6dvt/M9StT0PL9HJKd2SwsD7IObIY
1XV1ShA9U7vVn+vYkIpa9CHzolCG7GSoYV7j+yNok9dRpA1jYspAoPD4+CrwKS9Y
Bt/aM2B6VbdkZE5OeQRdGasxqiMHRMa23PyG7HMlalEVerk7qDzLw/rS9ZI1feuI
U4RK/2mRuKtfOenmrXwU1afSLF/1sA9OGwLNrdEJh4aLVmKQETh6FUggt7iAG9dM
FvMFAxsFvhThpavJ9t1VD9c34WE4oS5Wy1xnpp2eh8og8qdtzTYokUUDB/SLYbtT
mTHTelRhMv/MbJvrQvHn2/O5ZAsj+q1i9MkrPZ8d9RCpCiF/ihekttyQRDrYV9rU
C/3Dv/sSzx2dQGisWeUh9hXkzs8/I/YjgKZUsYa5USnD92KENDzPkNrEEFS9FJ6o
03WPJX5M81l8CR8xtVn/HPZj7WnvA3UEP++onW4uVTwJ5Qaz2La6DmtAiknNnx8G
NcW3XliMLlp/LpYchVjWYu9SUw/GcsaZioZMqd6U+2z3ihu4nB/gcAEkM4qJMEDH
F2VifKrOvEOKEFnI9z/in4zVvQ9JiOzIXWsnuO9AhUTRoKmKtuFFWi0OnAYMyysw
jXFDPcIjSR/lSWKE/g7iIAXdur++d1c1a466dZVGHzCY2mrnNayQbdyo1buMhX4m
K/ryqk1qsUBwp4DlTMrGElsbUeu6/bRPxQdUO6Ubm+WUY5Ej4KwsW1D+jHtVCH8P
9kvscRUI0rgCKWOJQncIdSWJKFqlSQoxuNixhtpYInCEw5w0fFamrBn9ltqkCpmM
kfQd/4qC1Wk+p5UQz6j5u5tTd480uXkaHR7d25kGMrvhvt6+8T8024Pi/6PaUpsJ
IfO2Ad0ndcWao8v4LiOPZtKRMb+/FCcB1seVjG84aUfgaEmM1/YDEvrTPau+8EZs
OfNaykrBtrYnayYO5zuUHx7gsbrmZtNkOmdovSmXYBcrq6z1dQT5UfFAR7vN9qXJ
eCgap++r9l+9IgpXqBjjOdsKC7oiMa8E2pW5yQE9SFaezAz+5JhMGq/xLYXunKn1
0Qy6s58CL4tknE7YGYUB+jzrLtQHseGutJZh+9eoQx8aadYC3HLtvluhW9M7OPxu
euBChAZic64BWeV6WeoafpDTxjS4o3sfnU9RIP2Q0fb1Gsh6JwnghN3ndMWDiSJC
MHRagYZ2jwxd8YpOPYg7srm3xQDFp8Sn+kM9CbJrqWFZ7DTd236qXh4pY6/2NcO/
RTS22WKg5XXZl23cBrtXKoKCXfmo6GbduxieP7qn/CAc7EmA6JTW6aiKCl4JlMsA
E/iudmODJ3PGQfVa/S/0cMuiUvmD8XjFPB2j+L4sLr4YNjaLzsybCmGil3/RXstI
jld5OQGzC02fMkvvDklLw4qiVOrbbERum5rFtQPxj1sBAXYR59/WSSH7JO7J/nA0
JtSLIhHAbrIwgsJKcmcgAQrgSF23+4tbrDWJI/U+/2MCpSVfRJxsvdcnntNzOPFL
8bhQWCHXSouXBv4AIPRrviT+UnB2TciHSFpsSzoG4aAYu++g/rUHxA21h8vxYRqA
GWBlnOFfiCNApRnI703T11ELIRxym+mfj23g11bvXIYUR9PE6wIN9eoTcYDncPC5
1qZHnrsk1M5lax9+vs2AVVUkkCTUt/3EAiHVXTz9FdAC2PVuvzcDyQJx3N8Ks4Ih
rejBYcPJRYLmWqxFADSA9Gx4JHRzh3Wopv9oRkSWLcp39P9nm+5osM8RJ5tJkFgG
OW0l7n26lfuw6Dw0XeuXg+9E4gsil1/lcTc/PFpi2Kwj5B+RiUVsoDs4MW7/Ujri
JDdBjv49P+ZsTXo+JzRfqBZlS6VDNcEEAOiFof5aS0vKDcYa86QNvIXG5TO288ow
qCFbwbuC4p+J4AXmwfLL7VWaqDaV++LlRUuj1ytb61H1vYoI6V+fk8JJY0G3cK0h
bXzzMUumhcDI6oBiW6faD6VAkxmFRITGPJ90C9a+y1DH2TOOpPSVieTmpU9y50Pj
OkE2QdHixfwm84ZX7/TcT6F0sQPO+XLMnHJpsYCcNye5gf+7n95PMRHderFM0TN3
T3wJZimKG4A8m/dFHJ4K1AryADBf45LICtbjweNfzpXquFmlzZl+18OqXMtaET/g
+SRXjWXtQm5jSwMNFxifzOPREHpV/Hx6mxmHCe3NP7lMlH6hxLqzJ21dNVg3i3Ol
BJmcvfUwd3BIAv94eFtnjOSjy6/bL5ITBstsqmNEKUKbbAgVZSwPbTxLNJtJwUyw
YomxAi3BY8uRyVC9821DdaHu7BvkGcGwIqiPRJBi20kWbPqa/t7fstvmuhSvtkqG
jexh0qqY9mzieuW0gyAUu4n5OYJ55Hzl4+bjhugvVLQNqiHNbjBkTK/63qJvJWNQ
XF9NxNbDdYRj4+M5OBx6lNnbvjQl4Jwin/get5RY001jKVcjuAvzXl4EHC+RWOJY
JyQe6vYT6NA2WqFWNb4JtuQSvFoI1cZn8mVq4qSCgCtKjYmyLZGeswUXxvOEkpWP
n2iIm5OxJRIw/F1H0KDp47jRDPZPGXyEYYlVtiujHaUSpRk7fUY7TMW1a8vIT3Gy
kkaGHy8ziVAd08aos6muC1f3i+d1lCSxVgqp8zFuf4uPBCWzTlC8DqFFDrhGasHP
f2HhDLa+CD6IIhJSk9VDrf9Z9+ELKNP9jiRVDrBLgE9r41iNDGggV5+1WCKC8sJO
kgoF/xlys0wvoH7YZb+ms1OyzP3IXGUmRxSGpXDK0JAJ1KGdRQx0Tr9a5bMCIHzq
BAtAdt1R4hP+dTPjGtqzq9/CeJg4hf7wjTFxlbjshV5/gErknBvl6CCmpfuBN7P1
NBjbaoHGfn35yuTY4UkQ/rE5wCHHq8E16EBKERY9lWeM8A9mQw4r9UBLvZqLTmsc
aOHXc3kDVcrWZXHEFw+B5jvrSk7KgKdsy7FwssPMaH2UGW7ex7Ci3YjfB+tIaAn5
Mo9XZh/YAFtemBVZ7TUXNKhKDaF9CC9fH8w2VpAAv2IF627rwaVIJnxf9JJLXuo6
wgQ/L5FhjPjfpHB9iFZyIQoF+/zbNsj8HNSSZ50eqdKUBv6JXM0rOFO+hfDT0K3P
1n6a5+STlrDmGSL+egRiAznPRnFyze3+acE5AvM+7Cnr1wLQNOIGj7E+8bZwK/G/
DUJ0iKNbk2+kcmUqARZKrZWK8A9BvEssA1ltD6AdGHzHjFWk1ZHSAHT4d/Cg4e96
`protect END_PROTECTED
