`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KOP09x8H0+lOoJSczBwKGDwwKj+hC2f0i6y/cZZoOuVd/ZHk2r7KysImvkGbVgSf
YQwXdMgWhTCjbuAaEoC5JRIFntJXJPMtHvKGf3pyuse7/dOVVEzbrxcZDy8EVw2O
OCdE1pygukyeBre3VZmNBMyvbmH6/uB9xLnnha7Y4Oj9oEcIekXOiWiUZY3P5ij2
m15gUcF0ylI9KRt9XXSVzlGBMMP7LWCQmewj3vO0Fs8s0xc88Et65kfSkIwowuSi
uVTkMI4pmNJPIX/w4VVVlCzMaRtE8xljAIWwyf7YlJ3vFyo+y0v1yZbOaNHSks6D
p7PsZlTJFkcoCWjYxBQp5W4CP6WneGN3zvqDfgWjTiVGqxMjxtyoAhW+S8KQ8SB0
m6NtSxenxOqpTS6uAATuOjM+znnMlGkWXr1B6Koza2ovncfuSNLiVAR6GJ8v6Bi/
dCNTr4LhfyXa+Rpz6UPFxGwLvmAOu4wrwtFQCH0UN+IzwJUm0Wkea216FsQQaY+P
DB1dbWgcfnNC1/qNOqPQMyVenENndbThts+Pe94dKcv9IE/ITsRnSWBKki8k//aL
qiZ5b1zQ4SQQxZ2fqFd9R+4dAZb5xhEoKdAG5wVJ8GiNI1FLhHhFr+6/G5nC6D5A
MfHuSKwEAkWbputP7J4ESH/k7znAmo7jz44sL5QCQEOpeuWBNWtbqL/GSPevxrce
fw4+2dR6dRoNsxd9pqedIl+rxQrpQkrgKC0CmjcgevV7FL526IgLq0wjc5OT1OFo
BO7jLALyamdjYOovLGY57tpvnnKW7/5UASs8VKb15mYBr4JG0WTM0Tf6euOA4+md
4jp+1ISPD58yFOs5/aBhbwWpmnj6qOg1mXRESK+tiP5/KmgKLVzJQ0HEpuZpxu2g
nzmshUGV0XCmWLx3q/UulLCHbWVmifOs8tIvbzRpyfh/vi4wOKm3WtWKS4DNwakk
O9YF8OpLD0VPgBuILmxWEg33kjTkIP3xFq6nKPSoT6NyZMfAWjTPa4e6TgJ5G11t
+sg31gxPA+OXGG9goL2eQs7GdyfVbGpG9aQlFZCR5tFLGr5FFWl/a/r5SI+XR5i8
RLmxqT/zbTbLJLjLLqudOS0bChHJ/e2GPXPROZ8MdEZ/w2A4I1WWjW9V01O8+qW4
bZmlQZA9NvQaxOpuxD34Wo85ue4+DYqHw4GDrrPYrt1o/9bqvIXorGC9glLjj2hw
sMJ8zMlNFF1M1vJF5MIyBXq3XkrZWionfDLDLq5fz+yKdV4QNyuEA/YdUz4/VWzw
mUvJVJVGvpq4E4a6v/E226gx15YAlfODSRw14tNj7SykYMQhdTnf0qppt1ok5McK
7BhUMUBCobo6vDGxf1KVYvUic8/OukSxUysC3JE0oIEAlsb9HHCDxY9P3GhdCvMz
ak3lq7mnEHSyrZNV1a/YUsYRw+7Sw90TgD8HhbGKQvUlSHiCtyWwl8pg+PYuC2Ko
JWACSjIzTZlMrVdEDmOZcKUB61NpOFeLPByMB3TmOEBtZxr6KRqwPFdG7OrX7sQY
CHrV4VuKcCs+J+9iQg9b/xz7qDwEN2BmgcoDggxjdABVdPl3Xy1sVHUbKUnsdOka
LCn/0oATvk+jgPnDh+9yeBIsukHy24vUa/yiHkhgCTXVHjbCjKpXMVV5OP7zzD0A
PNXH2A0eiBKC4bAJnGNibCTP5j5qrfvC2KFB8NmHBf+BrFZmRMx0IlIQqgpj/ia1
7Z3x6sCOBaigGjJyS57MmsUto3eudzzIuqABiFBGPJGhkhvkwnh3eoc8ZRsml3+s
xsj6SyrZcIx6eNGx75T2H3GNj7uYKkD4bUGPppTKk6KSR4ZNS0mzFMCRTy0BpycG
HjV8D1juaNpxrtPyvHk7mA/W8Bh8frsmxN07Shpr0WcEEp61oO4HsrZ0su7yh+do
3SAJJOQvgW3D09qVkZroPQoGTKgk06NBwtL60m3zg+kp9jU/pmv+TTSsRpiPwgn9
ytwxru/C6Y9ul/QtifMnNDJ/J1MOieZl8YFNsNLZ8TBPpEd/Z6rLharmxpb5UtZN
bTlgUTMHhlzYaPbFEzv7VbcilY0ak+9EBSbIBxFi2HLXRgtqYURagSxTANTBYUbk
FPecMYjT18rkA0Ig0RocTKf7IPCqqxptbxUQRGfgT2mKTgyg7sl9wdRj25UDOBWR
DS6fOT1W9ies1vyhz/o42l8ZzZEjZsCQobcdSttHxNF+zDmAe/yPgJh01BRy0DQv
P5uqHus1/7t1cKk4ut/32ZcHBPGaAApFQKOnLxZVqi0b1QRpGVugoI7ZAWVlGrpG
4Y3hjDjjVswMHpLe8+XZmSsbjkfRMnFurakcHJN5fw7c/7zI9MuicTWJLOPuuJMy
cnBjyWoZOlxrVez+0eqBzQXFX/i3x2Ko6S3TlTfF3E8se+0PTNune02LKRbvsstQ
j5uayLBDstDMd/Nw88t096zL9q13ZVU9p6rsYlrOUvrrQEXacENM0nQHNQ+T/iQh
wlJG5L09NZ9yuv/AlaP+cojjL6cdQPpnqNB1Ky86hyc4KGwmTAeFkpKb7JcREPaQ
bRQGkhzl8b5jZpXBS5L1MQVnA+nVlSFrmmJk+V4YCMv3KVG6ihjh5p6Vrjxr6JTA
dJuAj+WQGfFR8zfmhBX6XF321DffI28zCm4LsIsXRfQDy4sQZngBr/3KIk0P3ZAC
UyV6e4KufICbhxVwQaBkoGjRR8kYmvr+s9ETmYGJgwWDP+j9mefDb/E4jU1Y1Mga
Apzfbbr2qdcEV3wReg5oQIzKu/5wIs4DMCtNAlFHXtwdxYfHPqcBsUCjzH2M5Z71
biMN5ePxDJIHktETCbkbUyCA5EPGsjJykiXp+PdMS4wkcvUogkdm2BU/1dENKxun
rniXZpZQ1JnVBJKLNkL0z7VeI8BFEtIhTtNehNKdjyPQUotU9Z9Ywi9osgNdhNig
sF4CI7OPcpJtfkC4aIxPymSd4ORei1x/FGLtdc9WoY4VheNwtXwWpgbbssO78XPA
4Of1pAJ2hGdT/4XZAqmtrBTpdD20oLnlWTzZDYMlrROVQV5/a8FQ8xBd5g+0sont
oapsMOX/3IKvZoVDG/eMuvRPqMl6Q+sGnDP+Hpjqms3wIYc3X7mRPHfpwHXCtDYO
9M95mrWC0RcRqFz5u4SgUHiSbJt5uw91A8KizjKLo1WK3rw3kUPoGRlXo9uqwkbQ
EqfVvkOvVaRbSxzBk8TtdQYPqF+DT3787jUZiYPvIVwV8N98YqUTq6DCeZVfacHy
6yA5knZls8ee2A8p6HN/otQ27Xp/I3ILwG5LUHmCzz4+aaqbxMBOM4EBRXCyQYZH
5Cem3eL4pcxaNsWiXs0XaalzrOCh6a4JqAs4d8qkyY9b8wkzL3UccVnmePuLBdkS
FiVlIUYNUG/LzE2JVxPo4tq+yG9guE56EA1TqSmaZ7vEKOGlGAGrcntj/lpCQpbj
LGuFmfUDl3o5INnsBFj12wPOvIyHEbFyb/HVjoazrCmSdpyHhSbJ9VJRCBxhttr/
iTm6GYwB87ut2gYzF1bWsIbYG163lKDqWwZOuEQli6zgaA+Y0Ee6SGCTbx8xsNiw
KiGOZSp6RqYjbTwAH4CML13AsLQnm84eyG9e7kG/tbz0Ry4Zet2OOZLJ4xvzlXmT
p7dUOHcf4UDd+9Vzw+OyJyG55cofPgn+FZC5ep+fGBDvbs278PerQLSU14AZc37s
Em9BFaUkjL7IuaLKmlyLDeneS/CzZFkyXKrOHbNmorr3OkDBS0LVLOqDPmqE3Pho
WSmhRFC6CTHLEnQgEXWcwijo5dFII58/l37wolYMSVOpAJwGenMwhNY+ImjhTr4F
I9V789+sGmf6sjziV0vVxSR/c8d4XebOYMmsOSroRqXq9rLp+X5zX2Woeg5+GdhF
wVVd4YFTpE/DbMVxVPRfFg7bpaqn8t/0tbBD1N0MA2OeVMkxoJXu9k1jm8U/Tj/H
kZ7m6fUgcODZcOvW+1u2Zj+aBtlfb51o3PZeEHZ6gjKFTSY/7Lk/e9b/6bmhiyYx
N1yIKNkkizHXV7AIW68X7nKq5lV2o/98ODRA33zApAktJbu+Me6m+BDCOjw/1Bwb
CkYouK0KC3HiRHqNZ3ne2hljIykkJpOZt991SCFdeflthqOQGVtElsWVbjJf1kao
MO9/AHyfITeV0bFLMe6jBEXOeqYLymyTrSvkd/L6kpfV5PyP7yCBNHmLmv//QpOr
NnLoYr3IGmL/CKlCDZNrxzXDGjIdFkKUyUspNxN4EHsOcyUjSUSYptHtf4RNHnVG
xM5usok2mcCiKL/QDPLjF+VzbPkEXnWi8k6HaXEmAlDVPemwn7adlDkFwqPfJagN
DQ8i7YpgfdC+UPe7aBsRC/pXsL1NVf6citG1R5t7Y3wr+m3XyvHY9I0422/XjRwW
9SlOiG01EOJgpYqsVLguu764dGakW9sPETqGliOavDywbS5u3C2l7ua54qhf3ouT
FG0nHVByIWskEnc/xahebzOZlsHycuLhnMdvsDlXRvtDCsGGPNtl9lWocrPsPXF9
/TDvLlDBve/D5Qb9DCG1nt/BfNvUkHiMuV7QKl4NlNFjUWEVK3haSe6MJ/Heudyr
EbITWHIeN3zsWLd8xjmdaivwYxNYjbl+8XpG3v83upo3cFT0YY1uybgpbRmUuWS4
a7yBqu3zsQfyUwPxHZy36AU6PbHecyQnhv4+oPI9Q6PCvEeekq2ELGNcTv808yi/
pkdjCWmclYje0Tuf4Rbv8G2jsWoC/lcNSQAE2ipjwhg/u6F92JyXsraTVRwg67Q2
d0siyM/2RxHUerHmv9ztPb4WZeJGwYU09bbSTPOVDkdWxOgomNef1EmgMshUG39R
45Mj8Rlbj9DFaFxzGTivHIUqORNgEURZndAXtA2d+Q/pbgNoaBRT/xXYHZ9ZV1GZ
fJN+akeJIP/uAZCcUrS5GO6vgXserdU0wJ8DPH9TcEu9rk8AsLrDRJJk4csjfhdt
NYD0FfquD3wqxZ8tD9XD6UMQDj6kBvL3I9VFOkJu7V0kQvaA+gG8alI/ACDZUlxX
uDdHFOzJ1N4zGiis61ZGSUNTp9n5ASaGCCuwgtqObT90jR6p3c4xZH2i9vZ6MvQ5
anxX8st1AahOwcpC5yoT9x9l2dAh8itH4Cl/nkm8HVEEnnX58UJ1DAXkyFqmxh0l
hiQNL9Z50l3nYFLp7+GD8xy03m0SiBVEAX4eLBspCLL7pTaZ5/k9ZwSPsTDZTJfo
qU1Uzb8mjOBZ0qmVK6Norxf/GT+fDhzVSLSnNAVEFJI6NqqLtF637NbFjJF5B/IV
DEC9C3/zcyawHSALO3A0ekyFCvxG6bmSAdTb8PclsVm0kuygPowR1IqAs/1Ddfcd
R+s6IVN5E8jTO5cdPvaY3qR+n4Y7gOU2AzIvYwVKAcyulOSi7GTj/RZxEoGRr9aJ
UUhXy44YQ/aW+zv6ZcqZXHcnjbWMlwAV+bsQaaoBFcM1kOJCkOPZtfnO45QmMAWD
DO+WyTthrg1SghG6PjomAsjjytr7XVozcPZRgQbasaKTuE4KV0yZi6ceLAJ8tuFg
EXO7qnX60NmH1ZxhOmjLHpM/g7vID2E9B1gthev+GZW2TtjmKXBkB46Z0efxenZx
NPDKqf/mdu2KHa02sQwKEhCXDc9AqJZ7xnfj7ymFi1bHn1pos4wAcFrvE4Hu33pZ
IjyfDI8ZDgU/LcmzIgMM73KisH4/CytuohavyBy2ctcWwBLb4UT4CkHqgiyI6OF0
KuYBd5EpZ1ZrNuoBzNXCRe+tXlGQ3q6V80iIrNUjdtuMm7XmPnzJiX0BBKFLP2O6
Rf3WtyJE+Md2eKXY4n2MsEBH7xsDiNv2+p9YOlKyAFBGwWvK2NfaTjBL2hpGj/53
X4pbCZYVAO1RGEQ7QRAGqKwljyJAI7Rj2d2wWOcSi8+/hY80flvcyZFgRJccDV4n
ZrJTH59vPSmI33MwKXh0lh7Z6jzlLW5UxZoFeHKhelSxEo8jmA0JjcJv19QTHbXj
3SJYUchFSAYY+9TQRk4mfH/8di44rsJQxoqmrOQ7E0U8mfUcZ/QBrQ1niTJ/kzd2
YTC6stEIHigfxDPyHyQ5So+Zn4PBDkGatV3N5JXEN+gXKMa+OlnZw47JGFSCkbGw
3h1l4FL7sWkyYc32EB+Gi4Gbe6FHkcRbRsCl0wyipF2Q5LRicfPLiGx7uQ9X7YQC
xxMiKDoehFQnHKRaOAebrpF2EJ1GKeCxTAsYJYVZl6wuuM0A9RkJONIPF2R1aRvX
JwF1R/YcQFDrCDvSbXBbaZUfLgHCIb5qGSccILy6jc1jcHZSX8Qe1fiQvzMV7fQg
rPj5GY7/hSVInM84OHyYmzTi4jI7t7emQn05SJRq6ex36yGCQn8ayGMVa4w+xXin
1gj9MhMtS6vYBek6deB2KhXfOru5WfB40dnJFXS4AKpF6uCQSrXHwrHErfVRHG9E
QiA/2pYQd66eaL0VPYJ7p39SS8gv9l5aAXcQ43XIq4eEMhIh5lXdz0/wcPluVxe2
qXVegebIxafcmC6Q16jlZe5MWpfge2DBFqo80zcidiZrXhglKrfGVb9jype23kLt
RF1mqg+2eK3HciBP6Qeb5JoEh8cITdH8U7ytNeCH6ToW9wda7A4p26CFOtc6gDO4
YaU16jTFLsndh7jaCALcf2DP4TPiUdmOIlu55o4/B8iNpdtwproK943qKK6a46+E
ig2CUhu88UeisYM1NOX0Bn1CkGWWWzSGKNG6avmamf62RLto0579S7OX7vdiPaSG
RRVMIZTdMazA0OccOuLUb5FMIegBsgTnei/313p2zdxrPzRtHOapNJNizEzMV/Yg
EtP1IN+T+CHEu15uNwd5x7fZf3n+Jtssfn1WzAFKAWUtznl4Q4Edo1VatYtt0FuF
VY5Lp9HDYyd4gffb6pjZC1xi6PgZIxZvFOKOZ5AyLKCgYfK/J8T6XKMPXad1YWj0
+o/coK+RxUIFKn9GbaPTsVlVzmQo7hX6wHk3UMEk/mJtrjtJM4mT3LCHv/WIRGbv
k4QWgaPoywjMGc2XgCB6gppReIkJNefueGMcmPCXWSfdhqpASE1iJ9LUL2vZeht0
tplop+Iriy6fLRNjh06SWKbjzTDLBbEAbB81blcPFwBj64u4yuASjFnP/4O563EG
l3xzaVolX/axQnKMZ+tj9Zv8wsXdBCeKKbfxBRyUUb7XTqVxXpitoCABsAbAqohR
P9Buqof4DmoubAadvRHHAFVqbEX9mFUGVVhH6YGRg0dEBAUHo9A4PCieqSOn7tYL
2MB2WGWEPfpfbhjTn+2kwy46GLBlYyFawYqvIR2813z2KOwOV0hw5/NwRljV4V9K
Fs8X4thvKk98/DYUCc81bbeEhG3lSJNRYbYCscbewa4cOzHTQrrp+lZzPMPTNwjd
10yD8izm+r6aMSIhqvBZIbdCvLncMaCEGbkU456uLVBVUub1ELi5W1KqiXHkzfvL
t7wOij5PJp9yhXEU6imT+7oGiI3XwJSznGyLfWQEkj9jKAgwIvqZVvNL9ZfrP9ME
MPkz1Z1/sqOm4+6lRhzyi7nqkwdX5TXPDhtJc9/iDX6MxMRlSqw3vjxbIRJHCqoD
LITteAbxrg4eQVu4FtJRS4SX5mLs4trkMK6sLkbvB7fa+LGu/XVftjmTBx4uNUwp
VwUPXFzf5BtabnvmMfJjLc4mNLSvMyICE0h053p0xxcBMARzST4o93C5UrEY6V+Z
fsMFlYj75ch+zIzcvDbOuQ69AL3fpWCuxcctJQYsZbWhOxn6dkfJHyO8sBnSoZiY
4WVozToOp8CkfXfptdbEoI7qZF6Qfy7Ar4WqvzJTq+5SAoN9FC0R9ZjGsTxNFX1M
CkE3yqeC70BegKF33LM+F6TOiWeR4Psz2HMPmxxSW7S+X3DkTeqXWGJ72BlctvMd
U7P6BD7GhCW3i3E5Si0hi5czZ6SoMWdeXVyylYGwv3URw9RW6GboOHj1cWpb4eAi
81uUA5Q0qxC1eHkP+DdDJ8+Jk8zk6jUS3ocnJQdKM85/h3gg8JxE08NYd3xfhPgm
7l5c5z76HUR0W7BNF2za1iDTUrZ42lT+i+yTdE/WZAB9jWGFNiVWULrOsypgZWoZ
AALGTLT01rMA3WRYO11YX9ZW9avw0OuLsDqCm5qusZhBeqIzyZCThIgya3CpQXhf
0M6I4CVJdo2wORNBtd/Q+kH4nD0NR400gIgW+q4sF1+9LlxWpaWVDZ8xqSOAMZPK
+sEO0pOwu7DtBKnTBm7xJyQa46A4g29Ahud3RCDxL4p14n9CpixG8ZFpfwycMXYI
qYcXSoe23AyIX0RBrBHVORma80ti/jZo6JGkIM+jCUwvf0Bt86hskzgFodylMTp4
wqV9/GFUlivh/2k0yXL+AzlNI7msuGt8kzTD3abYhnfsiWalHOVIwl44OvV0EK2G
tH1BzNvk3rRBIdCPukseUZy9vpVAd5qy4ajrMl3cQmcst/BSQZZ8hdvdnLlZd5Kc
Ql8PoYERcrouOWufHT6zGieB/XrqdM4/tGOAoA319sqK+8MYwwj1b7vr5/MfXsD8
AnadDiVnY7Sb2M3e6r/eizpOq2N6kP5LeRx9g8tfluCOev3lvZNSBJ+FkUkutCat
nixA9BdFBCs5Qg7Ygz0T2ckC2r4HaSlkm95Cwl3BRiEE8x377/zNL+2M1wDSKKfN
+A52twqiRa8IjrysK2oG9iuj/HXjfCMM/a7KVgB8U6Ymvy+e4GuZtTP3RpRBEbx6
52uIwtwt87ja3X+fjPxXa3dTdwU092VstOD/KuIuU6TMXN3hDC0ffHbmoSCj9JjS
xfIXqhnEKA0KwDoKGXj9pOXQ1OmkQa5opqrIDRNw7y7hR3v2/B7Fl8RG9/0dPJB/
zBlPsxMjR1ljrOgz2mu4tI7r9C/LQq3NoSedhPZCTwus4TIaUiY35rbbRN6yS1Ta
zASACilV2cuiwqBekeWTi6vvX5+OmcIxU/30F/GqAczgUgJNmvx8ZJcy7YWTvyNU
l1oCEgwB8l9pQ5sREHM909G+syDngTvOx2O6kiWDfeLR5JPSIz3DGFRylSKXNA6w
EsKFTuVhDh5jGItm5Gsyhq4/Be3WspjjT2DiEnAbbVSKwnDSseRzNUGbsXj0l8WU
xRevrsjBOKnVAvB2ODSGj2UAcvV8Z+ZeLPpnxvOHtubmvQVD+qo2OYXKVuoqlbWw
uDXuenOAxf21W1TCPdCuI3IKPuZ7YGf3OKqwakZdevyfX/FIFiM0c0gQ4YiQ4C59
cA1jRxO5TlZI2/wUtunWStioMLDWC0bVE7cpILzE7i2i2YIjeGaqzO1WoD8nm7+x
uPgxfKMA8xCat12Su8891OPZGSRytTgxWX2taPY3BU8oaufaCc3lcJ55n5nYJ/6L
E+9XOgMfAmbeCcS8KFD5z+9kThA3cklxSDEKzajqVZWbfVIuUT6FrZOVOPaIKUZn
FifNYIbwOG+32zUuU4XJRnaa8mfAGPzfHZbPysXXgQcOjDfWxiHH4hietvxIf09d
5tEJELhoC8Qv8lhfc7w9J5vw5vBB1pw+o5jEA1MuDGz5E7FEpGYazK3Hgo2U2YlG
Ay/YM3sxxBZDHM4BTv3wAjsnV/TUxZtCxAVczarSTIprc5svT2aAse/QYYKOaUQe
lKN7EZc0amhqfjLE3E2BmOD9B/g8cJjy379Vug1bzdqptxNbbrH9gJyOJngD7abK
H5nQBRwIBbnzYkALoIzh/qznm5gjUQaUc3gWcHKsBSEmJR6IUm2qMGaKCucKgUut
i0yncE3zxVDEEvY/oApDz6RkM4NcO5okRFRlEnSdZhpdkjJbs3MDIVPDdyNsWQ2t
Mx+0cwy/Ba0OPnqTAB1FJAGX9ltoo+WvWW3KzWIW5nqqilHrr6bc6zD7mqk6MCuV
nk1WluZW0l68C/q1WLBXLlRpiFhon2HER7j9mS3tHoZbKAMwIvCmhBhMszIc+zmt
SXMkUB0QBNUjxaIXnMb9ypBP6NDy76Uto6pQwco+OMSWHOMRLt/5X6DTfRbsaRPl
lsoL33xREK8CUyIdfStVHSp2pHgQz3vfSEIxTusb3l+vrw/DSM46XzrApgMMGk7m
vZwOAW1Z6EwpTnT6EMERNfBsZ27ThFM8sFRPqo8vsvrBq7vJyhuwIKmZm5MYyJkG
b7zhxf9nhIpgmqlbz5GLGJcxpT/FYZNlQlk0V45UQxpBLLG9uyxwaeAYVfdFtidt
rMDYojsdT0VBsY44ieAmjzXrIA5BK3QwRNZEU1XWB4boMI0IjFwSpX9S4ZWakE3P
dGczeZcjSHwIr25YbhGcluaaves5Cf0gLygMafbzpaE7/p580ZtduJkHzKcBzpm8
VKGkIdUFYZmOFEzGMxLI/7/6iKKj2oOlyqGp8i6sZFqTWn8qVBZ7SHjRFEbtDcsW
YUr4u126VV4Wa4SxOOQSMLeBE5Aq8ZiWXolFQc6tzYQTyo3Ws4jM9zgavTMMUtCQ
W5R3Jw9iQfBiTeDpW/PY4iQjA+MVREuo6EjBvcZr4c61WP+yhXf7wp131qaPMda2
X5wvYqxYSi/CkJHI1ZktZMkl9IiRLLLtfIjw7Ny94IZb0r0GqlYoyGSBy8HQyCTd
CAuxD0s/z5uh4KQ2tzoNi64lFujGlgQs9paXW7Bk3GGGHsLgeAVO8R8Rj+hw6Xay
QuDsfJcWDG6+5Y3NKa03U07RTwHZnPYFNDpU0hhHM8jUTlSLir+AF2Ypf/2vNn0/
NKWneiGxSRvtiZVpzYIvUuxoNfjyV6DcB1C/vxN970v+6+TNEhpjSj9YbB899a8J
pg64P+QzTOoZ3e/B+knFM6jjf5z1TvpWhwBhnnmYRXghmsA9UO9hsO4UbeHNJsyt
QhurpqNabUDx4Ayg8pLJ7Pel2OHrvV/loMNaSUiCKm8d1ypqtSIg4XfUoTgQH5FX
vArDBhoMFeMC1YCQIlNxd5XI1ZWtRz8tO5isT6z5RjEdhMSHweF/V6nFMFuectGm
5EB+/AvZpfAskaAQl6TfTKvTsvNYLq0VWKvYiIFjNNoILeV8+zlxQKFzoyb67tQ1
fvh7dD7i0TNsfN9DKKNlLlTYNBAstfmWdw/2T3EjeUKT6YCMRo1FhnwM8wNTVS07
RFnR13K7WGr29Ly37dvXqCgMxZiKjsUEB7Y3hYHeKcsa++IWbDW/eImtivDWjbBB
s27SwPI+Z04Yq1dMYsQhXeAJhjb0OWbWUYVcNNP5e6uL7zLWfGuMjQpGUiFYo/Wa
rLmLkByZTSPQimuORwFZEUjxXS+RMu3LbqxiDkv0joSR2vpmyQDtGdI+xurMPflF
0dSafdCgEJ/WYUg9yncxyKA2DFq89bIiF64bfvNFH8qvCVIWrbSePfPjLjQj2ySc
QvxoGmQmvOFf+ZsHRmC7vxv+cUcLZm3bz59cZ7IT1OEYaqx0om8auOXv+AaMCN5c
d9OXZgxBXrazGX2EzB4Zue/Q9qEn0YlB+3stW1O73+MUyYBLz2SfRs6XyHgu86kB
xDw7TeOhc4e0NPm6WLCpFPGIoRW0wK8xTvqG8oFq0XSW1E3pbVUKeCHQ/AbjWWHj
y44qzlVXAE4ekqpskc98JsxWg+T4KMi6vTlTVP8cKn1iq5LC0sPwLFTjp102+4B3
llQjXajAZoi6BBsyJDWLNw944IEl8q5SSWTQ78sUxzW513YYZVKXpp5CKrpTkr1V
VkL4K2vvBVXRVK6lxcObSQOrgMhOIf1M8XgpTV3rkua6W+B1MVmv9FgC/yv8UTs5
Gw5r7dAdOnsgAeiahE+tjox8KRb225lN1Z4a29uhaWM5hOmhFnHKP006Y62gteGa
9UKuMx2SoDrATsV/6D6SJGzSQDhyF9f2/C/8B75yL5dVxZqBnWWQTDEdITYJQv10
/VO1hGA2SC/EYwQyb6ptGKApPszjLr/lUJVM6OyDeS1BDvwwzYtylQQP27A6Teqb
oWlvskhN1JOwGjOjGk1F1zefLlhtJfJUyYYcN/LEuWCPN/85GfdpJa49JTfWyJEH
RMXddiYv8p+zLh01GLCFOTN9INSKf95R8v1dO/ug1vqM8X1QbW4JBkSOdMg6kc1t
OLInhCJsnh0GJeqzHYL0BINFWxJzNAHXn9p3uaKjMKCP4y3KUd8s7iQ6WDLfRZ7U
4NaL4nc3qqFQMGsC2A2WhKiATsCpfrXcxImruq8x0QSGm5gdJtlBIDLohtKpydJD
woO3G35VLmtOnS1Qhxt/dRMhzFZzKJe83VtmFEpYl9UXs2t0BukxEn94YaH0751x
n247BHKWNd0s1cZGJYE5PBmgeHA3OavdliDrXaeoEybeqlSnMF5RH7+4bnyks3Fx
SeEA0C2L6sZZtYbbINYWr7GV/SKSuMo2UT6YIqktl1J6BbLX+RWXvXRldUT3ctgY
XQmmC5wx2meXGX9fy303XNVThUqauP6+fH8fBj/pLc+HEcnUv7c/kr0683upSB2e
R34OytolzhbOq6TSyA9R6wkQe6zIe3yNSWqD8C4MHl7iaU7E6upew+lwWmG7pwQw
/fXdAMZdxzjNgt7MlrNHBhCnMmMoQkd0oehrC4vvNHhEznCWGO2OY+bf+eb6ljR7
x0hk+RXfTx8ce1yarOr/wmbYydh6B1fGaV96Jw4hx141FoPXFaT3C+BEo91h1OcQ
ONmnjjxnkiCioFYe6OKa/c/0fjBAi4A9oYj0/dFhyURyLrb6nn4Jd+aMsm0TgnyD
/no7YvKeIOBApapg4R3MbYZneaa5WpzsqGPPjrr0QPIjx8En2ThzebXEx65avPAw
mf5x39PTKWsGke5FElKR7oxf1AXlMmCDNFaAN6euktQ82u6TRwDxMHuvah+LGFIG
TeuXau6C3ehqNOdWGJtM6Yya5ibiXrJbhvdDbzQBxwyFw9lrdJMIWUnV0+E3bStL
Tiak1JU3ryqbtCJZhKIkrPeDb0Bdc2WHKKkMCasZJ0arqvdWIMV4M2wC1JMTUSR8
0VnydoH7xd6kWwctjnzuq4HYm9aaNGSuPyzDEBb1+BYT3v74PEGP7fDE05Fb8IH7
torthkFcMeYO1JE6tk+qbuGSWkcKSBBMCaf+8SvN107ptzZsq4UnXqsSWmRa3nn6
wbepHbs9RhTI8NR2+8jwyY9uOq7RW98WF0gBTHUIMfbxHLjCBAAlaCiBj2Zzgh1w
+li8FMUe/ZXchcDZZDR+NasAgr79rqvBLrFjfuJHtcw=
`protect END_PROTECTED
