`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eYiJF11liRHBeq+XH/zSPUCemUjlAqL5rMRqV49U1aibkVtmb3V802wEVBZLv2CM
7mT0YqyE9cEKtEYoZ39gyixb8lLcnNWOpdUnnM2zJgJ7xVe6V3Fbj1lSlbzpX2cG
z+jPBbFWo38+gpQF0iyxEFEOJEVw15xlHc8u4fk8qcp76nnZIjUQsCatSJ16oz/n
6ZInW3CM97xEYLyur01Lr6FSH+UUZAKlAA4CDTj9tLFoLzxlMwWdv/DTvTB7Dhnm
P2z9oGxeNbdItWf3AL9EIa9ovXfXKg4r+Ewep9FTSHPB/N9eOJt706YB83SjlrJ8
PVG432S9hYOax7YL1bVx1UJg17AhUjplIyQATeFd14akxKbh6+aVdgEbjKMYIujB
f/8Y+ADRYP4Xljblp9wDqTf2J9iMDnuqUybPuPKJfoJLjreGVmjPAafCLLzSSI1q
vsgNI3qvN3f/fAvOERcJeJlLDyt6MaqdcQEhY6LlZa0aW12yAq0NG7prbPxtnhp0
datWHYjZo4FOIML2q6nOKAQBoifeYteg94firPr2OS5iWQPLCepRTIXs7j1Y3N89
slk+RqFOtwtnq9C8VGXEW87IoxelKTae0A73OHE9OVulT2uRXZeu2paiKBrY7XGO
RrTeDIbsSJ23Q2oVSClxVhkbJQVi0rxiRzmekwQBFKvN0L9hWIpWJtMer0K7pneR
88qp02hz5XYgCLq34/5QLg2oIu0ysKWzlUdC2Vg6YyevU2ar1DfuDnTSsr0p7yZ4
s5Wl4xsB034ccIswjVBkzvSgytHsClCWX8ChOSlWteUvQHfpL8ODlFH5BktTVXhp
YvbMW8SQUe4e26OPUzATTkuk247zE0BApTtaA2M5U4KKAyQ63HX5skzjOYDZCStb
061pScEvdK6kFSDscjNSmxB1svoo8jV6rl7OkQx2sFIdiN94LQjxmQNx3xXZcsFC
gXQVc474nv9ckYRdvg3sM5BLDMc0/lD+ZZMfKlV3Fl5dPihtLWyINeKWZSlS9yoI
bCWO3AfsVzl0x0WKImr94ul9xDefDGTkpSyFgZNNwje2I4XuIPCsXFLXnQkdMmbU
QgLEcPOeLXSIOWdVfcNMs5NXhGqytGAh5WznL/ZcgHehgWERugcWmn7nuxrUtOde
3V1tse98zEClNf6CM2XuS0qx1h6TgKQBOTGh4mRC4APp5WWXdowutCWtmz/DaYnS
w0AAPvU6XbZ5I9YDupmDfdJTGz1ccsvtUA4bZNT5WWN3vEL6Sa6spnjWO2roSgaX
y3W0toxRAAXWjFHB8YJCRqkMRy6ooyDlMvCOtPKKxDSwElUVjZkLm+cyXeITAE1b
yELHONyAtxe9nnsAV/a4pw==
`protect END_PROTECTED
