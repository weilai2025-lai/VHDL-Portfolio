`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
muiBRatIudmyEgrzCZ50dITOit9sOhAQHV81aMQbty494gBOVajObusRhpHgHDlB
FDlADy6zQUa6nZThquUijz/nXB3TqWUItlaYOtW3rjZTpNiPBMnc8cP1JUh1eW0k
iuS1nXyGlQeKnXfj2wunnM0ViDxq1izSCzGcQto07L8xtHBAS92tIUA5WTGkHHj5
xaG6hGtc6VIabxPf+qDRVSRpWhEdF8wDP4noQdyzCvz4lqflM17zTgAslebbZ76z
941aLiVWh4bLKeGV3zaeIahBUuq0EbPKPewh+Pj5MM8M8ieLHYrIjqnWC4JfvxLK
mngDaedxRbY92+iqf/qmCYDduR7ISvtJesEIqoWePenPA/oH1fgmoukBtAC4ANmv
bkeYNz0erXYstePnOUWP9SgEi2k+lb6QcSAK8h1Bd1c1isSXLUiTv0UIJ8eivhae
rwg4OqlWjeOakv3j9wfBkgg4e76IDHKmWEzy2+32oooJIEoKui3uK1EIwDppDwts
CjWFXKkz6EnSxx74vGXjmFjGGqUWQ2vwMobGWDPuBcIefLCtWEKBM9MLWEPxb+TF
ObyPRq40wFHFN6I2hlbUK0CHnc4ztvBJ2XSgLWReOOHTeRKptdrLA/S5lR8F0NqO
N8KT9NQVEDU2yaok5lTfB6nYulWsAlfTEQp9NR5Sb7FChX90Bfv9/qeimrO+7VsI
pZF41wQUDQK9gkz/yYI4A+5NJNd/C4MwOipL+RPWrwlqykXZrD/HUlXbYR5ezghc
xlXcZF8dlBEkweRgg5LPFuNrmKCr1o2MVlRDfN8BJ/1FY18HpxbLfr9a1A0abrXr
QDafwDeFIyljR8Jtd5mfiyqRKH458gsFWY/z6WlZuWkVW7v1qb6dmVLUDulM7lop
VU8e10tqqwfcItVR7yP3mwxzonauJaKy/jgInM5nMYP4rz3QLESX8qLmFWpJ4f55
uqwRzgEJPjU/5HzSsn6nL9phDFWjvf4j7RbpEKJGFLTpRdjT54C7ved0Qr6zS/iF
0I/eVCSFm4J6lyVGoS+4ETeq9tSKe4yqBS2wm7sXiiMNFSxFvoaacyjjOYoW/lyV
f4uQdhc53a1m/HxHnK54c3FIENrwmYcCqHqtpitge08LWN5LR50iFKaifE9s2Iar
McjwrIRMz4jVprlQAlU4B9HuCYBwc1DKINhAM+803Pw0+YBAhdiERVeEP7I9aJ9W
i3XokvYQJvwnEqZ/FIm+qVx/gRXqS5JJW56NkHMWm49UjdbL6DlyOru+vkVpsCWG
AfgSlXJzhs9vUdEdUcIHYf4x3Msa32jUxLwxN/DiupTPjqvMBqxTtuEeXoasNyBL
X+fSHhf0wsiRFzrCBP4p5P8DqS3UfBauxgbuGZ0TE6JIYZNXTqQVzNMBxQpUDRqK
fE3oo/OgwmXehgWFhKYZIH9zIgrgJ4P6gXikf5Y9MufB6mnnA0vEStkQQluzjuEd
r3nQRrdiz0hJ3u6E6Qr1dxU3nIX4frRmNwjFOoapY4W1jWz0rpO65zbDHgssR7C2
bdrUBQRjw7zpMo/crwky6YCzrCv9AXB5SedMl0Aw87s2bwc4y9e/bS8hK+S4CAmX
uHzWSQuSnSTPMxLgAxZ0EB5BcH/LO7xAVsda9bqX9s6VFZfPW9FFhZFy3PPdTZKE
F1M//b32t/1CiMIOXzSZLUvD7pAz9EySf1NY1EVNJ8s89Yq+wkcWOMygcVVbBtup
6B6qGc8VJuYb5xsSTOUS0sGXKvI5zTBFWDX1tXdr9lkADh9kE10Adzo9jd67Q8vs
yZVAFmKlGX3qQYF6VsoUUkpVx2/6WjX7uUXnZofDocMhCrEhRuZZo98zkuVFCo6y
hUeRHkYiEomh9emQeb5lTichEUeA0foGVqAtRIZyqi6yoUnVHGb6P0nDC79ub1uK
C3fEEeqEhQpnAvxRXYrPb0Zji3D/CbRph8LKgCB2iXiKaEdTA3RNTQ7yLXm7JcKy
ZZTetEOH/+2q0XxgKFJFZIddx60cJLQ4pQKXfKPetm9QTXwGwnzh3awE8o4jKHTz
jwY3E2R49KPYO29JA0cMOoSL8uCBG8Yb+zIg8OM+vplbmrCvgCKQkVosHTi5f1Eb
hIdL8VJAG+AzlzkvKhRBDAbLs9PuB6p6ZOJj1sWujkfcuaMTZ3ZQMsJnxFWHRpBd
ccYXk+4iYO4+UF+wKVH8nWwmCunQD9lsvBZ3Q1/yi7V6KwMRhbdYwgWjEiv9yPpW
SZK5Ozmr1xRlUm7Txlp/wXZFscT9yDaFjMiKDB84TjdMMkB9yQvW0olQMUY1CyWS
gBGSuVONqEiMUh1BfL0BLM9TOQt9gRE7Xg96x4uefBfdXS4ANqqbEfobJNFq+V7D
johpVR/3RBDRD+SWCw7Bx8J/+FKLOlOPjpLjc18MvVHFiQV2GZhc55EEBBWmGks4
mX5GIBCf9wESBmkYkknp9UqjiopumXKsfehAWHJsINdJyM2thXyyxi7JWqYc3XT0
69GLuedXQUm2/alefD0Fy5bUciAmHAgqgh/v5X3NZfZMRxEIH/MTs978iOibdFT1
I+R6SO5wp10y/laWMp16Bv6CucUGwvLbFmE3u1Fo3DmO0R6zq24yHO7qHquEjrvQ
WaHUzj3IbPWiG4yQu5+hki66bBVhOHs2mDayikjUXHCPFae6Aie8ltpLTbZitdRP
TV7vv8bHTj9eJ0fMx5BX5zsRz70lQ4P57LMRx73t37p73Z+In1o8WKB6d1/Lyh9O
FIn5NEbVSeMiLzFgi2GM0UDdVe3Hys3QGLxWZccIEA+YqSEJ4w49ZN37B8VmJAOR
hn7/+nStN/9wc6ZXMwdHQPQeOhTmHk4d2KJykvLlur+ys7rPQZMT+gGuinBweuPg
wQW//a+j4Z+oJBDmX3EwyWhS4ixuTOQ/TzhQRhdhG5qV3T9o47BAMFJY0CHqiAZ4
2OhbEXzX+3bNFKv7N7iFWUtcTc0pyNQibPK6pfzMW7Wuox95sb1KYF9YxNQ2My5M
K7Ra+PdVu2SKMjBjyc9lDuFaVBXryTOXFeu4cVI2gHQR22YMsY+khtYn+lEHgsIv
bML2M6oe3XYXDgjMZrfNZnbVulzVor/vFG8LRyxo7Tvm4ubJ214PdteCgT4uca/x
L5fLlcEOUzB+CYf7tjMHvSJ5t2HGwwV7Lg+hHOa9mOb/HY1ET+PLEdg8a2SO7+GH
BrnZ8BInTcWMlP8tCnIFP1kA9TtV9vAY3PfB5kZZ+FZw6d50KkDRbA1HOI0cizxr
5ukqTXW439UbY5wFmldl4royMUwEbhNUiQjkTFTu7vfN1ui+nr3be/GC1oEHw1nH
i8uTJZ/l9ty/w5Bp/by+0gDbQ+QMWIDusn3xXQf4VNKZr92ZKLMwcaOFkRbBcIzF
HfdXIWwPSjqhZHxZNjiUX8kkTJ5zbg/68bU+BseRaTuDKcLWtvmz+cw4uJOoVK/6
TN/rPYGpgKF8eXmU1tIVB0YkL0yPm3Ih52LdXiu+zYJcXXaOEoo7/lzSgnTvc9QR
7d4pY+84s24oABl4ovDZnfNcJh0okdlD0mMP+h6wEYlNzT1xqJNPc7BNxtt+A70E
JqPvcHCAbOxqr0HESbEKaYJCpDmnifd7vWhI1BH9fKgRJK8sLkuOYQ8/Kyc0LKBg
ZsSPP+uGBpsTtDd55IpcGw==
`protect END_PROTECTED
