`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrLjJBhth4MKomaTGH87v/b+Qr1IoI9bMoSRM4oYaMK4Cpshik2IDyl8+EDvl5v/
ZMwzrnRRy/Z3RYh0Yp0rCScoLXMnzVhh3J9mL6bH2tqN1uQG7h2mCAJu3SfXscF/
pXy8rcbtzYyGlebTUWS+MhF81S3BX8hKK1gRZAy/xzs6j4ccGpP43lHYRb00B0HG
VDDqhE5a589Wp2ICTbKxKheyZ9YiZZwfaVrXuDTM3QLgbDmj0qgRwUXbogUd+eVm
/v/QRETB9fNfQ+q1IY1QPu8n4UhTcuC2cpdvF8KvrWnrk9J6tN4UvjFbs9q68N7z
CJpnmCn7B5BB66JDVy8bBuWMGgSQ2V6Ba/QlpUyUC7+Z5225ZPtz5BuDDSooNHUy
McZz/zV8DIfFm5cu6Tra2sVyQnMFWFxqnJ1ODvhzbi/gU5weSGpO/5vV9nSjmSgy
CYSM2r6TjpH/TEUyvFPin1OVLtCWk7PyAMALPwrRUTY26DmKvwMnnmbaOkFd5wbR
n7xru36Qm6LGR44y0VEDk+e7TiquVJPuoUSdW6BL+Zi+/V1mIQuMLmVqefYXIo2+
XhyfKaFKN/UjUMkc6ZtDKtlvwXNAE4Sr7xy/RediaPQrFP5W+wlXxM1WcjAgbkvJ
NzYndNurbd0CHVqdQpztkHIl6vmYMoW+V4U08LdeLU1jjTiW95inlt7Hr82sBrwl
9LewDPJZCKoYzaWcYWgGTa227KYc6Q1D98bVYO4q25mqv3FStw7GEREmB1M7pR1H
k1A9tHD6/OFIJv8MNvbzMoXviwZ1T9yG8j/gRv218Ntyv1ecdK1PM8JCLwZNN4+L
hup8OpeF5SQvP/ehMnrmrPIQ7hwci0IFKhBxoatq7fXxD+N9ozSZqCfPPmyC2MCz
lJ9nspFbfWMV19k3HAY2nyMLmoJPGYJQPoKV5crFZF6RY2CdHny0cccTREHuXmWP
ZUNPSag3UscYXPMWWzrdKBI6zF71Ri39q0cS+hzKsrtA1GNZnT1HVp+RHgpwMF+b
yrIOVRKSpS5fkoePw3+2lfZ03k3XyMEE3EJOwcUQgU/hayNcU7sOXvyV7Y+43F0N
cnfNrRk1OGzO+V9W/u3ecIE24Hskl57AkkTpV71d2c+7kS//yMf8XrpR1P9hZeM8
Fj4qFuBh453B4WgLRpWTg1aGe6Apz+OFF09bMYs1JebOdHX3qLeqJ+8HAajZd8iG
xVuZmgzQXKtc4qW0OnPAwraS0rsgz+M4Bwc9YeKCi4Q9Kjx74CddSmgxiMaLXRy9
/pWcEnrdHDVZliW6XsBXaE/OZ7pXzqmr/RlotW90iSgn/OvvxfG6ha6z1NAJWXWl
/2qH4/kJ2ACQUf2iWMMcTx1wChhnUtOZsyqEliNMVUuquZHmEeKIT2mH81qtuWOe
2YFEK+9DZU+WP98WjFgSpaU1GDlQ26DvOS2/3OYkII9Ygbo3MY1a/wextQN/1ATQ
ZT4H4k8uuDHuk9vy4fOfXS4QzAlPOkOHWgfWeuNn0V+WHh7tttugCvFvd+FYCYBE
138gKPJZ2+WZHM+BUubRBLRmB6bVEfD0uorjM6u5sLaNpwCTQjHof9xSRZp3Apr+
ffZAd49J+L3ssQRgRq7Uf3nfnkkVQTmev4tsNH8jCbGRuQkIuxwlSphmT8lQroxC
6wE5fzPzpwyQNFiyFeViN8o8a82nCWA2QcvCLcIHffspXKpS/BYhXErWsVGs5TY7
1IXXSJyPVcft2rV/LCvv/gJxOgkAsNghwPmTROOjf2vSXGjMieePXw7WFbJZd65u
7hbjtegX8gvxqi5YVidWDjzGDy0bveoyrX1MQyaZu03u5DyhT1Se8livedA1G+gd
1OkV+1otxXC+xysHrMyHPKt8gNyKMUh5PKKjuq4w2PEbYAFMpiWKAX1Hx9U9yKp0
/6QvgWma2BiWxhH2kSkB0yzJy5QlCwfSLbj8+IkYrx03pQJ/IMQpGMCzyisKsHBC
gRZtJnvi3WCD7/WMuZJCmMvEUXco31iodYPlAmLcpDMnUXWN2Uob+LMVJNRIk0mn
jWBgmLzK8DnPOUpPQRlpMKYj51lZ9z+Jnxyib9WtXDhW+yu+bKaGagKAuboLAeLG
3OUbv0PrzPopXJoK50MmWogl3/IIQCxyFAOzLsASrFQnjflBE5GBGWgb1i9Hhi2m
TH7FVtZZUYJ8CfDhYqW4REYkfy9C7a8tKeH/WIs9PqsLX7Hz+Lg8ds//8xsO5n8E
PHD4+v3fYD+lOFNXMJCVqHlXfIUFY2UQdhh0j3Q/Ip1lU3q1gcBCka52m4E+Uc35
cyKJqb0xm4zmsAFne6hXb0ZR9rBATuycCqfzG78/ryi5snSCKTdgY4KIp9JVQf1r
1Wj4FyzHgk0c90nPuVqqhr3mo9RGuCX6paKzCcC3rtOo40kPl/+bdLwAxh0DGqlU
hvwqB1yrNYRhbGabefM7CduRRagQTYzvFyuuiXmCyaNs9gT/ZcJPg/4qC9kt8HPM
Fy3+D8aL+wDjmPMTHwhKJ+BlJ95kc6FK4G1BbbhdQMJc854SfsoQIWudLpvTMUSI
CuWALKluM6VIxu4nbwuTSQTfgg6miFKhi2Cd+gnU8zK2HOxV5Ild+24fYSy0roqP
+trl/7w1rWSxl0TnSxNiwsOKKFSx8g3kH+kiCYkz5f5+mVu8yh/irhXEyNusx1kP
tfE8nE2fP5SMfIE4UNINZVEz/Se9AY9UiPUUSvxy7NqF6SKl/bc9ALNSX8ZqUm84
ehVpnhlRcw9wgziczG501/9+o6/DviCEBqBFHHxPN5rrmggVAWoXgiNXbPHUexlE
HaGrNhkb67PAnU9R4UmXPwkI6oNZVjvM1rr2QfSD2oxPkjbA9oCF0KV9nsSDi6s7
JQX9dNrrFYv9oKwEXggNlx6r0wuICqXeGQKoTbmGBw2pKlOQ99WeaRaOz2Jg/ueR
J5FCeuArAryutPkxQ07WDobbrcZWtyvhYt3LCAsjNFiR2eJ56wEgnqK/ZpsMeU0a
yoxFfVby2ZE6LerKvwv4avoX2/Y5Dm2820jL3j3ZAj46wvHcAfC5b2WhZzAP0lPa
MRtF7gzkoMp+g5X5hKrzPyovBTXRiUsLvT+m5tdFkZZtRzINux7JWL273Qsko+Kk
21jEpicwDbQ0+VfwKtdptH8qtGXkmqZa0GVM6DQwy9GjVggE6dTvAfvNk6aIWRGJ
gMfDAy5WSWajYtBVE2ALCRVjNUa45HCMZaz0LyPJvKADenzF76D7zEcPmtAqcgDF
F1BnGMvDiDD11LPEipUSewiFo3YliKU73krouA9ccD8D6FDvcq/QBKlDDeXPqHfk
/IjlgW1uST6LtvgzGSkUzM+HOAgVeNG/8+7SIPKH71GafChFU2x1xkEJAsmUh9yw
Vk+UWXtJlFTAPMxTTIs6AoHkUprDRwv7pqe8lARGTpsyHiVcds6FSczHwr39RvCK
DTStZ8SBPSUeotSlEmS/1yHRXKF8/Fz3VOTX3JJX/TLaif0ZDRF9sZpCrR3WbWXq
fV/lE3PurkzvJtGIu0aYqBRidIJj8sYxj7emV8XRoy/OpptnZyq11B3Wn7qHXEBd
o1dzr0rre/JhzvkbdWTlEnmDHN5McSdb+vs4ZL5c3j3ksFF/dzo4bSYW4uf+So+B
qeafx7nCqsvq6BnHybhw29rtp574fed594lN7fYOlXQHvWtg5iJfxOTQwdu+xnc9
Pykc+IobDPX1KHQxlsNjuQ20Fvy+pBqmTmqNm8g+BJcXvFyd3tG5+QjgAYLSagPq
vYd7NfJTcxtzShPfo8ZYyEa57OxW+t2z97+NBmvRr9EmtGcv1fz+a5j6UAD3ZkJG
og8mdATl08OHQFQqEK3sz4uZmTusyK+hZQ7GMa/WqYxdlGkJFPblazu+jpxw3tAY
2aZabLc+7yIjZ6vXQIDvfjSBCzvU7qqDFMQ8EUdZ7VtbPRKg059GdWVwUpVcnZPQ
rBXTUU2y1X8rK07xAwZ2qQ1pC5IGQNErQ9O2s48Ppv8lKaGMhFX6L7Zc+RDSmymo
I671NlYmgyAwgr6yyzQ9h/JvT+1UndxjEQdWSOgzxIvHuGO3JmzTOJRt3Pf1rIqp
LZb0ZVyKFCJ0e9xLaW76cMPqkZtyU2HpyqafPUSR5S/xsFJwFmyhxuuLBTOoxYbQ
xWx4LINrYHoIY0UwulhgdhYny7VWf3KqwGSFQujbH2uDrgvME6jZdgC0j75E4e7c
ba5T5/dXJ1lv2znJbuODBlIpfmbAjz0l6uDk1XicJqn4/RpUT1JN3K3J9xLX6jAt
o4PSzFsM/M+UseTBqO6jm2j+TAvrWTOZMJdd4SHuECijakEytbKCq8BhZ7vMPJLZ
OtfOXCN/t7yfKGCMZTDJMTwIlEZS6k61FZN/+K/dDibD1nw4EP3zot9n9cl5wP5o
W+kF6fy66crOcZRGxmT/UPbAe3K22C1NszxarabXeS559HNZx17gF7B1mgRfV56g
WOOgHn4+H9ybCmBMj/h8i73tFRA9SzNyWd5nFpAhnP/TfDNJ6egDT/4EKo4CuNSC
cH90L6WTTZSC+Nm45e/HZiyeyEivtzKTsJrZaCw3GWrzViq32p+PwCHbhDerr6l/
ELv2OsXByEi2b1eRVD2QGsajjXw0SS35sUF4Knv3ZhZ06zic82d6V0MJMkzkcal2
Lv1kVTSoXEH4oxyf+kSCg2zZK0pgcDlP5VH3AZrUvkJZ3wixhk9X4zj6mUR8UWSx
NmxPkMazG5eS0NjbS3DqUQX2lwS2HM1/T2BfrDBA84zeNQRGFomIPKnRNnPTlRM3
ZP0hoPzOyV3WNwPiyCeBaSMJ8Eubs7+Cbp+LaI6wCbCJxF775ybBU8u47mJfYAmz
xdpvqm4Jk18tnT6qKCsnNDE4sPAYNlyDaATpKIGFnhJ/T/RB2fjnTGfEoRRe/i5z
zO68B4DV9k5vzpkmWCRs+P3/iZM8OvhS4zr4l9donRqbdWUzIHGA6Ctkh/qqW8dC
+imbI69Vh9vPWCPSWqTOq4nc1WlbwuE8yGDi4NT7BuQ0tK17yV6oyRkA0Xe8RePv
EsTSw6lCWl9XwP+n55srjE1MmLwGf3P7jwevYbOTs1d1rLaskFHDOsb34y1ptJzL
2a64j8SZDB+h7JQ++tF8FYVNh+9on5vcSHti1RHMEtNTFWeHogcogMtOY+0eloJD
Hp2gMO3/WlKpX4rU38hJ1EWAFugCqZqk+CmAbMyHyKSfYCUz4ddKddIpHRpBwpaw
AdEzEPkdYAhAzE2mBgZy7q2b/c+jD2/hH6XyMo19eZl1uE+Foq66fmjkjypEP1qp
7T4Zv1OAPdFzpy3LlI9EiiZgfTvl47cEUu0v2cR5LFSZL7pThVLyWyuvc4CMJK9H
+fxhVBxHghmyCyDN1pybR8ZI19y/F5Gl7QWleKcIs8Tl/O47ABwPe5hu+wfdGgTj
u3rN4kD5NG6uTr1XkkU5/02XVnPhxXP1QuwLd3H0YcjOP/VlL5MlHB7jDeYcO8Me
41PEb9gBO2pEAzKkyzbgeFFV8YhhdnxuYjSNRejARmr/EZF9OjMKu4OCgCGnsWC3
MBWppMV4uLM58Sb98mJZML8xlGOZgGebsC79tJ4tF+XmZ8xIpW1puPzx0yH6IlAq
kXWwZ5jxsPXvj0h0YKSBG0Vf9khzk8BKcIAoaWW9UWCG3yUVfiBoYh3HLwTjzTBj
35f1f54awTGQwDmJ/d57KwlFdoVVovUk8AcKwtNrNHnhx59cY6Fj9A/d6HE6W009
RluSYkWMVRtich+0G5eGmUCBw8jibxbwvMghX97VWE1IOW5QYC4TYW8m6tJDEwuY
B8sE4vCpWO5RKaIl8CWvE19LmLjXyUb+23lQEtTc0IeQpeqCOdgunEM0WTojPTuH
qyCiHDGYF1rEJ/4hMw5CBs6OkoJmzaadcPo7wyeD3e1XaXL9p5cXyRFjeWoFwhRm
eslmPFeW5zCYIM0GZnJL3g8HiG3iGDnrB0g/MX6kau6kBKXDl3+Zf9PBy1VnmiS/
KScN11NQXXbKCbTNr3dmTxIDZ2M6BsCzffWntQO1Wmv7kqOk9Jpag2ez6/B7UOlJ
FUApQbShKOH/x3HTeppwiX6bjeR3o0chr7gBUpwk1z0ylvCRfq/E4dOkgw+CMaSZ
V9hllGExjWAc43WCh9p7ttbL3J8gANfhnnlnNKnkeLUcAIdU9pJP1ciq9UmRdEgF
VYFMBpmZxv+3llvIQGikxzQIEHmdcChLOYOT4wCWlBe4FHiQCYKvnJilyykKGVc8
41hXnewOGs7wx0AYfdoVjdGULb2B5qDToPw3MDTRJhXlG2j+VgeH509TFqZHayji
cDuBgi40aYYwC4mBOAQKGyPgO3HuKJD3TSuBXIJtFEzT6ziATz4dDseEJQwRfzGn
uLaX6tE2BcTikHGSGGDjJHdO/8h9eatIKpi+zFYDrUGaO1tYRaxcOb6J5bFloIfb
sIC0vYgjq//FHour57jFCEYV0o3e95PtVnSEvOrHiprZTXJnR0N4og8cjrGmqQP6
ta9NV8sVW5MqwdQv8owCMAJKDYX2cHYSp6VC+z+5RYacmeHnCcfqTDYSUXr3Ajde
SXubi+iMVUBj62E00qUEXNbP+pebNRa9WxNHDUCTG2PwWVlRczMFlSJg2WEpthM4
Sp4wx9iRjjIxPTqCkqRvWuwHZPvU4LF32/F4J+lP4Wu6QwRB4Y2G085z2HAAZ53B
NCUxz9RpU7JsloeZZ1WfARNIEtorfINnE25o7gnswyV4V8XUhpJUhMZYVLjIHyVq
t5kswNgijIdb0AQ3qdhdxyqw8oABy86Cc93q7yBtbWzIcoZ7VXENazFEiMDnFt6J
wGZHzmMdgkfPwA7jj5SKKfbbLXAgY8JwMXiqE0RJv6/apOV4cGNrHq7O9uh28maB
nK1ryKrM9k1IgYQdMuikRQjKEYGw71OYR5qf66Vt/CO6fuF4dZXCxifDNWJ3Kdt1
HlC4kEOB0qcrT2mje7iqEonJn3i4FlpgyvOgE7iUV4B95n7qQzEwacUz3zW1dGxS
Wu4x7KNE/kYHJSUTQAKj0QzPhaqXqvTy7Du5imf/UrPMECd7n/n5Yn8Q9ET7xAnl
VAvbZYixCzD6eqBmNCPVEw+YfT6K4P2gx8x9KQ+mS4hWebDLAWq0hJLIHwoRsC/c
RnPiDyfWbp5MLI6cWP2syPIj7aECJJn5fgE3ox9G12A2N/hgRQdo0+ntqqwLyda4
T4esEVYxYH2uSF4ssN+0t6Yd59HYaG+wptxx5Bv5ftL3LjDnfuCc/VtF5d37s6iz
PPyLwdEGOqoBGmee6yUyLDWdTd6PJ4fqvbSrba6ZAZegcrW+ywOr/6nNPEBDsxm/
SJncE0WCSQjt1u4AcG6VwG6yQCUMeDsGtZRV0C//59tHCTRmGVCH7XloqTXklCcf
ZS3oyBbhOdND4Vg2WIlqCXiKBiQZMIzz2RicS2h0qo83ud5S2tOOBb9MBgqjCyx4
x7dNQr8QvKgkOmyfLWlNjJPc8+88Kh+hdZi9p0KWmQO682rPfL08jTpounw4Akgl
PgHi1too9AVuVQ8z+2P5snxXzpjSrrPT+pB4JYDrDn8KB7/+J6huNbHJB0XGZj5X
JS3lgNS6osMcBbd0ixrG1Ijv9/JbtAnzX9QWQbtSP+X3gigO59CDd5MF5UKnr8pf
BgNQyF+QZV00SHyHsQFcpYjLFEQTdsTbYnWMQoxtbN6jFrRBr/aXEGDhH48qhFkt
tlnSLqId4PIq7AzRslnEbqHQPoKoPpCLTjw6AnTFvWrPm7nCIrNSV/qf8V2o9FgW
zLlDtqsDDl5dEL0PM5PyDz6PM6kf6r16iakzj8osMyjKANHqiFPJxZP++iWoI6m1
l8tZC/cl33faI/ym6V2MVAGLwuKfbGKXJyEE3XQOsCcEikTw+Urv2FOIGhFURUiy
qZnLlDfNWkRv+m0hQctExllbkcg5YOEV69BylC+6ebUAYk9fpEcHR3XgCeGdvKko
kO6Q2MVR0pOm+ij1dk4qoTlppPWf7iDNIRrjYRSOYeEVHXh9J1wts/ZN2FQDbl+7
eYni4QDjSK6JuwXTFAQ9hb7wlQySmmc3DGWzDi0KDA9YQmkEYFOz6gwENW7PiD8n
CV73fuqwwHrk3QX9b4sW9AnHMkOp2xpSyRQC+I50i2zxqHJBZ+TFzrHjrhtUkP7m
AX2fXJNGwp6kLJ0VMVDzV7LDvIU/EGrQttTnXqOS2J3lR30Z7FSUfzb/RVWMv/4F
STQKFXvwTsFy+IgSCJG8xoxvEn193REkDp4+12cST9h7dhKLSGNwqHw9ZSWbsei0
G/dMKEI45ncLQDzoldjBjzcZ1iDV5dL96HURw8n8F+qAwL7pnICHiBa9N6jr2g9m
t+ujK77qGu/Uz+ZcCBTCpmjvSfc7KTgX8fb5/zTQG8HuzoRNZN+fKOcZdF2KR7RS
01h0N1yE0GcYbhfI5XXXt4h+tcEKm1jTkVmKU37SW2K9wXEmBOMSw/d4q+l7iD1A
w2DkCjBuiWz20opKe9a7K9Cr8xxOvogq37uSunV8hqryEn8Yg7/IYe8gVtHbBQxx
gyAnc8aJabbBdstOEKAhmE5MVhrWqKas1Kf8HJgIqPY4O8SuoVDae9XAMDZTn9Ba
uNrcPK4zzxWtUzJOO2qtqDxCMRV1XthUswY+mUdn4mFUaTfA2zICg03/5HZGJ2i9
fOJ7xz9bwE/rj87dx6m7AprFUUilyu1FFCwqnq3F//5i68k8CFkl2+ZNSew1wGA/
Zm5vqx5vLMQ6a108rLH40ab7d0+Q7lFm9BoxIPPiOhPh7nYYo5KqrXrJqBG25PsX
9Pzr4LzrZ1L3Xehdoc0d4TRNvW4qQtHg1QbDsoqXybeZoQd3V7NUftQxe4WRFA1F
y5L7skjElzqYNI5ZygM0n3XS48bVZiqCw8xPWMIGeOr4KSfx1GlCHruA0PVshCBA
wp7+4dBvgGrN7YbzN+lEVklZKELNKb2JMhSbzNCYN5gNwioubhwZ+yq8LiFAhyWn
rrj/tcOF0fgsUWVr3OWipwx1plglNNe8JKqDGgfyK9fGaPj40e0uXqRHtVJv2awo
HW73snJjoqV6G7g+w2fQlCCLCw6jOqQ3oZDu4Kz596QGrMpx9CSgUiTXycYAZwvc
dTE/p3cGN0T3GGlwe2O5el303Apa5r9pezK6ug7+dgrEgbSmWBsjqhvgwuRMBAgs
bwkuzQ4YiemoLtBsXuu/sAiwOdL02x8L+KSCDlmYEZSkcKbpfIZ1djVZix0y6nvf
zuhs03j0DbZHRfz7tvOCSe1stCYQs2n41E2vdyyDgyxi2jBk4ka21FNrMdCJzc99
gfHQCsbthvwe4fyjv/DvlkTI7qSJfHUhr8bNtwGN5T6lppY9/tClNUJZ8OeJJfQ+
XrfOmiMytFBRc5WPkYYhnCUbtNxECZ1ZBqqtHx9tPMMTkMk5MvQVj9tDOsFH+PdL
p4I/0rc+smrJ8wQQ1n9Hvashf1bQdZp1bYlY91WyX3yOI86qKjpYwiI9KR09Zz5N
mYNw1lkKdDx4zL3OYMUNGiRX1rHMjh60nOSX9cpc3dDtamoW3yQMYBVfvzc5BNo6
7STIdIqMNnYneOYGDqzkugnl/OIXGp81/WJMukstqrR4J9aQHocjm7LHqjoD6zj3
FG3S6GPQfBCyVWe2kg53bvfNtDVKBIeS9nnx7JVnN06ZpVzdwK7q7AV0GDAGXAc0
5Biysq63aCUghQD9mtZfp0naBDvL/oEoxaKSeg95Dy/eTiQJO5uI6myAjWTsqmvp
GXGxfaYylKx5p2bCze/Ls60HfHbq40Q7WfCNeWA09cqQFy+5gI9FfZmFiYDzj03j
a0U2j7HgPKbUqBR/69425rlTrilheJLYopiGhGDON5lJJleHbE2soWKRrcSk0UVP
DZ4MsvcVMxLBXfZjoeFkqDDKN/dzr33O/f9GekGmRvV9uluDejngfXghY0/8urOw
93oeLEaNmgZ4Ox9UDnZuH0plOUwFvE66qrgXn6t+1IY8LoIGH8+seGCEvmPonN/8
XQJcuICiqqqcA9Nf3wnLgHx4cn2SuXNH6+pUnuJWavauQFpXwtKXs3sa8uEOe/Um
AhtmJjGd9A4aSiI/Cpx5LvMbHOiiqT5FnUyx9gf0tJcK4qRa1tHFwdrrc2BKc4Me
BcHFByJ8PqhPo7F2wO0tSDPU1AiFjFAG25NrcUCJssqjiMTMaXLfA0b0KAuVBgmo
OicwIeMHytrhVQ0gScO041dPWw8JYftvqnFLUZ6WoAyKNR81m5pfUIAw96ZQgAl0
fnDYrCj9sxIF0zo4/XPY1Y7bKCkGS9GqMZHCd5MIWYRC46DV/5ciuTj41TO9Vd5Y
azT5qcK7urXhDIQZOmhYsbm8mxBaxETwwPuBCjBT4WkcNTFFkipWXTaJp2VT7dTs
UG0lsW7RKcaNESURZz2uwGJawO1d5h5HwJHeidW7X5wORKOMjoQOgcZByiOR0hr4
0CjmwTuvSWf8gX7M0276BJbFRq2DjWWNnAZ+l966xAsZ11jqgdO5R/gHHYJhOvIe
IkfDgSCRDC18Z+abvMRHcF5NbG9ZyBw7174L4BgbQHrn8Bw7bB5wyshrPuRmEJSK
CrXLVQhgY+P+QKG+UqD8feC/pFdCfi9wa3ec09c/tuEeeWmwW/Xine0vVqWgdpUW
bhEDMyw2oUJ8KZn3328IAi2iVb2znSaJQMja0UevLQ8lVqvj8H4eVjSzc/qAmfaQ
4CmMAQn2sRzmSWMhq9G7xgRPMQ4+MJv00i5/ogbcOnbU+bnX4TF+fbkJxcMUJxda
/I81n/l7fntaQyq2hlnXWRltrwbkPlbJE+5IQhdLdL4v4aDH72NIWq0zcHZyaJV1
Oi0DkvciWGyuPxeXJamZI5pp/LNlNzggYOAtmwm6t7M=
`protect END_PROTECTED
