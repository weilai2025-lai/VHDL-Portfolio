`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xdn7WfJk7j1mvqjvD5uyJ0xUgm7LC7l8s1aC0xw+SzslU3m9LwBvuX7PqZ8F5gPD
6MYIqsVhDevskOkiw8Cx6EsUAfx0SW/0EwBPwRHwnKy1/TBlJUb+xYXnWMFMNM6G
GIwkjsX/722qm9C964th1TJ0YiqKGn1MWA4nctQ0Ea4Kfqwi5M6Yg7ks2cSA4MwZ
`protect END_PROTECTED
