`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pwok9nOH1/AxuhE/B4L4OJk66VXJ+J3CGZ6PFvN6bHbc4/nWr/2GzvE16qVnOEzG
z+nyyhkgkyV0lyazQFJlitCgz7EWwIun3f4hTLEzZM77Kz8DMF3dx6Jksu4QcevW
kRRYypvrR2o5IjdYopO29Vpl6LjK2VFNaflvxK8jEFFTDQtENHQ1rWqGsYklAKD9
RIigaNMm+lnKiwVB9T4uY0PlcbTz/rVMs1mePqIV1YzhfwTpu2ReiyGBiGa//7I2
R5HONw3evYtMyvXFzsoRMXUvkPcY3fIwosWxO/4SGCirPn1yK47mbXeEUTiAG5GC
6Zmv36GqCwKfhw6G1744ozuWyMeaZ04EEWr3B0Sut0p18swaKPEiI9hM9ty4C53G
Hrg7KCSlYxdvw/U41FmCsQfW141H/48QfDKL8jwQUuj4DGM7W1f6m7tYverZnqhi
f+03/iL2qBUfBgjD0owGop6/67ncBe+vSushhOIDdxvAA47Fwmzt3gCGbEXPwT5X
BUzwhJPLxPJQzg/DAn7h1+5rSIrTR8snZCy+tOYJVxOBG5kC7vEKj4Qm3xGRiAEw
CPD4sKiu3VBeRGPr5TPDdIi/LOSZk0ZfzqViPaz2hDww1+j44anm1dyDe+JcH4ty
pAfDC89bI6beifsxHGlZHXE/26+KOMP3a7A0q3hEPX9pfOPClsZHxn+cmTyLFBS5
56Q+BQaJLMa02nX79wjCKDE5/1r4r3Ft+qJ511w7dnM3TV3o7fj0Ze8fXASRRrPF
uKys+zkPZhwOAGhbq6kmumODNWFN+GBE01eK5XdqGMG922cBS3JLaN0qW4vD6cOa
JnPUvJ51C/ooc75NVvjh7t+72D6PYTBySBEmv2v2AwTWaYRZBKKvWzZHYYUI5oTL
awwY2Lja5uVF5DnIukhlV8YcoR97OJ2766j4iZWWZjXtX7Ks9IBoyIOVACEtRtc+
E6GQ9zqCBI+j+XSPduZxkMqILxNSJ7td2jYbgALWLIBY7HGhfp5WYVjLmj0EXz9k
wMQj+HvpNfdjhStL/L5yoAPzmusjNyJulvRsjP5c9adtwFaVEsPQ/yK3c2cEbULE
ZdnDivEMjtZgTSxl+i7rZ79ZGCRTGopz2l93DcFuQUpwQr+hwGP/LgKjkLtODX2Z
vGs+dDgRy7IMxLCOEK5Rp5ZzlP3imQsM9xVSIjbXNRO7qLynKCkQFQGHrVDgRCGk
IRfGIkxUHl8XSVHdqHG9kUE84PNnzhoHQBcLEAT5YDUkb/7ef1qB1Tupwr+obo6t
NPXVBqIGa/Y2i62iP8nNwBV3MRXIB00xPrypg4tLGtqphqIqKq3FWPfJIZ43wI7y
HpBgHzzpyy41gRaC0/He2h8lxom79WWJDqAuxwgjf7bzv+ggBC8oPy4+CbdXCKop
ee67SQivc7oLb6SBE1ODy8I1Rv7Y6fDWneiGHvm+0UKpA3QRz6KRXNDmmREV8aTz
kCWDyJcSNAtHL+QlfKmB2PGmHwiXOEcP36JMNMa+wLj7hWLylkllXbw9V/hfx/a9
LhAETyYjGaBUkoecEKDCKhaBsH/Eo/gHiidaF12NEzQqg9b/2UTL+FutkFHW96Rv
OF6yLmXnmLV1mVt2+0tYRwznp4sYVeJwWC4ziYLP3c7+Ujd7P9pcbx9q4laY3Rac
MF4+VBKuGAlCO8MkIe3fQHZigTRkMTLR5KrtVZUlyR6zANkdydWhFgRPuaNihJlW
85GZoJ0mGdGbQqr81xcKEFGWRtjKUSem48x29tn6c5OpbOT6gCXteUNMUJLzVBBt
RjJSl8JiKoW7H+adM/gA/hwF2s/ksiJ60qzYA2SGX5MsChsZ87Xf9nQC7xbGZxY2
7rPkClLWiUU7Jm+5OMkg2UYwIundHKJiIsueajksrq3gjTjcS4JonHUmjDzG+Awj
DzDHl+raCdRWnN0cS/oHbdV2jaE7zmuwG+y5Ex08hvFs5ONPRBaRgyWLTi+hXTRV
GJTCfc/oBU9I8TkTDkJQ/n8tsP/O/OOB1IrPrIlHjki676MbMd40sLReS/6OcHzi
t73uRr0rKjPwchE1CYqwY4c2xq01qFzNMdLUNsKz8A9SByYN0wGfyahJ8tHrV2dh
EKI6AL05+utsCWhj0J4lrBBjAFUO2DOC5qivCxE8DnpbmKRvGsc89ziXkvOlxcK7
tqJEs4EKq+YOYTL/6LUyg1tbNwjc4BFoGSXDC2vR8ks0DgMLYzrT83ozNKLpz7YH
Y6DLbb8ZlEO2NBTFerJhJhYvPgYFqbtKErcfNgs0yGN60S56q9NTF7lEobTv3o+1
zt0QBm7nnLqzmJVLFDa7yHIcArDN48OHqQdteTkk1Al2wD05YWLPEKqvqvCGCRim
rg5iUpGUCca4LuvjgDMR5vWMHbUY/hflmV/RkWNYYquabb+quyPRZw2RIAYRyUNr
M4vvcRAkLgsNJxRkgNqHaxCRygoZoLQWkPrDICpcPmkzXiS5ymkm0oe2icNh81+j
sZR2CFZsCQNumI23JadJiA4OW7XsudxxDDw5qD8SNCc=
`protect END_PROTECTED
