`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZQHZMnlV3eip9JZirRWclGgE+rRoAyqZh5CsDsU9XdOv6KR1df0Z5iruxpZ/1dE
DGk3HERq/DwB8iMqAURV9fQyranATnsbPY4OjMYBRzV0BeAPwDY1dftgbHL2EM71
Jpw8F6WWDwVUm+mQRZF327yf5BqB/EBhfMbut8SOSynbPes0OPU7CojDRBrz1OzN
MjVYP4E/XsF7wS1B5+2VtPxV80+BM2AdWXLzQcI/uhQDzPEkOL2ja/70iTmqyReT
x5Z2T/PeUuAx+Toqddk9C76J+tL7W5x9m0Ydqf3poQUbFXPYydO9xyXOlJxM3m2Y
+6YhO7WrE+RBrNRnoONwGFjX0oT+O+Bw2ESTCkYxSlzR8O/F2PvLptNG7+JpoWQ+
wMGUv6wFBQewLowCoaYM3x8rgD8Fx2wgOS4HV/XVGgk1XzrnLky2tD01EUsTx3Di
5b5SVIJRxmyQ4Xc7gY/BLfFmspScZS80Q/wIuppUlwYzFjO3PN3h1gtJmY98qoup
di2iGpG2ckWi84kGh+zfPKhvcHFlfHjMpvh44ub3/WUL4sJaGKu/jFjM1/YYUCO9
ccijm0Xa/6v/YRWUBYE/rmm3iHZQzlviZdz8gLI6MZ9S/Ed59uPBOqL5mUX3N3bH
GqQ7JWQpgcoFaALpismIBig55nT2F8WXJxv5UCDNynP1Cpxe6dqySVWSZz7OcZ62
FTMA+R6Gfg7QfedWQ27fcgFEE9oEm8TGqPbkMraTDup0ZXWaNykV6v5eqBPtrrq/
yRbXv25s3AqOF1MjIKLFbzuXOpl6RTNTLsBkXkuGjO2IFVe3JAbeN1wJjcrQQeb+
8bPyXCr3fHPAAVeBk3nhPhJt7R9a3s9I9TmDOVVUyr/KVMBu2BET/7k9/dh1ABQS
zCWa4qVa/QccMlRNONT6wG1OAqraWnkOKpuNFSChjvWuAf5xnYiCrJ+x21n1tC7S
wx1sxihePc+W0FMa53KV+0J6xmVU3uoj9U1HrPfYNryHfrUEBNAsF67IRQKgIHyG
aC2NW9AILB0Uc9aQQqR2XNhh7wNuW/BNyR7918g0JIIBSWAy0hqmkz6YczyBnYDv
ONmdDb2NILwaB6hW6jWEhG9t5UIgddwGD0JRbRleUfn2UZDFlUiYU+BukuAiElb3
3ajETT1pY66KxZXcL6vRDKkuaRhC+lnttz2z+fN8bRIUmA3jgQyKxpcec1/EIYHV
N3zY6EifFpLmnHvQUjoxebwhVp/DxtI3wenh+5FxhFnP494dtEgwOozr/u55pb4X
VxYgF0JCb1Q+0CkH8TFTp3BsiuBJr4SnMln6PYKEoSbpTh5LuifM59RroQbSCweI
clxfotJF0Ap0BpFz0OC500cAWbX3fWwKdaBw7AjoqaG0+O1cGq0SnQ91UVdSB02w
Ew8z5OkHTo9RU6xw5pDsxbm9uJW9tCPDUcbS3eXti0hj1hkma/NCouZm4abyjzaz
lHGC54cd5rnoKY3LNOjW3K6G5+SPej+5vw500aE8kPjxgmMtFog2n7utjIn1zoCf
piQALWBYJ0UA4W5JaZCGo1lbAVb91xDqW9ar1ZC6qnQNimpN9NNGUtNIiu41Vsa/
YcN4FcyUejRHpZ4goOY5rgUxfZiPiPQiZg+rUaeQ8TKn2ywwMV3U9vhnMbUiKXfv
PjC+Ngk3xjIMZOscEXDGFT5IT3OSYrTu0/yUO73/LI1PMI0EE2nlB2lj9FLFyOtg
zv7kaotArt09wclaBYWiwH2Qgf27QUau+6nCvgox76O9sasPs8aNQLdPLvEVsPfl
Rnv4h6B4QXy1BIqzRydXp7f202P0l7KXShjygFZTP6h8rWAayKEWZ4/7dO1XYKf9
KL8l5b7AEnluvblreVjcLpDllBV+RIYZz4aA8CWgrqQakVgmAoXErpKkH48GK8PF
ib8lc+4ZfWPmgQ2J4X3kK0PyKVPakhAK62+xFqg8uXWgJMB1ks1xxnFkH4lrJNsI
vsBohJV3NHiVH06XZTdqRdgeA53LfBpWPDnt6UlGGCUwKxQ47VrV3g9l/W4wXYO6
EDXPyZwocUiMPfY7xlNsgnHIQmHqfDHBcC3pTe1O1sz4IvcGwwIkF1bmeebawOYX
04FviYs0nr+9TQfyFu+T8V0jTk1j9nYAfGMFFxkpQHBgySWW1i4kWKvuU/ygcg4w
vuwdx/0eH4Y8uzU3OLYb05Z8+DvItDfkqxT5WbuPHDqpwwWb7BYAPBWv4VnvdWBU
v3MVlDBbVlMiyiNUDWjICDGpCr9jgGZYk3YM0r/ar8KN/xyv86/MJBQkjhIUDXXQ
9lReX7ZAke/3Vzu5wzculJ8/VDmiLFYw1c0omHWORdf+NkPcRBi/aPdHZg9FFELA
oExY24aa33aKWvrR8euQO/TKtIiQ/wfPN4JxrDOnz+j7cFLzr4mFzsDpuHdnUxt2
QJqqOwJBXjDTsuIwlbvDw1amKaXJDEMzP30BFPwxxg+WkNY1MLzde/fpASq3kaN9
AV5yrtrR4u/+YhvMCsSoj2/d6lglxYsoEOc8qWEE7bao7WE17Y6HoRKsCgcS2na8
hC0ZJxSW4OJerAA1i5gVoVyl2RXukw7FeijuxY+4CblUjsuufFE5kbT9Iouq1hAQ
d+VS9XbT6EyzHOqg3La2/ey6ru/nHAaX4xLRgWk+yJo=
`protect END_PROTECTED
