`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/2tWX2RUmNojPEV7QvUtS3Mzqb9V8ccAYjXw4o+PmD7QUm+ravu8uH+esjbBMwm
NZ+K7TgWT8/IdRpkbh6qpzRfuypyrppc8mlmFGmt//3BJaBIjDBxdkyYEnn7HVn9
xMF4NeFLN2K/rg7V66ZwvqwtHt1hoy1GjyUAkuBu0skbGleEAfH6AYsEYiCRHaho
arDKk0z/QotNGciRDM++MzN/yuW/fsvG2B0w9x5su+ayM9HGBCsa9yJL8T1965Pb
OZKX2MMz0uOHftpgDd7I2jZz0foPzIQFLqfr6afgjwVTZ8EMfdJoom0TzxJj4BhE
MKOWZJe2CcaZEVmZgxahof/Tvv1wde4wNpaEjWNFDogYp1cNBGHsPwcAQ2pkhzOb
QhhcH3UbFy64Pi/NawcdI3I39M8FxwaPpWDfD2xQh3gEPOCM/IC7dO7vbzYjszKT
Q9M1bmBhQCQ2l+GRCzu8wPaV5dANQwyIFzVaiNz1ZJfyDifFw2WwGPVVmfvZMzBy
nPvO3KTr0CVE2eUvaRsVFtOnpIPhPbYb9Bj5Xr1cpCa8+2zCdCVew38KdozI5TfN
A/kibKyiluqIQMVXYG+cTHWQvT8Ootzfwr6Wji0fyWcsAfYjciLMkHkKv1mKu4sN
9SoQRZzjwttpj/mwJcSSot2kJOv/Rod66+z1p9Dwa0oNorWlhCrfH03T2a/ahCiG
C1slmiaYxmVWWvesnmupWY0pccIMU1UqqKOvUe/5J8HBKGmblZwWmlTVlGUFSV/W
ePjcrFNnrq/s4Oc9iWzNJ7OwI+quroqkq+OmFA10bwWun8WA8vnoHPvcAv/JthAB
QBf400LYPgEkeCuExibA4Ti3ojfqYJFHoR5h0jqhqfZBJ0uSRQ+25ocIHFs00sl2
`protect END_PROTECTED
