`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGishT1TP103BlqsJOS+N0/B/cCG2dNl9DcGhqvBHodsm6lsWylkKR+cmK5AQA4g
dDsY1xtLDZLy949gqPla6xtvognABR/xqJvbKjX55xXlq74q2R5kM5IfstSMBovQ
FB7q9rBv+VUANjl8sx3QC44YGA+pH2WGVwCfdhJazL4Yc0ELpgRrUd5tAnF+bLVI
3RUrtcp/xRLpnhy4zPO8Rkw/U2HYwlKKonXpBPYbPzSuTDVej5M8RZZ0Sb7b/e0U
lG8VnPqj02PJiA5Trwo+pwGIIizuR5mqj9bSYR+tyzo9qiKDhzFhHvscOgxEZFKY
0Nxnf+v3khc4Ln1bTQVmS93bRCia3DmFbg8jK/lLImmV4t/6aDxeL0gAsFBmX+wF
XZQD+DQqm7JRRfWlCD3vBHNxMLHqJY6bDQ9zl+6KD+tYQSD3NMPqzilOF0NX+iOC
bwINn+CqR/KBmq9FXLsNHM8eUFl3yZ+fFpfFy9zQXnU+f73ZvTIT0TLE/jmIzhz5
vEKiDbyCcV80TjjLWwspJCl6Nv/sHScwegxpqDMUCNUnGRtZLUUznHIvfogDZHOr
ZdxEOpApIevLJBJe6qTwkFtNJk3tt7PQM86UCku2/lGzTzJYpjdRnv5Bl4heiFZu
Z4QYSxDEcHEKJNQkK78CTv5DeifigvSLP7q/sv0zrYTjde0kqGVtuiAbc3wzXasC
j/f2Hh8O4xR4ZITPhaQyu/LRgCnbGmNlNwxUu1iSN8S4/2vnr/Q+fCTHHUmuYtDL
HCC7oK5rwar+ExTM3WtwJXoeFrzMg4ZjqW5QH6gQ9gBP9ytmUSJR5es5XdeV9V1d
TSvdfz/OSVSqTGhY6VNNQ+ZPu0Q+1+0zjTFWaAC5XzE2Jb3/6l2IaY3YqiXlTSLs
cBBTYD7M+O5PfaRrTcb2FJkf9kkM5cZ/ynQz2RcIXnWhpRevi6FBEQ6EcHZe63Fy
Kdv9LfqcmgdeUU7n+m6Krvi2LwpoqBCmMnC+EOkQfm6rNfPOb3DLm0ueW6G2RfHp
bG3ChM0uhbTZ/LnnJQ2E4UHJQcyMaZTUkRNZp8nR8PhmQGc6wgpBimVdgWn4l+0I
JqExTEcBfwq6zjkBialfPwMatxDIdQSh8H+9IYgiD7zWa8zaq8flLU5ZBga0TIi2
grDbsaF+kBPR477mEB9O3txqVqymAhRjBRCU8hn2hpBcPAQxedUjqf63aRG3VOXD
U50XtwbyYn9PgQ5lgEOibjUQ0gIC/5etLuH7CicoTSrmeRS7FXqW94hS1oJSBztj
pXv/MLdady1a0KAKrCkzncPvCcbd7LZc6fnPt72XMcoQFcsKnyRnCU1zaLReydhc
zpDOY7HWSo5m0zSpBtlX8Q1VMuTkrckZ19EH42RgGQdknZtfcgRdlkHrg12Dkk9S
sQCVVub3RZKtprp0/Y2nUXNxgXpaw39Wf1T+evqe/iuM8Atrq0fInxvzOzX6i96m
wsLfAk/OyE9Y+cZg1yxGkoyg/Deu4Y6PMMDC2euO9TURsOA6+RdoJRKxsBdJObsF
O8xsLwzPvFp391c5kWBmtSWSK6gJVAYk9+puXKqImypXvxoOjibLepXy44AoELAS
R7KvqMh+Kq9HtFcHXL9DYzvINpJP/pajg9Jij8Vdo/YZF9rCwRATuxvxR09SukTN
GwL7PxlFYWKIhKGZFTpZX/UUzcz8KEAP0uXfV9abWzwG7ylhxUD0YOEGEBBaCiit
DASVkdkwk1NogB5iVcvh/GPTiu9NoX5AMnNdvobInVk8u3b9Am7UcFdKalN7Oww+
8TUAt/U6IOJ8xN8NVCMaKHEhQAvhDE01oznNNdwf/x43MTE14lMyfRC6s4Q9X1GW
E+bn7KssWDWTD5+n+9/C6P+dQQSWKl2VmSWyuxUQZt2dRiO3A6z65SFSHfcK9EPq
wrPZn69CY/xS0nvhC1NBASS7BpGqz9QM1i4eiQz8qbYFxt7HQBSWafDlylph4Pp2
U3wQs0+ccUAxwUAEJKmLMYx1e68PmZmmsusF0Rtgkfs5M2OKQ2OvcSi3oqOXY8oB
wqErooYvDZcQq5DVk59w0P87k6r3vaft6pe3aguoTn+Nuv53x567PMFv8vJEhdbr
9tGYvoPNVeW/9We/Dv9DlGsVtGzFB2Chssqjt6OxEnRaF6pOGzN1KKz5MTCo1+I+
ni6AtLK3wcdsx55cObMWihR3Vznd3GtaW1BMp+ZW/GhbzKpiTz4r54Ng3d1j2l7F
6pw5MML3kh0qKOXHXUFH22kCGTfiWrCcRRAgPScJaheEoDjSu6Ggt9HWj9gL0XnT
Zn4EjubS2rcIp9zgOj9E9yqkUJGJz2ky50RGOzR6arOntA2kn4xjznwr1p42sQnN
H5pmSx8UJ6NMliev0BNgWg==
`protect END_PROTECTED
