`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LDpJT13A+ULX76E/vq4+r3A3NgFJh+6nYUHEy8u+lSGDee/yu+qb+TlKnHEYzMqt
dwQ8Lxnc8HKjFDXdzfRKQ2FuckjplEQMsWwliV5Sx8fogTLRDt/XS1U2UlE0nx/N
Y/5I8SqByWrqZm288bn1UQqiOj6qGJLniKeqyblVcugy6YUtEtFo/QlMiGZEEF+a
Lat9u5s04/O8H5+pd/VKB5VjAS8yy2lI0JSzzgd0kxIDJKDYLnQtsYuI72Bq1VaT
6jbxrdMM8SIhVBJIgvbiNErm7Eqqr/md7+amaOTJMrm6T/pFvcuF+RcFXJsXcM2/
fVHhtpgNW7VUPS1WZM37lMIDagUBYCIKESR0f5oZ2cXr+zJmMpbxfvqhj7fY8MxI
uiaPFd8Q2XKcVf2453cBTuZdDiTkqxkLVn/6A4b3eIsob3ZAmgr5c47gwPE1U7wh
tlzFJyucRwn2rc4Q9XfO0WMYPyPM1r/rEcURRuqAavjygvh3/phr6KauQm+F/1zg
FVn4UZP7ZEO+0QXrTwwjo4A5qg3qjbGBW1vDqchJpEpXZB2e6WttopcVVqwAxOwE
ODiuUEPAJurVgvF+hOsQ5uL8ZpFt/EVWf1QTDODx+6MxILqQnO31rxAvYn8aDsOu
dAusgD2YJz2jEoq86VyAUdGZjHcN6PH1h0mkhPh5hfbLFE8+qEiD0RAMHizSY7fk
yGP5XL2l/j3Gz0idEAcc737wF5IRielFA3NXfs6ATb791kZQVgKT0HxdR1goLcEN
3TSTdeOQrKjhc/HUkua+30t81gOpS9rInM2Bv3eGadHewPWzZh3/06u25KZEVoxQ
EgfYjYNAVGyUx8XXldPLuNvLbs+jQ0ikKygn0l3KveNEfGmmRVGkopggyJ884gKv
+DjPnyG9K9ycjbu8K5Cq7X3QZMdJ5M1vBFnCOEIZYPk0E+fIlC/TtCr9KEMmfSvI
DwA1qwdsVzXwI3X3qW5klhydXMhERTFkw50He9TgLmx+ilh47q3w1MMJfjchuCtF
5Xtjhe3DisFVmFCaBDhQoA==
`protect END_PROTECTED
