`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBa6KvpURYoSCIE64W8qiu/9AU9sNrBJYSbZzT7nBgfJOoWF2E360y7WyZ9SWCGZ
GuLXpIlIWaMOfYlGKjHjSTEcj209WZH8n9IkiBTQrNoVA8MidaIY9KWlUFCrJmrE
/V2r+E2vpBQH798iDUsZw2z3gE1/jsTx9h7Bl74clfJRBsBqN9fxFbJuaDZKSErb
goaEuum2RQqXEjOXz6Bu/0wTWeTRM+5uWpcF8LVP7LmQh8qUZ4F175X8uaPfjVWh
ApAVt3u1uTlkmHqJUTe6VHCwbQdPro8j3cMi6CtmMSK/Nq+LJ0565zq8i2/eBEeJ
iTo9Wb7RgWxdmy97KLuSc+V8xe1YnBzTV4rNhaEfBjT8NwyP/j0AzJomjJX6cncb
FZSIBmcD8ver4aXYwP0/k3iAYURSNlkQr2ArWK3FXPZXuE/CBPASPsV07vTQGs3w
hMPupgbTjS3dMRZlEU4UgFaCGpvGS91KXvYZ8OSjnvt3gzz0Ut5U/09Oyw3YpRJf
MrGWA6fI4XuLJwgRZxqVbl7WoysKa7I3BUbZOZTAF7nLZ+m+yzYSYieZKwQYstBc
ggAglDxX8BYJUcGcroPEj4LcS6guEtD/uQv2N8yGHvMLIv6/L5j3ldfOepezpDbo
FTGXYMdMzta3lQA7neFTTv3IBdFLWBXTFkYKHMGZwFSv+45F8Tb9CO7aV8oCOmiZ
3Jv/CM5s581Tj8egD3qqozij7WKj7XdtiYXr9MO4GWg8YnsiBANH1zwtJ7rW8Fd3
JXzsPoV2mb1r4GJ4cAdxL0VhPRdtHCiuAb0pHBBN5ZTyuIyWKCl+6j0rckRlyLAk
LShP2GnmOVGkGt0aVdNJL7zk53hqptW0Xsw/RRBvgLvq9oJgIzQ3Zxomudv4XMrt
mxh9SpbN0jmb29hVFbtx57JY5JXERuS0tVzQTxcHqTqdSyuKh957v2/hcD9JHiFY
biPc5tK0O/+IxmVmyh8lX9x+Nb1uTL8+g7117JbUymCXlion83A0QVJ96WxU3yXO
C1++puWi+Ik1wM5vNysBU/5sT8b6N0UCWML0BtrTVZdZt7au3a+JOuMJBBbfcZzj
vVBw9LETAzFA2hnG+WCWqa6PHM2BchgCg6yKzbFR0ayDoKLAboMAJZ3ZjYeF7UXv
opbBnGzoJKN3HAlv6mfl9f+asyzGUs7IZt+SB/mrmjiuITdfgOPJxTMumSJRV9/e
/d6Uxm3Nxwf7Be+3/uTaE4zR+bT4vPSN/+L0C3ROWgIrEj0t+huo2srKmdr9Z2G8
vmfTT8UtkIXKyT7UvCW4g+7uKB3ycIXAN89xfi06Gq4Jh14FZDbtKtqUK/dgJMa9
nIO4T4p6ch/nldM/R5X3dZ5MjcFDcPMN9DwiR4ZBo8ccY80RjthvqeIMEOb9/bvY
18BerrLSbjdWei24HZbiYSpQaQe1fcnLmP6QC7KTT+sIIbRifsKibwbB+rLjQanz
osptn5uIfHa0OU0KWqfleN+vuzI7HQaMYIrJqnfj5AAtfMmD6zNrp1W2VZanhci7
iCVyWEURKH2gZxgzwZ6gv23t8K1LDhb4tjUfQjKG72aP5Z8flbA1lJJxZRe3lrCL
FhcGb48CnxjHHEnr8JMdZqqA0NUwnF1zt/i1DPWxcWQahmxxhsv2r8neaoznzNXv
ekHAbB/5I/Y1dLhFlH7ey8XiHgn932zMbM5oi+LFV01oJ4Ehs77j/i12ZU5T2mcX
Y9EWoCI7Dvphxaxc0Awv43QHNV/6y5UNZVbWPp9KkPsf19JrndEpbGbMEklt6WZ+
JO1M6tQ13BXSGHb+PAHMJC2l5DZRfdhkncGv+8xVoHKV+sOkfcvyYwweZjx1fWZV
HWoRAI6IQDHdWOBNe2xIuw6jpZY/RrqwwJN36rUIncOSFAhhX3/cYbWOkw4Wd2Y+
k0Adsv1RWj3SyV1/cscKFpU2V1JAeaniu1G7OfXppN30e8FftEqw40u/UaZitnT2
ogLGtVdAwxKHI6k6zYO3Dy0sH/M/Oam5HeIOMOF6XncrFje4OfaFxxqVbMKsz29d
CUfGyXHmCZsa5CGtflESzdbvYMBW/kZC2kiL6RtY8I1KlBStSFV2/cSzUWlz382b
XTNHygxLbYV13XkpS11NUj2xDIIy218ONjLLyK4dhByk/4yMOAN4t6ZgPbGehutm
mxZfKTssZ/qEdnNllRni0x1NsCcWTZXK25EquiXUGotXF00rWyXn7HjWMa1NgeFE
bI2FV+rjkeAMrUWCk5Qxx7Ejlfz0N94CTDsyJHXcUlWPpYHv9A1srIJJR33LcUL+
0W50q1Ay/8iYhdfQ3Yz2JmP49lfBtHvYpM5tVvKNdjjlJkSGhAJXN1/4kdLYdTFS
vRrbJxYmtkB8VokJ2jJe76rCQPZX9RUV9G7CsZlIxqYdJxZk2SfQDAD5fC6nCtGJ
JUnjKWLfjDMjcKg7eW3y7zys0Dcwk2Ydy7xFApvRzYTRRYVVySyroaAJvr8Dt0RH
Gejr239Hg4BSjqa+M4oRqQpGS+Vpas8uCcVgOSeySJfPpWRjbqzVz1e7nq0MyKH0
iDyiwT4JIU/uB2GOGGToC09YTIt8NWWoeTyHDiPyqzmXGIooVnLPuznxjCJkR+7v
gKDYj+6CQUCWjhXwpt1N+eUHJHILSAwT8cJo02sQsPHIjYt0hnMLw9/qxSwZYPEu
IbSeZViVdy3cf17V97lLR42uT6QYDRluBrz1nwJSkD8Z0v9i5+Wbwe6jF1l5Y9Y/
bOVSzocxy7EvxNieNNdZ2R/DsbcEFiay5d3GJ/3K3mpyL/fxC2zVNN1EqnZDVnen
TS2Ke1Ff1GLnCU5nb7jUQOFC8x7++ym8EKFlWh95m2RkfpJhkXVaZu+KEV2FzShE
7NCniXbvQUrPcOSFVW3np7yhjy1XnAercEAxp2KsOK7GtDoL3wlg1AmDcq/xO/ZG
hLSRqzJzy1+RfSvzz8OD5iz7cDV1Qg0XopK/nTOPH6TNt2f8YsGPeuAZOguGAZqo
GdmwzfM/2p4KSZrF88PNLdqL8Pa/vGgGvOe/lFtZ64FFAGlnyMoHPfarI+KgtQJQ
g0a8mGMVILZ8CMfNjBXc9CiPyIOUZoo0+Yrexj3XSpj6WrIib5aKiQSALbI03NY4
Jqo8eeNmD+vPgfxcxlK7xKTUSkBDlBnd2NpTjPQHi32kR3tLwsYH/sisrM1sSXNx
batwDooC4Pe/Q5QjIRV4Ni8qy7db0el7Qa0pCPK6assx1MPtzJWUN5o4SyEyT77w
RpGeAugq4gWYcy7oGfHITDZGDlNW7zbLSI0duGOizJPY9BTaMWbSE7BdciBrSgLS
1lkrg5cRhRDGx3Zk3+OH8XCK9nThb6nQdDHba8qNBRpXp04ENA6A79m4yZJoQBoT
p4I7tuoZb+QegSj9uQn56Op3OrtpH5LKSXjBgRVtAJI0J8QfeSJqy4jkvSkTN+dL
comsZrYnk5UCuDsKbrVG8OB5aUXzYNaBuHPirNg61lw=
`protect END_PROTECTED
