`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HDM8h/7bYN2B/2zZJFxqo5Inf3Sed75jnE97jQvQF93BN2HinCiFC17JuHLAq/V2
aV8mk9bDnTT+MvWPTag9DDIWX1i6JQlDaoQG/kk8NIVZPE09RLtJA4OhDlyMT/cH
vZ0ioqQqZKmRpXK/2xut4GTOUlWm1M64StGoIpZ5Ljad/Z4cPwr127NRf/J9g2zg
fX6ceGbQxbXIQoxTRzJi/rXuVt6VDIX5LPculHYSZ7XrOt9A7abCoRcDJFOtA2rW
LzUXybuQ/nv5ZkQiKXyEAGphdJQexrsnWJZe9WVqTvzfHAm5IPRqHImx+cAhTeW5
vMVO9rXt9DgW+NET3GMnz6f4BB8ri+aSp+li7AwVH9gNwU/WZ69NGCIcv90oBD81
130fM2FGChS56UPXxAKHo1f/uVfeydJ0VQC15JH/Q0UO7m1GIGu+bgiqecrm4uE1
FAqtOz9sYXiEc9ncPCvppbjU1p+tO5U6vEsfTvGK0zk=
`protect END_PROTECTED
