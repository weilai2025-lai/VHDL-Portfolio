`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X773txTbmKpSWOa1SMYN4SgY9tfmY3ZADTtMYMLd4QpKf+vX/2o5J56DQoe/IWeX
8lJQpaShQ5sUwHte5bZ5BBfLyQPvj4PkkD6p20wQM7fgxYWqq4vErYLYMvcdUB70
84ZpHuUUvMHeTibs/YGFkU37i5Hot6rofVY7+8StBaBj6M3o74ToaS+iS6XUUlus
FDw3H+pQudW+zQCcRghgacbIAn+et7oHG9sA3zeIZwOihkDcIGD0PlhHIUdKXlo+
YP+DecMh6NJ52i16G8ulHOVcD3uynmZBY3sB0qEt1DCVNRxYfnY8Cl3CEhbL2gfx
Dlmy5Qitcjh0UzWv0HOocagtxUQJBjN0//nhwPr44wVGOrbJV4LrlgBdtK+D2OhN
cpIq0TGshIJ1acKyarl39nwzy+wMFIi8b9AgJNazB0W2XU8GJSb2/teic4TbE1Ue
cAHpHJH3dbXbZsnE3t7fr/tLRg39T/TbHOALUSBJDUgaT1b+3DPt1XvPBGGLBXR9
NZt/S6+SNTMfV/h2LnYNZjxpHN89BMOtltfCWKPTArRlDcKupkXI5btKp3eLdpeK
drviB9agsnkmDqu0bLulMT1/+FfIZCe7kPjcvqrMmePVeq1IDMbN5DPdZo5ybEwc
vTC+X9SopHgcQ8qonsMsi7T8+mSamloZlwaYeOqlZnfkAGq8H47mohgZFhDHantL
/Jfd92vKphnvEYU8e+Z0IAO+QJot1ySbEXs0pINCFwqNctUd8QVtoD4PYW3hvh0R
XIUIazVJ+s1ZellClEoD5cfWXEVTOdPKNaCVErcXF/ezcCObAORTRPhL1svfI6Yy
paPbI/FggoSzt9da4RsAPzzK84FxecG7c2ev1LhTM7UCiOz8ttx9URdSozMNYw5t
brmhHgjDqq/D6+aUwCU3maJFM0Yey2L6DV2YKY+fkPDN6CIeYyprLEozP20YOKZi
tsj9PfXFlhXNYbcNSuFs2PnO9WHGo4zH7nxCh3PNjPd36ZcsbYxPXRMYAZ9NKxon
C6SMmLh2MrBINWwRpWzbc5+v6OScHplNL5vltO+fvUsuBTDY+slduannZ5SnGGl0
CBr2QP83soLPkFLTcP3rcYiHDt6Ffmr/4Hmgj1sYaZeG6bWeYzwyvC38vy+49M95
w7gwaYigp7V0gh78RKstnkXgnkrRbcX8YhAtLhSI7TEOGJo2umQjOuxNR7J7K465
XlEHFsZp26eu2+oVFIhRBHXsMFheegzqOqN/6y9Ft2o6S8rYtDJ0EBPE0jSqkGxj
3nYxUlLkZSztpMv//QIGkI5EhP5HOpgqSATUQVsB8szxMxv755F9Ds8ZLTsWZ9ty
8xsB9N5gS9SKMUAmSHyfzbCxgbVlGcA/IuxtJQKk7MJpJdXwfgZPc9VXGPTJyV/c
pWQW9IKLYgzaEgCXLjYOjLLSHO2m1OBt2xcQj5Rk5ZRXDoxag2s7SGJMMiHQkxZK
ZfVFaDyEz1C5omoxRJSPecT47sRROKe2J8Y2s+Q7Mr5nUw5cqXXChPNBv7QU42ca
5RQ3rRR74wzyyvJwePsafqQwI6X7bG3eNXYdpADBMP2PFvbTMxCUTSPGLF9gUcUN
cbjD0m5DN6/JrdxI0p8SwCD5y+/T5UtOtdGPeyn5DvtMurspGhp/KfKXhNayRJra
hynAPeVXmJ6AmxEPfl8+PEDwd8J1GGOzqLE97D3sCUpqQu4za48phld6/aWlFwbS
TjM4K0/s4ctJpMsZe5HI+sCdzfjoYCMkvaI5OpR7y5YT1iG9lDxNMk3QKoK/xv2P
LLsGvJQywWiekScS6LDjeMT+/s/3o1QWcvnBGIsafJXagmDxCZ0Q4/+IsynP+1wg
4sZWftson+nLqFwudccfOTNGvBLVtJeAS9C0N1803zeNBCgax66OkHz6JnXPWUJK
41RPgx1t/DQnfLJQk6nQNkUNO1dObckahhZa/ogw4cEq8zVkfmCKkyDgDePlz+8S
IICOXu/tFz5BeBYyhNr2NIhf2iKpk0/0G7Rhv+YH0j6Ges3fIP84EbX4iAq9YoN5
PQG6iH8jxFXXYpLJO056tBnszwggf0LM4rjeVh6Wr45JB5Q1Sp5ulT1GPwtX8TzP
LxLnv5PfPGr/OwNGXbNJlcUS5hdbFg8Oq4NOj5NMCcBLoODlTt4t4oypqBZRX1ZI
GYN8nd2DTVqCj0bUNjSDLBfM3lyqHMtqkvrpbHq7pSK58vHwNvyN3JRAXFOtXZgw
hMij2e6eboq39E/VFMvG+HGmjwW6st+V5GxyJ1vGdXOqnY7bgo6PZ02EQD3ixd/H
ScLlLBFLl8q2luE6ygMPOgeC3Z2BsnnzEw51/brDYoau5Z+G99y+fo++DNF/ufZ7
kXcb6m0Owdy2Zeqn781TeJND5IGx/xIxKyTzVhnbohqHE7yp+3muLWOArQAmmfN9
F18SeqH9n0AaXnAzGJEN0kx3j00n/dJxLPhLNrkWWQ6rszy5hwJwHNJkdkbTXKCG
VpenhkgSxd0XpcmAlv3u6mn7J1Be/C9OieimgE8TNX6j0pOm+ePnjtqFlbPWLRah
QA7POhka0fuQikd+8xi9TxZL2XQd/Y2NkcctA81R63sb3+vurFBjp22xpQ/zsDYI
D9j6Aw6IK7fqX0mbjaDjKulQFaYjQd8qeIICXqOAV6Kfd78ny2slr0zfryTd/EA6
otrH19QlYAOZI/k2pyD+KHt7IBykiRIA+/9MO0NTRcbmb/K5EBSTASEaNIbwKEgx
q//7eSmzBzfr7ej7Gd2gF6rJOIDCLxdo6+F/K9gLBDRONie7Z6taAQDrlO1M/Mc9
r+O31t6aC0roVziEW6HagIVs5v5P/evbZnuLKpfS/Df7SO7x8oymdDPkbtN3MU9f
7EfdEqwwlSuQ9PxO8OF0tBRtNhVm9TLaB2P5QAB9VDzl++XKdS1Zd/nbLZ8Ba94b
Firz+cYEblPBTwYnTZ1PiX3ctuOe0ZD59uo9FNBC2MSnlMiv66GyfHGTlssZf4xh
bWG/sAr1gu9xpyoyFJg+9er636OSpyd+egbmg7YwePHvHTaa76ghQkzWzfXL6N+C
cu+DIAJurN60Ewm3JzFyYrLn45xYFlI2HAUfedLj/4rFNuc/BVkmiUopmESw3p/q
wWlYpVWB6XDARjR1levXZ+kE13Fn2WjHpX1abw9ubdHXnZWB6L5cPKBZn6bx44ic
4WgkC5+HcjTImRC9LPoKjvv+AZcjTJsAJJqtmnHWzEUZNtSl5LOgWt8X8hVyqjHe
AIWXxJlE4/3LWjYarT+lSzL7iGyXz5CNz6shvACKCs8FeI6Y8c3dtqHF0QoOyotr
q3RsqsR01AF2D6EthqOaKYNz+RF1/pg3LSpzwjLvN5bpujmH0ThPABaE5ozEGO5y
ba12eV8rTshn69k5y0alFCBt7RAOkbrY/nXXK0SCqS3u2z1iueOBrpK3+TyiZYXY
t1BwF5e2orxBcN8vj3B89HtkDOdPkAX3qyCIkI2OQxhphve8wDQRdduoLSql+/JB
MB4dqb4v6tZsLJ6uvo+GqxmL8ONhKnleixFypieqGyFDVCdAb+sZh3TMVDNFNc/+
79+iA/l6fXladt9NBpMTZzbS6aPobvykGMl9hkdnrKAypfBiuKxW/f4NnZjkHnhX
Ws+wsHxIXgJJPIRsaCXBl1fgK1DYVBRdE4/+P42RCohGui++B4JKbihHlb2BGvxX
Hr9PULwbVkYikGMtL+yOjgbWJ2tH8iWPeT6gLLwFC/lEgJFq863s9390e2/+aVSI
+4I/T7DhOSS6c696NGCPdpPq5jTzthJjoIv9/fqSGHbU/dppvT5V8xnf25o3w/ET
bd4Ygku55CYN7Ef5IUqQvzrt6nlFZHPaWG1tT0UcicIGN+GWTIyTf4lJNHvVjm5S
k+m9XHpWQOt40xvAsp3bGUzrVIxRZi0jtouXyNorC0tXwiMAa9eaCIkZpenWRc0w
Bqb/iR55Va8+7AqPh4ATcwqK2sfxGamHrv/y2WPLtwVv5wDFeKJpOssQwG1Q+a7s
YiC4OwvVEHOslTG92T+CdjVZ1Sx1LY8VRG11dZDqxAZZAX4NKfnb5s6CRxrJKjqu
wHBNIAZODgPXOjVrN7ITM9bEpxPCFRRcF1Zc96Cufv9mAiMddoW/DV6BDW7WJ5d/
VW5sSchwIMPc2O3MHBOKCNyGSH1rFRRLjD9n8dkgdEm3Uwg657zWoaHKbeKC1xxI
iLPUKHU7/OD2ZIhOVMMzZABe8kVtf6I9P18evsvniIF4gqmrd/aB/u/lW9vxPfEa
O56i9yKvgDVB9I09x0wRzDrMuAQnY3DvnesEblq83447HBOgvSZ4CfNdHVmtGeb0
2fFU03je57mUbVQskQ9L9JgimjKPj1GPlup2fNOBXJwNYEXOCZadvGDvvWGMJC+f
lacSM4x6TZHshSFqVY8tElgOb6M2L3aTFtf7jqQl8oZNT3YzdsrM6EKLteDwi+Pg
JeyQGgRL1xpPEdB5DetcPXDxZFGCULKUICMlQlsPlPe3XmWkpXU1dgirYuTblTn1
PlOGRLo+KGVBo/6mluqLmeU1Oanni04fe1QJdL6f+a1GSEssLRcsGLI7saEhN6yd
Rq758Sj0sKlJ0ZxW8WLVYl7bP37vZUZnvK0SjsRaIEedx/1ZiGoorcQMPcgAPSTh
3s5vQk1G547eULs6WLGqjN6kM+u5ym+temafR8B4k7ViNJEyoDR4t6lJ9K9scRMY
fD5mz+WnNVipqnKD35WHnXZMf0qd/eFfoXtuqAFdJqsB7T0GUhrhGzZOTJArZN+S
nWYc1JsbEYGah8GF83sK8AoAv2EZFhcMGEXUHh/wraT4lDACaIRZTEs9htcJZxnK
uVEGw3Fn4jsTFbYCEqRp5aO7T9IbckBR7tDv3tLmWQ6v+TJtl2Hie8TWhNnzIHFZ
bCpe5cn9KSnFSP5/Rsc5CrQGwJRntsjudxrMSTJcRanyP5DcW0zswe87dgRPZ8GO
x8Nps6X0RuYBasFQVODbLbm6OiRP7EdkQZ0VGCusT+w2YGfAP2nf+D/5EuYZ6US2
XcoSUy8nWHXPWdhvnTAZ003CiP2082VT7DDeo3hjmVO87rxrgf3X1alpy3Ms62HC
b9uBUM6BYIwKILGbkH63UKv6AO10rkfu/ergPlT1zz0+nYUwfyK7khnmv31eJ/KI
uXGuVj/8juZ4+n+1hNva5hOfzgwCeJYmkXyWF7W0gyGTm6Pjs9hWSR2F+rhCW26V
Q7VLzn4pV8k4XWoBEzyCnW4a/FmLfknIi8UFYFLiwIuAfS+Vp4RqwOAFROuS8+vU
ib7g0ST5KSRGbCPJgoLR64NBHnMl2eaYw84TP85h57GVOvsWMnVH9zQXb8+WVoeE
go3LeKxhic+4MtjjRpz5eFFdD1DssNSzQhonkh8MfRjBIT3A6Wu6YPEQsBd0ndE7
CxYjffk5iX/LLX8swSFRPHPGj/e/gxYA1VBqdzw/z+HguNN1FdiO764CrzqI6MAb
KhBgy7sf5uQvgFIJF4bavHBkztn9c3WXhqFF1x0HB9uIC9qh0EMNH1KeYmYAW3IW
T/4gL8o5UCFRhRCHNS97lWzFHXeaJNM0QkM5hj4vDbCAK+OzWmkYHQk9/tZKcIT2
rhPoS75yVEj94gpcoXaSv7WPSem/khcTeCdPE2BdV9F5yOXpwpfQQ1AM1h9zf4Zx
hONO2xpLVvpLDtgyLGLXsDwqGXEfmFRsWEx6dFBFK4vDemgQNEMAx8rdUsgBLbet
vQjVJtJBT0y6gNhbZ66HWC7GKZ0ozYmWGCuP0K5yE2b16dL9OG78Q+/Syht+DZ00
AXiv5FaK3MKOVIXX38tgXItmrRi7qHXWU+cHFX+h/FwAKtkwOg3k266Mna/+rRmY
K2tJ6nuJW+Aq+2yMzg7em9BuKsdH3ukIvY58a01iLxsEul85DoPhoms6o+5SWDA7
xJd54deJ5ZxHYgYcVVu7bMpq97VC6kjoxtN1Ni/X2egvo+ozqgfvIeVP/iMlYbvB
8CMhg7mPm0jTj6tWcdxPf2GXMnnbuHM2v4sTykmDZXHIt3kkVDPNQLfPJ233iBcX
Dts4W0HlMyIpzKBKhtAIUdX2eGIrElv+9qX1V46yZXGvUEtJFKPDx4RZC+MIcBly
M1GsikLD9g51qmZtww9vLD2o8vQ/cFPBA9ebOtOv2ElKT4FT5ZvQPprIpvhX2Anq
NYngA5gw1aoxEOG9qucQfYrp8jFgAm8sCi+OwLG8CisOcipm+y6x8J0AgnqEhb1f
iIsOKpxKYKtcJjZrWs65eiGMFcc0uZ4o1lo5jtDNjCMQHmYASWghq0zHG+Wi1fcB
G8bfJlVRQywiEvktB4LWGe9ibkfw65EOlAlhZB7u+AFR417sO7maw7jVa+7Y0jk4
2R2bgWk1cGie4LC7HJbvjjXRWjWdjeuty5Hvk3Gac2iBMXgWa5s2GJ4lXaM7u8eD
LS+HhUdNHS/Fn2JZxKeLBtbUPI1T8S57Y8rRE4SJY6uV/v6PFFeiVLL0zWJ3wg5l
ca82Bd1FJi279TLeAqQhHR63KKscFaSnrppMFwQz22Fp88kFpGJRfnS2FQARuqCk
lzHJxjU4ish7QDwm6NsGE8noUfEf04xkOgjYBaoAfYonaK3jb6nb7/Q55zfYTQAr
hN0VHJOIwLFFgUZUB+BUZSo0kUjoZ09Uf6pBuCK09o5JLDflFQ75wiyK7MnRe89O
EIzpj8YtW/uauR5v8Aozq0YAjzzTEcV8S/ieccQdS05kTPW9kLhYYYY/H2AN/04t
09U0DzjayADTX47dHAQaD74yKUdopz+7Au+qMMNWkCxm9cyISBSaEhkO0RHbOxr6
TMaLSBvYee8T/4NtmP53nYq+sx/LnZsSx8WcTfO0HxpjFHQkVWN29437K1M6rnyf
QZoLOFwuuuq4187xcNdIzUYHe/wQQt0ZYsvB8KyiaofUd/Eahb16vp64V8SFq4VY
ErdXj21Co/vIz+U0n0LFZBd3UYyH1vaZTvugIJnT4XuSOvSt9zpNtbx+zaV4vJ62
+Ygc/xDIwlZhA8RxAxOfgIyir8wJ7BshBtC6h9U1ubw+TeR9Vk0x3ZYr6vgQGPpl
hocBzwPP4qYyAwwgz510jbwyhfWoRx5ngqYl3t3Gzwg6EGbDiUP0nnDP+fGoQhvc
OcDTntg7aLbDB4r0TLzecP5yD3upgBC3RvycFZ/8SRwp2u6KthrzmPGktiorEiVg
LGqhe7GuSD4CE+FQ21Bpq8Q0GAI6FTGLqQBH9FylOgtuXKrZNdSTu6whA1JRn0WZ
2iLDjMAdxOObh/crnfoY3kvu3cfj/m7p2F1SLPbgPFADHoeLgzLg1VUy/3z1NvNk
HV0u35uYdF62IeshyXg9Chh2PBQzFebyOLghBgBv4qSmI7+8BQoUAL6siWGdz6r1
PscwPgOyzJALPCSG/nUPyB+MXFBUptIoeOBd6IzC9VPzlwb4CtrR3LLAOWZeltn3
98wXsfGTIMegzl05wX/z/4rwanSl0U24CA7QPiXDNVengb/4hA2mJmbqwkIquDZv
OJn+thaAimfoGsEq11JmK48Z4XG+CFYgqZ61BAcAsGof2cism2UJ3/IboEjuDb5h
/Xy3nrHu+X15whDCQj9yud/4oUMBbdXQh9dTnoVAkNu8JqBQGGOFaDFRDzcZHUVC
Xl9hKNu0KDT5ODTFrP24VZtvlxO5gx5Fd4YUw0zbnfHuklb60sI5WYj7L002PNiq
u3RujKplQpAC02FKOhfn3HbkojO+N0fX4ysibb0uZrA2THWKGmMZIo1WtNqOIiAk
H5UV1S1TZtSo+VVSi+8ng2pIewRnK96NnZbFnpvp4w6wEtZ9+qYQPye02mbI597H
MPj2h1dG9rrWFw/7Z5n5zcbD38yvvJA0ON+0ddQ4/rCsOorHEQHeZ321j3I7QAOz
x3DabelGy4LVhpFfsrdHtsRJZFwYs92utjiPwvrjOLgZyE3Tn35XTOeQwEvjsMyx
/kDAszKgDsS5v7BbTDewmYWZIRU4AnC+yXVJePyBXkGdfhexwqsPUej/ZU2EXad5
7ieJGZOTNopN3CmcqxAdEFJxdo+D3jJcPuhS63JdwubWI5tI6EDuO4KD9twr6/Ul
8hbGIdvANS9+1JGTxx0PyW7JBoCBCdqPZ51Tk0YV+CaDtJQhGjni7fGdXl3ENy4V
eZQ/OqzmpNlZz8o5qrVy6qE/xGkxpBWKnnDjtKDoavxbm0aybnGRHzqDPOr6Qr6M
Sn3w7O6ZXAj4NpxZey6XlCAVuobyVcN0c+TOAv0jWYdqn9s0deJ46rIne0Cf/m+8
AcxlzAFlmNa99f0iZEqkJ1oe6MaCBwc4xeL7E9KOPKQWwUA57Ig5ctj7P/+V4Uty
9eJKNTRVonC8kYnbeXV4u8G7dwbd4ypAOq9+TjLWUPri4h+APbPJdGEpcUvN+z5I
xd9wYL3t0tFASkuG7jASkXiHldKdABrtDbqWLFlPCUsr/tv3UIyrFL8klwZV69Wc
wDK2B2ZFPAhoT8fpy1vL0FXC+C/8w7TipaXv3GMBWgp+5RcbA2UYEi7KurEN8r9T
EGkIDKbH0NJBd0O/waZ7HMJmzlleDW+6krEURonHiw+Q1N41CffZm/xHkQEdK1WF
KsmdyE6ln9oDldo8TBaoZDFtrVoOSFfiJX/ed1QInt7MFoceGOjm7RTvRVDjB868
dfrA4WPpt2xigNTmkK3pE+TK+wRC9iPaO0+ysXotmNQL7EDKGN9iHUuTRk9lbwvf
Bw16FHbHHAhuw/HnV2l10ASydP97dA6I2byy7LanQ1b4FuZRiZ4sTeT8l8cTPrJw
1x5ikZe2E1a0bJMFNefDSOdjURPnppZAWk413pcSGihatkYBkItGelnvh9CBCcje
2z5zT7HNrvx4OXX7tryGSuVLEhVP2cS5Lfmp9Fd2+I7aq9t6J/WMYloyZZMu7wKQ
Mq+C0eFkqtEf7pRCo2MLgglbaUyCyzm+AJMDTviUluDIIyoZcwzhf867or/9uMpl
91CpnOmKXhIFtMa0hdqENI31BoRz+sXsK5UyKQTux4QK9LEP6e7mz/cGwE8aL7vh
IY2NMWlx0hUzi0xIOeB82hKvwNE2soxKYRulYZOdR7e/Tun8npjFmUW/VgLFb3MA
CfqwxaqQeoCib4dja7lj7+n/U5KGAAxtIkLS8bvj4SiaQcfJD7uhbAlXfOBitRZO
1btGv84xIerB7Ln38FTShOp+cd0tXgh+0UllVmf/B0UwtE8xr4tXfNdBRAUxefW9
hTaTXte2vHpbZvQLZbDczRNo5JzWqsa5bOwmR4ExCPO7j8VjAzz931GFlQAwcrJR
Oojns11jA4aBvJB8wm0g0gL4mSyFG2XXzDoywdSMNkVWQ90RieE8rTpySJpACyYF
`protect END_PROTECTED
