`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cvFQAgMYhFhTefBQLzQttvYsd7QDwB43FM4Qnr42K0aBoegAzJC0gj0mDYuGzdh
yn3AT5KR5Zm0MDJb+34kED0AGcYli0lARZYdnuHFsGWR/u8zn+n2DUY24h30vkio
YadWlx+HXp6dYGaaAjls5wM7AXQkCKIgUPIsfdj9oeHinJNKgPcUptffzFwqDFbc
HIzH1EeWX1bk1+RcrhMXN7A6z9NzxKbktkQ2sYR0+Qehct6OiTfebi5onjg4o5V1
O4Ga3abUiVjiQI/fP69Z2a/+akO/sNymCci10wYGv1zEKU0U+L+W1DT9YSVlSvKn
Wxh+kxIolBI4cDQJxbuJS6K5a6T3+uLd36P6sW2X2ycqxb7mHbUv3te0sxXyv9SW
bFKGyuqE14nCwK2o9L5nMUyvblayTQ9/NQXEvudr5KX+ZQswqm3TNJl5hRKMUmrB
JRMJo7Ey6GXOsL3WhBsTqHYHidmL9zz07zaZ4O/JSqARO6E54DKY9xHpL8EF8uBZ
1ucV6bIUcUWGOC/YcU/SnnY3HJcesC7GjJQaRaiN64CvoCg2CUBChr/aKXf6+OR0
JqcepRgDzXVvA16x02IzQ474hfT+5OKkanA9cq8S7kugDk/N5vzV0h51+an/WN8m
jdSDvy3vOEq4d2lRfNp2g+o7Mh2k6LmTRdzvtsnWjO8poSkw4VV9Xs5YHywoiMu9
nYTjpflMtUOknKYYi6Xsh7nx6cNY0m03/+cpaAIUQbneRobF1T3f7n3xvBTdOKdQ
GD1fOCNXNa9QDv8VqpKvbvpHJLWtJ3aRKfVcGF0Mlhg7sOVGRqeMHEreOzXCVDw6
cSi/7Fm+Q1rUBACQsqm+LskJH+yyevZJc8lOSMH704CYbuOaeSzdUZPzObgB9Grb
hoiGUYiV/S+b5Dbj53toTbBlSQyFKvbKwa927VQMEOtsrcyIhnN+9rBmlnv7CGj3
qT3o1UzIpnX9OKDZaaqxKtB0qV0TRljfCwSakUPUWBZOXt04DfIFrQkBfZ/xBfQ6
NvS/nPQVWta6y3CswvVkQ0DwtWFZY7l/ZgfBhqyPdwwGMB1sVsPYgC+ELpUqf6mI
zKKXPnAh/e/JgQsA1SsrNkhdq3s1xXpH9yh8/KkwtZmasGrKVxewNFaQNzR32P2x
pAlyrgEnGpm6B+bm5uJojjshelaoxq/bv0NHLYNVn524PshXgo1gqepxtgMJlR4j
6ouvAmRFbYRW3+Uh+zWZ9PLV8mhrXjoydVoH+ZRcurhF3wTXXYIdJBBQsd63wpH/
jxHkr2X3Z+iUAsvtFQXetbuWuZL9UxnVjp/wNVKEfHxRE5IBNrJ/Xeioyxb8jin8
hPY+CNj3ZitdF6ussjdFf+krP+m9XExDP49DRfdFrsv3l3NQzZQ1uPgdxHFH7+3q
FG6yfWACtsxWcwVFnWyIz0NFkQHKTWCRlwI0LeRhV32rJW7kIvCEiGPWMIuPgY2s
C2/VBItHEK/QwWjb7OM2ByIoHsjMUEoNBiZhZ9ad1LWL7roBlhWIAPImGbCLHbBC
Q3HSuW0eaN7F7kdfNcHoSOVDfpn21IjZV+25OX++5KluR8Lr/CzOghUV0aVbGa3K
TWBhKN9rdxy03GqE4tu5utFutO/iGaJ1YAgGIOSHHHgTmXk9ISQEOW2zdgy7QkTJ
qtaCxLbxS7/Z/0PSbKo9/Ipew7am0cHxN34EFenWot82YlZwlWr/qytiSSQ4SCIW
SzhO+JgZfs7BRM9bFKb1FN6L+/ixN9jUgGwx5jsdwNzRsLqo2iGd5rxyfXkiH45H
`protect END_PROTECTED
