`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mk1o4vvVNyn1NKZiZqGq8EkifhkL1c7sLIhfl+SXfmENcdnzLgefwEvhw9wtbnEh
4aBPsE0fQ4IfQOEKUzpZoSJTmJRRummVV6NP3kqe2o7lJvrQvWYxh2oylkjN1w+L
r7Ch0OSwUA1leVoF94VxaV5F1i9zwA2RQKXVfSwxkSWxIDUJLMbG7CtDejxWgQ6/
275aGRpqjYC8ngnlXHqt2NlzCjp2btW2lo+w4YxgxdSsxAqAxyeSfIc7hdfQlHHE
D4NFbBxEFndz2850LEV2YPgqbt6KFoKNRmJyaILkIcMvc7dro0p/gvtUUizPmmwH
W6UZkYcsuAyajUiPl9NveC3ky+qPkhBA4t4B0J5CDB01XDSFuoEySJ/Ny37e2tFI
IHaj/gxREWtR3wR9xc1UuhU+7llFWw8uwZ+JytWTW8dS2dmL5mVx1B5ObhVpssp+
b+0zoutPIM0hd2UB8gqTtYebs2X+grUgrLWRijd+ZUqWKTtfc0UXoJF9ZeuzcXak
ehlROLZsCtupLt0u1MRTLN8h2mkEVE52KaZRjQaDxrLsVtduJjhQasBcfjvI9Kbn
KRYK/3eo1XTrRTpKCo25Gxe8Q+SMVnKJhWGuYbnmPqVFTYR4jjl6ZwyN2LjkhLOG
t71s16znfkaCK6acdM/vTw2OE90VqaD1SP3b6xnQ8st3zdJwkaXmtbsXWg3POxbI
wbDtvKlggI897iWkmlO+kCUZdl86sONALD0D3uqzcnSHNYSblMxckAJol0FehcNa
Q66Fh+Ta/06iimx5f5vcnA5oVGuS8qmrF1rA7hdN3F/XZo5eo8N4v3vdd8JHzr3q
`protect END_PROTECTED
