`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3GFws/JzlCwIzmY1xOzSMDgG8i4U6142yXzF4FstqTODMRGGJhXpdAQG+f3pCgc
UubFAx6ajL52UOQvD2b6mmRUO0+kmSshVQgsgYwkClX902ijPuayt+7uzfHqRLPX
WOyOBQBAnSAgcvXrGklxt3+Jz7r9/sosqnLwuVNVuqLYgoBSw8R7Bq5OYqmPnWVQ
4Xebr3e0igWdhfJ0d/alOVpFVSmfQfgBgoCt+DVnW16s2GUnvBZsznR5JIec8T7L
/1+DiSzGpDEnbFSQRZi7Phwh+I1Zq7QjplSnIsT4CWs1oI1zCYjHkO2zVXhGgESd
nJQObGewnUaMWK1jOoI4q/hFfdGju7aoIsHx1cG4WzU8fKFIszf2OYy6u7Zf+jiV
MwLGR8WK1N/MKZp20m7XpwUSf6o5i9s0N+b9LxFqfXQsj4Ymx66MdBvGLIdzXu+Z
Nn37LjrUP8eLTGuoaVYcxgHovP8QENiRnIrv6KfqndcPrV5N7S9rcfELl6WjpG7m
djtiQ8KW/kqicgLT7rtLOKGBFATFkX2ILEOdEhhrzcoj1ZnCtiMqVZkelocV5+y8
Pp3x3T0D3xEpi5lK5WpACoGlqPRJiGFcLWJaKynoKznSqAl/ao5taZwifE7Eu7a3
dS1Y1WKPM5Ez4AfGggSkRUcFrYFAFKd06cmBdoFanSdzg6e8AaYEOtdCk+KNeKbf
bCeps6c5jTPLAcEdbU/GajWMhetPgCaw1bdP5zHxcbo=
`protect END_PROTECTED
