`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tSgwmspU6R4i8xWNikTV82EphlMZGy84ololYUeEaj6IxfYHW8xW9EpqSHD6K411
/QmWLKns5Lh2XGay+r5oIjrm7qdE3gqcPs0fRzn5laUFrgwZTwfXWtVPzXvhazyO
/KxoNHxv129naX96TsRPX/2uZfkBu+RnTSfo2J8RqoreoOEHbeL6642WbeMhGmcm
VdSEDb7SLVn0nxayYriFeBe9l8QjfncW7n10WTitismAz375ywwMWOgocmfJI4CS
ZtDjQgie64XesiB1VBwIXmEIMupQZo/mg/NDZPMjmd6sj8kBJ/iILTcCq1oyzQxx
TAdVd7KOUNhQgG0nyCS1UGo8QOIXazauCz9wJakRNZ9eEKalgPYj+HpmVsbbQxiK
OtXk8iXyEjCrDSGNOgDZpJQeVfsLrmZ3BXW8Pn97dRpl6BRwK/sudY/Fmq48gM+P
Ona3Yp/ohcjC6YU9DYoen2833Y4lBHVjpadMbBVO3nCkPumPqyGrLUT1hrW9RNeJ
EuhQJmTRkbjqzP7AhmbWUSzyw91r/WWJTybv1FeqCWv1HMKyoeOyuPsAtclamu5R
7XB2JEpHi5fDSgHcsChmux8gIu1FjYG8sY7oDw8h2lb+6T8aNXma+C98DbZ4O5xr
WB0N1EradCY3bPiOeT5lkcBSuZBYv3Cvs4pvJnv/5OxP1xHjekAbpDWBou0GQ60A
p4eKM3nTol6VsysZwCbSryztad014uXzZ+XsDnd0tBKyGYjLFc7utaxS305oeLvm
gIZGkKOQ79y59itAr2hMwkuVvq9LguxXl5j7sF5OWBNzJ8Kv5jzyXtT7gN9vHIzA
ug2t9j9+7yB6Lrrja7Fh1iYw5XO9SNE8LZIyZfsay1VJd7ug2tMfgGWhGaLDTq2Q
KCRENfH7wpZMtQQxgPfVgXNPad7ud28GMSItRaMe0GttN8KWb2ATwL3GXVkKr9au
QCLQjf26nvwuEE2z1371Tj/GLMLFG2ZBct24yX2P/Z7yLafxlSTvMWe43hd7FRp0
JSJn1Jyq4lSBazzg3s+qAC6xFKyjrh+MofvxcH1fkeE7puEPG8y8l/N8dbjuWYgr
eQSoAOYS/drxXdiCmjK0pN/t6/zSouB10VLjjeTDHzhkC5nkRLUQFT1RAUMoLyWO
pie3cZfCPP76bAnbM+TBRce7qJJvtr2wUvGA36MqiTt2VyWH8qkofQ93uGH1T/e+
Am7ZJlwpzNzLbg+k6wVh8ZQgi0wc/IIYI8VIiFUd0R6mvnLx5V9AH5G5+8cSE5PH
xfe0839FkYp/CKQDOAtAhvHwvNxoIMhkKFxC9zg8FxVtxFRSBRjr5YV5yLe9IjAL
Q/kbYkOII6CdtNMXo1FyFYEOFXaR6icI9KbcDAHHETeT5AuWDFMgDc3fOr4R0NhX
1mj8PScdVj0HtqL7Tq3tX4YykWYPiaXLhbUgc3Ki4MuEHRqxcLS9OsTkg70aaxOM
AegbFOlPb37G4yYhVERc/d/WVSbtclNKkYOvA/lUCFylbS3LZ5JWwE0/25NOkuaB
jGRHjxuFcrb10QZaBOXNzi1Tbucgg2pVlYBxkf0WaOuUE15A0WvOuASKEjqoQ1LZ
wTchIlCitPsfJuHlQ3uHCcOpZE2fAnn7PM061JJQxyQDLWZT1nHm0hCfyZpp/tyQ
Ufg8SWVCXO67Ih84i/uPHcltd1hNXDmnl/ttqVdq3ZeL5XIr4vQ0lwfD9K2m9o7n
v+plNSb8JsfvwJxglbIBCtS/uFIcEXxOD7ehczAQO9Pg6j9GHg6r8NoxgRrNZlNT
Bh/u4mv7WeuMylM6MeKvsSU4T/Xd5toRm1pe/WwKm6WwdBKf03IycU2ja9pVRPYf
7efxKwN4EfvYg7b14SvT8mQZD2wLDe+1sdFAbMm1W6N1ko/rGXnKISlmURLrKCvA
GBT8uLtNFfHS1bPRK8Zsk5U5lUjwlulEw+x9pyRWynXsRkdYXZwbhoe0PMpdSW8/
Fpxl49srVOPrNe8kq1247Lh2Q1F7CsV2YmLtm4nME2dpupVKwqp2Z2OWDvzuoC7D
5GGPo8U4T4UbXsu/TPjCnNKH1sgpCKXuKfhmkSeAcjcR9XDqLW+lF01SNBUhplzK
76swfNhYp1WDepUCprb6MMpWm/KIe0LXrbs0hfF0govgxxPp5opZ1s3yTABhDefb
vTy+ShPzlviUBEWfvK3Y4xRV8zVWw0ryYhVW3LOQVovuFqINGhx2Lexr0fJpYug7
KQV6dprRMuyXWjQhAogLi8uFgN+l4UyxEprCQML7ep75JCcBnJQQ+QROBN+5vYvP
Hea+AcaadqjFCCzKvScMN5QLSylUFw0FdLyT2Y6Se66yF0An+PqDT7bldWrQosEz
7cuyT7uBS8QQKh4ROWeqek7SUckGPXEX7Jlg2xMKWdSsxD1ga0p7OUWb1OqrwETG
HGHjL1Ffc0Qe3399LFeVNL5hu0BAODCG8bVpnMT8p3Hbmiry7cznrRuQTFULd676
4dddK6Q8of+1CyROtxHWHlm0OFRrTH6Z8udNiX3bIYtR8qya3kfTTTRvfLeyQdZD
NTpebl4upFoxHk0CQg30UYqORlbaimVS0tWZZ0HlinsUQCYkGoP6MP4EgHBcsZur
/8AxwIQhCckLXAFOVSTmEfwNH35m8nU/a53qansPb/FaNDxqmgyB3xioEER2yaXX
F6/jLKsl0OZ2zfTLSbwU162xTHFFvJVI2wfQJsgIoYeft686TeJwaJdzM8qn5Eq+
ynRhT/U+J+d5IXWeObPvpmo549eqTMktVU28fygT+HV/cEUsvFQPMzuoVb8K8WRc
NC28CWFTZ9MNi66Su3w7WRtN2gYkVSCXuJK91bCn75tUxzPyO5cxrfoAr5Bvfl0A
IpVrhQSVZFUfX6Wgdcm3IZGt9sAU7iuwZ+yOlYRQo2eplhwcncKF3FSI9Oz5Lo8g
IInrJo+bH1RA/ApZFsme0w==
`protect END_PROTECTED
