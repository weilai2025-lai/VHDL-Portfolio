`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1ThXQBbpOIizxiDj1s506qI/wdeUdGdGGoO3utswEjGXkehTi2R6XdnyTLKkuX/
HcoBYWBV5nqwt5Vlncl9928bteMbg1+u4OXInZ13HdpNFQEOJOU80uZTzHghilTv
b3KjYWAL0chj3DyTCqRBsVuh7FjhlvcRnE6O0vS0xmueUWbtTKjj5+T5Kdef/AhP
vY4znuXDIL1jf5CGXjv9Rd1zXBtabbBwkltOmO7NYVbjusQO2/O1JXLqncCasJsH
PzlgO4dDtRjTitOLcJ2tZ1tW6zJKLU1v/WsvQaMM54Eoa2NOjoMVcgSiED1udrrc
O2ULn/p79T2MyP9qhKBpdUsPP5snMw8iXJbdJVrQ27npQUhhAyYIy92VFxIQ+hdh
QrhdCE5zbyVoj7OhqikjaVRBOrZw2gy6jJ0vo9wyBxQAqmJy+JKYFxTDIMJT/o39
awuj8REZSzUG7ch2FkMSfg1Bl+J1d5+wcejvxj5ADgMs7BK5BIyFP30yLk/nvMDw
BSyneSFqda9G67LgMnme3O+3qWxVBwfl++iu+wXmEuNlo9xPxG7Ba9f3MFIDl7AD
SbA14pXXaarH1m3nBVs54O+9aYTUg+fNF1Av4cw3v7+2DcmzZzLqyrMARKGJygj4
4ej3TuhOTYonOhmBWF2hcNS6Mx1ZM7Fqsud36dmeRGcsBKkx5YipJt31AXNU2SAo
2RBaMFwDcZZGb96BuN/jiVWuvsJ/QL5lVa2iFkmiwVusGGJniRkrACfmIzfW8zAG
LLms+5LMBpHWqmXt3i/TteCYkiQxcdsnitj8LAkUmE0K5yT671EAxUWn3+4lHgbn
poOGpTWcPZnOGsvbdpkma3POYTIpw1FlOvtCE7y6gh9oqNaxqYSQ/Ap76wXXsz7f
qljXfXbd8is06wSmf69+jSz3ZrhV27Jzrm8WUGfFFEs=
`protect END_PROTECTED
