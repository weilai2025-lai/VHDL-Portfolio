`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3/g/29tph18M4sO4AwCcAi+ep45BlybaCo9T1V8rtS1VhjFHnKkTEXjFWyuaybk
six3M/SR2x0u8jdNiiV7pt4aOv3IHgSzKf5/iCicuycZEufgPFytR7HkuOdQaUQr
5WELo8exUHr8aR7/54bnOAYvaLLO+kVOtTEJ9lH9hq4ao9fzXs8x8nSlPsw7zjX1
JqRUNleiX6LrohCobY1f+p+99/z7K9jSSEJDgzyhHF/frjmB/eJj2gcKcjAkIHx3
4ngAfP2MxLs2/H3+mzJpQF8r8teR607Piz1st9+CX+WY8mN4B31xRjTKJWd31uZg
IwYw92hBWkJb4RPBhBw2g3CRfMTte8VX/T9TiG+FNe+Hq9REfhqU+O+Xf51iJi6j
GJlmgkcdgHf0PKOSRWuLI4B8VS/epbKpfuu72QVO24wsycniQJUA4p/TLPm+i9oA
LWR9dVeDxpNSBidUrm8XFFkQh42br0XNKpzYWdOCuNQWucTo3VI21U10vLvV9vU8
kFqOkZRriBcObnG0F+tDnEsUrJBYIDjk5doxnkQTEKeF73dbfl/VXSQ7pRNBfPQ2
LfKVUm417gnVbu5C912IKXu7qdyvSziXMEuQJ2nRKG69ukxbFzy2m0u7IwYIHgEs
1vqeY+qavfG/8UQatXWTk3numXm+dyxzcbEgRjAU49bbneSHT+P1RZMb/7mww+Sq
47F7GCNhuID6U6U+eEAIau1Xd8IQ634vgULQ4r2LauMLZvZAZrj7MUtzmA/zqcMB
0JORLVD7A3NAtUD4k9wwqKN+IU3xXN5k+cvnQcEKoE8iCTB9g6BPz1bYgPgs4Ttk
xXGDG43rZGmtqFXecloZ8IZghTXQBFGGJEhTxs7kiYwWKHDDJS7CrfsMyCibupbC
rjS0SoO4Q1exX3+FOqO+DaH3frtqZqjsbeF2k1ZGEtNh8oyGesciQ9RO8WY8sCT/
YXpTjo43lxklVGYGPNqzj8BacUH8jIZpSf1HLv5rER/ZX5hQUHxG75wSKQN5c5x7
/VR7QPbBPd2Iw1+JX91BTvTTJ+4yu5RTRxY8CASEQl0=
`protect END_PROTECTED
