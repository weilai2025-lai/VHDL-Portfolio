`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9jvnVnfowkeE8XXNNCuVUAzS2fGF4BtlhAm26OsoEtuV4FofmLJQKdWnIBwGTsP
LcOnK3AFC1H5HPyxs/0ar40H+XU78QPLWeYcfdsKKKrTc7gRx2ovcepXfbHSuMUf
FW2dcDIvNoALR8PX7mqhLyOqgMACc0RmHcM2JsqeawVSBPbuSXklhca0oTdsVaG0
Dybos70q382fpdjWEUC5DIN0bPj344xMOPjmCwWJRmbxr5GiALyiY0ZyXS1399ru
641qZx+4FDoWnQaIyAiFGn7OihiWJH+SCTcQoJS3AS6A/LZva5afFx53S9mIORoc
FnoldJC5/nn0Zd6AOTGRJUhHwS346eAmFEHnZZPo4/SkS3fbSSXoFLlkz4vfcS3s
OjzMBPNGeAWy9R5CDRejZq/GVztxUkG7gNZbvCtTSbvd3bs+/ZivpSe9RfIg2v1N
3Ecjs+8D2dBwiKtHDw8x3kGYMJ2t1JombrCDcBL6RdcC7TVMjM4JUtqImcLs9sOb
FJbG6rUyPghHFS61N3Nk1N8xV0a/WdL4sB5Y2qicbI6FJY0GAxqNAtvV/39qYGuT
IFjedZzVV86LUWgTGM7oRSC3yTxc/mXmppT2bgjgKTFqw+aCC3P00NuUntIQntzU
3dUkTh3uRTa0rXF1kcQD7PUJmcYR/uNyrzlUEaAj+rsYvujUJJzvvNqayNIa9jAd
j0EBYL9HNtqxj0CWfx0drCMws5+vkIMh5Gzt91N+FWpa1NQT/DPo3ths3GJIulK/
/tEPofLTpD7QrjKweyftVrfGYIH44ViHtEMI7XOjAS43SiojwjOGwCXb4bKik5Bn
`protect END_PROTECTED
