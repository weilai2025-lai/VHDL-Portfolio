`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6S5Cty8UooDlXptOWBYAbDNu5Q1+FyFEdkB13SrTJZ43I1We9a+lGfSge0oCto55
wCBD+p2Qq6xSMEHPrCUGUiliudEFfUtaUYO5Rj9g7sRkOJ/pi7c/+jTuQ70D+ioS
qdItFxPJ/OW1wjfyHE8rEipbi1RFDq94AXk2f+Db5p62MR7KbpEiX+HfAfDXphrG
OmzDjnZM8bOXZkTjs8iRoCYUQub3KgpKm88BLfw61i2ZInRYqGikMYjc4624pnZU
k8abzql8O8cFh89v7BzRQi+BguNRAoR3ZaZKJwnmvzVz7do9NSmWBYvZIlrxtHsg
xCs0GZeuS6vOgnA8g3aOhTaxGMNrr7Rn92dkUCGmfNpNZwzegmineDmFnuGJJeqt
/yCf0XAqMJBTsLiAQ1H0Uq+WI9EHJCdKumlkvk+gqsXqD2EPFpctDP6v8CzfqjCB
VQinny47z4gXwS/MirWT5g1aG87R1zYIiBtLS49nu14H6J7xt/oZVNgvYr39mkWu
KIAZynIfp8BrmOeL9jGlQTj6tGZKfhIdOg4LkZUUQt+PUxA0zHPePHYF+z9S70Wl
bx2+JlFEUz8GLwc9tgMBuqPQmpfDBVItWKuXfEO33mxkskzUMN6ZEeFFjZDqA6hk
c0qM/zEY/IEpzYg9h5hD7HMT7cJ1Oo1AIUi2O8km+SdTmLiokmJHJjLrdOLKpeY9
8Sn8YNft+QJxbMRhD97DQewNsvfYheH4x6HKegEuKJPivG3fds+gdusq2J3z4n02
QW6YgEb+PWJYgnZchMxnRg==
`protect END_PROTECTED
