`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6e6LwEADzqVx+8t3grEYPZYO+rK5SMTp9lnfnL0P0wPG2B63e72mIpOajrNT5rpD
iJpOBVvbMnTMxcKCdMg4qnp7LJ2YtRS4JVu86b/cLidIkSKTsMmJErj5Z8vWBd4u
2DnB/0/9tFjbHAX+tIoO9hHT1K2CpUWf3M6pDwYU2ozvC0irsFqiNh3ZoU7k8WO2
cXSg+hODR8Bzx+MgKMet+yZBWO2AihBXVil/8v4ita1SclGYh79fYj2J+2c2xBxj
OsdESGyp7vIu0tV1rOF/eYqEBfQlz/o8hQgbcfFcvRSZ/vJjk16nIPI+qJ8QntW6
z3FkO3j2nMOoAiNp+TgJOgmllX78dRKJJWw5+IZsihIevHQML0KEzq1TaRMBIZFC
esawUU8AuBLsbvD0ShqMOmrjfCDcAq3krERkAPRY4o1zHPcZEdDvjQZIF3SKuJhz
OvDOkwPZCjL5ig/kty0eVTqi6uq4e541xWBSZXgRG5PU9S8sk0BF4HmoVxAaIzzE
nQY73Afjnl8Yr2Qt4s8CXTCsrSKw9+J8hWnGfvTbzvbazQzUW8jbwknjHMX4a0OS
30aD4DenKHTv39i1pFu67q8z6CcZ2CWCUhPj13CATIiBKG4iNZxeQfV4i/PcvYg+
C72AvFzLzlv01i5+xyTchxb+BG561oNJrNRXmI12wIJwbfO5Ip4yH9Xj/f0pUIQo
2naMgcJhzBH6eXLR6QZUl6erRh3Hhhe7/P2CaB8S+L/ijb2nV47Y+R0kcJ+RDY3f
0zbzaPTEodlyj9+pKpEwOywy+mw/mN3Lfec97Et5o1uTMN9AnB797nI76HE99ISI
/MicGuigJ6xLwHHiKL2tEvrP6k42shWb/ny42wCO/YO1czoP6La8YqTQ7EKWUkOt
b+M6ElW+SVG/pXl7SWP7v+5oaQ5V01ihA06+Ij8fSv24lNVAJlfxr5dx04kpNK5h
oxSLf6SeqVsMBEbX5Wo+hasCSx5bGIQ9qmV2QzkKaFZ3iwWxpdti0bZIu9beIYYF
0q9A58Z0J2+6P3UKzRWPEhekOr09S9TNAmZLkZZL33y45MHO1QJ7/Gt7UJ3fkyE7
K+18qzerMna9/xMFuO1tdqOXCkTLRfpJBzB/MvZJ6ZLxkKFvx5guQoLeibCN/PQ4
0elhOYbHvt7uUPcrPGcVouIAot32bC5u1F80WYQPva0/9GrQAjiT2+QKH22ZyISj
Sx7fn9+fc8a4Z610w18BEzYNEBpWA90pM1xswwPR76p3WtjGgWBlHLWbGdxlE8M7
AKgVqCVhfilwJ6llFcBG/g==
`protect END_PROTECTED
