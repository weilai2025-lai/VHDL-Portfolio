`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgLFyYQ8MzO6ez2KHlPkl02Aj8DiIZGZv/iwYeuJK1rfDtR6TATYPmOPyjSwi19M
Q/xo96OvEQ0T3c9k7h670N7nM0X7UfpLPwCL+0zS/kccCBCQmh0NwciTt8OwJ2d3
1s2Oc876mH8GTS+TXRznMbCLC8+vkbGVpQ3e0sAkSpL0Y8+0GYKRxsIbI/a+7fp7
KXli284ODJbTS9JIVpOMv+HELIY9xGTYvAOtCeWh1OJTDOV+aZOXg1HQ5C4ieZCR
lDdc6ZgDSyOLYcYFF8n/sVRJhQTDTsdEyqFMgIPRomuWW/iXu52796y3LHJuUyzh
lT760r3P7O8MWEk6hUVNlaLEQojyctgFyCM2UqoTgEPibhG1CV7Io0wyhjsAA6XP
KzBLDlx5QzoJK6YZYVWIOfFQIDa0CHB9WE4ax4/LtefrNcHfJUNJ/DUp2OBDiOkW
TuPm+Li9ADPF2u8YICm9OcHeyVodKCaPtaVzADPPSB3md3GcFIUwY/hKs+qdc49i
4F/X31W+NMgxqVXULciZGR03lh3T+N8AALa71ATOBVE/tz8AFAdzJVChcSehNPtL
eLGKlcfF9AOxTE8F43bDCEgdjOreLX9GvDyTfd7v9u8zjIsNxCKaHOXRCGVy7yBO
AVRkDXZ+AxxpFTE65/B7iEQsKwyvRK5Gt3i+8Ao7BvYG8JtN+iqzYJsKbVo+/GZh
HdX7jKfG6Q/YRI+peAUU4BJRq/KoA6szC1auLicvfs6Rud3dMCJyWEedxwJk+ah3
Ic5T5c1LaYrwGaNRPGsARIComh4dTiFWaOgW4aLZhZYnS2Zz/x5xOIqByTueG5r8
UWbRSQezlrN0JUt37Ov0tTeO1mAIlmH6uQF1f23wgQ4T0pwMAR2ijTeyRrzGaTQn
ZNKv2ebJHzn8mUs58JOXS1ddn5KcRGp+xdQGUExyfvi1A8xwppcJZTUpjXBVr23h
yMWN3rpMS1DzaTS43BlNLprmQCjzO5wtvZd0/rMs9YAAzS5USZiP8WPbvtTWoEJw
fCWfuRQu9bofq9KPKK9Sv5evo31wCIr0/eaAco1v5bgRABTwSy/28ggif+clGSpZ
lep99EWlWngz3GHmXinv08Gk/KixS9EKzRCAZ42dNv+cV6/zA4FHcDNMdm7yr6x6
A5yyHrAJM+2wfEDQlCvKV1pjO+89DNSucB3PCNXB/cFZpeC9H2JB92uscYqvdN15
q7qtNod2Y0epKP2znj1zziWyINv02zP1X1ldTFV7UxnfknN1+vXUoLEzrbhjJLbJ
M8NNkzn+n0GXJBjk/GEbgC5yrCMXVyA7sdzzfoKaXMelnJxJ/okMgmFjT4DLbXli
Quo2J83ErvyBkkroCIoDe0hPByRdID+WSGkP82sWVpJ/P1qFoQgO+WXaiid8g4Za
k9uAq1/at1iVpFdP2Fvc7z62+mSP5HJ6NPI0Pn6PyWYIPk8jQzOKELJOaylRSgCo
mZEhHDqlJQA4SHIsyxCpfvVbQP/9hBMjtpWH4jeYiTk6fqp3PEn/9VVAARIJqV12
`protect END_PROTECTED
