`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yeWbsPcaTX49NWMt3kixPHrW2K7q1OyoBVHzgfWlsaoh6WwPE2Ju/6vzrfU0gf4i
UAi1bLMakkQ3i0oZWqwPP3ysKL01JOAFHktn/Q5x9X5DCAaXDtK4b8EjPh867iZF
pYCXJEhUUygQTqqd6nrJlQx6p/ueuSteOIt7PtkFKYuMRzsyL9cZ7kzl41+E5hIr
1g0Aj6I2d6DPQFWHClU9eLE3cUej7f71el19LeX/cIOKDbR+exFrKM1OzkptDL/1
UNBYTFNMuNHVOGfOdCke9pxphX7SdlGD97mcwXdG3nPoiWy0nh1HaVzyS9LEAVwo
zYHzgW93hdqzfR2v/cfMku32CwZuwY7RrIFppXq3dHmA3l/bzDIy6af/+kZuhhDT
jbH3/7vs8c1sLz2zWcwaSByb4z9pNEcGateon1ADpncwYK+cEfUP5bLcqO3+znAP
Q68jb2PVC6Ngv5ycRlheKqExQ8Z+BHa36EwEMeYiqo8H0L4FdohdmR9vC69+8k0x
he7YsHlFu3M5XwHNXKqrJFvS5rL32ynbiNLQjdCKNRuawdFHMhYWGVzj0b60hJJu
iL6k5peEDtN2nrc13VXUgjI1McL7CG7nsWiMhWnHUD0d6JNAkcr5AEicTaFNKrMp
`protect END_PROTECTED
