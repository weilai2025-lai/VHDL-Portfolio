`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3beyUbYwWpiZae4HBD2mkVpNrS4gwT7RDOmsz5Z+2YiQ/JaM8KwHpDVHaEy/7xOC
H8Xd4sS+VHJRW48egmjjbo58P8LtzfQ4FxpO8U74HJdeVS2VTcNF5A9IKG+74uxm
+4Z4cA5XmluB6ChIpfDpSw8sAVWaxJKU94Eq0OSnhytvTgBQNkfoZupryh+lS2gl
UrkmJ2qb1JAH7or3m0XhGs3hvDElJcdsU2kciQDlxtWVO6I/glxZA6rYH75bgWq1
pIbdrWLY4rdFfqWUZGMEHVFA1lO6oHDJrF+JvMJpGdrx9NQb5BmnmGffZDjUsAmG
6wbsvxA+24IRCc9f6NDd3R4XLwv3DboaIWiYvY5B8CaPzlz7ZiW7TFXNDHbeVPg7
TZZelyS9iy6IVHzXCVTHhCU3Pu8U0vST/szujTNrpFewmOb+B4Hto0c4wedRfiVx
W4TbRDFcBBYmTYma4qAEFxqzjwU9V0AzY8kekGIfO+R3wrM7nf2wLlc3LfvYcT6F
jzWOuZDo3+V+hT3Ba/stYth0laF1pvIdHNgEf8uBQYHyyyAAae8S/Ogv2WCU4rDU
sfVEvwhK7dE5qhbCYOAmN0t4PQIBhSA4TdQPvyL1QiOcgCPKnf4Q675nwT9LqRJI
1lO0d8BcxvG1v/rSNcNGNlqwlmD/R15kS6ftLi4s9FY8p3YcmAIcKVA/++8r75o9
6KjhMHN5Q01k2oF1sK1FsTb/RWNs/c9Y801Nma9vFgKek6PFgNKeNohAzqZKKPSO
VFm1JaTBfHXtXAJh1HsI25spgpIpUMpWdUlFWoG048DUm/TPfl81ZUwApPcfHGz9
0GL1EPHnEDNlRAKBuK7RLgA5NKK4Vxz6XS5CDI/dEA5nBjCHAHzp8RLLPoZIoRoe
zL4VKEt0k8JswSOqkUa3T4UQsHAmE9WXIfmIDH0oNPQ0yvD4BQzAueU5N1Q5ENqp
PjJc15m0kOfQVcQCqI7rGwiET/PMJt05AGUlf2trM3D5Gh1LaVe/heLl/Y97RrLR
oqAoCAAdV/B5qMkI/yIfxwmbfDBGKofnO+SoCfjl9Z4P8MtKvzxZkSec+BrcMq9+
ptlzlLWJFFV8CbJPoxNWXGhWcmrfOvHSA/TKcOpHua4kAFhLLR0enbNTahTdL/n+
1ISfVW2S593Yvf74nmKZh6yDtEcm82NiwV7WtDbCWmLC+8ZWA0Wfc1f3GKBCD9nl
Bi1VV0lv7VcCg3Znb3NyG/huW0EbxPzlrCD20j2s+1gTVGUizTvsfK7FlZenBts5
zWYED9TVXYlGCrnYtCsprJ8Ub5VTAQqbOvNor8cPaWtaIpLrZGL+EV4BYBjFIYFP
XBwGb1nvMAKHjF0h6YzYE9WQaVMkfQGvK2i9saiQbLbMS+So3Y9mPsikrM3wBd4s
3rO9BUxuMEDDtG28DR2W3g==
`protect END_PROTECTED
