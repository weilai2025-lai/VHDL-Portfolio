`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBkvOiPOZkCqzCqwBBCTT1YSwh7zoTQhS7hpZvy1vFINcJy4Oi5Crg9S49rt2zm+
iaR1HjqdMB6WZCS0RHFNHqjl/ck9Naa4SQm03gAcONIq45CR7xwyEfIxjNHCBCdS
dXqFxLvARe4LQStwJ7fF2cPmNnMgeE1PRSDbEaOEnjsVqVEjEh2HfT+y0YsoTTJS
yjPVVwU0/fVHOYoLSQL39Kp7jZO50xh33tQQAkxVCETo4ny+iiOL5RbFjXb20qBS
/VgdTbfg8FlkzCLsNPMlMM/2dSekEeTdGnz/dHSU836dCVtYx5YG4nqOPjisC01M
UjfNLDaijLTROHuUDmpFmvIHUoxclIouVXU6VNOpFZb3/2F8i91sWQJSlPDz2J7Y
nwVq9kfSmSmk0xo5iG+XrW0O+uO3JzUFs2J0Jmd7v48+o3iINBKy5egRnnKf88du
nflVfZdok6C1f9S+uegjxe99K2cnnsVBwapGl72yViWawNK83hlOkdCamvFFSdTb
N1fQm+G+W3CwdSGEiz/kEK4UgLpTki88Xptc/v2lq0GfXnUCWOuejzx+iUYX0Yuf
E6YHe4jMS9Y34NhXDaGVZ9OTTiz92zVthGNH6sphCe76Cd2QO+GvWoz63CCpWfRB
wj8Ixd4uBLKrgzlFa/QxTc112pbD0aS3PTMLPofI+t1IQqMLvl+6JKhex054NMqO
OMtTGiNwDkA0JNyc/9vOsKZYpw6oZttUvQD2pjeveJqCU+1snhR3NrLSuXx33VDU
onfeGQhgFTchSVyyLB6fldfWTeb/oXurWU0SFzD8VzF2r8O4738mzax/HNVp3Pj5
FhuY+88O+jNiRAprX9CBHVOYtBffvT6MIo3nLrDy4wG59fg9vCAMBmA/7eb4TBtS
/L914y7hFdN2R6C/0fuVTmBWkT4A32AJiEYyYNJw8uTixYJfopkomuGTQ5mIVYJK
qzuLee9tXkBNf8iUN1PfaulLbY6ahcKeFXtGoMBuRHdvh2hZliPNwAXMBa47U85w
ulBxyX4IZC1rZvEF7RGekdj3lZpnNO630WIwOdPORBiBns57L9fsYYtsJrErFKKb
zUS0jNrvAkpaJfa2NzpmIZVF6ImlMSPWQ8HilMAPXZ54kivg8NqVc8kiOIwNo1Ui
P8uZv9+pribLEb7GVBTzMQRq56qF2m4ZmLwFR0j61GrTqwX19chVwELDgXLwfPtB
ZEyXjYFnS2tpWg1txCsXzen6PrQdw3FpwG/c/+7p2DnAuetkEwXbB4rsE9CCEfv+
7q1iuqIFAG+qNkJWrzG3NM+SsE7rKZ64vxbxAGKCvJ4bBRPvqLEGFpJhPN9QAk1A
F0Dc6s4czfJqQNKoS5CUR0g/nkFRlVZOCh6jkfnqnY9zg8fn3zC3shMrHGRzwHj9
prvIjS0LBz/vrlOV9XXClyqAtHLmhkuib0qkMeb0zoRnDTycynrNHevit6RAN3u+
abCgjPjgAIvgvHxrDSfz49lrugtnqzrRJsj8I+xcWbY=
`protect END_PROTECTED
