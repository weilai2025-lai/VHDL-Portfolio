`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBb/HntsbwKJdiHqyFZVtFsLfj8Fsbg/vjiYEH9oejQJqtLk0BFx+YejObfvMlzX
+9TK0VjC++UgPLZBUF/RWjSw9/Pv4Nt38p9xIH9dfpg1Nbg0+39fOpRZdFejW6T7
ZWaavMQt/LHa3KLV9XRQgqZNI2El0vSpkdixZdu3fvHCNuXpsEM+I4dcS64Ny0Wf
ABPrhtGpkx673NZ/Un4AH50GVsBvduBjTNztnIfH2fGpxdG+kQwb+uRvyaE29c2O
fIkYdvmXmOxJyGUSUj7Nr5NIqOhmO8kw9HonqjaameZhhWSw0TSZhaS+VnNQPTk7
gutv3r5SG397vanxkCa1T6LsXgAsJbwiK4p9vdXMQXtWxZP59zK819WVvvFblh3e
SOuZTsawMxEd3Uoahnwd/QYo89rV3WyRonyUI7209J4Sqlng9+ptXWVs2sV9+V2h
iFQk5bDUPErTLLa3XXKVOW7GMLG5QhwGZbNsBmz24ebE1ME38SdQLmEN7ewPtEku
fMHzvz2cKChKBF9YPYFw6GhHmzcmQIeg3v5WlKgwvAc4i8FK6Y8uICzT9LDz/tfq
UjZVNztVRMCvZ2e2VM14K33FyDGSPjr56tqC7GP5oHhP4f4ZvNh7X5wU9K4v45nR
LyDWNTVlnXfK466cGg7CgCqG7C93qEIi/iheacp3L2l9Hf/RGeVIloFBZ6+Drmot
/BRp6vNWx+ggZQ3gsI+a0C4LQykJ8Zmnn+2UjjeTxztNotq7qA1lQYxogTE75JXM
IHW/w8Gak5CGEp9sJ3gXaiy9zSlI4srlpgk1jFo4Znwdsa6uUeFmnE6FsfW5RQ+8
k62nZMiVnXfT7hObD+yTjhPf8mb/7YsXZ0yTMy3QkoM+M6w3TVAIKspSVkFmH51S
spqIoqG8ilzZ+FahJNYTLRBJL7DUJyV8zpLdziMYTpbKazteVqDNqBtK5lmGqv0Q
/rdgR0fFrxveTV/3ceu1+6g3VXKjXQ03i9s9TCv/nI7MoPjwKT0TpFl8809an25g
Zx3ilHpVkMUPuOGE+XhqriQwzfU6ELC7EgcbMABuCrFY70HaS4YGn4XMQHW+30qD
G8g21tCNSxViyNM4y/e3wnFK5m57qydOZmZRRljB6Nd9JtennSlrc5GXxyIkN3nl
s2b82Q7yxuDHjb/laWGmchqQr+3GHsTHE0zfETku5h5Rc34Dq7FzPrg9VNBBzRtw
Y/KUeCJjzHkXgOI043F0m7kimW94FI15H8Ufxv05w8m8dI5/eVXo6eK1rvOjTxEB
mcteXf+qeBLFz45RrZWhgMRdH/32EK5762brvFC1hd9CBIJWG1F/G+3iS9/1yAD8
BddxpZ/S9oCSF/MtSkriOjVlczpfkN3PudFlcWECPa6HeqUWswyGxPAMjyif1vaR
c3J8LkJFtkJxOquWhR452cdqCQXlFsYdzxxiWjFQ7tuGFKk2WIBDU7uIvzwKRe66
SMPfmmosz87l4nti5qO6xEyZQTFJuPmIsRPDq5H+F6SxfXIcfJDl/jzTPQZeJbun
RxfSoNw1+je0885XMsEtDs7jy/PCP/foqEgKZo1K55gpWuovC2W1lwpb0sOqGQS8
aRtC8iVVHreMpjjtq856e/L+uUYP9EBciidpqVA6SZheeRXqh1kWuZNwU0fDc9r0
4oL7V/8wEoTtv5axeGkUzH+BFAnIwEcvkW0CKGJzC/viQmvCEjU1p+c1bmZwqzf+
ON7RytD7Hy4irExIee1CIARn5aFjrdqyQCV4fZeLc/Ce783FTSkOhfwDNq/JG0Fm
kTY+dYnHxPtbFyUlVSM6izEd2Z8jdkhqWqb35huuc++81UmsB8Msh8FuDMRoV59l
5VXaObEHBFFxGCDaznZhfTZHM0MUQXaSVxwwCquPUMCEMm8XE29SO22pyygc42kH
U1JC2CH11pUawFlV8y0fnvNmXTnzygcrHzuDgLHs1AK96iqXBBaE8P8jFgKpXT1U
RdV+onY9RHJsHomtX4w+50zXEPQTvjmJehXOIUda0iY7WUrN8OE9sdfgWRuxjbWL
s+Q1g7QjoCz+i24YC20BNk24U1IjA+cAOmIaOWQp18po2Asc0eY+GWiNEPxEn6zW
PvT5cs340O+oSI0Wj7rQFphLyhXr+L1FT0h7HItdMAj9sX5eVsdUuL8u/fc9CSuI
Ap2RO9sk+/hequDuDVLCrLjGMcTp43e/+7zgU4E6QvjhD0e9Wi1gzXmFHGLKm0NA
rcu5xd/XaGisQ/tkH41EYwN70MF4vk3fofC7d2owS4s3W+pUW0doSibpUcSGTKtm
KQi+zspv8pPbTyjJoiEcYE5YxrYEGtum9J4kAjrHw6JW+8NtEdSrA8fil2tnWxBO
QaN/he2bZhmqnYOwJrVsBnas1qSBvPegRmgNbV8nkmplx1CAyhpRjd45jeOlDQWp
Q9WSdp20DhYTAfHAgJUYAACFeaW5D/5jM+4tB1GRIjemE9yd8shafA677sv4HFkR
V+HGAeNuuIdxCaMpSeEyiQl1CZTVPvawEcOdCgm57hVigUL7R8acXKYrERksFEvY
of/jNrwoY6nzGOCJ1BvakCczhJbHrqCmMn3QftYoNzTQD7ydgCvj/dw/s8UnjnL9
BNzEn9DNtgzrH4Ade680E0BUEqlFc3br91/NHBCmLukmW0dxBwnyTRktWCOcZPFt
eib/gLYjBWqF6KxyhX+MAq1EwOiOyZ0toAfbnfTJ6+QB8lhkMsKCxqoTeD+6j8D7
HUrfERLsYE4AY1y9m4MRkKUVj3XRXZUxkLB9SKHMLgMPY9mQJmYGgsLN7Sqh2haT
ZCwljRD7537fUG+Lv7nZWZvvzyz9Un2CsGQ0ElZAHdgXbvyb2kazXBtbBymRPFH1
EmtpUyxM+BFqqjOZMCX/C4EyziX7tFINfQ56VlaXLQZmjdJPKhbtyx1DACYBZnwd
/o8xsWnzoT2BVgMZleuUxDTR6SnmAruhLJligCw65FvVsGsGxWwKvWuErq0nY82F
6bzq8ne087o2AoSLL1wt20Sz2o3aEBK1nI9C2mvhQ6BmoCnDbyw50q2VxzX0htLU
iUbX9gx/WFh0q86B9r9eFx9inbxLiVo8Ep+envNa6K67FyD1D5W4J33xeCSAcdiw
DFkWFkkyLlKFV6azHoJzWpMjmvqxZ8iyNkoRbSmYRyK6EcFDJC8wfzdQr6xhz17U
TBZY7mJ51bf90s8+Gq5bI4u496wXeIc8Nb2bs8iPjIXB2kBMeAuldnkufNLYDdl+
ryy1ujYWNusZqXOuBjlphJlFw95X62u3M7O/L61kuxgdJyAW0PJMdNiJio4Si6AE
gGDZ+7oNvlXP45f1Ua4OW2g8ECDLPDWRWESrk/rEM+jdc/VwcNERlnzzm2mLfrRy
/x3Qfq4vgX+07BYKpohOIZAUFdPbZ56qCTbl+xe6eYjGRBJoVlTPhaC9Qet418UH
/RkjbuBXaRk0L2K2n91rHhRTnFh1fF4CDKbYJOos/NmEL08dqafdeXXbylX/0P+l
WjUAJasJDGbramzb+NLG/VBpaYCYlk/NzzjgIppfyiMHy6iU0IbqmKsRXiGNj6Ij
tZEw0r7dLF61yNR3eilTXqR86PzwYMs4jpjgUWTTSArFPOicqhuvqFCYX8ZHPElI
mjwRBHUx9Z3dWD2DtmnSr9YCRbFfcbQ3+/V6PzThQNWS6nBOGMGlk8NSUOzfU2Iv
9vuizmtaGxsrPRZ+AOPvEp0l7hHKek9EZmY6zEsu+Btzb5wGPrvfRxucT6Cy+rlE
Mu97TdHZwLnpkGfw2uMbBZi3vHnb4sx++mf4ERPf432sAANCnyWrUYVwOnGfikng
sQA5MEiJpTYUX/300mkSB022Ufu6Y5RtutyuF3uDpTAuy8U1SDQPq5ZtaKPSOz4z
n0mnThifapIWXJzKcjAoTEkv6G57tK1Ft+N1P0GCrldzjP+CkGWZ3PmBEuh6QJsQ
aHv2G4S2lTcoyzFgvVepL8gqNSLGwnrNPMfbxOstx8Xh+yPZu1KuI24idDNyZrHF
qOrXL5NhwXfC+ZUUonDvD3X0KR3JTtzQI+piiGoTESbmfQHVOgMdv6PETbSDfD6j
DtcsJMl7E0bt1WK8UiPc2tgN88jEf6iXbtFkILj1WvrxyT26dpdSH7RTFxmgFe2S
bfjJghhXIEJzxb20J4utlF7AvTMF3S5i49lIj/U3+RCmcRdLTDYjn3VHykFMYZCr
5lKNAT4BjeajpVZIaH9cNpGyPB27+culpgLcgXigX0oIlPr+Qdd/NJlVCfVvAx85
yngC3Y0zpown3IFxAdvmnwwvBuxN25Ni0yOifGHaqeRAoz/yBoQZFYcMWeBB5pDD
xgq36yJEx+5V56/h7Am1KXf16xrWptyWA4iw+kueyzLuxmPW1515+b8+WkX/ofEP
FUFr6Eb/tafnuOj0hmPkZ4HFcZGF1bmKg6LNEqFnk0s82W6PLjxWHX6goZHRUgPh
7/w9TjQWfkudn4eEevFuWilt+SGsucaK+RiYkQ7nqWojIGxjOZqLNl6ug0938Erx
e4/hqAHlM94NQr5FkQdngciTwGCCn3VBjYSyGGlF1VlM7YNRq757Xc1/An6WiVYG
aV5hkhyvLbtGH7cQ0pnZUUzkXWZiDZRXqaDq8zzQ2dKFyQ5qPJXsQFHX44qgs+b+
UNm5RuP+v4QG/Rx1NnTxdGXKSdkxd/ndrYXIf6zqzCH2bSzZv8Quuc3hObGtnB4p
FMBFPxJ9+HqTaJN1acmrcxSHi2iuGurJ2gXXHY12OMCTV1QOOMjOCRFFa+RqACbF
ZUZMDwcOMnzFwR7w9+LwYbSobFxKJmwFjEH7KqZ5uBxmHs57vNVUrdqviS7RTQQQ
dQku/EC1XgWxS3Xij4tRkQ/e/l9fImNzu3UjRkFFPZMwD5Yb+t+h6JchCa9oQzu+
0ayZLDBa+FKhfXnUbphqb/HZJvouBdHOYqcXMABLDVSkHkzlTSeRkLpKvjGWu0H6
nlPgmTKdecFAnTLfGalwGacUy5OYs0PqUnAHhxLnc6ykgzvivTHng7D8GYVTgbHO
ayTqKNckCybJH7HXKOYJgEKGpDEIYcFxxQO53IpcA1SV11mSbpPMZY94pSF7bn5p
K/xzV9YS8fcz3UPYmfAYuf3viydLGr/9HoAVnr96Fu36aJMh9FNpx9KLVp41uS5u
mjMivT5YrLfsFI+r9bpMElNLvzPQ+iuZ3n8ykUASfurU36s7aaL7zeAfrelZBW3n
epSnf0gh6Ns+QgsdrfyUY2r1rMN5droxZ3yV9PNDkXXHOH+OHsp2US4QO9T9rXPQ
VOjcNzO9dhqQ+Le1OROhXe8/Q7zo7fmV+BG9LwCqdQGuVY7hHDoz5ENQC+9ghtOO
zoW1s15d0SUg/SMEhGPOK57vRtWKI+2kg0G6y5V72phpq2Pm2EQucaqEkg+lqduM
I1U4Q6AqC2i6v5vcypmu82uWCSz3eLB2LT2CW3YeIYO+4Gb4VWxyGuTKYMNk/U+O
PS0QnlvgpFeemCOlcRq2oMmD2s2i8tv5RU64Jy9mQAUWIYAlL8OVpy1KTpd7Bsm0
gnrFHDtOi1SMQ3O+AVq4ZH7Ih+cN7ZfAgLmKlhFPveoODNVezbUTaACh1vTqOITs
hyMSf8Rx5Ir5jBFv2iTpAAHjuozWHdbfpUzBrsPSKnWRS8i75XjBDnCA4n0JqnMB
U7S8bp6bEQFwREL6pDUELtVlS/lQ51OjXP8/zX2CBcmg6pNSa0u/Y/Fjg+dOzZBy
83BtZCw3kYUgvhX9xJQvC2Z2ouAXNy3BuI8/ouGo2CksgetUd/b4qJ40F82uIBon
rUwjBmxcS3yEBTNdGxTYNO4Gkodg3gsL0tYWqAR0e0I6L6scCUJysoGyyW8UrRqp
mtO6EUMm4VifiyX6V5FW2AXj5QunvM2dKhlQ3Pi2mujut1DWpN3w6Zz9R/gYU4x8
WQq06G8MbVQFanJNK9o8GSlLPtinfbehvgDuboj6NY0Y7l52qFOfXcw5JSG3z/JK
MK3vuEn1GSFWnUTGGc16ywIv0a7AkR0x9ZNRQrX9tE5oItxB2mylhWe/ebXptQCb
6hLzbz7ERhydEXw44hqfFN60ZUQPjRehA+JqSPwYFYLAK4HVvah8qEehicQ0vJRY
2yicu9hdjyHtNb+RcTRVqNrwP/zBq9aPwHixYjLAolJEBBF1EHOfczzddviNXqrk
ynCJSDYay04Q9J1PbW9kmR75kerZ1gLJWKFLDaWLmWP25OnrQGIoidy0QgLSikNv
1/97GtzAOAcDT19NudXFy1qXgxdoLXM8TxdF10vlxSoRl2EWuxJSrCB21MPpmrT9
aTof3O6Vm1T45Ufvw99RIw0I+gVMeESKhoSH4zy8WXq//DXsSY9e/cwXNejHAvOx
LrDpJ/p4Mlp4fgoEPQriVY1u55LJTDp0/Ap1/afO+UicoxrZvCUasefaUVkFAkwG
kSDR5S9S2MXzbqJUF8bDqpUeQ2b2BkUPGoj5kqOlv7ngDxxqdgQJ+FLOeBxB59A5
kSn1WU/xRzBlIUcIA0VD0JCe5Hh9LUp7vJPSzAObljFsY6xR5AcHPhtvQmVH1NNo
2Qrq1FXxdzpFMuprxh9N1gTEp07FZPBu6fwRhakeP8L5Wse/wjeo1EmErvJwpuc5
wCZ7V04jpi+EkAt2DgB9g5YTh3Pgl8sXnilZG6+CoWq2PHZFKeOjzs3fWvWhKJvE
0n9B4t4f8YLF59sh6ApfYgmetO0sopv1hZ61NgysDhmZZq+MBtIPpYue+0bS6gdZ
VB8V/ZUGUKL7GMgVJ2EsUXAWXaZ0+vQvsHZEk4SfocvDD2yPyHtZj+aZN4Jj3BXw
YoK0LuRqckrTCWaA0zvZcBmVFAlqms2mYm+Y7+oweLMR4EY389dDVP6p2uGbgheZ
tL/UxyiQeJdMM2WLQ2sXyO4nMV7ibrRkGzR8lDTTiGy/xpF6ccWH3tocG5ymDQUo
lM7jeJY/036nu4uFJwuzpWhNq9mKNGRgOWgsAFhPBdmyqvb2zUA9Xc/Dd4HCW1LI
zq9bQwipSMOlZ2PUeRGRazoIzi86e9B5j6xecYGddYOGUgsB1zNS60+y9JsZ8K9T
kv3N3hKeycSzSciVyKaZx27CHaH7t72MOOow+Cxc7q/xDi+3lXdNKMlCXwXQ3/jt
+ewKiYIGn8lqXpczM7EeESnyNhwIK5vkuVDCrW9QcOuIYX+aE2rfD84uKyiMUV2+
Yk/4iRmtLk47l5hBWNF4VScl44uEqUxlavXi/vVYBHeqNTP8ACOM8M2C38JsFuuB
l9zV/T9RVnQbBcIOIBCU/+sTzsI6ioteD9CgU11NRdd2jfGlu6tfg32Mfy6jkMSk
V5MnjMSCOInS/JuZ8tpJpDRBtspQPQlw0lj56yXZea6C2kOAs5q60X2riQvukMcu
rxKNfhGwN41DThiklq91D713PUu6ZoaKEpI887mO9U2FzN5n/PX6mgsFET5sbbon
+IvptXyDhQleWSYjIrXglEe3zxtrUny4pl+Ug1iAn4Y1A1GD0KIJSfBj0hRO27og
0OQUPtmUU5duLepH2xQMQuxdtJIsYJeDk4JRKXhlRWOBC7cHJJ1uNMWCD0BsfCes
cbdRqXYmpiQf3hHggbzouWZID+rP+HgxUkeLEPBMpNGXff0k5PE9w3Mbsm6iCK2Z
wg41gb9UbFqboJqQl+y4LaBz/4yuANwprg4B+Whq2hZkk/rD8t+fp6tYLFuJrpHl
3hA0L2SHFIMmdlHdQ0WL8pUM7Dg7eBbhdkbFWH5M+OBDIgOOtHdparyRBIyTqQJj
t7i1Fz/D0o7iHp4kXDFnOCfnPiC9+fHOU/Z4MV1A2N5RTEtgEFOSa9a4mYDXLNBL
M1izUf1vWCwRqUO2hZOxrRRVYFieaEIKNBy7QCbuc6F/QsnvLO63tM6cBbaxPlOU
uWst0pMgs3Wgy7d2f1FYtA6BUU+bnH3doqc/IVTFPExeDzOcJL5A7SCh2Ht4UWa9
W/DC34AGhtUYtgAHToXwcM9u0m1TFatjyPzQ9XkAdVyu1puYKnNBad2F6Z3r3V3+
CrvnRKBlrvDfDXw3OG500aN4m2tUrUCerxEG2VBbCm3EPtLpQNoWbgktM+dUpND0
/BSvMyzkrSDIwLi1cxcWsf+N/Pjk0UnWOHUMEJk7SdY5e/K6Y0X/P6OnvMl5FirO
lVZNx3gr/k5/AthL37ulBn0zt91/D93tzROpoWwRfxA55UsqaiFu3EGwFtu5U27S
UXM+lJET1CdNTyF63ohdpbSCVH4J51rUpMhfd1Z9x27pYlE1zWNIu4GzPUxaYnBq
Vo4GqQNkb/4pCrC29hpEQ89EGHiOC4k28oaIwjknZ6Gleikwh34ludU8LHjEUrTl
nQg9ovNv6bqB3E+ECAMc7bZbD7cn4vSY9B6tpvgsPN+mG3xHfhXPtRLf28FWvYrD
dD+QeupBjxsQ0seVutDja2h4HlVE/vi9DpytH6XZ7LBMRbjShFhlsJTUV0TTQbPA
s+RJOF/hjRkEqWpC9SUzyWYv7AC8YPGWJm0h7rI4UwtYo5ckh0M+fv0lhLS0allB
A/o1BSNxSCFl8RdAwY/+6vn2YUAsORipPfeN4HMvR7f2+rRGg6nHr+gxKSOp1sgY
+C++pQkCgXAmdB0AgbxdevwAZxLzCzJ01hQahgAaJfjdjhhf5UvryWzzbqNXHgwF
quwvHBYvCDuKxIkSPNR3WtECwXDGT/w/A+o1jR+4nEcmMV/3omjSJDx845IntjLP
9G9k5R6/gUrEi+pqHEXJWzxoDlJLQYZIsDRLeIhBCk0EkSKR464UozSs+I81tpmD
NqE04QpADi4FisXDQzVInT6/JQ5QEvRRjAyQvn/qeFwWEc6UWx6SEvLjGcDiTzIF
A8wTt8+ySnqOb8iG0oxnNLHwHAg/ChAVOpLR/rk295yi4A2Hp+ZCcznj7BGOs9RW
6wk7prnwE1+pLkNK+ZsF53U2lArfP9XAuoKobBCuIhswwT2oPkT0wYoVgY+PPNAj
I4fNr15GrsJJX5XlLgncEw+R++HoBUpE1/N1LikxUE3vTwm09iPnEwT6nSl4UZU+
wDbkx1blJSej0LzeRhzTvYACko4Xlew95pSLHih/NPlwR8rmeXFUnUB+mzlVPfUT
9z1zRYU0Hr3CIzc55830QmMRfvfk9uMnS5etG3lnrGSi7vaU0IvjlxJSXevyK0Iu
bxWG1XhQgIVeTGg0USadPlPFR918rNm44uf2mDWBueo7X4L6M6/lZ7XjN+8QpMco
89sxqPJhLT9SMV0Iba0UPyyJpGOVh6carkKgtgW2u2rZvT4ZZFwoEVmrUv2xFBH+
K2nJ61AK0wTmKJv/3ZIXHbeULG5EIf8BhZxiroeVmPO9a3+JZ9ZvLWLXvVmhUFZU
H9KvRQs3YEOUrLrT9bZC+9IwGwPfkypBx3UQ7pjvg7B6JsMMkmWoqECKbbiu6X6Z
q7G28sDTU/GCnUI0N78upaJ/vAbLrQeVG8oSTe7bTMmrOBYivv+ZWNE+BE0PxCD+
Me+7FM/8BxNCyYDuNfj7fYxh9Gf9H/AfDN20O+GSwhXE5HBziRYE6JPL8nDNROqw
HiTauZvwmi6/MU7nENwVJoJBDhParPz5jbdD1IurKrncjMJt/Woz/tvQZTqkqK+o
XyDuGbgyZDAb/HkUPxI/+xqVLCvrejiIt0aGdnLXlDK7CFURJL/ZmpfBwFZrgH+a
0oBYQMYhyA1GNnTxpjO72T2Vsk4WqUzh4RewRsXs/NtSsia6nrK6JuF1s9gkCawM
QKooZKzrD17/bCnMromgMTS2c14jscLvEWGgqOWSnte0Jh5ODVv3jGJI7ik6WS1F
qZUONOcWAT88A6yq79WvOkcSqLg/8GMSxdOq9F7A8FOn/SkQUY7Rz+iD0pdJccL1
YAQtUW+0K6RiYK7JpWZaPhzRH7DRlL+E/9l/2o51GscTrOjg1maq8zgM4b+6jb/P
9d777EhrRQwkWiIjA1JvzYa3NAeQv7hNP+9hy+bFybwCedo3h0ALL+TMea6pDIEk
MW+p1EMLffUDIARSteR37yJmKd4do5HVUdtRCIKXnsidBtWkh3g6ZBcFbMyfHUan
Rg0thD52K8pTX+jgM5I31/3ZohmiDAPaoLzX+S+2/kA/xTm3mtRqL7BJXdOVPdYi
4J0bAGJpMf2FDT7Al+6L+CSSW+KkWeGbUKSlBEcSCh1kFi5mfPOeZ+Z4mYXEicQq
H6cmhJ5MTKGKyyT5QJE8tE32HmBdbLOCp9MvRUOHbOKa30fhxkV9GtDgk1Frh+Ui
mNQlzlj/zc+KYij/o7cJHKRdxJ0K5QwhOXFYkGQMLKSoATZBg7fY32zn7dMvUoan
k+0CBLwVZ+BH6P36GMlEtTxzthdMJyL1vvV1PYuHxzZd4x6WpEEKDffd3l50ITKo
5ElnjDg5Y80ZHuWHmS359rWPt+7t4u0b3XLhfc5kyIm+EPDbY/i71+bqYU9G+Zkf
tXBUgkvFnrK+h/Bq3MKhNqXETYgbotZJ+zcRS1RzKUje7wurIJgeB9B/VF2vOHzl
VCr1NuOSdwHkscUoQmSaE1LOlfVIxpJncF/4VGYJXMvG9+I+MsK8Z/mHFKyaA0cB
Afnl7e++WFzl0nax9XByE4Ve8LdG8iBPuFMy0TEvgOCvQmw0/NChxTkqi9hoNNpm
mt/jtp0RG5YvGrXIBCvwd3EgW4PovO5+/DRSdSMFOZTtUdH38hhmOudE2C9wJsWo
I9ILHRgWln4pX62fZ7CzUVLX2f8R9f4RELXoARUbzb+yTdJqM/VKiitIEgDP47MN
Qa1XhckOwt2F08FmZIp9xZb0tamWcqqyAhoOj4RSgQvNhEwE2mTSDYs6PlnLeWD0
nBGS4usKBwGWzb61XbDAbHcL4IDqv4+XjZhNPEoVMeQ2U3vMawAYZW/RR7Zk/Wl1
0KoXxUokHjAiR9MVl8ZGkou1JXPrW7IlLtH7XH1ALg1utq9CQPQVq+JQWgfHT59U
vHytyaLlL/TWgBH86KpN6MpaSmY2rafaH2uWaMMYft2H4hVZCUZlKV8FEOschczx
4nvBl7Zd//odjH79gXmgMWZsxEVg8+E5bPawfSg4ZQR8kDMqmb0CCjF4pVypbI67
B1rDn3zG+ipTU5BltUn6UhXOxUWLtzuUB/uxdlYy6RddsIf1oACy9IrLCSdjraBc
CZEoXsSSK3AAOofxwjEqsaBwXyTX+XIHieRnspowcwxzMJ1MxUzTc6+GzW6das/q
tWw0xYg8+4hRuY3kZzo47plOb1/Auw74PnjTSNZf8thZdBXTne8MCmDixlsG9zBq
lr+FiUYDpaJLlBWES7pUrMtSWQ5e0P6f577YXEfrsDZSw9o8tA32r49vjRIzLLl/
OCNoYTctz/mYcK6IgC7WxF21ivHqRUQ6ycbYrkxhCMlX0gS6AveRE3sUUqU1lKfy
wjRotuW+rsUZPGN6Jsscusq4O+kjStfbwM92xsXMETLBIaoURJYldG7Nl2Mv0bXJ
2N/BgQ4PYMFH9uvcP4oGtI8AinXI/qxic1Ny/SiNs70zQnGBrpVFWvmLS3kkI/0j
ULLgtvCnZUQwPwBLqA59ouCRsY+7yADuvHI2JzMcasIlfXMSdyinRdipluSsyJlx
S47rUsESq8OZ9iFT8MN5LMPIQIIGtrEKsx7Pqn0HJVUFb4RsUBDHiOaNpF+6lmf1
/mZCuCVhMlqzz3saPcV56Z2n/OM38ugD986hw3uiurifQW0oAboMHhIeZLroLjVT
YylCDkuw+eLoP7tv09dUIVk2RtZdKiIkimzYnO8/doe5VHZVSW0IxgFZXfo8SYcn
GmyHnt+a7K65jb86wUOzEK8GlHX6cOveNNYDfLFKTKT9DzujcLCokZU8sChLU3Ly
HwxN1aE04/H7ytiwZTiCKBo3Co0rEK6zaPfLr8T2uMmYCNL4RdjMn+YNHxKZh+Ob
+SrWyH/0gFu82yLNe8VWpl4u75DqKWyCGRuCfkcbPOnnfWeEfv77WXV92JhiyzNb
IZiB1MXAmPKxhv0+gfiAe0FZYnwMdjYbHH04TpvzZimqNQtZPMB8wz3DziHeT//3
9rbZ2oHveHv11QjzD/Y/Mx6Dt2mY7RCUq20sazIAeDxVfHfT0tZRvT1ycOegxq2v
mwPoTMKfJxP/5ZaoEJrO3qiW77POx3lZjM/djd5ohiFzM+HI/gKvP+WcNUHqx96L
0p8Q1E2p6nKbBHuUFpLjvqr/ym6eNwIjwAe+17GNI9fTJy3qCK2z93OTyLPrJGHM
8HYRidT0QvOIoF3BhYCTG0Li2wnMlR+E33/HjCNdJ0FHAcfxxDgCfIloMxG6GQ7h
j8vPbbLbmfnA7b7Kt0dFnGrlKJF4vANyiUyfLvGve1iK+OE+unDwTkH1GBlcP95k
UYbesukavM433SOf9iCoUIU6bmyXaXY4kNsvXyl6mETQPe6sH4KOt0Z+0AmeeqHU
VJst1oYTgFXkSGmW9oO6BlbDhHnde25YKd/azjmyBrDTf5iB0uxQMNesXnFqXVPx
ErncJ3kSBaftc8VgTV2pI0T/mjOl/eeFUjG5kmYgzIg5z5ueIqdBpoz5+DwF+SLU
14PmaOjjhSIfAavmvcGCRukQgn81buSETnggPFwW+OOJUKVo7As1QBmNxAJBf5G3
pFPWn/BcaenkDCtUIuzSQPm5Wv6sY3G4IVBIxWMJyRhOt4cSRgbv5iD6ZVcjSN/L
UOlphVMnot8ON/NJgg56LyiPT+diqlKbTGneY+FMrg6bUzgJNzPXgW8OtDHK1763
4s+8MLuEwPK/D+5gt02k9gDsz+LWraXfa9lxA8fJDqU0S5PmeRfmJjt/4qiocx5v
UEo7yZdrC9y2xsWJWrHBBDHjYbsytqoyc9fhXOLhxDLCmDJofsjhXkjQv0SExMHt
3XF2dHfBOMsqmgHkG1wjpFtir3mGYOTGb1JH5CtGb5GoFBmEI3Q57WGbmZSwgVPu
WKiQuLhVRokuTsrLcICq7Hd94yIQ03xhViYLM2yTddYAkuNPOPP+fO7Jd48rEtor
/lxOqzMRx3o1vcFEevkLPzV7cX2u0sD/2uWWOuZjZOLZUtlrLE79g5STsX8E0uPp
NxzyebGBPxmgDCpi6eBJbCuhQmCKsMtpRMyUpkvxicEKQ6Y+IkntWsSNUzbnHv2O
5wn2NTa14LYNXd+YgFDDABQbkjYyp+00IeH/qkUcMO6YqsiM0Kq4cEYhS46KicN3
3LXCkvKNnsFRsL5H9mpW9T86+Utnfbltccm7A2W6w8pWRG2tUYAb8a8LBh0u03v4
n4m5TOvm6Hc0Ao1T/iXO3Q==
`protect END_PROTECTED
