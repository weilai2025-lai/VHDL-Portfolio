`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHWXwG8aepI38d5exB3YFOKOM0Tmk+nD5Pi5gbXRxQ2l5oOU1EPvwy+G5VGd8Cxp
7seeAlP5fBVe/ySTxZq3jaHShy+nP2WP8p0r720ehqKmNHkLl9WxpJp7eiq1h5Jf
344XeCkVIEN9yZZ65QnXVmQ6jW9lykswBk5wLTAT8lvjW6PFq+if4xTrhc8rRtne
Jdu0mkc2e00JKVyA6Dw5YkyhwbOdvTK2nVtCCTn+Mnw2CxTjnKDG08E5bshcAtwF
OkpfxHctr7+jsWuytsGn4dmiYQ1VWi+hOcxupr/HUEKguH5rJuI9Yk3Nq8jvboZD
thrIiJ42AaPr5Dr7+qYhoql0DpZWSYBzzg90wtDytSphYl4veLsGWZAKzy4cLtDI
lQS6OrYxaI4rDUFz5yY/8k6jSjjbf1nFR/l5CmzbVj6NqSVDd4NbwM3GZdC5pkN7
liXTbInKLJitH9XR8m2q+B01b9kdYkRH8k1wWr2CPTtx1x30EghPu1BnngMHch9i
PyyjxAmKib4g3tpMwHYcrCqnI1668DJA0AsWRzVRNNOSK7FmVZzapRx2h4Vvf5Oi
2Z1efC/c1C89vTiN+Cltl2hp6IQuEsTMgpkqWHoIcuo=
`protect END_PROTECTED
