`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iwF4JIxhQrRE5rye9WyO/WYa98pvvDZjBq+gCIBuKjZsORs98IyHf3e8V0Eke76c
/5EAiwZRI4Cw6dsWTt4PKJMwStziPJu5pZSjONDQiwKCfnU/DoPdMIP0QR9z0C6a
WMonNVC20Q7PvnM374GvQEKij6s7tivuJLeA4bwD3rUy0oeB/IN1otQTBmirIKQU
Hl4kkSnX7PkGY2FWVbtnoJmOITso6iOJg8hNwZSZ8Qk0n0o3xAnZogyAaCuq2WK7
ox70G50o67cMF3+VwASWGw==
`protect END_PROTECTED
