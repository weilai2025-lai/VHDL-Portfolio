`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bwa06DUIUR9Y4nBxiVmQv9MuwDUA9+wCtuC5LdMonRpeYR5ttMI8UV2Mz9IfDrnn
NvfqEO22r8Cj7RyUFPCyW4AzGOVj98uE9bRYAyyD6pa/AwSD1qLIEogErb6y6uSG
At351/MtGzF/2TUKP3v+K9fQBcjt1Ta4TBu/P0TWZkatLiAYNOotL8LnUUR+L9UW
QyAesAI7xUvLy1YFf9odYZZ+vvwIOVPS3jOKmkWKBdcj4Ub8fpiivkUebpWDHNQH
pwVtA64CnBja1X1Wuw52/IDLVuaS7FE52+D9Qw1veX6SvNqRMeFAy+vnHD+/DNTK
jWooaOJhBULAyRKDij3uP+14ZeFcAogFzRdriLK6FfG+0zRzuD4UYsaGceHJe1+/
FqrSRHei3HbA2r4QAKDkntWoEfwSUHwYYocDaDn5yf4hzYst4OJAd9bnh6ByjsXs
0jiifK+wdz0GbDvrevK3wTlvjInVBun+fVkmVCLtSix0AevBmPQuoGdIgdLdI4rV
JU5g4rTkBr8Tu5uQRhht3+qvSFPcPv5sJsjR6HfA7CKI7ovmujVRvhzUNblsQbp4
uCzaVqiPqC4uh9zzJM++79imgeIkIy9M7+FQugu2gbNmSxC8LvVWd1H87TC3fyxr
08RNh6oaY6LF8WRsS3FVeYWB5Sg80ezU9M1fppePwJIBFnKT4jTGJxzBmP4QsUbo
B0dui2UVjTIYJRowjsncfxyBpg+M3vnGnFQNjLQdaz6V1Dm9qUVjMHLm3mSEtBNk
9KQEUtH05yy2hYhAy8JvJIzRDAYg2KwcPi8IXfUCqx00+KoBHt0fza7gBWHitzvP
mPCcVtdmdhJ9WS1Yg8Iob1T5Lc4h9SaNXpLx4J8z414=
`protect END_PROTECTED
