`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rfa2j+lk61nZ+RiYxm55oqgGjzv1jIEp/UWbvIi5lx1qGfO/E1clxv9SaxuJYhYF
sC8LpiWpgP4lkXLSerXkUzUWVC8tt6jgeGQ6p9dz1KCe5j8FpximYRiSIvyOUUO4
3ZY9TfNe0G/T2yEtNuGHgUFKD8aQIGJzznD/DecYRizsKVi7usnkiXBw6RpgUZPk
Lr6xxKpINxd34KpRoYuaYNNs2M4JKlqslmKKmNT/bmWKZ+l4aJFTig/5VN9wuXiF
L2/WdpocS9kGbBH66pBx+yxA4Jf8KxXl9govpUP//LMtce3a+6VT8L+YhiQmxQEO
nfMZCKVNew2sXivXAA+/UhbaX9wNQY8tmI6RYBgL1QrUDdo3B2FxMKuHA+f+eVy6
a9p+ki9C1yRJ1hLqTlCFBo6KfWRA+kTanrZ3+E4RxQ1HuT82rZvd6e4yajjKUcuH
`protect END_PROTECTED
