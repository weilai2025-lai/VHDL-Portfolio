library IEEE;
library STD;
use STD.textio.all;
use IEEE.std_logic_textio.all;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.nn_config.all;

entity Weight_Memory is
  generic(
    layerNo       : integer := 1;
    neuronNo      : integer := 5;
    numWeight     : integer := 784;          -- 784 / 30 / 10 其一
    dataWidth     : integer := 16;
    weightFile    : string  := "w_1_15.mif"; -- 只給「模擬」用；合成改用常數，不再讀檔
    addressWidth  : integer := 10;           -- 784:10, 30:5, 10:4
    SIM_READ_FILE : boolean := SIM_READ_FILE -- 模擬讀檔開關
  );
  port(
    clk, wen, ren : in  std_logic;
    wadd          : in  std_logic_vector(addressWidth-1 downto 0);
    radd          : in  std_logic_vector(addressWidth-1 downto 0);
    win           : in  std_logic_vector(dataWidth-1 downto 0);
    wout          : out std_logic_vector(dataWidth-1 downto 0)
  );
end entity;

architecture behavior of Weight_Memory is
  type memory_t is array (0 to numWeight-1) of std_logic_vector(dataWidth-1 downto 0);

begin
  ----------------------------------------------------------------------------
  -- PRETRAINED = true：上電即內建
  ----------------------------------------------------------------------------
  ROM_MODE : if PRETRAINED = true generate
  begin
    --------------------------------------------------------------------------
    -- 模擬分支：讀檔（支援 BIN/HEX），維持你原本習慣
    --------------------------------------------------------------------------
    -- synthesis translate_off
    SIM_GEN : if SIM_READ_FILE generate
      -- true: 每行 16-bit HEX（例如 FC72）；false: 每行 16-bit BIN（0/1 串）
      constant USE_HEX : boolean := false;

      impure function readmem(fname : string) return memory_t is
        file f      : text open read_mode is fname;
        variable l  : line;
        variable mem: memory_t := (others => (others => '0'));
        variable i  : integer := 0;
        variable w  : std_logic_vector(dataWidth-1 downto 0);
      begin
        while (not endfile(f)) and (i < numWeight) loop
          readline(f, l);
          if USE_HEX then
            hread(l, w);
          else
            read(l, w);
          end if;
          mem(i) := w; i := i + 1;
        end loop;
        return mem;
      end function;

      signal mem_rom_sim : memory_t := readmem(weightFile);
      signal q_d         : std_logic_vector(dataWidth-1 downto 0);
    begin
      -- 對齊 1-cycle read：本拍取位址，下拍輸出
      process(clk)
      begin
        if rising_edge(clk) then
          if ren = '1' then
            q_d  <= mem_rom_sim(to_integer(unsigned(radd)));
            wout <= q_d;
          end if;
        end if;
      end process;
    end generate;
    -- synthesis translate_on

    --------------------------------------------------------------------------
    -- 合成分支：用「常數陣列」寫死權重（效果=ROM），不再讀檔、不用任何 IP
    --------------------------------------------------------------------------
    SYN_CONST : if not SIM_READ_FILE generate
      -- 依 layerNo/neuronNo 挑對應的權重內容
      function pick_weights(lno, nno: integer) return memory_t is
        variable m : memory_t := (others => (others => '0'));
      begin
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_0.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 0) then
          m(0) := x"FFDF";
          m(1) := x"FFF0";
          m(2) := x"FFF5";
          m(3) := x"0008";
          m(4) := x"003D";
          m(5) := x"0010";
          m(6) := x"000E";
          m(7) := x"FFF8";
          m(8) := x"000A";
          m(9) := x"FFF0";
          m(10) := x"FFF0";
          m(11) := x"0005";
          m(12) := x"FFF4";
          m(13) := x"001B";
          m(14) := x"FFFF";
          m(15) := x"FFFA";
          m(16) := x"FFD5";
          m(17) := x"FFEF";
          m(18) := x"0015";
          m(19) := x"002D";
          m(20) := x"002F";
          m(21) := x"FFFA";
          m(22) := x"0012";
          m(23) := x"FFEF";
          m(24) := x"FFDE";
          m(25) := x"0017";
          m(26) := x"0029";
          m(27) := x"FFAC";
          m(28) := x"0035";
          m(29) := x"FFE1";
          m(30) := x"0013";
          m(31) := x"0011";
          m(32) := x"000C";
          m(33) := x"0011";
          m(34) := x"000D";
          m(35) := x"001A";
          m(36) := x"002B";
          m(37) := x"0031";
          m(38) := x"FFD6";
          m(39) := x"0000";
          m(40) := x"FFD0";
          m(41) := x"FFFD";
          m(42) := x"FFB8";
          m(43) := x"FF83";
          m(44) := x"0073";
          m(45) := x"0029";
          m(46) := x"FFDD";
          m(47) := x"0019";
          m(48) := x"0015";
          m(49) := x"001D";
          m(50) := x"0005";
          m(51) := x"0025";
          m(52) := x"FFFF";
          m(53) := x"FFEB";
          m(54) := x"FFD3";
          m(55) := x"000B";
          m(56) := x"0016";
          m(57) := x"FFF7";
          m(58) := x"002F";
          m(59) := x"FFF8";
          m(60) := x"FFDE";
          m(61) := x"001C";
          m(62) := x"001D";
          m(63) := x"0007";
          m(64) := x"0037";
          m(65) := x"0017";
          m(66) := x"004F";
          m(67) := x"008C";
          m(68) := x"0135";
          m(69) := x"0131";
          m(70) := x"FEB4";
          m(71) := x"FB01";
          m(72) := x"FD45";
          m(73) := x"FE78";
          m(74) := x"FE97";
          m(75) := x"FF53";
          m(76) := x"FFEA";
          m(77) := x"FFF7";
          m(78) := x"FFE1";
          m(79) := x"0026";
          m(80) := x"0000";
          m(81) := x"0002";
          m(82) := x"001E";
          m(83) := x"FFFF";
          m(84) := x"0032";
          m(85) := x"0000";
          m(86) := x"FFFC";
          m(87) := x"FFC8";
          m(88) := x"0005";
          m(89) := x"FFF1";
          m(90) := x"0009";
          m(91) := x"002E";
          m(92) := x"0084";
          m(93) := x"00A4";
          m(94) := x"01EF";
          m(95) := x"0363";
          m(96) := x"0240";
          m(97) := x"0057";
          m(98) := x"FFAF";
          m(99) := x"FB41";
          m(100) := x"FB9A";
          m(101) := x"FDDF";
          m(102) := x"FDAC";
          m(103) := x"FC5A";
          m(104) := x"FEE8";
          m(105) := x"FFA2";
          m(106) := x"FFF5";
          m(107) := x"FF94";
          m(108) := x"FFCC";
          m(109) := x"FFDF";
          m(110) := x"0092";
          m(111) := x"000F";
          m(112) := x"FFF1";
          m(113) := x"FFEF";
          m(114) := x"0012";
          m(115) := x"001A";
          m(116) := x"0004";
          m(117) := x"FFA7";
          m(118) := x"004D";
          m(119) := x"007E";
          m(120) := x"01A1";
          m(121) := x"0423";
          m(122) := x"05D9";
          m(123) := x"046C";
          m(124) := x"052C";
          m(125) := x"FF5A";
          m(126) := x"FCD0";
          m(127) := x"F9AE";
          m(128) := x"FB86";
          m(129) := x"0197";
          m(130) := x"01E2";
          m(131) := x"FCFA";
          m(132) := x"FC04";
          m(133) := x"FD3B";
          m(134) := x"FE80";
          m(135) := x"FE46";
          m(136) := x"0063";
          m(137) := x"0157";
          m(138) := x"00E4";
          m(139) := x"0055";
          m(140) := x"0023";
          m(141) := x"0007";
          m(142) := x"FFF5";
          m(143) := x"FFF7";
          m(144) := x"FFEE";
          m(145) := x"FF43";
          m(146) := x"FFDE";
          m(147) := x"00ED";
          m(148) := x"01BB";
          m(149) := x"0174";
          m(150) := x"0283";
          m(151) := x"058A";
          m(152) := x"07B5";
          m(153) := x"029A";
          m(154) := x"FCF2";
          m(155) := x"FABA";
          m(156) := x"010D";
          m(157) := x"FF3F";
          m(158) := x"FFF0";
          m(159) := x"0484";
          m(160) := x"02B5";
          m(161) := x"FECA";
          m(162) := x"FE8A";
          m(163) := x"FD08";
          m(164) := x"FF7C";
          m(165) := x"02E6";
          m(166) := x"018F";
          m(167) := x"0098";
          m(168) := x"FFF2";
          m(169) := x"FFF1";
          m(170) := x"0007";
          m(171) := x"0018";
          m(172) := x"FFEA";
          m(173) := x"0129";
          m(174) := x"033D";
          m(175) := x"0454";
          m(176) := x"015D";
          m(177) := x"FEF2";
          m(178) := x"0177";
          m(179) := x"00B3";
          m(180) := x"FF44";
          m(181) := x"00AD";
          m(182) := x"FE3D";
          m(183) := x"00A3";
          m(184) := x"01CA";
          m(185) := x"FEDB";
          m(186) := x"FD60";
          m(187) := x"FF89";
          m(188) := x"00CE";
          m(189) := x"FF1E";
          m(190) := x"FFFA";
          m(191) := x"FF02";
          m(192) := x"FF28";
          m(193) := x"0245";
          m(194) := x"0111";
          m(195) := x"0074";
          m(196) := x"001E";
          m(197) := x"0073";
          m(198) := x"0059";
          m(199) := x"0025";
          m(200) := x"00A4";
          m(201) := x"0525";
          m(202) := x"06CB";
          m(203) := x"06DC";
          m(204) := x"01E7";
          m(205) := x"FCF7";
          m(206) := x"FF1B";
          m(207) := x"FF8C";
          m(208) := x"FC68";
          m(209) := x"FBD5";
          m(210) := x"F85A";
          m(211) := x"0123";
          m(212) := x"FEDD";
          m(213) := x"0295";
          m(214) := x"024F";
          m(215) := x"FFE2";
          m(216) := x"FFDC";
          m(217) := x"0249";
          m(218) := x"03DE";
          m(219) := x"0021";
          m(220) := x"0366";
          m(221) := x"0291";
          m(222) := x"FFE5";
          m(223) := x"0092";
          m(224) := x"0001";
          m(225) := x"0024";
          m(226) := x"008D";
          m(227) := x"FFDB";
          m(228) := x"0213";
          m(229) := x"04DA";
          m(230) := x"04BA";
          m(231) := x"03BC";
          m(232) := x"006A";
          m(233) := x"FDEB";
          m(234) := x"03F7";
          m(235) := x"0313";
          m(236) := x"0380";
          m(237) := x"00E8";
          m(238) := x"FCDB";
          m(239) := x"FF1D";
          m(240) := x"03FF";
          m(241) := x"010F";
          m(242) := x"FEA5";
          m(243) := x"01B2";
          m(244) := x"0390";
          m(245) := x"020C";
          m(246) := x"FEDD";
          m(247) := x"0393";
          m(248) := x"035E";
          m(249) := x"FF52";
          m(250) := x"0047";
          m(251) := x"FFF5";
          m(252) := x"0035";
          m(253) := x"002D";
          m(254) := x"0037";
          m(255) := x"FFF3";
          m(256) := x"01EF";
          m(257) := x"023D";
          m(258) := x"01DB";
          m(259) := x"0152";
          m(260) := x"00B9";
          m(261) := x"0017";
          m(262) := x"FF20";
          m(263) := x"0409";
          m(264) := x"01C4";
          m(265) := x"04B8";
          m(266) := x"FCEA";
          m(267) := x"FB46";
          m(268) := x"FEFC";
          m(269) := x"00F5";
          m(270) := x"0040";
          m(271) := x"FE81";
          m(272) := x"02AC";
          m(273) := x"008A";
          m(274) := x"0094";
          m(275) := x"0763";
          m(276) := x"0076";
          m(277) := x"FFA3";
          m(278) := x"FF77";
          m(279) := x"FEDA";
          m(280) := x"0003";
          m(281) := x"FFE5";
          m(282) := x"0025";
          m(283) := x"FFED";
          m(284) := x"010E";
          m(285) := x"00DE";
          m(286) := x"0396";
          m(287) := x"0362";
          m(288) := x"FFF0";
          m(289) := x"FEB7";
          m(290) := x"0285";
          m(291) := x"025E";
          m(292) := x"021C";
          m(293) := x"01D5";
          m(294) := x"FD6A";
          m(295) := x"FA93";
          m(296) := x"FAF6";
          m(297) := x"0470";
          m(298) := x"FF97";
          m(299) := x"FC01";
          m(300) := x"01CC";
          m(301) := x"00F4";
          m(302) := x"FFA1";
          m(303) := x"003B";
          m(304) := x"FCEE";
          m(305) := x"FB93";
          m(306) := x"FF67";
          m(307) := x"FFE7";
          m(308) := x"0039";
          m(309) := x"FFFE";
          m(310) := x"FFBC";
          m(311) := x"0027";
          m(312) := x"0007";
          m(313) := x"00E6";
          m(314) := x"0443";
          m(315) := x"03FD";
          m(316) := x"0145";
          m(317) := x"000E";
          m(318) := x"FDA4";
          m(319) := x"030D";
          m(320) := x"083F";
          m(321) := x"0328";
          m(322) := x"FF8A";
          m(323) := x"FFFE";
          m(324) := x"F94D";
          m(325) := x"FD93";
          m(326) := x"FC9A";
          m(327) := x"FD94";
          m(328) := x"FD30";
          m(329) := x"FC37";
          m(330) := x"FEC4";
          m(331) := x"FCE5";
          m(332) := x"FCA6";
          m(333) := x"FEC0";
          m(334) := x"FFE5";
          m(335) := x"FFE6";
          m(336) := x"FFD8";
          m(337) := x"000C";
          m(338) := x"FFB3";
          m(339) := x"0037";
          m(340) := x"0082";
          m(341) := x"01C0";
          m(342) := x"031F";
          m(343) := x"0218";
          m(344) := x"03BB";
          m(345) := x"0462";
          m(346) := x"0027";
          m(347) := x"037E";
          m(348) := x"09C3";
          m(349) := x"00B4";
          m(350) := x"FB71";
          m(351) := x"FB7D";
          m(352) := x"FB69";
          m(353) := x"FF73";
          m(354) := x"FDD9";
          m(355) := x"0260";
          m(356) := x"017B";
          m(357) := x"008B";
          m(358) := x"FF3D";
          m(359) := x"0044";
          m(360) := x"0081";
          m(361) := x"FF6F";
          m(362) := x"FEF3";
          m(363) := x"FFDC";
          m(364) := x"FFE1";
          m(365) := x"0031";
          m(366) := x"FFC0";
          m(367) := x"00F1";
          m(368) := x"0046";
          m(369) := x"0369";
          m(370) := x"0233";
          m(371) := x"FF3E";
          m(372) := x"FDE0";
          m(373) := x"FE51";
          m(374) := x"FC70";
          m(375) := x"027D";
          m(376) := x"04F0";
          m(377) := x"00C1";
          m(378) := x"FE53";
          m(379) := x"FD2B";
          m(380) := x"FE49";
          m(381) := x"00C7";
          m(382) := x"070F";
          m(383) := x"02E4";
          m(384) := x"02A5";
          m(385) := x"022C";
          m(386) := x"02F1";
          m(387) := x"01B0";
          m(388) := x"0178";
          m(389) := x"FFE6";
          m(390) := x"004B";
          m(391) := x"004A";
          m(392) := x"FFEC";
          m(393) := x"FFF5";
          m(394) := x"FFD0";
          m(395) := x"00DD";
          m(396) := x"00FC";
          m(397) := x"0354";
          m(398) := x"023C";
          m(399) := x"FFF2";
          m(400) := x"FF99";
          m(401) := x"FDA4";
          m(402) := x"FC0C";
          m(403) := x"FF55";
          m(404) := x"0051";
          m(405) := x"00F3";
          m(406) := x"FDF9";
          m(407) := x"FD52";
          m(408) := x"FE70";
          m(409) := x"04D4";
          m(410) := x"0400";
          m(411) := x"00D5";
          m(412) := x"0169";
          m(413) := x"0033";
          m(414) := x"0131";
          m(415) := x"009C";
          m(416) := x"005F";
          m(417) := x"FFE7";
          m(418) := x"00CF";
          m(419) := x"FFF1";
          m(420) := x"0029";
          m(421) := x"FFED";
          m(422) := x"0004";
          m(423) := x"014E";
          m(424) := x"0101";
          m(425) := x"00B0";
          m(426) := x"00BE";
          m(427) := x"010D";
          m(428) := x"0308";
          m(429) := x"FD68";
          m(430) := x"FEE6";
          m(431) := x"FEFC";
          m(432) := x"FC77";
          m(433) := x"018B";
          m(434) := x"FF5A";
          m(435) := x"FB5A";
          m(436) := x"FEC9";
          m(437) := x"FF77";
          m(438) := x"0094";
          m(439) := x"0489";
          m(440) := x"01DB";
          m(441) := x"FF50";
          m(442) := x"00FC";
          m(443) := x"FF49";
          m(444) := x"01A5";
          m(445) := x"01A7";
          m(446) := x"00C6";
          m(447) := x"FFFC";
          m(448) := x"FFFF";
          m(449) := x"0017";
          m(450) := x"001E";
          m(451) := x"017E";
          m(452) := x"FFA8";
          m(453) := x"FE44";
          m(454) := x"01E5";
          m(455) := x"06B6";
          m(456) := x"05CB";
          m(457) := x"0390";
          m(458) := x"01D6";
          m(459) := x"FFE8";
          m(460) := x"03E3";
          m(461) := x"00F8";
          m(462) := x"FC9E";
          m(463) := x"FBFA";
          m(464) := x"FFF3";
          m(465) := x"099F";
          m(466) := x"0834";
          m(467) := x"0602";
          m(468) := x"0120";
          m(469) := x"011E";
          m(470) := x"017E";
          m(471) := x"0104";
          m(472) := x"02CA";
          m(473) := x"0207";
          m(474) := x"00D6";
          m(475) := x"FFE3";
          m(476) := x"FFB0";
          m(477) := x"FFC6";
          m(478) := x"0005";
          m(479) := x"003F";
          m(480) := x"FEEC";
          m(481) := x"FE24";
          m(482) := x"047B";
          m(483) := x"09C8";
          m(484) := x"0985";
          m(485) := x"0777";
          m(486) := x"0476";
          m(487) := x"017A";
          m(488) := x"0520";
          m(489) := x"015E";
          m(490) := x"FC40";
          m(491) := x"FEBA";
          m(492) := x"0811";
          m(493) := x"0A31";
          m(494) := x"0467";
          m(495) := x"035C";
          m(496) := x"013B";
          m(497) := x"00F2";
          m(498) := x"FED9";
          m(499) := x"FDE5";
          m(500) := x"FFCC";
          m(501) := x"00F8";
          m(502) := x"FF7A";
          m(503) := x"000D";
          m(504) := x"FFE6";
          m(505) := x"0024";
          m(506) := x"FFEF";
          m(507) := x"0101";
          m(508) := x"FE67";
          m(509) := x"FEED";
          m(510) := x"03F2";
          m(511) := x"0775";
          m(512) := x"0756";
          m(513) := x"089E";
          m(514) := x"04C9";
          m(515) := x"007F";
          m(516) := x"0004";
          m(517) := x"FDB8";
          m(518) := x"FFB7";
          m(519) := x"01DF";
          m(520) := x"067D";
          m(521) := x"050B";
          m(522) := x"00E6";
          m(523) := x"027E";
          m(524) := x"019B";
          m(525) := x"02B0";
          m(526) := x"030E";
          m(527) := x"0263";
          m(528) := x"00E4";
          m(529) := x"FF8D";
          m(530) := x"FF81";
          m(531) := x"FFD1";
          m(532) := x"0015";
          m(533) := x"000B";
          m(534) := x"FFBE";
          m(535) := x"001E";
          m(536) := x"FF45";
          m(537) := x"002C";
          m(538) := x"0024";
          m(539) := x"FE7E";
          m(540) := x"FFB7";
          m(541) := x"0250";
          m(542) := x"003D";
          m(543) := x"FEF0";
          m(544) := x"FCE9";
          m(545) := x"FDC8";
          m(546) := x"016F";
          m(547) := x"05E3";
          m(548) := x"01DC";
          m(549) := x"0232";
          m(550) := x"00C0";
          m(551) := x"024C";
          m(552) := x"0397";
          m(553) := x"03E7";
          m(554) := x"019B";
          m(555) := x"0178";
          m(556) := x"FF21";
          m(557) := x"FEDD";
          m(558) := x"000C";
          m(559) := x"FFF2";
          m(560) := x"FFFB";
          m(561) := x"FFDE";
          m(562) := x"FFD2";
          m(563) := x"00B6";
          m(564) := x"010A";
          m(565) := x"FEA8";
          m(566) := x"FB89";
          m(567) := x"0071";
          m(568) := x"FE7D";
          m(569) := x"FD07";
          m(570) := x"FC2F";
          m(571) := x"FD38";
          m(572) := x"FEF0";
          m(573) := x"0012";
          m(574) := x"04CB";
          m(575) := x"057D";
          m(576) := x"FEAD";
          m(577) := x"0120";
          m(578) := x"0396";
          m(579) := x"01EC";
          m(580) := x"0237";
          m(581) := x"0032";
          m(582) := x"FEEF";
          m(583) := x"006C";
          m(584) := x"FF59";
          m(585) := x"0042";
          m(586) := x"FFEE";
          m(587) := x"FFCD";
          m(588) := x"FFEA";
          m(589) := x"0000";
          m(590) := x"008F";
          m(591) := x"00AA";
          m(592) := x"FEC9";
          m(593) := x"FF93";
          m(594) := x"FCDB";
          m(595) := x"FB20";
          m(596) := x"FC24";
          m(597) := x"FD75";
          m(598) := x"F73B";
          m(599) := x"FDC9";
          m(600) := x"FCB2";
          m(601) := x"0277";
          m(602) := x"040B";
          m(603) := x"03C2";
          m(604) := x"0414";
          m(605) := x"05E9";
          m(606) := x"0706";
          m(607) := x"06D2";
          m(608) := x"0349";
          m(609) := x"00E9";
          m(610) := x"0100";
          m(611) := x"00B2";
          m(612) := x"009E";
          m(613) := x"007E";
          m(614) := x"0055";
          m(615) := x"FFE0";
          m(616) := x"FFE1";
          m(617) := x"0032";
          m(618) := x"0050";
          m(619) := x"FEF2";
          m(620) := x"FF6A";
          m(621) := x"0059";
          m(622) := x"FD39";
          m(623) := x"FF43";
          m(624) := x"FB95";
          m(625) := x"FDE8";
          m(626) := x"FDA2";
          m(627) := x"0010";
          m(628) := x"FF83";
          m(629) := x"FFD2";
          m(630) := x"056C";
          m(631) := x"05D4";
          m(632) := x"075D";
          m(633) := x"0712";
          m(634) := x"0871";
          m(635) := x"0525";
          m(636) := x"0326";
          m(637) := x"0168";
          m(638) := x"0045";
          m(639) := x"FF60";
          m(640) := x"007D";
          m(641) := x"008A";
          m(642) := x"0000";
          m(643) := x"FFF9";
          m(644) := x"000E";
          m(645) := x"001E";
          m(646) := x"008C";
          m(647) := x"FFA4";
          m(648) := x"FFA9";
          m(649) := x"FF8A";
          m(650) := x"FF60";
          m(651) := x"FEFA";
          m(652) := x"FF9D";
          m(653) := x"03BC";
          m(654) := x"042B";
          m(655) := x"0325";
          m(656) := x"011C";
          m(657) := x"02B7";
          m(658) := x"0864";
          m(659) := x"07CD";
          m(660) := x"084D";
          m(661) := x"06A6";
          m(662) := x"05E8";
          m(663) := x"041B";
          m(664) := x"02BF";
          m(665) := x"01CF";
          m(666) := x"0059";
          m(667) := x"FEFA";
          m(668) := x"0035";
          m(669) := x"0086";
          m(670) := x"FFBE";
          m(671) := x"FFE8";
          m(672) := x"0000";
          m(673) := x"FFF7";
          m(674) := x"005B";
          m(675) := x"0032";
          m(676) := x"FFF1";
          m(677) := x"FEB9";
          m(678) := x"FE3A";
          m(679) := x"FC25";
          m(680) := x"FCEE";
          m(681) := x"FEC0";
          m(682) := x"003A";
          m(683) := x"01D3";
          m(684) := x"03CF";
          m(685) := x"0027";
          m(686) := x"00B5";
          m(687) := x"0582";
          m(688) := x"0665";
          m(689) := x"07D4";
          m(690) := x"0597";
          m(691) := x"0506";
          m(692) := x"0422";
          m(693) := x"01C9";
          m(694) := x"FF30";
          m(695) := x"FE99";
          m(696) := x"FFE4";
          m(697) := x"0001";
          m(698) := x"0023";
          m(699) := x"0001";
          m(700) := x"FFDC";
          m(701) := x"FFC4";
          m(702) := x"FFEE";
          m(703) := x"FFDF";
          m(704) := x"FD77";
          m(705) := x"FBE0";
          m(706) := x"FCD8";
          m(707) := x"FD70";
          m(708) := x"FBDD";
          m(709) := x"FE02";
          m(710) := x"011B";
          m(711) := x"00B0";
          m(712) := x"016C";
          m(713) := x"FF78";
          m(714) := x"FFEB";
          m(715) := x"043D";
          m(716) := x"0324";
          m(717) := x"0444";
          m(718) := x"04B8";
          m(719) := x"03C4";
          m(720) := x"0174";
          m(721) := x"0085";
          m(722) := x"FF61";
          m(723) := x"FF15";
          m(724) := x"FFB6";
          m(725) := x"0000";
          m(726) := x"0005";
          m(727) := x"FFDB";
          m(728) := x"FFF1";
          m(729) := x"000D";
          m(730) := x"0009";
          m(731) := x"FFD3";
          m(732) := x"FF52";
          m(733) := x"FE41";
          m(734) := x"FDA8";
          m(735) := x"FD36";
          m(736) := x"FF5B";
          m(737) := x"FE38";
          m(738) := x"FF71";
          m(739) := x"0101";
          m(740) := x"FE33";
          m(741) := x"FE29";
          m(742) := x"FEDC";
          m(743) := x"0087";
          m(744) := x"FF89";
          m(745) := x"FF66";
          m(746) := x"FF79";
          m(747) := x"FFC3";
          m(748) := x"0000";
          m(749) := x"0008";
          m(750) := x"0000";
          m(751) := x"FFD0";
          m(752) := x"0028";
          m(753) := x"0024";
          m(754) := x"001C";
          m(755) := x"FFD3";
          m(756) := x"FFD1";
          m(757) := x"0033";
          m(758) := x"0000";
          m(759) := x"0001";
          m(760) := x"FFE6";
          m(761) := x"0000";
          m(762) := x"000A";
          m(763) := x"0009";
          m(764) := x"FFDE";
          m(765) := x"FFFD";
          m(766) := x"0002";
          m(767) := x"FFCF";
          m(768) := x"FFE5";
          m(769) := x"FFC3";
          m(770) := x"FFC5";
          m(771) := x"FFF3";
          m(772) := x"FFF5";
          m(773) := x"FFC5";
          m(774) := x"FFA5";
          m(775) := x"FFE3";
          m(776) := x"0003";
          m(777) := x"FFD8";
          m(778) := x"002E";
          m(779) := x"0002";
          m(780) := x"0014";
          m(781) := x"0027";
          m(782) := x"FFF5";
          m(783) := x"FFC2";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_1.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 1) then
          m(0) := x"000E";
          m(1) := x"0003";
          m(2) := x"FFDB";
          m(3) := x"0020";
          m(4) := x"002A";
          m(5) := x"FFE1";
          m(6) := x"FFFF";
          m(7) := x"FF9B";
          m(8) := x"FFFA";
          m(9) := x"FFE8";
          m(10) := x"FFED";
          m(11) := x"FFF9";
          m(12) := x"FFD9";
          m(13) := x"0003";
          m(14) := x"002A";
          m(15) := x"0022";
          m(16) := x"FFD1";
          m(17) := x"FFBA";
          m(18) := x"FFE1";
          m(19) := x"FFE8";
          m(20) := x"FFF3";
          m(21) := x"FFE7";
          m(22) := x"FFF0";
          m(23) := x"0028";
          m(24) := x"FFFC";
          m(25) := x"001E";
          m(26) := x"0006";
          m(27) := x"FFE4";
          m(28) := x"0010";
          m(29) := x"0018";
          m(30) := x"0006";
          m(31) := x"FFEE";
          m(32) := x"FFEE";
          m(33) := x"002E";
          m(34) := x"0015";
          m(35) := x"FFF2";
          m(36) := x"000B";
          m(37) := x"FFDF";
          m(38) := x"FFCF";
          m(39) := x"0014";
          m(40) := x"FFFC";
          m(41) := x"FFE1";
          m(42) := x"0013";
          m(43) := x"FF9E";
          m(44) := x"0017";
          m(45) := x"FFEE";
          m(46) := x"FFFA";
          m(47) := x"FFDF";
          m(48) := x"FFEF";
          m(49) := x"0034";
          m(50) := x"FFB5";
          m(51) := x"0001";
          m(52) := x"FFF2";
          m(53) := x"FFFC";
          m(54) := x"002C";
          m(55) := x"FFEA";
          m(56) := x"001E";
          m(57) := x"0036";
          m(58) := x"0000";
          m(59) := x"FFE0";
          m(60) := x"FFE6";
          m(61) := x"002A";
          m(62) := x"FFC5";
          m(63) := x"FFD7";
          m(64) := x"FFAB";
          m(65) := x"FF8E";
          m(66) := x"FF54";
          m(67) := x"FE94";
          m(68) := x"FE2D";
          m(69) := x"FE5C";
          m(70) := x"FE89";
          m(71) := x"FE74";
          m(72) := x"FECB";
          m(73) := x"FF1A";
          m(74) := x"FF43";
          m(75) := x"FFC8";
          m(76) := x"FFF5";
          m(77) := x"0030";
          m(78) := x"FFFA";
          m(79) := x"FFED";
          m(80) := x"FFE5";
          m(81) := x"000A";
          m(82) := x"FFF3";
          m(83) := x"0021";
          m(84) := x"000F";
          m(85) := x"FFE4";
          m(86) := x"FFFF";
          m(87) := x"FFED";
          m(88) := x"FFE5";
          m(89) := x"FFE1";
          m(90) := x"FF9A";
          m(91) := x"FF47";
          m(92) := x"FE21";
          m(93) := x"FE97";
          m(94) := x"FF52";
          m(95) := x"FD62";
          m(96) := x"FB55";
          m(97) := x"FB05";
          m(98) := x"FD22";
          m(99) := x"FE22";
          m(100) := x"FDC4";
          m(101) := x"FCE0";
          m(102) := x"FB76";
          m(103) := x"FD88";
          m(104) := x"FF78";
          m(105) := x"FF76";
          m(106) := x"FF34";
          m(107) := x"FFF4";
          m(108) := x"0031";
          m(109) := x"FFE5";
          m(110) := x"FFEA";
          m(111) := x"FFC8";
          m(112) := x"FFF4";
          m(113) := x"FFF6";
          m(114) := x"FFE4";
          m(115) := x"FFD9";
          m(116) := x"FFB3";
          m(117) := x"FF9E";
          m(118) := x"0003";
          m(119) := x"FEF6";
          m(120) := x"FCDD";
          m(121) := x"FEF9";
          m(122) := x"0105";
          m(123) := x"FE9E";
          m(124) := x"FA58";
          m(125) := x"FBAB";
          m(126) := x"F971";
          m(127) := x"FAF9";
          m(128) := x"FC30";
          m(129) := x"FFFD";
          m(130) := x"FF8B";
          m(131) := x"FC52";
          m(132) := x"FC8A";
          m(133) := x"FDD5";
          m(134) := x"FFA7";
          m(135) := x"0081";
          m(136) := x"0000";
          m(137) := x"FFD0";
          m(138) := x"FFD1";
          m(139) := x"0005";
          m(140) := x"0004";
          m(141) := x"0003";
          m(142) := x"001F";
          m(143) := x"FFED";
          m(144) := x"0018";
          m(145) := x"FFCD";
          m(146) := x"0042";
          m(147) := x"FEA0";
          m(148) := x"0092";
          m(149) := x"01C0";
          m(150) := x"FFB5";
          m(151) := x"FC91";
          m(152) := x"FED7";
          m(153) := x"FE67";
          m(154) := x"FE02";
          m(155) := x"FBA2";
          m(156) := x"FD31";
          m(157) := x"FEBA";
          m(158) := x"026C";
          m(159) := x"FDB9";
          m(160) := x"FA83";
          m(161) := x"FD04";
          m(162) := x"FFDD";
          m(163) := x"FF9D";
          m(164) := x"FE2B";
          m(165) := x"FF62";
          m(166) := x"FFBA";
          m(167) := x"FFEF";
          m(168) := x"001B";
          m(169) := x"FFD1";
          m(170) := x"0022";
          m(171) := x"0013";
          m(172) := x"004F";
          m(173) := x"026A";
          m(174) := x"00EE";
          m(175) := x"FFD5";
          m(176) := x"059D";
          m(177) := x"04DB";
          m(178) := x"0535";
          m(179) := x"FF85";
          m(180) := x"04AA";
          m(181) := x"FF45";
          m(182) := x"FF3D";
          m(183) := x"F70C";
          m(184) := x"FA84";
          m(185) := x"FF8F";
          m(186) := x"0256";
          m(187) := x"FFB3";
          m(188) := x"F8D5";
          m(189) := x"001D";
          m(190) := x"FFD2";
          m(191) := x"FD92";
          m(192) := x"FC38";
          m(193) := x"FD63";
          m(194) := x"FF7D";
          m(195) := x"FFDD";
          m(196) := x"FFD5";
          m(197) := x"0022";
          m(198) := x"0011";
          m(199) := x"015D";
          m(200) := x"00CA";
          m(201) := x"FFB9";
          m(202) := x"0581";
          m(203) := x"062A";
          m(204) := x"015A";
          m(205) := x"099A";
          m(206) := x"03A6";
          m(207) := x"008E";
          m(208) := x"00BB";
          m(209) := x"FEEE";
          m(210) := x"FD95";
          m(211) := x"F6EA";
          m(212) := x"FBA2";
          m(213) := x"FEE4";
          m(214) := x"046B";
          m(215) := x"FEAA";
          m(216) := x"FC5A";
          m(217) := x"FA6C";
          m(218) := x"FF84";
          m(219) := x"FD7B";
          m(220) := x"FE42";
          m(221) := x"FE73";
          m(222) := x"FFC8";
          m(223) := x"FFE6";
          m(224) := x"0025";
          m(225) := x"001D";
          m(226) := x"004D";
          m(227) := x"0045";
          m(228) := x"0066";
          m(229) := x"FFB6";
          m(230) := x"0197";
          m(231) := x"06B3";
          m(232) := x"0AF1";
          m(233) := x"0B1D";
          m(234) := x"077C";
          m(235) := x"0161";
          m(236) := x"085D";
          m(237) := x"FEBE";
          m(238) := x"FC23";
          m(239) := x"FF5E";
          m(240) := x"F754";
          m(241) := x"03C5";
          m(242) := x"0182";
          m(243) := x"FF25";
          m(244) := x"0155";
          m(245) := x"FEC5";
          m(246) := x"032E";
          m(247) := x"02A1";
          m(248) := x"00C2";
          m(249) := x"FF8C";
          m(250) := x"000C";
          m(251) := x"FFDF";
          m(252) := x"0013";
          m(253) := x"0035";
          m(254) := x"003C";
          m(255) := x"FF2A";
          m(256) := x"0179";
          m(257) := x"050D";
          m(258) := x"0589";
          m(259) := x"05DD";
          m(260) := x"0133";
          m(261) := x"0766";
          m(262) := x"051E";
          m(263) := x"02D9";
          m(264) := x"06A7";
          m(265) := x"0499";
          m(266) := x"FACA";
          m(267) := x"FD86";
          m(268) := x"FC74";
          m(269) := x"0020";
          m(270) := x"FEEA";
          m(271) := x"00EB";
          m(272) := x"FF9A";
          m(273) := x"0649";
          m(274) := x"059B";
          m(275) := x"0464";
          m(276) := x"FFF7";
          m(277) := x"FE51";
          m(278) := x"FDF3";
          m(279) := x"0001";
          m(280) := x"FFE5";
          m(281) := x"0018";
          m(282) := x"007C";
          m(283) := x"000E";
          m(284) := x"0190";
          m(285) := x"01BE";
          m(286) := x"04FD";
          m(287) := x"0029";
          m(288) := x"FECB";
          m(289) := x"06EE";
          m(290) := x"0993";
          m(291) := x"0C25";
          m(292) := x"0D70";
          m(293) := x"0CEA";
          m(294) := x"FCFF";
          m(295) := x"FFA0";
          m(296) := x"0264";
          m(297) := x"091F";
          m(298) := x"0229";
          m(299) := x"00B8";
          m(300) := x"0271";
          m(301) := x"0352";
          m(302) := x"00BD";
          m(303) := x"00FE";
          m(304) := x"FB03";
          m(305) := x"FCB8";
          m(306) := x"FEBA";
          m(307) := x"0000";
          m(308) := x"FFD1";
          m(309) := x"002A";
          m(310) := x"FFA9";
          m(311) := x"0030";
          m(312) := x"FFA2";
          m(313) := x"FE3E";
          m(314) := x"FF51";
          m(315) := x"FC42";
          m(316) := x"FBF8";
          m(317) := x"064A";
          m(318) := x"01D7";
          m(319) := x"0D02";
          m(320) := x"0550";
          m(321) := x"F871";
          m(322) := x"EED0";
          m(323) := x"FEFD";
          m(324) := x"016D";
          m(325) := x"0648";
          m(326) := x"04C2";
          m(327) := x"0356";
          m(328) := x"00FF";
          m(329) := x"0309";
          m(330) := x"FF2A";
          m(331) := x"FD7C";
          m(332) := x"FD85";
          m(333) := x"FF1A";
          m(334) := x"FFFF";
          m(335) := x"FFF2";
          m(336) := x"0021";
          m(337) := x"00B0";
          m(338) := x"FFD7";
          m(339) := x"FFBD";
          m(340) := x"FD98";
          m(341) := x"FD67";
          m(342) := x"FF9E";
          m(343) := x"047E";
          m(344) := x"04FA";
          m(345) := x"0015";
          m(346) := x"0314";
          m(347) := x"0577";
          m(348) := x"FFAB";
          m(349) := x"F11B";
          m(350) := x"EA30";
          m(351) := x"FC4C";
          m(352) := x"02DA";
          m(353) := x"006E";
          m(354) := x"03F0";
          m(355) := x"FDCA";
          m(356) := x"FF57";
          m(357) := x"FEE3";
          m(358) := x"FFF2";
          m(359) := x"FCBF";
          m(360) := x"003F";
          m(361) := x"FFF9";
          m(362) := x"FFEF";
          m(363) := x"FFEE";
          m(364) := x"0007";
          m(365) := x"0063";
          m(366) := x"00E1";
          m(367) := x"014A";
          m(368) := x"F95F";
          m(369) := x"FE1E";
          m(370) := x"031F";
          m(371) := x"FDE5";
          m(372) := x"0322";
          m(373) := x"008C";
          m(374) := x"FBF8";
          m(375) := x"02BD";
          m(376) := x"F2DF";
          m(377) := x"EC92";
          m(378) := x"F18C";
          m(379) := x"F1D1";
          m(380) := x"FD03";
          m(381) := x"02CE";
          m(382) := x"01B8";
          m(383) := x"FB9E";
          m(384) := x"0480";
          m(385) := x"FFE7";
          m(386) := x"FD12";
          m(387) := x"FCAD";
          m(388) := x"018A";
          m(389) := x"000A";
          m(390) := x"FFBE";
          m(391) := x"FFFD";
          m(392) := x"FFE2";
          m(393) := x"0000";
          m(394) := x"017B";
          m(395) := x"0174";
          m(396) := x"FA3D";
          m(397) := x"044E";
          m(398) := x"0153";
          m(399) := x"01E6";
          m(400) := x"0346";
          m(401) := x"020A";
          m(402) := x"0AB7";
          m(403) := x"0190";
          m(404) := x"F0BD";
          m(405) := x"EDB7";
          m(406) := x"F992";
          m(407) := x"F9F9";
          m(408) := x"FD32";
          m(409) := x"FADD";
          m(410) := x"FF70";
          m(411) := x"FEB3";
          m(412) := x"FEA8";
          m(413) := x"FE4E";
          m(414) := x"FDC6";
          m(415) := x"0009";
          m(416) := x"0295";
          m(417) := x"FF86";
          m(418) := x"FFC5";
          m(419) := x"FFB2";
          m(420) := x"0001";
          m(421) := x"FFDE";
          m(422) := x"0166";
          m(423) := x"01A5";
          m(424) := x"FD8F";
          m(425) := x"010F";
          m(426) := x"0270";
          m(427) := x"04CE";
          m(428) := x"FEE8";
          m(429) := x"FD89";
          m(430) := x"0224";
          m(431) := x"F4D0";
          m(432) := x"E7AB";
          m(433) := x"F106";
          m(434) := x"FA8E";
          m(435) := x"FBF6";
          m(436) := x"F728";
          m(437) := x"F946";
          m(438) := x"FD69";
          m(439) := x"FCEA";
          m(440) := x"FACD";
          m(441) := x"FC93";
          m(442) := x"FF6C";
          m(443) := x"01BD";
          m(444) := x"038A";
          m(445) := x"FFC0";
          m(446) := x"0070";
          m(447) := x"0016";
          m(448) := x"FFFE";
          m(449) := x"0002";
          m(450) := x"00E1";
          m(451) := x"FFFA";
          m(452) := x"FEAB";
          m(453) := x"FC5D";
          m(454) := x"FDF3";
          m(455) := x"0209";
          m(456) := x"FE70";
          m(457) := x"F72B";
          m(458) := x"FAAF";
          m(459) := x"EA81";
          m(460) := x"EF63";
          m(461) := x"F987";
          m(462) := x"FC4C";
          m(463) := x"00F9";
          m(464) := x"FE65";
          m(465) := x"F9AA";
          m(466) := x"F9AC";
          m(467) := x"FF53";
          m(468) := x"FD73";
          m(469) := x"0228";
          m(470) := x"0058";
          m(471) := x"0175";
          m(472) := x"0119";
          m(473) := x"FEA5";
          m(474) := x"0091";
          m(475) := x"000D";
          m(476) := x"FFEA";
          m(477) := x"0018";
          m(478) := x"FFC3";
          m(479) := x"FE3A";
          m(480) := x"FE64";
          m(481) := x"FD29";
          m(482) := x"FB98";
          m(483) := x"FA30";
          m(484) := x"FA62";
          m(485) := x"F68C";
          m(486) := x"F767";
          m(487) := x"F592";
          m(488) := x"F986";
          m(489) := x"0071";
          m(490) := x"0024";
          m(491) := x"FF22";
          m(492) := x"FB86";
          m(493) := x"01B9";
          m(494) := x"FF12";
          m(495) := x"FF95";
          m(496) := x"011F";
          m(497) := x"02BF";
          m(498) := x"0296";
          m(499) := x"0402";
          m(500) := x"02FA";
          m(501) := x"02B8";
          m(502) := x"FFFF";
          m(503) := x"0038";
          m(504) := x"FFEC";
          m(505) := x"FFC9";
          m(506) := x"004C";
          m(507) := x"FE34";
          m(508) := x"FD8D";
          m(509) := x"FBD0";
          m(510) := x"F8FD";
          m(511) := x"F959";
          m(512) := x"FA7C";
          m(513) := x"F8BD";
          m(514) := x"F930";
          m(515) := x"0094";
          m(516) := x"FC85";
          m(517) := x"FFDE";
          m(518) := x"01A6";
          m(519) := x"FBC1";
          m(520) := x"F968";
          m(521) := x"FCD3";
          m(522) := x"0491";
          m(523) := x"FEDB";
          m(524) := x"FF06";
          m(525) := x"0537";
          m(526) := x"03A1";
          m(527) := x"029C";
          m(528) := x"FFA0";
          m(529) := x"018E";
          m(530) := x"0024";
          m(531) := x"FFE7";
          m(532) := x"FFDE";
          m(533) := x"003B";
          m(534) := x"0035";
          m(535) := x"FED4";
          m(536) := x"FEEB";
          m(537) := x"FFB5";
          m(538) := x"FADD";
          m(539) := x"FA44";
          m(540) := x"FB13";
          m(541) := x"F8CF";
          m(542) := x"0030";
          m(543) := x"FD2D";
          m(544) := x"FB66";
          m(545) := x"FBD5";
          m(546) := x"03A2";
          m(547) := x"FACC";
          m(548) := x"FE5D";
          m(549) := x"0085";
          m(550) := x"FE06";
          m(551) := x"022E";
          m(552) := x"01DC";
          m(553) := x"0115";
          m(554) := x"005A";
          m(555) := x"FEEC";
          m(556) := x"FF07";
          m(557) := x"FFF4";
          m(558) := x"FFE2";
          m(559) := x"FFCA";
          m(560) := x"FFFE";
          m(561) := x"FFE9";
          m(562) := x"000A";
          m(563) := x"FF6B";
          m(564) := x"FF7F";
          m(565) := x"FE2D";
          m(566) := x"FC52";
          m(567) := x"FCA3";
          m(568) := x"FE2D";
          m(569) := x"FC9E";
          m(570) := x"FEC7";
          m(571) := x"049B";
          m(572) := x"01C1";
          m(573) := x"04A1";
          m(574) := x"038F";
          m(575) := x"03AF";
          m(576) := x"FE34";
          m(577) := x"F98D";
          m(578) := x"F9F3";
          m(579) := x"FB4B";
          m(580) := x"FD19";
          m(581) := x"FEE8";
          m(582) := x"007B";
          m(583) := x"00A6";
          m(584) := x"FEE9";
          m(585) := x"FE17";
          m(586) := x"FFF8";
          m(587) := x"FFF7";
          m(588) := x"001E";
          m(589) := x"FFDB";
          m(590) := x"FFE9";
          m(591) := x"FEC7";
          m(592) := x"FE68";
          m(593) := x"FD89";
          m(594) := x"FE21";
          m(595) := x"FBCD";
          m(596) := x"FE1E";
          m(597) := x"0076";
          m(598) := x"0495";
          m(599) := x"05BC";
          m(600) := x"FF31";
          m(601) := x"013E";
          m(602) := x"FDFA";
          m(603) := x"02F6";
          m(604) := x"02C1";
          m(605) := x"00E8";
          m(606) := x"FF6D";
          m(607) := x"FD8C";
          m(608) := x"0029";
          m(609) := x"0017";
          m(610) := x"FFCF";
          m(611) := x"0274";
          m(612) := x"0009";
          m(613) := x"FFDC";
          m(614) := x"FFF4";
          m(615) := x"FFDA";
          m(616) := x"0006";
          m(617) := x"0023";
          m(618) := x"FFDB";
          m(619) := x"FED5";
          m(620) := x"FE72";
          m(621) := x"FF88";
          m(622) := x"01E1";
          m(623) := x"0105";
          m(624) := x"042B";
          m(625) := x"0507";
          m(626) := x"03E4";
          m(627) := x"FB5B";
          m(628) := x"FBF1";
          m(629) := x"01E5";
          m(630) := x"0235";
          m(631) := x"0660";
          m(632) := x"04C5";
          m(633) := x"06FF";
          m(634) := x"04C3";
          m(635) := x"FDA7";
          m(636) := x"FE3B";
          m(637) := x"023C";
          m(638) := x"0087";
          m(639) := x"00BA";
          m(640) := x"001E";
          m(641) := x"FFEA";
          m(642) := x"FFE5";
          m(643) := x"0019";
          m(644) := x"0002";
          m(645) := x"FFFA";
          m(646) := x"FFF9";
          m(647) := x"FECE";
          m(648) := x"FF54";
          m(649) := x"0105";
          m(650) := x"0377";
          m(651) := x"027D";
          m(652) := x"01D8";
          m(653) := x"0539";
          m(654) := x"0089";
          m(655) := x"01F3";
          m(656) := x"0045";
          m(657) := x"0229";
          m(658) := x"005E";
          m(659) := x"041E";
          m(660) := x"0023";
          m(661) := x"00B3";
          m(662) := x"004F";
          m(663) := x"FFA1";
          m(664) := x"FCFC";
          m(665) := x"0196";
          m(666) := x"FE4E";
          m(667) := x"FEB7";
          m(668) := x"FEAB";
          m(669) := x"0025";
          m(670) := x"0016";
          m(671) := x"FFB8";
          m(672) := x"FFE8";
          m(673) := x"FFE6";
          m(674) := x"FF9A";
          m(675) := x"FF8D";
          m(676) := x"00A4";
          m(677) := x"028D";
          m(678) := x"02C9";
          m(679) := x"FFD2";
          m(680) := x"02CC";
          m(681) := x"0057";
          m(682) := x"FC82";
          m(683) := x"00DB";
          m(684) := x"02F1";
          m(685) := x"FE49";
          m(686) := x"FBEB";
          m(687) := x"002A";
          m(688) := x"FFC1";
          m(689) := x"0358";
          m(690) := x"0143";
          m(691) := x"012E";
          m(692) := x"FF6E";
          m(693) := x"01F6";
          m(694) := x"FF83";
          m(695) := x"FE16";
          m(696) := x"FF71";
          m(697) := x"001B";
          m(698) := x"FFD9";
          m(699) := x"FFE4";
          m(700) := x"0016";
          m(701) := x"0017";
          m(702) := x"0024";
          m(703) := x"0001";
          m(704) := x"001A";
          m(705) := x"FF8B";
          m(706) := x"FF57";
          m(707) := x"0000";
          m(708) := x"004F";
          m(709) := x"0403";
          m(710) := x"00F1";
          m(711) := x"0170";
          m(712) := x"08D9";
          m(713) := x"FF9D";
          m(714) := x"02C3";
          m(715) := x"037B";
          m(716) := x"0251";
          m(717) := x"00E5";
          m(718) := x"07B7";
          m(719) := x"067E";
          m(720) := x"FF8B";
          m(721) := x"FE47";
          m(722) := x"FF56";
          m(723) := x"FF55";
          m(724) := x"0008";
          m(725) := x"FFAC";
          m(726) := x"FFE3";
          m(727) := x"FFC8";
          m(728) := x"FFF0";
          m(729) := x"0019";
          m(730) := x"FFFF";
          m(731) := x"FFE3";
          m(732) := x"FDD3";
          m(733) := x"FDB4";
          m(734) := x"FE43";
          m(735) := x"FEDF";
          m(736) := x"0194";
          m(737) := x"0177";
          m(738) := x"00F9";
          m(739) := x"0385";
          m(740) := x"0181";
          m(741) := x"FD06";
          m(742) := x"FF87";
          m(743) := x"0007";
          m(744) := x"0123";
          m(745) := x"FF22";
          m(746) := x"056E";
          m(747) := x"05F4";
          m(748) := x"0206";
          m(749) := x"00D4";
          m(750) := x"0036";
          m(751) := x"FFEC";
          m(752) := x"001A";
          m(753) := x"FFD2";
          m(754) := x"FFD3";
          m(755) := x"002A";
          m(756) := x"003F";
          m(757) := x"FFFF";
          m(758) := x"FFC8";
          m(759) := x"0004";
          m(760) := x"0030";
          m(761) := x"FFF2";
          m(762) := x"0041";
          m(763) := x"002D";
          m(764) := x"0002";
          m(765) := x"0001";
          m(766) := x"000F";
          m(767) := x"FF5F";
          m(768) := x"FEF9";
          m(769) := x"0070";
          m(770) := x"0072";
          m(771) := x"FD76";
          m(772) := x"FD94";
          m(773) := x"FFD5";
          m(774) := x"FF80";
          m(775) := x"0096";
          m(776) := x"0015";
          m(777) := x"FF94";
          m(778) := x"0069";
          m(779) := x"0023";
          m(780) := x"FFF9";
          m(781) := x"0007";
          m(782) := x"FFE4";
          m(783) := x"0038";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_2.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 2) then
          m(0) := x"FFF1";
          m(1) := x"FFD8";
          m(2) := x"0010";
          m(3) := x"FFAB";
          m(4) := x"002B";
          m(5) := x"0000";
          m(6) := x"001E";
          m(7) := x"FFF6";
          m(8) := x"FFCD";
          m(9) := x"FFD1";
          m(10) := x"0051";
          m(11) := x"FFFC";
          m(12) := x"000F";
          m(13) := x"FFFE";
          m(14) := x"0014";
          m(15) := x"0035";
          m(16) := x"0003";
          m(17) := x"0038";
          m(18) := x"FFD1";
          m(19) := x"000D";
          m(20) := x"FFFD";
          m(21) := x"0012";
          m(22) := x"FFFC";
          m(23) := x"FFF2";
          m(24) := x"FFF4";
          m(25) := x"0000";
          m(26) := x"002A";
          m(27) := x"FFEA";
          m(28) := x"FFE5";
          m(29) := x"000A";
          m(30) := x"FFFC";
          m(31) := x"FFD5";
          m(32) := x"0026";
          m(33) := x"FFED";
          m(34) := x"FFDF";
          m(35) := x"FFE7";
          m(36) := x"FFF2";
          m(37) := x"FFFC";
          m(38) := x"FFEA";
          m(39) := x"0029";
          m(40) := x"FFDA";
          m(41) := x"0008";
          m(42) := x"FFE6";
          m(43) := x"008C";
          m(44) := x"0002";
          m(45) := x"0000";
          m(46) := x"0010";
          m(47) := x"FFEB";
          m(48) := x"FFED";
          m(49) := x"FFF1";
          m(50) := x"FFFC";
          m(51) := x"FFFF";
          m(52) := x"FFF6";
          m(53) := x"0003";
          m(54) := x"FFFF";
          m(55) := x"0015";
          m(56) := x"FFDA";
          m(57) := x"0043";
          m(58) := x"FFF6";
          m(59) := x"FFEF";
          m(60) := x"FFF3";
          m(61) := x"FFDF";
          m(62) := x"0008";
          m(63) := x"0019";
          m(64) := x"FF9F";
          m(65) := x"FF6E";
          m(66) := x"FFD2";
          m(67) := x"FF96";
          m(68) := x"FFB8";
          m(69) := x"005A";
          m(70) := x"00A4";
          m(71) := x"032B";
          m(72) := x"0276";
          m(73) := x"002A";
          m(74) := x"FFC1";
          m(75) := x"FFBB";
          m(76) := x"FFC2";
          m(77) := x"FFBC";
          m(78) := x"FFE9";
          m(79) := x"FFB0";
          m(80) := x"FFEF";
          m(81) := x"001D";
          m(82) := x"FFCE";
          m(83) := x"001B";
          m(84) := x"FFE2";
          m(85) := x"FFF1";
          m(86) := x"FFC8";
          m(87) := x"FFC6";
          m(88) := x"004B";
          m(89) := x"FF68";
          m(90) := x"FFC7";
          m(91) := x"0004";
          m(92) := x"FFC4";
          m(93) := x"FEE2";
          m(94) := x"FE52";
          m(95) := x"FCE1";
          m(96) := x"FFBF";
          m(97) := x"FF4D";
          m(98) := x"FB2E";
          m(99) := x"FF6F";
          m(100) := x"01DC";
          m(101) := x"0076";
          m(102) := x"FEEB";
          m(103) := x"FEC3";
          m(104) := x"FF0B";
          m(105) := x"FE81";
          m(106) := x"FFE8";
          m(107) := x"0049";
          m(108) := x"00F5";
          m(109) := x"01E3";
          m(110) := x"0011";
          m(111) := x"000F";
          m(112) := x"002C";
          m(113) := x"FFEE";
          m(114) := x"FFF5";
          m(115) := x"0013";
          m(116) := x"0017";
          m(117) := x"FF8D";
          m(118) := x"FF4A";
          m(119) := x"FE6B";
          m(120) := x"FDC8";
          m(121) := x"FCD4";
          m(122) := x"FB7F";
          m(123) := x"FD24";
          m(124) := x"FDAC";
          m(125) := x"FEE5";
          m(126) := x"FB32";
          m(127) := x"FE89";
          m(128) := x"FDD5";
          m(129) := x"FDA8";
          m(130) := x"FC8E";
          m(131) := x"FC87";
          m(132) := x"000C";
          m(133) := x"0175";
          m(134) := x"0029";
          m(135) := x"030B";
          m(136) := x"03C4";
          m(137) := x"00B8";
          m(138) := x"FF2C";
          m(139) := x"FFAB";
          m(140) := x"FFE4";
          m(141) := x"001C";
          m(142) := x"FFE0";
          m(143) := x"0002";
          m(144) := x"FFFB";
          m(145) := x"FFE5";
          m(146) := x"FE7E";
          m(147) := x"FCB6";
          m(148) := x"FB5B";
          m(149) := x"FAC3";
          m(150) := x"F94C";
          m(151) := x"FC12";
          m(152) := x"FCFE";
          m(153) := x"FF82";
          m(154) := x"FBA9";
          m(155) := x"009C";
          m(156) := x"FEFA";
          m(157) := x"FB78";
          m(158) := x"FA82";
          m(159) := x"FE01";
          m(160) := x"03B2";
          m(161) := x"FCAF";
          m(162) := x"FFE5";
          m(163) := x"0449";
          m(164) := x"0394";
          m(165) := x"FED2";
          m(166) := x"FFAF";
          m(167) := x"FFD1";
          m(168) := x"003F";
          m(169) := x"FFE7";
          m(170) := x"001E";
          m(171) := x"001E";
          m(172) := x"FFBF";
          m(173) := x"FF68";
          m(174) := x"FD5A";
          m(175) := x"F900";
          m(176) := x"F5D4";
          m(177) := x"F864";
          m(178) := x"FDC9";
          m(179) := x"FDD6";
          m(180) := x"00EF";
          m(181) := x"00EB";
          m(182) := x"0129";
          m(183) := x"FB3F";
          m(184) := x"FBB2";
          m(185) := x"FD92";
          m(186) := x"FE79";
          m(187) := x"0358";
          m(188) := x"0520";
          m(189) := x"0136";
          m(190) := x"0139";
          m(191) := x"0537";
          m(192) := x"04AC";
          m(193) := x"FF70";
          m(194) := x"014B";
          m(195) := x"006C";
          m(196) := x"0005";
          m(197) := x"0018";
          m(198) := x"FFEE";
          m(199) := x"0064";
          m(200) := x"0015";
          m(201) := x"FED7";
          m(202) := x"FCFC";
          m(203) := x"FB70";
          m(204) := x"FA32";
          m(205) := x"FD31";
          m(206) := x"013C";
          m(207) := x"FBD6";
          m(208) := x"052D";
          m(209) := x"FAB1";
          m(210) := x"FD3A";
          m(211) := x"FC44";
          m(212) := x"FDCA";
          m(213) := x"FE65";
          m(214) := x"FCE7";
          m(215) := x"FCAE";
          m(216) := x"0497";
          m(217) := x"01D8";
          m(218) := x"0234";
          m(219) := x"02E3";
          m(220) := x"028F";
          m(221) := x"0026";
          m(222) := x"0360";
          m(223) := x"003C";
          m(224) := x"0048";
          m(225) := x"0003";
          m(226) := x"FFD1";
          m(227) := x"0042";
          m(228) := x"FF87";
          m(229) := x"FDF1";
          m(230) := x"FDDD";
          m(231) := x"FDFC";
          m(232) := x"FD8C";
          m(233) := x"FF73";
          m(234) := x"FB1F";
          m(235) := x"FC4E";
          m(236) := x"01CA";
          m(237) := x"0127";
          m(238) := x"0165";
          m(239) := x"01B6";
          m(240) := x"00A7";
          m(241) := x"FEE4";
          m(242) := x"FF70";
          m(243) := x"FF61";
          m(244) := x"02C8";
          m(245) := x"0571";
          m(246) := x"0483";
          m(247) := x"FFA7";
          m(248) := x"066A";
          m(249) := x"0660";
          m(250) := x"01F1";
          m(251) := x"001C";
          m(252) := x"0035";
          m(253) := x"0016";
          m(254) := x"FFC9";
          m(255) := x"0011";
          m(256) := x"FFA8";
          m(257) := x"FE55";
          m(258) := x"00B8";
          m(259) := x"FFAF";
          m(260) := x"FC31";
          m(261) := x"FC35";
          m(262) := x"00E6";
          m(263) := x"0091";
          m(264) := x"FDE3";
          m(265) := x"03A8";
          m(266) := x"05A9";
          m(267) := x"02DE";
          m(268) := x"0022";
          m(269) := x"02FB";
          m(270) := x"0396";
          m(271) := x"0142";
          m(272) := x"0157";
          m(273) := x"0520";
          m(274) := x"0399";
          m(275) := x"FE61";
          m(276) := x"0881";
          m(277) := x"061C";
          m(278) := x"FFF2";
          m(279) := x"003D";
          m(280) := x"FFED";
          m(281) := x"FFE0";
          m(282) := x"001F";
          m(283) := x"0024";
          m(284) := x"FF98";
          m(285) := x"FEEA";
          m(286) := x"FEEB";
          m(287) := x"00C6";
          m(288) := x"FBA7";
          m(289) := x"FD8B";
          m(290) := x"0125";
          m(291) := x"FC99";
          m(292) := x"FCB0";
          m(293) := x"0293";
          m(294) := x"0205";
          m(295) := x"04A4";
          m(296) := x"FCC4";
          m(297) := x"FC28";
          m(298) := x"0079";
          m(299) := x"02C2";
          m(300) := x"0100";
          m(301) := x"027C";
          m(302) := x"0367";
          m(303) := x"0432";
          m(304) := x"09E6";
          m(305) := x"088F";
          m(306) := x"0199";
          m(307) := x"0007";
          m(308) := x"0016";
          m(309) := x"0016";
          m(310) := x"0010";
          m(311) := x"0037";
          m(312) := x"0018";
          m(313) := x"FF49";
          m(314) := x"FCD0";
          m(315) := x"FD3F";
          m(316) := x"FB48";
          m(317) := x"FB4C";
          m(318) := x"FC4E";
          m(319) := x"FD15";
          m(320) := x"FC82";
          m(321) := x"FAAB";
          m(322) := x"FF95";
          m(323) := x"FB31";
          m(324) := x"FA0B";
          m(325) := x"F7F6";
          m(326) := x"F931";
          m(327) := x"FB56";
          m(328) := x"FEF0";
          m(329) := x"00A7";
          m(330) := x"FF68";
          m(331) := x"0171";
          m(332) := x"026E";
          m(333) := x"05FF";
          m(334) := x"01BE";
          m(335) := x"FFC3";
          m(336) := x"FFF5";
          m(337) := x"FFCE";
          m(338) := x"FFF8";
          m(339) := x"000E";
          m(340) := x"FEBB";
          m(341) := x"FD9A";
          m(342) := x"FCB6";
          m(343) := x"FD7E";
          m(344) := x"FE2D";
          m(345) := x"01FA";
          m(346) := x"00EF";
          m(347) := x"FE7A";
          m(348) := x"001D";
          m(349) := x"FFB2";
          m(350) := x"FD24";
          m(351) := x"F748";
          m(352) := x"F52D";
          m(353) := x"F03E";
          m(354) := x"EB98";
          m(355) := x"EE88";
          m(356) := x"F70F";
          m(357) := x"F717";
          m(358) := x"F9CA";
          m(359) := x"F934";
          m(360) := x"FA7E";
          m(361) := x"0051";
          m(362) := x"007F";
          m(363) := x"0030";
          m(364) := x"0009";
          m(365) := x"0005";
          m(366) := x"FFF4";
          m(367) := x"FFD7";
          m(368) := x"FE5A";
          m(369) := x"FE06";
          m(370) := x"FD2D";
          m(371) := x"FF6F";
          m(372) := x"026A";
          m(373) := x"012A";
          m(374) := x"0179";
          m(375) := x"FFC0";
          m(376) := x"011E";
          m(377) := x"FFC5";
          m(378) := x"040B";
          m(379) := x"F97C";
          m(380) := x"FE0C";
          m(381) := x"F8BE";
          m(382) := x"F22B";
          m(383) := x"F122";
          m(384) := x"F562";
          m(385) := x"F534";
          m(386) := x"F5ED";
          m(387) := x"F7B7";
          m(388) := x"F9A0";
          m(389) := x"FE75";
          m(390) := x"0002";
          m(391) := x"FFD5";
          m(392) := x"FFE3";
          m(393) := x"0025";
          m(394) := x"004C";
          m(395) := x"0053";
          m(396) := x"FFEF";
          m(397) := x"FF6E";
          m(398) := x"FD57";
          m(399) := x"FE6C";
          m(400) := x"FD5A";
          m(401) := x"01C1";
          m(402) := x"FDF3";
          m(403) := x"F977";
          m(404) := x"FC80";
          m(405) := x"FA76";
          m(406) := x"FCCE";
          m(407) := x"0039";
          m(408) := x"FE98";
          m(409) := x"FF9E";
          m(410) := x"FD4C";
          m(411) := x"F501";
          m(412) := x"F7A4";
          m(413) := x"F94F";
          m(414) := x"F8A8";
          m(415) := x"F8AC";
          m(416) := x"FA32";
          m(417) := x"FE8E";
          m(418) := x"0000";
          m(419) := x"FFCA";
          m(420) := x"FFDA";
          m(421) := x"FFFE";
          m(422) := x"0020";
          m(423) := x"FFCF";
          m(424) := x"005B";
          m(425) := x"0276";
          m(426) := x"046E";
          m(427) := x"01AD";
          m(428) := x"FF9C";
          m(429) := x"0409";
          m(430) := x"FF88";
          m(431) := x"FB34";
          m(432) := x"04E6";
          m(433) := x"FE80";
          m(434) := x"FFE5";
          m(435) := x"FFC8";
          m(436) := x"FDEC";
          m(437) := x"FC04";
          m(438) := x"FFC4";
          m(439) := x"F988";
          m(440) := x"F995";
          m(441) := x"FABE";
          m(442) := x"F8B7";
          m(443) := x"FAAC";
          m(444) := x"FB8A";
          m(445) := x"FF3F";
          m(446) := x"000B";
          m(447) := x"FFDC";
          m(448) := x"0008";
          m(449) := x"0012";
          m(450) := x"0027";
          m(451) := x"0008";
          m(452) := x"FF34";
          m(453) := x"02E5";
          m(454) := x"0238";
          m(455) := x"FEBC";
          m(456) := x"009E";
          m(457) := x"FB44";
          m(458) := x"FBE4";
          m(459) := x"FF5B";
          m(460) := x"0110";
          m(461) := x"0025";
          m(462) := x"FDE7";
          m(463) := x"FD94";
          m(464) := x"FB63";
          m(465) := x"FF21";
          m(466) := x"FDBF";
          m(467) := x"FCD1";
          m(468) := x"FC65";
          m(469) := x"FBAD";
          m(470) := x"FAC1";
          m(471) := x"FB02";
          m(472) := x"FC8A";
          m(473) := x"FF67";
          m(474) := x"FFEF";
          m(475) := x"FFD7";
          m(476) := x"FFE8";
          m(477) := x"FFF8";
          m(478) := x"FFCA";
          m(479) := x"0067";
          m(480) := x"0059";
          m(481) := x"0182";
          m(482) := x"FFD1";
          m(483) := x"009F";
          m(484) := x"FFDD";
          m(485) := x"0055";
          m(486) := x"FCEE";
          m(487) := x"FB7F";
          m(488) := x"FD33";
          m(489) := x"FF87";
          m(490) := x"04F2";
          m(491) := x"0379";
          m(492) := x"FEFE";
          m(493) := x"01CC";
          m(494) := x"FF8E";
          m(495) := x"FE06";
          m(496) := x"FEEC";
          m(497) := x"FB33";
          m(498) := x"FC50";
          m(499) := x"FD7F";
          m(500) := x"FDA7";
          m(501) := x"FF2A";
          m(502) := x"FFC1";
          m(503) := x"FFCF";
          m(504) := x"001F";
          m(505) := x"FFDA";
          m(506) := x"FFCF";
          m(507) := x"FF60";
          m(508) := x"00FF";
          m(509) := x"FD5D";
          m(510) := x"FFDD";
          m(511) := x"FEE3";
          m(512) := x"0036";
          m(513) := x"FD1C";
          m(514) := x"FE8D";
          m(515) := x"FF0C";
          m(516) := x"FE11";
          m(517) := x"FF44";
          m(518) := x"033A";
          m(519) := x"0089";
          m(520) := x"FEAD";
          m(521) := x"01C0";
          m(522) := x"FE5C";
          m(523) := x"038B";
          m(524) := x"0225";
          m(525) := x"FB9D";
          m(526) := x"FB54";
          m(527) := x"FB86";
          m(528) := x"FDA9";
          m(529) := x"0005";
          m(530) := x"FFDD";
          m(531) := x"FFD5";
          m(532) := x"0024";
          m(533) := x"FFEF";
          m(534) := x"FFFB";
          m(535) := x"FECD";
          m(536) := x"FF2B";
          m(537) := x"01C0";
          m(538) := x"0329";
          m(539) := x"FFCA";
          m(540) := x"0165";
          m(541) := x"FE9E";
          m(542) := x"FE97";
          m(543) := x"010A";
          m(544) := x"0070";
          m(545) := x"054F";
          m(546) := x"0537";
          m(547) := x"0427";
          m(548) := x"0571";
          m(549) := x"00F5";
          m(550) := x"FC0C";
          m(551) := x"047A";
          m(552) := x"0173";
          m(553) := x"FAEA";
          m(554) := x"FD3B";
          m(555) := x"FF5E";
          m(556) := x"0029";
          m(557) := x"00BE";
          m(558) := x"FFD5";
          m(559) := x"001E";
          m(560) := x"FFE5";
          m(561) := x"0010";
          m(562) := x"FFF3";
          m(563) := x"FE0E";
          m(564) := x"FBF0";
          m(565) := x"0071";
          m(566) := x"032E";
          m(567) := x"005F";
          m(568) := x"0372";
          m(569) := x"FF45";
          m(570) := x"FFAA";
          m(571) := x"013F";
          m(572) := x"0207";
          m(573) := x"00A9";
          m(574) := x"FE84";
          m(575) := x"FF52";
          m(576) := x"02A4";
          m(577) := x"03AC";
          m(578) := x"0179";
          m(579) := x"07E1";
          m(580) := x"00AE";
          m(581) := x"F9F9";
          m(582) := x"FEAB";
          m(583) := x"FF9F";
          m(584) := x"00EF";
          m(585) := x"0052";
          m(586) := x"0010";
          m(587) := x"0031";
          m(588) := x"0017";
          m(589) := x"000E";
          m(590) := x"FFE3";
          m(591) := x"FD6D";
          m(592) := x"FCE0";
          m(593) := x"FF55";
          m(594) := x"FE0D";
          m(595) := x"FF57";
          m(596) := x"02EF";
          m(597) := x"FF08";
          m(598) := x"FFFD";
          m(599) := x"01E0";
          m(600) := x"FF40";
          m(601) := x"0010";
          m(602) := x"0108";
          m(603) := x"06D9";
          m(604) := x"FC9A";
          m(605) := x"0125";
          m(606) := x"0200";
          m(607) := x"04D5";
          m(608) := x"03EA";
          m(609) := x"FD54";
          m(610) := x"FE85";
          m(611) := x"FE3C";
          m(612) := x"FF4B";
          m(613) := x"FFB6";
          m(614) := x"0015";
          m(615) := x"FFD8";
          m(616) := x"FFEA";
          m(617) := x"FFE5";
          m(618) := x"FFF7";
          m(619) := x"FF28";
          m(620) := x"FE1E";
          m(621) := x"FDF6";
          m(622) := x"FF51";
          m(623) := x"FBCB";
          m(624) := x"FF29";
          m(625) := x"020D";
          m(626) := x"00C0";
          m(627) := x"0297";
          m(628) := x"024E";
          m(629) := x"FF76";
          m(630) := x"01A4";
          m(631) := x"00E9";
          m(632) := x"0009";
          m(633) := x"0508";
          m(634) := x"023A";
          m(635) := x"01B6";
          m(636) := x"02A6";
          m(637) := x"0116";
          m(638) := x"FF2C";
          m(639) := x"FF59";
          m(640) := x"FFDC";
          m(641) := x"FFEF";
          m(642) := x"FFF3";
          m(643) := x"001D";
          m(644) := x"0026";
          m(645) := x"0032";
          m(646) := x"FFDD";
          m(647) := x"0041";
          m(648) := x"00BC";
          m(649) := x"FF0B";
          m(650) := x"FD50";
          m(651) := x"FC30";
          m(652) := x"FF36";
          m(653) := x"FFA4";
          m(654) := x"FFD1";
          m(655) := x"013A";
          m(656) := x"FF83";
          m(657) := x"FAED";
          m(658) := x"02B7";
          m(659) := x"01B3";
          m(660) := x"0173";
          m(661) := x"FFDB";
          m(662) := x"00AC";
          m(663) := x"0052";
          m(664) := x"018B";
          m(665) := x"003E";
          m(666) := x"FEDE";
          m(667) := x"FF36";
          m(668) := x"FFFC";
          m(669) := x"FFD4";
          m(670) := x"FFD1";
          m(671) := x"FFFE";
          m(672) := x"0025";
          m(673) := x"FFE1";
          m(674) := x"0016";
          m(675) := x"0024";
          m(676) := x"FF8D";
          m(677) := x"FE40";
          m(678) := x"FE66";
          m(679) := x"FFD3";
          m(680) := x"00A4";
          m(681) := x"0259";
          m(682) := x"0094";
          m(683) := x"FF10";
          m(684) := x"FEEC";
          m(685) := x"011C";
          m(686) := x"00EB";
          m(687) := x"FD9E";
          m(688) := x"FE3C";
          m(689) := x"0348";
          m(690) := x"02A7";
          m(691) := x"FFDF";
          m(692) := x"FFD4";
          m(693) := x"FEEA";
          m(694) := x"FFBA";
          m(695) := x"0012";
          m(696) := x"FFFB";
          m(697) := x"FF7C";
          m(698) := x"FFF2";
          m(699) := x"FFF5";
          m(700) := x"FFEA";
          m(701) := x"FFAA";
          m(702) := x"0030";
          m(703) := x"FFF3";
          m(704) := x"FF3D";
          m(705) := x"FF10";
          m(706) := x"FE12";
          m(707) := x"FE12";
          m(708) := x"FDFA";
          m(709) := x"FFBF";
          m(710) := x"FF87";
          m(711) := x"0154";
          m(712) := x"040B";
          m(713) := x"035B";
          m(714) := x"FD90";
          m(715) := x"FCD3";
          m(716) := x"0116";
          m(717) := x"0427";
          m(718) := x"01BE";
          m(719) := x"01EB";
          m(720) := x"008F";
          m(721) := x"006E";
          m(722) := x"0044";
          m(723) := x"0044";
          m(724) := x"FFE2";
          m(725) := x"FFD3";
          m(726) := x"FFF9";
          m(727) := x"001E";
          m(728) := x"0006";
          m(729) := x"0018";
          m(730) := x"0023";
          m(731) := x"0035";
          m(732) := x"FFBF";
          m(733) := x"0003";
          m(734) := x"003E";
          m(735) := x"000A";
          m(736) := x"FEC7";
          m(737) := x"FE5B";
          m(738) := x"FFAF";
          m(739) := x"0140";
          m(740) := x"0362";
          m(741) := x"01AF";
          m(742) := x"FEA3";
          m(743) := x"FF70";
          m(744) := x"019D";
          m(745) := x"FF5E";
          m(746) := x"FF45";
          m(747) := x"0064";
          m(748) := x"0075";
          m(749) := x"0086";
          m(750) := x"0014";
          m(751) := x"FFF0";
          m(752) := x"FFF0";
          m(753) := x"0023";
          m(754) := x"0001";
          m(755) := x"0001";
          m(756) := x"FFEB";
          m(757) := x"0009";
          m(758) := x"0028";
          m(759) := x"000E";
          m(760) := x"0000";
          m(761) := x"FFC6";
          m(762) := x"000A";
          m(763) := x"0047";
          m(764) := x"FFDE";
          m(765) := x"0000";
          m(766) := x"FFE4";
          m(767) := x"FFCE";
          m(768) := x"0008";
          m(769) := x"FFF3";
          m(770) := x"001A";
          m(771) := x"FFE0";
          m(772) := x"0018";
          m(773) := x"FFDE";
          m(774) := x"FF7E";
          m(775) := x"FFE1";
          m(776) := x"000B";
          m(777) := x"FFF5";
          m(778) := x"0042";
          m(779) := x"0004";
          m(780) := x"FFF7";
          m(781) := x"001C";
          m(782) := x"0042";
          m(783) := x"FFB9";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_3.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 3) then
          m(0) := x"0006";
          m(1) := x"001E";
          m(2) := x"0019";
          m(3) := x"FFFB";
          m(4) := x"FFE2";
          m(5) := x"FFD9";
          m(6) := x"000F";
          m(7) := x"0017";
          m(8) := x"000E";
          m(9) := x"FFF6";
          m(10) := x"FFE7";
          m(11) := x"FFED";
          m(12) := x"FFEB";
          m(13) := x"0020";
          m(14) := x"000B";
          m(15) := x"000B";
          m(16) := x"FFCF";
          m(17) := x"000B";
          m(18) := x"0010";
          m(19) := x"FFE6";
          m(20) := x"003B";
          m(21) := x"0006";
          m(22) := x"FFD7";
          m(23) := x"0018";
          m(24) := x"002B";
          m(25) := x"000C";
          m(26) := x"FFF2";
          m(27) := x"FFFB";
          m(28) := x"FFEC";
          m(29) := x"FFEF";
          m(30) := x"FFED";
          m(31) := x"FFFB";
          m(32) := x"002F";
          m(33) := x"0037";
          m(34) := x"0031";
          m(35) := x"0019";
          m(36) := x"FFED";
          m(37) := x"0011";
          m(38) := x"0015";
          m(39) := x"0036";
          m(40) := x"004A";
          m(41) := x"0010";
          m(42) := x"00A6";
          m(43) := x"0135";
          m(44) := x"012B";
          m(45) := x"00B6";
          m(46) := x"FFF5";
          m(47) := x"002A";
          m(48) := x"002E";
          m(49) := x"FFEF";
          m(50) := x"0010";
          m(51) := x"0003";
          m(52) := x"0003";
          m(53) := x"FFF7";
          m(54) := x"000A";
          m(55) := x"001F";
          m(56) := x"0007";
          m(57) := x"FFE7";
          m(58) := x"FFF3";
          m(59) := x"FFFC";
          m(60) := x"0004";
          m(61) := x"0000";
          m(62) := x"FFDF";
          m(63) := x"002B";
          m(64) := x"0016";
          m(65) := x"0026";
          m(66) := x"0013";
          m(67) := x"FEAA";
          m(68) := x"FE4B";
          m(69) := x"FD77";
          m(70) := x"FF50";
          m(71) := x"0032";
          m(72) := x"0000";
          m(73) := x"01AE";
          m(74) := x"0020";
          m(75) := x"0078";
          m(76) := x"FFDE";
          m(77) := x"001C";
          m(78) := x"0039";
          m(79) := x"0048";
          m(80) := x"0002";
          m(81) := x"0003";
          m(82) := x"FFD0";
          m(83) := x"0020";
          m(84) := x"FFDB";
          m(85) := x"FFF0";
          m(86) := x"0043";
          m(87) := x"0022";
          m(88) := x"FFF2";
          m(89) := x"0047";
          m(90) := x"0062";
          m(91) := x"0007";
          m(92) := x"011B";
          m(93) := x"0157";
          m(94) := x"0290";
          m(95) := x"FEA1";
          m(96) := x"FDA9";
          m(97) := x"FD8D";
          m(98) := x"FB2C";
          m(99) := x"FAAD";
          m(100) := x"FCA0";
          m(101) := x"FE8F";
          m(102) := x"FDE3";
          m(103) := x"FF28";
          m(104) := x"FF90";
          m(105) := x"0163";
          m(106) := x"01F0";
          m(107) := x"0165";
          m(108) := x"00D1";
          m(109) := x"0057";
          m(110) := x"0034";
          m(111) := x"0026";
          m(112) := x"FFA4";
          m(113) := x"003C";
          m(114) := x"0000";
          m(115) := x"0019";
          m(116) := x"0010";
          m(117) := x"FFD1";
          m(118) := x"0045";
          m(119) := x"002B";
          m(120) := x"01C0";
          m(121) := x"0400";
          m(122) := x"03C2";
          m(123) := x"04D4";
          m(124) := x"0185";
          m(125) := x"0185";
          m(126) := x"00F4";
          m(127) := x"F910";
          m(128) := x"F97E";
          m(129) := x"FDE6";
          m(130) := x"01EA";
          m(131) := x"FDE1";
          m(132) := x"F98A";
          m(133) := x"017A";
          m(134) := x"02A4";
          m(135) := x"04A3";
          m(136) := x"0362";
          m(137) := x"016B";
          m(138) := x"0011";
          m(139) := x"0040";
          m(140) := x"000A";
          m(141) := x"0001";
          m(142) := x"002E";
          m(143) := x"0016";
          m(144) := x"0042";
          m(145) := x"013C";
          m(146) := x"01F2";
          m(147) := x"03FA";
          m(148) := x"021C";
          m(149) := x"0250";
          m(150) := x"04B4";
          m(151) := x"04FE";
          m(152) := x"02F3";
          m(153) := x"03CE";
          m(154) := x"0139";
          m(155) := x"FD59";
          m(156) := x"F847";
          m(157) := x"03BC";
          m(158) := x"FA1E";
          m(159) := x"00CD";
          m(160) := x"FC31";
          m(161) := x"FE54";
          m(162) := x"007F";
          m(163) := x"013C";
          m(164) := x"024A";
          m(165) := x"012E";
          m(166) := x"00A1";
          m(167) := x"0055";
          m(168) := x"FFFC";
          m(169) := x"FFD5";
          m(170) := x"0072";
          m(171) := x"0036";
          m(172) := x"0073";
          m(173) := x"FF8F";
          m(174) := x"FEB8";
          m(175) := x"0175";
          m(176) := x"0016";
          m(177) := x"0094";
          m(178) := x"FF6C";
          m(179) := x"06B8";
          m(180) := x"03A5";
          m(181) := x"05F2";
          m(182) := x"0178";
          m(183) := x"0070";
          m(184) := x"FCC9";
          m(185) := x"FD70";
          m(186) := x"FCD7";
          m(187) := x"02B2";
          m(188) := x"FFB9";
          m(189) := x"FF8B";
          m(190) := x"00DA";
          m(191) := x"0450";
          m(192) := x"02DA";
          m(193) := x"00E7";
          m(194) := x"FFD2";
          m(195) := x"FFE4";
          m(196) := x"001F";
          m(197) := x"FFB8";
          m(198) := x"0031";
          m(199) := x"FED0";
          m(200) := x"FE9C";
          m(201) := x"FE1F";
          m(202) := x"FEA9";
          m(203) := x"009F";
          m(204) := x"00DC";
          m(205) := x"000D";
          m(206) := x"01F3";
          m(207) := x"05E8";
          m(208) := x"0314";
          m(209) := x"01A6";
          m(210) := x"03AB";
          m(211) := x"0117";
          m(212) := x"FC67";
          m(213) := x"FF4D";
          m(214) := x"FD80";
          m(215) := x"FA77";
          m(216) := x"FA34";
          m(217) := x"F9DB";
          m(218) := x"FC7C";
          m(219) := x"038B";
          m(220) := x"0603";
          m(221) := x"03B2";
          m(222) := x"FFC7";
          m(223) := x"FFE9";
          m(224) := x"FFF0";
          m(225) := x"000E";
          m(226) := x"FFF2";
          m(227) := x"FEF5";
          m(228) := x"FCBC";
          m(229) := x"FB91";
          m(230) := x"00C2";
          m(231) := x"FCD0";
          m(232) := x"FFE1";
          m(233) := x"01EB";
          m(234) := x"FE56";
          m(235) := x"01B7";
          m(236) := x"01DC";
          m(237) := x"08CB";
          m(238) := x"019B";
          m(239) := x"FAA9";
          m(240) := x"FFD4";
          m(241) := x"FD8E";
          m(242) := x"FC5F";
          m(243) := x"FBD6";
          m(244) := x"FFA3";
          m(245) := x"FF84";
          m(246) := x"FB99";
          m(247) := x"0362";
          m(248) := x"090C";
          m(249) := x"037D";
          m(250) := x"0006";
          m(251) := x"0034";
          m(252) := x"0025";
          m(253) := x"003D";
          m(254) := x"0023";
          m(255) := x"00C0";
          m(256) := x"FBD3";
          m(257) := x"F9AD";
          m(258) := x"FD0B";
          m(259) := x"FED8";
          m(260) := x"00DF";
          m(261) := x"FE42";
          m(262) := x"FC41";
          m(263) := x"06FA";
          m(264) := x"FFB4";
          m(265) := x"0755";
          m(266) := x"0543";
          m(267) := x"F6E0";
          m(268) := x"F2C5";
          m(269) := x"FB2C";
          m(270) := x"0114";
          m(271) := x"FFB7";
          m(272) := x"00AC";
          m(273) := x"FF3F";
          m(274) := x"FF08";
          m(275) := x"0340";
          m(276) := x"0800";
          m(277) := x"025D";
          m(278) := x"FFCA";
          m(279) := x"0018";
          m(280) := x"0009";
          m(281) := x"FFF3";
          m(282) := x"002C";
          m(283) := x"00BF";
          m(284) := x"FDD7";
          m(285) := x"FD03";
          m(286) := x"FA57";
          m(287) := x"FCF8";
          m(288) := x"FAB1";
          m(289) := x"FB22";
          m(290) := x"FA2B";
          m(291) := x"04CF";
          m(292) := x"FE13";
          m(293) := x"05E6";
          m(294) := x"03B4";
          m(295) := x"F596";
          m(296) := x"FC49";
          m(297) := x"FD0F";
          m(298) := x"0122";
          m(299) := x"FAC4";
          m(300) := x"FE35";
          m(301) := x"017E";
          m(302) := x"02CA";
          m(303) := x"050D";
          m(304) := x"04FA";
          m(305) := x"013C";
          m(306) := x"FFD9";
          m(307) := x"0029";
          m(308) := x"FFC4";
          m(309) := x"0018";
          m(310) := x"0061";
          m(311) := x"0144";
          m(312) := x"0128";
          m(313) := x"FE5C";
          m(314) := x"FBDB";
          m(315) := x"FA78";
          m(316) := x"0080";
          m(317) := x"FD33";
          m(318) := x"FB73";
          m(319) := x"FF6E";
          m(320) := x"0607";
          m(321) := x"0F7A";
          m(322) := x"0999";
          m(323) := x"FA1E";
          m(324) := x"FD64";
          m(325) := x"FC7F";
          m(326) := x"FC0A";
          m(327) := x"F9ED";
          m(328) := x"FC03";
          m(329) := x"019C";
          m(330) := x"0477";
          m(331) := x"0329";
          m(332) := x"028B";
          m(333) := x"FF0F";
          m(334) := x"FFB6";
          m(335) := x"0008";
          m(336) := x"0001";
          m(337) := x"FFFB";
          m(338) := x"0043";
          m(339) := x"020F";
          m(340) := x"040C";
          m(341) := x"0234";
          m(342) := x"FE97";
          m(343) := x"FC22";
          m(344) := x"FD68";
          m(345) := x"02FF";
          m(346) := x"06D8";
          m(347) := x"0EED";
          m(348) := x"0B36";
          m(349) := x"12CB";
          m(350) := x"0869";
          m(351) := x"FD7E";
          m(352) := x"FC79";
          m(353) := x"FE60";
          m(354) := x"FF3E";
          m(355) := x"0494";
          m(356) := x"FF64";
          m(357) := x"FE42";
          m(358) := x"07AA";
          m(359) := x"05B1";
          m(360) := x"FEA4";
          m(361) := x"FD72";
          m(362) := x"FFA5";
          m(363) := x"FFF5";
          m(364) := x"0032";
          m(365) := x"0000";
          m(366) := x"FF9A";
          m(367) := x"0378";
          m(368) := x"067C";
          m(369) := x"0539";
          m(370) := x"04C5";
          m(371) := x"09BD";
          m(372) := x"06E7";
          m(373) := x"0B80";
          m(374) := x"108D";
          m(375) := x"0C8C";
          m(376) := x"0F0F";
          m(377) := x"0818";
          m(378) := x"FDCA";
          m(379) := x"0454";
          m(380) := x"0366";
          m(381) := x"0077";
          m(382) := x"0319";
          m(383) := x"07AD";
          m(384) := x"045B";
          m(385) := x"008D";
          m(386) := x"05AD";
          m(387) := x"0284";
          m(388) := x"FE1E";
          m(389) := x"FE55";
          m(390) := x"FF8A";
          m(391) := x"FF60";
          m(392) := x"FFFA";
          m(393) := x"0031";
          m(394) := x"FFB4";
          m(395) := x"03FE";
          m(396) := x"0581";
          m(397) := x"078D";
          m(398) := x"09DF";
          m(399) := x"0775";
          m(400) := x"1402";
          m(401) := x"121C";
          m(402) := x"0A3B";
          m(403) := x"02A5";
          m(404) := x"01E0";
          m(405) := x"0540";
          m(406) := x"FAC6";
          m(407) := x"0252";
          m(408) := x"00CB";
          m(409) := x"0014";
          m(410) := x"FF4A";
          m(411) := x"FF9C";
          m(412) := x"011A";
          m(413) := x"FEC7";
          m(414) := x"017E";
          m(415) := x"FD6B";
          m(416) := x"FC84";
          m(417) := x"FF4B";
          m(418) := x"FF41";
          m(419) := x"0022";
          m(420) := x"FFD2";
          m(421) := x"002C";
          m(422) := x"FF99";
          m(423) := x"0192";
          m(424) := x"0662";
          m(425) := x"093F";
          m(426) := x"0D52";
          m(427) := x"0BC5";
          m(428) := x"0AAD";
          m(429) := x"0574";
          m(430) := x"0084";
          m(431) := x"FBE7";
          m(432) := x"008C";
          m(433) := x"FF3C";
          m(434) := x"0187";
          m(435) := x"FB98";
          m(436) := x"FD9D";
          m(437) := x"FED3";
          m(438) := x"FD5C";
          m(439) := x"01BB";
          m(440) := x"0007";
          m(441) := x"FDD3";
          m(442) := x"010C";
          m(443) := x"0021";
          m(444) := x"FC79";
          m(445) := x"FEDD";
          m(446) := x"FF6B";
          m(447) := x"FFDE";
          m(448) := x"FFD5";
          m(449) := x"FFC9";
          m(450) := x"FF4D";
          m(451) := x"FFAF";
          m(452) := x"0734";
          m(453) := x"09F9";
          m(454) := x"0CFB";
          m(455) := x"0651";
          m(456) := x"0337";
          m(457) := x"02B8";
          m(458) := x"FFA9";
          m(459) := x"FD58";
          m(460) := x"F97E";
          m(461) := x"02DF";
          m(462) := x"02A0";
          m(463) := x"FEAE";
          m(464) := x"FCFB";
          m(465) := x"FB98";
          m(466) := x"FA59";
          m(467) := x"FB73";
          m(468) := x"FE5D";
          m(469) := x"FA29";
          m(470) := x"01E6";
          m(471) := x"01E3";
          m(472) := x"FC89";
          m(473) := x"FE6E";
          m(474) := x"FF81";
          m(475) := x"FFFB";
          m(476) := x"0013";
          m(477) := x"FFEE";
          m(478) := x"FFBE";
          m(479) := x"FF3B";
          m(480) := x"01E0";
          m(481) := x"04B3";
          m(482) := x"043D";
          m(483) := x"00FD";
          m(484) := x"FE7B";
          m(485) := x"02E0";
          m(486) := x"FF6A";
          m(487) := x"FAFE";
          m(488) := x"005C";
          m(489) := x"01A2";
          m(490) := x"01A1";
          m(491) := x"FF69";
          m(492) := x"FED7";
          m(493) := x"FC9A";
          m(494) := x"0177";
          m(495) := x"FBF6";
          m(496) := x"026E";
          m(497) := x"020B";
          m(498) := x"03D4";
          m(499) := x"0438";
          m(500) := x"FE99";
          m(501) := x"FDF5";
          m(502) := x"FFA4";
          m(503) := x"FFF1";
          m(504) := x"FFF1";
          m(505) := x"FFFB";
          m(506) := x"FFE8";
          m(507) := x"FC1B";
          m(508) := x"FA4B";
          m(509) := x"FB36";
          m(510) := x"0169";
          m(511) := x"FB20";
          m(512) := x"FF18";
          m(513) := x"04AE";
          m(514) := x"0086";
          m(515) := x"0145";
          m(516) := x"FA24";
          m(517) := x"FC98";
          m(518) := x"003F";
          m(519) := x"FB03";
          m(520) := x"FD47";
          m(521) := x"FC2C";
          m(522) := x"FF04";
          m(523) := x"FB9A";
          m(524) := x"0449";
          m(525) := x"0342";
          m(526) := x"01F6";
          m(527) := x"0132";
          m(528) := x"FF9F";
          m(529) := x"FEE0";
          m(530) := x"FFA8";
          m(531) := x"FFC3";
          m(532) := x"FFC4";
          m(533) := x"003D";
          m(534) := x"0183";
          m(535) := x"FDF9";
          m(536) := x"FB77";
          m(537) := x"FA88";
          m(538) := x"FCF2";
          m(539) := x"F977";
          m(540) := x"FA29";
          m(541) := x"FBF2";
          m(542) := x"FE4A";
          m(543) := x"FDA5";
          m(544) := x"FED7";
          m(545) := x"FA17";
          m(546) := x"0126";
          m(547) := x"FE10";
          m(548) := x"FE98";
          m(549) := x"FF6C";
          m(550) := x"018F";
          m(551) := x"FED7";
          m(552) := x"02C6";
          m(553) := x"026D";
          m(554) := x"FFA5";
          m(555) := x"FDF7";
          m(556) := x"FE86";
          m(557) := x"FEE1";
          m(558) := x"FF97";
          m(559) := x"FF72";
          m(560) := x"0008";
          m(561) := x"002B";
          m(562) := x"0195";
          m(563) := x"FEF2";
          m(564) := x"FD9D";
          m(565) := x"00C7";
          m(566) := x"FD46";
          m(567) := x"F973";
          m(568) := x"F91E";
          m(569) := x"FE81";
          m(570) := x"FFE1";
          m(571) := x"FD3B";
          m(572) := x"FF35";
          m(573) := x"FDD5";
          m(574) := x"FCE2";
          m(575) := x"FEBF";
          m(576) := x"01E8";
          m(577) := x"FF12";
          m(578) := x"02D2";
          m(579) := x"020E";
          m(580) := x"FC95";
          m(581) := x"FFB8";
          m(582) := x"0001";
          m(583) := x"FD77";
          m(584) := x"FDAA";
          m(585) := x"FECC";
          m(586) := x"FFDD";
          m(587) := x"002A";
          m(588) := x"FFEB";
          m(589) := x"FFDE";
          m(590) := x"FF96";
          m(591) := x"FD4D";
          m(592) := x"00BA";
          m(593) := x"0487";
          m(594) := x"FFF1";
          m(595) := x"FD17";
          m(596) := x"FCAB";
          m(597) := x"FEBA";
          m(598) := x"FC87";
          m(599) := x"0365";
          m(600) := x"FDA3";
          m(601) := x"FB62";
          m(602) := x"FAF2";
          m(603) := x"0286";
          m(604) := x"0398";
          m(605) := x"FDBB";
          m(606) := x"FF0A";
          m(607) := x"F961";
          m(608) := x"FA99";
          m(609) := x"FE64";
          m(610) := x"FE34";
          m(611) := x"FCD0";
          m(612) := x"FE88";
          m(613) := x"FEEE";
          m(614) := x"006D";
          m(615) := x"FFE7";
          m(616) := x"0021";
          m(617) := x"FFDF";
          m(618) := x"FFDC";
          m(619) := x"FFFB";
          m(620) := x"FDC0";
          m(621) := x"FC94";
          m(622) := x"FC02";
          m(623) := x"F960";
          m(624) := x"FE8A";
          m(625) := x"FEA1";
          m(626) := x"FC22";
          m(627) := x"FFE4";
          m(628) := x"FE2C";
          m(629) := x"FFB0";
          m(630) := x"01EF";
          m(631) := x"0050";
          m(632) := x"FEE8";
          m(633) := x"FFBB";
          m(634) := x"045C";
          m(635) := x"00BF";
          m(636) := x"FF50";
          m(637) := x"FA6E";
          m(638) := x"FA5A";
          m(639) := x"FBF1";
          m(640) := x"FCB2";
          m(641) := x"FDBC";
          m(642) := x"FFF3";
          m(643) := x"FFD3";
          m(644) := x"FFF5";
          m(645) := x"0028";
          m(646) := x"007C";
          m(647) := x"00CD";
          m(648) := x"0038";
          m(649) := x"FE9B";
          m(650) := x"FCF3";
          m(651) := x"005B";
          m(652) := x"052C";
          m(653) := x"FF55";
          m(654) := x"FFA8";
          m(655) := x"FCE1";
          m(656) := x"FDAC";
          m(657) := x"002D";
          m(658) := x"0160";
          m(659) := x"FE60";
          m(660) := x"00BE";
          m(661) := x"049A";
          m(662) := x"FDE0";
          m(663) := x"00A8";
          m(664) := x"0380";
          m(665) := x"FCB1";
          m(666) := x"FC4E";
          m(667) := x"FB7F";
          m(668) := x"FDC1";
          m(669) := x"FDC6";
          m(670) := x"FFA9";
          m(671) := x"FFE5";
          m(672) := x"001C";
          m(673) := x"0017";
          m(674) := x"FFE0";
          m(675) := x"FFCF";
          m(676) := x"FDC3";
          m(677) := x"FDC9";
          m(678) := x"FCE0";
          m(679) := x"025A";
          m(680) := x"FDCA";
          m(681) := x"FD10";
          m(682) := x"03FA";
          m(683) := x"036F";
          m(684) := x"047A";
          m(685) := x"001F";
          m(686) := x"FCFB";
          m(687) := x"FB65";
          m(688) := x"0189";
          m(689) := x"FCE8";
          m(690) := x"01CD";
          m(691) := x"0417";
          m(692) := x"0385";
          m(693) := x"000F";
          m(694) := x"0191";
          m(695) := x"FFC9";
          m(696) := x"FE1C";
          m(697) := x"FEEA";
          m(698) := x"0015";
          m(699) := x"FFEC";
          m(700) := x"FFFC";
          m(701) := x"FFDB";
          m(702) := x"000D";
          m(703) := x"FFDE";
          m(704) := x"FDE4";
          m(705) := x"FDFA";
          m(706) := x"FEFC";
          m(707) := x"00BD";
          m(708) := x"FD79";
          m(709) := x"FEB1";
          m(710) := x"04CF";
          m(711) := x"050F";
          m(712) := x"FBF5";
          m(713) := x"001B";
          m(714) := x"FD6B";
          m(715) := x"FB86";
          m(716) := x"FEFC";
          m(717) := x"0140";
          m(718) := x"0420";
          m(719) := x"034A";
          m(720) := x"0340";
          m(721) := x"042A";
          m(722) := x"022E";
          m(723) := x"00D8";
          m(724) := x"0051";
          m(725) := x"FFFA";
          m(726) := x"0004";
          m(727) := x"FFEF";
          m(728) := x"FFFB";
          m(729) := x"002E";
          m(730) := x"FFF5";
          m(731) := x"0012";
          m(732) := x"0078";
          m(733) := x"0232";
          m(734) := x"01D1";
          m(735) := x"FFB8";
          m(736) := x"FF3D";
          m(737) := x"0286";
          m(738) := x"0482";
          m(739) := x"034B";
          m(740) := x"043B";
          m(741) := x"0498";
          m(742) := x"0263";
          m(743) := x"0259";
          m(744) := x"0301";
          m(745) := x"02C5";
          m(746) := x"01E4";
          m(747) := x"010B";
          m(748) := x"02C4";
          m(749) := x"0256";
          m(750) := x"00C0";
          m(751) := x"0047";
          m(752) := x"FFBC";
          m(753) := x"FFF8";
          m(754) := x"0030";
          m(755) := x"0026";
          m(756) := x"FFF6";
          m(757) := x"FFF8";
          m(758) := x"0018";
          m(759) := x"0012";
          m(760) := x"FFFB";
          m(761) := x"FFDE";
          m(762) := x"001B";
          m(763) := x"FFFD";
          m(764) := x"FFD3";
          m(765) := x"FFC2";
          m(766) := x"FF33";
          m(767) := x"0013";
          m(768) := x"0067";
          m(769) := x"0014";
          m(770) := x"FFD8";
          m(771) := x"FFCC";
          m(772) := x"FF82";
          m(773) := x"FFF4";
          m(774) := x"0097";
          m(775) := x"FFFD";
          m(776) := x"00C6";
          m(777) := x"0095";
          m(778) := x"00FF";
          m(779) := x"FFBF";
          m(780) := x"0015";
          m(781) := x"000D";
          m(782) := x"FFDB";
          m(783) := x"002C";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_4.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 4) then
          m(0) := x"FFF2";
          m(1) := x"002D";
          m(2) := x"FFE9";
          m(3) := x"FFD5";
          m(4) := x"FFC4";
          m(5) := x"0013";
          m(6) := x"0001";
          m(7) := x"FFDF";
          m(8) := x"0005";
          m(9) := x"002E";
          m(10) := x"FFD4";
          m(11) := x"FFD4";
          m(12) := x"FFE3";
          m(13) := x"FFD7";
          m(14) := x"0007";
          m(15) := x"000B";
          m(16) := x"FFF8";
          m(17) := x"FFC6";
          m(18) := x"0014";
          m(19) := x"0005";
          m(20) := x"0012";
          m(21) := x"0000";
          m(22) := x"FFFF";
          m(23) := x"001F";
          m(24) := x"FFCE";
          m(25) := x"000A";
          m(26) := x"000D";
          m(27) := x"000B";
          m(28) := x"0028";
          m(29) := x"0004";
          m(30) := x"000E";
          m(31) := x"FFE8";
          m(32) := x"0018";
          m(33) := x"001D";
          m(34) := x"FFF9";
          m(35) := x"0032";
          m(36) := x"003F";
          m(37) := x"0011";
          m(38) := x"FFEA";
          m(39) := x"FFBD";
          m(40) := x"0002";
          m(41) := x"0033";
          m(42) := x"0004";
          m(43) := x"FFF7";
          m(44) := x"004A";
          m(45) := x"FFFC";
          m(46) := x"FFE6";
          m(47) := x"FFCD";
          m(48) := x"0012";
          m(49) := x"0019";
          m(50) := x"FFF4";
          m(51) := x"001E";
          m(52) := x"0008";
          m(53) := x"0050";
          m(54) := x"0039";
          m(55) := x"0037";
          m(56) := x"0003";
          m(57) := x"FFEF";
          m(58) := x"0051";
          m(59) := x"0019";
          m(60) := x"0046";
          m(61) := x"FFFB";
          m(62) := x"FF8E";
          m(63) := x"FFA9";
          m(64) := x"FF89";
          m(65) := x"FF2E";
          m(66) := x"FED8";
          m(67) := x"FE94";
          m(68) := x"FEBA";
          m(69) := x"FEB4";
          m(70) := x"FEE8";
          m(71) := x"FEC0";
          m(72) := x"FF2C";
          m(73) := x"FEC5";
          m(74) := x"FF4A";
          m(75) := x"FEC1";
          m(76) := x"FEE7";
          m(77) := x"FED5";
          m(78) := x"FF6D";
          m(79) := x"FFB6";
          m(80) := x"0069";
          m(81) := x"0049";
          m(82) := x"0006";
          m(83) := x"FFDC";
          m(84) := x"FFF2";
          m(85) := x"001F";
          m(86) := x"FFE2";
          m(87) := x"FFF4";
          m(88) := x"FFD1";
          m(89) := x"FFB1";
          m(90) := x"FEBE";
          m(91) := x"FEB8";
          m(92) := x"FE18";
          m(93) := x"FE5C";
          m(94) := x"0068";
          m(95) := x"0131";
          m(96) := x"000B";
          m(97) := x"FFE0";
          m(98) := x"FF30";
          m(99) := x"FFCF";
          m(100) := x"0041";
          m(101) := x"02D8";
          m(102) := x"0275";
          m(103) := x"FFCB";
          m(104) := x"FD20";
          m(105) := x"FB95";
          m(106) := x"FBBB";
          m(107) := x"FCFD";
          m(108) := x"FE89";
          m(109) := x"0039";
          m(110) := x"FFD6";
          m(111) := x"FFDB";
          m(112) := x"FFE5";
          m(113) := x"0022";
          m(114) := x"FFFD";
          m(115) := x"0014";
          m(116) := x"FFA6";
          m(117) := x"FFE3";
          m(118) := x"FECF";
          m(119) := x"FD7F";
          m(120) := x"FD6B";
          m(121) := x"FD5F";
          m(122) := x"FF1E";
          m(123) := x"0205";
          m(124) := x"FBAB";
          m(125) := x"FA43";
          m(126) := x"FA52";
          m(127) := x"00D1";
          m(128) := x"01F8";
          m(129) := x"01C5";
          m(130) := x"0113";
          m(131) := x"FF21";
          m(132) := x"FF5D";
          m(133) := x"FECA";
          m(134) := x"FCFA";
          m(135) := x"FDB5";
          m(136) := x"FFD4";
          m(137) := x"0100";
          m(138) := x"00B8";
          m(139) := x"FFDC";
          m(140) := x"001C";
          m(141) := x"FFD9";
          m(142) := x"0013";
          m(143) := x"008D";
          m(144) := x"FFD5";
          m(145) := x"007E";
          m(146) := x"FDE5";
          m(147) := x"FD01";
          m(148) := x"FDA0";
          m(149) := x"FD27";
          m(150) := x"FCAC";
          m(151) := x"FFE8";
          m(152) := x"F968";
          m(153) := x"05C4";
          m(154) := x"0550";
          m(155) := x"0BEB";
          m(156) := x"0939";
          m(157) := x"0309";
          m(158) := x"FF59";
          m(159) := x"FBB9";
          m(160) := x"F798";
          m(161) := x"FB79";
          m(162) := x"FDE9";
          m(163) := x"FD73";
          m(164) := x"FE6F";
          m(165) := x"0069";
          m(166) := x"FF7C";
          m(167) := x"FFC4";
          m(168) := x"FFF1";
          m(169) := x"FFF1";
          m(170) := x"0033";
          m(171) := x"FFE7";
          m(172) := x"003E";
          m(173) := x"01FE";
          m(174) := x"FDD8";
          m(175) := x"FC5A";
          m(176) := x"FDE9";
          m(177) := x"F993";
          m(178) := x"020B";
          m(179) := x"008E";
          m(180) := x"FD23";
          m(181) := x"0756";
          m(182) := x"0874";
          m(183) := x"1441";
          m(184) := x"1241";
          m(185) := x"0926";
          m(186) := x"FD89";
          m(187) := x"FA89";
          m(188) := x"FD25";
          m(189) := x"FC46";
          m(190) := x"FF35";
          m(191) := x"FC92";
          m(192) := x"FDB4";
          m(193) := x"0047";
          m(194) := x"FF0C";
          m(195) := x"FF7C";
          m(196) := x"FFE5";
          m(197) := x"0048";
          m(198) := x"0031";
          m(199) := x"00C5";
          m(200) := x"0023";
          m(201) := x"0002";
          m(202) := x"FDFD";
          m(203) := x"FD76";
          m(204) := x"FBD6";
          m(205) := x"FC67";
          m(206) := x"FC1C";
          m(207) := x"F915";
          m(208) := x"F707";
          m(209) := x"FF3B";
          m(210) := x"0A16";
          m(211) := x"1388";
          m(212) := x"0C2F";
          m(213) := x"012D";
          m(214) := x"FE71";
          m(215) := x"F87E";
          m(216) := x"FF77";
          m(217) := x"FEAD";
          m(218) := x"FCF7";
          m(219) := x"FFC9";
          m(220) := x"FFCE";
          m(221) := x"0146";
          m(222) := x"FF40";
          m(223) := x"FFC8";
          m(224) := x"FFE6";
          m(225) := x"000E";
          m(226) := x"000A";
          m(227) := x"0119";
          m(228) := x"0107";
          m(229) := x"00DB";
          m(230) := x"FFA8";
          m(231) := x"FFFA";
          m(232) := x"039B";
          m(233) := x"FE7F";
          m(234) := x"FFA0";
          m(235) := x"FC88";
          m(236) := x"FAB8";
          m(237) := x"FE9A";
          m(238) := x"10BE";
          m(239) := x"15B2";
          m(240) := x"0488";
          m(241) := x"FD5C";
          m(242) := x"FFDD";
          m(243) := x"002E";
          m(244) := x"FFDA";
          m(245) := x"FFFF";
          m(246) := x"FFAD";
          m(247) := x"008D";
          m(248) := x"03D3";
          m(249) := x"023E";
          m(250) := x"00FA";
          m(251) := x"0021";
          m(252) := x"0021";
          m(253) := x"002D";
          m(254) := x"FFFA";
          m(255) := x"0171";
          m(256) := x"013F";
          m(257) := x"0240";
          m(258) := x"0153";
          m(259) := x"08EA";
          m(260) := x"0253";
          m(261) := x"0121";
          m(262) := x"065D";
          m(263) := x"FC48";
          m(264) := x"F7A4";
          m(265) := x"0279";
          m(266) := x"1473";
          m(267) := x"0F91";
          m(268) := x"FF12";
          m(269) := x"0147";
          m(270) := x"01B2";
          m(271) := x"0169";
          m(272) := x"FF4B";
          m(273) := x"FFD2";
          m(274) := x"0271";
          m(275) := x"04D4";
          m(276) := x"02C9";
          m(277) := x"02BA";
          m(278) := x"01D3";
          m(279) := x"0010";
          m(280) := x"FFBB";
          m(281) := x"FFFF";
          m(282) := x"00F6";
          m(283) := x"01FC";
          m(284) := x"02BA";
          m(285) := x"FE57";
          m(286) := x"05A2";
          m(287) := x"02ED";
          m(288) := x"FEE0";
          m(289) := x"FFC2";
          m(290) := x"04EB";
          m(291) := x"FCFF";
          m(292) := x"FE62";
          m(293) := x"0D38";
          m(294) := x"1660";
          m(295) := x"09DA";
          m(296) := x"FF6C";
          m(297) := x"00AE";
          m(298) := x"FF67";
          m(299) := x"00E1";
          m(300) := x"FE60";
          m(301) := x"00C1";
          m(302) := x"0445";
          m(303) := x"0595";
          m(304) := x"00E3";
          m(305) := x"0268";
          m(306) := x"0196";
          m(307) := x"FFBA";
          m(308) := x"0027";
          m(309) := x"FFD7";
          m(310) := x"0153";
          m(311) := x"0146";
          m(312) := x"0390";
          m(313) := x"FF15";
          m(314) := x"0897";
          m(315) := x"06A0";
          m(316) := x"0446";
          m(317) := x"0316";
          m(318) := x"0586";
          m(319) := x"02A9";
          m(320) := x"FE59";
          m(321) := x"0A39";
          m(322) := x"0719";
          m(323) := x"0535";
          m(324) := x"FD1F";
          m(325) := x"0285";
          m(326) := x"FB4F";
          m(327) := x"FDF0";
          m(328) := x"FF0D";
          m(329) := x"03FB";
          m(330) := x"01CF";
          m(331) := x"039C";
          m(332) := x"0256";
          m(333) := x"0056";
          m(334) := x"00F9";
          m(335) := x"FFFB";
          m(336) := x"FFF5";
          m(337) := x"001D";
          m(338) := x"007D";
          m(339) := x"0066";
          m(340) := x"045A";
          m(341) := x"0107";
          m(342) := x"024B";
          m(343) := x"0401";
          m(344) := x"FDAE";
          m(345) := x"04B6";
          m(346) := x"FBF2";
          m(347) := x"F89F";
          m(348) := x"F9C5";
          m(349) := x"FDBE";
          m(350) := x"FEA1";
          m(351) := x"FF73";
          m(352) := x"FD44";
          m(353) := x"0239";
          m(354) := x"FFF1";
          m(355) := x"0402";
          m(356) := x"FE4A";
          m(357) := x"02D9";
          m(358) := x"0291";
          m(359) := x"00A4";
          m(360) := x"0053";
          m(361) := x"0097";
          m(362) := x"0166";
          m(363) := x"006A";
          m(364) := x"FFFA";
          m(365) := x"002D";
          m(366) := x"0054";
          m(367) := x"00C3";
          m(368) := x"02C2";
          m(369) := x"FD53";
          m(370) := x"FE5E";
          m(371) := x"0004";
          m(372) := x"F31E";
          m(373) := x"FE46";
          m(374) := x"F9A2";
          m(375) := x"FF87";
          m(376) := x"0022";
          m(377) := x"FD1D";
          m(378) := x"0256";
          m(379) := x"FE1F";
          m(380) := x"FE43";
          m(381) := x"FEF4";
          m(382) := x"03C4";
          m(383) := x"0483";
          m(384) := x"01F0";
          m(385) := x"009E";
          m(386) := x"007C";
          m(387) := x"FBB2";
          m(388) := x"FE94";
          m(389) := x"0102";
          m(390) := x"00D8";
          m(391) := x"FFBB";
          m(392) := x"004F";
          m(393) := x"0036";
          m(394) := x"0046";
          m(395) := x"00C0";
          m(396) := x"FE89";
          m(397) := x"F6DF";
          m(398) := x"FCC3";
          m(399) := x"FFD0";
          m(400) := x"FF33";
          m(401) := x"FC6F";
          m(402) := x"FE79";
          m(403) := x"FCE4";
          m(404) := x"FFD8";
          m(405) := x"0248";
          m(406) := x"FDAB";
          m(407) := x"FD00";
          m(408) := x"FDDC";
          m(409) := x"FC31";
          m(410) := x"FEFA";
          m(411) := x"FCEA";
          m(412) := x"FD42";
          m(413) := x"FFAB";
          m(414) := x"FBED";
          m(415) := x"FA9D";
          m(416) := x"FDF6";
          m(417) := x"FFA8";
          m(418) := x"0031";
          m(419) := x"FFEB";
          m(420) := x"FFEA";
          m(421) := x"0014";
          m(422) := x"004B";
          m(423) := x"FEBF";
          m(424) := x"FFB3";
          m(425) := x"00A2";
          m(426) := x"FB34";
          m(427) := x"FA39";
          m(428) := x"FF7A";
          m(429) := x"FF08";
          m(430) := x"FC34";
          m(431) := x"FF15";
          m(432) := x"01EC";
          m(433) := x"011A";
          m(434) := x"FB8A";
          m(435) := x"FF8B";
          m(436) := x"FD33";
          m(437) := x"FBEE";
          m(438) := x"FAE8";
          m(439) := x"FB4E";
          m(440) := x"FF75";
          m(441) := x"FF83";
          m(442) := x"FC03";
          m(443) := x"FC85";
          m(444) := x"0065";
          m(445) := x"FE7C";
          m(446) := x"006E";
          m(447) := x"002C";
          m(448) := x"FFEA";
          m(449) := x"0051";
          m(450) := x"002A";
          m(451) := x"FE5D";
          m(452) := x"0131";
          m(453) := x"04B7";
          m(454) := x"FF1A";
          m(455) := x"FB97";
          m(456) := x"FBB7";
          m(457) := x"FAB6";
          m(458) := x"0019";
          m(459) := x"FAF7";
          m(460) := x"FEE2";
          m(461) := x"0266";
          m(462) := x"FC49";
          m(463) := x"FC05";
          m(464) := x"0114";
          m(465) := x"05BF";
          m(466) := x"FF01";
          m(467) := x"FC83";
          m(468) := x"FD20";
          m(469) := x"F7C9";
          m(470) := x"FE16";
          m(471) := x"FC89";
          m(472) := x"FEF3";
          m(473) := x"FE21";
          m(474) := x"FFFF";
          m(475) := x"FFF1";
          m(476) := x"FFE4";
          m(477) := x"FFEA";
          m(478) := x"FFCF";
          m(479) := x"FF4D";
          m(480) := x"00BC";
          m(481) := x"0365";
          m(482) := x"FE56";
          m(483) := x"FF59";
          m(484) := x"006F";
          m(485) := x"FD17";
          m(486) := x"FE9C";
          m(487) := x"FC82";
          m(488) := x"01A5";
          m(489) := x"0323";
          m(490) := x"01BB";
          m(491) := x"02B1";
          m(492) := x"00AB";
          m(493) := x"0196";
          m(494) := x"FFD2";
          m(495) := x"02EF";
          m(496) := x"FCC2";
          m(497) := x"F729";
          m(498) := x"FA3A";
          m(499) := x"FDE5";
          m(500) := x"FF51";
          m(501) := x"FEE9";
          m(502) := x"000D";
          m(503) := x"0077";
          m(504) := x"0031";
          m(505) := x"0001";
          m(506) := x"0041";
          m(507) := x"FE5C";
          m(508) := x"FDE0";
          m(509) := x"0193";
          m(510) := x"0292";
          m(511) := x"FADE";
          m(512) := x"F91C";
          m(513) := x"FD6C";
          m(514) := x"01DE";
          m(515) := x"04A5";
          m(516) := x"FFBD";
          m(517) := x"FF0F";
          m(518) := x"F7D1";
          m(519) := x"0451";
          m(520) := x"0075";
          m(521) := x"FCA6";
          m(522) := x"FFEA";
          m(523) := x"01DD";
          m(524) := x"FFA1";
          m(525) := x"FECB";
          m(526) := x"FDD5";
          m(527) := x"FEA2";
          m(528) := x"FE51";
          m(529) := x"FF07";
          m(530) := x"0040";
          m(531) := x"003F";
          m(532) := x"0043";
          m(533) := x"0003";
          m(534) := x"00DF";
          m(535) := x"FF08";
          m(536) := x"FFB5";
          m(537) := x"01C6";
          m(538) := x"02CE";
          m(539) := x"FBDE";
          m(540) := x"FAFA";
          m(541) := x"FB7F";
          m(542) := x"01B2";
          m(543) := x"FFFC";
          m(544) := x"02CF";
          m(545) := x"FF43";
          m(546) := x"FFDC";
          m(547) := x"FFC3";
          m(548) := x"038D";
          m(549) := x"00EC";
          m(550) := x"0371";
          m(551) := x"0351";
          m(552) := x"FF21";
          m(553) := x"031D";
          m(554) := x"01D5";
          m(555) := x"0193";
          m(556) := x"008A";
          m(557) := x"0075";
          m(558) := x"003F";
          m(559) := x"0017";
          m(560) := x"0012";
          m(561) := x"FFDC";
          m(562) := x"002D";
          m(563) := x"FF73";
          m(564) := x"FF9D";
          m(565) := x"0291";
          m(566) := x"0435";
          m(567) := x"FD82";
          m(568) := x"FDB6";
          m(569) := x"0065";
          m(570) := x"00C2";
          m(571) := x"0478";
          m(572) := x"FFA0";
          m(573) := x"0000";
          m(574) := x"02B3";
          m(575) := x"FFB1";
          m(576) := x"FE5F";
          m(577) := x"011D";
          m(578) := x"0285";
          m(579) := x"0497";
          m(580) := x"0173";
          m(581) := x"0237";
          m(582) := x"0426";
          m(583) := x"0424";
          m(584) := x"023B";
          m(585) := x"0208";
          m(586) := x"000B";
          m(587) := x"FFF9";
          m(588) := x"FFD0";
          m(589) := x"0002";
          m(590) := x"0038";
          m(591) := x"FFC3";
          m(592) := x"FFB4";
          m(593) := x"024B";
          m(594) := x"0225";
          m(595) := x"FE6C";
          m(596) := x"FA82";
          m(597) := x"FF30";
          m(598) := x"01F1";
          m(599) := x"0121";
          m(600) := x"001A";
          m(601) := x"FCDA";
          m(602) := x"FE25";
          m(603) := x"FF34";
          m(604) := x"FF98";
          m(605) := x"FF45";
          m(606) := x"01BF";
          m(607) := x"01FD";
          m(608) := x"FF31";
          m(609) := x"02F2";
          m(610) := x"0377";
          m(611) := x"010E";
          m(612) := x"030F";
          m(613) := x"015C";
          m(614) := x"000A";
          m(615) := x"001B";
          m(616) := x"0016";
          m(617) := x"0000";
          m(618) := x"0027";
          m(619) := x"FFCC";
          m(620) := x"FF97";
          m(621) := x"FFE1";
          m(622) := x"00F0";
          m(623) := x"0104";
          m(624) := x"017B";
          m(625) := x"FE24";
          m(626) := x"FC9B";
          m(627) := x"02B7";
          m(628) := x"0307";
          m(629) := x"006A";
          m(630) := x"01E6";
          m(631) := x"FF98";
          m(632) := x"01F7";
          m(633) := x"04B0";
          m(634) := x"031B";
          m(635) := x"FCE8";
          m(636) := x"FEFB";
          m(637) := x"0242";
          m(638) := x"031B";
          m(639) := x"02A6";
          m(640) := x"019E";
          m(641) := x"0018";
          m(642) := x"FFE5";
          m(643) := x"0014";
          m(644) := x"004A";
          m(645) := x"0012";
          m(646) := x"FFF7";
          m(647) := x"003E";
          m(648) := x"FFB6";
          m(649) := x"FFAB";
          m(650) := x"0130";
          m(651) := x"01A7";
          m(652) := x"03C1";
          m(653) := x"0343";
          m(654) := x"005C";
          m(655) := x"051C";
          m(656) := x"0415";
          m(657) := x"0792";
          m(658) := x"03E6";
          m(659) := x"042E";
          m(660) := x"01FA";
          m(661) := x"03F1";
          m(662) := x"FF07";
          m(663) := x"0186";
          m(664) := x"04A3";
          m(665) := x"02E2";
          m(666) := x"033B";
          m(667) := x"02D8";
          m(668) := x"026E";
          m(669) := x"FFFA";
          m(670) := x"FFD9";
          m(671) := x"001F";
          m(672) := x"FFF0";
          m(673) := x"000C";
          m(674) := x"0046";
          m(675) := x"000A";
          m(676) := x"008B";
          m(677) := x"FFFD";
          m(678) := x"009C";
          m(679) := x"004A";
          m(680) := x"0088";
          m(681) := x"0073";
          m(682) := x"00E4";
          m(683) := x"FD82";
          m(684) := x"FD9D";
          m(685) := x"FCE9";
          m(686) := x"0077";
          m(687) := x"01CE";
          m(688) := x"FE1F";
          m(689) := x"00FA";
          m(690) := x"00D8";
          m(691) := x"039B";
          m(692) := x"06B8";
          m(693) := x"02E3";
          m(694) := x"01A9";
          m(695) := x"0192";
          m(696) := x"0122";
          m(697) := x"0007";
          m(698) := x"FFC2";
          m(699) := x"FFE2";
          m(700) := x"0004";
          m(701) := x"FFE9";
          m(702) := x"FFF5";
          m(703) := x"002A";
          m(704) := x"0059";
          m(705) := x"005F";
          m(706) := x"012C";
          m(707) := x"032F";
          m(708) := x"0173";
          m(709) := x"014E";
          m(710) := x"FFD7";
          m(711) := x"FF71";
          m(712) := x"FF90";
          m(713) := x"00CF";
          m(714) := x"02C4";
          m(715) := x"FDFC";
          m(716) := x"FDA0";
          m(717) := x"02F7";
          m(718) := x"01FC";
          m(719) := x"0786";
          m(720) := x"0576";
          m(721) := x"0103";
          m(722) := x"0099";
          m(723) := x"FF0D";
          m(724) := x"FFE1";
          m(725) := x"FFFF";
          m(726) := x"0033";
          m(727) := x"0013";
          m(728) := x"001B";
          m(729) := x"0021";
          m(730) := x"0015";
          m(731) := x"FFBF";
          m(732) := x"002E";
          m(733) := x"00C2";
          m(734) := x"0095";
          m(735) := x"00A8";
          m(736) := x"FFD5";
          m(737) := x"0052";
          m(738) := x"02C0";
          m(739) := x"03E5";
          m(740) := x"0375";
          m(741) := x"042F";
          m(742) := x"0689";
          m(743) := x"04B8";
          m(744) := x"0560";
          m(745) := x"0104";
          m(746) := x"030C";
          m(747) := x"02CD";
          m(748) := x"0198";
          m(749) := x"001A";
          m(750) := x"0006";
          m(751) := x"FFEF";
          m(752) := x"0002";
          m(753) := x"0015";
          m(754) := x"FFCA";
          m(755) := x"FFF0";
          m(756) := x"FFEC";
          m(757) := x"0010";
          m(758) := x"000C";
          m(759) := x"FFD4";
          m(760) := x"001E";
          m(761) := x"000D";
          m(762) := x"0047";
          m(763) := x"00F5";
          m(764) := x"00E2";
          m(765) := x"003E";
          m(766) := x"0013";
          m(767) := x"007F";
          m(768) := x"0060";
          m(769) := x"003C";
          m(770) := x"006C";
          m(771) := x"0051";
          m(772) := x"003B";
          m(773) := x"FFDC";
          m(774) := x"0015";
          m(775) := x"000F";
          m(776) := x"0015";
          m(777) := x"004F";
          m(778) := x"0000";
          m(779) := x"000C";
          m(780) := x"FFCA";
          m(781) := x"0020";
          m(782) := x"0006";
          m(783) := x"FFE6";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_5.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 5) then
          m(0) := x"FFFC";
          m(1) := x"0001";
          m(2) := x"FFD5";
          m(3) := x"0000";
          m(4) := x"FFF7";
          m(5) := x"FFE5";
          m(6) := x"0037";
          m(7) := x"0004";
          m(8) := x"FFE5";
          m(9) := x"001B";
          m(10) := x"0014";
          m(11) := x"FFDD";
          m(12) := x"0024";
          m(13) := x"FFF9";
          m(14) := x"000C";
          m(15) := x"FFFC";
          m(16) := x"000D";
          m(17) := x"0021";
          m(18) := x"002F";
          m(19) := x"0032";
          m(20) := x"001A";
          m(21) := x"FFD0";
          m(22) := x"0015";
          m(23) := x"FFDF";
          m(24) := x"FFEC";
          m(25) := x"FFF2";
          m(26) := x"FFE1";
          m(27) := x"000B";
          m(28) := x"000A";
          m(29) := x"001B";
          m(30) := x"0006";
          m(31) := x"0021";
          m(32) := x"0024";
          m(33) := x"000E";
          m(34) := x"FFE7";
          m(35) := x"0009";
          m(36) := x"000B";
          m(37) := x"FFDB";
          m(38) := x"FFEC";
          m(39) := x"000F";
          m(40) := x"FFEE";
          m(41) := x"005B";
          m(42) := x"FF71";
          m(43) := x"FE8C";
          m(44) := x"FE2D";
          m(45) := x"FFC0";
          m(46) := x"FFBC";
          m(47) := x"FFFC";
          m(48) := x"000A";
          m(49) := x"0049";
          m(50) := x"0038";
          m(51) := x"001C";
          m(52) := x"FFD6";
          m(53) := x"0004";
          m(54) := x"003D";
          m(55) := x"FFE1";
          m(56) := x"FFF1";
          m(57) := x"0032";
          m(58) := x"FFF2";
          m(59) := x"0008";
          m(60) := x"0045";
          m(61) := x"001E";
          m(62) := x"005B";
          m(63) := x"0083";
          m(64) := x"0090";
          m(65) := x"0101";
          m(66) := x"01BA";
          m(67) := x"017F";
          m(68) := x"0133";
          m(69) := x"FF4F";
          m(70) := x"FDFC";
          m(71) := x"FC70";
          m(72) := x"FC26";
          m(73) := x"FF54";
          m(74) := x"006C";
          m(75) := x"01FA";
          m(76) := x"01FF";
          m(77) := x"0130";
          m(78) := x"00B9";
          m(79) := x"0080";
          m(80) := x"0025";
          m(81) := x"FFF1";
          m(82) := x"FFF7";
          m(83) := x"0025";
          m(84) := x"0000";
          m(85) := x"0015";
          m(86) := x"FFFE";
          m(87) := x"0008";
          m(88) := x"0024";
          m(89) := x"002A";
          m(90) := x"00DC";
          m(91) := x"0105";
          m(92) := x"01EA";
          m(93) := x"03B4";
          m(94) := x"032C";
          m(95) := x"0363";
          m(96) := x"0056";
          m(97) := x"F886";
          m(98) := x"F583";
          m(99) := x"F65B";
          m(100) := x"F673";
          m(101) := x"FDF8";
          m(102) := x"022A";
          m(103) := x"042B";
          m(104) := x"0318";
          m(105) := x"010B";
          m(106) := x"01B6";
          m(107) := x"00CF";
          m(108) := x"00CD";
          m(109) := x"FF9F";
          m(110) := x"0004";
          m(111) := x"FFF0";
          m(112) := x"FFC7";
          m(113) := x"0033";
          m(114) := x"FFCF";
          m(115) := x"FFB3";
          m(116) := x"0000";
          m(117) := x"0116";
          m(118) := x"01F6";
          m(119) := x"02BA";
          m(120) := x"04B0";
          m(121) := x"04EA";
          m(122) := x"039B";
          m(123) := x"00AE";
          m(124) := x"FD6D";
          m(125) := x"F4E3";
          m(126) := x"F182";
          m(127) := x"F1F3";
          m(128) := x"FA45";
          m(129) := x"FEC7";
          m(130) := x"007A";
          m(131) := x"0469";
          m(132) := x"033A";
          m(133) := x"0021";
          m(134) := x"02BF";
          m(135) := x"01EA";
          m(136) := x"FE69";
          m(137) := x"FD84";
          m(138) := x"FE75";
          m(139) := x"0065";
          m(140) := x"FFE5";
          m(141) := x"003F";
          m(142) := x"FFF7";
          m(143) := x"0011";
          m(144) := x"00C0";
          m(145) := x"0312";
          m(146) := x"04D4";
          m(147) := x"05B8";
          m(148) := x"0795";
          m(149) := x"0780";
          m(150) := x"0607";
          m(151) := x"FFD2";
          m(152) := x"F82A";
          m(153) := x"ED56";
          m(154) := x"EFD4";
          m(155) := x"F1DB";
          m(156) := x"FF1C";
          m(157) := x"050F";
          m(158) := x"0557";
          m(159) := x"024B";
          m(160) := x"0529";
          m(161) := x"02C4";
          m(162) := x"FF62";
          m(163) := x"0291";
          m(164) := x"0447";
          m(165) := x"00D3";
          m(166) := x"00BE";
          m(167) := x"005F";
          m(168) := x"FFDD";
          m(169) := x"0009";
          m(170) := x"FFDC";
          m(171) := x"FFE4";
          m(172) := x"FF1E";
          m(173) := x"0054";
          m(174) := x"0334";
          m(175) := x"0623";
          m(176) := x"0752";
          m(177) := x"02D8";
          m(178) := x"0425";
          m(179) := x"FCB3";
          m(180) := x"F598";
          m(181) := x"E98C";
          m(182) := x"F170";
          m(183) := x"0193";
          m(184) := x"015C";
          m(185) := x"0285";
          m(186) := x"FEEA";
          m(187) := x"FD88";
          m(188) := x"04CB";
          m(189) := x"011F";
          m(190) := x"FEB8";
          m(191) := x"FFE4";
          m(192) := x"0374";
          m(193) := x"0225";
          m(194) := x"0067";
          m(195) := x"00A5";
          m(196) := x"FFE1";
          m(197) := x"FFDC";
          m(198) := x"FFF9";
          m(199) := x"FDDC";
          m(200) := x"FF05";
          m(201) := x"0482";
          m(202) := x"03C8";
          m(203) := x"03B9";
          m(204) := x"04A0";
          m(205) := x"011E";
          m(206) := x"02E0";
          m(207) := x"FD54";
          m(208) := x"F255";
          m(209) := x"E774";
          m(210) := x"FBA0";
          m(211) := x"0536";
          m(212) := x"07C1";
          m(213) := x"06EB";
          m(214) := x"FFEB";
          m(215) := x"015B";
          m(216) := x"03C1";
          m(217) := x"FE4E";
          m(218) := x"FDAE";
          m(219) := x"FA04";
          m(220) := x"FCA2";
          m(221) := x"00A1";
          m(222) := x"0066";
          m(223) := x"0051";
          m(224) := x"FFD8";
          m(225) := x"FF9E";
          m(226) := x"FFB6";
          m(227) := x"FF2E";
          m(228) := x"0173";
          m(229) := x"0628";
          m(230) := x"0327";
          m(231) := x"009B";
          m(232) := x"FE90";
          m(233) := x"018C";
          m(234) := x"00DE";
          m(235) := x"FA64";
          m(236) := x"E848";
          m(237) := x"F163";
          m(238) := x"01F4";
          m(239) := x"02A8";
          m(240) := x"05F9";
          m(241) := x"080F";
          m(242) := x"FECA";
          m(243) := x"FF41";
          m(244) := x"FB91";
          m(245) := x"FC65";
          m(246) := x"FBCF";
          m(247) := x"F89A";
          m(248) := x"F9FA";
          m(249) := x"FE0A";
          m(250) := x"FEA7";
          m(251) := x"FFF4";
          m(252) := x"0009";
          m(253) := x"FF5C";
          m(254) := x"FFA3";
          m(255) := x"FF9C";
          m(256) := x"01E4";
          m(257) := x"0233";
          m(258) := x"FB56";
          m(259) := x"FDEB";
          m(260) := x"FF07";
          m(261) := x"00F6";
          m(262) := x"0149";
          m(263) := x"FCE3";
          m(264) := x"EEA1";
          m(265) := x"F2F3";
          m(266) := x"FB9E";
          m(267) := x"0999";
          m(268) := x"07BF";
          m(269) := x"00DB";
          m(270) := x"0089";
          m(271) := x"010C";
          m(272) := x"0289";
          m(273) := x"FEEF";
          m(274) := x"F992";
          m(275) := x"F9A9";
          m(276) := x"FC00";
          m(277) := x"FC92";
          m(278) := x"FE73";
          m(279) := x"FFDB";
          m(280) := x"FFE1";
          m(281) := x"FF63";
          m(282) := x"FF6B";
          m(283) := x"FEBB";
          m(284) := x"0050";
          m(285) := x"FEB3";
          m(286) := x"F6E8";
          m(287) := x"FF9E";
          m(288) := x"0183";
          m(289) := x"01F9";
          m(290) := x"FF1A";
          m(291) := x"FC33";
          m(292) := x"F962";
          m(293) := x"F4DC";
          m(294) := x"FEE5";
          m(295) := x"04DB";
          m(296) := x"0159";
          m(297) := x"05B6";
          m(298) := x"FD94";
          m(299) := x"FC8F";
          m(300) := x"FC38";
          m(301) := x"F986";
          m(302) := x"F8E7";
          m(303) := x"FBE8";
          m(304) := x"FECB";
          m(305) := x"FEB8";
          m(306) := x"FF12";
          m(307) := x"FFF5";
          m(308) := x"FFF0";
          m(309) := x"FF91";
          m(310) := x"FFA0";
          m(311) := x"FEC5";
          m(312) := x"FD32";
          m(313) := x"FF05";
          m(314) := x"FE07";
          m(315) := x"FC85";
          m(316) := x"000E";
          m(317) := x"027B";
          m(318) := x"0039";
          m(319) := x"F8B1";
          m(320) := x"F69D";
          m(321) := x"FCB0";
          m(322) := x"FD86";
          m(323) := x"0170";
          m(324) := x"03C5";
          m(325) := x"0137";
          m(326) := x"F9EF";
          m(327) := x"F6E2";
          m(328) := x"FB82";
          m(329) := x"FC80";
          m(330) := x"FC97";
          m(331) := x"FE1E";
          m(332) := x"FF07";
          m(333) := x"FFB7";
          m(334) := x"FFB3";
          m(335) := x"FFE8";
          m(336) := x"0036";
          m(337) := x"FFD8";
          m(338) := x"FFAC";
          m(339) := x"FFB2";
          m(340) := x"FE8A";
          m(341) := x"016E";
          m(342) := x"0249";
          m(343) := x"012B";
          m(344) := x"FC5F";
          m(345) := x"0241";
          m(346) := x"05F8";
          m(347) := x"FCEB";
          m(348) := x"FC6A";
          m(349) := x"0374";
          m(350) := x"FD4F";
          m(351) := x"FD73";
          m(352) := x"FDFD";
          m(353) := x"FDCD";
          m(354) := x"FF38";
          m(355) := x"FE55";
          m(356) := x"01FB";
          m(357) := x"0547";
          m(358) := x"01CD";
          m(359) := x"0260";
          m(360) := x"007D";
          m(361) := x"FE17";
          m(362) := x"FF06";
          m(363) := x"0022";
          m(364) := x"0033";
          m(365) := x"FFDF";
          m(366) := x"FFA7";
          m(367) := x"FF8C";
          m(368) := x"FFC7";
          m(369) := x"0068";
          m(370) := x"02BC";
          m(371) := x"FF7E";
          m(372) := x"FE02";
          m(373) := x"FFB8";
          m(374) := x"01A3";
          m(375) := x"FF29";
          m(376) := x"007E";
          m(377) := x"0312";
          m(378) := x"FD39";
          m(379) := x"FB91";
          m(380) := x"023F";
          m(381) := x"04CC";
          m(382) := x"01BC";
          m(383) := x"0235";
          m(384) := x"0253";
          m(385) := x"00A7";
          m(386) := x"03A4";
          m(387) := x"0416";
          m(388) := x"FE2A";
          m(389) := x"FE67";
          m(390) := x"FF52";
          m(391) := x"FFE0";
          m(392) := x"FFD1";
          m(393) := x"FFA8";
          m(394) := x"FF91";
          m(395) := x"FFBE";
          m(396) := x"02D0";
          m(397) := x"0453";
          m(398) := x"FDEE";
          m(399) := x"02AC";
          m(400) := x"01E3";
          m(401) := x"0297";
          m(402) := x"02D5";
          m(403) := x"0125";
          m(404) := x"020A";
          m(405) := x"FEF7";
          m(406) := x"0182";
          m(407) := x"FEF6";
          m(408) := x"0217";
          m(409) := x"0524";
          m(410) := x"FBA0";
          m(411) := x"FFC6";
          m(412) := x"FCB1";
          m(413) := x"FC2A";
          m(414) := x"0108";
          m(415) := x"FDD4";
          m(416) := x"FF50";
          m(417) := x"FF6C";
          m(418) := x"FEEB";
          m(419) := x"0012";
          m(420) := x"0011";
          m(421) := x"0000";
          m(422) := x"0097";
          m(423) := x"001F";
          m(424) := x"0367";
          m(425) := x"FE84";
          m(426) := x"0145";
          m(427) := x"057E";
          m(428) := x"0063";
          m(429) := x"0330";
          m(430) := x"02C9";
          m(431) := x"FCFA";
          m(432) := x"0428";
          m(433) := x"0306";
          m(434) := x"FFBA";
          m(435) := x"FDC1";
          m(436) := x"00D0";
          m(437) := x"FF63";
          m(438) := x"FCF4";
          m(439) := x"FF9A";
          m(440) := x"FA7D";
          m(441) := x"FEF8";
          m(442) := x"037F";
          m(443) := x"FDAF";
          m(444) := x"FD11";
          m(445) := x"FE8C";
          m(446) := x"FE73";
          m(447) := x"FFB9";
          m(448) := x"0003";
          m(449) := x"FFDB";
          m(450) := x"0072";
          m(451) := x"FEB2";
          m(452) := x"FDEB";
          m(453) := x"FDFE";
          m(454) := x"0088";
          m(455) := x"0324";
          m(456) := x"FF43";
          m(457) := x"0083";
          m(458) := x"FE41";
          m(459) := x"FAB9";
          m(460) := x"038D";
          m(461) := x"00A6";
          m(462) := x"006E";
          m(463) := x"02BC";
          m(464) := x"FF9E";
          m(465) := x"FCE7";
          m(466) := x"0314";
          m(467) := x"0806";
          m(468) := x"03E8";
          m(469) := x"05BD";
          m(470) := x"FE93";
          m(471) := x"0080";
          m(472) := x"FF9E";
          m(473) := x"0024";
          m(474) := x"FF92";
          m(475) := x"000C";
          m(476) := x"FFE6";
          m(477) := x"001B";
          m(478) := x"0148";
          m(479) := x"001C";
          m(480) := x"FFC7";
          m(481) := x"FE3B";
          m(482) := x"FCB9";
          m(483) := x"0057";
          m(484) := x"FE89";
          m(485) := x"015F";
          m(486) := x"0142";
          m(487) := x"FD19";
          m(488) := x"FD9E";
          m(489) := x"FD18";
          m(490) := x"FD76";
          m(491) := x"00F8";
          m(492) := x"FEB3";
          m(493) := x"00A3";
          m(494) := x"032E";
          m(495) := x"FC47";
          m(496) := x"006B";
          m(497) := x"00DE";
          m(498) := x"FB79";
          m(499) := x"FD1C";
          m(500) := x"FDBA";
          m(501) := x"FF57";
          m(502) := x"FF5F";
          m(503) := x"FF8F";
          m(504) := x"003C";
          m(505) := x"FFE1";
          m(506) := x"00C2";
          m(507) := x"02DB";
          m(508) := x"0104";
          m(509) := x"FF2F";
          m(510) := x"FDE9";
          m(511) := x"FDEE";
          m(512) := x"FE16";
          m(513) := x"02A4";
          m(514) := x"0137";
          m(515) := x"FE7B";
          m(516) := x"02A1";
          m(517) := x"01BD";
          m(518) := x"0020";
          m(519) := x"0013";
          m(520) := x"008A";
          m(521) := x"FE06";
          m(522) := x"0225";
          m(523) := x"FC51";
          m(524) := x"0358";
          m(525) := x"FFC4";
          m(526) := x"FD65";
          m(527) := x"FE76";
          m(528) := x"FEA1";
          m(529) := x"FF03";
          m(530) := x"FF31";
          m(531) := x"FFDA";
          m(532) := x"FFD4";
          m(533) := x"0014";
          m(534) := x"0087";
          m(535) := x"0137";
          m(536) := x"FEBF";
          m(537) := x"FC8A";
          m(538) := x"FD1E";
          m(539) := x"FDFA";
          m(540) := x"FA23";
          m(541) := x"FE83";
          m(542) := x"FD4B";
          m(543) := x"018E";
          m(544) := x"FBA2";
          m(545) := x"FD7D";
          m(546) := x"00DE";
          m(547) := x"0270";
          m(548) := x"028E";
          m(549) := x"FF33";
          m(550) := x"FFF8";
          m(551) := x"FDEF";
          m(552) := x"FFE6";
          m(553) := x"FFAC";
          m(554) := x"FD16";
          m(555) := x"FF9B";
          m(556) := x"0042";
          m(557) := x"0057";
          m(558) := x"FFBA";
          m(559) := x"0045";
          m(560) := x"FFEB";
          m(561) := x"FFCB";
          m(562) := x"0035";
          m(563) := x"006B";
          m(564) := x"FD39";
          m(565) := x"F8A8";
          m(566) := x"FADA";
          m(567) := x"FF75";
          m(568) := x"FE62";
          m(569) := x"FE75";
          m(570) := x"05C6";
          m(571) := x"00C1";
          m(572) := x"004E";
          m(573) := x"FC4A";
          m(574) := x"FDEB";
          m(575) := x"00BC";
          m(576) := x"036A";
          m(577) := x"FEFE";
          m(578) := x"0490";
          m(579) := x"FFC9";
          m(580) := x"FB16";
          m(581) := x"FF77";
          m(582) := x"FDD8";
          m(583) := x"FF34";
          m(584) := x"FFD5";
          m(585) := x"0026";
          m(586) := x"FFE1";
          m(587) := x"FFED";
          m(588) := x"FFD8";
          m(589) := x"FFF4";
          m(590) := x"FF7A";
          m(591) := x"0037";
          m(592) := x"FEBE";
          m(593) := x"FBF7";
          m(594) := x"FC11";
          m(595) := x"FF79";
          m(596) := x"0353";
          m(597) := x"01F1";
          m(598) := x"0435";
          m(599) := x"0292";
          m(600) := x"FBF5";
          m(601) := x"003F";
          m(602) := x"01C5";
          m(603) := x"FFC2";
          m(604) := x"0255";
          m(605) := x"FFEE";
          m(606) := x"020F";
          m(607) := x"00CD";
          m(608) := x"FD2D";
          m(609) := x"0043";
          m(610) := x"0112";
          m(611) := x"00DD";
          m(612) := x"003D";
          m(613) := x"0014";
          m(614) := x"FFAC";
          m(615) := x"001E";
          m(616) := x"FFDD";
          m(617) := x"FFE8";
          m(618) := x"0003";
          m(619) := x"0014";
          m(620) := x"0054";
          m(621) := x"00D9";
          m(622) := x"002A";
          m(623) := x"FE80";
          m(624) := x"00A3";
          m(625) := x"FF0D";
          m(626) := x"FEA4";
          m(627) := x"015A";
          m(628) := x"FD50";
          m(629) := x"03AC";
          m(630) := x"FEAD";
          m(631) := x"0231";
          m(632) := x"0016";
          m(633) := x"FD8A";
          m(634) := x"FD5D";
          m(635) := x"FF16";
          m(636) := x"0142";
          m(637) := x"0325";
          m(638) := x"017A";
          m(639) := x"FE8C";
          m(640) := x"FFC5";
          m(641) := x"0045";
          m(642) := x"FFD8";
          m(643) := x"0001";
          m(644) := x"0006";
          m(645) := x"FFE9";
          m(646) := x"0018";
          m(647) := x"FFE4";
          m(648) := x"0034";
          m(649) := x"00FB";
          m(650) := x"01AA";
          m(651) := x"FFBA";
          m(652) := x"01F7";
          m(653) := x"FF2F";
          m(654) := x"FCC3";
          m(655) := x"FE81";
          m(656) := x"FF3E";
          m(657) := x"00BC";
          m(658) := x"FE76";
          m(659) := x"01A4";
          m(660) := x"F989";
          m(661) := x"F9EE";
          m(662) := x"031E";
          m(663) := x"01E9";
          m(664) := x"03A3";
          m(665) := x"0501";
          m(666) := x"0102";
          m(667) := x"FEF2";
          m(668) := x"FE5A";
          m(669) := x"FFF0";
          m(670) := x"0000";
          m(671) := x"FFF3";
          m(672) := x"000B";
          m(673) := x"FFED";
          m(674) := x"0012";
          m(675) := x"FFD4";
          m(676) := x"FF4E";
          m(677) := x"FF9A";
          m(678) := x"FF62";
          m(679) := x"FEC5";
          m(680) := x"FE0C";
          m(681) := x"FE0E";
          m(682) := x"FCAF";
          m(683) := x"FDA6";
          m(684) := x"FCD5";
          m(685) := x"FFA6";
          m(686) := x"0287";
          m(687) := x"034D";
          m(688) := x"FEDE";
          m(689) := x"0443";
          m(690) := x"0806";
          m(691) := x"0109";
          m(692) := x"FC97";
          m(693) := x"0181";
          m(694) := x"FF24";
          m(695) := x"FD45";
          m(696) := x"FF80";
          m(697) := x"FFF4";
          m(698) := x"0025";
          m(699) := x"FFC6";
          m(700) := x"0008";
          m(701) := x"FFF6";
          m(702) := x"FFCD";
          m(703) := x"0001";
          m(704) := x"FFA2";
          m(705) := x"FF94";
          m(706) := x"FE49";
          m(707) := x"FD0E";
          m(708) := x"FE85";
          m(709) := x"FE70";
          m(710) := x"FD33";
          m(711) := x"FD4B";
          m(712) := x"FB4E";
          m(713) := x"FE86";
          m(714) := x"F8DA";
          m(715) := x"00AC";
          m(716) := x"FA1B";
          m(717) := x"FEDA";
          m(718) := x"0192";
          m(719) := x"F4E9";
          m(720) := x"F8FA";
          m(721) := x"FD7B";
          m(722) := x"FCCA";
          m(723) := x"FE22";
          m(724) := x"FFD2";
          m(725) := x"FFCA";
          m(726) := x"002E";
          m(727) := x"FFED";
          m(728) := x"000C";
          m(729) := x"FFF0";
          m(730) := x"FFE0";
          m(731) := x"001F";
          m(732) := x"FFDB";
          m(733) := x"0057";
          m(734) := x"FF67";
          m(735) := x"FEF6";
          m(736) := x"FE4D";
          m(737) := x"FEBA";
          m(738) := x"FE14";
          m(739) := x"FF71";
          m(740) := x"FC01";
          m(741) := x"F9F8";
          m(742) := x"FA55";
          m(743) := x"004C";
          m(744) := x"FB9C";
          m(745) := x"FC3C";
          m(746) := x"F932";
          m(747) := x"FCE9";
          m(748) := x"FD09";
          m(749) := x"FC90";
          m(750) := x"FE9D";
          m(751) := x"000D";
          m(752) := x"000C";
          m(753) := x"0009";
          m(754) := x"FFF1";
          m(755) := x"001B";
          m(756) := x"000B";
          m(757) := x"0011";
          m(758) := x"000D";
          m(759) := x"FFF9";
          m(760) := x"FFFE";
          m(761) := x"0018";
          m(762) := x"FFE6";
          m(763) := x"FFDB";
          m(764) := x"FFDB";
          m(765) := x"FFEA";
          m(766) := x"FF7E";
          m(767) := x"FF52";
          m(768) := x"FF38";
          m(769) := x"FFA4";
          m(770) := x"FEC7";
          m(771) := x"FF64";
          m(772) := x"FFEB";
          m(773) := x"FEC6";
          m(774) := x"FD62";
          m(775) := x"000C";
          m(776) := x"FFE9";
          m(777) := x"FFDA";
          m(778) := x"FF45";
          m(779) := x"FFE5";
          m(780) := x"000F";
          m(781) := x"FFE3";
          m(782) := x"FFEE";
          m(783) := x"FFEB";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_6.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 6) then
          m(0) := x"FFE8";
          m(1) := x"0005";
          m(2) := x"FFEA";
          m(3) := x"FFF8";
          m(4) := x"FFCE";
          m(5) := x"000E";
          m(6) := x"FFE8";
          m(7) := x"FFD3";
          m(8) := x"001B";
          m(9) := x"0021";
          m(10) := x"0002";
          m(11) := x"FFE9";
          m(12) := x"FFF3";
          m(13) := x"FFFB";
          m(14) := x"002B";
          m(15) := x"0034";
          m(16) := x"0038";
          m(17) := x"FFE1";
          m(18) := x"002C";
          m(19) := x"FFF7";
          m(20) := x"FFFC";
          m(21) := x"000F";
          m(22) := x"FFFE";
          m(23) := x"FFEE";
          m(24) := x"FFD8";
          m(25) := x"0007";
          m(26) := x"FFC5";
          m(27) := x"FFF7";
          m(28) := x"FFFF";
          m(29) := x"003D";
          m(30) := x"0014";
          m(31) := x"FFF0";
          m(32) := x"0036";
          m(33) := x"0000";
          m(34) := x"FFDD";
          m(35) := x"FF60";
          m(36) := x"FF81";
          m(37) := x"FFC7";
          m(38) := x"FF73";
          m(39) := x"FF67";
          m(40) := x"FEB3";
          m(41) := x"FF0C";
          m(42) := x"FF19";
          m(43) := x"FE8B";
          m(44) := x"FE9C";
          m(45) := x"FF01";
          m(46) := x"FF86";
          m(47) := x"FF43";
          m(48) := x"FF6A";
          m(49) := x"FFCA";
          m(50) := x"FFAE";
          m(51) := x"FF9C";
          m(52) := x"FFFF";
          m(53) := x"0005";
          m(54) := x"FFF0";
          m(55) := x"FFCF";
          m(56) := x"0013";
          m(57) := x"0021";
          m(58) := x"002F";
          m(59) := x"001F";
          m(60) := x"FFC5";
          m(61) := x"FFF5";
          m(62) := x"FF4C";
          m(63) := x"FEDC";
          m(64) := x"FEB7";
          m(65) := x"FEA8";
          m(66) := x"FE1B";
          m(67) := x"FD19";
          m(68) := x"FCFF";
          m(69) := x"FFAF";
          m(70) := x"FC79";
          m(71) := x"FDC6";
          m(72) := x"FD64";
          m(73) := x"FBA1";
          m(74) := x"FD21";
          m(75) := x"FE09";
          m(76) := x"FEB6";
          m(77) := x"FE1C";
          m(78) := x"FF4E";
          m(79) := x"FF86";
          m(80) := x"FFE1";
          m(81) := x"000E";
          m(82) := x"0059";
          m(83) := x"FFDF";
          m(84) := x"0044";
          m(85) := x"FFFA";
          m(86) := x"000B";
          m(87) := x"0008";
          m(88) := x"FFC4";
          m(89) := x"FFAA";
          m(90) := x"FF19";
          m(91) := x"FE15";
          m(92) := x"FC4C";
          m(93) := x"FB3F";
          m(94) := x"FD8D";
          m(95) := x"FD1F";
          m(96) := x"FE84";
          m(97) := x"FE52";
          m(98) := x"FF7A";
          m(99) := x"0082";
          m(100) := x"FFD2";
          m(101) := x"01D4";
          m(102) := x"0381";
          m(103) := x"0209";
          m(104) := x"FF64";
          m(105) := x"FD92";
          m(106) := x"FFD9";
          m(107) := x"0053";
          m(108) := x"0058";
          m(109) := x"00EF";
          m(110) := x"0046";
          m(111) := x"FFDB";
          m(112) := x"FFE2";
          m(113) := x"FFCB";
          m(114) := x"FFE2";
          m(115) := x"FFE7";
          m(116) := x"FF80";
          m(117) := x"FF56";
          m(118) := x"FEF0";
          m(119) := x"FD29";
          m(120) := x"FA4C";
          m(121) := x"F754";
          m(122) := x"FB87";
          m(123) := x"FD92";
          m(124) := x"FF14";
          m(125) := x"FDE1";
          m(126) := x"FD85";
          m(127) := x"FE56";
          m(128) := x"FE33";
          m(129) := x"FD16";
          m(130) := x"00EA";
          m(131) := x"FB9B";
          m(132) := x"FEDA";
          m(133) := x"0069";
          m(134) := x"021E";
          m(135) := x"0269";
          m(136) := x"00AD";
          m(137) := x"FF84";
          m(138) := x"FF35";
          m(139) := x"FF7C";
          m(140) := x"FFE8";
          m(141) := x"FFCA";
          m(142) := x"000C";
          m(143) := x"FFD9";
          m(144) := x"FF7F";
          m(145) := x"00D5";
          m(146) := x"FFDC";
          m(147) := x"FEB9";
          m(148) := x"FCE9";
          m(149) := x"FC0F";
          m(150) := x"FA8E";
          m(151) := x"FAC5";
          m(152) := x"FB0A";
          m(153) := x"FB1A";
          m(154) := x"F90A";
          m(155) := x"FB20";
          m(156) := x"FC8D";
          m(157) := x"FD27";
          m(158) := x"021D";
          m(159) := x"FB63";
          m(160) := x"007D";
          m(161) := x"02C1";
          m(162) := x"0291";
          m(163) := x"0156";
          m(164) := x"FF0B";
          m(165) := x"FC09";
          m(166) := x"FE45";
          m(167) := x"FF5D";
          m(168) := x"0025";
          m(169) := x"000E";
          m(170) := x"002A";
          m(171) := x"FFDF";
          m(172) := x"FFD0";
          m(173) := x"0329";
          m(174) := x"043C";
          m(175) := x"FFCA";
          m(176) := x"FE61";
          m(177) := x"010C";
          m(178) := x"FEF0";
          m(179) := x"F7B5";
          m(180) := x"FC05";
          m(181) := x"FF0C";
          m(182) := x"FEE6";
          m(183) := x"FCD3";
          m(184) := x"FDEA";
          m(185) := x"FD13";
          m(186) := x"01E4";
          m(187) := x"0065";
          m(188) := x"025C";
          m(189) := x"01C7";
          m(190) := x"0189";
          m(191) := x"FFB9";
          m(192) := x"02F8";
          m(193) := x"FFD2";
          m(194) := x"00FA";
          m(195) := x"0007";
          m(196) := x"0000";
          m(197) := x"0053";
          m(198) := x"0083";
          m(199) := x"0211";
          m(200) := x"0251";
          m(201) := x"0194";
          m(202) := x"0364";
          m(203) := x"00CB";
          m(204) := x"FE84";
          m(205) := x"FF02";
          m(206) := x"00BE";
          m(207) := x"F9D0";
          m(208) := x"FE85";
          m(209) := x"FD1D";
          m(210) := x"0072";
          m(211) := x"FB6C";
          m(212) := x"01B1";
          m(213) := x"FEE9";
          m(214) := x"FE65";
          m(215) := x"00D8";
          m(216) := x"0144";
          m(217) := x"FD3A";
          m(218) := x"FD39";
          m(219) := x"FF4D";
          m(220) := x"02AB";
          m(221) := x"FF0D";
          m(222) := x"0135";
          m(223) := x"0031";
          m(224) := x"FFA6";
          m(225) := x"00B9";
          m(226) := x"00FA";
          m(227) := x"0096";
          m(228) := x"004A";
          m(229) := x"FF99";
          m(230) := x"FDE4";
          m(231) := x"FE3E";
          m(232) := x"023B";
          m(233) := x"002D";
          m(234) := x"FCAC";
          m(235) := x"00B5";
          m(236) := x"0438";
          m(237) := x"FEFB";
          m(238) := x"FC95";
          m(239) := x"FE18";
          m(240) := x"0075";
          m(241) := x"0243";
          m(242) := x"022C";
          m(243) := x"FEBA";
          m(244) := x"03FC";
          m(245) := x"FF84";
          m(246) := x"0076";
          m(247) := x"FF82";
          m(248) := x"FFD3";
          m(249) := x"FE16";
          m(250) := x"00EB";
          m(251) := x"0031";
          m(252) := x"FFF9";
          m(253) := x"0112";
          m(254) := x"009F";
          m(255) := x"FF6D";
          m(256) := x"FE76";
          m(257) := x"FE18";
          m(258) := x"0077";
          m(259) := x"FE00";
          m(260) := x"02C7";
          m(261) := x"01C8";
          m(262) := x"004F";
          m(263) := x"036B";
          m(264) := x"00C1";
          m(265) := x"0139";
          m(266) := x"0031";
          m(267) := x"FDD6";
          m(268) := x"00E0";
          m(269) := x"03BA";
          m(270) := x"015A";
          m(271) := x"FD17";
          m(272) := x"0459";
          m(273) := x"041F";
          m(274) := x"0119";
          m(275) := x"FAC1";
          m(276) := x"FE1A";
          m(277) := x"0059";
          m(278) := x"0083";
          m(279) := x"02B6";
          m(280) := x"0011";
          m(281) := x"00DE";
          m(282) := x"000A";
          m(283) := x"01B2";
          m(284) := x"FFEE";
          m(285) := x"0151";
          m(286) := x"03A4";
          m(287) := x"FE1D";
          m(288) := x"FDD7";
          m(289) := x"04EF";
          m(290) := x"04C4";
          m(291) := x"03F8";
          m(292) := x"FED8";
          m(293) := x"07FE";
          m(294) := x"FBFC";
          m(295) := x"0181";
          m(296) := x"0491";
          m(297) := x"0384";
          m(298) := x"03EA";
          m(299) := x"0114";
          m(300) := x"034C";
          m(301) := x"0572";
          m(302) := x"002C";
          m(303) := x"0037";
          m(304) := x"00CF";
          m(305) := x"040A";
          m(306) := x"0155";
          m(307) := x"00B8";
          m(308) := x"FFE0";
          m(309) := x"0072";
          m(310) := x"0114";
          m(311) := x"032A";
          m(312) := x"0392";
          m(313) := x"0651";
          m(314) := x"04AA";
          m(315) := x"FF7D";
          m(316) := x"00A7";
          m(317) := x"0390";
          m(318) := x"01F4";
          m(319) := x"0561";
          m(320) := x"FAC9";
          m(321) := x"FFD7";
          m(322) := x"019E";
          m(323) := x"036A";
          m(324) := x"FC97";
          m(325) := x"065B";
          m(326) := x"0051";
          m(327) := x"007A";
          m(328) := x"0222";
          m(329) := x"FF68";
          m(330) := x"013F";
          m(331) := x"0237";
          m(332) := x"0014";
          m(333) := x"01A7";
          m(334) := x"0010";
          m(335) := x"0004";
          m(336) := x"0031";
          m(337) := x"FFEE";
          m(338) := x"009B";
          m(339) := x"01EC";
          m(340) := x"015A";
          m(341) := x"0206";
          m(342) := x"00F6";
          m(343) := x"0586";
          m(344) := x"0842";
          m(345) := x"02DC";
          m(346) := x"030F";
          m(347) := x"FBAA";
          m(348) := x"F792";
          m(349) := x"FF3F";
          m(350) := x"FF15";
          m(351) := x"005B";
          m(352) := x"0092";
          m(353) := x"FEC0";
          m(354) := x"FF06";
          m(355) := x"01D6";
          m(356) := x"FF6A";
          m(357) := x"FDB4";
          m(358) := x"0220";
          m(359) := x"FD9E";
          m(360) := x"FE06";
          m(361) := x"0264";
          m(362) := x"0152";
          m(363) := x"004B";
          m(364) := x"0013";
          m(365) := x"FFEC";
          m(366) := x"00CC";
          m(367) := x"0116";
          m(368) := x"0117";
          m(369) := x"FDB3";
          m(370) := x"007A";
          m(371) := x"FF69";
          m(372) := x"FB31";
          m(373) := x"FC04";
          m(374) := x"F91F";
          m(375) := x"F8D8";
          m(376) := x"FCB3";
          m(377) := x"005D";
          m(378) := x"02DD";
          m(379) := x"FD30";
          m(380) := x"011E";
          m(381) := x"01C7";
          m(382) := x"FECE";
          m(383) := x"FCF4";
          m(384) := x"0123";
          m(385) := x"FD8F";
          m(386) := x"FE2F";
          m(387) := x"FB44";
          m(388) := x"FE68";
          m(389) := x"004D";
          m(390) := x"0013";
          m(391) := x"FFC5";
          m(392) := x"001C";
          m(393) := x"0017";
          m(394) := x"0050";
          m(395) := x"00BA";
          m(396) := x"0272";
          m(397) := x"F9B4";
          m(398) := x"FAF7";
          m(399) := x"FA3E";
          m(400) := x"F73E";
          m(401) := x"F6D6";
          m(402) := x"FBF3";
          m(403) := x"F75A";
          m(404) := x"FE71";
          m(405) := x"FA98";
          m(406) := x"FD32";
          m(407) := x"FC33";
          m(408) := x"004A";
          m(409) := x"003A";
          m(410) := x"FAEE";
          m(411) := x"FF3B";
          m(412) := x"03B0";
          m(413) := x"FBD2";
          m(414) := x"FC8E";
          m(415) := x"FE3F";
          m(416) := x"FDA2";
          m(417) := x"FE85";
          m(418) := x"0080";
          m(419) := x"FFC7";
          m(420) := x"0005";
          m(421) := x"FFD4";
          m(422) := x"FFDB";
          m(423) := x"0118";
          m(424) := x"02E3";
          m(425) := x"0451";
          m(426) := x"01D7";
          m(427) := x"FD53";
          m(428) := x"FB3A";
          m(429) := x"FC90";
          m(430) := x"F75C";
          m(431) := x"FA52";
          m(432) := x"FD5A";
          m(433) := x"FB86";
          m(434) := x"FBEA";
          m(435) := x"0387";
          m(436) := x"FC3B";
          m(437) := x"04D7";
          m(438) := x"03BC";
          m(439) := x"04A2";
          m(440) := x"013E";
          m(441) := x"FA97";
          m(442) := x"FBDA";
          m(443) := x"FF07";
          m(444) := x"FD67";
          m(445) := x"FD55";
          m(446) := x"0179";
          m(447) := x"0020";
          m(448) := x"001A";
          m(449) := x"FFFF";
          m(450) := x"000A";
          m(451) := x"0121";
          m(452) := x"05A8";
          m(453) := x"0527";
          m(454) := x"01DF";
          m(455) := x"09C0";
          m(456) := x"0DBC";
          m(457) := x"0BE6";
          m(458) := x"00E2";
          m(459) := x"F942";
          m(460) := x"0154";
          m(461) := x"FD6A";
          m(462) := x"FAE3";
          m(463) := x"FCEF";
          m(464) := x"F7F1";
          m(465) := x"FEBE";
          m(466) := x"035F";
          m(467) := x"07CA";
          m(468) := x"0252";
          m(469) := x"FFF0";
          m(470) := x"FE5E";
          m(471) := x"0055";
          m(472) := x"FD22";
          m(473) := x"FDB6";
          m(474) := x"0156";
          m(475) := x"FFD9";
          m(476) := x"FFF4";
          m(477) := x"FFDC";
          m(478) := x"0020";
          m(479) := x"0059";
          m(480) := x"03CF";
          m(481) := x"079A";
          m(482) := x"088E";
          m(483) := x"0811";
          m(484) := x"0C08";
          m(485) := x"127F";
          m(486) := x"0A75";
          m(487) := x"0932";
          m(488) := x"0830";
          m(489) := x"0383";
          m(490) := x"FE38";
          m(491) := x"010E";
          m(492) := x"FE66";
          m(493) := x"03A9";
          m(494) := x"04AD";
          m(495) := x"020C";
          m(496) := x"01E9";
          m(497) := x"009B";
          m(498) := x"FDD4";
          m(499) := x"FC04";
          m(500) := x"FB4E";
          m(501) := x"FFA0";
          m(502) := x"0024";
          m(503) := x"0027";
          m(504) := x"0018";
          m(505) := x"000A";
          m(506) := x"006B";
          m(507) := x"0058";
          m(508) := x"01AB";
          m(509) := x"0389";
          m(510) := x"021F";
          m(511) := x"038A";
          m(512) := x"03BE";
          m(513) := x"0159";
          m(514) := x"0B02";
          m(515) := x"0FA0";
          m(516) := x"0856";
          m(517) := x"071E";
          m(518) := x"04D1";
          m(519) := x"0133";
          m(520) := x"0112";
          m(521) := x"0283";
          m(522) := x"0012";
          m(523) := x"0238";
          m(524) := x"0477";
          m(525) := x"FD2F";
          m(526) := x"FAD5";
          m(527) := x"FAC6";
          m(528) := x"FB7E";
          m(529) := x"FFCD";
          m(530) := x"FFC7";
          m(531) := x"0037";
          m(532) := x"0026";
          m(533) := x"FFF1";
          m(534) := x"0085";
          m(535) := x"FE3B";
          m(536) := x"FDA2";
          m(537) := x"FEB6";
          m(538) := x"FC74";
          m(539) := x"0441";
          m(540) := x"FBAC";
          m(541) := x"F8CF";
          m(542) := x"FA63";
          m(543) := x"FC54";
          m(544) := x"FEF2";
          m(545) := x"FBB1";
          m(546) := x"FB3E";
          m(547) := x"F957";
          m(548) := x"013C";
          m(549) := x"FE66";
          m(550) := x"FD62";
          m(551) := x"FBE9";
          m(552) := x"00BC";
          m(553) := x"FE37";
          m(554) := x"FBCE";
          m(555) := x"FB5F";
          m(556) := x"FEAF";
          m(557) := x"0089";
          m(558) := x"FFD4";
          m(559) := x"FFD1";
          m(560) := x"FFFA";
          m(561) := x"FFE1";
          m(562) := x"FF91";
          m(563) := x"FD05";
          m(564) := x"FAC5";
          m(565) := x"FBF1";
          m(566) := x"FB6B";
          m(567) := x"F9C2";
          m(568) := x"F942";
          m(569) := x"FCCB";
          m(570) := x"F626";
          m(571) := x"F7A7";
          m(572) := x"F60E";
          m(573) := x"F886";
          m(574) := x"F8E9";
          m(575) := x"FB67";
          m(576) := x"FCE7";
          m(577) := x"FD5A";
          m(578) := x"FBC8";
          m(579) := x"FD5C";
          m(580) := x"FEEE";
          m(581) := x"FF64";
          m(582) := x"FE72";
          m(583) := x"FE74";
          m(584) := x"FFAD";
          m(585) := x"0052";
          m(586) := x"000B";
          m(587) := x"FFF1";
          m(588) := x"FFD4";
          m(589) := x"FFC3";
          m(590) := x"FF73";
          m(591) := x"FD51";
          m(592) := x"FADA";
          m(593) := x"FAFE";
          m(594) := x"F975";
          m(595) := x"F67F";
          m(596) := x"F940";
          m(597) := x"FB80";
          m(598) := x"FC9E";
          m(599) := x"F53D";
          m(600) := x"F8A2";
          m(601) := x"FA94";
          m(602) := x"0127";
          m(603) := x"FF66";
          m(604) := x"FF51";
          m(605) := x"01C3";
          m(606) := x"0145";
          m(607) := x"FE08";
          m(608) := x"FEA2";
          m(609) := x"FFD7";
          m(610) := x"FF2E";
          m(611) := x"FE55";
          m(612) := x"0150";
          m(613) := x"001A";
          m(614) := x"FF98";
          m(615) := x"FFCC";
          m(616) := x"FFDE";
          m(617) := x"0025";
          m(618) := x"FFC2";
          m(619) := x"FEBE";
          m(620) := x"FC83";
          m(621) := x"FB9F";
          m(622) := x"FAAA";
          m(623) := x"FFAF";
          m(624) := x"FF45";
          m(625) := x"FEDE";
          m(626) := x"FE38";
          m(627) := x"F8B1";
          m(628) := x"FFCE";
          m(629) := x"FF9E";
          m(630) := x"FE85";
          m(631) := x"FEBF";
          m(632) := x"FD55";
          m(633) := x"0044";
          m(634) := x"FFCA";
          m(635) := x"F87A";
          m(636) := x"FB95";
          m(637) := x"FD86";
          m(638) := x"FEDF";
          m(639) := x"00B3";
          m(640) := x"0113";
          m(641) := x"004A";
          m(642) := x"FFE5";
          m(643) := x"0060";
          m(644) := x"FFEE";
          m(645) := x"FFE2";
          m(646) := x"FFC0";
          m(647) := x"FFBA";
          m(648) := x"FFB9";
          m(649) := x"FF1A";
          m(650) := x"FE2B";
          m(651) := x"FF03";
          m(652) := x"FCEC";
          m(653) := x"01B7";
          m(654) := x"FC49";
          m(655) := x"F8E7";
          m(656) := x"F9E7";
          m(657) := x"FC43";
          m(658) := x"02D0";
          m(659) := x"FF41";
          m(660) := x"FBA6";
          m(661) := x"0110";
          m(662) := x"FEDA";
          m(663) := x"FCCC";
          m(664) := x"FDB0";
          m(665) := x"FD8B";
          m(666) := x"FF82";
          m(667) := x"0193";
          m(668) := x"010C";
          m(669) := x"000C";
          m(670) := x"001A";
          m(671) := x"FFF0";
          m(672) := x"000C";
          m(673) := x"FFDE";
          m(674) := x"FFBF";
          m(675) := x"FFE3";
          m(676) := x"017B";
          m(677) := x"00CA";
          m(678) := x"0069";
          m(679) := x"012F";
          m(680) := x"0069";
          m(681) := x"FEFE";
          m(682) := x"FF6A";
          m(683) := x"FDC5";
          m(684) := x"FCD9";
          m(685) := x"0121";
          m(686) := x"00D2";
          m(687) := x"028E";
          m(688) := x"FDAF";
          m(689) := x"0389";
          m(690) := x"007B";
          m(691) := x"00B7";
          m(692) := x"0221";
          m(693) := x"0215";
          m(694) := x"015F";
          m(695) := x"01F7";
          m(696) := x"008E";
          m(697) := x"000A";
          m(698) := x"000F";
          m(699) := x"000C";
          m(700) := x"FFFA";
          m(701) := x"FFFB";
          m(702) := x"000F";
          m(703) := x"0023";
          m(704) := x"0214";
          m(705) := x"025A";
          m(706) := x"023A";
          m(707) := x"0428";
          m(708) := x"03DC";
          m(709) := x"0632";
          m(710) := x"016F";
          m(711) := x"03E7";
          m(712) := x"06F5";
          m(713) := x"0326";
          m(714) := x"00CA";
          m(715) := x"017D";
          m(716) := x"0429";
          m(717) := x"0081";
          m(718) := x"0459";
          m(719) := x"0119";
          m(720) := x"001A";
          m(721) := x"0086";
          m(722) := x"0109";
          m(723) := x"019C";
          m(724) := x"00AC";
          m(725) := x"0014";
          m(726) := x"0000";
          m(727) := x"FFFB";
          m(728) := x"001E";
          m(729) := x"0037";
          m(730) := x"FFC5";
          m(731) := x"0000";
          m(732) := x"FEC2";
          m(733) := x"FFF7";
          m(734) := x"011D";
          m(735) := x"02BF";
          m(736) := x"02EB";
          m(737) := x"0247";
          m(738) := x"FF77";
          m(739) := x"00C1";
          m(740) := x"FF51";
          m(741) := x"FEAB";
          m(742) := x"01C4";
          m(743) := x"0303";
          m(744) := x"05E1";
          m(745) := x"00A9";
          m(746) := x"01F6";
          m(747) := x"016B";
          m(748) := x"009D";
          m(749) := x"018B";
          m(750) := x"00BA";
          m(751) := x"FFD1";
          m(752) := x"FFE8";
          m(753) := x"FFFC";
          m(754) := x"0010";
          m(755) := x"FFF0";
          m(756) := x"FFFA";
          m(757) := x"FFDD";
          m(758) := x"FFF5";
          m(759) := x"FFE2";
          m(760) := x"0031";
          m(761) := x"FFC3";
          m(762) := x"FFEF";
          m(763) := x"0008";
          m(764) := x"0016";
          m(765) := x"006C";
          m(766) := x"00AA";
          m(767) := x"FFF2";
          m(768) := x"FFB1";
          m(769) := x"0014";
          m(770) := x"0020";
          m(771) := x"FEAB";
          m(772) := x"FEE1";
          m(773) := x"002B";
          m(774) := x"006D";
          m(775) := x"FFC2";
          m(776) := x"002A";
          m(777) := x"007B";
          m(778) := x"0076";
          m(779) := x"FFEA";
          m(780) := x"0003";
          m(781) := x"FFEE";
          m(782) := x"FFF6";
          m(783) := x"FFFB";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_7.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 7) then
          m(0) := x"FFE9";
          m(1) := x"FFFD";
          m(2) := x"002F";
          m(3) := x"0015";
          m(4) := x"0017";
          m(5) := x"FFAE";
          m(6) := x"0015";
          m(7) := x"FFFE";
          m(8) := x"FFE7";
          m(9) := x"FFFF";
          m(10) := x"0044";
          m(11) := x"0005";
          m(12) := x"FFD5";
          m(13) := x"FFF8";
          m(14) := x"FFF3";
          m(15) := x"003D";
          m(16) := x"FFE4";
          m(17) := x"FFDE";
          m(18) := x"0042";
          m(19) := x"0005";
          m(20) := x"000A";
          m(21) := x"0000";
          m(22) := x"002D";
          m(23) := x"0017";
          m(24) := x"FFE8";
          m(25) := x"FFEF";
          m(26) := x"000F";
          m(27) := x"0012";
          m(28) := x"FFED";
          m(29) := x"0025";
          m(30) := x"0008";
          m(31) := x"FFEA";
          m(32) := x"FFD3";
          m(33) := x"0015";
          m(34) := x"0007";
          m(35) := x"0001";
          m(36) := x"0007";
          m(37) := x"0010";
          m(38) := x"003C";
          m(39) := x"FFC0";
          m(40) := x"0034";
          m(41) := x"002E";
          m(42) := x"006C";
          m(43) := x"00D2";
          m(44) := x"0097";
          m(45) := x"006E";
          m(46) := x"0028";
          m(47) := x"FFDD";
          m(48) := x"0039";
          m(49) := x"FFDD";
          m(50) := x"FFF2";
          m(51) := x"FFF5";
          m(52) := x"0006";
          m(53) := x"FFE3";
          m(54) := x"000F";
          m(55) := x"FFFD";
          m(56) := x"0000";
          m(57) := x"004E";
          m(58) := x"0003";
          m(59) := x"0002";
          m(60) := x"FFE1";
          m(61) := x"0034";
          m(62) := x"0012";
          m(63) := x"0051";
          m(64) := x"0088";
          m(65) := x"0069";
          m(66) := x"0072";
          m(67) := x"00C1";
          m(68) := x"00B3";
          m(69) := x"0033";
          m(70) := x"00C3";
          m(71) := x"003A";
          m(72) := x"FF39";
          m(73) := x"0068";
          m(74) := x"FFFC";
          m(75) := x"FFD4";
          m(76) := x"000F";
          m(77) := x"0021";
          m(78) := x"FFEB";
          m(79) := x"001C";
          m(80) := x"0010";
          m(81) := x"003B";
          m(82) := x"FFF7";
          m(83) := x"0002";
          m(84) := x"FFDE";
          m(85) := x"FFD1";
          m(86) := x"FFFE";
          m(87) := x"FFF1";
          m(88) := x"FFE8";
          m(89) := x"0030";
          m(90) := x"FFEF";
          m(91) := x"FFDF";
          m(92) := x"FFFF";
          m(93) := x"0062";
          m(94) := x"0037";
          m(95) := x"FFD6";
          m(96) := x"FA3C";
          m(97) := x"F94D";
          m(98) := x"FBB3";
          m(99) := x"FB36";
          m(100) := x"FC2D";
          m(101) := x"FE13";
          m(102) := x"FE42";
          m(103) := x"FDA5";
          m(104) := x"FE9E";
          m(105) := x"00E0";
          m(106) := x"00A9";
          m(107) := x"0004";
          m(108) := x"FFE7";
          m(109) := x"FFC9";
          m(110) := x"FFF8";
          m(111) := x"FFE5";
          m(112) := x"FFC5";
          m(113) := x"002B";
          m(114) := x"0014";
          m(115) := x"003C";
          m(116) := x"FFF9";
          m(117) := x"FF84";
          m(118) := x"FF2B";
          m(119) := x"FDE5";
          m(120) := x"FD29";
          m(121) := x"FE1E";
          m(122) := x"FE0E";
          m(123) := x"FD73";
          m(124) := x"FD99";
          m(125) := x"FD56";
          m(126) := x"01A9";
          m(127) := x"FEAC";
          m(128) := x"02B2";
          m(129) := x"06C4";
          m(130) := x"FE25";
          m(131) := x"001D";
          m(132) := x"0158";
          m(133) := x"014C";
          m(134) := x"0207";
          m(135) := x"0019";
          m(136) := x"016A";
          m(137) := x"FF50";
          m(138) := x"FF9F";
          m(139) := x"003A";
          m(140) := x"FFF5";
          m(141) := x"FFE3";
          m(142) := x"0013";
          m(143) := x"FFD8";
          m(144) := x"000B";
          m(145) := x"FE06";
          m(146) := x"FE06";
          m(147) := x"FEB7";
          m(148) := x"FE4B";
          m(149) := x"FEDD";
          m(150) := x"FE7C";
          m(151) := x"03A8";
          m(152) := x"0411";
          m(153) := x"FD6C";
          m(154) := x"0311";
          m(155) := x"01AA";
          m(156) := x"FE29";
          m(157) := x"0279";
          m(158) := x"FFE6";
          m(159) := x"FFF4";
          m(160) := x"FC7B";
          m(161) := x"0358";
          m(162) := x"0210";
          m(163) := x"FFD4";
          m(164) := x"FEF6";
          m(165) := x"FF29";
          m(166) := x"FFFC";
          m(167) := x"0035";
          m(168) := x"FFDF";
          m(169) := x"FFD2";
          m(170) := x"FFCB";
          m(171) := x"FFB3";
          m(172) := x"FFF1";
          m(173) := x"FD13";
          m(174) := x"FF51";
          m(175) := x"0046";
          m(176) := x"0000";
          m(177) := x"FEE4";
          m(178) := x"0148";
          m(179) := x"FF13";
          m(180) := x"0075";
          m(181) := x"0305";
          m(182) := x"0063";
          m(183) := x"FCCE";
          m(184) := x"FD98";
          m(185) := x"046B";
          m(186) := x"0394";
          m(187) := x"05A8";
          m(188) := x"0298";
          m(189) := x"0473";
          m(190) := x"0592";
          m(191) := x"0152";
          m(192) := x"F9F0";
          m(193) := x"FB6E";
          m(194) := x"FF32";
          m(195) := x"FFE1";
          m(196) := x"FFE3";
          m(197) := x"0008";
          m(198) := x"FFDC";
          m(199) := x"FEF3";
          m(200) := x"00AB";
          m(201) := x"FF44";
          m(202) := x"FCE2";
          m(203) := x"FC5F";
          m(204) := x"FFDF";
          m(205) := x"01BE";
          m(206) := x"FFAF";
          m(207) := x"FCD9";
          m(208) := x"FD28";
          m(209) := x"FFB1";
          m(210) := x"FBD4";
          m(211) := x"072D";
          m(212) := x"016F";
          m(213) := x"0060";
          m(214) := x"0479";
          m(215) := x"028D";
          m(216) := x"FAC6";
          m(217) := x"00A6";
          m(218) := x"02E6";
          m(219) := x"0097";
          m(220) := x"F6F0";
          m(221) := x"FB8A";
          m(222) := x"FE8C";
          m(223) := x"FFD0";
          m(224) := x"FFAC";
          m(225) := x"FFC4";
          m(226) := x"FFFE";
          m(227) := x"FF4E";
          m(228) := x"009E";
          m(229) := x"FF05";
          m(230) := x"FF32";
          m(231) := x"01C0";
          m(232) := x"FFB3";
          m(233) := x"007F";
          m(234) := x"0111";
          m(235) := x"01CF";
          m(236) := x"FF65";
          m(237) := x"FEE5";
          m(238) := x"FFD0";
          m(239) := x"FE11";
          m(240) := x"0068";
          m(241) := x"FEBB";
          m(242) := x"01DA";
          m(243) := x"03AD";
          m(244) := x"FED6";
          m(245) := x"0197";
          m(246) := x"01B3";
          m(247) := x"FDAC";
          m(248) := x"F8AD";
          m(249) := x"FCA3";
          m(250) := x"FEE0";
          m(251) := x"FFE7";
          m(252) := x"FFFF";
          m(253) := x"FFAD";
          m(254) := x"0065";
          m(255) := x"002E";
          m(256) := x"FDE3";
          m(257) := x"0001";
          m(258) := x"FF3C";
          m(259) := x"01F3";
          m(260) := x"FFCA";
          m(261) := x"0060";
          m(262) := x"0642";
          m(263) := x"04A8";
          m(264) := x"FC34";
          m(265) := x"FA23";
          m(266) := x"FE1F";
          m(267) := x"FC93";
          m(268) := x"FAD0";
          m(269) := x"00D6";
          m(270) := x"FF53";
          m(271) := x"FF83";
          m(272) := x"02D5";
          m(273) := x"0483";
          m(274) := x"0023";
          m(275) := x"FFE7";
          m(276) := x"FB29";
          m(277) := x"FCB9";
          m(278) := x"FFDD";
          m(279) := x"FFF6";
          m(280) := x"000A";
          m(281) := x"FFD2";
          m(282) := x"001D";
          m(283) := x"FF70";
          m(284) := x"FF3E";
          m(285) := x"0080";
          m(286) := x"0030";
          m(287) := x"01A8";
          m(288) := x"FFB7";
          m(289) := x"008B";
          m(290) := x"051A";
          m(291) := x"FFC4";
          m(292) := x"FEC9";
          m(293) := x"FB4F";
          m(294) := x"0411";
          m(295) := x"04C6";
          m(296) := x"0632";
          m(297) := x"03DF";
          m(298) := x"FFB5";
          m(299) := x"06DC";
          m(300) := x"02D7";
          m(301) := x"0128";
          m(302) := x"008E";
          m(303) := x"02DA";
          m(304) := x"FCB1";
          m(305) := x"FC79";
          m(306) := x"FF74";
          m(307) := x"0008";
          m(308) := x"FFE8";
          m(309) := x"FFC0";
          m(310) := x"FF3F";
          m(311) := x"005F";
          m(312) := x"FFD7";
          m(313) := x"FEA8";
          m(314) := x"FDB5";
          m(315) := x"0253";
          m(316) := x"03C7";
          m(317) := x"062F";
          m(318) := x"06E9";
          m(319) := x"028B";
          m(320) := x"FE13";
          m(321) := x"FE40";
          m(322) := x"0651";
          m(323) := x"047A";
          m(324) := x"02F1";
          m(325) := x"FC23";
          m(326) := x"F9E9";
          m(327) := x"0063";
          m(328) := x"044E";
          m(329) := x"049D";
          m(330) := x"03B6";
          m(331) := x"02CF";
          m(332) := x"00B4";
          m(333) := x"FD15";
          m(334) := x"FF41";
          m(335) := x"0032";
          m(336) := x"FFF1";
          m(337) := x"0000";
          m(338) := x"FFA3";
          m(339) := x"00F2";
          m(340) := x"FF8B";
          m(341) := x"FFF1";
          m(342) := x"FD39";
          m(343) := x"008B";
          m(344) := x"FF19";
          m(345) := x"FFBB";
          m(346) := x"F8AC";
          m(347) := x"FC36";
          m(348) := x"FF26";
          m(349) := x"019A";
          m(350) := x"077D";
          m(351) := x"0939";
          m(352) := x"04D7";
          m(353) := x"0673";
          m(354) := x"FD7A";
          m(355) := x"01F4";
          m(356) := x"01C7";
          m(357) := x"032D";
          m(358) := x"FF08";
          m(359) := x"027E";
          m(360) := x"029E";
          m(361) := x"0096";
          m(362) := x"FFFF";
          m(363) := x"FFF4";
          m(364) := x"FFF9";
          m(365) := x"0033";
          m(366) := x"FFB9";
          m(367) := x"00E0";
          m(368) := x"FFA9";
          m(369) := x"FE8F";
          m(370) := x"FC48";
          m(371) := x"0246";
          m(372) := x"0386";
          m(373) := x"FEB4";
          m(374) := x"FA0F";
          m(375) := x"00B3";
          m(376) := x"04A8";
          m(377) := x"076A";
          m(378) := x"03AD";
          m(379) := x"096C";
          m(380) := x"00D5";
          m(381) := x"02E1";
          m(382) := x"048B";
          m(383) := x"0137";
          m(384) := x"FDEB";
          m(385) := x"FE5D";
          m(386) := x"01B4";
          m(387) := x"004F";
          m(388) := x"FEA1";
          m(389) := x"00E9";
          m(390) := x"FFE9";
          m(391) := x"FFFC";
          m(392) := x"0070";
          m(393) := x"FFDD";
          m(394) := x"FFB8";
          m(395) := x"FFAE";
          m(396) := x"0095";
          m(397) := x"000F";
          m(398) := x"FC82";
          m(399) := x"FD86";
          m(400) := x"FEA0";
          m(401) := x"FB8A";
          m(402) := x"00A7";
          m(403) := x"04C3";
          m(404) := x"0530";
          m(405) := x"071E";
          m(406) := x"FDF0";
          m(407) := x"0035";
          m(408) := x"0489";
          m(409) := x"02BC";
          m(410) := x"FE6D";
          m(411) := x"0209";
          m(412) := x"FF6A";
          m(413) := x"FC9E";
          m(414) := x"FCBA";
          m(415) := x"FA36";
          m(416) := x"FD6B";
          m(417) := x"016A";
          m(418) := x"0025";
          m(419) := x"0029";
          m(420) := x"FFF7";
          m(421) := x"FF9C";
          m(422) := x"FFDD";
          m(423) := x"FFF3";
          m(424) := x"FF7F";
          m(425) := x"FEF8";
          m(426) := x"FD23";
          m(427) := x"FEED";
          m(428) := x"05B9";
          m(429) := x"FDBD";
          m(430) := x"0168";
          m(431) := x"0291";
          m(432) := x"023C";
          m(433) := x"04AE";
          m(434) := x"0396";
          m(435) := x"044E";
          m(436) := x"05EA";
          m(437) := x"0880";
          m(438) := x"0348";
          m(439) := x"FDC8";
          m(440) := x"FB53";
          m(441) := x"FAD8";
          m(442) := x"FE72";
          m(443) := x"FB9F";
          m(444) := x"FD82";
          m(445) := x"01C7";
          m(446) := x"FFDD";
          m(447) := x"FFFD";
          m(448) := x"0007";
          m(449) := x"FFDD";
          m(450) := x"FF82";
          m(451) := x"FFE8";
          m(452) := x"FF46";
          m(453) := x"FFAB";
          m(454) := x"0256";
          m(455) := x"077B";
          m(456) := x"084F";
          m(457) := x"06D9";
          m(458) := x"FD47";
          m(459) := x"0082";
          m(460) := x"FEA2";
          m(461) := x"0059";
          m(462) := x"06BF";
          m(463) := x"05ED";
          m(464) := x"05A7";
          m(465) := x"00D8";
          m(466) := x"FC21";
          m(467) := x"FBE0";
          m(468) := x"F919";
          m(469) := x"F689";
          m(470) := x"FA7E";
          m(471) := x"FEBE";
          m(472) := x"FECF";
          m(473) := x"01E1";
          m(474) := x"0039";
          m(475) := x"000E";
          m(476) := x"FFF0";
          m(477) := x"000F";
          m(478) := x"FF95";
          m(479) := x"FEA9";
          m(480) := x"FE05";
          m(481) := x"FF81";
          m(482) := x"04A1";
          m(483) := x"00D1";
          m(484) := x"04A5";
          m(485) := x"0883";
          m(486) := x"08B1";
          m(487) := x"06C8";
          m(488) := x"065F";
          m(489) := x"0AC2";
          m(490) := x"0399";
          m(491) := x"0518";
          m(492) := x"0453";
          m(493) := x"FCFF";
          m(494) := x"F73C";
          m(495) := x"F710";
          m(496) := x"F9E4";
          m(497) := x"F976";
          m(498) := x"FD2D";
          m(499) := x"FE27";
          m(500) := x"0347";
          m(501) := x"006E";
          m(502) := x"003F";
          m(503) := x"FFED";
          m(504) := x"FFE3";
          m(505) := x"0002";
          m(506) := x"FF6C";
          m(507) := x"FEF7";
          m(508) := x"FD63";
          m(509) := x"0120";
          m(510) := x"04CA";
          m(511) := x"0213";
          m(512) := x"0229";
          m(513) := x"095E";
          m(514) := x"0A23";
          m(515) := x"0E6C";
          m(516) := x"1296";
          m(517) := x"0EAC";
          m(518) := x"FF69";
          m(519) := x"FF5B";
          m(520) := x"F8E3";
          m(521) := x"F9C5";
          m(522) := x"F683";
          m(523) := x"F739";
          m(524) := x"FAA3";
          m(525) := x"F9F9";
          m(526) := x"FC78";
          m(527) := x"FF37";
          m(528) := x"0318";
          m(529) := x"0007";
          m(530) := x"002D";
          m(531) := x"FFBA";
          m(532) := x"FFFF";
          m(533) := x"FFF7";
          m(534) := x"FFC1";
          m(535) := x"FF46";
          m(536) := x"FF21";
          m(537) := x"0198";
          m(538) := x"04C7";
          m(539) := x"01FF";
          m(540) := x"02AA";
          m(541) := x"079F";
          m(542) := x"0686";
          m(543) := x"046A";
          m(544) := x"02AA";
          m(545) := x"051F";
          m(546) := x"F961";
          m(547) := x"F8C3";
          m(548) := x"F863";
          m(549) := x"FB59";
          m(550) := x"F9B0";
          m(551) := x"FCFE";
          m(552) := x"FE15";
          m(553) := x"0020";
          m(554) := x"FF0F";
          m(555) := x"FFD6";
          m(556) := x"0083";
          m(557) := x"FF5E";
          m(558) := x"0019";
          m(559) := x"001A";
          m(560) := x"FFEF";
          m(561) := x"FFCC";
          m(562) := x"0005";
          m(563) := x"FE7A";
          m(564) := x"FFEA";
          m(565) := x"0031";
          m(566) := x"041F";
          m(567) := x"00AA";
          m(568) := x"FFB6";
          m(569) := x"FDF7";
          m(570) := x"FB6B";
          m(571) := x"FBB2";
          m(572) := x"FCA4";
          m(573) := x"F7BD";
          m(574) := x"F793";
          m(575) := x"F99A";
          m(576) := x"F7DE";
          m(577) := x"F86D";
          m(578) := x"FEB5";
          m(579) := x"02B7";
          m(580) := x"03AD";
          m(581) := x"0009";
          m(582) := x"FAFA";
          m(583) := x"FFD5";
          m(584) := x"FFB3";
          m(585) := x"FFE3";
          m(586) := x"FFFF";
          m(587) := x"0006";
          m(588) := x"FFCE";
          m(589) := x"003E";
          m(590) := x"000B";
          m(591) := x"FE7A";
          m(592) := x"FCE9";
          m(593) := x"FEB3";
          m(594) := x"000E";
          m(595) := x"FE7E";
          m(596) := x"FB90";
          m(597) := x"FD45";
          m(598) := x"FBAD";
          m(599) := x"F80B";
          m(600) := x"F8FB";
          m(601) := x"FB28";
          m(602) := x"FBB0";
          m(603) := x"FA3E";
          m(604) := x"0098";
          m(605) := x"0091";
          m(606) := x"FC75";
          m(607) := x"FEF3";
          m(608) := x"F9D6";
          m(609) := x"FD0D";
          m(610) := x"FC74";
          m(611) := x"00BF";
          m(612) := x"0083";
          m(613) := x"0062";
          m(614) := x"001A";
          m(615) := x"FFF9";
          m(616) := x"FFF2";
          m(617) := x"FFEB";
          m(618) := x"FFF7";
          m(619) := x"FEBF";
          m(620) := x"FDF8";
          m(621) := x"FD05";
          m(622) := x"FCC6";
          m(623) := x"FFB9";
          m(624) := x"FE45";
          m(625) := x"FF6F";
          m(626) := x"FE4D";
          m(627) := x"FE6C";
          m(628) := x"F7A7";
          m(629) := x"FD17";
          m(630) := x"FFE0";
          m(631) := x"FB3F";
          m(632) := x"FC13";
          m(633) := x"FADF";
          m(634) := x"FE7F";
          m(635) := x"FF09";
          m(636) := x"FF2A";
          m(637) := x"FFD3";
          m(638) := x"FF61";
          m(639) := x"00C6";
          m(640) := x"00DD";
          m(641) := x"0069";
          m(642) := x"000C";
          m(643) := x"FFFB";
          m(644) := x"0017";
          m(645) := x"0001";
          m(646) := x"FFF6";
          m(647) := x"FF44";
          m(648) := x"FD06";
          m(649) := x"FC9D";
          m(650) := x"FC8F";
          m(651) := x"0095";
          m(652) := x"FF89";
          m(653) := x"FCB1";
          m(654) := x"F717";
          m(655) := x"F69C";
          m(656) := x"FF76";
          m(657) := x"00E4";
          m(658) := x"FD0A";
          m(659) := x"FB9F";
          m(660) := x"0221";
          m(661) := x"02EA";
          m(662) := x"0478";
          m(663) := x"0491";
          m(664) := x"02E2";
          m(665) := x"0326";
          m(666) := x"0265";
          m(667) := x"0178";
          m(668) := x"0114";
          m(669) := x"005E";
          m(670) := x"0014";
          m(671) := x"000E";
          m(672) := x"0016";
          m(673) := x"0013";
          m(674) := x"0002";
          m(675) := x"FF6F";
          m(676) := x"FF1D";
          m(677) := x"FF2B";
          m(678) := x"FE29";
          m(679) := x"F7E3";
          m(680) := x"F8FB";
          m(681) := x"F8AC";
          m(682) := x"F9F7";
          m(683) := x"F975";
          m(684) := x"FFEF";
          m(685) := x"010D";
          m(686) := x"FC6A";
          m(687) := x"F82E";
          m(688) := x"FE43";
          m(689) := x"FB02";
          m(690) := x"00F1";
          m(691) := x"06F9";
          m(692) := x"0421";
          m(693) := x"016C";
          m(694) := x"FFE4";
          m(695) := x"00C9";
          m(696) := x"00A3";
          m(697) := x"00A1";
          m(698) := x"FFDD";
          m(699) := x"0008";
          m(700) := x"FFC7";
          m(701) := x"FFF4";
          m(702) := x"0004";
          m(703) := x"FFB1";
          m(704) := x"FFCF";
          m(705) := x"FFF1";
          m(706) := x"008A";
          m(707) := x"FE95";
          m(708) := x"FCB1";
          m(709) := x"FA59";
          m(710) := x"FD55";
          m(711) := x"FA47";
          m(712) := x"F92A";
          m(713) := x"F817";
          m(714) := x"FD79";
          m(715) := x"FE87";
          m(716) := x"FF9E";
          m(717) := x"00F7";
          m(718) := x"0000";
          m(719) := x"FF73";
          m(720) := x"FF86";
          m(721) := x"FE93";
          m(722) := x"FE21";
          m(723) := x"FF6F";
          m(724) := x"FFFA";
          m(725) := x"FFDC";
          m(726) := x"004C";
          m(727) := x"0008";
          m(728) := x"0012";
          m(729) := x"000D";
          m(730) := x"000D";
          m(731) := x"001A";
          m(732) := x"001A";
          m(733) := x"005A";
          m(734) := x"007F";
          m(735) := x"007C";
          m(736) := x"FFF6";
          m(737) := x"FEA1";
          m(738) := x"FCF9";
          m(739) := x"FBF3";
          m(740) := x"FE56";
          m(741) := x"FDDD";
          m(742) := x"FF7F";
          m(743) := x"FF5F";
          m(744) := x"FCC4";
          m(745) := x"0096";
          m(746) := x"FF63";
          m(747) := x"FE86";
          m(748) := x"FEF1";
          m(749) := x"FE92";
          m(750) := x"FEFF";
          m(751) := x"FFC9";
          m(752) := x"0007";
          m(753) := x"FFD3";
          m(754) := x"FFBB";
          m(755) := x"0024";
          m(756) := x"0013";
          m(757) := x"001C";
          m(758) := x"0001";
          m(759) := x"FFE9";
          m(760) := x"FFDF";
          m(761) := x"0019";
          m(762) := x"FFE2";
          m(763) := x"FFEE";
          m(764) := x"FFF2";
          m(765) := x"000B";
          m(766) := x"0012";
          m(767) := x"0003";
          m(768) := x"003D";
          m(769) := x"FFC9";
          m(770) := x"FFCC";
          m(771) := x"0121";
          m(772) := x"0089";
          m(773) := x"FFFE";
          m(774) := x"0059";
          m(775) := x"0022";
          m(776) := x"0004";
          m(777) := x"FFB3";
          m(778) := x"FF61";
          m(779) := x"FFFF";
          m(780) := x"004C";
          m(781) := x"002F";
          m(782) := x"FFEF";
          m(783) := x"FFFD";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_8.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 8) then
          m(0) := x"FFFD";
          m(1) := x"0000";
          m(2) := x"FFD7";
          m(3) := x"FFE4";
          m(4) := x"0009";
          m(5) := x"0005";
          m(6) := x"0000";
          m(7) := x"FFF1";
          m(8) := x"FFE3";
          m(9) := x"FFE2";
          m(10) := x"FFFB";
          m(11) := x"0010";
          m(12) := x"FFF7";
          m(13) := x"FFEE";
          m(14) := x"0007";
          m(15) := x"0002";
          m(16) := x"0027";
          m(17) := x"0003";
          m(18) := x"0002";
          m(19) := x"FFFC";
          m(20) := x"0005";
          m(21) := x"FFED";
          m(22) := x"FFF2";
          m(23) := x"FFD5";
          m(24) := x"0029";
          m(25) := x"0004";
          m(26) := x"0012";
          m(27) := x"FFEA";
          m(28) := x"0001";
          m(29) := x"000E";
          m(30) := x"0021";
          m(31) := x"001C";
          m(32) := x"FFE3";
          m(33) := x"0033";
          m(34) := x"FFDA";
          m(35) := x"0000";
          m(36) := x"0011";
          m(37) := x"FFE3";
          m(38) := x"FFE8";
          m(39) := x"FFBF";
          m(40) := x"FFAA";
          m(41) := x"FF90";
          m(42) := x"FFB5";
          m(43) := x"FFA4";
          m(44) := x"FFD4";
          m(45) := x"FFB7";
          m(46) := x"0000";
          m(47) := x"FFDB";
          m(48) := x"0018";
          m(49) := x"0026";
          m(50) := x"0012";
          m(51) := x"000D";
          m(52) := x"FFFF";
          m(53) := x"0036";
          m(54) := x"FFE4";
          m(55) := x"FFDF";
          m(56) := x"FFE2";
          m(57) := x"FFF6";
          m(58) := x"FFD2";
          m(59) := x"FFD1";
          m(60) := x"FFFB";
          m(61) := x"0000";
          m(62) := x"FFFA";
          m(63) := x"001D";
          m(64) := x"0015";
          m(65) := x"0068";
          m(66) := x"FFCF";
          m(67) := x"FF86";
          m(68) := x"FE83";
          m(69) := x"FE95";
          m(70) := x"FEF5";
          m(71) := x"FE93";
          m(72) := x"FD91";
          m(73) := x"FD63";
          m(74) := x"FE5A";
          m(75) := x"0068";
          m(76) := x"00F9";
          m(77) := x"005A";
          m(78) := x"FFEB";
          m(79) := x"0028";
          m(80) := x"FFFE";
          m(81) := x"FFD3";
          m(82) := x"FFC5";
          m(83) := x"FFCA";
          m(84) := x"0000";
          m(85) := x"0024";
          m(86) := x"001F";
          m(87) := x"FFEF";
          m(88) := x"FFEA";
          m(89) := x"FFF2";
          m(90) := x"FFE5";
          m(91) := x"FFD0";
          m(92) := x"FE63";
          m(93) := x"FE25";
          m(94) := x"FDFB";
          m(95) := x"FDDF";
          m(96) := x"FC8F";
          m(97) := x"FBF6";
          m(98) := x"FD55";
          m(99) := x"FB37";
          m(100) := x"FA39";
          m(101) := x"FDE3";
          m(102) := x"FC91";
          m(103) := x"FE63";
          m(104) := x"00DD";
          m(105) := x"FF7E";
          m(106) := x"FF3C";
          m(107) := x"FFB5";
          m(108) := x"0008";
          m(109) := x"002C";
          m(110) := x"001A";
          m(111) := x"0020";
          m(112) := x"FFE1";
          m(113) := x"FFF0";
          m(114) := x"000A";
          m(115) := x"000A";
          m(116) := x"000B";
          m(117) := x"014F";
          m(118) := x"020D";
          m(119) := x"0265";
          m(120) := x"02EC";
          m(121) := x"0238";
          m(122) := x"FF92";
          m(123) := x"00F7";
          m(124) := x"00C5";
          m(125) := x"027D";
          m(126) := x"0237";
          m(127) := x"FD8D";
          m(128) := x"FC9C";
          m(129) := x"FD31";
          m(130) := x"FAD3";
          m(131) := x"FEFB";
          m(132) := x"FCD4";
          m(133) := x"FCE8";
          m(134) := x"FDA8";
          m(135) := x"FF3E";
          m(136) := x"0010";
          m(137) := x"000E";
          m(138) := x"0011";
          m(139) := x"FFE3";
          m(140) := x"FFF9";
          m(141) := x"001A";
          m(142) := x"FFE2";
          m(143) := x"009F";
          m(144) := x"0271";
          m(145) := x"02E9";
          m(146) := x"03F6";
          m(147) := x"0554";
          m(148) := x"01BF";
          m(149) := x"0090";
          m(150) := x"FBF7";
          m(151) := x"F991";
          m(152) := x"010D";
          m(153) := x"FB7E";
          m(154) := x"0050";
          m(155) := x"FCBA";
          m(156) := x"022D";
          m(157) := x"0350";
          m(158) := x"FCD6";
          m(159) := x"00FC";
          m(160) := x"0186";
          m(161) := x"FD7C";
          m(162) := x"FD11";
          m(163) := x"FDAF";
          m(164) := x"FF41";
          m(165) := x"0030";
          m(166) := x"FFDF";
          m(167) := x"000B";
          m(168) := x"FFF9";
          m(169) := x"0005";
          m(170) := x"001E";
          m(171) := x"010B";
          m(172) := x"02D6";
          m(173) := x"01A1";
          m(174) := x"0634";
          m(175) := x"00B8";
          m(176) := x"01A5";
          m(177) := x"FEAA";
          m(178) := x"FB12";
          m(179) := x"FB67";
          m(180) := x"FFEC";
          m(181) := x"FE40";
          m(182) := x"FD2F";
          m(183) := x"FFCB";
          m(184) := x"FC86";
          m(185) := x"0226";
          m(186) := x"00E7";
          m(187) := x"FF40";
          m(188) := x"03BB";
          m(189) := x"051C";
          m(190) := x"0260";
          m(191) := x"FE40";
          m(192) := x"FEC4";
          m(193) := x"FFC2";
          m(194) := x"FFD7";
          m(195) := x"001D";
          m(196) := x"FFEF";
          m(197) := x"0005";
          m(198) := x"FFCF";
          m(199) := x"0262";
          m(200) := x"04C3";
          m(201) := x"01AA";
          m(202) := x"0180";
          m(203) := x"FDF5";
          m(204) := x"04F1";
          m(205) := x"FE9F";
          m(206) := x"FB0C";
          m(207) := x"FAAF";
          m(208) := x"FD44";
          m(209) := x"0269";
          m(210) := x"FE9C";
          m(211) := x"FFF3";
          m(212) := x"0344";
          m(213) := x"05B2";
          m(214) := x"0470";
          m(215) := x"0051";
          m(216) := x"03A5";
          m(217) := x"039B";
          m(218) := x"0478";
          m(219) := x"FF84";
          m(220) := x"FD9C";
          m(221) := x"0076";
          m(222) := x"FF99";
          m(223) := x"001B";
          m(224) := x"FFDE";
          m(225) := x"0003";
          m(226) := x"FFEC";
          m(227) := x"01B0";
          m(228) := x"02A9";
          m(229) := x"0119";
          m(230) := x"0132";
          m(231) := x"043C";
          m(232) := x"FD9F";
          m(233) := x"0256";
          m(234) := x"010C";
          m(235) := x"FD21";
          m(236) := x"FECE";
          m(237) := x"085D";
          m(238) := x"01DC";
          m(239) := x"F950";
          m(240) := x"0602";
          m(241) := x"0670";
          m(242) := x"FFF1";
          m(243) := x"0222";
          m(244) := x"02A0";
          m(245) := x"FCD9";
          m(246) := x"0213";
          m(247) := x"02A8";
          m(248) := x"FD34";
          m(249) := x"FFF4";
          m(250) := x"019E";
          m(251) := x"0013";
          m(252) := x"FFE3";
          m(253) := x"0010";
          m(254) := x"001F";
          m(255) := x"0152";
          m(256) := x"0353";
          m(257) := x"FF8A";
          m(258) := x"FD6B";
          m(259) := x"0148";
          m(260) := x"FB54";
          m(261) := x"FCC3";
          m(262) := x"F8C3";
          m(263) := x"F58C";
          m(264) := x"FD93";
          m(265) := x"0908";
          m(266) := x"02D5";
          m(267) := x"F942";
          m(268) := x"0066";
          m(269) := x"0281";
          m(270) := x"03F2";
          m(271) := x"0873";
          m(272) := x"011D";
          m(273) := x"005F";
          m(274) := x"06FE";
          m(275) := x"012C";
          m(276) := x"0122";
          m(277) := x"012C";
          m(278) := x"003E";
          m(279) := x"0000";
          m(280) := x"001A";
          m(281) := x"FFF6";
          m(282) := x"0036";
          m(283) := x"00C2";
          m(284) := x"023C";
          m(285) := x"FD98";
          m(286) := x"FAE5";
          m(287) := x"FD76";
          m(288) := x"FCBC";
          m(289) := x"FBD4";
          m(290) := x"FA6B";
          m(291) := x"FB9C";
          m(292) := x"0016";
          m(293) := x"04CE";
          m(294) := x"0666";
          m(295) := x"FA29";
          m(296) := x"01B5";
          m(297) := x"FC20";
          m(298) := x"FEE2";
          m(299) := x"0265";
          m(300) := x"FBBC";
          m(301) := x"FDB8";
          m(302) := x"0325";
          m(303) := x"0212";
          m(304) := x"FEAC";
          m(305) := x"FE34";
          m(306) := x"0088";
          m(307) := x"FFF6";
          m(308) := x"FFEE";
          m(309) := x"FFF5";
          m(310) := x"0000";
          m(311) := x"FEF8";
          m(312) := x"00CA";
          m(313) := x"0313";
          m(314) := x"FAFD";
          m(315) := x"FDC3";
          m(316) := x"FF8F";
          m(317) := x"F9A4";
          m(318) := x"F9AF";
          m(319) := x"0201";
          m(320) := x"047E";
          m(321) := x"0977";
          m(322) := x"0707";
          m(323) := x"F952";
          m(324) := x"F9F1";
          m(325) := x"FA98";
          m(326) := x"FBD4";
          m(327) := x"0019";
          m(328) := x"FB51";
          m(329) := x"FC49";
          m(330) := x"FEFF";
          m(331) := x"FEF6";
          m(332) := x"FC34";
          m(333) := x"008A";
          m(334) := x"01DA";
          m(335) := x"FFF7";
          m(336) := x"0011";
          m(337) := x"FFD7";
          m(338) := x"FFC1";
          m(339) := x"FCD2";
          m(340) := x"FBEC";
          m(341) := x"00A6";
          m(342) := x"FF62";
          m(343) := x"FD30";
          m(344) := x"FB83";
          m(345) := x"FCC4";
          m(346) := x"F9BF";
          m(347) := x"00E0";
          m(348) := x"0A53";
          m(349) := x"0CB6";
          m(350) := x"02E4";
          m(351) := x"FF63";
          m(352) := x"0479";
          m(353) := x"FCD9";
          m(354) := x"FF26";
          m(355) := x"0048";
          m(356) := x"FEA7";
          m(357) := x"FCC3";
          m(358) := x"FDAC";
          m(359) := x"F9D3";
          m(360) := x"FEA3";
          m(361) := x"00B5";
          m(362) := x"00F7";
          m(363) := x"0025";
          m(364) := x"0007";
          m(365) := x"FFC9";
          m(366) := x"0005";
          m(367) := x"FD96";
          m(368) := x"F836";
          m(369) := x"FB42";
          m(370) := x"FF23";
          m(371) := x"F777";
          m(372) := x"FE96";
          m(373) := x"FB88";
          m(374) := x"FA9C";
          m(375) := x"0448";
          m(376) := x"0781";
          m(377) := x"0AE2";
          m(378) := x"0742";
          m(379) := x"0131";
          m(380) := x"002C";
          m(381) := x"FE2F";
          m(382) := x"0351";
          m(383) := x"FF2B";
          m(384) := x"02E9";
          m(385) := x"FED0";
          m(386) := x"FB38";
          m(387) := x"FE23";
          m(388) := x"FDA2";
          m(389) := x"FEEF";
          m(390) := x"0161";
          m(391) := x"0119";
          m(392) := x"0033";
          m(393) := x"FF7F";
          m(394) := x"FFC5";
          m(395) := x"FD9D";
          m(396) := x"F7B6";
          m(397) := x"FC42";
          m(398) := x"F7D4";
          m(399) := x"F6B3";
          m(400) := x"FAB6";
          m(401) := x"FC93";
          m(402) := x"FD0B";
          m(403) := x"02C8";
          m(404) := x"095E";
          m(405) := x"072B";
          m(406) := x"0569";
          m(407) := x"0017";
          m(408) := x"FE37";
          m(409) := x"FDF8";
          m(410) := x"FDD4";
          m(411) := x"020A";
          m(412) := x"FF49";
          m(413) := x"FFE5";
          m(414) := x"FAAA";
          m(415) := x"FDC0";
          m(416) := x"FDB6";
          m(417) := x"FFE0";
          m(418) := x"0181";
          m(419) := x"FFE5";
          m(420) := x"FFCC";
          m(421) := x"FFEE";
          m(422) := x"FFD8";
          m(423) := x"FE16";
          m(424) := x"FAE6";
          m(425) := x"FBE4";
          m(426) := x"F8DA";
          m(427) := x"F75D";
          m(428) := x"FF25";
          m(429) := x"FF42";
          m(430) := x"F81D";
          m(431) := x"00AA";
          m(432) := x"05E3";
          m(433) := x"06CE";
          m(434) := x"0BD8";
          m(435) := x"0725";
          m(436) := x"FF6A";
          m(437) := x"022C";
          m(438) := x"00DC";
          m(439) := x"026C";
          m(440) := x"005F";
          m(441) := x"FB5E";
          m(442) := x"FE5C";
          m(443) := x"004B";
          m(444) := x"03E4";
          m(445) := x"0222";
          m(446) := x"0290";
          m(447) := x"003D";
          m(448) := x"FFFD";
          m(449) := x"FFC0";
          m(450) := x"0068";
          m(451) := x"001F";
          m(452) := x"FEC8";
          m(453) := x"FA9B";
          m(454) := x"FD72";
          m(455) := x"FCAD";
          m(456) := x"FB14";
          m(457) := x"015C";
          m(458) := x"0165";
          m(459) := x"0196";
          m(460) := x"0631";
          m(461) := x"05AF";
          m(462) := x"07FB";
          m(463) := x"07C9";
          m(464) := x"049E";
          m(465) := x"0053";
          m(466) := x"026C";
          m(467) := x"03EC";
          m(468) := x"FD02";
          m(469) := x"0138";
          m(470) := x"FECE";
          m(471) := x"027C";
          m(472) := x"02BF";
          m(473) := x"025F";
          m(474) := x"013D";
          m(475) := x"001C";
          m(476) := x"FFFB";
          m(477) := x"0021";
          m(478) := x"0023";
          m(479) := x"0105";
          m(480) := x"01B1";
          m(481) := x"FF6C";
          m(482) := x"FE6A";
          m(483) := x"FD69";
          m(484) := x"FE67";
          m(485) := x"0101";
          m(486) := x"00EA";
          m(487) := x"0063";
          m(488) := x"027A";
          m(489) := x"0685";
          m(490) := x"0A29";
          m(491) := x"0B59";
          m(492) := x"0186";
          m(493) := x"FF00";
          m(494) := x"FDE2";
          m(495) := x"00FB";
          m(496) := x"FEAD";
          m(497) := x"04A6";
          m(498) := x"0006";
          m(499) := x"FE73";
          m(500) := x"007B";
          m(501) := x"0142";
          m(502) := x"0063";
          m(503) := x"FFE0";
          m(504) := x"FFFA";
          m(505) := x"FFE7";
          m(506) := x"001E";
          m(507) := x"0085";
          m(508) := x"0301";
          m(509) := x"04C1";
          m(510) := x"FF62";
          m(511) := x"FFA0";
          m(512) := x"0406";
          m(513) := x"FFBE";
          m(514) := x"03F8";
          m(515) := x"FC78";
          m(516) := x"FD78";
          m(517) := x"032F";
          m(518) := x"0AA3";
          m(519) := x"09BE";
          m(520) := x"FD63";
          m(521) := x"F90F";
          m(522) := x"FF40";
          m(523) := x"FD5E";
          m(524) := x"FC1E";
          m(525) := x"00CC";
          m(526) := x"FEF8";
          m(527) := x"0342";
          m(528) := x"FF87";
          m(529) := x"013D";
          m(530) := x"0012";
          m(531) := x"0040";
          m(532) := x"0006";
          m(533) := x"0004";
          m(534) := x"FDEC";
          m(535) := x"FE63";
          m(536) := x"0330";
          m(537) := x"0450";
          m(538) := x"0184";
          m(539) := x"FFFE";
          m(540) := x"FF17";
          m(541) := x"0052";
          m(542) := x"FDD1";
          m(543) := x"F6F5";
          m(544) := x"FACF";
          m(545) := x"05A4";
          m(546) := x"0B0C";
          m(547) := x"0925";
          m(548) := x"FAB8";
          m(549) := x"FD9B";
          m(550) := x"FD71";
          m(551) := x"FCEB";
          m(552) := x"FE62";
          m(553) := x"FE45";
          m(554) := x"FDF2";
          m(555) := x"0285";
          m(556) := x"007C";
          m(557) := x"00D6";
          m(558) := x"0047";
          m(559) := x"001A";
          m(560) := x"FFDB";
          m(561) := x"003E";
          m(562) := x"FEF4";
          m(563) := x"FF9C";
          m(564) := x"01C8";
          m(565) := x"00F8";
          m(566) := x"FF57";
          m(567) := x"08E5";
          m(568) := x"00A3";
          m(569) := x"FF95";
          m(570) := x"005B";
          m(571) := x"FF25";
          m(572) := x"04C8";
          m(573) := x"08CA";
          m(574) := x"0352";
          m(575) := x"FF66";
          m(576) := x"F3ED";
          m(577) := x"FF8E";
          m(578) := x"FF09";
          m(579) := x"FF67";
          m(580) := x"038D";
          m(581) := x"0506";
          m(582) := x"FF80";
          m(583) := x"0264";
          m(584) := x"009A";
          m(585) := x"FEDA";
          m(586) := x"0037";
          m(587) := x"001C";
          m(588) := x"0000";
          m(589) := x"001F";
          m(590) := x"017C";
          m(591) := x"02B7";
          m(592) := x"01FF";
          m(593) := x"FD57";
          m(594) := x"FFFB";
          m(595) := x"00D6";
          m(596) := x"FB54";
          m(597) := x"FD54";
          m(598) := x"FEC8";
          m(599) := x"038C";
          m(600) := x"01A7";
          m(601) := x"06AF";
          m(602) := x"04D5";
          m(603) := x"FAEC";
          m(604) := x"F931";
          m(605) := x"00A8";
          m(606) := x"FC04";
          m(607) := x"FE9E";
          m(608) := x"FF16";
          m(609) := x"FE7A";
          m(610) := x"FEEE";
          m(611) := x"014A";
          m(612) := x"FE87";
          m(613) := x"FFFA";
          m(614) := x"000D";
          m(615) := x"0021";
          m(616) := x"FFB5";
          m(617) := x"FFDE";
          m(618) := x"01AC";
          m(619) := x"0215";
          m(620) := x"0257";
          m(621) := x"FE7B";
          m(622) := x"02FC";
          m(623) := x"039F";
          m(624) := x"011F";
          m(625) := x"04CD";
          m(626) := x"0512";
          m(627) := x"04B6";
          m(628) := x"064A";
          m(629) := x"049C";
          m(630) := x"FA4E";
          m(631) := x"FE30";
          m(632) := x"FCB1";
          m(633) := x"FF3F";
          m(634) := x"F967";
          m(635) := x"FDCA";
          m(636) := x"02AB";
          m(637) := x"FB7D";
          m(638) := x"FE2E";
          m(639) := x"FFE2";
          m(640) := x"016F";
          m(641) := x"006B";
          m(642) := x"FFE7";
          m(643) := x"FFFE";
          m(644) := x"0014";
          m(645) := x"0018";
          m(646) := x"0028";
          m(647) := x"FFE3";
          m(648) := x"00C3";
          m(649) := x"FEAD";
          m(650) := x"FD5A";
          m(651) := x"FE7A";
          m(652) := x"00A3";
          m(653) := x"0432";
          m(654) := x"06F8";
          m(655) := x"03FE";
          m(656) := x"0572";
          m(657) := x"05A7";
          m(658) := x"FB48";
          m(659) := x"F9F6";
          m(660) := x"F9C1";
          m(661) := x"F7E0";
          m(662) := x"00A5";
          m(663) := x"0356";
          m(664) := x"0113";
          m(665) := x"FE59";
          m(666) := x"FEAA";
          m(667) := x"00F2";
          m(668) := x"0072";
          m(669) := x"0076";
          m(670) := x"0025";
          m(671) := x"0015";
          m(672) := x"003A";
          m(673) := x"0035";
          m(674) := x"FFE0";
          m(675) := x"FFCB";
          m(676) := x"001E";
          m(677) := x"FF68";
          m(678) := x"FDC2";
          m(679) := x"FC70";
          m(680) := x"FD7D";
          m(681) := x"FEA0";
          m(682) := x"FDE5";
          m(683) := x"FFBA";
          m(684) := x"023F";
          m(685) := x"06C5";
          m(686) := x"00C3";
          m(687) := x"F910";
          m(688) := x"FA82";
          m(689) := x"F8A8";
          m(690) := x"FCD9";
          m(691) := x"FF81";
          m(692) := x"FA53";
          m(693) := x"FC59";
          m(694) := x"FDF9";
          m(695) := x"FE79";
          m(696) := x"00E8";
          m(697) := x"0091";
          m(698) := x"0048";
          m(699) := x"001B";
          m(700) := x"000E";
          m(701) := x"FFF5";
          m(702) := x"0024";
          m(703) := x"FFF6";
          m(704) := x"FF9B";
          m(705) := x"FFCD";
          m(706) := x"FFD6";
          m(707) := x"0100";
          m(708) := x"0143";
          m(709) := x"00B7";
          m(710) := x"0461";
          m(711) := x"0306";
          m(712) := x"06F0";
          m(713) := x"03E5";
          m(714) := x"FE20";
          m(715) := x"000E";
          m(716) := x"FFE7";
          m(717) := x"FCAE";
          m(718) := x"FC49";
          m(719) := x"FD5F";
          m(720) := x"FD06";
          m(721) := x"FE1B";
          m(722) := x"0043";
          m(723) := x"005F";
          m(724) := x"000D";
          m(725) := x"0006";
          m(726) := x"FFF2";
          m(727) := x"0017";
          m(728) := x"0005";
          m(729) := x"000B";
          m(730) := x"0002";
          m(731) := x"FFF6";
          m(732) := x"FFB6";
          m(733) := x"FFD5";
          m(734) := x"FFF4";
          m(735) := x"FFF3";
          m(736) := x"FFF8";
          m(737) := x"FF29";
          m(738) := x"FF2F";
          m(739) := x"003A";
          m(740) := x"0039";
          m(741) := x"0046";
          m(742) := x"FBCF";
          m(743) := x"FB26";
          m(744) := x"FC7B";
          m(745) := x"FCA9";
          m(746) := x"FDF3";
          m(747) := x"FE39";
          m(748) := x"FD59";
          m(749) := x"FD8E";
          m(750) := x"FF42";
          m(751) := x"FFD3";
          m(752) := x"0020";
          m(753) := x"0018";
          m(754) := x"0012";
          m(755) := x"0037";
          m(756) := x"0004";
          m(757) := x"0016";
          m(758) := x"0000";
          m(759) := x"FFF0";
          m(760) := x"FFE0";
          m(761) := x"FFC2";
          m(762) := x"000E";
          m(763) := x"0006";
          m(764) := x"FFFD";
          m(765) := x"003E";
          m(766) := x"FFE1";
          m(767) := x"0006";
          m(768) := x"FFDB";
          m(769) := x"001D";
          m(770) := x"FEFE";
          m(771) := x"FF6C";
          m(772) := x"FFBB";
          m(773) := x"FFFE";
          m(774) := x"FF7E";
          m(775) := x"001D";
          m(776) := x"FFA2";
          m(777) := x"FF94";
          m(778) := x"FF8E";
          m(779) := x"0020";
          m(780) := x"0031";
          m(781) := x"FFFE";
          m(782) := x"FFFD";
          m(783) := x"FFF9";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_9.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 9) then
          m(0) := x"FFA7";
          m(1) := x"FFBF";
          m(2) := x"FFFA";
          m(3) := x"FFF2";
          m(4) := x"FFE7";
          m(5) := x"0038";
          m(6) := x"FFC4";
          m(7) := x"FFFF";
          m(8) := x"FFF8";
          m(9) := x"0006";
          m(10) := x"FFDB";
          m(11) := x"0002";
          m(12) := x"FFF6";
          m(13) := x"003C";
          m(14) := x"0026";
          m(15) := x"FFF9";
          m(16) := x"0029";
          m(17) := x"FFF6";
          m(18) := x"0021";
          m(19) := x"FFF6";
          m(20) := x"0001";
          m(21) := x"0000";
          m(22) := x"000F";
          m(23) := x"FFE3";
          m(24) := x"002B";
          m(25) := x"0013";
          m(26) := x"FFD6";
          m(27) := x"000F";
          m(28) := x"000B";
          m(29) := x"FFDC";
          m(30) := x"FFFD";
          m(31) := x"0017";
          m(32) := x"000F";
          m(33) := x"000D";
          m(34) := x"FFC9";
          m(35) := x"0003";
          m(36) := x"FFFB";
          m(37) := x"FFD4";
          m(38) := x"0008";
          m(39) := x"FFF8";
          m(40) := x"FFDF";
          m(41) := x"FFDF";
          m(42) := x"003A";
          m(43) := x"0065";
          m(44) := x"0009";
          m(45) := x"0046";
          m(46) := x"0035";
          m(47) := x"FFF9";
          m(48) := x"FFCA";
          m(49) := x"0013";
          m(50) := x"0017";
          m(51) := x"0018";
          m(52) := x"FFF6";
          m(53) := x"FFE0";
          m(54) := x"0021";
          m(55) := x"0024";
          m(56) := x"FFF9";
          m(57) := x"0007";
          m(58) := x"0033";
          m(59) := x"0000";
          m(60) := x"002F";
          m(61) := x"FFF2";
          m(62) := x"FFF3";
          m(63) := x"0003";
          m(64) := x"004E";
          m(65) := x"0032";
          m(66) := x"FFAF";
          m(67) := x"FF46";
          m(68) := x"0034";
          m(69) := x"02C5";
          m(70) := x"0227";
          m(71) := x"0218";
          m(72) := x"00DD";
          m(73) := x"FFD5";
          m(74) := x"FFF2";
          m(75) := x"0028";
          m(76) := x"FF9F";
          m(77) := x"FFFE";
          m(78) := x"FFC6";
          m(79) := x"FFD8";
          m(80) := x"FFF5";
          m(81) := x"FFF2";
          m(82) := x"003B";
          m(83) := x"0039";
          m(84) := x"FFDD";
          m(85) := x"0033";
          m(86) := x"0007";
          m(87) := x"FFF6";
          m(88) := x"FFE1";
          m(89) := x"FF4E";
          m(90) := x"FF3E";
          m(91) := x"FECB";
          m(92) := x"FC84";
          m(93) := x"FD2B";
          m(94) := x"FC77";
          m(95) := x"FB5E";
          m(96) := x"FD74";
          m(97) := x"FF84";
          m(98) := x"FCC6";
          m(99) := x"FFE2";
          m(100) := x"0175";
          m(101) := x"FF8F";
          m(102) := x"FBD7";
          m(103) := x"FE15";
          m(104) := x"FC1E";
          m(105) := x"FBF9";
          m(106) := x"FD96";
          m(107) := x"FF76";
          m(108) := x"FFE1";
          m(109) := x"0032";
          m(110) := x"FFD8";
          m(111) := x"FFF4";
          m(112) := x"FFE7";
          m(113) := x"0006";
          m(114) := x"0001";
          m(115) := x"0011";
          m(116) := x"000D";
          m(117) := x"FF1F";
          m(118) := x"FE7A";
          m(119) := x"FD51";
          m(120) := x"FE64";
          m(121) := x"FFC3";
          m(122) := x"0107";
          m(123) := x"FB44";
          m(124) := x"FC26";
          m(125) := x"00B8";
          m(126) := x"FF7E";
          m(127) := x"016B";
          m(128) := x"0063";
          m(129) := x"FFB9";
          m(130) := x"FE6A";
          m(131) := x"FC8F";
          m(132) := x"FD96";
          m(133) := x"FD93";
          m(134) := x"FFD7";
          m(135) := x"FEAC";
          m(136) := x"FD0A";
          m(137) := x"FEDF";
          m(138) := x"FFE2";
          m(139) := x"FFE4";
          m(140) := x"FFF3";
          m(141) := x"FFE5";
          m(142) := x"003E";
          m(143) := x"FF8D";
          m(144) := x"FF50";
          m(145) := x"FEF9";
          m(146) := x"FE83";
          m(147) := x"FCF8";
          m(148) := x"FC76";
          m(149) := x"FFB7";
          m(150) := x"FF8E";
          m(151) := x"00D0";
          m(152) := x"0184";
          m(153) := x"0162";
          m(154) := x"FBC2";
          m(155) := x"004C";
          m(156) := x"FEF0";
          m(157) := x"FAE5";
          m(158) := x"FF69";
          m(159) := x"FEC1";
          m(160) := x"FAAD";
          m(161) := x"004D";
          m(162) := x"02A9";
          m(163) := x"011F";
          m(164) := x"FEB9";
          m(165) := x"FF06";
          m(166) := x"FFDA";
          m(167) := x"0030";
          m(168) := x"0043";
          m(169) := x"FFDC";
          m(170) := x"FF08";
          m(171) := x"FE7B";
          m(172) := x"FDB8";
          m(173) := x"FB33";
          m(174) := x"FE04";
          m(175) := x"FF51";
          m(176) := x"FD01";
          m(177) := x"01AC";
          m(178) := x"02D5";
          m(179) := x"FF6E";
          m(180) := x"0284";
          m(181) := x"00C1";
          m(182) := x"0219";
          m(183) := x"FBA5";
          m(184) := x"FE73";
          m(185) := x"FDE8";
          m(186) := x"009E";
          m(187) := x"FF8A";
          m(188) := x"FF65";
          m(189) := x"FE9B";
          m(190) := x"0131";
          m(191) := x"008E";
          m(192) := x"FF39";
          m(193) := x"FF5A";
          m(194) := x"0057";
          m(195) := x"0090";
          m(196) := x"FFF5";
          m(197) := x"FFE1";
          m(198) := x"FFAB";
          m(199) := x"FF28";
          m(200) := x"FEF2";
          m(201) := x"FCD3";
          m(202) := x"FC1A";
          m(203) := x"FE87";
          m(204) := x"FF8A";
          m(205) := x"FF94";
          m(206) := x"FF80";
          m(207) := x"FF5C";
          m(208) := x"FF5B";
          m(209) := x"FDF9";
          m(210) := x"01D2";
          m(211) := x"FE55";
          m(212) := x"FF58";
          m(213) := x"FD53";
          m(214) := x"032C";
          m(215) := x"0378";
          m(216) := x"0181";
          m(217) := x"04FF";
          m(218) := x"0217";
          m(219) := x"FF62";
          m(220) := x"FCDF";
          m(221) := x"FDA9";
          m(222) := x"0068";
          m(223) := x"004D";
          m(224) := x"FFC8";
          m(225) := x"FFDA";
          m(226) := x"FFD2";
          m(227) := x"FF4E";
          m(228) := x"FFF9";
          m(229) := x"FF34";
          m(230) := x"FF90";
          m(231) := x"0166";
          m(232) := x"005C";
          m(233) := x"00A8";
          m(234) := x"04AD";
          m(235) := x"045D";
          m(236) := x"04B7";
          m(237) := x"FFFF";
          m(238) := x"0458";
          m(239) := x"FF2F";
          m(240) := x"FA8C";
          m(241) := x"048F";
          m(242) := x"01D5";
          m(243) := x"03D4";
          m(244) := x"FEFF";
          m(245) := x"00B7";
          m(246) := x"FFD1";
          m(247) := x"0176";
          m(248) := x"FC5A";
          m(249) := x"FE45";
          m(250) := x"FFAB";
          m(251) := x"FFD1";
          m(252) := x"0020";
          m(253) := x"0023";
          m(254) := x"0038";
          m(255) := x"FE94";
          m(256) := x"FF3D";
          m(257) := x"FE72";
          m(258) := x"FF48";
          m(259) := x"016D";
          m(260) := x"FF0E";
          m(261) := x"0065";
          m(262) := x"FFAF";
          m(263) := x"02D3";
          m(264) := x"04E9";
          m(265) := x"05E0";
          m(266) := x"0209";
          m(267) := x"033A";
          m(268) := x"0444";
          m(269) := x"FE2B";
          m(270) := x"008F";
          m(271) := x"FF2C";
          m(272) := x"F9C9";
          m(273) := x"FE56";
          m(274) := x"0003";
          m(275) := x"00F9";
          m(276) := x"FE68";
          m(277) := x"FF5A";
          m(278) := x"0054";
          m(279) := x"007C";
          m(280) := x"FFF9";
          m(281) := x"FFC5";
          m(282) := x"005E";
          m(283) := x"FF17";
          m(284) := x"FE93";
          m(285) := x"FCC1";
          m(286) := x"FD5C";
          m(287) := x"FE00";
          m(288) := x"FFC5";
          m(289) := x"FE99";
          m(290) := x"FA12";
          m(291) := x"0069";
          m(292) := x"04D3";
          m(293) := x"0538";
          m(294) := x"0734";
          m(295) := x"0AD8";
          m(296) := x"023F";
          m(297) := x"04F1";
          m(298) := x"FBD9";
          m(299) := x"FC9D";
          m(300) := x"F89E";
          m(301) := x"02DA";
          m(302) := x"0000";
          m(303) := x"FF5E";
          m(304) := x"FEAC";
          m(305) := x"FF45";
          m(306) := x"0025";
          m(307) := x"006B";
          m(308) := x"FFE6";
          m(309) := x"FFFB";
          m(310) := x"FFBC";
          m(311) := x"FFAD";
          m(312) := x"FE9D";
          m(313) := x"FD77";
          m(314) := x"FD37";
          m(315) := x"FC97";
          m(316) := x"FA97";
          m(317) := x"FE3E";
          m(318) := x"FFCB";
          m(319) := x"00CE";
          m(320) := x"044B";
          m(321) := x"0627";
          m(322) := x"07A5";
          m(323) := x"0208";
          m(324) := x"0750";
          m(325) := x"FCEE";
          m(326) := x"FA9C";
          m(327) := x"F913";
          m(328) := x"FFC8";
          m(329) := x"04DD";
          m(330) := x"006B";
          m(331) := x"FD45";
          m(332) := x"FBBA";
          m(333) := x"FEC5";
          m(334) := x"FF13";
          m(335) := x"FFF1";
          m(336) := x"FFFC";
          m(337) := x"FFDC";
          m(338) := x"0035";
          m(339) := x"FFDD";
          m(340) := x"FF69";
          m(341) := x"FF2E";
          m(342) := x"FF2E";
          m(343) := x"FF07";
          m(344) := x"002C";
          m(345) := x"009A";
          m(346) := x"FB0A";
          m(347) := x"FEAD";
          m(348) := x"02FA";
          m(349) := x"01FF";
          m(350) := x"0251";
          m(351) := x"FD31";
          m(352) := x"0212";
          m(353) := x"FEE1";
          m(354) := x"F85A";
          m(355) := x"FA90";
          m(356) := x"FE7F";
          m(357) := x"02BC";
          m(358) := x"FEA3";
          m(359) := x"FD4D";
          m(360) := x"FFFB";
          m(361) := x"00B2";
          m(362) := x"FF3E";
          m(363) := x"0014";
          m(364) := x"0011";
          m(365) := x"0004";
          m(366) := x"0000";
          m(367) := x"000F";
          m(368) := x"FF04";
          m(369) := x"FE98";
          m(370) := x"FE7B";
          m(371) := x"FD1E";
          m(372) := x"FFC0";
          m(373) := x"FE6B";
          m(374) := x"F733";
          m(375) := x"F96A";
          m(376) := x"FBFB";
          m(377) := x"FFF6";
          m(378) := x"FDFE";
          m(379) := x"010B";
          m(380) := x"0587";
          m(381) := x"0292";
          m(382) := x"FD57";
          m(383) := x"FA76";
          m(384) := x"FD69";
          m(385) := x"FF62";
          m(386) := x"FC2E";
          m(387) := x"FCF7";
          m(388) := x"FFC4";
          m(389) := x"00E2";
          m(390) := x"0002";
          m(391) := x"FFEB";
          m(392) := x"001B";
          m(393) := x"0010";
          m(394) := x"0035";
          m(395) := x"0023";
          m(396) := x"FF25";
          m(397) := x"FE44";
          m(398) := x"FBB9";
          m(399) := x"FAC9";
          m(400) := x"FC28";
          m(401) := x"FD30";
          m(402) := x"FBCF";
          m(403) := x"F783";
          m(404) := x"FFB7";
          m(405) := x"FAA7";
          m(406) := x"0089";
          m(407) := x"003F";
          m(408) := x"0193";
          m(409) := x"FFCF";
          m(410) := x"FE98";
          m(411) := x"FB36";
          m(412) := x"F983";
          m(413) := x"F9AB";
          m(414) := x"F9FB";
          m(415) := x"FBFE";
          m(416) := x"FECC";
          m(417) := x"0112";
          m(418) := x"0101";
          m(419) := x"FFD9";
          m(420) := x"FFF8";
          m(421) := x"FFD5";
          m(422) := x"FFDC";
          m(423) := x"FFFD";
          m(424) := x"FEDA";
          m(425) := x"FBA7";
          m(426) := x"F868";
          m(427) := x"F8E3";
          m(428) := x"FB9D";
          m(429) := x"FA93";
          m(430) := x"FB9B";
          m(431) := x"FCA3";
          m(432) := x"FDEA";
          m(433) := x"0375";
          m(434) := x"04B6";
          m(435) := x"FFC1";
          m(436) := x"0080";
          m(437) := x"FAB7";
          m(438) := x"F1B4";
          m(439) := x"EF13";
          m(440) := x"F126";
          m(441) := x"F54B";
          m(442) := x"F6FF";
          m(443) := x"F8FD";
          m(444) := x"FD0B";
          m(445) := x"0124";
          m(446) := x"0142";
          m(447) := x"0001";
          m(448) := x"FFF9";
          m(449) := x"FFCF";
          m(450) := x"FFFC";
          m(451) := x"FFCE";
          m(452) := x"FEA1";
          m(453) := x"FC4E";
          m(454) := x"FA69";
          m(455) := x"F87A";
          m(456) := x"FA51";
          m(457) := x"02C9";
          m(458) := x"0160";
          m(459) := x"FEEC";
          m(460) := x"FD0B";
          m(461) := x"004D";
          m(462) := x"072A";
          m(463) := x"FE06";
          m(464) := x"FC8C";
          m(465) := x"F192";
          m(466) := x"EA53";
          m(467) := x"EDAB";
          m(468) := x"F193";
          m(469) := x"F4C0";
          m(470) := x"F846";
          m(471) := x"FB39";
          m(472) := x"FFB7";
          m(473) := x"01DB";
          m(474) := x"00EB";
          m(475) := x"0029";
          m(476) := x"0004";
          m(477) := x"FFF6";
          m(478) := x"0009";
          m(479) := x"FFED";
          m(480) := x"FF02";
          m(481) := x"FDE9";
          m(482) := x"FAA5";
          m(483) := x"F564";
          m(484) := x"FA0A";
          m(485) := x"FC63";
          m(486) := x"0008";
          m(487) := x"04C6";
          m(488) := x"0515";
          m(489) := x"FFEC";
          m(490) := x"02E3";
          m(491) := x"FB40";
          m(492) := x"F70D";
          m(493) := x"EAA0";
          m(494) := x"F1A9";
          m(495) := x"F90C";
          m(496) := x"F98D";
          m(497) := x"F8F1";
          m(498) := x"FB7D";
          m(499) := x"FCEB";
          m(500) := x"0230";
          m(501) := x"0342";
          m(502) := x"00D3";
          m(503) := x"FFEE";
          m(504) := x"FFE4";
          m(505) := x"FFD9";
          m(506) := x"001C";
          m(507) := x"FF9A";
          m(508) := x"FF1A";
          m(509) := x"FB7E";
          m(510) := x"F6D8";
          m(511) := x"FB51";
          m(512) := x"01E8";
          m(513) := x"02C3";
          m(514) := x"0224";
          m(515) := x"FC9A";
          m(516) := x"FD23";
          m(517) := x"FE23";
          m(518) := x"FCC9";
          m(519) := x"FC1C";
          m(520) := x"F5E1";
          m(521) := x"FA37";
          m(522) := x"0228";
          m(523) := x"0199";
          m(524) := x"0237";
          m(525) := x"FFA6";
          m(526) := x"0071";
          m(527) := x"0149";
          m(528) := x"03C1";
          m(529) := x"029A";
          m(530) := x"0093";
          m(531) := x"00D7";
          m(532) := x"000C";
          m(533) := x"FFDD";
          m(534) := x"FFAA";
          m(535) := x"FFBA";
          m(536) := x"FF75";
          m(537) := x"F796";
          m(538) := x"FAD0";
          m(539) := x"0194";
          m(540) := x"0276";
          m(541) := x"080B";
          m(542) := x"03F2";
          m(543) := x"04FB";
          m(544) := x"01F0";
          m(545) := x"055A";
          m(546) := x"FC25";
          m(547) := x"FFF9";
          m(548) := x"FFDA";
          m(549) := x"FEDC";
          m(550) := x"FFB0";
          m(551) := x"FF25";
          m(552) := x"03C3";
          m(553) := x"FF1C";
          m(554) := x"FF94";
          m(555) := x"0192";
          m(556) := x"0105";
          m(557) := x"0359";
          m(558) := x"004D";
          m(559) := x"0031";
          m(560) := x"004D";
          m(561) := x"FFE2";
          m(562) := x"FFE2";
          m(563) := x"011F";
          m(564) := x"0175";
          m(565) := x"FAB1";
          m(566) := x"0121";
          m(567) := x"FF1F";
          m(568) := x"05A9";
          m(569) := x"03C2";
          m(570) := x"037A";
          m(571) := x"070A";
          m(572) := x"089B";
          m(573) := x"FE4E";
          m(574) := x"0156";
          m(575) := x"0070";
          m(576) := x"0283";
          m(577) := x"0469";
          m(578) := x"025E";
          m(579) := x"FF44";
          m(580) := x"0201";
          m(581) := x"FEC7";
          m(582) := x"FF19";
          m(583) := x"02BD";
          m(584) := x"035C";
          m(585) := x"0305";
          m(586) := x"FFFF";
          m(587) := x"FFC2";
          m(588) := x"FFFD";
          m(589) := x"FFDD";
          m(590) := x"0023";
          m(591) := x"0298";
          m(592) := x"00DC";
          m(593) := x"057F";
          m(594) := x"0266";
          m(595) := x"FF97";
          m(596) := x"0158";
          m(597) := x"0155";
          m(598) := x"010F";
          m(599) := x"FD87";
          m(600) := x"FFEF";
          m(601) := x"FE78";
          m(602) := x"01C8";
          m(603) := x"019C";
          m(604) := x"FD9E";
          m(605) := x"FE81";
          m(606) := x"04A5";
          m(607) := x"02F9";
          m(608) := x"0343";
          m(609) := x"01B4";
          m(610) := x"FFE7";
          m(611) := x"02F8";
          m(612) := x"02E4";
          m(613) := x"01C2";
          m(614) := x"009B";
          m(615) := x"FFED";
          m(616) := x"FFF0";
          m(617) := x"FFEA";
          m(618) := x"000F";
          m(619) := x"0064";
          m(620) := x"01E5";
          m(621) := x"07B9";
          m(622) := x"02AD";
          m(623) := x"01BC";
          m(624) := x"030E";
          m(625) := x"04F6";
          m(626) := x"FD38";
          m(627) := x"FD3A";
          m(628) := x"F90D";
          m(629) := x"FBC7";
          m(630) := x"0397";
          m(631) := x"004F";
          m(632) := x"00BA";
          m(633) := x"01A1";
          m(634) := x"08DE";
          m(635) := x"029E";
          m(636) := x"05AE";
          m(637) := x"03EF";
          m(638) := x"FEC6";
          m(639) := x"0098";
          m(640) := x"011B";
          m(641) := x"0093";
          m(642) := x"FFF6";
          m(643) := x"0023";
          m(644) := x"0021";
          m(645) := x"001F";
          m(646) := x"0015";
          m(647) := x"FE30";
          m(648) := x"FD30";
          m(649) := x"020B";
          m(650) := x"02BD";
          m(651) := x"01B1";
          m(652) := x"FCB3";
          m(653) := x"00F3";
          m(654) := x"FC28";
          m(655) := x"FF2A";
          m(656) := x"0B2A";
          m(657) := x"02D0";
          m(658) := x"000D";
          m(659) := x"01E0";
          m(660) := x"02FC";
          m(661) := x"04B8";
          m(662) := x"0128";
          m(663) := x"01C4";
          m(664) := x"0030";
          m(665) := x"FF2A";
          m(666) := x"00BD";
          m(667) := x"0043";
          m(668) := x"0084";
          m(669) := x"006D";
          m(670) := x"0020";
          m(671) := x"FFFA";
          m(672) := x"002A";
          m(673) := x"0014";
          m(674) := x"0000";
          m(675) := x"FF10";
          m(676) := x"FF98";
          m(677) := x"00AE";
          m(678) := x"0097";
          m(679) := x"FC70";
          m(680) := x"FCC8";
          m(681) := x"FC24";
          m(682) := x"FA41";
          m(683) := x"FF34";
          m(684) := x"FFFF";
          m(685) := x"FDE4";
          m(686) := x"FF76";
          m(687) := x"FC90";
          m(688) := x"F82D";
          m(689) := x"00C1";
          m(690) := x"0322";
          m(691) := x"0460";
          m(692) := x"FF72";
          m(693) := x"024C";
          m(694) := x"0172";
          m(695) := x"009C";
          m(696) := x"006C";
          m(697) := x"004A";
          m(698) := x"002A";
          m(699) := x"FFDA";
          m(700) := x"0045";
          m(701) := x"FFE6";
          m(702) := x"FFF8";
          m(703) := x"0008";
          m(704) := x"0097";
          m(705) := x"FE8E";
          m(706) := x"FD90";
          m(707) := x"FD67";
          m(708) := x"FF64";
          m(709) := x"FE96";
          m(710) := x"FC39";
          m(711) := x"0029";
          m(712) := x"FFDB";
          m(713) := x"FEF7";
          m(714) := x"FF38";
          m(715) := x"FB53";
          m(716) := x"FC52";
          m(717) := x"003C";
          m(718) := x"FE89";
          m(719) := x"FBA1";
          m(720) := x"FE2E";
          m(721) := x"FFD4";
          m(722) := x"FFFA";
          m(723) := x"00A8";
          m(724) := x"0010";
          m(725) := x"004A";
          m(726) := x"FFE7";
          m(727) := x"0010";
          m(728) := x"0006";
          m(729) := x"FFD7";
          m(730) := x"FFEF";
          m(731) := x"FFFC";
          m(732) := x"FF84";
          m(733) := x"FF8C";
          m(734) := x"FF0B";
          m(735) := x"FE82";
          m(736) := x"FF63";
          m(737) := x"FF4F";
          m(738) := x"FE88";
          m(739) := x"FE97";
          m(740) := x"FC0B";
          m(741) := x"FBCF";
          m(742) := x"FC0D";
          m(743) := x"FB51";
          m(744) := x"FB96";
          m(745) := x"FC47";
          m(746) := x"FE07";
          m(747) := x"FE58";
          m(748) := x"FEDB";
          m(749) := x"FF21";
          m(750) := x"FFF6";
          m(751) := x"000F";
          m(752) := x"FFF2";
          m(753) := x"FFFC";
          m(754) := x"000D";
          m(755) := x"0019";
          m(756) := x"FFC3";
          m(757) := x"0025";
          m(758) := x"000C";
          m(759) := x"001B";
          m(760) := x"0003";
          m(761) := x"0028";
          m(762) := x"FFFE";
          m(763) := x"000F";
          m(764) := x"FFF5";
          m(765) := x"FFDC";
          m(766) := x"FFE6";
          m(767) := x"0000";
          m(768) := x"FFBE";
          m(769) := x"FFE0";
          m(770) := x"FFE7";
          m(771) := x"FFE7";
          m(772) := x"FFB4";
          m(773) := x"FFAF";
          m(774) := x"FF5A";
          m(775) := x"000C";
          m(776) := x"FFCF";
          m(777) := x"0024";
          m(778) := x"FFFF";
          m(779) := x"FFF4";
          m(780) := x"FFE9";
          m(781) := x"FFDA";
          m(782) := x"FFE2";
          m(783) := x"0024";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_10.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 10) then
          m(0) := x"FFC9";
          m(1) := x"0008";
          m(2) := x"000C";
          m(3) := x"FFE3";
          m(4) := x"FFDE";
          m(5) := x"001C";
          m(6) := x"0000";
          m(7) := x"000B";
          m(8) := x"FFD3";
          m(9) := x"FFE6";
          m(10) := x"FFE2";
          m(11) := x"0026";
          m(12) := x"FFC6";
          m(13) := x"FFED";
          m(14) := x"0013";
          m(15) := x"FFD9";
          m(16) := x"FFF3";
          m(17) := x"FFE9";
          m(18) := x"000F";
          m(19) := x"FFD5";
          m(20) := x"0037";
          m(21) := x"FFEC";
          m(22) := x"0005";
          m(23) := x"FFDB";
          m(24) := x"FFBE";
          m(25) := x"0031";
          m(26) := x"FFF8";
          m(27) := x"0016";
          m(28) := x"0004";
          m(29) := x"FFE6";
          m(30) := x"FFFA";
          m(31) := x"000F";
          m(32) := x"0026";
          m(33) := x"FFDD";
          m(34) := x"000E";
          m(35) := x"FFD7";
          m(36) := x"FFF9";
          m(37) := x"000A";
          m(38) := x"FFEF";
          m(39) := x"FFEB";
          m(40) := x"FF55";
          m(41) := x"FF7D";
          m(42) := x"0043";
          m(43) := x"005D";
          m(44) := x"00E3";
          m(45) := x"002F";
          m(46) := x"0015";
          m(47) := x"FFF0";
          m(48) := x"FFA3";
          m(49) := x"FFBB";
          m(50) := x"0038";
          m(51) := x"002E";
          m(52) := x"FFEB";
          m(53) := x"0002";
          m(54) := x"FFB9";
          m(55) := x"FFF7";
          m(56) := x"FFFA";
          m(57) := x"001E";
          m(58) := x"000D";
          m(59) := x"002C";
          m(60) := x"0033";
          m(61) := x"0011";
          m(62) := x"001D";
          m(63) := x"FFA2";
          m(64) := x"003E";
          m(65) := x"005C";
          m(66) := x"FFB9";
          m(67) := x"FF4A";
          m(68) := x"0054";
          m(69) := x"019B";
          m(70) := x"0213";
          m(71) := x"01E1";
          m(72) := x"01AB";
          m(73) := x"FDD0";
          m(74) := x"FD70";
          m(75) := x"FEDE";
          m(76) := x"FFA4";
          m(77) := x"FED1";
          m(78) := x"FFAC";
          m(79) := x"FFA4";
          m(80) := x"FFF4";
          m(81) := x"FFF2";
          m(82) := x"0006";
          m(83) := x"0002";
          m(84) := x"000E";
          m(85) := x"0040";
          m(86) := x"0046";
          m(87) := x"FFCF";
          m(88) := x"0019";
          m(89) := x"FFC8";
          m(90) := x"FFDD";
          m(91) := x"FFD5";
          m(92) := x"003E";
          m(93) := x"FFE2";
          m(94) := x"0118";
          m(95) := x"01B5";
          m(96) := x"0530";
          m(97) := x"044C";
          m(98) := x"0063";
          m(99) := x"FF61";
          m(100) := x"04BA";
          m(101) := x"072E";
          m(102) := x"0121";
          m(103) := x"FEFA";
          m(104) := x"FFD2";
          m(105) := x"FC7A";
          m(106) := x"FC85";
          m(107) := x"FD16";
          m(108) := x"FDE5";
          m(109) := x"0014";
          m(110) := x"0027";
          m(111) := x"0002";
          m(112) := x"FFDA";
          m(113) := x"0044";
          m(114) := x"0015";
          m(115) := x"0023";
          m(116) := x"003A";
          m(117) := x"005D";
          m(118) := x"009C";
          m(119) := x"020D";
          m(120) := x"069B";
          m(121) := x"077B";
          m(122) := x"06A3";
          m(123) := x"042E";
          m(124) := x"03DC";
          m(125) := x"0566";
          m(126) := x"0389";
          m(127) := x"038E";
          m(128) := x"03DA";
          m(129) := x"013B";
          m(130) := x"0528";
          m(131) := x"01F8";
          m(132) := x"026D";
          m(133) := x"FDE3";
          m(134) := x"FCAF";
          m(135) := x"F969";
          m(136) := x"FC3D";
          m(137) := x"FEE3";
          m(138) := x"FFFF";
          m(139) := x"0010";
          m(140) := x"000F";
          m(141) := x"0011";
          m(142) := x"000C";
          m(143) := x"003E";
          m(144) := x"0067";
          m(145) := x"0081";
          m(146) := x"0118";
          m(147) := x"037D";
          m(148) := x"050B";
          m(149) := x"05B8";
          m(150) := x"05DE";
          m(151) := x"0348";
          m(152) := x"04CE";
          m(153) := x"0279";
          m(154) := x"FF92";
          m(155) := x"FE13";
          m(156) := x"034D";
          m(157) := x"05E7";
          m(158) := x"04EE";
          m(159) := x"FF7E";
          m(160) := x"0528";
          m(161) := x"00CD";
          m(162) := x"FE02";
          m(163) := x"FD01";
          m(164) := x"FCA4";
          m(165) := x"FE72";
          m(166) := x"FFEF";
          m(167) := x"FFF8";
          m(168) := x"0000";
          m(169) := x"000C";
          m(170) := x"FFFB";
          m(171) := x"0097";
          m(172) := x"0176";
          m(173) := x"016E";
          m(174) := x"0117";
          m(175) := x"0404";
          m(176) := x"FD9B";
          m(177) := x"FF0E";
          m(178) := x"06F6";
          m(179) := x"0643";
          m(180) := x"FF8C";
          m(181) := x"07C3";
          m(182) := x"0721";
          m(183) := x"0240";
          m(184) := x"FE58";
          m(185) := x"001A";
          m(186) := x"06F8";
          m(187) := x"0482";
          m(188) := x"02CE";
          m(189) := x"FFE4";
          m(190) := x"01B6";
          m(191) := x"FE5A";
          m(192) := x"FEC9";
          m(193) := x"000C";
          m(194) := x"0062";
          m(195) := x"003B";
          m(196) := x"0033";
          m(197) := x"004E";
          m(198) := x"0024";
          m(199) := x"0139";
          m(200) := x"0236";
          m(201) := x"013B";
          m(202) := x"FFEB";
          m(203) := x"FF72";
          m(204) := x"FDBD";
          m(205) := x"FA2A";
          m(206) := x"FAD4";
          m(207) := x"074B";
          m(208) := x"039F";
          m(209) := x"00DF";
          m(210) := x"06FF";
          m(211) := x"0391";
          m(212) := x"0229";
          m(213) := x"0093";
          m(214) := x"FE9E";
          m(215) := x"0218";
          m(216) := x"FFDA";
          m(217) := x"FF16";
          m(218) := x"FE5D";
          m(219) := x"FEF3";
          m(220) := x"FC7C";
          m(221) := x"FDA3";
          m(222) := x"0082";
          m(223) := x"0033";
          m(224) := x"0039";
          m(225) := x"00AE";
          m(226) := x"0021";
          m(227) := x"0237";
          m(228) := x"010E";
          m(229) := x"FDBF";
          m(230) := x"FCC6";
          m(231) := x"FDC5";
          m(232) := x"FF0B";
          m(233) := x"FEA4";
          m(234) := x"0372";
          m(235) := x"004F";
          m(236) := x"00A8";
          m(237) := x"FDC5";
          m(238) := x"FDEC";
          m(239) := x"0121";
          m(240) := x"0815";
          m(241) := x"052E";
          m(242) := x"0060";
          m(243) := x"0343";
          m(244) := x"FC3E";
          m(245) := x"014F";
          m(246) := x"FDE2";
          m(247) := x"FE12";
          m(248) := x"FA29";
          m(249) := x"FF2F";
          m(250) := x"006B";
          m(251) := x"0046";
          m(252) := x"FFFD";
          m(253) := x"006D";
          m(254) := x"0165";
          m(255) := x"0088";
          m(256) := x"FD50";
          m(257) := x"F7AB";
          m(258) := x"F7C1";
          m(259) := x"F8AD";
          m(260) := x"F7AE";
          m(261) := x"F558";
          m(262) := x"F21B";
          m(263) := x"F28A";
          m(264) := x"EE78";
          m(265) := x"F191";
          m(266) := x"F7E0";
          m(267) := x"FECC";
          m(268) := x"0482";
          m(269) := x"01F2";
          m(270) := x"04DD";
          m(271) := x"FE5E";
          m(272) := x"FD09";
          m(273) := x"FEFF";
          m(274) := x"0241";
          m(275) := x"FCEF";
          m(276) := x"FC05";
          m(277) := x"014A";
          m(278) := x"000D";
          m(279) := x"003E";
          m(280) := x"FFF8";
          m(281) := x"00B2";
          m(282) := x"01CD";
          m(283) := x"005F";
          m(284) := x"F9D0";
          m(285) := x"F3A1";
          m(286) := x"F1CA";
          m(287) := x"EC67";
          m(288) := x"E552";
          m(289) := x"E82D";
          m(290) := x"EBAE";
          m(291) := x"EABC";
          m(292) := x"F1BA";
          m(293) := x"FE34";
          m(294) := x"FCE0";
          m(295) := x"FA3D";
          m(296) := x"036A";
          m(297) := x"077E";
          m(298) := x"FF42";
          m(299) := x"FE5A";
          m(300) := x"04E1";
          m(301) := x"0150";
          m(302) := x"FE04";
          m(303) := x"FA9D";
          m(304) := x"FDC0";
          m(305) := x"FF96";
          m(306) := x"002E";
          m(307) := x"FFD8";
          m(308) := x"0016";
          m(309) := x"006F";
          m(310) := x"01DE";
          m(311) := x"0053";
          m(312) := x"FA5B";
          m(313) := x"F426";
          m(314) := x"F346";
          m(315) := x"F39B";
          m(316) := x"F244";
          m(317) := x"F776";
          m(318) := x"F99B";
          m(319) := x"FD8E";
          m(320) := x"00FE";
          m(321) := x"005D";
          m(322) := x"0494";
          m(323) := x"04F8";
          m(324) := x"0086";
          m(325) := x"0554";
          m(326) := x"FDF8";
          m(327) := x"0122";
          m(328) := x"046E";
          m(329) := x"FFC3";
          m(330) := x"FD55";
          m(331) := x"FCB5";
          m(332) := x"FE12";
          m(333) := x"FEE2";
          m(334) := x"0002";
          m(335) := x"FFD7";
          m(336) := x"001E";
          m(337) := x"001D";
          m(338) := x"00E8";
          m(339) := x"0038";
          m(340) := x"FC3B";
          m(341) := x"FA1B";
          m(342) := x"F939";
          m(343) := x"FE58";
          m(344) := x"02A0";
          m(345) := x"02A9";
          m(346) := x"07E0";
          m(347) := x"07AE";
          m(348) := x"0666";
          m(349) := x"010E";
          m(350) := x"04D8";
          m(351) := x"00E5";
          m(352) := x"FEEB";
          m(353) := x"FCE3";
          m(354) := x"FF22";
          m(355) := x"0092";
          m(356) := x"FF65";
          m(357) := x"FDA4";
          m(358) := x"FEB9";
          m(359) := x"FCA0";
          m(360) := x"FEE4";
          m(361) := x"00AE";
          m(362) := x"0076";
          m(363) := x"0017";
          m(364) := x"0010";
          m(365) := x"0014";
          m(366) := x"00D4";
          m(367) := x"015E";
          m(368) := x"0028";
          m(369) := x"01C2";
          m(370) := x"02CE";
          m(371) := x"03AF";
          m(372) := x"087F";
          m(373) := x"06D2";
          m(374) := x"068D";
          m(375) := x"0584";
          m(376) := x"039C";
          m(377) := x"FFF4";
          m(378) := x"0379";
          m(379) := x"FE6E";
          m(380) := x"FE47";
          m(381) := x"FB52";
          m(382) := x"FFCF";
          m(383) := x"02AA";
          m(384) := x"05BD";
          m(385) := x"004F";
          m(386) := x"FB97";
          m(387) := x"FD84";
          m(388) := x"FF95";
          m(389) := x"0098";
          m(390) := x"0028";
          m(391) := x"0015";
          m(392) := x"0013";
          m(393) := x"FFD6";
          m(394) := x"005D";
          m(395) := x"0198";
          m(396) := x"0365";
          m(397) := x"0577";
          m(398) := x"0D7D";
          m(399) := x"0CF1";
          m(400) := x"0A03";
          m(401) := x"042B";
          m(402) := x"050B";
          m(403) := x"FF11";
          m(404) := x"FBC9";
          m(405) := x"FB7E";
          m(406) := x"0423";
          m(407) := x"FFE9";
          m(408) := x"00E7";
          m(409) := x"FE0C";
          m(410) := x"0130";
          m(411) := x"FDD5";
          m(412) := x"FE4D";
          m(413) := x"029A";
          m(414) := x"FEF1";
          m(415) := x"FEBD";
          m(416) := x"FEA4";
          m(417) := x"0064";
          m(418) := x"00CD";
          m(419) := x"FFE7";
          m(420) := x"0032";
          m(421) := x"FFFC";
          m(422) := x"0006";
          m(423) := x"02D9";
          m(424) := x"068A";
          m(425) := x"0848";
          m(426) := x"0873";
          m(427) := x"03F3";
          m(428) := x"FB6E";
          m(429) := x"006C";
          m(430) := x"FABA";
          m(431) := x"FC9B";
          m(432) := x"FF67";
          m(433) := x"028F";
          m(434) := x"FDBA";
          m(435) := x"FEE9";
          m(436) := x"FF7D";
          m(437) := x"F96E";
          m(438) := x"FCF4";
          m(439) := x"FD61";
          m(440) := x"F7CB";
          m(441) := x"FB6A";
          m(442) := x"FCFC";
          m(443) := x"FDAE";
          m(444) := x"FD60";
          m(445) := x"0082";
          m(446) := x"00B7";
          m(447) := x"FFDD";
          m(448) := x"000A";
          m(449) := x"0004";
          m(450) := x"0090";
          m(451) := x"048E";
          m(452) := x"03C0";
          m(453) := x"01F7";
          m(454) := x"00E8";
          m(455) := x"06D3";
          m(456) := x"FEED";
          m(457) := x"FD58";
          m(458) := x"FF6C";
          m(459) := x"0139";
          m(460) := x"FE9A";
          m(461) := x"FDAF";
          m(462) := x"0155";
          m(463) := x"FCB8";
          m(464) := x"FC5E";
          m(465) := x"FC75";
          m(466) := x"0169";
          m(467) := x"0088";
          m(468) := x"FB07";
          m(469) := x"FB81";
          m(470) := x"FD26";
          m(471) := x"FDF5";
          m(472) := x"FDC1";
          m(473) := x"0097";
          m(474) := x"00ED";
          m(475) := x"002B";
          m(476) := x"FFDF";
          m(477) := x"FFF1";
          m(478) := x"00B6";
          m(479) := x"0293";
          m(480) := x"000A";
          m(481) := x"FF86";
          m(482) := x"FE36";
          m(483) := x"FE0B";
          m(484) := x"FBAA";
          m(485) := x"FC33";
          m(486) := x"FA0A";
          m(487) := x"FE65";
          m(488) := x"FBE7";
          m(489) := x"0087";
          m(490) := x"FE7D";
          m(491) := x"FE9C";
          m(492) := x"FD89";
          m(493) := x"FCCF";
          m(494) := x"FB9B";
          m(495) := x"004A";
          m(496) := x"FC47";
          m(497) := x"FCCC";
          m(498) := x"0335";
          m(499) := x"FF03";
          m(500) := x"004C";
          m(501) := x"0379";
          m(502) := x"00B3";
          m(503) := x"FFB9";
          m(504) := x"FFFA";
          m(505) := x"0006";
          m(506) := x"00BF";
          m(507) := x"03BE";
          m(508) := x"FCA4";
          m(509) := x"FF36";
          m(510) := x"FD5D";
          m(511) := x"FF41";
          m(512) := x"011E";
          m(513) := x"02D8";
          m(514) := x"FDFF";
          m(515) := x"00CC";
          m(516) := x"FDD0";
          m(517) := x"0276";
          m(518) := x"FCD6";
          m(519) := x"FEA7";
          m(520) := x"0010";
          m(521) := x"027F";
          m(522) := x"FF80";
          m(523) := x"0262";
          m(524) := x"05BF";
          m(525) := x"040F";
          m(526) := x"045F";
          m(527) := x"FFC1";
          m(528) := x"021F";
          m(529) := x"032F";
          m(530) := x"0077";
          m(531) := x"0059";
          m(532) := x"FFCF";
          m(533) := x"FFD5";
          m(534) := x"FE2F";
          m(535) := x"02E7";
          m(536) := x"01F8";
          m(537) := x"FF80";
          m(538) := x"003F";
          m(539) := x"FDBB";
          m(540) := x"FA50";
          m(541) := x"FE5C";
          m(542) := x"FD0C";
          m(543) := x"FF81";
          m(544) := x"FFE0";
          m(545) := x"041A";
          m(546) := x"0246";
          m(547) := x"FF80";
          m(548) := x"066D";
          m(549) := x"0568";
          m(550) := x"FF32";
          m(551) := x"0388";
          m(552) := x"0224";
          m(553) := x"01A6";
          m(554) := x"00DF";
          m(555) := x"FEA4";
          m(556) := x"0060";
          m(557) := x"01D7";
          m(558) := x"004B";
          m(559) := x"0047";
          m(560) := x"003C";
          m(561) := x"FF9E";
          m(562) := x"FE1F";
          m(563) := x"00E4";
          m(564) := x"040C";
          m(565) := x"FEE7";
          m(566) := x"FFAA";
          m(567) := x"FB31";
          m(568) := x"FF95";
          m(569) := x"00F5";
          m(570) := x"FEF0";
          m(571) := x"FF1B";
          m(572) := x"030B";
          m(573) := x"0460";
          m(574) := x"02B4";
          m(575) := x"FC87";
          m(576) := x"0338";
          m(577) := x"FC79";
          m(578) := x"0377";
          m(579) := x"0000";
          m(580) := x"0084";
          m(581) := x"FEE1";
          m(582) := x"FFA7";
          m(583) := x"FEEC";
          m(584) := x"015E";
          m(585) := x"0122";
          m(586) := x"0040";
          m(587) := x"0007";
          m(588) := x"FFE5";
          m(589) := x"000C";
          m(590) := x"00B9";
          m(591) := x"00E0";
          m(592) := x"003B";
          m(593) := x"FFC8";
          m(594) := x"0136";
          m(595) := x"008B";
          m(596) := x"FC2B";
          m(597) := x"FBDE";
          m(598) := x"0355";
          m(599) := x"FC95";
          m(600) := x"FA9E";
          m(601) := x"FE78";
          m(602) := x"FE9C";
          m(603) := x"F934";
          m(604) := x"02D8";
          m(605) := x"0127";
          m(606) := x"0376";
          m(607) := x"00FA";
          m(608) := x"008D";
          m(609) := x"FE00";
          m(610) := x"FED8";
          m(611) := x"01BF";
          m(612) := x"01F5";
          m(613) := x"005C";
          m(614) := x"FFC0";
          m(615) := x"0020";
          m(616) := x"FFF6";
          m(617) := x"0004";
          m(618) := x"0046";
          m(619) := x"0055";
          m(620) := x"FFDC";
          m(621) := x"FFF0";
          m(622) := x"FFD8";
          m(623) := x"01A6";
          m(624) := x"FCF8";
          m(625) := x"F934";
          m(626) := x"FE7D";
          m(627) := x"FC8B";
          m(628) := x"FDE4";
          m(629) := x"FC9B";
          m(630) := x"02EA";
          m(631) := x"02A0";
          m(632) := x"FE1A";
          m(633) := x"FE72";
          m(634) := x"FBDE";
          m(635) := x"0115";
          m(636) := x"01B4";
          m(637) := x"FCDF";
          m(638) := x"FE62";
          m(639) := x"0052";
          m(640) := x"0001";
          m(641) := x"FFFD";
          m(642) := x"FFEE";
          m(643) := x"0019";
          m(644) := x"FFF9";
          m(645) := x"FFF8";
          m(646) := x"0045";
          m(647) := x"00AB";
          m(648) := x"0049";
          m(649) := x"0010";
          m(650) := x"FA51";
          m(651) := x"FC2D";
          m(652) := x"FCE4";
          m(653) := x"025B";
          m(654) := x"008B";
          m(655) := x"0032";
          m(656) := x"FE57";
          m(657) := x"FD5B";
          m(658) := x"FFA5";
          m(659) := x"FD26";
          m(660) := x"FD47";
          m(661) := x"FE79";
          m(662) := x"FB4B";
          m(663) := x"FC9E";
          m(664) := x"FEF0";
          m(665) := x"FFE7";
          m(666) := x"0166";
          m(667) := x"01CD";
          m(668) := x"FFCB";
          m(669) := x"0005";
          m(670) := x"003D";
          m(671) := x"0022";
          m(672) := x"0013";
          m(673) := x"FFF5";
          m(674) := x"0017";
          m(675) := x"006A";
          m(676) := x"003E";
          m(677) := x"FFFF";
          m(678) := x"FEC1";
          m(679) := x"FEC6";
          m(680) := x"011F";
          m(681) := x"0590";
          m(682) := x"FF79";
          m(683) := x"FEBF";
          m(684) := x"FCC9";
          m(685) := x"02F7";
          m(686) := x"0730";
          m(687) := x"010B";
          m(688) := x"FCF4";
          m(689) := x"FEF7";
          m(690) := x"FC13";
          m(691) := x"FCA5";
          m(692) := x"FE07";
          m(693) := x"011B";
          m(694) := x"0044";
          m(695) := x"0141";
          m(696) := x"00D5";
          m(697) := x"0012";
          m(698) := x"0019";
          m(699) := x"000B";
          m(700) := x"001F";
          m(701) := x"0010";
          m(702) := x"FFD9";
          m(703) := x"0000";
          m(704) := x"00BF";
          m(705) := x"0015";
          m(706) := x"FF0B";
          m(707) := x"FDC1";
          m(708) := x"010B";
          m(709) := x"0344";
          m(710) := x"0133";
          m(711) := x"FFDA";
          m(712) := x"04E1";
          m(713) := x"04DD";
          m(714) := x"02EE";
          m(715) := x"FF03";
          m(716) := x"FD43";
          m(717) := x"FFB7";
          m(718) := x"0132";
          m(719) := x"009E";
          m(720) := x"FE90";
          m(721) := x"FD98";
          m(722) := x"FF73";
          m(723) := x"001A";
          m(724) := x"FFDA";
          m(725) := x"FFE7";
          m(726) := x"FFF3";
          m(727) := x"0021";
          m(728) := x"0007";
          m(729) := x"FFDF";
          m(730) := x"FFEF";
          m(731) := x"0011";
          m(732) := x"FFCE";
          m(733) := x"FFD9";
          m(734) := x"FF35";
          m(735) := x"FE9A";
          m(736) := x"0177";
          m(737) := x"0171";
          m(738) := x"01E3";
          m(739) := x"0135";
          m(740) := x"FEB8";
          m(741) := x"FF95";
          m(742) := x"FEFD";
          m(743) := x"FFD2";
          m(744) := x"012E";
          m(745) := x"00D4";
          m(746) := x"FF87";
          m(747) := x"FFE1";
          m(748) := x"000F";
          m(749) := x"0008";
          m(750) := x"005C";
          m(751) := x"FFF7";
          m(752) := x"FFFE";
          m(753) := x"0007";
          m(754) := x"FFFE";
          m(755) := x"FFE8";
          m(756) := x"0032";
          m(757) := x"0025";
          m(758) := x"FFE6";
          m(759) := x"0039";
          m(760) := x"0015";
          m(761) := x"FFF4";
          m(762) := x"FFC6";
          m(763) := x"FF36";
          m(764) := x"FF3F";
          m(765) := x"0012";
          m(766) := x"FFEB";
          m(767) := x"FFFC";
          m(768) := x"FF9C";
          m(769) := x"FFAC";
          m(770) := x"0018";
          m(771) := x"FFDF";
          m(772) := x"0040";
          m(773) := x"FFF7";
          m(774) := x"FFD4";
          m(775) := x"0002";
          m(776) := x"0029";
          m(777) := x"FFF7";
          m(778) := x"0022";
          m(779) := x"FFCC";
          m(780) := x"FFF2";
          m(781) := x"0035";
          m(782) := x"0035";
          m(783) := x"FFD1";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_11.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 11) then
          m(0) := x"FFF6";
          m(1) := x"FFDD";
          m(2) := x"FFDB";
          m(3) := x"0001";
          m(4) := x"FFE8";
          m(5) := x"FFF5";
          m(6) := x"FFE8";
          m(7) := x"FFF6";
          m(8) := x"FFD5";
          m(9) := x"FFD3";
          m(10) := x"0007";
          m(11) := x"0015";
          m(12) := x"0000";
          m(13) := x"0020";
          m(14) := x"FFDD";
          m(15) := x"0013";
          m(16) := x"FFFA";
          m(17) := x"FFED";
          m(18) := x"FFCF";
          m(19) := x"0017";
          m(20) := x"FFE7";
          m(21) := x"000B";
          m(22) := x"001A";
          m(23) := x"FFF2";
          m(24) := x"001F";
          m(25) := x"FFE9";
          m(26) := x"FFDD";
          m(27) := x"000A";
          m(28) := x"FFF3";
          m(29) := x"FFD6";
          m(30) := x"FFE9";
          m(31) := x"FFEF";
          m(32) := x"FFE7";
          m(33) := x"FFEB";
          m(34) := x"001F";
          m(35) := x"FFE4";
          m(36) := x"FFEF";
          m(37) := x"FFF8";
          m(38) := x"FFFB";
          m(39) := x"0003";
          m(40) := x"0002";
          m(41) := x"0005";
          m(42) := x"FFFD";
          m(43) := x"FFF9";
          m(44) := x"FF5E";
          m(45) := x"FFDD";
          m(46) := x"FFE1";
          m(47) := x"000C";
          m(48) := x"FFFB";
          m(49) := x"FFE8";
          m(50) := x"0006";
          m(51) := x"001F";
          m(52) := x"FFBF";
          m(53) := x"000F";
          m(54) := x"FFF2";
          m(55) := x"0050";
          m(56) := x"0007";
          m(57) := x"FFFE";
          m(58) := x"FFF8";
          m(59) := x"FFDF";
          m(60) := x"001C";
          m(61) := x"001B";
          m(62) := x"0017";
          m(63) := x"005B";
          m(64) := x"0009";
          m(65) := x"0025";
          m(66) := x"FFE2";
          m(67) := x"0013";
          m(68) := x"002F";
          m(69) := x"006E";
          m(70) := x"005F";
          m(71) := x"FF8E";
          m(72) := x"FEA1";
          m(73) := x"FF59";
          m(74) := x"FEB1";
          m(75) := x"FFF8";
          m(76) := x"FF98";
          m(77) := x"FFFA";
          m(78) := x"0036";
          m(79) := x"002F";
          m(80) := x"0009";
          m(81) := x"0012";
          m(82) := x"0005";
          m(83) := x"FFDD";
          m(84) := x"FFE4";
          m(85) := x"FFF1";
          m(86) := x"0014";
          m(87) := x"FFA8";
          m(88) := x"0022";
          m(89) := x"000A";
          m(90) := x"0054";
          m(91) := x"009E";
          m(92) := x"FEE3";
          m(93) := x"FE99";
          m(94) := x"FD96";
          m(95) := x"0080";
          m(96) := x"FF02";
          m(97) := x"FEDD";
          m(98) := x"0169";
          m(99) := x"0004";
          m(100) := x"0077";
          m(101) := x"FE67";
          m(102) := x"FAF3";
          m(103) := x"FC17";
          m(104) := x"FE07";
          m(105) := x"FFC1";
          m(106) := x"0051";
          m(107) := x"00B3";
          m(108) := x"011E";
          m(109) := x"003E";
          m(110) := x"0020";
          m(111) := x"0011";
          m(112) := x"FFE3";
          m(113) := x"000C";
          m(114) := x"FFF7";
          m(115) := x"FFFA";
          m(116) := x"0020";
          m(117) := x"00A4";
          m(118) := x"00D7";
          m(119) := x"000F";
          m(120) := x"FF28";
          m(121) := x"FE8B";
          m(122) := x"FF5B";
          m(123) := x"FC77";
          m(124) := x"FECD";
          m(125) := x"01DD";
          m(126) := x"0161";
          m(127) := x"FFD8";
          m(128) := x"010C";
          m(129) := x"FE34";
          m(130) := x"F8E8";
          m(131) := x"FCA1";
          m(132) := x"FEDD";
          m(133) := x"FF9D";
          m(134) := x"01B5";
          m(135) := x"033E";
          m(136) := x"02DA";
          m(137) := x"007F";
          m(138) := x"FFDE";
          m(139) := x"FFFA";
          m(140) := x"FFEF";
          m(141) := x"FFF3";
          m(142) := x"FFE9";
          m(143) := x"FFD3";
          m(144) := x"FFE5";
          m(145) := x"FFD7";
          m(146) := x"0096";
          m(147) := x"00CA";
          m(148) := x"00EA";
          m(149) := x"FDA9";
          m(150) := x"FF2A";
          m(151) := x"FA18";
          m(152) := x"FD3C";
          m(153) := x"FCD2";
          m(154) := x"FCFC";
          m(155) := x"FD49";
          m(156) := x"FCA8";
          m(157) := x"FC7F";
          m(158) := x"F83C";
          m(159) := x"F8A2";
          m(160) := x"F9F7";
          m(161) := x"FE31";
          m(162) := x"00D4";
          m(163) := x"04C9";
          m(164) := x"0384";
          m(165) := x"01C0";
          m(166) := x"FFF1";
          m(167) := x"0026";
          m(168) := x"FFD0";
          m(169) := x"FFBE";
          m(170) := x"FF90";
          m(171) := x"FF97";
          m(172) := x"007D";
          m(173) := x"FFFB";
          m(174) := x"00F3";
          m(175) := x"02ED";
          m(176) := x"02DB";
          m(177) := x"006E";
          m(178) := x"023C";
          m(179) := x"FCE1";
          m(180) := x"031A";
          m(181) := x"0000";
          m(182) := x"FE60";
          m(183) := x"FA55";
          m(184) := x"F9E0";
          m(185) := x"FC44";
          m(186) := x"FAA9";
          m(187) := x"0003";
          m(188) := x"FF61";
          m(189) := x"0175";
          m(190) := x"FF76";
          m(191) := x"03D1";
          m(192) := x"01BC";
          m(193) := x"FF4A";
          m(194) := x"FF57";
          m(195) := x"0000";
          m(196) := x"0019";
          m(197) := x"FFFA";
          m(198) := x"0048";
          m(199) := x"00A9";
          m(200) := x"004A";
          m(201) := x"FEA6";
          m(202) := x"FE7E";
          m(203) := x"FFB0";
          m(204) := x"0020";
          m(205) := x"0242";
          m(206) := x"FE12";
          m(207) := x"015D";
          m(208) := x"02E4";
          m(209) := x"03E8";
          m(210) := x"0039";
          m(211) := x"FE7E";
          m(212) := x"F6BC";
          m(213) := x"F7B2";
          m(214) := x"F841";
          m(215) := x"FD9E";
          m(216) := x"0190";
          m(217) := x"FE80";
          m(218) := x"FEFA";
          m(219) := x"044D";
          m(220) := x"035F";
          m(221) := x"00F7";
          m(222) := x"FF00";
          m(223) := x"FFE7";
          m(224) := x"FFE6";
          m(225) := x"0005";
          m(226) := x"004D";
          m(227) := x"FF96";
          m(228) := x"FE69";
          m(229) := x"FEF2";
          m(230) := x"FEB3";
          m(231) := x"0070";
          m(232) := x"0194";
          m(233) := x"0028";
          m(234) := x"FF1F";
          m(235) := x"0253";
          m(236) := x"0497";
          m(237) := x"FD50";
          m(238) := x"0099";
          m(239) := x"0508";
          m(240) := x"FA53";
          m(241) := x"F2B9";
          m(242) := x"F620";
          m(243) := x"FA66";
          m(244) := x"00C5";
          m(245) := x"FF13";
          m(246) := x"FEFA";
          m(247) := x"002E";
          m(248) := x"FFC4";
          m(249) := x"FCD3";
          m(250) := x"FEFD";
          m(251) := x"FFBF";
          m(252) := x"FFD6";
          m(253) := x"FFFD";
          m(254) := x"FFF9";
          m(255) := x"000E";
          m(256) := x"00AD";
          m(257) := x"033F";
          m(258) := x"0021";
          m(259) := x"0133";
          m(260) := x"FF7C";
          m(261) := x"012E";
          m(262) := x"FF61";
          m(263) := x"FD16";
          m(264) := x"FA47";
          m(265) := x"FAF4";
          m(266) := x"01B4";
          m(267) := x"FA42";
          m(268) := x"FECF";
          m(269) := x"FF96";
          m(270) := x"FAB5";
          m(271) := x"F84F";
          m(272) := x"FE67";
          m(273) := x"0187";
          m(274) := x"FE82";
          m(275) := x"FF74";
          m(276) := x"FC48";
          m(277) := x"FCE6";
          m(278) := x"FDD9";
          m(279) := x"FF74";
          m(280) := x"001F";
          m(281) := x"0066";
          m(282) := x"002E";
          m(283) := x"FFE8";
          m(284) := x"0053";
          m(285) := x"01AF";
          m(286) := x"0226";
          m(287) := x"025A";
          m(288) := x"0141";
          m(289) := x"FF72";
          m(290) := x"FEC7";
          m(291) := x"FC6D";
          m(292) := x"F9C6";
          m(293) := x"FB34";
          m(294) := x"F794";
          m(295) := x"F9C2";
          m(296) := x"0053";
          m(297) := x"06A6";
          m(298) := x"02FF";
          m(299) := x"FBE8";
          m(300) := x"F863";
          m(301) := x"FF49";
          m(302) := x"FDCD";
          m(303) := x"F9B1";
          m(304) := x"F931";
          m(305) := x"FD00";
          m(306) := x"FE22";
          m(307) := x"FFF3";
          m(308) := x"FFE9";
          m(309) := x"0047";
          m(310) := x"FF7F";
          m(311) := x"00EF";
          m(312) := x"FEB3";
          m(313) := x"01C1";
          m(314) := x"04AE";
          m(315) := x"03D5";
          m(316) := x"FBF4";
          m(317) := x"0420";
          m(318) := x"0447";
          m(319) := x"FC79";
          m(320) := x"FFB9";
          m(321) := x"FE38";
          m(322) := x"FE15";
          m(323) := x"FE3B";
          m(324) := x"032B";
          m(325) := x"06A0";
          m(326) := x"0461";
          m(327) := x"FEC8";
          m(328) := x"FA69";
          m(329) := x"FE95";
          m(330) := x"FE01";
          m(331) := x"F898";
          m(332) := x"F60B";
          m(333) := x"FC07";
          m(334) := x"FED7";
          m(335) := x"FFC9";
          m(336) := x"FFF9";
          m(337) := x"FFF4";
          m(338) := x"0055";
          m(339) := x"0235";
          m(340) := x"FF96";
          m(341) := x"0193";
          m(342) := x"004D";
          m(343) := x"0090";
          m(344) := x"01C0";
          m(345) := x"0028";
          m(346) := x"00E1";
          m(347) := x"012D";
          m(348) := x"045C";
          m(349) := x"FD4C";
          m(350) := x"F723";
          m(351) := x"018E";
          m(352) := x"08C4";
          m(353) := x"05C7";
          m(354) := x"0640";
          m(355) := x"FECC";
          m(356) := x"FCFC";
          m(357) := x"01F2";
          m(358) := x"015A";
          m(359) := x"FC3F";
          m(360) := x"FE3B";
          m(361) := x"FE2F";
          m(362) := x"FF54";
          m(363) := x"FFFD";
          m(364) := x"0038";
          m(365) := x"FFDD";
          m(366) := x"004A";
          m(367) := x"0216";
          m(368) := x"020A";
          m(369) := x"FF5E";
          m(370) := x"0103";
          m(371) := x"0204";
          m(372) := x"FE4A";
          m(373) := x"00A4";
          m(374) := x"05C1";
          m(375) := x"048A";
          m(376) := x"FBC7";
          m(377) := x"F71F";
          m(378) := x"02D3";
          m(379) := x"02DB";
          m(380) := x"023E";
          m(381) := x"06CB";
          m(382) := x"0616";
          m(383) := x"02BF";
          m(384) := x"FF3A";
          m(385) := x"00D1";
          m(386) := x"04B3";
          m(387) := x"FF5A";
          m(388) := x"FFA6";
          m(389) := x"009F";
          m(390) := x"001B";
          m(391) := x"0012";
          m(392) := x"000C";
          m(393) := x"FF86";
          m(394) := x"0018";
          m(395) := x"0221";
          m(396) := x"032C";
          m(397) := x"02B7";
          m(398) := x"00F3";
          m(399) := x"0223";
          m(400) := x"01CB";
          m(401) := x"FF7D";
          m(402) := x"0417";
          m(403) := x"FE7A";
          m(404) := x"F8A2";
          m(405) := x"FBE7";
          m(406) := x"055D";
          m(407) := x"02B9";
          m(408) := x"034D";
          m(409) := x"0488";
          m(410) := x"0234";
          m(411) := x"052E";
          m(412) := x"FE77";
          m(413) := x"000D";
          m(414) := x"0401";
          m(415) := x"013D";
          m(416) := x"FE5A";
          m(417) := x"0251";
          m(418) := x"FFCF";
          m(419) := x"FFFC";
          m(420) := x"FFBB";
          m(421) := x"FF41";
          m(422) := x"0080";
          m(423) := x"037D";
          m(424) := x"0318";
          m(425) := x"FDC4";
          m(426) := x"FB9F";
          m(427) := x"00FD";
          m(428) := x"0003";
          m(429) := x"0136";
          m(430) := x"0213";
          m(431) := x"FA23";
          m(432) := x"F3A9";
          m(433) := x"0082";
          m(434) := x"0889";
          m(435) := x"0BB4";
          m(436) := x"0105";
          m(437) := x"004C";
          m(438) := x"0236";
          m(439) := x"FF02";
          m(440) := x"0287";
          m(441) := x"00B0";
          m(442) := x"024D";
          m(443) := x"FDD9";
          m(444) := x"00D0";
          m(445) := x"01ED";
          m(446) := x"FFF4";
          m(447) := x"0009";
          m(448) := x"001E";
          m(449) := x"FFE2";
          m(450) := x"FF35";
          m(451) := x"00CD";
          m(452) := x"01F3";
          m(453) := x"FECB";
          m(454) := x"FEC0";
          m(455) := x"01D7";
          m(456) := x"019D";
          m(457) := x"0053";
          m(458) := x"F9C3";
          m(459) := x"F4C7";
          m(460) := x"FE06";
          m(461) := x"0AC3";
          m(462) := x"0FD4";
          m(463) := x"05F5";
          m(464) := x"FED1";
          m(465) := x"0230";
          m(466) := x"0213";
          m(467) := x"0079";
          m(468) := x"04FE";
          m(469) := x"0066";
          m(470) := x"FA53";
          m(471) := x"026B";
          m(472) := x"0348";
          m(473) := x"01AB";
          m(474) := x"FFC9";
          m(475) := x"0000";
          m(476) := x"000E";
          m(477) := x"FFC5";
          m(478) := x"FF30";
          m(479) := x"FE8C";
          m(480) := x"01B0";
          m(481) := x"FEE5";
          m(482) := x"FDCC";
          m(483) := x"FF90";
          m(484) := x"00DA";
          m(485) := x"FD19";
          m(486) := x"FA4F";
          m(487) := x"F989";
          m(488) := x"0744";
          m(489) := x"0AD7";
          m(490) := x"07F2";
          m(491) := x"FF1C";
          m(492) := x"0056";
          m(493) := x"0453";
          m(494) := x"0200";
          m(495) := x"FD46";
          m(496) := x"007C";
          m(497) := x"008A";
          m(498) := x"00E6";
          m(499) := x"005C";
          m(500) := x"031F";
          m(501) := x"0202";
          m(502) := x"00A7";
          m(503) := x"FFED";
          m(504) := x"000B";
          m(505) := x"FFF0";
          m(506) := x"FF76";
          m(507) := x"FF70";
          m(508) := x"032A";
          m(509) := x"FE91";
          m(510) := x"FCC2";
          m(511) := x"FE7D";
          m(512) := x"FCEE";
          m(513) := x"F598";
          m(514) := x"F68E";
          m(515) := x"021A";
          m(516) := x"07FA";
          m(517) := x"046E";
          m(518) := x"00E1";
          m(519) := x"FE24";
          m(520) := x"028D";
          m(521) := x"01D8";
          m(522) := x"0300";
          m(523) := x"FD6F";
          m(524) := x"FBFD";
          m(525) := x"FD9C";
          m(526) := x"FD36";
          m(527) := x"FB29";
          m(528) := x"0087";
          m(529) := x"00FD";
          m(530) := x"0083";
          m(531) := x"006D";
          m(532) := x"FFE6";
          m(533) := x"FFE6";
          m(534) := x"FFED";
          m(535) := x"FF40";
          m(536) := x"026D";
          m(537) := x"FEEE";
          m(538) := x"FD35";
          m(539) := x"FFE9";
          m(540) := x"FBD9";
          m(541) := x"F9E3";
          m(542) := x"FBBF";
          m(543) := x"FFFB";
          m(544) := x"03C1";
          m(545) := x"065B";
          m(546) := x"01E6";
          m(547) := x"03F3";
          m(548) := x"02F3";
          m(549) := x"018E";
          m(550) := x"02CC";
          m(551) := x"FE8F";
          m(552) := x"FF20";
          m(553) := x"FCC2";
          m(554) := x"FA59";
          m(555) := x"FA53";
          m(556) := x"FF75";
          m(557) := x"FFA4";
          m(558) := x"0007";
          m(559) := x"FFE6";
          m(560) := x"FFF6";
          m(561) := x"FFCF";
          m(562) := x"0016";
          m(563) := x"FF19";
          m(564) := x"01C0";
          m(565) := x"0064";
          m(566) := x"FB92";
          m(567) := x"FC75";
          m(568) := x"F98C";
          m(569) := x"F6A5";
          m(570) := x"FC41";
          m(571) := x"FFC7";
          m(572) := x"0416";
          m(573) := x"0398";
          m(574) := x"01C5";
          m(575) := x"03E3";
          m(576) := x"05F2";
          m(577) := x"0622";
          m(578) := x"03B9";
          m(579) := x"FE4B";
          m(580) := x"00C7";
          m(581) := x"FB58";
          m(582) := x"F797";
          m(583) := x"FAF8";
          m(584) := x"00B1";
          m(585) := x"0049";
          m(586) := x"003C";
          m(587) := x"0014";
          m(588) := x"0007";
          m(589) := x"0006";
          m(590) := x"FF9C";
          m(591) := x"FEE7";
          m(592) := x"FF58";
          m(593) := x"FE77";
          m(594) := x"FB62";
          m(595) := x"FA69";
          m(596) := x"FCFD";
          m(597) := x"FC3D";
          m(598) := x"FC15";
          m(599) := x"FE61";
          m(600) := x"FF0F";
          m(601) := x"FCA2";
          m(602) := x"038A";
          m(603) := x"00B1";
          m(604) := x"0178";
          m(605) := x"FEF6";
          m(606) := x"FECF";
          m(607) := x"FD5A";
          m(608) := x"FDCF";
          m(609) := x"FBA5";
          m(610) := x"FB6B";
          m(611) := x"FFC4";
          m(612) := x"FFD1";
          m(613) := x"01A6";
          m(614) := x"0028";
          m(615) := x"FFE4";
          m(616) := x"FFF1";
          m(617) := x"FFFD";
          m(618) := x"FFA8";
          m(619) := x"FEEF";
          m(620) := x"FE02";
          m(621) := x"FC79";
          m(622) := x"FB3A";
          m(623) := x"FE11";
          m(624) := x"0293";
          m(625) := x"FE08";
          m(626) := x"FC2A";
          m(627) := x"FDE3";
          m(628) := x"FD2D";
          m(629) := x"FBF4";
          m(630) := x"0314";
          m(631) := x"FE9C";
          m(632) := x"FFE3";
          m(633) := x"01B4";
          m(634) := x"00A4";
          m(635) := x"FFAC";
          m(636) := x"FE6B";
          m(637) := x"FEED";
          m(638) := x"FDBF";
          m(639) := x"FEAD";
          m(640) := x"FF3B";
          m(641) := x"009F";
          m(642) := x"0004";
          m(643) := x"002B";
          m(644) := x"0005";
          m(645) := x"0024";
          m(646) := x"FF9C";
          m(647) := x"FE93";
          m(648) := x"FD3C";
          m(649) := x"FD4F";
          m(650) := x"FE81";
          m(651) := x"FF51";
          m(652) := x"FD90";
          m(653) := x"FB9A";
          m(654) := x"FA6F";
          m(655) := x"FA49";
          m(656) := x"FD8D";
          m(657) := x"F9BD";
          m(658) := x"0315";
          m(659) := x"FD85";
          m(660) := x"009A";
          m(661) := x"0239";
          m(662) := x"03CE";
          m(663) := x"012E";
          m(664) := x"FF02";
          m(665) := x"FFFF";
          m(666) := x"FEBF";
          m(667) := x"FEC8";
          m(668) := x"FE81";
          m(669) := x"FFF8";
          m(670) := x"FFDC";
          m(671) := x"FFDF";
          m(672) := x"FFCC";
          m(673) := x"005A";
          m(674) := x"FF7E";
          m(675) := x"FE8F";
          m(676) := x"FF60";
          m(677) := x"0041";
          m(678) := x"003A";
          m(679) := x"FC3F";
          m(680) := x"FDC0";
          m(681) := x"FD83";
          m(682) := x"FC25";
          m(683) := x"FC43";
          m(684) := x"FAFC";
          m(685) := x"FD13";
          m(686) := x"FE35";
          m(687) := x"FFB2";
          m(688) := x"0392";
          m(689) := x"FDB7";
          m(690) := x"0061";
          m(691) := x"03DE";
          m(692) := x"006D";
          m(693) := x"00A9";
          m(694) := x"0169";
          m(695) := x"00F6";
          m(696) := x"004F";
          m(697) := x"00A8";
          m(698) := x"002C";
          m(699) := x"FFF2";
          m(700) := x"0036";
          m(701) := x"FFF5";
          m(702) := x"FFB6";
          m(703) := x"0027";
          m(704) := x"008A";
          m(705) := x"FF7E";
          m(706) := x"FEFA";
          m(707) := x"FDF1";
          m(708) := x"FDF7";
          m(709) := x"FE6E";
          m(710) := x"0009";
          m(711) := x"00AA";
          m(712) := x"FF32";
          m(713) := x"0090";
          m(714) := x"0064";
          m(715) := x"017F";
          m(716) := x"FD89";
          m(717) := x"FB5F";
          m(718) := x"FD6E";
          m(719) := x"FCC7";
          m(720) := x"FE5D";
          m(721) := x"FE92";
          m(722) := x"FEE5";
          m(723) := x"FF9F";
          m(724) := x"FFD4";
          m(725) := x"FFF0";
          m(726) := x"0041";
          m(727) := x"0029";
          m(728) := x"FFE8";
          m(729) := x"0012";
          m(730) := x"FFD4";
          m(731) := x"FFE7";
          m(732) := x"FF75";
          m(733) := x"FF2B";
          m(734) := x"FEF8";
          m(735) := x"FDF5";
          m(736) := x"FE2E";
          m(737) := x"FCC9";
          m(738) := x"FA79";
          m(739) := x"FC6C";
          m(740) := x"FC4A";
          m(741) := x"F9CD";
          m(742) := x"FB04";
          m(743) := x"FE67";
          m(744) := x"FFA0";
          m(745) := x"FDE5";
          m(746) := x"FECA";
          m(747) := x"FF83";
          m(748) := x"FDE0";
          m(749) := x"FD79";
          m(750) := x"FFA7";
          m(751) := x"FFE8";
          m(752) := x"FFC5";
          m(753) := x"FFD7";
          m(754) := x"000E";
          m(755) := x"FFD9";
          m(756) := x"002E";
          m(757) := x"FFFA";
          m(758) := x"0000";
          m(759) := x"FFFE";
          m(760) := x"000D";
          m(761) := x"0010";
          m(762) := x"FFD4";
          m(763) := x"FF60";
          m(764) := x"FF56";
          m(765) := x"FFC1";
          m(766) := x"FF62";
          m(767) := x"FF7A";
          m(768) := x"FF48";
          m(769) := x"FFE6";
          m(770) := x"FF79";
          m(771) := x"FF9A";
          m(772) := x"005A";
          m(773) := x"FFF4";
          m(774) := x"FF1E";
          m(775) := x"FFFA";
          m(776) := x"005C";
          m(777) := x"0012";
          m(778) := x"FFE5";
          m(779) := x"FFDF";
          m(780) := x"FFF2";
          m(781) := x"FFF1";
          m(782) := x"FFE2";
          m(783) := x"FFBE";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_12.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 12) then
          m(0) := x"0027";
          m(1) := x"000B";
          m(2) := x"FFFF";
          m(3) := x"FFF5";
          m(4) := x"FFDF";
          m(5) := x"001B";
          m(6) := x"FFB3";
          m(7) := x"FFF7";
          m(8) := x"003F";
          m(9) := x"FFE7";
          m(10) := x"001D";
          m(11) := x"FFE4";
          m(12) := x"FFE2";
          m(13) := x"FFFC";
          m(14) := x"FFFD";
          m(15) := x"0012";
          m(16) := x"0020";
          m(17) := x"001C";
          m(18) := x"FFFA";
          m(19) := x"002E";
          m(20) := x"0014";
          m(21) := x"0034";
          m(22) := x"FFDA";
          m(23) := x"FFEE";
          m(24) := x"001F";
          m(25) := x"003B";
          m(26) := x"FFE0";
          m(27) := x"0008";
          m(28) := x"FFC4";
          m(29) := x"000C";
          m(30) := x"0002";
          m(31) := x"FFDA";
          m(32) := x"0016";
          m(33) := x"FFF2";
          m(34) := x"FFFC";
          m(35) := x"FFC0";
          m(36) := x"FFCF";
          m(37) := x"FFC9";
          m(38) := x"0000";
          m(39) := x"0015";
          m(40) := x"FF90";
          m(41) := x"FFBC";
          m(42) := x"FFA8";
          m(43) := x"FF68";
          m(44) := x"FF97";
          m(45) := x"FFF0";
          m(46) := x"0018";
          m(47) := x"FFA6";
          m(48) := x"0004";
          m(49) := x"FFCD";
          m(50) := x"FFDC";
          m(51) := x"0000";
          m(52) := x"0059";
          m(53) := x"0023";
          m(54) := x"FFE4";
          m(55) := x"000E";
          m(56) := x"FFF2";
          m(57) := x"FFEE";
          m(58) := x"FFEC";
          m(59) := x"0001";
          m(60) := x"0032";
          m(61) := x"FFD5";
          m(62) := x"0007";
          m(63) := x"FFB0";
          m(64) := x"FFBE";
          m(65) := x"FFC0";
          m(66) := x"FFD6";
          m(67) := x"FFE2";
          m(68) := x"FF73";
          m(69) := x"FF71";
          m(70) := x"FF9A";
          m(71) := x"FF5C";
          m(72) := x"FF2E";
          m(73) := x"0034";
          m(74) := x"FFD9";
          m(75) := x"0046";
          m(76) := x"0062";
          m(77) := x"007C";
          m(78) := x"002A";
          m(79) := x"FFDA";
          m(80) := x"0014";
          m(81) := x"FFF1";
          m(82) := x"FFF1";
          m(83) := x"0030";
          m(84) := x"0026";
          m(85) := x"002D";
          m(86) := x"FFE1";
          m(87) := x"0006";
          m(88) := x"FFD1";
          m(89) := x"FFFD";
          m(90) := x"FFEA";
          m(91) := x"FFD4";
          m(92) := x"FF5E";
          m(93) := x"FF99";
          m(94) := x"FF56";
          m(95) := x"FFCA";
          m(96) := x"FEA0";
          m(97) := x"FD7D";
          m(98) := x"FF72";
          m(99) := x"00EA";
          m(100) := x"037B";
          m(101) := x"04E4";
          m(102) := x"01E4";
          m(103) := x"0233";
          m(104) := x"033F";
          m(105) := x"00B1";
          m(106) := x"0030";
          m(107) := x"FFFA";
          m(108) := x"000F";
          m(109) := x"FFF4";
          m(110) := x"FFF8";
          m(111) := x"000F";
          m(112) := x"000E";
          m(113) := x"000A";
          m(114) := x"FFD0";
          m(115) := x"FFE4";
          m(116) := x"0004";
          m(117) := x"FFCC";
          m(118) := x"FFCC";
          m(119) := x"FFD1";
          m(120) := x"FF43";
          m(121) := x"FE2C";
          m(122) := x"FED9";
          m(123) := x"FF20";
          m(124) := x"FFDE";
          m(125) := x"00CB";
          m(126) := x"FA7F";
          m(127) := x"FAF3";
          m(128) := x"00CA";
          m(129) := x"02AE";
          m(130) := x"014B";
          m(131) := x"03C7";
          m(132) := x"FF96";
          m(133) := x"FD01";
          m(134) := x"FE1D";
          m(135) := x"0021";
          m(136) := x"FF6F";
          m(137) := x"FEEB";
          m(138) := x"FF18";
          m(139) := x"FFED";
          m(140) := x"0001";
          m(141) := x"0043";
          m(142) := x"FFBF";
          m(143) := x"FFD5";
          m(144) := x"FFF8";
          m(145) := x"FFED";
          m(146) := x"FDA9";
          m(147) := x"FCCA";
          m(148) := x"FF31";
          m(149) := x"FD9E";
          m(150) := x"FC27";
          m(151) := x"FDF4";
          m(152) := x"008C";
          m(153) := x"FE37";
          m(154) := x"FD2E";
          m(155) := x"02DE";
          m(156) := x"FBA5";
          m(157) := x"F92F";
          m(158) := x"FE04";
          m(159) := x"FDA4";
          m(160) := x"FE21";
          m(161) := x"F943";
          m(162) := x"FD20";
          m(163) := x"018A";
          m(164) := x"0071";
          m(165) := x"FEE7";
          m(166) := x"FF45";
          m(167) := x"0000";
          m(168) := x"0005";
          m(169) := x"0027";
          m(170) := x"FFD6";
          m(171) := x"FFA0";
          m(172) := x"FFD0";
          m(173) := x"FF9B";
          m(174) := x"FEA8";
          m(175) := x"FF2E";
          m(176) := x"01E6";
          m(177) := x"FC70";
          m(178) := x"FBC8";
          m(179) := x"FE0A";
          m(180) := x"0230";
          m(181) := x"FF96";
          m(182) := x"FE75";
          m(183) := x"FF37";
          m(184) := x"FF0E";
          m(185) := x"FDF6";
          m(186) := x"024C";
          m(187) := x"FC8F";
          m(188) := x"F9D2";
          m(189) := x"FF9E";
          m(190) := x"0399";
          m(191) := x"009E";
          m(192) := x"FF11";
          m(193) := x"FD6E";
          m(194) := x"FFE6";
          m(195) := x"FFF9";
          m(196) := x"0037";
          m(197) := x"FFBA";
          m(198) := x"FFB3";
          m(199) := x"FFED";
          m(200) := x"FFBA";
          m(201) := x"FE2F";
          m(202) := x"0231";
          m(203) := x"FE96";
          m(204) := x"FE4E";
          m(205) := x"01F6";
          m(206) := x"FC71";
          m(207) := x"FF15";
          m(208) := x"01A8";
          m(209) := x"049C";
          m(210) := x"0736";
          m(211) := x"FDE7";
          m(212) := x"0393";
          m(213) := x"05F5";
          m(214) := x"FED9";
          m(215) := x"FD9B";
          m(216) := x"FC82";
          m(217) := x"FD22";
          m(218) := x"01E0";
          m(219) := x"028B";
          m(220) := x"FFEF";
          m(221) := x"FE91";
          m(222) := x"023D";
          m(223) := x"FFD8";
          m(224) := x"0033";
          m(225) := x"FFDD";
          m(226) := x"FFBA";
          m(227) := x"FFE6";
          m(228) := x"009C";
          m(229) := x"0314";
          m(230) := x"05B0";
          m(231) := x"0259";
          m(232) := x"0584";
          m(233) := x"00F3";
          m(234) := x"00B9";
          m(235) := x"FF7F";
          m(236) := x"FFE8";
          m(237) := x"FE5F";
          m(238) := x"0145";
          m(239) := x"FECC";
          m(240) := x"F8E3";
          m(241) := x"007C";
          m(242) := x"00E9";
          m(243) := x"FA7F";
          m(244) := x"F905";
          m(245) := x"FB20";
          m(246) := x"FEEC";
          m(247) := x"FE82";
          m(248) := x"FFB9";
          m(249) := x"FEE6";
          m(250) := x"0047";
          m(251) := x"FF98";
          m(252) := x"0000";
          m(253) := x"0006";
          m(254) := x"FFC3";
          m(255) := x"FF31";
          m(256) := x"006D";
          m(257) := x"03B6";
          m(258) := x"0185";
          m(259) := x"FE63";
          m(260) := x"00EE";
          m(261) := x"FCC7";
          m(262) := x"FFFE";
          m(263) := x"FDEE";
          m(264) := x"0146";
          m(265) := x"011C";
          m(266) := x"0268";
          m(267) := x"031D";
          m(268) := x"02A0";
          m(269) := x"FA89";
          m(270) := x"FBA7";
          m(271) := x"F90A";
          m(272) := x"FC2A";
          m(273) := x"FF06";
          m(274) := x"FDE8";
          m(275) := x"FCF3";
          m(276) := x"FC9F";
          m(277) := x"FF8C";
          m(278) := x"012F";
          m(279) := x"0208";
          m(280) := x"FFE8";
          m(281) := x"001E";
          m(282) := x"FFD1";
          m(283) := x"FE46";
          m(284) := x"FF92";
          m(285) := x"0208";
          m(286) := x"FD25";
          m(287) := x"FDB4";
          m(288) := x"FD8B";
          m(289) := x"FCB8";
          m(290) := x"FD34";
          m(291) := x"FFD2";
          m(292) := x"0007";
          m(293) := x"0201";
          m(294) := x"0813";
          m(295) := x"0680";
          m(296) := x"0262";
          m(297) := x"F997";
          m(298) := x"F892";
          m(299) := x"FB57";
          m(300) := x"FAA8";
          m(301) := x"FF28";
          m(302) := x"FC1C";
          m(303) := x"FBE8";
          m(304) := x"FEEE";
          m(305) := x"025B";
          m(306) := x"FF9F";
          m(307) := x"009C";
          m(308) := x"FFF8";
          m(309) := x"000D";
          m(310) := x"FFDD";
          m(311) := x"003E";
          m(312) := x"004A";
          m(313) := x"00F6";
          m(314) := x"FBC0";
          m(315) := x"001F";
          m(316) := x"FFA0";
          m(317) := x"FEE3";
          m(318) := x"03C7";
          m(319) := x"FF64";
          m(320) := x"00EC";
          m(321) := x"0019";
          m(322) := x"05E8";
          m(323) := x"060B";
          m(324) := x"0723";
          m(325) := x"054A";
          m(326) := x"FDA8";
          m(327) := x"FD21";
          m(328) := x"FBBF";
          m(329) := x"FEE8";
          m(330) := x"FD0D";
          m(331) := x"FBBE";
          m(332) := x"FD26";
          m(333) := x"FD38";
          m(334) := x"FCCC";
          m(335) := x"0030";
          m(336) := x"FFFB";
          m(337) := x"FFF0";
          m(338) := x"0021";
          m(339) := x"0096";
          m(340) := x"FF38";
          m(341) := x"FC18";
          m(342) := x"F9B7";
          m(343) := x"01D8";
          m(344) := x"01FB";
          m(345) := x"FF39";
          m(346) := x"FF87";
          m(347) := x"0312";
          m(348) := x"072B";
          m(349) := x"07D1";
          m(350) := x"0061";
          m(351) := x"080D";
          m(352) := x"058E";
          m(353) := x"0434";
          m(354) := x"0487";
          m(355) := x"FBEB";
          m(356) := x"FD62";
          m(357) := x"FCA1";
          m(358) := x"FB32";
          m(359) := x"FBF8";
          m(360) := x"FE51";
          m(361) := x"FEFF";
          m(362) := x"FFEC";
          m(363) := x"005B";
          m(364) := x"0011";
          m(365) := x"0008";
          m(366) := x"0043";
          m(367) := x"00A5";
          m(368) := x"000E";
          m(369) := x"FE6E";
          m(370) := x"00B5";
          m(371) := x"07A2";
          m(372) := x"03DC";
          m(373) := x"00B9";
          m(374) := x"025E";
          m(375) := x"0231";
          m(376) := x"0978";
          m(377) := x"0289";
          m(378) := x"03CE";
          m(379) := x"062E";
          m(380) := x"078B";
          m(381) := x"0576";
          m(382) := x"0566";
          m(383) := x"FEC8";
          m(384) := x"FF54";
          m(385) := x"FF65";
          m(386) := x"FBBF";
          m(387) := x"FC73";
          m(388) := x"FE88";
          m(389) := x"0116";
          m(390) := x"FF5C";
          m(391) := x"FFA2";
          m(392) := x"000C";
          m(393) := x"FFEF";
          m(394) := x"0013";
          m(395) := x"FFDF";
          m(396) := x"004B";
          m(397) := x"FFBE";
          m(398) := x"FE0D";
          m(399) := x"0186";
          m(400) := x"01E8";
          m(401) := x"021C";
          m(402) := x"06A2";
          m(403) := x"0665";
          m(404) := x"0588";
          m(405) := x"0211";
          m(406) := x"FF75";
          m(407) := x"02FF";
          m(408) := x"0518";
          m(409) := x"0675";
          m(410) := x"0714";
          m(411) := x"028C";
          m(412) := x"FE35";
          m(413) := x"0131";
          m(414) := x"0133";
          m(415) := x"007B";
          m(416) := x"FE96";
          m(417) := x"0084";
          m(418) := x"FF5B";
          m(419) := x"FFE9";
          m(420) := x"FFF6";
          m(421) := x"FFED";
          m(422) := x"004C";
          m(423) := x"FF19";
          m(424) := x"008E";
          m(425) := x"FDB2";
          m(426) := x"FC6D";
          m(427) := x"FEC1";
          m(428) := x"FEC5";
          m(429) := x"FFC8";
          m(430) := x"0554";
          m(431) := x"038E";
          m(432) := x"FFDB";
          m(433) := x"FF9B";
          m(434) := x"FD74";
          m(435) := x"03D5";
          m(436) := x"06B9";
          m(437) := x"0BF0";
          m(438) := x"05CC";
          m(439) := x"FB47";
          m(440) := x"FB98";
          m(441) := x"00E8";
          m(442) := x"01E0";
          m(443) := x"022D";
          m(444) := x"FF4E";
          m(445) := x"FE46";
          m(446) := x"FF44";
          m(447) := x"0012";
          m(448) := x"002E";
          m(449) := x"0008";
          m(450) := x"FFF4";
          m(451) := x"FEDC";
          m(452) := x"00E6";
          m(453) := x"FCB9";
          m(454) := x"FB72";
          m(455) := x"FDFF";
          m(456) := x"02F2";
          m(457) := x"FE21";
          m(458) := x"033E";
          m(459) := x"049F";
          m(460) := x"FB68";
          m(461) := x"025B";
          m(462) := x"FBED";
          m(463) := x"FD82";
          m(464) := x"07AB";
          m(465) := x"03F9";
          m(466) := x"009C";
          m(467) := x"FC97";
          m(468) := x"0084";
          m(469) := x"FF63";
          m(470) := x"FC0C";
          m(471) := x"FF30";
          m(472) := x"FC1D";
          m(473) := x"FC6D";
          m(474) := x"FE4E";
          m(475) := x"001E";
          m(476) := x"0035";
          m(477) := x"0019";
          m(478) := x"FFCE";
          m(479) := x"FF28";
          m(480) := x"001F";
          m(481) := x"FC87";
          m(482) := x"FC47";
          m(483) := x"FAE3";
          m(484) := x"FFE0";
          m(485) := x"0059";
          m(486) := x"0948";
          m(487) := x"014F";
          m(488) := x"FC09";
          m(489) := x"04C8";
          m(490) := x"0231";
          m(491) := x"0203";
          m(492) := x"06B7";
          m(493) := x"FF9A";
          m(494) := x"FE60";
          m(495) := x"FCB7";
          m(496) := x"FE22";
          m(497) := x"F9FF";
          m(498) := x"FA79";
          m(499) := x"FDED";
          m(500) := x"FD24";
          m(501) := x"FDCE";
          m(502) := x"FFCC";
          m(503) := x"FFFC";
          m(504) := x"FFE1";
          m(505) := x"FFD2";
          m(506) := x"FFFF";
          m(507) := x"FF54";
          m(508) := x"009C";
          m(509) := x"FD81";
          m(510) := x"FC44";
          m(511) := x"F8DE";
          m(512) := x"F992";
          m(513) := x"F8F5";
          m(514) := x"FE68";
          m(515) := x"FF9C";
          m(516) := x"FA77";
          m(517) := x"039B";
          m(518) := x"0452";
          m(519) := x"013D";
          m(520) := x"FA02";
          m(521) := x"FDA6";
          m(522) := x"F580";
          m(523) := x"F823";
          m(524) := x"F6E0";
          m(525) := x"F727";
          m(526) := x"F7BC";
          m(527) := x"FAB9";
          m(528) := x"FD55";
          m(529) := x"FF38";
          m(530) := x"00CB";
          m(531) := x"006D";
          m(532) := x"0000";
          m(533) := x"001E";
          m(534) := x"FFD3";
          m(535) := x"FFD6";
          m(536) := x"00BE";
          m(537) := x"FF1C";
          m(538) := x"FB91";
          m(539) := x"F818";
          m(540) := x"F6D4";
          m(541) := x"F6A1";
          m(542) := x"F5FF";
          m(543) := x"FB61";
          m(544) := x"00D0";
          m(545) := x"0134";
          m(546) := x"0312";
          m(547) := x"FC5B";
          m(548) := x"F589";
          m(549) := x"F4D0";
          m(550) := x"F40B";
          m(551) := x"F9EA";
          m(552) := x"F6F6";
          m(553) := x"F72C";
          m(554) := x"F69D";
          m(555) := x"F908";
          m(556) := x"FCF6";
          m(557) := x"FFE5";
          m(558) := x"0040";
          m(559) := x"0024";
          m(560) := x"0012";
          m(561) := x"0022";
          m(562) := x"FFCD";
          m(563) := x"FF24";
          m(564) := x"FEFE";
          m(565) := x"FD98";
          m(566) := x"FA1B";
          m(567) := x"F837";
          m(568) := x"F887";
          m(569) := x"F652";
          m(570) := x"F685";
          m(571) := x"FD5E";
          m(572) := x"00A1";
          m(573) := x"FBC2";
          m(574) := x"0237";
          m(575) := x"FB52";
          m(576) := x"FC86";
          m(577) := x"F82D";
          m(578) := x"FB45";
          m(579) := x"F687";
          m(580) := x"F76E";
          m(581) := x"F8D7";
          m(582) := x"FB53";
          m(583) := x"FC1E";
          m(584) := x"FE4F";
          m(585) := x"0039";
          m(586) := x"0017";
          m(587) := x"000A";
          m(588) := x"FFF8";
          m(589) := x"FFF9";
          m(590) := x"FFCE";
          m(591) := x"FEAD";
          m(592) := x"FECC";
          m(593) := x"F9D3";
          m(594) := x"F89E";
          m(595) := x"F7D6";
          m(596) := x"FBD5";
          m(597) := x"FDEE";
          m(598) := x"FF5D";
          m(599) := x"FF9E";
          m(600) := x"033D";
          m(601) := x"FA96";
          m(602) := x"FACF";
          m(603) := x"F7BE";
          m(604) := x"FBD0";
          m(605) := x"FB52";
          m(606) := x"FE4E";
          m(607) := x"FB99";
          m(608) := x"FC59";
          m(609) := x"FBEC";
          m(610) := x"FD26";
          m(611) := x"FDB6";
          m(612) := x"FE50";
          m(613) := x"0039";
          m(614) := x"FFE2";
          m(615) := x"FFD9";
          m(616) := x"000A";
          m(617) := x"FFD6";
          m(618) := x"0010";
          m(619) := x"FF4E";
          m(620) := x"FD4C";
          m(621) := x"F6E9";
          m(622) := x"F718";
          m(623) := x"F9FF";
          m(624) := x"FFF5";
          m(625) := x"FF7F";
          m(626) := x"0579";
          m(627) := x"F93C";
          m(628) := x"FCD7";
          m(629) := x"FE1A";
          m(630) := x"003D";
          m(631) := x"033F";
          m(632) := x"0158";
          m(633) := x"012C";
          m(634) := x"0053";
          m(635) := x"FF7D";
          m(636) := x"FE23";
          m(637) := x"FE6E";
          m(638) := x"FD3F";
          m(639) := x"FDC2";
          m(640) := x"FEA0";
          m(641) := x"0072";
          m(642) := x"002B";
          m(643) := x"000C";
          m(644) := x"FFF0";
          m(645) := x"FFDB";
          m(646) := x"FF36";
          m(647) := x"FF77";
          m(648) := x"FC28";
          m(649) := x"F65E";
          m(650) := x"F655";
          m(651) := x"F9EC";
          m(652) := x"0044";
          m(653) := x"01F0";
          m(654) := x"0822";
          m(655) := x"00EC";
          m(656) := x"024F";
          m(657) := x"FF27";
          m(658) := x"FE7F";
          m(659) := x"FC6A";
          m(660) := x"FB14";
          m(661) := x"0104";
          m(662) := x"0001";
          m(663) := x"FE25";
          m(664) := x"FD84";
          m(665) := x"00E1";
          m(666) := x"FC62";
          m(667) := x"FD7B";
          m(668) := x"FF44";
          m(669) := x"002B";
          m(670) := x"0012";
          m(671) := x"001A";
          m(672) := x"001A";
          m(673) := x"0016";
          m(674) := x"FFE3";
          m(675) := x"FFBA";
          m(676) := x"FD78";
          m(677) := x"FB03";
          m(678) := x"F8FE";
          m(679) := x"FA27";
          m(680) := x"00CC";
          m(681) := x"0024";
          m(682) := x"0065";
          m(683) := x"FC58";
          m(684) := x"F718";
          m(685) := x"FEE2";
          m(686) := x"FE5A";
          m(687) := x"01F3";
          m(688) := x"FBEF";
          m(689) := x"FF54";
          m(690) := x"FD4E";
          m(691) := x"FDAA";
          m(692) := x"00C5";
          m(693) := x"FEC9";
          m(694) := x"FBAD";
          m(695) := x"FE0C";
          m(696) := x"FF35";
          m(697) := x"FFFC";
          m(698) := x"FFF2";
          m(699) := x"002C";
          m(700) := x"FFFC";
          m(701) := x"FFF4";
          m(702) := x"FFC0";
          m(703) := x"FFBB";
          m(704) := x"FF9B";
          m(705) := x"FF1C";
          m(706) := x"FE0F";
          m(707) := x"FD2B";
          m(708) := x"FFAF";
          m(709) := x"FF10";
          m(710) := x"FCCF";
          m(711) := x"FE8B";
          m(712) := x"FCBF";
          m(713) := x"FEAF";
          m(714) := x"0186";
          m(715) := x"FD5D";
          m(716) := x"FC4E";
          m(717) := x"012D";
          m(718) := x"FC83";
          m(719) := x"FA27";
          m(720) := x"FDE3";
          m(721) := x"FBE1";
          m(722) := x"FD11";
          m(723) := x"FE2E";
          m(724) := x"FF13";
          m(725) := x"FFDB";
          m(726) := x"002F";
          m(727) := x"FFBB";
          m(728) := x"FFE2";
          m(729) := x"FFF3";
          m(730) := x"FFE9";
          m(731) := x"0029";
          m(732) := x"003D";
          m(733) := x"0060";
          m(734) := x"00AC";
          m(735) := x"002F";
          m(736) := x"00C0";
          m(737) := x"016A";
          m(738) := x"005C";
          m(739) := x"0060";
          m(740) := x"01B1";
          m(741) := x"011C";
          m(742) := x"0346";
          m(743) := x"00A6";
          m(744) := x"FEB9";
          m(745) := x"FDCE";
          m(746) := x"FD7A";
          m(747) := x"FE00";
          m(748) := x"FDB6";
          m(749) := x"FD5C";
          m(750) := x"FF1D";
          m(751) := x"FFDF";
          m(752) := x"FFF9";
          m(753) := x"002A";
          m(754) := x"FFFF";
          m(755) := x"0009";
          m(756) := x"002B";
          m(757) := x"FFCC";
          m(758) := x"0015";
          m(759) := x"000B";
          m(760) := x"002B";
          m(761) := x"FFD8";
          m(762) := x"FFFB";
          m(763) := x"0015";
          m(764) := x"0001";
          m(765) := x"002A";
          m(766) := x"0031";
          m(767) := x"001B";
          m(768) := x"0029";
          m(769) := x"FFFB";
          m(770) := x"0015";
          m(771) := x"0003";
          m(772) := x"FFFB";
          m(773) := x"0019";
          m(774) := x"0015";
          m(775) := x"0017";
          m(776) := x"FFF7";
          m(777) := x"005A";
          m(778) := x"0045";
          m(779) := x"FFF1";
          m(780) := x"001D";
          m(781) := x"FFC2";
          m(782) := x"FFE3";
          m(783) := x"0005";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_13.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 13) then
          m(0) := x"0021";
          m(1) := x"FFF8";
          m(2) := x"FFC5";
          m(3) := x"000C";
          m(4) := x"FFE3";
          m(5) := x"0003";
          m(6) := x"0020";
          m(7) := x"0009";
          m(8) := x"FFE4";
          m(9) := x"FFAF";
          m(10) := x"0059";
          m(11) := x"FFD2";
          m(12) := x"FFDC";
          m(13) := x"FFF0";
          m(14) := x"FFF4";
          m(15) := x"FFF5";
          m(16) := x"FFFD";
          m(17) := x"FFF3";
          m(18) := x"002A";
          m(19) := x"FFF5";
          m(20) := x"FFE7";
          m(21) := x"FFE2";
          m(22) := x"FFFC";
          m(23) := x"0007";
          m(24) := x"FFE9";
          m(25) := x"0000";
          m(26) := x"FFE2";
          m(27) := x"FFDB";
          m(28) := x"000B";
          m(29) := x"001E";
          m(30) := x"0018";
          m(31) := x"FFF7";
          m(32) := x"FFFE";
          m(33) := x"0029";
          m(34) := x"0025";
          m(35) := x"FFFF";
          m(36) := x"0026";
          m(37) := x"FFFE";
          m(38) := x"003E";
          m(39) := x"0029";
          m(40) := x"003A";
          m(41) := x"0053";
          m(42) := x"FFF1";
          m(43) := x"FFD4";
          m(44) := x"0010";
          m(45) := x"0026";
          m(46) := x"0009";
          m(47) := x"0039";
          m(48) := x"002A";
          m(49) := x"0026";
          m(50) := x"0037";
          m(51) := x"006E";
          m(52) := x"FFFF";
          m(53) := x"FFF9";
          m(54) := x"0018";
          m(55) := x"000E";
          m(56) := x"FFE8";
          m(57) := x"005F";
          m(58) := x"FFF1";
          m(59) := x"000F";
          m(60) := x"FFEA";
          m(61) := x"0003";
          m(62) := x"0029";
          m(63) := x"00CD";
          m(64) := x"00F1";
          m(65) := x"0116";
          m(66) := x"01AC";
          m(67) := x"022A";
          m(68) := x"02F9";
          m(69) := x"03AE";
          m(70) := x"0396";
          m(71) := x"020C";
          m(72) := x"020F";
          m(73) := x"0127";
          m(74) := x"0000";
          m(75) := x"FFE8";
          m(76) := x"0008";
          m(77) := x"001E";
          m(78) := x"00AC";
          m(79) := x"0022";
          m(80) := x"001D";
          m(81) := x"FFEF";
          m(82) := x"0025";
          m(83) := x"001D";
          m(84) := x"FFF6";
          m(85) := x"FFF0";
          m(86) := x"0016";
          m(87) := x"FFDC";
          m(88) := x"FFFB";
          m(89) := x"001C";
          m(90) := x"01DD";
          m(91) := x"02C8";
          m(92) := x"02BD";
          m(93) := x"0345";
          m(94) := x"039F";
          m(95) := x"0336";
          m(96) := x"0780";
          m(97) := x"09FE";
          m(98) := x"0A0B";
          m(99) := x"0410";
          m(100) := x"03A8";
          m(101) := x"0494";
          m(102) := x"01D7";
          m(103) := x"01A4";
          m(104) := x"01B3";
          m(105) := x"0081";
          m(106) := x"019C";
          m(107) := x"0121";
          m(108) := x"0121";
          m(109) := x"008C";
          m(110) := x"0061";
          m(111) := x"FFEA";
          m(112) := x"FFD4";
          m(113) := x"FFD5";
          m(114) := x"FFCC";
          m(115) := x"FFEC";
          m(116) := x"FFCB";
          m(117) := x"FFE6";
          m(118) := x"0204";
          m(119) := x"02AE";
          m(120) := x"0182";
          m(121) := x"04A5";
          m(122) := x"045C";
          m(123) := x"0076";
          m(124) := x"021B";
          m(125) := x"003F";
          m(126) := x"0398";
          m(127) := x"047B";
          m(128) := x"FD84";
          m(129) := x"004C";
          m(130) := x"FE4C";
          m(131) := x"FFA4";
          m(132) := x"FDD6";
          m(133) := x"FFAC";
          m(134) := x"0421";
          m(135) := x"01F5";
          m(136) := x"01C6";
          m(137) := x"00F9";
          m(138) := x"FFC3";
          m(139) := x"0085";
          m(140) := x"FFD7";
          m(141) := x"0029";
          m(142) := x"FFF6";
          m(143) := x"FFF3";
          m(144) := x"0000";
          m(145) := x"FE8E";
          m(146) := x"FFC1";
          m(147) := x"FED8";
          m(148) := x"FE88";
          m(149) := x"0180";
          m(150) := x"034B";
          m(151) := x"FEA1";
          m(152) := x"FBC5";
          m(153) := x"FD54";
          m(154) := x"0007";
          m(155) := x"01D7";
          m(156) := x"FC42";
          m(157) := x"F9B9";
          m(158) := x"04D0";
          m(159) := x"01E9";
          m(160) := x"FEE7";
          m(161) := x"009C";
          m(162) := x"0018";
          m(163) := x"04A9";
          m(164) := x"0301";
          m(165) := x"00E0";
          m(166) := x"00DB";
          m(167) := x"0071";
          m(168) := x"FFF2";
          m(169) := x"002C";
          m(170) := x"003B";
          m(171) := x"FF5F";
          m(172) := x"FF65";
          m(173) := x"FE0D";
          m(174) := x"FE79";
          m(175) := x"FC8F";
          m(176) := x"FBD0";
          m(177) := x"FF1B";
          m(178) := x"FF7D";
          m(179) := x"FAF0";
          m(180) := x"FEB0";
          m(181) := x"FBB3";
          m(182) := x"0287";
          m(183) := x"0256";
          m(184) := x"04EE";
          m(185) := x"01D5";
          m(186) := x"0657";
          m(187) := x"000C";
          m(188) := x"0282";
          m(189) := x"01F3";
          m(190) := x"FFE9";
          m(191) := x"FD38";
          m(192) := x"0009";
          m(193) := x"FFEE";
          m(194) := x"FFD9";
          m(195) := x"0039";
          m(196) := x"FFE4";
          m(197) := x"FFEF";
          m(198) := x"FF97";
          m(199) := x"FED3";
          m(200) := x"FF28";
          m(201) := x"0326";
          m(202) := x"0088";
          m(203) := x"0097";
          m(204) := x"FF54";
          m(205) := x"FE87";
          m(206) := x"0006";
          m(207) := x"025A";
          m(208) := x"FC2C";
          m(209) := x"FC52";
          m(210) := x"0904";
          m(211) := x"03CC";
          m(212) := x"FE8B";
          m(213) := x"019F";
          m(214) := x"052D";
          m(215) := x"00F9";
          m(216) := x"FDB9";
          m(217) := x"02E6";
          m(218) := x"0447";
          m(219) := x"FE47";
          m(220) := x"FD4A";
          m(221) := x"0093";
          m(222) := x"FF49";
          m(223) := x"004F";
          m(224) := x"FFFD";
          m(225) := x"FFF2";
          m(226) := x"FFC4";
          m(227) := x"FE8E";
          m(228) := x"00BB";
          m(229) := x"0064";
          m(230) := x"FCCE";
          m(231) := x"FEF5";
          m(232) := x"FF9C";
          m(233) := x"00D6";
          m(234) := x"0193";
          m(235) := x"0096";
          m(236) := x"FEF1";
          m(237) := x"FD26";
          m(238) := x"01DE";
          m(239) := x"FE61";
          m(240) := x"FC60";
          m(241) := x"FEF0";
          m(242) := x"FC8F";
          m(243) := x"FCDC";
          m(244) := x"FB25";
          m(245) := x"FD68";
          m(246) := x"FEFD";
          m(247) := x"FD87";
          m(248) := x"F85D";
          m(249) := x"FC91";
          m(250) := x"FF49";
          m(251) := x"FFD7";
          m(252) := x"FFE6";
          m(253) := x"FFF0";
          m(254) := x"0009";
          m(255) := x"FE72";
          m(256) := x"0047";
          m(257) := x"001E";
          m(258) := x"F87A";
          m(259) := x"FA45";
          m(260) := x"FCD2";
          m(261) := x"FE62";
          m(262) := x"0517";
          m(263) := x"FC2B";
          m(264) := x"FE51";
          m(265) := x"FBE9";
          m(266) := x"FD11";
          m(267) := x"00F0";
          m(268) := x"FFBE";
          m(269) := x"F64F";
          m(270) := x"FEAE";
          m(271) := x"FB8E";
          m(272) := x"FD3A";
          m(273) := x"F9A2";
          m(274) := x"F8F3";
          m(275) := x"FB29";
          m(276) := x"F8C5";
          m(277) := x"FBCD";
          m(278) := x"FECC";
          m(279) := x"000B";
          m(280) := x"0011";
          m(281) := x"FFFC";
          m(282) := x"003A";
          m(283) := x"FE6D";
          m(284) := x"FD98";
          m(285) := x"FDE7";
          m(286) := x"FB0A";
          m(287) := x"FDDD";
          m(288) := x"FF2A";
          m(289) := x"00B0";
          m(290) := x"FF60";
          m(291) := x"FF9A";
          m(292) := x"FD7D";
          m(293) := x"FE6B";
          m(294) := x"0139";
          m(295) := x"01D2";
          m(296) := x"FAF5";
          m(297) := x"FBB2";
          m(298) := x"FEDB";
          m(299) := x"FC9B";
          m(300) := x"FA56";
          m(301) := x"014F";
          m(302) := x"FC3F";
          m(303) := x"FA51";
          m(304) := x"FD53";
          m(305) := x"FCFF";
          m(306) := x"FEDF";
          m(307) := x"0018";
          m(308) := x"0000";
          m(309) := x"0004";
          m(310) := x"0007";
          m(311) := x"FE8E";
          m(312) := x"FBD6";
          m(313) := x"FF2B";
          m(314) := x"FD39";
          m(315) := x"FC93";
          m(316) := x"F962";
          m(317) := x"FA6B";
          m(318) := x"FD90";
          m(319) := x"FEBA";
          m(320) := x"FD4A";
          m(321) := x"FB09";
          m(322) := x"FF85";
          m(323) := x"01FD";
          m(324) := x"0176";
          m(325) := x"FFBE";
          m(326) := x"FF74";
          m(327) := x"FE40";
          m(328) := x"FC3A";
          m(329) := x"02D2";
          m(330) := x"FF31";
          m(331) := x"FC4F";
          m(332) := x"014C";
          m(333) := x"FF0A";
          m(334) := x"FE21";
          m(335) := x"0039";
          m(336) := x"FFE3";
          m(337) := x"FFE2";
          m(338) := x"FFD9";
          m(339) := x"FF62";
          m(340) := x"FBE2";
          m(341) := x"FD90";
          m(342) := x"FBE7";
          m(343) := x"FB99";
          m(344) := x"FAB0";
          m(345) := x"FEE2";
          m(346) := x"FAA3";
          m(347) := x"FC66";
          m(348) := x"FC5B";
          m(349) := x"FA82";
          m(350) := x"FC97";
          m(351) := x"01D2";
          m(352) := x"0172";
          m(353) := x"FE0E";
          m(354) := x"FCD5";
          m(355) := x"FEEB";
          m(356) := x"0086";
          m(357) := x"00BD";
          m(358) := x"FC26";
          m(359) := x"FD86";
          m(360) := x"02A6";
          m(361) := x"FF6E";
          m(362) := x"FE9E";
          m(363) := x"FFF7";
          m(364) := x"FFF5";
          m(365) := x"FFF8";
          m(366) := x"0008";
          m(367) := x"FEF1";
          m(368) := x"FC24";
          m(369) := x"FC4B";
          m(370) := x"FAF5";
          m(371) := x"FBDB";
          m(372) := x"F92D";
          m(373) := x"FAAE";
          m(374) := x"FDD8";
          m(375) := x"FA70";
          m(376) := x"FC65";
          m(377) := x"FA3A";
          m(378) := x"FC3E";
          m(379) := x"F974";
          m(380) := x"0289";
          m(381) := x"FFF7";
          m(382) := x"0174";
          m(383) := x"0454";
          m(384) := x"FB99";
          m(385) := x"FE3B";
          m(386) := x"00B0";
          m(387) := x"0561";
          m(388) := x"0241";
          m(389) := x"FF0A";
          m(390) := x"FF5F";
          m(391) := x"002D";
          m(392) := x"FFDA";
          m(393) := x"FF85";
          m(394) := x"FF7E";
          m(395) := x"FF52";
          m(396) := x"00A0";
          m(397) := x"FBB2";
          m(398) := x"FC23";
          m(399) := x"FBE8";
          m(400) := x"F9B8";
          m(401) := x"F8D8";
          m(402) := x"FB44";
          m(403) := x"FD9C";
          m(404) := x"FD12";
          m(405) := x"FA9C";
          m(406) := x"FB39";
          m(407) := x"FB77";
          m(408) := x"00DF";
          m(409) := x"FC00";
          m(410) := x"0555";
          m(411) := x"00B2";
          m(412) := x"FE9B";
          m(413) := x"FF56";
          m(414) := x"0001";
          m(415) := x"0320";
          m(416) := x"016E";
          m(417) := x"0011";
          m(418) := x"003A";
          m(419) := x"FFD3";
          m(420) := x"FFFA";
          m(421) := x"FF2A";
          m(422) := x"FF53";
          m(423) := x"FF67";
          m(424) := x"037C";
          m(425) := x"0114";
          m(426) := x"FD65";
          m(427) := x"FD68";
          m(428) := x"FC28";
          m(429) := x"F518";
          m(430) := x"F7FA";
          m(431) := x"F886";
          m(432) := x"F7DC";
          m(433) := x"FAC9";
          m(434) := x"F84C";
          m(435) := x"FC1B";
          m(436) := x"FDB2";
          m(437) := x"FCB2";
          m(438) := x"FDDD";
          m(439) := x"FE9D";
          m(440) := x"01D4";
          m(441) := x"FF01";
          m(442) := x"FD20";
          m(443) := x"03B7";
          m(444) := x"0330";
          m(445) := x"0245";
          m(446) := x"018E";
          m(447) := x"002B";
          m(448) := x"000D";
          m(449) := x"FFBE";
          m(450) := x"FEDE";
          m(451) := x"0072";
          m(452) := x"03E9";
          m(453) := x"05AD";
          m(454) := x"041A";
          m(455) := x"05F7";
          m(456) := x"0051";
          m(457) := x"FEBD";
          m(458) := x"FCFB";
          m(459) := x"FD76";
          m(460) := x"F66D";
          m(461) := x"F703";
          m(462) := x"F9A5";
          m(463) := x"FC1A";
          m(464) := x"FD5E";
          m(465) := x"FC4A";
          m(466) := x"019A";
          m(467) := x"07AC";
          m(468) := x"0592";
          m(469) := x"0052";
          m(470) := x"00AD";
          m(471) := x"06B9";
          m(472) := x"0406";
          m(473) := x"03E2";
          m(474) := x"00FF";
          m(475) := x"FFF2";
          m(476) := x"FFE7";
          m(477) := x"FFD6";
          m(478) := x"FF09";
          m(479) := x"FFE8";
          m(480) := x"0526";
          m(481) := x"0978";
          m(482) := x"07D9";
          m(483) := x"0927";
          m(484) := x"0741";
          m(485) := x"0011";
          m(486) := x"06A9";
          m(487) := x"01A5";
          m(488) := x"FDAA";
          m(489) := x"F8BA";
          m(490) := x"FB73";
          m(491) := x"FF38";
          m(492) := x"0156";
          m(493) := x"03A3";
          m(494) := x"046C";
          m(495) := x"086A";
          m(496) := x"035E";
          m(497) := x"FD32";
          m(498) := x"01A0";
          m(499) := x"0410";
          m(500) := x"0243";
          m(501) := x"02EC";
          m(502) := x"0016";
          m(503) := x"005F";
          m(504) := x"0011";
          m(505) := x"0008";
          m(506) := x"FF84";
          m(507) := x"0092";
          m(508) := x"07A1";
          m(509) := x"084D";
          m(510) := x"07AA";
          m(511) := x"0B08";
          m(512) := x"0C79";
          m(513) := x"0BC5";
          m(514) := x"0C78";
          m(515) := x"02F0";
          m(516) := x"052F";
          m(517) := x"FD29";
          m(518) := x"FC86";
          m(519) := x"027A";
          m(520) := x"0572";
          m(521) := x"0C40";
          m(522) := x"06EB";
          m(523) := x"0543";
          m(524) := x"015D";
          m(525) := x"01F5";
          m(526) := x"0487";
          m(527) := x"04AA";
          m(528) := x"0403";
          m(529) := x"0160";
          m(530) := x"FFBC";
          m(531) := x"0034";
          m(532) := x"001B";
          m(533) := x"FFF8";
          m(534) := x"FFC2";
          m(535) := x"02D5";
          m(536) := x"0678";
          m(537) := x"0597";
          m(538) := x"0729";
          m(539) := x"06F7";
          m(540) := x"09AB";
          m(541) := x"08D2";
          m(542) := x"0697";
          m(543) := x"0DF9";
          m(544) := x"0EE5";
          m(545) := x"07AB";
          m(546) := x"066E";
          m(547) := x"FDC8";
          m(548) := x"0339";
          m(549) := x"0408";
          m(550) := x"0184";
          m(551) := x"016F";
          m(552) := x"050A";
          m(553) := x"059D";
          m(554) := x"0470";
          m(555) := x"05C8";
          m(556) := x"034A";
          m(557) := x"FFE2";
          m(558) := x"0024";
          m(559) := x"000A";
          m(560) := x"FFDF";
          m(561) := x"0035";
          m(562) := x"FF9E";
          m(563) := x"0177";
          m(564) := x"0395";
          m(565) := x"04F0";
          m(566) := x"04DB";
          m(567) := x"0023";
          m(568) := x"03B6";
          m(569) := x"02A6";
          m(570) := x"0560";
          m(571) := x"03F3";
          m(572) := x"0B49";
          m(573) := x"05D0";
          m(574) := x"029D";
          m(575) := x"017E";
          m(576) := x"04D3";
          m(577) := x"0252";
          m(578) := x"01BC";
          m(579) := x"02BE";
          m(580) := x"05C5";
          m(581) := x"FE74";
          m(582) := x"FEF8";
          m(583) := x"03C3";
          m(584) := x"01FB";
          m(585) := x"FF5D";
          m(586) := x"003B";
          m(587) := x"000E";
          m(588) := x"FFDB";
          m(589) := x"000B";
          m(590) := x"FFAC";
          m(591) := x"002B";
          m(592) := x"022B";
          m(593) := x"0296";
          m(594) := x"FE06";
          m(595) := x"FF69";
          m(596) := x"0216";
          m(597) := x"00D8";
          m(598) := x"FC8F";
          m(599) := x"FD7D";
          m(600) := x"0568";
          m(601) := x"05F3";
          m(602) := x"07EA";
          m(603) := x"02D5";
          m(604) := x"0022";
          m(605) := x"0487";
          m(606) := x"040B";
          m(607) := x"0535";
          m(608) := x"039A";
          m(609) := x"FF4E";
          m(610) := x"0194";
          m(611) := x"04F3";
          m(612) := x"0099";
          m(613) := x"FFBF";
          m(614) := x"0057";
          m(615) := x"0029";
          m(616) := x"FFE8";
          m(617) := x"FFD9";
          m(618) := x"0005";
          m(619) := x"FF94";
          m(620) := x"FE25";
          m(621) := x"0017";
          m(622) := x"F7D9";
          m(623) := x"FC6C";
          m(624) := x"FD26";
          m(625) := x"011C";
          m(626) := x"FF16";
          m(627) := x"FBA4";
          m(628) := x"FDC3";
          m(629) := x"FE20";
          m(630) := x"04C0";
          m(631) := x"024B";
          m(632) := x"073F";
          m(633) := x"0138";
          m(634) := x"FEDF";
          m(635) := x"FD42";
          m(636) := x"035D";
          m(637) := x"0307";
          m(638) := x"012F";
          m(639) := x"0357";
          m(640) := x"005F";
          m(641) := x"0006";
          m(642) := x"0000";
          m(643) := x"FFF2";
          m(644) := x"002A";
          m(645) := x"0000";
          m(646) := x"0021";
          m(647) := x"FF89";
          m(648) := x"FCA9";
          m(649) := x"FC82";
          m(650) := x"FD61";
          m(651) := x"FBB5";
          m(652) := x"FCFC";
          m(653) := x"FFEE";
          m(654) := x"00A2";
          m(655) := x"FDF5";
          m(656) := x"009C";
          m(657) := x"FFDA";
          m(658) := x"FF89";
          m(659) := x"0175";
          m(660) := x"00F6";
          m(661) := x"01FA";
          m(662) := x"010F";
          m(663) := x"028A";
          m(664) := x"0433";
          m(665) := x"037B";
          m(666) := x"01CA";
          m(667) := x"023C";
          m(668) := x"00C0";
          m(669) := x"0062";
          m(670) := x"002A";
          m(671) := x"0008";
          m(672) := x"FFF9";
          m(673) := x"0017";
          m(674) := x"FF9E";
          m(675) := x"FF74";
          m(676) := x"FE3A";
          m(677) := x"FD60";
          m(678) := x"FDBE";
          m(679) := x"FC41";
          m(680) := x"FF9D";
          m(681) := x"FF15";
          m(682) := x"FB0A";
          m(683) := x"FD5C";
          m(684) := x"050F";
          m(685) := x"032A";
          m(686) := x"0293";
          m(687) := x"0432";
          m(688) := x"06DE";
          m(689) := x"05EC";
          m(690) := x"0337";
          m(691) := x"038C";
          m(692) := x"0439";
          m(693) := x"0236";
          m(694) := x"013A";
          m(695) := x"0180";
          m(696) := x"01FB";
          m(697) := x"01B7";
          m(698) := x"0042";
          m(699) := x"FFE9";
          m(700) := x"0024";
          m(701) := x"0013";
          m(702) := x"FFFB";
          m(703) := x"0006";
          m(704) := x"FFA7";
          m(705) := x"FECF";
          m(706) := x"FEC4";
          m(707) := x"FE47";
          m(708) := x"FBF5";
          m(709) := x"F986";
          m(710) := x"FB6F";
          m(711) := x"FD6C";
          m(712) := x"FDA1";
          m(713) := x"FD33";
          m(714) := x"FFFD";
          m(715) := x"0121";
          m(716) := x"FFA2";
          m(717) := x"0074";
          m(718) := x"FF2E";
          m(719) := x"FD96";
          m(720) := x"FD46";
          m(721) := x"FDF3";
          m(722) := x"FEA3";
          m(723) := x"FF83";
          m(724) := x"FFF9";
          m(725) := x"001A";
          m(726) := x"0044";
          m(727) := x"0019";
          m(728) := x"FFCC";
          m(729) := x"FFE4";
          m(730) := x"000F";
          m(731) := x"0001";
          m(732) := x"FFE1";
          m(733) := x"FF96";
          m(734) := x"FFB1";
          m(735) := x"FF6C";
          m(736) := x"FEE8";
          m(737) := x"FDBE";
          m(738) := x"FF5F";
          m(739) := x"FF3F";
          m(740) := x"FF63";
          m(741) := x"FE6D";
          m(742) := x"FD54";
          m(743) := x"FDAB";
          m(744) := x"FE21";
          m(745) := x"FE2C";
          m(746) := x"FEA1";
          m(747) := x"FF48";
          m(748) := x"FF22";
          m(749) := x"FE3D";
          m(750) := x"FEC6";
          m(751) := x"0012";
          m(752) := x"FFBE";
          m(753) := x"0011";
          m(754) := x"0019";
          m(755) := x"FFD5";
          m(756) := x"000C";
          m(757) := x"000E";
          m(758) := x"002C";
          m(759) := x"FFD9";
          m(760) := x"FFE5";
          m(761) := x"001B";
          m(762) := x"FFEE";
          m(763) := x"000D";
          m(764) := x"FFF9";
          m(765) := x"FFFB";
          m(766) := x"0019";
          m(767) := x"FFAC";
          m(768) := x"FFCE";
          m(769) := x"0006";
          m(770) := x"FFF6";
          m(771) := x"FFDB";
          m(772) := x"FFCF";
          m(773) := x"FFBC";
          m(774) := x"FFBE";
          m(775) := x"FFBE";
          m(776) := x"FFB0";
          m(777) := x"FFA1";
          m(778) := x"FE9F";
          m(779) := x"FFCF";
          m(780) := x"001F";
          m(781) := x"FFF5";
          m(782) := x"0014";
          m(783) := x"0000";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_14.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 14) then
          m(0) := x"FFE8";
          m(1) := x"000E";
          m(2) := x"FFD3";
          m(3) := x"0027";
          m(4) := x"FFEA";
          m(5) := x"FFD9";
          m(6) := x"0016";
          m(7) := x"0009";
          m(8) := x"0000";
          m(9) := x"FFFD";
          m(10) := x"0013";
          m(11) := x"FFF0";
          m(12) := x"FFF2";
          m(13) := x"FFCB";
          m(14) := x"FFE0";
          m(15) := x"0007";
          m(16) := x"000B";
          m(17) := x"001C";
          m(18) := x"0000";
          m(19) := x"0000";
          m(20) := x"000F";
          m(21) := x"FFE2";
          m(22) := x"001F";
          m(23) := x"FFEC";
          m(24) := x"FFE0";
          m(25) := x"0002";
          m(26) := x"FFC3";
          m(27) := x"0010";
          m(28) := x"FFF8";
          m(29) := x"0019";
          m(30) := x"FFCE";
          m(31) := x"FFBD";
          m(32) := x"FFF2";
          m(33) := x"FFE1";
          m(34) := x"002E";
          m(35) := x"0051";
          m(36) := x"005F";
          m(37) := x"0025";
          m(38) := x"001A";
          m(39) := x"00AB";
          m(40) := x"0101";
          m(41) := x"00C5";
          m(42) := x"FFCF";
          m(43) := x"0025";
          m(44) := x"00FB";
          m(45) := x"00BA";
          m(46) := x"001F";
          m(47) := x"0016";
          m(48) := x"0019";
          m(49) := x"0002";
          m(50) := x"0037";
          m(51) := x"FFF5";
          m(52) := x"FFEC";
          m(53) := x"FFD6";
          m(54) := x"FFDC";
          m(55) := x"FFD3";
          m(56) := x"000E";
          m(57) := x"0036";
          m(58) := x"000A";
          m(59) := x"0018";
          m(60) := x"FFFF";
          m(61) := x"001D";
          m(62) := x"0072";
          m(63) := x"004F";
          m(64) := x"0093";
          m(65) := x"0053";
          m(66) := x"0079";
          m(67) := x"01A2";
          m(68) := x"0157";
          m(69) := x"00A3";
          m(70) := x"0169";
          m(71) := x"0151";
          m(72) := x"0280";
          m(73) := x"0353";
          m(74) := x"0279";
          m(75) := x"01A0";
          m(76) := x"00DA";
          m(77) := x"0052";
          m(78) := x"001D";
          m(79) := x"FFF1";
          m(80) := x"FF9E";
          m(81) := x"FFB7";
          m(82) := x"000F";
          m(83) := x"FFCD";
          m(84) := x"001F";
          m(85) := x"0034";
          m(86) := x"0010";
          m(87) := x"0008";
          m(88) := x"0010";
          m(89) := x"FF98";
          m(90) := x"FFFD";
          m(91) := x"006A";
          m(92) := x"FFD5";
          m(93) := x"01E5";
          m(94) := x"0230";
          m(95) := x"0157";
          m(96) := x"FE13";
          m(97) := x"FF0B";
          m(98) := x"0502";
          m(99) := x"032C";
          m(100) := x"05F4";
          m(101) := x"07CC";
          m(102) := x"07C2";
          m(103) := x"0427";
          m(104) := x"0166";
          m(105) := x"0176";
          m(106) := x"00BD";
          m(107) := x"006C";
          m(108) := x"FFE9";
          m(109) := x"FFFE";
          m(110) := x"0010";
          m(111) := x"002B";
          m(112) := x"0002";
          m(113) := x"FFF7";
          m(114) := x"000D";
          m(115) := x"FFF0";
          m(116) := x"0008";
          m(117) := x"FF10";
          m(118) := x"0103";
          m(119) := x"00D6";
          m(120) := x"F986";
          m(121) := x"FF16";
          m(122) := x"FD4E";
          m(123) := x"FEF3";
          m(124) := x"FBCA";
          m(125) := x"FE04";
          m(126) := x"0303";
          m(127) := x"FF3A";
          m(128) := x"0575";
          m(129) := x"09BD";
          m(130) := x"066B";
          m(131) := x"09B8";
          m(132) := x"07F8";
          m(133) := x"0388";
          m(134) := x"02E9";
          m(135) := x"0101";
          m(136) := x"0035";
          m(137) := x"0000";
          m(138) := x"FFEA";
          m(139) := x"0028";
          m(140) := x"FFF7";
          m(141) := x"FFE2";
          m(142) := x"FFF7";
          m(143) := x"FF22";
          m(144) := x"FC8B";
          m(145) := x"FC0D";
          m(146) := x"FE3F";
          m(147) := x"F952";
          m(148) := x"FD33";
          m(149) := x"FD9A";
          m(150) := x"FF22";
          m(151) := x"FB64";
          m(152) := x"FB14";
          m(153) := x"0018";
          m(154) := x"FE92";
          m(155) := x"FF00";
          m(156) := x"FF9E";
          m(157) := x"03AB";
          m(158) := x"0547";
          m(159) := x"08F6";
          m(160) := x"0D67";
          m(161) := x"072F";
          m(162) := x"0461";
          m(163) := x"0267";
          m(164) := x"0005";
          m(165) := x"FFDC";
          m(166) := x"FFD3";
          m(167) := x"001B";
          m(168) := x"003A";
          m(169) := x"000E";
          m(170) := x"0054";
          m(171) := x"FE6C";
          m(172) := x"FB8C";
          m(173) := x"FC71";
          m(174) := x"F65E";
          m(175) := x"FD60";
          m(176) := x"020C";
          m(177) := x"FE33";
          m(178) := x"009A";
          m(179) := x"0123";
          m(180) := x"02BA";
          m(181) := x"004D";
          m(182) := x"FCE1";
          m(183) := x"0233";
          m(184) := x"FE8D";
          m(185) := x"055F";
          m(186) := x"03BE";
          m(187) := x"0899";
          m(188) := x"065D";
          m(189) := x"05E4";
          m(190) := x"04BB";
          m(191) := x"02A5";
          m(192) := x"0135";
          m(193) := x"001D";
          m(194) := x"FFE5";
          m(195) := x"FFF5";
          m(196) := x"002E";
          m(197) := x"FFCC";
          m(198) := x"FFCF";
          m(199) := x"FD46";
          m(200) := x"F921";
          m(201) := x"FE42";
          m(202) := x"F85F";
          m(203) := x"FA1C";
          m(204) := x"058C";
          m(205) := x"060A";
          m(206) := x"063F";
          m(207) := x"04BF";
          m(208) := x"03E9";
          m(209) := x"FDA8";
          m(210) := x"00E4";
          m(211) := x"0141";
          m(212) := x"0093";
          m(213) := x"03AC";
          m(214) := x"0436";
          m(215) := x"087F";
          m(216) := x"08FC";
          m(217) := x"082A";
          m(218) := x"062A";
          m(219) := x"0479";
          m(220) := x"02DF";
          m(221) := x"0116";
          m(222) := x"FFFE";
          m(223) := x"0005";
          m(224) := x"000B";
          m(225) := x"FF7F";
          m(226) := x"FF76";
          m(227) := x"FE9F";
          m(228) := x"FB5C";
          m(229) := x"002F";
          m(230) := x"FE37";
          m(231) := x"0108";
          m(232) := x"0383";
          m(233) := x"FF6E";
          m(234) := x"FB7D";
          m(235) := x"04C3";
          m(236) := x"003D";
          m(237) := x"FC81";
          m(238) := x"00C3";
          m(239) := x"FCC0";
          m(240) := x"FCF3";
          m(241) := x"FF74";
          m(242) := x"05D8";
          m(243) := x"05B1";
          m(244) := x"0B58";
          m(245) := x"085A";
          m(246) := x"08F2";
          m(247) := x"0639";
          m(248) := x"03CA";
          m(249) := x"01C2";
          m(250) := x"FFD4";
          m(251) := x"0012";
          m(252) := x"001D";
          m(253) := x"FF3E";
          m(254) := x"FF48";
          m(255) := x"FE92";
          m(256) := x"FA8A";
          m(257) := x"FA52";
          m(258) := x"FF39";
          m(259) := x"00FB";
          m(260) := x"02A5";
          m(261) := x"020C";
          m(262) := x"052E";
          m(263) := x"0255";
          m(264) := x"FD0A";
          m(265) := x"FA18";
          m(266) := x"F0DA";
          m(267) := x"F266";
          m(268) := x"F8AA";
          m(269) := x"FDF2";
          m(270) := x"046C";
          m(271) := x"05BB";
          m(272) := x"0980";
          m(273) := x"064E";
          m(274) := x"0815";
          m(275) := x"0841";
          m(276) := x"0361";
          m(277) := x"007A";
          m(278) := x"FE74";
          m(279) := x"FE2B";
          m(280) := x"FFEF";
          m(281) := x"FF5D";
          m(282) := x"FFAB";
          m(283) := x"FED1";
          m(284) := x"FC3A";
          m(285) := x"F9D7";
          m(286) := x"0219";
          m(287) := x"05D4";
          m(288) := x"0B75";
          m(289) := x"04A6";
          m(290) := x"0198";
          m(291) := x"FA15";
          m(292) := x"FDF4";
          m(293) := x"F707";
          m(294) := x"F476";
          m(295) := x"F5F1";
          m(296) := x"F702";
          m(297) := x"02A7";
          m(298) := x"0908";
          m(299) := x"049C";
          m(300) := x"0396";
          m(301) := x"03F6";
          m(302) := x"03FA";
          m(303) := x"01DD";
          m(304) := x"035F";
          m(305) := x"FF27";
          m(306) := x"FECB";
          m(307) := x"FF73";
          m(308) := x"FFD2";
          m(309) := x"FFAB";
          m(310) := x"FF1C";
          m(311) := x"FE58";
          m(312) := x"F9C3";
          m(313) := x"FA45";
          m(314) := x"015C";
          m(315) := x"034D";
          m(316) := x"FF82";
          m(317) := x"FC04";
          m(318) := x"FD9C";
          m(319) := x"F85E";
          m(320) := x"F9FF";
          m(321) := x"FA99";
          m(322) := x"F832";
          m(323) := x"F8AB";
          m(324) := x"0A06";
          m(325) := x"0FF1";
          m(326) := x"0C68";
          m(327) := x"0372";
          m(328) := x"013B";
          m(329) := x"0247";
          m(330) := x"FDE7";
          m(331) := x"FFE8";
          m(332) := x"05FC";
          m(333) := x"026C";
          m(334) := x"005F";
          m(335) := x"FFE2";
          m(336) := x"FFED";
          m(337) := x"FFCD";
          m(338) := x"FEEC";
          m(339) := x"FDF1";
          m(340) := x"FBB1";
          m(341) := x"FD89";
          m(342) := x"01A0";
          m(343) := x"027E";
          m(344) := x"FDE5";
          m(345) := x"FBDA";
          m(346) := x"02C6";
          m(347) := x"FF4C";
          m(348) := x"FF95";
          m(349) := x"FCFD";
          m(350) := x"F4A1";
          m(351) := x"FA33";
          m(352) := x"0370";
          m(353) := x"04A5";
          m(354) := x"03C5";
          m(355) := x"FE74";
          m(356) := x"026A";
          m(357) := x"01E9";
          m(358) := x"FDAA";
          m(359) := x"00B8";
          m(360) := x"0070";
          m(361) := x"FF33";
          m(362) := x"0029";
          m(363) := x"FF8E";
          m(364) := x"0001";
          m(365) := x"0016";
          m(366) := x"FF5D";
          m(367) := x"FEEB";
          m(368) := x"FA6E";
          m(369) := x"FEF0";
          m(370) := x"FF93";
          m(371) := x"02CE";
          m(372) := x"0447";
          m(373) := x"045F";
          m(374) := x"022A";
          m(375) := x"FBED";
          m(376) := x"FFF3";
          m(377) := x"FB55";
          m(378) := x"F840";
          m(379) := x"FEBF";
          m(380) := x"FEA7";
          m(381) := x"04E6";
          m(382) := x"FC5D";
          m(383) := x"021C";
          m(384) := x"FE07";
          m(385) := x"FD98";
          m(386) := x"0086";
          m(387) := x"FE21";
          m(388) := x"FC4C";
          m(389) := x"FE22";
          m(390) := x"FFCA";
          m(391) := x"FFA5";
          m(392) := x"FFD6";
          m(393) := x"FFD7";
          m(394) := x"FFC2";
          m(395) := x"FFD3";
          m(396) := x"FFB9";
          m(397) := x"FFC5";
          m(398) := x"0339";
          m(399) := x"08C6";
          m(400) := x"02AA";
          m(401) := x"056A";
          m(402) := x"0576";
          m(403) := x"01B0";
          m(404) := x"0024";
          m(405) := x"00C8";
          m(406) := x"FA33";
          m(407) := x"FBB2";
          m(408) := x"008D";
          m(409) := x"04CE";
          m(410) := x"FFF3";
          m(411) := x"F562";
          m(412) := x"0004";
          m(413) := x"F756";
          m(414) := x"FE14";
          m(415) := x"FA91";
          m(416) := x"0006";
          m(417) := x"FF79";
          m(418) := x"FEBA";
          m(419) := x"0007";
          m(420) := x"FFE7";
          m(421) := x"FFD7";
          m(422) := x"FFA3";
          m(423) := x"0000";
          m(424) := x"0354";
          m(425) := x"0347";
          m(426) := x"01AA";
          m(427) := x"06E0";
          m(428) := x"004D";
          m(429) := x"FF06";
          m(430) := x"017C";
          m(431) := x"FC75";
          m(432) := x"FE27";
          m(433) := x"FD83";
          m(434) := x"FC59";
          m(435) := x"FF89";
          m(436) := x"023C";
          m(437) := x"FDDF";
          m(438) := x"FF6C";
          m(439) := x"FBE9";
          m(440) := x"FF2E";
          m(441) := x"FDC9";
          m(442) := x"FC28";
          m(443) := x"02A2";
          m(444) := x"0015";
          m(445) := x"0088";
          m(446) := x"FF96";
          m(447) := x"FFE0";
          m(448) := x"0011";
          m(449) := x"0036";
          m(450) := x"FFC0";
          m(451) := x"00AB";
          m(452) := x"02F5";
          m(453) := x"0686";
          m(454) := x"00ED";
          m(455) := x"FB65";
          m(456) := x"FCC2";
          m(457) := x"FEB3";
          m(458) := x"FE95";
          m(459) := x"03CE";
          m(460) := x"0328";
          m(461) := x"FD05";
          m(462) := x"FCF9";
          m(463) := x"0127";
          m(464) := x"FE62";
          m(465) := x"03E8";
          m(466) := x"FEF6";
          m(467) := x"FF99";
          m(468) := x"FC24";
          m(469) := x"FABA";
          m(470) := x"FD6F";
          m(471) := x"00B3";
          m(472) := x"FE8A";
          m(473) := x"010B";
          m(474) := x"FF82";
          m(475) := x"FFFF";
          m(476) := x"FFF9";
          m(477) := x"0007";
          m(478) := x"0010";
          m(479) := x"00FA";
          m(480) := x"0150";
          m(481) := x"0284";
          m(482) := x"FF7E";
          m(483) := x"FE68";
          m(484) := x"0390";
          m(485) := x"0128";
          m(486) := x"01DA";
          m(487) := x"02E9";
          m(488) := x"FFDF";
          m(489) := x"FC76";
          m(490) := x"FCF2";
          m(491) := x"0045";
          m(492) := x"018C";
          m(493) := x"FE3F";
          m(494) := x"02D6";
          m(495) := x"FCF1";
          m(496) := x"FDBC";
          m(497) := x"F780";
          m(498) := x"FAB5";
          m(499) := x"FED0";
          m(500) := x"FD0D";
          m(501) := x"FF2E";
          m(502) := x"FF25";
          m(503) := x"008E";
          m(504) := x"0018";
          m(505) := x"FFD9";
          m(506) := x"FFE9";
          m(507) := x"002A";
          m(508) := x"FF66";
          m(509) := x"FFCD";
          m(510) := x"FED5";
          m(511) := x"0158";
          m(512) := x"FDB2";
          m(513) := x"FE62";
          m(514) := x"02BF";
          m(515) := x"FF90";
          m(516) := x"02A9";
          m(517) := x"000A";
          m(518) := x"04A9";
          m(519) := x"0479";
          m(520) := x"02B3";
          m(521) := x"FDB5";
          m(522) := x"018B";
          m(523) := x"FE01";
          m(524) := x"FD69";
          m(525) := x"FB52";
          m(526) := x"FCD0";
          m(527) := x"FEA0";
          m(528) := x"FDD1";
          m(529) := x"FECE";
          m(530) := x"FF73";
          m(531) := x"FFC9";
          m(532) := x"FFD6";
          m(533) := x"FFF8";
          m(534) := x"012F";
          m(535) := x"01FE";
          m(536) := x"FF5F";
          m(537) := x"FF2F";
          m(538) := x"FF4B";
          m(539) := x"01AA";
          m(540) := x"028C";
          m(541) := x"0198";
          m(542) := x"033D";
          m(543) := x"016C";
          m(544) := x"0030";
          m(545) := x"03C0";
          m(546) := x"0050";
          m(547) := x"00A2";
          m(548) := x"FEFC";
          m(549) := x"00DE";
          m(550) := x"FE2E";
          m(551) := x"FECE";
          m(552) := x"00B7";
          m(553) := x"0560";
          m(554) := x"00D8";
          m(555) := x"FE8A";
          m(556) := x"FBA1";
          m(557) := x"FEE5";
          m(558) := x"FFD7";
          m(559) := x"FFE3";
          m(560) := x"FFE6";
          m(561) := x"0011";
          m(562) := x"0124";
          m(563) := x"0247";
          m(564) := x"0185";
          m(565) := x"018D";
          m(566) := x"FF8D";
          m(567) := x"FC76";
          m(568) := x"036E";
          m(569) := x"FCF2";
          m(570) := x"FF1B";
          m(571) := x"0149";
          m(572) := x"01B1";
          m(573) := x"0229";
          m(574) := x"021A";
          m(575) := x"FCF7";
          m(576) := x"FEAE";
          m(577) := x"FD49";
          m(578) := x"FD84";
          m(579) := x"00F3";
          m(580) := x"FC31";
          m(581) := x"01FE";
          m(582) := x"00EF";
          m(583) := x"FB8C";
          m(584) := x"FBAA";
          m(585) := x"FF62";
          m(586) := x"0019";
          m(587) := x"FF99";
          m(588) := x"0011";
          m(589) := x"FFE5";
          m(590) := x"0003";
          m(591) := x"0085";
          m(592) := x"017F";
          m(593) := x"06BA";
          m(594) := x"0416";
          m(595) := x"0473";
          m(596) := x"0269";
          m(597) := x"FF5C";
          m(598) := x"01E5";
          m(599) := x"03F9";
          m(600) := x"FF9F";
          m(601) := x"07E5";
          m(602) := x"02E6";
          m(603) := x"FEDE";
          m(604) := x"FE81";
          m(605) := x"04C8";
          m(606) := x"0208";
          m(607) := x"FFCD";
          m(608) := x"0141";
          m(609) := x"04C7";
          m(610) := x"0097";
          m(611) := x"FE3A";
          m(612) := x"FFC6";
          m(613) := x"FFE3";
          m(614) := x"0016";
          m(615) := x"0023";
          m(616) := x"0005";
          m(617) := x"0015";
          m(618) := x"002B";
          m(619) := x"FFC6";
          m(620) := x"FE60";
          m(621) := x"0205";
          m(622) := x"02CC";
          m(623) := x"0114";
          m(624) := x"0150";
          m(625) := x"FF93";
          m(626) := x"02C4";
          m(627) := x"FF40";
          m(628) := x"FC66";
          m(629) := x"0406";
          m(630) := x"064D";
          m(631) := x"009E";
          m(632) := x"0144";
          m(633) := x"0492";
          m(634) := x"FEBD";
          m(635) := x"FBAC";
          m(636) := x"FE77";
          m(637) := x"0440";
          m(638) := x"005E";
          m(639) := x"0257";
          m(640) := x"0101";
          m(641) := x"0026";
          m(642) := x"0014";
          m(643) := x"FFDD";
          m(644) := x"FFF2";
          m(645) := x"FFFB";
          m(646) := x"FFE4";
          m(647) := x"FFE8";
          m(648) := x"FE90";
          m(649) := x"FEAC";
          m(650) := x"FF32";
          m(651) := x"FF67";
          m(652) := x"0016";
          m(653) := x"FBD2";
          m(654) := x"FF4A";
          m(655) := x"FC6C";
          m(656) := x"FEA7";
          m(657) := x"FE2B";
          m(658) := x"FFA3";
          m(659) := x"FE15";
          m(660) := x"04B0";
          m(661) := x"FE0C";
          m(662) := x"FF97";
          m(663) := x"FF5A";
          m(664) := x"0344";
          m(665) := x"039B";
          m(666) := x"0225";
          m(667) := x"044F";
          m(668) := x"01D6";
          m(669) := x"004B";
          m(670) := x"000F";
          m(671) := x"002C";
          m(672) := x"000A";
          m(673) := x"0000";
          m(674) := x"0042";
          m(675) := x"0008";
          m(676) := x"FF21";
          m(677) := x"FD54";
          m(678) := x"FC60";
          m(679) := x"FF54";
          m(680) := x"0165";
          m(681) := x"FE97";
          m(682) := x"00CB";
          m(683) := x"02A0";
          m(684) := x"05E9";
          m(685) := x"FCC7";
          m(686) := x"FC15";
          m(687) := x"02BD";
          m(688) := x"0233";
          m(689) := x"FEE2";
          m(690) := x"02CB";
          m(691) := x"01A0";
          m(692) := x"03DF";
          m(693) := x"0302";
          m(694) := x"0168";
          m(695) := x"030E";
          m(696) := x"0223";
          m(697) := x"0009";
          m(698) := x"0026";
          m(699) := x"FFD1";
          m(700) := x"0040";
          m(701) := x"0028";
          m(702) := x"0021";
          m(703) := x"0024";
          m(704) := x"FF2A";
          m(705) := x"FE27";
          m(706) := x"FDAC";
          m(707) := x"FE30";
          m(708) := x"FD89";
          m(709) := x"FC91";
          m(710) := x"FBBC";
          m(711) := x"0201";
          m(712) := x"0277";
          m(713) := x"0032";
          m(714) := x"0059";
          m(715) := x"FDAB";
          m(716) := x"FE25";
          m(717) := x"01FB";
          m(718) := x"FC6A";
          m(719) := x"FCED";
          m(720) := x"00B0";
          m(721) := x"01F1";
          m(722) := x"000C";
          m(723) := x"00F6";
          m(724) := x"00BB";
          m(725) := x"0028";
          m(726) := x"0011";
          m(727) := x"FFF0";
          m(728) := x"001F";
          m(729) := x"FFE6";
          m(730) := x"FFE5";
          m(731) := x"000D";
          m(732) := x"0049";
          m(733) := x"FFEE";
          m(734) := x"0033";
          m(735) := x"FFF5";
          m(736) := x"FF27";
          m(737) := x"FF0A";
          m(738) := x"FDA5";
          m(739) := x"FE5F";
          m(740) := x"0241";
          m(741) := x"0239";
          m(742) := x"014F";
          m(743) := x"FF04";
          m(744) := x"FFCD";
          m(745) := x"0204";
          m(746) := x"FFFA";
          m(747) := x"FE79";
          m(748) := x"004E";
          m(749) := x"010C";
          m(750) := x"001D";
          m(751) := x"FFF7";
          m(752) := x"FFC6";
          m(753) := x"0029";
          m(754) := x"002E";
          m(755) := x"FFEC";
          m(756) := x"0017";
          m(757) := x"FFEC";
          m(758) := x"0039";
          m(759) := x"0002";
          m(760) := x"0004";
          m(761) := x"FFED";
          m(762) := x"0078";
          m(763) := x"0106";
          m(764) := x"00B7";
          m(765) := x"0009";
          m(766) := x"FFF5";
          m(767) := x"0012";
          m(768) := x"00A0";
          m(769) := x"FFDF";
          m(770) := x"FFEA";
          m(771) := x"FFBD";
          m(772) := x"0059";
          m(773) := x"FFB1";
          m(774) := x"0003";
          m(775) := x"FFD9";
          m(776) := x"FFCC";
          m(777) := x"001A";
          m(778) := x"0031";
          m(779) := x"0004";
          m(780) := x"003B";
          m(781) := x"FFEB";
          m(782) := x"FFFC";
          m(783) := x"FFF3";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_15.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 15) then
          m(0) := x"FFF3";
          m(1) := x"0006";
          m(2) := x"FFF1";
          m(3) := x"001B";
          m(4) := x"FFF6";
          m(5) := x"FFF9";
          m(6) := x"FFCF";
          m(7) := x"FFD8";
          m(8) := x"FFEB";
          m(9) := x"FFCA";
          m(10) := x"FFE2";
          m(11) := x"0001";
          m(12) := x"FFE8";
          m(13) := x"001B";
          m(14) := x"FFE2";
          m(15) := x"0009";
          m(16) := x"FFD7";
          m(17) := x"FFF9";
          m(18) := x"0003";
          m(19) := x"0020";
          m(20) := x"FFE8";
          m(21) := x"0006";
          m(22) := x"FFFD";
          m(23) := x"0005";
          m(24) := x"0008";
          m(25) := x"003C";
          m(26) := x"FFD0";
          m(27) := x"FFF9";
          m(28) := x"0004";
          m(29) := x"000E";
          m(30) := x"003D";
          m(31) := x"FFF2";
          m(32) := x"0007";
          m(33) := x"000D";
          m(34) := x"0009";
          m(35) := x"FFF4";
          m(36) := x"FFA0";
          m(37) := x"FFD9";
          m(38) := x"FFBD";
          m(39) := x"FFD5";
          m(40) := x"FFA0";
          m(41) := x"FFED";
          m(42) := x"FFEF";
          m(43) := x"FFC1";
          m(44) := x"FF7E";
          m(45) := x"FFB8";
          m(46) := x"FFBF";
          m(47) := x"001F";
          m(48) := x"0025";
          m(49) := x"FFF1";
          m(50) := x"0021";
          m(51) := x"FFD7";
          m(52) := x"0038";
          m(53) := x"0009";
          m(54) := x"FFF1";
          m(55) := x"0013";
          m(56) := x"FFEE";
          m(57) := x"0032";
          m(58) := x"FFE9";
          m(59) := x"FFE1";
          m(60) := x"0024";
          m(61) := x"FFF0";
          m(62) := x"FFCB";
          m(63) := x"FF23";
          m(64) := x"FEC4";
          m(65) := x"FF41";
          m(66) := x"FEBA";
          m(67) := x"FE64";
          m(68) := x"FE7C";
          m(69) := x"FF00";
          m(70) := x"FF60";
          m(71) := x"FECC";
          m(72) := x"FCCF";
          m(73) := x"FCE4";
          m(74) := x"FD9E";
          m(75) := x"FEAE";
          m(76) := x"FEF6";
          m(77) := x"FF91";
          m(78) := x"FFBB";
          m(79) := x"FFBB";
          m(80) := x"FFAC";
          m(81) := x"FFBC";
          m(82) := x"FFE4";
          m(83) := x"0029";
          m(84) := x"000D";
          m(85) := x"005C";
          m(86) := x"0006";
          m(87) := x"FFE4";
          m(88) := x"FFE6";
          m(89) := x"0004";
          m(90) := x"FF0C";
          m(91) := x"FE93";
          m(92) := x"FC8C";
          m(93) := x"FCF5";
          m(94) := x"FCCF";
          m(95) := x"FC74";
          m(96) := x"FB80";
          m(97) := x"FBA1";
          m(98) := x"FC82";
          m(99) := x"F9E5";
          m(100) := x"F6AF";
          m(101) := x"F9AA";
          m(102) := x"FAD8";
          m(103) := x"FEBF";
          m(104) := x"00C4";
          m(105) := x"FF30";
          m(106) := x"FED7";
          m(107) := x"FEF4";
          m(108) := x"FF4D";
          m(109) := x"FFD2";
          m(110) := x"FFD0";
          m(111) := x"FFE4";
          m(112) := x"FFFC";
          m(113) := x"FFCA";
          m(114) := x"0011";
          m(115) := x"FFC7";
          m(116) := x"FF9F";
          m(117) := x"FFDD";
          m(118) := x"FF5B";
          m(119) := x"FD7E";
          m(120) := x"FDB5";
          m(121) := x"FBB2";
          m(122) := x"FB4E";
          m(123) := x"F9E7";
          m(124) := x"FB60";
          m(125) := x"FD8D";
          m(126) := x"FD10";
          m(127) := x"F621";
          m(128) := x"F603";
          m(129) := x"F8E6";
          m(130) := x"FB4B";
          m(131) := x"0040";
          m(132) := x"01F1";
          m(133) := x"016D";
          m(134) := x"02CD";
          m(135) := x"0138";
          m(136) := x"FF5C";
          m(137) := x"FE3E";
          m(138) := x"FF8C";
          m(139) := x"FFE3";
          m(140) := x"0025";
          m(141) := x"002D";
          m(142) := x"0022";
          m(143) := x"FFBC";
          m(144) := x"FFC8";
          m(145) := x"01D5";
          m(146) := x"02B5";
          m(147) := x"00B9";
          m(148) := x"0433";
          m(149) := x"016A";
          m(150) := x"008C";
          m(151) := x"FAE9";
          m(152) := x"FCB8";
          m(153) := x"FB79";
          m(154) := x"FC6F";
          m(155) := x"FA6F";
          m(156) := x"F9A5";
          m(157) := x"F9AC";
          m(158) := x"FD03";
          m(159) := x"F885";
          m(160) := x"FBB2";
          m(161) := x"FBA9";
          m(162) := x"001D";
          m(163) := x"FF42";
          m(164) := x"FF20";
          m(165) := x"FE8C";
          m(166) := x"FF5E";
          m(167) := x"000B";
          m(168) := x"FFF3";
          m(169) := x"000A";
          m(170) := x"FF58";
          m(171) := x"FF39";
          m(172) := x"FDF7";
          m(173) := x"0381";
          m(174) := x"0854";
          m(175) := x"04D8";
          m(176) := x"05F0";
          m(177) := x"009A";
          m(178) := x"01EC";
          m(179) := x"0032";
          m(180) := x"0238";
          m(181) := x"FCC7";
          m(182) := x"0193";
          m(183) := x"02ED";
          m(184) := x"0364";
          m(185) := x"0414";
          m(186) := x"FC13";
          m(187) := x"FBDA";
          m(188) := x"FC28";
          m(189) := x"FF8A";
          m(190) := x"FDE5";
          m(191) := x"FA8E";
          m(192) := x"FD9F";
          m(193) := x"FCCC";
          m(194) := x"FFCD";
          m(195) := x"FFDE";
          m(196) := x"FFC6";
          m(197) := x"FF5C";
          m(198) := x"FFDA";
          m(199) := x"00F1";
          m(200) := x"FD11";
          m(201) := x"FD34";
          m(202) := x"0556";
          m(203) := x"01A3";
          m(204) := x"FE47";
          m(205) := x"022E";
          m(206) := x"0476";
          m(207) := x"020E";
          m(208) := x"02E8";
          m(209) := x"FD9C";
          m(210) := x"FCB5";
          m(211) := x"FEF5";
          m(212) := x"0123";
          m(213) := x"0493";
          m(214) := x"FB73";
          m(215) := x"01DE";
          m(216) := x"03C7";
          m(217) := x"FE3C";
          m(218) := x"FCF1";
          m(219) := x"0062";
          m(220) := x"FF13";
          m(221) := x"FF0D";
          m(222) := x"0124";
          m(223) := x"FFE9";
          m(224) := x"FFC9";
          m(225) := x"006F";
          m(226) := x"0136";
          m(227) := x"FFC3";
          m(228) := x"FB53";
          m(229) := x"FE67";
          m(230) := x"031A";
          m(231) := x"010A";
          m(232) := x"052B";
          m(233) := x"039A";
          m(234) := x"00D2";
          m(235) := x"02C2";
          m(236) := x"FD07";
          m(237) := x"FC56";
          m(238) := x"FE05";
          m(239) := x"0191";
          m(240) := x"FB16";
          m(241) := x"FE83";
          m(242) := x"03B4";
          m(243) := x"0108";
          m(244) := x"017D";
          m(245) := x"FE18";
          m(246) := x"FF99";
          m(247) := x"FE32";
          m(248) := x"FF65";
          m(249) := x"FFDD";
          m(250) := x"FF47";
          m(251) := x"FFFF";
          m(252) := x"FFE8";
          m(253) := x"0005";
          m(254) := x"FF03";
          m(255) := x"FF2D";
          m(256) := x"FC8B";
          m(257) := x"02BE";
          m(258) := x"02D7";
          m(259) := x"0026";
          m(260) := x"0079";
          m(261) := x"0040";
          m(262) := x"057F";
          m(263) := x"0614";
          m(264) := x"FEE0";
          m(265) := x"0078";
          m(266) := x"FD85";
          m(267) := x"FD3D";
          m(268) := x"FC92";
          m(269) := x"02FA";
          m(270) := x"05D2";
          m(271) := x"01D5";
          m(272) := x"005E";
          m(273) := x"FF49";
          m(274) := x"03C9";
          m(275) := x"FC60";
          m(276) := x"FBCD";
          m(277) := x"FBB7";
          m(278) := x"FE67";
          m(279) := x"0028";
          m(280) := x"FFDA";
          m(281) := x"0047";
          m(282) := x"FFFF";
          m(283) := x"FEAB";
          m(284) := x"FC2B";
          m(285) := x"007A";
          m(286) := x"0051";
          m(287) := x"FFEE";
          m(288) := x"FDC6";
          m(289) := x"0397";
          m(290) := x"F933";
          m(291) := x"00EC";
          m(292) := x"05F6";
          m(293) := x"03FE";
          m(294) := x"FE3D";
          m(295) := x"027A";
          m(296) := x"FCFA";
          m(297) := x"FC7F";
          m(298) := x"FF24";
          m(299) := x"0662";
          m(300) := x"FD93";
          m(301) := x"FCD9";
          m(302) := x"FDC0";
          m(303) := x"F84D";
          m(304) := x"FA32";
          m(305) := x"FEF2";
          m(306) := x"FE51";
          m(307) := x"0011";
          m(308) := x"FFED";
          m(309) := x"0019";
          m(310) := x"00A9";
          m(311) := x"0091";
          m(312) := x"FA55";
          m(313) := x"F9ED";
          m(314) := x"FD75";
          m(315) := x"0214";
          m(316) := x"FE44";
          m(317) := x"FD82";
          m(318) := x"006A";
          m(319) := x"0633";
          m(320) := x"075D";
          m(321) := x"FF16";
          m(322) := x"0408";
          m(323) := x"0850";
          m(324) := x"05F3";
          m(325) := x"06B8";
          m(326) := x"0505";
          m(327) := x"04A9";
          m(328) := x"02A4";
          m(329) := x"FEEE";
          m(330) := x"FCB8";
          m(331) := x"FA8D";
          m(332) := x"F92A";
          m(333) := x"FE01";
          m(334) := x"FE3B";
          m(335) := x"FFF7";
          m(336) := x"0000";
          m(337) := x"FFF0";
          m(338) := x"0086";
          m(339) := x"FF92";
          m(340) := x"FD09";
          m(341) := x"FBC5";
          m(342) := x"FEA3";
          m(343) := x"0591";
          m(344) := x"053B";
          m(345) := x"0096";
          m(346) := x"01C5";
          m(347) := x"0750";
          m(348) := x"FDAB";
          m(349) := x"FAA2";
          m(350) := x"FB09";
          m(351) := x"096E";
          m(352) := x"0916";
          m(353) := x"FF9A";
          m(354) := x"06A5";
          m(355) := x"0889";
          m(356) := x"01C5";
          m(357) := x"FFB2";
          m(358) := x"00E2";
          m(359) := x"F909";
          m(360) := x"FAB9";
          m(361) := x"FEC9";
          m(362) := x"008C";
          m(363) := x"0050";
          m(364) := x"0000";
          m(365) := x"001A";
          m(366) := x"0085";
          m(367) := x"FE1F";
          m(368) := x"01A1";
          m(369) := x"01D6";
          m(370) := x"025D";
          m(371) := x"048D";
          m(372) := x"FFF8";
          m(373) := x"FFC5";
          m(374) := x"099A";
          m(375) := x"0002";
          m(376) := x"FBA9";
          m(377) := x"FAEF";
          m(378) := x"035D";
          m(379) := x"064F";
          m(380) := x"05AD";
          m(381) := x"03B3";
          m(382) := x"0194";
          m(383) := x"00B2";
          m(384) := x"023A";
          m(385) := x"0573";
          m(386) := x"FBF6";
          m(387) := x"F83D";
          m(388) := x"FED1";
          m(389) := x"FF9C";
          m(390) := x"FF50";
          m(391) := x"FFF2";
          m(392) := x"0008";
          m(393) := x"FFE7";
          m(394) := x"006E";
          m(395) := x"FE8D";
          m(396) := x"003D";
          m(397) := x"02A1";
          m(398) := x"FF4F";
          m(399) := x"0323";
          m(400) := x"0361";
          m(401) := x"FE4B";
          m(402) := x"038C";
          m(403) := x"00D6";
          m(404) := x"FD68";
          m(405) := x"FCD5";
          m(406) := x"01CA";
          m(407) := x"031D";
          m(408) := x"0469";
          m(409) := x"04F5";
          m(410) := x"0465";
          m(411) := x"0812";
          m(412) := x"06CE";
          m(413) := x"01F2";
          m(414) := x"0345";
          m(415) := x"014A";
          m(416) := x"FEAB";
          m(417) := x"FF4E";
          m(418) := x"FFDD";
          m(419) := x"FFE3";
          m(420) := x"0026";
          m(421) := x"FFDC";
          m(422) := x"FFF6";
          m(423) := x"014B";
          m(424) := x"008E";
          m(425) := x"020F";
          m(426) := x"0246";
          m(427) := x"FF79";
          m(428) := x"0263";
          m(429) := x"0245";
          m(430) := x"02FA";
          m(431) := x"FB0F";
          m(432) := x"F9E5";
          m(433) := x"FC92";
          m(434) := x"01FE";
          m(435) := x"06C7";
          m(436) := x"01D6";
          m(437) := x"0516";
          m(438) := x"02DA";
          m(439) := x"05A4";
          m(440) := x"038B";
          m(441) := x"00A8";
          m(442) := x"01F9";
          m(443) := x"FF8E";
          m(444) := x"FEE0";
          m(445) := x"FF33";
          m(446) := x"0041";
          m(447) := x"FFD2";
          m(448) := x"FFFB";
          m(449) := x"001D";
          m(450) := x"FFED";
          m(451) := x"0161";
          m(452) := x"0384";
          m(453) := x"022E";
          m(454) := x"0305";
          m(455) := x"0463";
          m(456) := x"03AE";
          m(457) := x"FD75";
          m(458) := x"031D";
          m(459) := x"FEB4";
          m(460) := x"FF3A";
          m(461) := x"FC89";
          m(462) := x"0487";
          m(463) := x"066B";
          m(464) := x"03BD";
          m(465) := x"06E3";
          m(466) := x"0976";
          m(467) := x"011D";
          m(468) := x"01CF";
          m(469) := x"FA28";
          m(470) := x"FB02";
          m(471) := x"FDC7";
          m(472) := x"FCE6";
          m(473) := x"FF2B";
          m(474) := x"0000";
          m(475) := x"FFEB";
          m(476) := x"0034";
          m(477) := x"0007";
          m(478) := x"FFCD";
          m(479) := x"FFF6";
          m(480) := x"01D8";
          m(481) := x"00FB";
          m(482) := x"032D";
          m(483) := x"0303";
          m(484) := x"FFDF";
          m(485) := x"FBAE";
          m(486) := x"FBC6";
          m(487) := x"FF71";
          m(488) := x"02A9";
          m(489) := x"FD48";
          m(490) := x"027F";
          m(491) := x"06CD";
          m(492) := x"05D5";
          m(493) := x"0A07";
          m(494) := x"0820";
          m(495) := x"F9D5";
          m(496) := x"FC67";
          m(497) := x"00DE";
          m(498) := x"00D2";
          m(499) := x"036F";
          m(500) := x"00BC";
          m(501) := x"00D2";
          m(502) := x"00FC";
          m(503) := x"0012";
          m(504) := x"FFE0";
          m(505) := x"0003";
          m(506) := x"FFEB";
          m(507) := x"FF04";
          m(508) := x"0248";
          m(509) := x"00CA";
          m(510) := x"0439";
          m(511) := x"0479";
          m(512) := x"03B9";
          m(513) := x"002A";
          m(514) := x"FE53";
          m(515) := x"FD8A";
          m(516) := x"FC2D";
          m(517) := x"031A";
          m(518) := x"099A";
          m(519) := x"0797";
          m(520) := x"066E";
          m(521) := x"060A";
          m(522) := x"FD95";
          m(523) := x"FBC4";
          m(524) := x"027A";
          m(525) := x"07FA";
          m(526) := x"004D";
          m(527) := x"FDE9";
          m(528) := x"FFE2";
          m(529) := x"0041";
          m(530) := x"00A8";
          m(531) := x"FFDF";
          m(532) := x"FFEC";
          m(533) := x"FFF7";
          m(534) := x"FF9E";
          m(535) := x"FEB0";
          m(536) := x"FFC6";
          m(537) := x"FEBF";
          m(538) := x"FF49";
          m(539) := x"03A2";
          m(540) := x"0206";
          m(541) := x"0162";
          m(542) := x"04AD";
          m(543) := x"0302";
          m(544) := x"02BB";
          m(545) := x"016D";
          m(546) := x"03F1";
          m(547) := x"03A2";
          m(548) := x"FEBC";
          m(549) := x"FB31";
          m(550) := x"FC98";
          m(551) := x"FEC7";
          m(552) := x"FFA4";
          m(553) := x"FF06";
          m(554) := x"F797";
          m(555) := x"F9F7";
          m(556) := x"FEBD";
          m(557) := x"FFFD";
          m(558) := x"0008";
          m(559) := x"FFE9";
          m(560) := x"000B";
          m(561) := x"001B";
          m(562) := x"FF42";
          m(563) := x"FD5D";
          m(564) := x"FE6F";
          m(565) := x"FD4D";
          m(566) := x"FCB0";
          m(567) := x"FB2D";
          m(568) := x"F94F";
          m(569) := x"FC55";
          m(570) := x"FD75";
          m(571) := x"FE37";
          m(572) := x"FD33";
          m(573) := x"F7C3";
          m(574) := x"F72F";
          m(575) := x"F495";
          m(576) := x"F9D0";
          m(577) := x"F57F";
          m(578) := x"F840";
          m(579) := x"F7F6";
          m(580) := x"F51D";
          m(581) := x"F2F1";
          m(582) := x"F47B";
          m(583) := x"FACB";
          m(584) := x"00A9";
          m(585) := x"FFCE";
          m(586) := x"FFEF";
          m(587) := x"FFAA";
          m(588) := x"0043";
          m(589) := x"FFF1";
          m(590) := x"FEE9";
          m(591) := x"FC25";
          m(592) := x"FEBC";
          m(593) := x"FD2B";
          m(594) := x"FA92";
          m(595) := x"F7C9";
          m(596) := x"F32A";
          m(597) := x"F759";
          m(598) := x"F5CF";
          m(599) := x"F2D4";
          m(600) := x"F42D";
          m(601) := x"F346";
          m(602) := x"F242";
          m(603) := x"F111";
          m(604) := x"FC4D";
          m(605) := x"F608";
          m(606) := x"F33D";
          m(607) := x"FB87";
          m(608) := x"F9DB";
          m(609) := x"F835";
          m(610) := x"F964";
          m(611) := x"FB14";
          m(612) := x"0008";
          m(613) := x"0032";
          m(614) := x"FFE4";
          m(615) := x"FFCF";
          m(616) := x"FFF5";
          m(617) := x"001E";
          m(618) := x"FF10";
          m(619) := x"FD4E";
          m(620) := x"FD79";
          m(621) := x"FC01";
          m(622) := x"FCC9";
          m(623) := x"FD8A";
          m(624) := x"FDE1";
          m(625) := x"F85E";
          m(626) := x"F959";
          m(627) := x"F74B";
          m(628) := x"F75F";
          m(629) := x"F8A6";
          m(630) := x"FEF1";
          m(631) := x"F99B";
          m(632) := x"F867";
          m(633) := x"F9A9";
          m(634) := x"F9FE";
          m(635) := x"FBD0";
          m(636) := x"FD02";
          m(637) := x"FAB4";
          m(638) := x"FD6D";
          m(639) := x"FC88";
          m(640) := x"FEE1";
          m(641) := x"FF6C";
          m(642) := x"002E";
          m(643) := x"FFF2";
          m(644) := x"FFF4";
          m(645) := x"0002";
          m(646) := x"FF28";
          m(647) := x"FCDB";
          m(648) := x"FBFA";
          m(649) := x"FCED";
          m(650) := x"0076";
          m(651) := x"03D4";
          m(652) := x"0290";
          m(653) := x"FC46";
          m(654) := x"FD4F";
          m(655) := x"FD75";
          m(656) := x"FAE6";
          m(657) := x"F892";
          m(658) := x"FD06";
          m(659) := x"F993";
          m(660) := x"F9BB";
          m(661) := x"F891";
          m(662) := x"F7CA";
          m(663) := x"FDB4";
          m(664) := x"FBEA";
          m(665) := x"FCAB";
          m(666) := x"FC97";
          m(667) := x"FC36";
          m(668) := x"FE85";
          m(669) := x"FF65";
          m(670) := x"FFC9";
          m(671) := x"0024";
          m(672) := x"0009";
          m(673) := x"0001";
          m(674) := x"FFFD";
          m(675) := x"FEFF";
          m(676) := x"0002";
          m(677) := x"0464";
          m(678) := x"0061";
          m(679) := x"FF7C";
          m(680) := x"FE65";
          m(681) := x"FA99";
          m(682) := x"F679";
          m(683) := x"FD10";
          m(684) := x"F8D2";
          m(685) := x"F8AA";
          m(686) := x"F7EA";
          m(687) := x"FAAC";
          m(688) := x"F707";
          m(689) := x"FCA7";
          m(690) := x"F95A";
          m(691) := x"F994";
          m(692) := x"FDD0";
          m(693) := x"FEAB";
          m(694) := x"FF98";
          m(695) := x"FF7D";
          m(696) := x"FD9A";
          m(697) := x"FF84";
          m(698) := x"FFFB";
          m(699) := x"002A";
          m(700) := x"0017";
          m(701) := x"0000";
          m(702) := x"FFE3";
          m(703) := x"002B";
          m(704) := x"0205";
          m(705) := x"009E";
          m(706) := x"FD70";
          m(707) := x"FE37";
          m(708) := x"FAF9";
          m(709) := x"F9CE";
          m(710) := x"F79B";
          m(711) := x"0245";
          m(712) := x"FA64";
          m(713) := x"FC12";
          m(714) := x"014B";
          m(715) := x"FCA6";
          m(716) := x"FDE9";
          m(717) := x"FC97";
          m(718) := x"FA3E";
          m(719) := x"F85F";
          m(720) := x"FE45";
          m(721) := x"FF44";
          m(722) := x"FF57";
          m(723) := x"FF97";
          m(724) := x"FEFF";
          m(725) := x"FFE5";
          m(726) := x"FFFA";
          m(727) := x"0010";
          m(728) := x"FFDD";
          m(729) := x"0018";
          m(730) := x"FFDB";
          m(731) := x"FFFB";
          m(732) := x"0001";
          m(733) := x"005B";
          m(734) := x"00E7";
          m(735) := x"00D8";
          m(736) := x"01CA";
          m(737) := x"02E8";
          m(738) := x"0146";
          m(739) := x"00EC";
          m(740) := x"FEAC";
          m(741) := x"FE23";
          m(742) := x"040A";
          m(743) := x"FFCA";
          m(744) := x"FE1A";
          m(745) := x"FD4A";
          m(746) := x"FF86";
          m(747) := x"0076";
          m(748) := x"0012";
          m(749) := x"FFD9";
          m(750) := x"00BD";
          m(751) := x"0018";
          m(752) := x"FFF1";
          m(753) := x"0002";
          m(754) := x"FFD5";
          m(755) := x"FFBE";
          m(756) := x"000E";
          m(757) := x"FFE7";
          m(758) := x"0039";
          m(759) := x"FFEE";
          m(760) := x"0020";
          m(761) := x"0007";
          m(762) := x"0029";
          m(763) := x"FFFC";
          m(764) := x"0029";
          m(765) := x"0053";
          m(766) := x"007C";
          m(767) := x"0019";
          m(768) := x"0037";
          m(769) := x"0044";
          m(770) := x"009A";
          m(771) := x"00A5";
          m(772) := x"00DA";
          m(773) := x"009F";
          m(774) := x"0111";
          m(775) := x"0051";
          m(776) := x"0040";
          m(777) := x"0085";
          m(778) := x"0092";
          m(779) := x"0026";
          m(780) := x"FFDC";
          m(781) := x"0004";
          m(782) := x"FFF7";
          m(783) := x"FFF6";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_16.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 16) then
          m(0) := x"FFFD";
          m(1) := x"002A";
          m(2) := x"FFDF";
          m(3) := x"002D";
          m(4) := x"FFEE";
          m(5) := x"FFF5";
          m(6) := x"0033";
          m(7) := x"000B";
          m(8) := x"000C";
          m(9) := x"FFE5";
          m(10) := x"0020";
          m(11) := x"FFEF";
          m(12) := x"000D";
          m(13) := x"0021";
          m(14) := x"0002";
          m(15) := x"FFD4";
          m(16) := x"0001";
          m(17) := x"000E";
          m(18) := x"FFC5";
          m(19) := x"0005";
          m(20) := x"FFC8";
          m(21) := x"0026";
          m(22) := x"FFE1";
          m(23) := x"FFD4";
          m(24) := x"FFF7";
          m(25) := x"FFFE";
          m(26) := x"0000";
          m(27) := x"FFE0";
          m(28) := x"001C";
          m(29) := x"FFBC";
          m(30) := x"FFD8";
          m(31) := x"FFE6";
          m(32) := x"FFE9";
          m(33) := x"FFDA";
          m(34) := x"0010";
          m(35) := x"000F";
          m(36) := x"0033";
          m(37) := x"001A";
          m(38) := x"0000";
          m(39) := x"0046";
          m(40) := x"FFD2";
          m(41) := x"FFA4";
          m(42) := x"FFCA";
          m(43) := x"FFEC";
          m(44) := x"00FF";
          m(45) := x"0051";
          m(46) := x"FFF3";
          m(47) := x"FFC7";
          m(48) := x"FFD7";
          m(49) := x"FFB1";
          m(50) := x"FFCD";
          m(51) := x"FFA9";
          m(52) := x"FFE8";
          m(53) := x"0010";
          m(54) := x"FFD8";
          m(55) := x"FFD9";
          m(56) := x"FFE5";
          m(57) := x"002F";
          m(58) := x"FFFC";
          m(59) := x"FFF7";
          m(60) := x"FFFB";
          m(61) := x"0001";
          m(62) := x"0011";
          m(63) := x"FFAC";
          m(64) := x"0034";
          m(65) := x"0092";
          m(66) := x"0076";
          m(67) := x"003C";
          m(68) := x"0070";
          m(69) := x"0000";
          m(70) := x"FE97";
          m(71) := x"FCC6";
          m(72) := x"FECB";
          m(73) := x"FC39";
          m(74) := x"FC44";
          m(75) := x"FD16";
          m(76) := x"FEA3";
          m(77) := x"FDE7";
          m(78) := x"FEF0";
          m(79) := x"FFC0";
          m(80) := x"00A0";
          m(81) := x"008C";
          m(82) := x"FFF4";
          m(83) := x"0019";
          m(84) := x"FFC9";
          m(85) := x"FFDE";
          m(86) := x"0007";
          m(87) := x"0019";
          m(88) := x"FFEA";
          m(89) := x"FFF5";
          m(90) := x"000D";
          m(91) := x"0034";
          m(92) := x"0135";
          m(93) := x"0156";
          m(94) := x"0393";
          m(95) := x"03C2";
          m(96) := x"04A7";
          m(97) := x"03C3";
          m(98) := x"FF94";
          m(99) := x"FD5D";
          m(100) := x"02EF";
          m(101) := x"0160";
          m(102) := x"FD0D";
          m(103) := x"FC33";
          m(104) := x"FDC1";
          m(105) := x"FCF5";
          m(106) := x"FD43";
          m(107) := x"FD19";
          m(108) := x"FEB4";
          m(109) := x"0083";
          m(110) := x"FFE3";
          m(111) := x"000D";
          m(112) := x"FFF1";
          m(113) := x"FFDC";
          m(114) := x"FFE9";
          m(115) := x"0025";
          m(116) := x"0027";
          m(117) := x"0017";
          m(118) := x"00F0";
          m(119) := x"025D";
          m(120) := x"0611";
          m(121) := x"0541";
          m(122) := x"06D8";
          m(123) := x"08A1";
          m(124) := x"0702";
          m(125) := x"04B5";
          m(126) := x"060A";
          m(127) := x"08E8";
          m(128) := x"0115";
          m(129) := x"FDC4";
          m(130) := x"FF72";
          m(131) := x"FE50";
          m(132) := x"FE2C";
          m(133) := x"FCFB";
          m(134) := x"FD0B";
          m(135) := x"F82D";
          m(136) := x"FC86";
          m(137) := x"FFD8";
          m(138) := x"006E";
          m(139) := x"FFD2";
          m(140) := x"0019";
          m(141) := x"000C";
          m(142) := x"0036";
          m(143) := x"0015";
          m(144) := x"0011";
          m(145) := x"0092";
          m(146) := x"01C7";
          m(147) := x"033D";
          m(148) := x"06EF";
          m(149) := x"07CE";
          m(150) := x"0BED";
          m(151) := x"05BD";
          m(152) := x"FF9D";
          m(153) := x"001A";
          m(154) := x"FD05";
          m(155) := x"FB03";
          m(156) := x"01A3";
          m(157) := x"003B";
          m(158) := x"078E";
          m(159) := x"018A";
          m(160) := x"FD28";
          m(161) := x"FD97";
          m(162) := x"FE09";
          m(163) := x"F94F";
          m(164) := x"FAEA";
          m(165) := x"FF71";
          m(166) := x"FF69";
          m(167) := x"FF8A";
          m(168) := x"000E";
          m(169) := x"FFFE";
          m(170) := x"000B";
          m(171) := x"FFFE";
          m(172) := x"0030";
          m(173) := x"FF64";
          m(174) := x"024B";
          m(175) := x"074D";
          m(176) := x"0A7E";
          m(177) := x"0F88";
          m(178) := x"0CA8";
          m(179) := x"00FB";
          m(180) := x"FB9C";
          m(181) := x"0147";
          m(182) := x"F95A";
          m(183) := x"F718";
          m(184) := x"023D";
          m(185) := x"0375";
          m(186) := x"042C";
          m(187) := x"009E";
          m(188) := x"FD8D";
          m(189) := x"014C";
          m(190) := x"FFA0";
          m(191) := x"F8FE";
          m(192) := x"FAF2";
          m(193) := x"FFCC";
          m(194) := x"FFDF";
          m(195) := x"FFCC";
          m(196) := x"0008";
          m(197) := x"0084";
          m(198) := x"004E";
          m(199) := x"00B9";
          m(200) := x"FF9A";
          m(201) := x"FF07";
          m(202) := x"0244";
          m(203) := x"05D3";
          m(204) := x"09D8";
          m(205) := x"0DCB";
          m(206) := x"0651";
          m(207) := x"FFD8";
          m(208) := x"FEAD";
          m(209) := x"01A5";
          m(210) := x"FCEA";
          m(211) := x"FEAE";
          m(212) := x"0581";
          m(213) := x"0380";
          m(214) := x"0549";
          m(215) := x"0256";
          m(216) := x"FD8E";
          m(217) := x"0419";
          m(218) := x"0167";
          m(219) := x"FD1E";
          m(220) := x"FC8D";
          m(221) := x"FF15";
          m(222) := x"FF6E";
          m(223) := x"0035";
          m(224) := x"0012";
          m(225) := x"0012";
          m(226) := x"006E";
          m(227) := x"0090";
          m(228) := x"FFEB";
          m(229) := x"FF3E";
          m(230) := x"FFF2";
          m(231) := x"0252";
          m(232) := x"074C";
          m(233) := x"0FCF";
          m(234) := x"0BDA";
          m(235) := x"F8AF";
          m(236) := x"F95A";
          m(237) := x"FA7C";
          m(238) := x"FFCD";
          m(239) := x"0209";
          m(240) := x"06E2";
          m(241) := x"0477";
          m(242) := x"02B1";
          m(243) := x"012C";
          m(244) := x"FDE3";
          m(245) := x"0249";
          m(246) := x"FDCB";
          m(247) := x"FBF7";
          m(248) := x"F93A";
          m(249) := x"FCDF";
          m(250) := x"000B";
          m(251) := x"0004";
          m(252) := x"FFE7";
          m(253) := x"000B";
          m(254) := x"001E";
          m(255) := x"020F";
          m(256) := x"012C";
          m(257) := x"009E";
          m(258) := x"00E3";
          m(259) := x"00E8";
          m(260) := x"073F";
          m(261) := x"0BB3";
          m(262) := x"059B";
          m(263) := x"FAF0";
          m(264) := x"FC8C";
          m(265) := x"FC8C";
          m(266) := x"FB9A";
          m(267) := x"FD42";
          m(268) := x"05B9";
          m(269) := x"0811";
          m(270) := x"04F3";
          m(271) := x"0514";
          m(272) := x"0345";
          m(273) := x"0197";
          m(274) := x"008E";
          m(275) := x"FD21";
          m(276) := x"FCBB";
          m(277) := x"FF92";
          m(278) := x"00F5";
          m(279) := x"018D";
          m(280) := x"FFF6";
          m(281) := x"0039";
          m(282) := x"006A";
          m(283) := x"019D";
          m(284) := x"029B";
          m(285) := x"034C";
          m(286) := x"0306";
          m(287) := x"02C2";
          m(288) := x"04D2";
          m(289) := x"0921";
          m(290) := x"0416";
          m(291) := x"030B";
          m(292) := x"FCE6";
          m(293) := x"FA40";
          m(294) := x"F679";
          m(295) := x"FDFC";
          m(296) := x"043C";
          m(297) := x"097A";
          m(298) := x"0875";
          m(299) := x"0284";
          m(300) := x"0736";
          m(301) := x"0394";
          m(302) := x"02B7";
          m(303) := x"FF55";
          m(304) := x"000B";
          m(305) := x"013A";
          m(306) := x"01D6";
          m(307) := x"0051";
          m(308) := x"0050";
          m(309) := x"0050";
          m(310) := x"FFCB";
          m(311) := x"0222";
          m(312) := x"02BD";
          m(313) := x"03A3";
          m(314) := x"0308";
          m(315) := x"0489";
          m(316) := x"06D4";
          m(317) := x"0669";
          m(318) := x"FED1";
          m(319) := x"01B2";
          m(320) := x"F81C";
          m(321) := x"01D6";
          m(322) := x"00D7";
          m(323) := x"FCBC";
          m(324) := x"FA7D";
          m(325) := x"056A";
          m(326) := x"0464";
          m(327) := x"03DB";
          m(328) := x"006A";
          m(329) := x"019C";
          m(330) := x"0727";
          m(331) := x"03AD";
          m(332) := x"022C";
          m(333) := x"01F0";
          m(334) := x"0129";
          m(335) := x"FFC1";
          m(336) := x"0001";
          m(337) := x"FFE8";
          m(338) := x"FFF1";
          m(339) := x"01A0";
          m(340) := x"01F1";
          m(341) := x"0402";
          m(342) := x"0309";
          m(343) := x"033F";
          m(344) := x"0410";
          m(345) := x"0501";
          m(346) := x"01AC";
          m(347) := x"F3EA";
          m(348) := x"F23B";
          m(349) := x"FB1C";
          m(350) := x"F9FC";
          m(351) := x"FC45";
          m(352) := x"FEFB";
          m(353) := x"FE1D";
          m(354) := x"07B4";
          m(355) := x"049F";
          m(356) := x"FD1A";
          m(357) := x"00E7";
          m(358) := x"05F9";
          m(359) := x"0336";
          m(360) := x"050B";
          m(361) := x"05F1";
          m(362) := x"0215";
          m(363) := x"0020";
          m(364) := x"FFDF";
          m(365) := x"0002";
          m(366) := x"00BD";
          m(367) := x"0114";
          m(368) := x"02C0";
          m(369) := x"0428";
          m(370) := x"0448";
          m(371) := x"001A";
          m(372) := x"FCDD";
          m(373) := x"FF1F";
          m(374) := x"03BF";
          m(375) := x"0010";
          m(376) := x"FA0C";
          m(377) := x"FBF9";
          m(378) := x"0007";
          m(379) := x"F8F3";
          m(380) := x"FC50";
          m(381) := x"FFFD";
          m(382) := x"05E4";
          m(383) := x"05BA";
          m(384) := x"FB4E";
          m(385) := x"03A9";
          m(386) := x"07BD";
          m(387) := x"0797";
          m(388) := x"095F";
          m(389) := x"05C1";
          m(390) := x"0139";
          m(391) := x"FFF7";
          m(392) := x"FFF0";
          m(393) := x"000F";
          m(394) := x"0046";
          m(395) := x"0071";
          m(396) := x"022C";
          m(397) := x"02ED";
          m(398) := x"06A6";
          m(399) := x"020A";
          m(400) := x"FC96";
          m(401) := x"FFD3";
          m(402) := x"FE9B";
          m(403) := x"FF29";
          m(404) := x"0151";
          m(405) := x"FB89";
          m(406) := x"01E1";
          m(407) := x"FED3";
          m(408) := x"FE16";
          m(409) := x"01DF";
          m(410) := x"0537";
          m(411) := x"054E";
          m(412) := x"FA18";
          m(413) := x"0020";
          m(414) := x"05E9";
          m(415) := x"073F";
          m(416) := x"0544";
          m(417) := x"01EC";
          m(418) := x"0212";
          m(419) := x"FFF4";
          m(420) := x"FFFB";
          m(421) := x"0018";
          m(422) := x"0021";
          m(423) := x"007D";
          m(424) := x"015B";
          m(425) := x"02F1";
          m(426) := x"024F";
          m(427) := x"FC8A";
          m(428) := x"FEE8";
          m(429) := x"02FD";
          m(430) := x"03F6";
          m(431) := x"036F";
          m(432) := x"FD80";
          m(433) := x"00D2";
          m(434) := x"FA9B";
          m(435) := x"FC37";
          m(436) := x"FB5A";
          m(437) := x"FFEA";
          m(438) := x"0046";
          m(439) := x"FF14";
          m(440) := x"FF7C";
          m(441) := x"FDD5";
          m(442) := x"039C";
          m(443) := x"0372";
          m(444) := x"05C8";
          m(445) := x"04FB";
          m(446) := x"03F2";
          m(447) := x"FFD8";
          m(448) := x"0020";
          m(449) := x"000B";
          m(450) := x"0089";
          m(451) := x"0115";
          m(452) := x"01C3";
          m(453) := x"FF3B";
          m(454) := x"01CA";
          m(455) := x"01E5";
          m(456) := x"FF4F";
          m(457) := x"0618";
          m(458) := x"08E1";
          m(459) := x"FDEC";
          m(460) := x"0140";
          m(461) := x"0007";
          m(462) := x"FB81";
          m(463) := x"FC41";
          m(464) := x"FE4C";
          m(465) := x"0442";
          m(466) := x"0334";
          m(467) := x"FEFD";
          m(468) := x"01EE";
          m(469) := x"FD02";
          m(470) := x"014F";
          m(471) := x"02DB";
          m(472) := x"0555";
          m(473) := x"0403";
          m(474) := x"0190";
          m(475) := x"FFFA";
          m(476) := x"FFD1";
          m(477) := x"FFEE";
          m(478) := x"00AF";
          m(479) := x"0085";
          m(480) := x"005A";
          m(481) := x"FE83";
          m(482) := x"020B";
          m(483) := x"FE88";
          m(484) := x"FE56";
          m(485) := x"FD5E";
          m(486) := x"FB68";
          m(487) := x"FD27";
          m(488) := x"0334";
          m(489) := x"02D4";
          m(490) := x"019F";
          m(491) := x"0224";
          m(492) := x"FEFA";
          m(493) := x"0301";
          m(494) := x"FE7D";
          m(495) := x"014F";
          m(496) := x"0058";
          m(497) := x"0185";
          m(498) := x"0337";
          m(499) := x"016C";
          m(500) := x"0396";
          m(501) := x"02D1";
          m(502) := x"00AE";
          m(503) := x"0090";
          m(504) := x"FFFC";
          m(505) := x"FFDC";
          m(506) := x"0068";
          m(507) := x"00A7";
          m(508) := x"FECD";
          m(509) := x"013C";
          m(510) := x"00B5";
          m(511) := x"FCD0";
          m(512) := x"FF8A";
          m(513) := x"FBAD";
          m(514) := x"FEBC";
          m(515) := x"FF25";
          m(516) := x"0377";
          m(517) := x"00D6";
          m(518) := x"FBDC";
          m(519) := x"0214";
          m(520) := x"FCA3";
          m(521) := x"FE8A";
          m(522) := x"00C5";
          m(523) := x"00AC";
          m(524) := x"FF8C";
          m(525) := x"01EB";
          m(526) := x"0425";
          m(527) := x"048F";
          m(528) := x"0475";
          m(529) := x"01CB";
          m(530) := x"0072";
          m(531) := x"FFE3";
          m(532) := x"FFAD";
          m(533) := x"FFB8";
          m(534) := x"0051";
          m(535) := x"01F2";
          m(536) := x"FE59";
          m(537) := x"0150";
          m(538) := x"01A2";
          m(539) := x"FF96";
          m(540) := x"FDCA";
          m(541) := x"FA37";
          m(542) := x"FBF9";
          m(543) := x"FA37";
          m(544) := x"0314";
          m(545) := x"00C6";
          m(546) := x"FE8B";
          m(547) := x"FE21";
          m(548) := x"FBD5";
          m(549) := x"0235";
          m(550) := x"03C0";
          m(551) := x"00C0";
          m(552) := x"00F1";
          m(553) := x"02DC";
          m(554) := x"0462";
          m(555) := x"0349";
          m(556) := x"01E0";
          m(557) := x"0123";
          m(558) := x"FFD7";
          m(559) := x"FFED";
          m(560) := x"FFF4";
          m(561) := x"0050";
          m(562) := x"FFF3";
          m(563) := x"0345";
          m(564) := x"006C";
          m(565) := x"FF18";
          m(566) := x"0041";
          m(567) := x"0285";
          m(568) := x"FD20";
          m(569) := x"FCDB";
          m(570) := x"FED7";
          m(571) := x"FF58";
          m(572) := x"0098";
          m(573) := x"0428";
          m(574) := x"FDB0";
          m(575) := x"03DB";
          m(576) := x"0267";
          m(577) := x"FF4B";
          m(578) := x"FE84";
          m(579) := x"FF0C";
          m(580) := x"0356";
          m(581) := x"02A8";
          m(582) := x"0420";
          m(583) := x"031B";
          m(584) := x"01D7";
          m(585) := x"00F5";
          m(586) := x"FFFC";
          m(587) := x"0025";
          m(588) := x"FFD0";
          m(589) := x"0034";
          m(590) := x"0065";
          m(591) := x"01D2";
          m(592) := x"010B";
          m(593) := x"0031";
          m(594) := x"00F4";
          m(595) := x"FF9D";
          m(596) := x"0057";
          m(597) := x"FF83";
          m(598) := x"0173";
          m(599) := x"FBFE";
          m(600) := x"0006";
          m(601) := x"FDD9";
          m(602) := x"03A4";
          m(603) := x"03D3";
          m(604) := x"01D9";
          m(605) := x"FEC5";
          m(606) := x"0070";
          m(607) := x"032B";
          m(608) := x"03F0";
          m(609) := x"03DB";
          m(610) := x"02AC";
          m(611) := x"0169";
          m(612) := x"008E";
          m(613) := x"0062";
          m(614) := x"FFD9";
          m(615) := x"FFD4";
          m(616) := x"FFBB";
          m(617) := x"FFBE";
          m(618) := x"0006";
          m(619) := x"0044";
          m(620) := x"011C";
          m(621) := x"01A1";
          m(622) := x"01D3";
          m(623) := x"0154";
          m(624) := x"0167";
          m(625) := x"028A";
          m(626) := x"0175";
          m(627) := x"019A";
          m(628) := x"0260";
          m(629) := x"F9C2";
          m(630) := x"FDD5";
          m(631) := x"004A";
          m(632) := x"FE4B";
          m(633) := x"FB17";
          m(634) := x"FFDC";
          m(635) := x"FEFB";
          m(636) := x"00A5";
          m(637) := x"018E";
          m(638) := x"0188";
          m(639) := x"009F";
          m(640) := x"FFE5";
          m(641) := x"FFCB";
          m(642) := x"0023";
          m(643) := x"FFF1";
          m(644) := x"0003";
          m(645) := x"000A";
          m(646) := x"0036";
          m(647) := x"FFFE";
          m(648) := x"01B4";
          m(649) := x"00A4";
          m(650) := x"FD4F";
          m(651) := x"FEB4";
          m(652) := x"FD25";
          m(653) := x"FE9A";
          m(654) := x"FC2C";
          m(655) := x"03EB";
          m(656) := x"01A2";
          m(657) := x"FFC4";
          m(658) := x"FCF7";
          m(659) := x"FBF7";
          m(660) := x"FDD1";
          m(661) := x"0359";
          m(662) := x"00E0";
          m(663) := x"FCE6";
          m(664) := x"FE14";
          m(665) := x"FFF1";
          m(666) := x"006E";
          m(667) := x"0051";
          m(668) := x"000F";
          m(669) := x"0003";
          m(670) := x"FFFF";
          m(671) := x"0013";
          m(672) := x"FFFD";
          m(673) := x"FFE4";
          m(674) := x"0028";
          m(675) := x"0073";
          m(676) := x"0206";
          m(677) := x"0387";
          m(678) := x"02C6";
          m(679) := x"000E";
          m(680) := x"FE24";
          m(681) := x"F720";
          m(682) := x"FA60";
          m(683) := x"05FC";
          m(684) := x"0184";
          m(685) := x"00BD";
          m(686) := x"0544";
          m(687) := x"FFEF";
          m(688) := x"034F";
          m(689) := x"0753";
          m(690) := x"004D";
          m(691) := x"FB52";
          m(692) := x"FBAE";
          m(693) := x"FE15";
          m(694) := x"FF25";
          m(695) := x"FFBA";
          m(696) := x"0021";
          m(697) := x"FFFF";
          m(698) := x"0006";
          m(699) := x"0023";
          m(700) := x"000D";
          m(701) := x"FFE2";
          m(702) := x"0032";
          m(703) := x"0022";
          m(704) := x"0126";
          m(705) := x"026B";
          m(706) := x"03DC";
          m(707) := x"0417";
          m(708) := x"017B";
          m(709) := x"0057";
          m(710) := x"0101";
          m(711) := x"0035";
          m(712) := x"FE6B";
          m(713) := x"FE45";
          m(714) := x"0092";
          m(715) := x"0060";
          m(716) := x"0143";
          m(717) := x"01CC";
          m(718) := x"01E8";
          m(719) := x"FFC0";
          m(720) := x"FD97";
          m(721) := x"FDF4";
          m(722) := x"FDE7";
          m(723) := x"FF37";
          m(724) := x"FFEB";
          m(725) := x"FFE5";
          m(726) := x"FFFB";
          m(727) := x"FFB4";
          m(728) := x"FFDD";
          m(729) := x"0012";
          m(730) := x"FFF6";
          m(731) := x"002B";
          m(732) := x"FFB5";
          m(733) := x"0045";
          m(734) := x"0069";
          m(735) := x"0076";
          m(736) := x"0151";
          m(737) := x"011B";
          m(738) := x"02C5";
          m(739) := x"0282";
          m(740) := x"0028";
          m(741) := x"0207";
          m(742) := x"FF02";
          m(743) := x"FD92";
          m(744) := x"FF34";
          m(745) := x"0092";
          m(746) := x"015A";
          m(747) := x"00A5";
          m(748) := x"0034";
          m(749) := x"FFE3";
          m(750) := x"0019";
          m(751) := x"FFDD";
          m(752) := x"003B";
          m(753) := x"0007";
          m(754) := x"001A";
          m(755) := x"FFE1";
          m(756) := x"FFFB";
          m(757) := x"0016";
          m(758) := x"FFFF";
          m(759) := x"000F";
          m(760) := x"001D";
          m(761) := x"FFFA";
          m(762) := x"FFF2";
          m(763) := x"FFB5";
          m(764) := x"FF89";
          m(765) := x"FFFB";
          m(766) := x"0072";
          m(767) := x"001F";
          m(768) := x"FFF4";
          m(769) := x"FFD0";
          m(770) := x"0027";
          m(771) := x"FEF9";
          m(772) := x"FEF9";
          m(773) := x"FFF9";
          m(774) := x"0017";
          m(775) := x"FFF4";
          m(776) := x"FFDE";
          m(777) := x"FFF7";
          m(778) := x"FFF1";
          m(779) := x"001A";
          m(780) := x"FFE9";
          m(781) := x"FFF2";
          m(782) := x"FFB1";
          m(783) := x"FFE6";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_17.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 17) then
          m(0) := x"0004";
          m(1) := x"0017";
          m(2) := x"FFD0";
          m(3) := x"FFCC";
          m(4) := x"FFE5";
          m(5) := x"FFE8";
          m(6) := x"FFD9";
          m(7) := x"0033";
          m(8) := x"FFDF";
          m(9) := x"0023";
          m(10) := x"FFB6";
          m(11) := x"FFB7";
          m(12) := x"001D";
          m(13) := x"002A";
          m(14) := x"FFE6";
          m(15) := x"000E";
          m(16) := x"FFF8";
          m(17) := x"FFF2";
          m(18) := x"FFD2";
          m(19) := x"FFD8";
          m(20) := x"FFB4";
          m(21) := x"0014";
          m(22) := x"000C";
          m(23) := x"FFD7";
          m(24) := x"0023";
          m(25) := x"0013";
          m(26) := x"0040";
          m(27) := x"0002";
          m(28) := x"0028";
          m(29) := x"FFC8";
          m(30) := x"0008";
          m(31) := x"FFE2";
          m(32) := x"0008";
          m(33) := x"FFED";
          m(34) := x"0003";
          m(35) := x"FFD9";
          m(36) := x"FFAC";
          m(37) := x"FFD8";
          m(38) := x"FFE1";
          m(39) := x"FFD9";
          m(40) := x"FFB3";
          m(41) := x"FFB3";
          m(42) := x"0006";
          m(43) := x"003B";
          m(44) := x"003B";
          m(45) := x"FFBC";
          m(46) := x"FFF8";
          m(47) := x"000D";
          m(48) := x"FFDD";
          m(49) := x"FFFC";
          m(50) := x"FFD8";
          m(51) := x"0013";
          m(52) := x"0023";
          m(53) := x"FFFE";
          m(54) := x"000E";
          m(55) := x"FFEE";
          m(56) := x"0010";
          m(57) := x"FFC6";
          m(58) := x"000B";
          m(59) := x"FFEB";
          m(60) := x"0004";
          m(61) := x"0048";
          m(62) := x"FFD0";
          m(63) := x"FF76";
          m(64) := x"FF8F";
          m(65) := x"FF0E";
          m(66) := x"FE6F";
          m(67) := x"FEEB";
          m(68) := x"FE3B";
          m(69) := x"FDE5";
          m(70) := x"FE45";
          m(71) := x"0061";
          m(72) := x"007C";
          m(73) := x"FEC6";
          m(74) := x"FEB6";
          m(75) := x"FE6E";
          m(76) := x"FF0D";
          m(77) := x"FF62";
          m(78) := x"FF9F";
          m(79) := x"FFB9";
          m(80) := x"FFDB";
          m(81) := x"FFCE";
          m(82) := x"002F";
          m(83) := x"000A";
          m(84) := x"FFE4";
          m(85) := x"FFC0";
          m(86) := x"002F";
          m(87) := x"0024";
          m(88) := x"FFF7";
          m(89) := x"FFEF";
          m(90) := x"FFB9";
          m(91) := x"FF07";
          m(92) := x"FD78";
          m(93) := x"FBAF";
          m(94) := x"FBF4";
          m(95) := x"FBD3";
          m(96) := x"FD43";
          m(97) := x"FCDB";
          m(98) := x"FCB3";
          m(99) := x"016A";
          m(100) := x"0112";
          m(101) := x"0018";
          m(102) := x"006E";
          m(103) := x"FEAE";
          m(104) := x"0008";
          m(105) := x"FEE7";
          m(106) := x"FEAC";
          m(107) := x"FF13";
          m(108) := x"FF5D";
          m(109) := x"FF5E";
          m(110) := x"FF56";
          m(111) := x"003E";
          m(112) := x"FFE6";
          m(113) := x"FFF2";
          m(114) := x"FFEE";
          m(115) := x"003B";
          m(116) := x"000B";
          m(117) := x"0001";
          m(118) := x"FEF8";
          m(119) := x"FCA4";
          m(120) := x"FC83";
          m(121) := x"FA22";
          m(122) := x"FB36";
          m(123) := x"FE14";
          m(124) := x"FD3A";
          m(125) := x"FE9A";
          m(126) := x"FCB3";
          m(127) := x"001C";
          m(128) := x"FE13";
          m(129) := x"FC26";
          m(130) := x"02C9";
          m(131) := x"0225";
          m(132) := x"01D0";
          m(133) := x"00C2";
          m(134) := x"FFD0";
          m(135) := x"FCC9";
          m(136) := x"FD86";
          m(137) := x"FEB5";
          m(138) := x"0025";
          m(139) := x"FFEC";
          m(140) := x"FFFE";
          m(141) := x"FFF5";
          m(142) := x"002D";
          m(143) := x"0022";
          m(144) := x"0126";
          m(145) := x"0338";
          m(146) := x"00F1";
          m(147) := x"FF3D";
          m(148) := x"FD8F";
          m(149) := x"FE95";
          m(150) := x"FECC";
          m(151) := x"FBA7";
          m(152) := x"FE38";
          m(153) := x"FC33";
          m(154) := x"FD1A";
          m(155) := x"FC88";
          m(156) := x"FD0D";
          m(157) := x"FADE";
          m(158) := x"FB6B";
          m(159) := x"03CA";
          m(160) := x"FDAB";
          m(161) := x"FB9D";
          m(162) := x"FDDA";
          m(163) := x"FC1E";
          m(164) := x"FDBE";
          m(165) := x"FE60";
          m(166) := x"FF90";
          m(167) := x"FFE4";
          m(168) := x"0036";
          m(169) := x"0030";
          m(170) := x"FFD9";
          m(171) := x"000A";
          m(172) := x"0172";
          m(173) := x"03ED";
          m(174) := x"0415";
          m(175) := x"FE92";
          m(176) := x"FF59";
          m(177) := x"028C";
          m(178) := x"02C5";
          m(179) := x"FF71";
          m(180) := x"FF69";
          m(181) := x"00FA";
          m(182) := x"FFB8";
          m(183) := x"FDF7";
          m(184) := x"0188";
          m(185) := x"0111";
          m(186) := x"01F1";
          m(187) := x"05D0";
          m(188) := x"038E";
          m(189) := x"FFB3";
          m(190) := x"01A1";
          m(191) := x"FF90";
          m(192) := x"FE69";
          m(193) := x"FF39";
          m(194) := x"FFB1";
          m(195) := x"FF95";
          m(196) := x"000D";
          m(197) := x"FFFF";
          m(198) := x"FF89";
          m(199) := x"008F";
          m(200) := x"0306";
          m(201) := x"04EF";
          m(202) := x"03CA";
          m(203) := x"0085";
          m(204) := x"0127";
          m(205) := x"00E7";
          m(206) := x"02F8";
          m(207) := x"FF12";
          m(208) := x"FDF1";
          m(209) := x"FFF6";
          m(210) := x"FFA7";
          m(211) := x"05EB";
          m(212) := x"01C3";
          m(213) := x"02F4";
          m(214) := x"039E";
          m(215) := x"0818";
          m(216) := x"0627";
          m(217) := x"FE27";
          m(218) := x"0162";
          m(219) := x"001B";
          m(220) := x"FE08";
          m(221) := x"FD70";
          m(222) := x"FFF8";
          m(223) := x"FFB6";
          m(224) := x"0013";
          m(225) := x"FFDB";
          m(226) := x"0010";
          m(227) := x"0135";
          m(228) := x"04CF";
          m(229) := x"04EB";
          m(230) := x"030E";
          m(231) := x"00C8";
          m(232) := x"01E7";
          m(233) := x"01CA";
          m(234) := x"FEF2";
          m(235) := x"FE10";
          m(236) := x"FB97";
          m(237) := x"FC8F";
          m(238) := x"0406";
          m(239) := x"0837";
          m(240) := x"032D";
          m(241) := x"036C";
          m(242) := x"05BD";
          m(243) := x"0175";
          m(244) := x"0300";
          m(245) := x"00C7";
          m(246) := x"0390";
          m(247) := x"FE08";
          m(248) := x"FDA1";
          m(249) := x"FEE8";
          m(250) := x"00C0";
          m(251) := x"0008";
          m(252) := x"0013";
          m(253) := x"0030";
          m(254) := x"003C";
          m(255) := x"01D1";
          m(256) := x"0307";
          m(257) := x"0132";
          m(258) := x"FFDF";
          m(259) := x"0000";
          m(260) := x"018F";
          m(261) := x"0076";
          m(262) := x"FDCC";
          m(263) := x"FDEC";
          m(264) := x"FC79";
          m(265) := x"FE3A";
          m(266) := x"FF66";
          m(267) := x"FE5F";
          m(268) := x"0466";
          m(269) := x"0195";
          m(270) := x"0330";
          m(271) := x"030B";
          m(272) := x"FF74";
          m(273) := x"0201";
          m(274) := x"0631";
          m(275) := x"0086";
          m(276) := x"FD93";
          m(277) := x"0204";
          m(278) := x"00F7";
          m(279) := x"013C";
          m(280) := x"FFEC";
          m(281) := x"FFDF";
          m(282) := x"004E";
          m(283) := x"0158";
          m(284) := x"FE53";
          m(285) := x"FB99";
          m(286) := x"FCB1";
          m(287) := x"0142";
          m(288) := x"019D";
          m(289) := x"029D";
          m(290) := x"01BB";
          m(291) := x"FF12";
          m(292) := x"0008";
          m(293) := x"FDCE";
          m(294) := x"FA66";
          m(295) := x"FD52";
          m(296) := x"FFD8";
          m(297) := x"0058";
          m(298) := x"052C";
          m(299) := x"02E0";
          m(300) := x"00C3";
          m(301) := x"FE51";
          m(302) := x"03DA";
          m(303) := x"0034";
          m(304) := x"FD6A";
          m(305) := x"00AA";
          m(306) := x"009C";
          m(307) := x"0007";
          m(308) := x"0005";
          m(309) := x"000B";
          m(310) := x"FFFA";
          m(311) := x"00F7";
          m(312) := x"FE99";
          m(313) := x"FC33";
          m(314) := x"FEA4";
          m(315) := x"008E";
          m(316) := x"05B8";
          m(317) := x"0268";
          m(318) := x"0032";
          m(319) := x"FDF8";
          m(320) := x"0152";
          m(321) := x"FF0A";
          m(322) := x"FE03";
          m(323) := x"FCAB";
          m(324) := x"FE96";
          m(325) := x"0071";
          m(326) := x"FEF4";
          m(327) := x"FA5A";
          m(328) := x"024E";
          m(329) := x"FF4C";
          m(330) := x"03B8";
          m(331) := x"FFB1";
          m(332) := x"FC4C";
          m(333) := x"FDD2";
          m(334) := x"0075";
          m(335) := x"001D";
          m(336) := x"0003";
          m(337) := x"FFDF";
          m(338) := x"FFF6";
          m(339) := x"FF24";
          m(340) := x"FE7B";
          m(341) := x"FF8F";
          m(342) := x"0312";
          m(343) := x"0231";
          m(344) := x"01E6";
          m(345) := x"FE12";
          m(346) := x"FEE6";
          m(347) := x"FA72";
          m(348) := x"066F";
          m(349) := x"0B17";
          m(350) := x"0A7A";
          m(351) := x"0833";
          m(352) := x"02F5";
          m(353) := x"FB0D";
          m(354) := x"0174";
          m(355) := x"0031";
          m(356) := x"0200";
          m(357) := x"01C2";
          m(358) := x"01B9";
          m(359) := x"FF84";
          m(360) := x"FBD6";
          m(361) := x"FEF1";
          m(362) := x"0079";
          m(363) := x"FFE5";
          m(364) := x"FFF5";
          m(365) := x"0032";
          m(366) := x"0068";
          m(367) := x"FF68";
          m(368) := x"FFE4";
          m(369) := x"FF4E";
          m(370) := x"017F";
          m(371) := x"FDC0";
          m(372) := x"FD55";
          m(373) := x"FD5A";
          m(374) := x"0011";
          m(375) := x"0140";
          m(376) := x"0665";
          m(377) := x"0A96";
          m(378) := x"0312";
          m(379) := x"06FE";
          m(380) := x"06D0";
          m(381) := x"035B";
          m(382) := x"074D";
          m(383) := x"01AF";
          m(384) := x"0084";
          m(385) := x"017F";
          m(386) := x"FD20";
          m(387) := x"FD36";
          m(388) := x"FD24";
          m(389) := x"FF68";
          m(390) := x"FFAA";
          m(391) := x"FF73";
          m(392) := x"FFEE";
          m(393) := x"0070";
          m(394) := x"0058";
          m(395) := x"FFD9";
          m(396) := x"FE66";
          m(397) := x"00DA";
          m(398) := x"00D6";
          m(399) := x"0028";
          m(400) := x"0275";
          m(401) := x"FD95";
          m(402) := x"FDE1";
          m(403) := x"FB2D";
          m(404) := x"0659";
          m(405) := x"06E6";
          m(406) := x"07A6";
          m(407) := x"04B5";
          m(408) := x"03B7";
          m(409) := x"043F";
          m(410) := x"0317";
          m(411) := x"033F";
          m(412) := x"0014";
          m(413) := x"FF96";
          m(414) := x"FDB5";
          m(415) := x"FDC1";
          m(416) := x"FCC1";
          m(417) := x"FE7E";
          m(418) := x"003E";
          m(419) := x"FFEA";
          m(420) := x"FFE5";
          m(421) := x"00D3";
          m(422) := x"009D";
          m(423) := x"0001";
          m(424) := x"FDEB";
          m(425) := x"FE7C";
          m(426) := x"FC51";
          m(427) := x"FF8E";
          m(428) := x"FE19";
          m(429) := x"FB68";
          m(430) := x"F9B6";
          m(431) := x"FC42";
          m(432) := x"03D7";
          m(433) := x"0594";
          m(434) := x"05F2";
          m(435) := x"029E";
          m(436) := x"0476";
          m(437) := x"02B9";
          m(438) := x"FE24";
          m(439) := x"FE3A";
          m(440) := x"00E9";
          m(441) := x"0009";
          m(442) := x"03C5";
          m(443) := x"FF54";
          m(444) := x"FDB2";
          m(445) := x"FDCD";
          m(446) := x"002E";
          m(447) := x"FFFB";
          m(448) := x"0022";
          m(449) := x"004C";
          m(450) := x"00CC";
          m(451) := x"001F";
          m(452) := x"022C";
          m(453) := x"FBCE";
          m(454) := x"F8FA";
          m(455) := x"FE3F";
          m(456) := x"F7CF";
          m(457) := x"F80D";
          m(458) := x"FAD4";
          m(459) := x"F67E";
          m(460) := x"0082";
          m(461) := x"05C6";
          m(462) := x"0083";
          m(463) := x"04F6";
          m(464) := x"0276";
          m(465) := x"0042";
          m(466) := x"0094";
          m(467) := x"009B";
          m(468) := x"FCE8";
          m(469) := x"FDE1";
          m(470) := x"01BB";
          m(471) := x"FD48";
          m(472) := x"FC44";
          m(473) := x"FCBC";
          m(474) := x"FFED";
          m(475) := x"0013";
          m(476) := x"FFD7";
          m(477) := x"FFE9";
          m(478) := x"00DC";
          m(479) := x"0194";
          m(480) := x"0081";
          m(481) := x"FA7D";
          m(482) := x"F62B";
          m(483) := x"FAF5";
          m(484) := x"F965";
          m(485) := x"F95C";
          m(486) := x"F346";
          m(487) := x"F307";
          m(488) := x"FAB1";
          m(489) := x"007A";
          m(490) := x"00BC";
          m(491) := x"FCCA";
          m(492) := x"0276";
          m(493) := x"028A";
          m(494) := x"087D";
          m(495) := x"00C4";
          m(496) := x"FA92";
          m(497) := x"FFFD";
          m(498) := x"01AF";
          m(499) := x"0013";
          m(500) := x"FA6F";
          m(501) := x"FDA8";
          m(502) := x"0036";
          m(503) := x"FFB8";
          m(504) := x"000D";
          m(505) := x"FFC1";
          m(506) := x"00BF";
          m(507) := x"00E2";
          m(508) := x"0002";
          m(509) := x"FA0D";
          m(510) := x"F755";
          m(511) := x"F9BC";
          m(512) := x"FDDA";
          m(513) := x"FB7C";
          m(514) := x"F74D";
          m(515) := x"F796";
          m(516) := x"FA64";
          m(517) := x"001A";
          m(518) := x"FB5F";
          m(519) := x"FA51";
          m(520) := x"0014";
          m(521) := x"04E2";
          m(522) := x"03D5";
          m(523) := x"0035";
          m(524) := x"FEF6";
          m(525) := x"014F";
          m(526) := x"FE7F";
          m(527) := x"FC2A";
          m(528) := x"F9ED";
          m(529) := x"FEB8";
          m(530) := x"0014";
          m(531) := x"FFF3";
          m(532) := x"FFFA";
          m(533) := x"0013";
          m(534) := x"002A";
          m(535) := x"FECF";
          m(536) := x"004C";
          m(537) := x"0069";
          m(538) := x"FACC";
          m(539) := x"FEBD";
          m(540) := x"0082";
          m(541) := x"FC19";
          m(542) := x"FCF8";
          m(543) := x"FF1B";
          m(544) := x"0358";
          m(545) := x"FDEA";
          m(546) := x"F746";
          m(547) := x"F93B";
          m(548) := x"00DF";
          m(549) := x"0588";
          m(550) := x"008A";
          m(551) := x"0144";
          m(552) := x"01C9";
          m(553) := x"0235";
          m(554) := x"FE17";
          m(555) := x"FA06";
          m(556) := x"FDA9";
          m(557) := x"FF73";
          m(558) := x"FFCB";
          m(559) := x"FFD0";
          m(560) := x"FFEF";
          m(561) := x"0000";
          m(562) := x"FF50";
          m(563) := x"FCE5";
          m(564) := x"FEFC";
          m(565) := x"FF1B";
          m(566) := x"FB83";
          m(567) := x"FE20";
          m(568) := x"0117";
          m(569) := x"F7FA";
          m(570) := x"F460";
          m(571) := x"025E";
          m(572) := x"02EA";
          m(573) := x"0218";
          m(574) := x"0677";
          m(575) := x"FB57";
          m(576) := x"FF04";
          m(577) := x"FE6E";
          m(578) := x"FF54";
          m(579) := x"02B1";
          m(580) := x"01E3";
          m(581) := x"FCCF";
          m(582) := x"FD13";
          m(583) := x"FAC9";
          m(584) := x"FE87";
          m(585) := x"FF27";
          m(586) := x"FFE6";
          m(587) := x"0000";
          m(588) := x"FFE6";
          m(589) := x"000A";
          m(590) := x"FEC0";
          m(591) := x"FCD3";
          m(592) := x"FECD";
          m(593) := x"FF89";
          m(594) := x"FD01";
          m(595) := x"FC59";
          m(596) := x"0017";
          m(597) := x"F717";
          m(598) := x"FB80";
          m(599) := x"FE59";
          m(600) := x"FE9A";
          m(601) := x"024B";
          m(602) := x"051C";
          m(603) := x"FC71";
          m(604) := x"FF0D";
          m(605) := x"FC8B";
          m(606) := x"008A";
          m(607) := x"0380";
          m(608) := x"0094";
          m(609) := x"FB18";
          m(610) := x"FA9F";
          m(611) := x"F9C3";
          m(612) := x"FF3D";
          m(613) := x"FF59";
          m(614) := x"FFAF";
          m(615) := x"000D";
          m(616) := x"FFFB";
          m(617) := x"0008";
          m(618) := x"FE8C";
          m(619) := x"FD89";
          m(620) := x"FFB1";
          m(621) := x"01ED";
          m(622) := x"FF97";
          m(623) := x"FC2A";
          m(624) := x"FC4A";
          m(625) := x"F9E9";
          m(626) := x"F7A3";
          m(627) := x"F9ED";
          m(628) := x"FB28";
          m(629) := x"00F3";
          m(630) := x"0065";
          m(631) := x"FF7C";
          m(632) := x"FF90";
          m(633) := x"03BB";
          m(634) := x"026C";
          m(635) := x"0505";
          m(636) := x"FECD";
          m(637) := x"FC14";
          m(638) := x"FC5F";
          m(639) := x"FB29";
          m(640) := x"FE52";
          m(641) := x"FFB5";
          m(642) := x"FFFB";
          m(643) := x"FFFC";
          m(644) := x"FFE6";
          m(645) := x"0026";
          m(646) := x"0019";
          m(647) := x"FFA2";
          m(648) := x"01CC";
          m(649) := x"02F5";
          m(650) := x"FFA2";
          m(651) := x"0002";
          m(652) := x"FDDA";
          m(653) := x"FDD4";
          m(654) := x"FEBA";
          m(655) := x"011A";
          m(656) := x"FDCC";
          m(657) := x"FEEF";
          m(658) := x"FF20";
          m(659) := x"0116";
          m(660) := x"0273";
          m(661) := x"0524";
          m(662) := x"0070";
          m(663) := x"FCC4";
          m(664) := x"FFA7";
          m(665) := x"FE9A";
          m(666) := x"FC03";
          m(667) := x"FC5D";
          m(668) := x"FEAB";
          m(669) := x"FF35";
          m(670) := x"0006";
          m(671) := x"0000";
          m(672) := x"0005";
          m(673) := x"0014";
          m(674) := x"005A";
          m(675) := x"008B";
          m(676) := x"02BC";
          m(677) := x"03F8";
          m(678) := x"020C";
          m(679) := x"02AD";
          m(680) := x"FF7C";
          m(681) := x"FF35";
          m(682) := x"0146";
          m(683) := x"0090";
          m(684) := x"FFE5";
          m(685) := x"FFD6";
          m(686) := x"FE3B";
          m(687) := x"FF9E";
          m(688) := x"02AB";
          m(689) := x"06AF";
          m(690) := x"0377";
          m(691) := x"01DD";
          m(692) := x"026A";
          m(693) := x"00CC";
          m(694) := x"FE7A";
          m(695) := x"FE9B";
          m(696) := x"FE0B";
          m(697) := x"FEE9";
          m(698) := x"FFB2";
          m(699) := x"0000";
          m(700) := x"FFE7";
          m(701) := x"FFF8";
          m(702) := x"0020";
          m(703) := x"0011";
          m(704) := x"00ED";
          m(705) := x"01D7";
          m(706) := x"017B";
          m(707) := x"0247";
          m(708) := x"044F";
          m(709) := x"06EA";
          m(710) := x"049B";
          m(711) := x"054D";
          m(712) := x"07CF";
          m(713) := x"056F";
          m(714) := x"03DC";
          m(715) := x"0221";
          m(716) := x"FF23";
          m(717) := x"FFB9";
          m(718) := x"0209";
          m(719) := x"0335";
          m(720) := x"0265";
          m(721) := x"00F8";
          m(722) := x"008E";
          m(723) := x"FFA9";
          m(724) := x"FFB4";
          m(725) := x"FFA7";
          m(726) := x"FF9F";
          m(727) := x"001E";
          m(728) := x"0024";
          m(729) := x"FFEF";
          m(730) := x"000F";
          m(731) := x"FFFA";
          m(732) := x"FFE9";
          m(733) := x"0041";
          m(734) := x"0073";
          m(735) := x"0187";
          m(736) := x"0106";
          m(737) := x"0224";
          m(738) := x"01C0";
          m(739) := x"005F";
          m(740) := x"FEDF";
          m(741) := x"0029";
          m(742) := x"01A8";
          m(743) := x"00C8";
          m(744) := x"00EA";
          m(745) := x"FFD7";
          m(746) := x"01B5";
          m(747) := x"0132";
          m(748) := x"0051";
          m(749) := x"00DF";
          m(750) := x"008A";
          m(751) := x"0002";
          m(752) := x"FFF2";
          m(753) := x"FFF2";
          m(754) := x"000A";
          m(755) := x"FFBC";
          m(756) := x"FFF0";
          m(757) := x"000C";
          m(758) := x"FFF7";
          m(759) := x"FFF2";
          m(760) := x"000C";
          m(761) := x"FFF9";
          m(762) := x"FFF4";
          m(763) := x"FFDA";
          m(764) := x"FFD9";
          m(765) := x"0006";
          m(766) := x"000F";
          m(767) := x"FFF4";
          m(768) := x"FFEE";
          m(769) := x"000F";
          m(770) := x"0017";
          m(771) := x"001C";
          m(772) := x"00A5";
          m(773) := x"0047";
          m(774) := x"00B8";
          m(775) := x"0020";
          m(776) := x"0020";
          m(777) := x"000C";
          m(778) := x"0023";
          m(779) := x"001A";
          m(780) := x"0021";
          m(781) := x"FFD2";
          m(782) := x"FFE6";
          m(783) := x"0010";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_18.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 18) then
          m(0) := x"FFDF";
          m(1) := x"FFA9";
          m(2) := x"000D";
          m(3) := x"FFF3";
          m(4) := x"FFFD";
          m(5) := x"000B";
          m(6) := x"FFF5";
          m(7) := x"0019";
          m(8) := x"001F";
          m(9) := x"0000";
          m(10) := x"FFE5";
          m(11) := x"0008";
          m(12) := x"FFDE";
          m(13) := x"FFE2";
          m(14) := x"004B";
          m(15) := x"FFF0";
          m(16) := x"FFFA";
          m(17) := x"0063";
          m(18) := x"FFF9";
          m(19) := x"FFFE";
          m(20) := x"001B";
          m(21) := x"0001";
          m(22) := x"0033";
          m(23) := x"0020";
          m(24) := x"0002";
          m(25) := x"0007";
          m(26) := x"0012";
          m(27) := x"000D";
          m(28) := x"FFCA";
          m(29) := x"0028";
          m(30) := x"FFFD";
          m(31) := x"001D";
          m(32) := x"0037";
          m(33) := x"FFFC";
          m(34) := x"FFF5";
          m(35) := x"FFE9";
          m(36) := x"0016";
          m(37) := x"FFFD";
          m(38) := x"000E";
          m(39) := x"0005";
          m(40) := x"0067";
          m(41) := x"0009";
          m(42) := x"001A";
          m(43) := x"0041";
          m(44) := x"0031";
          m(45) := x"005C";
          m(46) := x"FFFA";
          m(47) := x"001D";
          m(48) := x"0044";
          m(49) := x"0034";
          m(50) := x"001E";
          m(51) := x"0015";
          m(52) := x"FFDD";
          m(53) := x"FFF3";
          m(54) := x"FFFF";
          m(55) := x"FFF1";
          m(56) := x"0000";
          m(57) := x"FFF9";
          m(58) := x"0014";
          m(59) := x"000D";
          m(60) := x"000D";
          m(61) := x"FFFD";
          m(62) := x"0013";
          m(63) := x"0073";
          m(64) := x"007E";
          m(65) := x"0059";
          m(66) := x"00D5";
          m(67) := x"00C6";
          m(68) := x"00FA";
          m(69) := x"0146";
          m(70) := x"00CB";
          m(71) := x"012D";
          m(72) := x"0169";
          m(73) := x"010C";
          m(74) := x"012E";
          m(75) := x"00D5";
          m(76) := x"0067";
          m(77) := x"0022";
          m(78) := x"FFF0";
          m(79) := x"0019";
          m(80) := x"0024";
          m(81) := x"FFFF";
          m(82) := x"FFF9";
          m(83) := x"004C";
          m(84) := x"FFF0";
          m(85) := x"000B";
          m(86) := x"FFE5";
          m(87) := x"FFEF";
          m(88) := x"0022";
          m(89) := x"009B";
          m(90) := x"009B";
          m(91) := x"0118";
          m(92) := x"02DF";
          m(93) := x"01DB";
          m(94) := x"0023";
          m(95) := x"FE15";
          m(96) := x"028C";
          m(97) := x"0493";
          m(98) := x"013D";
          m(99) := x"0342";
          m(100) := x"044F";
          m(101) := x"0336";
          m(102) := x"03F5";
          m(103) := x"02B0";
          m(104) := x"0051";
          m(105) := x"FFC2";
          m(106) := x"FFD3";
          m(107) := x"0056";
          m(108) := x"0075";
          m(109) := x"004A";
          m(110) := x"FFE8";
          m(111) := x"FFFF";
          m(112) := x"FFE1";
          m(113) := x"FFB1";
          m(114) := x"FFF6";
          m(115) := x"0015";
          m(116) := x"0058";
          m(117) := x"01AC";
          m(118) := x"020F";
          m(119) := x"02FD";
          m(120) := x"04B5";
          m(121) := x"02A0";
          m(122) := x"0409";
          m(123) := x"0279";
          m(124) := x"0170";
          m(125) := x"040B";
          m(126) := x"0322";
          m(127) := x"0394";
          m(128) := x"02C6";
          m(129) := x"FF51";
          m(130) := x"0304";
          m(131) := x"0577";
          m(132) := x"03FD";
          m(133) := x"0451";
          m(134) := x"01EB";
          m(135) := x"FF3D";
          m(136) := x"FEFC";
          m(137) := x"FF8F";
          m(138) := x"003F";
          m(139) := x"000B";
          m(140) := x"FFFB";
          m(141) := x"FFD8";
          m(142) := x"0021";
          m(143) := x"002B";
          m(144) := x"0124";
          m(145) := x"02D9";
          m(146) := x"0458";
          m(147) := x"06A3";
          m(148) := x"0355";
          m(149) := x"01B5";
          m(150) := x"0246";
          m(151) := x"04AB";
          m(152) := x"0158";
          m(153) := x"02EA";
          m(154) := x"FED1";
          m(155) := x"02EE";
          m(156) := x"0466";
          m(157) := x"093D";
          m(158) := x"07B2";
          m(159) := x"0A19";
          m(160) := x"07ED";
          m(161) := x"033B";
          m(162) := x"037B";
          m(163) := x"010F";
          m(164) := x"FFA9";
          m(165) := x"007E";
          m(166) := x"0026";
          m(167) := x"FFD1";
          m(168) := x"001F";
          m(169) := x"FFF8";
          m(170) := x"FF9E";
          m(171) := x"005E";
          m(172) := x"014A";
          m(173) := x"00FE";
          m(174) := x"04A8";
          m(175) := x"07F0";
          m(176) := x"0402";
          m(177) := x"05A0";
          m(178) := x"04A2";
          m(179) := x"065B";
          m(180) := x"053C";
          m(181) := x"061C";
          m(182) := x"06E1";
          m(183) := x"0DCC";
          m(184) := x"0CB7";
          m(185) := x"0BED";
          m(186) := x"08CD";
          m(187) := x"02EF";
          m(188) := x"0268";
          m(189) := x"FCEC";
          m(190) := x"FD13";
          m(191) := x"FEC0";
          m(192) := x"FF6F";
          m(193) := x"00A0";
          m(194) := x"0017";
          m(195) := x"0043";
          m(196) := x"FFDB";
          m(197) := x"0030";
          m(198) := x"FF5B";
          m(199) := x"FF76";
          m(200) := x"01DF";
          m(201) := x"00A3";
          m(202) := x"0332";
          m(203) := x"02D2";
          m(204) := x"021F";
          m(205) := x"027E";
          m(206) := x"05AB";
          m(207) := x"04BB";
          m(208) := x"0BA8";
          m(209) := x"0942";
          m(210) := x"0AEE";
          m(211) := x"0626";
          m(212) := x"0071";
          m(213) := x"FA4D";
          m(214) := x"FC76";
          m(215) := x"FB4B";
          m(216) := x"F908";
          m(217) := x"F892";
          m(218) := x"F9CC";
          m(219) := x"FB7C";
          m(220) := x"FEA1";
          m(221) := x"FEF5";
          m(222) := x"FEE0";
          m(223) := x"0014";
          m(224) := x"0007";
          m(225) := x"FFED";
          m(226) := x"FF2B";
          m(227) := x"FF74";
          m(228) := x"0008";
          m(229) := x"019F";
          m(230) := x"0010";
          m(231) := x"FD80";
          m(232) := x"013E";
          m(233) := x"0767";
          m(234) := x"0955";
          m(235) := x"0402";
          m(236) := x"0535";
          m(237) := x"01DD";
          m(238) := x"001B";
          m(239) := x"FB79";
          m(240) := x"F6A7";
          m(241) := x"F845";
          m(242) := x"FA98";
          m(243) := x"00CB";
          m(244) := x"FA1F";
          m(245) := x"FD39";
          m(246) := x"FD50";
          m(247) := x"FA14";
          m(248) := x"FAA0";
          m(249) := x"FF06";
          m(250) := x"006C";
          m(251) := x"0042";
          m(252) := x"0004";
          m(253) := x"FFD3";
          m(254) := x"FFBB";
          m(255) := x"FF8B";
          m(256) := x"010F";
          m(257) := x"0017";
          m(258) := x"00C0";
          m(259) := x"01B9";
          m(260) := x"FFE3";
          m(261) := x"01C4";
          m(262) := x"FB6C";
          m(263) := x"FF05";
          m(264) := x"FD44";
          m(265) := x"F79D";
          m(266) := x"F8C3";
          m(267) := x"F822";
          m(268) := x"F4E9";
          m(269) := x"FB4E";
          m(270) := x"FB7F";
          m(271) := x"FE4F";
          m(272) := x"FB4F";
          m(273) := x"FDF8";
          m(274) := x"FFA1";
          m(275) := x"FAA6";
          m(276) := x"FB87";
          m(277) := x"010B";
          m(278) := x"0000";
          m(279) := x"FFC4";
          m(280) := x"FFF2";
          m(281) := x"FFE0";
          m(282) := x"FFF9";
          m(283) := x"FFCB";
          m(284) := x"FFF5";
          m(285) := x"0023";
          m(286) := x"FF2B";
          m(287) := x"FBAB";
          m(288) := x"FB10";
          m(289) := x"F992";
          m(290) := x"F861";
          m(291) := x"FA90";
          m(292) := x"F7E4";
          m(293) := x"FC41";
          m(294) := x"FC2F";
          m(295) := x"F914";
          m(296) := x"013F";
          m(297) := x"FF11";
          m(298) := x"FEC8";
          m(299) := x"0154";
          m(300) := x"004C";
          m(301) := x"001B";
          m(302) := x"00DA";
          m(303) := x"FC82";
          m(304) := x"FC86";
          m(305) := x"FF26";
          m(306) := x"0000";
          m(307) := x"FFD1";
          m(308) := x"0021";
          m(309) := x"FFF1";
          m(310) := x"0023";
          m(311) := x"003E";
          m(312) := x"01DE";
          m(313) := x"022E";
          m(314) := x"028C";
          m(315) := x"FACD";
          m(316) := x"F936";
          m(317) := x"F817";
          m(318) := x"F9A3";
          m(319) := x"FD7B";
          m(320) := x"F9E7";
          m(321) := x"016C";
          m(322) := x"0503";
          m(323) := x"03C2";
          m(324) := x"079F";
          m(325) := x"02AC";
          m(326) := x"016C";
          m(327) := x"FD06";
          m(328) := x"FDE7";
          m(329) := x"0056";
          m(330) := x"013C";
          m(331) := x"FFEB";
          m(332) := x"FF99";
          m(333) := x"00CE";
          m(334) := x"0145";
          m(335) := x"0029";
          m(336) := x"001A";
          m(337) := x"0000";
          m(338) := x"FFAD";
          m(339) := x"FFB1";
          m(340) := x"025B";
          m(341) := x"01D7";
          m(342) := x"01C1";
          m(343) := x"FDE9";
          m(344) := x"FA86";
          m(345) := x"FA5F";
          m(346) := x"FC62";
          m(347) := x"F983";
          m(348) := x"F802";
          m(349) := x"FDC0";
          m(350) := x"0653";
          m(351) := x"FFEE";
          m(352) := x"03B7";
          m(353) := x"0629";
          m(354) := x"0212";
          m(355) := x"FCE3";
          m(356) := x"FCAB";
          m(357) := x"FC50";
          m(358) := x"FD2B";
          m(359) := x"0132";
          m(360) := x"FF88";
          m(361) := x"0015";
          m(362) := x"FFD0";
          m(363) := x"0025";
          m(364) := x"001B";
          m(365) := x"FFF6";
          m(366) := x"FF81";
          m(367) := x"FF73";
          m(368) := x"FE49";
          m(369) := x"FE03";
          m(370) := x"0060";
          m(371) := x"FEAA";
          m(372) := x"FEAA";
          m(373) := x"0043";
          m(374) := x"F7F1";
          m(375) := x"F6F2";
          m(376) := x"F957";
          m(377) := x"0008";
          m(378) := x"0389";
          m(379) := x"0038";
          m(380) := x"043C";
          m(381) := x"02D8";
          m(382) := x"03DD";
          m(383) := x"FCBC";
          m(384) := x"FE4D";
          m(385) := x"FD36";
          m(386) := x"FD90";
          m(387) := x"0018";
          m(388) := x"FE88";
          m(389) := x"FDFA";
          m(390) := x"FF42";
          m(391) := x"FFFF";
          m(392) := x"FFBA";
          m(393) := x"FFBA";
          m(394) := x"FF84";
          m(395) := x"FFF1";
          m(396) := x"FF16";
          m(397) := x"FB98";
          m(398) := x"02CD";
          m(399) := x"0221";
          m(400) := x"FBA8";
          m(401) := x"FAC6";
          m(402) := x"F9EF";
          m(403) := x"F4B1";
          m(404) := x"F5D6";
          m(405) := x"0316";
          m(406) := x"0666";
          m(407) := x"0320";
          m(408) := x"0236";
          m(409) := x"FA5B";
          m(410) := x"01ED";
          m(411) := x"FF20";
          m(412) := x"FEBA";
          m(413) := x"FEA1";
          m(414) := x"FC54";
          m(415) := x"FEA0";
          m(416) := x"FFF3";
          m(417) := x"FFD6";
          m(418) := x"0005";
          m(419) := x"000A";
          m(420) := x"0053";
          m(421) := x"FFEA";
          m(422) := x"FF6F";
          m(423) := x"FFD8";
          m(424) := x"00EC";
          m(425) := x"FFBE";
          m(426) := x"0287";
          m(427) := x"FF24";
          m(428) := x"012F";
          m(429) := x"FCE6";
          m(430) := x"FB01";
          m(431) := x"0008";
          m(432) := x"F75F";
          m(433) := x"FF94";
          m(434) := x"04E6";
          m(435) := x"FFA0";
          m(436) := x"02DC";
          m(437) := x"FDE5";
          m(438) := x"0033";
          m(439) := x"FF83";
          m(440) := x"FD66";
          m(441) := x"FF8D";
          m(442) := x"0076";
          m(443) := x"FF0F";
          m(444) := x"0027";
          m(445) := x"00A5";
          m(446) := x"FF2A";
          m(447) := x"002B";
          m(448) := x"FFEF";
          m(449) := x"0001";
          m(450) := x"0000";
          m(451) := x"0180";
          m(452) := x"02A1";
          m(453) := x"FF5A";
          m(454) := x"0072";
          m(455) := x"FE0E";
          m(456) := x"FD02";
          m(457) := x"FF42";
          m(458) := x"0020";
          m(459) := x"FECA";
          m(460) := x"FB98";
          m(461) := x"FFB5";
          m(462) := x"02F4";
          m(463) := x"FF3E";
          m(464) := x"FCFE";
          m(465) := x"F8E6";
          m(466) := x"FE52";
          m(467) := x"FD27";
          m(468) := x"FE47";
          m(469) := x"0010";
          m(470) := x"FF3A";
          m(471) := x"FE69";
          m(472) := x"FFDD";
          m(473) := x"005E";
          m(474) := x"FF2F";
          m(475) := x"FFF3";
          m(476) := x"0005";
          m(477) := x"FFBF";
          m(478) := x"0034";
          m(479) := x"02DD";
          m(480) := x"030D";
          m(481) := x"FF94";
          m(482) := x"00AD";
          m(483) := x"FFDD";
          m(484) := x"FD27";
          m(485) := x"F937";
          m(486) := x"FD33";
          m(487) := x"FE6B";
          m(488) := x"001A";
          m(489) := x"FE6A";
          m(490) := x"0195";
          m(491) := x"02E5";
          m(492) := x"FBA0";
          m(493) := x"0068";
          m(494) := x"0139";
          m(495) := x"FC9D";
          m(496) := x"FD11";
          m(497) := x"FFFF";
          m(498) := x"FC6E";
          m(499) := x"FD27";
          m(500) := x"FD7A";
          m(501) := x"FF44";
          m(502) := x"FF6E";
          m(503) := x"FFF4";
          m(504) := x"0000";
          m(505) := x"FFFD";
          m(506) := x"0054";
          m(507) := x"0341";
          m(508) := x"0289";
          m(509) := x"FE95";
          m(510) := x"FFD6";
          m(511) := x"03F4";
          m(512) := x"0004";
          m(513) := x"FD22";
          m(514) := x"FAEC";
          m(515) := x"FE08";
          m(516) := x"FE93";
          m(517) := x"FE95";
          m(518) := x"FF7D";
          m(519) := x"FEA9";
          m(520) := x"0492";
          m(521) := x"03B4";
          m(522) := x"039C";
          m(523) := x"FE3D";
          m(524) := x"0171";
          m(525) := x"FEF2";
          m(526) := x"FFA6";
          m(527) := x"0040";
          m(528) := x"FF4E";
          m(529) := x"FFF3";
          m(530) := x"FF91";
          m(531) := x"000D";
          m(532) := x"0044";
          m(533) := x"0027";
          m(534) := x"0018";
          m(535) := x"0226";
          m(536) := x"020F";
          m(537) := x"FE66";
          m(538) := x"0154";
          m(539) := x"0493";
          m(540) := x"02BD";
          m(541) := x"03DF";
          m(542) := x"FFE3";
          m(543) := x"0270";
          m(544) := x"0163";
          m(545) := x"05A0";
          m(546) := x"0413";
          m(547) := x"FF05";
          m(548) := x"0633";
          m(549) := x"0200";
          m(550) := x"0185";
          m(551) := x"0095";
          m(552) := x"012E";
          m(553) := x"FED6";
          m(554) := x"02DA";
          m(555) := x"01A7";
          m(556) := x"0166";
          m(557) := x"005A";
          m(558) := x"0021";
          m(559) := x"0009";
          m(560) := x"FFDF";
          m(561) := x"000F";
          m(562) := x"0050";
          m(563) := x"01EA";
          m(564) := x"0221";
          m(565) := x"FFD6";
          m(566) := x"0018";
          m(567) := x"0434";
          m(568) := x"0902";
          m(569) := x"0655";
          m(570) := x"02A5";
          m(571) := x"0171";
          m(572) := x"FEFA";
          m(573) := x"01ED";
          m(574) := x"031F";
          m(575) := x"FFD0";
          m(576) := x"02BF";
          m(577) := x"FC64";
          m(578) := x"02BE";
          m(579) := x"0401";
          m(580) := x"0374";
          m(581) := x"0365";
          m(582) := x"04CF";
          m(583) := x"0265";
          m(584) := x"0183";
          m(585) := x"0026";
          m(586) := x"0038";
          m(587) := x"0008";
          m(588) := x"0015";
          m(589) := x"0005";
          m(590) := x"0066";
          m(591) := x"0222";
          m(592) := x"01A1";
          m(593) := x"022C";
          m(594) := x"024E";
          m(595) := x"0320";
          m(596) := x"0631";
          m(597) := x"06F1";
          m(598) := x"0342";
          m(599) := x"0123";
          m(600) := x"0140";
          m(601) := x"0338";
          m(602) := x"0622";
          m(603) := x"03C4";
          m(604) := x"06FE";
          m(605) := x"01DF";
          m(606) := x"03E5";
          m(607) := x"0173";
          m(608) := x"043A";
          m(609) := x"038F";
          m(610) := x"00BB";
          m(611) := x"02AB";
          m(612) := x"0263";
          m(613) := x"0057";
          m(614) := x"FFAB";
          m(615) := x"FFEB";
          m(616) := x"FFED";
          m(617) := x"0009";
          m(618) := x"0004";
          m(619) := x"00EF";
          m(620) := x"03E3";
          m(621) := x"03ED";
          m(622) := x"02CA";
          m(623) := x"0401";
          m(624) := x"02FA";
          m(625) := x"05EC";
          m(626) := x"01DE";
          m(627) := x"FBB6";
          m(628) := x"FB97";
          m(629) := x"036E";
          m(630) := x"05FE";
          m(631) := x"003C";
          m(632) := x"05CC";
          m(633) := x"0305";
          m(634) := x"007D";
          m(635) := x"FF43";
          m(636) := x"04FD";
          m(637) := x"FF5A";
          m(638) := x"FFD8";
          m(639) := x"0304";
          m(640) := x"0204";
          m(641) := x"00C9";
          m(642) := x"0009";
          m(643) := x"FFF9";
          m(644) := x"0011";
          m(645) := x"0007";
          m(646) := x"FFF6";
          m(647) := x"003E";
          m(648) := x"0285";
          m(649) := x"03E5";
          m(650) := x"03AB";
          m(651) := x"0379";
          m(652) := x"02A7";
          m(653) := x"0256";
          m(654) := x"00D4";
          m(655) := x"FB60";
          m(656) := x"FE2D";
          m(657) := x"01E4";
          m(658) := x"FE1F";
          m(659) := x"01F8";
          m(660) := x"046D";
          m(661) := x"02A9";
          m(662) := x"0204";
          m(663) := x"0083";
          m(664) := x"0352";
          m(665) := x"000A";
          m(666) := x"0257";
          m(667) := x"0236";
          m(668) := x"0193";
          m(669) := x"001D";
          m(670) := x"0038";
          m(671) := x"FFC2";
          m(672) := x"0036";
          m(673) := x"FFED";
          m(674) := x"0040";
          m(675) := x"0009";
          m(676) := x"00D4";
          m(677) := x"018B";
          m(678) := x"04FD";
          m(679) := x"05EC";
          m(680) := x"0473";
          m(681) := x"01BC";
          m(682) := x"0199";
          m(683) := x"020A";
          m(684) := x"01F2";
          m(685) := x"01B2";
          m(686) := x"03D3";
          m(687) := x"0686";
          m(688) := x"0018";
          m(689) := x"007E";
          m(690) := x"FF94";
          m(691) := x"FF0D";
          m(692) := x"FF2A";
          m(693) := x"FF16";
          m(694) := x"FEDC";
          m(695) := x"0109";
          m(696) := x"0092";
          m(697) := x"FFF8";
          m(698) := x"0049";
          m(699) := x"0012";
          m(700) := x"FFF9";
          m(701) := x"FFE3";
          m(702) := x"0001";
          m(703) := x"FFD1";
          m(704) := x"FFFE";
          m(705) := x"0167";
          m(706) := x"02D1";
          m(707) := x"02D4";
          m(708) := x"0457";
          m(709) := x"020A";
          m(710) := x"FFA2";
          m(711) := x"FE4D";
          m(712) := x"02AF";
          m(713) := x"0162";
          m(714) := x"FF65";
          m(715) := x"028F";
          m(716) := x"02CC";
          m(717) := x"0072";
          m(718) := x"01F0";
          m(719) := x"04D1";
          m(720) := x"0212";
          m(721) := x"FFD5";
          m(722) := x"FF0A";
          m(723) := x"0009";
          m(724) := x"0020";
          m(725) := x"0001";
          m(726) := x"FFFA";
          m(727) := x"0056";
          m(728) := x"0036";
          m(729) := x"002D";
          m(730) := x"FFF5";
          m(731) := x"FFE3";
          m(732) := x"FFF5";
          m(733) := x"FFD8";
          m(734) := x"FFEB";
          m(735) := x"FF34";
          m(736) := x"FEFF";
          m(737) := x"FF4A";
          m(738) := x"0078";
          m(739) := x"FF66";
          m(740) := x"FF61";
          m(741) := x"0068";
          m(742) := x"00B5";
          m(743) := x"02A7";
          m(744) := x"035F";
          m(745) := x"0366";
          m(746) := x"02BC";
          m(747) := x"02D7";
          m(748) := x"00F9";
          m(749) := x"FFFE";
          m(750) := x"001B";
          m(751) := x"FFEB";
          m(752) := x"0032";
          m(753) := x"0028";
          m(754) := x"000E";
          m(755) := x"FFF3";
          m(756) := x"0016";
          m(757) := x"0022";
          m(758) := x"FFD3";
          m(759) := x"001A";
          m(760) := x"FFEC";
          m(761) := x"FFDA";
          m(762) := x"FFED";
          m(763) := x"0002";
          m(764) := x"0033";
          m(765) := x"FFE3";
          m(766) := x"FFAC";
          m(767) := x"FFD1";
          m(768) := x"0017";
          m(769) := x"FFE3";
          m(770) := x"FFE0";
          m(771) := x"0005";
          m(772) := x"0026";
          m(773) := x"FFFE";
          m(774) := x"0013";
          m(775) := x"0014";
          m(776) := x"0017";
          m(777) := x"FFCE";
          m(778) := x"0027";
          m(779) := x"FFDA";
          m(780) := x"FFF0";
          m(781) := x"0008";
          m(782) := x"FFF3";
          m(783) := x"002B";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_19.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 19) then
          m(0) := x"FFED";
          m(1) := x"0028";
          m(2) := x"FFF7";
          m(3) := x"FFE9";
          m(4) := x"FFFC";
          m(5) := x"FFF5";
          m(6) := x"002B";
          m(7) := x"0004";
          m(8) := x"FFCC";
          m(9) := x"FFF0";
          m(10) := x"FFFF";
          m(11) := x"0012";
          m(12) := x"FFE5";
          m(13) := x"0011";
          m(14) := x"FFE0";
          m(15) := x"FFF1";
          m(16) := x"0015";
          m(17) := x"FFFC";
          m(18) := x"0000";
          m(19) := x"0000";
          m(20) := x"0003";
          m(21) := x"FFF2";
          m(22) := x"FFE2";
          m(23) := x"0014";
          m(24) := x"0004";
          m(25) := x"0037";
          m(26) := x"000A";
          m(27) := x"0011";
          m(28) := x"FFEB";
          m(29) := x"FFCF";
          m(30) := x"FFDD";
          m(31) := x"0014";
          m(32) := x"FFCF";
          m(33) := x"0020";
          m(34) := x"001F";
          m(35) := x"FFEF";
          m(36) := x"002B";
          m(37) := x"FFF5";
          m(38) := x"001C";
          m(39) := x"FFFE";
          m(40) := x"FF5B";
          m(41) := x"FFC5";
          m(42) := x"0013";
          m(43) := x"FFC6";
          m(44) := x"FF39";
          m(45) := x"FF8F";
          m(46) := x"FFFC";
          m(47) := x"FFEF";
          m(48) := x"002D";
          m(49) := x"FFE2";
          m(50) := x"000E";
          m(51) := x"FFFB";
          m(52) := x"0008";
          m(53) := x"FFF6";
          m(54) := x"000C";
          m(55) := x"FFEB";
          m(56) := x"FFB4";
          m(57) := x"0000";
          m(58) := x"0000";
          m(59) := x"FFF9";
          m(60) := x"FFE2";
          m(61) := x"0004";
          m(62) := x"000F";
          m(63) := x"005A";
          m(64) := x"008D";
          m(65) := x"011C";
          m(66) := x"0173";
          m(67) := x"014B";
          m(68) := x"0145";
          m(69) := x"0184";
          m(70) := x"015E";
          m(71) := x"0139";
          m(72) := x"0164";
          m(73) := x"0104";
          m(74) := x"001C";
          m(75) := x"FFE4";
          m(76) := x"0020";
          m(77) := x"FFD7";
          m(78) := x"FFD3";
          m(79) := x"0018";
          m(80) := x"FFD7";
          m(81) := x"FFD1";
          m(82) := x"FFD4";
          m(83) := x"FFDD";
          m(84) := x"0023";
          m(85) := x"0022";
          m(86) := x"FFD4";
          m(87) := x"FFD2";
          m(88) := x"0004";
          m(89) := x"FF75";
          m(90) := x"0030";
          m(91) := x"0086";
          m(92) := x"009A";
          m(93) := x"01E4";
          m(94) := x"0100";
          m(95) := x"FFC7";
          m(96) := x"FF64";
          m(97) := x"0058";
          m(98) := x"FFC4";
          m(99) := x"FF85";
          m(100) := x"FF04";
          m(101) := x"FD62";
          m(102) := x"FFBC";
          m(103) := x"0180";
          m(104) := x"FFF5";
          m(105) := x"FF38";
          m(106) := x"FF83";
          m(107) := x"0036";
          m(108) := x"0042";
          m(109) := x"002F";
          m(110) := x"FFE4";
          m(111) := x"0029";
          m(112) := x"FFF6";
          m(113) := x"FFFC";
          m(114) := x"FFF3";
          m(115) := x"FF9C";
          m(116) := x"FFBF";
          m(117) := x"FF62";
          m(118) := x"FF43";
          m(119) := x"FF41";
          m(120) := x"FEF5";
          m(121) := x"000F";
          m(122) := x"01A8";
          m(123) := x"FC9C";
          m(124) := x"FF2E";
          m(125) := x"01BC";
          m(126) := x"03C5";
          m(127) := x"020B";
          m(128) := x"FF1F";
          m(129) := x"0065";
          m(130) := x"01D6";
          m(131) := x"FEBF";
          m(132) := x"FEF1";
          m(133) := x"00A4";
          m(134) := x"FF82";
          m(135) := x"FE01";
          m(136) := x"FE34";
          m(137) := x"FF4E";
          m(138) := x"FFC9";
          m(139) := x"0018";
          m(140) := x"003E";
          m(141) := x"FFC6";
          m(142) := x"001A";
          m(143) := x"FF41";
          m(144) := x"FFFE";
          m(145) := x"FF52";
          m(146) := x"FDFF";
          m(147) := x"FCFD";
          m(148) := x"FEC0";
          m(149) := x"FD0C";
          m(150) := x"FEB0";
          m(151) := x"0082";
          m(152) := x"0531";
          m(153) := x"01D6";
          m(154) := x"03A9";
          m(155) := x"02C3";
          m(156) := x"044F";
          m(157) := x"0432";
          m(158) := x"044E";
          m(159) := x"FF96";
          m(160) := x"FEB7";
          m(161) := x"FDA2";
          m(162) := x"FE27";
          m(163) := x"FD99";
          m(164) := x"FE18";
          m(165) := x"FED3";
          m(166) := x"0003";
          m(167) := x"0022";
          m(168) := x"001F";
          m(169) := x"FFEE";
          m(170) := x"0015";
          m(171) := x"FEFB";
          m(172) := x"FF76";
          m(173) := x"FCB0";
          m(174) := x"FC85";
          m(175) := x"FD9D";
          m(176) := x"FA90";
          m(177) := x"F9A0";
          m(178) := x"FEB5";
          m(179) := x"0217";
          m(180) := x"0032";
          m(181) := x"FCDC";
          m(182) := x"04CD";
          m(183) := x"055D";
          m(184) := x"055B";
          m(185) := x"FB69";
          m(186) := x"F9B0";
          m(187) := x"F567";
          m(188) := x"F52F";
          m(189) := x"FD9A";
          m(190) := x"FDAF";
          m(191) := x"FC26";
          m(192) := x"FD93";
          m(193) := x"FEDD";
          m(194) := x"000F";
          m(195) := x"FFF2";
          m(196) := x"FFFB";
          m(197) := x"FFF5";
          m(198) := x"0027";
          m(199) := x"FEBA";
          m(200) := x"FF1B";
          m(201) := x"FD5B";
          m(202) := x"FE72";
          m(203) := x"FEF1";
          m(204) := x"FAD8";
          m(205) := x"F6AE";
          m(206) := x"FC38";
          m(207) := x"039A";
          m(208) := x"FDF1";
          m(209) := x"FEC1";
          m(210) := x"0866";
          m(211) := x"FF48";
          m(212) := x"0073";
          m(213) := x"FDC2";
          m(214) := x"F9E5";
          m(215) := x"F447";
          m(216) := x"FB8A";
          m(217) := x"F956";
          m(218) := x"FE22";
          m(219) := x"FDA6";
          m(220) := x"0187";
          m(221) := x"FF99";
          m(222) := x"FFE1";
          m(223) := x"002A";
          m(224) := x"FFBD";
          m(225) := x"0025";
          m(226) := x"0026";
          m(227) := x"FE48";
          m(228) := x"FC2A";
          m(229) := x"FD59";
          m(230) := x"FE98";
          m(231) := x"FF7C";
          m(232) := x"FC24";
          m(233) := x"F8B0";
          m(234) := x"0001";
          m(235) := x"FB86";
          m(236) := x"F80A";
          m(237) := x"063C";
          m(238) := x"0784";
          m(239) := x"0830";
          m(240) := x"F9C5";
          m(241) := x"FAE5";
          m(242) := x"F92F";
          m(243) := x"FE94";
          m(244) := x"0420";
          m(245) := x"F9D3";
          m(246) := x"FE12";
          m(247) := x"032C";
          m(248) := x"0136";
          m(249) := x"FFC1";
          m(250) := x"FFFC";
          m(251) := x"FFBF";
          m(252) := x"0020";
          m(253) := x"FFF3";
          m(254) := x"0007";
          m(255) := x"FE6F";
          m(256) := x"FC75";
          m(257) := x"FE9A";
          m(258) := x"FB23";
          m(259) := x"FEEF";
          m(260) := x"FB8B";
          m(261) := x"FAA4";
          m(262) := x"FBE6";
          m(263) := x"F9B2";
          m(264) := x"FDDD";
          m(265) := x"033D";
          m(266) := x"06CD";
          m(267) := x"FE6F";
          m(268) := x"F73B";
          m(269) := x"FD3B";
          m(270) := x"FAAD";
          m(271) := x"FDD7";
          m(272) := x"026F";
          m(273) := x"FC80";
          m(274) := x"FF3A";
          m(275) := x"0077";
          m(276) := x"FE53";
          m(277) := x"FDBC";
          m(278) := x"FF3D";
          m(279) := x"0006";
          m(280) := x"FFF0";
          m(281) := x"0011";
          m(282) := x"FF6B";
          m(283) := x"FEAA";
          m(284) := x"FF53";
          m(285) := x"FFFC";
          m(286) := x"FE22";
          m(287) := x"FDF7";
          m(288) := x"FDD4";
          m(289) := x"FC56";
          m(290) := x"FCED";
          m(291) := x"FEED";
          m(292) := x"0109";
          m(293) := x"0712";
          m(294) := x"0067";
          m(295) := x"FE9A";
          m(296) := x"F96A";
          m(297) := x"FCE7";
          m(298) := x"FB95";
          m(299) := x"FE08";
          m(300) := x"01E7";
          m(301) := x"FF78";
          m(302) := x"01E1";
          m(303) := x"FD53";
          m(304) := x"FCE6";
          m(305) := x"FDA8";
          m(306) := x"FFDD";
          m(307) := x"FFF8";
          m(308) := x"FFC7";
          m(309) := x"FFCB";
          m(310) := x"FF58";
          m(311) := x"FF28";
          m(312) := x"FF3C";
          m(313) := x"01FF";
          m(314) := x"FE6F";
          m(315) := x"FFE1";
          m(316) := x"025B";
          m(317) := x"FF4F";
          m(318) := x"FE18";
          m(319) := x"FD02";
          m(320) := x"006E";
          m(321) := x"FB3D";
          m(322) := x"F988";
          m(323) := x"F91F";
          m(324) := x"FB7E";
          m(325) := x"F928";
          m(326) := x"FC51";
          m(327) := x"02F5";
          m(328) := x"FDBF";
          m(329) := x"00EF";
          m(330) := x"0044";
          m(331) := x"FC6A";
          m(332) := x"F939";
          m(333) := x"FF5A";
          m(334) := x"FEEC";
          m(335) := x"FFDC";
          m(336) := x"002F";
          m(337) := x"FFC4";
          m(338) := x"FF74";
          m(339) := x"FF50";
          m(340) := x"FD03";
          m(341) := x"FE72";
          m(342) := x"FB4C";
          m(343) := x"FE42";
          m(344) := x"0597";
          m(345) := x"029F";
          m(346) := x"00C7";
          m(347) := x"0281";
          m(348) := x"02C4";
          m(349) := x"FD7F";
          m(350) := x"FE22";
          m(351) := x"FC5D";
          m(352) := x"FF0A";
          m(353) := x"F89B";
          m(354) := x"FE01";
          m(355) := x"FE73";
          m(356) := x"FA2E";
          m(357) := x"FF92";
          m(358) := x"0099";
          m(359) := x"FA1F";
          m(360) := x"FCE4";
          m(361) := x"019A";
          m(362) := x"FF4E";
          m(363) := x"0006";
          m(364) := x"FFD4";
          m(365) := x"FFC7";
          m(366) := x"FFBC";
          m(367) := x"FF37";
          m(368) := x"FBFD";
          m(369) := x"FBFF";
          m(370) := x"FF76";
          m(371) := x"FDFA";
          m(372) := x"01B6";
          m(373) := x"0080";
          m(374) := x"023A";
          m(375) := x"0132";
          m(376) := x"04C6";
          m(377) := x"FFE6";
          m(378) := x"0252";
          m(379) := x"FDC6";
          m(380) := x"FBE5";
          m(381) := x"FE45";
          m(382) := x"FE42";
          m(383) := x"FC56";
          m(384) := x"FC8A";
          m(385) := x"FDE6";
          m(386) := x"F9E0";
          m(387) := x"FE6F";
          m(388) := x"0227";
          m(389) := x"0130";
          m(390) := x"0116";
          m(391) := x"0114";
          m(392) := x"001A";
          m(393) := x"FF9B";
          m(394) := x"FF72";
          m(395) := x"FFA3";
          m(396) := x"FEC5";
          m(397) := x"FCE4";
          m(398) := x"020C";
          m(399) := x"0229";
          m(400) := x"0075";
          m(401) := x"00A7";
          m(402) := x"FC98";
          m(403) := x"FDE9";
          m(404) := x"0463";
          m(405) := x"FF76";
          m(406) := x"01A9";
          m(407) := x"0118";
          m(408) := x"FE58";
          m(409) := x"F838";
          m(410) := x"FEED";
          m(411) := x"F9E5";
          m(412) := x"FEA9";
          m(413) := x"FE50";
          m(414) := x"FEC0";
          m(415) := x"FEB0";
          m(416) := x"FF1C";
          m(417) := x"0227";
          m(418) := x"015A";
          m(419) := x"FFFA";
          m(420) := x"0018";
          m(421) := x"FF3C";
          m(422) := x"FFB4";
          m(423) := x"015C";
          m(424) := x"FEC6";
          m(425) := x"FC0A";
          m(426) := x"02C0";
          m(427) := x"FF5D";
          m(428) := x"FFA3";
          m(429) := x"0789";
          m(430) := x"0194";
          m(431) := x"FFEA";
          m(432) := x"047D";
          m(433) := x"03AB";
          m(434) := x"055A";
          m(435) := x"0134";
          m(436) := x"02C7";
          m(437) := x"0540";
          m(438) := x"FCB4";
          m(439) := x"FE8C";
          m(440) := x"FD59";
          m(441) := x"FFCF";
          m(442) := x"FE45";
          m(443) := x"FCC3";
          m(444) := x"FE5F";
          m(445) := x"0388";
          m(446) := x"00CC";
          m(447) := x"002A";
          m(448) := x"0003";
          m(449) := x"FFA1";
          m(450) := x"FEF3";
          m(451) := x"00B4";
          m(452) := x"FF71";
          m(453) := x"FFF7";
          m(454) := x"0418";
          m(455) := x"05D1";
          m(456) := x"02A2";
          m(457) := x"093D";
          m(458) := x"033C";
          m(459) := x"FF58";
          m(460) := x"FD84";
          m(461) := x"FD11";
          m(462) := x"0149";
          m(463) := x"028B";
          m(464) := x"07E2";
          m(465) := x"0ADB";
          m(466) := x"FF48";
          m(467) := x"023A";
          m(468) := x"0074";
          m(469) := x"04E4";
          m(470) := x"FF69";
          m(471) := x"0356";
          m(472) := x"0383";
          m(473) := x"05E1";
          m(474) := x"0264";
          m(475) := x"FFE7";
          m(476) := x"002A";
          m(477) := x"FFB7";
          m(478) := x"FED1";
          m(479) := x"FEFD";
          m(480) := x"02AF";
          m(481) := x"02A2";
          m(482) := x"00D1";
          m(483) := x"FE63";
          m(484) := x"059D";
          m(485) := x"011D";
          m(486) := x"FE01";
          m(487) := x"FB17";
          m(488) := x"FD8F";
          m(489) := x"0283";
          m(490) := x"06A6";
          m(491) := x"0329";
          m(492) := x"03D1";
          m(493) := x"FF8D";
          m(494) := x"0505";
          m(495) := x"00B5";
          m(496) := x"021D";
          m(497) := x"00E8";
          m(498) := x"00BD";
          m(499) := x"01BB";
          m(500) := x"003C";
          m(501) := x"0432";
          m(502) := x"00F1";
          m(503) := x"FFB7";
          m(504) := x"FFE8";
          m(505) := x"FFCA";
          m(506) := x"FF43";
          m(507) := x"FFA8";
          m(508) := x"02FD";
          m(509) := x"0631";
          m(510) := x"0156";
          m(511) := x"0053";
          m(512) := x"036B";
          m(513) := x"FFF6";
          m(514) := x"FC9A";
          m(515) := x"FE74";
          m(516) := x"0578";
          m(517) := x"083F";
          m(518) := x"08EE";
          m(519) := x"02F6";
          m(520) := x"FFF2";
          m(521) := x"FDD7";
          m(522) := x"0672";
          m(523) := x"082D";
          m(524) := x"0418";
          m(525) := x"0343";
          m(526) := x"030F";
          m(527) := x"04D5";
          m(528) := x"0511";
          m(529) := x"03C7";
          m(530) := x"0048";
          m(531) := x"00B0";
          m(532) := x"001A";
          m(533) := x"0002";
          m(534) := x"FFAA";
          m(535) := x"0011";
          m(536) := x"01C0";
          m(537) := x"036E";
          m(538) := x"02EF";
          m(539) := x"01F6";
          m(540) := x"FE20";
          m(541) := x"FF9E";
          m(542) := x"FA57";
          m(543) := x"02F3";
          m(544) := x"00BC";
          m(545) := x"0575";
          m(546) := x"0382";
          m(547) := x"0AFA";
          m(548) := x"028F";
          m(549) := x"FE92";
          m(550) := x"02FC";
          m(551) := x"0742";
          m(552) := x"0535";
          m(553) := x"033A";
          m(554) := x"0593";
          m(555) := x"05B3";
          m(556) := x"040C";
          m(557) := x"02EB";
          m(558) := x"009B";
          m(559) := x"0061";
          m(560) := x"0024";
          m(561) := x"FFF0";
          m(562) := x"FFDF";
          m(563) := x"00C2";
          m(564) := x"01A5";
          m(565) := x"01F2";
          m(566) := x"034F";
          m(567) := x"0270";
          m(568) := x"0079";
          m(569) := x"FCAE";
          m(570) := x"FAE1";
          m(571) := x"020A";
          m(572) := x"FD29";
          m(573) := x"FA06";
          m(574) := x"0584";
          m(575) := x"0131";
          m(576) := x"0738";
          m(577) := x"02C1";
          m(578) := x"067F";
          m(579) := x"0323";
          m(580) := x"08F3";
          m(581) := x"0845";
          m(582) := x"04EE";
          m(583) := x"03C1";
          m(584) := x"028F";
          m(585) := x"0115";
          m(586) := x"00AB";
          m(587) := x"FFC3";
          m(588) := x"001E";
          m(589) := x"FFFC";
          m(590) := x"007B";
          m(591) := x"00EC";
          m(592) := x"02E7";
          m(593) := x"035F";
          m(594) := x"FEC5";
          m(595) := x"FE4B";
          m(596) := x"02C3";
          m(597) := x"FC5B";
          m(598) := x"FE7E";
          m(599) := x"FC39";
          m(600) := x"FD12";
          m(601) := x"FCD2";
          m(602) := x"FE30";
          m(603) := x"FBBC";
          m(604) := x"06D1";
          m(605) := x"049C";
          m(606) := x"09C1";
          m(607) := x"0622";
          m(608) := x"036A";
          m(609) := x"0507";
          m(610) := x"02CF";
          m(611) := x"0493";
          m(612) := x"00CA";
          m(613) := x"007E";
          m(614) := x"FFE1";
          m(615) := x"FFC4";
          m(616) := x"000C";
          m(617) := x"FFFE";
          m(618) := x"0095";
          m(619) := x"00BF";
          m(620) := x"036E";
          m(621) := x"0389";
          m(622) := x"FE08";
          m(623) := x"0045";
          m(624) := x"00AA";
          m(625) := x"0051";
          m(626) := x"FDA1";
          m(627) := x"FC0A";
          m(628) := x"FE02";
          m(629) := x"FDC2";
          m(630) := x"F972";
          m(631) := x"FBE9";
          m(632) := x"0140";
          m(633) := x"044B";
          m(634) := x"0323";
          m(635) := x"0473";
          m(636) := x"032C";
          m(637) := x"037B";
          m(638) := x"FCB1";
          m(639) := x"FEF1";
          m(640) := x"FF39";
          m(641) := x"FFDC";
          m(642) := x"0000";
          m(643) := x"0000";
          m(644) := x"0007";
          m(645) := x"0034";
          m(646) := x"0022";
          m(647) := x"FFF7";
          m(648) := x"00A4";
          m(649) := x"010B";
          m(650) := x"FEFD";
          m(651) := x"FE6E";
          m(652) := x"FC92";
          m(653) := x"FF4B";
          m(654) := x"FEA2";
          m(655) := x"FF96";
          m(656) := x"FD3B";
          m(657) := x"FA14";
          m(658) := x"F9B5";
          m(659) := x"F8BC";
          m(660) := x"F849";
          m(661) := x"F6AA";
          m(662) := x"FAC0";
          m(663) := x"FBCB";
          m(664) := x"FFD2";
          m(665) := x"FEB3";
          m(666) := x"FC3E";
          m(667) := x"FEF5";
          m(668) := x"FEA7";
          m(669) := x"0079";
          m(670) := x"004D";
          m(671) := x"000F";
          m(672) := x"FFFC";
          m(673) := x"0030";
          m(674) := x"002F";
          m(675) := x"0023";
          m(676) := x"FFFB";
          m(677) := x"00C9";
          m(678) := x"FFA6";
          m(679) := x"FE1F";
          m(680) := x"FFC5";
          m(681) := x"02DC";
          m(682) := x"0093";
          m(683) := x"0257";
          m(684) := x"FA78";
          m(685) := x"F562";
          m(686) := x"F9E7";
          m(687) := x"FC7C";
          m(688) := x"F7B0";
          m(689) := x"F597";
          m(690) := x"F74D";
          m(691) := x"FB8B";
          m(692) := x"F9AE";
          m(693) := x"FD1E";
          m(694) := x"FC78";
          m(695) := x"FCE6";
          m(696) := x"00E3";
          m(697) := x"00D2";
          m(698) := x"001C";
          m(699) := x"0010";
          m(700) := x"FFED";
          m(701) := x"FFE2";
          m(702) := x"FFC9";
          m(703) := x"0005";
          m(704) := x"FFA9";
          m(705) := x"FF32";
          m(706) := x"FF3F";
          m(707) := x"FECE";
          m(708) := x"FF1B";
          m(709) := x"FED5";
          m(710) := x"FF21";
          m(711) := x"FE1F";
          m(712) := x"F977";
          m(713) := x"F7D8";
          m(714) := x"F910";
          m(715) := x"FD15";
          m(716) := x"F4AC";
          m(717) := x"F77D";
          m(718) := x"F68A";
          m(719) := x"F610";
          m(720) := x"F9EF";
          m(721) := x"FD41";
          m(722) := x"FF95";
          m(723) := x"FF22";
          m(724) := x"FFC1";
          m(725) := x"0056";
          m(726) := x"0050";
          m(727) := x"0009";
          m(728) := x"FFC8";
          m(729) := x"0022";
          m(730) := x"FFD8";
          m(731) := x"001A";
          m(732) := x"FFB7";
          m(733) := x"FF69";
          m(734) := x"FF49";
          m(735) := x"FEBB";
          m(736) := x"FEE2";
          m(737) := x"FD41";
          m(738) := x"FE22";
          m(739) := x"FE61";
          m(740) := x"FD9B";
          m(741) := x"FD8D";
          m(742) := x"FCF0";
          m(743) := x"FEFA";
          m(744) := x"FE23";
          m(745) := x"FDEE";
          m(746) := x"FD67";
          m(747) := x"FDFA";
          m(748) := x"FDFB";
          m(749) := x"FF43";
          m(750) := x"FFA3";
          m(751) := x"0024";
          m(752) := x"FFD9";
          m(753) := x"FFF1";
          m(754) := x"FFF6";
          m(755) := x"001D";
          m(756) := x"FFE0";
          m(757) := x"0010";
          m(758) := x"0031";
          m(759) := x"0024";
          m(760) := x"000D";
          m(761) := x"FFFD";
          m(762) := x"FFFF";
          m(763) := x"FFC5";
          m(764) := x"FFD0";
          m(765) := x"0000";
          m(766) := x"FF96";
          m(767) := x"0008";
          m(768) := x"FF92";
          m(769) := x"FFC9";
          m(770) := x"FF90";
          m(771) := x"FFCF";
          m(772) := x"FFF2";
          m(773) := x"FFCC";
          m(774) := x"FF54";
          m(775) := x"000D";
          m(776) := x"0004";
          m(777) := x"FFE6";
          m(778) := x"FFE3";
          m(779) := x"0021";
          m(780) := x"0007";
          m(781) := x"001F";
          m(782) := x"000D";
          m(783) := x"FFFA";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_20.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 20) then
          m(0) := x"FFD2";
          m(1) := x"FFFC";
          m(2) := x"0000";
          m(3) := x"FFC2";
          m(4) := x"FFEF";
          m(5) := x"001C";
          m(6) := x"0001";
          m(7) := x"0041";
          m(8) := x"FFFA";
          m(9) := x"003F";
          m(10) := x"0013";
          m(11) := x"0012";
          m(12) := x"FFEC";
          m(13) := x"000B";
          m(14) := x"FFE2";
          m(15) := x"0005";
          m(16) := x"0021";
          m(17) := x"FFD3";
          m(18) := x"FFF5";
          m(19) := x"FFF0";
          m(20) := x"0007";
          m(21) := x"0006";
          m(22) := x"FFE9";
          m(23) := x"0005";
          m(24) := x"FFFA";
          m(25) := x"003B";
          m(26) := x"FFFC";
          m(27) := x"FFD7";
          m(28) := x"FFEB";
          m(29) := x"001B";
          m(30) := x"FFC9";
          m(31) := x"0035";
          m(32) := x"0000";
          m(33) := x"FFDE";
          m(34) := x"FFBF";
          m(35) := x"FFA0";
          m(36) := x"FF7D";
          m(37) := x"FFBB";
          m(38) := x"FFF4";
          m(39) := x"FF8E";
          m(40) := x"FF66";
          m(41) := x"FF9A";
          m(42) := x"FFF3";
          m(43) := x"FF6C";
          m(44) := x"FE52";
          m(45) := x"FEF5";
          m(46) := x"FFDB";
          m(47) := x"FF4F";
          m(48) := x"FF61";
          m(49) := x"0003";
          m(50) := x"FFD4";
          m(51) := x"FFAE";
          m(52) := x"FFFB";
          m(53) := x"FFC7";
          m(54) := x"FFDA";
          m(55) := x"FFE8";
          m(56) := x"FFF4";
          m(57) := x"FFF3";
          m(58) := x"FFE9";
          m(59) := x"FFE7";
          m(60) := x"0001";
          m(61) := x"0011";
          m(62) := x"FFF4";
          m(63) := x"FEDA";
          m(64) := x"FE33";
          m(65) := x"FE2D";
          m(66) := x"FE30";
          m(67) := x"FD8F";
          m(68) := x"FE33";
          m(69) := x"0063";
          m(70) := x"FE4F";
          m(71) := x"FF8E";
          m(72) := x"FE85";
          m(73) := x"FD5F";
          m(74) := x"FD8F";
          m(75) := x"FEFE";
          m(76) := x"FEDD";
          m(77) := x"FF5D";
          m(78) := x"0000";
          m(79) := x"FF6F";
          m(80) := x"FF56";
          m(81) := x"003F";
          m(82) := x"0013";
          m(83) := x"FFF7";
          m(84) := x"FFF2";
          m(85) := x"000F";
          m(86) := x"0030";
          m(87) := x"FFCC";
          m(88) := x"FFD5";
          m(89) := x"FFD4";
          m(90) := x"FCB6";
          m(91) := x"FCAA";
          m(92) := x"FB42";
          m(93) := x"FBBE";
          m(94) := x"FDB3";
          m(95) := x"FCEF";
          m(96) := x"F9B9";
          m(97) := x"F83B";
          m(98) := x"FAAC";
          m(99) := x"FEA3";
          m(100) := x"FE45";
          m(101) := x"0265";
          m(102) := x"04D9";
          m(103) := x"0080";
          m(104) := x"FD24";
          m(105) := x"FD2C";
          m(106) := x"0045";
          m(107) := x"011D";
          m(108) := x"004D";
          m(109) := x"FFE2";
          m(110) := x"FFA5";
          m(111) := x"FFF8";
          m(112) := x"FFC6";
          m(113) := x"FFFA";
          m(114) := x"FFFF";
          m(115) := x"FFC9";
          m(116) := x"FF97";
          m(117) := x"FF92";
          m(118) := x"FCE7";
          m(119) := x"FB5E";
          m(120) := x"FB8D";
          m(121) := x"FCC8";
          m(122) := x"FAE6";
          m(123) := x"0021";
          m(124) := x"0489";
          m(125) := x"02B0";
          m(126) := x"0024";
          m(127) := x"02A3";
          m(128) := x"FF5A";
          m(129) := x"FC77";
          m(130) := x"008B";
          m(131) := x"FDEB";
          m(132) := x"009D";
          m(133) := x"0358";
          m(134) := x"03E2";
          m(135) := x"0524";
          m(136) := x"0192";
          m(137) := x"0024";
          m(138) := x"FFAA";
          m(139) := x"FFE9";
          m(140) := x"000D";
          m(141) := x"0035";
          m(142) := x"0019";
          m(143) := x"FFE6";
          m(144) := x"00D4";
          m(145) := x"039D";
          m(146) := x"FFA8";
          m(147) := x"FD20";
          m(148) := x"00DC";
          m(149) := x"0246";
          m(150) := x"0007";
          m(151) := x"01FB";
          m(152) := x"0427";
          m(153) := x"FDD9";
          m(154) := x"02F9";
          m(155) := x"01BB";
          m(156) := x"FF7E";
          m(157) := x"01B4";
          m(158) := x"0413";
          m(159) := x"FF6B";
          m(160) := x"0246";
          m(161) := x"052D";
          m(162) := x"087E";
          m(163) := x"04E4";
          m(164) := x"0293";
          m(165) := x"006E";
          m(166) := x"FFE4";
          m(167) := x"FFE2";
          m(168) := x"0018";
          m(169) := x"000B";
          m(170) := x"FF8F";
          m(171) := x"FF49";
          m(172) := x"FFCF";
          m(173) := x"01A3";
          m(174) := x"0054";
          m(175) := x"FEBC";
          m(176) := x"04E8";
          m(177) := x"03E7";
          m(178) := x"0585";
          m(179) := x"FD0F";
          m(180) := x"060D";
          m(181) := x"FE6C";
          m(182) := x"03B8";
          m(183) := x"050D";
          m(184) := x"FD90";
          m(185) := x"0598";
          m(186) := x"0542";
          m(187) := x"02BA";
          m(188) := x"04BC";
          m(189) := x"0515";
          m(190) := x"080F";
          m(191) := x"095C";
          m(192) := x"04F8";
          m(193) := x"0153";
          m(194) := x"003A";
          m(195) := x"FFFE";
          m(196) := x"FFEE";
          m(197) := x"FFDA";
          m(198) := x"FFE4";
          m(199) := x"FFE9";
          m(200) := x"FF49";
          m(201) := x"0509";
          m(202) := x"0284";
          m(203) := x"FF8D";
          m(204) := x"FFD3";
          m(205) := x"0014";
          m(206) := x"01F7";
          m(207) := x"003C";
          m(208) := x"0151";
          m(209) := x"02C7";
          m(210) := x"0265";
          m(211) := x"02B9";
          m(212) := x"01AA";
          m(213) := x"0327";
          m(214) := x"045A";
          m(215) := x"0424";
          m(216) := x"0458";
          m(217) := x"0304";
          m(218) := x"0524";
          m(219) := x"0A5E";
          m(220) := x"035F";
          m(221) := x"01AB";
          m(222) := x"014A";
          m(223) := x"FFC1";
          m(224) := x"FFE6";
          m(225) := x"FFEB";
          m(226) := x"0029";
          m(227) := x"010A";
          m(228) := x"0241";
          m(229) := x"03C6";
          m(230) := x"02B6";
          m(231) := x"00AA";
          m(232) := x"FFD0";
          m(233) := x"01C0";
          m(234) := x"FC23";
          m(235) := x"01AA";
          m(236) := x"043C";
          m(237) := x"0113";
          m(238) := x"0068";
          m(239) := x"FD87";
          m(240) := x"0095";
          m(241) := x"02A9";
          m(242) := x"0840";
          m(243) := x"FEB0";
          m(244) := x"FDA9";
          m(245) := x"01FE";
          m(246) := x"0424";
          m(247) := x"04B8";
          m(248) := x"0464";
          m(249) := x"026A";
          m(250) := x"0102";
          m(251) := x"FFE8";
          m(252) := x"FFF8";
          m(253) := x"0006";
          m(254) := x"001F";
          m(255) := x"0091";
          m(256) := x"0042";
          m(257) := x"0033";
          m(258) := x"0570";
          m(259) := x"02AD";
          m(260) := x"03BC";
          m(261) := x"0382";
          m(262) := x"024C";
          m(263) := x"0602";
          m(264) := x"FF3E";
          m(265) := x"0350";
          m(266) := x"F9CB";
          m(267) := x"FE32";
          m(268) := x"02C0";
          m(269) := x"00DB";
          m(270) := x"0342";
          m(271) := x"FEFF";
          m(272) := x"FBC8";
          m(273) := x"0231";
          m(274) := x"FF15";
          m(275) := x"045F";
          m(276) := x"017E";
          m(277) := x"0471";
          m(278) := x"0338";
          m(279) := x"02F3";
          m(280) := x"FFDD";
          m(281) := x"0012";
          m(282) := x"FFCA";
          m(283) := x"FF80";
          m(284) := x"FDD4";
          m(285) := x"FE29";
          m(286) := x"0348";
          m(287) := x"FE67";
          m(288) := x"FED5";
          m(289) := x"FFA9";
          m(290) := x"FD63";
          m(291) := x"FE59";
          m(292) := x"026E";
          m(293) := x"0152";
          m(294) := x"FB55";
          m(295) := x"00DE";
          m(296) := x"04DF";
          m(297) := x"FF36";
          m(298) := x"0396";
          m(299) := x"0827";
          m(300) := x"0123";
          m(301) := x"FC6F";
          m(302) := x"00C2";
          m(303) := x"0108";
          m(304) := x"02A8";
          m(305) := x"087B";
          m(306) := x"0141";
          m(307) := x"00B6";
          m(308) := x"0029";
          m(309) := x"FFF5";
          m(310) := x"0044";
          m(311) := x"FFED";
          m(312) := x"0094";
          m(313) := x"0180";
          m(314) := x"00B6";
          m(315) := x"FBD6";
          m(316) := x"FBB6";
          m(317) := x"FFA2";
          m(318) := x"01F1";
          m(319) := x"FEBA";
          m(320) := x"02F3";
          m(321) := x"0325";
          m(322) := x"048D";
          m(323) := x"05BD";
          m(324) := x"004E";
          m(325) := x"FE2F";
          m(326) := x"01E6";
          m(327) := x"0237";
          m(328) := x"FC50";
          m(329) := x"00A3";
          m(330) := x"FFEB";
          m(331) := x"FC79";
          m(332) := x"FD0E";
          m(333) := x"FDF7";
          m(334) := x"FFCF";
          m(335) := x"0073";
          m(336) := x"FFF8";
          m(337) := x"0008";
          m(338) := x"00A5";
          m(339) := x"00B1";
          m(340) := x"0306";
          m(341) := x"00A8";
          m(342) := x"0126";
          m(343) := x"FF54";
          m(344) := x"02A4";
          m(345) := x"0510";
          m(346) := x"0275";
          m(347) := x"FF13";
          m(348) := x"02FB";
          m(349) := x"02DE";
          m(350) := x"FFB6";
          m(351) := x"028A";
          m(352) := x"FD28";
          m(353) := x"FB1C";
          m(354) := x"FFDA";
          m(355) := x"FE34";
          m(356) := x"FC57";
          m(357) := x"FCED";
          m(358) := x"FC4F";
          m(359) := x"FB85";
          m(360) := x"FB84";
          m(361) := x"FE8C";
          m(362) := x"01DC";
          m(363) := x"00CA";
          m(364) := x"0012";
          m(365) := x"FFE2";
          m(366) := x"0052";
          m(367) := x"00B7";
          m(368) := x"04C8";
          m(369) := x"01BB";
          m(370) := x"0286";
          m(371) := x"03D3";
          m(372) := x"044E";
          m(373) := x"073F";
          m(374) := x"FCF6";
          m(375) := x"009B";
          m(376) := x"0188";
          m(377) := x"FAAC";
          m(378) := x"FF2E";
          m(379) := x"FC9C";
          m(380) := x"F9DE";
          m(381) := x"0445";
          m(382) := x"FDDC";
          m(383) := x"FB3B";
          m(384) := x"FE10";
          m(385) := x"FB88";
          m(386) := x"FC36";
          m(387) := x"FB0D";
          m(388) := x"FDF6";
          m(389) := x"042E";
          m(390) := x"FF48";
          m(391) := x"FF09";
          m(392) := x"FFD4";
          m(393) := x"FFF1";
          m(394) := x"0016";
          m(395) := x"0111";
          m(396) := x"020E";
          m(397) := x"FF39";
          m(398) := x"FC37";
          m(399) := x"0016";
          m(400) := x"FFFA";
          m(401) := x"FD4E";
          m(402) := x"FD00";
          m(403) := x"002D";
          m(404) := x"018D";
          m(405) := x"FA26";
          m(406) := x"FE2D";
          m(407) := x"FD60";
          m(408) := x"F819";
          m(409) := x"068F";
          m(410) := x"F731";
          m(411) := x"01B7";
          m(412) := x"FCAD";
          m(413) := x"FD4B";
          m(414) := x"F989";
          m(415) := x"FA92";
          m(416) := x"FCE0";
          m(417) := x"0126";
          m(418) := x"FE92";
          m(419) := x"FFEF";
          m(420) := x"FFDA";
          m(421) := x"FFEB";
          m(422) := x"FFED";
          m(423) := x"FFFA";
          m(424) := x"FCD2";
          m(425) := x"FF6C";
          m(426) := x"02BA";
          m(427) := x"05A2";
          m(428) := x"0282";
          m(429) := x"00B9";
          m(430) := x"FE39";
          m(431) := x"04B7";
          m(432) := x"FEB8";
          m(433) := x"F6C7";
          m(434) := x"002A";
          m(435) := x"0487";
          m(436) := x"FD1F";
          m(437) := x"025E";
          m(438) := x"FC5C";
          m(439) := x"FC81";
          m(440) := x"FA1F";
          m(441) := x"0073";
          m(442) := x"FF8E";
          m(443) := x"FF90";
          m(444) := x"FF52";
          m(445) := x"FC8C";
          m(446) := x"00BD";
          m(447) := x"FF62";
          m(448) := x"FFF9";
          m(449) := x"FFF3";
          m(450) := x"FFBA";
          m(451) := x"FD89";
          m(452) := x"FE3D";
          m(453) := x"FF18";
          m(454) := x"FDFD";
          m(455) := x"0102";
          m(456) := x"067D";
          m(457) := x"FF8E";
          m(458) := x"FC13";
          m(459) := x"FE87";
          m(460) := x"0488";
          m(461) := x"00D2";
          m(462) := x"FA69";
          m(463) := x"FE58";
          m(464) := x"F97C";
          m(465) := x"F8B9";
          m(466) := x"0077";
          m(467) := x"FCE7";
          m(468) := x"02B3";
          m(469) := x"FDAA";
          m(470) := x"00EC";
          m(471) := x"00E7";
          m(472) := x"FC77";
          m(473) := x"F9F0";
          m(474) := x"FFB2";
          m(475) := x"0004";
          m(476) := x"FFD3";
          m(477) := x"001B";
          m(478) := x"FFD9";
          m(479) := x"FD48";
          m(480) := x"FD1D";
          m(481) := x"0217";
          m(482) := x"003F";
          m(483) := x"01B7";
          m(484) := x"018E";
          m(485) := x"FF4F";
          m(486) := x"FBD5";
          m(487) := x"FF75";
          m(488) := x"0082";
          m(489) := x"FF3A";
          m(490) := x"FF00";
          m(491) := x"FB71";
          m(492) := x"FD95";
          m(493) := x"FEDE";
          m(494) := x"FE2A";
          m(495) := x"FEEE";
          m(496) := x"FEC0";
          m(497) := x"FD38";
          m(498) := x"05F9";
          m(499) := x"06CA";
          m(500) := x"0450";
          m(501) := x"FBF7";
          m(502) := x"00D1";
          m(503) := x"FFCE";
          m(504) := x"0005";
          m(505) := x"FFD4";
          m(506) := x"0066";
          m(507) := x"FCC5";
          m(508) := x"FE68";
          m(509) := x"FECA";
          m(510) := x"00B7";
          m(511) := x"FF11";
          m(512) := x"0258";
          m(513) := x"FE36";
          m(514) := x"FD74";
          m(515) := x"FEEC";
          m(516) := x"FD74";
          m(517) := x"0416";
          m(518) := x"F95B";
          m(519) := x"FCC4";
          m(520) := x"FA53";
          m(521) := x"FB8B";
          m(522) := x"FD3E";
          m(523) := x"FD2D";
          m(524) := x"0541";
          m(525) := x"FCF1";
          m(526) := x"00AF";
          m(527) := x"0011";
          m(528) := x"FCCC";
          m(529) := x"FB2B";
          m(530) := x"0082";
          m(531) := x"FFC3";
          m(532) := x"0053";
          m(533) := x"001E";
          m(534) := x"0086";
          m(535) := x"FE79";
          m(536) := x"FB51";
          m(537) := x"FD77";
          m(538) := x"FFC7";
          m(539) := x"01EE";
          m(540) := x"011D";
          m(541) := x"0091";
          m(542) := x"FCA5";
          m(543) := x"F8BA";
          m(544) := x"FB82";
          m(545) := x"0406";
          m(546) := x"F970";
          m(547) := x"FA63";
          m(548) := x"FDE0";
          m(549) := x"FB20";
          m(550) := x"FF69";
          m(551) := x"FFA0";
          m(552) := x"0155";
          m(553) := x"FF43";
          m(554) := x"FC7E";
          m(555) := x"FDAB";
          m(556) := x"FE58";
          m(557) := x"FCCE";
          m(558) := x"FF28";
          m(559) := x"001F";
          m(560) := x"FFF7";
          m(561) := x"001C";
          m(562) := x"FF98";
          m(563) := x"FD7A";
          m(564) := x"FBE9";
          m(565) := x"FAE7";
          m(566) := x"FF08";
          m(567) := x"0059";
          m(568) := x"00AD";
          m(569) := x"014C";
          m(570) := x"FAF9";
          m(571) := x"F7D0";
          m(572) := x"FECD";
          m(573) := x"FD66";
          m(574) := x"FDA7";
          m(575) := x"FE4B";
          m(576) := x"064C";
          m(577) := x"0230";
          m(578) := x"FAF8";
          m(579) := x"03EF";
          m(580) := x"03D7";
          m(581) := x"007A";
          m(582) := x"FF58";
          m(583) := x"0385";
          m(584) := x"048A";
          m(585) := x"009A";
          m(586) := x"FFE7";
          m(587) := x"0009";
          m(588) := x"0048";
          m(589) := x"FFFE";
          m(590) := x"FE63";
          m(591) := x"FE32";
          m(592) := x"003F";
          m(593) := x"FD28";
          m(594) := x"FDFE";
          m(595) := x"020A";
          m(596) := x"02B1";
          m(597) := x"00DB";
          m(598) := x"FCA4";
          m(599) := x"FFDE";
          m(600) := x"FECE";
          m(601) := x"FCE7";
          m(602) := x"01C3";
          m(603) := x"0266";
          m(604) := x"048F";
          m(605) := x"03A0";
          m(606) := x"050E";
          m(607) := x"098E";
          m(608) := x"092D";
          m(609) := x"0553";
          m(610) := x"05F6";
          m(611) := x"0554";
          m(612) := x"0693";
          m(613) := x"0087";
          m(614) := x"FF8D";
          m(615) := x"FFFA";
          m(616) := x"FFE4";
          m(617) := x"0029";
          m(618) := x"FFD7";
          m(619) := x"00C2";
          m(620) := x"0432";
          m(621) := x"014C";
          m(622) := x"0529";
          m(623) := x"05FA";
          m(624) := x"0946";
          m(625) := x"0540";
          m(626) := x"0012";
          m(627) := x"09AF";
          m(628) := x"0553";
          m(629) := x"048A";
          m(630) := x"07DC";
          m(631) := x"052D";
          m(632) := x"0A93";
          m(633) := x"083B";
          m(634) := x"07DE";
          m(635) := x"091A";
          m(636) := x"05CB";
          m(637) := x"0840";
          m(638) := x"0760";
          m(639) := x"0788";
          m(640) := x"03AA";
          m(641) := x"0023";
          m(642) := x"FFAA";
          m(643) := x"0034";
          m(644) := x"FFF8";
          m(645) := x"FFF0";
          m(646) := x"FFAB";
          m(647) := x"0098";
          m(648) := x"0591";
          m(649) := x"0631";
          m(650) := x"07D4";
          m(651) := x"09D8";
          m(652) := x"0B01";
          m(653) := x"0A1C";
          m(654) := x"0820";
          m(655) := x"0C1A";
          m(656) := x"0973";
          m(657) := x"0BB5";
          m(658) := x"0E51";
          m(659) := x"0E7A";
          m(660) := x"0DDA";
          m(661) := x"0E69";
          m(662) := x"0BAB";
          m(663) := x"070C";
          m(664) := x"03BF";
          m(665) := x"02E4";
          m(666) := x"0308";
          m(667) := x"037B";
          m(668) := x"02D3";
          m(669) := x"FFF6";
          m(670) := x"FFDE";
          m(671) := x"0001";
          m(672) := x"FFDA";
          m(673) := x"0026";
          m(674) := x"0012";
          m(675) := x"FFFC";
          m(676) := x"0225";
          m(677) := x"0458";
          m(678) := x"0647";
          m(679) := x"0864";
          m(680) := x"091D";
          m(681) := x"0AA8";
          m(682) := x"0838";
          m(683) := x"08D1";
          m(684) := x"099B";
          m(685) := x"0DB3";
          m(686) := x"0AAE";
          m(687) := x"08C2";
          m(688) := x"0480";
          m(689) := x"0405";
          m(690) := x"04D3";
          m(691) := x"017F";
          m(692) := x"01F1";
          m(693) := x"0185";
          m(694) := x"027F";
          m(695) := x"02F2";
          m(696) := x"0051";
          m(697) := x"FF3A";
          m(698) := x"FFC1";
          m(699) := x"FFD2";
          m(700) := x"0027";
          m(701) := x"0006";
          m(702) := x"0003";
          m(703) := x"0058";
          m(704) := x"0140";
          m(705) := x"015B";
          m(706) := x"01D6";
          m(707) := x"0280";
          m(708) := x"040A";
          m(709) := x"05E2";
          m(710) := x"0326";
          m(711) := x"0299";
          m(712) := x"02F7";
          m(713) := x"0402";
          m(714) := x"0394";
          m(715) := x"0359";
          m(716) := x"0131";
          m(717) := x"0022";
          m(718) := x"FE79";
          m(719) := x"FE23";
          m(720) := x"00EE";
          m(721) := x"013B";
          m(722) := x"0092";
          m(723) := x"00E1";
          m(724) := x"007A";
          m(725) := x"FFD3";
          m(726) := x"FF92";
          m(727) := x"0019";
          m(728) := x"0014";
          m(729) := x"FFC7";
          m(730) := x"000A";
          m(731) := x"0011";
          m(732) := x"0025";
          m(733) := x"009D";
          m(734) := x"00D3";
          m(735) := x"00AB";
          m(736) := x"00C3";
          m(737) := x"028F";
          m(738) := x"00E0";
          m(739) := x"005D";
          m(740) := x"008F";
          m(741) := x"0091";
          m(742) := x"0082";
          m(743) := x"005F";
          m(744) := x"FF76";
          m(745) := x"FCF2";
          m(746) := x"FD9A";
          m(747) := x"FCE0";
          m(748) := x"FF5B";
          m(749) := x"0026";
          m(750) := x"0014";
          m(751) := x"0001";
          m(752) := x"FFF3";
          m(753) := x"002D";
          m(754) := x"FFE1";
          m(755) := x"FFF0";
          m(756) := x"0034";
          m(757) := x"000B";
          m(758) := x"0015";
          m(759) := x"0004";
          m(760) := x"002F";
          m(761) := x"FFDA";
          m(762) := x"0032";
          m(763) := x"0033";
          m(764) := x"FFD8";
          m(765) := x"FFD5";
          m(766) := x"002B";
          m(767) := x"0029";
          m(768) := x"FFFD";
          m(769) := x"FFFB";
          m(770) := x"FFFF";
          m(771) := x"0006";
          m(772) := x"0041";
          m(773) := x"0039";
          m(774) := x"00B0";
          m(775) := x"FFD1";
          m(776) := x"FFC3";
          m(777) := x"FFF4";
          m(778) := x"FFED";
          m(779) := x"FFDA";
          m(780) := x"FFFE";
          m(781) := x"0023";
          m(782) := x"FFF5";
          m(783) := x"FFD9";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_21.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 21) then
          m(0) := x"0010";
          m(1) := x"FFD6";
          m(2) := x"001D";
          m(3) := x"FFD1";
          m(4) := x"FFD6";
          m(5) := x"0027";
          m(6) := x"002C";
          m(7) := x"FFF3";
          m(8) := x"FFE7";
          m(9) := x"0002";
          m(10) := x"0004";
          m(11) := x"0001";
          m(12) := x"FFFF";
          m(13) := x"000C";
          m(14) := x"000D";
          m(15) := x"0011";
          m(16) := x"FFFD";
          m(17) := x"0003";
          m(18) := x"FFE1";
          m(19) := x"000E";
          m(20) := x"FFE0";
          m(21) := x"0023";
          m(22) := x"FFB2";
          m(23) := x"0024";
          m(24) := x"FFED";
          m(25) := x"FFD3";
          m(26) := x"FFBB";
          m(27) := x"001D";
          m(28) := x"FFCE";
          m(29) := x"FFDD";
          m(30) := x"0007";
          m(31) := x"004E";
          m(32) := x"0007";
          m(33) := x"0057";
          m(34) := x"FFE3";
          m(35) := x"0005";
          m(36) := x"004F";
          m(37) := x"002D";
          m(38) := x"0032";
          m(39) := x"0042";
          m(40) := x"006C";
          m(41) := x"009C";
          m(42) := x"0033";
          m(43) := x"FF74";
          m(44) := x"FF29";
          m(45) := x"0024";
          m(46) := x"FFFF";
          m(47) := x"0089";
          m(48) := x"0059";
          m(49) := x"0046";
          m(50) := x"FFEC";
          m(51) := x"FFD9";
          m(52) := x"0013";
          m(53) := x"FFF0";
          m(54) := x"FFE4";
          m(55) := x"001B";
          m(56) := x"0015";
          m(57) := x"FFFB";
          m(58) := x"002E";
          m(59) := x"0002";
          m(60) := x"0031";
          m(61) := x"0016";
          m(62) := x"007C";
          m(63) := x"011B";
          m(64) := x"00E9";
          m(65) := x"0069";
          m(66) := x"FFC1";
          m(67) := x"0023";
          m(68) := x"0092";
          m(69) := x"0006";
          m(70) := x"0015";
          m(71) := x"FFD8";
          m(72) := x"FD62";
          m(73) := x"00FC";
          m(74) := x"0098";
          m(75) := x"FF80";
          m(76) := x"FF51";
          m(77) := x"01C0";
          m(78) := x"007D";
          m(79) := x"0008";
          m(80) := x"FF07";
          m(81) := x"FF36";
          m(82) := x"0002";
          m(83) := x"0006";
          m(84) := x"0040";
          m(85) := x"FFDB";
          m(86) := x"FFF3";
          m(87) := x"FFD6";
          m(88) := x"0029";
          m(89) := x"0018";
          m(90) := x"00D8";
          m(91) := x"0063";
          m(92) := x"FFB2";
          m(93) := x"0095";
          m(94) := x"0098";
          m(95) := x"FFF3";
          m(96) := x"FE59";
          m(97) := x"FD0E";
          m(98) := x"FF4D";
          m(99) := x"01AB";
          m(100) := x"FD6F";
          m(101) := x"FFA2";
          m(102) := x"0322";
          m(103) := x"0161";
          m(104) := x"003A";
          m(105) := x"0020";
          m(106) := x"007E";
          m(107) := x"00BC";
          m(108) := x"FF7A";
          m(109) := x"FF60";
          m(110) := x"0015";
          m(111) := x"FFD5";
          m(112) := x"FFDE";
          m(113) := x"FFEB";
          m(114) := x"FFD8";
          m(115) := x"FFFB";
          m(116) := x"FFE1";
          m(117) := x"008A";
          m(118) := x"011C";
          m(119) := x"FF78";
          m(120) := x"FFBF";
          m(121) := x"018B";
          m(122) := x"FE1D";
          m(123) := x"FE89";
          m(124) := x"00B4";
          m(125) := x"039D";
          m(126) := x"04F4";
          m(127) := x"0294";
          m(128) := x"01C6";
          m(129) := x"021D";
          m(130) := x"FC45";
          m(131) := x"004B";
          m(132) := x"FD5F";
          m(133) := x"FF39";
          m(134) := x"FEC9";
          m(135) := x"005F";
          m(136) := x"FFD0";
          m(137) := x"FFE2";
          m(138) := x"0027";
          m(139) := x"0038";
          m(140) := x"FFF6";
          m(141) := x"FFEC";
          m(142) := x"FFCC";
          m(143) := x"0014";
          m(144) := x"FFCD";
          m(145) := x"0129";
          m(146) := x"0150";
          m(147) := x"0198";
          m(148) := x"0325";
          m(149) := x"0125";
          m(150) := x"01E1";
          m(151) := x"04A1";
          m(152) := x"0363";
          m(153) := x"0163";
          m(154) := x"0117";
          m(155) := x"032C";
          m(156) := x"009D";
          m(157) := x"0456";
          m(158) := x"0485";
          m(159) := x"0652";
          m(160) := x"FE90";
          m(161) := x"0042";
          m(162) := x"01C7";
          m(163) := x"0255";
          m(164) := x"02B6";
          m(165) := x"011A";
          m(166) := x"00AB";
          m(167) := x"002C";
          m(168) := x"FFCE";
          m(169) := x"0003";
          m(170) := x"001F";
          m(171) := x"0020";
          m(172) := x"FEFB";
          m(173) := x"FE74";
          m(174) := x"FAC8";
          m(175) := x"FAE6";
          m(176) := x"0173";
          m(177) := x"FB95";
          m(178) := x"F810";
          m(179) := x"FE19";
          m(180) := x"FFE9";
          m(181) := x"00F5";
          m(182) := x"FE0F";
          m(183) := x"FFC2";
          m(184) := x"FBAE";
          m(185) := x"01F4";
          m(186) := x"005F";
          m(187) := x"FFF2";
          m(188) := x"01C2";
          m(189) := x"0446";
          m(190) := x"02F6";
          m(191) := x"0541";
          m(192) := x"05F5";
          m(193) := x"02B8";
          m(194) := x"FFF1";
          m(195) := x"0005";
          m(196) := x"FFDE";
          m(197) := x"FFF5";
          m(198) := x"003F";
          m(199) := x"FFE1";
          m(200) := x"FE80";
          m(201) := x"003C";
          m(202) := x"FC05";
          m(203) := x"FE3F";
          m(204) := x"FE08";
          m(205) := x"FD13";
          m(206) := x"005A";
          m(207) := x"FF51";
          m(208) := x"FBCA";
          m(209) := x"FAF3";
          m(210) := x"FCFA";
          m(211) := x"0002";
          m(212) := x"FFA1";
          m(213) := x"FFB1";
          m(214) := x"037D";
          m(215) := x"008A";
          m(216) := x"FFFC";
          m(217) := x"0138";
          m(218) := x"009A";
          m(219) := x"03D9";
          m(220) := x"0344";
          m(221) := x"0384";
          m(222) := x"001E";
          m(223) := x"FFFE";
          m(224) := x"FFAD";
          m(225) := x"FFF4";
          m(226) := x"0096";
          m(227) := x"FFD5";
          m(228) := x"FDCE";
          m(229) := x"FDB6";
          m(230) := x"041E";
          m(231) := x"FEF1";
          m(232) := x"0127";
          m(233) := x"FE9B";
          m(234) := x"FC2C";
          m(235) := x"FF1D";
          m(236) := x"FDDC";
          m(237) := x"FDDF";
          m(238) := x"F984";
          m(239) := x"FF1D";
          m(240) := x"037D";
          m(241) := x"FFC2";
          m(242) := x"00E1";
          m(243) := x"00A6";
          m(244) := x"01E9";
          m(245) := x"0083";
          m(246) := x"00FB";
          m(247) := x"0396";
          m(248) := x"04EF";
          m(249) := x"01B6";
          m(250) := x"FFCC";
          m(251) := x"FFF9";
          m(252) := x"FFE7";
          m(253) := x"FFEB";
          m(254) := x"FF90";
          m(255) := x"0023";
          m(256) := x"FE8F";
          m(257) := x"FBCB";
          m(258) := x"FE03";
          m(259) := x"FD18";
          m(260) := x"FD29";
          m(261) := x"FD16";
          m(262) := x"FA99";
          m(263) := x"FCA6";
          m(264) := x"F7CA";
          m(265) := x"0035";
          m(266) := x"0300";
          m(267) := x"0471";
          m(268) := x"FF8D";
          m(269) := x"01CC";
          m(270) := x"011C";
          m(271) := x"0339";
          m(272) := x"0466";
          m(273) := x"0570";
          m(274) := x"FFB8";
          m(275) := x"00DE";
          m(276) := x"058B";
          m(277) := x"014C";
          m(278) := x"FEA4";
          m(279) := x"FDC9";
          m(280) := x"FFF3";
          m(281) := x"0008";
          m(282) := x"FFD8";
          m(283) := x"003D";
          m(284) := x"0164";
          m(285) := x"FEB3";
          m(286) := x"FBA5";
          m(287) := x"F912";
          m(288) := x"F592";
          m(289) := x"FD99";
          m(290) := x"FB09";
          m(291) := x"01C2";
          m(292) := x"0686";
          m(293) := x"0AA0";
          m(294) := x"0983";
          m(295) := x"0591";
          m(296) := x"0336";
          m(297) := x"00C5";
          m(298) := x"FB5C";
          m(299) := x"00B5";
          m(300) := x"FF06";
          m(301) := x"0399";
          m(302) := x"015F";
          m(303) := x"0368";
          m(304) := x"00F2";
          m(305) := x"FEB0";
          m(306) := x"FE27";
          m(307) := x"FF8B";
          m(308) := x"FFDA";
          m(309) := x"0013";
          m(310) := x"00C3";
          m(311) := x"02D5";
          m(312) := x"04DB";
          m(313) := x"03B0";
          m(314) := x"004B";
          m(315) := x"06EA";
          m(316) := x"060D";
          m(317) := x"0D02";
          m(318) := x"14B8";
          m(319) := x"1687";
          m(320) := x"1D45";
          m(321) := x"0F18";
          m(322) := x"09B0";
          m(323) := x"055C";
          m(324) := x"0047";
          m(325) := x"FFE0";
          m(326) := x"0055";
          m(327) := x"03E1";
          m(328) := x"FDF0";
          m(329) := x"00D8";
          m(330) := x"02B5";
          m(331) := x"0459";
          m(332) := x"012C";
          m(333) := x"006E";
          m(334) := x"008D";
          m(335) := x"FFDD";
          m(336) := x"0030";
          m(337) := x"0028";
          m(338) := x"00DE";
          m(339) := x"0494";
          m(340) := x"0734";
          m(341) := x"0C8D";
          m(342) := x"0D76";
          m(343) := x"1719";
          m(344) := x"1EB7";
          m(345) := x"22E3";
          m(346) := x"185D";
          m(347) := x"0E04";
          m(348) := x"0215";
          m(349) := x"FAF6";
          m(350) := x"FF43";
          m(351) := x"004D";
          m(352) := x"FE34";
          m(353) := x"02D4";
          m(354) := x"FF1A";
          m(355) := x"0359";
          m(356) := x"00BE";
          m(357) := x"0009";
          m(358) := x"03FE";
          m(359) := x"03F7";
          m(360) := x"026E";
          m(361) := x"FD29";
          m(362) := x"005B";
          m(363) := x"FFFC";
          m(364) := x"0017";
          m(365) := x"007A";
          m(366) := x"0046";
          m(367) := x"04EC";
          m(368) := x"0AAC";
          m(369) := x"11CF";
          m(370) := x"1598";
          m(371) := x"1943";
          m(372) := x"14AD";
          m(373) := x"0A97";
          m(374) := x"FD59";
          m(375) := x"FB55";
          m(376) := x"FE97";
          m(377) := x"FA99";
          m(378) := x"008E";
          m(379) := x"0408";
          m(380) := x"0246";
          m(381) := x"FE72";
          m(382) := x"04C8";
          m(383) := x"0493";
          m(384) := x"05E3";
          m(385) := x"FED2";
          m(386) := x"FF20";
          m(387) := x"FD78";
          m(388) := x"FDA9";
          m(389) := x"FC5C";
          m(390) := x"FF6B";
          m(391) := x"FF90";
          m(392) := x"FFE7";
          m(393) := x"0000";
          m(394) := x"FFF1";
          m(395) := x"059A";
          m(396) := x"07FC";
          m(397) := x"0980";
          m(398) := x"06CC";
          m(399) := x"04FE";
          m(400) := x"00E2";
          m(401) := x"F5BA";
          m(402) := x"F894";
          m(403) := x"FC88";
          m(404) := x"F8A0";
          m(405) := x"FB5C";
          m(406) := x"FA67";
          m(407) := x"FC14";
          m(408) := x"FBC5";
          m(409) := x"FFA5";
          m(410) := x"FEB3";
          m(411) := x"FEB6";
          m(412) := x"FF1A";
          m(413) := x"FF8C";
          m(414) := x"0036";
          m(415) := x"FDB0";
          m(416) := x"FDB7";
          m(417) := x"FF5E";
          m(418) := x"FEAA";
          m(419) := x"0020";
          m(420) := x"FFF2";
          m(421) := x"0002";
          m(422) := x"FFEF";
          m(423) := x"02B8";
          m(424) := x"03E5";
          m(425) := x"0084";
          m(426) := x"FD30";
          m(427) := x"FA0F";
          m(428) := x"FD45";
          m(429) := x"FAFE";
          m(430) := x"FB14";
          m(431) := x"FCDA";
          m(432) := x"0216";
          m(433) := x"FF8C";
          m(434) := x"0214";
          m(435) := x"FF50";
          m(436) := x"0049";
          m(437) := x"FF52";
          m(438) := x"0024";
          m(439) := x"00E1";
          m(440) := x"FB4C";
          m(441) := x"F9AB";
          m(442) := x"FE5B";
          m(443) := x"FC9C";
          m(444) := x"FBF9";
          m(445) := x"FFA5";
          m(446) := x"FE7E";
          m(447) := x"FFEC";
          m(448) := x"002C";
          m(449) := x"0009";
          m(450) := x"FF5D";
          m(451) := x"FEEA";
          m(452) := x"FF6F";
          m(453) := x"FCFF";
          m(454) := x"FA78";
          m(455) := x"F8F4";
          m(456) := x"0248";
          m(457) := x"00CF";
          m(458) := x"01A1";
          m(459) := x"03CF";
          m(460) := x"FB02";
          m(461) := x"FC98";
          m(462) := x"FBB2";
          m(463) := x"FF51";
          m(464) := x"FF70";
          m(465) := x"00D6";
          m(466) := x"FBA8";
          m(467) := x"FA2D";
          m(468) := x"FC6A";
          m(469) := x"FC06";
          m(470) := x"000E";
          m(471) := x"FB5B";
          m(472) := x"F9E1";
          m(473) := x"FD7F";
          m(474) := x"FCF8";
          m(475) := x"FFEF";
          m(476) := x"000A";
          m(477) := x"001F";
          m(478) := x"FF28";
          m(479) := x"FD2D";
          m(480) := x"FB44";
          m(481) := x"FABB";
          m(482) := x"012B";
          m(483) := x"02A1";
          m(484) := x"0279";
          m(485) := x"0007";
          m(486) := x"0261";
          m(487) := x"03BA";
          m(488) := x"FE3F";
          m(489) := x"F9AB";
          m(490) := x"FAF4";
          m(491) := x"FAA1";
          m(492) := x"FF97";
          m(493) := x"004D";
          m(494) := x"FEBB";
          m(495) := x"FE57";
          m(496) := x"037C";
          m(497) := x"FF56";
          m(498) := x"FB99";
          m(499) := x"0035";
          m(500) := x"FF96";
          m(501) := x"FE10";
          m(502) := x"FEC9";
          m(503) := x"FFDB";
          m(504) := x"0052";
          m(505) := x"000B";
          m(506) := x"FF9A";
          m(507) := x"FC94";
          m(508) := x"FC84";
          m(509) := x"FCCB";
          m(510) := x"0187";
          m(511) := x"022D";
          m(512) := x"0042";
          m(513) := x"FDE0";
          m(514) := x"0056";
          m(515) := x"0503";
          m(516) := x"FFEC";
          m(517) := x"0047";
          m(518) := x"FD4D";
          m(519) := x"00E4";
          m(520) := x"FF17";
          m(521) := x"FFB9";
          m(522) := x"FF61";
          m(523) := x"FF1E";
          m(524) := x"0383";
          m(525) := x"01D4";
          m(526) := x"FC8E";
          m(527) := x"FE34";
          m(528) := x"FF56";
          m(529) := x"FE36";
          m(530) := x"FF96";
          m(531) := x"FFDA";
          m(532) := x"0022";
          m(533) := x"FFC9";
          m(534) := x"0065";
          m(535) := x"FD63";
          m(536) := x"FF83";
          m(537) := x"FD58";
          m(538) := x"FFE2";
          m(539) := x"0053";
          m(540) := x"00BB";
          m(541) := x"FFE1";
          m(542) := x"FD77";
          m(543) := x"01B3";
          m(544) := x"03EB";
          m(545) := x"FD91";
          m(546) := x"FF4A";
          m(547) := x"011F";
          m(548) := x"FE82";
          m(549) := x"FEA4";
          m(550) := x"FF2C";
          m(551) := x"00BD";
          m(552) := x"0109";
          m(553) := x"FD2C";
          m(554) := x"FC18";
          m(555) := x"FF03";
          m(556) := x"012B";
          m(557) := x"FF26";
          m(558) := x"FFDB";
          m(559) := x"FFD5";
          m(560) := x"000C";
          m(561) := x"0003";
          m(562) := x"0029";
          m(563) := x"FB57";
          m(564) := x"FDEC";
          m(565) := x"FEE6";
          m(566) := x"FDCC";
          m(567) := x"FE8B";
          m(568) := x"01EF";
          m(569) := x"FE89";
          m(570) := x"FDAF";
          m(571) := x"FEBC";
          m(572) := x"01C0";
          m(573) := x"0358";
          m(574) := x"FC7C";
          m(575) := x"03C5";
          m(576) := x"FC87";
          m(577) := x"03DD";
          m(578) := x"0123";
          m(579) := x"00B8";
          m(580) := x"019E";
          m(581) := x"013D";
          m(582) := x"011B";
          m(583) := x"0091";
          m(584) := x"025D";
          m(585) := x"FF7E";
          m(586) := x"FFC6";
          m(587) := x"0003";
          m(588) := x"0002";
          m(589) := x"FFFA";
          m(590) := x"FF4C";
          m(591) := x"FBF4";
          m(592) := x"FCAF";
          m(593) := x"0030";
          m(594) := x"FF93";
          m(595) := x"FE7E";
          m(596) := x"FB65";
          m(597) := x"024C";
          m(598) := x"FEE1";
          m(599) := x"00D4";
          m(600) := x"FB52";
          m(601) := x"0249";
          m(602) := x"0368";
          m(603) := x"FDBA";
          m(604) := x"01A8";
          m(605) := x"010C";
          m(606) := x"FEDA";
          m(607) := x"FEBA";
          m(608) := x"03C8";
          m(609) := x"003F";
          m(610) := x"01A9";
          m(611) := x"FF43";
          m(612) := x"0029";
          m(613) := x"FE40";
          m(614) := x"FFD6";
          m(615) := x"FFDC";
          m(616) := x"FFD5";
          m(617) := x"0001";
          m(618) := x"FF3F";
          m(619) := x"FFA6";
          m(620) := x"FD2B";
          m(621) := x"F944";
          m(622) := x"0279";
          m(623) := x"0047";
          m(624) := x"FFB0";
          m(625) := x"01D1";
          m(626) := x"0185";
          m(627) := x"FDBF";
          m(628) := x"0007";
          m(629) := x"FEF0";
          m(630) := x"FCF0";
          m(631) := x"0011";
          m(632) := x"FC8D";
          m(633) := x"FF73";
          m(634) := x"FF7B";
          m(635) := x"FCD6";
          m(636) := x"FFCB";
          m(637) := x"FF8A";
          m(638) := x"FFC5";
          m(639) := x"FEDE";
          m(640) := x"FE14";
          m(641) := x"FE76";
          m(642) := x"001E";
          m(643) := x"000B";
          m(644) := x"0018";
          m(645) := x"0007";
          m(646) := x"FFD5";
          m(647) := x"0060";
          m(648) := x"FEEA";
          m(649) := x"FB3E";
          m(650) := x"FA78";
          m(651) := x"FC1F";
          m(652) := x"FDD1";
          m(653) := x"FBA4";
          m(654) := x"040C";
          m(655) := x"00FF";
          m(656) := x"022F";
          m(657) := x"FB0F";
          m(658) := x"0078";
          m(659) := x"FC9F";
          m(660) := x"FFAE";
          m(661) := x"02A3";
          m(662) := x"FCFA";
          m(663) := x"FDA3";
          m(664) := x"002B";
          m(665) := x"FE6A";
          m(666) := x"FF6E";
          m(667) := x"FF54";
          m(668) := x"FE46";
          m(669) := x"FEEA";
          m(670) := x"FFFB";
          m(671) := x"0006";
          m(672) := x"FFFA";
          m(673) := x"FFF2";
          m(674) := x"002C";
          m(675) := x"FF4D";
          m(676) := x"FDC0";
          m(677) := x"FE7C";
          m(678) := x"FDAC";
          m(679) := x"FCB7";
          m(680) := x"FF81";
          m(681) := x"FEA6";
          m(682) := x"01BC";
          m(683) := x"0065";
          m(684) := x"00B4";
          m(685) := x"0437";
          m(686) := x"0688";
          m(687) := x"FF48";
          m(688) := x"0321";
          m(689) := x"FF45";
          m(690) := x"018E";
          m(691) := x"0108";
          m(692) := x"00A9";
          m(693) := x"01A1";
          m(694) := x"01A4";
          m(695) := x"01EC";
          m(696) := x"FF7E";
          m(697) := x"FFB5";
          m(698) := x"0005";
          m(699) := x"000C";
          m(700) := x"0004";
          m(701) := x"FFEF";
          m(702) := x"000B";
          m(703) := x"FFEB";
          m(704) := x"FF49";
          m(705) := x"FF1D";
          m(706) := x"FE2C";
          m(707) := x"FEEF";
          m(708) := x"FD5B";
          m(709) := x"FD1D";
          m(710) := x"004D";
          m(711) := x"016A";
          m(712) := x"FDD0";
          m(713) := x"02C2";
          m(714) := x"02C4";
          m(715) := x"FEB1";
          m(716) := x"003B";
          m(717) := x"032C";
          m(718) := x"03F7";
          m(719) := x"0075";
          m(720) := x"0192";
          m(721) := x"0491";
          m(722) := x"01A2";
          m(723) := x"003D";
          m(724) := x"FFE8";
          m(725) := x"FFE8";
          m(726) := x"FFDD";
          m(727) := x"FFE3";
          m(728) := x"0006";
          m(729) := x"FFDB";
          m(730) := x"FFC1";
          m(731) := x"0017";
          m(732) := x"0024";
          m(733) := x"027E";
          m(734) := x"0225";
          m(735) := x"FFED";
          m(736) := x"00A0";
          m(737) := x"01F3";
          m(738) := x"003D";
          m(739) := x"FF2B";
          m(740) := x"FDBE";
          m(741) := x"FF86";
          m(742) := x"01B1";
          m(743) := x"00C2";
          m(744) := x"00F7";
          m(745) := x"023C";
          m(746) := x"024B";
          m(747) := x"0192";
          m(748) := x"016E";
          m(749) := x"01E5";
          m(750) := x"00FE";
          m(751) := x"0019";
          m(752) := x"FFF0";
          m(753) := x"0032";
          m(754) := x"0026";
          m(755) := x"FFF9";
          m(756) := x"0001";
          m(757) := x"0000";
          m(758) := x"FFE6";
          m(759) := x"0009";
          m(760) := x"FFE3";
          m(761) := x"0001";
          m(762) := x"FFC7";
          m(763) := x"FFDA";
          m(764) := x"0008";
          m(765) := x"FFEE";
          m(766) := x"000E";
          m(767) := x"0017";
          m(768) := x"000D";
          m(769) := x"0028";
          m(770) := x"0015";
          m(771) := x"FFD8";
          m(772) := x"FFDA";
          m(773) := x"FFEF";
          m(774) := x"0089";
          m(775) := x"002B";
          m(776) := x"0087";
          m(777) := x"0022";
          m(778) := x"015B";
          m(779) := x"FFFB";
          m(780) := x"FFC1";
          m(781) := x"0024";
          m(782) := x"0006";
          m(783) := x"FFE6";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_22.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 22) then
          m(0) := x"FFF9";
          m(1) := x"FFF6";
          m(2) := x"003E";
          m(3) := x"FFFE";
          m(4) := x"0000";
          m(5) := x"FFF1";
          m(6) := x"FFF8";
          m(7) := x"0006";
          m(8) := x"FFD5";
          m(9) := x"0028";
          m(10) := x"0011";
          m(11) := x"0022";
          m(12) := x"FFE5";
          m(13) := x"FFEF";
          m(14) := x"003A";
          m(15) := x"FFA5";
          m(16) := x"000B";
          m(17) := x"FFD5";
          m(18) := x"0014";
          m(19) := x"FFD1";
          m(20) := x"0013";
          m(21) := x"002A";
          m(22) := x"0026";
          m(23) := x"000F";
          m(24) := x"FFD0";
          m(25) := x"0001";
          m(26) := x"FFF4";
          m(27) := x"FFDE";
          m(28) := x"FFF9";
          m(29) := x"FFCC";
          m(30) := x"FFE3";
          m(31) := x"001D";
          m(32) := x"0021";
          m(33) := x"FFFB";
          m(34) := x"0009";
          m(35) := x"003F";
          m(36) := x"FFED";
          m(37) := x"FFFE";
          m(38) := x"002B";
          m(39) := x"FFFD";
          m(40) := x"000D";
          m(41) := x"0013";
          m(42) := x"FFFB";
          m(43) := x"FFFE";
          m(44) := x"FF60";
          m(45) := x"FF87";
          m(46) := x"FFE9";
          m(47) := x"0006";
          m(48) := x"0005";
          m(49) := x"FFEC";
          m(50) := x"FFE5";
          m(51) := x"001F";
          m(52) := x"FFE6";
          m(53) := x"0039";
          m(54) := x"FFEA";
          m(55) := x"0019";
          m(56) := x"000D";
          m(57) := x"0001";
          m(58) := x"FFF5";
          m(59) := x"FFD1";
          m(60) := x"FFDE";
          m(61) := x"001E";
          m(62) := x"0024";
          m(63) := x"006A";
          m(64) := x"0049";
          m(65) := x"002B";
          m(66) := x"001D";
          m(67) := x"00B7";
          m(68) := x"009C";
          m(69) := x"FFF9";
          m(70) := x"0063";
          m(71) := x"002F";
          m(72) := x"000B";
          m(73) := x"006E";
          m(74) := x"00B5";
          m(75) := x"004F";
          m(76) := x"001E";
          m(77) := x"005B";
          m(78) := x"0063";
          m(79) := x"FFFB";
          m(80) := x"001B";
          m(81) := x"FFDE";
          m(82) := x"FFF1";
          m(83) := x"0031";
          m(84) := x"FFED";
          m(85) := x"FFD2";
          m(86) := x"0017";
          m(87) := x"FFF8";
          m(88) := x"001F";
          m(89) := x"001B";
          m(90) := x"007C";
          m(91) := x"FF75";
          m(92) := x"FF83";
          m(93) := x"FFEB";
          m(94) := x"FF84";
          m(95) := x"00B9";
          m(96) := x"00F2";
          m(97) := x"00B4";
          m(98) := x"01CB";
          m(99) := x"01A3";
          m(100) := x"0119";
          m(101) := x"0066";
          m(102) := x"0125";
          m(103) := x"00E3";
          m(104) := x"00FF";
          m(105) := x"00D1";
          m(106) := x"005B";
          m(107) := x"0025";
          m(108) := x"FFEB";
          m(109) := x"FF9A";
          m(110) := x"FFF0";
          m(111) := x"004C";
          m(112) := x"FFE5";
          m(113) := x"FFF6";
          m(114) := x"0014";
          m(115) := x"002C";
          m(116) := x"FFEF";
          m(117) := x"0017";
          m(118) := x"FFA4";
          m(119) := x"FFE7";
          m(120) := x"FFF8";
          m(121) := x"FFBD";
          m(122) := x"00D8";
          m(123) := x"01C7";
          m(124) := x"0479";
          m(125) := x"04CB";
          m(126) := x"0527";
          m(127) := x"03E8";
          m(128) := x"033A";
          m(129) := x"0248";
          m(130) := x"01CC";
          m(131) := x"0298";
          m(132) := x"0230";
          m(133) := x"010E";
          m(134) := x"FFA9";
          m(135) := x"FF57";
          m(136) := x"FFA7";
          m(137) := x"0016";
          m(138) := x"0010";
          m(139) := x"FFF5";
          m(140) := x"000F";
          m(141) := x"0015";
          m(142) := x"0001";
          m(143) := x"FFF1";
          m(144) := x"FFBB";
          m(145) := x"FF26";
          m(146) := x"FF36";
          m(147) := x"00E2";
          m(148) := x"01E2";
          m(149) := x"02DB";
          m(150) := x"0193";
          m(151) := x"033B";
          m(152) := x"0391";
          m(153) := x"04BF";
          m(154) := x"0B20";
          m(155) := x"09A3";
          m(156) := x"0BFB";
          m(157) := x"08C2";
          m(158) := x"0612";
          m(159) := x"0228";
          m(160) := x"FF2D";
          m(161) := x"00A3";
          m(162) := x"FFB2";
          m(163) := x"002C";
          m(164) := x"FFEF";
          m(165) := x"FFA4";
          m(166) := x"FFD3";
          m(167) := x"0016";
          m(168) := x"0013";
          m(169) := x"FFBA";
          m(170) := x"FFCB";
          m(171) := x"FF7C";
          m(172) := x"0029";
          m(173) := x"01D1";
          m(174) := x"01A2";
          m(175) := x"0200";
          m(176) := x"019C";
          m(177) := x"0199";
          m(178) := x"02AD";
          m(179) := x"02D8";
          m(180) := x"05DB";
          m(181) := x"FFB4";
          m(182) := x"01EF";
          m(183) := x"004B";
          m(184) := x"004C";
          m(185) := x"FC6D";
          m(186) := x"FAC3";
          m(187) := x"02B7";
          m(188) := x"FA9F";
          m(189) := x"FEDA";
          m(190) := x"050A";
          m(191) := x"07AD";
          m(192) := x"02A8";
          m(193) := x"0099";
          m(194) := x"FFE4";
          m(195) := x"FFEC";
          m(196) := x"0014";
          m(197) := x"003D";
          m(198) := x"FF4F";
          m(199) := x"FF02";
          m(200) := x"00BC";
          m(201) := x"0270";
          m(202) := x"0210";
          m(203) := x"0567";
          m(204) := x"0091";
          m(205) := x"FE83";
          m(206) := x"FD79";
          m(207) := x"011F";
          m(208) := x"FD9A";
          m(209) := x"FA46";
          m(210) := x"F695";
          m(211) := x"F489";
          m(212) := x"FA87";
          m(213) := x"F910";
          m(214) := x"F95F";
          m(215) := x"FCB9";
          m(216) := x"FE4A";
          m(217) := x"02D2";
          m(218) := x"073B";
          m(219) := x"0945";
          m(220) := x"04EB";
          m(221) := x"0215";
          m(222) := x"00BC";
          m(223) := x"FFF7";
          m(224) := x"FFD7";
          m(225) := x"FFF9";
          m(226) := x"FFB4";
          m(227) := x"FF16";
          m(228) := x"00D7";
          m(229) := x"0066";
          m(230) := x"0293";
          m(231) := x"02A9";
          m(232) := x"FCE2";
          m(233) := x"FC74";
          m(234) := x"FFF2";
          m(235) := x"FC44";
          m(236) := x"F807";
          m(237) := x"F805";
          m(238) := x"F56A";
          m(239) := x"F6C7";
          m(240) := x"F61E";
          m(241) := x"F995";
          m(242) := x"FC66";
          m(243) := x"01C8";
          m(244) := x"0219";
          m(245) := x"0115";
          m(246) := x"05CF";
          m(247) := x"088C";
          m(248) := x"0610";
          m(249) := x"02DF";
          m(250) := x"0026";
          m(251) := x"0004";
          m(252) := x"0019";
          m(253) := x"FFFE";
          m(254) := x"0023";
          m(255) := x"FE24";
          m(256) := x"FED2";
          m(257) := x"00D3";
          m(258) := x"FC7A";
          m(259) := x"FD7A";
          m(260) := x"FC61";
          m(261) := x"FA43";
          m(262) := x"FCF0";
          m(263) := x"FC3C";
          m(264) := x"F9D2";
          m(265) := x"F8EA";
          m(266) := x"FB39";
          m(267) := x"FA8E";
          m(268) := x"FC8E";
          m(269) := x"01F0";
          m(270) := x"05CD";
          m(271) := x"0716";
          m(272) := x"0306";
          m(273) := x"030C";
          m(274) := x"031F";
          m(275) := x"0944";
          m(276) := x"0536";
          m(277) := x"01A0";
          m(278) := x"00A7";
          m(279) := x"FFDB";
          m(280) := x"FFE6";
          m(281) := x"FFDF";
          m(282) := x"0023";
          m(283) := x"FE43";
          m(284) := x"0059";
          m(285) := x"FEC3";
          m(286) := x"FA7E";
          m(287) := x"FC8B";
          m(288) := x"FC04";
          m(289) := x"F6C1";
          m(290) := x"0138";
          m(291) := x"0052";
          m(292) := x"00E3";
          m(293) := x"FFFE";
          m(294) := x"0326";
          m(295) := x"0843";
          m(296) := x"01E1";
          m(297) := x"04E5";
          m(298) := x"0275";
          m(299) := x"0000";
          m(300) := x"FF48";
          m(301) := x"FF4C";
          m(302) := x"023F";
          m(303) := x"0407";
          m(304) := x"02E8";
          m(305) := x"010B";
          m(306) := x"FFFF";
          m(307) := x"FFDA";
          m(308) := x"001D";
          m(309) := x"001D";
          m(310) := x"FFA2";
          m(311) := x"FE12";
          m(312) := x"FE08";
          m(313) := x"FC58";
          m(314) := x"FC2C";
          m(315) := x"FE88";
          m(316) := x"FEED";
          m(317) := x"01ED";
          m(318) := x"0739";
          m(319) := x"FC17";
          m(320) := x"FFE5";
          m(321) := x"02B8";
          m(322) := x"0054";
          m(323) := x"02DD";
          m(324) := x"FCE2";
          m(325) := x"FAFF";
          m(326) := x"F9F6";
          m(327) := x"FC6B";
          m(328) := x"F971";
          m(329) := x"FCFE";
          m(330) := x"FECE";
          m(331) := x"0027";
          m(332) := x"FE7E";
          m(333) := x"00A1";
          m(334) := x"FF73";
          m(335) := x"FFDE";
          m(336) := x"FFEE";
          m(337) := x"000A";
          m(338) := x"FF9B";
          m(339) := x"FFA4";
          m(340) := x"FBE8";
          m(341) := x"FF6D";
          m(342) := x"FEEB";
          m(343) := x"033F";
          m(344) := x"0437";
          m(345) := x"00F2";
          m(346) := x"02FA";
          m(347) := x"0041";
          m(348) := x"07A1";
          m(349) := x"08A7";
          m(350) := x"0297";
          m(351) := x"FDFC";
          m(352) := x"0562";
          m(353) := x"FB54";
          m(354) := x"FC78";
          m(355) := x"0293";
          m(356) := x"011B";
          m(357) := x"01D1";
          m(358) := x"0337";
          m(359) := x"FED5";
          m(360) := x"022C";
          m(361) := x"0102";
          m(362) := x"FF4A";
          m(363) := x"001F";
          m(364) := x"FFF1";
          m(365) := x"FFFF";
          m(366) := x"FFD3";
          m(367) := x"0031";
          m(368) := x"FF8F";
          m(369) := x"038A";
          m(370) := x"0161";
          m(371) := x"01D0";
          m(372) := x"0211";
          m(373) := x"FF62";
          m(374) := x"0151";
          m(375) := x"000F";
          m(376) := x"0344";
          m(377) := x"FDAD";
          m(378) := x"FBBD";
          m(379) := x"FBB4";
          m(380) := x"FFE5";
          m(381) := x"0158";
          m(382) := x"FFA4";
          m(383) := x"0338";
          m(384) := x"01A6";
          m(385) := x"FFB1";
          m(386) := x"037F";
          m(387) := x"02C6";
          m(388) := x"038D";
          m(389) := x"0117";
          m(390) := x"009C";
          m(391) := x"0002";
          m(392) := x"0002";
          m(393) := x"0002";
          m(394) := x"FFFF";
          m(395) := x"00A5";
          m(396) := x"0180";
          m(397) := x"08CB";
          m(398) := x"021B";
          m(399) := x"04C9";
          m(400) := x"FE38";
          m(401) := x"0391";
          m(402) := x"00BE";
          m(403) := x"0519";
          m(404) := x"057F";
          m(405) := x"01A8";
          m(406) := x"01E2";
          m(407) := x"FA62";
          m(408) := x"FF34";
          m(409) := x"04E7";
          m(410) := x"FDEB";
          m(411) := x"FF31";
          m(412) := x"FB72";
          m(413) := x"0088";
          m(414) := x"05E2";
          m(415) := x"054E";
          m(416) := x"0438";
          m(417) := x"0130";
          m(418) := x"005B";
          m(419) := x"FFE8";
          m(420) := x"FFE3";
          m(421) := x"000A";
          m(422) := x"009A";
          m(423) := x"0218";
          m(424) := x"0271";
          m(425) := x"0496";
          m(426) := x"022A";
          m(427) := x"00AB";
          m(428) := x"F898";
          m(429) := x"01CE";
          m(430) := x"0362";
          m(431) := x"FD35";
          m(432) := x"FFC3";
          m(433) := x"01F0";
          m(434) := x"020E";
          m(435) := x"008F";
          m(436) := x"FF9F";
          m(437) := x"FE57";
          m(438) := x"FEAD";
          m(439) := x"0347";
          m(440) := x"FD44";
          m(441) := x"FFDE";
          m(442) := x"052C";
          m(443) := x"02C8";
          m(444) := x"0271";
          m(445) := x"022C";
          m(446) := x"0061";
          m(447) := x"007C";
          m(448) := x"004E";
          m(449) := x"FFEB";
          m(450) := x"FFF8";
          m(451) := x"014A";
          m(452) := x"0150";
          m(453) := x"064D";
          m(454) := x"0496";
          m(455) := x"0028";
          m(456) := x"0006";
          m(457) := x"FF46";
          m(458) := x"FD18";
          m(459) := x"FB9C";
          m(460) := x"FE75";
          m(461) := x"0235";
          m(462) := x"03C5";
          m(463) := x"07AF";
          m(464) := x"056F";
          m(465) := x"0255";
          m(466) := x"02F7";
          m(467) := x"05D3";
          m(468) := x"02B7";
          m(469) := x"033B";
          m(470) := x"FFF2";
          m(471) := x"0280";
          m(472) := x"02DB";
          m(473) := x"0364";
          m(474) := x"00EB";
          m(475) := x"FFEA";
          m(476) := x"0002";
          m(477) := x"FFEC";
          m(478) := x"FFE2";
          m(479) := x"FFEB";
          m(480) := x"02A3";
          m(481) := x"06E1";
          m(482) := x"0632";
          m(483) := x"FE21";
          m(484) := x"FC6A";
          m(485) := x"0022";
          m(486) := x"FE94";
          m(487) := x"FF32";
          m(488) := x"FE8C";
          m(489) := x"0266";
          m(490) := x"03D3";
          m(491) := x"FFF1";
          m(492) := x"0174";
          m(493) := x"0230";
          m(494) := x"0164";
          m(495) := x"FFC3";
          m(496) := x"FD00";
          m(497) := x"FE8F";
          m(498) := x"029F";
          m(499) := x"02CA";
          m(500) := x"01B9";
          m(501) := x"02BB";
          m(502) := x"009C";
          m(503) := x"FFEF";
          m(504) := x"FFF7";
          m(505) := x"FFB1";
          m(506) := x"0004";
          m(507) := x"00F1";
          m(508) := x"03C6";
          m(509) := x"0820";
          m(510) := x"07A8";
          m(511) := x"0145";
          m(512) := x"FF37";
          m(513) := x"0151";
          m(514) := x"FBFD";
          m(515) := x"FDBC";
          m(516) := x"02A1";
          m(517) := x"0011";
          m(518) := x"0055";
          m(519) := x"005C";
          m(520) := x"058A";
          m(521) := x"015B";
          m(522) := x"01AE";
          m(523) := x"FF29";
          m(524) := x"FC00";
          m(525) := x"FF87";
          m(526) := x"00F0";
          m(527) := x"0284";
          m(528) := x"0300";
          m(529) := x"0103";
          m(530) := x"000B";
          m(531) := x"0030";
          m(532) := x"001A";
          m(533) := x"FFEA";
          m(534) := x"FFC1";
          m(535) := x"028B";
          m(536) := x"0586";
          m(537) := x"0689";
          m(538) := x"0627";
          m(539) := x"0363";
          m(540) := x"FEA1";
          m(541) := x"0156";
          m(542) := x"0107";
          m(543) := x"FF62";
          m(544) := x"FA18";
          m(545) := x"01BC";
          m(546) := x"FDC7";
          m(547) := x"0010";
          m(548) := x"026D";
          m(549) := x"00FD";
          m(550) := x"03B4";
          m(551) := x"FE04";
          m(552) := x"FFA1";
          m(553) := x"FDD3";
          m(554) := x"FF1B";
          m(555) := x"0190";
          m(556) := x"0080";
          m(557) := x"004D";
          m(558) := x"0042";
          m(559) := x"FFF4";
          m(560) := x"001A";
          m(561) := x"FFD2";
          m(562) := x"FFFE";
          m(563) := x"018E";
          m(564) := x"04B6";
          m(565) := x"030C";
          m(566) := x"06EA";
          m(567) := x"081F";
          m(568) := x"06FA";
          m(569) := x"05B8";
          m(570) := x"0619";
          m(571) := x"049D";
          m(572) := x"01D1";
          m(573) := x"019C";
          m(574) := x"F94F";
          m(575) := x"FCA3";
          m(576) := x"FE5B";
          m(577) := x"FFAF";
          m(578) := x"04BA";
          m(579) := x"FE17";
          m(580) := x"FD27";
          m(581) := x"FE4D";
          m(582) := x"FCF7";
          m(583) := x"0033";
          m(584) := x"FF57";
          m(585) := x"FE8E";
          m(586) := x"0024";
          m(587) := x"FFE9";
          m(588) := x"FFE9";
          m(589) := x"FFDA";
          m(590) := x"FFD1";
          m(591) := x"0062";
          m(592) := x"00EB";
          m(593) := x"022B";
          m(594) := x"0420";
          m(595) := x"0687";
          m(596) := x"0A3F";
          m(597) := x"0A69";
          m(598) := x"0637";
          m(599) := x"0BA6";
          m(600) := x"04D4";
          m(601) := x"056A";
          m(602) := x"FBCB";
          m(603) := x"FD3A";
          m(604) := x"FDF8";
          m(605) := x"0127";
          m(606) := x"04A8";
          m(607) := x"FF57";
          m(608) := x"FC75";
          m(609) := x"0185";
          m(610) := x"FF17";
          m(611) := x"0119";
          m(612) := x"FE77";
          m(613) := x"0045";
          m(614) := x"0058";
          m(615) := x"0001";
          m(616) := x"0023";
          m(617) := x"FFFB";
          m(618) := x"005B";
          m(619) := x"005E";
          m(620) := x"FF9C";
          m(621) := x"FF49";
          m(622) := x"FF5D";
          m(623) := x"018C";
          m(624) := x"04A8";
          m(625) := x"03BF";
          m(626) := x"002B";
          m(627) := x"0694";
          m(628) := x"03A3";
          m(629) := x"0807";
          m(630) := x"0036";
          m(631) := x"0392";
          m(632) := x"019E";
          m(633) := x"0684";
          m(634) := x"0751";
          m(635) := x"03BF";
          m(636) := x"FFCE";
          m(637) := x"01A1";
          m(638) := x"FC63";
          m(639) := x"FCC2";
          m(640) := x"FEAA";
          m(641) := x"FF6C";
          m(642) := x"0026";
          m(643) := x"0000";
          m(644) := x"001F";
          m(645) := x"FFD5";
          m(646) := x"004B";
          m(647) := x"0009";
          m(648) := x"0011";
          m(649) := x"FEB6";
          m(650) := x"FE1C";
          m(651) := x"FE1A";
          m(652) := x"FF6B";
          m(653) := x"01E8";
          m(654) := x"FE2C";
          m(655) := x"0076";
          m(656) := x"01A1";
          m(657) := x"0184";
          m(658) := x"084B";
          m(659) := x"0807";
          m(660) := x"0677";
          m(661) := x"0638";
          m(662) := x"0A40";
          m(663) := x"0300";
          m(664) := x"FF2C";
          m(665) := x"0255";
          m(666) := x"FDA2";
          m(667) := x"FCDE";
          m(668) := x"FDE5";
          m(669) := x"00FE";
          m(670) := x"001D";
          m(671) := x"FFD4";
          m(672) := x"0000";
          m(673) := x"0057";
          m(674) := x"FFEB";
          m(675) := x"FFA8";
          m(676) := x"FF0F";
          m(677) := x"FEC1";
          m(678) := x"FE7F";
          m(679) := x"FB75";
          m(680) := x"FAA2";
          m(681) := x"FD66";
          m(682) := x"FB4C";
          m(683) := x"FF12";
          m(684) := x"FF2D";
          m(685) := x"0182";
          m(686) := x"050A";
          m(687) := x"0088";
          m(688) := x"0852";
          m(689) := x"0639";
          m(690) := x"07C1";
          m(691) := x"0168";
          m(692) := x"FBEC";
          m(693) := x"0104";
          m(694) := x"0004";
          m(695) := x"FDE7";
          m(696) := x"0083";
          m(697) := x"00F8";
          m(698) := x"FFF3";
          m(699) := x"FFFF";
          m(700) := x"FFFC";
          m(701) := x"0002";
          m(702) := x"FFD9";
          m(703) := x"FFF5";
          m(704) := x"FF6D";
          m(705) := x"FDA8";
          m(706) := x"FD26";
          m(707) := x"FB3A";
          m(708) := x"F98B";
          m(709) := x"FA0A";
          m(710) := x"FF04";
          m(711) := x"FEDD";
          m(712) := x"FDA7";
          m(713) := x"01C9";
          m(714) := x"FD2C";
          m(715) := x"FE82";
          m(716) := x"FA91";
          m(717) := x"FB7B";
          m(718) := x"FC1C";
          m(719) := x"F83E";
          m(720) := x"FB6F";
          m(721) := x"FE23";
          m(722) := x"001D";
          m(723) := x"FFA7";
          m(724) := x"FFCB";
          m(725) := x"FFE8";
          m(726) := x"FFFE";
          m(727) := x"FFE9";
          m(728) := x"FFF4";
          m(729) := x"FFF2";
          m(730) := x"0034";
          m(731) := x"0026";
          m(732) := x"FF47";
          m(733) := x"FE86";
          m(734) := x"FE42";
          m(735) := x"FDA7";
          m(736) := x"FE62";
          m(737) := x"FC88";
          m(738) := x"FCA9";
          m(739) := x"FDEB";
          m(740) := x"FB73";
          m(741) := x"FA76";
          m(742) := x"F639";
          m(743) := x"FA3B";
          m(744) := x"F948";
          m(745) := x"F995";
          m(746) := x"F9B4";
          m(747) := x"FDA1";
          m(748) := x"FCE9";
          m(749) := x"FD4B";
          m(750) := x"FF5F";
          m(751) := x"FFEB";
          m(752) := x"FFCE";
          m(753) := x"FFF1";
          m(754) := x"0002";
          m(755) := x"FFFA";
          m(756) := x"FFEB";
          m(757) := x"0015";
          m(758) := x"0009";
          m(759) := x"FFFD";
          m(760) := x"FFC9";
          m(761) := x"FFF0";
          m(762) := x"FFD6";
          m(763) := x"FF86";
          m(764) := x"FF7B";
          m(765) := x"FFD6";
          m(766) := x"FF8D";
          m(767) := x"FF5F";
          m(768) := x"FE60";
          m(769) := x"FF77";
          m(770) := x"FED9";
          m(771) := x"FEAE";
          m(772) := x"FF11";
          m(773) := x"FF4E";
          m(774) := x"FDFB";
          m(775) := x"FFC9";
          m(776) := x"FFF6";
          m(777) := x"001C";
          m(778) := x"FFBD";
          m(779) := x"FFE6";
          m(780) := x"FFCD";
          m(781) := x"FFFD";
          m(782) := x"FFA2";
          m(783) := x"FFF0";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_23.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 23) then
          m(0) := x"FFDA";
          m(1) := x"000A";
          m(2) := x"FFFF";
          m(3) := x"FFFC";
          m(4) := x"002D";
          m(5) := x"FFD8";
          m(6) := x"0011";
          m(7) := x"000E";
          m(8) := x"FFEE";
          m(9) := x"FFF5";
          m(10) := x"FFDC";
          m(11) := x"0022";
          m(12) := x"000A";
          m(13) := x"FFC9";
          m(14) := x"FFDB";
          m(15) := x"FFD4";
          m(16) := x"0000";
          m(17) := x"0001";
          m(18) := x"001E";
          m(19) := x"FFE3";
          m(20) := x"0012";
          m(21) := x"0032";
          m(22) := x"FFDE";
          m(23) := x"0013";
          m(24) := x"FFF1";
          m(25) := x"000B";
          m(26) := x"0002";
          m(27) := x"0000";
          m(28) := x"001B";
          m(29) := x"0028";
          m(30) := x"FFFD";
          m(31) := x"FFFB";
          m(32) := x"0016";
          m(33) := x"000E";
          m(34) := x"0017";
          m(35) := x"FFEE";
          m(36) := x"0020";
          m(37) := x"0000";
          m(38) := x"FFFF";
          m(39) := x"FFE4";
          m(40) := x"FFE7";
          m(41) := x"FFC7";
          m(42) := x"FFBE";
          m(43) := x"0032";
          m(44) := x"0009";
          m(45) := x"0000";
          m(46) := x"0000";
          m(47) := x"FFEA";
          m(48) := x"FFE0";
          m(49) := x"FFFF";
          m(50) := x"FFBD";
          m(51) := x"0001";
          m(52) := x"000A";
          m(53) := x"FFF5";
          m(54) := x"FFA5";
          m(55) := x"003D";
          m(56) := x"0008";
          m(57) := x"FFF4";
          m(58) := x"001E";
          m(59) := x"FFE3";
          m(60) := x"001B";
          m(61) := x"0002";
          m(62) := x"000B";
          m(63) := x"0034";
          m(64) := x"001B";
          m(65) := x"FFDB";
          m(66) := x"FF95";
          m(67) := x"FEF2";
          m(68) := x"FEAA";
          m(69) := x"FDD5";
          m(70) := x"FEC3";
          m(71) := x"FF2C";
          m(72) := x"0007";
          m(73) := x"FF9A";
          m(74) := x"0040";
          m(75) := x"012C";
          m(76) := x"0050";
          m(77) := x"005E";
          m(78) := x"FFF5";
          m(79) := x"FFF8";
          m(80) := x"FFD7";
          m(81) := x"0017";
          m(82) := x"0005";
          m(83) := x"FFD7";
          m(84) := x"FFFF";
          m(85) := x"FFF4";
          m(86) := x"FFF9";
          m(87) := x"FFB4";
          m(88) := x"0018";
          m(89) := x"FFFB";
          m(90) := x"FFF3";
          m(91) := x"005A";
          m(92) := x"013A";
          m(93) := x"010A";
          m(94) := x"000D";
          m(95) := x"FC51";
          m(96) := x"FE43";
          m(97) := x"009F";
          m(98) := x"FEB8";
          m(99) := x"FF73";
          m(100) := x"FE2B";
          m(101) := x"FCD2";
          m(102) := x"FEB5";
          m(103) := x"02B0";
          m(104) := x"FF41";
          m(105) := x"FE54";
          m(106) := x"FCE9";
          m(107) := x"FE8D";
          m(108) := x"00DA";
          m(109) := x"0025";
          m(110) := x"FFF9";
          m(111) := x"FFFE";
          m(112) := x"FFEF";
          m(113) := x"FFFD";
          m(114) := x"FFC5";
          m(115) := x"0019";
          m(116) := x"0055";
          m(117) := x"008E";
          m(118) := x"0095";
          m(119) := x"FFE5";
          m(120) := x"FC0A";
          m(121) := x"FBA8";
          m(122) := x"FC6C";
          m(123) := x"FE62";
          m(124) := x"FF19";
          m(125) := x"FAE0";
          m(126) := x"FC9C";
          m(127) := x"023A";
          m(128) := x"0192";
          m(129) := x"FBA4";
          m(130) := x"FE51";
          m(131) := x"FFFA";
          m(132) := x"FE94";
          m(133) := x"0327";
          m(134) := x"018F";
          m(135) := x"007C";
          m(136) := x"0177";
          m(137) := x"00DF";
          m(138) := x"000F";
          m(139) := x"0023";
          m(140) := x"FFCB";
          m(141) := x"000E";
          m(142) := x"0018";
          m(143) := x"FFBE";
          m(144) := x"FFF6";
          m(145) := x"0448";
          m(146) := x"032C";
          m(147) := x"FF4E";
          m(148) := x"0218";
          m(149) := x"0475";
          m(150) := x"0647";
          m(151) := x"0489";
          m(152) := x"FE9B";
          m(153) := x"018D";
          m(154) := x"FB63";
          m(155) := x"FBDB";
          m(156) := x"02DC";
          m(157) := x"02D9";
          m(158) := x"0391";
          m(159) := x"00F9";
          m(160) := x"0310";
          m(161) := x"0233";
          m(162) := x"0368";
          m(163) := x"0302";
          m(164) := x"FEB5";
          m(165) := x"003C";
          m(166) := x"0037";
          m(167) := x"0000";
          m(168) := x"0004";
          m(169) := x"0000";
          m(170) := x"0066";
          m(171) := x"0011";
          m(172) := x"0039";
          m(173) := x"0620";
          m(174) := x"04CA";
          m(175) := x"0278";
          m(176) := x"0182";
          m(177) := x"02DE";
          m(178) := x"02E8";
          m(179) := x"0023";
          m(180) := x"FF90";
          m(181) := x"FD3C";
          m(182) := x"0152";
          m(183) := x"FD60";
          m(184) := x"FFEE";
          m(185) := x"FF1F";
          m(186) := x"011B";
          m(187) := x"03E0";
          m(188) := x"01A0";
          m(189) := x"0387";
          m(190) := x"04B3";
          m(191) := x"05A6";
          m(192) := x"04F7";
          m(193) := x"036D";
          m(194) := x"0136";
          m(195) := x"0013";
          m(196) := x"004D";
          m(197) := x"000A";
          m(198) := x"0024";
          m(199) := x"FFE9";
          m(200) := x"FE34";
          m(201) := x"04F0";
          m(202) := x"00CB";
          m(203) := x"0077";
          m(204) := x"01F2";
          m(205) := x"0007";
          m(206) := x"03A1";
          m(207) := x"0351";
          m(208) := x"00E6";
          m(209) := x"FC43";
          m(210) := x"FF01";
          m(211) := x"02E8";
          m(212) := x"06A7";
          m(213) := x"04B8";
          m(214) := x"0513";
          m(215) := x"047B";
          m(216) := x"09F6";
          m(217) := x"05E1";
          m(218) := x"FF17";
          m(219) := x"0302";
          m(220) := x"057D";
          m(221) := x"01FA";
          m(222) := x"0149";
          m(223) := x"0027";
          m(224) := x"FFE1";
          m(225) := x"003D";
          m(226) := x"FFBF";
          m(227) := x"FFA2";
          m(228) := x"FD8E";
          m(229) := x"0181";
          m(230) := x"FCC9";
          m(231) := x"FE95";
          m(232) := x"FBF6";
          m(233) := x"0216";
          m(234) := x"0133";
          m(235) := x"01CA";
          m(236) := x"02A8";
          m(237) := x"0295";
          m(238) := x"FE4F";
          m(239) := x"06B0";
          m(240) := x"0482";
          m(241) := x"010F";
          m(242) := x"050B";
          m(243) := x"069F";
          m(244) := x"01CC";
          m(245) := x"FD05";
          m(246) := x"FE2C";
          m(247) := x"0191";
          m(248) := x"01FC";
          m(249) := x"FF68";
          m(250) := x"00E1";
          m(251) := x"FFF3";
          m(252) := x"FFCE";
          m(253) := x"002E";
          m(254) := x"0030";
          m(255) := x"FEAD";
          m(256) := x"FFEB";
          m(257) := x"FFE0";
          m(258) := x"FE17";
          m(259) := x"007A";
          m(260) := x"00F3";
          m(261) := x"0065";
          m(262) := x"FF26";
          m(263) := x"01D6";
          m(264) := x"00A1";
          m(265) := x"F59D";
          m(266) := x"F3FE";
          m(267) := x"F649";
          m(268) := x"F7B4";
          m(269) := x"F594";
          m(270) := x"F907";
          m(271) := x"F6D1";
          m(272) := x"F634";
          m(273) := x"F484";
          m(274) := x"F747";
          m(275) := x"F8DD";
          m(276) := x"FE77";
          m(277) := x"FF8B";
          m(278) := x"008E";
          m(279) := x"001A";
          m(280) := x"FFB9";
          m(281) := x"000B";
          m(282) := x"0016";
          m(283) := x"FEC5";
          m(284) := x"0052";
          m(285) := x"012D";
          m(286) := x"FF9C";
          m(287) := x"FD9A";
          m(288) := x"FF0D";
          m(289) := x"02ED";
          m(290) := x"FF1C";
          m(291) := x"00AB";
          m(292) := x"0156";
          m(293) := x"F8B1";
          m(294) := x"F1FD";
          m(295) := x"F03E";
          m(296) := x"EF0A";
          m(297) := x"EA83";
          m(298) := x"EA06";
          m(299) := x"E8F5";
          m(300) := x"EF90";
          m(301) := x"F3E0";
          m(302) := x"F328";
          m(303) := x"F214";
          m(304) := x"FB7E";
          m(305) := x"FF7F";
          m(306) := x"003B";
          m(307) := x"006E";
          m(308) := x"0003";
          m(309) := x"0053";
          m(310) := x"FFF7";
          m(311) := x"FEAB";
          m(312) := x"0127";
          m(313) := x"0161";
          m(314) := x"0080";
          m(315) := x"FB70";
          m(316) := x"FF85";
          m(317) := x"0027";
          m(318) := x"FFBF";
          m(319) := x"FD9F";
          m(320) := x"009E";
          m(321) := x"FF26";
          m(322) := x"FF4E";
          m(323) := x"FCB4";
          m(324) := x"006F";
          m(325) := x"FCA9";
          m(326) := x"FAAF";
          m(327) := x"F8E8";
          m(328) := x"F436";
          m(329) := x"F7A7";
          m(330) := x"F3FE";
          m(331) := x"F6FC";
          m(332) := x"FA8F";
          m(333) := x"FEF1";
          m(334) := x"FFEF";
          m(335) := x"FFDF";
          m(336) := x"FFDA";
          m(337) := x"FFD9";
          m(338) := x"0023";
          m(339) := x"FEEF";
          m(340) := x"0270";
          m(341) := x"0144";
          m(342) := x"FFFC";
          m(343) := x"FFAD";
          m(344) := x"067F";
          m(345) := x"0215";
          m(346) := x"0252";
          m(347) := x"0428";
          m(348) := x"0025";
          m(349) := x"039A";
          m(350) := x"00C4";
          m(351) := x"FE0A";
          m(352) := x"014E";
          m(353) := x"FA15";
          m(354) := x"003A";
          m(355) := x"FF2E";
          m(356) := x"FDE3";
          m(357) := x"FCE5";
          m(358) := x"FB27";
          m(359) := x"FA7F";
          m(360) := x"FAE4";
          m(361) := x"FF14";
          m(362) := x"FFCA";
          m(363) := x"FFE0";
          m(364) := x"FFDE";
          m(365) := x"FFF6";
          m(366) := x"FFF8";
          m(367) := x"FFA6";
          m(368) := x"03D3";
          m(369) := x"0529";
          m(370) := x"014F";
          m(371) := x"02CB";
          m(372) := x"FEE6";
          m(373) := x"FC18";
          m(374) := x"FEDD";
          m(375) := x"0294";
          m(376) := x"05F8";
          m(377) := x"03C2";
          m(378) := x"FFD9";
          m(379) := x"FE09";
          m(380) := x"FC6F";
          m(381) := x"FF64";
          m(382) := x"FBCB";
          m(383) := x"FD79";
          m(384) := x"FCBC";
          m(385) := x"FCC4";
          m(386) := x"FDF8";
          m(387) := x"0004";
          m(388) := x"FFDE";
          m(389) := x"FF26";
          m(390) := x"FFD7";
          m(391) := x"FFFD";
          m(392) := x"0015";
          m(393) := x"FFCD";
          m(394) := x"0055";
          m(395) := x"FF9A";
          m(396) := x"0309";
          m(397) := x"009F";
          m(398) := x"01F2";
          m(399) := x"02D0";
          m(400) := x"02B4";
          m(401) := x"FF47";
          m(402) := x"011A";
          m(403) := x"FF10";
          m(404) := x"03D9";
          m(405) := x"FD92";
          m(406) := x"FFBC";
          m(407) := x"FEB8";
          m(408) := x"FA25";
          m(409) := x"FC2E";
          m(410) := x"0196";
          m(411) := x"FE02";
          m(412) := x"024D";
          m(413) := x"FA2A";
          m(414) := x"FF3F";
          m(415) := x"0368";
          m(416) := x"02E0";
          m(417) := x"FFA9";
          m(418) := x"0010";
          m(419) := x"FF91";
          m(420) := x"FFC6";
          m(421) := x"003A";
          m(422) := x"FF7C";
          m(423) := x"FEEA";
          m(424) := x"FF33";
          m(425) := x"FEBE";
          m(426) := x"FE8F";
          m(427) := x"FE59";
          m(428) := x"0168";
          m(429) := x"02AA";
          m(430) := x"074C";
          m(431) := x"FCDD";
          m(432) := x"0263";
          m(433) := x"FF26";
          m(434) := x"FB1B";
          m(435) := x"FD0C";
          m(436) := x"FDE1";
          m(437) := x"FFEB";
          m(438) := x"0110";
          m(439) := x"012F";
          m(440) := x"0260";
          m(441) := x"FEEB";
          m(442) := x"FB6B";
          m(443) := x"0286";
          m(444) := x"0491";
          m(445) := x"0004";
          m(446) := x"003D";
          m(447) := x"001D";
          m(448) := x"001B";
          m(449) := x"FFEF";
          m(450) := x"FFBC";
          m(451) := x"FF2B";
          m(452) := x"FEA3";
          m(453) := x"FCD7";
          m(454) := x"F8EF";
          m(455) := x"F958";
          m(456) := x"FC68";
          m(457) := x"FB5D";
          m(458) := x"00CA";
          m(459) := x"FDA1";
          m(460) := x"03F4";
          m(461) := x"02D1";
          m(462) := x"0345";
          m(463) := x"01F3";
          m(464) := x"0021";
          m(465) := x"FEE1";
          m(466) := x"FEF0";
          m(467) := x"00C9";
          m(468) := x"0363";
          m(469) := x"00EA";
          m(470) := x"04D3";
          m(471) := x"04ED";
          m(472) := x"039D";
          m(473) := x"FFDE";
          m(474) := x"004F";
          m(475) := x"0041";
          m(476) := x"0016";
          m(477) := x"0023";
          m(478) := x"FF9B";
          m(479) := x"00D7";
          m(480) := x"00FC";
          m(481) := x"FC48";
          m(482) := x"FB7E";
          m(483) := x"F95D";
          m(484) := x"FB84";
          m(485) := x"F9B6";
          m(486) := x"FE3D";
          m(487) := x"FC8F";
          m(488) := x"FBF6";
          m(489) := x"FEDD";
          m(490) := x"FD85";
          m(491) := x"FBB1";
          m(492) := x"F786";
          m(493) := x"FD2E";
          m(494) := x"02D3";
          m(495) := x"FE9B";
          m(496) := x"FF35";
          m(497) := x"0112";
          m(498) := x"0152";
          m(499) := x"037D";
          m(500) := x"01F1";
          m(501) := x"0041";
          m(502) := x"FFEB";
          m(503) := x"FFE9";
          m(504) := x"0003";
          m(505) := x"002C";
          m(506) := x"FF98";
          m(507) := x"003D";
          m(508) := x"0525";
          m(509) := x"00D2";
          m(510) := x"FC7B";
          m(511) := x"FF0C";
          m(512) := x"F911";
          m(513) := x"FBD2";
          m(514) := x"FA83";
          m(515) := x"F421";
          m(516) := x"F546";
          m(517) := x"F44E";
          m(518) := x"F52D";
          m(519) := x"FB7E";
          m(520) := x"00D5";
          m(521) := x"FE23";
          m(522) := x"FDC5";
          m(523) := x"0286";
          m(524) := x"011C";
          m(525) := x"026C";
          m(526) := x"FD14";
          m(527) := x"0197";
          m(528) := x"02B2";
          m(529) := x"006B";
          m(530) := x"FFB7";
          m(531) := x"0005";
          m(532) := x"0007";
          m(533) := x"FFEC";
          m(534) := x"00E1";
          m(535) := x"0021";
          m(536) := x"0585";
          m(537) := x"039F";
          m(538) := x"FD51";
          m(539) := x"FBB0";
          m(540) := x"FE38";
          m(541) := x"F94A";
          m(542) := x"FAE2";
          m(543) := x"015C";
          m(544) := x"FF44";
          m(545) := x"F83D";
          m(546) := x"FF7A";
          m(547) := x"FB67";
          m(548) := x"016C";
          m(549) := x"0116";
          m(550) := x"0056";
          m(551) := x"FFBA";
          m(552) := x"04E4";
          m(553) := x"017A";
          m(554) := x"FDE5";
          m(555) := x"0020";
          m(556) := x"052B";
          m(557) := x"0138";
          m(558) := x"FFDE";
          m(559) := x"FFF4";
          m(560) := x"0000";
          m(561) := x"FFEC";
          m(562) := x"0075";
          m(563) := x"00A0";
          m(564) := x"051A";
          m(565) := x"0740";
          m(566) := x"FEB0";
          m(567) := x"F6E4";
          m(568) := x"FF71";
          m(569) := x"0372";
          m(570) := x"FF17";
          m(571) := x"011C";
          m(572) := x"01C2";
          m(573) := x"0414";
          m(574) := x"FE7D";
          m(575) := x"00E9";
          m(576) := x"0028";
          m(577) := x"03E3";
          m(578) := x"FFBE";
          m(579) := x"FED9";
          m(580) := x"0296";
          m(581) := x"01FF";
          m(582) := x"0126";
          m(583) := x"05D8";
          m(584) := x"03F1";
          m(585) := x"012C";
          m(586) := x"FFDC";
          m(587) := x"0000";
          m(588) := x"000D";
          m(589) := x"FFA6";
          m(590) := x"FF20";
          m(591) := x"FF66";
          m(592) := x"049A";
          m(593) := x"084A";
          m(594) := x"0015";
          m(595) := x"008D";
          m(596) := x"0183";
          m(597) := x"FF4A";
          m(598) := x"045B";
          m(599) := x"01A5";
          m(600) := x"0299";
          m(601) := x"0127";
          m(602) := x"04FF";
          m(603) := x"03DA";
          m(604) := x"00A8";
          m(605) := x"0477";
          m(606) := x"0336";
          m(607) := x"01A8";
          m(608) := x"06D9";
          m(609) := x"0400";
          m(610) := x"FF3B";
          m(611) := x"0682";
          m(612) := x"0304";
          m(613) := x"011F";
          m(614) := x"FFD7";
          m(615) := x"FFF6";
          m(616) := x"FFF4";
          m(617) := x"FFCB";
          m(618) := x"FFD8";
          m(619) := x"004D";
          m(620) := x"02F9";
          m(621) := x"022A";
          m(622) := x"FFE0";
          m(623) := x"FD88";
          m(624) := x"02D8";
          m(625) := x"02B9";
          m(626) := x"FEFC";
          m(627) := x"0074";
          m(628) := x"FEA0";
          m(629) := x"F93B";
          m(630) := x"0397";
          m(631) := x"FF3D";
          m(632) := x"FF86";
          m(633) := x"005F";
          m(634) := x"0216";
          m(635) := x"0189";
          m(636) := x"00E5";
          m(637) := x"0113";
          m(638) := x"02BD";
          m(639) := x"04B3";
          m(640) := x"0038";
          m(641) := x"00BC";
          m(642) := x"002B";
          m(643) := x"FFAB";
          m(644) := x"FFF8";
          m(645) := x"FFDD";
          m(646) := x"FFFD";
          m(647) := x"0096";
          m(648) := x"01D7";
          m(649) := x"0115";
          m(650) := x"FFAE";
          m(651) := x"FBE7";
          m(652) := x"006D";
          m(653) := x"00B5";
          m(654) := x"FEB9";
          m(655) := x"034E";
          m(656) := x"032D";
          m(657) := x"012C";
          m(658) := x"025F";
          m(659) := x"FEF6";
          m(660) := x"FE1A";
          m(661) := x"FCED";
          m(662) := x"FA47";
          m(663) := x"FDCF";
          m(664) := x"016A";
          m(665) := x"0032";
          m(666) := x"FF89";
          m(667) := x"01BF";
          m(668) := x"0110";
          m(669) := x"00DC";
          m(670) := x"000B";
          m(671) := x"FFFC";
          m(672) := x"FFF9";
          m(673) := x"FFEA";
          m(674) := x"FFEE";
          m(675) := x"FFE9";
          m(676) := x"FF3C";
          m(677) := x"FFD5";
          m(678) := x"FEE0";
          m(679) := x"FFA3";
          m(680) := x"FFB5";
          m(681) := x"021B";
          m(682) := x"018C";
          m(683) := x"0034";
          m(684) := x"0325";
          m(685) := x"0291";
          m(686) := x"020C";
          m(687) := x"00B4";
          m(688) := x"FE9E";
          m(689) := x"0187";
          m(690) := x"058B";
          m(691) := x"0226";
          m(692) := x"0243";
          m(693) := x"0061";
          m(694) := x"012D";
          m(695) := x"0039";
          m(696) := x"FFCD";
          m(697) := x"FFF8";
          m(698) := x"0015";
          m(699) := x"FFE8";
          m(700) := x"FFF3";
          m(701) := x"FFEB";
          m(702) := x"FFF8";
          m(703) := x"FFE2";
          m(704) := x"FF2C";
          m(705) := x"FEBC";
          m(706) := x"FE06";
          m(707) := x"FC40";
          m(708) := x"FD59";
          m(709) := x"FF00";
          m(710) := x"FDEC";
          m(711) := x"FFE8";
          m(712) := x"0233";
          m(713) := x"01B4";
          m(714) := x"0019";
          m(715) := x"0164";
          m(716) := x"0013";
          m(717) := x"020D";
          m(718) := x"03B9";
          m(719) := x"0459";
          m(720) := x"0222";
          m(721) := x"01F3";
          m(722) := x"021D";
          m(723) := x"00C2";
          m(724) := x"0088";
          m(725) := x"0007";
          m(726) := x"001B";
          m(727) := x"FFDF";
          m(728) := x"FFED";
          m(729) := x"FFAB";
          m(730) := x"FFE2";
          m(731) := x"0018";
          m(732) := x"FFF7";
          m(733) := x"FFD1";
          m(734) := x"FFA5";
          m(735) := x"FF94";
          m(736) := x"FF94";
          m(737) := x"FEA6";
          m(738) := x"FF19";
          m(739) := x"0087";
          m(740) := x"0124";
          m(741) := x"015B";
          m(742) := x"016E";
          m(743) := x"0276";
          m(744) := x"025A";
          m(745) := x"FF77";
          m(746) := x"FF78";
          m(747) := x"0065";
          m(748) := x"009B";
          m(749) := x"015D";
          m(750) := x"00A7";
          m(751) := x"003B";
          m(752) := x"001D";
          m(753) := x"FFE8";
          m(754) := x"0036";
          m(755) := x"0019";
          m(756) := x"000B";
          m(757) := x"FFEC";
          m(758) := x"001B";
          m(759) := x"0004";
          m(760) := x"FFFF";
          m(761) := x"FFFB";
          m(762) := x"FFFE";
          m(763) := x"0029";
          m(764) := x"FFB8";
          m(765) := x"FFE6";
          m(766) := x"FFF1";
          m(767) := x"0039";
          m(768) := x"FFC9";
          m(769) := x"FFEF";
          m(770) := x"0000";
          m(771) := x"003C";
          m(772) := x"0028";
          m(773) := x"0018";
          m(774) := x"FFDF";
          m(775) := x"0001";
          m(776) := x"FFDE";
          m(777) := x"00A9";
          m(778) := x"003F";
          m(779) := x"FFDB";
          m(780) := x"000B";
          m(781) := x"FFF4";
          m(782) := x"FFEF";
          m(783) := x"FFF5";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_24.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 24) then
          m(0) := x"0057";
          m(1) := x"FFD2";
          m(2) := x"0012";
          m(3) := x"0035";
          m(4) := x"0027";
          m(5) := x"FFDE";
          m(6) := x"FFF9";
          m(7) := x"FFFA";
          m(8) := x"002E";
          m(9) := x"0016";
          m(10) := x"FFD4";
          m(11) := x"000F";
          m(12) := x"001D";
          m(13) := x"FFF9";
          m(14) := x"FFDF";
          m(15) := x"FFF0";
          m(16) := x"FFFB";
          m(17) := x"005A";
          m(18) := x"001F";
          m(19) := x"0022";
          m(20) := x"000E";
          m(21) := x"FFFD";
          m(22) := x"FFFE";
          m(23) := x"FFEA";
          m(24) := x"0015";
          m(25) := x"0022";
          m(26) := x"FFE4";
          m(27) := x"004A";
          m(28) := x"0010";
          m(29) := x"0002";
          m(30) := x"FFD5";
          m(31) := x"001C";
          m(32) := x"FFE8";
          m(33) := x"FFC3";
          m(34) := x"FFF0";
          m(35) := x"FFF6";
          m(36) := x"FFF2";
          m(37) := x"0014";
          m(38) := x"000B";
          m(39) := x"000A";
          m(40) := x"0008";
          m(41) := x"FFE2";
          m(42) := x"000D";
          m(43) := x"0075";
          m(44) := x"003A";
          m(45) := x"0023";
          m(46) := x"FFC7";
          m(47) := x"FFEA";
          m(48) := x"FFD1";
          m(49) := x"002A";
          m(50) := x"FFEF";
          m(51) := x"0000";
          m(52) := x"003E";
          m(53) := x"FFEF";
          m(54) := x"FFFA";
          m(55) := x"FFFA";
          m(56) := x"0003";
          m(57) := x"FFDB";
          m(58) := x"0009";
          m(59) := x"001A";
          m(60) := x"FFF1";
          m(61) := x"0002";
          m(62) := x"FFBF";
          m(63) := x"FF91";
          m(64) := x"FF5E";
          m(65) := x"FEBC";
          m(66) := x"FE9C";
          m(67) := x"FDF3";
          m(68) := x"FE1C";
          m(69) := x"008F";
          m(70) := x"FE2E";
          m(71) := x"FFB9";
          m(72) := x"004F";
          m(73) := x"FF79";
          m(74) := x"FFB6";
          m(75) := x"FFCF";
          m(76) := x"FF3E";
          m(77) := x"FF49";
          m(78) := x"FFD7";
          m(79) := x"0013";
          m(80) := x"0016";
          m(81) := x"001F";
          m(82) := x"0033";
          m(83) := x"0001";
          m(84) := x"0001";
          m(85) := x"0024";
          m(86) := x"FFEB";
          m(87) := x"FFEA";
          m(88) := x"FFE3";
          m(89) := x"0033";
          m(90) := x"0073";
          m(91) := x"019D";
          m(92) := x"02BF";
          m(93) := x"FF4E";
          m(94) := x"002B";
          m(95) := x"FD2D";
          m(96) := x"FFF5";
          m(97) := x"038B";
          m(98) := x"01A6";
          m(99) := x"0217";
          m(100) := x"0180";
          m(101) := x"FE60";
          m(102) := x"FF04";
          m(103) := x"00D8";
          m(104) := x"039F";
          m(105) := x"01CA";
          m(106) := x"FFC5";
          m(107) := x"FFC6";
          m(108) := x"0058";
          m(109) := x"00A2";
          m(110) := x"0026";
          m(111) := x"0009";
          m(112) := x"0003";
          m(113) := x"003B";
          m(114) := x"FFC1";
          m(115) := x"0013";
          m(116) := x"FFFF";
          m(117) := x"00B7";
          m(118) := x"0079";
          m(119) := x"0225";
          m(120) := x"04BF";
          m(121) := x"0336";
          m(122) := x"0237";
          m(123) := x"FF1A";
          m(124) := x"FEC3";
          m(125) := x"FDD8";
          m(126) := x"FFE7";
          m(127) := x"02DF";
          m(128) := x"00B2";
          m(129) := x"FDF8";
          m(130) := x"029E";
          m(131) := x"0002";
          m(132) := x"0394";
          m(133) := x"06D6";
          m(134) := x"02B6";
          m(135) := x"0113";
          m(136) := x"0413";
          m(137) := x"01E7";
          m(138) := x"0025";
          m(139) := x"FFED";
          m(140) := x"0007";
          m(141) := x"FFF6";
          m(142) := x"FFD9";
          m(143) := x"00D8";
          m(144) := x"0067";
          m(145) := x"0274";
          m(146) := x"0188";
          m(147) := x"0364";
          m(148) := x"00E6";
          m(149) := x"FEE7";
          m(150) := x"016D";
          m(151) := x"0113";
          m(152) := x"FD69";
          m(153) := x"0350";
          m(154) := x"0295";
          m(155) := x"0398";
          m(156) := x"0282";
          m(157) := x"01B4";
          m(158) := x"02F7";
          m(159) := x"0090";
          m(160) := x"00CA";
          m(161) := x"007D";
          m(162) := x"0192";
          m(163) := x"0295";
          m(164) := x"0405";
          m(165) := x"01D1";
          m(166) := x"0060";
          m(167) := x"002C";
          m(168) := x"0020";
          m(169) := x"FFF8";
          m(170) := x"0001";
          m(171) := x"0143";
          m(172) := x"01D8";
          m(173) := x"0447";
          m(174) := x"04C0";
          m(175) := x"016C";
          m(176) := x"0110";
          m(177) := x"023E";
          m(178) := x"FC40";
          m(179) := x"FC46";
          m(180) := x"00A6";
          m(181) := x"016F";
          m(182) := x"FF81";
          m(183) := x"FDD4";
          m(184) := x"FBF2";
          m(185) := x"002C";
          m(186) := x"01F0";
          m(187) := x"FC34";
          m(188) := x"FEF2";
          m(189) := x"FF6D";
          m(190) := x"0133";
          m(191) := x"0360";
          m(192) := x"0480";
          m(193) := x"01A2";
          m(194) := x"006A";
          m(195) := x"FFFA";
          m(196) := x"FFD9";
          m(197) := x"0005";
          m(198) := x"004A";
          m(199) := x"0174";
          m(200) := x"028D";
          m(201) := x"02B6";
          m(202) := x"02A6";
          m(203) := x"03E8";
          m(204) := x"0227";
          m(205) := x"012C";
          m(206) := x"01FF";
          m(207) := x"FA75";
          m(208) := x"FBDE";
          m(209) := x"FC86";
          m(210) := x"01C4";
          m(211) := x"0583";
          m(212) := x"FDC7";
          m(213) := x"0195";
          m(214) := x"FD31";
          m(215) := x"0147";
          m(216) := x"FF39";
          m(217) := x"FB14";
          m(218) := x"0088";
          m(219) := x"0136";
          m(220) := x"0122";
          m(221) := x"FFF8";
          m(222) := x"00C5";
          m(223) := x"000F";
          m(224) := x"0022";
          m(225) := x"000B";
          m(226) := x"FFA8";
          m(227) := x"00C7";
          m(228) := x"01A6";
          m(229) := x"033D";
          m(230) := x"01A4";
          m(231) := x"00FB";
          m(232) := x"0141";
          m(233) := x"FE65";
          m(234) := x"028B";
          m(235) := x"01B8";
          m(236) := x"FEE7";
          m(237) := x"FFF7";
          m(238) := x"029F";
          m(239) := x"FF98";
          m(240) := x"F94B";
          m(241) := x"FA3A";
          m(242) := x"00ED";
          m(243) := x"00C2";
          m(244) := x"0210";
          m(245) := x"02AF";
          m(246) := x"022D";
          m(247) := x"0020";
          m(248) := x"020B";
          m(249) := x"020F";
          m(250) := x"009B";
          m(251) := x"0034";
          m(252) := x"FFD2";
          m(253) := x"0008";
          m(254) := x"FF6A";
          m(255) := x"FFCD";
          m(256) := x"FF86";
          m(257) := x"FE9F";
          m(258) := x"FFE1";
          m(259) := x"0123";
          m(260) := x"FFA0";
          m(261) := x"FD6C";
          m(262) := x"FFAD";
          m(263) := x"0133";
          m(264) := x"0168";
          m(265) := x"0466";
          m(266) := x"0977";
          m(267) := x"02F8";
          m(268) := x"FE01";
          m(269) := x"FCAE";
          m(270) := x"FCB6";
          m(271) := x"FBF6";
          m(272) := x"FE02";
          m(273) := x"FD3F";
          m(274) := x"03CB";
          m(275) := x"FD27";
          m(276) := x"FFB6";
          m(277) := x"025A";
          m(278) := x"009F";
          m(279) := x"0019";
          m(280) := x"FFFB";
          m(281) := x"001C";
          m(282) := x"FF9B";
          m(283) := x"FFDC";
          m(284) := x"FD35";
          m(285) := x"FC3C";
          m(286) := x"FB60";
          m(287) := x"FCDA";
          m(288) := x"030A";
          m(289) := x"FFE6";
          m(290) := x"002F";
          m(291) := x"FE44";
          m(292) := x"FFCB";
          m(293) := x"0914";
          m(294) := x"0B13";
          m(295) := x"04CE";
          m(296) := x"05CB";
          m(297) := x"0285";
          m(298) := x"F894";
          m(299) := x"FDDB";
          m(300) := x"01A1";
          m(301) := x"FC48";
          m(302) := x"0114";
          m(303) := x"FF92";
          m(304) := x"FFA7";
          m(305) := x"0205";
          m(306) := x"00A5";
          m(307) := x"001C";
          m(308) := x"0000";
          m(309) := x"FFAE";
          m(310) := x"0045";
          m(311) := x"008E";
          m(312) := x"0006";
          m(313) := x"FE3D";
          m(314) := x"FBD0";
          m(315) := x"F8A1";
          m(316) := x"002C";
          m(317) := x"FA39";
          m(318) := x"FE02";
          m(319) := x"FF85";
          m(320) := x"FAB8";
          m(321) := x"FEDE";
          m(322) := x"046E";
          m(323) := x"05BB";
          m(324) := x"0937";
          m(325) := x"0D5E";
          m(326) := x"005F";
          m(327) := x"FFE1";
          m(328) := x"01F9";
          m(329) := x"FC42";
          m(330) := x"FE91";
          m(331) := x"FDFC";
          m(332) := x"FFC2";
          m(333) := x"0070";
          m(334) := x"0097";
          m(335) := x"FFF6";
          m(336) := x"FFDD";
          m(337) := x"0020";
          m(338) := x"FFB0";
          m(339) := x"FFF4";
          m(340) := x"FFC4";
          m(341) := x"FC93";
          m(342) := x"F9FB";
          m(343) := x"FAC7";
          m(344) := x"FD12";
          m(345) := x"FE2D";
          m(346) := x"0073";
          m(347) := x"0245";
          m(348) := x"00B7";
          m(349) := x"FC1C";
          m(350) := x"0491";
          m(351) := x"04E0";
          m(352) := x"0742";
          m(353) := x"06D2";
          m(354) := x"0514";
          m(355) := x"FD8A";
          m(356) := x"02DF";
          m(357) := x"FC04";
          m(358) := x"FE64";
          m(359) := x"FCDA";
          m(360) := x"F9F5";
          m(361) := x"FE39";
          m(362) := x"FFEF";
          m(363) := x"FFDB";
          m(364) := x"FFF3";
          m(365) := x"FFD1";
          m(366) := x"FFF5";
          m(367) := x"00A8";
          m(368) := x"FF8F";
          m(369) := x"F9A4";
          m(370) := x"F873";
          m(371) := x"F981";
          m(372) := x"FF5D";
          m(373) := x"FDF3";
          m(374) := x"FF16";
          m(375) := x"002B";
          m(376) := x"00B0";
          m(377) := x"FDA8";
          m(378) := x"0478";
          m(379) := x"02BA";
          m(380) := x"08EC";
          m(381) := x"082F";
          m(382) := x"003F";
          m(383) := x"0513";
          m(384) := x"00C2";
          m(385) := x"00E2";
          m(386) := x"FCB7";
          m(387) := x"FB2B";
          m(388) := x"FBFE";
          m(389) := x"FE2B";
          m(390) := x"FF46";
          m(391) := x"FF3E";
          m(392) := x"FFD8";
          m(393) := x"0066";
          m(394) := x"FFFA";
          m(395) := x"0021";
          m(396) := x"FE91";
          m(397) := x"F7D5";
          m(398) := x"F4C7";
          m(399) := x"F4FC";
          m(400) := x"F9C1";
          m(401) := x"FF69";
          m(402) := x"FE63";
          m(403) := x"FC12";
          m(404) := x"007F";
          m(405) := x"023E";
          m(406) := x"088A";
          m(407) := x"0254";
          m(408) := x"03D7";
          m(409) := x"033E";
          m(410) := x"FE69";
          m(411) := x"FED1";
          m(412) := x"FE59";
          m(413) := x"004A";
          m(414) := x"FFBD";
          m(415) := x"FE6F";
          m(416) := x"FE54";
          m(417) := x"FEE7";
          m(418) := x"FFAC";
          m(419) := x"0025";
          m(420) := x"FFEE";
          m(421) := x"003F";
          m(422) := x"0064";
          m(423) := x"FFCA";
          m(424) := x"FF1A";
          m(425) := x"F82A";
          m(426) := x"F517";
          m(427) := x"F473";
          m(428) := x"F380";
          m(429) := x"F599";
          m(430) := x"F542";
          m(431) := x"F806";
          m(432) := x"01F2";
          m(433) := x"00C0";
          m(434) := x"045A";
          m(435) := x"0755";
          m(436) := x"052D";
          m(437) := x"FFBE";
          m(438) := x"03FC";
          m(439) := x"0045";
          m(440) := x"016A";
          m(441) := x"037E";
          m(442) := x"0210";
          m(443) := x"051E";
          m(444) := x"0170";
          m(445) := x"FF0A";
          m(446) := x"FF95";
          m(447) := x"000D";
          m(448) := x"FFC1";
          m(449) := x"000B";
          m(450) := x"005F";
          m(451) := x"00C3";
          m(452) := x"0210";
          m(453) := x"FCD0";
          m(454) := x"FD35";
          m(455) := x"FC0A";
          m(456) := x"F9C4";
          m(457) := x"F836";
          m(458) := x"F2FA";
          m(459) := x"F0E9";
          m(460) := x"F86A";
          m(461) := x"F983";
          m(462) := x"FF7A";
          m(463) := x"028C";
          m(464) := x"FB8B";
          m(465) := x"0041";
          m(466) := x"04E0";
          m(467) := x"02FE";
          m(468) := x"0290";
          m(469) := x"0227";
          m(470) := x"03F7";
          m(471) := x"04A9";
          m(472) := x"FF32";
          m(473) := x"FD00";
          m(474) := x"FF25";
          m(475) := x"FFF8";
          m(476) := x"0007";
          m(477) := x"FFE8";
          m(478) := x"0052";
          m(479) := x"02D0";
          m(480) := x"00D9";
          m(481) := x"015A";
          m(482) := x"01E6";
          m(483) := x"0321";
          m(484) := x"F9EF";
          m(485) := x"F732";
          m(486) := x"F53F";
          m(487) := x"F241";
          m(488) := x"F323";
          m(489) := x"FA07";
          m(490) := x"FB9E";
          m(491) := x"FD4C";
          m(492) := x"FC9C";
          m(493) := x"FF66";
          m(494) := x"0070";
          m(495) := x"0306";
          m(496) := x"FE11";
          m(497) := x"0169";
          m(498) := x"005D";
          m(499) := x"0448";
          m(500) := x"FBA6";
          m(501) := x"FBF2";
          m(502) := x"FF9D";
          m(503) := x"0011";
          m(504) := x"0038";
          m(505) := x"0015";
          m(506) := x"006B";
          m(507) := x"0505";
          m(508) := x"015C";
          m(509) := x"00E3";
          m(510) := x"03AB";
          m(511) := x"015D";
          m(512) := x"01FC";
          m(513) := x"04FB";
          m(514) := x"FA7A";
          m(515) := x"F6EE";
          m(516) := x"F331";
          m(517) := x"FA25";
          m(518) := x"014B";
          m(519) := x"07A0";
          m(520) := x"FFAD";
          m(521) := x"0035";
          m(522) := x"FBA5";
          m(523) := x"FFB8";
          m(524) := x"023A";
          m(525) := x"FD72";
          m(526) := x"FFAB";
          m(527) := x"FF9A";
          m(528) := x"FBB0";
          m(529) := x"FDEC";
          m(530) := x"002E";
          m(531) := x"000D";
          m(532) := x"FFF4";
          m(533) := x"001B";
          m(534) := x"0019";
          m(535) := x"02A5";
          m(536) := x"007D";
          m(537) := x"0276";
          m(538) := x"0304";
          m(539) := x"0084";
          m(540) := x"00DA";
          m(541) := x"FFF9";
          m(542) := x"FD16";
          m(543) := x"F9EA";
          m(544) := x"F981";
          m(545) := x"FC63";
          m(546) := x"04D2";
          m(547) := x"0554";
          m(548) := x"0364";
          m(549) := x"0518";
          m(550) := x"0078";
          m(551) := x"0123";
          m(552) := x"0318";
          m(553) := x"00BF";
          m(554) := x"01ED";
          m(555) := x"FDA3";
          m(556) := x"FF65";
          m(557) := x"FF33";
          m(558) := x"FFDA";
          m(559) := x"FFD2";
          m(560) := x"FFF6";
          m(561) := x"0007";
          m(562) := x"FEF3";
          m(563) := x"FEEC";
          m(564) := x"00B5";
          m(565) := x"0332";
          m(566) := x"0238";
          m(567) := x"FFFF";
          m(568) := x"FEA6";
          m(569) := x"009D";
          m(570) := x"FEBD";
          m(571) := x"FC6A";
          m(572) := x"F655";
          m(573) := x"FC6A";
          m(574) := x"05F7";
          m(575) := x"00A0";
          m(576) := x"FFE6";
          m(577) := x"036C";
          m(578) := x"0223";
          m(579) := x"0109";
          m(580) := x"028F";
          m(581) := x"FD10";
          m(582) := x"FFD6";
          m(583) := x"FEA0";
          m(584) := x"FE88";
          m(585) := x"FF28";
          m(586) := x"0011";
          m(587) := x"FF9C";
          m(588) := x"FFE4";
          m(589) := x"FFC9";
          m(590) := x"FE19";
          m(591) := x"FCD8";
          m(592) := x"FECB";
          m(593) := x"FF33";
          m(594) := x"FF3F";
          m(595) := x"03AF";
          m(596) := x"02E5";
          m(597) := x"0000";
          m(598) := x"0026";
          m(599) := x"FC5B";
          m(600) := x"F8D1";
          m(601) := x"00C0";
          m(602) := x"0627";
          m(603) := x"01D2";
          m(604) := x"FD8E";
          m(605) := x"FE8C";
          m(606) := x"02FB";
          m(607) := x"FE22";
          m(608) := x"01F5";
          m(609) := x"FD14";
          m(610) := x"FBA5";
          m(611) := x"FA1B";
          m(612) := x"FDBB";
          m(613) := x"FF35";
          m(614) := x"FFC4";
          m(615) := x"002A";
          m(616) := x"000A";
          m(617) := x"FFF6";
          m(618) := x"FE46";
          m(619) := x"FE3F";
          m(620) := x"FE36";
          m(621) := x"FC11";
          m(622) := x"FC41";
          m(623) := x"FCA0";
          m(624) := x"FEAC";
          m(625) := x"FCE8";
          m(626) := x"FD78";
          m(627) := x"FBAE";
          m(628) := x"F913";
          m(629) := x"0150";
          m(630) := x"047D";
          m(631) := x"01FA";
          m(632) := x"FE8C";
          m(633) := x"02BB";
          m(634) := x"0334";
          m(635) := x"01B3";
          m(636) := x"FC6D";
          m(637) := x"FC52";
          m(638) := x"FC35";
          m(639) := x"FBAE";
          m(640) := x"FDFE";
          m(641) := x"FF17";
          m(642) := x"0033";
          m(643) := x"0044";
          m(644) := x"0016";
          m(645) := x"FFFA";
          m(646) := x"007B";
          m(647) := x"019F";
          m(648) := x"02A1";
          m(649) := x"004F";
          m(650) := x"FC73";
          m(651) := x"FC76";
          m(652) := x"F8E6";
          m(653) := x"F9C2";
          m(654) := x"FA11";
          m(655) := x"FCB4";
          m(656) := x"F77B";
          m(657) := x"FE84";
          m(658) := x"02B3";
          m(659) := x"026B";
          m(660) := x"FDC8";
          m(661) := x"02F9";
          m(662) := x"03DD";
          m(663) := x"FE6B";
          m(664) := x"FD60";
          m(665) := x"FC6D";
          m(666) := x"FBD5";
          m(667) := x"FC9D";
          m(668) := x"FE8C";
          m(669) := x"FEDF";
          m(670) := x"FFF2";
          m(671) := x"FFFA";
          m(672) := x"0027";
          m(673) := x"FFF4";
          m(674) := x"006A";
          m(675) := x"0130";
          m(676) := x"01EE";
          m(677) := x"018A";
          m(678) := x"01ED";
          m(679) := x"032D";
          m(680) := x"FDD8";
          m(681) := x"FB55";
          m(682) := x"FA6D";
          m(683) := x"FE92";
          m(684) := x"FFD8";
          m(685) := x"02F7";
          m(686) := x"FFF0";
          m(687) := x"FD6B";
          m(688) := x"01F3";
          m(689) := x"06C6";
          m(690) := x"003C";
          m(691) := x"FBDD";
          m(692) := x"FE05";
          m(693) := x"FD1B";
          m(694) := x"FD5C";
          m(695) := x"FEF3";
          m(696) := x"FE9E";
          m(697) := x"FF6F";
          m(698) := x"FFDE";
          m(699) := x"0005";
          m(700) := x"0015";
          m(701) := x"001A";
          m(702) := x"0011";
          m(703) := x"FFE6";
          m(704) := x"001C";
          m(705) := x"00B3";
          m(706) := x"0128";
          m(707) := x"0301";
          m(708) := x"03C8";
          m(709) := x"02CA";
          m(710) := x"025B";
          m(711) := x"023F";
          m(712) := x"0449";
          m(713) := x"038E";
          m(714) := x"003E";
          m(715) := x"FEBE";
          m(716) := x"021E";
          m(717) := x"029A";
          m(718) := x"02CF";
          m(719) := x"03A1";
          m(720) := x"022B";
          m(721) := x"014F";
          m(722) := x"002E";
          m(723) := x"FFB9";
          m(724) := x"0016";
          m(725) := x"0005";
          m(726) := x"000C";
          m(727) := x"0032";
          m(728) := x"FFF3";
          m(729) := x"FFF4";
          m(730) := x"0011";
          m(731) := x"FFA9";
          m(732) := x"FFCA";
          m(733) := x"FFD7";
          m(734) := x"002C";
          m(735) := x"009E";
          m(736) := x"0018";
          m(737) := x"00BB";
          m(738) := x"019A";
          m(739) := x"017C";
          m(740) := x"0063";
          m(741) := x"0109";
          m(742) := x"0192";
          m(743) := x"01CE";
          m(744) := x"048D";
          m(745) := x"03C7";
          m(746) := x"01BA";
          m(747) := x"00B6";
          m(748) := x"00DC";
          m(749) := x"008C";
          m(750) := x"002E";
          m(751) := x"FFFE";
          m(752) := x"FFDB";
          m(753) := x"0014";
          m(754) := x"0012";
          m(755) := x"0000";
          m(756) := x"0023";
          m(757) := x"001C";
          m(758) := x"FFEF";
          m(759) := x"FFE4";
          m(760) := x"FFEB";
          m(761) := x"FFA2";
          m(762) := x"0004";
          m(763) := x"001B";
          m(764) := x"FFD8";
          m(765) := x"FFF8";
          m(766) := x"001C";
          m(767) := x"001D";
          m(768) := x"FFB4";
          m(769) := x"FFAA";
          m(770) := x"FFBB";
          m(771) := x"FFFB";
          m(772) := x"FFC1";
          m(773) := x"FFF8";
          m(774) := x"FFF3";
          m(775) := x"FFDC";
          m(776) := x"FFCA";
          m(777) := x"0025";
          m(778) := x"0032";
          m(779) := x"FFE9";
          m(780) := x"FFE9";
          m(781) := x"0000";
          m(782) := x"FFFD";
          m(783) := x"002D";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_25.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 25) then
          m(0) := x"FFEB";
          m(1) := x"0014";
          m(2) := x"FFB8";
          m(3) := x"FFE8";
          m(4) := x"0006";
          m(5) := x"0005";
          m(6) := x"0031";
          m(7) := x"000A";
          m(8) := x"FFD0";
          m(9) := x"FFF8";
          m(10) := x"000C";
          m(11) := x"0011";
          m(12) := x"000A";
          m(13) := x"0025";
          m(14) := x"0009";
          m(15) := x"FFFB";
          m(16) := x"003C";
          m(17) := x"000C";
          m(18) := x"FFFC";
          m(19) := x"0004";
          m(20) := x"001B";
          m(21) := x"FFF2";
          m(22) := x"FFE2";
          m(23) := x"0000";
          m(24) := x"001C";
          m(25) := x"0008";
          m(26) := x"FFFC";
          m(27) := x"FFED";
          m(28) := x"FFD7";
          m(29) := x"0009";
          m(30) := x"0003";
          m(31) := x"0020";
          m(32) := x"FFE7";
          m(33) := x"0026";
          m(34) := x"0012";
          m(35) := x"FFFE";
          m(36) := x"FFF3";
          m(37) := x"0021";
          m(38) := x"006C";
          m(39) := x"001A";
          m(40) := x"0060";
          m(41) := x"000F";
          m(42) := x"FFF2";
          m(43) := x"0001";
          m(44) := x"0056";
          m(45) := x"001D";
          m(46) := x"FFEB";
          m(47) := x"0045";
          m(48) := x"0037";
          m(49) := x"FFF5";
          m(50) := x"0010";
          m(51) := x"000E";
          m(52) := x"FFE2";
          m(53) := x"0029";
          m(54) := x"FFE3";
          m(55) := x"FFBB";
          m(56) := x"0012";
          m(57) := x"FFF7";
          m(58) := x"FFE6";
          m(59) := x"FFCD";
          m(60) := x"FFFB";
          m(61) := x"FFF9";
          m(62) := x"FFEE";
          m(63) := x"FFFB";
          m(64) := x"0016";
          m(65) := x"FFCF";
          m(66) := x"0021";
          m(67) := x"FFEF";
          m(68) := x"FF8E";
          m(69) := x"FFD4";
          m(70) := x"0024";
          m(71) := x"0040";
          m(72) := x"01D0";
          m(73) := x"01C0";
          m(74) := x"0146";
          m(75) := x"0032";
          m(76) := x"0002";
          m(77) := x"FFF8";
          m(78) := x"000D";
          m(79) := x"004B";
          m(80) := x"FFF3";
          m(81) := x"0009";
          m(82) := x"0002";
          m(83) := x"FFE5";
          m(84) := x"0019";
          m(85) := x"FFEA";
          m(86) := x"0047";
          m(87) := x"0009";
          m(88) := x"000C";
          m(89) := x"FFE8";
          m(90) := x"0010";
          m(91) := x"0034";
          m(92) := x"00E0";
          m(93) := x"0068";
          m(94) := x"01A7";
          m(95) := x"00CD";
          m(96) := x"007E";
          m(97) := x"0158";
          m(98) := x"0090";
          m(99) := x"0403";
          m(100) := x"045E";
          m(101) := x"03C4";
          m(102) := x"033C";
          m(103) := x"00E4";
          m(104) := x"0153";
          m(105) := x"0194";
          m(106) := x"00B0";
          m(107) := x"00B0";
          m(108) := x"009A";
          m(109) := x"FFFF";
          m(110) := x"0012";
          m(111) := x"FFF2";
          m(112) := x"0017";
          m(113) := x"FFDE";
          m(114) := x"FFF0";
          m(115) := x"0029";
          m(116) := x"0009";
          m(117) := x"0097";
          m(118) := x"0048";
          m(119) := x"0053";
          m(120) := x"01BE";
          m(121) := x"0322";
          m(122) := x"0468";
          m(123) := x"00DD";
          m(124) := x"FDEE";
          m(125) := x"FD07";
          m(126) := x"030F";
          m(127) := x"067B";
          m(128) := x"040A";
          m(129) := x"01F0";
          m(130) := x"02AA";
          m(131) := x"FF57";
          m(132) := x"FD13";
          m(133) := x"FFC1";
          m(134) := x"FE73";
          m(135) := x"FE97";
          m(136) := x"FEA4";
          m(137) := x"004D";
          m(138) := x"003D";
          m(139) := x"FFF3";
          m(140) := x"004B";
          m(141) := x"FFEA";
          m(142) := x"0000";
          m(143) := x"0023";
          m(144) := x"FFED";
          m(145) := x"FFDE";
          m(146) := x"FE3A";
          m(147) := x"FEE3";
          m(148) := x"FE2C";
          m(149) := x"FC43";
          m(150) := x"FC85";
          m(151) := x"FB12";
          m(152) := x"FE25";
          m(153) := x"FCB2";
          m(154) := x"FE2D";
          m(155) := x"FD72";
          m(156) := x"0097";
          m(157) := x"0394";
          m(158) := x"0574";
          m(159) := x"019F";
          m(160) := x"FFD8";
          m(161) := x"034F";
          m(162) := x"0255";
          m(163) := x"00D8";
          m(164) := x"0022";
          m(165) := x"0072";
          m(166) := x"0032";
          m(167) := x"0006";
          m(168) := x"002D";
          m(169) := x"0040";
          m(170) := x"FFD4";
          m(171) := x"FFE1";
          m(172) := x"0075";
          m(173) := x"0180";
          m(174) := x"0037";
          m(175) := x"002B";
          m(176) := x"FF54";
          m(177) := x"021F";
          m(178) := x"010C";
          m(179) := x"FE5E";
          m(180) := x"0102";
          m(181) := x"01CE";
          m(182) := x"0420";
          m(183) := x"0460";
          m(184) := x"FFE3";
          m(185) := x"0045";
          m(186) := x"0294";
          m(187) := x"003C";
          m(188) := x"FE20";
          m(189) := x"02C5";
          m(190) := x"027F";
          m(191) := x"009C";
          m(192) := x"0381";
          m(193) := x"01A2";
          m(194) := x"0069";
          m(195) := x"FFE5";
          m(196) := x"FFFE";
          m(197) := x"0017";
          m(198) := x"FED9";
          m(199) := x"FFCB";
          m(200) := x"FE8D";
          m(201) := x"0074";
          m(202) := x"FD3E";
          m(203) := x"FEEF";
          m(204) := x"01DC";
          m(205) := x"0044";
          m(206) := x"04E1";
          m(207) := x"FE89";
          m(208) := x"FD49";
          m(209) := x"027A";
          m(210) := x"0430";
          m(211) := x"03B7";
          m(212) := x"00B7";
          m(213) := x"FE56";
          m(214) := x"FFBE";
          m(215) := x"FCC1";
          m(216) := x"FEE0";
          m(217) := x"FFEB";
          m(218) := x"FFD2";
          m(219) := x"FF5B";
          m(220) := x"0346";
          m(221) := x"01AB";
          m(222) := x"004A";
          m(223) := x"0002";
          m(224) := x"0030";
          m(225) := x"FFC3";
          m(226) := x"FEDF";
          m(227) := x"FEDE";
          m(228) := x"FD2E";
          m(229) := x"FFE8";
          m(230) := x"FE89";
          m(231) := x"046D";
          m(232) := x"01D4";
          m(233) := x"FE01";
          m(234) := x"FEC7";
          m(235) := x"FE01";
          m(236) := x"0304";
          m(237) := x"067B";
          m(238) := x"04D8";
          m(239) := x"01B5";
          m(240) := x"0090";
          m(241) := x"021E";
          m(242) := x"FAF6";
          m(243) := x"FD46";
          m(244) := x"FC81";
          m(245) := x"FD3A";
          m(246) := x"04D6";
          m(247) := x"01AD";
          m(248) := x"0238";
          m(249) := x"0269";
          m(250) := x"013D";
          m(251) := x"000A";
          m(252) := x"0007";
          m(253) := x"FFED";
          m(254) := x"FF79";
          m(255) := x"FEFD";
          m(256) := x"FEA3";
          m(257) := x"FCF7";
          m(258) := x"FF00";
          m(259) := x"05B5";
          m(260) := x"0199";
          m(261) := x"FB4A";
          m(262) := x"FFFE";
          m(263) := x"FFCC";
          m(264) := x"0242";
          m(265) := x"010C";
          m(266) := x"0669";
          m(267) := x"05DE";
          m(268) := x"FF68";
          m(269) := x"FE79";
          m(270) := x"FAB6";
          m(271) := x"FA5D";
          m(272) := x"FBA5";
          m(273) := x"FC5A";
          m(274) := x"0281";
          m(275) := x"00F2";
          m(276) := x"012D";
          m(277) := x"0331";
          m(278) := x"0199";
          m(279) := x"0015";
          m(280) := x"0009";
          m(281) := x"0003";
          m(282) := x"FF9D";
          m(283) := x"FEA4";
          m(284) := x"FEE8";
          m(285) := x"FDBB";
          m(286) := x"0200";
          m(287) := x"0121";
          m(288) := x"FF8C";
          m(289) := x"FCAB";
          m(290) := x"02C0";
          m(291) := x"FB6D";
          m(292) := x"00F6";
          m(293) := x"0824";
          m(294) := x"0C35";
          m(295) := x"0CE2";
          m(296) := x"FEA0";
          m(297) := x"F79A";
          m(298) := x"FE7A";
          m(299) := x"FC93";
          m(300) := x"FEC8";
          m(301) := x"FEB1";
          m(302) := x"019A";
          m(303) := x"FE71";
          m(304) := x"01E5";
          m(305) := x"0139";
          m(306) := x"01EB";
          m(307) := x"FFDD";
          m(308) := x"0027";
          m(309) := x"0032";
          m(310) := x"FF7B";
          m(311) := x"FDE2";
          m(312) := x"FFA5";
          m(313) := x"FE78";
          m(314) := x"FC10";
          m(315) := x"FC5F";
          m(316) := x"031C";
          m(317) := x"FF3D";
          m(318) := x"FA1D";
          m(319) := x"FEC1";
          m(320) := x"FEA2";
          m(321) := x"FF34";
          m(322) := x"0FC8";
          m(323) := x"08D9";
          m(324) := x"FBCA";
          m(325) := x"F793";
          m(326) := x"0045";
          m(327) := x"FC15";
          m(328) := x"FA82";
          m(329) := x"FDD6";
          m(330) := x"FCDC";
          m(331) := x"FDED";
          m(332) := x"01C4";
          m(333) := x"0251";
          m(334) := x"01BB";
          m(335) := x"000F";
          m(336) := x"FFFE";
          m(337) := x"0000";
          m(338) := x"FF87";
          m(339) := x"FE60";
          m(340) := x"FDA6";
          m(341) := x"FCB3";
          m(342) := x"FE3A";
          m(343) := x"FFCD";
          m(344) := x"0016";
          m(345) := x"00F2";
          m(346) := x"FD00";
          m(347) := x"FF5B";
          m(348) := x"FAEE";
          m(349) := x"071C";
          m(350) := x"1622";
          m(351) := x"05DF";
          m(352) := x"F95F";
          m(353) := x"F873";
          m(354) := x"FB2C";
          m(355) := x"F9DE";
          m(356) := x"FA10";
          m(357) := x"FD71";
          m(358) := x"F9DC";
          m(359) := x"FC24";
          m(360) := x"FEF4";
          m(361) := x"02C8";
          m(362) := x"0044";
          m(363) := x"FFBD";
          m(364) := x"FFC4";
          m(365) := x"FFBF";
          m(366) := x"FFA1";
          m(367) := x"FE56";
          m(368) := x"F926";
          m(369) := x"FF25";
          m(370) := x"0089";
          m(371) := x"FCE1";
          m(372) := x"00CB";
          m(373) := x"FA80";
          m(374) := x"FB7E";
          m(375) := x"01E4";
          m(376) := x"03EB";
          m(377) := x"100E";
          m(378) := x"0F00";
          m(379) := x"03FB";
          m(380) := x"F92A";
          m(381) := x"F728";
          m(382) := x"02C1";
          m(383) := x"FB25";
          m(384) := x"FF97";
          m(385) := x"FB60";
          m(386) := x"F8C2";
          m(387) := x"00FC";
          m(388) := x"0142";
          m(389) := x"021C";
          m(390) := x"007A";
          m(391) := x"002B";
          m(392) := x"FFD7";
          m(393) := x"003A";
          m(394) := x"0053";
          m(395) := x"FE7A";
          m(396) := x"FBE9";
          m(397) := x"FCA6";
          m(398) := x"0069";
          m(399) := x"FC4B";
          m(400) := x"F947";
          m(401) := x"FB93";
          m(402) := x"0046";
          m(403) := x"033F";
          m(404) := x"056B";
          m(405) := x"0836";
          m(406) := x"0668";
          m(407) := x"012A";
          m(408) := x"F5FA";
          m(409) := x"FC02";
          m(410) := x"FBFF";
          m(411) := x"F70B";
          m(412) := x"FAE1";
          m(413) := x"FBA1";
          m(414) := x"F926";
          m(415) := x"0032";
          m(416) := x"0333";
          m(417) := x"0176";
          m(418) := x"FFE3";
          m(419) := x"FFC4";
          m(420) := x"FFE5";
          m(421) := x"00D2";
          m(422) := x"0041";
          m(423) := x"FEF5";
          m(424) := x"FCE6";
          m(425) := x"FF0E";
          m(426) := x"01BB";
          m(427) := x"FEC9";
          m(428) := x"FD80";
          m(429) := x"F991";
          m(430) := x"FD84";
          m(431) := x"07FE";
          m(432) := x"056F";
          m(433) := x"05CA";
          m(434) := x"082A";
          m(435) := x"03C7";
          m(436) := x"FCF7";
          m(437) := x"FD1F";
          m(438) := x"F9B2";
          m(439) := x"F70F";
          m(440) := x"FA7B";
          m(441) := x"FCF6";
          m(442) := x"F9BD";
          m(443) := x"0415";
          m(444) := x"0659";
          m(445) := x"021E";
          m(446) := x"FFB4";
          m(447) := x"0014";
          m(448) := x"FFF0";
          m(449) := x"0056";
          m(450) := x"00BE";
          m(451) := x"0150";
          m(452) := x"FD7D";
          m(453) := x"FC7C";
          m(454) := x"FFE6";
          m(455) := x"FF4F";
          m(456) := x"FFB5";
          m(457) := x"0167";
          m(458) := x"FEFE";
          m(459) := x"03CB";
          m(460) := x"0733";
          m(461) := x"0940";
          m(462) := x"0915";
          m(463) := x"FCDF";
          m(464) := x"F9C8";
          m(465) := x"FA57";
          m(466) := x"FCBC";
          m(467) := x"FEB8";
          m(468) := x"FADE";
          m(469) := x"FE9B";
          m(470) := x"0061";
          m(471) := x"05F6";
          m(472) := x"0547";
          m(473) := x"0144";
          m(474) := x"0034";
          m(475) := x"0017";
          m(476) := x"0000";
          m(477) := x"0012";
          m(478) := x"000C";
          m(479) := x"0372";
          m(480) := x"FF21";
          m(481) := x"FD94";
          m(482) := x"FE58";
          m(483) := x"FE5F";
          m(484) := x"FBF7";
          m(485) := x"FF78";
          m(486) := x"FFED";
          m(487) := x"074B";
          m(488) := x"07B5";
          m(489) := x"08CF";
          m(490) := x"03F0";
          m(491) := x"F620";
          m(492) := x"F531";
          m(493) := x"0110";
          m(494) := x"FBF5";
          m(495) := x"00AB";
          m(496) := x"003F";
          m(497) := x"FE32";
          m(498) := x"FE44";
          m(499) := x"0345";
          m(500) := x"003C";
          m(501) := x"0078";
          m(502) := x"FFD5";
          m(503) := x"001D";
          m(504) := x"FFD6";
          m(505) := x"0039";
          m(506) := x"FF9F";
          m(507) := x"03C1";
          m(508) := x"01E3";
          m(509) := x"FEFF";
          m(510) := x"00A7";
          m(511) := x"FF2A";
          m(512) := x"FDFE";
          m(513) := x"0186";
          m(514) := x"FFBC";
          m(515) := x"0471";
          m(516) := x"0354";
          m(517) := x"02E7";
          m(518) := x"FE7A";
          m(519) := x"FB35";
          m(520) := x"F8BE";
          m(521) := x"FD8C";
          m(522) := x"FAEA";
          m(523) := x"FC23";
          m(524) := x"FF9C";
          m(525) := x"FE0C";
          m(526) := x"FF12";
          m(527) := x"01E0";
          m(528) := x"FF94";
          m(529) := x"00C1";
          m(530) := x"FFFF";
          m(531) := x"FFD5";
          m(532) := x"FFEE";
          m(533) := x"FFDC";
          m(534) := x"FFB0";
          m(535) := x"03C0";
          m(536) := x"033C";
          m(537) := x"03A0";
          m(538) := x"0227";
          m(539) := x"00F9";
          m(540) := x"01B1";
          m(541) := x"FE11";
          m(542) := x"FD7E";
          m(543) := x"0321";
          m(544) := x"073A";
          m(545) := x"06C6";
          m(546) := x"FF43";
          m(547) := x"FD17";
          m(548) := x"FE54";
          m(549) := x"FD44";
          m(550) := x"0165";
          m(551) := x"F9BE";
          m(552) := x"035A";
          m(553) := x"FF8E";
          m(554) := x"0013";
          m(555) := x"0008";
          m(556) := x"FEDE";
          m(557) := x"001D";
          m(558) := x"0019";
          m(559) := x"0022";
          m(560) := x"0010";
          m(561) := x"0015";
          m(562) := x"FFE1";
          m(563) := x"0241";
          m(564) := x"048F";
          m(565) := x"00D4";
          m(566) := x"060C";
          m(567) := x"05AC";
          m(568) := x"05E9";
          m(569) := x"0151";
          m(570) := x"FEDA";
          m(571) := x"FF61";
          m(572) := x"02A0";
          m(573) := x"014D";
          m(574) := x"03BD";
          m(575) := x"0580";
          m(576) := x"FF11";
          m(577) := x"FE40";
          m(578) := x"FFA4";
          m(579) := x"002F";
          m(580) := x"048E";
          m(581) := x"013F";
          m(582) := x"FFAC";
          m(583) := x"FFC7";
          m(584) := x"FCFF";
          m(585) := x"FDD4";
          m(586) := x"0001";
          m(587) := x"000B";
          m(588) := x"0028";
          m(589) := x"FFE0";
          m(590) := x"0089";
          m(591) := x"01C8";
          m(592) := x"0325";
          m(593) := x"FF8C";
          m(594) := x"0246";
          m(595) := x"044F";
          m(596) := x"02D4";
          m(597) := x"0083";
          m(598) := x"FF86";
          m(599) := x"011A";
          m(600) := x"FDC0";
          m(601) := x"00E7";
          m(602) := x"063B";
          m(603) := x"0612";
          m(604) := x"FD17";
          m(605) := x"FE8C";
          m(606) := x"040D";
          m(607) := x"FFE2";
          m(608) := x"0291";
          m(609) := x"007A";
          m(610) := x"002E";
          m(611) := x"FF5C";
          m(612) := x"FDC1";
          m(613) := x"FF79";
          m(614) := x"FFD3";
          m(615) := x"FFF8";
          m(616) := x"0027";
          m(617) := x"0000";
          m(618) := x"0046";
          m(619) := x"010B";
          m(620) := x"0257";
          m(621) := x"0540";
          m(622) := x"0687";
          m(623) := x"022A";
          m(624) := x"FBB5";
          m(625) := x"00FB";
          m(626) := x"007A";
          m(627) := x"FE0E";
          m(628) := x"FC33";
          m(629) := x"FF40";
          m(630) := x"0817";
          m(631) := x"043F";
          m(632) := x"056F";
          m(633) := x"014D";
          m(634) := x"0320";
          m(635) := x"FF3D";
          m(636) := x"FFA7";
          m(637) := x"022A";
          m(638) := x"0099";
          m(639) := x"FFF1";
          m(640) := x"FFEE";
          m(641) := x"FFD2";
          m(642) := x"0022";
          m(643) := x"FFF2";
          m(644) := x"FFFA";
          m(645) := x"FFF8";
          m(646) := x"016C";
          m(647) := x"0156";
          m(648) := x"038E";
          m(649) := x"07CC";
          m(650) := x"08CB";
          m(651) := x"0082";
          m(652) := x"FFEE";
          m(653) := x"FFB7";
          m(654) := x"FE5C";
          m(655) := x"0257";
          m(656) := x"FDF2";
          m(657) := x"013D";
          m(658) := x"0011";
          m(659) := x"0130";
          m(660) := x"0828";
          m(661) := x"04B3";
          m(662) := x"03F9";
          m(663) := x"0280";
          m(664) := x"0187";
          m(665) := x"01A0";
          m(666) := x"0122";
          m(667) := x"FFBC";
          m(668) := x"FFF9";
          m(669) := x"0063";
          m(670) := x"0015";
          m(671) := x"0009";
          m(672) := x"0025";
          m(673) := x"0001";
          m(674) := x"011F";
          m(675) := x"016B";
          m(676) := x"021F";
          m(677) := x"01E5";
          m(678) := x"0076";
          m(679) := x"035D";
          m(680) := x"036F";
          m(681) := x"FAC6";
          m(682) := x"FC4A";
          m(683) := x"02A2";
          m(684) := x"020A";
          m(685) := x"01BE";
          m(686) := x"04BE";
          m(687) := x"036A";
          m(688) := x"0313";
          m(689) := x"01FD";
          m(690) := x"03D6";
          m(691) := x"00D2";
          m(692) := x"FFB6";
          m(693) := x"FF6D";
          m(694) := x"FF21";
          m(695) := x"FECD";
          m(696) := x"0123";
          m(697) := x"FFD6";
          m(698) := x"FFBB";
          m(699) := x"FFC1";
          m(700) := x"FFF0";
          m(701) := x"0034";
          m(702) := x"FFFC";
          m(703) := x"0032";
          m(704) := x"FFBA";
          m(705) := x"FFE8";
          m(706) := x"FE86";
          m(707) := x"FF7E";
          m(708) := x"01D9";
          m(709) := x"010A";
          m(710) := x"0620";
          m(711) := x"0111";
          m(712) := x"FC01";
          m(713) := x"014A";
          m(714) := x"FB3A";
          m(715) := x"FECE";
          m(716) := x"FEF6";
          m(717) := x"0042";
          m(718) := x"FF20";
          m(719) := x"0136";
          m(720) := x"FEE8";
          m(721) := x"0082";
          m(722) := x"0248";
          m(723) := x"0260";
          m(724) := x"016A";
          m(725) := x"0001";
          m(726) := x"001F";
          m(727) := x"0007";
          m(728) := x"0033";
          m(729) := x"FFFD";
          m(730) := x"0026";
          m(731) := x"FFDB";
          m(732) := x"FF58";
          m(733) := x"FE92";
          m(734) := x"FD2B";
          m(735) := x"FEE0";
          m(736) := x"FEBF";
          m(737) := x"FD1D";
          m(738) := x"008B";
          m(739) := x"020B";
          m(740) := x"0112";
          m(741) := x"FCD8";
          m(742) := x"FC5C";
          m(743) := x"FEFA";
          m(744) := x"003C";
          m(745) := x"FE73";
          m(746) := x"FEA5";
          m(747) := x"FF49";
          m(748) := x"FF68";
          m(749) := x"006A";
          m(750) := x"008D";
          m(751) := x"002A";
          m(752) := x"FFF8";
          m(753) := x"FFF9";
          m(754) := x"000F";
          m(755) := x"0002";
          m(756) := x"0000";
          m(757) := x"FFD2";
          m(758) := x"FFF4";
          m(759) := x"FFE4";
          m(760) := x"000C";
          m(761) := x"FFC3";
          m(762) := x"FFF2";
          m(763) := x"FFDB";
          m(764) := x"FF95";
          m(765) := x"FFB9";
          m(766) := x"0007";
          m(767) := x"FFEA";
          m(768) := x"FFD0";
          m(769) := x"FFF6";
          m(770) := x"FF55";
          m(771) := x"FF10";
          m(772) := x"FF40";
          m(773) := x"FF59";
          m(774) := x"FEBC";
          m(775) := x"FF79";
          m(776) := x"FF5F";
          m(777) := x"FF76";
          m(778) := x"FFE7";
          m(779) := x"0019";
          m(780) := x"FFEB";
          m(781) := x"FFCD";
          m(782) := x"FFFA";
          m(783) := x"FFF8";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_26.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 26) then
          m(0) := x"FFF9";
          m(1) := x"0005";
          m(2) := x"0017";
          m(3) := x"0011";
          m(4) := x"FFF6";
          m(5) := x"0000";
          m(6) := x"003C";
          m(7) := x"000F";
          m(8) := x"002E";
          m(9) := x"FFE9";
          m(10) := x"000F";
          m(11) := x"FFF3";
          m(12) := x"FFD9";
          m(13) := x"FFEA";
          m(14) := x"0011";
          m(15) := x"003E";
          m(16) := x"0000";
          m(17) := x"FFF8";
          m(18) := x"000E";
          m(19) := x"FFE7";
          m(20) := x"FFF6";
          m(21) := x"001F";
          m(22) := x"0017";
          m(23) := x"0043";
          m(24) := x"0023";
          m(25) := x"0009";
          m(26) := x"FFF0";
          m(27) := x"FFE8";
          m(28) := x"FFF3";
          m(29) := x"0019";
          m(30) := x"001C";
          m(31) := x"001F";
          m(32) := x"FFDF";
          m(33) := x"FFEC";
          m(34) := x"FFED";
          m(35) := x"FFCB";
          m(36) := x"0027";
          m(37) := x"001F";
          m(38) := x"001F";
          m(39) := x"FFEF";
          m(40) := x"FFF9";
          m(41) := x"000F";
          m(42) := x"FF85";
          m(43) := x"FF89";
          m(44) := x"00D5";
          m(45) := x"00A6";
          m(46) := x"FFCB";
          m(47) := x"FFF7";
          m(48) := x"FFC0";
          m(49) := x"FFBC";
          m(50) := x"0011";
          m(51) := x"001B";
          m(52) := x"FFF1";
          m(53) := x"FFC0";
          m(54) := x"002C";
          m(55) := x"0016";
          m(56) := x"0002";
          m(57) := x"0015";
          m(58) := x"0014";
          m(59) := x"FFEB";
          m(60) := x"FFE7";
          m(61) := x"FFFF";
          m(62) := x"FFE6";
          m(63) := x"FF84";
          m(64) := x"FF92";
          m(65) := x"FF45";
          m(66) := x"0010";
          m(67) := x"FFC4";
          m(68) := x"FF15";
          m(69) := x"FEC2";
          m(70) := x"FE51";
          m(71) := x"FDD9";
          m(72) := x"FF9D";
          m(73) := x"FEF7";
          m(74) := x"FE22";
          m(75) := x"FDA4";
          m(76) := x"FEA9";
          m(77) := x"FED2";
          m(78) := x"FF79";
          m(79) := x"FFC6";
          m(80) := x"FFEB";
          m(81) := x"000A";
          m(82) := x"001A";
          m(83) := x"0037";
          m(84) := x"001B";
          m(85) := x"FFF0";
          m(86) := x"FFEF";
          m(87) := x"0013";
          m(88) := x"FFDB";
          m(89) := x"009D";
          m(90) := x"0065";
          m(91) := x"001D";
          m(92) := x"FFA0";
          m(93) := x"FF74";
          m(94) := x"00A7";
          m(95) := x"FE96";
          m(96) := x"FEF7";
          m(97) := x"FFB5";
          m(98) := x"0047";
          m(99) := x"0142";
          m(100) := x"0108";
          m(101) := x"0153";
          m(102) := x"0062";
          m(103) := x"FBBB";
          m(104) := x"FE8C";
          m(105) := x"FC5D";
          m(106) := x"FD00";
          m(107) := x"FF2A";
          m(108) := x"00CA";
          m(109) := x"00F3";
          m(110) := x"0009";
          m(111) := x"FFF0";
          m(112) := x"FFF9";
          m(113) := x"0002";
          m(114) := x"FFDE";
          m(115) := x"002F";
          m(116) := x"0022";
          m(117) := x"005C";
          m(118) := x"FFC4";
          m(119) := x"FF53";
          m(120) := x"006A";
          m(121) := x"01F4";
          m(122) := x"00C4";
          m(123) := x"FF8F";
          m(124) := x"0181";
          m(125) := x"0230";
          m(126) := x"FEA6";
          m(127) := x"FCE4";
          m(128) := x"F9F2";
          m(129) := x"FB68";
          m(130) := x"034C";
          m(131) := x"00F5";
          m(132) := x"FE5E";
          m(133) := x"FCC5";
          m(134) := x"FD90";
          m(135) := x"FF8A";
          m(136) := x"0215";
          m(137) := x"004A";
          m(138) := x"0000";
          m(139) := x"FFAC";
          m(140) := x"FFC4";
          m(141) := x"0030";
          m(142) := x"FFE6";
          m(143) := x"0000";
          m(144) := x"FFD5";
          m(145) := x"006C";
          m(146) := x"FF50";
          m(147) := x"FF2F";
          m(148) := x"008F";
          m(149) := x"FEDC";
          m(150) := x"FC9F";
          m(151) := x"00E8";
          m(152) := x"0109";
          m(153) := x"050E";
          m(154) := x"FEF1";
          m(155) := x"0215";
          m(156) := x"01D1";
          m(157) := x"FEE7";
          m(158) := x"0146";
          m(159) := x"FD78";
          m(160) := x"FC33";
          m(161) := x"007C";
          m(162) := x"022E";
          m(163) := x"01DF";
          m(164) := x"01B8";
          m(165) := x"FF62";
          m(166) := x"FF3D";
          m(167) := x"FFC0";
          m(168) := x"0000";
          m(169) := x"000E";
          m(170) := x"FFF3";
          m(171) := x"0003";
          m(172) := x"FFB6";
          m(173) := x"FF89";
          m(174) := x"FD6A";
          m(175) := x"FAF8";
          m(176) := x"FDBB";
          m(177) := x"FD94";
          m(178) := x"FE62";
          m(179) := x"004A";
          m(180) := x"03EB";
          m(181) := x"0046";
          m(182) := x"FE1D";
          m(183) := x"F833";
          m(184) := x"0100";
          m(185) := x"00AC";
          m(186) := x"03CE";
          m(187) := x"02BC";
          m(188) := x"023D";
          m(189) := x"041C";
          m(190) := x"0395";
          m(191) := x"0165";
          m(192) := x"02EA";
          m(193) := x"0067";
          m(194) := x"0083";
          m(195) := x"FF6E";
          m(196) := x"FFE2";
          m(197) := x"0023";
          m(198) := x"FFCF";
          m(199) := x"0036";
          m(200) := x"FFC4";
          m(201) := x"FD8A";
          m(202) := x"FD3C";
          m(203) := x"FAA6";
          m(204) := x"FA27";
          m(205) := x"F8E1";
          m(206) := x"FB81";
          m(207) := x"FD02";
          m(208) := x"FEE2";
          m(209) := x"FB97";
          m(210) := x"FE59";
          m(211) := x"FB6C";
          m(212) := x"FE39";
          m(213) := x"FCA4";
          m(214) := x"FE52";
          m(215) := x"FF2C";
          m(216) := x"008F";
          m(217) := x"F9C6";
          m(218) := x"00BA";
          m(219) := x"02A4";
          m(220) := x"0334";
          m(221) := x"01ED";
          m(222) := x"0202";
          m(223) := x"FFDA";
          m(224) := x"FFFA";
          m(225) := x"008D";
          m(226) := x"002C";
          m(227) := x"005C";
          m(228) := x"FF4B";
          m(229) := x"FCFF";
          m(230) := x"FEF4";
          m(231) := x"FC8E";
          m(232) := x"FBAA";
          m(233) := x"F724";
          m(234) := x"F92D";
          m(235) := x"F613";
          m(236) := x"FAC9";
          m(237) := x"F7A0";
          m(238) := x"F9CF";
          m(239) := x"FB05";
          m(240) := x"FD96";
          m(241) := x"FC04";
          m(242) := x"0314";
          m(243) := x"028B";
          m(244) := x"0585";
          m(245) := x"025D";
          m(246) := x"01A4";
          m(247) := x"0194";
          m(248) := x"0337";
          m(249) := x"03DE";
          m(250) := x"01D9";
          m(251) := x"003D";
          m(252) := x"FFCC";
          m(253) := x"010C";
          m(254) := x"008D";
          m(255) := x"0150";
          m(256) := x"FF47";
          m(257) := x"FEE0";
          m(258) := x"0140";
          m(259) := x"FD87";
          m(260) := x"FBA6";
          m(261) := x"F7DB";
          m(262) := x"F636";
          m(263) := x"FA99";
          m(264) := x"FEE2";
          m(265) := x"FA65";
          m(266) := x"FDE0";
          m(267) := x"FDDB";
          m(268) := x"FF2F";
          m(269) := x"025A";
          m(270) := x"FDF3";
          m(271) := x"FD48";
          m(272) := x"FE2B";
          m(273) := x"00AD";
          m(274) := x"FF5A";
          m(275) := x"FDF2";
          m(276) := x"0442";
          m(277) := x"058E";
          m(278) := x"02A8";
          m(279) := x"00A7";
          m(280) := x"001C";
          m(281) := x"00B7";
          m(282) := x"00E2";
          m(283) := x"0285";
          m(284) := x"0090";
          m(285) := x"0173";
          m(286) := x"008C";
          m(287) := x"FE8F";
          m(288) := x"FB67";
          m(289) := x"FF97";
          m(290) := x"02F8";
          m(291) := x"0235";
          m(292) := x"0022";
          m(293) := x"070F";
          m(294) := x"0464";
          m(295) := x"067C";
          m(296) := x"0625";
          m(297) := x"FB3C";
          m(298) := x"FB8B";
          m(299) := x"FC4B";
          m(300) := x"00FD";
          m(301) := x"FDB7";
          m(302) := x"0018";
          m(303) := x"0229";
          m(304) := x"0445";
          m(305) := x"06C5";
          m(306) := x"015B";
          m(307) := x"FFEF";
          m(308) := x"FFE1";
          m(309) := x"0040";
          m(310) := x"01BB";
          m(311) := x"033B";
          m(312) := x"03BE";
          m(313) := x"0355";
          m(314) := x"FE53";
          m(315) := x"0150";
          m(316) := x"046B";
          m(317) := x"03A1";
          m(318) := x"00EC";
          m(319) := x"03EA";
          m(320) := x"040C";
          m(321) := x"06D5";
          m(322) := x"02F3";
          m(323) := x"07C7";
          m(324) := x"FEB7";
          m(325) := x"01EC";
          m(326) := x"FEFA";
          m(327) := x"0286";
          m(328) := x"02A9";
          m(329) := x"0106";
          m(330) := x"00B9";
          m(331) := x"02CA";
          m(332) := x"017E";
          m(333) := x"030D";
          m(334) := x"005B";
          m(335) := x"0030";
          m(336) := x"0000";
          m(337) := x"0020";
          m(338) := x"00D9";
          m(339) := x"01AE";
          m(340) := x"0183";
          m(341) := x"0256";
          m(342) := x"FC33";
          m(343) := x"0321";
          m(344) := x"044E";
          m(345) := x"02E6";
          m(346) := x"025C";
          m(347) := x"0248";
          m(348) := x"0810";
          m(349) := x"03F8";
          m(350) := x"0298";
          m(351) := x"044C";
          m(352) := x"0455";
          m(353) := x"0264";
          m(354) := x"0186";
          m(355) := x"FED1";
          m(356) := x"FE34";
          m(357) := x"FD53";
          m(358) := x"FD6B";
          m(359) := x"FC55";
          m(360) := x"FBDC";
          m(361) := x"003F";
          m(362) := x"0090";
          m(363) := x"0002";
          m(364) := x"000A";
          m(365) := x"004A";
          m(366) := x"009C";
          m(367) := x"0239";
          m(368) := x"05ED";
          m(369) := x"0665";
          m(370) := x"01FF";
          m(371) := x"FDF2";
          m(372) := x"FF27";
          m(373) := x"FD6E";
          m(374) := x"006E";
          m(375) := x"025D";
          m(376) := x"0764";
          m(377) := x"0003";
          m(378) := x"0181";
          m(379) := x"FF78";
          m(380) := x"0294";
          m(381) := x"FD3A";
          m(382) := x"0233";
          m(383) := x"FDE0";
          m(384) := x"FA2F";
          m(385) := x"FB20";
          m(386) := x"FB3D";
          m(387) := x"FE40";
          m(388) := x"FE9C";
          m(389) := x"004A";
          m(390) := x"FFB0";
          m(391) := x"FEFE";
          m(392) := x"FFF0";
          m(393) := x"001C";
          m(394) := x"004A";
          m(395) := x"028A";
          m(396) := x"0357";
          m(397) := x"03A0";
          m(398) := x"0443";
          m(399) := x"FF14";
          m(400) := x"FD04";
          m(401) := x"0136";
          m(402) := x"FE69";
          m(403) := x"FF9C";
          m(404) := x"016D";
          m(405) := x"FBBE";
          m(406) := x"F98F";
          m(407) := x"F7D1";
          m(408) := x"FD87";
          m(409) := x"FFFA";
          m(410) := x"00E7";
          m(411) := x"FDC8";
          m(412) := x"FAF9";
          m(413) := x"FD4C";
          m(414) := x"FE17";
          m(415) := x"000A";
          m(416) := x"0170";
          m(417) := x"FEDB";
          m(418) := x"FFC8";
          m(419) := x"0011";
          m(420) := x"FFEC";
          m(421) := x"0014";
          m(422) := x"0050";
          m(423) := x"00F5";
          m(424) := x"FFF5";
          m(425) := x"00D9";
          m(426) := x"02D0";
          m(427) := x"0151";
          m(428) := x"FE9B";
          m(429) := x"02AD";
          m(430) := x"F88F";
          m(431) := x"FABB";
          m(432) := x"FBFF";
          m(433) := x"FB7B";
          m(434) := x"F9CF";
          m(435) := x"FC7E";
          m(436) := x"F867";
          m(437) := x"FCD9";
          m(438) := x"011A";
          m(439) := x"06D5";
          m(440) := x"0213";
          m(441) := x"FEF0";
          m(442) := x"FE38";
          m(443) := x"008D";
          m(444) := x"001A";
          m(445) := x"FF9F";
          m(446) := x"00A5";
          m(447) := x"0042";
          m(448) := x"FFEC";
          m(449) := x"FFCE";
          m(450) := x"FFF3";
          m(451) := x"010C";
          m(452) := x"009F";
          m(453) := x"FC32";
          m(454) := x"FD6B";
          m(455) := x"FC48";
          m(456) := x"FB4E";
          m(457) := x"F331";
          m(458) := x"F28B";
          m(459) := x"F66C";
          m(460) := x"F852";
          m(461) := x"F95C";
          m(462) := x"F940";
          m(463) := x"FDE4";
          m(464) := x"FA7D";
          m(465) := x"FDE3";
          m(466) := x"02D7";
          m(467) := x"026D";
          m(468) := x"046C";
          m(469) := x"FF60";
          m(470) := x"000F";
          m(471) := x"FE28";
          m(472) := x"FB6C";
          m(473) := x"FDFD";
          m(474) := x"0004";
          m(475) := x"FFF4";
          m(476) := x"0012";
          m(477) := x"003B";
          m(478) := x"FF7A";
          m(479) := x"0275";
          m(480) := x"00FD";
          m(481) := x"FF60";
          m(482) := x"FE95";
          m(483) := x"FDF4";
          m(484) := x"FD25";
          m(485) := x"F94F";
          m(486) := x"F78D";
          m(487) := x"FAE2";
          m(488) := x"F8BF";
          m(489) := x"F66C";
          m(490) := x"FE98";
          m(491) := x"FF59";
          m(492) := x"0417";
          m(493) := x"01DA";
          m(494) := x"000A";
          m(495) := x"FE1E";
          m(496) := x"FF24";
          m(497) := x"FEC2";
          m(498) := x"FEC6";
          m(499) := x"FD00";
          m(500) := x"FDA3";
          m(501) := x"FE0A";
          m(502) := x"FFC6";
          m(503) := x"003E";
          m(504) := x"FFE6";
          m(505) := x"FFD3";
          m(506) := x"0001";
          m(507) := x"04ED";
          m(508) := x"03C2";
          m(509) := x"0472";
          m(510) := x"0133";
          m(511) := x"FE5C";
          m(512) := x"082E";
          m(513) := x"067C";
          m(514) := x"032A";
          m(515) := x"0580";
          m(516) := x"02AF";
          m(517) := x"0450";
          m(518) := x"01A6";
          m(519) := x"080B";
          m(520) := x"0379";
          m(521) := x"03DE";
          m(522) := x"006C";
          m(523) := x"FB64";
          m(524) := x"005A";
          m(525) := x"FF81";
          m(526) := x"FEED";
          m(527) := x"FD8C";
          m(528) := x"FE63";
          m(529) := x"FF08";
          m(530) := x"0027";
          m(531) := x"0003";
          m(532) := x"FFCD";
          m(533) := x"001B";
          m(534) := x"001F";
          m(535) := x"05EF";
          m(536) := x"0671";
          m(537) := x"0502";
          m(538) := x"062C";
          m(539) := x"0465";
          m(540) := x"062A";
          m(541) := x"0372";
          m(542) := x"020B";
          m(543) := x"0150";
          m(544) := x"0531";
          m(545) := x"076B";
          m(546) := x"0159";
          m(547) := x"0378";
          m(548) := x"FDE6";
          m(549) := x"FF8F";
          m(550) := x"FF3E";
          m(551) := x"FDB1";
          m(552) := x"FF71";
          m(553) := x"F9D3";
          m(554) := x"FC37";
          m(555) := x"FCF3";
          m(556) := x"FED3";
          m(557) := x"FFB3";
          m(558) := x"FFD6";
          m(559) := x"0007";
          m(560) := x"FFEC";
          m(561) := x"0037";
          m(562) := x"0012";
          m(563) := x"023F";
          m(564) := x"01F9";
          m(565) := x"013A";
          m(566) := x"025E";
          m(567) := x"FF9B";
          m(568) := x"0536";
          m(569) := x"054B";
          m(570) := x"0476";
          m(571) := x"0569";
          m(572) := x"04FB";
          m(573) := x"096A";
          m(574) := x"034F";
          m(575) := x"FF82";
          m(576) := x"FACC";
          m(577) := x"FFD6";
          m(578) := x"0152";
          m(579) := x"FF28";
          m(580) := x"FAAA";
          m(581) := x"F8B0";
          m(582) := x"FB83";
          m(583) := x"FD22";
          m(584) := x"FE6D";
          m(585) := x"FF58";
          m(586) := x"FFCC";
          m(587) := x"0000";
          m(588) := x"FFFA";
          m(589) := x"0001";
          m(590) := x"FFD1";
          m(591) := x"FF4B";
          m(592) := x"FDC9";
          m(593) := x"FC48";
          m(594) := x"FC81";
          m(595) := x"00E9";
          m(596) := x"0688";
          m(597) := x"0089";
          m(598) := x"FDD3";
          m(599) := x"0212";
          m(600) := x"FC51";
          m(601) := x"000C";
          m(602) := x"FA75";
          m(603) := x"FD20";
          m(604) := x"FB85";
          m(605) := x"0093";
          m(606) := x"FF94";
          m(607) := x"FCBC";
          m(608) := x"FB02";
          m(609) := x"FAD4";
          m(610) := x"FB55";
          m(611) := x"FD43";
          m(612) := x"FE85";
          m(613) := x"FFE5";
          m(614) := x"0010";
          m(615) := x"0009";
          m(616) := x"0032";
          m(617) := x"FFDF";
          m(618) := x"FFCA";
          m(619) := x"FF1A";
          m(620) := x"FFA6";
          m(621) := x"FB9F";
          m(622) := x"FB23";
          m(623) := x"FF5D";
          m(624) := x"0062";
          m(625) := x"0555";
          m(626) := x"00E9";
          m(627) := x"0150";
          m(628) := x"05DD";
          m(629) := x"00DC";
          m(630) := x"007C";
          m(631) := x"038A";
          m(632) := x"FBB7";
          m(633) := x"FB26";
          m(634) := x"F8F0";
          m(635) := x"FC56";
          m(636) := x"FC9F";
          m(637) := x"FC0B";
          m(638) := x"FDD1";
          m(639) := x"FEFD";
          m(640) := x"FF67";
          m(641) := x"FFE3";
          m(642) := x"FFE6";
          m(643) := x"0000";
          m(644) := x"FFB4";
          m(645) := x"FFFC";
          m(646) := x"0000";
          m(647) := x"013F";
          m(648) := x"0192";
          m(649) := x"0184";
          m(650) := x"FE5B";
          m(651) := x"FE53";
          m(652) := x"00EF";
          m(653) := x"01D4";
          m(654) := x"03EB";
          m(655) := x"0470";
          m(656) := x"FEB0";
          m(657) := x"F965";
          m(658) := x"FF49";
          m(659) := x"FED0";
          m(660) := x"FCD6";
          m(661) := x"FBD0";
          m(662) := x"FBE5";
          m(663) := x"FC5A";
          m(664) := x"FE33";
          m(665) := x"FD77";
          m(666) := x"FE3A";
          m(667) := x"FF6D";
          m(668) := x"FF6D";
          m(669) := x"0003";
          m(670) := x"FFC7";
          m(671) := x"FFF1";
          m(672) := x"0030";
          m(673) := x"0019";
          m(674) := x"000F";
          m(675) := x"0159";
          m(676) := x"0077";
          m(677) := x"022D";
          m(678) := x"FFCB";
          m(679) := x"FEAA";
          m(680) := x"FE66";
          m(681) := x"FA37";
          m(682) := x"F7E8";
          m(683) := x"FD6D";
          m(684) := x"FB5F";
          m(685) := x"FD58";
          m(686) := x"03B5";
          m(687) := x"FD48";
          m(688) := x"FD33";
          m(689) := x"FF4D";
          m(690) := x"FE85";
          m(691) := x"FE67";
          m(692) := x"FE8A";
          m(693) := x"FEEB";
          m(694) := x"FF11";
          m(695) := x"FFAD";
          m(696) := x"FFFC";
          m(697) := x"001E";
          m(698) := x"FFD6";
          m(699) := x"FFC8";
          m(700) := x"FFE4";
          m(701) := x"FFC8";
          m(702) := x"0002";
          m(703) := x"0018";
          m(704) := x"002F";
          m(705) := x"002D";
          m(706) := x"FF89";
          m(707) := x"FFA8";
          m(708) := x"FD2C";
          m(709) := x"FDE6";
          m(710) := x"FDC2";
          m(711) := x"0094";
          m(712) := x"FF5F";
          m(713) := x"FF6C";
          m(714) := x"017B";
          m(715) := x"FCE3";
          m(716) := x"FF16";
          m(717) := x"0015";
          m(718) := x"0097";
          m(719) := x"0048";
          m(720) := x"FF97";
          m(721) := x"FFC1";
          m(722) := x"0025";
          m(723) := x"FF2D";
          m(724) := x"FFDE";
          m(725) := x"FFF5";
          m(726) := x"FFF9";
          m(727) := x"0017";
          m(728) := x"0001";
          m(729) := x"FFD4";
          m(730) := x"FFEE";
          m(731) := x"0034";
          m(732) := x"FFC8";
          m(733) := x"0052";
          m(734) := x"FFD7";
          m(735) := x"FFE9";
          m(736) := x"006D";
          m(737) := x"0096";
          m(738) := x"FF70";
          m(739) := x"02E1";
          m(740) := x"0375";
          m(741) := x"02AE";
          m(742) := x"FEA1";
          m(743) := x"FD82";
          m(744) := x"FF11";
          m(745) := x"0022";
          m(746) := x"0007";
          m(747) := x"0068";
          m(748) := x"000D";
          m(749) := x"FFFE";
          m(750) := x"0047";
          m(751) := x"0007";
          m(752) := x"0006";
          m(753) := x"FFE2";
          m(754) := x"0020";
          m(755) := x"0005";
          m(756) := x"FFDA";
          m(757) := x"0045";
          m(758) := x"0039";
          m(759) := x"0007";
          m(760) := x"0007";
          m(761) := x"000F";
          m(762) := x"0021";
          m(763) := x"FFC8";
          m(764) := x"FFFF";
          m(765) := x"001A";
          m(766) := x"00C3";
          m(767) := x"FFE8";
          m(768) := x"FFE6";
          m(769) := x"0051";
          m(770) := x"0031";
          m(771) := x"FEF6";
          m(772) := x"FF49";
          m(773) := x"0004";
          m(774) := x"0031";
          m(775) := x"000D";
          m(776) := x"0005";
          m(777) := x"FFE2";
          m(778) := x"005D";
          m(779) := x"002A";
          m(780) := x"FFD9";
          m(781) := x"0005";
          m(782) := x"0020";
          m(783) := x"FFCC";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_27.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 27) then
          m(0) := x"0026";
          m(1) := x"003A";
          m(2) := x"FFE3";
          m(3) := x"0011";
          m(4) := x"001E";
          m(5) := x"0008";
          m(6) := x"FFC1";
          m(7) := x"0057";
          m(8) := x"FFF3";
          m(9) := x"FFEE";
          m(10) := x"FFDA";
          m(11) := x"FFF2";
          m(12) := x"0030";
          m(13) := x"0052";
          m(14) := x"FFFF";
          m(15) := x"000B";
          m(16) := x"FFEE";
          m(17) := x"FFF7";
          m(18) := x"FFF5";
          m(19) := x"0004";
          m(20) := x"0005";
          m(21) := x"0030";
          m(22) := x"0002";
          m(23) := x"FFE7";
          m(24) := x"FFF3";
          m(25) := x"0026";
          m(26) := x"FFE5";
          m(27) := x"FFEE";
          m(28) := x"000C";
          m(29) := x"FFD4";
          m(30) := x"0007";
          m(31) := x"0006";
          m(32) := x"FFF0";
          m(33) := x"FFD6";
          m(34) := x"FFEE";
          m(35) := x"0019";
          m(36) := x"FFC4";
          m(37) := x"FFE9";
          m(38) := x"0030";
          m(39) := x"FFF2";
          m(40) := x"FF84";
          m(41) := x"FFE2";
          m(42) := x"FFEE";
          m(43) := x"FF51";
          m(44) := x"FF88";
          m(45) := x"FFF6";
          m(46) := x"002B";
          m(47) := x"FFE1";
          m(48) := x"FFE0";
          m(49) := x"FFCD";
          m(50) := x"FFD1";
          m(51) := x"FFFE";
          m(52) := x"FFF1";
          m(53) := x"FFEA";
          m(54) := x"FFEA";
          m(55) := x"003B";
          m(56) := x"003D";
          m(57) := x"0009";
          m(58) := x"FFF6";
          m(59) := x"FFB8";
          m(60) := x"FFD4";
          m(61) := x"FFC9";
          m(62) := x"FFDD";
          m(63) := x"FFEC";
          m(64) := x"0000";
          m(65) := x"FFE4";
          m(66) := x"FFA0";
          m(67) := x"FFC6";
          m(68) := x"00A0";
          m(69) := x"00B5";
          m(70) := x"FF8F";
          m(71) := x"FFD5";
          m(72) := x"0066";
          m(73) := x"FF08";
          m(74) := x"FEF2";
          m(75) := x"FEDB";
          m(76) := x"FF33";
          m(77) := x"FF1E";
          m(78) := x"FF86";
          m(79) := x"FFAE";
          m(80) := x"0065";
          m(81) := x"003B";
          m(82) := x"0019";
          m(83) := x"0028";
          m(84) := x"FFF2";
          m(85) := x"FFF5";
          m(86) := x"FFEE";
          m(87) := x"FFDC";
          m(88) := x"0027";
          m(89) := x"0038";
          m(90) := x"FFFD";
          m(91) := x"007E";
          m(92) := x"021C";
          m(93) := x"017E";
          m(94) := x"01D4";
          m(95) := x"0010";
          m(96) := x"0226";
          m(97) := x"0161";
          m(98) := x"FC58";
          m(99) := x"FD79";
          m(100) := x"FDF8";
          m(101) := x"FDD2";
          m(102) := x"FD9C";
          m(103) := x"FD39";
          m(104) := x"FC9B";
          m(105) := x"FDC4";
          m(106) := x"FE25";
          m(107) := x"FEC2";
          m(108) := x"0040";
          m(109) := x"0103";
          m(110) := x"0039";
          m(111) := x"FFDA";
          m(112) := x"FFEB";
          m(113) := x"FFB2";
          m(114) := x"0000";
          m(115) := x"FFF6";
          m(116) := x"004C";
          m(117) := x"0038";
          m(118) := x"0065";
          m(119) := x"020B";
          m(120) := x"0491";
          m(121) := x"04B8";
          m(122) := x"041A";
          m(123) := x"03AD";
          m(124) := x"052C";
          m(125) := x"0047";
          m(126) := x"FBF3";
          m(127) := x"FABF";
          m(128) := x"FDBA";
          m(129) := x"FEAF";
          m(130) := x"02DB";
          m(131) := x"FEA1";
          m(132) := x"FC03";
          m(133) := x"FD24";
          m(134) := x"FD82";
          m(135) := x"0030";
          m(136) := x"0391";
          m(137) := x"02F8";
          m(138) := x"0118";
          m(139) := x"001F";
          m(140) := x"001D";
          m(141) := x"0024";
          m(142) := x"FFFB";
          m(143) := x"0042";
          m(144) := x"000E";
          m(145) := x"FFB6";
          m(146) := x"FF99";
          m(147) := x"01CD";
          m(148) := x"028C";
          m(149) := x"029F";
          m(150) := x"04C1";
          m(151) := x"0469";
          m(152) := x"0458";
          m(153) := x"00AE";
          m(154) := x"FCFA";
          m(155) := x"FE8C";
          m(156) := x"FEC3";
          m(157) := x"FF76";
          m(158) := x"FCD0";
          m(159) := x"FAC8";
          m(160) := x"0010";
          m(161) := x"FF20";
          m(162) := x"01AA";
          m(163) := x"0201";
          m(164) := x"0229";
          m(165) := x"0229";
          m(166) := x"0079";
          m(167) := x"002B";
          m(168) := x"FFEB";
          m(169) := x"001C";
          m(170) := x"0001";
          m(171) := x"0034";
          m(172) := x"FF3D";
          m(173) := x"FE94";
          m(174) := x"FFA2";
          m(175) := x"01D1";
          m(176) := x"0450";
          m(177) := x"076C";
          m(178) := x"03F5";
          m(179) := x"04C4";
          m(180) := x"0846";
          m(181) := x"020C";
          m(182) := x"FB92";
          m(183) := x"FE5C";
          m(184) := x"01A9";
          m(185) := x"055E";
          m(186) := x"02C3";
          m(187) := x"0185";
          m(188) := x"03A1";
          m(189) := x"02EC";
          m(190) := x"03C8";
          m(191) := x"0393";
          m(192) := x"01C0";
          m(193) := x"01DC";
          m(194) := x"00FB";
          m(195) := x"006F";
          m(196) := x"002D";
          m(197) := x"001C";
          m(198) := x"FFDB";
          m(199) := x"FF27";
          m(200) := x"FE75";
          m(201) := x"FDEF";
          m(202) := x"FD50";
          m(203) := x"00E4";
          m(204) := x"052E";
          m(205) := x"0380";
          m(206) := x"0683";
          m(207) := x"0175";
          m(208) := x"03CD";
          m(209) := x"FB24";
          m(210) := x"FA79";
          m(211) := x"FCDB";
          m(212) := x"00E9";
          m(213) := x"FD59";
          m(214) := x"FCDB";
          m(215) := x"0241";
          m(216) := x"02E4";
          m(217) := x"01A6";
          m(218) := x"FF9C";
          m(219) := x"FFFE";
          m(220) := x"00DA";
          m(221) := x"01FC";
          m(222) := x"011F";
          m(223) := x"0064";
          m(224) := x"FFD7";
          m(225) := x"001A";
          m(226) := x"FF69";
          m(227) := x"FF24";
          m(228) := x"FE83";
          m(229) := x"FF5F";
          m(230) := x"0087";
          m(231) := x"0511";
          m(232) := x"02D8";
          m(233) := x"007A";
          m(234) := x"0333";
          m(235) := x"056B";
          m(236) := x"01E5";
          m(237) := x"FD9E";
          m(238) := x"FAF4";
          m(239) := x"FE8A";
          m(240) := x"FD3E";
          m(241) := x"FDC5";
          m(242) := x"FF05";
          m(243) := x"06D6";
          m(244) := x"04EC";
          m(245) := x"0080";
          m(246) := x"0165";
          m(247) := x"00E8";
          m(248) := x"01C6";
          m(249) := x"04C7";
          m(250) := x"0236";
          m(251) := x"0041";
          m(252) := x"000B";
          m(253) := x"000D";
          m(254) := x"FF6E";
          m(255) := x"FF7B";
          m(256) := x"FF23";
          m(257) := x"FF20";
          m(258) := x"00D9";
          m(259) := x"01D5";
          m(260) := x"0413";
          m(261) := x"01EC";
          m(262) := x"053F";
          m(263) := x"0889";
          m(264) := x"01A0";
          m(265) := x"F9B7";
          m(266) := x"FEA4";
          m(267) := x"0473";
          m(268) := x"FF61";
          m(269) := x"FF8C";
          m(270) := x"FF34";
          m(271) := x"FF97";
          m(272) := x"0069";
          m(273) := x"FE46";
          m(274) := x"012F";
          m(275) := x"FE07";
          m(276) := x"0240";
          m(277) := x"0454";
          m(278) := x"01B2";
          m(279) := x"0039";
          m(280) := x"0018";
          m(281) := x"0005";
          m(282) := x"FF33";
          m(283) := x"FE96";
          m(284) := x"0088";
          m(285) := x"0022";
          m(286) := x"02F0";
          m(287) := x"02A7";
          m(288) := x"02E1";
          m(289) := x"0657";
          m(290) := x"0732";
          m(291) := x"0468";
          m(292) := x"0124";
          m(293) := x"FEA7";
          m(294) := x"00E2";
          m(295) := x"04A8";
          m(296) := x"FD09";
          m(297) := x"FABC";
          m(298) := x"FE5D";
          m(299) := x"FF97";
          m(300) := x"FECA";
          m(301) := x"FC80";
          m(302) := x"0205";
          m(303) := x"0399";
          m(304) := x"0406";
          m(305) := x"0145";
          m(306) := x"0166";
          m(307) := x"000A";
          m(308) := x"FFEC";
          m(309) := x"FFF0";
          m(310) := x"003A";
          m(311) := x"FEBD";
          m(312) := x"02E1";
          m(313) := x"0274";
          m(314) := x"006F";
          m(315) := x"FEAB";
          m(316) := x"02CB";
          m(317) := x"0217";
          m(318) := x"0015";
          m(319) := x"075B";
          m(320) := x"0558";
          m(321) := x"FB7D";
          m(322) := x"03E2";
          m(323) := x"059B";
          m(324) := x"011D";
          m(325) := x"FEBF";
          m(326) := x"0053";
          m(327) := x"029F";
          m(328) := x"FED8";
          m(329) := x"FD1C";
          m(330) := x"01F5";
          m(331) := x"0295";
          m(332) := x"02AA";
          m(333) := x"01D6";
          m(334) := x"01D3";
          m(335) := x"FFE8";
          m(336) := x"0004";
          m(337) := x"FFF0";
          m(338) := x"FFA2";
          m(339) := x"FF20";
          m(340) := x"0102";
          m(341) := x"FDDB";
          m(342) := x"FCF6";
          m(343) := x"0194";
          m(344) := x"01A4";
          m(345) := x"0104";
          m(346) := x"03B2";
          m(347) := x"03B8";
          m(348) := x"FE79";
          m(349) := x"FFA6";
          m(350) := x"01F8";
          m(351) := x"085B";
          m(352) := x"011D";
          m(353) := x"038B";
          m(354) := x"0002";
          m(355) := x"074F";
          m(356) := x"0186";
          m(357) := x"FED5";
          m(358) := x"FFA4";
          m(359) := x"FE99";
          m(360) := x"FD6B";
          m(361) := x"002A";
          m(362) := x"00E9";
          m(363) := x"0002";
          m(364) := x"001A";
          m(365) := x"FFE4";
          m(366) := x"FFDF";
          m(367) := x"0084";
          m(368) := x"FDBC";
          m(369) := x"FE49";
          m(370) := x"FCA5";
          m(371) := x"FD92";
          m(372) := x"01A5";
          m(373) := x"00D0";
          m(374) := x"FFC8";
          m(375) := x"0655";
          m(376) := x"0250";
          m(377) := x"013E";
          m(378) := x"004A";
          m(379) := x"0C52";
          m(380) := x"06F0";
          m(381) := x"00B5";
          m(382) := x"001C";
          m(383) := x"04C9";
          m(384) := x"075B";
          m(385) := x"01E7";
          m(386) := x"FF29";
          m(387) := x"FF9D";
          m(388) := x"FD62";
          m(389) := x"FE4B";
          m(390) := x"0046";
          m(391) := x"002D";
          m(392) := x"0001";
          m(393) := x"FFF6";
          m(394) := x"FFAC";
          m(395) := x"006E";
          m(396) := x"0059";
          m(397) := x"FAE1";
          m(398) := x"FC47";
          m(399) := x"FBC6";
          m(400) := x"FCF6";
          m(401) := x"FEEF";
          m(402) := x"00B8";
          m(403) := x"0249";
          m(404) := x"FB70";
          m(405) := x"00E9";
          m(406) := x"0696";
          m(407) := x"0B42";
          m(408) := x"07D9";
          m(409) := x"028A";
          m(410) := x"0349";
          m(411) := x"013B";
          m(412) := x"00F5";
          m(413) := x"FEC4";
          m(414) := x"FB8F";
          m(415) := x"FF2F";
          m(416) := x"FF7C";
          m(417) := x"FEA9";
          m(418) := x"0134";
          m(419) := x"0005";
          m(420) := x"FFF8";
          m(421) := x"000B";
          m(422) := x"FF91";
          m(423) := x"0039";
          m(424) := x"00A2";
          m(425) := x"FF01";
          m(426) := x"FB44";
          m(427) := x"F6EF";
          m(428) := x"FB42";
          m(429) := x"FE4C";
          m(430) := x"FDDB";
          m(431) := x"00D9";
          m(432) := x"F9CD";
          m(433) := x"0060";
          m(434) := x"0E83";
          m(435) := x"0BD7";
          m(436) := x"0255";
          m(437) := x"FE39";
          m(438) := x"0285";
          m(439) := x"FF56";
          m(440) := x"FA50";
          m(441) := x"FA94";
          m(442) := x"F75E";
          m(443) := x"FD89";
          m(444) := x"FF44";
          m(445) := x"0071";
          m(446) := x"01FD";
          m(447) := x"FFDF";
          m(448) := x"FFE7";
          m(449) := x"FFDE";
          m(450) := x"FFA5";
          m(451) := x"0130";
          m(452) := x"00D0";
          m(453) := x"FC67";
          m(454) := x"FBEC";
          m(455) := x"F7CE";
          m(456) := x"FB82";
          m(457) := x"FA27";
          m(458) := x"FEB7";
          m(459) := x"FB84";
          m(460) := x"F947";
          m(461) := x"FBE9";
          m(462) := x"0A0A";
          m(463) := x"0AA1";
          m(464) := x"0289";
          m(465) := x"FC84";
          m(466) := x"FC86";
          m(467) := x"F84E";
          m(468) := x"F6C8";
          m(469) := x"FEE2";
          m(470) := x"FD72";
          m(471) := x"FDC6";
          m(472) := x"FD68";
          m(473) := x"0014";
          m(474) := x"00E3";
          m(475) := x"001C";
          m(476) := x"FFF7";
          m(477) := x"FFEC";
          m(478) := x"FF78";
          m(479) := x"0275";
          m(480) := x"FEF7";
          m(481) := x"FF83";
          m(482) := x"0149";
          m(483) := x"FDCD";
          m(484) := x"FB8F";
          m(485) := x"FB9C";
          m(486) := x"FC78";
          m(487) := x"FD61";
          m(488) := x"FC8E";
          m(489) := x"0242";
          m(490) := x"0814";
          m(491) := x"064A";
          m(492) := x"FEBD";
          m(493) := x"FAA7";
          m(494) := x"F876";
          m(495) := x"F9AC";
          m(496) := x"FC6B";
          m(497) := x"0333";
          m(498) := x"FBB2";
          m(499) := x"FC57";
          m(500) := x"FEBC";
          m(501) := x"00C1";
          m(502) := x"001D";
          m(503) := x"FFAE";
          m(504) := x"FFF8";
          m(505) := x"0006";
          m(506) := x"000D";
          m(507) := x"026E";
          m(508) := x"FEF5";
          m(509) := x"0015";
          m(510) := x"01FC";
          m(511) := x"0335";
          m(512) := x"0206";
          m(513) := x"FE7D";
          m(514) := x"01C7";
          m(515) := x"02BC";
          m(516) := x"FDFC";
          m(517) := x"018E";
          m(518) := x"06F7";
          m(519) := x"FDEC";
          m(520) := x"FBAC";
          m(521) := x"F7DA";
          m(522) := x"FD76";
          m(523) := x"FCC2";
          m(524) := x"FF08";
          m(525) := x"FD09";
          m(526) := x"FC7C";
          m(527) := x"FE14";
          m(528) := x"0045";
          m(529) := x"01B4";
          m(530) := x"001D";
          m(531) := x"FFD4";
          m(532) := x"0026";
          m(533) := x"0010";
          m(534) := x"001A";
          m(535) := x"0144";
          m(536) := x"FDCB";
          m(537) := x"FEC8";
          m(538) := x"00C6";
          m(539) := x"0308";
          m(540) := x"01BE";
          m(541) := x"FEA9";
          m(542) := x"FBC7";
          m(543) := x"FDB1";
          m(544) := x"0034";
          m(545) := x"02D8";
          m(546) := x"FECC";
          m(547) := x"FF8A";
          m(548) := x"00BA";
          m(549) := x"FFB3";
          m(550) := x"014F";
          m(551) := x"FF95";
          m(552) := x"FBBA";
          m(553) := x"FBB6";
          m(554) := x"FF60";
          m(555) := x"00B9";
          m(556) := x"0204";
          m(557) := x"0235";
          m(558) := x"002B";
          m(559) := x"FFEE";
          m(560) := x"FFE3";
          m(561) := x"FFDE";
          m(562) := x"0012";
          m(563) := x"00B0";
          m(564) := x"FE44";
          m(565) := x"FF22";
          m(566) := x"02FB";
          m(567) := x"FD2B";
          m(568) := x"FEFC";
          m(569) := x"FFEC";
          m(570) := x"FA53";
          m(571) := x"0066";
          m(572) := x"FD05";
          m(573) := x"FCDB";
          m(574) := x"FA89";
          m(575) := x"FD5B";
          m(576) := x"FF51";
          m(577) := x"0039";
          m(578) := x"FFCE";
          m(579) := x"FDA9";
          m(580) := x"FE00";
          m(581) := x"FFE1";
          m(582) := x"03F4";
          m(583) := x"0478";
          m(584) := x"0274";
          m(585) := x"0215";
          m(586) := x"001E";
          m(587) := x"FFFD";
          m(588) := x"0006";
          m(589) := x"FFE5";
          m(590) := x"002F";
          m(591) := x"FF71";
          m(592) := x"FF30";
          m(593) := x"FEE2";
          m(594) := x"0218";
          m(595) := x"0192";
          m(596) := x"004E";
          m(597) := x"012E";
          m(598) := x"03B5";
          m(599) := x"06E0";
          m(600) := x"FA95";
          m(601) := x"F951";
          m(602) := x"F5C5";
          m(603) := x"FBE1";
          m(604) := x"0219";
          m(605) := x"0328";
          m(606) := x"FDCE";
          m(607) := x"FF8A";
          m(608) := x"FEEB";
          m(609) := x"01B2";
          m(610) := x"FFAD";
          m(611) := x"0241";
          m(612) := x"02A9";
          m(613) := x"0164";
          m(614) := x"0007";
          m(615) := x"0019";
          m(616) := x"0005";
          m(617) := x"0010";
          m(618) := x"FFFF";
          m(619) := x"FFFE";
          m(620) := x"FF3A";
          m(621) := x"FC5C";
          m(622) := x"FEB5";
          m(623) := x"0469";
          m(624) := x"030A";
          m(625) := x"014F";
          m(626) := x"021A";
          m(627) := x"0217";
          m(628) := x"F8D6";
          m(629) := x"FAB7";
          m(630) := x"FBB3";
          m(631) := x"FAA8";
          m(632) := x"FF47";
          m(633) := x"FB1F";
          m(634) := x"FF5E";
          m(635) := x"FFEB";
          m(636) := x"005D";
          m(637) := x"FFF0";
          m(638) := x"0033";
          m(639) := x"01B1";
          m(640) := x"0268";
          m(641) := x"0140";
          m(642) := x"FFE6";
          m(643) := x"FFCE";
          m(644) := x"0018";
          m(645) := x"FFEE";
          m(646) := x"FFE8";
          m(647) := x"004A";
          m(648) := x"00A2";
          m(649) := x"FDA5";
          m(650) := x"FD0C";
          m(651) := x"0095";
          m(652) := x"030B";
          m(653) := x"04E3";
          m(654) := x"0321";
          m(655) := x"0193";
          m(656) := x"FF86";
          m(657) := x"0066";
          m(658) := x"FD52";
          m(659) := x"FA40";
          m(660) := x"FC64";
          m(661) := x"FC73";
          m(662) := x"00CA";
          m(663) := x"021F";
          m(664) := x"FEEE";
          m(665) := x"FF56";
          m(666) := x"0126";
          m(667) := x"0216";
          m(668) := x"025C";
          m(669) := x"00F9";
          m(670) := x"0008";
          m(671) := x"FFE3";
          m(672) := x"0001";
          m(673) := x"FFE4";
          m(674) := x"FFE2";
          m(675) := x"005D";
          m(676) := x"002C";
          m(677) := x"FFC5";
          m(678) := x"01A0";
          m(679) := x"032E";
          m(680) := x"0340";
          m(681) := x"0223";
          m(682) := x"0230";
          m(683) := x"00D7";
          m(684) := x"FF59";
          m(685) := x"0014";
          m(686) := x"FE9D";
          m(687) := x"F87F";
          m(688) := x"FA15";
          m(689) := x"FE72";
          m(690) := x"FFAE";
          m(691) := x"01C5";
          m(692) := x"01B2";
          m(693) := x"01AC";
          m(694) := x"019F";
          m(695) := x"016B";
          m(696) := x"010A";
          m(697) := x"001C";
          m(698) := x"000E";
          m(699) := x"FFFB";
          m(700) := x"FFF7";
          m(701) := x"0009";
          m(702) := x"000A";
          m(703) := x"001F";
          m(704) := x"000B";
          m(705) := x"012B";
          m(706) := x"0138";
          m(707) := x"00F3";
          m(708) := x"0014";
          m(709) := x"FFDC";
          m(710) := x"00B0";
          m(711) := x"FFAE";
          m(712) := x"FFA4";
          m(713) := x"04EC";
          m(714) := x"0125";
          m(715) := x"00CB";
          m(716) := x"01DB";
          m(717) := x"00AB";
          m(718) := x"0158";
          m(719) := x"035F";
          m(720) := x"01D8";
          m(721) := x"00AB";
          m(722) := x"0140";
          m(723) := x"019B";
          m(724) := x"00F0";
          m(725) := x"002B";
          m(726) := x"FFE7";
          m(727) := x"FFEF";
          m(728) := x"004C";
          m(729) := x"FFF1";
          m(730) := x"0014";
          m(731) := x"FFF6";
          m(732) := x"0032";
          m(733) := x"004D";
          m(734) := x"0002";
          m(735) := x"FF5C";
          m(736) := x"FE7B";
          m(737) := x"FDC3";
          m(738) := x"FE91";
          m(739) := x"0030";
          m(740) := x"FF54";
          m(741) := x"012E";
          m(742) := x"01A8";
          m(743) := x"0087";
          m(744) := x"0211";
          m(745) := x"00B4";
          m(746) := x"016D";
          m(747) := x"01A5";
          m(748) := x"011C";
          m(749) := x"FFD6";
          m(750) := x"FFB2";
          m(751) := x"FFF2";
          m(752) := x"FFF3";
          m(753) := x"0009";
          m(754) := x"004A";
          m(755) := x"0000";
          m(756) := x"FFF3";
          m(757) := x"0006";
          m(758) := x"0014";
          m(759) := x"0004";
          m(760) := x"002A";
          m(761) := x"0013";
          m(762) := x"001E";
          m(763) := x"0097";
          m(764) := x"0073";
          m(765) := x"FFEA";
          m(766) := x"0008";
          m(767) := x"FFC1";
          m(768) := x"FFE3";
          m(769) := x"0014";
          m(770) := x"0065";
          m(771) := x"0066";
          m(772) := x"FFD1";
          m(773) := x"FFB2";
          m(774) := x"FF88";
          m(775) := x"FFF5";
          m(776) := x"FFC1";
          m(777) := x"FFF8";
          m(778) := x"000D";
          m(779) := x"0006";
          m(780) := x"FFE6";
          m(781) := x"FFF7";
          m(782) := x"0003";
          m(783) := x"FFE2";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_28.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 28) then
          m(0) := x"FFE0";
          m(1) := x"FFF5";
          m(2) := x"0006";
          m(3) := x"FFDD";
          m(4) := x"FFED";
          m(5) := x"000E";
          m(6) := x"0032";
          m(7) := x"FFF7";
          m(8) := x"003D";
          m(9) := x"FFF4";
          m(10) := x"FFF5";
          m(11) := x"0028";
          m(12) := x"FFC9";
          m(13) := x"000C";
          m(14) := x"000D";
          m(15) := x"0000";
          m(16) := x"0028";
          m(17) := x"0005";
          m(18) := x"000C";
          m(19) := x"FFD3";
          m(20) := x"FFDE";
          m(21) := x"000D";
          m(22) := x"0016";
          m(23) := x"FFFE";
          m(24) := x"FFBE";
          m(25) := x"FFE9";
          m(26) := x"FFF0";
          m(27) := x"FFF0";
          m(28) := x"0023";
          m(29) := x"FFC5";
          m(30) := x"000E";
          m(31) := x"FFD5";
          m(32) := x"FFD4";
          m(33) := x"FFEE";
          m(34) := x"002A";
          m(35) := x"FFFD";
          m(36) := x"FFD0";
          m(37) := x"FFF5";
          m(38) := x"FFE6";
          m(39) := x"FFE4";
          m(40) := x"000E";
          m(41) := x"000E";
          m(42) := x"002D";
          m(43) := x"0081";
          m(44) := x"FFB6";
          m(45) := x"0011";
          m(46) := x"0023";
          m(47) := x"FFFB";
          m(48) := x"0028";
          m(49) := x"FFF1";
          m(50) := x"0008";
          m(51) := x"FFC3";
          m(52) := x"0001";
          m(53) := x"FFE4";
          m(54) := x"0010";
          m(55) := x"0025";
          m(56) := x"0013";
          m(57) := x"0003";
          m(58) := x"FFF9";
          m(59) := x"FFCC";
          m(60) := x"0009";
          m(61) := x"FFF6";
          m(62) := x"000F";
          m(63) := x"001F";
          m(64) := x"0005";
          m(65) := x"FFFE";
          m(66) := x"0004";
          m(67) := x"FFE0";
          m(68) := x"FFCA";
          m(69) := x"00C0";
          m(70) := x"01A8";
          m(71) := x"044D";
          m(72) := x"03D0";
          m(73) := x"018D";
          m(74) := x"0123";
          m(75) := x"0124";
          m(76) := x"010D";
          m(77) := x"008C";
          m(78) := x"006D";
          m(79) := x"002C";
          m(80) := x"FFF4";
          m(81) := x"002D";
          m(82) := x"FFE1";
          m(83) := x"0012";
          m(84) := x"FFFD";
          m(85) := x"0006";
          m(86) := x"FFC6";
          m(87) := x"0004";
          m(88) := x"FFF3";
          m(89) := x"FFF5";
          m(90) := x"001A";
          m(91) := x"FFDB";
          m(92) := x"001F";
          m(93) := x"0031";
          m(94) := x"FC4D";
          m(95) := x"FB56";
          m(96) := x"FCD2";
          m(97) := x"FD2B";
          m(98) := x"FCDF";
          m(99) := x"FE56";
          m(100) := x"000A";
          m(101) := x"FEA8";
          m(102) := x"0648";
          m(103) := x"048D";
          m(104) := x"FFC7";
          m(105) := x"FFCA";
          m(106) := x"0102";
          m(107) := x"01A5";
          m(108) := x"0157";
          m(109) := x"0028";
          m(110) := x"FFEE";
          m(111) := x"FFD7";
          m(112) := x"0011";
          m(113) := x"FFE2";
          m(114) := x"0005";
          m(115) := x"0008";
          m(116) := x"FFE9";
          m(117) := x"FF3F";
          m(118) := x"FED6";
          m(119) := x"FE32";
          m(120) := x"FDEB";
          m(121) := x"FB6B";
          m(122) := x"F877";
          m(123) := x"F8B0";
          m(124) := x"FC49";
          m(125) := x"FE3E";
          m(126) := x"FCAD";
          m(127) := x"FA3A";
          m(128) := x"02A7";
          m(129) := x"FEB3";
          m(130) := x"FD78";
          m(131) := x"01C6";
          m(132) := x"FF1F";
          m(133) := x"FDDA";
          m(134) := x"FDDE";
          m(135) := x"FF47";
          m(136) := x"FEBF";
          m(137) := x"FEF8";
          m(138) := x"FF8F";
          m(139) := x"000B";
          m(140) := x"0011";
          m(141) := x"FFF4";
          m(142) := x"FFE4";
          m(143) := x"FFEB";
          m(144) := x"FF40";
          m(145) := x"FCEE";
          m(146) := x"FC18";
          m(147) := x"FCB3";
          m(148) := x"FE64";
          m(149) := x"FB76";
          m(150) := x"FB18";
          m(151) := x"F9F9";
          m(152) := x"FB83";
          m(153) := x"F96A";
          m(154) := x"F953";
          m(155) := x"FEC3";
          m(156) := x"FB72";
          m(157) := x"F9CC";
          m(158) := x"F957";
          m(159) := x"FE6D";
          m(160) := x"FE20";
          m(161) := x"FE22";
          m(162) := x"FD14";
          m(163) := x"FE8D";
          m(164) := x"FF32";
          m(165) := x"FEB3";
          m(166) := x"0022";
          m(167) := x"FFDD";
          m(168) := x"FFDD";
          m(169) := x"FFD5";
          m(170) := x"0033";
          m(171) := x"FFC5";
          m(172) := x"FEBB";
          m(173) := x"FB17";
          m(174) := x"F9D5";
          m(175) := x"FACF";
          m(176) := x"F7F2";
          m(177) := x"F823";
          m(178) := x"F9A5";
          m(179) := x"F5CE";
          m(180) := x"F932";
          m(181) := x"F783";
          m(182) := x"FB07";
          m(183) := x"FD3F";
          m(184) := x"FABE";
          m(185) := x"FECD";
          m(186) := x"FBCA";
          m(187) := x"FF56";
          m(188) := x"003C";
          m(189) := x"0118";
          m(190) := x"FE39";
          m(191) := x"FEFD";
          m(192) := x"005F";
          m(193) := x"00D4";
          m(194) := x"0019";
          m(195) := x"0034";
          m(196) := x"FFC6";
          m(197) := x"FFD6";
          m(198) := x"FFF1";
          m(199) := x"FEE4";
          m(200) := x"FF5B";
          m(201) := x"FEB4";
          m(202) := x"FA13";
          m(203) := x"F96B";
          m(204) := x"F82F";
          m(205) := x"FAFB";
          m(206) := x"F8F6";
          m(207) := x"F714";
          m(208) := x"F636";
          m(209) := x"F6C7";
          m(210) := x"FF5B";
          m(211) := x"FAD0";
          m(212) := x"00ED";
          m(213) := x"00DB";
          m(214) := x"FED1";
          m(215) := x"FDDE";
          m(216) := x"00EC";
          m(217) := x"010B";
          m(218) := x"00C9";
          m(219) := x"0020";
          m(220) := x"0059";
          m(221) := x"FF75";
          m(222) := x"FFC1";
          m(223) := x"FFFC";
          m(224) := x"0006";
          m(225) := x"FFD6";
          m(226) := x"FFA7";
          m(227) := x"FECD";
          m(228) := x"FE92";
          m(229) := x"FF0B";
          m(230) := x"FF3A";
          m(231) := x"FCBB";
          m(232) := x"FBDC";
          m(233) := x"FD87";
          m(234) := x"FC6A";
          m(235) := x"F4AB";
          m(236) := x"F38B";
          m(237) := x"FC84";
          m(238) := x"F7FE";
          m(239) := x"F447";
          m(240) := x"00B0";
          m(241) := x"FFCC";
          m(242) := x"F638";
          m(243) := x"FCFA";
          m(244) := x"F929";
          m(245) := x"FCE2";
          m(246) := x"FEE4";
          m(247) := x"0160";
          m(248) := x"02AA";
          m(249) := x"0117";
          m(250) := x"FFF4";
          m(251) := x"FFF3";
          m(252) := x"001E";
          m(253) := x"FFBD";
          m(254) := x"FFCB";
          m(255) := x"FE55";
          m(256) := x"FF9D";
          m(257) := x"016D";
          m(258) := x"029B";
          m(259) := x"01EF";
          m(260) := x"0161";
          m(261) := x"031D";
          m(262) := x"03B7";
          m(263) := x"FD2D";
          m(264) := x"F787";
          m(265) := x"FB43";
          m(266) := x"F5A3";
          m(267) := x"F1F4";
          m(268) := x"FD4F";
          m(269) := x"F7CC";
          m(270) := x"F4FE";
          m(271) := x"FB3A";
          m(272) := x"F8FD";
          m(273) := x"FF9A";
          m(274) := x"FDD8";
          m(275) := x"0143";
          m(276) := x"01E5";
          m(277) := x"0039";
          m(278) := x"0028";
          m(279) := x"FFF5";
          m(280) := x"0019";
          m(281) := x"0020";
          m(282) := x"FFAF";
          m(283) := x"FF5C";
          m(284) := x"02CE";
          m(285) := x"049C";
          m(286) := x"05E0";
          m(287) := x"084F";
          m(288) := x"06AD";
          m(289) := x"0A1D";
          m(290) := x"079C";
          m(291) := x"019F";
          m(292) := x"012D";
          m(293) := x"026D";
          m(294) := x"FA53";
          m(295) := x"F353";
          m(296) := x"FA6C";
          m(297) := x"FB36";
          m(298) := x"FEED";
          m(299) := x"0116";
          m(300) := x"FE0D";
          m(301) := x"FE44";
          m(302) := x"FBE6";
          m(303) := x"015B";
          m(304) := x"016E";
          m(305) := x"FF2E";
          m(306) := x"001B";
          m(307) := x"0036";
          m(308) := x"FFF6";
          m(309) := x"0016";
          m(310) := x"FFF0";
          m(311) := x"0082";
          m(312) := x"055B";
          m(313) := x"0849";
          m(314) := x"087E";
          m(315) := x"095F";
          m(316) := x"0879";
          m(317) := x"08F7";
          m(318) := x"0947";
          m(319) := x"06D9";
          m(320) := x"07A3";
          m(321) := x"0C0B";
          m(322) := x"09DF";
          m(323) := x"01EC";
          m(324) := x"03DA";
          m(325) := x"FEA0";
          m(326) := x"FEFB";
          m(327) := x"0178";
          m(328) := x"FEA8";
          m(329) := x"017A";
          m(330) := x"FDD5";
          m(331) := x"020A";
          m(332) := x"FFF8";
          m(333) := x"FF00";
          m(334) := x"FF8D";
          m(335) := x"FFFD";
          m(336) := x"0045";
          m(337) := x"FFDB";
          m(338) := x"000C";
          m(339) := x"01DA";
          m(340) := x"060C";
          m(341) := x"0753";
          m(342) := x"06A7";
          m(343) := x"075C";
          m(344) := x"06A8";
          m(345) := x"097E";
          m(346) := x"0784";
          m(347) := x"0848";
          m(348) := x"0101";
          m(349) := x"0362";
          m(350) := x"0E9F";
          m(351) := x"04FC";
          m(352) := x"0099";
          m(353) := x"0347";
          m(354) := x"FD7B";
          m(355) := x"FE71";
          m(356) := x"FE5F";
          m(357) := x"00AB";
          m(358) := x"FF8E";
          m(359) := x"0695";
          m(360) := x"FFC2";
          m(361) := x"FEF6";
          m(362) := x"0015";
          m(363) := x"FFF1";
          m(364) := x"0035";
          m(365) := x"FFDA";
          m(366) := x"FFA1";
          m(367) := x"0173";
          m(368) := x"03EB";
          m(369) := x"02AA";
          m(370) := x"0630";
          m(371) := x"030F";
          m(372) := x"FE64";
          m(373) := x"0248";
          m(374) := x"0107";
          m(375) := x"020E";
          m(376) := x"007E";
          m(377) := x"022F";
          m(378) := x"08C5";
          m(379) := x"03F1";
          m(380) := x"0084";
          m(381) := x"FF5F";
          m(382) := x"FE1A";
          m(383) := x"FFC5";
          m(384) := x"00EC";
          m(385) := x"0009";
          m(386) := x"047E";
          m(387) := x"072F";
          m(388) := x"00A7";
          m(389) := x"FF2B";
          m(390) := x"0018";
          m(391) := x"FFEE";
          m(392) := x"FFF2";
          m(393) := x"0033";
          m(394) := x"FFA6";
          m(395) := x"010C";
          m(396) := x"01F3";
          m(397) := x"FF8A";
          m(398) := x"04B9";
          m(399) := x"FCEF";
          m(400) := x"0150";
          m(401) := x"0552";
          m(402) := x"022F";
          m(403) := x"0394";
          m(404) := x"024C";
          m(405) := x"033A";
          m(406) := x"069E";
          m(407) := x"0554";
          m(408) := x"0539";
          m(409) := x"009A";
          m(410) := x"03AC";
          m(411) := x"0198";
          m(412) := x"03BE";
          m(413) := x"013A";
          m(414) := x"05EC";
          m(415) := x"025A";
          m(416) := x"FFF3";
          m(417) := x"FFF1";
          m(418) := x"FFF8";
          m(419) := x"0038";
          m(420) := x"FFDC";
          m(421) := x"001A";
          m(422) := x"FF89";
          m(423) := x"010D";
          m(424) := x"FE7D";
          m(425) := x"FEBB";
          m(426) := x"024A";
          m(427) := x"015C";
          m(428) := x"04A6";
          m(429) := x"0157";
          m(430) := x"0082";
          m(431) := x"06C0";
          m(432) := x"0639";
          m(433) := x"0650";
          m(434) := x"0454";
          m(435) := x"FE31";
          m(436) := x"FD45";
          m(437) := x"0043";
          m(438) := x"0246";
          m(439) := x"0565";
          m(440) := x"013C";
          m(441) := x"FE23";
          m(442) := x"FF2A";
          m(443) := x"0160";
          m(444) := x"0067";
          m(445) := x"FFB7";
          m(446) := x"FF89";
          m(447) := x"0003";
          m(448) := x"0037";
          m(449) := x"FFDB";
          m(450) := x"FFC5";
          m(451) := x"FF95";
          m(452) := x"FD63";
          m(453) := x"00EF";
          m(454) := x"041B";
          m(455) := x"0165";
          m(456) := x"04C1";
          m(457) := x"FFCB";
          m(458) := x"FD74";
          m(459) := x"0485";
          m(460) := x"049C";
          m(461) := x"0673";
          m(462) := x"014F";
          m(463) := x"0128";
          m(464) := x"0250";
          m(465) := x"023D";
          m(466) := x"0154";
          m(467) := x"0174";
          m(468) := x"FDE2";
          m(469) := x"FCD2";
          m(470) := x"FF2F";
          m(471) := x"0214";
          m(472) := x"001D";
          m(473) := x"0061";
          m(474) := x"0005";
          m(475) := x"0023";
          m(476) := x"0023";
          m(477) := x"FFE7";
          m(478) := x"FFC7";
          m(479) := x"FE34";
          m(480) := x"FCA1";
          m(481) := x"018F";
          m(482) := x"0325";
          m(483) := x"FF74";
          m(484) := x"055B";
          m(485) := x"00F5";
          m(486) := x"0520";
          m(487) := x"064D";
          m(488) := x"052B";
          m(489) := x"07AC";
          m(490) := x"0647";
          m(491) := x"0586";
          m(492) := x"01D9";
          m(493) := x"FCDC";
          m(494) := x"0334";
          m(495) := x"0424";
          m(496) := x"0383";
          m(497) := x"FE95";
          m(498) := x"02E0";
          m(499) := x"030B";
          m(500) := x"FF09";
          m(501) := x"FF11";
          m(502) := x"FFA7";
          m(503) := x"0018";
          m(504) := x"000B";
          m(505) := x"FFF8";
          m(506) := x"0012";
          m(507) := x"FEDD";
          m(508) := x"FE4C";
          m(509) := x"01F9";
          m(510) := x"0226";
          m(511) := x"FE94";
          m(512) := x"00F5";
          m(513) := x"04EE";
          m(514) := x"0030";
          m(515) := x"032E";
          m(516) := x"0535";
          m(517) := x"0742";
          m(518) := x"02FF";
          m(519) := x"FE2A";
          m(520) := x"FB20";
          m(521) := x"FF24";
          m(522) := x"FFFB";
          m(523) := x"02FE";
          m(524) := x"06DF";
          m(525) := x"00EE";
          m(526) := x"013E";
          m(527) := x"0174";
          m(528) := x"0024";
          m(529) := x"FF67";
          m(530) := x"FF63";
          m(531) := x"005C";
          m(532) := x"000C";
          m(533) := x"FFE1";
          m(534) := x"FFC2";
          m(535) := x"FF97";
          m(536) := x"00EE";
          m(537) := x"0056";
          m(538) := x"FE4B";
          m(539) := x"FF15";
          m(540) := x"01BD";
          m(541) := x"0433";
          m(542) := x"FCCB";
          m(543) := x"04E4";
          m(544) := x"FC72";
          m(545) := x"03A3";
          m(546) := x"FF12";
          m(547) := x"023B";
          m(548) := x"FE30";
          m(549) := x"FCAE";
          m(550) := x"FDCA";
          m(551) := x"00FF";
          m(552) := x"0099";
          m(553) := x"006F";
          m(554) := x"FF7F";
          m(555) := x"0157";
          m(556) := x"01B7";
          m(557) := x"0030";
          m(558) := x"0073";
          m(559) := x"002B";
          m(560) := x"0022";
          m(561) := x"FFC1";
          m(562) := x"000F";
          m(563) := x"FE9B";
          m(564) := x"0161";
          m(565) := x"FEA7";
          m(566) := x"FD1E";
          m(567) := x"F9F5";
          m(568) := x"FD44";
          m(569) := x"FFF4";
          m(570) := x"FDA8";
          m(571) := x"00D9";
          m(572) := x"015F";
          m(573) := x"FC0B";
          m(574) := x"0370";
          m(575) := x"FFDA";
          m(576) := x"F946";
          m(577) := x"FEAC";
          m(578) := x"FE24";
          m(579) := x"FD0C";
          m(580) := x"0159";
          m(581) := x"FEFE";
          m(582) := x"FFFF";
          m(583) := x"010C";
          m(584) := x"013E";
          m(585) := x"003D";
          m(586) := x"0046";
          m(587) := x"FFF5";
          m(588) := x"0007";
          m(589) := x"000C";
          m(590) := x"FFE2";
          m(591) := x"FF47";
          m(592) := x"0068";
          m(593) := x"0074";
          m(594) := x"FCF2";
          m(595) := x"F974";
          m(596) := x"F835";
          m(597) := x"FC88";
          m(598) := x"FD3B";
          m(599) := x"FD43";
          m(600) := x"FB25";
          m(601) := x"FE30";
          m(602) := x"0223";
          m(603) := x"FCAE";
          m(604) := x"FD6D";
          m(605) := x"FE12";
          m(606) := x"FEFE";
          m(607) := x"FD03";
          m(608) := x"FEC5";
          m(609) := x"004D";
          m(610) := x"004E";
          m(611) := x"011D";
          m(612) := x"00ED";
          m(613) := x"0051";
          m(614) := x"FFEF";
          m(615) := x"0000";
          m(616) := x"0016";
          m(617) := x"003C";
          m(618) := x"000B";
          m(619) := x"FF93";
          m(620) := x"00AE";
          m(621) := x"FEEC";
          m(622) := x"FABF";
          m(623) := x"F929";
          m(624) := x"F7F6";
          m(625) := x"FB8E";
          m(626) := x"FFA9";
          m(627) := x"0280";
          m(628) := x"FE15";
          m(629) := x"001B";
          m(630) := x"FDE3";
          m(631) := x"FE24";
          m(632) := x"01E4";
          m(633) := x"FE02";
          m(634) := x"0380";
          m(635) := x"00E9";
          m(636) := x"0332";
          m(637) := x"00DB";
          m(638) := x"FFB9";
          m(639) := x"01AA";
          m(640) := x"FFFE";
          m(641) := x"003D";
          m(642) := x"FFF7";
          m(643) := x"000E";
          m(644) := x"FFFF";
          m(645) := x"FFBE";
          m(646) := x"0039";
          m(647) := x"FFD4";
          m(648) := x"FFBC";
          m(649) := x"0022";
          m(650) := x"FDE2";
          m(651) := x"FC78";
          m(652) := x"0195";
          m(653) := x"0339";
          m(654) := x"FE43";
          m(655) := x"F6C4";
          m(656) := x"FD82";
          m(657) := x"FE8B";
          m(658) := x"0020";
          m(659) := x"0039";
          m(660) := x"FDDE";
          m(661) := x"0207";
          m(662) := x"03E4";
          m(663) := x"0379";
          m(664) := x"0452";
          m(665) := x"FFEF";
          m(666) := x"01C7";
          m(667) := x"0166";
          m(668) := x"FFE9";
          m(669) := x"FFEE";
          m(670) := x"004A";
          m(671) := x"FFE7";
          m(672) := x"0000";
          m(673) := x"000C";
          m(674) := x"FFF1";
          m(675) := x"FFD2";
          m(676) := x"FF13";
          m(677) := x"FCFC";
          m(678) := x"FD2C";
          m(679) := x"FD7B";
          m(680) := x"FFF2";
          m(681) := x"0567";
          m(682) := x"042D";
          m(683) := x"0024";
          m(684) := x"01CB";
          m(685) := x"FD04";
          m(686) := x"FEEB";
          m(687) := x"FFBA";
          m(688) := x"0158";
          m(689) := x"FFB7";
          m(690) := x"007C";
          m(691) := x"0554";
          m(692) := x"03BA";
          m(693) := x"0212";
          m(694) := x"01D6";
          m(695) := x"012C";
          m(696) := x"0057";
          m(697) := x"FFF1";
          m(698) := x"FFE7";
          m(699) := x"000B";
          m(700) := x"FFEA";
          m(701) := x"FFD6";
          m(702) := x"0004";
          m(703) := x"FFF6";
          m(704) := x"FF1A";
          m(705) := x"FEE8";
          m(706) := x"FF4B";
          m(707) := x"FF4F";
          m(708) := x"FD31";
          m(709) := x"FBAF";
          m(710) := x"FB24";
          m(711) := x"FE34";
          m(712) := x"FEE8";
          m(713) := x"004A";
          m(714) := x"00F6";
          m(715) := x"FE4B";
          m(716) := x"00A2";
          m(717) := x"FFCC";
          m(718) := x"FE4D";
          m(719) := x"0005";
          m(720) := x"024F";
          m(721) := x"023C";
          m(722) := x"00F5";
          m(723) := x"FFFB";
          m(724) := x"0014";
          m(725) := x"003E";
          m(726) := x"FFB1";
          m(727) := x"0009";
          m(728) := x"FFEE";
          m(729) := x"FFE2";
          m(730) := x"0005";
          m(731) := x"FFFE";
          m(732) := x"00EF";
          m(733) := x"01B0";
          m(734) := x"00FA";
          m(735) := x"FF04";
          m(736) := x"FC8E";
          m(737) := x"FC94";
          m(738) := x"FC84";
          m(739) := x"FF59";
          m(740) := x"00FD";
          m(741) := x"005B";
          m(742) := x"0078";
          m(743) := x"FFEF";
          m(744) := x"FE4E";
          m(745) := x"FFA8";
          m(746) := x"FDF6";
          m(747) := x"FF42";
          m(748) := x"0033";
          m(749) := x"009B";
          m(750) := x"007A";
          m(751) := x"000E";
          m(752) := x"FFE5";
          m(753) := x"FFF8";
          m(754) := x"0027";
          m(755) := x"0046";
          m(756) := x"0003";
          m(757) := x"0011";
          m(758) := x"FFFC";
          m(759) := x"001D";
          m(760) := x"FFD0";
          m(761) := x"FFD8";
          m(762) := x"0051";
          m(763) := x"FFF8";
          m(764) := x"0034";
          m(765) := x"FFB3";
          m(766) := x"FFEC";
          m(767) := x"0031";
          m(768) := x"0032";
          m(769) := x"FFE3";
          m(770) := x"FFDF";
          m(771) := x"FFE6";
          m(772) := x"FF7A";
          m(773) := x"FFC7";
          m(774) := x"FF80";
          m(775) := x"FFC0";
          m(776) := x"FFF5";
          m(777) := x"000E";
          m(778) := x"0052";
          m(779) := x"0000";
          m(780) := x"FFDF";
          m(781) := x"0004";
          m(782) := x"FFE7";
          m(783) := x"FFF8";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_1_29.mif
-- Expected length: 784, input: 784, padded: 0, trimmed: 0
        if (lno = 1) and (nno = 29) then
          m(0) := x"0027";
          m(1) := x"0019";
          m(2) := x"001F";
          m(3) := x"FFF1";
          m(4) := x"FFF4";
          m(5) := x"FFE7";
          m(6) := x"FFF1";
          m(7) := x"FFF9";
          m(8) := x"000B";
          m(9) := x"000A";
          m(10) := x"0022";
          m(11) := x"FFF8";
          m(12) := x"FFE4";
          m(13) := x"FFDE";
          m(14) := x"0027";
          m(15) := x"FFB4";
          m(16) := x"FFFA";
          m(17) := x"FFF9";
          m(18) := x"FFE4";
          m(19) := x"FFF8";
          m(20) := x"000D";
          m(21) := x"FFC8";
          m(22) := x"0001";
          m(23) := x"FFEE";
          m(24) := x"0007";
          m(25) := x"FFE7";
          m(26) := x"000C";
          m(27) := x"FFE3";
          m(28) := x"FFFA";
          m(29) := x"0018";
          m(30) := x"0010";
          m(31) := x"0016";
          m(32) := x"FFF9";
          m(33) := x"002D";
          m(34) := x"0002";
          m(35) := x"0002";
          m(36) := x"FFD7";
          m(37) := x"FFD3";
          m(38) := x"FFDC";
          m(39) := x"0087";
          m(40) := x"004C";
          m(41) := x"0032";
          m(42) := x"FFEF";
          m(43) := x"0005";
          m(44) := x"0015";
          m(45) := x"0007";
          m(46) := x"FFEE";
          m(47) := x"FFFC";
          m(48) := x"0039";
          m(49) := x"0031";
          m(50) := x"0001";
          m(51) := x"000C";
          m(52) := x"FFEE";
          m(53) := x"FFDA";
          m(54) := x"001B";
          m(55) := x"0018";
          m(56) := x"000D";
          m(57) := x"FFD8";
          m(58) := x"001C";
          m(59) := x"FFF6";
          m(60) := x"FFF7";
          m(61) := x"FFFB";
          m(62) := x"FFA6";
          m(63) := x"FFCA";
          m(64) := x"0004";
          m(65) := x"FFD7";
          m(66) := x"FFD7";
          m(67) := x"FF90";
          m(68) := x"FFE9";
          m(69) := x"FFA2";
          m(70) := x"FFA6";
          m(71) := x"FF65";
          m(72) := x"FF04";
          m(73) := x"FF97";
          m(74) := x"FFAF";
          m(75) := x"FFE9";
          m(76) := x"FF57";
          m(77) := x"000B";
          m(78) := x"FFE4";
          m(79) := x"000B";
          m(80) := x"FFFB";
          m(81) := x"FFDD";
          m(82) := x"FFF5";
          m(83) := x"FFEB";
          m(84) := x"FFCF";
          m(85) := x"FFB9";
          m(86) := x"FFCE";
          m(87) := x"0077";
          m(88) := x"0014";
          m(89) := x"FF93";
          m(90) := x"FFB3";
          m(91) := x"00A9";
          m(92) := x"0062";
          m(93) := x"FF84";
          m(94) := x"FF60";
          m(95) := x"FEAB";
          m(96) := x"FDA2";
          m(97) := x"FEE7";
          m(98) := x"027A";
          m(99) := x"01A7";
          m(100) := x"0094";
          m(101) := x"FCAE";
          m(102) := x"FAAB";
          m(103) := x"FDCB";
          m(104) := x"012F";
          m(105) := x"FEFE";
          m(106) := x"0014";
          m(107) := x"0119";
          m(108) := x"0044";
          m(109) := x"FF13";
          m(110) := x"FFD5";
          m(111) := x"0007";
          m(112) := x"FFE9";
          m(113) := x"0005";
          m(114) := x"0035";
          m(115) := x"0014";
          m(116) := x"0009";
          m(117) := x"FFB1";
          m(118) := x"FFB3";
          m(119) := x"0019";
          m(120) := x"002D";
          m(121) := x"FEA6";
          m(122) := x"FDE6";
          m(123) := x"FF9E";
          m(124) := x"FC3B";
          m(125) := x"FE58";
          m(126) := x"0017";
          m(127) := x"FF24";
          m(128) := x"00A9";
          m(129) := x"044A";
          m(130) := x"018D";
          m(131) := x"FD1A";
          m(132) := x"FF15";
          m(133) := x"FD6A";
          m(134) := x"009B";
          m(135) := x"01AC";
          m(136) := x"FEE5";
          m(137) := x"FEFB";
          m(138) := x"FF65";
          m(139) := x"001E";
          m(140) := x"000D";
          m(141) := x"0040";
          m(142) := x"FFF0";
          m(143) := x"FFD8";
          m(144) := x"0099";
          m(145) := x"0034";
          m(146) := x"002E";
          m(147) := x"0088";
          m(148) := x"005D";
          m(149) := x"FD35";
          m(150) := x"FDF3";
          m(151) := x"00AD";
          m(152) := x"0085";
          m(153) := x"02E8";
          m(154) := x"FE98";
          m(155) := x"FE98";
          m(156) := x"019D";
          m(157) := x"04AA";
          m(158) := x"049C";
          m(159) := x"0197";
          m(160) := x"FF3C";
          m(161) := x"FF9B";
          m(162) := x"FFF8";
          m(163) := x"FDB3";
          m(164) := x"FDE8";
          m(165) := x"FF03";
          m(166) := x"FFE0";
          m(167) := x"FFD9";
          m(168) := x"003B";
          m(169) := x"000C";
          m(170) := x"FFD0";
          m(171) := x"0007";
          m(172) := x"008D";
          m(173) := x"FF6F";
          m(174) := x"FFAF";
          m(175) := x"0043";
          m(176) := x"FDBE";
          m(177) := x"F8F0";
          m(178) := x"FEAD";
          m(179) := x"FDE3";
          m(180) := x"FE1B";
          m(181) := x"0264";
          m(182) := x"01D2";
          m(183) := x"FE61";
          m(184) := x"FEEA";
          m(185) := x"02A4";
          m(186) := x"015C";
          m(187) := x"02B6";
          m(188) := x"029D";
          m(189) := x"0222";
          m(190) := x"0149";
          m(191) := x"FCD5";
          m(192) := x"FB60";
          m(193) := x"FD84";
          m(194) := x"FF2F";
          m(195) := x"FF75";
          m(196) := x"FFF1";
          m(197) := x"FFE4";
          m(198) := x"0002";
          m(199) := x"0020";
          m(200) := x"006B";
          m(201) := x"002E";
          m(202) := x"0192";
          m(203) := x"01B9";
          m(204) := x"F850";
          m(205) := x"FC13";
          m(206) := x"0183";
          m(207) := x"0046";
          m(208) := x"018D";
          m(209) := x"02E2";
          m(210) := x"FFDF";
          m(211) := x"006E";
          m(212) := x"00D9";
          m(213) := x"01C4";
          m(214) := x"06E4";
          m(215) := x"0885";
          m(216) := x"0254";
          m(217) := x"0172";
          m(218) := x"0090";
          m(219) := x"0225";
          m(220) := x"0291";
          m(221) := x"0194";
          m(222) := x"FF67";
          m(223) := x"FFEC";
          m(224) := x"FFFD";
          m(225) := x"0005";
          m(226) := x"0004";
          m(227) := x"0004";
          m(228) := x"FFE6";
          m(229) := x"FE2C";
          m(230) := x"FFBE";
          m(231) := x"FD05";
          m(232) := x"FAD8";
          m(233) := x"FD36";
          m(234) := x"FC45";
          m(235) := x"FEA7";
          m(236) := x"00A2";
          m(237) := x"FDF2";
          m(238) := x"00CA";
          m(239) := x"0038";
          m(240) := x"0734";
          m(241) := x"FE19";
          m(242) := x"042C";
          m(243) := x"057A";
          m(244) := x"047F";
          m(245) := x"FD6F";
          m(246) := x"FF51";
          m(247) := x"0014";
          m(248) := x"FFA7";
          m(249) := x"FDBD";
          m(250) := x"FEB3";
          m(251) := x"FFE2";
          m(252) := x"FFEF";
          m(253) := x"0007";
          m(254) := x"FFF3";
          m(255) := x"FFBA";
          m(256) := x"FF42";
          m(257) := x"FE36";
          m(258) := x"FF13";
          m(259) := x"FD94";
          m(260) := x"FD7C";
          m(261) := x"0000";
          m(262) := x"FD69";
          m(263) := x"F966";
          m(264) := x"FC49";
          m(265) := x"0058";
          m(266) := x"FBA0";
          m(267) := x"FD04";
          m(268) := x"00EC";
          m(269) := x"FD7B";
          m(270) := x"0244";
          m(271) := x"05A7";
          m(272) := x"0B83";
          m(273) := x"FD8C";
          m(274) := x"FDB3";
          m(275) := x"0346";
          m(276) := x"FFBF";
          m(277) := x"FCF6";
          m(278) := x"FE8E";
          m(279) := x"FFDD";
          m(280) := x"0006";
          m(281) := x"FFF9";
          m(282) := x"FFCA";
          m(283) := x"FF9D";
          m(284) := x"FE94";
          m(285) := x"FEC3";
          m(286) := x"FDC5";
          m(287) := x"0141";
          m(288) := x"003A";
          m(289) := x"00BA";
          m(290) := x"FAB4";
          m(291) := x"FD2F";
          m(292) := x"035D";
          m(293) := x"FD45";
          m(294) := x"01F9";
          m(295) := x"0489";
          m(296) := x"01E4";
          m(297) := x"00DD";
          m(298) := x"006C";
          m(299) := x"01F0";
          m(300) := x"04E7";
          m(301) := x"053D";
          m(302) := x"072E";
          m(303) := x"04C1";
          m(304) := x"004E";
          m(305) := x"FD9B";
          m(306) := x"FEAA";
          m(307) := x"000D";
          m(308) := x"0016";
          m(309) := x"0003";
          m(310) := x"0011";
          m(311) := x"FF6B";
          m(312) := x"FE8A";
          m(313) := x"FD53";
          m(314) := x"02E0";
          m(315) := x"019C";
          m(316) := x"FEE1";
          m(317) := x"00B6";
          m(318) := x"FEBE";
          m(319) := x"FFC2";
          m(320) := x"FC95";
          m(321) := x"FDD3";
          m(322) := x"02C6";
          m(323) := x"FDD1";
          m(324) := x"F70B";
          m(325) := x"F538";
          m(326) := x"F795";
          m(327) := x"FE9A";
          m(328) := x"03A4";
          m(329) := x"0217";
          m(330) := x"05D1";
          m(331) := x"026F";
          m(332) := x"02DB";
          m(333) := x"FF95";
          m(334) := x"FF7B";
          m(335) := x"FFFB";
          m(336) := x"0014";
          m(337) := x"FFF8";
          m(338) := x"0013";
          m(339) := x"FFD6";
          m(340) := x"FEE7";
          m(341) := x"FFB1";
          m(342) := x"03DE";
          m(343) := x"FEDA";
          m(344) := x"FF9E";
          m(345) := x"0207";
          m(346) := x"0009";
          m(347) := x"FF98";
          m(348) := x"FF21";
          m(349) := x"03A4";
          m(350) := x"0079";
          m(351) := x"FBA4";
          m(352) := x"F792";
          m(353) := x"F7C8";
          m(354) := x"FC78";
          m(355) := x"0277";
          m(356) := x"00D5";
          m(357) := x"FDF0";
          m(358) := x"03BC";
          m(359) := x"04A9";
          m(360) := x"04F4";
          m(361) := x"00F6";
          m(362) := x"FFF1";
          m(363) := x"FFDF";
          m(364) := x"0022";
          m(365) := x"FFF5";
          m(366) := x"0010";
          m(367) := x"FF30";
          m(368) := x"002E";
          m(369) := x"0046";
          m(370) := x"04AD";
          m(371) := x"0163";
          m(372) := x"029E";
          m(373) := x"0189";
          m(374) := x"0443";
          m(375) := x"FD24";
          m(376) := x"FF72";
          m(377) := x"0068";
          m(378) := x"FF92";
          m(379) := x"FB8E";
          m(380) := x"F82C";
          m(381) := x"F92A";
          m(382) := x"FDD5";
          m(383) := x"FE9B";
          m(384) := x"FBD4";
          m(385) := x"FEDD";
          m(386) := x"0284";
          m(387) := x"0527";
          m(388) := x"02EB";
          m(389) := x"0110";
          m(390) := x"0007";
          m(391) := x"FFE1";
          m(392) := x"0012";
          m(393) := x"0005";
          m(394) := x"FFCB";
          m(395) := x"FEAA";
          m(396) := x"00D3";
          m(397) := x"03E4";
          m(398) := x"03DE";
          m(399) := x"048A";
          m(400) := x"0417";
          m(401) := x"00F6";
          m(402) := x"0004";
          m(403) := x"FF61";
          m(404) := x"FE52";
          m(405) := x"00F3";
          m(406) := x"FF60";
          m(407) := x"FC56";
          m(408) := x"F885";
          m(409) := x"F845";
          m(410) := x"FD0A";
          m(411) := x"FF64";
          m(412) := x"0092";
          m(413) := x"0130";
          m(414) := x"0153";
          m(415) := x"0402";
          m(416) := x"0248";
          m(417) := x"00B2";
          m(418) := x"FFF1";
          m(419) := x"FFB5";
          m(420) := x"001A";
          m(421) := x"FFE6";
          m(422) := x"FFFD";
          m(423) := x"FDDC";
          m(424) := x"FF4B";
          m(425) := x"0486";
          m(426) := x"00E5";
          m(427) := x"03DB";
          m(428) := x"05A2";
          m(429) := x"0334";
          m(430) := x"FEC9";
          m(431) := x"F87A";
          m(432) := x"F9F7";
          m(433) := x"FE28";
          m(434) := x"FC3D";
          m(435) := x"FC59";
          m(436) := x"FAEC";
          m(437) := x"F8B0";
          m(438) := x"FE78";
          m(439) := x"FD9E";
          m(440) := x"025D";
          m(441) := x"FF6C";
          m(442) := x"011B";
          m(443) := x"03E0";
          m(444) := x"00AD";
          m(445) := x"FF58";
          m(446) := x"FFD7";
          m(447) := x"FFF5";
          m(448) := x"FFEF";
          m(449) := x"000A";
          m(450) := x"000D";
          m(451) := x"FDA7";
          m(452) := x"FF99";
          m(453) := x"06F3";
          m(454) := x"01B6";
          m(455) := x"0399";
          m(456) := x"0363";
          m(457) := x"0358";
          m(458) := x"FB67";
          m(459) := x"F6C7";
          m(460) := x"F6CB";
          m(461) := x"F8D2";
          m(462) := x"FE21";
          m(463) := x"FB01";
          m(464) := x"F98A";
          m(465) := x"FE96";
          m(466) := x"FCD0";
          m(467) := x"FDF3";
          m(468) := x"0281";
          m(469) := x"FEAA";
          m(470) := x"FFBA";
          m(471) := x"0014";
          m(472) := x"FE0A";
          m(473) := x"FEC0";
          m(474) := x"FF95";
          m(475) := x"FFF2";
          m(476) := x"0019";
          m(477) := x"0019";
          m(478) := x"003E";
          m(479) := x"FE27";
          m(480) := x"FF34";
          m(481) := x"0588";
          m(482) := x"0196";
          m(483) := x"0276";
          m(484) := x"0331";
          m(485) := x"039E";
          m(486) := x"FFC1";
          m(487) := x"F752";
          m(488) := x"FA5C";
          m(489) := x"FE53";
          m(490) := x"0028";
          m(491) := x"FBFB";
          m(492) := x"FA6B";
          m(493) := x"FCF2";
          m(494) := x"FB49";
          m(495) := x"FF46";
          m(496) := x"00ED";
          m(497) := x"FBD2";
          m(498) := x"0179";
          m(499) := x"0015";
          m(500) := x"FF03";
          m(501) := x"FD91";
          m(502) := x"FFE5";
          m(503) := x"0044";
          m(504) := x"0013";
          m(505) := x"0025";
          m(506) := x"0015";
          m(507) := x"FDFE";
          m(508) := x"01FD";
          m(509) := x"0166";
          m(510) := x"00B2";
          m(511) := x"FD75";
          m(512) := x"0682";
          m(513) := x"0856";
          m(514) := x"0146";
          m(515) := x"F84E";
          m(516) := x"FAAB";
          m(517) := x"FD19";
          m(518) := x"01C1";
          m(519) := x"00E8";
          m(520) := x"00EE";
          m(521) := x"FED6";
          m(522) := x"FEFC";
          m(523) := x"FE3E";
          m(524) := x"FE35";
          m(525) := x"FF36";
          m(526) := x"051B";
          m(527) := x"005F";
          m(528) := x"FCA9";
          m(529) := x"FD96";
          m(530) := x"FFF8";
          m(531) := x"FFD9";
          m(532) := x"FFC2";
          m(533) := x"0035";
          m(534) := x"0021";
          m(535) := x"FE01";
          m(536) := x"FFD3";
          m(537) := x"FD3C";
          m(538) := x"FF0B";
          m(539) := x"000B";
          m(540) := x"059B";
          m(541) := x"05BA";
          m(542) := x"FD65";
          m(543) := x"F7A2";
          m(544) := x"FF2A";
          m(545) := x"FE34";
          m(546) := x"0159";
          m(547) := x"FC51";
          m(548) := x"FEB8";
          m(549) := x"FF2E";
          m(550) := x"FFE6";
          m(551) := x"FD60";
          m(552) := x"0067";
          m(553) := x"036B";
          m(554) := x"04D4";
          m(555) := x"FE39";
          m(556) := x"FCBB";
          m(557) := x"FD24";
          m(558) := x"FFD1";
          m(559) := x"FFE7";
          m(560) := x"004C";
          m(561) := x"003B";
          m(562) := x"FFD8";
          m(563) := x"FF63";
          m(564) := x"00C0";
          m(565) := x"FCAE";
          m(566) := x"FCA0";
          m(567) := x"0414";
          m(568) := x"0510";
          m(569) := x"034A";
          m(570) := x"07D9";
          m(571) := x"FE0E";
          m(572) := x"FFAD";
          m(573) := x"0160";
          m(574) := x"FAE7";
          m(575) := x"FDC3";
          m(576) := x"FD95";
          m(577) := x"FE20";
          m(578) := x"FF29";
          m(579) := x"FF05";
          m(580) := x"FE5C";
          m(581) := x"FF65";
          m(582) := x"FD92";
          m(583) := x"FBB2";
          m(584) := x"FC68";
          m(585) := x"FE06";
          m(586) := x"000F";
          m(587) := x"0012";
          m(588) := x"0018";
          m(589) := x"FFDF";
          m(590) := x"FF62";
          m(591) := x"0020";
          m(592) := x"0084";
          m(593) := x"FEB2";
          m(594) := x"00B5";
          m(595) := x"036F";
          m(596) := x"0158";
          m(597) := x"03DE";
          m(598) := x"0685";
          m(599) := x"FF71";
          m(600) := x"FDE4";
          m(601) := x"FD53";
          m(602) := x"FBB5";
          m(603) := x"FFF1";
          m(604) := x"FE70";
          m(605) := x"FAEA";
          m(606) := x"FAF1";
          m(607) := x"FBB6";
          m(608) := x"FF6F";
          m(609) := x"FE8F";
          m(610) := x"0002";
          m(611) := x"FDE0";
          m(612) := x"FD4F";
          m(613) := x"FF42";
          m(614) := x"0001";
          m(615) := x"FFC5";
          m(616) := x"FFF6";
          m(617) := x"FFDE";
          m(618) := x"FFF8";
          m(619) := x"FF9C";
          m(620) := x"FF03";
          m(621) := x"00FD";
          m(622) := x"0163";
          m(623) := x"0060";
          m(624) := x"04CD";
          m(625) := x"04F3";
          m(626) := x"03B1";
          m(627) := x"00AD";
          m(628) := x"FF75";
          m(629) := x"FEA0";
          m(630) := x"FDE8";
          m(631) := x"FDC3";
          m(632) := x"FDB6";
          m(633) := x"FFE0";
          m(634) := x"FE78";
          m(635) := x"0029";
          m(636) := x"FDA2";
          m(637) := x"0027";
          m(638) := x"0050";
          m(639) := x"FF66";
          m(640) := x"FF54";
          m(641) := x"FFA4";
          m(642) := x"0003";
          m(643) := x"FFE3";
          m(644) := x"001E";
          m(645) := x"FFF4";
          m(646) := x"FFE8";
          m(647) := x"FFC5";
          m(648) := x"FF62";
          m(649) := x"011E";
          m(650) := x"03B2";
          m(651) := x"03E5";
          m(652) := x"0390";
          m(653) := x"056E";
          m(654) := x"0697";
          m(655) := x"0265";
          m(656) := x"00A6";
          m(657) := x"FFF1";
          m(658) := x"FCCC";
          m(659) := x"FE02";
          m(660) := x"FFEC";
          m(661) := x"FF83";
          m(662) := x"F998";
          m(663) := x"FB75";
          m(664) := x"FBEC";
          m(665) := x"FDDA";
          m(666) := x"FE8F";
          m(667) := x"FECC";
          m(668) := x"FFEE";
          m(669) := x"FFD7";
          m(670) := x"FFFA";
          m(671) := x"001B";
          m(672) := x"000F";
          m(673) := x"0004";
          m(674) := x"FFDC";
          m(675) := x"0020";
          m(676) := x"0097";
          m(677) := x"027A";
          m(678) := x"01A2";
          m(679) := x"0017";
          m(680) := x"FFCD";
          m(681) := x"01EE";
          m(682) := x"04BE";
          m(683) := x"01A6";
          m(684) := x"015E";
          m(685) := x"FE52";
          m(686) := x"FC5A";
          m(687) := x"FE67";
          m(688) := x"FE3E";
          m(689) := x"FF14";
          m(690) := x"FF63";
          m(691) := x"FE66";
          m(692) := x"FD40";
          m(693) := x"FD9A";
          m(694) := x"FF1D";
          m(695) := x"FF4B";
          m(696) := x"FFBF";
          m(697) := x"0019";
          m(698) := x"FFC2";
          m(699) := x"001E";
          m(700) := x"FFF3";
          m(701) := x"FFE6";
          m(702) := x"0053";
          m(703) := x"002E";
          m(704) := x"002D";
          m(705) := x"007B";
          m(706) := x"FFDF";
          m(707) := x"0101";
          m(708) := x"002A";
          m(709) := x"FFD3";
          m(710) := x"FDB9";
          m(711) := x"FDE5";
          m(712) := x"FD1C";
          m(713) := x"FE16";
          m(714) := x"FE43";
          m(715) := x"FE04";
          m(716) := x"FE5C";
          m(717) := x"FE0D";
          m(718) := x"FDFC";
          m(719) := x"FEC8";
          m(720) := x"FEE1";
          m(721) := x"FEBC";
          m(722) := x"FF12";
          m(723) := x"FF7C";
          m(724) := x"FF97";
          m(725) := x"000A";
          m(726) := x"000D";
          m(727) := x"0017";
          m(728) := x"FFF4";
          m(729) := x"0037";
          m(730) := x"0028";
          m(731) := x"FFF4";
          m(732) := x"0034";
          m(733) := x"0009";
          m(734) := x"0035";
          m(735) := x"008F";
          m(736) := x"007A";
          m(737) := x"0060";
          m(738) := x"0026";
          m(739) := x"FFE0";
          m(740) := x"FFA6";
          m(741) := x"FF79";
          m(742) := x"FF62";
          m(743) := x"FFF0";
          m(744) := x"FFFC";
          m(745) := x"FF5E";
          m(746) := x"FF91";
          m(747) := x"FFED";
          m(748) := x"FFB4";
          m(749) := x"FF4D";
          m(750) := x"FFC9";
          m(751) := x"003E";
          m(752) := x"0008";
          m(753) := x"FFC2";
          m(754) := x"0006";
          m(755) := x"0036";
          m(756) := x"FFFB";
          m(757) := x"FFFA";
          m(758) := x"0013";
          m(759) := x"0005";
          m(760) := x"0008";
          m(761) := x"FFBF";
          m(762) := x"0009";
          m(763) := x"FFEF";
          m(764) := x"FFED";
          m(765) := x"FFEE";
          m(766) := x"FFEA";
          m(767) := x"0026";
          m(768) := x"FFF3";
          m(769) := x"FFDA";
          m(770) := x"FFFA";
          m(771) := x"FFE9";
          m(772) := x"FFED";
          m(773) := x"FFF3";
          m(774) := x"FFDA";
          m(775) := x"0000";
          m(776) := x"0036";
          m(777) := x"000D";
          m(778) := x"FFB0";
          m(779) := x"FFD4";
          m(780) := x"0024";
          m(781) := x"000E";
          m(782) := x"001E";
          m(783) := x"0003";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_0.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 0) then
          m(0) := x"ECAB";
          m(1) := x"0863";
          m(2) := x"1612";
          m(3) := x"13D7";
          m(4) := x"12E6";
          m(5) := x"F683";
          m(6) := x"031F";
          m(7) := x"F20A";
          m(8) := x"E8C1";
          m(9) := x"FBA8";
          m(10) := x"EC7C";
          m(11) := x"F400";
          m(12) := x"0D58";
          m(13) := x"FB5B";
          m(14) := x"12C3";
          m(15) := x"1209";
          m(16) := x"F6C4";
          m(17) := x"FFEA";
          m(18) := x"F752";
          m(19) := x"EE23";
          m(20) := x"0C13";
          m(21) := x"0A4B";
          m(22) := x"F583";
          m(23) := x"1C76";
          m(24) := x"0070";
          m(25) := x"EE1A";
          m(26) := x"0670";
          m(27) := x"006E";
          m(28) := x"F9EB";
          m(29) := x"0D34";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_1.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 1) then
          m(0) := x"F89A";
          m(1) := x"F94C";
          m(2) := x"04D0";
          m(3) := x"119D";
          m(4) := x"04FD";
          m(5) := x"046D";
          m(6) := x"F77D";
          m(7) := x"0451";
          m(8) := x"EF88";
          m(9) := x"F3B8";
          m(10) := x"E9CE";
          m(11) := x"0010";
          m(12) := x"FFA0";
          m(13) := x"01AB";
          m(14) := x"117E";
          m(15) := x"0381";
          m(16) := x"F544";
          m(17) := x"FDDA";
          m(18) := x"FD0B";
          m(19) := x"F4BC";
          m(20) := x"FCC2";
          m(21) := x"129D";
          m(22) := x"FA04";
          m(23) := x"0560";
          m(24) := x"FD7E";
          m(25) := x"FA5C";
          m(26) := x"FED6";
          m(27) := x"0202";
          m(28) := x"015D";
          m(29) := x"095D";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_2.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 2) then
          m(0) := x"0353";
          m(1) := x"15DE";
          m(2) := x"FB9C";
          m(3) := x"E3F1";
          m(4) := x"F904";
          m(5) := x"F3E1";
          m(6) := x"1120";
          m(7) := x"F440";
          m(8) := x"0FAD";
          m(9) := x"0EC7";
          m(10) := x"202B";
          m(11) := x"0672";
          m(12) := x"00BA";
          m(13) := x"FEBC";
          m(14) := x"E25C";
          m(15) := x"01E8";
          m(16) := x"145F";
          m(17) := x"0B9B";
          m(18) := x"0995";
          m(19) := x"0DA5";
          m(20) := x"00AB";
          m(21) := x"DD66";
          m(22) := x"0051";
          m(23) := x"FD30";
          m(24) := x"02D9";
          m(25) := x"FC0C";
          m(26) := x"09F8";
          m(27) := x"FD64";
          m(28) := x"F772";
          m(29) := x"F3E5";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_3.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 3) then
          m(0) := x"FED1";
          m(1) := x"030F";
          m(2) := x"F2DB";
          m(3) := x"F948";
          m(4) := x"FE3A";
          m(5) := x"FB38";
          m(6) := x"03FE";
          m(7) := x"0607";
          m(8) := x"034E";
          m(9) := x"1607";
          m(10) := x"FBEE";
          m(11) := x"10DC";
          m(12) := x"0902";
          m(13) := x"0187";
          m(14) := x"F9D9";
          m(15) := x"116D";
          m(16) := x"02F5";
          m(17) := x"FB19";
          m(18) := x"027E";
          m(19) := x"0901";
          m(20) := x"08FB";
          m(21) := x"0388";
          m(22) := x"0334";
          m(23) := x"EE11";
          m(24) := x"FB32";
          m(25) := x"E725";
          m(26) := x"EC9F";
          m(27) := x"FDED";
          m(28) := x"001B";
          m(29) := x"04FF";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_4.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 4) then
          m(0) := x"FA91";
          m(1) := x"F0E7";
          m(2) := x"FDD0";
          m(3) := x"0A5A";
          m(4) := x"1B76";
          m(5) := x"DE25";
          m(6) := x"0EFE";
          m(7) := x"0042";
          m(8) := x"F2E7";
          m(9) := x"EAF8";
          m(10) := x"05B5";
          m(11) := x"F8E1";
          m(12) := x"062F";
          m(13) := x"F7D5";
          m(14) := x"F365";
          m(15) := x"1426";
          m(16) := x"0CEB";
          m(17) := x"0BDB";
          m(18) := x"0DC2";
          m(19) := x"EBB7";
          m(20) := x"FBCB";
          m(21) := x"F7F7";
          m(22) := x"EAF5";
          m(23) := x"FBEF";
          m(24) := x"087F";
          m(25) := x"F259";
          m(26) := x"0AA5";
          m(27) := x"0435";
          m(28) := x"F256";
          m(29) := x"0159";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_5.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 5) then
          m(0) := x"19EB";
          m(1) := x"FCAE";
          m(2) := x"FEBC";
          m(3) := x"0E74";
          m(4) := x"0592";
          m(5) := x"F353";
          m(6) := x"EFB0";
          m(7) := x"FFA4";
          m(8) := x"0B13";
          m(9) := x"EF15";
          m(10) := x"06C5";
          m(11) := x"F816";
          m(12) := x"E07D";
          m(13) := x"0F6A";
          m(14) := x"12B8";
          m(15) := x"E23B";
          m(16) := x"0590";
          m(17) := x"EA3B";
          m(18) := x"056B";
          m(19) := x"0AC7";
          m(20) := x"CE45";
          m(21) := x"FA88";
          m(22) := x"07F2";
          m(23) := x"005A";
          m(24) := x"05F3";
          m(25) := x"23AA";
          m(26) := x"124C";
          m(27) := x"0ED6";
          m(28) := x"F3F2";
          m(29) := x"FEEF";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_6.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 6) then
          m(0) := x"01FB";
          m(1) := x"0023";
          m(2) := x"07E5";
          m(3) := x"F267";
          m(4) := x"FFC7";
          m(5) := x"F168";
          m(6) := x"0CFD";
          m(7) := x"0744";
          m(8) := x"0DB4";
          m(9) := x"1313";
          m(10) := x"14BD";
          m(11) := x"ECA6";
          m(12) := x"E59A";
          m(13) := x"EB92";
          m(14) := x"FFF1";
          m(15) := x"EB0F";
          m(16) := x"05FE";
          m(17) := x"FC10";
          m(18) := x"03E7";
          m(19) := x"FDFE";
          m(20) := x"FC69";
          m(21) := x"F5A1";
          m(22) := x"0130";
          m(23) := x"0BE8";
          m(24) := x"024E";
          m(25) := x"0F7C";
          m(26) := x"0403";
          m(27) := x"12D0";
          m(28) := x"0128";
          m(29) := x"EF5D";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_7.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 7) then
          m(0) := x"0EFE";
          m(1) := x"016A";
          m(2) := x"F357";
          m(3) := x"00B6";
          m(4) := x"F027";
          m(5) := x"08EE";
          m(6) := x"ED86";
          m(7) := x"1758";
          m(8) := x"09FA";
          m(9) := x"089A";
          m(10) := x"EEF5";
          m(11) := x"0EEC";
          m(12) := x"E94A";
          m(13) := x"FC95";
          m(14) := x"0B36";
          m(15) := x"EB45";
          m(16) := x"F601";
          m(17) := x"FA74";
          m(18) := x"FDA4";
          m(19) := x"F28E";
          m(20) := x"EE05";
          m(21) := x"079D";
          m(22) := x"0802";
          m(23) := x"F049";
          m(24) := x"FB41";
          m(25) := x"FE32";
          m(26) := x"E9A4";
          m(27) := x"0A02";
          m(28) := x"0636";
          m(29) := x"FB1D";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_8.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 8) then
          m(0) := x"F33D";
          m(1) := x"FB6A";
          m(2) := x"0A23";
          m(3) := x"FB2A";
          m(4) := x"E4FA";
          m(5) := x"233B";
          m(6) := x"F494";
          m(7) := x"F8C7";
          m(8) := x"F6B5";
          m(9) := x"0AEA";
          m(10) := x"FD5B";
          m(11) := x"16F7";
          m(12) := x"0DB2";
          m(13) := x"0C2C";
          m(14) := x"FA5B";
          m(15) := x"FF34";
          m(16) := x"EEC7";
          m(17) := x"FC74";
          m(18) := x"FF19";
          m(19) := x"0FF2";
          m(20) := x"054F";
          m(21) := x"0E42";
          m(22) := x"0DCD";
          m(23) := x"FF2F";
          m(24) := x"F9D1";
          m(25) := x"FD7D";
          m(26) := x"F2E0";
          m(27) := x"EF46";
          m(28) := x"1904";
          m(29) := x"F1A5";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_9.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 9) then
          m(0) := x"073E";
          m(1) := x"1EEA";
          m(2) := x"0F25";
          m(3) := x"EAAD";
          m(4) := x"FD7A";
          m(5) := x"F5D7";
          m(6) := x"158E";
          m(7) := x"F26D";
          m(8) := x"08CB";
          m(9) := x"0687";
          m(10) := x"1B6B";
          m(11) := x"FB66";
          m(12) := x"FD50";
          m(13) := x"F980";
          m(14) := x"FA02";
          m(15) := x"0250";
          m(16) := x"0BE6";
          m(17) := x"077E";
          m(18) := x"FFEE";
          m(19) := x"08D5";
          m(20) := x"F59B";
          m(21) := x"DFE0";
          m(22) := x"FFE7";
          m(23) := x"17A7";
          m(24) := x"052F";
          m(25) := x"05BE";
          m(26) := x"1120";
          m(27) := x"0D68";
          m(28) := x"FEC6";
          m(29) := x"EDF6";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_10.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 10) then
          m(0) := x"F028";
          m(1) := x"0107";
          m(2) := x"F4F2";
          m(3) := x"FEDA";
          m(4) := x"0A1A";
          m(5) := x"FC1A";
          m(6) := x"FC6D";
          m(7) := x"00F5";
          m(8) := x"F79C";
          m(9) := x"F95A";
          m(10) := x"F663";
          m(11) := x"1088";
          m(12) := x"16C7";
          m(13) := x"017C";
          m(14) := x"FAD4";
          m(15) := x"197E";
          m(16) := x"0C4C";
          m(17) := x"007D";
          m(18) := x"EBE6";
          m(19) := x"F6F2";
          m(20) := x"20CC";
          m(21) := x"06E3";
          m(22) := x"F85C";
          m(23) := x"F96E";
          m(24) := x"FCAD";
          m(25) := x"F3A8";
          m(26) := x"FE2E";
          m(27) := x"E986";
          m(28) := x"F13C";
          m(29) := x"1F17";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_11.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 11) then
          m(0) := x"0189";
          m(1) := x"E518";
          m(2) := x"F8B9";
          m(3) := x"105A";
          m(4) := x"019E";
          m(5) := x"067D";
          m(6) := x"F187";
          m(7) := x"0AF6";
          m(8) := x"FA4E";
          m(9) := x"F6CA";
          m(10) := x"E9BD";
          m(11) := x"06D0";
          m(12) := x"FE3B";
          m(13) := x"FD59";
          m(14) := x"0A83";
          m(15) := x"FED6";
          m(16) := x"F4A9";
          m(17) := x"FBBA";
          m(18) := x"0935";
          m(19) := x"F89C";
          m(20) := x"F16B";
          m(21) := x"1488";
          m(22) := x"F16B";
          m(23) := x"F1EF";
          m(24) := x"FC5E";
          m(25) := x"F6DF";
          m(26) := x"EE11";
          m(27) := x"FC04";
          m(28) := x"0E50";
          m(29) := x"FE6F";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_12.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 12) then
          m(0) := x"08D6";
          m(1) := x"1511";
          m(2) := x"0650";
          m(3) := x"ED79";
          m(4) := x"FDFA";
          m(5) := x"F69A";
          m(6) := x"0AD1";
          m(7) := x"F9AA";
          m(8) := x"0685";
          m(9) := x"03E6";
          m(10) := x"1492";
          m(11) := x"F83B";
          m(12) := x"0194";
          m(13) := x"F966";
          m(14) := x"FBF9";
          m(15) := x"0121";
          m(16) := x"08B6";
          m(17) := x"0380";
          m(18) := x"FAC8";
          m(19) := x"05D1";
          m(20) := x"F22D";
          m(21) := x"E591";
          m(22) := x"FBE5";
          m(23) := x"1047";
          m(24) := x"FF3E";
          m(25) := x"0198";
          m(26) := x"059E";
          m(27) := x"0B56";
          m(28) := x"FD26";
          m(29) := x"F439";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_13.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 13) then
          m(0) := x"FDAA";
          m(1) := x"21FC";
          m(2) := x"FA28";
          m(3) := x"F92F";
          m(4) := x"EDFB";
          m(5) := x"0F16";
          m(6) := x"FDF1";
          m(7) := x"FAEA";
          m(8) := x"F9E0";
          m(9) := x"F324";
          m(10) := x"00CE";
          m(11) := x"1762";
          m(12) := x"0EA7";
          m(13) := x"F717";
          m(14) := x"F795";
          m(15) := x"0C79";
          m(16) := x"0020";
          m(17) := x"0A10";
          m(18) := x"E3B2";
          m(19) := x"0457";
          m(20) := x"111D";
          m(21) := x"FDF4";
          m(22) := x"1451";
          m(23) := x"0298";
          m(24) := x"042F";
          m(25) := x"ED4E";
          m(26) := x"09B3";
          m(27) := x"E911";
          m(28) := x"F5BA";
          m(29) := x"108B";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_14.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 14) then
          m(0) := x"F44B";
          m(1) := x"0011";
          m(2) := x"1401";
          m(3) := x"128D";
          m(4) := x"F997";
          m(5) := x"17A8";
          m(6) := x"FD02";
          m(7) := x"F0A3";
          m(8) := x"E661";
          m(9) := x"E7E5";
          m(10) := x"E594";
          m(11) := x"0024";
          m(12) := x"0AE4";
          m(13) := x"0A2A";
          m(14) := x"2470";
          m(15) := x"066E";
          m(16) := x"E8ED";
          m(17) := x"F5E0";
          m(18) := x"EC6F";
          m(19) := x"038F";
          m(20) := x"02D8";
          m(21) := x"113C";
          m(22) := x"0863";
          m(23) := x"1ED7";
          m(24) := x"F9B2";
          m(25) := x"0403";
          m(26) := x"058B";
          m(27) := x"F589";
          m(28) := x"02DC";
          m(29) := x"0169";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_15.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 15) then
          m(0) := x"FCD7";
          m(1) := x"0039";
          m(2) := x"0C3F";
          m(3) := x"0505";
          m(4) := x"F3A3";
          m(5) := x"0826";
          m(6) := x"F752";
          m(7) := x"F166";
          m(8) := x"F67F";
          m(9) := x"F132";
          m(10) := x"030D";
          m(11) := x"FAA1";
          m(12) := x"0601";
          m(13) := x"0B23";
          m(14) := x"0026";
          m(15) := x"F55B";
          m(16) := x"FB6D";
          m(17) := x"F9D6";
          m(18) := x"007C";
          m(19) := x"00E4";
          m(20) := x"E69D";
          m(21) := x"FF7E";
          m(22) := x"0092";
          m(23) := x"10E3";
          m(24) := x"FA18";
          m(25) := x"1012";
          m(26) := x"13F9";
          m(27) := x"F89A";
          m(28) := x"02BC";
          m(29) := x"0045";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_16.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 16) then
          m(0) := x"FFF7";
          m(1) := x"09F9";
          m(2) := x"066E";
          m(3) := x"FD45";
          m(4) := x"2405";
          m(5) := x"DE20";
          m(6) := x"085A";
          m(7) := x"FBCE";
          m(8) := x"FC84";
          m(9) := x"0847";
          m(10) := x"FF3A";
          m(11) := x"F092";
          m(12) := x"F0CD";
          m(13) := x"FF80";
          m(14) := x"04C8";
          m(15) := x"EB04";
          m(16) := x"1007";
          m(17) := x"05DA";
          m(18) := x"1752";
          m(19) := x"E98D";
          m(20) := x"05A4";
          m(21) := x"FDA4";
          m(22) := x"EE53";
          m(23) := x"101E";
          m(24) := x"FEB0";
          m(25) := x"08EB";
          m(26) := x"104C";
          m(27) := x"1299";
          m(28) := x"F1C5";
          m(29) := x"0AE9";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_17.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 17) then
          m(0) := x"13EF";
          m(1) := x"067D";
          m(2) := x"0310";
          m(3) := x"07BA";
          m(4) := x"0181";
          m(5) := x"FA90";
          m(6) := x"F7E8";
          m(7) := x"021D";
          m(8) := x"0AEA";
          m(9) := x"F55E";
          m(10) := x"0891";
          m(11) := x"FAA1";
          m(12) := x"F08D";
          m(13) := x"0E46";
          m(14) := x"09C7";
          m(15) := x"EB84";
          m(16) := x"04B4";
          m(17) := x"F05C";
          m(18) := x"0049";
          m(19) := x"084A";
          m(20) := x"DC19";
          m(21) := x"F68C";
          m(22) := x"0647";
          m(23) := x"079E";
          m(24) := x"FC60";
          m(25) := x"1EAE";
          m(26) := x"10DD";
          m(27) := x"07BD";
          m(28) := x"F83D";
          m(29) := x"FFCF";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_18.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 18) then
          m(0) := x"FA33";
          m(1) := x"E9B8";
          m(2) := x"0BB1";
          m(3) := x"0C26";
          m(4) := x"077C";
          m(5) := x"03EF";
          m(6) := x"F737";
          m(7) := x"F501";
          m(8) := x"FFAC";
          m(9) := x"ED23";
          m(10) := x"F909";
          m(11) := x"E8DA";
          m(12) := x"EF0B";
          m(13) := x"E927";
          m(14) := x"045B";
          m(15) := x"E639";
          m(16) := x"F015";
          m(17) := x"1053";
          m(18) := x"127D";
          m(19) := x"F6A2";
          m(20) := x"FE5B";
          m(21) := x"0EC3";
          m(22) := x"FAA1";
          m(23) := x"0855";
          m(24) := x"19E7";
          m(25) := x"1700";
          m(26) := x"0342";
          m(27) := x"0B55";
          m(28) := x"0F51";
          m(29) := x"ECE2";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_19.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 19) then
          m(0) := x"06E1";
          m(1) := x"0F56";
          m(2) := x"F197";
          m(3) := x"F798";
          m(4) := x"071F";
          m(5) := x"F308";
          m(6) := x"FA90";
          m(7) := x"0781";
          m(8) := x"0E94";
          m(9) := x"0322";
          m(10) := x"097B";
          m(11) := x"01E7";
          m(12) := x"088E";
          m(13) := x"0DD6";
          m(14) := x"F86F";
          m(15) := x"00D4";
          m(16) := x"0DB0";
          m(17) := x"FDA2";
          m(18) := x"FB24";
          m(19) := x"034C";
          m(20) := x"FC32";
          m(21) := x"F09E";
          m(22) := x"F9F5";
          m(23) := x"F7F2";
          m(24) := x"EF02";
          m(25) := x"063E";
          m(26) := x"FD62";
          m(27) := x"F88B";
          m(28) := x"F153";
          m(29) := x"189D";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_20.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 20) then
          m(0) := x"F9AF";
          m(1) := x"FE36";
          m(2) := x"0B89";
          m(3) := x"FAED";
          m(4) := x"FC0D";
          m(5) := x"09C1";
          m(6) := x"FF81";
          m(7) := x"F863";
          m(8) := x"FF73";
          m(9) := x"049B";
          m(10) := x"006F";
          m(11) := x"0103";
          m(12) := x"0255";
          m(13) := x"0440";
          m(14) := x"0491";
          m(15) := x"FC5E";
          m(16) := x"FA91";
          m(17) := x"FC55";
          m(18) := x"039A";
          m(19) := x"0658";
          m(20) := x"FDB4";
          m(21) := x"01ED";
          m(22) := x"0538";
          m(23) := x"09E0";
          m(24) := x"022E";
          m(25) := x"034C";
          m(26) := x"0358";
          m(27) := x"0219";
          m(28) := x"0368";
          m(29) := x"F7E7";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_21.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 21) then
          m(0) := x"05CD";
          m(1) := x"045D";
          m(2) := x"EFBA";
          m(3) := x"0094";
          m(4) := x"02DF";
          m(5) := x"F78A";
          m(6) := x"F74D";
          m(7) := x"06F6";
          m(8) := x"09F5";
          m(9) := x"FF14";
          m(10) := x"039F";
          m(11) := x"01E5";
          m(12) := x"F521";
          m(13) := x"F9FA";
          m(14) := x"FDA8";
          m(15) := x"FC67";
          m(16) := x"0374";
          m(17) := x"02C4";
          m(18) := x"F9D8";
          m(19) := x"FDFE";
          m(20) := x"0A45";
          m(21) := x"01FE";
          m(22) := x"0977";
          m(23) := x"F42D";
          m(24) := x"01FB";
          m(25) := x"FF99";
          m(26) := x"FD37";
          m(27) := x"FCBB";
          m(28) := x"F84A";
          m(29) := x"0CCA";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_22.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 22) then
          m(0) := x"0791";
          m(1) := x"FC5C";
          m(2) := x"FB69";
          m(3) := x"025F";
          m(4) := x"F66C";
          m(5) := x"01E5";
          m(6) := x"FFB8";
          m(7) := x"F90C";
          m(8) := x"FD4A";
          m(9) := x"FD56";
          m(10) := x"08AB";
          m(11) := x"02D1";
          m(12) := x"F79F";
          m(13) := x"FFAF";
          m(14) := x"F1F6";
          m(15) := x"F558";
          m(16) := x"0124";
          m(17) := x"041E";
          m(18) := x"09E3";
          m(19) := x"02D0";
          m(20) := x"F389";
          m(21) := x"FC56";
          m(22) := x"00F7";
          m(23) := x"F67A";
          m(24) := x"04B3";
          m(25) := x"01EF";
          m(26) := x"0299";
          m(27) := x"F929";
          m(28) := x"05C7";
          m(29) := x"F926";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_23.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 23) then
          m(0) := x"0981";
          m(1) := x"070A";
          m(2) := x"09C9";
          m(3) := x"EE5F";
          m(4) := x"F6D8";
          m(5) := x"0FB8";
          m(6) := x"F6DA";
          m(7) := x"F7A1";
          m(8) := x"06D6";
          m(9) := x"1DE6";
          m(10) := x"0907";
          m(11) := x"02A5";
          m(12) := x"0AD5";
          m(13) := x"15D8";
          m(14) := x"FDB5";
          m(15) := x"FB1F";
          m(16) := x"F82D";
          m(17) := x"F253";
          m(18) := x"1194";
          m(19) := x"19E7";
          m(20) := x"EE3F";
          m(21) := x"F3F1";
          m(22) := x"0B59";
          m(23) := x"0225";
          m(24) := x"EF96";
          m(25) := x"FB70";
          m(26) := x"EFCF";
          m(27) := x"0263";
          m(28) := x"11AD";
          m(29) := x"F371";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_24.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 24) then
          m(0) := x"E88D";
          m(1) := x"FF79";
          m(2) := x"12F9";
          m(3) := x"007E";
          m(4) := x"FF55";
          m(5) := x"00A9";
          m(6) := x"041A";
          m(7) := x"F8CF";
          m(8) := x"F8A1";
          m(9) := x"157A";
          m(10) := x"F752";
          m(11) := x"F8C7";
          m(12) := x"FE0B";
          m(13) := x"F767";
          m(14) := x"0FDE";
          m(15) := x"04B4";
          m(16) := x"ED1F";
          m(17) := x"FA53";
          m(18) := x"FA16";
          m(19) := x"0014";
          m(20) := x"13EA";
          m(21) := x"0A10";
          m(22) := x"0731";
          m(23) := x"120F";
          m(24) := x"060C";
          m(25) := x"F4A7";
          m(26) := x"FFE8";
          m(27) := x"0AE4";
          m(28) := x"03A9";
          m(29) := x"EAA6";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_25.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 25) then
          m(0) := x"FC3E";
          m(1) := x"E819";
          m(2) := x"EFAC";
          m(3) := x"0353";
          m(4) := x"0A41";
          m(5) := x"EDC5";
          m(6) := x"FCB7";
          m(7) := x"1003";
          m(8) := x"05C0";
          m(9) := x"F166";
          m(10) := x"0677";
          m(11) := x"F7E6";
          m(12) := x"F241";
          m(13) := x"ED9A";
          m(14) := x"F66D";
          m(15) := x"F8EB";
          m(16) := x"FF87";
          m(17) := x"0B4F";
          m(18) := x"102A";
          m(19) := x"E790";
          m(20) := x"FFFB";
          m(21) := x"FEEA";
          m(22) := x"F2FC";
          m(23) := x"E8BB";
          m(24) := x"09B6";
          m(25) := x"0111";
          m(26) := x"FEF1";
          m(27) := x"071D";
          m(28) := x"F725";
          m(29) := x"FF97";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_26.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 26) then
          m(0) := x"08C7";
          m(1) := x"EB21";
          m(2) := x"EAA0";
          m(3) := x"02C3";
          m(4) := x"FE62";
          m(5) := x"07CB";
          m(6) := x"E738";
          m(7) := x"1DAF";
          m(8) := x"16C3";
          m(9) := x"17BB";
          m(10) := x"F65A";
          m(11) := x"0D3D";
          m(12) := x"0277";
          m(13) := x"0BAF";
          m(14) := x"FE90";
          m(15) := x"06BC";
          m(16) := x"F5F4";
          m(17) := x"F1AF";
          m(18) := x"052D";
          m(19) := x"0B8E";
          m(20) := x"FAF6";
          m(21) := x"17A0";
          m(22) := x"00C4";
          m(23) := x"E157";
          m(24) := x"E9FE";
          m(25) := x"E531";
          m(26) := x"D460";
          m(27) := x"0723";
          m(28) := x"0F08";
          m(29) := x"0226";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_27.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 27) then
          m(0) := x"EB2C";
          m(1) := x"F30E";
          m(2) := x"09DB";
          m(3) := x"05C0";
          m(4) := x"0756";
          m(5) := x"F409";
          m(6) := x"22BB";
          m(7) := x"058E";
          m(8) := x"FE04";
          m(9) := x"FEFB";
          m(10) := x"009D";
          m(11) := x"F410";
          m(12) := x"F576";
          m(13) := x"D48B";
          m(14) := x"F73F";
          m(15) := x"14CA";
          m(16) := x"02A6";
          m(17) := x"1181";
          m(18) := x"0180";
          m(19) := x"F9E7";
          m(20) := x"1A0E";
          m(21) := x"0C5D";
          m(22) := x"EF85";
          m(23) := x"0732";
          m(24) := x"2946";
          m(25) := x"0771";
          m(26) := x"048A";
          m(27) := x"0F90";
          m(28) := x"0137";
          m(29) := x"E9AF";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_28.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 28) then
          m(0) := x"084B";
          m(1) := x"0314";
          m(2) := x"F256";
          m(3) := x"FF59";
          m(4) := x"F2E2";
          m(5) := x"0813";
          m(6) := x"F6BE";
          m(7) := x"04AC";
          m(8) := x"057A";
          m(9) := x"FA04";
          m(10) := x"0221";
          m(11) := x"041C";
          m(12) := x"FBA5";
          m(13) := x"FA60";
          m(14) := x"FAAD";
          m(15) := x"F87B";
          m(16) := x"FFD3";
          m(17) := x"FE58";
          m(18) := x"F406";
          m(19) := x"0182";
          m(20) := x"FD32";
          m(21) := x"0583";
          m(22) := x"0A44";
          m(23) := x"F706";
          m(24) := x"FDDF";
          m(25) := x"0172";
          m(26) := x"FD88";
          m(27) := x"F58B";
          m(28) := x"FF95";
          m(29) := x"05CA";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_2_29.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 2) and (nno = 29) then
          m(0) := x"F6C9";
          m(1) := x"F37A";
          m(2) := x"05C6";
          m(3) := x"FEB2";
          m(4) := x"F3CD";
          m(5) := x"112F";
          m(6) := x"FA07";
          m(7) := x"FC60";
          m(8) := x"FC94";
          m(9) := x"088C";
          m(10) := x"FC8F";
          m(11) := x"062B";
          m(12) := x"0450";
          m(13) := x"0036";
          m(14) := x"FC49";
          m(15) := x"0230";
          m(16) := x"F327";
          m(17) := x"FC75";
          m(18) := x"FDDB";
          m(19) := x"0A27";
          m(20) := x"04CB";
          m(21) := x"0818";
          m(22) := x"003B";
          m(23) := x"F997";
          m(24) := x"FFC1";
          m(25) := x"FB83";
          m(26) := x"F2F2";
          m(27) := x"F758";
          m(28) := x"0BB2";
          m(29) := x"F89B";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_0.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 0) then
          m(0) := x"0919";
          m(1) := x"057D";
          m(2) := x"F596";
          m(3) := x"12E9";
          m(4) := x"FDA1";
          m(5) := x"E977";
          m(6) := x"F0BD";
          m(7) := x"FDB4";
          m(8) := x"E655";
          m(9) := x"E756";
          m(10) := x"2464";
          m(11) := x"010B";
          m(12) := x"EECC";
          m(13) := x"104A";
          m(14) := x"FCF0";
          m(15) := x"E9F6";
          m(16) := x"0479";
          m(17) := x"EADB";
          m(18) := x"EEC7";
          m(19) := x"1244";
          m(20) := x"F6A2";
          m(21) := x"13DD";
          m(22) := x"F4C0";
          m(23) := x"E4D6";
          m(24) := x"044C";
          m(25) := x"13B5";
          m(26) := x"1932";
          m(27) := x"060F";
          m(28) := x"035E";
          m(29) := x"FC35";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_1.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 1) then
          m(0) := x"11D2";
          m(1) := x"088E";
          m(2) := x"F17A";
          m(3) := x"ECFB";
          m(4) := x"08D8";
          m(5) := x"03B5";
          m(6) := x"08BC";
          m(7) := x"FD3E";
          m(8) := x"EC60";
          m(9) := x"F29A";
          m(10) := x"1F23";
          m(11) := x"031B";
          m(12) := x"F317";
          m(13) := x"149A";
          m(14) := x"0A0E";
          m(15) := x"FDC4";
          m(16) := x"0BD8";
          m(17) := x"FC6B";
          m(18) := x"1DAB";
          m(19) := x"FEFC";
          m(20) := x"FB0A";
          m(21) := x"0E20";
          m(22) := x"FF19";
          m(23) := x"D77C";
          m(24) := x"FDAD";
          m(25) := x"1CCE";
          m(26) := x"E81D";
          m(27) := x"2294";
          m(28) := x"04EC";
          m(29) := x"F60C";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_2.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 2) then
          m(0) := x"1509";
          m(1) := x"FAF8";
          m(2) := x"137A";
          m(3) := x"F3A7";
          m(4) := x"2A28";
          m(5) := x"CDE4";
          m(6) := x"0653";
          m(7) := x"DA3A";
          m(8) := x"FE79";
          m(9) := x"0F9C";
          m(10) := x"FCB4";
          m(11) := x"F5A0";
          m(12) := x"07A0";
          m(13) := x"DE38";
          m(14) := x"F9CB";
          m(15) := x"0D8D";
          m(16) := x"2AB6";
          m(17) := x"E353";
          m(18) := x"158C";
          m(19) := x"EA55";
          m(20) := x"0A1B";
          m(21) := x"F00D";
          m(22) := x"03DE";
          m(23) := x"05E9";
          m(24) := x"1726";
          m(25) := x"FCCD";
          m(26) := x"D240";
          m(27) := x"2803";
          m(28) := x"ED27";
          m(29) := x"0098";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_3.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 3) then
          m(0) := x"FEED";
          m(1) := x"FC81";
          m(2) := x"FC9A";
          m(3) := x"EB2C";
          m(4) := x"DFEE";
          m(5) := x"F2A5";
          m(6) := x"09B5";
          m(7) := x"051E";
          m(8) := x"2919";
          m(9) := x"071F";
          m(10) := x"ED19";
          m(11) := x"FF07";
          m(12) := x"00B8";
          m(13) := x"0B77";
          m(14) := x"2298";
          m(15) := x"0C4C";
          m(16) := x"D417";
          m(17) := x"FEE6";
          m(18) := x"0AE9";
          m(19) := x"E866";
          m(20) := x"110C";
          m(21) := x"F9DB";
          m(22) := x"FB6F";
          m(23) := x"113E";
          m(24) := x"1B6F";
          m(25) := x"E7AE";
          m(26) := x"F1FF";
          m(27) := x"13FB";
          m(28) := x"0704";
          m(29) := x"10DB";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_4.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 4) then
          m(0) := x"12A4";
          m(1) := x"127E";
          m(2) := x"E7E0";
          m(3) := x"0120";
          m(4) := x"0C8A";
          m(5) := x"F9D6";
          m(6) := x"CE05";
          m(7) := x"F51D";
          m(8) := x"19E2";
          m(9) := x"DA13";
          m(10) := x"1BBE";
          m(11) := x"1A28";
          m(12) := x"E45A";
          m(13) := x"F1B5";
          m(14) := x"1135";
          m(15) := x"0F2F";
          m(16) := x"F216";
          m(17) := x"F6A6";
          m(18) := x"05FC";
          m(19) := x"0021";
          m(20) := x"023E";
          m(21) := x"FAA4";
          m(22) := x"FF4B";
          m(23) := x"FE3E";
          m(24) := x"F044";
          m(25) := x"06CA";
          m(26) := x"0C95";
          m(27) := x"D56B";
          m(28) := x"0476";
          m(29) := x"0D7C";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_5.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 5) then
          m(0) := x"0559";
          m(1) := x"F2DD";
          m(2) := x"197C";
          m(3) := x"F7D1";
          m(4) := x"FED6";
          m(5) := x"0EBA";
          m(6) := x"0AA9";
          m(7) := x"E77A";
          m(8) := x"E0DC";
          m(9) := x"25D6";
          m(10) := x"079E";
          m(11) := x"E54A";
          m(12) := x"1ED5";
          m(13) := x"1987";
          m(14) := x"09A3";
          m(15) := x"119D";
          m(16) := x"0543";
          m(17) := x"1894";
          m(18) := x"DC8A";
          m(19) := x"1C08";
          m(20) := x"FC63";
          m(21) := x"0360";
          m(22) := x"F8E1";
          m(23) := x"F84A";
          m(24) := x"F13E";
          m(25) := x"F194";
          m(26) := x"E0CC";
          m(27) := x"EABC";
          m(28) := x"02ED";
          m(29) := x"EC74";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_6.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 6) then
          m(0) := x"FAE4";
          m(1) := x"E992";
          m(2) := x"1EE6";
          m(3) := x"1B61";
          m(4) := x"EA1B";
          m(5) := x"D0F7";
          m(6) := x"01B1";
          m(7) := x"F4DA";
          m(8) := x"096D";
          m(9) := x"0A69";
          m(10) := x"091F";
          m(11) := x"EC57";
          m(12) := x"0827";
          m(13) := x"1236";
          m(14) := x"F490";
          m(15) := x"EB47";
          m(16) := x"F4F7";
          m(17) := x"E258";
          m(18) := x"E5F4";
          m(19) := x"0E73";
          m(20) := x"0274";
          m(21) := x"0684";
          m(22) := x"FE13";
          m(23) := x"18DC";
          m(24) := x"1403";
          m(25) := x"EB06";
          m(26) := x"1033";
          m(27) := x"0A99";
          m(28) := x"0024";
          m(29) := x"0B5C";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_7.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 7) then
          m(0) := x"1357";
          m(1) := x"019E";
          m(2) := x"0C67";
          m(3) := x"E9AC";
          m(4) := x"1386";
          m(5) := x"FFA6";
          m(6) := x"0208";
          m(7) := x"0845";
          m(8) := x"0360";
          m(9) := x"1052";
          m(10) := x"FDAB";
          m(11) := x"0F2C";
          m(12) := x"0DCF";
          m(13) := x"0A31";
          m(14) := x"0108";
          m(15) := x"110E";
          m(16) := x"FCAF";
          m(17) := x"048B";
          m(18) := x"F335";
          m(19) := x"0AA7";
          m(20) := x"FFF5";
          m(21) := x"FE5F";
          m(22) := x"05B1";
          m(23) := x"1046";
          m(24) := x"F435";
          m(25) := x"099C";
          m(26) := x"FD2D";
          m(27) := x"DA36";
          m(28) := x"FC60";
          m(29) := x"FCCA";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_8.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 8) then
          m(0) := x"22DE";
          m(1) := x"106E";
          m(2) := x"DFE4";
          m(3) := x"FB7C";
          m(4) := x"F589";
          m(5) := x"169C";
          m(6) := x"05D2";
          m(7) := x"135E";
          m(8) := x"F537";
          m(9) := x"F6DD";
          m(10) := x"F91C";
          m(11) := x"16C0";
          m(12) := x"FF8B";
          m(13) := x"D71B";
          m(14) := x"1728";
          m(15) := x"FC92";
          m(16) := x"F4B9";
          m(17) := x"0B27";
          m(18) := x"00E8";
          m(19) := x"FA83";
          m(20) := x"0479";
          m(21) := x"FB65";
          m(22) := x"F2C1";
          m(23) := x"1ACB";
          m(24) := x"0E79";
          m(25) := x"F1B6";
          m(26) := x"299C";
          m(27) := x"E4C7";
          m(28) := x"F970";
          m(29) := x"0482";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_3_9.mif
-- Expected length: 30, input: 30, padded: 0, trimmed: 0
        if (lno = 3) and (nno = 9) then
          m(0) := x"DE42";
          m(1) := x"EF92";
          m(2) := x"172F";
          m(3) := x"FDD9";
          m(4) := x"FE75";
          m(5) := x"16C7";
          m(6) := x"1503";
          m(7) := x"181A";
          m(8) := x"0B86";
          m(9) := x"FF37";
          m(10) := x"E347";
          m(11) := x"0E2B";
          m(12) := x"01A4";
          m(13) := x"F9AE";
          m(14) := x"CB7A";
          m(15) := x"FEC3";
          m(16) := x"001F";
          m(17) := x"06DE";
          m(18) := x"1147";
          m(19) := x"FCFE";
          m(20) := x"FB8D";
          m(21) := x"0896";
          m(22) := x"109D";
          m(23) := x"0F36";
          m(24) := x"ED8D";
          m(25) := x"1113";
          m(26) := x"117A";
          m(27) := x"EFF1";
          m(28) := x"0EB3";
          m(29) := x"0576";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_0.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 0) then
          m(0) := x"181B";
          m(1) := x"123D";
          m(2) := x"AC6A";
          m(3) := x"CE16";
          m(4) := x"3614";
          m(5) := x"42E0";
          m(6) := x"B6BA";
          m(7) := x"02B2";
          m(8) := x"FB59";
          m(9) := x"C756";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_1.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 1) then
          m(0) := x"E431";
          m(1) := x"CB16";
          m(2) := x"3DEC";
          m(3) := x"287A";
          m(4) := x"C86D";
          m(5) := x"C0E7";
          m(6) := x"3399";
          m(7) := x"CEE6";
          m(8) := x"EDEA";
          m(9) := x"22E5";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_2.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 2) then
          m(0) := x"F3F0";
          m(1) := x"A60B";
          m(2) := x"AE0B";
          m(3) := x"D6C2";
          m(4) := x"BAB7";
          m(5) := x"4965";
          m(6) := x"1535";
          m(7) := x"002C";
          m(8) := x"0EF1";
          m(9) := x"0BE4";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_3.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 3) then
          m(0) := x"CF7E";
          m(1) := x"2786";
          m(2) := x"27E4";
          m(3) := x"E501";
          m(4) := x"FE62";
          m(5) := x"2101";
          m(6) := x"B486";
          m(7) := x"ED32";
          m(8) := x"A099";
          m(9) := x"414A";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_4.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 4) then
          m(0) := x"341B";
          m(1) := x"06AC";
          m(2) := x"AAE4";
          m(3) := x"47CA";
          m(4) := x"080D";
          m(5) := x"DDFB";
          m(6) := x"3A73";
          m(7) := x"CCD3";
          m(8) := x"F521";
          m(9) := x"C9A9";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_5.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 5) then
          m(0) := x"C470";
          m(1) := x"0DD3";
          m(2) := x"2152";
          m(3) := x"253E";
          m(4) := x"B648";
          m(5) := x"12AE";
          m(6) := x"C73B";
          m(7) := x"E831";
          m(8) := x"3A4E";
          m(9) := x"9A11";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_6.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 6) then
          m(0) := x"B5F9";
          m(1) := x"C9B2";
          m(2) := x"D7C5";
          m(3) := x"2660";
          m(4) := x"4F6F";
          m(5) := x"D49F";
          m(6) := x"B7CE";
          m(7) := x"0BBC";
          m(8) := x"0965";
          m(9) := x"032C";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_7.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 7) then
          m(0) := x"408E";
          m(1) := x"0295";
          m(2) := x"158F";
          m(3) := x"E18D";
          m(4) := x"D4B7";
          m(5) := x"34C4";
          m(6) := x"47D8";
          m(7) := x"F111";
          m(8) := x"B4FA";
          m(9) := x"D38A";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_8.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 8) then
          m(0) := x"060D";
          m(1) := x"3EEE";
          m(2) := x"B9FC";
          m(3) := x"D4B7";
          m(4) := x"BDF6";
          m(5) := x"B9B7";
          m(6) := x"D959";
          m(7) := x"D1E1";
          m(8) := x"2526";
          m(9) := x"3302";
        end if;
-- Auto-generated VHDL snippet for pick_weights
-- Source: w_4_9.mif
-- Expected length: 10, input: 10, padded: 0, trimmed: 0
        if (lno = 4) and (nno = 9) then
          m(0) := x"185C";
          m(1) := x"05B2";
          m(2) := x"5F36";
          m(3) := x"ACC2";
          m(4) := x"2E5C";
          m(5) := x"AD88";
          m(6) := x"F07E";
          m(7) := x"DDD5";
          m(8) := x"1F2B";
          m(9) := x"D0FA";
        end if;

        return m;
      end function;

      constant ROM_IMG : memory_t := pick_weights(layerNo, neuronNo);
      signal   q_d     : std_logic_vector(dataWidth-1 downto 0);
    begin
      -- 也做成 1-cycle read，跟模擬/你整體管線一致
      process(clk)
      begin
        if rising_edge(clk) then
          if ren = '1' then
            wout  <= ROM_IMG(to_integer(unsigned(radd)));
          end if;
        end if;
      end process;
    end generate;

  end generate ROM_MODE;

  ----------------------------------------------------------------------------
  -- PRETRAINED = false：外部可寫入（保留原狀）
  ----------------------------------------------------------------------------
  RAM_MODE : if PRETRAINED = false generate
    type memory_t_ram is array (0 to numWeight-1) of std_logic_vector(dataWidth-1 downto 0);
    signal mem_ram : memory_t_ram := (others => (others => '0'));
  begin
    -- write
    process(clk)
    begin
      if rising_edge(clk) then
        if wen = '1' then
          mem_ram(to_integer(unsigned(wadd))) <= win;
        end if;
      end if;
    end process;

    -- read
    process(clk)
    begin
      if rising_edge(clk) then
        if ren = '1' then
          wout <= mem_ram(to_integer(unsigned(radd)));
        end if;
      end if;
    end process;
  end generate RAM_MODE;

end architecture;