`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dy/2iy6PseKiN/Xn+TZlVmCmZK1Vp8I++uDJEYDNtTXJi3fTbTUN3n//0HKXWAOW
OcEKSpcXdDAfEDN3UOUM+AGWenziX1bYmtDvPlyk1Y5Jt8agcBwkZiLTTlE2lEVv
ovOV6p5skAnqu7DuAbrMUwzdy8RRPLnL8kZvXvNVOrJ5PTVz8NSfM11psYbCNnKr
1JlVTKsab6WkFdVCbIRW5/X0FBRZMTK9BjTd24Nn0xW5D4c1dwEZVZXvX854X4ke
SfopQ2VcjozSYpNcmwF9bWAHjsZpc7lj42FkOwegHxgBp27UiJvGDWXL0iHU5ikK
EvjOF53y8MeWcKai7jfym3QRSZWwcAIqSNdVEIM3Rl+CMPbMWKnKDtZLczwjO4Jw
4s+SvvYnbarmAv44+Ebdh20wnXFX0vjZnX1edh6DZop0hQG9MWvG5x2HG2TwC836
U7heJ6YLfazKO/YwU5b6q0DBnXc6el2kMbPeo6YzOV1dLZqNf5I77l0+NY1OWOBT
fzatCwayJcLrDj2JCkysG56sF3xfMhs+kyK2kovgx9IxY1MnV97o2HpsU3P7N9E3
kSDT+An3ovA7ZimBQg05UBwM3AZ0b2i4nF/Vnl3FQK2yHkd/YFqtrex0Q1CdziRm
QdZLDojp+9gUPf/+WIxB9rcnPRwg5dJB1x3LGa3DrQF8uGAsrSLob8H5kiv9uGZY
+s3q+svF2ZOSRHnG0F65jv6C9AFuBUhrrEbVSKq+4z5q6exr9bcNSaIvyHYt+AOT
lpVc2ChWURZIM4tMLoXot6CmJSUPdCtRIurpI407Rrw4QOzB4eG3VRixYmWGV3jz
3fI9FteLMpiFR+Y8uRRa1Y7FVqoJCEVS8GjiSCDSq0e94GGIlFFMc8uR7Lyin1ob
Ij3h5V4s1hIxqR2iuZcl/sMoXYxgnk/hTwbwgl1UGvjtzHLYVNxx4mXGEQqIrJES
NGiXz8Mtunvmp3JIHA+PfL3eSit9vvW0yPh/18ap4VnEw+OB3lL4VVSCvNC/s3eB
H2ScEtDiqbAfniqwcF/HNG28gWWLiKKoiLpllEI63S89axmRwPviOFA/i/cN69LB
lC2BSRERtx3LhjJ1DKEwjeBaSiEFiInDhwzpMld3zb4m+4nfxJWToblNPq4sCtv4
E7AcyZ7tSPJuu91RynCzbwldGS6Dj5ZJdaNAnEkW38fWxK9cnhLh2dCCsHTH5lcF
Qf0db9Wnx7oT1w5a9cNdtmXZ/cCwiCqEuEsIJLhFHfY=
`protect END_PROTECTED
