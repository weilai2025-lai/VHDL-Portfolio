`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/iLgXMDVHjJk+63WZKZTcVraSlcIRsHjj5F33jf5yL/Dq7TBlyPMhimumqpK6PBF
pcU7WOcJqyzLPMnyg6y5PPKOywwJpUV9O5tWcoHoTYogaEWCP1jzDRgmduV0hWLD
vL/96lI+WoBsbrFjPwELlHI2P/qt8T1OhnlhRih8mdWZxTWz11HGCouoS0FEsumL
QaNzbXyqfiCPfnmqCGklLaFns6iEm1RS4uor5KXIozn1n5lwcuyoAjfsezhIcl+S
TX8v6SZBW5TxB9ujZlZq4LvuUbY4RkLT9NerLw53aWAwIMTp1atH6s6W75MlY/cC
gwKKtVwdDNvYDjS/YLlvPCkiYT2Yvoa6DX9Bu8bra5ofPs4wtHsR3gFIODaPXSjp
cnhZz5n97jEluu6t7DWSShzkZfVXcCxXBCX7XElLo0d07CBLueqhfub0lmaDbdtt
Qf6uDT8WSnua5TeK8Zf4vucuFDlOZLUURAFMXhGr49GolPmy6kEFqCFQAgHJ23mo
fllJQba93FxQhT5Q0eR/vby3ZgzXAoosxR321vGXKIOZkc7IM1K2aFx99I7E/hfB
WW6XdnBHr5JqaLyP86BR+EPpN3kH1gmr9qzyUuWN5TMEuedYUzfrNrRyyHGgPDWI
+btzKdiSRd5WmJqQN1jpmvsemoVfWHQt0nWll5jsl8pmst1B5ofphQq97DijJKU6
xYMmettITODzL/DYx9j6LqoYw2pJCVhALBAR5wiSnfJs27iyIj/0jmzovnOKUpMt
QTsw51loe9hiONnKBQWydnk+lNs6BYwbecbP1ZLII71rjUG75MOxvoMAI1RlMKZv
YMRlyebQR4BejOGN4gHpFw58SJUg+jDJrAjeSX4Rv7TzDx3ZH9Y97susB64yExuv
p7BwzFu4z36mzCdm0AoR3T+Yk90Dsm117SDt4GJ/ooReqO3B0+ysdCQGMowPcFyO
b8yfQXReQ6le0+oeIqPCELaf/sXaQlQc63APu6QWcvyEiOW3zth/oM3bs405nwvJ
7FTMuWsZXn0GU2Ic3uhCPJI736LxjGCQN6IbGGhvyxDZzEzDh0F1kWObwhCnzPZb
+arkGrKWKjX4o2HlVLledldRD4Tc3/fjK8qiFxOcvTko5StmRl4UblGPJqZBDcWp
MO4OosAr4iFdNHyqcRg4B57mxL8MEAdoMLoMQjT6EYGXQFSylnjFcrnNn0Iiam1q
2Xb39ywlQdo9jzPwPEgk7vpqmpUvf6o5xQBGeZmbmlG7dCHdU3xbG/CqX3u9up7t
Wynr1yS/9+TP/gEWvmUDAoNkaEzkIiCk5ks/vezUcpSAFdwSHVhIyM7zQqSkk0qa
pJ8RAxH13nw9bgBdzdMTGM2HfWj92rOge9E9mE0XVr1O3F3WCVcKJYo8Jpezjy28
NlIVWGJ+uCnMpeH8/fgsUGXG5Z7XBNe7OpAVfL8rSqRTH0YL51ORcshFuLdAOgA3
1ec1VjCed8XRwEZMZZ61s4aJucfMj4NpDZQTxaiF75ANWcYlmeaSYHmkCqYQjWBl
EY4QDMjbBR1e1osu+HdfI6tMcCNHUpr+sT0Otym3D9WaIReezh5QlzSpPO9Rjnfp
1wAPweluIacHIRTsDTVfB7HsSbUifIyif+bEcCXq3BswsB7g1IPEQemPneTM5WLI
FPKe8bL0VHM5v45r3FjAnL/L+WkXmf2VCVqPibCkTvoNaSIG29AA33mxKAEkAlDb
VnjK82TFD8nriloSV7Vj7EOuhuNfaWjVOvJeFBC3mC1iiR6nhGUbGItIkWFtCyfB
EY7EHxZOiluYC1wAmK3V95e74h0RP3lzbdtRL3hnZZgm5DUiuHAC1W/+31ALp5kY
jzGf7hUvj8bff3q2K5vgT9w/QEEqu7A/oHVGJzT2dTLjJz6CYeciIjntJrN/7dM1
ptfRyUaH1IU8dy/zicMyRJLUbrctzr9zw5/myfflE1EZSOqfgZD6dX7HcUYlacdK
2W2oFhgSeUrz/Quk3+GsDytPAygaR4zyZzNRIv9lcCL94AhyQhdoHg2lxB2QQGsX
f9qCk53HfwVYjb3Tj3W5hfR1hg5SSOesHMYEu/3asqnE9Tg+R9wKjfnJatR+cI6K
cVI6xH1GjFNRByNA9cyEp4Bk2/xZyWHPHjh4d1XlEV2LRNXo75pG5foGadcsRM2g
8PZ1XjyVijQiuaioORsF4KGphva1c1UyNXUBpCGclR+UVhP2HWAz4EnR+nkRg7If
szx/ETAH/RYnuh/laxm2d5Ly+PpOjbnjEZ/EcKoHMyBTu42KvKlBofWg2h0FLs7u
emtNKnK6644ZwEht2UxC6KGoZj+YhxHSI1H2Vpp3op+9UjnrmAQa1ZwQjoE9KQrT
NOsbD1JY25+IyKdLQ69I7uoMeLZDFRsXLkB69nmwCVmd9uQJkRfmNsrFxmfMuA3w
tHMjvFmcZ15pKuObfPxfdBu9mBG++LGjwCUR9Tc/WiTaN1/TVxLyMdEMdgyEQqxE
vQssgYoy7mx8Vp9ZAxZQ0s4MPeX5AiXRbPdXE9WgMSE=
`protect END_PROTECTED
