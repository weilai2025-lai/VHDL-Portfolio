`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJ5DyU0JXIMsGXw7AzoH4M7C5+rT1Xuehe1G1r2l2zTjEJCzd/h8e5/Kncl0Au/X
t0XQAqEtNmLi20ELjQwcQyxb+OC/1s/trNIgXBdLGKVOTgx4O18SYbttN06gW/za
qYvIZ/GD/Xk9Q0GTvYIv2bDb9EGGlxa7dt++slEGBAlowAghGHBRZyg6oyLt6MJJ
1RE7ETDdrzM+FYVZs95fAf+Bw40UzG1DLfOr8JFPzcsNg+CjG6JQ0nV3mQ+opik3
lI6ADuXN4DgPqgtD3sBQm0KtZkqWkllNYCirVajQMwdXdKhJ7gXCwxrwZnHbz1yv
jXrKWOexOeRFdra7Tj+vZXeo7agNZSVXAcu6Lb2fwoWP6EzNszJeyUf6EQb1kcLA
RTgnJX8spBDuDEp9CBUNRqCmldUTomd97JrK3btd7RjRKmzH80tK7WTjpUihiRMs
lrECxbpptL6/gx8QKayj2mIW5x4ikrvCPweFbQlHPmzQYKw3nlM768DYIMZ0p0sU
lWprD1PzlyBkUDYFpnVnxlA4QB3ZCE1QqyTj4TRYTeUO0pXLxF+5ZNOKsGSLDmz5
GbRCwrWvc1hndXWI7PaWlRpgmeE+4HRa3yeJGxsx/56Titb3phd2yqiPI1EPRDnx
t2D90zc9t1X/Nk1p0gyE/uTn3Kq42J99TskOYsx6jRwLTWeda5FqfYmWRXTJ0ba9
t5Afb5UYKSennfbUAom2QtKhlFr/4NPlfYTwMJCVdtfSmSte+8lvfTbieCjyB2as
KHdLwZSPqquJI+5csTAmW5J/8zW+eECg9FkmzywVWrUYlqD6EmYz8CCGFONA30wz
s95yDtX65padWp6+eoWiynxgAzXstycz7OkWxH+qrcNcdjdhLCnWL7TRBgG3ZJec
jCtOAQIJbP6HQQ5p2mTyZVC2RSDob7Jjp+gZhA2M/1e7MveI9ivGAQZNTpm2mLpI
hz0DpbYYmaticsPwvdXtDq9z51+g0tMGBznrtK6VNWMTgrA4GmignAFTajZsex7q
YJWY0NsU6mZF4hAHFEbi3NlL2/OFaPy5vehOvFt9Xn5IHBFLhFzoGbLAESz9cAMT
XYKJ2cyEsM42dXUfKI5mRDqU8j7l5Dh1lygKYbVVG5Y7N+5R4zLIATPyPzTwj6de
6varR45Wzn7N8o6mtSrtpJwMEvcFet5R7xP8QWQ0B+ZqMG231eolMofBmbx8NQ45
YCOOk/4eve/gOF3rREYDtputUst/jJTlun2jbW833Q5zLfYiS5lgwntNSxDoo9Sq
Bm8V9KXtWolSjdmnZR8thkiJhn918aIoQV9unoNEFgBL9nuZR1VQBCW2e7A9CJ8c
Edb7J28cLF+/3YcTFKLbE3iObzvimCNZAJcANKisTJI81OdrsYNxljiheaxok0+q
xDdSHMn6jrJPgRxQYkbCf0DV4X1tlVWlcHgyPDqA+i+g2rfDaWdgRnAUtdE3eO71
MJMHW81dp2efVkGVkyJHX4BzAfMMqn/6DHCdalKrqODZRYp3kTh2Uqt9kywWQfm+
HUKEcPKcpArrG69HzuLVm1kIev8W2dLqUdnCWXQXZjQwsYB1nyJO3KVIntD3Z5FW
XZzhNbWmV3PcF/2QwSSwbce4XPfztl1RhqOq4SrRyCdUKTcme6wwOUJQ2nwXaPua
Uwak/2mOj5LiDO7DWQhito8uCVvv9Efv2fqdCfUhno4IQftlCXXyv7r1cjs9mp25
gH9MgmBsEE5EFYBzWWVtFPcpofLen7PljYUPD+sWT7MTn0585lT7nNpqnKrAnPfr
1hl9FiFzE80H9N2bfkxFdGPSbDOu92ZpY4lGV/lGUZOsaT0YApjFlLz2Bnf6dYLV
`protect END_PROTECTED
