`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x8Qq6+h+ifRc/NMw/yGtWsxs5gXR2FvnAVBBWXC07mtVF71Kr5uLphCqSbeTauJ2
kofGDuPssFqX1H75J9EzwPCl6nyy/MCeWvl9Msv6XFUf/PNQdh01mj0VYZkOMqP7
hTolzNQ7n5u5eKCDAIvDEIJDj9QtFOrRBSh7lffcMUfZPY0H+FdGHoiTJkWDiwfo
0dkO19mzpj/Ouq60MXqBkHrW1QTFzXtSdz2WKLhVQbX1KEDrkrkD8EDZ+nqOFroj
nMYLB7XWwE9RkFzNjrV2n4pyqMT1iyyz5esKMkJXB7sel2mSFJM4zhEKNrdlWrVd
VAwQYJb83T4CXgOCExDtONXcIWQP/F9YBqstjRXIZwU1XEKLOlqirpeWEQsbA0rd
iQFEoEGPfsdieJZerAS96BBdxS8blE0vdnkdgDTvkDzUiBABn/wNotwRjtNjlQdA
tR9vf6RD/wcn1NkMHIJidZ+LR/HmlVe50IU9PAaakccxzy8LTVrpOQzWbTQfq/2+
1XBK8ET2BXCJ3QrjqKcXpCf4kr91J5FFdJs5iwMoVGQSjFE/fN8+Puj+hwcVyBxa
bGXo483MFUYdK1cTWzYXt2XUN2VhHStJ4ADqUYK5JPqT4UdT2Yo7hm4eM3GC2dYh
z4k79Z/ef+qMd8pHg7R0QWixZuDhtajKa1Vv4puxOodMJUi63HHYeo8BuJ7wWI1o
XyO1+ZRk5/oMy2vhgE8/YoRkxKM6hy9XGyiAUXkBmzcYJvTyfqHLmJayLZF/yAWA
ysVb2UATt57CDkOfHhooURbx4UPFtc1MoUV1gAVSURyqKzw62jymucxpNKdr1Bum
t3erQNsjn48iyVvNGjrjucqFqLzVqwG5AJSJ0/yql6YZCKq9kZomJa7P49+9l4w3
e8UuxL33GsELRMMjXyD9wKYHIabYZmXdzyYZ4UJMK4OFg2lyybOkq+L/EJ+M4r2U
X7aRaQDWGeytYDmnj3Np2XkvR23wRzUAhgdKOpUjUAWq5FUEJrGo8nPWnuL8dBFU
whzSxNDzg2n3KX/sYBvGtto/Pg3Vj76c4ZLDcE0F6F5uTd6RV0Se9GKYCqo6uuTr
7cbUVHpySsY6djVFMrSR/FceNFmvdTshM7fliuT51j5eyQK8vwXPMiMF6Of9UmgJ
2VYXk+T+9R4UKnitZPT5INubnlMMK2Hsuy29M+XglITDJF2tdFsCN+tYZPN2gZu/
pmp/HuQ2xwceby7aUbPWjiKeJglnfaJP1TiF+HlOqSc4FCH2SURc1vTbmk00G9zV
k+EmKq5skbopTht6KpOxZv4CFq/0C4JRI3DdBsUzSr5gCDGlCIYla1PyeKaKxCNH
XaIusBXrGGZITmup6utcC8jYFumPmWlpJcGS9o3iNEePS6gzSgnlUpDc/mtkgGnh
P8lsoa/j9tZLJd+iiG+TGEGx29KAiRpnbDGUi0KuD61GkxjlikGhDt7AzzOXu8hV
6WlHI4TsotzqVYZliHzN46r8MSW+ESz8z14yywSFyZiaYZr7y857Ir2HY4618HoS
fi6C9wqwJnqB46AabBxguEr+KrqaYzCE2Gce+58nDLEhAZOuy3jUcT8beP5pA7s2
eyDoWneCDia+8CY+yoCBC+fhplkyuL5aiT1/A7DV/VcceakxMM8OArGr+O+rzo1K
Ok8xGJpsULWNbS/CEMeBeVjtw/1Fe1AgvubFeUYlcxbzdqiD+RSrZjCcYjhBVymQ
C5I+VvhsJFZVm+cS9MuEAewEdbgaE0JyUCm9fiHcJrgxz3hlivE/OqP188W3AApI
JzjpFVs1wfKybnxQ57fTUNcLXrsajQwa+ZIyJam7I2W6dTmsWBlv9h+fLbAxiBEr
Teb362qBzqav1L3xuAt+MIQn9ugefGz7l6r81ixRRoz5XMYo15N/p5vbya+7Ao4R
oAvpyrwnOaz57pzsRBMJR7AcS915JqjZM2M22URzDcYeyFGEUUxLSFu8aLM6+iWl
WxHn8sE2TMBj3xkL+R8V3RaB4niIEGQCakz4/yzS+eI8KMCzE1YjiqD4sR2Bcoh4
+kWHxwdkMhDie/bSHkiqIhUkIq6sPOYxTlMmhb4pEjfGUyRgTDCdzBTH3zIWTykE
HK5WXjIr6OutuovQb+mGbZOA4tYltWbejQCdj8K8loGsSqBZsqmnDdbh5/I6m5cP
1AcSBtIf5ZWpbLVqmwriaMnZ+3UfkicxFmdUfAk/D1Z/Tt/5NIA2S6r6uVsskoNH
5xFI4+UrSGvGbuaPQFIaMi2bzvtI6MSCsAcq3ZePjI2Q37vLe+CNZ+Vii7ZV86DY
gzTfygMJA35VB01otxRSxVeuy5jKNU7Y8YpvE23rkAoab5dPoUzK3u48fin9x7rw
unedjBbM60I/c8FuQZpPhyaxEL6wbyaebtV0vXuAvs8tcOlMXuiYfzRv/n8ieMJ2
oRw0MMsBmOTZpLX1tc/9kb3GvtbYmBBsMXALWqd7hHz2LGZv0MMyS9Oceu2x17m2
e7iw+As5x0G/paG5nouhGE/GNoSQ41fE0YduYTTdwGOS95n7gQcMWyZSJcyUpFJo
tPj43J7WVTDzmAcnlDqtRHdcdwCufmMQDwY3MyerCLOCIYO6PLUWSUoQrfKsSV/Q
JZ/9VshVuWGIDJdMpM/63jPgVr61jhfgNL1nZBj6kM29/Nin4OgMI2T5AB36Y/Rh
OZ2ZEDU3+/vfOUM03UHrZIGNsdfeNiaDQNHkJfm6HqC161Mx2W2aEHECQDm+YdOH
1/C5E/bg5U4Z5Mnp892TgjGxuIDwT5Syz33YvYl5nyOJc0Ue845brbkA8cJiqH1u
g74oNrXlVeyU8y5RRlSgb/JkSM1mTGtiZx2TgxFUz18TH8ksOpxhv7PbISk66uU/
8FgEps5SeaECfZS5GWo/C1ZG32d3znUq+h1Y+wJrFZxty0JTpxrawRB4djfOKdS/
zqKoCMrJ4xP7XkH3btyJW8dYgP2iSHAcyY4A8OHW+sQiaofn2LocrBPzv66F8A+Q
MU4NH9HoffY/9l7iqwV22yNRPz/bC9O40k4NYjUVR9In1lyBx4apUCaN1PgQdoTR
2175Se6VNgUv4/t997h80dGhWyDYvACqueyONipEJXkxz2IqefV/5FTXOSrL+ImW
3nkL9MRjCbS2Mg9odqLMR18imsS1SYDuPViqlPZXDtZV/9MjqzQe4lT16hMZH/wR
3c5T8U4SptDg802wNwwpkcOfvBQyjTydvk+AIByxikKCPrk9CDW2f8XKINLt1KOW
lTvYpvDAqHJvxwSbz9GWsk9Yb2WKY+VP6kxbZd7HHjDQadNnSgiXAf0SAa7v5liR
VdszAw4vMJNzSFbEBg0as8b7HZUdOz/C9rtpJzRhRwlqZXBK4+lym/PQA6EDVCux
DdEfj7CpBRkEYzTjF3krxmtE0+6GN8gRJ5v+hCPDHxAwx52bPLi3gtIFG3/CHL/n
xcgE6UekdXcWzBO9Bh+cqeUuWjWBXjdkmEfg6oI83UjHRXLxNjnOhJj4EpyHCke0
2Su9gSOKHvYpPUwDyKbc/QJIt+5QUFLGxK0/Q5nw53ZauUKcoi0HaDRwzjdKWE/V
A2goyndmofIFjwD56nLQkbrmq1TZKm+TAIpz7gx5igAYEasKQyhcG8hWpBKBqmbc
u4MG9Q87puHcZNvqtMhCtK2wd04DKeQmGsPlEPSHoV1PTslIJbnxnzeEG2STT10V
5cUQDcwdTzziJ77GLMzkoAAOPGe6mN3dGnNRhtGak5nS6PtniHxzWLRve/h8TF/M
pKBc7qK06ouYz+9MpxFuwqfGuaolTN8HF509PRsArf4O1WXp2DUeoTRqW7vla+cs
VszjQ8dxFw/2XrK2KS5fsXfJedoG9x9ATSXQcVMbup9Vslegr9GQVOgzdvZrJmRK
CFEqYNfHNKafWJVMX0e04jPALmOCroSLde6wGcWMC5HmF9znLrUM52RTYqGGT57f
1Jb9+3D55i5A2IorjIOFI+8D6pZ2XnydIrPKRru//Lbn01n4D2gmQ6Lb3I9KXf4Q
AldvhQN7GWItzNwX/ozgMfp0BFwmAdvgN1jTqOMytCIPHa6hwVv97HGiHaaaDDf7
m/pz7DjrKdKdAIFDddZ9wKR2oUpQGB84jE5tZ8AayBKDvPURnxHTbc2W9OqFegAp
xDtxw98fIT2S/NIb64pbGn1ADfuapQm2gmpq99YMCGAtv8jNzDqXYqGJ30NuQ6fb
9aHo1xehHjxhhRexgCeT/OUW3muA7fVL57mIaVoIXOSPE6fTRWQ4aOZbmxa3ZMrs
oH+cNqEeTkSr2iQfRWmrmEuN2iQF9poEw5AefNnBj8a861u2M92bgCMDQL6ZiHEq
kMSR6HwIYehzt/LUxfmkyjxhS3JqDGTmGlXcuBwHgwwBQpLe6d4ZBa4kAFjsvemm
lCJPdgqHPTol+DPHNwyfwJdsRq3OA2Iivjvl5x9UbHXt7OOuSlnWEmFzgG1XjpE+
xPng0SdNX1XrwaSmr3yRqr6tarzDiEiw52YqSIto1gU0VA+aT+/4S4w1TCnWXBeM
l9fmLSyYQyJV3kMTri/IoVA6wYibLrH7CQ3TBvRaNQ7ojw3rWuLS97lz5uJz8leU
QygSIjmSVbyM+47zOQRY1wdDXITLUD5bLiRDQ+pz+tTBeoJ6z0d1+EkrcYCXvsSV
XfxbUB2ianCFGMP1fyK0XuRi9l8C0Aw3ZqaNuMAf0WS1NosM7jy/GrjR3U64Qcn+
qTPlElm1oJAXpfXkYM3bQQGRd9IriVQUhEmls3pmQgzI5CNHLvWwtWXC8hTst/ur
YJinh8XWJBM7mP3y06YZOQG517AbT8tWmdxRPA6aYysOKgnyIa3dx1wnnXqenrhy
SEtqavGvwyG7bGxBNa1PWw3TdhFtX5zdrN6g3thPftdhYaNjq5Rd1j6aqYNAeE1S
2tMzkO1CpsfbkZl4rtA0QNkKFVeB5wLmzupYhzVraxlYrHHsu1i6r7ZcK85HhLkt
Wb+EDvp2/BW8NbikDmnMFpf0vHoijWvM35DWzFm+7RnqApzvwrTkfeN9zc3J1wPP
SEVCl0lKQsOMwed+SuFYFtLzXVpfjz9dZow/KnxuWl5H2/bm49SgpRd8u4oQTwlq
4EmjBtdlxEg8l53UhWCl8tQyZdbXpgo8HXBNfGXKZUA+FSTeRbfX0sJrAuq8N+2b
ksG2gSosojdSL9fD+Lj5DJz3na8NwiWIP5Y4q4LaZ4PGZypcHWcQ8obsi8aOcnaa
zhchZEB9aEFWroTUQWegvF/6qykul4+sVSQAxCZDaEAm99tS9n22PMTnHBDW9Ppo
o7koMc1nUI36eLqCf7PM4dED+wqVWqGdZC/W5zGbZV+GyKy8INmN1tx30a3uUBq7
w7f0cugbqN1ywApmsClk+L7Mvv5Grx3CjTiLeR3O5l7FpEywc0KR1K8rAFeEVp3B
8rgV9z+9S6HJNRmgdATw4Xn+LU1xxAx/C9q0vlFb22nEBUsGocgzVInwmPW1hSE7
OAlWIctAg5JPBgbQFCO6WG02x31zkPRWYErz2YJQNJI=
`protect END_PROTECTED
