`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7Zw2n/C+rAb4TUe+tZGBDSlfdfeMeNoMaXeLQmluounSi3SDQhYFppKy3LzbFCy
kotyRvrAVQsL7z+punsrTyuvwlRgLqGuMXq/h/KfaK4XnE8p5mucD9VoageNmHPe
+BuX6K1Ri5DD/knUbBPtBJg1gMeNnEvYSDfbcvYdTcdFo77G8RFv5w+XwNoD1TGb
DdodcqgvK+Ke4GRHhSf3/Anuo98yQKv0LkZoozMx8Km7SC5YEtNy1UYsx9+UvzLW
6fcF174oSyI6PnyltwyiGirhKRhr6Sm2a1uyrINISC2CwRKU0SIRWnF2+WEcf+gY
Nzf5tpbb6F3reGaNnBHGM6BRdVeJQrIim8cXSS7YDzKD2pZJpujHkuTPXKKjorv/
5cZinVqFRIhbcN/XxoLz10CoY9ABkdIuaN2xaX4vuH04yOi0MvetzngB6MWni/Yf
LIRe1LXOmdy4dOxtmKIbLUZI2sGr8AAeMC9CTDhNAHb3rEx5tg4DJLgb5GixZdNI
kStji/PlQLip0lsKdhUt9pi+mkEtV944uKVHa+xil5/mPMsL92DEu48JoTScuJDk
KTA4OvjRgfruntRKU0a2qjGkSc0y4YFFaHLxRDGROctAfPug1GX725EodUzwr4I+
w0IXcYvbbDgwm1VuMQwCr2rDJiVrru3AW7klwXdbMTrTTlwp8TFdOr6Y1auQPQMy
T/NgcQnN36uoFJ3iaZUNTHdSEfixA/1D7Tc+hphsj/KGhkfNku630aT91aesthwi
RpqzjMQOXUsVwLeinWZH6fydIoBVPANyWhdc32/kqFTxsSBtCuvsqtJCyAYV8uyp
MNJ/d+6oVgaiPcTxljBeYmycKjufJvNuurEqJ99BGnMtwUJKzKKd6iqZ9OE8FNsw
tI8G5RjP8HIKt2K8WTYmYyirmNkzEhlrucqVjKuZtf449ux3o0Durb1iIGD30RS0
J7htjsf/oIRVAFkn0ajNDX9zNxStPunEgU7quuSCkItp1k5OdvXTkwtscMLdQgNd
OW6gzkOMHQ2IcHUEU6hTlt2/PBAAiKgp+7inpIxl9UdGouFOt7AE2/A0bg7d5JOj
6/GU6Xvi5ILJqBZ+XJad5pVm6HYq/hJ+kxqMfuY5hOzn5Rzh914VQI0TPCGAlnSW
q47w7cd0QIimfzAg3LHqbBINbjcaKtk011za1CSkx2JkJMg5oTXf3Ld40p2mXiwG
IV6NK00mvZw9EF5/Tm0t1dkKyYo7s72w4VSBulS1Xy+dNuAdSc96JHZ9grZKMQYk
ssLgkH9eI1YBpx5bIJWgsqqPdOoZ9VF82cwP6RnvpdHAmo6vJWoBT9r9vkIfuM2b
X6op5kOjOroZCFvu/dnYkhmKY8E9LBwAgvIOv05whsd5JFYSe/91AkKX3fH8l/qb
Ost/gqXquReLJewEvfEnh8EOy1KRRpDL1u2Kv4UR4FfABg5pjcG1MwsyzX2NIxjF
B1+mPX2t6hNHjlGvWeFrn3C8rfqVnj5RNg+/YEzdDubZ9SXEFhK33TN5wDkYBF9H
3zGAU9kRZY+BckW5kbQNOp/a/gj0zoq7W76Miu804fYGhkvNXVLeliHVBk4byD8L
BZVD6Sxc4EuZ2BFr4vTJFq9WqY8vsMHTRaATsfW3/+KGvOrOlr/Z5qHLp9RAgezQ
RdW6hzIkzDxO2ouaRn4G9s5IheMCI8fEJddjDnF8+Aozz0Ob/8GDhrtbXRTIkqWC
8PJY5HIeSlA9MOo2j2HSOz8NRB/HDf9HORDgI3QRSUZ2NOPbEImz8knJW2WZsNsQ
rVUXNg0bzswVOdKViYGacdw+2KGPjuEgj6GFGthaJVhh/pw0oMPw+UmqjYim3TKC
KbXKATBmORDlSP+CAaRFRLyYz7T8tangFq5C/ts9J1jwyDJkp7yAWpEVNtDvR7yk
QYt0rFaASeVlGWiOF0SZ1Ei1izsRRp3bFwskxoqebtKRs1qyevFux/M7m/AU8HIS
BmrN4e4KUKFW2rWj5ca7dkyamaNMa1FaHMizusYVtMaJJS3VN9PkVkjgFIHehKvm
XfW7ul7xBOTJiTn3UzZ9Kor9QmJFB8hAeBSk3ipfps3kV6CFsSVmT+VxxZd+UOLc
wasUKXNIbsDOPRH500FfsCwT0IU4fXL7c1R5WZD1mwV3bVVjdCAkifRaQe7OqBeT
QkxtJMbh2DZLPdJPRzGB8GwrsYf2nHWjqmmMWHTMjtvfiaP1nV47rNmH/8VUv6bO
13G7ZoL6zMlhr485s5o0MfAs2VRlPaFjyVa/9oa5fS4IHStMeQBV8eIzmAO9YARU
LiMBSNvZklieWaTwHR5irHbwMllR+sTdBlME8dzjy5g22jTkTMAMz1Bvdm1hW72c
DOV1DfI4IAZ+wg69WyyzZw3ERLMAKRRT6u0YDqDtv6iW7EZXWljH0VrP0IdYMNIW
q/hGC3EZu5yMFz1ao6ns4M6c/EU3sNh9JUO6Z0PWoUON1yj//qkSMBrkCDZ9MdYg
Y5UI4zHQ3Sn2vz9NELyf4sDbKFHkQ5IfGXZbFkzf/NSfpgvvsWW6usoJtdzXz2OP
v2BpuNYK5FjUqSQ/P0BT7q8CogBwhqZRktACxpjE/Pc6Glg858x3bc2fNS1ey3fA
zZi8eEujdaJ/cbSmAA2tTPDQxuKWcBG+YuGUcHba8GY0OiHeGLnqCiIBZQhxaOub
jX0SYQwXhLQFIoLRy6mL8tLoQKGmnY7YmLDamKGZcaOhezS3T6+pIzokERufW8FJ
`protect END_PROTECTED
