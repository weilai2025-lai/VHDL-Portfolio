`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODfDneBHP1nPDQ3fYslhW9IyBSMiq62tZnl1LV4NGdJ1PETXnDLQSt7n6zAlzAg7
j+AbDaR8LrDlPr6o2b8wqq0EIldmnK4VFUui6F4zDnXTq6f/iFvX2LAk4DIjsCp9
Q96EEeh+Pobj+NhyiAfxPH/l/stKT8aFuYV0UeMu7hzeTsiruVsiwkeM9tAMx7C7
JUMj+R/agXe8kWIIVvWg9XiXrIOeNEEG0geopwtZZ2SUf+/Fmo46H8TMoBhjsnYD
yK4qjBnXxpQwycmRp/QwUjXuKs1MXmQUFzT5wtibK7N92g5/CxGE5vkdczDaqFfn
aoQg9W3k7XxqR/ZNGieVbHBu/KMtkm9z0iesPLLhXqM9CpS+6NZAIM/F8UgmUdfu
jAAVANikZK65OU9RecG7A1WCnFvhBE9+Eju0Zog4AFt7bw2PceghDJHsQlU8Fd3W
BR2aMnPzD2vdGcgfjMwmuSy84uVpHmzXqnv21/Mh4tM9y00N+o6IeGaeYJJhELgj
v8xVaYUfljVam0lli0FAWMGfGIoMPV+AM2Ba3vgLpwINcglwO4iLm317RXv8kmE9
WrO/ec0Y+M4RXG7o1iGqR40wupTGyPfU1AnAhuiKfKd7TG1Fw1bXsiUhRE1VG5mD
j0hYMKcaZGv/a2rrFt6ljYOZJ5L5gE4uOzAzZ1dxXMC2i6eyE4ksgJdBYw3usLDM
Aisxl0vUiELrGx/KFp8IvI5N5hMytAGly7aIYK4F/NIw2xML2CHzuGtI46mG8M6/
UQtoZjePm8vEPCSe0V3gYVnafJvXfUoFMZklEjgNe2abpuzP0ssnHp8j2M0D5nh0
aspHHiGf7NbTorCQMVqzPrXn8I0xMx6l2YgffudbjfYxuRhCKHZm3pP0Pk8XVssI
tW/eqfqzZDMUfUTTdlYVUFLGG3L5yec85PQ+z7TnUjavQIcM9i+ffcuw4iOgBWtB
/C+KqOInZd7Wet6qhEafifgCFZXuAaDRZqcbXNez3uG2XaY2n3vceA9EM6w55jTl
OHlrAToh6QIYuxM/Aht5AVcqZfrmUk9w4KPkrqovKBSsSwvYm6Gu3yOnRzS1PxNm
EnSAFgYSpCI0RI6dUbc1p4zRh1D0OyS0pw18wVI5ZnEKXSMbarr5ZlhKlPn0km3c
iSyl0Zf9oR4+ftATZa+Ynk3BnLtfrn6DctCct43UmRcX6iHGeGhPkPT2YWKlY/Co
rwkNFJJBw/NWY9tfK2AYWVd7aJTOy4iOcOeULLyWTpcydvVKikc6A9a0ml3Q2rOZ
QEvCB0hyisBwoiuu6CaORgTXGq8oG6fJiZ+ryfOnmZnA8hUXPRY0muxa1X/CdwYW
7cb1DhDsd7Sr3mspFwLMo6nPgbUauG8yiRFNKzsyfMqLTSUnnEv59ld6/+BMC0Zx
786cGhNfnBFjSycQI20nLJnBXc5KuUgcH8wlZqKdThiWAHnP02vRAv1zIQ/8AJ29
aYZdCVtXwQFqKDGUhYocpCUJ0+ezNbwogmiIBeQ79HjD/uhb+JVQcPQ9ejIvcmJo
k+9+cYxkj+c847k044k9QKgxrLgQXt+AOHk3jPHvY5K8Ps28zhZbulbfONOY8eyZ
Oo26bZ+GlRxjTf9h1A0Uhi4vSu3lj4GBWK1IGx22u74l3Yy3a8UfTDta6TPujWYd
Uf3kwjxpY/8QsY5NmtTK3VpgiQ+i2s386Bi+ajbwv6+iRgyDDIcCa/I0i4gvxvyv
8NIXso/0k8I526w5INXo4x3XvwpSaXGzhyMG1U7vEHDUFPmm84edTXc8l5yIrvZE
CkFR3Cz/nJPvl3kgHu4TGng4xtiXzeWJGu2Qqx94U7Nqay4zr5lW5HEe3ndWxs6V
zsqvTfA+F+vtkgEY0VYbc8wPzoFmM1qHD7Wyb7keN/Yf+JGhcsKEsRr8ZmI82Njq
7AktVEJIkSj9IvXVwAJKZoDoctDhkh77GgxceTOEVIFy2Op3cac3Ltef1QxepMb2
c4E+nJQKmgcwacbmjg+SSkyicWlXgBbMd93MBXofjKQjNlkFWngMhswEr3DXCFMj
k+x5sp27UHv09wLmvegFcxDLGL5Q4K9Gh51/FSk+yYqCTOnruBL0A+DowHN5ndqw
lFH7+XJ/bOymB+KO3Umc+ZaaoNBNX0TUmy/X24gOAxuATjj5tGvflUXH7mH6HE5A
YwEknsQhw3rqaVcYBOTX6pPi2VVwQfA7nxQ6BaOguuDRAETnVU1dgjWDcXbkvNCg
561XWEnQuOs6z+J9pMQRS8UCILnWuG2YSgcBZDf+jPgPOscuA6c7hAjWNSYv3Ehc
omYHCA+3U+TY0t6imfVfQcf99v171rxTv0etHqyC/R2vgyX6WvvZEyCukANbMbFU
K0BdyLLjTENcYtwczr50CiH16MvANt5NI/Rp+92ORqaliiyywi1tfp1Gdz9DdnhA
ThL5u00EhmZokQeGeZt9gdBLuwBjffOp+SCVoFgOMlcMphnQiIPoXc+Z4XDxWXqX
5EQKqafZOP39hWEijt8sMkTF7csQO+0bHsxYZ+ZW+eTaczOG9/NAt+z1v2UxL8YG
sNeVuEiL94U+tm3R+Pm36RtS/Td0tQTzUZfSuRVnZtNLUJHKngFw3gpNRB/0kTbF
KdnDhGVJB9LMXaX2E2Jy9ZNnf9n6o0k26PkADbp7wx3zq2+qNZuxTpf8wQAs/WmK
PBINy8EeUv7DYQBJr3Jho++arGFXjClZhYXbkFOQs6m3PwASbh1wdgSl0mBt3tKm
akB0wxjPV21Vx3iGIhOKkLJU2Hhp963WexcKXFKDGTGtSzVmAdm5HmCs5LrGC/g3
p5ZJjpYObD+7usjgt3P1WZAYgGJO7oc1SKfmtbWW8oSBPfS7vRnL56UQ5Gv5jEL9
9mByC7wgZ76n6WZUYSIH52+hJXychbrGYvmd8aVF4Lrs32Ecr8vndsXlpxh09Esx
NJUo6X0Y3TJL4guIocLL1UqUqh2Vcd5JQDP+TnsNnwH7a67wEzcNEsHEbL/3OQTN
VYBIygXjGcCtrnZW7gpwbBVT+0uq22h6ooGrDMc4uD6RFsC9n0fUySlTJYLTrVv5
E4ZPHPIFCzCKrKBW7oazLyAVBbB+8dkrP+gJi+TYMBFeO44tRJmD+WOKGJrG5TdR
k78QmksHeN/1sTkdduvMkre01I9WVTEZLP6U02IVqIwAEZeQJ2dXpeHSmQ7NMc7C
QmDUkQwT8ltWABRu7qP/O2rzApxND6ixq/oZ9JD1DONg5lmHzonXLIJrhdD/adA4
AMjkuclh8ZM9uBANglCtdKOJ+/mc5KOsi7xS72hSYMn8Q2T3HC8Vo48LWtNrY1aT
fn9TtvOZLOAM+HlIfB27AVbbv+inIEYO/wUULNoh7sKlD6w69jI0fH9ZY5nXPLoY
W2X8mqzFSPpnGHGZiskmiZ/ihwGKYbCF0Id+mVWTanw/XKhTeqfY4I3QLgsJgL39
CnevnDFBxRZR/DVeMiH/sVkfSJN8wC+SFL0UrzuZUDFz4BvU6SvuyarBlFJVx8HY
IklwlnF6yZjc5KcirgBfbaBTBGe31FkvFCPg/NCdjNjD3Ll1dHTrgQOsujK1R282
9T+HD94ARv1tCcMD1eNk175XGavxAUjzO9aslNnvXDz85yWT9H3VynEXbGbXqplN
OrGWfQ1YuST/1mFAxg15WUu4IUmh6jBY98QPh4mawgMRGdQbwbqY/v6Qti0ZR0Jr
cAlXide+54kz5mpD57QNOiqLQnGQznXAb8t9pMHFbrPVZg0qd7YvPy8DWr4fSAZL
VpWAxwsLFDHA5FlLLIc+vxLDHEe2ykf+7YcgtO9UzSfKPBDoYuvxcwVPsuJYIYUI
/4rs/964VIReoN9SJHetJ1akRKJj/UGPXeX2eQlz0z3vCjIucT8knUNcraRYZrzw
o8OHDCXwH87rYsm2WgPEFnT4+UNgj92qqN3THByxg6S3W1XHU82pPxW2dEGB/V2X
LQU6ZA/b36ulCpQXqwEzM7pUPpb+ulj34BsCXwkXwlmr6M7A1R/7DftMjtrHe2yj
5jVwAaegyEfW70s1Mr/3Phkx8LG6EyzhSlwvSIVpaRBc/XaZvWCelSevUmT5eER9
WQV8Nv2YuFjxZ0k1j34lwFEmsSN0cjnxuCWmnRwf3opLgcSOVMSdhdagGw+EsiVN
`protect END_PROTECTED
