`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYN+AwE2T2YyfNZgP6QVsIYQKFuFnrwGRz4eUEL2GCNfUgoBt6FGRLrONrB38UxW
4Ti9zmnpaPCvbV7qU5JYIgSUsl0RdGyn0gcWVPdKVzJUHqz+D+Y27wYMCK9n5I5/
a+LXtQ+iykY9yFyiYYoLThAbOOG/FCxTFPyilO1z/kpiR4xcCqNo1NrG/woYjY0i
5N6Mxmvy5Q0TdgQej7Lipv0277BFemUEBRvm4v95Q8G3iktvPI7hrq+XCakvj9+9
x8B0tqJqA3B+aDbaLdMuIh1D8c5F5sOR64fwsTD+CJ4dY3MYfzquNds528TE9OEQ
mpAX8VEE4GPyTfma7oB+taTPnuur/1vZN5o6rpTPJ0MVUrw9IE66vMi6evo2m2O2
SyQITTc60IbSj6lxx1QTnBPAQ705Om4soaVsd0nbH7kn/FAznBF+qzG57ng65B2/
TnUe085bg/5EO/Hw5f07nWaqDa6IrIrF2lPdw6u5vOcqcMg8RmMvsXTQaxlUEXfd
hzHMrEHxku1w7rKtjG77hBvUjUqEkQdbpRutc3FTaXjrYtGc8WBDzB5wPmqf3Aji
u0iuRHimLC/dK+ECcikaCueRzG0Qq0+VhDn/Ok5AsNm8sfNKjsUR/qD3ylz0jGOX
MTE49bE0TJSAon94GfuV2FHERq3RLj4/TtM0hLSqZexBkgKf2heNAKRK/jfLS3k3
KWxhYegB8aTJwkwQP5ONHgUdGs/dw9w4PLRMo1+YA2TE63yUVn9WUNBq8eZrnnUT
P+Oieyc2XnCYH2UXT17h1VWfo91ASof9hTBn8VaCnnIz3kVFxMFpMaIWaa/swm97
bCAyvQISwvvFDcYHvcBu0eEqAvBI4nH75bCoTAEZBpCFsg8Ji/M3K0jA4FfzogOV
YA98B8K6iogGzKuJbhFRB2TTEWCrixNi4oASabSzn50vFbfc4MGfmFkYyjDcVuLw
f77e4fM/rwDpBT6IKzAFQyXyO/oCz6FiXC7kmoiR/TThUI8EQYkHFcazgyPwyIYd
mSycnZOo2UCdlYsN9ojEahFfYeMvEcr5kiaHUbrR2adhEdXeM9Nz7veaeStMrUmn
jEAZ5oXgc7VxpjQ3I72PdUz3HRPlTMfHgcHfUOeeLczinlTlf4Z1v041ZMbRUCdV
xyvo2sH4+2QWSQtol1QX4pq7CV6eRkvvb23NFfOwC59m2nXt045Zupk2sH2y9lfo
n5q+QJnHW/spwucxJNkH3E5XCZCY0w8DErPhmWDX6msmk6PXuSYG35JRGsMcuTfB
EFtG6ba8zHJLGZ1qs2mpt2LaggjmJP0FIOmMNcNDoiOMyV/d7V/dFtQX5Ia9Rw4M
xcauQRTC88hJKFdYGrfD/AlVRvub9BNim7f/aNE2BIGCr3HXQtzBYR5Lfo4dUreg
eA+th9poMQpGcmg9CUAb8dN4+2JlqnTDzm8U0mzry9YHbP4TVlylyYipQg3SX38G
+ptDyTUL5kB3VgslR6uWrqVLGNvINuNZo5LUBT6+H6V5SXJsdiX5WJUOcTw3P/gr
9/yyYhNNAZxvSUfkELR2K4EqltGLBkupE86eXqJQdr3Dh139AsZvl2xlyogaxi1h
B8tegabzbqL+QLPDwDpyoCfwe02YQpJZci5+y1LP0PY35Hk4mfO1cC+0RLvbo3rz
oTzxi7gB+AK9Kzs5jzTzypST5ODj8R5LHmufTMJ4aB8aH7RA3Ud2oLZHaFBUDdMB
G8JUGNCq58vIE3ZwVpLTctxI/kyuUnnVJMtVek1M4cs+m9gwktNEFoQh4hOCxImj
hakwhkzx4MuMNgMEixOHrXIU4Q0ToANg1bzqYjsXyn06BJqa24SMy1omH4ywcln7
d1daatUixtJnv67+Luuk/VGM8dO6Zpdby0CQmpXdFM40n7Fn7s4R+JIEhBADPshS
W1N5B/bGJpW4SCmzXXysl805pOQCynKRdEQ1fzIkakpiDfxGX174K1D5PdhKKPk8
Lm5AcOrpZRZVHDG4FYrp79dwQrEKLBf87CVC58b5QKo8xf+LA9lr49Nonj8/2v4E
9LQ9dKvFJpRVhxc6dGiciGkFaFopij6tzYu35ksvpOWfZdV4U5TNFSM1yeA+SgPp
i60eBWUyCKU7gasT+SDDfMQyoC+mlmFqNRUsm9xH1smv891h7eFy52tzQzDnKwae
gNVC5GNLt8FgfwlD8p4aBoZYVZbu0f2+CVZUX4luELDR1n6v2aQ2MHWCQQi0qAfQ
J3cQ/ezUe6/ETLpJmW0x+nzok91AEMwi7iqm92zGte5M0PWMy3BbrkmQoLvaPct4
nhJVhs8o7rRZjczAh5LuIs0yi4CPsEOHoyBdpl9QLnTKrPygprZ1wIYc5rzbreP+
Fzm7Z7mCHirpguYDro1/n1P9tr+g9vqtVDBD1QgRC1YpGwJbnVWkI5YPwnCKPEEx
qjHA3Up6oKyKR644GXoV4nbJ+vLsgqmBU+3q/8mmxeb5590N8iJW4uaP36dkPw2z
c35+WhJdjG/dbkUcipcUiv7bpueOJWJDLa5EezX29Q0Y3NHVwW8AXAT6rHpsq1Tp
WSTJoZibQEZcYk7+EZZUCRBGFvc3oTFqAezJjFUL2ugIOCkec51z5xn6XCURBHf3
7ncknqgiv8pydXUMVjK7mBGNftvca7/8VEofs8ZJxh3b5o20NtOmzV/T/cMbCac2
4Q7qENuF6Hmt5SHxVruU9pF3Dx/9fAlUkQoBawGkmkPlTbB17KGnfPsUIU5Wv0c8
zDlKeTfG251RfE0v7fJWpTIcC+f6DCAl1huO7yOpA6u2WP15OCKcAX9+FbHMRnA6
y48fTSsgaR1IFzRPHn+cAHumQYP4/qPte1w8ofxNhiiExOx3+o5Jn5QyMjYKaCjw
6adu4vyYsXFcRJ96xWA8sJ/lWHrskRZLoUYBjUBs9ML/EHSD3cwZAsAU4l5B9R9Q
8ym0ANTQWHJi5U40yM5SY6WsMSNKqVL5xQLd6OL5+cLVHMrYrQJmZq2w8U1yKnTU
GtQPxHdQL797imcp7pXcW9cSsi7LINlu/DKS9fJ//mQHe6OkWUc2+z50lByb4zzH
WozBWKdPfHcw6b+tMPUD0Raor/GqE2iZQrIjbIbvMhnZuSeCG5vOFy/iSa7ZrVhR
KxnbhquKgfJcE7evEA5FLQNcfNL0A0BP83zcRsAG3fvqPHcjzujrlIfHja1/IYDG
WU+Vj3wGDdQgDcvnJE0zY6bBCIhsfvViKsOPFXmsXnhkux4LY9HIemwHqFpW9bgB
8cPIJ/LTnrYqoaLCYDGy0TF8PvgoV+IzGvr7YW31F08zreRhXzxLpQXzYzYAeAnH
3MxuK1RngxcITCrnHGpsxHpX9LcyXph1Yaro5KJ2N3CCoRuXDJ6jHxx1p5SnQyQQ
dEarafKFmJQyhy+LmDFofNlAbQeA4KtLoUw6qQrz18ptM6ufipC0Al+AhPP/0Dxb
suEM7nOXyB21VnMvoIcHDGWloJdsjJ4ugFbw1O3FS1r7c/PCCFd8D7EnThkqeodG
hIKeDDfx4a374jtDC6XYlKHnQ8QC1uM3i6ahnc+Ysuab0miG2z5GmPc5gR4pC8qv
9yEYsoYNUUz/A8obSbCKf1YtjKCf/mI3KG1r/UX+HXUh9Mdp5pABzroIrVi7L4oD
q7elKD6DIoDt08LOaUAZ87mKV38/nx2L/Kb5X+4ZYDjAeyLejPccQIfFPMWP1xdH
Urp6cQhgGYxmXf+aixXP2/ycVfRW/PBiAeAnYkzvFm6sXySzxt8cqITFzqiDko5k
rma2oYWrV3feXIEKqqr4dzt4KYfLv6eLxwwIBN5UIemt+mh0SxLqq5fO0UOvBDtZ
hk77tuRbFJUIhkCG2a1moUmx7EbnfabUTfl0SVo+S8f6kwtr8IX4N/eTKD/gjWx4
+RmF1W3C23lzto3S/yKquLZWCDdcpvbpbQf52YSJvCyzELpkQoweT56wdQac7EB7
aFOYRxZVl01/KnZqH4u+ec9cxyovtW9Dr27IwqjOAmHQKOQMQQYePn3G9Yp82PO8
bAmVoHT4l8y2aP9kp9b1PU0lzDkoknbQX3PmaYyLtoxvYj6pCaFpZ6OakIzHajyz
+uawRObtRaf4V1aqxKkhvqXorRem1Uo3tLF/trjVgtzjj30whYMyAO0FmgQQfeDa
2bsmCJY+rT9EevWqWFsBPK63tYUprFTlCPtXmS3azoz6+kQ63cD/udLahXW4owII
0fNqiqzQXjobB0yjRYUlAYI03HLqCboeBKUNfOh/E0+rHCEVzFGz7sOMQesStcqi
B4iekmTPnLxYOBLiGpnRKIlPClaci0k7F0e+dZJ3MaFY1uCfOyWNAfO9BWo+jgLG
XRep7uSMoRB2BgOdI2ahohzxFV2HaSbDpk/gjGXd/bn4R26wJtnAM/hC3aNbIIx4
kqffAbE+h4O+6Tha0ENPAFbj85OBtkYuD4Vusx9rEXIc77qRpiH676XZ9ZPnsYQK
0NBxwIj7r2Wveq3XLTTT1XWfckcIaxVIIqpYOYUM9NLAYGvV1u4lDbyvXgSSMuLw
+mYn6tqiQM+hRtReEmTPlvDIITzNa3ythLp6T3s3gmWwOCNi2OzP7i7yoHkuGc5/
JVIVpVnGkqtKrAuXixF0vcaNkLAFJ36pDpGM5qVnnmxrnEUtuEv/HlwULtVqsky9
CF9e7g90m1/9+uc5MnYAldETq/vB2OCDfBdm+ydpuvuTy0eeX8W6oJ1PnWq2asn4
ymsGviKXhMTiTy1Bzz7ppLErqvmdPtex0buSlhtasz2R/gQX/IeHOWfgkWNUUHAH
XFq+KALOMUbWifFvdbdra/WoTevsqigfx17puhNyqyLiBo/+Qt49jZ/eIslfRz9l
+HZ2HThVNFIorLxRNwplOVG+UEedZOkIv7UjFjhb6LE63wJhe+LOVLqgkg22s7Ec
L0BI+6Djv6vMCb9dVhCqhZjg4pcD9F2sPO5MEgANFae451h4prTM/fGHHgQBp/ur
nAJ+h/4oo7ODHWqYJkNBsgIvvuBAHnr9LkUVv/l4j/nQUMrI1vd8xfCsBM1+EaXS
0OejNjotr+WdqWEYir3ixoosjhwqtqgb73ysbpup2eE/0c8wnKdQ7Dn7b7ZJ58em
SYvLqi8qIgOWP5DIJC+15KlRDFJSuixuVQk8T35kJ19Ij5AXct4R1FqWAPbL6h5R
Ke9c7VZnDjpUNjpY/IT/OZ0/nu497jsP2ent1enG4Qby9A5lypf2EJkd5t714+cG
dwqxy8rShBlUuwOfic8BDg==
`protect END_PROTECTED
