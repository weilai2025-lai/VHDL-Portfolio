`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xu3IKnpi8tv57Pmm+9Q+AT2IZ2TV54kSPG7C5fuiYa/HGyU+Fpax9otV+0z2ktQ0
wr0UHUP8LohhWpyPvoIpaAohOfbmqYCOw3YBfxZ+n53DnJF0KXAZAIw3oaVV2K6h
yktGlDbJPhrG8yq2Lwoq+N+MhkF5Sv9hA1XIMr7QjKJwtOF9rnzV9GDEw+hIp6fz
pkhW38MZNOeYKuT1i4vFyLl27cjUPg1jlx/28NXhKXpGRB62mdsynij5SRwk5fCg
Jy3aTKORcvM8Vgp/6mlzOhlF/3q2/RBD11AiTvO/URXv3ysOM+Wo+p8iPEVRB0EB
pdRbqywMUeN6NYIQJuaUJJkZnoZXBJYRtIz/2kAtzm8NnzYEnRFyjlv93KCvU8zx
R57vWV4oOdpwnIs3P2S36jFTvvX2as5jO6RIPiReunR0RP4Hewsp8snWiTmU7YiN
QDnDLrSwp82DK8t4y0NpwCHl42OwXqHv+KhSQqCgK8K+Y3vvKWxEllvgkblmlEHd
Vgh0Kd/6pseeLjnTkYg5T5QEJXEPzXE1r2UwLKKa4jYpWfxgDT/+DpHWrpBh4Zik
wQaiX8Ii7EfckpxOfxIayxqV35IidQ5ayLdfDgn81POTbOITGsLWfapdt1KJT7O8
5C6j7suTRekAvYksRQPXWg==
`protect END_PROTECTED
