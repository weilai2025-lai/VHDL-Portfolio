`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJIs7XJHbe6C8fj6MhW0io6yB86kDm+ZJvAJb6MfnMNMHIE+uf8uXutjEHe+iBYQ
gnh/XfJs8d81JI2wJWe/zMwicUo37IVP3usB8cluJxcvKP9rqcMiFdvKjW9mUsCF
GXio6feIgRez/F7MwhxZhJuiu8KGD1CBEmbfHgvmp1jCwVHmdx8AruTFXwsgAo0K
fKev9MljlWYxV72slxDEhtafK5qmxLrfb9h5di3guyPAQn/qGkff6EXPRvSwz0GJ
OjL0jbX54JMi1l8Rnzy8N0pet0QE4Z58VozEQ1kZi31RBwWCGbeQkwX4Yc7ianms
aoGblfL45nxbAmnttWSEHCu5o1+ddhTOCfa4MmEb7TOGA74PJGsqqr8NAB2sFCy+
4o/6QIWexf4YEnQkr52LY1FzeIFm7fa1gI8ffmlQ+aanetjQzsTnWvZMd4WBJQdz
i/K9WyWPeB/10/Ahgom90m159atrwPhZ4pW0xyLgKeeLIjBuBmZzKZ8kbTKvAVTV
DbBRDXR94QiuBUqAsAbUVscDpMumNgOt679pg4Fm2WjrUO4rOLJtuD4Uk8SbF3Q1
73W37Oeb3I5AZMRy0C19Ixb22O+NaniJ4aRtQn8Vh87LkpBovYThytqkJ3nEXhu6
Q0mQzXCuz06qos3yDevWYkQ0fLGCuF7KC0Rsn8m4m5jmmCL+Exx9tr/mcvqZCS2/
w1IP5FM8IseqsaGK8gThaLM8TrXzUK+IKIsfnYqsFgU=
`protect END_PROTECTED
