`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
buzdTLBT2O3PQIOvBTR/BwBroJoB8Fmcn/M9LV8ou9cI/8BxEjQKl7YcVc0V8BM7
hIk6vjdTGUPCSSHkwosIjK7xkfbepUM44eL/m7zouT7gUWh0tr2BEivVBh1IwtzK
Jv4B7Z+amxEGydXb/IlhSAa63sPIPUm+1vv7GSgYY0yjPDdXRCmMUu9wSxHeOlVk
Vymw/kEv3lFsgloGy8JXias4M6fnbUcGVVBTmlNnnZL4mxABYRRh8voWewdU4lr/
ln8bcy6g5JbQsWGzmrssqBehwdV7xmNYaJl/U8G/rVBxU8J2hAuKFlOFcywID2aa
f2QmvgOwPml12jCX5dvHSS3DoirX/5XP1Vw+kV5X0+ocqtTOv5BBFH8qjqaGNncG
C0bC2wk3W76WB/+5OHi8Bnxfm0urhyhx3859YbPrfs4Sa84o2BkH9i6PGtSMW1SM
uMVyWEt99JNCA3pOwnBpi5whiANE3X1AY+rii1gtN0hpbYrE7eEzdP3eEsrIf4Js
nAO4o7Hx2uGBvW7Or4vWlVSV6yYE0IWR0KJXTleknrn2KdY52k7LH4rvtPhSNRdm
nV6hJofoFTmeeb0+ZVZXeo8rx/BIvQakA8Dj1gBjRlPoVB1zx07z59f4aTJ6PGbg
3iAMmafrDSk8KmSRaa1uILiG/LVtzyIJhhWiXlgWY43vMUvVo+xCmm8LZgKSthc5
zGVZsVNTjUrKY1ByUG+HSqqg+CCZ6PYiMlyeNaQ4lH/mou+rdHLAZAFG2QvFr9wo
7QycGkzuSqfqwhY518IfRlLwignBurYsIti12AjzlnIMSryrdoIUN00aQsZCVPjA
tDMBkSER1lPRg9LarQiobfX60sVH1YQlWgvs4X7l4jBUSUhSYfdwT3O0BC2BmJuZ
qkGKaAR9QIiP7AK5W0YbIMbUsyqjWsRs6uWT55JszpZcyrho4uoXNwfmgwQ4Pkw4
U9rYX+iMhODzaj7+EvyG/PQcd1HFpBRwZGzFtXtLr/nMCh365McY7R+VxiRok2pR
bBqXSM0RqkQBKmP7VdzoieLTCV4azxo5ox0Jy2YiW/aflY3wCPVRcpC2f0WtTnrk
kfN6zJk/Jf6sv5bpcWGWnktwggaLiQyuPj51y9wesoaPHnTYf496L/5J3BhAG07B
sr8G6t2cC4fDySsA8MBkm/Nmvz4ya6YLa965KvEGFId6vhbZ+5RJG9DpSAAMU8i8
6mufPCQfdtqNFHMeJdvGQ4iSI7b76kTXMRaYqKzdcGmTgDq8+hIt0c5tMnbmHCYz
J0/Kz3WhpQbL3A87d+nfnP4PcEp2r6VnjNO2DuPK2jvrKU2Tpwv2JZE9lrniTVhB
G7Uo9QXksBRBcj9glXPL3d+QpkqLm2Go3zacZiQAgknj59cO9MGXGb11DN8Ui7ca
J5Ljt2Brg0jiiWxJZvnW3uGIgVfCJG+O9V0dj5RxqueW+ToObaZMu2SK0LWL/WOo
9/SE0Za2r38S3CpK3nLeE3N/VQoo1bDETJQQTHBlCWBx4uWkGI3Whwb/KG3c+aIm
DyRfNP3fXLEt5KkhtD3o6GQTmjeeG1HyQyoxwAnAXS1JzTft95uKLohtfbtKVCm1
BSosurgz/f1R6XGIR7JNZCfY6bXgPmqEiOJy2CiRijlkXSzgGb3mKR/dfNNYEdqR
i9meWRo+zhZU6eK0snfymh9Su+5W7EdJl89LIX0BRhRDbpxpVlcXaAhnOD9tea2b
OuWiQlPL3x0eId8Bx5EpWZJq1EWBUjwcBkc6NUKD+lEUVkl+hVt2d4rsFiT7M/S3
utaOwu9zXfdB79V5UW8j8fB01onPd0e+9q1N5t2pSoR6j+hF5gCGpp4Pwv/+7Oai
jHLhJQHv+9Lu1PfqHGjMhAv/jO3W4xOyAXOPQTjSPyhJ7phVNAwJnlQDZKPsTiWg
LAAiF9/GFW6xrOhwsYBdJrw7WnqDsgZaOrYG4K2tWpGLHWl4kuHiDfafDoNI8Bbo
SwngeAtf6S2vDWvr9fgTR2PfH6uUFE3Aue01PAZk93iKvxCGADJvTAvbAkzewrL4
Ahbk2wYmCILDeGeNzPh5vCVw6G4koL8LtuPSRr2OZDiceBDkOkrx5vcn736D8Axi
fErybYpk5BHrgRuF7oMO0SByOPVxzs6PBRamCX0NzV1PgUem2HT3aFY+zri650ss
E+p8jP4H/OkEXmObC4hfsRG1z0mhjTUNAdQTayvgND/YyTiBSrQddbLqnOYsE+y/
f6AX76VBkfamdIiqT6N/OOYzoRYb9d3X7ertNzgyL2MsJ9pS67rA2JkorWTpIb4x
VmKS6lGaYmov3rE9qxrFkwtUrW95yOTP8JtxII2TWRMybujeXxtYbCeQM/0DcB9X
Xgn0YPWwalz7stOiB7F9hKuv6dM/PqMJnsQ6YwRJJ5TDAyjBMZK+RLYddM3g2iua
VyKj4KNCQ23WXHC8O5NdPCE0XBmbucyWTyLDSb8nuoHxHNSY+GGgak/cu/a8gEjX
8egmGSoL+AiekGPlM0iDkBtVtMaNsyxWzLBncoLNSYzrgqebOGGaRoac183UpEvx
roKMQJ2gjki53WaY3kg9gZd9DJFNtwNLQrrDWXM5Hr5lFDVIqUbVkeF3S+EjUECT
U16s+zZnscLmQv/10pCmn7v5uQ6EVyDvpiwBlk7wAAHngZzVUpOagTHyJzP0UJI6
d2FrJNGV/LPpEDRuB0lOTeVzn+Qph1kbJYwnJFCvDze8j29BaSGFL9f0szJ7nerW
5Y/ggSJvV0RBMul4vahPuehFt4+pbrE2wn7SRvRWxRGNCp4vugjE2mrwHgBgfT2f
gOwp4xPbPaUo/ph/7UiPCZQeF8bJnOOkx/G/hj8YfhLtcFPROeGWSCykMMhBaL3W
Qbo7YPiq4RJEm52pvD9VdHbJIwTFLzTHPf+FFYAzedPHB6JfLfjJWbnvwAh7emll
beqTx5lcfrbTaihfuhGhT/4OpWOzcHVedHfnb874KqOEa+rbuxaoqD6vVGrmFNJu
gdyi9CoY9hXvHpOCT2q9Gd2joPV3nLz5H/A+gy7XYF//C+wpwJrUqop+vCZ8/UJV
AOd2N/rfyhYce4XK3j5j9uB9pS3Ti+gMDtFKGtL+uOc0xvDZSLLiu9S5OUGZyVe8
dlYX4EflspmqVex0YPAkBfTdD6S4mG2d11g6fvW2N0X4YeL35sggYOhjS/SJxAz7
Zt2vFaInORyhcV8XiT8UR4i0b39I136jrKqlWYD9oEJK1YUmRpNxOcOVBMRP+Scy
C+lAhAyN2adIsmEFMc/nFrGb+Zyby+y1cpboNOakhPo=
`protect END_PROTECTED
