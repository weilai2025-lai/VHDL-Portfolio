`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PumJQY3QYNMG001D2blMGoVQlRw703eyFH+nAadiLPA8Kckt9TZLNVuBMsU8G6l7
VDci9ZZdZg1mUe22OrBK97J8BS5xLMh15U+2LzYUpYNJeGevgpHwlz5yoiIfjSoA
KvKdQN3UxYtEdheFNjMzL4LnUNy0IZKbXvh+O1vH2G3VFASICxtNODzBzTXzcKhm
BWA0MN2AUY3HLDO2qthd2tuCYj+mcWOWqVKNgMZiJO+JSK+/cXQn+124+MDXFI1w
BsuqcLBGEW9SBJ35qX4f13n95U8BX25H+K0hL7D6AGzuswmy8tNnv7d2MwRkkzf6
M+GhLrh0F1AxiN/XaljasuYNvI0HCCvEZ0vHVqDWE3/xFHlrhDTT9thWXhIdS2bL
744AKzWprEQNo6T1fkBBbC6SAgxu/RM/OPjO/s/6yGzVQK02xwSKwzCtifVBUSNs
YRqqJg2clE/o1pBOcf8KGncyqNz0AHrxc3neqCPWw4JoYY/81FXs0SAtsDv1ex8v
vMM0xewjveQnuLaObd6a/qbjdahyGxy04l8U1atjVSWdz/qS+o4qlWOrqHBZEaWC
Xd5+mi010BFonrvj08oCw6HsOyS5BSRit+dgZKc16IFpuBR/ls6e48gB5KZIZEim
4zUqwOdNNEizTcc64SKhVIdnQCTN25arj/KYnKrBebBWQYelSHhHUhYIOjrM1hyk
jYJ4NEmRFAYhsTdmom4DgQPQU1O3BWTrFOJcO0b8q0qdAcXdEK7GNmWiSUzRO/Ju
QqjVkhRH3sQ3ikQEW6WnZy3yMyU/78NNSPNEmB4oQQa7oHYaeCYAYZ90oQ5siFrS
NYPjgBDUeIkLDyHrZc5p1QH09XXRwBEsV0X44/5kKY9eoZ5dqnF5XVKDOv4ECnam
x57qtojVrRWKXmD/cm2XSixrq0y6diiqB5h/2133nuKFN2sS5CicIJywM9C2kYW6
aim00axWGbop2L/eNPozP4PYjclIHpELjPa1sC6VRM/nGLUK2Yw2NoLarbuKMIlc
kZ/0bX+n5LauV5WhdnbqwYLvq831OT7s7x3Oiup50d1El7PsCuPLfIsucGJxrrsh
xCG1nwqk21r5nBGFKClW9IMKz123Hg1Jxv03zsg+B+TdK++udv/Nc4ev+rg9EYQ1
xcvcMUmkH1PP1uh1pOUqX/uNYL78nHEPx/Q/PbLAAQRhdDCi2tOtCw6iC83p3izk
Aou1EO7JuwNfGAiYmlyOq8WtRRIhgJFur42yNOhJjhjQP6tyV0EIHf6/4XjQNVyj
Y+mA+cowR4dL7gdez+qydwqRUSvP5s9O28X+FMSzHTBQX5cqObahALI/rYCo8Qq0
cmKtIUvzPybcz1xp4iLL+IsYeE5k2VxPEUSmTDBa/dpA4fx2TC9vh2tT2a43cIKb
41CcAEn8GuLzfZWky81V8ucpgNYCrObPWN49D48gV17a8crUgyCeF2AmeA1tzFh3
p8fzwZEdgkKLLxENa6FNL8U/aB+A8RfaKqgLPg5PrrQQUBXTjzgp+TDs++Z68BNR
utwznFvAHNDhVtbe8HpGRt221QZvwo2/kwN3TLG/UIYif2rE8JGpvV6ebey+K54Y
Qeg7OUDKHBk9uRTgyPjP1TKdM86Ec8+a5Qyhij4NdI/zhYztJjgwtJDmK4Yx1Z+t
8H5RGg0tE4AeD74+lo131pVOdmlqo9bVrzUWGlTrIAT7syEFhqcCt8bSIGOQQKBc
BZEkzfFUleN5KMVqzJpuUFM0XEZAr4x3GczJQK6/1LPMBO7EgMOozz2Tj0/ONeZu
W8z663Fr6R71J38XaNaCXS5wrsg2as264h5VzgqB+ArgxrIUsCJqw66RaskkGZm6
rsUjbhQf59P/LVNwTAl+m44Pp2eIaS9csWUxPndhkgxXSV4LFSl1xz7fUIFLSd+H
eY5yVz4iNQN47gT4jlzEpyj2CLes/sY3U0XeUIykTJgxybfXX2bpry6BoIBKJ8Eo
Y3DnVTobvgq8ylB6ZvlOr0QkrDIrKhjNJtRdf3VNpyHfPRKBlHnixqDfZe+tIqKK
izbf76vO63wc1mcmAQrfiJH3WCq6MgbS1Ilue/2PKm+XZeTd81NSADw/2BD2jqEk
xhHW0yKZjVXUeM0vG9r+Fi7mUppPNvKIoMlggvbFaTd8N4boQLgMGE7Ek3cmwEsl
lIQkeqQr8WMcr6GKm6k3RR1uM/O6/14FchomcBtvddbvprwH6pidwOazGNjECFu3
l/rb/jX8nR6V9r9eAOy3KRb5oQ+kH8y0GWlCrPhUKKtAQM2yyuQ+loBl6ex3N2JA
GfTAojHalcFcQOOyhg5bFAfGzpTb0FkfSQgUvaf4wOHUMYL4kl09n6dmNYJVtmi5
MyM6/IOYidQmehcepwsNz62kNl5/8MI/m3UmD5L2z3Bb9XILh37VsRSkFYfBpwxX
IGhL7HL76OO0g3p2D9KxkBCrRL5qP14E9xSr0T4yqXO3oT1TJ4Gl0Ae8/51GbskS
W5eEa20uAOMbJWlkEQSA1z0+439zn9sSLr9/6PZfJiTuStcZhpN81UuUccHca5Bo
OMBl1uLxTR6xIt+Pbzlg5ZftLyj9cjME9UIKXOxwKu/81PQxTEL2SefBzJq9Eds5
1eCvR83v7PstmHe14lo9jDsyjmQemqj//1WSv0vHKvaJknN3bdflI/l/hiayt1ib
HTUMp8BfZqjFX0OEep1rY7Jndoi9MmYSaFQlw58YpTd92H5y+ZBWfT5Exyf3D1MT
nNF0V1BiBODSFsHsw4nRM+GkBJ2jUzCQGAuNq7ZbHlHFZAY0BXFtMzNNM7wjpqoB
jjCg7fJnW6UTvN7wZwBt9qzFjAApzh7pOZtgil6XqYZh+2avQZGcJKU8VOilC+8s
LLBrAuzfjP6BG+R2koOKmfUcg/lchfExjbI5BhfnMI7vxj5XQCev9SC3YOL5Apf2
++8C5cYG4TUKZhJeKDqjaWSRJaf9D+XrmfyLBUMPs8PqH4/QUB3Vic7xeOFi/5EN
Cmt98oD6cry9RJDbI/1hw9EQnKOOaCJSnFuACTerzDmb1VmVgAYo5jcJQXEFU8jN
hBVvUrB9ukhPnM5hzxqL7yINQmZEk0sAm2iuXS2F6JmdxbFrWRNrRpbhaW5Cy11/
+A/ux5craxzy1Ir9IfnoWpT5Y5Ifk+QjE+XqSLyGcyXNiQZPqIYm5UwCpimcUSe2
TEEcb2brwlyXy4yoqzBRt/1qPdbS00zGnlCj57uYbvZ56aa5MGQ/Jy92Kn+2sDQv
BwBtuTrqY9niCeeSJgC9LasPVO3IEbROF/V6/ili7Mi/VRgbJtl4GNJQn+EekmwO
js5sj3rsPlXIFoAOSnvtC2MaIEZ/zWNrZxfKPXd44l7bQJlsUDgnKCv4PGhiM485
hALMIDE8UYT0rpYqy0qBl3pwrUBKTYaIDzfm8G1eScWwr500+x6HrKiDVqWjHGed
D3L5xjrhuDGAe/NDbA85AQM5G8tUYPZAMaSXy/Bzf4uihDaFApolvotqu0pGZJjp
g7z/hYTfWPfLlvYUu6yYQbmCA8h4VM+8E57GtXpuuwZ0zftL8EJ0JxY35crXw84x
c1gPVDsVEnUFP4FBJRiixdokisIcfA2mLOBFY4JwoUu95GYmw0+Z+XZSiUt8wdqd
ZITDrjilpQ0IbRj3d5HZ1L2WgvbqpXporoP3XJVTXp7WPxEYheFtnoYVdZxNgSWt
ABN1O/OY67NzvjdMLFv6/fNN1aaJ4EuPwJhWyfmoRW2Nzh/geBAXJExSAw9ajp8h
FCdVNJjC98lIgzwA2vyuVdkuBPjG+Xwvooysb8b5Qq8drRv2ciYjy9AdAYJVhODs
kVavSdBBkLoGZZ/G2fr+WSteuAU8y932Wi4iERwfVmrsiu6xQV5O94g1lAxSCUDb
aCU50ao3GcSazQvsQqJ/FR9Jc+jiihU8nR4vilVj6jXmPY4yJBsuQJdKhD9pbRMo
MYYX7+vRtuCYpRnd9fiRAYuSx1NDo3t4AQkjqjCcfB2hCGJBD1EdaThL9HdXOg6a
qDXQwX3ZDUmarJF+Y1S3biH2wU5r/iwMHPIy2PYLTSSVuhgMegF3oJVpr+5Nd/Hy
/ePaIgJ9dhlWlzPECjg/RAYcaR5U+fuYauWOsFQi/OA59Ww91HEZJlW4GViEW7hX
AzYeAIYPxme0eoZWi61n69mHp4slOMyDG2/wGFSsQwcQem7Oi7B/Ag1iV49PPYpL
haITBwsqWzNbKkgFmkR80zZefBpdoyEzob/fJYIRub3TdSnOhACHlEa8lMXGXQLU
6KqAfc1KDuOXntqIDSACaBllGn+9QGkAaSQgKGTZwVJkidp+dVrU1eYz8TeQi8K4
3i/GmdYH+tjwGPGlqLXwAaKaEzPLwsWkYgB6fnZcTET78o6hzf1IUIdAohHaQNw8
NlMUDa3OdcSCYsvIk24BY2DyLPeyg9WdMU+WSsiOrE2N8ttRjtQznKLYZQFOtNY0
FzQFVv9gADLEUYzbY4GUf1yQ/M/z9Bb6qr/ibr/uwmGDtsBN4wnxK+6T1aXTjUAs
UBOBi0zoY+tKE4aKDlKD2xtg5aKJ2GH0mP+7WHFQj/k3+cCY0koc3eVLOpw0m/18
Itp94Jh+YLrak3t/3+04LLfIZFEoAArKVWsdOW6D+YbsRMw4xo31/pO2e+CWBlVm
gN2RYhA7mSF/qRtKuGCJsyPa8mYb/TzKy+WZWSRTB6ASePCt04eMRe3coeozRDkx
cCeaOX5k7CFTViWZW32R6jyWV0OI53/70kXR+toN9URpYm0F26SieG6W2gJ3bmn5
YdKFm8ulof7NXhJdCVKQuWyuCWhOsLroVePGs3DOC40E280AMl7dcVHO2nSD7+Ai
pl4ToHeyvyarMXJUo8a+eyryO1MRkfr1/0ioUyphGgLaJUN2pAIfbz7qxCXR+XqC
XvXaWF4XoBn9LDrybZ8CQtip44ttURYl6MxRjxislzgQ3RAHcPmfSlEqGNtKKOQX
TEej88nEqWCZueQPngpMQzgbPaypcpPiii6+R7NTbkmCqHLI5sc+w7KxTwuGNOKH
i43FGb9jAVLCbbgxCZWs9rLsnTZF4FnVJzxV+hOavknqKNczeMvz2MEFoSS0im2w
7YHPf6M0FrRiMnHAnQ7/UYI59Wz9JvMAMzrf2B0hQpG6ykaPZ6ELMROER2N931Td
YjAKtqmqSQo5GeZePv3XQLlmaX3UmbXEbcxCSkotBK26Ak71MYs2w8612C7i7jhy
RQZ1FbIDsOzje2qmfSHIDaOA7EyDRVkKLHdWWQRk0Xo/jF0xrZs5o+hwLqErfTxA
6X2KV38PIIJgMNblTpvfzIrVoRLLzKHjwPFevu8NeJ6npxa9ZflO5qKpUxkdWZS8
5IDwbvCWZbJ47CYUeJwAYDAP05w+TLpIsHNKl+xhyAscbuhYx4zWEkfl6I1hD4ul
pCydlBFfVVyVpcVlWKIojT/vjzjV5lSFeO1aVql9oT5+bn1ktkb7Yqt8rSg7Su9x
ebginZq6XLGPVoHD3B5oUSk3jbEVA6jK7JJROEW3odfnoGvGNqbGAVz2CvW3rUpe
ttGbSKohy3UqH4MhN+zZgg0EMFx6e3G7jPvnKmQCgf+ytg1dVUvEFEZUnDgZ1/qA
LpG7wetoXrTgK7yyejG24yqtxMsSI2n9T9zqlRvmgG9zmlCAQFl6X1I5SmpiZzXJ
Za5mewOOfsmPCIFCSsJPohWUctVfUEw7oiiFatQFfl/RhkaPkTg00hQG5RPyvPeW
LRzFt2uiA2FedMty9nH28PCagzlCnwODNeJFvkWrAuR9OCDVxbDAr3E9QpHWrgw0
vLGWFrldwVUyVoGlpKvWGDDS5tUUe2eonuRgN7Bw51raX2qvkdOztUhAO8qZVSAa
oKHwBhVo1lX+DEJ/3jq27P036tmE8M3q7tTePWjFTHTllskY1l1Iy9/2L8eTPeSv
SfxUpv2oVwu+8DxiNtdnO/TzJPWqFnEt3xL6gRjY1XoIIiZMprg66khJ4STaVMRa
pwMT5km1XXsZsmMhn+J6l5ri6crBwAAhnI/vG+pmOJrtG9ojCTW9GTjTOHV4Id+3
NxSXazpDYXT9kEgCdQVJK9AH90w2v2Y4JJ+IOYjrP1kdDrZfAL3OteRH+WJu1Bag
mtu61W3kVolYhyVMmWk6LeTk55OBSoepONgsU12rai7K5xZRO5FvqUMmsAHygfOF
NBlbcSo0IN+w0fUgaillTyPryjU962G/D90smpoxSSdGj+6laNYGo1qbjRKH3Uv5
LtQpLggV3gWAKCew1rP2u0SCvQ6vTiPPhwi8ur/aAVvn52CzIbD5B5rD6slMBAyw
Jkp5uijinF49IwOld96mtXhVfVbui//bkHzw9cr0KV6UN4kKleTqOvV+oMJrUrEg
uEDiZbQHBThq5BxFM7M6HP92R58mp5DGREJ8lmW7kpN+1OoLUefixOtIrkjRQNTR
xmDzjhhgZG+W0x6qWvJmIVKRzywGtykaiRt5S/XNmyv3W+ggTW0pB7SJ/+3TjMw2
w2xTxxCuTSFy0uqHVSbJDigawRu2rAZN1Bo8Sjwc8AOosJxbv9tf0PBbxD6XnKv2
INBlTHAEHfluOlK/rUZ5vn7s/tfS+ahnZV2PtBLBoaDs0cVjJA+PWHWGs5z5swjo
03K2iT3gPlA0uE3tBzsfe/dRpqfulWU2fNclvImZlfLv6p+hnlka6Sj9zUdQgh2F
GMsKVAyjDLZm2a2Md1Hk72yfEdxLxeaTnltZ1m5JVmcmQ36YxNxBSlBa1Ymc76UO
uwENxS/K8kA3d3Ope8dXO7WH6HyE1NDNO1dHOU4V8jYMszrOOHCbudpLxWrM2Biq
jItmMxxTqYN2hm1jCB6LNbdGliLIb9nDI6prHfwTCcaRIjWd/c//5ZEVAlgsrfuc
+tdTmE2h3g7IPKEOHC/uf082miRKo0sF3uhB0GM4DAE0co66+/vrB+0zJRwC4N4t
cWFv24xmNMjz71y5UQsq/sda0fnihf7A2mS1VvdWgaCbf925ptmxAGv61blYrkej
zWFjkyN12ss3n2IIktZENs86X04gA1AsV5weJYPYkbn9KO+imdtHa9o8vO5EIbMZ
8L5nO4i7IT/G63Oatl77M2sRgbQ3VFCuCP8ApziVCI6jMi2u95gRFgIhw5T3iDsQ
43YhCNUgCjZ13Sz0yCWvTmsdwC4JU5ttWlFNLGx67JcgOdwliS792JYXPHgdbF7S
j+WfZY1TJ2bPHlxVfgABjf6btA8VNNK8u7HosX49N7ZnHJlVSvPlqKB43hSSZIPx
+iP4wvvXOsKWR1d1ZA/MRq272mfzxbsvm2jROTgQer8P8dcPaJ2It5gm4uHBxFbe
GiVDvAqneyQDRcjnmsC9SEWNS+pBkBmzP7GFX6s+gQteMyKFNiawsxTU54pzQmcq
dHBo7MZ91gfLnskIq7nBAIn5yP8EAEImXbZ5hvT9Lq8hprDlG60IV1S4D73ZByUW
3z5ZV8EdoCwZ5+3slp5S2AKKnhbJ1+O8voAdhkHAmD0bLCQ/9NmV5m0lfeG6eysp
iI+a7attNpizfbR66xi9wZFhCg8hKBmz4BPdRGIQEFLG30GzbvNVJQlEEeLbOBng
mPZCqG8GApu0AIzhCsrYUEbpd0PDjeZtIu7DB6WtikPYN7oo+SGINBUW075RJ5K6
ee8xQ0vTYxc+TGcJ+CAHvVyllNonTIzQLbNmN10WYg0WJvF+a9d8flvGeK73aKa0
ejm78JbvvAvCUKkwGClWWWGB1c2BtPD9CCZoWDbRGul73ZwR8mUEjUwYVamxW0+j
1v/qRkRoQncZZTzoad4R/iR7MXtmVMGkrWgNbTGY8PAS+4FUvSSkKoUpOieLfLHw
qj9Lea1ANas2ARQivLQOl4uhtDVi/JyDZuQLRT+ZsyrRiepbVlr6WrJpZANZLDnm
3x79HgkynQPvowGmg3Gur3RN4uJCjNncw0tcKpyMBsyRX7BV4/om3OnRkOHVdgOO
555ChcR17rRc5eqyRj+fB1Vh59Nj55KOjDaAIDAZJH56m6MKMeNtZnDylvJXwn20
ZJpAXA8PyQyS/ZeRc0Hiyj+GLSJu/aV9K03tu8g/AMOhDhauVezM+NIu4YkLCZ5q
OBrOFwp2Q/ObsfM/9bhQfxJSuVg3robnwcJufeVvyTzQiB97lxd2Okwu2zQNJgQs
gGrzpEwj4md0BptfJmOFpxUpELc3uJUgU1YGr1NFMarpErwwFccPltQoUa+ItZ+o
NJMf1yM6Q2N5yLlhQKOIBRTOPAi3pjq2rHyKxovPLsEgcdvZcFRe220g77pDaeNY
PUV6+gK0hEZXqcFWfXEM2XHjJRkO32gUeJGDQS3zXUkKddMaaV09f/5TSJ+76g3X
zLBxMzQImSpyxATpxdzj6Vd4FK5r+rvUtpABvg85BkkErbeTQEt96NuFiN+s4nrR
p1R+XDEh7M9ieYP99IqJKZlDq9N0ovZ2v36hIhfvfqpW1R8Sdt0dd6RsjTwbYSv9
jQjQwdQVupSp7D62RLSUQcMomiwq1lXGVVOZhQA5CvONng1a2zvGz5d5P7H0Mg+D
jETbrnGglpTIDH8TP70IhOYZlsWULcbyHGF+MtZnU/uXshcuLaRqCJOglFw+Oygm
AjJ4ATmWKVu8gXP+/ELMLxM9dXWH0DuMIEOlPdF8Yosnq3S6ihsF4z6jfBpHwbUk
Xw/2qxWwVqgjIiH6QKZFqGLAmcnU+JcrQd3WOSYY1xfyqRU2QzkNX+dAnSQaZL6R
xPwtNYVYjEqqn0tqbhyXS0lutcZz5pne9nDRe9ZvPh1fUbSKnHEd8v9oSNplUnmH
A0YyuxF2xsQlQ6zXw2PEkb56dLfZzgZm+UJZubggC2u8BDF1qBDxbNBe9UAWiNQ9
jQj/Y2YKPkRDfzIyZnoLX83d4KvNTPI9XXxyIM5V1lfRSObLvhgb+YdLAoT9iyGc
/RVeX4FjrxIcpoUrMW+8Tebx31nVdUfx2tCOO4v3TDaCS3z1rsmvzq8S53NQijTu
Z3dNfrzOCytMRtQedXSu2j68puluYAKkfA7LtSo4mK85SmmURLy29Ahr6sdAZCe8
/qHybkMZY4icMFXpBUYHVliK1b7Nwb0hzPM/mvrrmRiJzURE6dOyezpAO6nhO8Pl
HKvLXpjjRutc4IImejnNNvrr6i/ktgBtaW1UyslkIkAmYipmDInMzQxS+yqut/z0
RSNRgDPU3S+URwGUusySDwqoWhLTu8Jmqv8MJ3ig/2cQ/vOBtsnvCjTXdmOo0Dsa
885N0mvx+ziytV+V4Y93hNkZXB/VpLhXsfXN3ogt+yVbHfTQPQCZbmp3kU48JMQu
TLqxbGIyz0jYYY1aODCfHPISriCqEClxtBuqbgTW0GscbUc5peWksD+lCqMsIR8t
GZ5ghGRkYPyokzT1FLn0ImCK+dHPxjUuXbh2DtX1t3XUQwq2bZn/lFydlrLxuad6
AM1G1bD48QvFNFfYET3IQyo7jrPwRMlAMR6ELeGVitB2OjgxhgzrN5lptQKPlM7g
fchBW/zW5VrdOcigdQBBhSoUWyVqoQFK3ThbcRSreZG4QQj0jWg2Ww97RRzhaqa1
fCEhU6fIfNmtECyigd0FWXUlrXQ200gSPPWK6P0OuWMemyPvK2hv3clnGkZNjQEI
`protect END_PROTECTED
