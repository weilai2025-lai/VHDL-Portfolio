`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rsRFexsf6QmGg5+K+EEp7snDRclUZw5oKTb7POGHq6XmJsQfNRhnA+bi+slA2LTz
FK0DWBZLPMMKGxwcEHh/nov0xTQ+m9DMKanbl7noRCUwhdERKTNHI1FtAMVp+bqc
yfHs1hWL8whtqG1+ABPVqbBG/3mTV1BnP+KeYhHDoVd4Yte+eCAH3g8sECfGbKeP
ZCnaJ45EpdZ1Y7tAWGflp2lnv1UwYfTSkkC+2o3H+JLWUzxAMJ0zQungKrX9QRPs
FHpyfUx64cxSO2DI5qDoqhZOzpsv/6VHxQZdti7fmfOW8Zdzy1YoU3Uy7NhoqmzS
kfXQvN3f/MhAqsUDW9uVUsE2Sun9ViT8W3kbnLOzXF7C+BYXl/V66XMT0cxu4Vvl
vGuWAU7JRrVUjjYX4uoXA0dELWViXWZNT+hDYHs2sTPxufPu0a16e6eCcgldhAuU
61Jf+v2q/EFGBfNh5uV+Y6iZbrvPTXOtj0hHvY8sM2CasxwQ69vUHKsSN8Y1AEpa
m0L67DzTf7zWhzZRtqgRlUvuATyGEeCN62gW9MX4sEc8b6GYEN9iBi0fSXMOrd7E
GFKz+fvZpRQlg/NsDiO2IszZt0EjkTWCb9UO1lp9L8OOkIjqr3SqmuKCtpQLsLXX
dwo9EGEQjrQ8q58A6WIJpL1mq4FV9aAft56QwhwNFcuBbqEEXgtpw8LnKkwcgJnM
0zBn36tOzGm9KSJcZJB99xYhbo+Ou8M54pYihabw3Ol1Ffrmkbo+CLT5A6VNRBxx
YC8d4YBzOGMR8ZbfIiNHXCGbzN3PUev+LrLynwfEGGdBc+oa6bFT2/1KpSR+cmks
+IV/aaUdLxRthZszLT+6qZUjCOCnupnhhhPRPVhnlkoDhZOnLhFsUTgXPg+8V75g
kQ7kFe3OW539rRb1s3N/w3t9Cfnm7loLOxgyKHuqEw0eGhWKlzZf97EmCBULtnQy
eC2EFxZRmeXQwUZfU1djo2e+bm6oahalDdhVHaUqtseMkN0J1OEVZzx9pPG10PD+
mSKgIKZd458XOc444FkibqCIDOCrL16xjMauTf2ekNpsffM4CdCnW06r1L7QllIM
1caMd5Heu8g0d4D4bvI4KGm+9sgyd8VwF+fQ4YgeUEi2ohQfyHYHhZP5szGzfxpN
ZhDXHDH1AeEZo9WODdthfr/3lHZ6gg3TZGTFhte0sgKen7lsKoP+Twn6iooLHoGS
pzqfjSvKuJw6ABTLE+SWcKh8ugV6w9dNnH8aXKXynSpviHWrsrdU8Kp5iYmBLYLZ
VvkbmAek+GTt/88JEL7jntxtJ/kPrJ4qV5cSjbWgrfdhSvsib/vOnL1Teas3/yro
HaTideW8MOnhtv4E+GnwEx4T65cykXKK3hNwMGER8Lse+sXSQFcSgym9MWkDMIYi
0N0J8AI59Wb3BwUNwcrkYkdXp3kIQJfmuYisCUcjpnaCsbmyAl/dk/ga+8N7g+Cv
wrgZLKfQv24Nd+duFIE49ePSZlwk/uw3xjpfFDCvz4msmc90XviRgC3syxsjEp4R
FlR4kuIG4O4LxVjBsjXxRVySeYmTO0Kfh0nPJUnR5pQuzoi9tWlIo4NL13ACa0kD
Ni8iiWnRfGCbqIMOqfIsdlc2yy5FuNzH4ffboWvL+czKYteSieue6SCJTqzk6q3m
u6XDDzjHQCOunEZ6izKN3uyXCz6ZbYN9WKnqWsJ/9Rrz8yUlXzHwQvHqUAuuZgBF
`protect END_PROTECTED
