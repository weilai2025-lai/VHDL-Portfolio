`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jcDiKRMndhWiuaufJ8hgKcvcc1E/IQMumu7OHGrYjSgszzt3Aa4Vq9TqlZNLjbI8
VRpXr3c3e9YRvfPxlpV7fak1GRC9BjDgclTepn5B7IfqluIUBSOCPKkFrdoQOeq1
FMWfs23m+G2EPJm5dPSQgtj2VvaVSY3mTfsSpkZnZYSWGeUqps1S1P/bUr8D1CxA
bFNJ+WNoQK3J4rTZf4WwLCCS/IwKkNdx/4zEXJJmY3SmW9cWs7oHJYa8A+SgSE6D
5Hwj4x8dJwHl8iuk9Ht0Ah4Jw+L1tME6CS1hy9vKZonqVH8CINXNTbFC+rKaB+OT
ZOqGULulCxdoIUKS97JAMxGxjYZsacgw42hscbC8BGEpDtwwOdNWu2ICNoyR2epl
QHdtFYR1kwEjmHad1ySX43+sYbrR8ggZvJceUsQjtLdE6tnVbpqFklXLLmY8Gagb
o7E+gwOYH42bLvvCW1o5mCz3kfyGrX2ew0M5nbnKe1m4uHpjAXs2bTTffCK/BELz
lh0UAdzH27PmV424hkHqDpHWy6RcJwbZoK038QfSMNV4BK+aMVLYT3Z2r31l0W+A
Ai1ON57JVDXAmhBY9k3z4ajHEvttmwBJfTl6ZIZTqM9s36/NuF3j/Uv5MRjJMnPe
vXNbm18UCRacAy8aWQERb65sTm4tn4fRKlmM26c/BaHs1tnYOhFQOcDTXSGSJkCc
p4smjM72uA1Rv2CphxQONg==
`protect END_PROTECTED
