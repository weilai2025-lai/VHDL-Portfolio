`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4etefD8FjNdn4/eZ2vkkIEsv5gnJ68TTlk3TYpk6su3Yb7dK+FtGpOOz3jIZh3U+
N4sM6OmF7kO+4xSEG7AYINtbhX/6blkJsvwQfTtc/xvgbxOKSV0uQEpaOrbTLFcM
tY78nZjLCQvqT/J4kQsCc2XSQzfQRI+HV1I08g0WiwdTdti43ZBKxGFrokfvP9Cz
EHs/yLeKPmYJ85Blcl6uwO3yn8cCpWyKcZFFzaxUp9ZBrHVkwLfXAI/5krayF7td
UtcDGteMOMCTS10cFZZP7LK2ilryu8lc8cSW+OgRpgb+78yw09QHsT/wBljiCJvI
rquwKvd3W3Px3Tw3TRB8+REdFVKt4o3SD9nehZ8AgksFJC7glflaz90DSO70+bmf
ECkgCUOEC1TGpnMUklKkMVT9YCBe/iKyphAs4sM8xyHOCxgnmVO+4DDO+G0gzAG6
vznjMOxMVzji0R9m9OnvSvj13f5uCTI3WtvkJdd48YuOh3peoBfQ4ZDJpi0h1X4n
kWD3ao8kWl/lNFWIjH5SlGVkHibXtfalx5N3wQToHkzyDJ/Fn4lwsQoMe5cz5W+Z
c/nUZ5seaZMylhLqAmV5XIh11p0GFucYwjWjnxFhSvQo97F1BM0KOKA1zAMh/ET0
wSlaCtRGRMFu1DYnI7rUjcrFr1ZVUkVaaf/pAKTUnFa4Wnj6l4yeb6awZsTJ9EKw
3/jdeXgNTRMovP1jaE1V+AlBT0jLcfemAzkUC+11vTGT+j+qI3VjHXnlq9uzL7KL
hKMgdoIXCqSEVLedaKmE5qWUoSorahI2/NdYzh6WBfVxR8UMDdIOy4m50yrB5WUN
Bqh6qpH3oMOl8wdcOGxk1yREOX6QEHN7gU/XaJvo8JqNQmkSlmQ14n9R1iFIZwTB
9LR3nmaBXMyiCou/22m6ojHLYtKDO2Dl196cjgxYDa+SASjYDGM0whsc7K2oGcz7
lh1ju8381uHEKXlWW7Jo3u8y/W78xQZnUUKB9MqyysRKB4t4jOZbQfBSeF1q9Dn4
im9SIDXTH3ppqweQI91b4CGslMCUuKtrGfnajts0BxCJX8ovsoIU0E23sR2/E547
nLRvWEzWY9HF9D1Rdjr0BywhkxynUP7GLro9MrFlFKwBnSWyKAYr6uJ+l4DU0iYq
XFdtEGnVRytHuYpeoMKV6QO+LawGSBT4AMSHw352I+o2Xiv5afRVPnmd6bUE0WUG
QKekO50Tnfj/nmRShM63FdybSdZOtwzVMchB4mp6L1niywbCIaDfsGx9f22NaaP1
k1J2NCCV0agL+pZM80FMTXI0pMMXCERN/4DewG5zN9WVafO4I3BTmWLMOEoVE2Bd
kgkhL8Xmhkw0ZcgvY018Gg+/GrJ7HXA1S8HJ/pp1db9LOGNihuCuJoZ6v8BUemdS
9tSiUMf8Kt3cSyE5CX46FYvhALkWsy2zvNJXwvvgue/pz1dfogfrhvb+yXuWzVlw
42YW+JZ9lTQd54hOU+8hl0TZ/yvXcHCWXeohrIhrxHA=
`protect END_PROTECTED
