`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+anHxplzvleKZV0xGeNGkkk4nabGnTo39EHqSCGG+nvrcz2gUkvK2sVgbQAbHr5A
B+KyVfu6SCCq4SYOAnSCE2CVfBJp0yUsWi7lJ21GE/pWuwdqq6u957VPBwRs6XWU
5pMb7mbcAIF/nG1cxUm2hE94FEyAgp1zp9EnWJMG30CMAYcoFi+B8GCk0aAImtzz
+XV9UQ/8skWku1lwQkCFnZsXDYj7qYpBC0AsMymFXyz/MVy9u3n0tF6LeUViw7FR
8bfr8iLC414zymvGioiog+AWCQrSczv3+LqBNIpdTEH4Q5wR0sFE7PXM7Qq/J1f1
syAWCv8Y8h0jJmLzUChNIJ+vaKRdljydZUVJS9tejinFh6Kde5Dh503llAIWtbTK
LPY8I3Zn1KxIlKIW53Zz3LJlzTKalfq6KQn9uDrxnrnZ8tLCsTiKWDfhOdzjlInF
1x8/Yzr1YCfRCEmY0ifAo/Th6Nr7h1DU4P+khMe4g7gc3GK1u8kWugfYGnsTYiEx
5kSBo62mQt0LiOZ5QVJFuOUvifdR899BGThjtWdUM0M1uY6FamdG+7f1lhS6tmRw
5XKYK8SFVqUXdSooULhfRg==
`protect END_PROTECTED
