`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fsHv3rKP5FWwu7tu9Oj/orXMHIc3/LBMPCe4LnZ37I1SByvSxDaBS8UKzJR8fS/L
uNg6lN3Byk1R5WLB4CiEAeYX7opyFGllVwFB4p/DB9/LFaF3JH6e9fh2a7U8plZF
tuH+v9dzvHrG9LlrCKvI6qVAnf2iBdndOgEVmHMb2G9EzGGkqqygW+6qYV5vp7g+
DLciX9vFDfSJJEpAIzEeCveT3fx1+2s/3831mbQJoO8cBNVmluWS8u6vqmcL5TH/
82MxgohgOFyXKG1Ln3OjaW+S+94FXT1WX5eO7CWsadgVcoHI6hwCMhM6WwpDN0+3
vUNrnsE0TGU2/ruNjNIF5TVKyTYnn4syNT26q5F5xdViNmC7kbMKfJygNp3loKoZ
GuKUcc8CjBsc73AyGmkxxjLfwNGkUU1L0Y4visoj4iSaXkZ0IJdrDBsomzBkrGLh
U0o4mLBoGZM0XNTgFbUJTAfePBYQo07eGO8/YNfIcHPyoG8UTDbQJu5YNjntcNcQ
mbqSu75WBJy1e0E7+QfCFdquYgwmeaqZv6JL+9of0PmDGZqhWJT23/RBwB/rDzrD
CgM9+/PeTJE3cOfCogiO318b0ASGSHgnHiHFgNM68pBPlqJic+9njlzNVcrKGAil
LMmJ3ZHLrjmvlix+nOLLh9fkjRBmwOopw+fBqh2l0hvuibUJEUErpNb/iJWw+Q2V
G7AGNeFLWP8YmaTLw+U7R1lh7AofrPsGGOPQn9nxJIYp0C2J7b1+ubjOvNjDrfxa
KtXJerMQRcAiZcMWhSK6Zub3etQvv3erA4IGynAeObW+ibNcv8uCPd/LSIEhD9wa
C4TIrcpyepBDq1tyVxc/uTIRY+vwt5kJiekbONrjY5HT2kU++GQVYWW3Eq8z32J9
/zVwTapviAh3pvn6BTTiFRHJf01sJdZXgVmPXZJ5YMyZJ5LAdCI3D7IUL5pkv5S6
BolgGRvyxj3zcEWrg31Trr1lZGBHOwdSdLvLf6u5AlI0RdiQ5ac0wOtwHVstyJm3
uORBPseJukukIMPYQRDoebDM5/U2dh5JLCzp1RyxaRLxWLvG1/LH7H7jxPoxKIQq
kPpIDLehqeY7nzpBwlKg8imto37TZIMDZXpIkO8o8Jmnh1JTO3pBa/7Yn4qS7MRa
dOHgNH3+tEQaG1Q4Y2iCM5ifhB3oa8Qr4tIJkkZ0NxCIVEK2Bpwg8gZ9HIlSOisS
x0wHamPPeaT1BlTdqTIQG8q9+A9wEmT7V6GDgsXlJowfP4KwsUteijI4jxTdftSF
nV0Mj2qBnBlNfdbtry7ZiMP92uljOG0z0MhVrAyQ/XeyFUzKm5Wj/LnJ69+g5qtA
5569NOwTvnKbsDeyH7aQxWjXdcAHfuXkvVITyAcZOXMEWjXzLevupzlbjfPQiAd+
TUiR1oZPdUO2zYG3YB7FE19WjTySqxNqUi+coQMh6zZdLV2+VcCAF0fiu0DBVm5L
ulAZr9IXe+W9t6DFzcFUbXSP8rahu2COh/6xQDfPS7lh4VYRWqpXm3toTWKM5pa4
nKTQ0Z9A6CGomIEXX2w7s0f+kq+zT0FM52OUAUbjYlndI8HnoKdXI15kbzkMvPJp
Bjlm1LScKhf2RvjvmsDIeBdSu5aFZ5BdbC9GVq4VsoTVcfB11dLSbOl+DY9Q64yb
zmbcGpxdnK3TFLhyDLjg1psq1/wJdv4XX+8Ajr/dOMf474lWDKuJGWKvG4sP30gy
mOIwOEBKo3lH73y4c9hDsKspL67eywwRxJGMHPIOg8Jn1rgToO0wLIOPKMxWewGZ
5PLnU6GcA9Aqtv7kwwjTISAyWAlXDbGv1QeEffk46NZMRE4ZMonXxBLN+ga/6pm2
TMhNpm0Yyj6wcJ4d1DOa7I3UI8VVoga+k7eSvQDF/OqMNC99BngzmvT3vfkqpq9z
TTlI1Inai0a2EuaY+TIUBd7lCSW5L46ChNW4Zph6NaU4iyQ/4Y2ZVBGz+Iro3aF5
BXDqmiKb0RyW9Tr7+5zoeq4SFc9GuSdePtmsIQkaLFIg5SOHSR+0+FNtYN0jHfFP
CZXJGYMT/C7bgffrIUNHiizI5qpeR2jWy144xKv9wF5SRPrz1Fh1RL4NqNlxvmCv
Kyxbp+ezjAVwkEIhLXhgzcZrPmdPtNV1ePAWAG2dFmPhHptX2kqNljjBZ8QaM5op
j7BocNS3veFj04nA7Qx3TrgK14T5NxXNN3dor3y8AeJBFQtEzisuuksgR/e1CNnf
g+km5QBqpVUfluLcXcSL4uiXbUVmFPEJ0brJbTDCf27VGrOTTHjME6yRPZRup4eY
A9oCFPM/uC5JLXJiJ1iyg734h87pzG8S2I6NEUL8Z0PvQZ8g0h0FT/nlVMbAnzxy
+XYYoQ9TkqUsZc483TXs8b9wI1KVZCffykf8Jz6Kg2ZqkW0aFUwlJ7dZfTJXUB7L
65p1WirMXXab1ZrnwT3RET7qNnWcIH9BOoNxLh1rwsR6DlTGgftGQKxsKaCIiKkE
naGZAfKF1E1M+pQPxIXfMMOzW+xTb4F55iXQnaAwLQCCaMrKF1mGvkalNbo9aSFR
2LecQDqbaqmDMH2yaIHumlrYUZQ7CtD6+VWGfvSjXU0NQdPWB/TsC7w6s5JNPYtd
URUYMeBX1aS/65IqpS+cORfyrW44kgdsQCsb4HkGm8F6+CoRk04DvOqCaIWBsGoI
UpkpjecekVRJQhM7/poeLjUvqkLfopHcySniFQqNXC0NwQOgWb+a738R9mynrMcx
R9jNrE3zTalrbIXcQ7CSqWTOD3HDf6y2bToxvTRcz6MJ9TE116iio5xSHiJLaC9W
2Rtu/9e6ZmO3/WVeH4TCGvA8A+GBA5/gjcIJQVCIGiU2z8j+b8qffkzcBYLAU7EP
ctxrNQmjxAZu7dYz4n7f0DC9jjKKKJVfzjDAPOgTtvah3miF2mYFKbRpFg9OkBlS
FyIaR+CoVR/ip2Xt9lJ/IO3WYFGJ523JSuG5BIL3yUAmm5Bx/TyU2dGTKCU9CAks
UqILZ0ueI2NQW+ofPi50H7gUE5yPVM+DoBIX6uV2je3wM/2qM8C72Qan6YZbStcs
SSqOQJBjVVgGr8J+sQz7Sd0vjEpUr1deQtbSqf/3mbkyFpgUfu0kv2MpSYUMy+2D
3RQG2zw7MsRq7M70VS4IiG5Qxq0SHqaMjiKiI/P5dMmduGlvhKfh1oUXN53W6GMl
J/Dx1+HDSX9mD0rUg/ljNGgQA8KquTovc3z2EtU/L6aRquTnEIRu66Ojz7J1Ho/i
WQX6JelhguHf/urFmffgWDWrCkmtMjKE9barReefGwVaaTkTRHkB51+Zcn2Pa/Ap
PieOaTkoXUq55gOPjloo89pt/bGc4c0BdOjcXU0W4I2zzElOGE0r8adMQS2a+aY+
QDw7LxYZhDvQSfiFR+MvfoDXt8JI19QiTqI2M8AsM19lF1xAU5hDt9lTUXjZ9dJK
2w6t+LZCnYkbdyXFl18EWcSpxAL6aV1ZR7L+zBYERduzsNAPL9B7yu1l29QTeBbt
dF2Nnf3ORHuqjWu65ommcfGln9LTbsUmXtsIGY2Ttoa0z5JIlcAQpPIW8bmtco8f
rQzRO/P0vhFM9zZIQXUDhpAiAaRUOEbODNwUOv7KMi4=
`protect END_PROTECTED
