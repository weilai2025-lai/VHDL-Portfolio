`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7N/JJcXuFMFpUrT5q83w8tb3PEWBuYf+QgoyoeOnZlsBz2YtYFjMndO1jETfvOg
xiZ6dtcudneJXLC/Dwx1pyNQ8d/cRzxI15KCkBTs3T4Fw4F0SMeGHBeucfPAQ9n9
eCGn9u3v5M267kHddeD+FuwL3U31IAAirvL5DHzxVQ4nMKDxxFPUljV79MwBbA5P
7SL9Vkz2mG976jHtq45F+MSxqW9Owu0dt7/74KjPyw4vHgOT8bJ9fMuZf4O5FM+/
f5siq9rPal+tcmL62F2Rldh5qFECIaqG3WAaum0Lj82ImSP3uQ9cuSx0YT6w+XcR
QhItm16MsO8EBUow3M8P17V80XshbecYD2rg7qpSyzH1vzsM97cBGON56oDrNRwc
HWCDzZ7/T0MdJNiBVI4tmKNFN7LSbM9bLvvOPSok5tJyGeTG+GEVqkK3tdzuk4rq
hyZbrub/G83A221G5AS2D3E6rUlQkD4it+4xvLu1qPddV13Bd7YOVTRmUYpkR04I
`protect END_PROTECTED
