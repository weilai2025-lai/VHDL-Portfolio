`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gBpQCyi+PQBqeLjAbPQJaqgwg9q9slJ8VyruY/tegWBWHrjVAjAGqzwaq9ZGjyH5
claDBP+S6E7udtMLY3SQ52v9meqixp59FDQ4FFKAdmi9EVQFbJgK5nhoBaagf/1B
YE3W76sKbMuPi2vjUjnvQI5soB5nTfPobRyqDrcFUtzB5FAfb+Jbwl5v3z+D24D9
d7OkCZ9+lOHfelz1dQAgvMJra8tIdEdCdHLKtWx5G6laHgSvNzRAK9aSI3ULoTmV
ULO9b+tQr+VhA0gwpUJhlsOFhv1qE4P3E+4pcZSht9rTF1LRy+XfE0fKU5aqr6EI
BQFORD1TqLGV1yCCBjUD5Ygf0PKDnsVQ9yvE2hzi/9KN8QRMDGP7vJ2s5K1MIyAR
7w/DCfQSkzGvnExNQf7GFOZhTGFpokzjA0oN7HLGRgFROxBYDypUe2otbV0d00vZ
Q23YxPIOsEZ9+nibbdX3pkWwikASrLZ9C/FXlH2lcvD0BUL8yKBLao0Axon6VbTH
29FJVJwMe5IdkOUQ2farKyIvEREbuQTTa2SrUG5aB6UCxiBjAI0MtmrjxdtmmTr5
ePBKSEajYuTIBx1TrmQfkb8oMHM1LKmD7d3cwGeUOYoBhdwY2YhJNcjXwF5MjDQ+
Xs3q3PbtKTTV1P339igMvqbdtFZlXXZDvY3cFMAPAF7FKBcABXfZpyfnFx0NsHiB
+C+pbZllE5IhFpW87xeP9Nb7uXmsYcb2vH95Xb46DYQxyEg9Qyca7RWWGW8QAqy8
gIsmuMrHuwfPodK3kBBwzz8dEnvzBjN9Tb7X2knL3ULOitT609251lShP5L8rgSd
H66c7xvtxq2Gf+b5c1wjzRmkuX92u8FuFFfsPhyrnz6/HrNc/gmu2vsgHS2hAO59
um3g7RFLzbXNdzU9lOzU1Uozz2sfXEhbU8UoLrImKgqYaGPd/dKxJgwC1l5RuP7C
QnUtL1Av05qJ9+rSGMoNP5YSGvCy0BciBuH2eNcPlTL9VRjmszkP46NFJtJDNK41
27yNrIhgs4x676P8XBeA6sO8T4siCidLKBcfNzgOjIYmB5Q5hd7zGMEVkOy+t3UC
jLIp+gZjT/7H7am9OIQr5Pqctog8HhATeARJlgj3Yz/93nKgzo8WRzILh5Q2FQHI
fqlIs6OOdMcyBhMou+srsPfzST1Tv9042ogbUNTpLfEAHV66cDkfCZsoREVPIclP
Q+4plgkh+/02MFPF5JogJxgJvQzj2SsojdlaihXSiqgIqwixsgmfOc4dZLFG0Qk+
PM/gN0u8lWKYXvyLedCrjCD9CW+9PCgezE83lBhIsvutWSuO1N3AwBjaKPuETx7M
ZpQe9Tv1xsPiNw8Y+WvXhFoOeLMxWAb+xAJ7MnIR15d0HmB5U6stPU9Zk1JzQAQk
jo9bNS1jnt/DtO3GXahi+f+blhNBiJ5i4PbbvXZDx8YVK7CWWgpAu5ENgpZhUASN
+m7GGzhuWrI8paB5ooo89dD7PdW2sSPQgLcxjbyTzW82LlIlJEdC2fbe8mrUEtqH
1f7khJVHl24qhM653R4EbDlvv+m/xzrzVLxCrxBEOWIloJKfLUyjR9BzouwotO13
fYcPCBZpDcs1nIOUgMmcZDhMRoT+/gC6KZeqIBfxOBarQTep6Zjo9KVIFKwq7HUF
LLv8jtoUaVlDy5xSMchDKJiPhAd4sbftWzzCeKzXYobQj1qY6GB3ioOLxeTXDeXg
6FSHvg94g5snwkub7Zr77OQvk4kWraEbUEJLX/71Zqm7ZRPjwRwcgyRUF+tHl966
`protect END_PROTECTED
