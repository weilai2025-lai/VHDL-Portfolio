`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIz+y3ZyVmWHDsg9aHwcpJjrkGgzd93aDI+qhA/1CL/s6sPy3s4XVLwX2RKkITJv
6Rq68abg+jTOImv/pKNb7HtC1mBc/iVheEUj2oB9WVGKSsFLUKr72LAQ5L//0EHl
zGtMpjQyj/ej4L9DWP4rxldTeeH0pBE5neeCG5ueqBIcmxe2lCCLFbpNbk89NENn
/DLHhEmvzT6pVyMhknzLWTlAUAd3HRW/lEau3fq8ZOtkQbMGQeo33dk1Y9bOAoDS
sDjVa0qYD4ALrgkfaDrg6MVvWYH5S3Iqo5WeQv72fNLmQojojHtWmTzXdlm8jdmJ
vhys1J7EEgLiAEHuKollpxC2UywV7hPTOTm3/6wKbGgEKi/SJo35W34O2Eic6Wpi
q/VAaa8uPExBsIHVDO33QcQOoUPhXB5bsmlc1RjN4D7KH+SWvYIZXOFPgA5louhZ
bH/C8TAL57q5jkHX2/9uXM7jZ2pDoLqTSsKe3ekbfBgSXrK76QaP1eTKW22ig+8j
uXlQABMW35iMP5Xdi11p8rv70kUp67d001aYcpjVM/g2dVFymwof74mtEDzwj9as
uguRzNDI9FeNAH0lF9LmiAcqq9wNvVoo+v/bfVnZ1WXzIPIOdFhL/1D6DURmcsYG
8hH3h8wof9BAtTF1sgANmleNKV7299RsgWacHy9ipQh8lf+MUpM3BJnUQDAq36vE
SaQbmkMA9ks/8v+FAZ21Qi9uE5mft7Bx+fkGL3T2OYPxzYmZReW/G3AWBsz/ho5D
BxbyIGD2K1/AdQYF+ufCl+sQFVkDtIuQhD42XfwQpWvPdm44djq2NMZL4qRoLT7I
DI4pAAEeHZATjiU/zqjuxn2wwWgUfQc4/M8WLArpfdFFy/R2/p0hIoZnPf6PBNZ+
BRMlaEww5DmQuXEIP7lBfhXsSyII1nSmdkXiLykL1oiisibuOY04N8+L9nOqpipE
OTEMwTe/U9XYx7I/ZDkUEB5NNTOPDczmPXAQ3Aktjf6ylmDfQ6YEJOIEU8LO+k4Z
QEaPwWW7FlITY4HTpoDblkm40Q47TBow60jWtRXQzpRdGjb0CPwzF1B1mvl9jgz8
fcvzmImLDuGqUB7CevFY02/o6dM96VKJDXvGPgAXxrkpydFB8rBAoEXgrf79GQKw
Jl2tmBsQgU2eJoUHnkVuHN4sW+0WZRm3qwsJKDniqdcT7M2VDr7ofLJGKlDjZ38U
vk5NYi3LS6+hy2n8rcgzHJ25Dixoy65KsEiQWZ4x7lA6o8r/8WiFyL7EZhsaJQ6Q
02NpCgZTea0DJ5ssM5cLONX+MndUB4PuNrk2ZsHGDbSIH4JftZY8uzvXYsLtYISu
Qr5rykNh6DOOPApwJ9P/b9v/lzyJ6NnkKs4Fr0DPKlTAFsktPZYUNT2/xm9ECkfl
xn8QjOm0YMBETrUFkg+dys1rD/Bnr+fPq2Jy59CYqwzDe/0Yj+/TLCMfscVWTNfL
BHHKuMfMwWznugFYAnCSLz5L/fRYln+Ik691E54lvEw+UWtutQ1TpI24bnuXVWul
kJG2O86j54RXjC5RZbsQOdqiBBcqBJf9NRcyJcerBilyjLJ9yOjjs2YtQgBPrwpa
pDdt35lak/j8q2xcBhfmNh7xIfBUM+mlejcW8e3lEg6KxVDQBqfJQ/xHk4XA/Zgr
sbKSR3V+ZGqwlTdPgJt+v7fxEQsTKnei0CUqLm7+fRQr/2kDb2DrEFbLnlMWLez3
MlqKBKb9rnenPIWAfSgNwanlokfB3oYy7mAhFiJXeShZk27ibfgwe0UlcO3czIOc
ZiVw7tsE3YMiSIHX65OklRb7jANbyHLx83UrKMLqcQN78FuATISMlzlCvgastLwu
cWKTFvqhe75nhn18MiJZzsqQiUtScUaB0aOkrhr4RvhhWclLHdVQtnvx0ceD8mwn
HhjjZDJXT7FEu5Q3LQ2PlEo7PKnKSF64jfB7K8bUCOcK9GvQxwEg9sVaITJJrCKw
y5bi1LAsetpXOw6xG5OCAkqCTAa1oFaiqJDQh0eDy5hAXRlnHrobXDrHeNhHeIgN
BxFJyv882tkdY++VAlqCYHVY7j/kucTKIn0iAezDbn6UcWNGflnUVzXRjDhMcZPQ
aLB4shNCGCOPGgW7dn5xlCXCRNWqMXbowybu3fZth5zdsh9nIDzJL8HyzYgY/syQ
vrKtP9Aw3v84SwGtVDBvOkbD5k6PQdI7dwQhQf3pB7+v+KkKWNqAoirMhGPu9X9h
W3K+nMZ7QRRVidUgjJO0V98VXO38cIkFPJMNCjq5gTY=
`protect END_PROTECTED
