`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHrQJ3NkIplJZ06fZgNlvqTotHzeort3h8h2ULoG4n+sYYGl0yFoUZWbloe/h13C
8XsQ1QM9U0vQdLyxYFSSZCh+Y5Og8kfhb/H1htSN5UdfQ4UuAoQqvvXFdCXGrS0U
84yKMnbeGTqzukat5R21s+FFinvgDNuuyLHo0zgenL8UjRcPXoKY2wG0sNfyxTvY
ncrSQBU1kJcR3/sglNKm//0uZNppwM8eBZMk/ltvo+nX7pPCjPqjfHwJKCkbAfQj
CLu1WKE8RI6MkFXY5PGV9rTumN6hxXzA44iorkozaaqwIKjubp+XiWdt5abT78Nw
ZI5dfZubqfpXKUzhT2Iw10pn5+4rLBKc9zISD+eDdXWQGdxmp0K87i5ccbJUnfD4
5aexZpInL9NrZUeDmq4QRQNB9zDQhslf9ufJcTc4vu6XrwRYAmHmfB84eyCe3YTB
Q7nOZcbTUvYEndEl72KheySeyj6GzUTS8kjxVowmC60pL3zeeQcSBjTqfGyqgPvP
VyVbwEUhI5H2+jhpQwclwc+bQhGKu35DdsRYYGVm9CbykQ1Rv310lP/kWxkbCJPN
b2X/JdeD3Ph6frdUDAPJED8ta7zC3gZMU/Jpx81QeToYxkVnXCm3IKzf1k0oxXXO
p5Nmh92sJUSLDs9g3qGXk/3cWjyY0dbEIK5X7acHrApkU0vGPcsfChMaLhcOjpL9
wyGj/oeIyAsf8O0WRwxTpHLekxutKQ/2Fy5IaquXyFnXI1pYtPvOZTgTCguJi4VG
DMrg9ln5o9cmNTYAJtXMdA==
`protect END_PROTECTED
