`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7iujFKtFnRVGUHR1/8nNWUcwaI3pq37AfYCj01uP6stOS4SiDeMvcUB0F3DHOZL
/l0/dctdlaoaxHxqAAfxnnUS9x1/DiyGeQmdR68kUM2mwC4xXGOanWIGu3Yxd+BA
zBRQ8dfxcSWqCvIrjMnhyaSI6XejdlnfUky97UOzE3VW3AEcnahA+P74yi8IFsMR
g6+lEnnauxcVNrDDbDItVW5J2edyZmb3e5mMM5shg5Xi87nXXvU23bzpLT3ZnHB0
uWVgAYAD5gEYNmygaK6+8VxR8j5jzwFPewdadNtwqogUraKimDIMe0olfKNWMT/R
174Bm70PBVoYDae1XtUQgDNrcVz2OvWXM8l1fSy9dXQufqAQiwW9aDv7SW0fYMZ/
W48uYQzBZjvFlqNQsMdnLL9uXVwdTc8Bca9fAYDjt0FfCfeUyFaEqWCw2EHwu/zE
Kk5ls3UeBE/4ZKaRQwWHnw==
`protect END_PROTECTED
