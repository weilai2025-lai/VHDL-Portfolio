`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9rHS8pjeP5hgA4dwNMGalecEJQXp7UHdJ7VtpYvwKx3JliZHq1+BkI4JamNReyv
DjNk/SF5M9rzFQhwNK3OVAEhJVCLkzCMBVb1Ut53zQE+Z2/jIb3uQLVxtu3j6Blw
6ntcwYiYIyMdwT4nRFRmiroP1onoDIgTLiqm1o+9+4OTI2FGWE9N0ChQ6/vqlUwQ
z4Yyga9W6FBcruqvmkl1PRftjriNbjF4eW4RauVMCiSF7uKiFxCwGgmzPO5CReKm
5c6KpxHRpVjWLM7nlRbhpq4GOaK09ywKjYIb6KpOF7DFnfyrtSun6Gwx3q4v9a2+
N+Q6lBF4X2Knhvmtj/QIjVCV8IHXvDsdHSI14MyuJ5pq31qTEMSvOutGrTwgQgPf
nyDpNmMoZ0mQMhcR/AtOTby9nsUwfiog7o7D3NESf5vgkd66EyB1naHkDzq15GpD
gOCC6o7S8iQrqTIN3qkcTofhWUKgavwPMS9ffIrVRfu24FOwLujNnRKtbngG3gOs
XKRRSHUx67BEc6sq3/tt/7If/feP0gewSqoVLjxMPk7Qn/glEEjaBofn7cw6UAZX
CQVBjZq7J1tY/up6gtrBSYfrRpFHaNMN0ZM+kqHvN19zP28ekOOHGfnRhrYlQN/p
OWkCecaVva3jQ/oEQI63j+VCZ25sotUuUlhRZC8CNo0hg2Rbb5hxhp8fbVKr2MDh
na8GmJGPAJ8vDX1V2jgRrM9RhwIErQ8dlXBZ227JnJNzYDOm5XVbQLnA27Da27Fy
YkiT7zmvEY/Jdy4VCmqYrB5JZB6XDPMIR3EZVFeAt/qANwkZQN+rB2Rc5HI4b6oP
qFWU9Vqr2hWhRqd+EZZVStYwNZf98bm4virAYAHCtguyJLUP4330rHwcSoFpZDLy
jmigzkg3/2/xZfNegbBv8r5OJlJUCOpNu/fi01gtUBv8m534v05B8qH0mo2TtBqr
OELMlwPVGN89bUWtE3s7LmoUwMdHs8DANOW101uh1VcF0oP84MwZ6/JrUn48KIe/
rylUI494JJRVaYp0mFmGkyJFMaUuXx2TQ2guA5y6SzaTqvBsPdAo7TE72kV6kd2G
fLpt/KW+gn61TJSsmwzvxXY6GvrrJvKh2cWu0RxHu3t2of2N08tG4KnQ6KLnKqcB
J6D+n4MCyOU/jAOBuSOW9yc3YLBM8JvzzdR/+D+I8ZTVb11kHLkYGQUELJSTMHdR
L5YBk0KrpfxpgBIdWIrjIWcfJey/TEcyhmZjwRkD9gimurWWx1rmFbAkTD7oZzzJ
0fwQAr27330hja+0LziqTVpGQIp76iS85PwLmzsapPGX9+cVx4ZKKSuxo1TQitqS
dhdircQsFNgj8UM2+WpaCPKlUHhDGyqe+DQnZ7BSARMFiDPM9eO3LgbpGRaliFOH
fxZIfC63SNwA4UM6du2TeKX6jJBKoMw7Q1C1AKuNQvPl6mqpT3WTJq8AUJJeV5r+
7YxLbVnpyBXOX4112gxdvV2sr2YGZCMErdvAQ4ZiltYpLYvJrNrtqECySRW2G3uz
ZCq/3piYJmD3aFZyHvVZilbX9jD+62ugGFgS1XwA+SEAAGlyKJXZr/P8pwC7uvKv
XQaC5ylF383dwFYhhXBB6hiet5WvNP7h2K5SHqgnUmHArp3F9TWrVbB04nfcCzIt
+UAMFYEKbXjhv3lEEk9fcY6gMNEsK1p5JFQ0WaZA9M5DWslmtdqLEGtZNTAaFqFv
sweywJdB0X6wj1pL4P8w/xW+5NdqkWo5Fny5v7D0K8seo2A4FGdNu4ZbZWkF4HvE
HmbvLKLr6PU1SG18TFcZH+7GqkKNsr/TswA6JS+VBb/rEL968eNELWnd9Ovf6gD5
QJoX2W9+EmCiMUGxE49boCQCfxqQj6C+dv6iKc/yYrEuF13+ibrNGOm6hz7e/arU
aQb1B6R2LAnooKiRkTPe83vRUjHYLZ3e5+hCtn52e2LLHTCIBcyCPM4cUAxf2Srz
mOmcinXb3Q6fP1cpi8a7DB0H5zHGuU4g7zv2K07lfFP0iQQTFTPsKjqNr3pTH/eC
xVyJd8dsyT/KmsRAfOgwrvIlcjgCXjhHT+dWt4k5+ZcJpjW0jYZP7HR/5RiPFPY5
ibwReRQD5+8qFWNwdzc70SY2O63WpokK2axBKsuqAjRypT0RX1hNbne2n9L2V/DP
HPme+DSXN3yXzuxXAfivXxa/ocE6UNmp9pjadYLrNUJxmByHhEWDYf3q6kW8ETWC
MN+gYZ6TkX3s+tPILticuex5/+XKf4wJldjtnLWLAiBYeR7d61sjRE6fu+IpDopS
wVBzgUdFSXIDESNs8oXNK4wCsH+oE1UQIsAnZ+Rva2LYrqWip8pRW7pqH9VyesBI
+WOG5D4zugZ8q+pTr/Lo8o1h8JSTTT8u4vYkMMHvzyTnWpBl6Vmckv/3VdJHwPxn
xG9AiyxCysXjKghBffMn3Dqb6HZenacoOnGfj9FfhmiQZu8UjQ8k2aRIm8daVhEb
7uyZj2aC9reLotmc8hW1PAVUopVTdCChyvKYlnul5WYwjtnXCmoquFiS/kNi2sL5
Mb18sDnFXFkoAmxE5Xgb1jk93PNAHRInOipHlILkj0sXhAKRglBH+BOYRNXmBPVm
KWEJQDi6oMqM8IFA8vf1g+gODOcXaPJXRc1AsR5oCyiI5e3+rr/FXnsMvln3emQ9
gbg571aqpON+EbqRNs5BuozQbeC52vX1+qRsfyWWVGipP9ngjkHiIbD6Qwlk8uCp
MKdqKEpMplFg+OySsbArVI+BeaJC9eUVSggg68MxQQcoL4PsuhWfjkwoPhkbISWm
lsyarGI/QSL6UFPYwftVh/zLbxy1LXrjsDZJkuZRt2cdJA9zvvFGBI/kd6ziGgFq
QynEce+BFL+ajzvmkOR3m0uh5gCX8elLd3rlNUTxPiRg+en0O6WKrzoSWUh5Dayj
V3r2d41EmTqIen4HALqmfjiiTS5H+xdxib0k3xGmyT//LFHJTyX0ESjRc2N/3SYL
P7NThNwaat8Kv95aklrMPUUEp7S7ixPycmR8iJoZ4JK4awn4ME2wMugThS618hcb
JwHxTMDW+BHc8DYhPN/8NfAOK1tVxjI3zxPy9NL6jKI4HV9hDQ/nUVmyQYgv/noH
tRShyrNmaL3ZY5OMWAXeWoAcDTxFYqv2FQ0oaRCbhMR1R4xWLBWht2ypdF9rVNlF
yNoJDuaXJc7gDixjyW5AVT1ML1oNXg6U00OdEh+kL2Prvpjrp62mN6ON2gkQcfjh
7He2Wf1v47Fv4BSPOW4dOxrB6UQUBKAWQFyff/KmNRkS11jk3PHThdRYMHaCeyax
m6NSFJXmWHoaB8CCD/LNE8bftrcHzMiWrprLe/h0s+m8Nb9OueP7isW9yP40RE6P
dO0A+GtAmrpECFV9s/XME5SXuqGH2ZpAtQYfNwF4HdSI7Y+zPB8rbHoLkY7rNht1
/1aTd1q3pFontxHtPf/A03T8e1YyMJ+JYYHe3TOtJAM9z1OVKgWByzhHhUua+wEc
VtTbEdOl1sBe4EEYbdubEYYwQSzwKR65Jf0MchnCBmI0NfG5g789bbzNP0dWRG30
ARz2dcO6mX//j2J5SYkdVA9SzpcE+QcNbeFKX9vajb8ih9Xf7HT1f/Cfo5DOgiu5
0OPXaqD3dlkE248/1onNGYWoVYVB7bPgPL0/l9fq403BOO5HZIU0tkhWRrVe/dBs
IRQwjENC4vDb4xM65/vj7sP90ph95Oho48slaE1834VokxfNv2+wq8IroIafPH3r
ChjK+rok409F7jU8s9u8bkT5Eg5jdDWsypjE8yIee2wpVs2rW4uo5TIp37PPw5sA
+WA5ZV78Mj7zhrJG+1lQHtEYetjcOfn2XWB3bk0UzoyRbyOZfCBCiVSGFLI/TgCe
xJN3c2LPAzR2COt5FP9Bk3cE/yB/T6Tny5TdUcEhw2D1LZOykOK2oEu272iJtZ1h
Nvy9aBzCgPpjpXrTe9yYYwrnku/Eo0YN2gD1g8wy/sijr6bayk+62ApUIA3f6esc
0yruXE5SAxrROGdcKwHJgXtaNGEmR8DBi4VgBrQYBRq1PExfHkjNsJSJTZGKHVIG
rmSKTlU+cuwi+qg+jCam0pxj+yD+9BHzOinIoLscfjaQXuTz59eeMLEzasqod9f2
JvUCHjiBpEH4F/+ZiVQ05/Z9jnFrcOuIi/bLjmWuDICXmb+vyhBLzXtzqGGYAviQ
38siAezor2Dmd79CyDP0OBvy1vacOKWHrESv+CdwdmfaXUUW1vYnBDQLXQPBvzQb
MdYcIX13wOxq2AQBQnOQ2B53QlPNgqcSfBbQ18ScDGLZz2+63y5hI3e8KB4YDCXZ
DL7Tf2fUBoPZK+YmtCRP4dIj2+BUvaM6rkx+zB1vF/tLf6MkrStA/ILUaMix5byf
8q9kNnNPcW5U828EupXZifeOx4kRdj4YY1EiRLBFbx+ljE4pe2oQoesyM/Z/906c
tJPW0TMkPGQ/jAuwsDJi3x4/l+D0iGHzoS24HaxkVW1Lro/1Ov9BYHm60PL1ZOv8
Y2abNQeYphscqsDnMwEwAUDp58fnkG72Wqnt/DCNOtWHUV5KfXuGtHpOQpT9GVsU
nsU5cI9U+R7p1V2T2XvgvDJPW67lqSGnQ7W+VbePmb+7p7OQwnXxNwGmCBDYhqG2
dNTtG3OUDoNoRE1zPxnTQ8d1lSqL/YgHLgf/ADInUjHUX2R2JTJ3rwZqP1ZTS01R
e0uUVbiNIrQ5e/LJwQLRMCFtFEZ/HHFYECyARHdzeqrHF80qjyNTCT4ioN1GgvF5
KbjjWe9z1fvIQ6c7uZP8Mfci6kNvMWOI98Lji2pER1XyUIIcQjUOI6+ZEMet1jEj
AC6dEI9yLHSzdwB3qiNI3ZPJoiEI3ZPW1QuP3wSX2Fs2i1zL/T+wsMtQaO6rokZ2
JzILFdTY6zd4epbRwPAcEBleHgjyiBC/sVeobqbhFYMZvK40L89e5Okjw8P2baoU
YqdFXh/J0iE/ucogN0SPL5BqfdqfB1CGzqBnmtuF+/gSWzMGqPiXw3DU+5yho+0L
R4sqJ36IzJ+l7795ah6UHm3p3w4LR4ZGSCiq/GB6wisbivDXWP21b0c77Eao17zU
oAl0UtMjHqrnU0fClecSa1v4MRyTHpasfgxSlgF4jJO4aFq+JfxN+j/pxwuqE6ya
5EJTQ01+JKGdICwyKIqqkw0kzJfFGsqx4ezh8MTI7hKNUIzBBUe4jrh6gy3pf2wi
B2U18dDR3oTuFTayUSQDYdnOZxf6kFOlP232uVz8su3Be5ocFzACk0+j0sOxTJnC
lcA6BfGk4Ge9lwvRAP5CEQojfhWwKQmXSf0J6fDnxt1q/SNz8IklXtdc0TsNZgaR
52LgQVPx4FdkfmTLr4oR6RMTfdiHixEfMitGMe5Zm8vdhb8I/ndBAtAnsmdRNIs3
AVfnngIa+HWIuJ7DIvgmauJoOiNaoQ/mk0sm5wsohbXIk0v0qCOYOdDBAfHzKqcA
EQ1JxdlR1yYrt5R7DQhMrXOYHPvjx+wFPe/ICDxGxAyFflioSPRFpO46RoaR6fnH
GZTGZSq3cGWlo6R0fpdBa+Y+igKb1+333AeMA388t/PtW700HfTmb28FaauKZr5J
hzSWojsKRa2y4tI8JwH628OqQHHrA7RvHylS/AKJfaciMppoLKylmoXdTwGLNpEB
vPDBexWRJ2XoOoPcBUsvjaeG+OHMAr+p83RgVhE26iYJl/KXqzB3RQM41Pkk5PL1
OUzxgCB3IW8NBuvpY70wBb/zWUa2ALVtXToYVRf3esLvYvzPDvD71Ap8qm5JRE/8
fi1040tSpkkDSeWtpm2lxgw2e2Y/kzwo3D9zkyXpVimSX4GbGmU5Q/YuPhVhiQAt
NTQhQtaDnNkSkyHeZFLDGybEkDvnXtU2Pggf4he9DPbA7LWkUr0Ve1cABiygL1cc
7X5yvG6CT5cCTWa6xWRgWUzhZfHqLGXu6nl1AX8Wbe37CdFBI4v1G1ZsgsutUF30
lovmnDPqK3vZkOarMyTI3gxjnmvElWAlV+L8VLuELyMkR7JTFWgwGV4E4IWcbaH2
NCuJvsFsVh2TvVB31TaIzNBRVFRj/+KqpRoUo6Nevuj8YEewl7lQRrY7czbMa9JM
h05QVNMg0oFVyG29l/PD2n80XJ51lz1YuP5YBJEdSZgHNyAyCCKjR+eJnBlQEeTr
ToRb2jGtfJ7xZiJEipzENiW+Co4g+R+rFZt8jT8ZQYYqR/X/SoFGO6EesCgUYq7m
LEHp+ZE1vk2a+PZ0hbIpQCuRUlltUbUNUR8OuvLTOyQJEuGy8Miw9wgfdXddV8RN
dv3Glgi/l6gFMZRRQTf5xycKZjWnkrVx81NoiO09qKuaewTXOpiqhUkLSWKUvRbU
ytKf2K8WEHucyB6Xt4lYOQwDYS+FObrKuqWCTjthof5TaWXhNoMnMeKsCi2Befof
PK+2eTuMLpD6O05hvu4t02dOlzd86xeABQOG61L8YK4ZShtVHon6Za8fUU/QQnFn
+7cDNnARRjRevv4qfAPN1SHSL15aDqkXQWm877Vp6T01p4xOLOgw+3UKLsYmZCgR
GKjZwXDAzW43RALnAI+qnNuPmXzIRPmzMRFv0ukkhLI2XIFM/K3tdP9NgBPRpNiJ
VB0URTqQYRjtw03ehLPH4uOY1ZlRjTtqAPLHLGhRUg/PRj6CHvbFgLwLQG+6Djle
XYlpwuKC1TMx5nrYAaSSdp5FxbZdb/wUwE4SX4x3u+pz8FSk15aiEmJGR4J+xnRG
0imTck6jApuwn+wawb66HUx8W4ha2/3dVwn6up0k8Q/UrscZaPAxvYigKo+fWerX
XYU3blOUC+2sZPyox6WrNSPYkeFgPrlcB6WFOUCqM0kNXLuJJ62TwWLhlTWWfhwD
VI+49O23EZcCaIdbljDr7DEbcLIMA1uKdOq8pfGuZN3Qi4aOnrLRAoXD1nk4Lu6h
o9A/pRpXxxUi4qIzLCVHZJVX5fMFKRaBHs8vKwrdhkEp76/kfLadxz6CYxBQZt6B
shQFORDH01Zf68QstNAaSN4ePqYMvRbjwFe46TAMilA5Kcz3TgSftJfAXMzbP3uQ
dgu1uv9FwyFHCklIUoO9B7B9/YpS/BQGtLw0uUPWCQatsM3tcAuFWA8npDbKj/sp
fLO9ASrB+9PF1NNUpWQGhHzD3BNDlx7kbiKlLQWierChXNl0iBBAnkbLjJTg5H+0
/gJ+2AX213ixYQDuGRa6ssi6cHektkQa3B+MUtR7EP07sCl7HXZ5oz65FG9e2Env
hu31YTGImFjPFppNRd6TPbFfSxVnk4Z0XM8yorl2jTs6PcIOZWiXBVF9tX84CAaS
IOiDOfIep+ws1efF0Rs/RnDUQiNiOVK28plWPK2JjdZU1HoiVIehN4i1NbMEz5yh
+VqEZ1OMucZdB/iIwh13oKe5DVRQoccjUIdqFdxX2vXMbg+GC7mnI1m2Cj3U8Tr7
degIQImAxTZ1Zw4CyncU586Sz4j3P/4qc3eXnZ24YCRyY5xmO7kriYNk7GuWrn2/
O96zWI6rHdzD8uCgcKYvxLyWwlp8m670czgGHf+B8FgZaUWJn/XaO5DCCbiPoYvM
V+a2uOooGUEbBMqWAWsO30lU3qRScQ8rtSDOhx7IKlTdFAU+2iCNmikrdgo7S6lg
cBSfR6FG48aN7bh34PwJgoZDBsUdEyQxqjXqTpOtT27nTBCcmxvvqqLX23dJHmxq
9teNJ7dKye2CBwWKDCsGuGpm2xrGItGQR1amL6NOwZYSVvzMK3j5Z1TnvzFMcZDy
ym2OISxFHx5hpHOvAAOmIH3d8aGPHt3PMcLXTF9SBJkqbAvTLafwIwBmRwxEvUcl
lyjOQ1PbCOHyCoAmI3dsKZWnbehJksPKknV2v+grT0p5Y9tL68tVuz27IjeFxLh/
SXyvj6h4zAbAhpxmKfbrfulKoKccIZMniQ5GGcITQelE6xVHUYSVXTeoyVSUKG/r
ZIFYw5nmEf7+3+8ljtpSKTrycruvbhUy9BsojJBmGlFSWzJlEYrilCi73da6MOLz
qRzNmXIoh6+NoBwVS6/PVtpjOowXlKhALDyXd3mvfE6Dwxh+j4Ag4X1PachRdM8T
7cP4PbvLbM/IrNcKn0P0SqpQ2WDqfOhufYZy3qGEZFyM/75tQUtWu03eYea1YxgS
2YWuTQiyHzc3NlU2MskGMQLjAVqspk9SCdWQQZZ6VEJpLKnIOsys8Jxuy+T22x1h
naAEwFHNlfu02KPlSINNPYM3RIqscKY9J0d4FPN869iBnYezqKJAB4cA4/8twsDQ
IkNdHCsjJ+J56lnuqpuUOXBaC5u+ZCUW8eoge68uIWMOXYp8gvYSBZHU81ToX7Y5
hmQq1FpNzUSqQv7PmYJYjaSRIFHVA9PqSsSOryjXYw1UnKDR/+m2IACVG7L7r3/5
X2QDD/m5URqz8z9/poY+X4wHnR+OIDGiNEuT4U7lLdIdMdKxZaJ66PMGD4CLkU4D
Ee167EBn4Y4y0O2NUlAMJxXLwgl5Zn0maNXTt67L4p6QjoAs1CXEhrFeFoMYC1e2
7x3w4r9YBbn46tN1xrLGbKWapFTmPuQ9PGC2euS6D5X8oNN4CQpYn2Y+X8UPhhA2
akkIUKkZkcClOrcOJs9505DzSP/HO1d0+2RLMKNjk5Wjr31DtlJ/eTKDyJRTpoSw
4+GwVupzLilghrxnfJ9ea+fYaMKIoriz0EqGi4QRIWR2v/QLlfUygZ7x/AGnxbgO
B4//VjPhxyAMsSUAuvchd9fdRhXq/x7Ep5wVfy7QYLFIi43HVhgLGnR+rKjzZ51i
UkE7bg+HDk88QFpltXk81QPQiKgFDt18RMCKCM9VihR+xMFXHtuxbWhHkPcjojQV
GE/plDqUSU8J7nyG4rqMHmUSqIZc9EF3A89GAgHkFi4C5P1RWiKEGXoxEQcz2+k+
sy07P5zkW3imu9mvJSc3BtnmK2MFT6dUhM66jf29jaVfts0ZIM+wkzstJNmSmAqc
qPBExSdsoF1KJHu9tUyOLIPaKmLFCbROX2zLtt1NW1cwLAHu/wd9yU7hYxsN4ex2
npG0GE+wa1NQbWBbTyoRR2lvjlW0d5MCtCN+KmdK7yxVIPqOqVUb5STR4rzJp0I9
NVkqkQtOnQ8CjdXFdCS5M+n+hDy7eHzoavVS+MwvGonAXlBMvRioVhuOXGFSRtCK
0MjNFHCirzCpxcOjsnrrvwyWj6kFvpr2Z2UL2bwn8n2J3DDZy9lvwHVHi9W/EWGt
HEfJKM9ugZIlLXoJ1Zcn8x2QW3emBp2fI0wfggyub2CHlCw6ml5qlilDrfOsfnon
f/TbSwDOoE8glR0Sv8h7PrxXay+P666y0caAmiG87BxPIDGS6AKrvMNNGG+6dfh9
cYD957E6A4mQ8EZ/PQoImBvwmcgL64KgPWutbRBL21iCWDDdfnpCj+XQqQFHngwg
y88AGTR5mMGm1+KRmHhLyk1Hrsq/PGO9J7XX2sLKaMyXRLQqz1v45UJ5uGUfMsfk
PggPodFBBersto+3Yu+G58b8wD4LJO5TysJyLG7LH/ZX+JvnRR5LzAY86xZV2kQP
bjZwGaOcTkR+vpkHHm7hrzXd/s8wrKT4/wX/9K8SR/OVup13nFc+7DUhwWejsiNm
5JHTnJjD0J1KPWRTdkGBA2wrvfXLvY+abuhzOFNObqSP6FZGHWeEyFA07JqdvrCp
GnSv71RAXqBAZmlSxSbG/v7oF3teAXLIPpO0b9HpWGRefJCEQZyoF0njGKSgv8DC
X9SEb82l6rUzEQwR3Wlx3D4MRVrKmQJgImz+x2PAGx7a/71AJwofdlqE6F/SYyKb
+Mu/bmpoZhKeL40Qm3jB1xxncUicwHgxCTojwWTz8unlO5Cgp6Yrzx482ZOseYtK
FdtrdKtqRTtJy60PJDDYWjm1Bu0UfKlFpCnvMa5h3qluGnXHfQiXESX79Tv6RAtJ
PIi1bZxprhpe5sXJtTdFw4PES3aoHi91Ws6YiAE0GZM2cAbBEdg3BdcTC1h2RjtZ
gTrss42wiRptL3hByvvtoV4O9J1C4HL7MeWr0qzZXSmHjnmM6NCgJG1gIpcD5Rwq
2GLQK+OLKl1LaRctFsBVr59ntL9+0x4wrDrauR03gOFLGRyfrwjLPdmA3f0Tgaik
LuFwL3BcCD2GAY7jrHSPcS65GkeMZOzeSlTR8t2TAqTe35RedpQUjRYF4oY4D6p6
nZFiAYZP1BFKbp53WfcReU8JyXPYWcsfepRdplp0/6PMKyHyCuRWKR0GMTupKqKV
QWTO2bIu4gytAmNXbex5Wl1V5BKv6VDSOF8QraazrgLDSG3zU2edAHAjs9go7nhO
615CB54t02bKxLFTy5uJDIpaMx3ZVJhPqWRjDR/RsZL2x8AZbQ3W05dQa/U1W5SO
gGXU8a8yVHuBhnK7YryfgOnZi7x0K8midemOAViFnqsEAj6RexJbN+MrYZBYD+6t
DzoV3KJ1UmnjHR6jxgJDGL+LFOaBbsUxzEnLCaXCg5a1ge3IC41Hwrv57hSYiyQG
/KF6zvLXojJlJ1rbbqQqQEJBOtUrsbnGO3mMUCI+s5D+aLX074OdFwPaQN0ifK2D
7AiWXSJPQL47bG4jYrqeV1oRYTq/eKDd860HFl0xHyClP6e+LiHKHqxpiCPIllNo
jFLIU/cuB1N9CjSWKYXk5SgzbBat8Rnf0q3m5HEKW+IPIBaZ+dhVmhyjjd30mynH
l63KpF0uYVb3b5Zu/+DF1QXe5VU7BGyQ3N3a/3VguojvUowt0antXmOBr+edxT3G
Frkhzv5EZkv+e/CBn3MbFvM3ii7/u/7/ffuDreGc4ZZOpXu+f2RMv31Mc5emy35t
KkMpSMguw0al7Qx4bcJ5jwuK5Vk/MVbMucMukG3YdhhjxjyEn6YH11BmvAXEYwTi
1f04Gk53d4K3uvvzwVXi/I9KK3Oolc83wrus+gEdo5s4p7pDLrUYdLY80ZLt8kPH
w1AOXP/xr3xgk5c+syBmkKcJ21YORAtH5/1wYzPhwbsxQEu8KDMKOtv/1ZEbNbtS
MtdNnqfj1A0bGrL9aJ7rflpFf/M9U7mMvAbLZMP2AIJ1kcGZlZeeqbt3s026JX1/
ElAJyeGUzT6BllOVyQJfHiek01lGPUxkkFDpn36gYLS1Z1hsz1GGpFJsC0MxUwyv
FBnK52/M04AVr4aq58EOfYJGXwYUCkgWcH9uQaFy0s7nrllYVF1uJTX0F0fJsNBM
c+aDx0tSZ7KAC3OZgKkcPe8ukcTREUOc0K1HiuRM3tt8y9hpXKEzIiXv8wPy/72O
mD/8JIqTstlGgUvq8w8fJnb4hmxFsEFAV1xq/KB6cZdzHmqjGhhe7cwKrnjeoqSp
7F9Oaf1MnwbpSOoqDne0+wj8jo5Luri7p9KX2E0sDyPMoKKQu7sEPnmwcD1e50Pt
FAsn2Dw3hk8NYfPc2Gont63VY5v7rrB+8OLittNApihbrH8tenmNPfd9YmA9YJ0l
XQdcTCm8fvxTqjccJXuKOzlLszAEkx/BXlacZ4RDlj94OJ8FYVKQUfBsMW0x89KF
fiT6ulJA/eeiopOUpiTFmcr2l8jdR4lwk0OmHYkLOEG0omMw+q27qabNrYmss4rw
+oCxDkZUe7Mq/B9GGNkohn1UL+tEtYotwdzQf9i0ZotR6nU1UurKxP4e1kR48Pra
bifGu4X9Z5j1ygWJfvMki+FGrx3dMO2BIZ5mwx/3R1COlMZ79DNyE4vGMWZlmdRA
MEXK29WRRYXziQye2bmXYdyDh+u+YaXUjdRMdhrG2sykIvhXUoBhPkhGF7paqDD4
oBCAS6Oyyb45M02n38eY/XqMun/0kpfj02ZbcdJA1ATtrgHnyHehL8WYE+QXE2im
Nv+iy5kdfD/DS5k4wEANBgyRpJ8GDvC2nqoMVkzS8KbOJHvnbbReWFkWt7FoFtiU
VKJaLKvD2iIPJCIqQwpN2sc2TKQcuO4H2gUMMHOy36d+1tGo2+hSH+hVQWrShs1y
kfi2yBmQeyT2D+o0J/g1TpoXyG2PVmaBpkXKAAwyBPyLLbPMU8yQ7SVu/iOK9mCd
t8f3J+0wiV/cAuQsW+988RY5akzkRkgTxKxLv202P5gIRhIeoBGe+4nzG8vbWpeP
jUEApncKLFQxphppfl8XqcDonJxO2jU9BQssAIHV+BpibEhDIBdYnlnvgyFjG1SZ
9Tumx5b2K9Bxn4Ma32tvXsckEeRF9Nu96ULhStHVPoOqcBijeCApKWJ2mUn4p1iU
GZXBK3bUiECK2Mee1GcZVwZMEaZt3zKtJwazmMrpKXGfdnJNUnw7xNP3pNLiwJKs
bfjEWlRQMOBVsnZ8RizTgDzISoQ+tN8zx0vMkBKueZEJCUTLwYKQUUBvMxJoGDGL
0sooU2dOaZSBVgYMGU985tRtiLU+ZKE2KT44n1rE+e5Ps+8r0g07SuR9+B4D1Bwv
NGVCQ4LHpfyYxZNqMuuX8agAMOpy9OUeqH5WOpKYQqnr1W6552X1vkPKlnafB6bg
V69HZ5ThMhzgzPQIZbc7e1erDqMbRpMxHpiCbl7f9f8EsPfPpMZ7XkoXICjK6ffL
O02LuorbZjBsKGutVgEBeR+vxIf36C6y0WFP/8YN4i3Wm3vr918+jVZ+XBBNP6wi
BhugvD33JCUtzNLq3QC/enPEbJGOBx7V5dANmMKtECTMXu0JyodEpaDXtDxrKbNv
MW8p5aFjyQ5yBqY2VNGi1JIEB5jdPNS9k1oT6mGQCOJrHo0dsd0um3YFP0reP4br
CjFSBBgBOUexZRMzl9Kgc6Gw5v+y7TOAy32Na5W1k165KR/xqVDsCjEgbSg3dZQG
fHJsjLQTeQjqFfq3U1Z37JA70fqBmj6deJ/FCg1OWfG2D+DoXFyV+r3r9G/7NewF
+yVsJUkarD3T9QvFJkLN13Nn1ewcPelqvazjgX6SMZBxzvCQ4j05f1LNMnLaw5Qp
Cce/81XRHZO4Pl5vX4maZBsa4Lgo1XXmftsBWSlFiHyw6Oo4mdjmro0ymX2bF++j
SFVtcHMj4wKLsSlUBAXJjaaasQF6zyBQz+D7cM1Zq6+JcGJw4oniwvSf+qFnswVR
CIt3dGVO+Xny3ffrQNZd3IsN4gP0s96RAN6fkuSVI/JiFah6Sn0nTqTxRP8fIlg5
v1IbxlC7G16YHj5slmdziWg+GD6Fd0ro3SPR+0bPhT6Ck59ym0SX3FqPNZHiVKyD
`protect END_PROTECTED
