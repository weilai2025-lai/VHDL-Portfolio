`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IuwmJUZ4D17YQiKEWHhrJvlOtkCrU7I1IEGA4lcIIalYOSkD4A3bHsYDjk9DcLK2
7xHSVE/RDGPYEqiXlxrNjyJtZ5H4kUX5bv8NOha9lXoMl6yTLMVNiSS8onN4WNBd
Fr1gFSyEHlbzpWYxs4fgMdMk4tPap2ydQAaFNPFWbr3NXN9YVzHMx09dU9+NXoU2
27XBoG+KGeP2P0hok7TBaGgU9LLZP5CUWyfNj7E7dqugswxFQS/uENSXObxCR8Ob
uJHrEmMAQrMVIAN1+4E41/S9w8MBbMnemYvPDicWHoSe/NAbLDbozAb/FEI9NAeC
N+gWDYYQIdSU77eacpqfeBUAthwyJYSRbYl06fRMA6URh/K6lcyIybDYOQof8+0K
M+sm31Oh2kLo1qTLFfzrUza27oliojIjbNhh1kLyZS9rXTtjYQUtXMUUDlV/8TFm
mrloGJ9/zYf0aoe2X62rCsK2UAU2kNPsf1yAplMq1v6ink5zijPwYZl7HTSNjgsX
FJ+jHTB9skjGJYpwbRSa6JkvymhS3PvsQ+xczWjaN+ZCR8KUO5xFuV2ikiCek9c6
VHFyaawsUPTpeG/hB5TKSZJ0yjWhKFS6PEcdWwukWl0MkGCqxmBXJoYdk+17eh5g
L++79A6L4i4irBKRwqniBaFTnRRbPRDnEEKMkyRhp855gj6f+L0DpcIg5DpIbR8x
fs0adasUQGOikNy/eZ9jQpm0pYUFjaKmIoG0ljARmQ3EQOad1cyvMaYm+tC7GmBj
lEKIe4nP+vBhld9vq/Z3vcVyiKVNO7VusDXRVgUlUE9cPuv2zEYmY/wS6XVbrM2H
aojv5cozO1uzY711WGYc7W122uENnvN4JdlZHx9kBsclYavz40r3ZgZXV76SFKw+
BmHz9rcdzUcWerynHh7695hKjko4TdyqxKNVTVryYW7PDtt/0Ocsuye3zF38oQdt
n0afxqbxHE7Iy3HME+xpGSnFdiI5Ks/YaOWMggLeyk6kQj09CQNlWpBBwY3ruSon
NKGhe4+Kyiu0rL/Ddb9oQ0GmST03ymTw21HQvKtQwEzJpD1p+sVKZCh18TG7FxxO
hd4kpT3M9i4myUTyEGbMLw==
`protect END_PROTECTED
