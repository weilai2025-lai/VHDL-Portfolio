`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NuKDkAZFJ9uqIRR9Qw4d+g43FGZ2+OO/CnCoT7tZPJbavTHEYOFKL0HwBeB7h6Cj
ZeYU8RcT5QyMsUoh1Z8VT7act/ym5AdShRjFxDqp9oBorJCww0ZHT09kVPD/dWQf
1r/wUfE/T7/Ar0Gu8qwrpN/py2NgJnQOcRj5rl5yZZYXUg0du5jKuE3dfJuDKWXp
RWnsBvLKCBxJWgN91sbmkHXlU9RhX6qpdv+lfZRzi+DQgthQleRCITtPSSMWLnFf
4/DypF9MuMhTLIL9LvbIs9XBZgYUAJXr9uWK9jx8yBR/5Vu4iyhkRe8i2pMk5Opx
vz8ip5l9uoJ9LaXRQzC1K9jLa8iSMvomveRdhJ1aATtf+F3T3z5s7dewzmmFq+2J
`protect END_PROTECTED
