`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gqcsAFhMpRpaDKSHXGNK3tj/J5QfyZV6uBRNbjwrPCXv2szo6DeevVKM7JlE8H3
LK+Qz7q2vHeGoa6Uf4Un91SwD4cNg0sNaFvemrUL8N9jZIq1tikpdvlbD1UxYlkd
hL1R2L9vg6iVIl/qawwSaGy2gCOHWkY0XK6OZOfzS8wfhDPOA7HnMrkl/AwSjY7D
T7RWfxYMnxZrdcuU2JZ+IilM321lTp3SQNawMvoTxK6AHPfMCQDcrYuej4eYthU9
JGjEYSVivDzjVc80hid4UiYh60M3Ejgdq5f0R74lqQk/4CUy8ji8gRGhKcG6+Rvc
WUo1PLwEEDi/7GbqOrm8bxpGywX07eqS7zLV5PloT12O/SHxkvC8dnraue4+fxq7
/Kxw34A9PatDvpO/Aq0CKktwkGR46fRfRmNeGhM8JS4Beoawp4AcWTFHTBil/nos
3i/8mtYODBumx5h7ITbyLRKBz1F6LNUJmmf1yBWKTzvnX1iFPeG4gJnSeA1hxso0
0ZJQ9WwFH+40Ivcaif/qsJHDX1cwISE2e1LLPHdmsoshJG8BHGPD5gVfQp+mxSHW
3lL9mD7qNp5N5CuiSoyY+jhHW3ms2kyXjVT+mkl7a3ZzEas8VMJAYzgIhbrwXeAG
JvShZISfaU7A9ga2fuiZGfUuvQTGSDBTlh9drkOYqo7Ht5NawCr7Ec9U0F/BtLu4
i79Qmjys/JmUH+onkQf5eY5wEJkkQ8hq+dBCQrlwsOrwrU0phgDQ5h4mS6de4Bnh
Jt68h02QIZrwqlKnrJsJWtPItBFtunCKcV5Eog0L2Z+NzhmN9r0NUMKSWAE2nJdV
+Dxe/2hepht9RQL0VJrR8GfvSSQJg4T1aSmQ2jRIn7SaZ+g/gyhlcKRmi86xMaOw
F4ftf1AY9UcrZONcDG7BVkq3DpB/I2DY7ky0QbPM/cNgcTIJ1ESIMa3XMn72Em/z
n8K84fjsZtfQs5o8uSKQuWrbY5cVN8BXkoMLHUZ58wbeq+CxmdAW5NKUodao+uAd
sxZw+1Yby1q6lWZIiCUCbZ5FhxylGtnTK/rrr3cR3J84zZa5tgvE8smMX0G665/S
Tbiy6swKf8fk8tIXAHORe+G43I6VdE9mY+26cimAMRd1Gre0xG+3f2Ibtmt2epKK
7TU1lBfbfwBKPNXiY+Wvaqpo+rtdSnHRQx3vdn4lLSIhncwp+4evDEQ9yrLxvqIP
PAnN0Fk4F8chOA/wGrv+WegdbT2jjiVhK/j9EySVfh/rg2Y/zUUVhz1UHOaS3/rF
pIhI6oyPppqHVPzcCKPlHN+gecLf0Oq/vge9bEJaKq3q8emgeyVuEkib+4cP509u
srdLa5HBXgAfkPyW1dVac8vQbp0kW2LGsn2n0KpVG9zGRGzY1s89/RDVxrp096GG
w/crq40RRQZvk9wn7JNrgI06v8EuEphH6nEtFJ4r6WvVOSZ7hmTbO8WWaZVHqmJR
B/8powmZYeYwNwhrUFWCEdfrJw6LVDHbaQBt+ljK/lkgRiDoeepz2nZIy2DdHwA/
zPSs7m9WmRGll2Yy84LIGAFIz1A+2qDVZifAjl9rhDLxgHX+OqChXrOduWCzNBQS
UB4V9Yvp+/UdOtbDTDPFKcv0GcSECd7hUPrWr4rJs6rgbMxEjoIR0FLTiNeUlb7D
UF+4IIxhOEAXscusTAVFuL2biIlnD9lOz6cykWjkCqJnqP0sDS84NNT2QOz3bh+F
z6Gcz5qq3O1GSD+Ldm7mUUkShl6qJeAHF7fxPce24E2nZcyv3ojAUkiysuu+ccRg
Aaw/0Ff9+WyFhUJFXElqJEoL4UzPltUrcnmngmxq2cR9r3N6/E6XBok8YyQ/NnMl
+4Fdhgr6C4S2ITGr6xcRr24cYQqMPtNXpyChE7Ql+N75bxpH/9fCRA1DDgiYO79H
Hg8fAuMMar83A4XEg7p/y4BnX6U/Y/JagmdMNmXuLujj3VhEx4u8M3RMowzR2E5P
gHn39RxJoWZqwnE/yNaKrWFtVXTT5S+ax1xOBsVdqCphIAt1CgzYat8Fp5uSpYpA
N4X9wcWD5dfH0vwBT3W5NenJ+sszwohbjFMC2BN1GjG+uGaqSOLXdpFHGyMsykjc
QUs6TxjIEjDPJiCNRaphNhCAMVmbP8/jYviCUgqednclueSSrTHZnirvuB/ca2t0
/u99s2yDTZvIzSjGV1H0Lg4BlUfVA6kgxXOfNwwxQ+2B4ukH3/VyZILSY/ShIf//
tzRxO4VxWzxufrtymO/d57zS23RV+ytYm8c2bCLqUI8fiubVOVEuTbRlDlsH4ql0
9p0paiUbbqlHu2VtxYLZLKXuuqATuhZ3l2o5UW4BHzxHdQ23edBG9Oa7/FOUHCDw
UvSU1CcCqtfq7FvIpUYJkY49EmMwVKYoVrbEV3jaU38OkROVKQgJDpK8LcCN9GbB
1fgQS3bujIaJnmQlaGnoUgzAGULdOdcJZh8ItyDIQROsMyuDMyNB9s2QoBC232Gi
Ie26uZYG+JF50z2lPENFYA/ftSNkvKa5N0L8VO+3+kI2EXQZHInuCxZW03Hxc4b+
ZJwCS+qkCVR2AV8wOEt4rBf0E685iU1bWUOot3QFzMowBz9tU5JHLw2L0V4WMDv7
VV+7KuGrlhBZQVhv0/L/VVkt8KXcjwEJXlY2/LSLpcyXGym0PJjnY3qv3KX4uBAt
je8ijQzy+ML0g3uxy6r4Jnl8wDz7CseDFESMRAWoLr0xGWymuPG5Jlu+rI4w+98U
YSIaSjx2+1NpFFEQ3pyaxF+h9BFKJgsLsvMcO4DpZL1ls5SImTm1/hx2SnMM8nhJ
kcm3HQ11wIeMqfChoJsh1+kH27iSBW8D6ZVTEn7CWulIqP3mdLZDkZ0av0qMW+Y1
LsuCp832qQboKoUBl+3jG6DOmdldH1ueu1O+0AoGezs=
`protect END_PROTECTED
