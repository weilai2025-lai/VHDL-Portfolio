`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKR+lDwRxLqyCZ26/dHNgzf7AnPbygbSKj/67aoct4LKhr3iJRx+bTVh//BHjwIg
5yRtuKxS8jC87MbTqJHKay2yrBIOPK7le2MOC7gzZsOUWN/UWpJwydiiLHcFReR2
egREjYYmy22b9vOyRCaxNuiNGouMYi050wvFe94btynKhqR5GrKxRGo8SBngIjl0
x6qmeM5R1IO3EL6UBjhoUujlEk6oaFYB+hmG0EHK55p6dxsLtvQyAuEzfZFOjaK6
Q/ZWGw8mkTYh/OpA9kV61Wu/L4pMUImuZ7cBEZ/Gv6MhRjV1BS6WFTW7RU9rhr0e
0ddUP2N9PijwIHB0JMaOqAuKLBGN5mMwxWd7JXpccRjda6EwijtGKIUUpWzyLU43
VdszwLT9cnT6nMuRBg6peso8Jojp7w/MrJeeT6MAvJ2Fu4xrNd4vql6sdZOalyoZ
8t76BDg656Qn8zw00JBwcWNiUaCc+4Q4dmm82DHaBJnCoJkf9qdOrMG5gBGLOdNw
BE04r6VC3Ussn1upizbqRhTtNCC28yTmTeziWq5cd79Jzk1szkkXDOWfMaIxeA7j
V6IT+UTb/GL7JLIITBmsOpBJJvna/F2n49fc+eZypZf7FgEoTpwJZK5OAqVIV6XJ
PAxkEPBzwL2M5DzkOXhl6ajDigqRkKupaHHjIs5HGMK052cL9e3XqayiaOHsQi5s
hTeCj9UTSJLdYltKZBNYb0nQUUp3MjuE5CgF3wVYZCvaDho2MZHc12cBXDNICNqd
`protect END_PROTECTED
