`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWPVO03SAHPoL5A1eKtuR5SqS+r5FX1ViW28mZ1wUVUtE6ECMBE/OdHJ1rocp8TD
WNHU+E7Em14xuKfBT1bpiHa6jHiAg4kvEP/ZjCV6pBhY/SnvB3rTFMTnnnMbpsbv
EG8r3LW3OkBP6ELyaJmIOdZ41/TAxwCp/oPtxPcXMpLlxCHicoZ0+/fkWSQxIlVW
T4CCI8DIDFg+aNVLpiGOQynAglyxHb9qXSwcQjWXNDI9ml8ZmstxdOI6pDySoI57
5wEo+deqxgacnePchKWZQ6ddEZHXx2gSNBPJpqNWPM1SCqyvBbKun0r/NYr+2OAD
wruuqEIlVM1VfvzErd6mt9wxYVskZizyqz76H+vJtcHePfgoMW6hOpTrF80NtCo1
bf3Uzcke0Sviw1ms2mPtPT0zgD64VNEELSR1kohqpkg5qGbdj7gqv/VQskkB5JeP
UFXz+astjmcjkVJzu2Ki1O8OO9MInEpeIPd3tUEopoVkxmVGE2uDx0eeF094ggGh
Jfd1tAvqz5l73BjErKynB3KlAknKgJKv3zcKvKTIsSh+ceTVWzk/+UIxKEqYgimV
NewUSxFVqBzLNETR+Gke7JBWIXnvo7X9NtL1gJVWZej5NEc90hw45WYC2MP3Wqdh
DDaCA8HBWfj6wR2z6GZ8Ixt93ZOIL1hcVAguxGrGs2QAhus/G4xCTjoYkAKTggDK
VH+B1lbIRemtRejpbJ7vPFTZhBzkoTObyU0cTh6l4V/thdcdG03dT88f5pYnwlzm
0tcaOUfwdXJcVRhRiEtxzFqTEn5AJB5PtKl0bIIwwzHz66q6znm+ropASAAbvn9J
eRQuNVp6QkHU9hKTZnCtX/xsLJI3eQChTVyrIMEHLV1bnL1AYTM0nFHLVeS3QR9b
BG5rZzf9GfTO/Qrl4VBSh3IxxKvajrwBsURLhnDgO4yQi/yTnEhm4bm2B8ZlYO9g
rSAl9n8mQJfyTeJv+qUuIUyh9t8iANx9lMOdcBl5XNlP6mQSKIPFagPdlsVek/9v
W5+DYV3yr0dtkSf1U0hHCQPIHUecgTm4Ct5F1zIyZTY=
`protect END_PROTECTED
