`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tif8NA4rcl3CfUgBqzVCAqwkP4gI0AkXaXOJgehEYpmVPDRBr68GcDQW/yFgIdqb
jOUhWB3uWJTrWakbMEFLO1TqznmZjV/zluNpfhmEKlIZETioLKDV6aMBP3uBeDrM
WF10sBrh1eeeuITrGw25dHYb1jH1+K6e8TtNJI7Nh3GlQLgbVZOS/xfLzo9IPi6J
KqDu10u/JWjQnqRkTuAAUTmxj+HvE5bmeP4SqtXTz1o0Ix9a4PdgF+Fdw/4I1p7i
rgYoNDJGeNW7R6E5UKWtzDiT0KB4fndn5N+g2NiPiWzIyS0PgecEz+ghQSU9Q/AD
YVBUjK3wmOfMjUMOO3i1kTXeyLKMukFDbBotGPqUb0ukqxzRZqpG1Tl+U81aqVbd
2VGY0b/WjwcgvTHHIw4P8e2dVGDq87OZ2X2SskiqkzYiGW00L0oIFiy/8f73bVyz
h+KBWJDaVulcsxVX2DXMzlUYtjnuCbPFlQ7LyW0bt4tRpWfjjSYRXTHKR785iMzd
mcblVztoD17wAWFgc8qVHjLYiA1TBQUo6SKh26mFXiTXUi/DW7BqqqvpgREmLBCn
accw3eP1kI4HyU50UTMaXxws80iVTI37ABhds36HJa3Ssyp8OYIYFAwxGVJSNJ8X
shhtONkq+BL/Mcw9Lq1Gzw==
`protect END_PROTECTED
