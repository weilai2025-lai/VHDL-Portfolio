`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTJm9yleiUU7c2nrr63R084iT9YUpwxXJA/kO1PeEbpkKgsGdYBhsosv3cuQ7I2h
AvsZV+REG1Vh7Cvp2hRNkULRlHNEbNBll1OA/azIaqgbNDck4ysqOIOJ/R9us8wO
E49OJil7xdIuQ/gmW/V3BcptxlhjFL+/Q/CcyHN+y8rq7wY37Jo5/7H/2coB7dU8
Tyy8mAjCaOZPKE9C8G+JiWwX95VIV7RIZnRpIvtakcjposW2mc1ocQdNrShulL9+
POEX1AleCLbDpupHAq3IOiwmiK/agDk2bO0GFrM7PFPKn+xiwvAF+cUDyhdeXoBY
4h4RqY7jdUDA3pVPi4z6kQLIDNQ5Xy8311He2ucufD6miR0kIcZE/L9pYqbUStlg
VHNl4/mIIix2pUOnRUU8bZrN2VZowb9GV4JF8tR4sbCA2ON0JOK1L8El4X2QQidL
0ftI82ISUESExjO1KYpcAYfivMZEDlyqPNWqjZuV8R8O3MvLfgtOxpLMdXOERvCu
XEA24B6qy5bHjgWC8moXJXSHKrHlMMNR1D8a3r+TDCB+07fknOmnDp5wNhcprUXC
S8lKtlQS4vHz4ZaV4mF3eD4pksHelP3edqrXq+qQL+xS357VE+Z90QTi8QMEnB0p
`protect END_PROTECTED
