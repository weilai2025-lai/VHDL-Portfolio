`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBGfPkq9nKXUQO8AHQbmhTjFWWBEK4VwLGSiEJjO4FokyV+/Zy0xd9ZVAEAZyGFT
J0eQZydVraEYbxgVKJrP0x27OKOD7gTVWEPoJvvGUuzbuRv9AQEpmJd4UKuEXN7O
y2hqX3ojh1R+FnTpgk5ZLkLEWk0OV4jQ+oGUvawoD684kyUAeWIxBsJtPFD1o5mj
3kh27ZL/3y7GHnm116KpYexiRth9PwLcEACyrFEmC7Sv8s5HLhS7FqGAKUEQKucS
U88Nk52C0Ij5syX26Dw5v18S0/ylDnRkSez+rQ1/2UIMD5QlYviaTOz86Nl3ybYZ
kUzxHMMwP8K1hRnNvWnI5bVkyKyjVTwOoXK760UpkNRR/fkLffQ8KnfI30ENqExZ
tiMZ6KQTRWjEvBheteLcnoUm1SlYlkj1SvFHoqXA/Xv9atz8DiwxBKW01CvAUFyA
Xchj2qxjvw0sHfNE7tZBcZj85Nj3afG9oFixE9ewiJa6Hap7n9A+KPiHYdwZxNJf
GW+j+uQBUDngP22PmHvMN18vPFRxW7CLSG2iwsS+tU70wf/Yx6plxq268j9TI6Yi
KgJD1ofE/vInyBbWGwMuzM4HGWqu/zm1ztyae4GEJT5cpp8NKEixJJmuPEOBiU9t
xZ0a9n6TeM334Zdv7QL1odbSc0uqckR3FLd2jHaYuZxIK6fifAEg0CLw0DDA5fAw
l/Yh4OD2a+KJJx0mi+eif44eOBDrzPKxV9qoqrDprfWnttZ+esSJcaOzrZEoX1oJ
F/5JuAUyMcBxF3LJxDIFjZ6UuCJ6kFoZO3pIJMHNrRVpAlL3dXa+tSnqFz+VsHnm
+xZ9l1ZT6f1MhSOFOhc3XChRQkLLv/m6fPAcypTDdxjSvBi4Mj/+JadGC3Czn+Sz
jcf1PSORiy6KyqiyVwsfBMkzyovyOPLwTEDGV0txw61OvwM3MxYPUN10fWTFnLye
ve9m5kse2sruhXvGIqN5N9O/uz0uPDoz9+jvOIOxstuxEu8mfeuQJGCPrxFUai+a
QwCb8TEC0cKfxXu6PP+MSnoScGrdTbClD5ldqdMO92pdZnrueJOQ8OuO/yvw/eFS
azqIocMMtrAvGtwue7vvlEtaDYGO/H0NfH1jvIcu5oKWaLGsx4XFVXQQLBXuIwu2
0TxulLwOUEeozCoOdpzR4H7NQzZDEHOSLYDHLhY73EcsefrpY1W9zsUawXot7h1z
2Mw5epFvPLvkKYDY71IL5ZWDnYVNbZpo5k4JRhj2PtlJ2NN/45wqLflsI1LZRmiL
Vf74S3AXsOnziCuoINFWvPuCTE5qxnqxhQME/vN8A/je+61PdmMQxAKBbFgIf2sx
o96Dy45YHotmPWcqM5GhqzW/utJdduZBKambySQNRhwpT2zLmMxx9oNki2qyMuTi
cQfLeknsoy+9QBeRMZFwmAFo88gTPKEGtB7h8qd36DUsoMik1hurG+EInBEoGbLc
8ZcrrxvJ8TDua3yT1wBZrenWhSJe01MRmOzu7LT8UcTpHKy3rCv/Vyne/9mHpOhE
iMxRZ4SepyW4Uc2mExs63QKJPqlRnPsOLfvQLsVJZHU=
`protect END_PROTECTED
