`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rx2brIKwv8JcT86uiEDLalFx8TnQ1o5GxcoXqo/62ZzNJlP5wdpcD8Vn5TktLmv8
jhY0M2wWY3B038TwDnZsfh7tUFTEcNdz0HUj6zyqPrkPEdu4vBwaC+2/l+aQqflA
Y8hChZdw9E52Qw+lA3ifXslEI5p+IQgwb6MX9Sq44rXJQg6TAggNWaOpIf7ecVFH
NazGs07DS574tMZ/U3Szfi2q0WfRDKM2UZmmogLlNguqYsPcV6N7wBE2GWEPo8ka
K8Vx5/pMdW44xmpsw9wE6TNMLtWN3DkwvQiJREdnWUfndkJaBGfQJlY7qf7rIVmS
fiLRCbd7ypPReHm00P8X9Rl/5lDDHychun2e9lPl4OqPN8j8yEyKVPlwE0MDmGJ+
VVJN8jrOFrAagzTJYm7077JOlN09f+FpyF5ieE4voxeoKD5jRRIBEZIm9Ny0n4rV
jloI6LgfcOsnXgLJ1dqVuuvC3iBepFYwCwBmHhLUmsqeQUSNY8PF8df8FW0EsdGF
D8TmDk7t+IZt7rfuQSuAVL3yuXfmLPSrpeiEV0+0qsm5vnrGAJjwzgmEdASatuLr
00BcF602u6xrn1Pm+Mj3ZkHRaABXnsF+90P0Kwbs/YAFTqJ+WzEVjHUZSVAGJ42E
lTrluEByjlpw27cTNUzLg6Grx3gdx9tMYvJ4JFGlJK4aT1gb8lGP/qIsh/5JjuUF
HB8+GKImcfJ2uwsB+PnjEw2A3joc6NLQxe+iSXlWpkoflUuVNsJmnOOwhVJt2rJ3
nXDuZBmfWDAfK1ilkguwwpxtxhT/V6xP8Is6LP2/hG2vewKh+6R2Z2WFhqZMJr+f
jEmMTgcQetG4n21ZH61oVg==
`protect END_PROTECTED
