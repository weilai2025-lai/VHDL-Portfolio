`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5H7Un134fyo3vsbJjSIsJUzek3pDLOoy2icN2kvs8IR6xS0jj2UTTKvv7J/z31Co
g9Fdhp01eYO1N8lKWcdv00qEu4DZ1W7yG3n49q3Kfq4/P4AE30tEaw9qmSKzBqiC
UaXb635zA/F4G1RxRSSb8gEGle3Ot92nVRiDTYJzxuCPBKJ3HXQyx2BQIqVr0/W/
`protect END_PROTECTED
