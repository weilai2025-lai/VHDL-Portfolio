`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sVxbvMn4POz1o2CXiN6vly5UdmwC0qn7FuEo5atA5BT80xre7VfWzVal/UPidUS7
2aakhRxujbDntdm0/nILRklW8YyF6YErRZIB2zzxNRUWJEvahO6/EnpxgbjLWBla
vGaAikGhvy0Ouhs3v1thCDrF44t60KtQnkbn68jJd1dy2I0seIX/lMDuN+fsKe5U
aUD3nGoWX+D1urG7jWhtEw==
`protect END_PROTECTED
