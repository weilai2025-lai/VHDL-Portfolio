`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNR0mMHGgF7nYsqiUNjnLAfx6g1Z5ZK2L3JGFGpMV1LRMpqpjYeMx85Q7VetKdrv
bSahyQ/DzhCB7wEEiSU4YFt3EKQRmQXKZHXwFY8SZVAGq17so/+MLzyhoBvsI/Se
4T8U3nyzHQIiym51vJDI41CexdxAgU9Pao0ZeUyb8oG402iN9WvzbRA1rpyURkcA
SK5th9avD6knhXs2t1Fn8htTFEwfXOWh5sSxOr61Hzc8HLly3WrztdmfACV0WPi5
XeVdHj9YqaHrokmfN8Xap7h8fEGXuT5SbaouM/w5XoyuSIAJgLGA7CA4j3c349VT
VWF9dc1CsjcChIEiWEQxW0sNJNCxUdz1ygyGEHp6AMnDfip7JJ+mb8sGJ69uJpau
ZgHzTjetYtOq0dLrF5l6YP/FUWkyxI1bDpik/PqZ2oFPynt8kzx2YuNDrmqAFWA4
u3cSlLHQ6VWOK5z2q7SEp3BDCW2HyqI2+VSNIKSF3TZodqJqJZifZoPSwhDuSEJI
+8tbioyUlKubmXiDSEvT4BkWTWepfTm1cok4FvdbpvdAKvu1P/4szu4Cg+Jx8DHR
LqVt+fwQJVKq+zCKYdiV9vjSnr7mS2bhFE/RgSexG60T05/NAvX9xu7EcuS8jOuP
QRHr6UlkavB2N7siobt1g9PrlvVce5qsTW7IpjBcCwoj9+PyCMEgJI/Zl1eMpfrH
5//J7rVCFEy044oZMEDW9IsJvthRK0iNuRk5pxF3uVMjGw859lUSpcuyvOczW6vT
94wSugcgmDJXJ4LSNPShwRyZTucHZmgC10F0wYV7AeTqlzqpuaxXuDxBJIZtf9WC
YtFT3Wp3bj00Ys3LFlfIRM8puonTL2A5DY+GgFCeqiOBA40lj3qak3FwthqAb6/V
EaWyJdsSiZOChaPh1+la+BNo0asgMx9/2Rq9AGr2xXG27wTm8U/a1etywr/sbn82
8PTxQQs1TvfgIbfrLzyFJ29fXsO7L9ft6L0tI3JS6P90gt8+aKo7al0LPTUzIdue
qQTC829Z/bXB/8zZ5YYvwZYM3ILPt12lI57+PHDxUuAKPmEyeLPcm+2vAuXmPtS0
/TAW4kKp/rTn+QuKUprxtPd8rcKQKeLYgcCx/6Xl+nXxfShSiDGyewAELC9a/z7X
S5nMaeihtOhBlPpUzM+teGjK7So85Yw0xvfNBYa6tbXCKU2NBo6zlzlmSqNvz+VY
UvLpRYq8qDkgnF0VrUUOqCzvJNr7PzxUEGpA2U7ok1pzwCzW1nT6r6gry4Qdd4Ct
Es/WNLyL3no556ZjeVLJlaYqtPgXdObufes/vFI6knuf2Ka9HCndio3YRoy9+O60
eAqRVDFVpFDMneeGG5WVtmIzoWjFF+EJzeq8yAc7TLdNAIyLxN4AYpyyP6DTCKGc
cRtuYRnIc7AoaqELB57rYlzzoCEaoNZtXiY7zEXCVdiLDX88cacM2yswxmrMduOO
XBRgRl2oPCrOv0CqGoJDP45Ns5lGVinQ57QUb3LJ2UUkZISS9KsSq6zObu0k/gLD
oXTZnEe+r1cND5wsvFduFNHGQotm3SHfFtif5pSj8iWI1pMTJWU/mZe1/o6s38o+
m0OaF/RMj32aZ29JOI7WSQeTC1kthWCw3aY3swDlsMHbBz6j6RKFzCte8aVNqyGa
NXW7KxIajwENw9ZitkGCzt5ttL413Q4Y/v/+NuBli/8puaRQEY6i7zPRExaHYCfN
378PjZBeCTftT+x/yicjmTHg9pegL3Urg9ujVwCFv6hHCyuUPCscNyqa43QDs93X
wwdO6b1zoba0rktG6VAP7tb9kBATykp2APiPZolMe1WZceISG3Vt+ggXBpRwpzoc
NokPok3E9cvNvml2DP2eT/J4lQZ8UgmGLkqGPZ1Q7OwwjX6pPE/PN7gWj2Zq7KCA
7eE3dwwSUZFStw3JWaQioKx5/1ucnzRKwGBCCezGLQfQHOUgjm0hDub1kgk+lwt2
5DbMH67yMx/1Kqfd/2ufFtu0LZvb/qB2iN0c/j6R1BDSNrbo3E1iCsmPgzN/fmeW
r3jnbQAiTe6ySlHJrwS+d9uWQf8TJvDKJaaAtFU0xg09n5k64miwCqHx5HCeeEnN
xs4KJSqWhMeKNoZaQzyWM1UKP8HEU//0jMPXahG+AmDsj5HOyV3RNefjzplRs/73
w+eDJHE6lu21ISTkJ13ntLfXLAIEWDPYQ9REkKYta/K97Qn2j1hL6vWVHq/vfZnZ
xldKvpElVy8rzAfYyKdUFe/IGlLfKePECaB70wJK5QDW8z0bzvZSptMBY0DBlxWw
5y03PcUoAn2Tnbe1ULbanP2CVZoXHxlIMP1kQ2VviS/5gtfKr6VyMhEGcIpSUM2t
q3wtOr2VYg8ZcMZOoREUillkaVPQQAChYjWkQmWJZQzhbhlHX+j3+eZoApn36FNo
LGF9MdeYT8b1NlK8PRXZwN73Indc9jZS1JyUrPIXg+QBjoTJCxge1p9yrhHjOAfV
kufiuO2gRA5AGMOoAE24S4fDYK+8Y5lwJsW05TYxoQxv/KVJCpjf2GseVadRIqS4
fvOuUz0n+/0JO4F6xYyk4auH97yk9smLOhA8l83Ha/hL2cdQHvPZVecbTGzBPc8X
rFYiRzFwlfCuLHt9rjnP2z849fXDvU50mVb+MsDmR4S9k2OBlvIsjt8l7lIvo3Ap
EQwqwA76/GTIpNG5Tv9W2CStaV7bcAKmeTWKmCViJLKojETU4t3uxvDLojax6rgP
ZEdPYlF7tkOX45qOa130Rbg2QweHJ6FKhwKbbnvvv4buBq9U91soOgtTQlC1kUiU
x7a652eOtFOnaIF0cXNy4aV5bmJx0lf2Z0x1r5dGRgWtnyoaz9z2hzi49lWN1BIJ
vmQhayCv6xRq+eoZtV0tpu7LFOjR1oz22/YcdjLqlCswy8caoGcC087RSGvML3si
zz4bE11K4kgT9EPDsDIyCD61G5V7VzWpypi99SSH4gpkfQBFRSPLyaDhayNhoA/N
QVtk5WSiY5uesVqNjsJqBob9TlsFf0Q6bPjUIzLyN8TTytj7ZOMePP2U5do2MPWI
cEwN8sDhCsW8FLbjw/5G3XaHo/yLVAfsYRrXMHNRfN/96dKzXZT5O1DfCScfVBQz
7bfJBh4cB5+46EEFRwdG62VlsXHOY4jO9ZH+v3uWPk8Q160KZs2qXjsOFw0nCO/e
yFxmRYYLdlcu7L1hPEYvZY2hu9POH/qJexBFN76b1V4XyBTw5EUyGIsmVDDm1XdI
IHcwam0h/qQyK0HWKICvxKbXH4/DqcetQxTYH5o8So5R1XaR4IJiXYUtLQxA0z/B
XhIUA3AFXBEMzekpX2IIfWHCmt54LG0xeu/vTOanE8xgan4vz0FqyW05pcnM25t/
lfKT+43cLIJZBubMGJEotJknvzRRSyUcrGVuLKrDYgTpZL9rbbVtnRRiG7OaBqSw
9UycDjiJirIVt5EpHgJX8UJs5YdMe+MrGgeBhSbStaONIiY6bzzzejn2yfSlCRi1
bAc0+WNEYs17NXpHdyHPNcYiE6xhk727LSzQ62EHm2yL1cud0iiv47mulP645LM4
m7hGFwPslJi58XEYHGidEGhwXZNttUWOM0QO6FH1thJPC3D6y67w6hlzXnNu3XU8
u8Ybv6QuEqbXOZe9MEqLROLUdqX9YnI+iR9MQffr9Wo4LVKSQ6DfNh8e4gv8nkOo
EOlvepwNWY8E2czVQgut0nUTrANKlhkeP9nWHbM+ySt/shJMbt8zS3U6KbGRAVo8
P5qK/VOL73krBSN2UIZEHLvXkbxhdv1U1lCVMBuajuyRWKVCWziYe/Flzkr4Fz51
qVeMjvL1BHCvvyM+59zbn0wnSbSeBuwNzg2YmBBOz0h+vaaJtjS7nS0vHGYmjQry
nXwX4f+xwT7f/Jn3SGvvrklT4w1tu+MGkj4PZ/WW0K+jZNRdB/VjvA7fsyUNcT6c
jmpyNbN/1wpYTS+DCvfqT4lOlbofGy+6BVthy/L40dkWYr93NPxwNkKQnXn8+Shc
7ekBJsBUGVXxomfty9f/iZcCBSix5sjlhttTgTkEu+uRA+r7nA7Ie8/3uRN08LwE
9H+UbhDbVMhOBBO2GzkbzqD9P0y3iFQg8kkBVWtS+h1wNipHEZJ2nvmAqNOpR0Tt
cQlSlwg1M3AnSxsuGAhQz2lp9yruQVmNasC8XL7kVQMI5SJJ4ae0Q1Ou8axXRrhw
cbXsWKfJap46YPdoITyIzYP3RkyVXQr59K25nA9xYH6MZTCFyfVtk8gDilYts32G
PuZncZq35XB/42BtLQPD2Mnn1+SS5NLSAtxmcDK+yktbpu0HMStFH9grV2v/a4hU
ll/k2AHmVqetHYnRe8sAjuyIZEz3EDMkd/Sd0GSpLGHXuccs2aWyjUWokAmN2wpl
nERFivnfRe86n3CbR5t2gN4Im8EhGWShUr6gixdWF7JvqzBRB6WAvAUTYJmZ09dP
iCy+R/K1DLKJwU+bcm9Tbkp8HDkHRPPAXSAfRBfItjADzN+sZEe7vjcAzP2QtSiq
dzKqhSRgDUQoRnNh+CQqHkTHLn20FARQLKOmdfarw1P9QVOsGcMy/XcYjamRTIgt
wWvu+XWROkQmfe+tBqxPKF3+w9c/sj+Ec1sWGJUzSxKvOzbk0JIS1Dd+dATiR47w
N9pc/OYZiQG0cq1j0CdbWJ3btedl+Yj9MYXiV5QRKfyUb6GvS878RVdsx2TpIzT5
du0m7m95RWMzEcoSZg/ZtawFY1zn1g1/451jl8Ck9jDKVgfXDfLCxK+nTd+U5Epp
bDfBavSWhMONZ2rcXkoDRobWDpWl4hWoF4UowdgK1IsJG/YR3HLq/EYsG91PtgtK
lT7ZzX0ACrMe/uyJkl7c4gZI7kDnciumuyWpBGBGpN/k1A9Ikv20Xz+YF0cS5Mql
Z357lNf5JqnFZk6r28As0a38VaDnDKEwoMz+8rpaJrurnre9UYhOz+1QQfFHQJoC
sepbM7TUnSxUbsrLtQWxkgwMsXA+aSde2uhUAdPKK5p2t9EA4cqI/TKO30JutYmz
EglWeNzyu665AbUa96Yb2d9+XytYajcZeAmaB6mkA/7+0s7tEmaQ0mFLAFd9iVag
Hc/tluL8eLJ/OoXmOhbv3++wnbQOaCw/MfVPCT1yYXZ3v07P3x+VE7RFlbl+4ozo
2BOtkezGnmsOvtglNjYhqF4e4ESgI7lVXBtk4hxvAhDpssyx6NLW22X3iqOA2qnm
2VFmY0+SS07RsBZUq4V3D/5BksJxg85eeJxK8MV82VPS84hv/ui8tqdsOem6lmKb
bDavbQX2oHfiNY9XepB8i//s3qZjqH6PNzw4vnfODWLqjNjl1UNyZa4m2BpxyDGM
+1na3l4AF7TsnfnEPVlbNCJQ50krUG2PGZLlXVLnzFJl15WbRpHQoqpNxASpeHL4
guaCk01sOGmpjUS/Miu+VVr5SAWGCkYN3UymtmYvimVmU9Vl9DW1SOWQCKUFmTJ+
8s2TqgYL1GbeS9L+yBbEeLlvcLRLIy4b8ecQsbWLuwpGnOd9sI0+J+1iHRV4WxlV
/oJn5zzq6a5cSq79JSr4SaCbYAnzpYWRuVhdsPIR6pQN56JiQexIQsWWKfT0WoSW
pT5Yyoss6s8PmQzls3MXFVubXthRSRBcVT/CnTNftN/Mia2j//2RQ531096I30KS
rSrJHx0nFAWvG0sUNOgfL/saeNCQ9xrtmPV8NGm09Q8UGeNoaN8DYZtcmCnXHoHa
i3PqXwy4JU3oV4japezzTwEkM7LKjg3SUi/IPj6qkLD5v1h6VYDOKP3TPpeWUQdk
65Q1YvRdcGTz4SiQ3HKladgRdnYb3iC6GqwruO5hzQd/URIoI5A62OtMWJ4ccxQk
AWh/O7Nh/ICgYp9Av7qCR/SKd0WLfMp7ul1W//dHZwMwpcpuJzkKXxuoeUKZRCFB
Kgtu0SB6wjLCKyTrMW+Ivzdw6Bz5n9Nd6cLzfWC/m4twIbYyNfjiL55pnuGAKbSH
uFTlz/32+maLUMq9qcJG/T1WEbUI+RcH8HdraALos5j7SJ2JhA3K+4az7kKOwBgB
VxzUw+v8Q94m85xCqjDildPdf5EOx0Skr5KYD7Ml0nXgqXCUfLbrQnXf8ldIb34O
10mFD1PKV+6oeHQRvYsxk3GNMmE8lhTyJ4OUqQRVxZF/ELFwwZIW/d8WDdRuCgKs
vK+lOKPeUEXLUFZihMDD099UMaTmuO/6JynGi1Q/haMU1laoPmtwo9FFMbAGVCp0
yqF6YniSlmBKPj9f9tsOd1tgptfmBENdfgeqKbcvqpgvPALfoth09nItwqulAlNT
45JUP2hKB79UM7ORyMRvCG6dQvc2xs/05rurv8E+qvvn1ISD7iCJelOVQ5hHrbx4
VXSf1FOUh149RujGnSGgWBzgykifxnWWPPIlHTAZfsADBlTrDrNFnBUo0DhC90jJ
9M55s5N+eC+8FzRzQx5f5FijPNS08+ZcBSQJp1KWLNxNYLhvXulUZfcDCY6xShfg
ER6mGrq7FCymiOC2PSPnlDYdG0AaYKkp0AEwruQeJZXt2J9Ue8GqzPS96rx7AEx/
Mz26dQr52Y3/FW88ab/b0zNFNADTmaEDcwGZ4bszC8m5gCPJVR1QqRDkaEOu2BaL
wcfj/1V9swkZfdJG4Ifn67FAFVJy04v7fgZkBoOCKhRPAzhaVlK5c6zLXlBwiez9
JkHtBc6QLUdAJN9EM8q11Z3fGRny1AmSEw31WRUNhTJgt+sCtx/fFTHUuhzvFLro
i3TbvOR70M5l+ufS1tTJhsFegzQOqOpbtk2dynutimfIS4+yg9XkBM6dheEcFuJH
koGfyFcY8yJJSnrkT/o2NYAuuoJqXL0zagySTQ4zO5E+D70xeCqlAByK/Q9sPrsM
ahOMJ9W/XVX8KnP3XolNuluoBTaMuFjPIxfL2spQyM5qO3UZAQjKQyefIc4ZCxB9
hqsu6MoTA7Mpi2eUYn26CC+o5lTuVmNhRWkwIcUUBEyGvZuR6tCkQkFruWdujfbJ
JZkc+OGsh1ehng5wotTI9a+JpLs1eccc9f7sdAsRKSMUv3kzDeHjARFsA4s3yPFc
8lVVZ6wByebapQI0TDZJ5F2rYnK3PI9dXOZgcTCRmVZhfaQX0dJgKMfuqGmt9nCN
nWnJw14EX2hgAY2ZMp6bqg3Ibcl1RdlGzzVx5GmfvfkrAkUgrdibc0viv53RbmPY
C88/BbOXT1XFU0gPGw7KJ1k6NOuHbRJ0hN7Xl9kuErNezZ6jzj2fzUR1Id5/leKV
E8ZhZF75O+jVw2e/EO/p8gFopFGRKpp6gOXoCq2oD2fV8a2gNw0cgstpFfcu/dId
jqq9JrYCDD6b/o2lsIHip6Cf20prycN+JUTgc7tNnZh8kYlzNFlCs0SYDKXEVvud
jxCf+BkaxRdRGm9GDZuY5pdlglervIn0ltj0YPl5uuOZUIT7boqeDBjx+ilLxF/b
LkBMpJeeOU07Z+OoSGdE1IHaSEx4fyP4wOtgtEw2PYp2+Rt+mCtRr6O2j1hD1Fm2
Hi33o4XCEx0pSETRETHZkhJnevLckmJwGlOOUwSSenRlqlIoPpNfQUMVQ06TA186
aljZ1eht1no0SU2E2fs2yWLB0dJDGqbRF+rOIGPVZ570+OzhWu7u3cagxmiXrzHq
VSMZTfOfeYa3Ufze/dPCOwKEeGkYjJ/oc+/2bikDmYrBeSrv85Df2LbZi2+kWnBR
qFDvDr9Bw75ZL3inpBTMWHqOFvPv3BagEYxA1c1/N7MpuM3CILVGGZcYjRsp/5tz
bRJyCqc7gnq9w+z4vBgozzEpa3Utt3TfAMdMf6VVgjCg5v4l3GUwbgsx2dzE4Niq
9HcxVqTDRGob7ObzhIDpIrG67GTREyjXGoayrpQN+lA5X2VEma4uxtV+aVvMJ+jQ
ofEc0unx00kL9VsPTlypbEU+i4x5CnOzErCDMHb+foaoVqc59nO2EBz423Xr19G1
0QBSUjrAg4N6lyFdIb8Tl/HHYcwDg7SXy/hLGjZQIjDRI8QsJIVM6d9Zm099SmqI
QVYHMS2RKd6ohTBpLsK7oFpUwj9BDX96LuM55ZVJeM8ExXizYB+0+p1Pvhvq0LFR
ZqkLd7gyYoCmE/toFYVjKgRj77BaQke0HWextVtbJYfG6mzl2aALosUvY6U75mh6
8EF3rkWc0UJUaWnkAn/A6VMhMb/unkB8gKm7BQj8o5rmrCRUWN3TbZwGTMiThAgm
lXVvgG3eOJnLC09hbTAHgdL/SwTo3NeXs+zi4rCX8j3M0kYdISVhVcn0w7kURzcL
F2za9MjWbkuA1GDVGejj654Z+ov3dLr39kRq9uDrrOI0tXaz7YwbCxEd21FsHHn+
MwOZS0+KEITdInpBjvtFl0dM6GpY/337I/jCF9fMMMEG41VBZU4MBTaC9Hxdlw7b
ydcHT8LvANRt9/yVLVvTPJ2NULFCLBJ1l2/l3H4n6bHWcVY9Txjxza9mU2QWbEj+
SCMquFZNMlakNsEWfquAtXKupX3t8xhUrOqkTVjPinHrXLpTW5jQ2uB5Nm6Xjs2y
I8lBcIDMVxTxb0ZkS0EkCWxxELBsxPFpTKPrfcOU2Qi6JJWrbmtmgxeQg083y/70
1p3eEFUCRFBswOp7sRYQVZeQH2YS2Q6nmNISP8MXN4nrq4pI/RHAKLXC0mBREIbu
fJs7liAY5Wcyji1+b8XTmQs+yXb89MxxozmAZ/iwFBq08bMTYnNsiQyYzt1Q4n86
WLsquqfq4V4zvDJ1ApkVUFS+f3cREFvVvEYhOutNQ+/flfQiWwpq9ySjgc8eACnM
mlvO+ECZX6ZPDrsdr90+M1coanZ1+Sxmm/k71gTlIxHZzlJoUrpM++Y0Si1A11PJ
PG0BC9fSJoXhr1cVAFvPWLfKxU5CCjXKOc4o1+gyfF7IkvapCuIOLTRERx8yF/7W
fj66hjJkm5CsZJSVF0Rd2KXfSQ853LTEcGE5pTO/LdpfZopKdPxF8kCTBprFivhl
vp18An45TfL4RdPEkx20pRWlWlszsuvyfmlgcBp5m3rwoxPCln1SYOJMbTI7suZ4
pOfM9vmlKwcLgK7jb4bLGxHHf3K9OlzVm8vh9iO1mlSRdctVSkCMYrW1MOc/Bmao
zLkhgu9UDLaEaMYtcbpX27ZR3zz/xJ7FpHsCvrHZVlY906GQ4RJdKERK9bFX4MK+
bLhUzEnxUy3TG7fmxh22BYjT4bJHSrEzGfApT+Be9FUgI4IXTe2wvGq180tGp9QQ
VSb7HCvm37qZK0VxchmTjDH8UYbRBK+S4oBn3QfWuMYMz480GktQhNcIn5FVT+Gt
f9jKwa7TWIAmEvUNM6Y7ztxvJ+JtiXPZxl+2PkUS8vL5QZDAJsP90rlG7K389wbj
N5wf1p+2fBw/F8vzNAGFzNMairopOKF1cnm665euo1TNeQG5aOR8j86POArwxw5M
2k6nu4F/4d6UxStPBlm26FBucFhFD2vsoghuI9+9vV0HbtVS9YjtecB1TfpIBW/2
tfWQj+gH1qZf5NHikuAQSVxTkUhkHKHrhi/db/ThdbhXtga/+0xnUP+GnDxWZ9zy
bEMHwmWyC83oDS4heriih9m7eYeWmzk42W0h0b9rX1m6JBtAqHny4oxiwxoGzljo
xbI8DM5hTkdEzn6YxYDdSGSekza7+E3aV1CGL0MkYJ7gteA/i8ehOEK/OKn/ibU4
mNnCQD4SVlyHg8e427a4gw5+1QXMaIINiaeMVmq8c/0VuCCHB8tzcjauiocaHEZi
pz/j//GuI8dZB2OfgLf6upamkhwEcanUjqLqwEvwPKVXITDz5N10xfG5+7doMcOR
Ey+uc4j2fEZBNZ1mUFawRb4xfWNImt5ix1AYI/JQVWtT1B/Gg5HAAFn8MKYeixZm
BKccfY/eeUC91AO0qIZq38OV0Bl5xY1qzvxE3dL1HZtdrzHRxDLNBBDyl1HbS8r2
lC5Y2S8accwDOBIDMqs4TWffM8a1AZYf3VCYYD66KHkQyJ/v8DUmtGEIucP+maXf
JHRNQ+6PWHCBa1ZI6caAPjHwjJr4+0FPOL2wUScF0I7SJLjrYvWo7/D0rA8LVPik
POTrOWOmGQOEQVx0i0wJa37lawsfRd6cfONBpQ2+nxcIfykPFC5L8HTjeJJ4uW/d
4pyKD8h323VPX/QocMlRf0hNM+V2r/Jze1P5T+vwXy5gWTmijoHl96ZMZfjxCqw9
vccH6vdWWFycSLxU0e6ODk/eWwagXmNBO7l1fXWTQFseX3pIDCmMiUcIsZx4WJed
60J4TLgy8RZ+Xw1c8CY6dfKLycch6Kdzfepu7e0TEdsuLr/DCj+iKyRkXSLH9FQe
RBbN+UMCc7Q6DwCQkGSfbvhlVhi4CZTqkbKYINU0gaDqB0tH5E7nYeAZGzj/Lly4
9tQi1JtGatqoBoAhxB4tCXXZ63TMqddoWw3HpLxVDFsVl4dmWmP+FS7mzgLIsVU0
Mp/AVOW4nvX9xyzPkK3UjSR57EmPju0uxcfIlQAkscXzYjtnvBm2dlQ/LYLonzpJ
KeF44yd6r8lAbhLnfn92PAXy4ApxpEvBbTZZKERgvZtd9mbTJUeY6N8MZyoz0XTH
DnkRSz+9RUUpR09RLIPAVqu8hzUGP5w/sXnvqHmmro5swsNFGtc3fQAOy7KrLWaF
2xpRne7mAttfIyR+9Y+PJuPXAHw6EWI79UGDPIxkfv9bxaxPdbRrYUjKEp3NojO3
Wm1iJX6ruDBN7mjgQ7/Aiy77rVhj5jJVM6S5qXATw5gauwxOhC7o2P7pH1Datd0b
sAPtHl2HBpr/7NI8TY5vIEcvIQOKp0RmEeGcTwHcOdj8RzxOlA8TDSUW2KcsqvCB
xxPYXaD4YyKn6ek7pUtqG7z/dbBtBQQo6kKcKtZmja4rmRHiE1wHHs4ABEVS4L6z
ozklZMWiNpfOneHjJcdr62jKew5jzuBmKlvF0A154qmLP2iubRNlJHNO+TCHtEkT
fLUBYvtOVCLmeKfj8fee/CDHQYCvmEEo85Oh8byOnNqGLqYIqb798hJNwxHllruf
cdVarWhh0+BXTPKwKvchg5F+d6f+bhCgST7wILLMxxdVu/aeM3gSWb7BNw5GAT+K
uNBgWaAMUJ71E97nb1Hx67TzZUnvGZCzOmaaejM3Inu14Q3M11xbcuUufDjBkMn6
LeqPTUV8CZZ6p4aXDCxIOVE2jfL2U3G3YZGggMC0VabEVRtS/Hqc+XiDjh3CZh4j
Ivb7mR7NTbjsT3r0X0J6m4nfVxg5Hen9ck8SuZAoHiSPBV+mSB11zJSU4yTE9LAz
NHKXFaIJjVyJTv/Yt0RyYK5a07keQ+G7N3rOJtfRd5+xLvroD3/JOlU8XwpclJyA
x2AY6O7+hjF4d3clDJlBdeMcuX0zeWs8gIxCFkygL9GaG7n6/7GldzgPa6C1mgNL
znigGU2G4OxKDy4ipQTyhTkJhKVoWmSsIsDoerfQox+YvbdaLf8euw7vymFlpZpQ
e/Z6QPTu841aEek/h2v+xGxMl6tsRwlyPK6XFJ352sypIjlmqRoGmW+6SMM8fW7b
4Mk/BEClIF9RnXSBaho7OfwUuq8sjH8ecZCIE5534rq+WvFv5UpjYpOZ0QPmOq6U
NXjZSN2G3aVl/WQkcT17I1p4ep0XSn90Z3LdJw/acaZQjJ1Zq1fH60h6/Fdnla8A
svy/e6hCUOveF11KA4P4fLXTgnjEhIzJ/D/JX83WI/M56nxam3KAnRteHomYdQve
ZWBaMtX9z41xCPCOSipmtTSYG8yAwjDIUMpAQOB6u5g8Ju3iAF1/t/dbH8/1LNys
5eCv07dytJAzwgM/zyo2HLoURddha3Ne4WOZHHuEDyOFqVxg552LqLB0Q/pwzNIH
kzPM9I2/cB+0XHkyOWto9r4e1HbPlNrm2P6P/BBIv5l15RUpfuJKUiU95qG7WY91
tpj/VjTHNKXSsHDWZSUIzysodSJHdVaijCSRpf84yZIAOOmbbrx4x7883nLY2g+H
kmN/cp/MEku0jXFW8bCaC2OhZWYsu1jCcqeyHA4gkTWDZ/Qn4l1yyYPkP41oG0v5
3CB41YC/nm6zTcHoy31y7oddLtSBk7ThBEuNVKNxHq9GnKX2IbEpKvhzgsSGTdz7
/2LiEFMaecJ5mqTP/ZS1GI2hnbJJWXbDLbpdqovovxOoUwgrV8i3ucJDgb6uAyMq
DZwBR9ZeIodXLBp5Iz6XHgplVR6IXsGhlJcYSgzdqLo9e56l+4zpGeAu5YfHX56c
VfoFOYQBRtCBeG4JPSByKKgeLQycD0shTOlhGyLy/xCaznk7wzF2Z1UOaYC7d/ub
/yhsoNFWncbsBwchigL+xGZRFVqOCUKaP+r30hXOFXafPyT0mx7rYbHme/E8TqeC
xU26n6Pq7oZbVGC1U7cpNQXlDAATjrhfY7yubGUaEZPUSPYTnaHry7hmMcCkGTkX
3l2dxPdGmeEK9YCJymNzsodRjFI7u5Q77Tkw799GR0XM9nWm1w2Ct9tFJ70lforn
I8v2Y5evUrS6nJG6/cgulfCEVA5rDHzRu2WVt344Dau+7ntiTWwMpn+kaqn4EQET
WXFWfwbowSOKr8yWbxALRGJrIJNvYqArm+3jvN3EsQMuAPB96vCseoNpaZX7QZX8
VTw1HtyKan7dF3hDqgVF+3gRSsdT1Gw46t4j9ODpTI1K/tM65o80S6vNrwOXxmYD
wm+I3Tc6bvWagvBrl+mYs/y+O7G1GozNceBmHUVK0RwsFMEjGEyA7ojZ99W0j6Ug
QPl8ehKoloFE5LIN0C/P4IdchfueerxGrMIPaw+Mr5ZzEy1olyWq6sqV/pPHxiUM
dekUduiSX92MWmZ61JtkwKlf1JmPTUkAwiEzGumeL0FR6nm0+8i8+/39h1RB3fGt
D595tUkhCUV8RMiRiz7P2kZg09IxFCGwkAA79hROvpVI/H93qgNS5RMV4ToydMbQ
r55I9cAhutZWz4bq0hWtgsGDxtagcS8YBJpuBOvHzRIQz2TAY8+I024H7N4rcOMQ
jsqtyyy5zqx5KIQQPWtGPoB+5mI6Jnugen9N7lquUyAvAc4zB3J99lcjUltmMp/g
BEocu5Nj9WAdX6iFUoZFD0agcrf2zl2ImtEXbVkHALKYRj4UXAUD2W9Ao7CQS8ix
DwUuAQyQZnzhY64RqZihijgbsvvZHj55WAqWiUfVDqjbZGr88Jb62JeY89sOiLAv
RRrU08FHA7mWyNVyLtKQRgnyx05LnxJe6QCjwTNA10/FfQ81yUhKKdISj0GSyoLP
l8kdmGdLmbrsWV+ilEHYJYgId47IrqXyOzz/M9UbuS+VOeHeGre85/mJz54Olgu4
9yawJqWYBTicDazcKyDArNEfEOjMWfqUEledOEwC06MW8yN7Q3PtC+CNTW/nTMFo
r9wM7H686XQrQ7F6ZbU0j81P1+gmUDyIATsyAKrONTGA2zEWuVtTqf4UYEp/FfO5
CAUq6P1gswC1wfCP6B3hhD6AvY9bI7PPYhnoU3+rjoP8/NdpMmy7ZovYigkpvGFf
88+vT1GnjHVUVyp7476ziG7jD61jVjnpscqHYQ5fE7qL11kmrOi8vFB+1W2iqwDQ
0rJzEKytdabQB8JSMHH+8LEnnd/xcKn/8a3e70jfkHEJtVT9r2EiMS+U7X/Q0dj4
iGrAmKPvay1twq/+ciKyPFbP8o2LT3xc74VXbh6mj2DFcEaRyNrIVd56dO7sAUdK
Hl3WqMZAFb9tYztN6dZj52odxGX/yLAoNiJizayNX48zkIFur9orKARYLFOYI1GL
waEim/YAqflmcN/I/3OFuaC0k2HV9SKq6IpGgzAJwh05Dcrly7uzm8d6f4ed0baJ
P7Jwy0PxuZbcu+8ouxI4wL9m2zBt1V7j4OcbzJWY03hyGzqAO6pvTJbMbD/sRq86
86XF3SeZIbkvziamqpXzhbX3Ju+FFGAGu/+X4lJLLW+KnUcPEvBF5x6AzMOpH10f
bemHvDH21lQTOh07e0wFV1cYRQI7FWcaXViULzJvW7MM1uqH/umB9BFLx0E4sZ1G
dqBqbx8bjdFPPafsHhnfTUmDomWAi5UTThrjHrUgiWyGhBUQuhSH+/vOQIbpGkoL
wX/tj7dqo4LCsyphunNAIYGuSch4+61uFHMQj3MGerq3Pwyu14xgWNinH+oUKrZf
tH30iEDbkTVGJ7ovBoZB1K86MipzWyFRtoESFMOwXqwLemPK2+rRLU5LrnYais7g
GvoC8ZH8PESev8s4QWjxvPd3B+oySf3RKEeHkvx2S8Pe3KT9mTohdc313g9xxCq2
Kf5Rtg4JIeh5OLKZzhBDeJhO17YL/3SCM8AGYRvx8JyqW8qOah+dYWM0ZBQOizPb
UfyPL5DxQLJJ5VlxzAqZhiCcmPBH7XSxgNMZVHuOGFYsJmghEaWQC/e0aB1YYXBi
eZFkjg0nlp+dikTXZyZShUxDP9PKBNLds3MyfZ3jElPgPJdOmcA6yaYcoqvNwyK2
gb467RI7wdhzh3qIqWnmSrr1T3x5OmXTbG0ZnP151/0x0y+1JaHSd78cemB9nOwZ
m/yZgb6nuqQ0cSlifOi3polTW2pBaYA1mgtxPUiLVFHRBwCdfOIC+zP4cITTb412
UisDlyEQdEsRio8arex00d2JcxL6ZlxRMie2/15+pTQxSH87/U97Br72yv+Zu3wu
WdGF1LdU4CNzxkfC0KdyVbLwxd3rMns6922C0oYtuImF2my2Naz0Ge4FZY6jGDza
9AKvU0OQcdYiBRsgsrv4X4vL8ofJmum760tsPvZaAmd1FdSP9teyxt9JUN0pWzYs
1iBy8s52udwwlS/Vm8CkwF4AP8stURdqAWVixcTPnUhU/Nt5dbzgs+PHMM0cEe3R
nkQWmInIJ96lxHMz3y7mqDW1dYwYP0Ax+lJnSZMba+SIWRtkc95I1mzinHWBuagW
VCe3xTdJG5RuDRy0aCq9HfmX+L+iKEXPIIgErGQG3hXYuHhowAYiKns43Pckhvsw
mOrskwPzf3zaLmLfHCf0j456Wsn7Z1jrKxaPxxcY6t3LEHLtFvPS9PwFXfb+05zr
9JIqAsXDGuJs0c0q/ALf4bKkow9tmOV4/1hqM3cNY8lpBEa/kA+u42MJSUWtfkYu
nK0dEmqoUVkPLfUMMRYXLMFWGpZ9tg4UA2H4H4IE4HUKzT+ChoQhAFzsxxD4NgN0
1Vjq6Yf3sRACdXI37AiaRgutPcaeIZAWgJIEBC1DOS1bDWIWK2rvGikNF20jlxlY
lM8gXoslXdC3qucXWwTbH6JthIUG1BApfbUZcbMryFA0c3IwXJwG/D0bjQ4TOez4
c62e+iJUxDBtZ6xpNweEg1l2+W56e52RJ5pPdIOwijtPU7QXcqAFMFexVxPahbeg
8jh9qvuH+NuBp25dLhuCPqDGWd3IdrePW6lfHyFdY2Ugq0iAv1rofDgrCqdrWBfo
wDddowhIDv/2UDqqAt5x3sKMK5j5dAAfboK/0p7UhAdWMe4ZpnYzXKfxs+f2QVu5
Qvsfp3RRwn2t5dN5sXA+qkm5u0mniqVvufUG9OYfQyBoirNFj5XP9XJxbrY6BFj0
sbYAMY+STRiKG0deE4suPiNG3FiFIlAXE+Aj84yi7VkDy40Nfa9iiASHoTIpTFBw
ma8g6O5VGTnRWGPYwXI12k+mDr7CjDXFSA4VNpDYBMA1Ow30ae6cjOxnKWCadUiw
uhzTgyYQIkngHJoOh/WD/KRo6IqVMBr24lQ8Ybfp0FD9jaGMMlzOOvI9XKmKIDrU
6sxQeNtRZllPZcL5vV9pN4ChEbval/VzLPXpvx7Lt+hrUXxcHg9uL8M+SYYFz2DT
m1AXcHMhNwtStfUMSTD4A0EBjkah2fjlkHoTsgdh3sbBlPbaHxjwg2+SAvRDJHSX
FGKm1Kn/4DGgXfRgbHqreOl1Z59X1zCqTz4wEj/2WmnmC0W8lPgTH2W5ygV4Fydb
ngtAfC/Go+twReP5QXPVkYrf2sO/8/mIJA/rgjm7R0PZwlRb/vSmVQazihs8TDas
tBnBR88Xbm192y7dqVKwDhr66rfZiHawh9fNjRM71+GYqeTT6AzE0Cu+sSqG8syd
/tiIw+10Dv9KBDKdT0NwuvGpOepKZGDzluBDVw77YjKF3g8motf6W8WxPqqUzmIe
1SBnSgJD+ANma9Fj9qQiISXs6So/9NGYj6oaM+eyrNBbq81W7BA2zF0meYbv9jcU
kM2SAdkJHh638CgdeeKuCoJ09+ivKVbbFvVi0HzCYTFd4E+XYNgEk/Q2mZEjijho
jFFANcemHsXVPm3VzuodsyhHyUwk4AfFcQX1YI6wNeQQSTJ+t6hQ/Vb9cN+lD/0L
b4/JbLsmYZt3aUkH7FL+KEuv1AhpfYjH2SlhjQNOa3qADo5rkiyNiDUvS5WiqEHr
iACTx0n8TSm22uTGTlT7wRpvMoDXu2ddV1dfkmXJmifE0ktccGM9hi8xNGAzmy9J
ltZ68Df92ZB9oR+MX+QNCSw8J4lhoehh90/li2KaFT06ISes0lokofPLoahg/KOp
f41zi6MkS5C7mE8XH2sxDFcExnGjQ0gnrarj9M/TW5ddHFlHyXnTrNjTYqdBgEjK
XQhs7f1M1czQ4MS/jTtENcQReAr7DGxM7OJKIpcVnwYQz0viUhe/HNNH6y/fhZDt
Q2AUJmsD5yXQ82t3Dr1xQHlIyB9kH3M5w09sACYg04VrUBOFCj7Uema/aCUV1VKY
aZkMtzJYif66JTxSPrZZWqe0T8d2um5bSofjzuTVOjZqDE7IRh9ZCwdk/r/cYBix
Hk+e2MER13/Mi7AwXWxhjG4FUQGELKcOtol74y4HNOVtDt6oLjWfmA/TyvBix8DZ
ButpEDHHNt4KUaiLNHPTmLcFrCFlE/AbvGYCKVT/AvkgCDmfMLD9/p70bSR8LJt7
3S4He6quFaXedCtbYGzUwiPz9wjUw5YOetOq74i9WgxsikzyRpFefmlWEOF28eOq
9gsmxjVUcvK/OV3rTogqdnKJ3QJih3YlDuGNXZNzfEbGxW3w6SCvOSLCfTAY54eo
HfJXuwH8qCt3eSOE4CclB6ulTFNPpvkyxe12wkO3dYG5I92ms9BaeNqGgSNUlroN
n3SUPacxiPrVltNbcVvwoPfTCVrwyU/Rjc4164s63VFVkM9sKJ5kUPt452GFo+u5
W9bBv8KQNeiZ75qZmkOVQM4OvI4WzmkY5JVy5FF7+ACGUMhHoKxqk+wXNXaVzpGj
cHSgGIkvvUbniIUBjzBTEIsvemkgQFGLmQTXgCKm2xQY3QNvG2DvHT74eHYPFZL/
382c9bxXtwKLNC5qMaReiuH6CQyJ3pr8dUpDWzSakWJkI4xMXK/onAJcac66bKCe
PXR8jvd6GG1VVCCFGkf0D69GywoeHKCq70l9CwjR3jI85Ye5lk8bhwVH2L/KFFpM
whfWRuJQ8v99eLFqDBwo1CfgSCKmBw96vNMnM9wuYuFa1oIWGgjmQMMc6nw12Xnz
fo0j0tDNrg/SjZwN/ZMBGf7olgSVRIxW1GxuuTr2pSN3fpOZ0aGFK81C9v4ssoqO
x/gA0/ILD2JPa65TQ8khxsBayWdkxsMMeelDdzXNXWxQ4USODwJtVUOod+GAMrtI
bJdH/jDcJHJ43gy3ztF70rswyvP5mhfc67V65srSdQ9RRBsT/si7QDhO6PbX+aqZ
UINedfIv7OjvtPIrvU53sZTgzsxxQVzOAMuG9wsXU3vmlVwedCRk2eqn3vGn428p
gHWrQBg1OsYsJHUpu68l99JdnsZfetETWx4nX2H9vK9QilIOz8NMsfVrSRPhZPWy
Epn+SnCqL+NkGfhyFGvaEyE5InDBObtsY2qIqXABfNWVQGZSK8Afj22dhP2AmYm+
6zfiik83I/oyhVUpZMm8TAzPixqIq1pI5al9ZjJqmdcdUEfieu4hNdcNBxQ0RdoZ
zHhJvJVGPbPRY8IyYyEzJaAGzVdai1uB87v+01NAnt5UhvEYu8sWH6h1EYrtzUqd
j1OQ3IWh5V7vGgVh5hwduNgsGE0RwcIYaqK+23ideBNv0qM1B42p0HcJ4NZhbBFk
7qimNoxI0Lot6koo+lroMoaPhBjJRxeQK8Cv2OAqMiVTCQzkF1z1UQyJpBojhJy+
9Al0pSRo/0BmfP5EWtGW5Hilt3fp6qSZlTs648HmqQhUbL0qaXUeK7zdyzL3cPb1
4H2slKLpehOTOnMpQOnzo6BXnBGblHaZndaf8WXF3CaNeV8taWNLBaCwgjpoGN46
rDfhAjeUL9H69rwxOcne2IHCB8QF/9Pj+h/BoRL0VcIH3Ycwxgbrf5eE+/3Gmoll
aZrOa43Y2deutKm15J9ZGvZxQO2kyItGw7pLJbkpRttOwm2rCAv/NNaQKvnvZZ/v
dY/8et5R4qMjB128k44sLtw+i52B6Adq1RiTbu3CnqwnSjZqS01ZQkJv3+27KKSp
sP4gxbIGTNJMln4SdJyMi2aoMC3wSCyG4YtYKVqMO4vPjyWGRjt+DToRQEJwxhSV
Ava1aERQfpXWWTP/VKguALw75FMSCWzPEqWG+QaWIfD20wTW3e/jqK8lesxG9LUf
dMo+oCn4l4d7sFLLITW+8SUkAMHFGUGXw0SuP5TcchrULF4KbN0bwM1b3H1wRECW
xXnHyn+bnJwfjfhjlw1Xdkz/k22plDNF2+gnnhRVM0xWuH4/F4kOw3tPdVSLowpC
tgkyZ1pbBf5Ixo3F/DqOe7sz/oLmHaVH/vsoR3m9osuJKRTlP3uiZSQpo+3SYn4b
3YS2/HFg/vHOHcSWdjlzmQrlVCWFIciyedg0ejpDKPe+tkONCWd5B1H4z6B9z9OQ
QZBDkSikCMwRGlhsDnLrvKmBqpOXfR07erDCMRbR8mk6Rh2Rx6hlDnRExGyYlUDJ
w4xWsfqdXvAy4hLMPem1C0YnercIKJr6A9hGTodJGiNvbey1GumLsX/PgaAsjhUa
rX77hTIwlAzLHugYNApI2WQ+kb+b3yI0wKFrlLAcE7n1gs9tXn/hGlMJDNzbDPyu
WrD4ktNoo01sBrqE3ayJ7968ifZuYNGQwsHoRaV4KVhfBA5+r4JZUX0YYA5AIr9I
OkPb0XCAXMAYhqFfhpuGygOZMPqighN69bCSbKC1Y4cwjjIfdX4GQY2i6Vl9EN6h
bc+shdth8D+MPZbzwpYFFYX16FRH2/P7DGpIk3kH5Pk2aHXPiFRR4LM0BZe6mDzr
U2PcsCFoo/8xD6yZ4xR7q+7f3BFjzlreOQjCJVd1eM2sb1k4X0WhjKnR0nLQzLim
6LwOjWuf8pqEPCcJiAg4i2vvi+xlGXIeI9R9smz5wb4eThWaCQVWWaMobgFTOPBE
EHbEXbgscWAKcSfEzGK0fmrTrxEDc2mv541AiOZi/Kn2ztYNClIq+4DQ15iRt0ma
55eHjj0V8XfrCRQmUcqIbW3EtLnlg2zueh6Lm1YZaXIslqdVaah2uLbXFDNc6tAK
xhLYvvuSlFnIz04osmPyrETsMIhBlFkX5ERduUgefs+7D/DE5EA1yQH9EvGOuDn6
L0O+mREcFA/FzYhurfPhDDEHhiIKRum8LzILRpHTrepOAivYkG6psjoc2Pw7Fvfv
bmYTyjP3U5Yql222mHVtxm2PHoHnIaCFunaAAFYDk7V5dvbFzf3rGkxTzJHj8eCM
4rCY4t7H3K6sj8ZLlkUZ5xN8RIPIZ6eCNAmYM+TIaaXM7r7YUL8fGldDIrToceAj
p5DvNHFGe5PdKukBRiZkk+t85glccOQAVD6fntNF3gCMA4c220CxuX7YPD+fx8eZ
R0anGncgsUajvsZ533yPlT5q5/V/RWYDwTAUKA5Hf7jLio7Igr/TNQurFy5t8DT1
PLcMakBwYToHYtwVZg6F39YWqIhWIoJM63qtS5hbKYGatl+bjBYeyzSgCCVIdTm6
ie/4S03MT13JINsQFWIzI87rDOPkGRb8MF2cepukLnCN0kC2t1JjkaYG7C2oq9ug
2xLbwV3ISMrexHvnMcZyX46ybprH4HYRaiOzCNGQQA0i2iqiKpfRhlG2tLEuG/r1
PzLPI4YQACw+Zqf89m3TrYFzEjTo51m5BVL+z2aWCQHZqu2IQp7ZIKg0f3GIXDUB
OzyFkU7WhJK7zI30byyHStKOsK2nU5rZG8sOlLKkm50JODXaVyFliq9XYA92xcD6
E56JfsW3Al2pdc0mxeoVA96Fw9PYM1cVfrALa1ETYPAI/4bbT1vu0P9lVnjVr+vu
WSl06JAMXGTMPZVR25axeWNfwMFPwra8iJW5jgoS/fgKhfHFVfnZIMjTXH0QAK3e
RwqFA4SRGGWi3P17IpeyBlB/p+vdT974AM8AgkgjyGgcm3ZzOO8FkKm4H7Aqt50J
KEFahrGylOwyK1eOZQlrQNOceHRxLydsbGPQTrhsFcWHR8oIfU+ZmbXLBcNfyagT
BsQg6UMAkjM4CFaZEKtbiSw5vCDUN7TfWLbxZ25Uo9av/3LmYImJiprTjaDsduSf
7NCcXHWYNnF7WJCoKKo0b0QQhYri1e0KqB864EhjRZ2Wmdl72ZdGONpMT3Dah3Zk
wfrz+/6ThtaB0g2gAqSO8dSxUu7WZVrMZjQYzaJhbWZmhQ4+SgZnO2KqgMLDrYXN
gxxMkdYjtjHWu4tpMYLNU+3FOD0WXc/L0I1rfkCgz6g7pO/MTq30uptoUYgHueYZ
RH70+ilrubmxLUP+0zjHik/qiazGlApfHzCMRAfqmLzHH+4vqyfi25e+FVS1P2Bk
92XnV8BCijCn4ZFycwepwtg168P7cuKd8QYUzS5tAiJyfy2AHzA9MYvenotttfM0
yJVRFsMGi2n8bbzZQx4TozkJAazpbswdQCVB4DOl+WfsEHx3vnG66daSr3H/6ubB
ynL2j3/PerBSNya6zw3vpbj0i541KLjH8e4iEmCr4K9O1eJa9JkRjDEzYshpKWUA
lJKj+Mcr5mQamDa2gBMIZhwfTwFA9fDIQiPn5sdsvMLYFwEP6oKtdKetSuYT0pND
x8wNTyqVmg+Mz6G+jv+rPpFTdwqPXREvtt/ukC5bJvujhBc+hc5bXoQ/DBl8qbDC
L5wqMNaeKwfTPp1hhAtW6iKXK9roW2AwkFGf9SDkchprPYYVhcBCgrwuaLdQaYI8
cmdwwYvEv2Knq+KSoCo4O1+UJ2IilwNQ2MJ7u1uKDw2ZpLQ581qCzrlQOPzrzUhP
7JQS2mlZ34iC8oxyvarpUmlTlvgNWTC5gJa8PObirAqknNKZW0pR88Jyo2eJpfCn
nYhbuKl6xTu+H0nJ0J01/iozfIPu4wM2Pv5sRUVf6Hdqo9TV1aqAmI1N/JI4aXsQ
myeepVbH8nSfzF76fPYpKZgwrH1uf9haO8801hPZaDcr9K/9VdrhQ+Mmz5mXORi8
PlqvQmqQtZCT8KKEwIw5D6yg5fWKb5EZS+BAyXGKBkkbiW97I8q547V3m+ubDjur
dY82bolnQG/VsnPzrX4rVYQ15wfRwjN5rSEVNd2Z9o0i5eciaIvcrfJTFkRrq16o
zkHQvChf4RuCwmyaI25Al7ByAN2whwL01sgO+IC7VMZhU+4oTkiEKJHSEvtY14rS
0JftxQiV6llYKvAFC1SJHLLh5d7OeSyo+H787mfTRIIuZsJm1xJm+H3KsnStcnNF
/3bxru7z2/5W2R2cReiAslxgS2ovcsahWnERjTbaFAxbaw6JIcH8mx0OCcxJjbCZ
GcDLvOY1DpyKszDH7odYwTZsIbmZJrskcktlZeMXUx/lkFS5kDPqBb7j8xkWektG
d6OA+Vs3ZWEzHlZvOd5eHCQBmvqPzx8ddSV77Rv0EMY3il87Em8UuVtZiN0u+DXq
HK8iau8N6+yvQ7TvrFjU/j2CPrJw3g/8W0u6nF7njmfBWMC/zTyyU/4ntU2jtTc3
d0rYXRNtTNgIsmzlbBtSXcDWYSPkQ/6ifrTq+K90wB4/yuT744vTyF0Tq7oBrP/8
3ifx7PUjfEtvdrzLA1a1DXAAtBryiiwDwaFO0RN10lAOXuCXsULYm7P9L1rkXDnn
RPYWZV4eu3V9Is4/hXi0EhsBqEkBY0z8fNXMScI5owvA3N2iEMqj5aX/1PrSjUnw
tKRfjUsDjopq8v35OjfYL3+fBACVSCwAdJEA7OQH9NZ9Egmoqj/nHozbj0cl5Fck
PgzrocDNBcOWMYiQRIpPGRFHvwZMIYUq81lMV4QmyEiEfjRcpF0KN66pWFTFaKKj
YbkJjceoVnFaJ72HVYeF2WWlxmfDwWkLaxB9RX1yFDj27YRkfu54hTiSfCOJMukM
lopsj6wOJyUhPPWLsaX9Q0PyJgd6QbW9pb8MOdmJYnn45xUTjoYjNWrIl7KNokjd
WlNadXYq+LjETFnOg5l3AOxxvXUvgkpK03LGUcXzSXK7hJEKr5PnfHFRIf4EundY
op8VmKRkkIBXNWIbOQtLlbByCd9V63PpNb7pZ3xf/s2n1241KT0joqzklX6Ln0OX
SoOTXYrO3pzaNFDlWs9Hi45e+eNn0J6uwx/r6+xr1z4vp7A/i9/M45lYSNOdsbID
ABTrqEEBbXMiSOACe5wWzgep87OUmmCGtPMsGNlHsqpOpPhz2TSPwYbeU7gsGpQX
oInbaMrd/MMOxi4IpIbQnUzAROTQpmiXuwIY8DrFm4LPbZqTHymXZ05zyykPXAgr
Jtx452zNvQY2QuMlLM0zjDhW6LUdjmooxvMzR5ooY7g8vxiqKreOy/bR7MjWHZFF
ZqColjJNojuIJwAHtA0gTbZwr7WlOUbwX/bDotpu9+5LNY1iH602tuPgbVJJ5Y+U
+T40kioLMTUYNZsVFgmNfVL+3aAPFGkabVf+i8ADSPO4IbR8c2C1Se3LZgRWjTN0
jUWNpmH+DmPD9KxTjr7Cllw5CoDAnPFFM4gWI0kyXIWkDAYlcu/Rp8KeA7om0I/q
47Lpq7Bb7cQW9J7sC5F9q0qO9aZ5atHAZT0pcA3u8KpXNz5fcBB+idNQ9NoYYYr7
aKQb4Wrz9XBvNa1NGpxH3omefYkuzw151e0Xs6OEa3mjRuOaXSc+ymM3JPnxdOKd
Pmmztjm7YOYPthFwiJDbb6V2SzOAqQIFWIAOBqosYMumi684nONwNvJcXL9eVc/v
uXgFDh1xwcvG9b3XnSNm895MUWXbq1DiIYhCAXWvNNEvkArU0EQcqZs4Yfu7YEdN
OLNturflf0LiQ8uzIuB1ABNSZc2ka/fEK+apQ2YvxrdjhG7vIflx/PN+h0RhQE2g
I0jTkm7SahUveAYiyHFhtTYDkRPQQkfcSeBPv1tR/+TZNc80InVaHyK9jm3k7HGU
U/cStldhSBqZBen1o6CzwAWpleigoElgFKoswVN+gbquCfcWK6SBO/OYU6+3nM3F
Nrdyy04lFsEyJjfrZcG+xui3Q29+e3zk1vxO2xJbgaT+Z0+wOSeCegibN6cQp9Du
oGZxjpV4/90bhsPERMz1Ui4eqHKYoEt/FuvdiXbPCqoC8ePtdOS11ggXuOWilvH2
KjqamAEBejYySpm0XCT8THrH8HgkvUGOzHeSYfpd+Wmzb7dXDb1U2prBRjNFfHR2
dscdeg9VQIGhCAyQGw+Nq8vqinI/q91OuEoNIrWfjLnSlvB4g3+uYmoIjTiUFQ2I
IdSIYbB+S1GElXvmZp7kDPzE3RhjA16RTypblTOKMKU+zetBd5ND1ffDY1EQlsSf
gm/XAKeahvmzmLsrOkdlQYbbtREeLym+RnlW9RlVrOFvDsgZ85R/ccawIb8GFi3z
ZvvSaSI52KzBrdyWSvssVIc8j7o3sopvcg0Jmd73rIgRPiIRz3koDbWkgiZqQivP
q5LRa+KhCvog14THrymL9gIHBUGldlcoa6uTyF+reYyxlL50wGKCrd4V0InD3wBD
t37BXGT3IxMMS2XDxhayL0+QrkafJZwbGfqYd+PvEfZtXGjRZ9JhlnSbfaMT4tuH
8AAYI9m1Zx8l9wGSFhyCiHslwqfkWo3sdN+qmFfMVf8=
`protect END_PROTECTED
