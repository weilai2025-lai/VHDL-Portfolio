`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P30o8/NWJWZt9l47XGQicn4Buc7UWyMvu9tuXjLeC/AOBWJXvLU34Xfgu7HKpkhJ
P6Ari5FSSKHM6Kir4j6xhSPPH0svNnq2Ud/21rouVDSeijf4JsvQTtUKREGOMfMD
kOLsyFP9749A1zXK2JyuWJMq4pzhLADivSU68xSQSeWxd1EcHx6QtiUt/petzsAn
8hsy6AuXBWH9xuQ181ZpzNU5lgJ6p9BUV936fg6ope5GtLm4R7rwLJew8TTnXv3z
oJyw+g9rdlMPAwqJuOfNPNit9Ju/kVewqkqfApDNwuGvL4LpSSQPoGZ2cOVB98CP
tOxVCIe7htd5Da01WL9gGlss0P3AaMR5vU68Z56BvILp5iYZ+TOJgWtpQ9DOkxSy
jCgci0/ecElP5u1vK2GEKlVj/QFwXSImUmzhgEBr7vj+x6Xb29FBoIrwtW0C2ZV5
Hdp1fHW6dvL+CWBjCUW6aO4RopnjkirCA8CSJfrsIxvx0Y1XKWZwXoFns4CELEkU
Dpmu44dUmD4t33uum43SEfitTvs2i0yYyGtm5lxLCecy8xC1Bx/SFW9sgc9me3J5
sR0a/y1liXtR2GpunrlcPjdEku1Cx6/vF6bCwNcIasxFJqq5PqMsa2c7e7ThhZhZ
cU23RnJGJmtKcTDO5HAnviwKx69WHy2kzQMW+YxwyjoLybNXzPCtFLh4v51ZWjFY
T1T4rXzCDCB45VH35HX6sErIHDJ+Wr2Lm16vanNldnYSWCs3pNODG61vZuXATlnU
13xKTm2wFwsr8ZZvrb9IZzDFQGUtqkvM03HaVJa7D6kRDMLVaeXNB6NAVLRG4nuv
xHXCuhF6pgOpciIibtrMVFIHX+xwBv85jb3IiZRvyW1O1n3PrxcWYGAkl/hZer6x
Ddx9wgODEaBoamgL/umJ5mDDFs8LgHGPnDfPuD2dAj45BYanI14r4MkHP75KguBi
TPMp/F9m9M5rcFFZd7o4KmDfzGVfzQ4VotX/bzArTXGW9/lispCZuOb64SP34QBy
f0h078Gm8MfuWwf+kbGPDB/n6AjQB9RfEbqEseTPiaEy0OfJsvqMG7ZFjER/YuhV
aHwoM+K628xgNzjNIO3WL/RV4fZefrIDdIokeE/HjxG5gh5Tv6Fx+vNVes2Wy5Ah
lx23nWnZZmlmYFyUQ5+suR+vZo2zN0jyMDJQ+Cl5uLDiakZV6EzL3bHbtSwVxYiq
MQkRAv8L/ha6vYO0osrmKGJRWGtPnwFLWUHhhbO772gAfCGmhoSp9uA3lfmlc74v
iCCxHSVO3HggPWd0y5+p3HLHvzD9fWmOxXZQYUtXx7a0YX3KcLNUfwqHlqeshd3f
v+Nhxc09KwZYEgEedfSKcjNPyw9utFDJhyLICKRtmUi5LX0QGT4wQh5Bvv0VE3LD
cX0FX1KC64f+6lQBJ0Fw0/f+INLMfRJtB/olZ9bypIy+egPYPUWF7N8mN2tq/w8O
ZKATpgMkAzpHPX3iV70Io5O9tXInoOlg/qGUVO4wCKcGYffUet2B5F46PYRD3+f+
G/CVsgXEXqg2XGIiC+3ajXN77i+awA04B+84GgY5H1Xg52kdvq+j62peHZ1mGfuh
rcCZH7yT0tMEVEF4zhhP+06z5ZIZnXakku4HD0mL4+k=
`protect END_PROTECTED
