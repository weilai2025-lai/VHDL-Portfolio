`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egrwR8ZGxnEUtdIXLukxX8aPMcEZqUTnMyacEgnC5rBFL+5r3ujRYgy3OmOfNyCC
ev4DJCyQNT9umuzk/NNNM0N63P//qNDuiBumnk0nPgKa8bXbSuFZPv/EdQAou6ao
eotpib4TvDTSNume+LHmaKdkfoKMxx0Tjcf9Onq8qYE8QnuzcChZwjUEvuLUJrKo
j//YZJIblYpY3frRC2a9hKc9xdOVRxJ6MzKZkt/t2mtYDPw7nkBOmQOUpehGRVlz
FG3GUPiQMICsJhJHx2ZoO/L3pF+T/YrNPExmc2RuNjMRR5vmoQD81xbkfLeKGt0U
Dk8tmf4G50zHAF//W9gm+iQHikBn6lrLYgnS3hh2lkBl7TgOrvS4S0iMX/VEkdH0
Yf3HTy1a9YQsC7w77SIG88aoqZkDSjPuUGUNGWvhkbWWfUcueFsON/H5Kc/IpNKY
8gPV8uAJVRdH+pUwvWRpwv+yIFd+P4kaG4tovEnl2bC8eisSPQMTG8ywotZnD+6S
uDKjOWVMmYL6RatF61IQd9FxUi5DVKbHEGSyUQws5s0a54XOpUHt0wha8/DZjg3W
uS+2T4dGwbnxCY6CrB2eedtEBCBNLuJidFECPq/YucWVrthyF//kaUx86JIrzyW4
5fjJ4d6XZFygHhfyC0RVWhhtAY5PSerB0h58rp9LJDou/NxXG3pRmPl65M+q4dFT
B2/VwhrF3zKTfMm5ukKjQK+sZ53KWDvyy5Gjw9xCwwRL2L53nSARBR3BeEx0biIZ
1RTdLWmmzbxLmN8T0Hphs4aTJ7UrZ5flH1b86OR8r65xpP0X6pxv/IpPOKfhm6e2
XWS6FlYuntaZDPUV1Ef9J++44AM6+0DvBz4v4NyNMIJfNHOT3JdsWdneV/zT3Nz7
cxQ5a3Xt+B2leyLAEJwUQlACT0cRcCRFGKt6SltjLEEDTMWfsj9N7Nox72cM4rF+
r7UJaLWCaAUh6jyNriZHTSDEnjC6pciB3rmPrkyCXMa6b837mEDddB0g1Bt3piAl
d75erChY9940z1lQvqUiuU1b0xz6f02XvHWolzbXpPtcQ2elR0LHCpZkAe7HXAvh
MSjVG/j/yrqYTIp6F8bUr/5HMnHgwBSiZtq/TRVqdRAURu+Z6Fk3TfHBz5GG9BVn
ap+oljKePkHCjkLDO0/ezBcX9/r378ZydUTMQ4502T651un/uaFZTKItBB7EQ6Ij
oH3bXwlXvXH0IB22zlUMG1mVK5mRUGYnjez29nl6KhjH107UXHsw/2oCzxE3ma3o
fqK7affJtvGbmS2WezsbAFa9jW/m8e3MN+6b0cKllIrFefPadgEFRg0Z1BIcBH+K
23q0kf2FhaQtddsfT3BYVSaBIoURqISO+fz13s4+egGHbMQck8iVGvuoWPTyuRcp
woR5J9fO9y1WVxlWStcmb8+ZSMVcaw5HLhMfyJiB7Lzk6eYq7bHkBpiPXBoa7o48
sBI5+MOL5vIMLNR7d6+VNUOeesPn8G/LmHvuYkcF5AwQlQf4zEwLmQczEVGB8tIW
gukhfDGC3Fr6VxNlq+5i1dNcJgGSFSaT8sOpo0Zno0Wvbq2M5aAtvlBcxJ/BVFdF
O11NHzLbrRvr2JEBategCirQk9s2i564VDTgO78aX0IgrH6f4C6RNMGWyFPylSQ6
b86K6TC7erwdY7E0y+VGoCt7UUBIiJ9PGNVDrm6sJ4Cby9WbPFvlGvjb7ODd3MzS
jp60R3Gn5lRUaL7MGB+BYV8aozsW5Spk+CmHqybTFIMYLbJrtuHMxRPR1egYJI2L
HTj00QmvPvCOfWUFfQHXxDPtWYsn9UU7t+K/LTQfoU1MD3Y08f376yjMLPGkLQMb
WgkPjWm4RC3px0/7JpQLu4Mx8o7bkBv3cY4seoWONBIi2uVMjbBzsBT16TRX8r2U
dJxJsVejCPl90ZPD6dcTEbcbrxhvOCn9edMck8aAJMgnY5Ve0bSpHn9Iz5OXzeFg
FNjrwNI7zzL5FStJsk/6C4LhcAQu6OJYq9of4kL6sC3mxHOhxWBf97t0ftXUFGsj
tGULRgzOrGsooOpZwhLTKVsQJJQtE2EhWgA70L4yAAIoFnwH2mhQJZ7hz2XHbVpv
AvwsjU02j58C58jtY5CuKiNMQb0SdXugpo7eF0sSkNnn6OLtUe5P7+DPncUQYhTf
c+JEEpTVl8zBL2n2I3dZCkFDJfddq2bLOgvXHX2VonDjqskL4l6SzM5BYVZzg4I+
7tWRRusf8beacl5q/7bd19M/q5J7nHC9Jv0lFHMhtdGjMNj9o6mj9s6io3Q2Unl9
phcu19NobaUGjlCI+ksRu1OFpgjo7cH9VwqtNjDednfphwC+FsNMoU9qAwnf8b5F
I+u+eDTbS9iXx10yUGYKhopRIGwR4d3U9QKytw6onh06kIuzujRGjdgIqP1kCS5b
zBGv92t5jiZHph13RXKqwkpJJXQjN2U8e1xhyXKanaNOmjxK8o1Efpa230zjwhDc
pmAm6yduZYtMv6K5Wh6CiicBt9wqjH66yCJ4InuIlYxUoOB7/RmOyxDTspen9kxH
XCEPnThAvcfIJPEGieePBPr6ik2x3K/ZRfQCjWzPZbqkDhFTgb7/Ty3GAxn0hF1L
YuP4xHgnCEoiL57Tep83l9MC8d3MtWPZvFxZc5dewPJYn6VOUx8tqVBYXZTGrgIA
GVj18MmglrXMyLl83ZAB8PkMAZmfi2effZacyzxrRiIeYSU6aAkd9tsAYuOhql/7
YwKjuyUl6Q/B9c1TbxxdavdXalA1SefETrBa26cWyTLkv4ibYrt7p76p+AYdNlV8
FVDCuySbb1jgJsIeiOX3EJzyzLNWjnNuqHSgrm9aVPaQFmpu4O34LOpNAf2eUuAX
Gopsw6lkF8FLvA9EqtxPrIp02fbiE2UJtvHh6FS91XFTDvrmIsdfqOE6YqDslFez
1WNvBL3z05GYrQg43xqLUjMnCYoXPe8HUdFY1X98sALVfwMfnVfPWwLp2/01GutQ
I9vvLMABMQcvHFwDn+0GEqDMVRp3VDXDQfuOQg5aQh5MlB4nMRPBIVTzkSZd+tEJ
LAUMy4cehSdKydPj+jpDLiccMXDaQanZxCmPgq9ZP8NFcRKkbsr3oUOgcHE6CCvJ
+5uXjR8Bc1acHpiNhH8krSt6gc3PdbjZqFyrQdiFonN3oD6LewrvpvzcMzHgwLwx
8nBSlSgWc25z0K1/M2CsZbC2j3ZQzFXZ1jhbH7nb4WnyIDyUj+zRq6DSmu/kE6al
JnX22Xeh1SHQn6fgYfUHSgW3RAHfVcHzVluVndldOYl/pJ7R7NifgM9aEf0/ZXvz
LRvqgDU9a3APWcU7Rf3VidN4oTDmP65t2ac8duhQJQ165YqJU3eOdPJ/Kv22vtt9
6Uc8hwXqxn6kXikdAYgSiGHHfy13jYnkNFAWj7GF4x+vrSr48owLyRrSqIi9+M7u
f648mEtoy1JzdC1Qs3F3u0XP9lKEma3VNPBgEdY3oG7TbDDSlzy+0XdetdAYLGXA
Sp3EJBQjqLDUEYZ0GhyVizAEefdqaMNafXySEEsx5YkG+q9m8u3tGsPtQFKRIMRS
HDjHfNScuT54rhLfVRbiWbqAYzkCUBcEMTQeg0UkXxeDsVqEeYfh/yOQzTFB4YgK
SYkNDjmSfQHGVrQcUYXHSLRuaJIWs+QOdAGf67Zn6sja1uk37o+BTNelITvNnBKy
hWrwB/VlMRcc7W2qwCfRmmnaldXAD5MDBK+nCDhs3JmdOg0WeyBK9tNwSBu8Khtw
ftODHIhGRQniLbZahRDpVTPM875QmKX3dgMOpulY87K6l+Kej4JWSwilXPQviJky
pSrqs87ISM2RcAvrtvSS/unxj+Y0K2SMGnnT0pRsKKZk3DY79QqCctGy7qcX5hGc
2vFxQIKJLDHRxurhDIx5oTghOtrv9/7xOROJJHmROoiDCQIzC6QeTwRnbuyErIav
vpWI6Htzvbs0radXwKBLI2bw2O8fmAaO2WzceRdwE3I/TjBWP05W1J/Xsjv+ZuKZ
w0JkUHl2se3tBDrxpoK/Dwrga0XoBfv7pEAcEH2fPJ0o7T7x3lsVrMEYmBpDA6Pm
rk5u/uFN1ZQMSeF5kCtVrdJuKU+WUGqxSxV+yThpN9AtFW/5lEP7Zlfj9Tl4LZGl
IxpPbWcp78ubz2C2rAeBCwqlh0C9z+LpYc4CuTakCAOhhzH+xojUlmZP32BJYKVz
KD9+JZCUsThcFOwKFxGUrZb4RcYsN3WPORRA2i8s+LZQpTholDMnIZL7OKh0pUSB
YH3dw28zuqPh5k5AoPPUbCByAIbME1qNN/BaMC16GgDhFK4YIamcInsZZkijr3P0
ywMztgybJ3G9xkkyV5v5TLAsE15QPoo+m9SxT8eZWkgnzZGLoz8PTIW2jJb224om
aHYpk7CXqEEB/3enGnX+7qtGPPzniFkkTJXFOId7Fr+ZcyvvviO6V+CksqfCJXXM
vRWYt9bt+3dqPkgdT5D1xVhZLKO3+3achSIT4YBhnVl//zIuNz0OXmzIW/y29E8n
N5oFExhMGTm+Av79l6uayEYqpv4gKhEREXTOm/wMNyyANSqP8y+h63yc8SU4QVqN
Le+KFaQVu+ozEy6Cw0i7U3wgbdE9VUY3TMTZ6RRgUYE94NshDifOUeY7+FRIq6ya
D9JyTXiWglPTVyLCJXvkHf8FlGcAf/Pm/z0AXdlXe8gRyXq33QwcQtXVP4Utl8IH
bHzPevcXOunHWh6DdRIuj1Aqo7qT/KpojwH+Aqd+fC+aLJqw7e8rSJlzijPb3fXc
jRvAo3SE1NuwTYQfTcv9qIfqLYI3j+yxJYVvvVDaNSmrZG+PN8tbwUJLTTfcZHGo
Xunby9wooloFdYMW2aR1Hu5XUDNtlV+EBLTgDhfwdhWn8t/epraAL/hhJlTwW6dN
1hONphHg74girgXgKzLvzvg2WluJ3IDysBJHE1s+jSUhfyRqX7qbwYq5wMMHGIPb
lUUiWRKj/Pl1qvfNEw04zidmFo8UILO0OeooR6TmzelLwn7ZIg63s3JmNQEhbYqI
65aEe8GJW9mG2RM0AsZIiZSwEMjtukQ3FfMnItP8I+RKtZoRXyOrkXdcKRuuLTJF
D8QgBaUlljRnf+V5ekVp4EcIadZER6wSKysA/uEARGT5uHlM+CQa/0VU8pezq++3
M30PCtoZI9cqFxzH6cH7vzbzNRM2IynyMaMBH1OhsiGjkNSdEcvicgNUCMAIHjF6
gouv1usbIZwI/QSPLHgDr3kDtqjdcTbBpXT3vRzD+Ob6rV+VTfNCiPFcu2I8iRIt
cHT5QxLJ05kIHlRt5aBkJ2gdWEtLdd/Ap5Ay+4bOrWZodFPLRr9gxNkMuh4ZAHEI
FbolPSoK1FCiJDUjLbm++WreAg251DLiXc4lcKwYswD7ZBvoya7z0eRNuALE7tdQ
gZ9rrQTaT7bIcvJRo5tnlx1m44OqzrwaHlEGOhU8dGqEHUuyvbkkV+k4IqNAiZJQ
UVfYmq2zzbG7F4gUzYCmJv2LLi8oyBPl68QEYZsNUlSyQrv+k/LQ5nz1+gE+bjS0
YREsZlPZRacJ0aTRSWHZjPB/IUHfA/7WA8KhHxQIQeJ8SvTqRWutvaWtElluX92d
spBnWYx1wnLgv1AFJCbNgw==
`protect END_PROTECTED
