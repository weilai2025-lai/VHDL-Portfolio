`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KiMXnXHI5vxyI5qMRhLy4WapGtEGQfGKw5E/UaUEBMW80nArmjTzHumGa3pCntvd
3Ee9tLNYYyqkt62joIGa8OdFKx+gwMl8z7zhdtxZdfnevMzE62ijEpBhr7TKIFJX
HRiupJ6ufHkQkVPh21a6OJ6MvWSaKk2kl5k+LbOXPiGyRdoCi9Gt+MJs04lLRlzB
cKqj6w338X8XFbXoNHCZRNrh0xM+CQKqYgrBjJhCJ9spWkhdO+q5F1r8cLCKxKWT
w1k+FCc0NCnHRgVf4mL6S3IPW4n2ih8sNalu1uXX9F63MlZCfmEf09I0BfQVxu3M
o8AMypDbgMsPVhpR0Yn0m0ljyDwWtC+qdLMewwh5eQl+51Lx6xeDpkFBNlfo8PQe
W9t0k+sEQwqdhbyDV7O/YHfRFI11QkNzdJA56hh1VSEFSURFYV0yZlH0VxiIGM7U
azKbrfj5kc0wqUeOP8FDQYyd+zDrRgTzPCoghn7kSkYuGoVsPZtNKe9B9T3F3KT9
BV7dIGIGY/UTnsgZ2vPpwuJ5s24+CmcTVoa7ZqVKQWOM7m0y0IrMJyO0vvxe3fPH
XlNunyCnV8f3DaSNlS2giAWXYkb044heXmSBmhjYyY/oludZhRV+7qChSBH+cI/q
HvUbngq7iOdOPd7ATjfOs/+WSug4l4oASpBx8MVbpvSVrklVXpmeUdBsAaBnLIg3
Zw176/4Wz3xVdEB/aojSZ4/iWrXizT3/38pv3YzZ+7izi2JeRgBzSmoyt4RzN/hn
gSmJvERAyvpdybrU062dQjXoytx9P135oeGUwKYNXqhS2KWPQfaQIRFngUyRMiRZ
OINz9mC/t39H7lnKi0/SIr1JRnO0xqA0nk57vXCASX3oS305ovcLhvXX2UaE/5XI
mZauN3Wu5c+cfPzjpFXB2rScP1cniBGpFA3/mmCKHkwUZQwZzkr8FLNehlsuKGBy
IAaGSA4yqXlJhgxxdBHb31FhySIWmTqsaO3JhJZAby0rJ10uOT9bs2j0+hjAwGV9
+2EaMKppfMLOlRtyofUUndGyLCTfNjHXGGaFCGI/4QcbaazwC0UVXRKhNGds/e2b
T24fMLm4cJwnOkax6kg4f+GYeJZ838pKKtMhLL73mMY4V57f2g2gxP09RFPMfue+
xT0WArIZRQ33TUFR/wRxmtL949xMkZsZv4/KU+KDDzQbb4Ggm+HA8Lewm3oF+wB8
oL0vT1ixW8B38WXFwKvQ+ezBlbuXjzAzAqRCTaWp3jBfRpcla7YuLYLwejWjYRJ0
hBAHOcDRm9228F5NTZAUxdTZRKnwl1RhF16ksyS1r4Lw4XP12VVKDePonK0zSctf
aNCEOSYHDGuaQZfnjqHK5UIJwa/pnhC3qSgig7JpqtBJdjc9afCMJyGYlkOclPGz
UcdHe6TuyU9buLZYWKqqL96bx/jDA+PJlJ+mNNkbU3lKthEBc7LkHrzapWn5cQM8
ZDNv85+pDv/xZ9Yj0g4Q0mzqHzGDkMTvzCu50Yq0gPkDA68WmR9PL0ymow5sHvlm
qBQwCGUmXl67BweVpdLWldDYc2/IEpAVvdAIvZRr4NR3ZcOZ7XoB/YuzhYaBIlub
cixKmAAZDj2I5JIQFLMvSKIA8yhKd/1mEKovuaaaeSqG5+BwSq4Ks6x0nV8iwKAJ
bOjtZgORr0HTAUpGrjqiUGk4j27Cja+fUngN2eGDNciqO/Eiqi9QID5SKSKdX5iK
KmferFF9P3994nAbuiH83eiOwDrKJGKOmZJGXoQOQDnpEjL83arzxHqnj/E9j5VQ
Y2+AE+RhSXjVlEJRKLnSOer+jNRdiyV5L/a2puO3myW5DiUCR1UacSlViTA2V514
G38d+hKG5bccpTQqljyJ9fcZZ9zuLK5kgoouVgk3W91U2JAxbd2Kr8jnWV6hFhZ8
Y3z/BrjPURf6Yf+xx42WV+iXFxWkejDEeO6+hkrRIeXG+cP2qYC2rFTO2U4suiyH
E3Jnet+9W07ka381OZLzQRuBuXxuFcMeehVmgEaEK/oLUfpyU8tcyZkXuF39oVNp
Jy3YTeo4Ebqjz/B/zs9uV6Td1OZYlv1ifs8Y8gEBZ0M+vZ3AXVhfpC8JrQ47fHTI
WzrO2A+U1MSFHb8Gi71NQejUW1jqhapjJmjAWo6W/uMnINiEWpTHR2s2wp+YZuLl
nJD3B52w9Ny6nPQ9QfcREBTiDZRBB0XsZlZXfYFr/njy7pzVhsMTHZXDxPKCrMDb
2IlOb/6TrljO2wn8gpRFlzbcTqe9rUK5/MTe7y5zyjCrVrBhrUsjf9PldYViLTFE
jXBscOvXEGbsPZqtDC+8Bpq/6Mh12c+9TDk6lpT0ra0P8zF2unDFo7dR5jUxfu4H
UMs8eqe2NfKSP9DEOESL05oXng5ABocYYznU4oPIHIqataBudj16wD/MJR8dpgBu
Wqch1rZUiRaYHD/DJUCErIqhywGxd0vL8OHaybISdAgp6xtnWM/tamGR0mVconLU
9W4mYpoet0Ztgj9lJyKisbOqrEACFo37pCM9Wg/jOX4JwkZn4TA8GeYpZvgQ3p3O
yIlBCA/p0kq5rIFWVf/XjydnLhpNWHtByESLF4eYqFTHWSXAaxJm34q01ok9tAKz
ky3gRt5s9ITpsyyOci/lJw9/2Q2lO8AcN6Ez/VYcn6CZgyKRJ1LJCU9PjI6P9CeW
BonLYiQmMYyB4Ue0QMCKHtejNfwlV0dQlwskzfPUkcmm8F+kVsLn51UZM6KwMfa0
P1vmNiAkOSt5yb8iQB2JdOh1eGRXOXo5YXIaKof8s6tysklrX1EolivJmpl3Ynr6
UKR5tivISFQ+xWbJqg3Xe/Q9YigDMGnEianPgFcPNTrMapvsOcJ7Pam4zo2ekC5Q
Si5/nWboHHpYfylPnkhEcHIWGY9HCCXXBEjo4xHlE5CH78PMVTBcw3pusE1XVUYA
OA7TXQj7YqQhi/0d9Vzqi7Q0Obu1o5eZh98a3C0FkbuhkdM+rPwIBBoIVHK8lFuG
vwl+oDELltDCQU6QrbP7KZizDc0hCS+clMGsueHy9JJFqo/594XYsP2lkfnLcbFV
t6HjdudzZ6K1mGLA5zYGOzmzl10o4e//ZCUvzGJ+F3vg9xoktiT34lHIvy8DU+H4
TdFrfOXQISc2wtrW1+GKch7tYuONcqczti2lt37Z4KMrEd9OmTuUTNBd393ViSY0
ZXyNsLhDceQLDfXVAPlZLA2bSHaAmTUn0M5T+qZxgvx5vPUbPhycSios8zZS09Uh
qJQAJNS14ePSAXc1yY1qlxZ3Kiy2BDuvbjF2kcFzkvBMOuBTO6OjzAwLcpymPeig
y49um6u+xaDzcWYE2sKirGHkLDV+Q+Bh3fKJLlbh/WFSvo4zq148PgymtwABluX1
0b04uKVwHHFwd6WKk7QqcwnJNOM5omENTgt0lWX886fS68grT46iVMfg6XzkzFeW
RoO0X1rI9nxlnCb74UvUYRu0A3YdQdSRxYK3zSTZErdwW4CGOy/zUWVwc9HLHgPf
OwNHBQ067h18uV/5diPL4hief5m/XkXDj0uejfi03I7l+xrpr2DDiWqioCbmWaKw
6UiBeWxe0d6Hdg8ddGMrkfsb4E302eJStx8dMsogsiRIp7iSIOG0PZLHJRSiV8ze
bM0DSrPkGvLRvrVGnbUXjhY4trV1fjFZDkcui3MxSN4S9uKYHo1Gb/BrEGa71gY0
yTBR+Sx/AB1aJHxDsUt5mcfT6PS2Xfa28ju0psIloonbTBCJIWCpXOp42p+bvvVd
5H5Qyvy1voIqWC6qYeJTev/BRA9ySSTiF20nuJ5BnhuypLVLrySZ0ENz9etqcQGe
AHeLpey1lx4mWbAVzmhkQvWHDJGQWNPYc4NlpptWHV/mUYxk8qCA2uiUeoDURYy+
0S7jX8KDWr8lpPX3DmwHc/6z06cAKl8KrjDX2YxRYhj/ac7bgj9hzONBiKxWX6DG
SoAzXg/HOsdoArNv8Ar13GpRApJQlJBxg8XusrJdkZffOw7GWSuHeP7hDlSsdCG/
iwXEuJhP8FNMP89v6PkaMFso/YvcqUqfaLcDP/Vqrx+O7N3wjSzpP6FeKjMt0gF7
9Y/ttsoHPH2BIA6kXTWwvKTdylNeuEH8UrFpMWvY/+TP7Zh/77x9mo4jC80A1qYK
iXyZdVvSymmw2KmCYmDFQQPtkaSLc+upz9eywa0KQe2WqnxP93c8BNXu720zPI9Q
hIhT/iVRCZeaO6HtjMfzDrXfSGiV2tIGPUaJsFmNYWFe9TL1r5YjIeW2iIaYDXXF
WzFlDOIISR1+PbpVudeC1qLpKvNesphQtDHaN9ZnqQPAGmAlZCAZJLEYRR+pJggB
+S+tgExv8DfscF3wkmBn6eQwLmk4dcJnRdsBLZ0Kd7rR1YjQhg7xTu37/cSGoNsN
/gPMIhYQXRRGUinXGqCBB7UdVpCqH/8gDIV8bmLHWVi2KKkygYhxDB3oXr+QLGRY
gVK5nCHEkqArT8NlW+ehMxxYTlwd9hX7+olAyKGrgWuIvGePq9tQMfVl1KNE5PPF
smk3NAhjLKRlNGlvf0QAVzyvJDmOKLDycTppxGb4RGxWd0il2RwJChQqSi2QZ2f1
+gVT0KYK+Qp34/MZdr6IqAzYfA+2BkODbA1+WOY8lcqPl14cHHvOSOqt2iwtV/Y6
5laY8I1Ws6q09O7atpjIZuzwlhHS0Ve1UbEp4KWqrWrBqltbCB8CUeLzyLFLfjVV
4t444c1QK+OVMLhCjTYf8LZVnIZteJXKqC9Rc1hcnWrdJINQxlfhR2GzxrYBR40/
tFZPBRKQnfogf0XTvfb/KvQGw5Gb25x0BFG/gYParoFHLQTjAupIBiWFTdD3eunc
bYoLKsOuXtQyNDjCJ2rvGg1yz2mbGM0rCZAztzVFE6OR+UXKnMTcRR/FiydRfs3/
Vj1ac8NOXfRlWmDvlMhFMHkn/zaFrsK1HnpXPyYonk4P5l7sZhf9Vggi+Jc69Jkr
yd7Tm62DSyFu9MZJA+R7QPhH1GXtnDUzwCzGChnxOfVvZz9qt4R2Z8wYU2sXlKpE
chOs2h2kCvtIUzFlFopIonhBdsCCmo3HRH6jxUqMS8//SUC0zwx6FHPF440tVoVU
WXpSFkzG4FBpXKgvLBd91rRD9assSkx3Hbt+S6pR8xqETTrtMb212lDn6hYRVSbM
SrfYj5csYsMGg3Atf6qs+UhJUyjC1vcP7De70Ma0o/Wb5xJqbtMwSIpykWjPKO+U
7vCpXXnA+FeJkKwI1nqwn6FmFrKRU/3tJPTYoYKUhwhsLvOqh1MKwYf68HdBVpuU
XKvWZKxMX5JaB0+mEyCIcQRPXeDHfg3e11ujua744gqB0hoY9E0PfiQlbYWVPnnB
GatmHFmi03R2cjh1CFBBRej/0CXnu55JGvrmRs6WKlr2fDBNc9PimN7c7kDDjBuG
KaCsb30uCHx81mHn5XohodrSk5Yu5pFi2wR6/ffzABYjYHgYea/+See3F9N4XPEQ
MWchm94kzn0ET0/c66hgU6tfXhPx9dOILCCbbKCidZ4pm3DXf2j+KlmVQUWAkcBj
w+Epp/LqbB6YKniSBUf6rqYhvFA5KY8zCptPfPLkYyse0yaYBK662Ph/JfjHDshq
AP0pSQLBkzgoluTPOnj6lnHOv7LAzau15K13XA0P6iaHjH98Emaer7ev4YVysL0/
nj2o/YCsmg1jfcRhy9YDPWAFpqw38szGbhIlcZqn+WA49J4hDasz9HuXL73BNzkw
bNuwHNbmtlOW3cn5i2NisDLl/2GpTtf+qm4tq50JSoUiMe2xhyjW8EQ+W9zcnrK7
05mQHGkQAp2T/eCPCIX8nBKZtjfFeSxQ5t37RvflxjVVudlQS+9D1FhAIFYlFqmq
vuqO4rTBf8vwQ/qjxrSvgzZ3X/X8SAh+zmf1jzOSJlYo6iPZKYQBAcaG8HQOWnbf
x+ELgGPW4kSk2eNLMtp6oLhtONYQtOtkaNr/csR5BOhafoLx5MZyoVvETKLzoCz5
9YJo76aIvKeDbnJQ6kRih3ae7Dh4uZuudxqqCfv0yS6nc4Guo9g9i7CoBVPHd3Tm
K9O7d574epjPsI97MnrQNgFn+Yx2sareN5yHk4MUaIBdiJDPdw/e2vJb5CFj/Xdm
tW6kFuvt8LWuvjy301r0P0OUpzzr1fVvIPhFgnAqTVLo08F3xBcrRl+Clmf19qkF
d8THooLjk4WBM/6M+WgByGuh2Zw6b1/6wL1CBgB0bd3yg1l1WmWNhXSjJPrHNAat
qcpFRJh/1ntvs90Mkb8innunOFyitTbEZkYVZIaF3W383p2FxLhQUzikWvYpdqmK
lAcyhea1loWwFoczqVSEMkNFOgtO7gkR/AnEaNhKo838we8aoyoVbFVfmq0Jie1M
2THwDBkEOOXY9aQdP+/Ayor2TjXdYn/wFO5i5HVfYumIzJygcMN5Jpihnq9ruS/x
xSxOtiA1yzEmDbHtlJYOlyazeFHphl1Sh/5DCzD4ZzHghp9nFGrFRP1cVZOxDIh2
89HmAOaOB8WtvyukWocZamLj014FSLfVzlD7ZNP/cAYHb0U1Bdq9RnC8mVltcFs2
fSMtvIAm6ajm4A3/sJoAJ7UtPepa3tUkKfoUQ2UL+Y3ZkvO3uGT2b8ECu3SehIlI
+NVNido27RDJwjpd7KgpDTFdoeCcxNQ2Iq7ZtY2N0FLNydHclYj8/QYYdZNSiB73
QaYJft8ijAOHBPjBeZ10Ozck8GerHiytUDfLRAxOong+dpgUCBA0n6zQZK17MTaC
9enbUciOj8dLEvdumY4dM78AnBrY9zIUdZH4j6mRTvQPZQ6H8wEbk/6ffxPKbfwk
1xNSI3tysZXk233RB0dDF9Z61JfSjfgnGhVAzFHiRaMu2QNbDOERZQPFYmFYmJ+p
usCeNIj6TqZngqN3uQlW9SVV94OQfNu1oWfHc61ibozgm2nUO6QZvFL4R2R9y+f+
TQMvZcg4i+VX99UvONJPg2SLbTyXnowJ5UAbFizIkCMexZBXXyg3HhciXsDL4Qa0
7izhtAXGgwQvPedFUOn0Py6w6RNTJCyAvUCGPQDYaC5r91UOoC1E8wxgpbd1G4pr
0AyTGIRwG4JJC4lKSKozUWmtnbkI/gmhyh1d0kq2AIeSqsp7XP5WsJhweSSr5l5J
H1Vjzj2MkaGRDMZQKE9sBR0RkXlfM4u5zVajxn/Pk2OpEHw1uhhtjxzqPGt8I2Eg
B+ciy+n11+0/X89Wu6fxf1aSmLN89hfeDj1LlSMe4fJtjSSXqXIKgLX8ZCD9vx/f
vOsFsT0uMTcnoNsxJU8T6hrfmDI67WeNIaKC9P7yhM29gmtIoMGPWzqIc5GDFyWk
6bYdBqZ56iozQR69U1MK6SHqjtmVDTVdcVluSEfyrYTHoBBK+EMJcJxD3CMhzvTe
gP/j2nnK1HmNkmPvhRgwkRdaXddByvU75ah3jMQXrl+bRkDHvf+JdA2adOG7gEmL
8qjESfE00PgYvf3JEbqwZiifTcuBMNJG3ICEp1XRHAQE1H3Ys3orMmlxqyckQE4x
UEXuJ3rjvH4637Hc0Gw8mPk2YT4UMkWU582amRktTc66bnKDOQtXqwsxsCiX0yqT
WxvUnmgpLScN6q0Sr6N6klUCu/FczLe0bAvMWKsi5Fo81VKCzXywLuEWdSOwvCVz
WF7k2rCbUIIYgV1ttYP4HGogfmpHji5eqH+yK2b8018IA6IexKA+dm0qmFuPthMJ
oA2gLqLeaSEBQjKT4BY6iQ2n/6V2KOK1Fvzp/zflPhNVQjWCbafzd2+73/XyM7QZ
jyrXMEuSypT7ns6O3aNzdfptbRQzr2uMeTqwKFG5u2vm64WHq59jusMTC6fsgeIT
haT+QjgSsnuO97VCjvsuK/PNhjK/9Eqcem5y9O9fbH7zYus3NjW8MMjjl3RRjYhk
tztjLHwu02maitudBsK6/1DINFcypR3Q02z/Cv752SYaphyfCZ1d6fE1U8VeYfTv
/Mlj5tyw+amdOiEiJOOFTGLhBhd+dTCNO7irB//r9LqRo/47kguq7l5117381DPl
uBxdnANb0PAYRZ8DUGsNVupEIcofKYvB0ECvczb2/s/O9/fDxsWcjIi1L29//SzL
/wOHXdbc1ZUyNEW4Ei663vy+VZ4TjUrFS1/oiOZ5rhkZ2JKCmn1D0gQYUZeEiBX5
1c2MrYm2fmZNdZMShRzhXIKYBQIUIP5Zi1IplkeK9jvGBja7pfLVkZb9apx54BWU
ufdrvRdYmIozpkeDUQmvqjDj1vdl1wa4JiEkoioZfoAQLcUtYOqmxAIkldgaF73r
4NZHR9uNqR/gft0g80JiFJdHXKzI/Sqhcw90oFBCBEdWGjScVX7KUwVsxHiDByh2
MVlHDP6JFF8dqfAuiricLYlr0xOmH66VfBTOgU3oiaBtbupKI79fhIPl/lA9APpD
zEuFuR+2A2vfciJzo7uVmp+M8oF1ZfpwCgfZRnYP/O/X63i3ZdtNANG96rabHzn2
etSGTzUl5C1Jf1lZqaIQGkVz9MBbuhZc7EePI0jXs37yhrparCco3k2xFBxzAjhM
3CGp6UUFLXJPDfBZK0BRcEZXxv1V34dzD6+2kvZacStUnh01s6xd0Wl9cXs+trfp
yroErDcIVbzX7mLdcsZcEklYXvg1SGAPPLmgT8rHOv7HU4r0vpd5V4IaRJVmw71U
M88jQmBoYKqt+dcGC1l+q69osaYXHgdQTi0irU/hI/WDwZoNXXkGl4esmzTVS3lW
m9X5a+Js+F+aL1tmwuAXPWFWtriyRk5VPxRR9BKQT+fp7VJGwLFu0SLxPcJqnzU5
2pb3PBG02sYqrkUCEWt2qbtf058XYn6oYSBR9hat3P8ve0UZ4KoyrgUDu+h2WPm3
5ne/wFdH1c4JGgfFJcdtqPObGVnEcRkCzQFd5bRsQh+5pTXFQ/nRkKZh6aCXXUWL
jT6zHiDrzDJw0ZfOWbGm7Tm3Win+7ce1/FhhoE4ydGoFtrgrj4pYHaOLDjB3RwgA
/h/ro3Q2We3Ak3lHbpDoqTyImtouVCLs3073naAN51PhXj03Tr7CQv/cc2MFUU7I
k7JAxPvsgxp40/IGP09sSlzNyeW6V4m7O38DbXF/pFEd5HK9/xJWNl8dmCVDm5ks
SJpLrGmDwNV7503oW33ZIbWFH5swLJkRujS4JDuWEanxN4DjoQOsX21CIcYWRFuG
5LRHjKNDdG5azO/wfoK3mTZYIFNvYRHwpxm98hetjp7TQlbjs0dJ1cQVdyzyj38S
uVlTEg68YJ3nxLp+JzNbMJFSJjghtNkFltseazBdHnvqGNwDQXXg6wUap+MjbRL2
slrmuABhsqxkSQjckizTiG5OvW/8GxPc3d1j9Iy0BoQRgdh0/7o8y5F4CSpEdEpn
CrRu4c9Rx7YSbNidIin/Rng78hBsdv0cZcEbitvL5kfmrJ+SQ9GHJT5OSypaFTj2
T/vvohsRVlzKDWreDde7vROhOFd/pLyziw04WmI1DdUjP0t6mHqSGDKSB/yxtPj9
n1YOnrcBcegavwq0OgT9nHev1gggAMDbGksW7GYvOkWDbFS4/bCNJ//LFGVT2GoP
zLbCId66vexiUK7PeHv6lxhVWsxu6xpW7MdUjwxfCL/lScJ6Nva7VXyWDRbxingc
vpYdZrJW5EwJgNGh1HQ2nXiiq3y9ECr9rcRDd5+D5FsQnsS2OAkPch8t3wa4DPkC
AZ918G9wYhvGjCiOOBlLmFgPRpVd/TzRndNv5eEMrqzAlUP1+0rUjE0LNQwhipSL
vU2ql+2HfDG17ggFaH1wwL3ecPxiYryjX6vIfZ9ZY0xbIEha166vj6vhXbl4v/u/
22GFYzWk4jEK00ffAFSYmTUSbwP9l0tWiWW6rKCywEhOBGbSYveRJJb5FVHehoUr
t18WrmmgKmRu8URsKf6P6rkMWyhSXTaomssQ4ExHN9bnbHWRyjr727C5ToGaFSMx
+SfgZscwbF7Thlr9zO3RHMh3OzpydwOdt9UH/ym4JOnuJXn1L6u64gIadskp0BJs
p2ME9mi0MSmtARaugMnEUbND9TzlH9FCgvWeyxSKLAFGVRLXBn+26nkylulywxWN
YIAKNER18YF/PABcuHH5Os2NSjklDoFQnvF1pzdjKDl5Rd7XpAyIaWvOKtFx4O6P
Ccc/QL2U+ACRTYvb0ZyJ5dNAXUBcx6p8ixc/Drl6DHEozQYqJqImYG+Nx0Sr+pzw
xlsl33gH4jyEIbhJBfGwApafYl4P2mknFdihB0McPKTD3vD4LtkI3+Z59CF547f+
tzCd5QvnczWYzJM9rrVdHOmvXw6bF7cBuRBXupYIYg/mWBVGft3MbKtZNSWKXjD4
OX/MPzIBLpq4nKM+srjXyDent6nINvdFCVRJTABs0rORU9ysZ7zKVHp0PEPt1PcW
vKu7uIrtNJCR2M4PgtxqLZ4eLXgp8PVfRbi48u7xigEohDmemrrbJM69a7WN7V6L
wHwzWUlSdwgi8Kkzf5F0RbJMY2Ci5u7AwaAOpt4/6cm4T+xqqgZvdzh3gqmEwoVq
8+/ktA/9SKtxNyldYID/M0/KjaRYScl7sOOiEi5Bf1O0vrXA3Nve/UHW1VlLetME
1d4KrME5xnePsJWCX7fIrz/6RwaGm1N4+9l6P+lNiJQmmCS59YZo721tz4pXv9qP
CwztmZ/dx4a7O1C+/8OmqmWqPs02H7KHY9+vPUKeD/5z7Y9ujMcti2K7YYlBhDBn
+RnPKhK7W4YhUa7DnR+wq0cEZ/OELArB2AWRd/jpILBRMJ3Vsac5GTneRsazto7i
QUE1ygxrpbqE6BFjIW10pROPdrwpEF6ObyhqWoZNjWcywU9BYKvDOjYNOZYfDSGM
LLrbhKLBs6QCCK9ibLLDgv5d9LWG58ogcZdblF9VrfkbS8OwJmyOlTjMTQuFRy+0
vBatK7N+pq92B+WyCtPVKiO53E6+pEX6L5vHSRIDieI5oFR0znuXmK5QNYv5xowA
2twxfEX2yjV1WcamWnS/jTtANy7R2TQEko05taj0zkNlujFRctPQ97dQg0qfpTM6
OIj2M6jN2drkZ5RSO0DjFpeXpc6odPQpyaCSlU2gJDW5PppcZje/Z0XOnkb40xrC
4YQXF3yjbzdtGTxdg0zL/TAZqD34J80mDyo5woZ8EYWdfk4j+eNL8n9WcqpYJGDj
be7o+8l3Z2v1h06p5qU5ZIHOMPQ/MBSgjtq83xazCWXcX0X69DSbrKd50H/5lMYz
f6Ps1gW3ahq9FPMUIwDtrcgcnGCGkJIvbA5Y9OwXjyaFTtbpxcjx/UGKVrema6XH
BSx7+CuCp95mBsh+t055EB88pl17qg4LkzzG6YAnwTte/0nbVeEHeTeExIyI1McC
RWZ+fdq20+DJrp3ffKFBUNY7fceVQFwJJEiIuKAL0bbGfawJAoUVBBi5dWM7lvID
SxOaDHiPXEStNg+XLdIs6Ehpi7ExPR1jggqftodJbEYThj05sKV4EYHg6SksV3by
6A6MrIJ1xiS2OcEOI0AJx2hI9+f2zgI3+uHuniF3xFfaoWR3ANf10SOoE88J5CS0
oDZFFO4/pfMZMMFw5d9tmHNOSunX1Gf4zhq/arpxVzz5M1N3bv11WjeqSXX4dYTf
rXOnLuzgHfWMZk1iQEAAhfv+giaGjrJi6G9g04H75JnjhlZ1g+YqS3Rl8UgnRkYW
tZvZnWxsYNDFhMXnoymi8I+1j9HdJGElkgVaOvDDHopRjkhrRq976wSvef9Izyuc
fRpO//uFJi+SRKzVYqTrExSFLpNGA9+F2rvcxb6wVUY+WjJLbqy7kVIQweVm6Ghf
kK4jeEv1OxnpLROoD88J9udiFJCQTIniYnbv/OnFAkYbzOp6Zll4KaHS4WU7XSJg
96OQ+e9fJbwLsAMfHeHWYQ5FUUgyCcL5dTYBXYLYcMyXmva4nY52/F/W9SlcPNfk
B2RSUgu6SJpfSbFfo9xZHDMaOq+qW1smuWtuB44coQKR1gphAfkS2BFLgumEe2HX
8+3rDYBoJfiIe5XSIioMS8fQ7Lu1FOlFa95fH4MA+/WJ6ReGo2VJ/hd4Chx82eJU
nTrwGxEcPju1edhzI3A74TZCH2Ut3hdKhLuKyPKTgKOiUYwgRY1A4ZsyX5NSddZQ
+TGPahObJFfMXyW4RxrUBkIbGP2EpnsPB4YQbudf/5ye/m99v0pXGT6UlXYUTRh+
KjL3OL9rlBjXwbwCFkxqAaYQziIbPVbObsf0QPedNXaSGKpXbMzI+1mNe+QoF8Fi
53AfdBnCxTDBVY233UwgFpbTW+MhANCjO9yTSoQzu22Ex0AkhePF+gqFT0U+6qO/
KyGdZmyElTKVTgcFaNq0j9bvW+oZbSZINRuHSoj22GoVVgy9MvVuwe9n/plVvsnp
YPObENc/hfwFFJhwDWQ3gMe1UyPYGk7MWy0R+yRrlwYPZCEEeUc7qZ6n1RHLgKm+
OChuN+Lt5EnPXM9bMcgzwwFk4fb0tpqHkeDUcOmsmvTmifjVrSAT2XoYTYzstaOh
RNg5t4mS5+j/7LW+AqBFXZxd/sbX9iuAElzsfBlciOvRHRcvvm+5SQ0fdFmB8l6U
JRSEX3KF2gHmQRb1KIdI47UVpPIEA9a+jDl+PiCXP8o1zTXCJSAL/lSBPIAbXriH
QweJnuZ2m7koqChvl3NWvIz8wq7uoOyACANOgxz7K8Cuf4y6+xwn+68gl9OFXvsB
6ZcLmiDhmWOa2faj7IgjifnigXCzGeJTg94CEOnCjFpr5AUzPpMsgEnuUaKiE7iu
h8dNchQsjTC7ZupNnnzqBDFWjbj+c02MpUtYbzE+zyYnCaiuq8gq6ZrW3I2rq8y/
lIv1CD/Vsi7JUPbvWwRGHX+g+uJt9JKwRudDq6LGT2WqiIZEg82jXOQZhKgwLHuP
2zYZ4xH1cDq3hIe2VdP3IQ1nurE2GS9koYqzSWY+Lj9gPz9+QS/cpTdRVWt6DHHA
ka2N9NhekaJxJzFgmon+Vh8sobccpvzbv70NPGn0d9YJlykw5PxJj9VTmoy5LR9Y
EgLQ/2XEuZL4TVsvNIxi1OskbJEd57+ihLI1vOOpczQENPgH0f/+Hy5pyYeOjSYQ
WzkXY7LKFETAFTj7AzTOmBCeItBNY557VkqAkWwOlwfQ4Rk4wLcjrKWcrM/39JuQ
VrJ47zeEnXBvDy54L9so4BS8bksccrie404JHVts2/elpOY9R97RXvt7MsqLS5LF
yisa5D78fsayqXP0qIYHLw8yZn1e14Xio9RavRvwGYE7RuiaPwI4Dk22hjaMoSiy
F+7ioGUycKtJz+3KoPU0juqS9H6Y6ma1CJ1vS7oqg5FOws/40VOKB4JOdw/Mjbkf
cdRaVfevyltq4BLDC5mdz+6MEKp0kJMRSP0nQrquOopjD6VC/P4tAP52mej7ZPqp
Mhba0BoKi1POP7/AjRmkZ4qIXy4CSNmgwrg5TIy5Tr4j7MoxAobWnS2IxYXloee1
FFvVrEzonKka75OvE34IG4BSQ0wdAMElcHEwHVQufDyqdJxWf24/JEoCg3HpzeWU
BIkmMpj6x47MoYhUuSrQNsaSxWDYkTPG5AYbdMjb5YIuF9IPl1BrknCKCur8JprW
5BQZYGvd+fFsSDGHOOzRfaMdfsbkG5VCB5AcYBReRX/rZXYQTwOhIjDICLwPkBtb
7t3vOr9c8L5IMhUssuCcD+zt6LaHVzP9TG8Nv1nMvdqs2u1ro3gMLWcnJFzMpXEA
dBYXcX5rLz1MfMgSz2VNYiGi1OLbh/FJqJyJvDt/ycJ1l5822Ro+B1HracKtZngl
LLc2jYv+oVEopaLlKiFzsmMyDfaQvj8AUAgxpOmwzpdNWvE204ulJ/0x7YMYwNQ0
DZFVWY1kgQsLayX3lKJq69V8gBA0NeLrXzJ213ouznKoLcKAgFKhQmwMyOH1tbNz
OsVRBCIBT6L05KPfRg7hzNNyaQpswkEYuP1kK8siN2AQQdriYP34mv1wWpCWg1H+
kh3BWaS4oQNchc+hKJ2UluFPsF/pD7sP8uWNH9lgo5J4hBnFaW3bwNqLEdnPPWLJ
JW5UCJVDB7VpJ/aiJ+dIS+Td2p1NHX3IQ48Me+dxq82DVvxNsD/TkkRdyYgExM+n
hAK08KsDA1s7kqDF4yFWSJYDpwcy53eLAwc6rmf/6vXVmHuonn5dWU7TaCRPuRe8
ACH10AnVmawayjmYY6o1suib78TMpMBBYyS5rPDg+B2eHplc8Is9UCHgnxkrxp46
Ne3OEeKTnK+KSE+/hKFUZXUsArHk/CJcLYJsdDi2dXKznoT/guyUQKo2WdA/LkMj
t22frgVeoSZqD4U+S+fJb/PPA1MmDPwV+Bq6S42hRhO9KEML+6rUuHPweKVVw2pH
t4BumbixvLn7QntkuvmOcWCg5Caj+2/RPJ1IopaMoYcCbP89A4E+U2gzSUbHSx7F
XLJdLtPQwGQLb2pBqc8LKBqYRFq8CmU/x+EwjTQ/ak6BRcluh9iWVuxiPkYeY+h3
I6qd+zHP4jauwHKP6ryyZnwTusdoWI6bPkXZbivZvAi3oJL0MBN9Cc6mXRqBtxHB
kY1P5IsAZ/15NSAqUrZUCDh8Yk8pGkGrdTO4l+QHLDpVo62zV4YeSHG29tss19JE
jy/am2A6TEcs+k253b4gESzl/E4kJ5edo/p12dqC27aYqIhwARCwmfur0HzFoWNA
bcnknyk2who4DG1tsipRiqH7VqFcqX6oua6hAA7yIdJ2D8SoHbBJ0cEMoVbRwdsD
aLunqiWDMdDVoM3kt5ooUoHj1pBaYgw/A/kdzfQwglQeR444G1b+BtXOLTlNdH5t
UPGtZl+t4HbIFiUZ82K1w0ruwFkGvxTEY7elf+JKgNXKtzRp/rrWlQ6EECA1hh8b
zArjd8PQJOjzHqOiyw4mTmBsRfp7AKkwhWZwHfk7dXqMhtbv4ebVKnTPRMp7n+wV
Wq03vtNuY1QdTQG141g6sWlU1ckhTzFGWm79mHA61hFazwT3EJIkhG3aXdmitHBd
FwShU5vV1JurDwgo/xyKgFs2Z1xFSy8HFRd31jj0OgJNkf6JsltBtc4OzzqXZVyJ
N4VQIgLej4nTprk9mkCT63ncB8VS5F17N8PrI6E4TnqujQyybtbWzkANSQ5/oS98
KwlzVNcqNxLvVgVCtxcXTc3LIBOJGrdG+uxMgw5qX1aOzg13OkcYWjfKNTt8eHcS
zyLPvYnfIB/iM1Z71IcF5r6Pv84NRiUtV+QCpU6fYLXVExgg0HlNVjXYOqJrMasu
PfnqLXyab3WV0lbMxeYeohxmArIbQa+X8YIzQkE29ZP+xuS2s5Pacy7yPEMuH4dU
kxRXshvQdAwhAtDUcKGhCuH4ppjO19fpdEx94zrY3sHR3iMp3/S0/0evjkrHPsIR
aptDr0U/BGsG9MCMlJIEahqJ3HlGr2/0ILIzZPxnYGO6a9h0A6GggJmvL6BdGYUX
x7+fprmxXbYhXw6kzyju98BJay2/l9djg5rwb2RS62+gTeY9THo2nL3nYaRMjJXm
98yi+CDZES6Br9BbmpeJjuERiOQ8A4Dn0PuIi7/srCsy9C53q7V+I0gKtnASB6ko
cmPx1dZFNHR0aFeiDwhlP9no4rTUiUQqHOBwJWG+g7/q8VIRO44UNxHvyCrq3NyT
P6RC8CRn+nTnVydkZGqhHz7zyjHYNVNJrvZM99rTqu8=
`protect END_PROTECTED
