`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBOgKRC+Vh/zMQ31cUjipLbngh9oyKJTELHF90mrbS9RHlMipciSjWZvCPuuszjS
B1kNN11/CioGg/HZ/V7R9NJSXnET0lLk1GcA0b7jzdV8c92e6EaDa+V696ZRYcUo
Fr8AssQRjvkGoKQBJ1DBKPT8OMw+w9+D0vXZQhIXb7yl/oGq/a5yXJQrBq0EbCpX
p9GBnTjXxoHg67qjqQkpMCBUcZU12yBkZPbDvcP788L43MHTxef06w6BWWcsxkTl
FKS5MKohuC1qoaWWuQiEpddWUL5Lsb3GTnp4EUTzvGVrqPSkq/7T9VKq0KNnT+7L
C9zQoHQvuEG9+v/VlVyxahhYvFeCqtpAxDhPbKh9EZyp8w+tyY5fSBz/bZSRZRc1
T3PoaSsttH1dlJet6o+hgN0ooajNpTBuXC+J0P/DwJ91+HxfERtItgw2FRB3XMj3
qL/QMzEIxxz7UKIQ4ZcgDmV9pEL99IOlCH4zeq9tf/qLHzplP/cIZLIw7ADxyMx7
ZwzDour89CdZcsP+giCK49g2+DbkskLRmHITWtXwT1h3cjoim5Ilyp4wt4kf+Tth
4bABW4rQO2zkRf71+AHTfWy7gezo0X06gRqq6kcmN1Mq3uErnwIxsFFzUxy6QNWa
2Sxkxh7M3swSJa5YtDa3M9wpaWDzhv2EQmfMOhDsfjX+Z/Ll21x5olS5bCNB94QI
glSkTrtEwCk9NvRsTTr+nvCp2VqXS9vRXglZ5lqdf18i5rue3wHcp1m4JovQhZkn
lrQy9FOXyj75LTskj4ovZu8DlMd7S9ODMlVeg+PW2PI0rtFfVpz+5q05sr90I81V
XMsqcek/LTOs0CMebt7PhmMuoWZBbLRgXILiktLDPLglD+R8tPoKNBmpg1+lfHAi
dqAUJfrXlDtKBazWrqs3W53jouoVvacJtRgVc18fYQGvRrFmMVVITWhlBuYhn2nD
CLVgELC6ScY1NF+9tqBcN54R/nDvH2Ab+J8Waw6XPWMBdgC0rCb7L6Ju+ykGCqko
k8HbI1RXWZy47qfZJ7VvRNDU30jiz824jXLu+jJqyKlolkzqw58FhYgwiExFsgbh
4iHqjs4nfL/M833uo9CrCzIbS/yLWyZD2RtqZWfPqGP8t7q3XqsiDi30r6LYsvJt
+RYSe0UNjxK96Zzo9xXRyYw0Tfe0Y5Z90HqHARTTGnOcAROP/HUNecukM9LC2PdI
hJw9RbJf0ivQgYz67Z9jQDBy4XL7vgMzLY6hMksXeuTywVArB05iFmBzTUWtJu+U
C7J/CF38wPHtd+WHPmWpryg4EGkANuax8qdEl3RHKeN8hy/+Vxdb6fSzNi3Fe78E
Mh00Pug5ilKTl12iel9teSe1P4gRpR7n4ATo4aOHC/3MmSHc4+eP4Rp86Gsy+toK
WtVqtvBHuojyh9hHNeBObVXj8cpFiPeWA36jXYQmd2QyrZAfWBAaBjidNILMowMv
8pk/wLLaCuPu6E02DU32cBeOGjDZCtbb1snoTgCXKgJEz60XkhsNs2aSUK4mYUtL
53BIcUXBGu3VNPQMtaAgAcB6paq8EKRUOmzwxggYE3C21D0ueMW1NCMS8WlxT4Js
aPzHVLyMfxMe96Pl3I2oPLCdf3/MQ1butl7c9S4xU+Q3dYn6MVrPGj0l10Qaj8IO
EGdaTYfRWKmWP9QwQaRjS2H8958QXLmLHcHnHrJ9b97sfHKoIK0UsV4aEomvX9Iq
q051jPkYtAU7MyMss8Ip2Lk9NRXldCavFFxtn8igmLeYDrC53P1YUBl9JVWz1vfL
4/8H2Zju+sNP8223W25awtmV8ybYQTJU6dWjN6WSEYqRVkogej+awirRFHOGgL7z
woCmiDriUpDcV36WUCimvyeh9r30MdHO2/1AWU7eoY0asMp7fwuRPmHUjR4LyyQG
uaMrX4leZtOltz5tMSMQxQd+VX78Gy36TRVIa3jY67STjJ2na0RqZQtfIx1RkImU
ve4w9d4k5XKoVOoa//mm+SQZU3JyV20UihVFt/TiehymxQYnFPnsnChQMbAvz0MB
BuFln3+gGVdn3t/rSqx4DCwTeYL68tWjDXF99PDs0AABTOGqawhrSsNr/3JIXUFh
uo2Inc5KALuDLsztp51lP4xBST5BwUkZF09DJv5PsSNhPwyhk3w/A/9EenTkzwMd
Ho0tyf9NsRCIJPpcufnV2IOMEUeXdLxT4uy+nFO8UA/RuuD/TSDQWf/SUab8E1fn
RBn/gewyrEphvdUnhkVcvWPqZ42Mk2mIq6SbU9KWNAE6ttSHGNm4q7ALo0fpim4q
tLO0xIfHmQS9mgSYYOdSRDZKcHjUjkea4NflrxZsw/X8cwfxsc1UtspiXL89epJs
ekPIpac2zo+W8SlOTfOMKzam0R7Mn5eSn4znX9cJVPYPBpFKndrdL2fRLuIktogz
3OtJEMG4B3yxpWONfFBIUzaHSGr4bnBcm29cs0CI7SFAzzvDEp+lhMaUMKCFla0u
zeJJmlL/pw9ONiYveM6tnM2sXIpwSdKfxQS1APSzFaBCWWszndmywdk8X8LnlcZe
ammo7JAOBjkIf/k4nXMvMd5UtYQ+Wr2WVakaH4KmVu96QUUhfHY5nmWjwqRIJjhl
bfFLNb0AJYe5OcPe+c9t54fbXgghVpQDJjruLjg/acMKjRIvZQGWT4/pgApe5IaO
eNUrvw8CuKCMNkfM8mbzVAAQplDB+ENqNfFfBw/3tKj7o+WMbD/SN+NfijU0rYoR
4xXTF2KUJNH/b1XRkrxpn6oyG8Gu+u7dil2gFI6B4Tsou37tF+BCtwcwZRTlqMxr
QmF8LHOSUFHqeSJp6yh6DDHi0iDS9NtQBj2lUKBmgzb5nJopN6Lp3shoDB63HDDO
sitzrn4OHhidtXX+8OlSlXWq/HJCXnJsQREdOSPCuM4KsxEsO54HqYr0P8BK9WlQ
TYph71b24CeEyfNvcfSr9rgCAuMBhmPC8EywKbaQ4e65l3mjzlYKlGrnfCcjQR62
3lMWXj5JpatM3cvdDHJ05KcYDIP6Y9t0DgcryJ6KgrvF1XMWlABWddTUfBo4Z6Tv
E75lqvkSX/dj2yyOagSnZGsFyKmfuTGhsC7CiU/xfDm0rGc5dOI1Rhev4Vz7Idz7
TjiwGGLsD+7IbuLaHDvuTaVhCrnQPXwjuh9RHN3qeuFOypclyCBkyY8ENM8nRbpO
jCnhnyup+piIawpZCQfLV3XSu1SJFO5aHQAN1x4SyILWpZUjZclLYezCkAA+FFDU
meuLrNmhnR8CocgzsLEvybbbVB/GO04gVIu1VkkAmmoCFzIV+rXRuhKWQKzjKajN
F4QSPV7evL/ZuZSDQKg9qw==
`protect END_PROTECTED
