`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FAUQCcvjDRUKNBgMUtJDiiuNi2sO3mpPks8BVaUJbb9NzDfxabIKD7Cwrtf7xcxV
GIK/Y8PXm1ZnihWtcmdMdS46otXrY55bmSSSJon0EsScJGuGghHrMWC6DHq5n7mo
3s8sCcPRVyQDvDxRV3iGg7jOzpA0a4Edqts/y3p6rvL2A2w/9luW71fKXr15ZSA9
Vtv95K1bdvGSEBpM+7jEI16Al4W5jMgVymhq8EJciuc1bpvNI2Drj49YICv/gY4O
9YYO/Tx0ugDhpNcb4vvXTiYGl1JdWDczSLnqRf9NMTkh0ICB+/56zpfSNxXRNJ5C
/2gofCn69Fqcb8u1m1YqXn4K/FdJy6EYKYJESrTPFLHbs0x2HHCueWuSqCzOjLQ6
2d5HmUqRrNrNFSFIckpNdPbbCyfuwyKaxEfMdRMjtz6+7kvC0KiY8ig2DhL3uUey
PHq2+PKKBNr5zZjCyBNrNpagZp5Qqcl99qg6ZenyH11TmA+EGa/IN+smB0rNRFM1
TBCM8x+8jlNf4sHots8a0w/RcuPoRZ6PdjmP+Ins0BIFyDGYFWJaq4z+jN3xDbdW
cfYW3jqLQ7+VzHkdHqID318+/B17IixmwHNDA+vdxHEUxB0dNQIBphbvwsLMSxvZ
CZG4EfUqjeIlBEzVPKn8FEVoUcuMh55Jrq//l0s+r9WGejXxfJNStSyD81UnSdyw
aju8anlgJ8do/Xyt3md0B9LgKZurgTKBy0y2PMr4GFdc339X3lJ4dklT4IvqxBEj
PCdA/GnS+xf+aco1GB92nFGMGjhRwBrYCtoYl6Br9qSZXqPNk47AfR0Bi9LVv9jy
PAnMs0NXBV9YfQ8DayLB5ymH/WmaajCHd7E+73tGNwOcQwuUZ0DmhRDz2/hdt1V/
wpoWXwb1dAe2yldhmNAEEmHMmiTCVt43z0cvcnMO1DykQL4gcQ/hYqWXUFBU4shq
/lk/SsrRlgBnKCJHJOyHx5hMbvruPQDY4E3TppfKPWkzGb6cbeCnN8EI8zY0HGcI
t6hzHbUqKfkz/db+fKwpkrV06LNGWjQFrzXLuwIhknZH65HaBHTlefZ1k263v3Mp
IyGWswzxflJqx591MQm1UaDSrUWOhAXgUfMO6Clt3fjQvGstUqZolkHC6X5iLaGm
Qoa+pSK5lLS90jZsQz4Ha35FEMr33gzKRO0geIZg4VkXu6U+db68X1O2dIu2lDiF
Zzbicj/OQGPK+NypjdXxIRbBMrIHQbU7Y1q1C8pUESkVqj2v6ApWyhLz/tQGyFMG
gNvgjpRtWXtW/FimtNx1+qfeTFAFz5spb6tEUvgxr53IUqDYVKwc04EiYSiaaUpB
yEr+eYLjXuXI7ItsxffVdNViz+0R7tidggelQGrfX8xYc2D3G2M6cm5a7fhzYX37
7qH+KQDWrqA+9r1xMknSug19gB9/f3uPtY2KzoqAn9k2aPViw+EG88huYoJ3lKan
YGs/hb5j3RQtjtHOSX8ewreC82X+Sbppau7u4ZVpww65Tx5gy3eoWIC48eSSeKvo
tMwHCoLXLHa0dm12SfqTOmunPrfc7pDnG1/PZhJxpMCV7/EYdDQwr7gp1+9q79t6
+IIVyXYvDf4rBrReKpZSM3/ac4CRCSp4B0RP0oKlbcAt+VXnQgvy9rndLr38f6gM
usU3v7M5iH1aPPyRMbs9IYVd+COpe9RxHVpCBxF20DVoy9W8uRltayClGQUKrgF8
5GyLjDTpVIu8BZWEvfICFxLZC0qhEcCv5Oa9Z1y1IJOjcdpH/0X3R3eTPCSNhR+3
CGIclsS77KKoelKZbBTdAdwQqhVrwvQLM1mcoJ1OdTbnhjG8j2P0I58CQVXODKEa
xNva9lhTqEuCjLjrnJKGYn2vINOMI9DIDk54+2lOfMuDxsD9lRhImMgc8USnaQTp
ymRYKZLJl/Qum/1u/7v+Ty6T/vPcGSyKkWNVEbW7CqOpX71h9/SndbKxtvGZEhHR
vS2uaEIcYYAiejfYNSwEwXX+1RhZf2Fq08cnO+DDhU1vacnSbSRt2AWORHTSjihx
693829cbaDFZ1KjP8ZX4+wNekYeaDUXw1WWW2ttn8NwSPdg46hY2naTUbiMCNzud
7kLa5KIbP20ImuR+qH1/fy6GiMPYzO4krRNGYIfBcSNIoUxRQnTwKWv7o8qwpVVO
71uZKWq6hsLCRaHNzNX4G+dM2D3WNtR0Z368kzPm7Qyfg3JzZTeXNHU/SZ+M+dlo
hVyEtSzLCssAy+COPp4Vm83LjUrEaN0y/jMg//AO8jOmq0FmJqP1JmAEUTol5ApM
D2h/id028HilYN3cT49Fy+OtCakBqklrpG0kJoNxK1kBq2W/BSdsc6NOsLgwQGgZ
JvgIKTrkijj2ITf7KECfSQz793PQcQrrwjhke/GoIblJl6SPZDqrNUkjCthsvmKT
GldG9n61OmmY0hLZITndGpRbqO+t2tcLm9Kr8nQYdZSfE8uiSsbcE1RBPJLg+kUw
H+ZgXuOxd2fyuaXlzBqpN3/TvDr4IvfNqWQIja3UquATjVWsi4zgFTPdG/KF95g8
/cKfX1KcFB7QK4nyH4FblIlriv4a/z1l58Psie6lN3kulDkDb99DxsvDPeNiSX+O
9WH49UcPQrpttT980K6IlgB+46rxIvMILTs9UKnPCrQpzSDirHyQPoIunUNZYhv/
tVkcfozHy1dZplOkGIoO3KXNbMw5IDahhvZz3lhokDEPaHD39J4r/T626iY28A3j
o0RLegYwuiDjex0QLcJWMqzQemKar12n5vFf17ad3HgrdBibSUnrunVBTQkLmFEb
8ji0sE1OkrGBd8zN6O2p96M+HcNPIGffxOZcW+Jc4kqrWH1M8HDXP2HgMAsAlO9l
zwDbVuM38whC2fIfGGqvpW95xCC6btNxp+Cs8ga3TZpvCyZoAScEiuInQKsQ0RXt
i847UYplx0mpXknkoFivRFJR6J8vYaJ+V9JrpqZHu7Ao+fp1mDZtwnnNuLYuNCgI
TdlXjZzw0kKb0Yi5GVsoT1X8rBpi0syVqpoLNreDQqOCkKnHVuYaR+0La0yVYnSF
lwaIr9woRk43B63xnvWdOKzldZYGmu+St65hzjCq3wnd+wfXvQJnN9HKEguwtVrf
al1pmB/gBbn2KMFYCu/nLNSgZjMnSEyAUf0xtIe44s/zfwCENHsPZ9jL7CEdMH6n
Z2k/fBhRwEZ0mdEMbbVaWBHVHMfmOpjK2ispWDJSpIFDhBLIC9hobvkKOWcFzzma
1pJ3WYDyzTBBY7NC6WCUaBsdndtiwyb6vw+f637HpVkZXIJy13NsCXqp/SwCDclB
+xxZC8MdI6A/ous1LcKmpxpblvMUrobujlLNfqHdx78FziwvVpn0mxZSsVSdND92
iE5mm0OK0Qchvw8LuczaLbjLuJi4WW4iLGanojTRBOFPxjgDsAL6XF5r/qytmb00
sA8R3VImlOrsnOOx5ChqhN14OOl+7WKaH2QY76/wBaKlk/UgbiuTtJ4ema4t33OM
o5JXOuvTARvmD//lcdfn0Ebochb8yYtKNgrnpSZDt8c24lAFMTxeUflUe7n/Qsca
O91CxYdpXRCnm48xfqk9n+rpcA2mwUVgjjizNnjip1V5JRQEV2z7I/fzqfDaF6hR
helQsTmvt6wYIcsRo3NVtlfUAq+/Mvuf9paju7oOtzmSWqbBJ+J9xWlI7urL7vhN
gC3H/1Fr7aAKoh4N0/4awERmoprRA44JYG7m61U8RbzxWdjaDBvZ0E8DySCaJEPD
Kypqk8ADdNY8GUIF+EjZ0mCUDIjeZUCpCmh6Ap9iVwD1U9Yk+8z2DYBw2EXLa8Ud
fiX/e5pgeruo+qKtXddvziWGyLjpFwCVqGGKbA8q7QMGECUHzAbQfuDiZIWtplTT
BCrtH7cr+fZkQFruWX/hlLwraqLcRiUGm3ar77d+aiTWQuthHn2kkKo0HsPtaVNy
q/Bx+1sD6dirx0S773Kczrg5pgh/wexxbHnQ1v40e1rYYBHsEg3oZOO8OQ1l0rl/
1mK2A7m8GViCcwz+1iD8bLE19BiggEogQvEZ8qkf0S1l0w37z//0XQZjQuAFXGTe
/OGEoWIeOhaZQKDLR1AQb17bFAVyOnBOtGEwqANoWU1o69zrXu/EDVEHKCRt63cN
w2y51wx5TqoqbNkKzhv1IlCW7olWPci6tDtna0NOIQY45YivQOMnZDYT8+ExVSPi
P/45IgMk9KfdYZhlOuE1UnN1/+23FWy1FX7L3O1olJJ2WYJa5eIKFdDZRNKPKQ55
QqLr8mmHZlKW96Q+w/MMWkyvkLijMhA0gzSAyyGXZzKglWIea1/fRC0qidaUrnDh
mOgo3kHbaxGLUvIRUfxK+LZduVEeukB1Eq3tHbJPoZLwb+o+e6wFsWEGpmrQUry9
aLNQMqQhnpXz4aBeTa24ItfOgPZ+zf+92l6VEH6rd6Gx6IEDly2VN9TpaVeJOk8+
0RMegNZxgxqdd+R63AIkBFtPaN4ttyaGIaQNQRr66WDTbYS8x0wI10Bu814f21pW
b8/qrraxt6vrChaRuDR1NFtJ+/tR/+FoICK97Lq/Ke4rHGVgG66xq8IOfrfsvQ8u
/lskFk4Du15Wwmh4qkna38Hio8fyNM2M4GMjNC/Qouk5xOSCnjhZutXMb1hWLCWE
hUZcGp14JdaSGzJfKnk7uhAEfvKE4gqaMi3idKqlFnoTUrmQY6j9H/3lpeZQvb1I
CrdwryU+zs07SfsbSVOkLaVdUMpt9xjyIwxzew1DwDKq5RFr8c30TgZ5vM5I0kai
bzf7kktJJ0Zzcr9V4RjncXFM7RAV1nAvmBn9b7NfPLtFH9eILH/KOWNVG7MDdD1D
JfPV8mqSjdkNfeEFQ2ui1zvYSrBg788GRsgbkhlhgfoLz0LdCije4pY70+BdA+0Y
ABR26DmtrdQWOZm9oVx9Kxjom4Qb/nZHVRJ7KDdBBLNOZRnSN0Qrq5QOPdAs6tvN
NSdq9k7yVgv4tb6N4O2fkdwL5dF7JvqEBj0OoKwQ/J/sWyY/mX2BGmvzI4+PaUiy
rajG2yuLkheiTAFe6vCpo7EpFhuY+o3FdGewW9oX87UqOAQNr272xr5PRJc3uERh
n8Gq5Wtq+FKR9gztTV08mkGoA+8iHcy2QwMyNAZwaIfE/NFqzrQrtgvaYXBtYzZo
vZR/u6rcU/CDU2G3GKMjKotLU8gb+IBd311lH+VioViOA44Uei7ez4c39UtES9N9
HKJ2/y4gEddu+oda0zKiJg0jaP8KV9wEL13BIDt9DLfGY2QRt5lzYyXT9CeXatkx
na78QvJdiOtQSRxur2uQ5hgmqxjBwAi0JoQgwlncDpFVfPanNmJYeLf4WQCEcnaa
0gxdogAa+EzhhB9NXSIoxPf6Tpi7g5HHGl7jDymkIdoHKoa67oq5ND0hk33NNrbb
toICSYNUiINGL58sKoDOZF29T6iCg07Jha/iDnSxLdOTdhFtG6boz4p0IIlerlv1
1kc8d3xxyaVfRHWcMcyEWBvqrkyd6XRz3b/HbYInSUHQQJgCD2iTdjVvzJRcJKv2
NUpJW8bFlWz30Jwe1ocspb9GCL6Eu7SiR7yoHg5i3/VBRPeKlca/3y8SB2rO413z
FmaQ+0w5OtwFhsSjkIWU1niQTwPaDBqeimTYX5xSzlCMSJzkk58PkUkDCZT7wzQ2
EjhifBborAvjulwRsZi2v6EMaYWykDUEwsfjB9S59JqQoAtPqzoGTizGpXUWGBlt
nH0repH/6shNBcIzYqKH+QMX0XmFsF8ywYquBLGvEkm1re9zFaKDJ2fbJzzEXNBH
jb0GMvj37ObeyR+U475Bz+Y1TpM/q4F2kDiohWIumWiQ2rM2pZcmsPql1Ci4KKIW
OjYmCsUCt/fF3TcwfZCG9sbFtlaXzHnbkTO9JWpOHHM+UfrKI+335uxRij8iSSwd
U7O2ua7p0chlmNaoWLD0rIgaeFtjsgCFytdV9AiClJEidAAQJkOuAEMb5zWtHKW3
yl5zSWBl7xw402dqLL3imVEhYXr176qH8TXibBPe0fyW4Mdy8cRpRwSjyGMIH4ek
SnYayrKkvAOHW/8iZijiryymrgrH2xlKgWKRbMielzjhYfZr3kqlrrPJXgEfc8ix
vHWAjhGlMI+yEhQ5ymDJij8unjBuzSVlyPbr/8Tz6Ztpqf6zoV1dwwlLg/+stOHT
P3rcTqhllMrz4qqbJFxanI5G8WYK1RcuZO4kyABRdKMm2GOA/OtAkN5O8BszplfL
DuzZ/w2MXua1LYxzZcLYSHLxdpOWS8SgW+AexUeUeCbtowkdpI+WBipMnY2jFouo
C1uM1kZ/1j0S5M17cp9KrjAesOxbXQ1D6MpFzuirMQZSvrc3y8iC+1YWD0h6m+ov
+k3BqqxnBGsmaaUfhYwRmjLBIbehS3KZ9lE1TSUje9XT/pLmgGEG57nVlRpNtzoD
ZfXvrDkm43+kT1jdTYTuXlkTwxDrA3WMxhUFX+cgkP9GJ21mW04xSkM7fIqrsdG1
DwgwpymMZ1NP/SSw6zjYjbpNoJLV4nTZEQGZVKO/DkPJIqyXAI6hrjuPedQywLpc
80fWbERBykgSf8206GAZnAQoJqrnEpTtUfIK7ps6aodAM1GonEezqtAjsyUnqMcQ
ypnQ9nGkReiTYAMf6ovtXKu2GjKE/u3zA6X2zrSdtGMK6YRUTeJo9DOrIFl72Ftb
3pG/IiEyQK0wYoBMfC5J8hlxKzhHS+cyhFZ/KyWz009FpS29t6tjTT+heQVA0EX+
mRxnPVoZkywTLEh9GradmKOlwZmlerdb7zCjUmgUJfKQ3+oQRmJ8LRzG82BrfF7V
aLlT04kq7VACItYWT6/xnVqUzyEQ6OdRnFBffm+RnwDpE+Cd7mFn771z/SwRIW6v
pveL45/4oczdMso1aTCfZKGx7nsqm8N8e8DPLyROGK9eHQ+i5xvTxRrQqlrC0WNA
vapW48GFG7Xs/+DBD7evz+EEysoCnftlCn6ewCeO9ud5TAO28jdNN6CQN6umr3dv
HxvFNZZvht+K8p0vDDOi+W45RrZAiKHs/Wr0gyOd5pngjOeCaX2FVlz5hhCTzpmU
bG+OvIGSSasmsYaxHuC7g1HaEzsatx15XmQTWxRKwBlfn/7KP5nrT3rKYH4dYfEw
hqJWOfcLckHtsmALfzgoSsInHinGHlHVndvfUqfq1QbiXuMzgYBKn9ljdrP5yxAE
rdm7wUmU54yv3QAwFj/Pt3RYRTGCXIojJYTo8LlSqXousJqGjs0T99T3yiXAZhnD
vETzXd4gmNZ7JFwJABib7V1jiYhC0Bi3mbBk4i9OVf3FbWbNLPFXUn+JUZ3FFk1j
ed4470nL9Ds35mwwRUSqBk9mak9xzdKlk8jN1ru+2ruw0NdT/3cTVGMYaaW1bflr
eNbE8t36JiZJn3vjOELiL+aoSOekhZCA+XKtGe/m8XUQSB9+Gc/NyO/tqxN1hjTi
yzhnHTHlNYLXEAj9OjzBe4UpW1eRvk6Ca9PeIdBEyvm+GS7DKxe3+47Xz4Qt39Fy
rLMIRyd6YXJOP78lW+9KVsXQUR/9e2KQhB5LXap0fyP2jbvm3WO78x2HB5PYOVyf
gQMUFSRw/y6wa49oDzHrBT2gRpjeCscd/HmBF4jTTMLtMCD/UQflOmhE6+yPCJPR
O2evGBZEQDIZwAmyElmFgYs7hyC3YH+96KdfKkaaiF2X3TeZJGcqQYwzeL1/Zxko
FluTBVgq4wxxPIsKHqCh2yPo/1iYeyaGmLloF7LCA6pvU26B4Qztlq3giU2Mt8I2
jTHRyEsCnAx6RPP7e6CxZJQ9nGRDMojm2g0wUyKk0N7x/R2GKGYXNk/7NK2fJZPV
9XSLPSYk5bC2a2owBb56WmBSgVBEvaLXxcmB+GysYHg9JO9OGY/b9WVtAaIMH5nx
GQFsrf5Hn4xcz8NyD8JAZ/cL8V3liYDw+6UUsrluZA5X1xvBUZQLTYI4YB/SUPQL
r9+LLQetTXb0O6r6US38Gpye/WqvmMGoCqWnRq16ZOT7KNAAeApCMfCjCMFF2+tL
0js/V5lO78k4URxv2YE+uXZwUJhoGBjupPjjkmbkFJoOe4i4Cmvqx/pi6ZFRFkzv
QDzlQ4JXEHENWiBYzhh9ZnrMp2Pp77nYKbNEZYtyBVOFr2Ic3IPzz3zWdmjyyYpm
+R430EogJeymHM3pRv1nsuTwDZeqY0RdIEHLc/YZ/vC0iBHruvx33xnLIV5Dlho8
pCWldmb6hde95QgAMTwgj9jj1+1/N2GGenf4UIRpnSf+U61RZhZrjxcQIO1yEeMq
ngxGp3kBeuiMurHJOkrcc5MW4vX6NEZzzjzEniPRubpjyorO1QD4ZVD8GiaDkLeC
OSPU0521kRN4vVHMdKMR/Hv8PnRgkqxW/DEY1ZjZ9q3rGPl+Dvn79fujR15pxcpK
mjTdDadHNVt7Tpbd8OWfgvWUQuynTezIvnMxRg3rm3Wwxca80FS44QHd+Byn8YHq
6+1dZ0aW2K2XbmVjI8KaPfrm/1gJ5cOlAbojQfpL0SrFWtHAeOUAlq505BinalUG
jpGxcDBK9JgnOcp8ngy9UHS5GPK9N4IzXla+cmrgdYs3+qTIF7c1aPswyY71gjXA
hphWXP2fQdieutqqXUJKTKmU+Z8r6fll5s4WEhUCPsOxvqAKQyIhXaASqieeFBJC
TuCuShc8GuFcoX9XrD6nM7Qh08XiK56WoTRhAtoYx9jjQ+0K02ALICoSOM/uBT+g
FOeZHcmAUVUcgVQr4AuRe4u108yGGKoiV0DSHL0YAHiPybwP2JmUxs9g5CChfK3V
2ET1xtBrMjfdIpoX1z0/0UPli+kQn8bY+vKwZM78JjqCFknK4orp4f1R/syxYrDf
OpSkKMUX63gkNzzgbGK+CxQcm1ISo0NpslqRHfiNBOEQmXzPi50snnHWgy2hBiEP
kP/rShWfEIfNR0ohHCL+rY5nI4e8kpXtW0LO4ALEKvRhEjEXNPKfhnxkJdcQsvY2
4x0mb9qbWcTvT7sKMzMNbOQOL4zuUTeZILKt90manH3sFx91hBZJnXzRUS3fByvn
9NiBVlHoxhJ0AYlihyeiVCbcHuvecuOL9E7HyZxHozo242T/+w4l388U5ZD36A5O
vcE9QjT9Rj5zeGQXcTo13DY6rEGmvFvBuYqKAfL7MtTo74Fj1uh05Er8p52QLPFi
Bglco+Z6RFK7S5ikF6qAQ0xuXHs6CceF1Ib5cHMW8/04jOOQ5/ovzUD09nMPmjjv
o0cjR2mDfsTwZfXkzBfXoZLHINn3WOjyUJxpYdLGSA4FvO5awImf754CPaJDeRoR
VM9je0Wh33hKf8HHAmC+SWRS5FB71db2RbhtuTdecdoayFUJowRym93kWZBaP3Yr
HycNcclipZecJ3DY0dmd+CO9HArd15/7bUolxKV8G8KEDUtFwALR6yuMqT1Kv7jg
2ysiMAPAz4luabMZ+9DAxb/RZAYWHhXzXo0irGACtvyR+OjaYPG4LciJPb1XiLhJ
16Je9Kt95tUbqoNs1qH8pUmzr3soLl3SGksA7WZqB83wy//rrM+3PNmjHiGCOuOj
rH47RUFS21kMedCX25ITrAAToqT0QoNc9wBSd2Jr3Zccpdvr6R0bCzRU6o5mJ/Wb
EiWfiNeo3ZQiLTDPA7HWSDmUOdu1nhzafT6aPMMXDFkCY/7euRw2v48HY7xT0oMT
K4Wp7kYeJWdXSlfCK0yGekEakSfR+zZx6CwHLNlawbmVtBzJ2054/uSNowy2Lo+K
yqVuJBwpQ2WIF8gQ64SxRbvuyFOAJsNy5ooF1NWIEoHJ0nMWrfZ6PONc818QhivO
JPjE6uVPYUh1T4Sv+6V4I6tYLCPY4yxW3CiEF36t+RKH7ukELfdyB8Q0R2bld+Uy
82d6m+czdc5nKWyKu6DxW10rC9LVmwTPkInDopAG9ybpl+CL+K8N8ryY4jw11cxO
SmhTn0tSHSK6oI6+NHW+XZY5IJNw6Fd8GzODpHfUvJZfHZeQav9BnsMkCP0lMryi
uC/EajbSFgqLu7THH0jgDY+aPsP/qVN6olfjcpinqdf9i6zZpW5WnhpdI54VfZFl
NDP8u86I9MXO3Jx1BPVm1C01xxQTeB/ay7gItPY4igKWi5UcH+yWapoYS7/TngUo
BpX/9tZr1OWUv4yTeKF+TGNYe+ZPUDZ8v5HbWn5UCocACDWIZpykSiN01Joi4r/H
nom0UE44ebOf+LAZfOBB2o2MTGYG9xnxWWS92rJOKZzjAP/IAvxHlyPVDH69uT9G
ctA3byj0IUGI3HbU629sxVZD8cjE6e4BMRN6x3fIvdHeDFI0JAnLr2NQcYPe1TvI
N9HAe8r6LWl7sEsbGxCGH7m23Sth89a5odbfPxFLSQgbdG0mBRpWPViDhYz5EKy0
qlwwQx6nuQGM+ymfL+FEe6j7MOIgQKsRX6vxrd37QEilCjmm/8gMQ5c9vIAM7Wz1
0qrlrx3vcz7cWWaL6oLEOXqUTR+49tWOeRt29x6k4NuUQT0fGwM9Ac1rTl+xWAU3
PZX+JVExF8PIBtWCq7l14TLNAVXp0eAJAt1uJbR9eatRqynbM8jaR+B+qt8ZC5kV
J40jkk0oXwUC5iG7MwUCivxwm9TeHLrRvVG+wzMkC6hVB5EDCgUi4uA2e+iiEBZa
HvUenwzdzWZjKxXpLSg/CLwO40utLtNz+6tvmv7MXs5IkRkL1IOMrBpLFMfQVpDa
U0k6fEiAoQYldZeo48/rAUiUqhvV4F1xY6euWm0i021shylJ0t4/0tJoqWSfAe+5
qjWi02ArbGRreCZNVDmGJm3FtU4VtWXKhcUISbwu4q5VrlLIiCXhuKHIfgFhQPkS
gGnQmTvDYif1/XqnWv9rgYU4a7fxOJ7p2NBpD3E2Qsg8so+L0WJdFRdwB1/wNdHi
ho1SaEUL5NHID9dOfCiWPfXmzlr+tKkgwwScX8D/qb24coc89otFXWoDxRuNQ9qQ
SNg/DQNRrrLhhqDfjsCd3zIk3tHblKU7QZFugz0Bj+G4dIMoV9QShljXeY5Rpdhd
PA/SH3SHDg5MtTigH1KIyCpkqH2U1n+RRVMDtlH8uCp5V2BSaRHtzmvfjJUw8YsJ
4Fou+8XeVtvVHFzGwxZsglxVva2diXWXTGgA6i+l92/2dtYxYgL2YzWyKbCEbUGV
iTV86/hTdIDQGZibsdqvxuCF5XdvAuDLrunPgQVucjCQT/eXLLB64z04UzRrBGDA
POG8/yRkOtO5VfuXJWCIcAXQy4csw12lmspGzj+19teyH9Icya/LlmHY8dQHJTAS
x7dTZ6ALpRwlHZlWlu1Ffo3uQhlDuuIThWZrvhxbsqdzCKmaIl6x4HYQA5UWxR/3
BFIZUsO/H1ffdaYLLtU/ykpSolH4JbPL5KwttprfvIjWqezGzJ+niS51ZvoXpoQ2
xpmOTwubfRxDm4NpKvBPJiT6EUn7DLULBiFpJe6AXv/wPzC0/poZULYYf6wrsD/t
FKrQDD8sBzHEIYkPJEH4voNOKgUq6oEgAkRBJ2sMkTtLiiG54YAcH85wytoVCAbN
259cOLUWP1OjPIuj0wvPtGl0JkUkCHofcyj9Bxaa+d17v3SHYbFRdyLWsdeWiB0J
zHA0TCL7kHCnyt1P9vIxmHACHymBVb5mLtPNzogGYAycwbQOuVVmkhMHCv4gNL4e
XaN3SA9c53PZpcxgBhJuUplcvnhrZNkJU/bBqJUZRfJPk9qqEOlZWe+MxGdDry3T
/YhwuE+I2w4AYKgcB63aAaQgWwG+4G2nBc0l7N5LwkWFqLceNDYCNy2ZmHIX7d9T
8M0Emuwm4VR7Zil1lHBE6jOZCzXnCiUEL5td5wr9lWe7i6amkocnmD1CKYQ0JbBt
RtGgS1NH73ZSSrRZ4Q++88DSLSV+dSIdsTS8PqYXXyyamz6czatEi9YZGz1wjicM
TVu75cfuzs2guOqwLq9XugJ1upJVkKedKZuXjd2JDOvSRV8RfSykq4g9DGq2rOFQ
cBtlkmvu+DAhufDh6PhjvGeD6ysx86NcQ3qwDDj5hPue1vKNtUQDLc+utWCdEFaq
vIYpoy1crVU+ZRnHkI5hHeSN8ctVZVj1b5wiFByyurtfJ5UX+dZi+XmsDvCMfrBE
mnxljTMWli9NonDmYZWGdqFPwaEITMJEegCZ3AUMEbMZdq1egcyQKjJDibzjsykp
rw+NqXPDvD3ke6kRmhhMMCWdDTriIyldnRa0dhcovdgoevqiIuJWXAeoNNGbtfsU
U+7dUFmbBtuWJBl7YLcL2tbQD9WeGMSTWG5i0cYV+lfnJPNMtgiykvaeFPCBOwpU
CNcoVDs8WEH2Byk7n9R1VhaxpYE8AJml0/hU4ruH8aiJ2lrC2N+Si+yfvT2GixJZ
GTyRM4pS/uu/0oqWpOY6172pXEvhKz0s92LVF94M6LQpPYYEOfZsurZfNP1lwF3O
K+vVPvaPNERs8MLaareSUKr+S8ivj/MG3Uzr8yisCaTrbwDgk84S4Mmay4mgr7D7
JLadwyJPCtyTNEGguZK/pzNV4PT8CQGHh8ZfnrJMG3J+CNDuqJCjscvHZjmGTTvk
6oqIlmN+DYk1atxML2w+nPDdFsuwSm/8QLXIo502A0NpZeF9ZP0h8U/guf/DPUD6
f2UCjJdeDcIvSHyDjGAECCIWn6/KUmXjwboWj+HeH2KLD5onD5RYQbvkkf7evC3/
pcRuZUNWHKFTz1gbsoYtdESBz7gJppGaU1HrNmi3bJChYCED6LLaT9r+nbb4eOym
U67py+Zeh9rj59grNQ4x9Fr+fcAKLntSH6XOOFN3Eaf0qNIA+Oyrh4H2orWSJIAW
BQSh1ohdgEI1QxaxFlDHwnNoxXh0SdxDLateBOjXdpjeCsOhehsJOYb+xrjR2aHm
qEYONi+VEOvrM+cAADZVShyjz+AgBQEpNrrO9In0tqM2LcFQgeUy5gGWVncrXaAJ
/s97fvTHAjsdm+yRWAAPC1NitUYeHohpaTIWsGYBo5jcMKlFjFZQP6duV6+oQv+a
zPjCRY5nSXxZ9B7Sqp/vaGTZZmv8veLSHQz7BxVgRmARywIcCO8CA/din1nT1dCK
mSbcl6/gIJpg3WOAM870BdlgAgn4zVnQlzakUhk0X4Cw0wHWHSz0oy0yVoErAMqz
rgHmpBHdW8/yUIxeOXHGSRTAKdIMaXIYmtAEtQoQ+/zEHtHQD/GiXd3I4T2S8ubX
TlzV0YhddLRLZw7UkPJ2d3g35B9DFgIuZenRLg4KeOn5jdleSFU5UczZl7P8n5UQ
YSsZq/oh15j5mIK63/nXGRyn8gFvGrjtJvehO5BEjA4Nu7QDC5M0YjIDtBayT7Po
DaY+o21w1HCmUMpvgIditSMxzecgndXIh41aUcyZxg/eAmXz3p54stoxo4cywtE6
gTZIPkurgvjT6+aED9t8QIoLOESNmBaDVZxUZMwp7aQemoIBYwvZF3Ja/BPdeV0d
5DF1boRieHUj5hR2s+grGIF7hIW8AmBsyZKYj4joxa/z3O+BgIndQOZCB2A0QCr1
MCixJrw331EyszG6ntaWjVh8aCoKGC2FEepY2kvyPdyp03xJbefhIjAO2bJzADaR
Jk7UO6JEwI33hA1Ujy1N/TyU/Jd13PA190WStGJdaLhUobYVj5yNXIcj9HoLvUp5
5pFzVyPk2zSSBbQJ4rZy1WhbTax6lfmcosGmjDUk8m6w8tKUY8WZUjEvsCpZAmr7
LdhwdWbJwSGR6OfQfxr2AhthrfX/VwdT6RVmQIDboVwP3eHICxAXCVHt9RBx2CBd
Ruk6iUBt4NMK7d/C6ugB+vpHi5pzQc1HOTQrtcgTxVPpymcS+azOIwliBA1PUdq4
PvVoNRxyVj1VvXWtav7He+28z4sJVWH3WCNnrt0Fv3sFxAQqbkfD4deQ5F6NEyeq
3lzgTgbUgjedAWT69NZJ+XX71V4n1l5VDdLLYEr9bMrI9Ja6yoRRlQW4kV2Tlcrf
Jy4w9NY+HAECTBbVzvcKGHu03jqZEtNxGj/bftrfj0PdG2Bpe6AgZSjWi5l/BU//
4QuApWN1OZBsLVEvvwK6h88CqCgbHC8QC5yEqMCRg1PERLl/IzKy/2dFa3i//NVY
diNZDwAoWGT+BI8KXFq8I03ODsIRdv8A24k7mTZfd7BbsJ16D1NszPv338ZJjMph
hO2Cxi5q+LOzAmGt625M8A5E3+H5Rup2Qbd/KfSniK4CsXOKzaRCU8tNLNxdzYst
4wyago3Bod+TeDWoKp++qUhAGPxi222YkPSpPqu7AbsCS+jqOXMBT5bY10v/o8QV
fbUOX1t06DK9hEj3tw9spyUBAnBoiTx9fSy6iwd8iql0ZRvs7pR2DI5BTZW6pXUS
v/BfdlJQ+jW31lY3tGDlCQSBJSPuKhcyUZp8xuuRX3FeG2+XAnQeS+KJsj8vGd9w
5WR4j9VSm/YosZJIRjoMab7h1T13oFDmcJ9dDoZTySsJqnxJhaGdKrvTi6xtUQG9
CYWXT2d2y5HWZUO8xcsB37XB1FvtHXbHIx1alsKQ6Y5fZLVmDWCLz/C2loeIE/Pd
BXeKMrE3P5gAjSERpCn4UJh87uXJ5OMe77L+tmc4GDYZli5/ADVL/x9jRNiQkiKU
b4rcA7WJ0KyVOwtzWNre2N1XoIXA2ymyJnHLJxDrxEJ5uFKE7avpwDln6ftOyvRd
EvSMGUaNj/qCn1kPSxijRqpUsa2aRCVPHkazQey+ELSjZbjQUj3Ug/R4HPclYyy+
fN9B1l2PzMHp9SQ7h/o7GgQVjvFzxbuQcqITohQGJ+vdvrVl99L1T3tmOAyaDgkQ
19PRoK1Q6/KOEi8887RSK7MIGO8JtHKF4f7x76nmU7NEeCQ8BQvkwOyM+PJQkR+m
bxtx6LAJaS/cIO6EKLsM6MfTCd/umRsc0Jq+6e7DQhXh3t1fXUMvx0NwZpzeJYc2
Ppb8xUpzm65LlkN7qHHtmP97n4Z+1gG9kJgRnfsdWrJ8oFqzDhnsoO0hmGo6jZJz
gVruw+8Ci3QaHvQoWofcauHXVh+VhpgUsY/y/+bC/r/VTL2xfyqEywdtmcG3YipU
ecNWHOZ+8RzffWjD4A7E9wzO9Bq9P5bL2Yp+0yNW3OlNH/20W/p8tbzI+EZ5EZrP
q7vC0GuzAdSj2lSy0ym29RIFLY5YBuMbVADnaRF5QjlgxiHpONLigupW5NvKvHJL
F0HArX2BYIywzERD4ALshkmL4as54NcgV3GLrOqRdzGb+OwY9Yz4xbPY0R4pJQoQ
PEhYhyK+NFZuzsXqruFjbRoSYDkgGF2V0rMyvlbMxkjU27YeQVG0j1utlGEoYElc
w/dTlZfekbSZz41Q+e4deCr9T9msWsJBfNd6zaJCx3CSU9jbHG2lbd6fXf+aFiWe
5BFaWSbBu0pPVD5zNju9qYlFWMnzDdQ+1c0piDjGOEM=
`protect END_PROTECTED
