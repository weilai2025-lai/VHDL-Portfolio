`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cl35ph1TAV6UeN7l+th3CjjDvcRKkFUQIxsOEa/a1/XTben/EP2j/5aivPUjZTqp
dP2AU4+Bqx/X0KzP/2/DHOj8St8i1iq4eYswaYPrxAVYPFUcHxJn852Ftlii3ONR
he07iTDaVVn08emyHv/s033dPzvTSME2Np5adYjD/nlyNA1JJmibr0oSybQ9rggg
U09Jfj07QjJ0arlBm0Z4BNLGQy+rAywXjrAo77ys+XV+qKJtk+p31/mB/Yp++ZWz
qmftUnBZyGlEkuLT01z+vOn5UqbjHz/tUBOEeFYgk30RdG7eXZGua5/PlNNCQ85w
K7L5ZJ0O5Jl5FG7Vq2qqvv/7B1s1EvehGZw7BPZ2qLcSpHam5Mv/7B9drf39W6AU
Q3ktWucmF1QBjiTgo2jBRinwuXdmhX+52FRb9f3+q1v1ZJGVrqFqOLTtt9yR+gBF
Li/bdk3HGxySSfjXTd1FIspfRKlz8uwhm+78kmM5nyi1tDa7SA6q3S0rtMPt6ocr
4eqT5q525DQyOP7oNMb0KPM1/cu97aP1xhdmAnPJk2Zs4n0E21O5ayYpL4bZWINm
9qXip0n0/BNXwANAjEPvIt9EqEh5Ps/GHHDQiMGP/RXaeaRq2w74x/fThEDeV6A6
R+cCIW0PEIuSftPkGz0BAO2k6R7BETklVKUU0vU1mgEnXS0r3wMyKnSydSadQziN
unqL/cUDt5CdEdGueT1JnYjPJQnjhkC5RYjJT6O4RAfq3nLRERFiR11tVChUJMC+
vhKBFKMtSfZ9oYbIS2YUiiLZTH1PaYDHmNUnao9qMKPvTGgx+XTdsaPDuAhKHgc8
uX2+pr7koQJ4IY4Zz6c7YFvawnGYFDEvXUdUX9yt/tWiJ2OcFAfs9lxf3ZtooOdX
CQt1FEG/SZUxO8h1zX+jVxfZhh5QH2uTt7P/7y+C38d9wnM+Pes2FbmAwlsDl+A2
lcCJ1smZUSYjVv/8d5N/nNBe3nw7bRa9Qi1MrT305vNif9s9JJuhLpV6HKG/QS8C
hqGuEWxjY9zI3ayycb8h78Uo0UGs6kduzvLVarSnVkXiXobbP+DOsCI0IL1Ygll+
UQUCaVaiDPU/aATf5OjFkMSnSjbx22ZzXyfU/FHXiM3ltP8f2mKLqtMmIjLc7E02
Q/ro5sF2WJHkUeqvhb08Q8s/Nv71y2N31QPc5sEEBFauToFp87wiLI1gA89XILQl
KUBfDO8lwqN048w6gvbyZ/VzIYVObgLEyXBhfErrVxSeFbOuBUhzoMwxLvwuJNPd
jAJ9G7uUtZ4HTiZXCCIrocoMtNlOAxBX3yV7CEi85tIVyNyhggHO5+0L5fIKABDI
F3S3+eFUAZHBdPe0mny100v+K8Jx489SWRYK1sE9yZAvjcfiTqAjFEeaNzAdAq7h
7eC7sctMbLYK+9AbWc1/TpXumv3Ogrk/G74ihIYpQ7jq+hreQvbiaPb7eQ7N1ucs
Y4Ggbgj0RnDdE5LPrTQ+LRUvrxG/Gzlr+2N9zd+Omko73GDqEcE9Kl3ywSuuwXqc
CmhqBABgezzNNSY0ew8B5taBt87VheigxI8nqcrexhgNre7L9V14DCbqvbM4Wy2B
rAwcfYNAEE/yfgJQUssJXny0+3k5Bo4AauDpJwmzEiu2yuCkoDUX2YebuAHvkWfH
S1d2KoDQfXGhcfX9FzZ9wdEP8lRUW8IEzKiNvYPkIYkUSRKTDCqCB8Gy8o7TvyPd
P50OaaAp9chvUOu99li3rfjiGXYcmxiEMeZz3FZRg4rkAmxtvlrFMNERjfmRtVVL
V53425bHVlXofL72vjytRIy/hnl7GWwIWSa8qfMf79YtzAvkK6UFUyReY3TKce1+
UoKk8p430XThSspFlQZl7DL5G1BSLs8auSI4Iznzs+jpHMgbTjWhbfs0/S5qUNE9
/5OCaKf1c0U3jqUhGK3Yj5ncPMTAeyg3piYFzSRvx+UZsyvlVEPDcD2SjHNN5VLL
OOQYsf9JlS4MfTrmB17VE520PAJ1wpQsvtAkMbSxPJWboDPWzh41zCvxUlKXTSbc
oHGp8CYYAoKcy0opJMIDci3axeVa0h2i8hpZ8pldGR2kgjqOlDOubqzGr1l5KHoE
jENt8Uimv0byG2z0eZBVVjr7GNfE8hjKUgmew1xEsKf2MugHz0Uu4C97GUurj4Si
H1MwrNYLG8pGiAw6vDqlqGXLkyEA8dbeRXYHFNUuq979R3yIiqfe73MnD4UMqllw
RcjUneYiZ/yO3LyyaWHhsx/JZIsSaM+kdUoi6VSvXt4RB58CMO+Kvcdx2CVE1GBO
RXqgy4AC/klykk00J5F/MfmdH9TxRBX3wiM1AJ+5pr+N8cTHuNU1Vbw4nxBhInjf
LxoDDH3oleTf094562pz+l9wFN6pVuM3ualQkFv0lEd6dBHVk4ZU5NbpOFosHqhd
AeEhaF5YYF2lfsUO32TLkHgfd1Oj6Wy8ODUf5f6Z9I5pcabZmrWNFyoAMBUedP2h
ZgSr90GI53ujt1lAFfoBv8zIFIyCqrD/huQwco2ABMEbWz5NPcPAQrekWVM4rjk8
Ip60xCfJX9Hv8yAlW6BuudX2aiwnS/5+lD+U8mS/Wjdr2iuXfkM5pZff9KyLk3AS
EVGsvxMPhERhN82d4Wf6CI5WoB5QG13+BvA4Xy2mkt2PovtKK6weHMhmvxRvvtNO
ZJoj6dly+LlkRHnaAN4fCLbbP5jL1Ys8JfYt8rr+clYi26tnHeRjeMFaR6DzcJ4J
RL2ZdAXaauE8U2wf3XgF3qKlea5i8iD39bj67rh9xezBwPoB3mU+jE/MWNz+Do9W
EFIhvF9Y/ulpG+7xVvvjxdlkGxqgZcR5vmNCLyv3N/uhW3e1RxrgoAyKVOHIYCqZ
D02q6vYBipqabE8D9ZMk6R4krzMdHq12dwWAMBH8mPm5TAyjUD8wO3SNlMm4U9MT
hbUCNLphiii7jMPk/Q04DqrOSUg1v74y/g6A4R1w3BszxsfaiiFzhV71IvRHeIHw
m5m+fsU0TpuJTc6Oy6G93U3V34CSLUafF/cYd6ygTFTw/W6pgTXeLhlvxhWWkYR8
Jrgwpq6Sbrzwy4IxGRpIOnkhw4Rbpw8QKcCsM/0wmYsrqSTrWVrQzOkif5S/dc2J
sRUvWFTnRz+anXezDrgkgeGsDDsBxFS+O1uwubNNP1pvERvOXLaUFTNTNS4nsin1
u+mcnCEIXMnDeUaSPMlQ5+oOWYlWw17Kn+dnefnd3YRw9R4Ee7TNMZMRUjDIUc2k
aTUY3S88Gq4mzP1Stvrks8kYtkJqaMA2Z7S1QgLrM3CBk+GjhN4xUgDEVWkkgr35
/lkcO9EYRhEPzM/hthQWLOZ/l8nKJ+XdT4biT4aSnR62Y5KxFpMLmZz+RsYcwz+V
Qu2XfUrumECYsjmSBS2chF0ABhuwnfyg5UJsxX5aDj0sh7Iv74X3c4BYrvRn2Rjb
X49yh6Yo+K1iMJAvhvRo//dviBs2zyHmxOWIdui339Vdd3UW34nuzGEYRXAOjdXN
UI500ht6A3jMGlOtrKX5jh2zEOrEoJzTydG5r393RXuZcCkGtmAGCAZX2lxwUyZF
v0GoZz67a0aQt4n3y9KmQBu4q0ggerMMKEml/5NRfbRH7+bjtJYDxFoMPwuTqSb8
+da+uTxjotR7In9u8VWOytsgaj4yse11fzN/SoHhuojrhdgLalx2gCImwIo7pAqZ
hs679s1guG+NGVoDX9VE/qISHZRLcVL95i4/rabfYBWeZfxmwYlj3kcNMfsyouPA
B5QAge9C4I8NkO4EK/l5DTfIx4RpnydnSN3ERc+WUVRPCiQ50F0DyAn9jHeY5mSx
F4CVcZ0hL3bX29DudNGv3Ys/inkAID3V1u/d6Bkh/iXgbFmyU3yQlNOOT7lEmY5e
0W4fYTWbFgyswVFQFdhd7jmWqxGlkF6LwzTcSwLZFepX/E6h6POJP4BPvl5XaXrf
po1FBsyycTouSzCQtOU76uYxGBUg3ANbvqZMkuH1nvtE0zMeOvvbkBRajaK7wJ5C
opNQchmvQvL1C2gzzdbfsTc05JSBAzHsO3yAU3mRUdOYLLpyIF9OVvyiwnJCk9wv
hX6Gfv+YKnIkCMtgQ329ulmfIg2gCwmh6mvVKwSIp46FFgxAGx4V6MM7tDBF86p1
Vdql/4EO/DNP+c7QsqMeHLVHErwO5gkL1t80wlmjJu0b+PjKNumqR/w7iYMUU4Ei
zvbXkrq0fSK4SzCNDAcr5YfwpUvuwouPBYW3+ZfAxoH84Z2na+kq7xz1ObQEbw+d
CQheqX8iysggXQM6Llqf4J2Yvxd43wJdmc1hiPK289alC1c/yWyZKZyJRsTPPqKm
A/TVuhNn2rD0Y0xcU2YJF3wTTLxI203nMm/szFODLMN4xCdmUjK502UkXkEA3awb
wLma3lCGzLwI7NqQ8MJ3NkOlSomN9rcFfcq7UnsQgPHnvJ27bpTpUxYgN47bLtOB
1639FuqyyPg7qygS+SW1VrXAc5sQgB371aVA/zezNI+AISSQnetVkIdL53hdi2bc
CIUuvEcEEGJ1of3NDgB4izs8GBTNhfm2/EUGJtz0qxrVGnlO26zz5sW+o5yjm6CG
+c6Cj6qD3f4LIEOETR0XfZB6NZAINLh7ZxXr5MBX/wc1o/FiCsgpaMfUkD9pifWq
aquWKrI2cjb5SPdTkv57xCgnPOjNt5ZkH2X3t2eLiIaCIRRZv+rqLHas3FmPqsrt
vZQsB10RuAYgYrBaypiY6wlmbNJBvBndbZS6jzwC2da86HmbKZYWUjd2Kz8O7/L9
H4Z3v63g1PsMHNswUpbNS09komQFJ9t1cFPVOv33dYwG3db9WpenGZqR4yy8YMfr
YZjZvU7f+tCxLPmWmM3GIsqX76g+VpP0r8twS7uzD/+mKO43JmBLDmdyvep0a8Q3
uYAMSsUVamTJWl9E0e+5khO9nFKklefTH10W6bnBwK7TzRNP1LUBxjHmOm4Hdf8O
6kHqsnGiMyhnOt+OqUvK8O+VUnNfeGP2heAI+F5qQE2bJ+UsXYVSgLL64iI86qoF
Dyki8gPQDNu9kPy+JaL3F6DkLNMRpM9gAfA/VMVJPHePT6XpnSgxhZZoBJ0RFcvl
7RKRJkeb8p6MrULBBE76iGKawBwCuK4QS+29JfBLS5qaVWbmfeoUW3/SgVbX+fGw
RKn3aSnCVgw1p2ygRbligdeFeXBDUcPzqNkhubad40fyw5YZBcOilxYYmSlxFmTZ
0jT4xaJtcKSjanWPRtceGhop+T5GhkBzCWwCKnj9KgnwGuMiklcyBCWFxcqS2e8A
lvLIbPy/fYHEbHGCudugzMhqVDTJEd5D0jimt21gM4rCZrooSsVaw/8YsNI41QqP
Z06tD9xBMRPc/PVJjwE1jO4jHVE9jHQ9OoxIOfEz/B990BHu3aTX3oSFePl38+1K
9lEyLFW8JTSa1YKzKTIW2M3erI8pMpcZ/U6jYctcKbs2PRFs+Jtoy4LuhANPcEZI
rzV6dR66MQL46a2BezJSHC2ymJoHIHTb7u5AfeJC/aAKVpu+KRbNj/Sws28PoRPD
g+c7pZIHlxMDJ8vSwaIgKl+MOs+zR3SFDM+b3LkwibKLfTgiMeeSGZaS14gEMLc0
8YpLKeZ94HYPocAK7fMiiw05g++5kkOUQmQivL5I30KsXZ8rIc1w9bdaUIpKCQaE
hvntDaNXoNwA5dyHNUOIbTGjRMinZz5I7dQCBZnpxuuTHA9hQRYJGl9sgbfLnOxz
FwPzxndNgNRHA2nvm/Hkkgc6eiEGenTyGTQaWSSGoGrGYnG8CyxVYxm3o4rJeb5y
rU5vvtzIyaC3WtTcoLVvLxvTb3p1OphqbnPzqpRgZouUfw61MoHv9go/0PU8CIoV
Gv0fMJop0DMDiYQA4Xwdvsn89R0f07riI5xlrtdo2LYfzIB4Hij7r62UZGfTYgCP
x6pOsjD5byGZSkELPIaq2bL8EQ9D+Ky7Yu0Je1eEpkdjWADSqV0LZOq2yjsHJfXN
fAGj8kyx6X6dt2oswW8vhNc1duRyO6mamktufQKM1uMx45k3Xi+UyzInKKA3VSQ8
4gS5u5c8OR/QpYYQPwfiXdGBe5qHkeeCiPS7zLbyuKsU/mBUinZqzEl/1kMycV/m
QYonVjoSIgOf9LCNmP30QVYBBo/z1QGJEBU9T0yOg1SK8CrKqytBDnN/GvmodtVS
Reuek9L7jhwfjJWP5PnUl7jbQd3efEImE5bArbrakIC4EzYSf7CTjs4WLGYqzy/q
DSB7DbO5tro/trNzVOegKGhmX4hRqF3TYRWx1ORH5EF2C9ZuM1HuWXhEIkAAWHJ2
GKGJFwVj2eoGwhS7+Q2eXWBTE3DdAhJJf+ElF2hXOMyKMrY0kM0iZTv3e6fi1kMf
3+RuOS82Vt6H1r6XYk48oLPwfKGm3wQXL4tlwsUSXrowyvlBjewep7wCETo6UJVr
pzTV775FUzWfXaCRsC8As+a5VG82/orgMhfIivlomlfJMl07cEjiBCtg6NYt6WV0
oD6NJO9vDQwZq73pNNnA8LdMO8lhwrtD9jsPvU4ukuFkyVFHpPxoldu4eHkD8g79
z2KU+AjDkVJkP9kw/+jF702EwE6lBpPemLbFkYuqFgbX9fKSt+3VvxdW+mr9k9bQ
bxaDGLCxGolHcpj2gnNw/SleNqLTY3jrgcY/uDALuxE62YCjsCOfeV1BsoJ0Ybl0
hRK6KA72IFAHMnu/VbD2mkyhghIX+SmcFG2OA5mEMAauVeQyu1kOEomcsyBWNrvk
2BCc9obVhSF9KT5lOVIBf7h81FeYZBi1bWftjCESF6G2mgGw1gMQXszHzH1uxDMB
u72H+T1/5pRxqUjLAD9IZQgbV5ZA75FNj2GDw89izcaFqQqd/gxs8feBEGM8QrKq
E8vu10Sl0hZCHW1y1sb2oiaOArK/1R4qTNS5b9xgmTiEbYzi4zVoErhMVa8U1q7W
g0eJxVujlx8DS/2DebLkuDsbDPztqFLMlQaeUeYt7/X7xV5TQgyhW6UWjATOig+w
vUus3t57nhmo1OReaiVyw7b+P3n4DiqexMFd2RkP+fB+CAx7q/iY8Ddny9JMwawK
NQmEWiFa5uy8mOF0nPwik5flsf3w2f8ft2sdmlLIv5esR8/dOfsE/xvPKS6Wwx2D
lrB10oSJgJmtGMGvHksp/2x7oj3CGKYWjZOOxeneC5QsqhYaaMYLEk8Bh15YbxXo
kN27yJkhL0UaekH2ecsBhBgGsSCJ98jyZtod5+Wj+HlQjaR6y9CvgucaOr7YlEB2
JZL36aKM4EcAXCx4p5YFxw==
`protect END_PROTECTED
