`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQYPvGCH9xNqTMedB2mVZl7HViuSqs//GtVAWdxLna8ce0VL2fI7iedxi0PDYjfc
S7azimEJWRoZADmk2Bulo21ZHr4p8ACnBz0kCqWjAOJEgllMpicjvzuZzvZsNnw/
eP9w/PhFHgoHTF04O8UGA8Uawl9ir7X6u1k5Iqlgyp8ogRyEN+RS0JcVmYj+4tpD
9boiWPKvH1BFmePhz/8OWReX9QaZGcb9bnJpWurMzA7zxiwCK8pn6ZUxg4jz0stQ
dQ+OA4VW9hkiOy58RuqQiblIi96FxmCvKAaktOT6wjpW0OBXZ0ZLjitzFaiXc7uk
wqXdyI7s8v1al+zfEu0f7HStFjkOt0YSlWAAUIwEzw7hTZT8mboLBTUxeCavWSpM
Rn5HsK4z7QP8Z2l71IJfF5Jh0Nl+ow86/y1s0WTfyE9xCMvU64VE5HK2qdTx2mud
j7gXG/cujiIh9S9FJtuJkCs1B1tUYgp00h6xng3ssnRqxiKC/WJDd4D6lt2Zm8hJ
DemMmmgSmTkXy3KhAVjhZadEWCxFENADfpQdtzZHzuFS5wAucsMsZjkLSRTvhVbK
aA6U/+3V70RYwCSOEre0wZEy0knwhFC8uT9V8OtCZWIbPceRWqzc99nWIBA+bmd2
2GDpikC1HHI1RdPOO4s7l0qc0geHDlB+pEmP7k0/YRELGDftDO7i2RkVbOLPvqPA
Vq2TMsGy1zp7rznvIaLL8uzEErbGGe9ReA8e1T7hSa7pr3fWvAM8dDRK0EzeCPPF
PzcJ0gj8HuETAOOPO5tsxRRUpKMkzS0F77dZn+CZKOuJ3Ha2Emchz9WW8ugAjqOz
P6Dr19KHGleKUnQSXuw04IS2YeF2Y4Cro0ThFbhs15irJcyQEr8Ji6wiENprCzSh
6YNsArmrm56ZUxYcYXxIAcbU8GspO36E8fPGPc0VOsvePP9YTCv3KGoUSxWEZIp3
BFLoXFGMKBYMpFPLCH2DwHQlfPcsEXJOz/VUWuYUhOoWvAVP/635wuTmZY9rSbe6
i4plFhdIksX8qLbDRQ+DmFhG03kA2rcdmsQlJihwteM/gmBxe7+UUULO4PYQcoG3
uB5HdnHHFdKcr5KNI+V48f86Xpc3adxwMc1+SFF+vG7nFNrbuJdhN03GdJKzpOhJ
xf1JIuTi9w0opvO4mPyU95blocmG9HSxi/nOpFKab7NqnONeobT2K6KY3Pi9Ww5b
ia9jV5VpbcI6i53OIF0oZAFEDdPrOowovMYpvD5raqM9kJIIq2PtxY71YvS1FYhy
4a3/bgPPZ21Tv61hDhvZcToVZxNDldCbCFcejYdzEu2MHRme+pAACzIl8/xjdQZq
/gTrQKWbmoqYlkVla1BOOpKRt7zwnxR9KmXgkrLmtpDnZEa7TINVp7tYqBE0hpfr
eXqakackqoWJwBxO7V6i/rK9l9RNJs//lCFTXOw79ZfJHub6SgLKmKkrZe10q0Ov
SZwSk4/oAP0SyyjH9ghhYRldiU89IX3BeEg850/qV18ZAIS88D4rwlyOlm0TPTV1
kue+eaSaI81A4frFH1/BOq6601tL4dYLtsQW1R4kRmeFo/h13wfavMVEaVrmQZmI
0KHJB3DOucjGb+Yg4tcDdGVoDo5cMLeil6OO4rhcrQf5r3Qg77uzmokhODRlwvZE
Yh5OXsJ6RDRfnd+13Tt+/6zubdMg6iHcXMOKwN3+3Mai6YWAQOffA2xBw7kL57qE
OOejEusMtSMMicXKDQTIJwqFDe4HQ93ujLn8H62MFmqljRy0Zq+zO51YK9xEVEpU
r8zKP18KIePvfGfj+QG354mLzVvxdCKfIywG95TMtGNmXDVlyOjvi4T5ZGvksJfL
1uEDcMM4ae4uLBU8I1sYoXfR4RsL5SIuKfNC/AUiZoFoVMEmpQgMokMJjns4mBKS
D2DNIu8UiGZIfJmjV2N/ob8yORZJDUHKcGOVlmJv1iO+0BTeQguqNfpufjfY/F4Y
QuSBC3hIPuaaszo2ngSnv/j04VJeS0idpzvxSvF0MdtDgfTtXilVYAnZnzkUV9qL
r8Hc1+AKsdhLm8Nm3SkCv49HLLqcJGPU8pRTpxw1tFTbZzVeshz6i84kqfJpVSho
6wK7TXozR5J13SOQfnTfJN7YQrQmTbAsmXmt+gQJ0TxsHnr9ys2HTX6/QOAjKFJA
GJLM9hpbI2+MFMkoZo1UYYP47GHP4FZMc7PWcgWqvkiwVEpdNHdj0WrmZEvCp7HM
oyCDWhutpVGc6tP4qAaGHR3ziWmUtkjTg1psst7RPhTraOIqMjUXOy3DuXmC8/Jp
P4fcdKGpMut8aOFVGd7NQ5FjQ77QH8wJJ39aB7xWtCpKOKXYLXktgMgbfCPbv/OD
zoDyUgFsU9dXJqn0d3Af2MAQ151mKQrPdxi3YfbPz8GmMABRhwStGcVpbRfy96Io
0xiwcNTE1rqGtGgDz5zIjpWsJxALxc6q9vCoBtPUPXz1jAnPLgwt3lsgjcZy4S5Z
2YovCwXOt4D4baoYQ5GILvU4pJoviuqV7szDREJI5UrLPWAbnRybXxBpNU+iYqGV
PQSCGouLM2ms6vPFFWtGQru094OztaYVQVY+Zzj+ltWDzg54X8wbHNlkbiCkJaaV
84bVXTd8mFVrN65ZJmPXopfiBTVEI6YEjy9uX9qpibC44uJ/n0iw4qCmYUvpHDW6
YJf+Y2paFbZERPLzYqpby5Da0Afxm5qm1DHI4uP3nSUxWLebbUnv1PTr7R4wkgK4
AH/YJOg7COupeYD184B6qXKGlqOHy4UWwRWUkZEDHKQuyfq9JB5OSDfRudbmmmG8
xLyOls8nEBJy2m9pJU4vzxMO4H++q4L7yQJatEIjl5Vj8n0c4ytOe9oxsK/QG+He
MXn/evtNb79gQsFlBFOi5OvghLaheYRsLYgIvdTvCL4iWTlJEWhsUmMvBiXZflHj
XzFGlLxUMJ5ZpbfCU2OQPicLnoPWEN7q+txwP/P05WWCdL7jRwtvunzl7ME5WJKk
DtTdp5WvCOirzaqZoscKKuYpg1UMpOBdZVre7w69zfPw8U4pGcV0TaEyNgSozYSp
0m0upnimBfnWkYKD1UW/oAtsOjvzFVRvit2Dp/J6tqQLmcLipU3fGxcQ8ksPTXMs
KfDLr/2pJEIaJ5q7kyYdhVYbx3oOkoWq77nDbhoJCTnrN4YDcYfkFa4ZjhLn/H2L
PpUsNb/LT9MmjhHMAm+KsTTOsEV7iGrCu8P+EVX1U3kjki3jy/WcGJBqee2GGUin
SFdUrSRP9iY45WhDnk8X4B6paklUXXe5Sj5fm2okQRPo1vvflwSc2FHybfQEpjnA
EmhSvrgBm4sf4NIfqPcVCZRty/8qeXKw8k5z3MXfilR3/0Vtm1f/ex00IGuDDAOK
nlCA51Dq9tPHrCX1vA60xYBPjH2TlMVvMKu0izwsbML6zhHUgIXrjATQKzNnOiHT
y96vgAvfSdhrpIx4kHtjL7/Xq2HV0+82mz+2Za3IOw+MIvN3QzO3J/0UurfNNQ68
A7Qx4cKTeEYKtNVv/72hMNvDX7ZT/f3bs7XlXHvCgFQ6esn2zK9S+WljbDklqHfK
52+emg4uq0LpayrJKh/P0LD2DIFPgdK9+seYHRCgXw9Ciz1KmvxFb3QkeaD7XiIv
hAsbtqP3E0p+dJLwTEtr3d4e3j0szOdR5RpjW4WKldJGAWQrsoUbKBs3bskg/2f9
5fLcFjkbWg86joulSWFB1g9TNRDB2YQv3BCaI8pyPxSSXaIwiPJkoPHdKW7LS0CD
jHp4kErpiYs/6MXlgjL4qKtueO0Rzwxdxn26TaRuqUhXs61vsDp8j5isPYjIr0EQ
bDQhOP+9cFMogwQwo0HrrYkpwUvLINxoVjS1ncSOi1mrOHtU/6NMRzXYzG3xQnjl
QtWMdBBRlF+2vbVPDW5jkXu1p+4/6fY2gOKYinvmHO7sQWP4WQMYC/riEKdo38ZQ
jNC4l0dVEtibbtiE4P9Yaa3IsdVIce3KxxWAea+j5iK6gbOmasTdONwQ9LuSRVDr
MLr8C9G8TbMgFVpfYKU1qaTyV+q2vXd9EXwkvfdTT5dzeq3wwKpx/w4ALTBhlUVk
lDBZx6VDmqbZXOrPFbux9l6XSxgrgRxF6qfevS12P5TRcKH9l8CNLSs+KYeRg3BH
pFKhhsHffz5ECODtyi6HDeSadkP4Y2f4rUeaoZH30dV+oh1QeUQ324+U2Ri4L5p8
A4XLOILOxyc/QsPl7Zx3J+SN6B8Jw28C6fQ1PuhcjfAPEpE4B/L/yaG0effyHfK1
toGXNxgRaUOtQYesAW/n4Gic052ZMg85MfF90a1ark61jxfZvO2M5PLnTCCLdhM5
yHsS0875+gaIcGhPdu/KQGBJ8gQ5fwStZ9Bjnlk7a5tbhopsApVfmv/Hg0yvfZc5
7epp/nLT5PXsIfww5WAqNNOql9M0kGJvbAZL8rx6CLnXcSqw2LDdag1b8Q8uHHx4
2FNaSJfz/0KY2N4Zi6CttM/TDi6F7ifFF10sNakkqTdV/D8u0H6XeBXaX3Gx/I9L
aqFgd7n4w6Ex4ObNl5Js88+irjxGEm3EO7STm1V/nXuJ7vm7Q70tZ7I+2Y9IeSKZ
c8LN/9ZH49dPcgOABB02c1+nfjfPanE/VdEJKDqoT0CcL91uV7u+SP/smZicVmCC
Qh2gYy14m3BZ5UkACYMQ9NQQPTwwAYKDW8ovw7OkvWsgzRn6p6/ocP8drm/J/bG2
ovHItCOR0cbTX/+ydQl8etRgfFD2yvKptIIr9rtyOqAOcWV0w4USu5U6ISmex2qT
kwjwHuAfseCGPzoafWn1DA4rD/ytbTpeAmfPGeJ3TsjY5BnCQu8QnS90QiXeME17
k87K7IanaTpCkBUxNkTlhEeu+Sf1huI/BQc/MYaJAt4fcZMfwQWLSDhBBIHe3UxS
xGshZ8fEunUUbvNBzDm5zUeMIf3b2czbbkBrr680KCnGsSKUg5KjFD8qK6RoKOQH
EA8C32QE+Fl05YPTf0RvglNqwyxgIRo3HT8QKSwYuvjMucexng6EtI6EYfsAd3gE
sugymvV6kwzoTbDSWdGuuV5kblT7bdfYzSnRBOV2NW8Blr17kMJj65b5R2uXdPZd
fUvOG/ynwoNj9UiCrbQUuo1bkSlmwytTOZ3aLJOGZLtSSDZu64lmBWV92cIAhyMC
gUZlJQ42ozSJIOgt0HNSCVr2uSCfAyFODTxONtWzMmsjd2GdhQC7uxDjZ02TdWxI
8xhQk+UqBfm5sKDKZY0ToMC3hdbVfBy0bP+rFBg5KD2SKIY/X2ea4pIhFFCD9Mn3
56a/XE9HmWaSUEsPVMHKLZDPY7W7bPKtX+6n2YLOBecpixg6jsHeDPAVxDh6L9O2
5IUEBxrskaW1PbfkTspWoac4/8gXaqdlw5PehKVbSXbMkgvB73oOVrl3omEGLtsA
jW7pOJviltiQN1bR4KYk/s8gV++TQoH/H6fdG83xWuVkkxTTnHgu8oDmPq7a8M1X
sVVuyrDe7xJzl6gBVpSTniKRN9iBAHLPRWsoFxoQCJkXEXHFqJmm/8UCj8X3ne+j
OqGLEpZjla02AB7aPsu92qtlVlXTGXROrdGbWZ5dGgGxjMGYnzNVf3IiQFpO4Wsd
i52LDU1BWCWPSPJJHg+7vI/V1qxyjNvv8ZMA5Q5Hh9Ww8E/AADeuX7wN2EFRprGz
+9nA7tG2OankQ6Tz7cfZa4Q4vQ0SxhPxyD4o76nEwpga7MzLGceoB2mIEKcg3OKB
ndEfD1k4t2KvdcYxQ4NGL1ptcaJbCqNLGmTAqufZB5P4XLhEnPjhXcKO0r/v5CP1
s4F1wPX7pK5ys96lT280EltLqrVMUIPhiJo6VPTW+DjWkht7FhNsiH6Q/i5JZdZm
jkTPK6j85xHTsUjIdQhGyZzsdKz1ddVoK1cUTp2CvXlsaumisRMH2hjUDse48vsk
k+JDzYCbsO8M6htJ5+NTHnPpGIGg7+cBg/6mqjCI82D6X5xT/W6G/3SlWEVDu9qX
8WzhloI4CbdjS97q3ranJXpOfv8f4JN4oXrGW20oN5uOQWyN+foIAVEiTn2XeEZS
KfO2ilMC4XLbDt7Py6DcyJbaXi54HJl+Wrf5aJQV6wds56ttW4SpwVJyppe8cbd/
3I0aVBhl7GJwFmtc//JCj7d0/l4ntbo3dYZeX0zSL4F4rLwQmn+rJFRE3BvuLU2h
Czr7Bcv6iFQSSqegrsA1yy/tneOLwlmbJWqwR3dNZG43VfdjT1ABnjlVV1FYt5eQ
Nekr1X3Ps3tsJyemRo5/NLRjspqGKuqwkttW68mbTN399CDx4SrKoNzwD5m/3xx3
5rDqlu9/iH9jJKyDEGT0iFSmmAzIBGyLGOE0Zidkhbvwt5WdaOAxAbVq4RKvNS7C
KYoEIDeDT7Ul+fmomHwyBfX26W7pz42f+ic3FWMGY4bbVB9Fac0o9WzbytXH9tNf
/UrES+K+Ud3tbS7gtjAt63MVuJAZ2rZZe3mDIEd9+vpXrFwuA1qKSWAUvfrClTlb
e+AhtlOQpB8hufcqVllseHHXdQ+HRiO/OZ4ScZ7/9fX6HLZmGi2CYJ0nZ/m6Ljjf
6XrOqOP9/158xm9dVXzys+TAyD/MtTCxi4WC8NGbJXd728u2svTTf66IViQqZ+Gs
ZdkuecWG8q/nRSq8YgBDno9yXaSctdh4kJDtWD5NpLx7iQbeFlmR7hMCsUNwa9eL
iNLXDDzihWF4sNzK0BJD/54QuVpWdDBJ0iK9aXId2lIEPSocPYM1Vbd/7a9UWDqW
Dqdz+PaoBrarYgCswIB1oR7Y2nwJYrBR8Y0HXYKAspZXRabB6VO2UqoU7w2mLr0o
YD0kson4+ImZHUFKwuPiTA47QmcrlN/gIT8UFadbKwpgW8XooHwTM3oBZ2UQKPw9
0GqnQ4ahpdBVLOgx/MfYCaUUzLaciTwHoL+6xZUVn+WknLSjIzMZLKWSvhJMwF32
eGfZKq3mI6Q8uIyAulHzByQ5G70kAwsOsa8RJ3wlUeTNYyFinWXjvpNLO3O1l6Gf
Azfg0d3uza4ZUpRkoms73d5lvZh1Zyw6Q2NJyj/XafOboZEu8KMyzQajvqGqgt7K
g6SQyr/XZ71GIVuoYGc3FRXEyWtrhFAjOWebADPRnm5sSnyAoQa1DNBsqsg/01Bm
NesTXGV2wum9kGZLLKQ+cuWO7/LF5oB5ZQA6PaUljfvsvmBJ0SOiTwgDwAysR5cR
5ZbXswZNnvILm1QPN6jE26SVuV2/zktMu3PppKL6J87SKB0n922H8mGnnZfc6wsi
Fmp5+J/FCXoWtu/Kx4RWEm1VxgLrMjiZEDNfNzlTJSkMtC8NXsDYNCQQTbTtcbVK
kg1yqTttYda3ObL+EKfRmlMyA1VZP4GrBN2yQ5m/M3OaRbiOA7XAeEeFTUG3g2wJ
RiztD953tIVxn0uV0BvN/UqiUPJ25Is6W/UB2ENkpSWlcarrj4Dls3EvomGaULtG
MHpzJ8dZqt3EOjbNlgXkoWDnMunsY0Y7yve76DOrYh55xXs0ylbg5EHESbrLCaiy
uO6HLmMq0Q8mivLciyN5qCyOpbbkOIu6mqq7j5VS3UOPzTbcqNpQoShyb6U2Ons0
UbUEC4BbkAONETf/pJm2V0VvBA/OdjvqGhyeBEXxSlDIqQpUYVcjLQya5OPonGsX
fj3rdSGdkHbQXcsX4pL4l6Sz8PWx3PTBIUKyYsAZZ+iMDZc6HHOXGxMesZ3klgvd
nE33q4jfAc3GdMXPTXyfwRa1Yr0HxqNrApoKpfzo4MdJe80eB3BY3Zasr4bz5anv
3Kc5DQ3XloZ8zbL2xjgg9m4hPA5Z31j1bVsAMZpPjJuY1wGZzFMDXENQWlcKgtIv
KMJLmMVvOw4UucAGeyQVO7QcISfoj/sF44M4yExf0RZbY3I2CPwk8/dqz7wBjM3Z
hMZdv9htR9u4ct+jvXG9T4bAgFaukUw44bUeZ+duYZmyRs6wk80X+BIc0hg38M56
x+YPVFras8CdoUC+2WDAwAf7kLU/eYSo9D8oTcU0LlCLzAPw5vLWr1pMTzHKvgxn
uWIGv7vbLFTQYN3HWwHNWUK0zjTGHOyUWXwQNWXIwPzDaiWFssEUYlfs88l+eRjr
c3mVf31ju5Dw3zi2CME8bL3PFadrX+4S/QoeBETo+7PUmFYeu4FrE9b0Oxr19Xtq
LLqX7EQGOvswS7Xp55EliFt5RxefsLBZljXEU7RYrv/g82iM2gr1w10LOYFn3i5X
Hgt9esNrkCDii/a17puavxBEvKXR3IOS/QotSC/sDoIZFiR6ws8f7ry3CmS3UgLM
OqZ2lNhLFYOxefgfAffhsrrZXm8bh7SANaVji4S9//CJh4oO9Kecr7BKFgAbzTR4
uoStVXSC7o7+zb4lj/P29kLS+0IRB6ep5eWNckZHVtq28fFyF5J/hvcC7+UU/K2y
fKbjrQCF5AztMYzHp8k9ZQ7Hr+iTwZZ1R3BA2iFVCDHoibdIrYLrFpBBJdZLw8ME
e4ANlemRn7DosJOKbKlI1SEtA69WEujqED/U4/t4BspgYASCUnL5+5j303sWRfR8
jwgcnmKOTTM5sLq2RQ+nimY2LUWvjO9HejhrcFUXLDlYOL5lhiP91SWbg3yPfdWQ
Tx2wkLa67/bk34HGlgcvH459kB1KM/Z2eWd5lqQoD8tl+xhlbddFqou6kqOaKkhK
RznKTU3at4Hvz7YKnm19hXIT1J/ICW7aKfqavt6my8KbLTeNt9bPJ4Pa0h1p6Pfk
ZfGReMeBZmk+VqwG7IqOlFrhrclQL0f+ILA0VGYURiBljzSsJRtwRIQrsvNYI/0+
V3fATY8jHoKEbvpUfAkf4BmdhLFNJkeI9kgl1pMRpB067OoRxfN7MIeLx1l5NSXy
zlUfzsKcvFcnCTIL4Rl2jLDCc8blpzKall9QumR+YaDuy68udzuNPdNZRK9zYrVe
D/9nMxkun0zU9BsfL9ScUeIqp5n+v2kUBUpolGKZ23MdKr7RI2n6erLjGeiG8zjP
OvNuOXvOg/ITtM0w4XbWvawUQ5x33oWqkH+Ec+QjaBdAirJnO18pkySZ4T5rQg9c
ppFZ1tyvC89M5skHHF4/vVRnQKe4FPQAI6mVV3J2D1eh4bEWppSphWoT3Z17CG7A
rXT/BU/zzpULTpoAljw+9blq0liklPbW6e6r7uPRsFFUa8qwIlZaa0dsKmkC3j3J
38JRAZV4DZBRpfgQSu4u3BhsreGFwWfZaI0WpLtkgn7/RD1L1iQ/wqcc/vh2VqoV
KnKgVJSRZ+X2IAstURIljvAaCYUo1sWmMpbk1KLnestNYhu/Q7aQyd4jilkaaU9N
53I0bY3uFxgUtg7llLKkWU6YNorZ5DEsFwsdef99W1mN2ixOyhvYu4c/CP5n+3Bz
AmrN46WQLfZk7eGtPkBChwgYDXVeq4GTeUsVljSiFusghJjLFntH0XJXU1F2XJXW
1oT8Y/GcZUezN9Gi9AZVPX368tkD6Lkx0fzkzDgqobkcmA0DSsd0yCymihl1kLIE
spnQ11wXZ/OwIMvgdz9c2UFhlOAyEei2SjxDSlWIFHP3RiKJBJ4FVKCZ9ot6DyFD
nLvk4ZTJD4tPAhejn5WsPGpg8g3sPP/yampxaBsdZcLEEzJaHfVbrfxIeJvT6U2f
k8JcHb4lMXuXRRn4lDKN6pFdFdirAgp9EztOYu081j/WjqbbzLmZptSoTJtEEz/G
Ti9fZ2ShJj0uIyTuqw9UYBr2sI+9e9m93Ma2hL2l14sbVuD3OastS4JHujaScP9k
jtv3ByGLeE0svL3WFLxYsClFoWqGPnHAzZFNLmPr6iS92fK523g1Wp8TMAe+8wT9
qiybPPWnW0MEJRqNuOGbMj9VWlQdY+yo2NVusL1MY3qtsLBYPvYb2ai77AOIr7g+
sFGEUMqkdkO1x1qhhp2Ryx0I5UjMQGpetLbSRCNA2tcVIJs+3hAGdqVcGngyGpQw
2JQqw8oMygqBsH06/s0nSjwlLoHpcw6gUOXAYHZL4VukErhnLgRpL139EtNNr2a1
tg661tm+TBJfwq2tPs/CjtBdpAr2dngU28ozdZ3rypvIG1X1OY0mul4umrbUIY74
OpUj4gGs89g9n5A6X5zVbHD0vo69ASceRdsol01lb2nTgQ/r1Rd4ZmE5WpcQ2vb5
YXQtnpHNx2RtDs3mTKWlCZ+zhryHQUHYQjmApBbBXhqTnJuo3fNogsUVoX2dY1gq
jo0lcbyRElo6VUYW7AeZP5FEl+Uv/e6AZNUWRdRQbfEKbT10kw4myQoR+yFaXMdA
cKqFXmEaoPKpfFZfwOR6qWtRCsHNWkaXJzVGgxiX+U8Zh/bkdS5dp2BXshTheF1k
FTkPWLZQ67LY74UMgYN6oYlffx9SKVp7tVp0ZsdmkwZidMRWhMNRvtwonCw19izS
lLmwm790O/s5jVHQD8+kPH21OV6CIWD46A+a2MwMJyKQnnZNXpM0j9C/WBQUMdtv
Mc1dFqCIpuu52TKAnGE73KXLb+oAk4ixSaFSDhe6GSDveoWSeJ2SW4974AnTBb9Z
oc+ckUd/XJnQPyjNqbQrPIwEtn4YmWnDt+K9APjGyA+Rvg4Oz9Mgc1+UUHsoK1+t
A+QyHAQwTgIDfURlY20/h5FN6LjowKehw6pX46bNFBuVLY6aR3k0+uvTY22NoKsu
G2pxTsp2nwd+P2W2RYf6uo0NMwUkvvwRyXLXm3qJmwbRzOo8yGPNVKmSNsIaHdVx
XZeK9ql+vbq6v9b9A4Fe0Q1Fa5DkKv+5xqDBdCpUMcn4owDAT7wqf4m+9OTz/ZD2
n+kQ3ZfHvC7fFpXbT9lBwioKInyYzi0+jRjV6jkwFLUX9oHTypVRskpfzJlmV9xf
Pfteu0o3QzKSmQzhVDKMHHDsGf2hYACIOtqMPBIZokqPz01DqOLO+OUeYalsCnL3
eJLh5UtsNE4VOxi9RVPlS4hr7swxQ3iUN3nIgH8SJ2go4fWJ2v4U5P1aMNNvy56J
jWDNvbTmtbPNgn+fwT1imrIcSUX4bEOAjlyBFEKVJ6t2OYajMJFI2OgMVhW45TwR
XKNmkRDAOXkWnlUG1i0m3LU9fFiOZvEncjps0IWNaFyQnRoU+G0MEWC7eSLwPa0L
SEF4ZRx/6CNWxrrTvZFPMltt0TrnE6Qvjo+BYbe0opCL8YSHMOKYWjVXKOaqy5tr
P4SE+j/6UjW3Wf0TP/FRBte5jX0/j+RMaqGX8cs5gbnC4dlKhB7fO0W4LI45mi6R
pouXklteaRFcrTg4T4O/3zJv8ErlpiF8r2rj1jSYEos+HXlJGigPTCxSNaKc//T/
fmmpyABbFfDHjUiHzIqzt3PMohR9kIVcw8TwbY42YKPCCB6Yfq610elTQOmpE1XU
TWes68GIv81Twj+Su19FQWPCThslDKSbcGMDH46nHUpbCFhG2+MYTTJvTqc0GfOa
8c0ijlkmVRl/pE6IXe+7fFvfmUTFRgJNm9owVKXlKlUfg10iANRhSMzPIVkjtOiC
MrRSMpmYUgv/zwqCAK6xWx1X5QWkpSkWOXJNKtRrssKm6eAFeuNphGbyKlDsHY3j
G2rxOIYaTdc513OLPeNTkM1Ubn3yHpeRHB300ADMHYSbaNG0wVtbgKAdajmdKqoo
6AExW1IX5s/0dG/Vi0cJ4ic7SOrTZPsON91iCF+hfuhDs0fbGwCjXZUzfaScoTH0
bBbOp3he4c4Seot3sXcUfDPSQLdOVQ63veD3P23aQyaAkFnidOd640Bu2J/ZQqD0
Uffzh2AYk7th6ye4/15O99DrwovuB4Bh+N4D0/fW3aTLNLimL2/qgvrCbzXEC47h
qPCyc2zzAOZdQO47B1i36uAESyDkUvGs8kP5LGlAsV/x3NNKbXjbVyO16+4liq3f
nreKfEEZfC0YTf2F0pa8XrDgOq78GjI04ytBtL+peE5coC8R/+wrzun91HHsiqhh
6nOd7IO3IqRRoSjMK0RK/g7fHe+GsFlRWD9gUjHPlVLOzEAHSWB16/uA9eG/ZzQq
OflJ64No6vPKnvJUVceJtMIjhtQVA+DgHuklEOAedNpQcmvx4rucKbmqfBgKK3pB
lYATW7zCc8BJk3hVOflbzq0jbyQ4EXjj0UhX5F9q8HxLiI0GwLZoGUKfYWxHKr+8
Og804993xvZnyfrxuw/Tpo8Y5TqeBWrtDqp22ResTFqEYTRxA1jyVb2zfGbqrOkN
4Xlh1j0WEap2zFi70OrX/eqZ/j3AgjbVPRWzax/f9G53Ssi4mhNP5itJvGHhxwgF
/MBo74kYydvYjUaEsZWk2F31xjvlP3pnIKSSweQJro4hfORZcU4Hq+QAsRH1bS3F
RPIGZWwSvodIbdUMfK0aOAXhKfrAgfyZ4ogX6zTOe3b5LPy37E+01X++/gTnPxEb
b1unBGdf1PA0rVwE2IP5JZtrsMlkZGPicNmkLDaFewDB9vbvKkQjuLLYf4GzczpF
mt8XWSdAU75bT5NGpoOS+A+cJsLz6Yb4xYCzFrdZ3bWRa1N/yfRXN5u/aJMBMqGO
I3BlC9enWyT6/OLOHn7Q0eqG5yiFvyaP8ZTiR4qVwLKSYlcuXwSc792lchbC3ILU
UxslZmyTDqpoykYA9GUf4szg6DkfYEHTAFX6S05QHtw+zAfMRx0NVImz3Q6H+i8w
QQrT7CgdZKd3JFrDor071Q==
`protect END_PROTECTED
