`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bPv/w7nFLgMKceQBfAiif+shyZJTK43rEHLYoUK4Z89sUgFUPH1GDWWI3cSh/Ici
iNJCv5dFZv8nv30f3i5gSj4PAkkuV1YAr3uyg/pfROQmHMQLbZN5UZPurGvqAT20
DzlrrfezX1p9PDH1Kw9UvJ8j+gl1Pp7Wg3xgN41z3DJjm6s5Pi10k5Lohs5o1yH6
ujs3WXQsbWvkbvkXn6Drq+d45cjgh0uw8az9+4w7PqX7buYe+pYQKfwnAfWYba48
oeWcHzIDEq31AKlMFUaJisqA3aJCKeIuiYRDfQ6Brm5rh0TSuLsJ5pirai/VK56h
UxDiGvqByml0LMbRZTKTFhr7XOTz0cvOwpuKnxnSpZuWsyM+2XSnC8ESYK/CJObI
0ZXp9ZJQ9kSs9ws0gIVj5XYI4kzs/RECKVmpjtAmj/6EEYt8ZXPuuF5FSuk+JznH
eodyhkiBVIiYRwcisRCPVkX94fKhsrECb/Y8jt/Sqj8uZytBfQdnfJUo/iRHbY2X
pYHsaekuMi+DLEYphBvR0kSZcFzA+AAxdlFUqUC/AAmCIIX8QA+bciVOw2ax4u4l
VclAzGxyZG2xTiU/CTl1XNaq7hBVYrAjzrZlymjU6QC6wY7gWqegJESsSqCKa1s2
MlzmwYMPlJ21WYHoX7eT3IaDHWQ70IzdbN/zyMxtaiIobAoDlZYOUpic4MKUBBl/
4z3gsH155IO7EttzbkyR5NypiM5NRvFT5LZL0dNseIhoY0RufuXoie3fVX16IFZL
KGwEf3dFMFfMDbxlY4Wy0dwFP5GXIjWumv7Z9PzaLegW5bJMqDMkV8QXoDWXJOPL
XhJOCV7OoyL5kf4S2vlhNSgODrjgGx0548XVBV4YeztTmC1A2tUHq3E4NmG/Fm90
Ac713JwlUYcjR5483zA7rSsEtoZApYl9jeeNaZWUOQDHKw/0IUD2E146AZJ0O5Px
tsYFLaVhszKH3I4yG3Mxv+EjT9ugxoF2fGxMDV8jgptut69e0krSqLLVawVdhH9D
Evsz8enizjLqbpNPezrx0VTaHzkzpbKisG6fLpiYUZpIRAWiYAph8ZGaQDxO7d9Z
W04LhA6GfEIDX8lPPpMT3BH1cR1zrNn/bnJpliwrSi/G7VtKNfqYx4woil6Ksv04
`protect END_PROTECTED
