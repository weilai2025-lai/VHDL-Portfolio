`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oI71O1eiIHffKFNLWovY1x/OFD3/0MWBPBSyUuG2q4LyevfuFbSQV0w8VQid/naa
lM6ijt1hEgkqlJfVF1MpZB+pvN/6BOWz09KdDWzMEnLTBYgHZgtYghj5eVC2Ja7X
5GLT0N+79uToWqGSAaoihEAJpsyUKy2hlcpyLqvzzwa3lJ6SzFU3m5FkclcvQ1+p
`protect END_PROTECTED
