`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTIEQXjKnYmxKmjwsS+9NrOE0WXyEwV8vZTdIU68EkdMDtesV0zzN1gYWV+1pAKH
PGGz+Q9uEkt+hf3o+uj9itYvT5QWhvCk6CLIyjPzvbf7AI01OYKcKh5wwgB6WX83
t7xIRV+epAo3SO1QomR0AseLgTEVIpUSGyLg6iXGN4bmZq3KvkYcPYHkQ1NE10Bp
fc/dlMRNKGCXURXECidBId/YbxfbLF2st81u7p0vxujP1UQ4L5lkKZ0v98f0KibO
albJ6nnwnoD4Jr2kYLBd2aYjhBmk27/5ZneUBlXMNWHKxkm5VZ0W82hl8YQVI0o6
P2yoWNYJ5wy3V8TeJNjoGgBkGJRS3+SqntM+9nnZWOPnO8ov/drbVGqB2a5TO700
+yW3f0DL+CoLNHpYdkK6OfARzl0V1NO7yb3OxBlxBRJcgxFbxZbe98eHrESkXDWb
K+wr2EeCDoxxpCXrNbuuuATxNSoq4tfKYqrJ2p3bDIWNB44HUmhQwPkQWjQqWa6/
Ky1GfPkIVysoq/z2ikNIB5DtiVGZLEgkrH7II3UlzaB7mzBGmfp/NWhn5jXp/lng
Facrox5+BvnnVOT/ZviC60B5EyTnpeXsR8qnjnkQToKTF0k/eW5g/rEH6SnXBKdd
eXFR7dReXVIBafJJ8rQ+mFNB7kddOl7RQHRwAqo86aKqZm3YEbKsxHTfr+piwshG
N0oL9yKbn9Jnw88pcIW0W4y1U3s3sJeDb/XwKx28UkL9cZtGihmYGWy4bF12/wW0
tvlJkHnzBf1+AL7+T2PUji5SIJdy+zh2P8wQj+kpzd6xh+TPDI0orqbG6thrd50K
+po1RUWSwlGCpZBcq2rls1EKKIkcf9fGg7C5jtLILaZI2C4Smr8v2nmntRGBSuy5
LFf3zaZNMiMgl2ygiIqrsPBmVtHcCiqUmFsqqlJVqfKEzoLMofXglDTvHjz/sJI/
TpW+dD212TRDNL/1700EsVHP3FTMMFmmqXLDiUBhb7SL48Fow7iCjpN0gfI1L+/t
YS0pa7ZJpLbB5raOeGXLv8pD1/0ZM1IPYq59fjVdBluoFFnDtTSmIF9Xi8JCGdHN
4Ey2Hb5uFpkJhAvx2BZQCWHOnmlACdWQeOeK0OMO5h0zneZXF3890sNVK/EniEUS
MB5R3+DPTIZKbOjAwbUSom9AITOA+h0K90yETeDRJdMcxzZOyhJxBQsoJirEfdTK
r4AJvR0DxNCmDuamHylQCr0aGe4oaj+0IIHvXG8sltHfBgmmPuxtB8G4XlvV39NR
7rAQPyLVlmFdK6yOZsYG4waUXBel+zXR1fH9ZiQYPT02WBZNIRcXJa/Kdlg2dRm0
vASnC+0orR1cnliw9R+xDxPmyAuggR7X29Q6kb0b8w8EdyQi2JzSt7s4IQ0YqWRc
d2cZ4g7oAcIUPUeQDRQk3xjKMBiwuYZi5gs+786dGVyHlexhBiNJ4uQ+GP/zMmWy
fcG5Io3+EAJ6K2PpQwQ3uUt5PLSWnoN29WxQfqjcFtCDqRPml5bHS4S2ew53qEMq
XY/YlyQzClJMz2mKcDuwGr/8AcK8gQ1izatWEOyVnIuujq4m8DXvdAPQhGkKXMkq
ZS7h0FWHCgF5Abht4az5vqP79noa7aaHWlU+G4IwfgE98csMqbb4l3mvCpxt0j0T
lA5mVzZjH03rRiLhXL+pWkkrcNrbob6iR4DK94E/7PYnelDV8NLPiiJYFmoqliye
7qnVARIQvEo6eWI3L/gv8bOCrGNUnDMOhxSMuEt/Zfh8vmIaj/dY8LnZHu6HbBMh
LXwYi+tLObr7Lv+zKHXAiRR9j9OZh0KEH6BjwrOQy8OjxeyCcDCf88KIkqze6dnT
bevZJldPSwSBxSoH6PsTiEPOQ4n68q4WQDHD3qJuIBewqf0Q/8OruOGAI44l5rRA
W6c4n4CU1tCHvBIYjplfAPe/D+LzU5k+t2K/9GWGsXbf7U1yIlB5Z6LwBzo2h5zi
+7TEOf+lxYHWhaH528BMOPHx/s1FF+/4/+3EUmCx3BA1IgD7I3BK4+spjz49E2jb
wP3We++3xMkuFkkO70wAJ0el7rHMr8KkAutj1OFZeMdPiySWmXFS63fO76TWaE/g
bDWDr4O/ybSoVy8VfnqyZ4T/HXfloE0qaAqm0kj62ObwDnj/MJ4f+yduGmV6VMNH
H+q7KPIrWu0ubfOHXWdD9pEwV4zDJb2D9OJkAaKpRJ8woOqcPee6X0+3CG41Eeal
X41gh0jq7Eyfy+f5CTiPwQ7kHm/Oew66G09yoq8xVIeG7JuTIYUS2JRlDE3KLLRg
1ebe/VtDLVZycPW7+WhVZyidksCN3N1YoZxtkiyzW8qXn3OecnEzvOzWMTaz7H81
UN6B6SK0m82lHrxG92xCgjZ3PVXmhlK3+6EFuKj8L7c=
`protect END_PROTECTED
