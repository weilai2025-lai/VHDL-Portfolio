`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJv0tIj5Rp4EMa8FixJYpkq+kDBy7qwZjFOnY75QPEG7sx9ct0wVC2Z+kxFbqKQM
qvUsV6biI/s1Cfhl0DXCvcjLg/sbiwzodnTE+cN0tTmnzywWR3sojz9he6LljWi4
sNKdPGp3jF+kaN2nXsUtyz+pqzHWVAZySAzZdSP8vs49miYpYRX4Shq/ewqhbLnk
3gI816oOy2epFkGgco/Sry5CQQNW0X3EfO0+PzlCikqFRZhs3AGAK8xzQ8jU6iTq
3pJ/1e6dbNnmCdP5m4SDL+CsL0cCOt45TzvQKFRJw9YFEyxU8h/iu/3qduwymjZS
dYvcAyoifc6hTIqJ8ZjUTHGrga3kpy4Tlt6/WFmhaBcIFpaIolVFmYm8KMRZQ/C1
zrdqHSpmBaj60KyzeYmKDNOkwuqAUscyT7gE7ulby0r5rx8/S3xnOcGs83BbezIo
iSpiJOfeoRF9lMrprPQ6InAfWT5vvrA2+U7mQZA+rU68ow9QaXO/CB82fvr17qwc
sEuv+R2fA/qFVG98kJswknIUx9quNwy2wHxMEFrSAIP6c7BGwO3/6Ig6asFYDXrm
dCXsj+HUNuRxsnUZk9wpuAJ6ai95FMg7h/9wqOQ+6x9YMfz8kWMkq2KHRYjILn44
j6GfF6hx00fV/dPIMX4kXuTtuV7LRO6BEyH6RjxYEn4dj/eZuEeXcODzmNmKPEIv
gTaIrrCAsmOJ/E8+WxTh+dGSGBKJriFysTO311sa92cBmkO8P40rlX/jB1FpLSnj
AnJn6rwaYldqRrxJyptI6A==
`protect END_PROTECTED
