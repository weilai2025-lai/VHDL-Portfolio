`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0GU4YEiLHigVSbCgA0gewaojPz01fC7qO0GYE2VfQaxQmMK6rdz2KL+1c9rC3xLI
KJxpxwmBXHvH2uK09aN87zqwxBC2qGtWLHyMbjj0KMFYJqD4ZghR+ac8Eb2m4gZI
o13sQAbYIegVTz7T/T+JmN1aLcL0OcPmyt+JSocQxCT6yObXyaZOtvElckLdbMZ5
zjnI2QFvTkARSi6ASuxQSw/IQt8PfS7k+SgAmEGiQtgdDHEXFmbkmYpGl6IVWDUW
TAUcP3JOEnNzLzDGYU2CgSTOeuPKWpSTYcSb/ewkXC63qV5OT777s+hJpP2FRJk4
i91ZKyPvfYDEZsYCsPRLyddwE+mAjqOqsV9rK/tT0NHE1cKyufx6B5AbD6lbqRlI
g5RqaFRphsyW4x0khDk/VClAVw5CUkB5SczkTxDx1ziLLwcLJm1wEUTRr/40KEwY
iEy8oMiCkCGNi+EMM+rnkEu1JFuEFHHW5d+TLQgjuWvf4CGN9xLNfQ3/tXi1826G
GJi3iyKRu2Glt8yYL6SxK3UjHsgFIAbVnh9XcG+Wop3/x1Oro+rDdTSiHbIFpWDe
WSaPLgiKs9FWdFLyDMaNKk5+/lExBJHrZB0XtPK0jjOUMzl2MiMLcRsDtjPphxGC
qR/HqYfZZ4WueUc012UQjK70gKRo73Ox7YS9YDj0Ns8ojFYgCHbnrwAOUdQxC+uH
Enw3QklRKFsolkIR/irXdcG9MyWl27TQTaCSNGKO7hs8tplL5OjSjIeBWjkfYgXG
uHW26HSxDrgPPMZ7spVyx6cOxMOqIv4QhuRdt/J9UZeaIYN5gVv38ll3gBUII60P
/o4L+X8Js0wtkFMLQTz5oUP9GASsmxWcDb6EpK1LLHCxrSVdlM5q7majqYA6+P4t
9dKy7MtVDE868bseIQyIdYezcDvWbE3mZJn0wVZLxtWYE/JCkLxYbsczdVbv/gUc
RxAKSTysLRQHFFF7l93JKLKGbKCwjA+RlBT1ON5RVIKsKoArL4EYNoJij7H24QGE
v51pxEe/O0e27avgpsQ436FAZonM/IaAFad1zmcd192vYX5a30p5A9NLsPzzEPum
vVVPSMGKEOOqZq34jSXqgaTde8vOA11/aUzRNTpUJTZYbrhzSldf4gbl0L3CQJyd
FkWexM0D01GNzZ4JIxaO6Ccuwstnes222FJFjGqjZI2s70r0k8rcnt2iqVL4/YuH
9h7m+bT5D07cCdeaBrEfSyLMeqIR3GtXSknKTtf101g=
`protect END_PROTECTED
