`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsC7TnWvZ2kpmWEmAdsAWspF0efXK18reGzrL8Wdd7Vqj0rveGVE0FMC+7pzfE0c
nHN3KqGwA9fOyGdxkJ8Bpr4i8e4DWtx5yVFiEM2GPHdTncj7usQHmvryBqy/MnlK
W55geSMcreV3n2RuQE5U632B4E5t1kgXNX6UeDLULEj1jul6V7VLBN15m9DwZj6b
Oij3U2DxYQYTTuBs+wxifehsPh611ISSHJ90Eh+nkaSucRqEWSb5WLjfs1U6BA9A
KIcdHN+mgjYzVH+Hwoomi3osin5jUvD5IBNdthCPi7r7ngicuDT1JZqJafBDeM/x
hr4QRRz6lmGp7zHh56L0XMu7fdqyW63s9EAme1CuYIgvwXDB4FwZtthO5KsuimfL
fofIeIB9APVQw9VdUD2u7fY8rGitPcPSUida7GZXxXKkYzD+d0mSucAe2ix1zdlp
6B1pbMT8zuJluTkDjKcE0qO9TtDYxUSfctgsYtBXOthM9aeyOZwNYjSmUMH5k7if
u6qS12ElYnYw4DldDuVuVjfZ9T7IBjx1JVgpD7HZ/6rau8skqcOjchHVwS3Ub4qK
XMXjAKU/rR30fG8k7vJS5mJKfeo+GASOvI96UCrRjWKXow58SQT6hhGQGNjq53x3
98XO6uDDtuZJfbNYDMUJbDlTOTJjuV3towFxEBjLdLG57mc/O2+zXLT1zJ5oQ6Xf
bo1itGlK3bGh0F4T0MuzrNFL3vTtWZKtdbhEcQOlSG3AJ6X/nMbglVoCrAabAOdz
YvmViPW2zsh+LT9NeBoMKBtVsBFo4nIjj7PrrvIe1mLfqjTz+nRonjPdcG4/juH9
eySyzQRVVealaAhYyqc7c5DsbjwIlx6HcrhDpd8a/E78msJWGdgDCupC30hm4Jiu
Hab8CNmBJzXgmqsyp/Kzp6BCb5SyE/YIAZkTLQyOs1fhdZt/PL/jGId8/EBO3PCi
H2yiPRlMYRqHK5WKtuBIKDwP2zp0gYkvSQkYe+Y5rlNLxUw+zo6JGK4rTr6F3nJn
JLcrVXLcJL0OHy5gzERgKkRa8QSNfznuSAH4Xrcvr3HmAqpsfWVLo+Zk3mtGxJ+d
M2KNGcRURvYSEIsPtwlTKhhNkJioMlr3Y3DDpL/f8kKX6Q3va5JINC9m3rMP3XIi
zQWGkHOzkckKfmlkq5rU3bQMDnhpx3tkAaJV0ehiA9ljA7ng5MFi7wt0Dh3OXNN4
4Xy8falFgdjTwuw2TD+SN9h94sZ1uCbysMzNVLryuC9SHIhQF2+FNNTGAXuivqCd
FTl0svr1Y/roaNioXnlLI2DQDDm9GiakvDuL9Acfc7IfbYaNhh6kx6O96IBjAI4z
px3kVCjjwjtShKQ/1DNPILrWlVcbJG8D57bEIIAjDBvOlIyEpHBHW8wIAopfr+Jn
ozL7TIbBE0VWjSHUX5aUpZvnPCf9/FXx2CDIh//A4X+ihB3vIyrwyRCw3YIYgW1X
Rzwvhr+DZ3Wm2yIvqoYqn3Wu7tfPXdldLKFvuyVttl8oBWqmWouQyTodml1GZ0As
qVbl64Cb6TEJVtaoueL65yxlIVK9xysCcgH22z8CjwuEy87z0A/jZY+sMcFn7vts
iF87AH03Yc1HX6bl5quIXKq1nBKvbI9fVJyOXFbQ02MRHvJ4LdLhUUV6F/3OrgOq
in8gPoKVswNdj0ndh+7zR4ldCjzMIkxJK7gHgWARoX2gg5eddVY55E4gg3BukM+a
nDw+4XCzmqbokrlaEFpcJ+W5U9Kmo94UZXT8kl3pXyRyDVcvvQ1KwW4vYKCrinoK
lJZZd3QywE/FjmOfMT/guVsUAzSSLe/oIaXhD6MfykFb/nahU/CeHQ/NP2hRPNLi
nyh3CQfSCGTc3oezSkKUpZroGApOVMmv4fjcT0LLa7Rr3mx0wkNH84KtBl/5O3RU
K1HY871gC0DMxThJeXPf74ST027LRvuguEEwhSKuAkuhEyAbMWN04rAxavVFJmZ5
S484dGa4xQZZEmhUnEdoitaaDIhHLMNkLTU83/vkYKbAmFjxbhpj7puVuj8S3q3g
GV4Uki8DZkcXjM34RKi9xg==
`protect END_PROTECTED
