`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/p3WlBSh3VqAUhM6YCA3amKXoJNmurOeL+10ueSTeNl23IMG+1mh7WKIqFVSXmmy
KN3unWKAaEhsH+Vdpvz+J3bmSKjrY7BKLQzA/Z6em6vLfFrfmPokbJOTKashe1R2
r8u9B1tYQW+SsGZEhTQK0eB9bBkZlkxbGa65pxJnV6nBPVW+qArr+GChfSZcp83A
T5zL4HYp9hCFZFJMq+zgh+3SG5ytwbI8sm8MneiV3MfOppMgTOCwSpaGi26Gin41
urCKip7SIzK7/Uwz+242RTZb7GPdxg2Jhgz9afP117v+zmV5/vhU7NomTfBkMy1H
/tnPBl4PEs+/2ktibJ1jMmyhs0af4L80NLtRj4OHfAmn8Wj6UwPCBIP1HD7VDnYj
lKPXJKK/pkgwpcdb/YznImvE8UpVRB6iJZEFzBSL3l2/1d0S3zp5jT599wA53k9l
9FfgBD32Odp3ngYUxvmBOxGbcbj4ybwxvHlyLPPxDow8cwW1cW5LrwBmvhC28ocB
84qGQzgs+JgrF3OWIv3XA+KSuMbiR6eXUkaMoHcNKW1l3f2pIIhcExIbPpqNsl7V
ggY4J4zcFCm3fi4DQl/9pAueCmJOI9UFpafGXwqg5Lcq3O1+Lq8s39v3W5ppgafW
i2IJ8FLLsKVa0M0Cw0ALcXY1u9Gj7eS2lNzh6vNpCRCmJ+U/pbtuVLGC1uFAnfjN
bWRg8iN1XPzi927RVynu+KcQ5DWp7fqJi+I8XAAn33CXLNaeyNlEamvieTzunv4l
byZdcoxouezK555mcJIPUNZ16IOdD1QfFJsIUvMh0WayAS1IicIK3GtjvxZ2tJph
JTR/gII0a0P1XBxPAm4ffCA+T0Y4b4DxZ4K/TdwRT/x1c4EFA8V8Bz18qHQc0IuM
/9xV48qHO5KQjF558XpQmdKDLK5UyrKyfOxUMf+9mqELuUdbwUycbcu2pjhmVkN6
eqMyVGKt8JtZY/6LQFwbj9pZrURhNcXA3Su5SNxbJXNX0taj5kOEnkYlK2Ah39B9
CSxMb/EeASuFlyRhBsLcE/hxgTIXXqsZVI06GpLXgasnE7AcBH6bG0MgTIpYxUbY
qAafdOtiKZyclDdbS07T03RoCMG0D5gVsrnOz0mUlLK+C/f2uDf4ciWKzr/uwDun
5Y3+PDL9USG+oc3wYGM83GT9TI94RUarFVXPr3+D40PpuBCj0jCjSQEKQYIImuXe
tvEiVd6KkxpsVXgtmUKJdXeRGv44YH0PSPI40EPSmR8UVpTeE0nmS8MkQDSXCmoM
mRg8EWVhS+hUGqGECrW5zRIEXqcI0pBl9auo6uclOnH4oWyOfBfCSkmPCyc71w7d
9BTCuYj3scC0FOJx/a2NEJEEKH7azyCNj89QQlyd1bIqOVd0MDhOU5CdHgx8zydW
uzQoF8zheAMNpwcVxvaARywUFsVjAmRMjbDmDMqq8APbiHARVP7ruB0jgkcQ65T9
9/3CYXfk7ulQ6HiR6ZOwJukVxQCRb+yKWHbwZHTnC8Ra62TrJEfOd0K0XKuBDLBf
34qHaYzuDnKRmLmPNzWMiIKvqffhV0pI+ksYOt1coR9UEIepslwxUJhfaaBdox9F
lqsYQYAf1CmT1bP4JDkwOM07VvbgIyBtaQpxbvF5K55YYRNS9jxohA8Xpi5YElxq
yMuU1HsuXv/t7lOoTVrro8HPntgUBah1bG0NI6gGC18B+XRsaUV60xWrMdTvwH/M
Dd0LgM/wZVcOD3QnE0ynCdljzDbAXVr0zV4fl5DUo5vClH6E3tGqDL12K4j/IS6+
XkWwhNEfEYHIuCTYy6CUdxbcHXcvUD8A4SLAmhwmiox/gQR/pD8LI3pa4uoW1gE5
EP96pNBYEeOgYTSKThLm/jrSjSzLUy0exYMYN/WdsNpCVq4QO9wk61O0azzcP79p
R0k83XKXc0Vk5ONDR9vTy5osdVNaJT9wYgQtW3n4yvj6grGTbyFlSUxfJ8mY9YvJ
pChvpSt9f99itrI1RIR8siI5q82jy7fHGIy/dxtwGs/nLC1DYh/mCDNR0yJMrtnG
FkGleUTZ5NvDVrCs82m7HPaHniQT5c7oVrhT4T3fPptUUYlca291z6pPsL/n3kvU
0lkW4wHcc5xpuUml3T88/uqmIS3j7w0j54oBnl6v9bhCiC9fN54x/egNZ8XFmA7n
GZabS+ojr/s2I6jwbmqQfFaTDhhL85DqH91CRLfiZRgxc7unU8lpDiobYg3L+ews
NfyZWS129msWOPSj3r1OAJ4b8mlxJVqmH7h9LXK6KwcWWvRtrMDAfTdBotxYwOL1
XLbLlIU0N07icMP/ILD0R03AyFJrRwX+5DePfWYxT4pW/+Gm/BQLfrAK3qpUaS/U
nF3uEyqCMFNoJCKl7+kHkz9wKakvjhcsh61SACwFA8ai63apiIiXRDG6sY1HokUq
`protect END_PROTECTED
