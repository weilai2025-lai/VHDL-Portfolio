`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8hv1Z9y6NThPr3/l5Jt7x+nIo+mI8McO6kL9oAWhmEExDKZizkwf2nQsLZPumtmr
k1gyxEN0EmEQcU+3mhLnFYZWnaUaH0sz+tLYlDbFmM6ik2dwBlc+uCZruCMOm2rY
07iGGdG2MJW5hMovtCR38kmm1Mb3MvPtjiqYBPOuxdpN2pMUm6ZzQE/q/3e1Dqas
vApMudhuq0ZhQsOrVViwF9cq42xI/NZ9XR5AGDP1VWdz63tNY/qM0715w49HYMNG
nrhMRk8jYaDk+22aWTp5qlD6C4dfc2PqKdm3vaoeGzj7LMBlKb6pnNt8GH076e9/
vYxZ6mJVcC2fxY4ywlqQHk8us9pL3E3RVtn9onlhQxSaUZhjd5LZ/4ujwdyT02wS
327LGya7Yy00cZye8tDGeC/6Y9sLwjRhq+lfrUgXMc6niSqDZ0Dv1pK7I/3ydN7k
IH/ylLxPPldSfYXLMAfNqRcrfxSFqTYNoyPR50ij8ze4QYkElr/O4v7bGyqWA3yH
Zq3wDa9Y2KLyv9mr+/4M0ZUFByNN0Vp0WnMOZmMaFEbRImHxtTjpeQIh8hR3Dvss
owOzcmRlivZIdgabI4g80E+Yv3blAQSw1UjFRbeXsbbCvdSTOfdLXgitQ3tWBJ+M
8OxRleSDfeQDNBm1zBLwomH/ifZlYilbF2VnqJI/mG9OFbFlZkBvp5GhCF/i7S7O
up+G7IZ45ujj51cxd+9usSDG1Q86IrEnTKecbRBjpdfk0VBBNlmtCNXrpFXFroTa
+eqvMCyEQff2zBhq7ap0yuu+NoIPcVP4rF+dDySLPtxoOSgiyFzlis4NMhUwPlY6
EaC8Lvip/l6sf6B+saqotoxOx0OgsaOW2Y17+L6OMjRLt656M8/0h5H9rWryw4RB
zZYkp3j9ftFVznaDrtQeBL5UKr1htm8F1RqqT/ijWgVqbJbK+RkzPeDsbwm6w3Cr
uC7WUHQkMyV5SKQEo3WN3pnsdsoXqSLaMY9Js1Yj2DhajS+g/m4iD89WXGyr4HT3
LLg1QHqXt9lfa2/MscDB7LFB87eXX3IANYxZs/zUzxIiVr5ak/wiMMQOkrhLFC4C
deNhdqzS39R94NSZA+WcikcwDoSK0HSal1n6h5kW3cK+pBns1TqhdvpKF5ie2yG9
be0B0UFwd6LP4mgeXWKHY43SFSvsptHx2Go8voJBfce8IUWABn2ecz93OH4O7cfl
gETHaChwvukTT7Rz7VLVVpKzWCZhVS7dU1mbufthmxQjeyKFMOByVYKfd74zX2Mt
dbxgwnl215ixRvL9u7nZgB2OzHDP3o5BVuNKMCqQBsvEJEbuTj/0dujzm4+kXAX3
TyXsHyuqkiEs4uSFk2enHJNSAymR9TzfjLF2VpB46HAfT4gK7pm/t3w0jt+v40DY
AyRj9Df0ZiEaMSNAqJlm9wjK838zl8VGYETa5HNApOI5Dgaa1WlEWmGGptDRfAEZ
M9IHAjU+enOTyc+kxNzhG3kjjhqn2YkD6VIvfc9oKorzCD90VljoBaAILkRd8DnX
93jcfZWd8hM9KXkBvqom/vJxLhR2EsKTnJ2UbfowVh50cELyjG8R4u9B2NJW7ZDD
herX1iQaIhUZjk03wpEkO9CIuffsDtKKc/4NJrTyb6iUFR0mymmeJVEFRai2q9dS
XltfEmI5uonFM6cv40RSyZjNz5dHgCaPDhD15xBNJWYhtLqNwmVZqdz4veaj1aYM
ieKgR9uH5TyMue12c0MmmF3+tNSuXmdLIyrMKdT9xv9ZQedSwdx1SaDE/0UDqPGG
cFEopEic9xY7oc/FesFfc+G0OXG8JJbEv+IJthbUK1/YJ4hWJU7HJwvDEHHUabQg
YpUkM2E0vteDOGqUbXPLnpF2Tchytikb7Cf0X4gTvZ5ljqKt+5wVQlzX7maMfBIo
6sTh3ugUvrPEMO11WPGqMG2qMnXm8HhcAb76RKrRpKQ2QfZzDKw5Nr+eavJ6IeMl
yhgIXVWNepvjexjMkq4qXjlHdqulggzlYEdH5AU5LfsS0Wtn82HrjBwqhhoZijuX
BjARikQyyrDRPRC9bmvz/GN+ZgDXuLaAoEajEHe7xE0iLcxHgWD/cZYiNgdkgXjI
pITb2wkBjqeeBzHCL+EWTP6fvEqiQOA2y4ngGbuZHxnyafG9kdhlxNu44Xokn29R
IMTbwonzwmyRNXWg15qJLsPTXp/I/eUjCjfbWbZDxYIdXI11To2L9LPVhaQvZMox
IGIh9IJKZCFcoJlEv39XsMMFThjQezMTrgsdGQ3NGJFJiLvUi2IHH7LNt0off3QY
3sf6db2UmBWxfGSu3b2CrQ5DufCnSG33f2JfU+OtVWO/bNHa+caQw4kfMn+6C0Sr
ad8zGIGrC08JUKg4FQmEncYoOSyeJnEQ+xn8mnxf72nA+LwtSECjPVKO2an5gQIH
+khTwpM3VT6JNxu8WJY3Zl5jXSpdi//83i8q0ADH3q1wxJjV/m/NBKNTEopR/nF6
SRDH800kZZGNh4jHHAybti8A9A4jYz7D12ghkwJfyESpjepXF7Jri3SKVV/1AuPx
RrTnfeWIBtgTtlp1A+tcYWy6Jgrx0YZxcq9fYNibH6qy1f92RXNiANj5cgJLDJrb
YQgl/GVK2OAKvkWax+fGV4dszaPSKrPuFSwKR+zdHXEXf+VP8AbDWjfZ9XWa8zI4
N78Cut8M9K6PSRpl5ORHwCHLnx6PAwzXcj7OKy/1GV6yOSq2hivvir4F6xQFmL3C
ja/myrxBOkq9FRu1pZqY4Dg9bUP5YY07FNfKasZIlyC5JleqdFW4lo3Bx+JrpHGj
sWhF91pysAd/qcdDBAWw6xC4n+r6afjpViZ49UhaN4kvf6DdeNmX2jI2Zy/SlBOw
TnVyODPcLoLC7AFR92klDkgD7fOvp8oYodrwPCtUv0qa65vkxz8F9i5+kVXOWzQ1
AqYYW2/TH3tWZryq+sJ7TZ4ZbHsUbAw+t1Q7KO1WpfZQsPV7zRFgdIw/VMoDGMnZ
ssjBk1J7WAiMPqQoNRcY5cHd7dLTUCLTzAimLX3oOnTPGAMRrkbmoNzkEc7S/sKn
Y5AsvBQnV6UZAG+am78WJWrg2cV5MCy+sYa2S+XCfMAGnqRrhhWrHBX951917JoH
QKO4gAlIW0Ro/RPQkBk2gtW9IA4tVraMU1rwvghD8HcxCVCBhtwTTpS41yKsdEo/
NnVhzzSpDNs6A3zRHPpT1mWWgi+SomhvVUHv9Qs37HlKBANChF/eJSAg72tal4gl
RCncrNl5J7WjmkmCr+suPfr618ylyjonnV1qiH9eJZ+NsdcJsoCF4x/pziLJGmTU
OLBzthoaHiAD+aqba0vEj3zw5QkMasEgbehJ56fv+oXMr36aB42ni0/zN/Ci/1Ej
JgEsvlH7XLMLrdxYzG7yUqaNhhr4u2qSvsXJl0FYmPyCEnCALyDGcFOGJk2aNfLX
yu0mA/OUbq1bdE7FJBmrfyCY9TMf8PC+71faPraQhNqNWA9QJtgqn2X8o2aoKEk6
jt9O1IQyKEMI0863cyhwU4OsF531/E1ndUq0Vbzqpg7p2F85ark4fcpYtaMPxT47
TvAdSdtwJjJnHRALk+m5xatn5V+tYXoAMHCQuGnzSog5Wm912EJA1FJEXdktDdul
D9cXaFzaHbZy+tiQV4Ka0sIYF9bhPwDJbraV5M/jiVDs6t03sq3uJlxWwm2lC/ik
hoQx52JC6RQQHjI0oP2LXDyKcYq7ZcsjN44IhtvioWKSkTFGrLtYidK/Ix3mrdsg
uVTNGYOp7UPEoKnAlyQnDTNTR2TAH0k3qPZGRmfKeUi4wQdGSbqGu2wUFnmrMw3k
aZDMWFYykN+ZOtjesetBINrdT97O79eBvKMHlWTSyAwgowkP3nB1WYzrK8Fq58v7
xVNOWCSMDY3MIO1i3ZVcxlJVUbA0ohEsXZMXM65do3GVAGEWeXxVcoDvlPpkswqh
W9joek5OBZFg86FYQrtWqjdo4X1T/fS4R3jDTG4aKUDhDfTVz1+wljSdQRGaeW7o
BpL5iHNse0yrZRj2vrKgixJj1eMlOLQlSh4Bend5ymstL+H7dUSlRcnxKrIDXzyj
yneG2s9geyWJKQPEcE48V53YA4oa80TedXaQAZ78FWIvSiyxh0KqopqeDnFlUqAy
zZrJILjpI0sO9mYCI8XvEa2rlRV0k1Nl1uqPBxrymc80kJ67smExrODAtlOeB+4M
+nL1ZSqRMpKBQmrR/jyx9tdmm5chA2r9cdzvmmoPaV8x35TeaR2ObHMwWAnFUXWx
7D3JzT++RaOiiEtG0gGkT/h8433UfB4sOiQt6p3H/yTPV7peDOaJdiJ1PuD4vmtc
jZNfNBeewyOVF2jpajo561ZmRHlSokWlOLYEp10l8XgVfLi++xE2QbpO/avjJaAD
MweKUXTZdxmuWjTDdJVnkAAhrTzHLtzAFpZ1SrTIweAce624UyMEZLWfXe0I0X1I
rb9Izuug2ELKk/1EUNY1FaoD4K9mpZ8Lhu5WP50TYqOI5GkykMUxmtW+9ZgRes9H
KedYhsxjIuDvhixLI0sBlSL4ksnzlNwIvo/GGnstkh0VvGOFoWEGS+wG17AaJAZ/
`protect END_PROTECTED
