`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F+sgHXKpURmpsTouplvU4npGbfVP2/NAmIHX/7boBvYbQmgLusV2vlqioNop+7E4
bxkemDGGlXaJ+U0AgydywAeHIwCsbo+l9SnCnjGKu4V1vtmGoZ3RXum2hkH09p1u
XfAX1gLo5Dg/NCR9wfWTG3itzrD0nN4QrCwuuUtxbvSlyrKtUZx/5Z0Rw2xsDVTW
+NXkx7i3Dz5D3EOYq2GOECahFJp/VMthXtyoJVKd97nmyOX4HPmfhUviqjtFGwKp
x8rS8XYBuU+ZEfhr1iAINsR8Tix4vakywW8E/RM/CFdYc9PObPBEWNiCwRlci3bz
m7nJmFaR0KqW8Jy28wS0VeET5LvOgV9+ABGHwwTciaRGz57v8wI7W10huFunDFoj
rnJKGoxApsMb8/sV4zdOg4rh6bOmGDxB09Mqfyi7cmUO/qr6ybz60CW3I0EylPmo
5x1CdilWHWRrFCEyQ3w6+nNjEX8oruy5m/MhcnXTHoQGNOuXcxg3wBczCZn8DD9W
VCi+ZgvP/N37U3nnyf4a4E9vvD6jpp3MFPh4/PyjsxyvfUtdGx/IayVguPU/x+Vd
ZkDlZzpqubac5CEsl1OMkhGZTLLtaMF0HfFVv2Le3eM7ow1t4DqcjUx6O7Bu1rLh
DZlJF3Qq3cFqaRjf0uUWvRyeZhMytURHt9IHrv5jEFlapOfDaFWx4j23bd83xOwR
uG8OisB+K7xmITmq9yJummYBrlg0ASthclZfFEIkSix7j2WZ692A1Je1CPqxeRYI
LkW+1inxFkvBeDpzknLA747S7htksA50UqSkj7Ca1KDQ8cao5gv7/H3x9RRFY71h
K/qdAoQjj6K6dj+jQgk7HDYyCK3emHPfFrke6dBRA3RSMilSbldfxJbNomaOqM13
CF4R9MmBdgI6OZhsdS35YrLK5NhB+3bDzWFHSgiCRYYBp7CyWN+Subo/QmHk+sMD
KlXsfLhOw0sE1X8remyHS6v9J1j1hLUfbR4Pew+I5b7u47PJwE2bVvEgMbesRBK9
H4C9rNcp5f9slqXX0nMVNTLvw0Xt+DkMYg3LSmLkgMAIK3r68FAKF8/AH147wNWF
HrngMn8WdFAWg7WxEpuc4HLhbq2Y3hVvSyqT3nJkkCUXVsDLEcAou4O+gi6MrdJV
YdVS4dz5QbMxvo3bLidpjIrbT4qmH8CIFwIqYtswSmDps6RsjzXYZQB/moVclePG
SZK2PakBu7PxwfV4uOKq3/ZZrq/IrWP+PLVhJJ/mx76d7bogEBSfbq3WQsWLr9GJ
K4HS8503q3WaYnmT/igLWNFNbBAn/ZLb1Z0Zg0OgoTtLYuqjzpp3yaNiCNfZMtAp
YGwYxJWcKm9j3u3l3HhNZ02W0DaLd1rs2liV0I0w6M8ZIradfonlvKCxeA/73FTO
5pXCnXXXXdjQS5jUt3wf9fsLvjPJmD4dJd00jxFhtj8YeB8DM0Jm+L3mRfP0tgb6
MH2W5Oo1+SmmgjrBXQUvg55C6RVZowtkbCBk1e0Of10nltH/qYG6K3FEMInm//ja
lfT18trP5g2ClLitBYWNgkdo+2/PIerD0hH38pMtrx2+I/6tJgr+eVqPF7jW7QWk
raIPc5eNP5dueu0+2ssUW/4B/8QF63fp45tDpD0lVS+R+BD7+ti8zjq2qNUmQ255
sQ6jz2FuHJNQ8icGg1n9DH2FZMZ5Eno8h5Z4JxxtbUKZjB1ZXkGhaMn+SjeAkR2m
RyKp/2YpYonj3IO7Xyx1oA==
`protect END_PROTECTED
