`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbKj8Eo9S7MhHwpNecp9H8fU2Lg8X1iZnMzxPtVYbJJszUqemGF0jiV4445R7sXy
1eKXMHh8pRSIk9hlwATYZP/6DEXeFebzSgPP//sCbdAt+6UNpxRQS67Zv3puK/v/
jiTQ8lpuFeUYgjzwBfkyJRXrMCAT/Pjn8oZjUn4MA3sj05oxAC8V5WHbQAQ9cn42
uAlQAjuzlKLktpnbMJWI9zZJY+mCAj9Xhl4dZ8gEvyA33ypxpJF/IqhOkWhq2ELd
GnRhWtZcuzIPC61HSHDrLJg8v/5n4rH1265UV+EGtAVyq3TNVCcdeCKO8Z+rSuKl
Wzh7IWrdOuB0k0WqoYyOzBhMZGG0VOUFjl68VDVUG5JeAE/nH2hnJfjr3jLaUMuY
EW7TeEFHeEvARYNd/Outn8qrOmW251mapB3YEcOz2F0d2IQh/ZxDkJoIbiH3XSeL
gmdZtT6LiLE4USYO83NkmORBUxJ59BdnW1p4xp2ttdDub7d3xjxoW69L3ms+uKKF
yyyFVsAzssis9ArmQ8uyLgM0vg93q+lG38yNxTzbyV7/i2IJ45QvZV0BFvXL9ZK4
dGYkxdV77BEfHWCCet89GPT0qWGLViWhrPvSFCrtG1kyvs7GpUfjQTTkZUBEpUEI
T0VHftKNKQWPPxnjg/t3RQWCRT0siubzwoM8GjHcqe2ssrrvKipIJDwzXMkvvp41
3YNqvhVqy+fQ6WlfBJcIohxzI23l0ks0HXbTJ6Fg827YhhpjL+dZwDVZjZaMa4yT
Y16sIUA5HgH0tf/3TCPoPBWxu0azEonhiiNqzcypR1CrAD0BWK17EYxusUssLEyl
lRJ4wdTh/UMlYoWTQkFZQ9znBHX80dJKh21Rhq3UHbI3ZVO64Kdh73l7ZSxSzyrs
kHNsv6RP0MzS7tgLf6eIiWiEPUgAaxb2edEcqxhBCm3J8Z/l0oI9iwhIh8bUIBDC
flXvbfIAPULErndCLNlEtyNAdGHGULEJpAek19tNrcp0Dq4MJiJy3ruAwunfOeAp
q8P9zLbxgiViy2+HKm6B3RZyhpT2FnMCLOdh6FHoIQgjowtTyesrb9EsBmv9LbSa
7f90GCk03EiGLe60pcewP3lBkizzNYKbwP9wgV143kU=
`protect END_PROTECTED
