`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpgpA51rcj5ACHnjuQYZdvSRIIxsIijfPbmavLtriMT1vqb9+Nll6bLaCjk+j+Kp
A/76USHrnIMyPVl0cesaI6qcNhMoGDz2JVkVSTsw0XeSg1TcqehZUUVE3bOjqLnm
8m4mIdAvlEwb4w+eWCEzR84XH7wt4iO2gKJpCw0wqL5z7XP2yAih6JfcRujRljLp
uAnqP+GhmhytSZ3nr1RTGeC6xoduKayKejqq5UcudwY3yuSBeccd9EHIZkCSXRNV
RjZM7vFZwxOG9AyJRGzuU/sgsT8OgjIaa/fKEvAllSVSfSebdw7Jceo82p6cJVCR
B4gzwMgz3qy6N9m9M2urQYYhQST9lfTVpYa8Wdlz0Swasou9CP7lRbTeHG9byyAW
DNQ3xSXUW0sxAukobMeluoI+NfI6kfg4ncSiTVBU7AtkBQ3vx0Gcasu49F3/CC/3
XmWNgGt6sRNTCREI1BloIbaMuZqnxiybUtIHjOQ6OdqJV0iKSU9qwKJUqf2DI6h3
KywY/JBRyzNuL9mG8s4IbgEwW+KqzU2Wq8WSpPEZoELMeYzPLYp/7OfNVX+dSaZh
yMdmAJoKey2lPhaFqHPx4weCo9bRQ5UcTHyYKpVB8y4/5SzMry4Gk4AJibEjfdzn
Ozaw1BMASj4f/NYiIq26LaEQsti3i1tJwvLXWABvQ7m8ZGdX6OwQFn3iCsMQIRjK
ffs857P645OeZdkmIBPk3kgZV9p43RFMr8KVH6+0sLT9q6X02NN6Dton8pSFsbQj
Xano2qOokm/ZonTbkUUP7KBscB+FL4+4URruxkFFRdcczDfq3Nx0H7EE3Imjkczp
/pgDJf36pip4sgvn/o653vxT25kIALevHP4YuOkLmc4AChH/RV8QUFN8y1ZMvgv/
6dwSWdAxndTKmp/aNxB37kBBrVQ/oJAPJc7ojtlLl/n7ts2E2CvaBPLA0ofgWA1M
iheTr31GC+gCZoTfOCTgSiDWeaRoXKOA96VQOM4klHB/bqdL+wvz0EDNSf9bg87b
6K9+ZA+XEtFcR/oyTeoZ1ECZydbTx38osz8p11pYK9mTlHl1BcFEdodI+9b2ilSj
OZXFUJ93vinDzzS3OWr2ZrMArxOU90u4khtzNGWbKUqg0FC70CuGoqsIkSaDTgD7
5wNB44SKnJkid1tsCM7dBFzK+BCEG4TNgfyC3WdwbxR8cIZ9ianfUX0LQTniRwvB
nYRr3yv1ziJRUUF7uGu3D14KSnaD8Xp57Yv2iKU1tS6e2SrLia2pYf68jmlnAGoB
HZC8mYdYRdB/lnkH5C0AlgnZvUv99Y9gCy1kGrqmq6VO3jhLc0KwcTNR4AGKGSA/
eccl4naEpZWdrErxJaBiii3WRzDvWU+d/c9riqZMMdBoycC2gpr1PMp8c+TLtyQY
i/mosHP6JbrgtTvoxR71HZXg1KTIWMccnc7+oZP/UJJXmAT+TwCzvdDQmpUNeVOq
M98zvn2MjliFqiWX9TjxMyEfxA50KxuzmuUSoS/zYKSXuf/c/ZiKYd9jhtbqqCxi
vD+KcXE8s309I64Ojqy/GVyL0guzqglHGOUjxDV5fQudWzJuaP1wp0FepHzoB0+Y
kXDQBCSEd9amyZidQ5ANHPTuZqIQmVr8w/ZR+2s04BI+S36LlWUl/0EX/YwhibVz
X+xl0Sg1I/tkKABZMGqFzPwsczKNJqFYUwapWIdSgA2fajChFz5w20QyakhYDdjJ
vAeqXJ+U/rpfooYJ3kaiR4W79GLozjh3ZUtJ4a3lZ1eRJ8IPRmA254z1RQBw9adt
sz77RaZuEKlhtJ4x92afCIH0IJI/DGgw/BJRggdlu/iBVO29l9BVAwbW3SOQneJ+
hvDroZ6bKhtkjFrnt1uxtcDvk7TJWPGRRiva6stT9qZjWJ7PMeIBcX3jPO4Ky7vf
bN8rxwagP9SXNSIwbSiGXcQR9KckNsLxaYlOnVJxVeUvDF0MxDPOViAx/yHYpFh3
6JfK4ODcOvHHpeOw32CcDAR9sSdGOoUXyELaeD8uCWb7+0prgkdQp3UgtQuGCNgK
/MfhUh2WRyen28gchijv68e8bQOVbb3Ptfq4j7DMzYyT7CymIcWdUJBIVC+Za13h
mjpACielp8cIk/VFuatal/f7YvZXzIEpJcUeuNbXrio904PtDMzmPBukddxdBFiV
hxMysamkeTvhmKQ6HYbzZbW5MK+Eh8HuUequR3IoBSejWWaVdgT230qyyjlukyap
BpuifKgUGzfHxaG7a0kQVng21w76+FYpI3JHSQhf0nbFrBp9TTk2Krd9eCq6LLFB
wolroiWxLhhphJ5fCAU9NpRwmC80u/EzOqy5128Ny5L8VcmLW/mEayLDxMjj3CyV
X26GhMVxHeXRQlr/p26ztzB/pXcsSb5Ge4yMzowfnj++95dHFntFkKEBbC/qapkd
d/K+RR9gN0iqIavdaJhnlpoB4/7rXtC53CBYwpIXvuLBaDnBbJi6c+MTp+isvf5Q
vrrmVxS8DAcP3RWJz3HCQDlZttK/TWUUYHx1MJ9jZl/59L5+4qiWrP98rdXOM8HJ
8ovumV6O85Ue2w0i8DQbKiw3ASGCFRtvDzBVoot5w4tSmARZ6AEPwSfhPtD5zsph
1L12XmsjEg1tdQb6WsaOBBqZKlp02nI1uCbJJSjVY35dUK2RWEZ69DypERD4JsR4
mdwDmrrbzoyjdlwM6OfIPbF7r6RuO2ICYNih5imJhdHrMCUZTbL/K2ZrDXXMweZK
HzCg7EGPIIgQ6/jNCT3Hfb3Jb18wcW1Jssj8gl+vI5vvsbXj49NNqnVD2zRfoL/p
OAJncbAdaO7rMTOIpmvVbxpLQKXAEl1qexrWsu2g1KPOxK8ewhIi9y3r4aqTJwDJ
w3k2ouxp1kenvm6fWJUwPxhc4xVANJhBqrIuLlk9Sw5VpzHpOllaKKSI98dhPfcP
XlWM5yiY3kOPrWtLtWnGAC8JiPwVMiF5y4+HD/W92iS2HsDc5lq7mDhzjS6C7um6
XQPvzuuWi8hZLcqixbsdus1lQUzL+X/+1LMeQTR16LftbhjuEpco5t4cPyZJzBgN
noyhCl9/hdoZjdOIpmRzBXf+NPcxDzminOmN8zhE43f83jN+RUg4lc5zNdoK5roe
QDoOsDiKOR8xp41p0Be9qQIqheyf+HHWihkGX0L+Hd83sMXQKTGdxPdXSJ5r13NI
T3JadnCnEay5ysz1M3Eg2nUEHSzblQj2FJE/mM1mE+7eVkUaQSYUv1GP2xFxs+FR
hIixZ9iiCwktH35XjlEmDwm3k4kWVwjbHHWPPtK70tgntmnn28yZFSz14R7S1RIO
XzySvsDLqCq9TpFbMjD2TRPhfdV9qbFi1P8XE83XHKX1CMYi65rmE0kesEG4kLFA
CwZrejmqOgN7GCSjYUfFUHa12lwC1gvMnyYIVXMbHWXsmwpeIASj1k/DWbL3pOx5
88j7V+r6fNOhifjLfoHWEQ==
`protect END_PROTECTED
