`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h0hBiLSWkuyfHca1lVz5fVyCdaRgNKgcCltTpAq69z77elzxCLsmiJXVkglHmP32
D1uGKuUkMB/3/2rwLVsmpDbse8X5pMHkp1ySPjmUpSTItVtAcdHsXnPzSJ6N2I8c
94xt3XN8qtS6cSvqaH2kCnXpdaWJD0I1qMprK30sQF05+eJXY7YDL6cUlrr1E7FI
7tAmMaAxb9mat5x7inhnp+8NZKtYgbU3i6eFXn8Ifh2Y381iS8yEV44JhxBG5BTE
VcjLhWkapXiKd9Lo83378VQaF998QYg4IK+xLSWTahVBzbjg5HKCzCB4HIT/51yV
rQlYDa5x1rzcB+p/++Uyc8Cmk35tDsd7vceXjcPeiDoBKX5IHdwdW96l8eRBDZoa
L/OZtIVeQgKE3wiM7O3ew8oyUm3BVN/KR7lFt9hRyzTTNTOxG40LC0wNO+bZHo9g
cl7rmo4hWXHZdpkzQuOktkV78CNpxRDrszW+I0cdhBte2adboD6dXEzfxwJ8gCkJ
Oo+8bMqJ3DJxjVfV+prrNJUaNVErV7jRCiK46WRgmhCS02BG1icJrkkE0NMaM8Z7
76J7GUc07YL5SlheziGtq/2BmavCASihOLCXg7HYuoaSn24i2kUWaVmF29soivoa
7LoI45GuhTMqrW90HGxdfHm4RosHmRKyFRJuplojXCGej9d/ZK42u4+03kJ1fCSe
Esg5+cUzsP33MBF8c+4FjLQVngzQz7rjaZVvmxlidcEMYqb9DTOEdK1EwK+JMw2t
d465unBKNrr8tgrkiSi3UXJbyWj6pf5Gon/pw8XO8p9xSSpnlAX3fpS31OL2shCw
68canpkbfG/kui/J/u1Urlbi9izibzyap4I04Vn0k3GfEuPebqyjOZqru/8LdcjH
lrV552tAv7nhGI64U19PRCpsaXfyH5DerJVmFzU5jn+XEKKfuQs/O6dQ18zAgQvi
bhxuGuqPhMrTMG0PdA/kipS5TMV7xJ8KpYMPDzUeDbsYTNHFWQ1zufbAreSv0jRT
HGw/EiAhn6Z2J08tJ+3oltwsACiAwCL9I9V5mRYyteiJSADeVqIKJeMyG9s22S5w
majKiBhTuM3pRMSqntI3v/paHxWUV+sR73Lr9aBXYY6AtWirKBtjNkhiOh6EwuhH
u9QA/rXvqhNa6UCUBvPnP5ksABXc/yNx+Dqlw4NqwKbAoklsSy7ruChhiQIi/G/0
TfY8VCNLYa7CVl1/f1Km9g==
`protect END_PROTECTED
