`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZY1V2mSYulZCeop3vRcAdAuJNmuFtWoBnw2iIky2FX9ElDD1y391mBDSHFz0ZZK5
rg9vAh1sZX4lwBhTgQz7Oi1WVPx8sYpy4ufqZ+YaOEz8tLNepcmR/F3naTM+hoeI
4as5Y51mcU4yQvMe0+gDwXXV1lZnJXNtPB3HWG8y8pprv5BUuUcLs0NfD721gohy
h1h/awdvZwyO+lMMVYqQJ9Sl7Oday2n4osd8mrJKpB/U7m9D0T65xX/JmAN+8vLa
FY8C1Z1GqhGIb9Un3Y+nTlCrAMhaW+ugv2cP7EtQ683dkL5Vjjo61bQAXVXsCvQX
4jM4kbpe6v5jsYsKJ6dOGyvTD8WMLKcKs/Iq9sL8rQ5gMhRvFJTq+diq+J58hqeg
MPh9QXVHWq//kz69WyxxHrWzts5L+QK4vnLgmK65YcjAJZM7XdRUWhnC9occeuJo
/5nnyllw0MYd6AsP+0augr376xv/WJeFLyAY1xYHGx580Md1LzlqPRi88VUNQj4T
Vgh0wLV7gETFMXFAVUo8XpaT5mTFGeNj3VgJwPd3k8m1rb3dlWiaetqk0FRlQdJ8
J9u9bW8xV/KeIK5JdFPm2G/HYUt5VFJ3Z0G3tO3c6gaoRhktDTEcvrbRmcFxxVAu
COOMNFBe3X5hmoKFAB4zBYZZgzUlLk0vNgF7bO6YAu3xHQNHDW9SiCg5qTwbcQmg
gYAtKin6n8+wY56dCRXlF/FUJOO5GacIX3MAr8GyoXaiAFg3KsUIhP3x2NU67vNw
I5aHuZpf5y4otnw41V7odUfWv6DgXGXl3LH217hnVb6UxTGt7DYyFRY/YDXg8osg
EocwoZtIvpjRpUZusMrMr206A3lTVSf6wq5PQjmpzaYDAbhVPCVR/IkcZTh7jNF9
re4dJPXx7AMSsWx62i6e8g==
`protect END_PROTECTED
