`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SpeL3oEMNqE4o3J5IH0yu3TY2bCnT7mXE8epCL164Du5KY4tVl0hlp+N8gYfJRr5
V5DUR/8zxpZbCLNkCIViUPVnjK1TaPij3VKeu/t0rMOf89fEQpWRO+zagjTLLus3
NMUs2vVbM9ikU+UpdbWLjxOEdggDfRqbsI34NeBmy/9CshTI+210+Ph5kzcfXTNB
ADWdiLD4s8y+l88Bq1m7Ald4ncMACa+AgXqc2IPR9fGFgzY1OyEGRvVVDO0r+qr/
j4uS0iJ7XWzSuQynriYoEiD3uQ/K+xryLByoSR5ElioW0UsEs2YzK9R1J4bN7LmI
d988fuxh+GXCzsaOhzmi2Xqh1M6OLNiJjV3xi80uFuCBVnUyw0ZxXB5pG1eOp+uk
FbfkwA/G/sts6lnO7oohq3BA+iqyHfPFgCZ/q3XFdz9A8t6mbAoYRiZ+rcaGV7vO
Wbu3CLkb5jYs2PiN2SHCVMN5IGaK9t7Z7em68Vyq0NYWHDu5YWnsYph6RQp38G9v
ibsjtYT/hOdfC0Cpw4CUpKG6KBfRiqqjP/iADXpa8UlLvv9svnWkxrFUBmaYilks
4OShK6nK6POCGRbE5pQYMPP2Ow2+hWyGY+KzpOxmQFQS5mj//JCZE/9xqVUE3Jkk
+eYXwECTB8s4dq+Ju5dKeL7mved7RwHdm2sz3l/x2Olw+9cHGzbbMMWS4MWPr3ZR
+oQEt9gtYEOx6yhjKI6+SuDMNQCsDeXSkFipqNEBe3TK77QvGFhEKiM8Ra/5nG8P
IBON/FFlU0apCqFlpKW98FHIRkAdyIaX78SjIR/p//uqhiOPm/tZc0bdQJVfEzc4
DuNo2Nw7t8Y2EQAAyxVwWXGILCbPch2FjMZLEAKOETH5v7nWGZcvfl7tK9GXtnWX
GsztBMUzO3uhD8tu3x9bKZ/YU6UjCOKzUjt8EJChKZYgjpIYiFZ7UYG/ZL9qNJLD
jqWNla01slphNLbqZdcFCmUmtrw3pH76UQp7uZ3NC6wSyR0pVbcA8BG/f4vhjwDN
cZFeH8gcOepKhK8P1hJvR05mBPM9asjmkbDFratClMKPaplfRbE6g43bkfj/TKnN
zYASakMxXZ5A3/ndcrL4F6/0reAyaCpYE7xYDJ3v4dGjhF06zXpu4ehxVCtvYums
oIzTzoMlYjL7/C7vTS6bpyvb+DtstY7f70lzqETFc0Z5WIEwsj52zg4xaO144Bv+
c8X8BpIwFXb8Ggol26c2ghpHPnaEaq8apSSsFoJGhoyumW7yu+E6z7Oc15yyqAHL
pEfpBWUwFIG7+49UrEM8dyfI5tZGptzyju2wfTWsszuJmIWfTemcJ571y/P/Wbt4
3di7EY7QW+0bkQvGzwLcrcfYIO/Nig0p2JH4cc3BEHOMOe7CXmcOSNpy+bKxuotS
oh8YZSgw8SBsGwb4i0R+h7e0wQTSCEAD+9eHxEFcqZ2tPf7zYNrK/aqnqV5JycAA
cw1QIarvwUgXITsz7YcVG53kdbwdub0nWJw/ZOCKMsFIKPPOEzAWdMgh+xdrsQtc
5d7DXgIzGKMFkpOFUIF/GYc2sXCP4FK8RYowAIqIDgBVOJ98/aY3Mt/fJ3e9iT0z
7+rTCfCmTmI4UF1rk0MSxmo/LWEiuoYHNer+rXQfRCLNpJRdAR/2xbQ8CF3icnn6
Z9B/BHdPjhMakkkGkBoeF2yPPYtWp7BPgzEFl7xaoxeU1DJ/KnYscheGNSGnJJEu
Y79arWgzIoENG3lpnhx3ou1OmPOnm1Lqaf+fol6xMhpNmk7uj6axttCywqf/XzAz
23k27FYV6u+v665NaQC5kR/zByFkkmeaA3j9sQLHpWpGlOAnsE6kH9LPN7ou63ov
kawAtRjKeqrkvgF4JivEi297/q2P8O78Rlp8dexDHkI/B/NKkLk1Kprt8DiKIPJz
`protect END_PROTECTED
