`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7o/r/G/puKTJzC0N506NFNVOuT35k5yLz34+x49L/p/4AZRhOLzs+YlC0qxEpWyQ
ceAK2yTIgSexb7cp7ASETA1aD8O/akk5RTQ95ZKYWkhHGaQzTM0mB7/caT+BP3m6
KtszExhBqqfRc2HiAByt0YvckF6neGYmEmDSj7xIkgblA3nYkacUjQf25sEqJgs+
6CAix8KnZczHC7Qju9ntcQ49sQjGh+LsZYTA1P7lcou1+nHH4cP6gZ6KuWFfeB3P
EgFNv+2Z1jWCFGOjUZR52wiKuPGXiiwUprxVGofnjdRoht7MjUEMJSfHnyuiB2vO
f2tdFvCbVzeTmuFsFxZPcNy5MXcLFJDTHkQPHGSxk2iWWjxQv9cMbFVo/orp1QYe
hSCV35Eb2t//5knARZijKm5yWIGP4Nbbp26P7RN07sDsSieBJWiyyegmaAGLeQeO
oVW1464khx6T8Mg7yfWDFNXsiILROT3+0WqOtrZYKsIYEQ8PbsJv/wxOFajVtieU
C7oKm2nFe6Oy6fPwxq9UkYnCtGneyHRonACZ3Xpjv726vZ12UdnhLE3UxjykDqy1
wbvFTqaNTO7AbOSGWBbr5nzNmgwGA7S/qVT18Suv2hcftjyCLCyESagBBR7zecsL
nDgOX1DaIcuWcxocYh9gVOhuVhwKsMCJbfqdWCttvfUWc5wYTiXNDXt2zeh0baGr
RpkQAXyfjnhAVu8lB+VcoE+LTeW0WV0j+hnIVE6SP3ev5oPxwYWOvvVV41bC/fad
uEPk7vLUzgdtEqwfm4dpCEFbfZc64mqz/PyHvTgT8OH78l9hi97lQ8GPGbZEUkZu
VCXAEbJFwdMHm/dI3lXxr35ToNQFRxsFgswLiukEVe79q+HOv9syObDKCC64uHav
NmxbBc3VOLUGj3987qciFbmAN+V3D+2Qa9wOsmnB2oCVviPV5SZ/F0vMs/Ww3wcN
mMNzxMdmvCBByN+n4vAjnOs/IH0lt9VadiD/bqZPORjA6RosD6WMyUgyr2jJ1kkf
Gxo4cvsMAcvAiRbnlQhs9NQG+4CRKbXVfR+WveY/kDXbVehELrUKpT5P4ZhBNd7Z
gi7ZGxqpjuCccguUWa9mMA/JYhNkfGASIQRJ2XVTI0LcHvXMbRUyghgbo/IvJMnx
pdBHQkQKrMQi9HSgWDG9d76NXTD+rarNpB7tjbe94GenkjVkGLMnRP58GN6a5Sxc
sl08p4KlAnBtIjGEEPQ1JgbjZmdDvZchFz66XJlWDwb2H+Vk09Us7qK6kBXFF22p
G2wqs0f/wXpJ3Bx0l007/c01em4hD5qcoOZjU6XOt8xl3/Kta+5aaJ7Fsj6v/IPd
8nb7gIPcF1ZCooiVjtDJJ5u8ZhgTUl2iMZbWAzSNCqL5RY5q0Da8sRhjYANhP8aX
REkZZaxT5cO3odzf/Uro7fW2w+eInUjGVm5xe2k0kEwTUtQkeWJXC0of+lYIOWjw
6xBpISzUTmv6xmDsOiaj1tOEnWs7ga8WQuxNhO0edDZmFJQ0G9UtS6C/A7LJzz34
8FI6fAydAhenySkD2bD1Z8JO1doU61DV7+YZM9wtbIpW+ZfK94g2QCpycjyCrfhA
BjeiJc6ZNkmNqlW2JceCQtwVWmYYuSzq1xGkjC/8tzbnSJFWHMo9S5V56B6l+t/Y
NNj3Mx27ad9IEXTre4YHz0OjDDZjYPEqJM7OM8k9IverMOimwKlrXrlRmQBVoWLu
bzWHil4aZgkc7EnB6YQN7NQS6PPLyyznQ036S77M4u/GnjEUs1q3/qKFG7WomCsg
MoZYpPH/pstOviTFs8CiXHGOULrE5H23CjDTll7MlGrbWB8i/hoO9o7nv/Vyjrw3
3cKgnFjXNSgcEQDKYK1p6yrP8wWQ8iNDtAGeWFxslsnKowwwAtMbs8IzCuAo3zmB
axOgn7wIqsjR3Ov4zHXHTeVP5k5EYbxDixAn+w90EHuapJrwd2XeigaUxpOsBsnA
kSSebeGuTrHbRzbk3ogZ+Igh0lbsY8V83aQ+CbaU3ex+1jsUk28K/wcj24j3F4Tn
u63KiCSy01/AGmoPBLRxc2cBMSc2Hv5dc/R9bH/SedjgZsiwtB2VER/26gjvMyCa
a1SAFv3hjLluTIouM1gWDGRwXIqiYs6NE6jLqxKBLMcm9BgofVSLYBRWgdjgRt0a
LWsnyg11M28keZHFwZfeiRl7zKA8lANrxo0GUsFSFL88GIurPJG8AlXhNlD55ZBg
mJ9bR5yrA9AeudPw7v95vkl4WEy4LU7uSl2OOlagKEdQcEO5P2KASRtTA9tstB97
Gxm/xItod0Oai6/qR0c26qSJCzicPelVl3tj3UvJ4UB8wEibudhicN47dcVAX7hE
nrotGECCS+Vk8r8tqSlOYIhJVyUZZPHDoOelmmZB4VlsGL4lSdHo1AWbFfEBczUc
0ULbsn3newkQ0p0hPhkbb19j0LtVTnTd1VIDQiBUQLcZQ21rcB+IMg6ahMLWW6CT
7L/ekZ5OckoWo4/KE/3sadVx6/qAza3M/maipUg/gKTISfMvOdeezWh3PAN+faBf
BAb2+SjtnBJyRaRWYXDlUC7FEopdZaTXjz3KS6X9iG5qZ305LcKFusFeEg6CeD7h
oDyyaY9Mgp1JhZIkNZZeMvefdTZtEoYjZBa2eA72QbxNdJAJFHTq8ryTy7zmq2Sg
KqDaB3x0AwLa733bgAB4Nkx2fzvvR4nebdhM+hl4nwBbgosjl7G7/C9YZrIhrCQA
FrOTbsSH1I9567zMHQg2pN8RcBSLoW3p9a3D3MV1KBg95agCf3aLUSYcv5EG0hEa
8hCuCjrallqSBlH9xdx2hyG09Rb5gotB7jn8mFlu+3gLPg/V5HPmpS4k9k9HvHtX
vwlnyWDF202IFtS4bbeYwhr6oA1p3jmNs25KCXdJ6pUUDfI7d1Ccm+7mo/zXr5Gl
sq0oyc5hJKti+iJye9NSJMBMJf2eoqsdSz4S3e78iwmxw9WjG3g5lGKBEYpS+Nru
01Fo4eCQIaGo2q8de6pCtftYkgCyS8ZOlF0oMH8xiDstx6XTFL55TQpCik2IGM8V
KQuTEquBHQ2VvKKtvVODPQvoljPzLVoAeXaPcVSgHWGtcKEFwKksUh+pwHgKV/4R
1XNiewdal5wP/Y/ydV7od56hSUTXO17eb0mScHEMfXM/9Mk4PQl1bvQ78efxy3u9
SLoUJ24YW2iuhoBwoBhtz3pT5aCvx6R144CXUejOKThNRU3oOgV8wn+154b+ME2K
kpYUoaBDTD7doFQMSrCiIpPKwXQpep4bC+KYsusdi/tmEwNU5J5qYkHfm+eN64F9
oZVGLBDVbL/b6K3fggJlG4KHJetloJb3T6ENM2Ffps/6InoXEX0P8lLklNl77eax
siTEDmvYApqujawxmc9DBE+vD2A7lA8Ap3vkAyGwoQw4CVPSv75u2g8ld8yqG2d4
GdAxoXt6k8clyH1L7FCXGA3WCylB4aHntVx5w/b9Ybemx6IT6ENsUcxa0aTs++Pj
Zz2kozPiHe4ufHPpbuen1v+/b4L3RO1GkIHwBKZ2x7wECXDy0+8fP5+qP8yBTqI6
+rfxcDCkKc/K8fzVNe40dAVn5d7j+2+Q8BqOcRvd+mMER9iyhPDdi9stFozOI8GC
iLsMrc2wou1Nr0mtLiip1DB81pD+pD0HMkF4pXKiQ6tbbHzEgwD7HfdnwA6FLF7d
e0fwPfPYpaYPjh0Fck/6RTleUvtFfflLgJ6tbOkCvO9b/TPcwa+Kn1rIfwNQqx9K
AzNDuisvkwJCz0JRVQhx4VdyG5CcWoBv2bdRQNsu+rinuAhLj0MFf+0Z4MJflz25
9VF65nt0/Yg4D7n42pRaKA5NJjMbvh1aBTh9UgksC2KbwKfnOtYUa1pr5v5lZY7C
Sn/WtknbZJ5wxTmPqOoQqo7rWdZq+0T7T8dcWWojUOorL15EXAlubGbYB+4ep7Ne
vH9UrdiqmNPw1qWH6Ca2sODqU3z2H3zmxiJeJQkklb3DQ5mNpERATSr4Da30h/84
beVJGUaOlehr3/jYn5Fbc0o7W2i0LX+6ykhMAefSBTuBO/LQ6wNv6ewjUZ7hRyaN
tduQ/Wh/OTPkIb9Ek9NfO6mwGy19mhhIMGEwCZaYZXWszYopcEsz55bqGTRJDOm6
Q+OegjMVlO7G8HT6NMsJqVkXdxrhBk6ZS/j0hMqERjTrZfybrByAKkmCRFbfhZe5
+/AmgkwU10bNITu2FjGJ5g+lVrhFZsCP6a8epENLQVv8EnF/DOF9pMmy/qt01f4z
Yo0aTFm7kFvNBVFG9+wDuLgERyfpIzdKnZd4BQyzzE8ECeaOworSDKzSLvDTklGy
86rFm3He59ty6AueDRv335K6qzhpUDNX4BMtpolCyFhChyvzPFOIk+Erd0T2pARv
PjzobGkk125qf/UDZ6w7JqceFIpjizeCihCpzvGwuRLUyIYL09G2fJe/AswjQfRW
aeLGHZx9NRMX1g/ig4UwPxxQPQ2mq3YcS6mZYsuq9KkY2sQVFE+Axbt6r1xvNGdU
BSKUe0LuzWH2gtlSwEydMEyIaxL9vYD5rr5PRQa8tlooglTeF7xrmhvIreBmIUlq
7hDWYa0IExKKaRVZAhKoXxL6G/i1MdmSbBEEbSEh0K4CUiKBfVbNozrdg2lB0ZA+
cUAk0uOhiARUrhyhj8vFmpjq49CgBHg6IcnIqC57ye/2ViFZRVyVCZwnluIgFZ+f
QEFwSLS3B3tzmraxa5wn77KvPAkctuHpWxb21OyfmvpSoQLT9XPbsvP+zrQeKjab
Moxvam4DplaEq7oKpQU4iMOwv71F50M4ivIPA6C4+AK8OrbnPG1mplDRq5k6mEZW
Bv9Jchq/RQuYbq23zOd8ok+G38+klI6j0KObmmqBPHVIJ4tE8y68TV49K/QB1li0
+EC8huVwGtT0TqY2vniJkiCIWewiMsTnseFs3Zpxl6JlW/oBrWOjZYWFp/bVomrZ
KwNcJgPhccHNczIYZLScqtgbyU5XdR5cBoEIcmbsrE+SptNSyALK7g9tQNdrm6Lz
yOV4pMggCanQWOwfMQpUC+rZXN27kEanK4L/47S3r4DI9N0CG5+zct9RADLrB6yx
qRGt3qmErt5xQzLjvrVkK6vOFhjjwWKOiIFxFOFnElQ+Nr1zP37+0/W+8CcEei+f
n1RoYuqq00jUeOIfeXw+o4Ri6ene0z7+Lal40dhyQtbzqM7hIKjte1sgf6m/NSx4
W768iOY8xUSH6lRM67Akq4AKTyt0jgpsmJdmR06ILTnPOxaMajX4szFoOBEBmE0r
MNPXNA3pkJms4gFOZyIyRIpPK7LOzxTiD8V4u9TlhcvVYnobm5UIQrGt8o5TQe6n
S5kDX3m610Vi9SINgO5aNM2AAoCJD5KFA7QADxa+4/C36YO7P2WOpVBeLerFgxon
ezUsI74IUCOFg1M9lGUbzArxsD48MmFk/hDPaJfksW0jemosh4zOhohGS8Zu9RR0
ZQW7U4as9LgvIyW9MkKQyn0csFrkTEUAfzgddpsSGePUVZYVZ1BJpnISOVsgntxr
sEAX4U4L6xxRa3P6kD9w4Tmjn4GrsQPmtxRCfjNRGvVGIhMebBBx15Yr0SfRj/M7
3Bch0sV111SXOolC9IzKfniYJZXhRO/besjS04fQ4BPyvwc5Aubc7JVp5BjAjswC
bqCo/mAkNnB1PQS0B8r1xLb981Xak6ONsh/IkwSpGbJDc4xN7PcvohgHjEZ4a5CG
GchB3Gf/D+eTV+zdNsgZUh+tMCeflUpHNHZd75T4nIB8LoOHI2GYtrVeO0I0sg6p
0NBjP7Xx4zljXF5/lj2rFbLXuTa0B1542E2jGIC+JWAmD0fzMsf1L1ReHzS9gHqH
alB71FPWRqQZJv2hrA0GuE+i+GbjVO6Z9uxOs/SqNieShHx0y0imgku4p9nPeVjC
EgxYB5gcCjyN0vygo1rBMWZ3eYcQPX6kekW6NVMMjqqddjgL1NUgJ7H6t6mqBD9m
1buLOft47hyFg+5pJ7SCUn4aU/1yhgCglFhhGtX9K1HEShU9pcVv9mOnKy+nsDT+
SGxW3GBLUTYpw/AApdp4kiElPFEQ5+Y+2DX0jmAA4lmnGsOtvrky7wS1hl6uGHWB
I8pO2H+VKZ5BGQxFNt+Wta6yM2jIFu2mgWc1zwnxqa01sj/XCiDyrnKeH8wEyMu8
7imE2ReT5j7ZF5hPcAvT41I852SCIFMqoDlYMMHkI7tXsZoM0Axt+rMzRiQg2pty
rgQlhXJmPi6Aqm7C75H4RPLewjt7iUVvqeEb4SlLeNXjijscayHfEIq5pbWMPBO6
Aob17cKoDupRHD2M4kp9hZ9oHL1+Z/qLp+baxl1vY3xYjqCRjSsx9dWuwCneAVX4
lIKcKmhawOfVkXq8WfoBXZaZKSFJ5PXGcH1UdXctvT72UU4oXtmS3C7dQcIhwcUx
DFB2jCG1hxvlP90LbBBgxr3DtLVRuMGlihbS1FyZvdvqGeJJ/8wAG7alfsC8Ssd2
olsphV1wLb0PCoBoc3bYf2rAT0Uj9FiELNSMIxnizM78XzxXeJX8NfCrjf3wDdnk
c2E/bDwMfpPm769jQgk4bDBTJVADD9i3789JFmBwDOppD0B7Yjd2Iv4k4zsnrwOs
j9CC+MX3Cjsb72P1cBsdnGqCxBjjJIX+R7sD6ux/dNcmc9mqmovdj4l7RxFn19xI
1113mCvSYYs9J/XV+phnHR2jq2nOFgoVI2PNeFDf6xy5LDtt07i/bOY2YSAsy+q6
WOAQDijBmT+lOQcXxa/UQeHc/0hySbhj192q7pnJwGCqs6MsQ98ZIbsyryTP/peu
FVNSEVbwhcOpx1xnLSeWik9UKdlknCgpaEhoFRZWbxZRPDgTVGMlNurds5t4WvlF
NLzUiTWZmpDQzSMrVtn2vlBrtN5aWjdM4s5rSddmJGN8Q5TbjAlM/nQhUqu0lIYO
cwDxRHadIZ3ReNORre6SZIqy5V6THV9hEXqUuXWRz+ELv9kyqCr+BCs4SsSKLB0z
NmhW1S9nZt/HmqRocUaPbtlgTgNiq4BoAlx9M+p0GH86p7Nz8B9q0TlQo55amZ3T
MgT3UN8Sltuc3GJkS3Z3Z/K50u45hqtjHOHv6+WEbcf5ps96za2ll7X61wwjWVtN
MbU5MIejpA/USSjTKnIxfHBGgmGnKD3frltCa1a20YqzRjP9E+xRDWpOwMuCH6rO
uCSaIjxvMRc9JsaZuEKHXqRCttE6oj1q0aLTygBDQ3zQkfcWA+B2C/yRQlLY7vTM
79fvfQlqrAy0OlyiKFJL1S8vJ70r5fBuhx/BLeaoNofbZd/7XbMuW2KANkFb+Bjm
5JlpaYR/pshTKQJVQPlilzEEIlyyp44gJJpZqHbjZUkcsSjcie2ySBwheKaaPxFr
bp/By+6e+x9LptHgIHgn1LBgI8z6PMu6UWTSvFwDNpemhIYR00EO0xihHs+snRvi
xI7L3wRvy7btXWtHfZGRnMrTcO/rwvTYdA4YU14HQXXo9N68CmFxJzwgQs6j89QP
caApgVzwiiJIMoECuZZcsM4PzDPJkAjtblq2ZJwc9Q/PKJ7aNBkViSSPG2Hg7Egx
FZ0QCpqcOIjReSgwzUsqxP1HM+4Uc7IW87EAtp9Axy3ATZEN8EUPN5EBjxcadibn
88bwy17SmQZfEG6p6ZqGIF9rOoBB0oSgXrhofur1TXZGNufF6OZxB6gVlBIGwiUe
UkCx+r4Kk8pKIAOzYuvhvc+WKDuMdEKwj3CvF9+HBKUmJasC+udV56voLrZeI+Fj
aqLH+RnBbLQX4SUSNd18cxh2hchPIB/ytPn1Ug+4ojEG1IJ2d7KnKYuFDqMtebyf
TwgR3+xw2JyhiGJaoJpbF+8TFiuQIGO7DvZUyYtqhwndHyLydMnKSW6nBCk2wgRA
/6lhBKZSb0+KJdLgydN8Yv7iIv8yoZKwPISQRtYl1vM/fuGT2ymTG6XTIN2gq04e
xppS8Uke5B0YQTnh7iUWgcEjws8inGeNyhWZQbpnkOujCrcOZFxacyvUZsVsbz+d
XXpBNrqCuwjoYq65OMbMO9QI1X/1F88r7zP8uHQQa357U7u+/1EK2WkP3zIgc1Ue
8ekDQ8Ts5Qumm6ly13Uamy169J89AWkmYkiDWaaZOpaPKl1DxQA0V+H567nI/k09
L7qFa+gHY82K2Xa2TQ9qYkS/R8FD1HoX1+y9fciXu5WF6VjniVHSwsaC+dsvxdq7
Gug9EpnlfGCwaa+RofZsZe5amp+vruEalEZKeZFePggYWQganff4VI7OsG6nTJh8
FC/PjTKq5Rjy0B673RCD0KI5oyNNjYfpT4vkZbVA2ILCXjI3R1bem1/4xEeCi6DB
w8C1awOoKMcpa59aRZ7RaSB9sWyDtWeSE346EFhXcSvNtTPYVbf2Z5mnCojqGHas
+UYEwKGcqi5pgs+JgZlAGtAp1jaL4URC3TgpuU/W/0kYsC0O+uWbSHJB7U4r0YjO
dqk3yn9WM+XWGY2EqINnRw47cT42kFTziIcVfnIIgnsT7Z1iwpLGU97e9nA1AhW5
cd42hQGKtr4luLJJqgzKiy1vzGpnd421wdK20Ow0KNVl1NjHb1UBGkDzltDXASuv
O/LtXpFVPlcAQw0oZQgbuUU6Qor1SOD01lvZSCarG1o0kIHGfnRFBBJLyiOKeIcH
vrgN93JdCIL3wpljm7zf9guO4qIxZx/9POvZOlVtORpHYDTbbd75yOxO2hMEoRqC
R3N5sms++UnAt4/FlTM7w7vr4pOgC+88CYNbdB31WhNwZShHXYmIp30D47E54wIv
zxDZrsKC2+nGJLibn+h2X4irt+RE8cIdtFp/1qLSi4Ffn49U4xIqGafIgTU94fg/
6+ijBnLgFIIhj5DotKGcybtJ0w/bCFEfSi2Ll/zgnd8AGHPf/mLxJIS1jscxWvt4
IcCJEONCNihCdoaGniz4rALqaFpz37ptncVt2esDTQ0/KrV+dmx7WeQ5a2ScQUnP
LR0rBa5GfnYZErMb0SB4sUtRRpC7V7GwANODqTwbKGXW9/m2CBdi1vkfYxAfnDj+
+tlq4GpMsNRMPpPB5YHCd8f6Ousrsu57LF+nady7mhqcTaijFa1ZD64MO0KPG2/U
jztYuCmOM81AD2qeb7kiwmeP4u4W0H5op/a5EneBBOhcT8ECWCPbZ4ohdqAbWSVF
g/pZYKZTRdey01fmEyt3SZZEpRuMFQ1CnxqkEEFTWkqOIa9+FvelEWmTuWWbwZqs
Ar0caMMQyHHw/nw/off6pw40PAXSh+pOIgjbcA3HbKGes733Mlf8tLNo/5mXGjwT
oSSxPplxJU5PSrXYUMrZ55qyOGedZuCX47dQRG9psm8Hw2KenzXc7OjvoNfFd32s
tdxtRLEzcsAuV5rhhGmSwgzxDW9fzteqpcb7UgCUBev0A/Ak0TdFAD/BeIL9bOyX
iaFEEb5Kt1qXuy5e4VtC8XQcQUAFIYxxtGfAndSwVDwvDRhhbqQIQWR6NMcbzrx0
f/9dilBiE0yZmuv7gO+tQqxAbVZsyIs6iq6dffONLrzWZRBaaGd8CYNpfi31u6uv
UT8pAK8qZc9R5Ag2SvdqrUA0Hc+TUZ5Vs8/+XVy2feO3dT722RdElKooFOToW5hq
q0rcEh05RSUQaD98lm9+aLpBNhZeMhWAiFzsg84C5Em/gCxOTO5DopBuGrwv8sn4
bjOoZ5Qd0HCLSuW0uF4fsvQpmBzIei3N0nXb5SMi+3zKvEg3AH5Hj/AKfDUuYfo6
cXd3VDNU5v46xCi8ZPzXQ3sQTBZsZagUV830zAlnjFCvseSOVG9vUkxZNyLUPn4s
NjadlH6Y/peQWWjpAaMQCVx02FuzLhAzwgv8HexBuysUDe7dhZsq6yJUGsqoiBSJ
cSjFcpFEQD1ORQs7WbMMF734mkX006OslDvTSpPO6O+Nq+bcPbF91KRD/vA4kO9/
01cSvGwub+ActTo2pavOp26icDDhteSzMMiVvtx/w5+I5OnhRr8LROWN3/dy0dea
TBJ5Wfo2lidUZ42aCnI0NjrVnhRQWy0nlLlbDHYL6hgzOXCYx+MmgtRu/DsTP7Qx
o5IqMW0iSFRevP+91g3xiDh5U0HR0AFgCt3VxXzzDhkjstNBks5Gzw85e3K3djTm
YTnp+kVDlvGbBY2/jsKyfmj84LWPCBWoluQpuAjVwW3yE5pinCPs4szVgL4j6n5L
EkHqMA2V8fQUz1mC1dKmFoESQi6I8tSN5QCq5pGzb6NcnRJJKlhrZiDPAkiA7/OK
B5tYxHB7imsGJGKIh6vZSd4hkiMQA868HAXpVz4r12QDmRw3yU/0KpQfOtL3/ZpR
mz3+8NWWaKjMkv3Bt5GXQNfteMp5D/FWam3vNLs79534BFNlJzbmhYRN/0BOIMMc
JyoUJP7OJhs1Wy2Trdc+/iyOWHwBK30wInMENqVntEEDooXokkaLYXYfWH2PtuXU
EJWNaSB8rYalfHAnCpxaJwU+jrnCKiyPH6VFOgrvEIncOnMGp/vHMw27+B46Vewx
dpQAFX8FCkctb+r33KP91OlBx4FsPUruX+RF8+4eOWOhmLvmY5CVhcGLfC7m7ORy
S9x0gz6H33PUrp4pgniPDBnzsH83gyPzgc73Ble+PCwBhjdOppFjKJf6O647+Kga
VhTG/nUpIHQwYkp+t5gl/i2X7paaxKfCtaY/oie/jGHjCVeImM/PGErX+Msj6iKf
L+LDsLi4UuIUeZoiBH3TdSrasnTo1oLH95kvd4lsWwCoIjVnjXGD1ENq2Jl6flUV
e6EAy+ObPl5u+8DDOrwO6IzlJUlSje1i0p+Yn6V/EwUhnjg56LaEPC1DK4f1Eika
+7ASAeTX9XbiKzQniRb/aCF0yCr7NrpMBqyQxZ32lRmVpByTCx5qPubNOj7jgrFU
fRrAugPOwo+t+9a0utr4MmXc7sE+yQ0VNKZhLOIZ2sUKDaZmXWHiO/GWXqZ8NzDZ
yFb2m7iJJY0J9UtZRCU4AUU0OL2J1Ix5oZAMm6Py4QPiqHFGebMjThYKLhN0salV
dDzsf1Sv3t6ZnfL/n4/ZgIxbyMZtHABdDyRnwywaoslD/JvJStGYegmLfz5yl4GD
bg7b9U93KjsdqJdCY4l5pvEG8CnKNjMyp+wmc6GzxbBzB70V8VskF9ZhTH1KxNja
deA0iBtZNvySnZLgpDNcPB/CpAY8TcIf+Li2yVMeiO/JqNbSlEX9CouZXM/GG3vv
vSbAUNaEhfp/tlkC41Bu5iGx95gMed16iTPdEzf758zbJDmU6/z7hjl3vWYqugU7
azGeC/F0dcGg1EPLtJXL6lO4Tf3GTSphA+FBrWYX0GUlxtEo5B/sPqyqvYK1ifqF
AERCfRU9L1HSkoQUWfCBN+FRKLhjykWVfc64N9+XsadWrAEnKNqPUyDXeob504qP
emyLuv7DQ8kqBlrCQ7yWaXatZV/O1WYamtPb6sUwQ3d4N1mf/anKDjO2H6+qjT6c
7H4qrIQT9lIx73l/Zr+sk7YwDnWZe8iG3EiFG+pdw2fG78xEwsAxbF008E4XrKfw
RcnIo9zqEVRVoZKpHIClBbjFxtUHs+fVoy5D8oUQU3dlKp/K8eYf06ruYqDO/X8/
n4U8h06YBmDZvTa+Jv44BlHwumC5JWXdY/JJ6JBVWD+Dia3JjoQP7ZOVceoV3wh3
28JLn4L45h+rrtCqG9ZrVOdFQLKYa3UFOxBkU6n8u2AfpnYxz6OR7m6YBhdpMed5
mgLNPFBQqHSh/aD4BcxNXpmV2WVv6/CbJrjKWB3+xmDefQ2CL799G1jvUdp+dfHD
d7dEOEhg67nSIsS/Ac4zcHt5MZ/TycRFTlQARxu6CpO/fnIbitQZjEqnGnjgQCou
aTjfRnA0GTekyAVuLV/jp3cPQGpNe/IIhwV/irLG34An5YuDi0YG51Y7fsDduBXJ
8unsaPzcwA0FX0u6OPoymHGrYVXgo7KKcIZg5QZRgEU+tGSjGkKUd5FjKy8VxliS
kYUvPkJG1dsVfvi0A5MCZhTnKWQ9PJV2BJbQyyRBQW8wBMSMGvMTsBObjWGVoxrr
NFz4JSu/A+iw9vID8GQYJ4vXDoj0FIe/CnUlGpn6In+HEgbm7g3d8CFi3MdTSi1u
Uh0V6+2bswMogVzW/vr68iDhgKaaSjncNDrSG2qBklGXz75JPq8Vm7ua8/7THheI
NppRp9ykl5EIYyAMmzK8T5NGfuqTMMwIsIP47AaC5NMo/r8YVs45as6X2QKRZ2YV
vAv+VGgXPsNLaaL2WKxQkvGDypyvse88eSfzZQeeSnfYWomVGXAZS/bZe0fCmOdb
JUjgVE3GtgybW9WSkyM2Aglt1iYnFs7fNC9XTsFhaz4nClqi014cRwbwOv4h539u
LoNjUuqGJ3J0SV1DjyH+8LszWyukAJbsgAxHuDFdVnzc0kHNLhjxF1SgJ9wSyTaE
aAKLkV/ii3WA8zOS2FaCQ0/cOIwhHEWrF7XxsuZPJPUzQPMakvV4EQOdxZ+Nih9H
vepa+YshhhpKNqM/biR4lQETRLp87V1txzETZF8lJoTMq9RWwuNwBC7PYiKDbsVF
iOU+nZTUfJ89xsGrmCR8MsVO5QLCjVj+tRL06hDzRfYzzYs+lRNr9PNEZALlyhKY
6W2zgiJiDXWJzL+tyDf+ameQ2kocyuLcnwedZ9Hr0JN5Cr3t0QS0Mb5c/+sOx5gU
C9RwWBNph44+vWQIQ7tzJFil29MVLScwUt1z2uFYMWcbEucqpQhA9zexxUwTDGN1
lnZOx21wjySPl7arWi8aMG+7Zc6SMwTbW2zLEc2+CWi1dwcIpYwBYWjUrF7A4Urh
ieX/Um324SSUynPYkryh9LFfhP8l/G6J6NlV4mZTQdtFXw2PFkw7tfusSs8sc7CU
VRvP+WCJQHrB6RlWm3VPfBtKal+kgWcObskOfXrg4QeN8kv4WHptIx9CP5socvT2
IYZ34dRx1ozIskCmB0gdyUwEUHP0PZyjwnOCFRsK5pKjNsjxVRmmsxFv+yyPDZGB
KacjAs78xhrRrfiWplIe36+9F5jd47FUelddbs1P9oLihZxTmKv1MlkOK9NGB7MX
Sm3NIHuc00aH63/L0qeqydLXmw8ebTxt13HoJJJXkBl/nyK2KKE3pyt3Qk3KLpUU
9YFqxn23Bg91dXXQszjdgfUKxhh6t/SXlfDXbeUStWMr1g2zwb+GfqE37sH3cIj0
DGc+Ftpj4to1FSeeNVaYKGol7Sp8DuBB86MIXCwvLzVMstBG1wlhsb7k3xo7DgJP
D7yOkf0mDHrdqWuzzuRTHLZpKfH3hzuidPL7PHs20NadiI86hS21+frnBPN1PnQw
Zj8TMLFxbFjQ6Dx0pSF+GZsbh3/ChyG43gGP4fMMBhA1PDVIQ2EWA6j209vPDh+u
fe9irMZycV2VOobCApidhcddt9oEh0a+QK0OiN/ZzXoXYDncF7CYYzO6m7hgBiWD
Zb96dOUB++zhQpsXHYzewxoyzW23OZajbDJ+cztBQxlQGGiURbnMHAh7ibiQGwf6
A/m0CeD7BHGIYe5MFb2l7hYZ+rMP4TzWnuiR9308h82uC2Vy20LXvBL7cCybydyL
QYafibzuS6+Lcd1lCcNbIKjbGIJAdrkJvh7zdChPplcsqTQeDwJHmB2ix8yu6aCM
NaoSbPBRxBwi6NlwIVPGcR/Aq7o5OnKwAfLj8mq0ecgh7NcBMOb9eVXFYygPXk34
PDWrGYTWQjNOgAFyFh6rCL4xzK/WRj+V6G9BSGOUOGohSFtT0JLz0a9nJO60w4Rv
oKzhuQRIeo5CVw+aStvTplXxqJn444WqeLMPgRp1kuAa66NpfVIqmKPHIwxHqcVp
Nbh4d9Rc4D14+txqmHGo55WSzkkIwUj8ck+K9tkxTbNqoauEYkmo+nT2lD8zgdvE
1CLouTob4yGGrcbnuPSLNVxhNkNRsY9bgVvRox2uLR7iLivzoVMzD9iQzrn+ex6e
9SI2iVb7x+4sfbzamffFrtmaVq4qgn6V/VuIy9zt3tFVQbwpKWVe7BqyE1QPk8eT
zcy/rV72LaQ0+TTsdmTPXwOjdVticCF81RNz6zBA1FFP6qDkJN+whw2WbHKM2cld
Jy6YuU0W7DkqleWvE1CK6ocngHMRBTXlc1wrYwsTxQmC6pnpNt8H1EGu+k4F6wir
7qEgoXKC25Q9SithJ/kzMkIpcSKDGumNEGZrYOhLGmlhoIEbdq1CS1W49br9xiap
xBFdQC6elK/gJIKR4OwFaf+8TNTx5Xoa99UjuQyv6OMAFYd7TeAH3j4WnPwXONJj
Yhd0HKMBWV/qPoJPVWt80DEtBZ9dCmfd6H0ouHdkgOX5ko+sl5bMWIDTtr/XrJuO
Rea1GK2I8cHXkIqtUCkojnB8GbIg7HJPhYedfu+WguZxZy0V0LR9sciYa1r7zTLc
WhV1dMxhsXlRmaAaF3l6DKJPA30I+03hI6FSKs35Z77UzhqWPACtXtgo+sgEPXHR
XuQmbGuF6wTQ6kjZ0rQtqMeJrklk3pZcb4Oe5uru6zY+/RAJT5EhtlXHKAP9KIhx
TEamcsbD5J7iWt2cbhQk96B5VzktBZ+h32SyYyuH+mf3W7ppAcbKAA7qNhGKVQAW
Khq8a6jSGjqGA/C6+0jlb7K7jEqkcV6nO3+iFA4YxQTrmRqfN63/V0u2CUJeZJuW
We4hBMPm2bI/87PB/o+eKCCgAyNU9M5Uj1iyB2MBLZvYo939nkTvrASUNoL8Pjq2
kLuwS2M40ZjWSOYTwtUlKhHvzmg36LR9Z6PShiMkEsJjHRWoznNKAI1G5FNmiaGL
8oHlf607f0uKZBDZUwTKJzaZ+azuAXrDM13LsqVDlv70TyUmdWU7b8q5jYf4la/r
+K16yWFbeyJfh3M/nSndv/M12K59XqBZFHNvydpa7m/jWOW7RPC9a1H1DnLyacJS
C30z7ENj67JfcJ08YiqVE14+ESzkddLEi1jRDnzuhdbw3at8i0T/laGCf3iCDhey
6fOtMyEzuTtvnwR7khKAHkpjeWkrcyYiRTe4Azr4oxjRIeLGZ77X1048ir6g7wMS
3NiV+FEbBRY8x1hDSGHqplSCvqXyV2n7B5ZcH1AYWHKmeahnh0v+WX/Iy1o3Zs4s
IBf0D6OGHLtG3UXJp5wyy/boaVHp7/I3aRSBsXDez2cyPMXZettMzJbUIhdo1oTN
MSFOakrtHWRUbRY+A09uy/VjTq18G1HbqD1HjNrwYHJJaplPPSMnj8+fWaSYbXN1
xlGVsOaBdEzmNF2IKdiKorwhnYh8YJlenGf2Csw22/yV+VD6T80Jatdz8A31WuTh
iZk12wHKyj+cSbk5uJQGnX2SCsBRqIpBJRvE+q7DlqBJBFDKTGDQY7ytwaO61Fr8
5KJEETrDsZvJTejJWLawrESkORN6+Sl+lXvDRfPAZdzrbZo2onxYPOF+1Hn8rbM0
LRi15Aj/aSTafhvzBLW+Hy9JCuKuz2hmRIiWtagrQDpEHFWLLVi/TUOq1cbbhPrD
jqweh+DU97hs+eBC2DoaNhvUQ9cd0+FX/TgYBlg3Ud+0pDM4ochNpeVyVN8UXjX3
zFpdkh/gMKlulwQV8fIuToBDYvLu+zGYsPe1hU+0VsDyphghSoIIhCdp7bffSeE0
vdG02o3sGSHU32aIhhcbzYyiGgFhhcw+8px8f457xn4URINOFLWT42C0xArNsYjd
DHQLX1RJfRo1VxxfAXUWAyJ/gmGbKFLyNGAkvancreMrKCbHSV0U34KQhhSUMnIn
si1XjTfkS2XqW26Q8/sDqDjZAnBeim8HluCKXOL2req7AEinzSHmf34E8swxLt+p
wSUJHk2X4l9LcM+rIepMs+tojcV+Xzd5Ultd4ELUVGinME5fW4qpWDsd5MR3wNqD
efDVV54NyZcOYPN6E8QQDMEVyKO9aWK7aZNyKnVOzZp8dh9RlDItFaz/G/5p2UBk
iIDHAKHPKrRwm2l2jhCqbCO4Akm5f/p7FPJ6AeLL0v5Vthq5lk9LxYjegePRazqO
sbdzIMEpAIKdCld2H6qBZEbTM9ST3qSR2A6utxnZGpiVjjCfIs+51B/kRj+qX+Np
/BzLp0iADuyng+Mr3jgsEcxr9ujOTfZQadVGswVX7MoSTromJN7cFQZb6DpRfgxd
yyfeA5NgCctYQ/XLIFh8g5OwbfBKrksfSfdAe4X7N7aUNU3uZTMxVX/g9wrUyYlH
U326ZvAAmpuGtaEYL57jzMDGzDYgWLc4c3GBtq1/TU/sbUd9vTX7bltbMkpDhTIM
oBG4V/8HpnEsfA1UeJgsjW+A9Fn79dNFtXRh3X0TdhWAVf1ElM3fRz/FnurT14Nj
wi7ZJg3sIDo2sTRix1xGSMOIK6gHNzo1wnocD1Xa2APcqCKVEY9EVQ9wFNqq8s+e
Nlnt0b1olba7RCu2FxsRYvCvrNIlORkKouJ/eGacChtePDI0UZpnVyWqeiXXr5Oq
b1k+j5L7MORDombS+MOuJuYcedCp0aRk7fSqP0M03hEJXEGaGV7SZXIxV5Ltepth
Ci0ZDbSW9zxCJxYKc1sgd14PQho20b3dULXDQUxfybSsbk2ny49q8L171IncNLr4
GY7IJCq35HX+4cTNZuTT0W9sgJ75/NqWjzj7vQjLawfkqu88VfzOonlsAub5Ed4y
1UpGmMfZt1zFjnx3MNYkaBbDBH5bWSJGQMc5kLTm9rGVZAUCXxGxFTUQqbKCMRss
6HN3oLv1YZrFQe2aGDtukwY2WPvCgcVEV+GkZMxC59qXMP1QbzbitFOIxpyqA57s
kOhewBZYAp8ep9qFDo7/alLRJzKW8fpczBEqS1uuOPpf2G7NMZBN+c2RR52N6hu0
oHsytrJvK6nLHbbBp6cp3Mf+//CIUZqLxAcf6PEIgVeJ2knZXcxcrBjtmr7cShUb
dD92X0vADouLw7+GYYuiZ81+TvTipvLHbn/8+DK4ZvY1mR/n0FL0EcWwCHuV0iXQ
FvjMQP7cfabPN6S+NdqsgAfE1yGBadBwzxhvr9vtZTeLPPRA/ZVA27Gdhj3dr85G
xGhRRYnJzTUEjE27OxL1M7cDLhS7CI/a5ahoQQJAvFeIHgPmn6uoxvcL/PmK5sNv
kATDYFhvLZVGsLX0vGwiwS71PtDhDanI4QSPcuy71+8cvpW12/topvdwlrHLtylu
gBjJYNRO88mCjG4pvkdSGjbOqMKbvE2kGE2pv/RXvSGiYwDgjbpuSUYfSIXEK/Ln
PHlMKj80p75v72oEvsycXkY424FkfPOSxFyJ83oxnU0Wdiw22aVp7y+gMseuVRv+
SM/Y3g51fjOo5MpmHY/gRd1l/2KFSTFbP/IvpHTtJaozkoasW+EEfkAb3/WSEidj
+dDbR2jXQCrN4g/pxS44IZi1U4UvPkzAhIIQQ/M+9LwtVWpenDR2iDJdc8B6+S6x
AQfHS8f8Ry5T0pTwpQv3gdCp+yyTLBR88sIjp7p3PUJQ/ZRTvIJmcir+mgIb7kON
91llaHiB5FQqAH9aZ2yVRcjdwBsO1jxEi0JEgivD9kdDwc8AtcP7rJ7Pgg9peWQI
9cttvaW2si6S8rDrLDORKGg6/hJqNLkPQI/1FwlTFOgbnkOZgwoNspqqvsN03tDC
sJ5Jh0Fau76Oa+6I8p3yf2hjCL+w4CdpcTwVl8+CDwsA5hOFCCxv462vfAtgERmP
jJI3YQyhiOd4E9QHBSX3LFVWcVJ+T5+V/WkXuoIpnsIJ/jwF4xLfVvHivkvR+g5J
UQJmWFN0Jb6CmWGmbA0OujATA9XYpfUjIgcBMyQfk2wiAQW9klwvVE1f8lyR8fQn
xO6rD+E679RNtT940Xj8AkSdAsPZ+4NX9rZEIOekTf2nMMFSMs42m2NGkeuZCHEb
JvbxKI7fUr5MuNIEb5fl0/nOzPeLoqATtj6RLRGv+/R4t9eFiqsuL++PcNBB6a02
nuohMcTRsWhok+fqdNnNBPaARCu8azoVnqrjVc/emIfOR4yJfn86v0CusN/pEGWr
B89XvvVpRkkWVHXs+bax+DxC4I7TQFBdH8Qcv1QDTJ61rm7rc3NyjGScVVxoKCLS
I7kBLwl52jp0L6Nk6rOWsbSC/ItuwMSne7X8cPe9XSDSfL1hEWcCp2Np6MrSaM58
8jbcykTNl7kv1GO12cw/wAa0a9CkgKAi0zgF14F7/YRWDl/ma9JCjptuIvsJkoi1
fZaWTfA2AHtp/S1pup5ORAkAX697fBnl0IHl4u+P9zk73HV4fOfEcaspVTbKZl9F
GjbVl27JNwPDerU+DRihziSsPAOPI1+DGjmD4FaB3Ith0QFSdbtmJMqI4SDGQUjy
h2+YvUw5XEPJ4xtKa/VgpO5rvmzC9zkrGIfAMxE50HtycC9Iu6Zoybx1IJGnX0d6
jUVX2lcJlB35rVKWKwhMzIIy4DaW+c7ZNu8pP11s3ywUCVi1MBnSIX9fP1huEwPu
nPsX91/Jhjej9jvhsB1NqQZthCv5lwk7JYWe2oBE6mtz86noBcM114rLqHz10vEO
6vEtsx8oxlUmzLfFGhWE+AXGPQGGQjKWD9Skwk/lkX3QyRcdPv3yqrPDQyU0p+qu
82cpmFMFP/y512xVX6ekvTpmv2AdjyYZz0yHIXyhraT1PcP2foX7egOGma0XPtYO
m3byGr2hqLiVjklaKywAosu3YG/CAjj+sPHVQpr/0bS4UhqoQagnw9arhN7Z8NFU
nmgxoaEXdsLON7gjxGelLHD+9S9U7h+npMdHjo3XoimnohsvAey+8Fr1Ylz6BFsC
b/58LNQWub7HY1uTEEnhQWuUHilHjgToHZ/++XY52HTUwzu31BTXbMnjOCrp0oO7
RUwWpcuhKmgKrPy6h2dld5hPRsK0a56qP6u7nXDLCCO0TxzpxpUUtk+QoVRrE3rZ
oCiFCw7V8MLedsRgwlcxZuShhDQ/Ahaoqfn/tdYbEbt/9vNo9rsqMFZN5KkwVrd7
OE22ivYinv5Y3rHRbq0rBhIsOOqIVIp8A5O1ylA6f/vFzOolXIiVFmExlddEG/0p
0hLzU6Rz5TDTMCa7m9EPgqbTZo+uKTJmtzj/8TX0UUaTlE/SCJc15GdSga2n8sMo
dTzJjaajJuiqEunJUpvKuwPpwW53sav2V7bnvajVTd8ujpUFaEEx3bWLhEkVqrzc
7oTkRNptOOWb8ix44HvWSIIawjlN3JlZtYicvFpWtFccwTCf9eu62qpRlzEO9RGP
Q/vEpkUXU7yz2r4GIzL/GOrvrPMNVL1hgEkAXeV8AQ36MKpq/CD+U9NdgYxddzdR
P8KL4faIHF+JGs9sjVMrT9YAmGXvC+fL7st0w00EdJ6i1B66tQpk17jf0lwB2nvh
HkzDdcT+sZTqu8TUmG/KBSiveEcnWsFPG069Hq/jBJL8KOo/K3c7AzDt81Q6DO/E
VQgku5kYyrtwwxLDiDHB2O2k/xF/uyz4UwSRuimyFskLiOheW6bmMOzxXXkoFKPF
jDw6dmm50wiPerzNWCir5q6YuXsPhyRVPzOe2ZafguJJ7gcjmYa2mA+nKHTzD4cl
tj9nmtRFKC97ImxWu+gmvYGRaqxZD+2d2aCedGzmRjvvULt8ULdTax/TC8aSWxms
buvitRWEasp5KAbPebzqwrORFSuItPh8jhwkWQxmmAXu3/lLsbjOsOpbJri22SyB
0vEgNswZa7WyetAJzD5jWWa4cOJpy0yLmeHlCeAx6D/p6Orfu/YNZzQwOj/THysI
A55GSZHh7g3w065VfAFLJA77LViZe2T4VwziZn4I64+WuJyBM3wNcY0eeYditvw6
+PgqfjYxqgZmQQfo9ntFAnXS+NjaiiQNY39grjXSYXmwQwtiKdVh9Y2fP+dfqalI
pN7OqsQsCgqBEyDFyL1j10dPGh79wRkH4APNbborWdqV/2v2BKBpRjrutO/tAjQV
59xnDdttgCPJj124CLkkIycESSJptKD2Q2zhRaOk1hR2uT6XEG7XBqigzncb+HLO
T1VO9JQJ0TN/LKshLkwmlKwuG03bUoPiwzbceGabYbjAIuiLy9Yocve/6xbIx51U
T7fBxlQY+bBZogzyCtz7ANz4uI9tYcQrHm4PqrAHd59htyLP/q2WKpB6yw0i+vfV
CO/T7Tg4lJQ8D2nYaPbFhIq5yMBCQKB2Fg6rw33cAiV/gENPrVTXPZcrmOUXY8UZ
Xv4PO8fCDfKwExAlXkQc44Fc7Rab4y2/Ll+4lUVqXDooAmofDIa52Jr8OJ7N0Aei
qCJCQ7Hs8xh69q01hKqn83qZmXTbYSbSoF/vfK6D9RUp28tx8GMV68hPlipeFL8l
gJWfiBTlEs2oJyAl26dMUuH6cL4Izmnuxrkv7llxNqBpGJNflwaQQx3XSDuJrBHI
3UENgSo95TxahUdhfBi5SmqHToLG97eYc4OXIFYCafDw4Su0xd5OArfOLBb19KpW
8J0OCZLWIi/A8mEqLpcE246X1NNy7utgD5STnjM3fpTOiqT5xEUD/0fc/z53uaNl
a/HgNSZIU3nQl9pF1TXAjl8BAKNASE9c/x8dYuN4AdDaGD1CRz0aqRsYplSDbAKi
HymTo3q2Abm2EIxKEfeUpoo3R+3iliVExDGzGgb+OYOjOxotkiZ7PfhXPQwMm44u
iGScFs3KDf+Ji/xsxqJWE4jUPts7QzwM61Ab9VyGOXopfbxF+1oVU964ghwUtFz9
X/a3+AXQzG1t5rPEOE3sPFTBMf9Cjy5E8W/pjCDGB1EXZMw6j91B3sV5BH76gIkD
awECbHgF+VlqfhhopX5xvTyM2wyYohwfbVTpIOzreIU/ysIH103W1YzgMZyVyTlC
gqA67XtMF5WIQPN5AGy/7Nn6VRlFCcKrQSyOwFGDNaTyVroSLYH6ILrj1jOdH3uW
2KxWweb8H8st9X1CnAPI9Yl5waQWeqpG8/neQjS0A0e9wdUR6ns4GmB4iR8vIZH+
uAVySHQpP2PwPVuo7FEVP96zGenOo9CdvSsT+la5qRVRpHSYK6/HfnO7w/xem3k6
yym0mSvJBmVhN24iu5fiyMPRFS/k4NeKUS8ZUrsapzYFmA8bCDgzR8607XERuFH6
Yn5gKOGjtZsyylFPGrdng97DITC+sqRfTjDzvNKxrcdHFtUjyL6aC6Kn+iaQFMGH
1unG8iKl8r3BiMu/AjSs7vlYAh2NTFmEMdWkrLSnHBMjMciZZx0AKWqGavlK7CvI
S+Y8vlGqzEbcmom+bwV8pAAhgGQRRCH1xXvr6JB+G85wO5WZJ68lXIKsHOJ8M30U
X0ODEZByAFLcBYtqGpFVQg3hJe1cTuXQDM13ZUtlcej3ZmjZSz6liiGS4hC9nxG0
Vd6zNp1GrT1AJ7QDaVZazwaB1/NczwbHIlV5aF0ySS/Wm/KDTiPWYb0qeuLTzSsw
7KiRXvGqTekaR6mnr+ufn8+/Eadbn1ZY3D/f5ASxTZyvH7i3JQFCdKZbnkpGF7GQ
syTTQwryJFYHBvxDxSExWoxXZ18BnMf3MzsDTrWGtCyO+DNht4cxbBJ1mwALfPXz
DBMzsikUh4LY1pKrtcFHhVz0JUD9gHKjWkO61Wm4tMNFNUT5x6/4ohGGgRUnvfn5
kBas+vsTKuOQVGaYLItXEpJSPbjisDBkcZOko8lddV4pAhBlZ4C/97LzmKQXkO1t
Pq+ezZ0A1pJMWdBovBsBbJU+ijaZg/9tuZAGM05eue3HYNUA0BV5kk34A6tvUhK0
yYBQfCwB1p2+/pX8V2IyjUCXYwf/C4r5UmWfbsyqYRLv5/y9kL3WI+q8DybnmOJq
zGLyhx6n3p84InU5QEiOv2KtrT111y/DIQMghObei4iCfgHzevDREu1Ac+Fu25Ot
KeC5e5NYCOGf75/DxljDXCRjd/yu4AtLf/HdG5JLUZCCOxeyCu3/0ZuQjk/vIPDa
I5nmKNBSgdjh1G870CdsDzFaKRH5E+3d/T5E3LRippKu47Qr7gaPWwWFbgSFzf0T
rPxqtCtYp7AqUjxYSWJQKs3h2t9f+rEO5dYm9ZY+u8c5AMfzm/DdSRGdGiCeuY/W
wS7HYcLlgmz1ov6m6awlIMnArQVPsoupdVmW9CC2MuPaZSDECdxe9yhJUzhqGeOF
HYHez6sc3PMHpIqQ9XAxetBws85Fco0ioyRh/jCk58FmvvU8bSdlfsga/ekVQyqt
PQVFxNK98jD2VLrP4Q6MiNo8BuCBb4BohYpgJ3sFW0OatMC7Tj+FlmUK6Cpp8a0w
GH+ZNJyQGRIB5JfKCJ/zs7es18ibxEc6jFzSmQRQPZwpnIJJjlJr+IF0l2hXeW6j
UxOHYKanuMxyBNZoboSI+J+Am2zAf+HzYNL/4t+5BZ2jtlPQeWCWY/WBVhezWMRJ
FLRcT7BKzOxwBisDX5qomPTGckb5Jodq+7Oxiwg51pprDOtrHRNN98aMtEH/SDrF
zG6xXMQ4pp67HTnbO3+zVS7OTxQG1aVEBM+nqSPjKh20pvr6zSrNncbNTzkAZItM
bvtPoXao4NvxUuPQ/9FDUvVtjUeNq/6nBA/TZEnNUf/gI4cDerI1t8WotQerI9N1
zelEcckhiB72bij99GK39qj35pALLZNtxpvRE76IWe6fZ2A4Pn2GMrs+1Uwc/SF4
J4z5E5lGuL9JSmXGObcRYCUoVxKjlVOwvCLMHG1TKoQI8o/id2kqyku/oSDXylfP
hXeBkbcqCsieCCc5qA65xslc5wMExdGr/il5CGP97cUFecL8fbOoZ9mX5vfq5FzS
zG31sUx3MnAdEJ9BpwUcTSplQNpZuHlDim2PtVhP9PI/O8A5CLIMiYiRLBINGtiN
QWcXm+FsAyfkL+y87dG9vfq0LEk5NWL03lZ6f+PIIorfkpoEuq1Ab0jmQVy8ouJ6
SrYdc2po3o/qj5GLOfbbOGxOEniBUCHZ0Cmp8rpOIl6Md/6SiAahppcW6fGVY6CA
cE1w4azJGVFRYVSyV25CvIPUFkNDfQYjsZhHCZGCeOIZRE8ZlYfZ6PdvJJE77kks
w8RJzcgPlKIlQlYA7UiHKCTjamhxld3BawTpSRnyy1JYQ79/erDoy73BgKin4JUc
WmcuYVwiED5dKUb8xxTpsHekB1SHTKMSyoikG4tPg7L8HP8b37xFXgBsgYWiQkbA
rDUEWoO1dI6YaLV4FRr17NOKBlf8TloS+bcL82jNgMFJzK1v++wnmMPWuqwwyUV+
O8lNyz3Nkf+Z0L/xICkRuSgZfuOouLERdCkyA2au+itVVHPFcJLaG7E+QbxCjclu
aDuT+rb5JW2x3G9NI2c9UW30mklWZjiGtnK8vbgzQQ7fj4UDZZT9zSF1H5R5Lfdg
cmhd9S4l2JY36723ATA9UW8OACp+cfg1OaWRRolqrG7FvrFHsJn6HaxE12P3irxV
a5nMUL2KsnCy+fI0GYylpEFuOGsvNcQR/aVTnp1Ir2hw0+28rbOTJQvgpjqwIR9c
o2vAST50uW+cIJYbJZ411RUXPVrVYhqp/rA9VaypBflr8XysKzpPRiFSe72M51ci
z6mHVa74Dz8TDbzU9JrkEq+lGk+q9BI6d7KDMdQGKcBHzILA29zufNOlH2mGnZWU
TGMXXyZvPAAPimIO4sizMCY8Q6mwktaPILZVsmP6ec3/6KTUjq7YvpVZFK1xxjrj
0hc+Db9XxY5UTXvsiqx1pIK3p/pLqvXwUon5PsKCkJCh66JRqxevZieDnw8FxQ6Q
Uyc+uKZ897ZaAEvwOfdUlu9tYpJTrkiisBp8AISpoNEf3meC/1Kx48zgfgnBVIUr
andY+Qphn3+p9ggqpOaHsyRk7DS1HPcq/53eBwcXhw0+kfg+7+wp4OK6jU7FnxYQ
zskUBE5K4heeF5YX9C4yDvgA2RZDHBa7ifN6IhLOQVKpk5UksGFlmJHsl2dI0nTk
TfbHN641eExMtPZfp9lteQ3Uq+67/KJPpeVC4tDpkeX0x9YfWjiMYMlbKDeexfhz
FIXwDt+Bvkz4XTWCa+qF9nIUV4PIuA0KLcoX4L1liKwdnt9Ahof9dJ93uItmoLDu
Yram7rRUMFor4iQs2KyMabeVGwvrW8G70rb5rJgakTmd7KZTCs3wg8P9VNyPGPXx
R1joYJcskVw/A8i+vhLn1UZ1nZJs7t3q1XCX1KkPgd6f+dNZR7/0fSNaCLTAq1Ri
aqdUxvZvEFI0duuTLUcCi5nArshHk31lJuZzjBgDlGSb/QBOSl3x+f9xBHHnrj8M
+cGdCbMgQUggXU1M0mkLgHheo8PgntmZcxMhUtfds1WVj/14oKBY/vsvENtrdV8P
HfJAOlNXKudVSEwvieDat2KmpgBMjHfYDGKcjzZff2RxmuDZOYo4boORaRvBwRB1
PQCmGdBdAXY/MiS7SKr3rM0H4lVodZKvhqx4QDG/BqDmsSWn5oXhUBy0rzc9JJor
n9J8V/ea1c+ZJD5XjEIZiEOpXXEAPZLT4oufTPESWMTvkFwpfpyRzxCjtPU8Ilbq
QOnCR2cYoldzra9+B2vOqySEd+vnx5uQAHHfrRvkPCXLZMtH99SBeJRCSQXSFyMO
fzsr3VWzowNLoHxKfHyNiUlML6VEIhY3qWJsp2xYOEmT5S1X09FJ3hkTxYRym8R5
CJ25yxPzh8FLFCSlgtYoFhDvjf09aEx5/yp+4qIjrVGkiz7ZWYIrNLPJt67frgNK
f5CSljabIEMc0bIbyUec98DWD7pc5qDfRRCUxPSYPWBghrSObifQVmuAf5YBLJzt
vZ5fa8nsAfdKFYb5BsZApb1OdCRj4rWwK4w/sqkx2+a+s9L6MrGQVg79ZYXMQafG
jMV/3Wc9woMlQl4Cm5/QsAAo2gAeQOgjNTLDc78mFhU1K7wJyycENX/nMdMiK+0a
Vvgmz9i9C4iy4B3s0MXsWwNUNeQ/GNJNt0ruT5rIfoQ0r4aU8FJKefyB955bZZxk
wK6tBzPSF0GoIV+t34vp8TlYa8vMsczfEl4deNqdmuQ9fqGoo5a9mvzSulTD9Pyw
Hhpsk3gjwJvdBGfODRZqhnnzFI69dHGIaopYjly3/t09mCmpcwyPDr/4vQ2hkIe3
mQkbSOt5mHA8SQVvCDrp+dEfg4sl+5XRINNI4/KJupoIX3mvpoJX/1+eyq8QwLN1
PnYI+eBynJmtEA9f1oVnvTSNXIrqAI94o0xEIR1aqsA10eIhOWHmsiM8vIL2zagp
e/bnqmWv2ApcWDwm6RacWSKJsRXsQeKEHIB7+vHcjbGKcx4wVzn1f3DElCEX69gp
Rr6TwQd9aFfFU6oEFatZdD9hSOZyUqXeIaixDhPAP6alyRJm7Oa3jVUha6/Wj84f
fwWCYQCo/L6Lonid5kHrjsQaiCQ5APLq7bUbqXfKx7isHd2ZtwN5TxbEE1DMkRwx
dWYmd6qCtKigwbwToOVBfgaZh++WUbUcTLK0knljeOBh+Xrh/18r6IA003Ev9R0b
K5q9wjxydpUmDYbIK5bDsOAddi0tR28Up4HZC9EmR9ZlhfqQXtQYNk54SZX/g0Zi
klTYoBThE4mJgRVa+HHIH2BjotJJ8Iap9CY7G4fheU4/nvz/gL5Mq8c34mn+yhoF
VT0bIf6hkZxfIDi0vwUPMJtdKoIsIcyhuhbBkXLQ3LuOP/9r8/IE+zkr6cElOl5n
XQYhweGGfNY2sGCS+P9M53kPJ43QRo+OybKPsDZlHajyaNfGSd7q5ZW8fM/OyKiu
9JiD4gHi9S8MBz/4atxefgypNzWlTyQO8X3gaG0hQeFzTYaKTZmpBg69oORCD3/V
Ytlad+ZvgrXW+Qh2e1Z07Vt5nGaobOIhCV+r3CuhH4/JUq7zTwKHKLtO+rsA2pfi
rA4IaTR2iR64XqTzUG/VMlkh7xqZreBKZztdLKNh0FybKq4Z3kupR80zwKdniJEE
VX5Le/wU936JtOiLgiwx4BlqjYDAuv5GIW+pDP00zzI5GpMhFAVc7H6wZ0zD+WxB
qyVyZ6TQbGTw20POQZ2UjHjyLy+P9Y/5fnXxLIbWT65gMSmVgGTNyMcNQ438on2z
d9ZSZ5+VqoB992fiPdNOqf6V2yiT/anRpZdT2mWUogLo5+M3hUHbuZPXnMuhGB0L
t0zQ7B1t8s64c12B1y/atDJyGcl9fXUjZfd194w0J8x8c444hHrl8kjt+tIT90pn
GUgQEngpzLwWsgx8CTwLek89MPnGjPWpIJJePKgWeVcN5U6zlJLNSsUNeXv4uOC1
0Ru65M1eMRqGFkHYtYufPaKZYNn+q+a2IyLAtO8D4LTyBGkpA8OoaThFiDi3AQ27
v5QYJcGflFdFZEZyTC4G8XBQUJj7Trzn2zAqUfFjb9sL2lCmxosmhKLZx+X8JbtP
RSg/OdDUepl4QysyWtxfd2MMHcsi+sKPPj4Kb+L2RhD/Ukami3GXsxhPPGECq5yC
DHCKXsvQtE+Ccl/dy4xvY1DX8ph8XiAtloIrqCHB082Cl8i+ltPAxpwalCc5+LGZ
I45+QpS9Vx5q/rvDY7vkGWwCs9FJu+vEjdDWkU/A7ZbiVGKOHITrvwZnTNgTQQ0B
YyRtapTDPTaTEHp+VGbMQh3BnDlQtBKjYeR2IfluXBNK6AU0/F4fr4zeKWd45R44
S1nGkI9kKEcnE2X+SFSXkKWqqR55Ap/CnT/x8p10D1G/rmxJkHtTQ1fjShZe4CdD
bguEV84g2+/olw/YA+ih8AFB5ilgnUwsQLgZMYYeH/dvYStBBOd204V8G2McTcYY
g6yc3U89LE4+n22odAshx4IBVIFP+P5wbM31OannM/tmM6bvuzl5859JqxC70iN+
DbmnV0+GaUktooQJNMZoQ5DCMfDK/PFc47MNlhJVHwvwppxkqcyJh1LZK0vrM99V
+KNAFTtQ6BwMRvuphBIjGGzirOTVYLlm3DxEa9IdvkSMDfIWBpUcoEHrQj2bt2dw
T1yCVUEFO0cXXfeQate9gXqqSiqZcptxN0i+TPyn+LcmAT85QkSENCg7mtaQnUrW
nn+KNW5nrhV/R6jAdGPYxPOoVaSeYJtssKy3KDO4UDe+q2fqYTQfR+GEWQQr1pjf
/K6tIuDxG7Aas5IndXAo/Ru4jzb/wNtH1hvJHj4dM/K/uJNemio3AF5++2X8dA7J
YPlsN8auWzs2evIAPKEpB+l2+SoJzBsoaS5asPsARJtw41FYPys6N28LZgWsfaXb
zJNNBvWIhF+e6c0Na5Xn2J+Tv3afCdYdbvjNN/Fi0+/R+mFjuUdoPagq52+hlZ7n
8GXalq1fBlOLlMOQUX6saVwYiE0DBiaqZNt47fITNu+bmSias3PDPGb1siDkq1Yv
4uJxR8rYwfAlsJRF4xhmqMSK33pKYhCCZrWfSCFluCPVORLFSWPJISO+9NYf8iYn
fbbF7rvwgQtebb9m41ccLb6TT4sZmxlo0g9E1L59k1z2vEamqyJosuW3F/doF/s2
yhDvuglnG3hYndSu2HN0/+Fe4nSNKyTg6aBWwCgh7Xxn53aofwIZvbVpBFOFHlbt
uuepredNf6G4YBRGP3Kowes5+fPbRebR0fnovCnyy0QG/YW/NSbHKgPEZTKDPEic
Zd0MPDiKPGLbVKSVzi3YhImBPnHoekKhGnWsGjKTJRPqZwG3UHo4V5iWxPfzO7qV
7vaiFaNPso7j3tEgYMYq8QGOC9KYskw1R/HAcVMT/ulwi0lnxdYtqOeDiHf8PgfS
cHgS5Tc/zcNVD892n2Iq6UOUseZ4YvYtLCkb0Rx1PPs1mnl0pKa2KOGmPKpN/19t
wFb1Z9a3T7uD2kUJixRZCXrr3IrVLsFKehYuqb1fFaB8C3vLvZglV6V39BCF4Jrc
EOl8AZgRydxJ0gLROpkueGuEUIkB+oDaVYQyejVK/NOCXPh6vq5S9uI9z95ufidq
JPQ78pnXnADVoLYDVzruA+Xt4HU9bZeNwYOOO7k4M+mUWL5fLV20yETLjMJ1WxBr
AOVuLlVGzzvHshF2NdjxzAPcutO+GcGdrNv2pdN8BEVW+bE9EI5ekedIIfZbAUBr
6UfmZ83J7yLlq19UCj3ucdLb/M3JjS99kDYRVlrXb1nYDEQARkB+oNYJQyufPUb+
oVZHLto3BG0CtbC38Cp++LUxt4473W613NPzrRJWAY/NgTbeh4NwCcfsetrouzU0
kqKOTDg1cQpC0FD99rlzoIk6zpGkZUeODlknrzZK7YejQ/G5eEWKy3yamHsfYYpO
vesAmzm5zZ7QNMW8tOU2JbmxH1jIHrCMaLgrivcQzfBt3+EwF9wSYsY4kYewjC4q
bNHRUfqkGYuD9aZ+mhgLsK2XxujXfa1+Y46mHPm/T7Tg9gjJSLo21CMkiNHD2rRh
aIOo/pEwBalkOy3t9sgzddxI+YzZF2gs1IrLNSgGok7bJsrDpMhfDto6NsqvN6u8
5WR7QKC4oI5yWiCOi8OOyMmUK61o+EvbaUwjFAPBs7vnuwcnPvqFYa0E+0hBoPAn
S9SKXVsM1ebR4ada1K2vsdSZwEDn3HBX2QbFo77ZT+MsSgvT0G7o7K+k6Ox0a9Bt
dWfCPZYJEKo5ddCiLAH5Vg9LxH3rZqjjAQcJYGyEIXx3H2vzJIssD3CzrDESOkZK
BI6Oo0S8QeePFUhfN2p97vOt5lInHcP1WNU6utzoxzuSnFrVTpaGvVPlKXdp46VK
/kHoYedsQhHyOfJCbuTzEYN1aoDo6w6+eZfT6poUE2uMgRBTykKul0GUSscXjv0J
dm68K9Y5VZuVZc4A8tJFJYDH46cNZncUvpNdDj/hrCphxo0CN8GLPK+1rhsdV6Q5
7FFcQ6V29dw0dEMbKQn2YDzqbEAeYt6NaBUe8w3YPTCa5ThIk8d1HifCpNSILJ/6
qrL0w3Ie0ijQKlNvZmyrIDLz09KTsRxy+wu45F16q2RIyZJVF0l0j+BAUtRTZxw6
4yTslnV/6olYISvVYY2ZLNflfs8zQjVEKlEun6EzU20iXw+NC4Q6CmhIB3NgbKC7
Uueh4S7OTo3iSF1c1g2+BudtIBu4wnS878r58U6/P5XjiNZNEpBieTnnjXC932f6
VKVrcfBk9KGswLGF0ZYb8Nms7mEhnfS5gOEp7LaWxIXDj3yF+kpf0Y253sg+3loq
yT3CggypocIMV9nyZw/oWB+DEsy5vuoHe1dGEIIDcIXT8gW+yoznvlEXJkn4JIz3
R91+YIBHme7g7+XycmhmuUBjvCP/BFSu9HhYs2ANXhybjZltDuTW1wYIwvdl84a7
B2tcfQhPAURhRLBTfNxJu/3WV0BGJo7HrJJvbY6SfvFP4b33ZgcQzI37I2+SG47+
SedO8g04W0Yf2BVhe7TOTUFFbLpDNDcsAvtnPX90ogKs6DjIB5KMaJpCOebK+xpb
/PeoCpaeNYFWxRUn+odf3jSwK5ueqdxcRa+VgTlkIA3nsGlHWLuW4vIERXbWbGC+
QpjWgMxhf6HZDcV1jG1lWpjceux5oiZK7/HVpNV9AidON7vQ4lb+zUxGb4vGWRf3
zZhXPZHaxqhw0ycKMDjbv58sxdwp4FYkmiR8Tx/H4IvOJt1iXa66HVo7ud4Pmr7e
cHd7mcBYFc9kVlpn0S28gFq4dkMK7yl87Y0Q2Ox4y6Cke+npZYlVSIUzo/uEQpi5
KPlgfxSSGyZ8cpKG8cuOzw2zm7vv/Y6bLAMNF7wCXzSHp3XsYWkaUNlD0KS9cQKH
9z9GP07eUjpxJix9ku/Dh2W2fwoqKk/4P3stgqYU2Wpxx3iREU5GvzOF41vFuA5T
4qDv05795JIwgBr8eMGMmS66KiN5RPp+PT+JthMB+HHekhzXXlNitwePFilWtTu+
5llWB+rQ2uIyUKRQGzlY/nvTVKnWkFnKPiJlaYZE7kbzHnhY0ScPNLiibqzFNip3
Mai3QyQ9yP2adbUzOWJYtUMLan749mRT2cQ7D7UtkrF+Ugrh2zRx0QvnGfU8HJO2
Fb7e0ny3XZnDB0tGgLV6QsrWAQToe/EBPiF1vwHVAs44FU67ABno/6PLRKDqJ37v
+UscWdYRv12+A9R+he3gdz/z0LoTgMDSLhlYPaDJ6JxtNrwJ6JbAZaLoBartHhNB
D7j0E161jyNQr68gW7uG/ineHrHjEUP8ws8tb5whtwJPLKGHzavkANd/i9OFOhVQ
gI/xKFgDrZKpVWQzV5zh0QYR7CP275iM2hoXUNGzPlx3GNrqNgjiinBAMRjKj1S1
XFVoqkC0BMmuwJ3C9Uc1RofOp6XKj5Mu/Z9T28wJ3xki9peietk9p/7SbOi5Jtux
/Qrb4gSWJ87BSGuWdF0jlM1kS923u03LfTDIjA/bRkmAoM/EcR1hUDyO/Bkuqp8Y
40SX5LJJRKEkXElhxb4kSM8dNuKnlJmxeWk+ZlJ9QXCI0XQX/I3xuZduO1vFUXhm
VxFGUDkreEiQB/qOiyoSrBFXa1N20gHTSt2UPc/VvK1MdpncEMz4nrYc1REXBStn
oH5yBTgCkSIlBFLGI2FPcwY6EW117eg2YW9qm/5p2Wo6UuZfKEjri0tSYJgQ7CNu
4I8H/66Dkkk51tEbtzFrO57pNLqEMD9sTZkOt1gavj/FOQ01Gi6IAEsMXi189fpu
sOaug12i1Yav0qptTmNO0t0Q2SMgIV9VnyfaZANM+7F7n2CBJAqbFxjuDBzxVgUT
X7dos78ujAjLzu0gSqRldrWaljeY+k+/cKtgYmzWQ6gQKMJf45dHt5ZH9tMoPf5o
oieu0lm11TNUI/TdIcHA0U7yGU9knuxIqbPR/6tiGcAA+dyo0mLsR13oFuNR1r1m
UN7lyRbrleuxcQRvQ2JbvnzCRK8z2HmrzMH3+3skKDvc5GF5sDJ+a/3CStnud0Yp
re9nBpizqOkf67dRsfUZ2DszU71zZBmMwKsGedf3nnxpi1CprcX8tSTadMHWovJP
4SurH7sxBJKjHHacedTmxxh+Nv9ZwQ/wK9HOCx1xpVYsSg9mmb+ZH2EGzKko1Hkt
7+u0jZ/ZYbqEm6EUDa/AxgcVCeGNQX8Ri/mPEgdSXx6VrWaavivw9ZKgSL8XqOnq
nDDJQ1+VbuFPeUyvawLJXeP4m/b5c9Q33stKR4eCG/W0bHlX3HyccPLtGSEioeks
vL4j1+ymhTqtB0Qn3squBKfBL7bfN1crBz5ttveK5Tcun49idBvtFd8Vj0hBr3kc
kYkUr6rFuO0rhBpR55/07415zO5AEMSvETveMx4wbC2gVJcApv/BTnGdOcANxQR+
mM4U3POWanCohr+bGi4eMkqUMuRx3FAAf7LeSsxbTHXeXLM1+Rj6RHmDMk00OVdE
GFgDi1/jGry+yZekk2vOlxL/nMb1ipSGXtLTfwMGJPW25qWeQwXgGUEJbfw2clgi
2fTQng+rg1fSJum6x1cpximS2VGH9h46pBvdKTWkBhjZy9nDA0RbODkrvVOg/dHU
bc/8NRd6VdNoClsLensa8gTubJaabXM1jGpmZYP5N0mpYVfbsiMv0Wo1EtYR43Q/
sk4IyxmncSTGx0HAyAucSuPHt2Od4sSWySh4724wXOWvv7q4oZSapZ6CjRDu/YER
94coh9I2ya+LfQ5s/ViY5JhS3axb2iOKWnh4wYl4SeD+YlBdU4ieHMKuQGmKsgrW
IifxHxEQzofY189oxT9As58l/lFpNVlAuRE83HMnuvjYGMhi9cT6EiBSYJ66cMDJ
yTAW1kLxJHsXge7X9hTnVvYqKlejTM+s/pWS/KhnKWx2WvRBPuy1xPVjj9QbHfAn
99KiTbtyVgxDqE+wamda20iXJseXcEFdpuQbl42EEKulyo/6vnF+FFUkz9QRZEFr
DUvxi2uVSR6CepMxtjjNML+nrEBjTYA54TNEJxO0iApX0KkStTUKz9A+8cjMZOJV
TUj1hn9l4KAiCFqDUHkCWT4jFW+387XwfFn4mSvRssS0r7BqRy2PNJh4u6MGrtLO
gkRn0pp6YTgyWnE4tFSmYy9aZF5sp9JL16oDcitSucoeqv7VMS5UHcGtMwV+aVR/
pszP3b8/tDFz8KQDWq4DRx9zJe8Xa7NitOoKGhhzYGtw5KeLjcTnoHKNzS1TVZFy
Jq31eDbbGn7NJd9DPidws5G0isPA1xHcxYDonQBO2ilBYz0p/4ilNUlwdpxlt2fh
/MYttOdC4ht59j8WRxZkFcw2GA7+rqi3UwagDEyETAZeQwd2SxwLpC6ViFbmuPYP
VH2DJqejjGHa4tEeA2uzi8bJS2ic7EZh8QzLVplybUG/R+NssYcfB2kE5xunMm03
PGUKkNxtlccJ4k1RGTx4h9rXhvC38OMBqnZYa+BSZ4ppcEA5jEnQsuwmkw9p9bJr
TEsxv6g8yHIrKvG0CB3QhnWIBQIWu578W5vbvCVGpPQTmipxwLuEEcH3CluJvVlb
aKBslv+cRJNVNLfjpJ8jXN2qLNIxruVhLCtTJ+Ak6hix4nu16fIBttM9gSF+2OpL
idyuCafkppC1yLqGrZlNLTaTF6DrPuGx7IEsXoEzAy8J4xO5NoFrqdjVTph6Qk4c
G+PKJ+Vpe2Jkv3Jc4rvlQUGF55ufmMc5zVYKvQhnrib5qvi95WBsCJuIvALFhIHX
egI/oBGhqRhm4SsIs9PjySc4NMGyz41amGV0IVv5BX8S0BZSbKMOU6szILphmprP
SMzPQLzvWmjG3FWZkrsZOwxaNW5KZDIu0fUJm4gmcKTOcWDdofSgzQw7dvaY66KK
ZpcVnoBzuDWhoUZY+JOtkwb3IfihcT5RhxeAXnZ/e1jxBlYOegjACbBvnhFEJlkE
Y3F+Mtd/ECH6IKMgIoi+igq9kjVK6KMguV0I5jT51PPrl9ODQQAIRLRrCPIGj2yT
o0UsbuuXV41jbbaR8pzyxyad70j5Z2+ZgoD4PMiMQBlAVLG8R36g80XqTcX0ynFN
B/CKusopiFNmGtFtIdgFGV6jghFjyTMKr8aZFyoGK3n+NuccxgEELyKD+RclrW50
M/SHbIkL/rb2fQG+6YRN3xwNxx0MEWB9mBenIHcwj09Lo121+9ltc+YX44mvQEpv
DHx9qm2HAizi4PcxYqfJNAU9p2BOMkscilv5c1K40aANqWAu/tB1ENUnAdTx+++I
HSPvr0FEMaTUJeEd4bSH9O3+32qOij71KpAWBH7tVUM4ol4S7bxg5O0VQz2kD3uf
V8kIJ7jKALPJgKxNNpeADniytOAh4wvcG6GjjAiPaMbUTpihOFQEc45MdAxqkTRh
+bXdLmfo0gh46uijgAt5LoGioFDH/nsDRhGviXb0q9Y5CAJBj87/nw1P0pqHR5/q
rcrIw3P1zmMYZOu9ZANHs6MHVhjYwZN+Z9oxNAG29cTqEPCjfUUBkCSZwmxdxsI5
pCll1pCGiWAxmszuMT8YU+STN/Df1wEGbtgyEDRPVh63kyju2+X6XGp6y/gyyj7q
aCduwPzAGL4ZlOAxrM1VP2LRFJB+cbHz6p+OwsshY8fC43biSTgmaWfhlz/GJprf
cs5Gji2Ai//xAQhPvt1+yXYHwFGTbUdgQiVcl9PKdVOs7WhuCxPssDpHb7JMWmqR
vO2CTE//IQKobwOynSbQxg7qE6Pfx9Q1/H95glOHxHFTMTYHqlLYWWpRksiOsJQd
YLQn3tzQVGJZisOWgbYBZ+wnohcwbC9GOVoM/iEzmOsUFlb4dG/Kw4bxYXfh1nDf
dhr7VOQj37YGmfdck7A3cGBJRBem03RPdXbM95OqDVZRmbevKDFzwVyJCOdxdcj7
/fGRdKQJwcx9SIFJDSco949HDCrZdInHzc8okStqnCKD53mj8q92agydN5+36lib
EHu9GocxzMJ6hXTcS05/uxJ+5HpEUTJDZ9k/QKeaj7wX5FZ/ms7Aec2i3PnQPfIB
nrfIxsGUV5oR4/rLnBqNHB+a9uFPfprJo+Sc8g90/m0aSoGA44DJXKnVGFp+5xfq
hOhojz8vHvTx5bnfk4s7tq2PPfEpx83DbfH3ekSe3XiEsBkG4nmYe4qh/Up8QKj/
GusaGulgcymAdrJvtAeI8kaGpL72fuxqzgK2yCoq3fmy8L8/2IszXFQZkVTCH1/G
sszUkXCsW4gQ0tES6vc3lNhWDea7NGw4ilSswDRC+5D01hp1TGPQ3V8DuOXsDEUB
iUig2NUZ8aaEhxjNEQR7MlsD6kax1x9rhn15Gf01jm7rTUjiUTR0rAX+TfnjT9a+
JIqprkQn00AJ8M1ZvlT3/6KyP8AHC5ZJHrx1JVew+BiEd79rYdc8EfT1qMxa3tor
+UAPCCc6tqHEwjHi5zE/31wY12seURUh10XXM48NL9HbG8rtAWklizO4WKASKZNO
nGHX5RnwBqg/wPRfrEz5vvfvUoLcPhN0mfvu4xO9y8wWIPgrjO09aMXaTBKlNfSs
n8+fLN3j+DaXYfG/QB746Qd9i2ZdTMI6Q6HlJ4T2Y0HyyC1PMtH7ToemptFc2Bjq
ePQN6M6vtQXNM4+iDZivSaJTrgdbxMY7qRR3SxoLse75HhdVcn4/Wm0cLleARElt
7BovriB++KzLgJbfRPiwi8WtMuqUKv88PXcbP9y8Jd0ZFSze26aaPGu1MIAsYJ5S
OJoDuwSrCLdRQBzQkPsgoZdP1s9Khq8mtE7dtjm6P9C6kWfiBQkVGQbXLzkU0LDS
6BSiENKhn6lL84Jj+tvSFgkN7dmt5vfgEnDN21/3/Bb2w7CVkh0r/kdAht7pBVMV
xSUybOtucdH5O4PaBxpFUTVLQoAJMTUl4Z2d1yLIiMyiY8y725eURnlKdEdqoZRU
5g2LiVRUv6G5GMW2phPB/YtJawqNZTYggRzrHuxEWQldhbLLnY+KqjF2RTeidHvu
iEEQYWq2SVw7pYFnWP/PCL4pMmC/U8bqtvZRexG/QJ+wwt0kD4ekH5ZBp5XWi+a4
OlHbQuSUeCL84U92CIXb0W87BvJvH9Y02GgMtbdKTRFvhm9NPam09CFj996KlN6c
Yk7Quovi+6lco2bzUj7zgitSiLp2HwR6YlLquca6/tJdhy1yP6I1jEEVy8ko4Spq
FVcdxgIhsy9P2wVJkKvR3d3BUN4GBwz7jnfxxDVriWeOnYESQMJxLEa9VIaqa4Ng
q3/eRy8m8o+/EG6nNX/ZlEwtM0S9Pz1jQceQfNZQkm3U1aIEa8f6v6YLAJJugSSo
Dr7yHnuhpL57C6W8fSMFKLhYZMlxT02OEqb96PQXBrGFMy/ImSqIgneOHPaYYndT
2u70MH1sybcirpAjsQle8utFfGzrU/UIBuG+wAt7dWhnfHWPWYf9GcPjPzUPEXrS
CQnTwbvCCrMBv6m9jqld3FAqsTfIGs1umK47n55O7XHsx5tkcAmCpcgEg++GlkcS
PNQsBAHzwSjb1MwUYvC2GzAsc3NIHryyYRoy85400WVD0aMNHa5K+Sas4YcUPKR7
4dsjUPUiP1O8FEe3rN9H9t9zOtPmYBXT1HsAtpkh7WLSh1GnzmQOO3vMyY8097op
U56UEu61TsIT5YJ2OxhP6HbTgBaTQxNq8CCsvsV5yDms/PaSkxfjC3UJbgkJA32l
YbMusyxqWVRBTv8fsnRUY0FhK94VNKAwmRCZqFEMXvPDaiauCJJ3kXJgqkqn/Cbd
C7xTol+2Lq9o/n7PiTPmfzO4jtExyIFxO/dFBQ3o7Q5bMjz1b0n4RuIdFfpNaewc
mfoCH4sdKBYznn91OcFIgmdVDenASDXCV+QP+nyEqVyjTiH+kaWhf+UvlAT+XjPX
LM/oAC1PrzB5WcpnFH9s3b4VeEE6uVijLVcU6YV4b64syb7KIAIL31zQIzb0uxjy
rTwSepfpvkj75K8WlwRVckDUpZ/3iebpKZoxcHJqARYP7QTVu+zvtREq3JkRIm0B
1fo/hW41IVMKyp1TCasymjAodTSBkrhBKxAD9j8mqfV+/e0GN1GeG2rfr8c/aEFe
aGLmlvZa8vSbTvWLZA2i9hlCQzh4N/+JHs0M2pZr/24DEqtktvxii4AH1i7Z5kf2
gWrg6FGpNH3t1jM5Rxh8hhrNw83Q8eHhFD/leQKkoT1dQrf/LKzshrpmwkbZJTVc
dA8xDyf9hXqli5TCYs0XpOYW/SvDEMXRoHs/Me1mrAqA94qNNHWpXOMq3XjGIHvB
NStyAi2UyTbpwobbTr6Oc8yb/bQFGwkgjl3XPbRgeqZuuqORbbsTkeyjRKz6JMAh
T0tp7jDPtTwU0iuBS1W+Eomcqz41dspmmsJCCkfefi6fw7w3EiU0bxElUDtaZiFH
Hqv6pdTijlcGaRqwMfCBLFyQFVkQabXKj3sEUmbqYRy6+lmXIL0O5kK5Wh8aBaCB
CQ2e8nkWjiZ4s2DYnifQB1Ei2eFMJHgjWf9LO1j64n5+2Ii5epO4FTFdccHnM0dN
Iueu8yg0VLiteCxx475S9GYZwQvxBJS/Mj+GkjEOCKjf3tKU9LVkXdPidqOTEKZw
jCCsESvvFLlWVP2QkN0DH74fmdaYlqLbA+bKq6X1C4f+Fta2r0fuugjzQ8ACfgQC
8ZTTtD2U+CiOK5gl/2F+48F3D+Hl4AmBOz/xHgVhcP4UYzGv7oH2HgS79+H3E9hx
XN2lW7rnjsYeMwc1iZ/O4o9ImuMpP1P3+hXWOh6sXT1IDdZn6QgNrkrT8PFdAHxT
upwnyqur6rHzzK70iBkRdSrwSavCfdvGtvaRFlcdts4X8fxqGOi8yntbz8gg/XUL
D7iCvmkf5OCl5QSnR5R4GbDMlBed4cOCfcdxRM7t6uvy+olD/WAw74+tFaF8WLpN
KhdTdxeYOJU6BYIr4pVqDpJGga3ejxWQu06i5a/fKOaBSbjkcFWM97FMcIX6I7ax
+LCzNssJZ3XHu5NOyLaHexfZg8G6Nr5p6AfpKGJVDP0+8CnSC0LdL4zb+lSXcw20
ZLMPuMJV+xO3QoYeV2uJni/ejJhvTHbSatOLNs6Plztb4UdetbIQBWsz9jCU/4rY
VcURkss8MNpbNgi9stYmie+I/gAvr2rx0+bsPLh5zM1LYXLLz2iChFy75YByPuBl
p6KPTkkJ9pMQsE4fitSBQ2j2eUQ6HcxcsYDpLwtR/CF7caO41VR1Ij7diMl5lcBe
jr9nBsQ/ztm/+owCUn9sNL7qOJjKx+VUzDhwa/tle5mcpYE2zZuuEWMFoQHf8F7W
diLSzpTBuIT8CVEPioYW7bc4qjJn94/jkNmFGz0w4rSfORM/CqZhjBhr1iAX+iJR
KXjkLKwCKLFui7o0SCX8sFp/7aF2gAtbvTE4QthTtIU4rdH7wiymcLJ7wZE+UIXw
C8Gg3a0uvW5Ve9nc8cbTmzsszaFiihoAaH/56x7eE4ocntY7+QwDWP4UbQyO2dDr
xrJFoHzGLx7TUbGeAzQJD6/BydTcpYL79mxx4ZRbNY+cUfEVhB/wtynhBaxhj6x5
owrcA5s73yEQucmMvGPTzysY5E39mURXd/42u5MUNeEAZcikvYbyqn0VH7Sj7hLg
e+5Fs0UvGnzIyl7YLhlIiVTTtyElR3JGYJoXHw/NIhWtcBQ/gqVC/cFFDNH/uD5b
FgvExmD5IlixIhnRQVaWIzZNwbiiKVsDLhMA701k4mj6CRUpP+Z3yid4WM/IJ7NM
II7fhpNflNsfIrfwmLuPminwnbj8VAKf6rGlSm1J6lgGAnpdUuesnXYAj6U/OQ4g
D+U9YDm4mKWy5fYiuamuNv7O0XGxKYS5vTJXGbU9dMn8UX4Q6S4wzvqxyQtmZskv
LiJ8Qec1mQyd5zh4dF1MbAkPfQ88bGY4XW3xgW/Lfz8IeZMBA5ecRVB5IHaGQUdg
1MaLKdYLiVzFrcARrwwuc9J+e4rJojsbGffPAxQY6moIYGgsdpmFNxZLpnOj+oM1
DgN8qkAxuclgVvxNzg75YgzcNhzK4SmIRSrAZ7oTzaLuNyTfRmaoGsEaLDYGxk6e
iUNhJFJeXmTLWiQFi00cboH/5gKqyEBrU7XUtNIU4uBoQvlnvOrVyqDxGdlv4eac
3qGqBtMHoja6xC9rlbxgCcWWqNs0w8qGmfcL+7sGtPVReUQiuguoMgp68oUiXcuj
RN3TP0Tvl116J3ORkrw4LD/AminxaRyFH/WQ9rwpFIqRTP/XRG3ixnGcvXBjLBe/
+DbY/7yXHAsDzuzS/c4rqthjkVahoUlzRCEjn7sMki9dcTGzmy3TLuQy/bMPGIrj
tGHE6ZyiWihtY8bAddQMD55/kskXH0INCqnId7Lo8KfSBzT3YArlz/iHI4hLcRcZ
BWmhXjDKuCmdwGSQ2zC8VbY0UKKUzcVOMAbyIu0zCeg6CcMcelUftacel0yFBUKy
GK/OxWi90HwVexM8YWktsOgVeGng7ablbMNqpUlUSKVfsmX/MRm81mMpXvDXLXht
1XpUgtIQWMz93Jec3dX1wsWWhNjxekO60SKYJys6XuTvLFKpwWxFg30IVJC2l+FD
sZGoIvsyfSPKQSkkZGmNyZh2WezAslYKO2h7b8qnZfFQYIgMbPvIBfBgHeLkXcZY
IisVfXXq1UxPk8RXi2SMGPnbIR74VmGXh+4INZ8swQ6N7MIfb0rXFGeRTyBm7g8j
Ge99IUwGZuGVDH2GqINWrMF916FRimIVqXk05jbCG8bS0e7blBwqYDi63B8KcD65
gT3GQd8IW/LfcMtYWpZHmtoo52b40V9RxotsB9gjPBG/i8CRNU3HJ7fRMwG0gfN0
AegiBu2nRWXL4rn105+xxxyX8K63fsxiYpg1zGqqWIhR2b+p/ie8/kHM/x1OxkB9
85e3+RkTf2DOYzlVSdbwEI5QBpSk97JNdK/kkdXlKWpyWaVZVIG2yf/ciiNQhC7n
bCg9k5Yk2iaow6zd5jsb/q0NIUeZqvmxu/u/ZnCQabkmwHQGB8dSi8paAKSXM+lA
GYZpkmHTBOmxj+y4v98uFvOBVq1EPPOpx4F831e0dsM+hYtjWSeRqXVuITutRbO2
Ut+Eh2RbInaE5IUU4SR5TIEf88MjL5sIa6GonG73hNCNUksYb7ary1snMhWJQuYJ
hqp+9qDV5osrBPpJZQI/mbIksTlalLPJcuzlQrrUEJ0l8L30ezKsGLxx0ge68AxN
zXoonVaWfv3Z6cDRjUpadhgMVKBO+rIeQX69fWK+Ee9w8LEeLt8ch7aNpRydgZLe
W/8mMLuAE/TGl5MIKbZHr7FG8XyXZJl4ITMjmKHwaGhu3Ef3JHRO9wPDFWg1hRrh
XoArF+P8KbNBxoP1aO7qqQ40SyofxZZGXpuG4e770Y9h8QwXdCKpfJxtXBRJtcZK
KiVkdP+UeiB//MGg42Nf9c+OhWGB/w0H5LMvc2wRS869g7WfNh+QW88mcC8Dwawo
JrrBh6kirQxu2Rzv4TZB7uKWfNtxQY4J/jH9YUXHQVtP1Y2AZVbKOkCW/3gRpHR2
nVo1UeFXLnHGn0e6NXxmoNc31fD/qmnYtp5r3L82Yrq/oNx6aMBSc2XCjB4pWqbT
LDwH/BDKbfnDE/BTz3oIpqACc7Erl2NrELb1YLMOqSqJMagt+Sr0l/ETOY1a7trc
iaCHv4T/CoNXv5vKbKsYJIsZPnIHZEXJi2IrvTLJHNMvF+DSfeivESLSCRc3Jgec
u/mfsVXRLeLpr2hQYNDSJjVn3e1VQQs401LAaBoI3LenXFfYbcze8bkZ/mxGkkSV
ZicE0qwk7iOPOpSyp7HkL1sTL7bJD4oir6EVGyHEXYRHHhEBJA7KAbYZeR3mNxR5
2vrnW5D5iCVxbGMT0RfoHe8Nfq197e3zS3mhMDXPx7vRJRBvfQW/oQ5JKOy1AN4x
9JyGA66jojf8qKksPmP7XpuPc1oQLDeJqoigCetoAqt5sMY4O2AkFhy1p6wJ9/F9
bx6iUhDxCTkwR76lUTetSH0WG9dBiA8xwVZaFrKi8jWsW2v4ssVHCgUXRZXpCcAX
29AODcgzPwqat9wija2LGry1Q0YNhIKO0VTQH0HrC9/bnkYaYA0tjECA77dvyTy4
Zz1FxELt0g1gKQYUjOj9o8qAkqNMVaevpgJcSctSrJyabrKNLh7LHh0gUIyTRNk4
v09pQzkwvq6mg0qa6aEEYJKCJerEgTO+DrJqzDpNfD2hYDqqYdWExZlgYbTodNBa
dXQSgW/50yArvOcyCSM6Uy6w+j9QaFRQ344qgSepBxSzqNMTWfy7M/9JO0JyMOXs
+Cuawxhbcbg7h7whjEEXCEBappH94jKaA55bLJ4w+MMtpnlFZPwpr4qjppL1lrVl
v8MG5qrfjXdYiGlBg3HhOHGMiKLBfBRkw8fhzNh9O5F02iLJaCJ+05FhYTDiAjUR
5YCto0Epf4EIS3SquSGaNYHOD2Qd5bPyhKE9Mr1i9OvZaTGuL9jx5EVlj8h49YKD
EYGZEnTGacB3yw1j5C1+SX7ua2WaoMJZa0p/bg+hlFqu4RvGrpSpS5yXvU9SQSKv
RzHAoxXzM7ZfKGBV9mhWJOiIE2jzJySGWQIt6pE/N2UwQN7qiq8n1wC1AoJu23kf
hfpIh51+j5PjqLOha2YJ5sCLE46AhWbegN3afTUtcu0wJ6mzLkQpEXAkqBQN9kwQ
bOEwB5LXBfMtnhGwOIdYHXvykz/SGK0UDliaw2pxEscwBdA4LquU3DXIESbEG/ek
XPV7+7ApzcWnZNFBdAfPGClsor8ciAOTt32djAW21dF7oVwo9W+bdJf1oAG8Q5j1
ruMZmotXo8YzCQ3RxEO7C1ZmbBqU32x5N/758utx+AHHxSUL3HBgGd+CjpwR5yxK
1qAg/3VFcx/npIhvq+bjshLB92p1XHqP0+sGy88BmTH3tWsCY4ff9YtGN3eNv7zf
/9wvBDxAAyICpzAs0Vh3P/B0ttN1drhllNR/FVGCfN9oaNfxbZsZtPeAm3baKcPH
jpxEdOTZJXXVZoXag+H2fGHlrBSNVUexlf3MqMv3x77cqd8h2+utB4R1Rxp3eW6O
fX9qrnmq3SC9XuqiqAEdNAHgDdTjkHyK8marSTLQ1RqTPFyNkPtNROw6kAfOxivS
dHXGtl8TylrdVF+CvSVCElGfVb/BtK6YwiXJKGteej41wDVt46f5Jbr2ZYBCJZ5M
6uP4v8rKrFDzn5Q2Vc9av42n0w9e+qlvrGW4kYvbnTLrMOYHYcCMxUzdoDSYV1cp
Hsv7aCAYd9Sw/GDNPdXVO9OFm3Yh3EcjM41hshsVrBtotAsBZHWQPVCn49wfCzgB
bC86+TChiG9P/BI2QJiAbyo91SmARoQrBdq7lJhrNzcttkOQg+wzTYzmCYlCTgCs
4Xft/KpYmsVORfxMsfvv0AcRL0CWe3HvfGddxUKPVmUmvp6nTSb+RzuPMX4fKx3J
PGHWY9ODw+i8FKNiukbVjFMDGvegIRk3NsF9KiC59DDJpatgqRSMkDREbOaZpaL3
khD01r3r9CZF6iTMYUGLR8e7RB8JjXoZmiJd2L0OEwBpOBojrC+jul+DtLOQ+6xu
DEj+F8iADKhrZSSQerNU4yLLww9XN5Rvbcm+T636kcWhQ7/XZMxbJvNWecXXWVlj
Q1cR+gPQ73TcdcZeM0l53OWNsPUoLGt0aSHSrPE0SRN/IJEuaPmtLjC0M+wpdjPd
F78+QXIB6SuLducYBMcgNYgjHVO8AJKb/I/uY/DJBH2YI3qbj0l+p1evtkOWd9eE
ItN2Tbp22J3lfZnX6w0/Ao2JWDvGhMxisWgK2szC+te9nQoxi6ggLENWuoiSVgn/
VzP9/a92xpR3yWBJBW6rE8ZiiaCT4WkIuWPnHae2IHWdwV46ET00Uv1rAnxzIDmN
olE9Sd3E4t7XHKM7a7onQh+B+xK4/LBrFMZiM+PUK8gITK97lJxpA2uECOAZ9X1L
5eMUP7YIYwO6xz/B0QaesqJDCEk/i6Hnr+w8jk+cdVbYgusAFJ1TbwdBhexZiF35
5WODj75Mh60q9cUrvLWCb1NKdLt5ZcbFr9BiItGX0xGnKenJIUzsbetr87WXk+bq
ZD84bIYLzLXc0BrrrpHj3pOp8fsHEmw2P3I1hrApWsncj6l9lyWN6lcO0nDNoafI
MgqiH1pNeWrMeb+cGWina7bwLq91nPUxNZnuvLU4OsJOu53XN5z5YqmKwa4yU/Lo
QmeOlsZi3HYAWmBMmngZDpyBtSK8QcPuRUgo31TBqDtg/UTz9t54QisY+DxrR0Yp
EUA77g5nJNv7sDlXIag1fjPSGRMUhEbXj+ntwHeHtp8/dRn2jWWIZsqtx3NbRVLN
6pp6VaKZe0TgJtEXhG0kQyiSGKqmkfi3cVcG807xwpkainD/NPGogH8tE7RA7AKS
tItgu8InH/kuNgjM7G4kRCR1/YPOZnFO4Aqf+lPa/vVCwaRzBSJYfL1XbosDfBSC
3Cw6a6ZWqWLvRtCZFrloNAmvYV56ygLnB3rUpDdlMKy/JfH9tmoKLQKW6QbkZyjm
CemF+0eGmgEfl1vPhBhvnT+Oq6GxpmattBRWwwVTo1HtyM8BRGGTSmdu7IC8jjMZ
xfJ2O/fBvK4+y7ztdn6F6QM3hEfQmB9TkTC4N1/HtQCIm8A+QKbR+qlyGfCKKIS3
gByER74hs/R+xPRa1M9ZWffmdq4zVEl6ByuUFhtrZJ8XG4yhZZpcVRQugTfN6OB2
xcvYdVNG/kJ4Le0qK6xBicn5G9xRC0bzRKJmTqu4503dvBgcQj5TLYaght9YaeTz
n3MXrzh6UN4ar43IoekSuR+KAq6FXIj51g8PaBjpvyEzOYT1jQquu3tp3VbcMZ4S
uqwmSHZzfzCQYOEWycdThu7t7n3H57NXBmNgTJPxK5Knlore0oPP8NsUcV3/uLD0
RJYlxsDPmNnndgOoSyjfnPpLaaoWMkPX0fOag9ryoyZhtSIE8Zn40dpb/7jguOmv
ELkxJGOYMLhlwLqiaVpBeFy5EkO+ddvnH4Z/XPmcX6r+CUxNBgDhwt4/wf60AwPr
gaEj9O1PiTG6jYCuSHv1GDL4Eu6ysVr1RGdL668LvSxyAg7E7vQdljszpFg35Z7S
H98m+PIyN3w3cBwgmwX+/+z73KayhPIMYkGhMLHmODFuEysvSJOoUD6Fx9F1Q2Yn
RG3HTmwNfIIzlMG7aFReln0BLbM82ImcBvNUHVLmoK54BBVznDB2tjvzAqbwh9QN
tjC1DsAZRouJ4HjwyNbjk5XjRRMzTAIS4UYwNzu3McW9WyNJ4xFB5QFhWstc5Xay
DS8aVgMg/BYbz3zVYmszpb8goJfLrFl0reiekbVxnLkxV1/X05Vdg82cCwbNMH/O
CoBdrmff+rsqVH9EZyS+bSURTG7ZcPwMfemmezlEz/UGCzXfz4ifdFC3uwlczB7Y
WD8IgheXqujcn3oiF8bt71MluO4YI8zwEth96ry+k8eyEQ4Nd0U4MFkuwF9xOdra
MI+rJ06CxLkeZhEHtdQNP+mVQHUvKSkoxuGheCtYYddLvW6X/XAUOHgyya2m+Vpv
9AQ6UGAD3a7O8AvAmyVHRFiCmya7pbxzT8WMwr1SZgBanuuU2wMFrwyg6qZHjq0x
vHHmoqfk1xXG9mcoX7P6V4HmFL5vsdfahOW5XKo5CuSAi1mFjhwE2gBZCtA+Q0kk
RE5BsGfMImCzih9XtXpZOcyuPNITg7qcYkdH91XF87tkHqgMRA+GfbVb0Rs1aE+b
Vq9qOHAjUgHc7PPTzIbGMtXGcGRfmBHo+rjnohejlGQhS/Z8GmhIwN5ObhH5Q1ub
O6tLCQh/j7EIrkdDxzAI2qmWkM3DxKYNYUxN5JTKorDsDiEtQdl52kRNezAgTD+U
Dw/Qtj1GXvsAZuTMbOEoS71QfpJ4SEpHb0mDK9XEvYVp/8qU0j1TvNHmYKDHTEjo
/oupB5yWIGscLr7XtVrFAVGRxtTCYFtdaRPm69tK0kBda9Vt2pvJeaEoLkO0SYnr
GL4gJlayj8z8ZLltNSN6RIVoEfkNGfCrAoQEl/CyuRJw/Sh10vsRe6NpEY4/LIcD
Jr1o23Y84ORGquIMKAnXCTFAGeBKt2YAghdTJ5J5rGgE0AmihF0zrLqZp2pySGmo
FD3k2ElpZrQUHmYpuUmoMTKFN4bmyL7rvT+ZQSeobt77/mX9Bp7b2bVlwdi7Lo0w
crB/U4oBkShQx+oQ86fFVTn/ZgTXuTcvIoQ0Psvp1TuL6yVKYcUBOB4aFG48Pybs
CGfYpG0rHo3TI4AjIAbIkgzeaRCw5ws39PMFEIK7RrWb6ZWhDuDC2jeeyFQddoDA
+dEzIGJm8NkO+93CJTLzDnKv4Dr+72reZRLpnOCKcacO7GyFiMn5CLzPxTzLs1z6
TIRsaQ0GVw+IXI9TeAhIitevAFbzH6/W8YAcFRu7ioIY4Y4dt26JoFg9bba7geJC
Fe1yT8rzd7af0AYsLyihL206Ynz2Hf/IbIm7VPP03t7qWfkWYVqBZte95RtdZ+V3
FT44wt9C2OX5E7LcSjL2WVoGDyZVudSj+4qUC3SZfeX56axgodLWN1yQ1cC+iAw0
/Q82DQz7Rez5xGFhTp8VWa+LWobg0EGUlDrPLnSJC33BpwX9dlHzKQo2Dw613x5v
zpOKAaAMjCsWdT2hXjw+ZDUvrd1AXNxqFdddwJVd7M1gCdvfvhtL7kbt7im8kEgz
KxGqTxzISLRMG9w2YktCxT5PPnBLh/OObeIovQVpKYqxMb3eQ0EBFakFj6xkMxsO
4Yr0xHPsO2ZW67he0/CmX+KSefeSG41uKVpRcicqXdUmy5t+hI+kvOwnSiKDoARZ
Cm060XGQuiRM7OC7qGODD15mBoWt26o6c2ReUGE/QeXQdMrIG5tjRbo3u0Zr7gzY
/DBu0RNlZJAte83v5YrfhLzIXiEbFK98OizoONcbJz3ZP6NkNWHsPWpJ2BeunKAl
AYD9WaAFCb4Pmul2PRvhTm1tqIeKxOzZ7PXuH1xYBKwajUvn7p5dr0gylMWErPUP
Tip9rgf5Q+NTCKjKt/17DlY9UQeGbQkzzeQdplPvx7ch7IbQMjObs0e6fy+CZZ1T
OMv8AOpueMTccdh1Av1GBJ+cyfEiHwYySOckY23glKt/EuYC3I55AReZUnbBBcnN
dWISrmNugBVJJIqVzwPZnjtmNk/zCXPyF1GqSB6V2Os9lhVXjr7HnXIq8Y8P/M7P
OcGaQC2OZYxXmqdXPf8wtP2Hg1tGrEZFIslF8IDSGM90RJx23ubhzLo9LH7nqKjc
yRGJ0F3bVdd+wO6kJ5ILvYkKLXskF7f7EtkMdZwrj0n+ehWAuE4w02AaLJj3InCj
hydm4GRIK4A3YMhoByrD1CEqrWoYpc3SvzDN+EoO7f5OeDZsg8vkNkbkxPldbRYI
bVT2DTmLmGzqhaX8VLZTMyeXeN8ajqzD6pFCaOxJiDC4OgtcihaY6oADC7emCN4w
D+s377NI5CAyZ7HGIDMNO1OX1t487rdg8QvLcqKU2UR4yxa1Ro9V3C6Fvf0Eq6+d
NF3r42IPWouBseLEZ36almcNBawjGx5qWHux59fjJQ+TNS/Ra3k1PrraS7y+BqI6
LKAZrSofqkpDSnypKDBaCJO+rk1cbng+Zf/xz5HgLgqzfJTMtu07hFXmSyZekSuh
Sa5BCPpZ7G2mdW1/rQ5IuUt9oiFIOvCBxNFQXelcmwFsp7yRrzkAQw3lNp8pzCFe
oZJLuzhAWOlijva1Sqk6RL4XGXAVYKlmitxphGsiSO3T5vh9Z0DQavrL31UgnWsV
Lw7yB0L3AGup38V2pklH9zkqDwqCNHPE72TjM5tbwz0kJfYwQB2LCVpPVyu8VrXM
j5QSLZPQwCkN2/gsk4nuOnzvQFQT7RDAcKdpAa9o43thrlSxKbPtJ41TJNGoCnKZ
ajuzJK/y2r/e+YQYTg/4gBjOw0KjEAocdbp630bZz1LIxfP+1N+HzVVrhpbw3P5Y
YRUl0ohaljU8pft3oC8D4Wxt0esAJ+ZLjt/aR1OLbgBn2Kw+9FC+iBHzyViM76HR
/6SzbFGkwhEWukhDcZg/h3VFFYE2KF6FNyaBupe5FyI43DqqJrnkxoGyJSD0NU/B
fT19apbOI+Q4VmVoZf5xuv1goHzMja9gMnW5pfClAamFxaYoInyUVjg5W6sTTFPw
bLCyuTi0lcgPfp3TpTfuITLw9dtP0oaSyA0MjIvsKS9F/pqL+HlNhBjSEyqAvLe6
SBB6a7pqRttnth0hthXqKvvPOVMANI3WHkpJ1K2E0WyOxe4bMDjYdRp3IooFvBl3
UJvqDAGdhZnBZvb6uk/mSSteko83V+h7KsjaeBRNQj/u8r9IppEJtvwWKvI/OCsw
UZjeYR3ap4iAgeNT/vQ7PxHCXaNntgLkBtQ4Ce2e2qrGF2p9s9yNtwsYru4fgymr
YRlwCgqGv6/aikmqPmEXCWH5R7QFD7X6SL7/AyBvD9aHi1J3bEGya87bOceqQPS4
VwGqtmWvy8ojhL9HhSqitkBMbd3xGzuFajL2R/CsMJxBX3WVjQlYtMsDlNWE+qRH
g3ebgbcrJW+pn3LeZkuCJqAlNEcusHyLYZngXlVhHlv4G4cOa1h1dabOiiuLeUfk
wja2hcQZ4voTN7Nz+oH/Er+JLfhTgqAZ7mRVKFywyYluOfS3FLcbRVuNkYD4EdzX
b/fwMm1wN5xuIj4hEmtKyXsimGQZuIFn3gLT/kLZM9LlAJqK9M028/KS+X3JhiHb
ip53HtnBX9vx14dH+riw6JRBC+NjdNKKCA6sE6ihA0ai2FmuRh1LzdLmHtjXXb25
zUICUNheUvwBIL+ULIR8fvGT8RjFLpnthjKlhLpYJcPiggVosKSiBxcHYE5YSY5z
DRYzLwTbEZZhIvSZyBFszBXAD8VHN7j5zFj4rEqea9qTTsXi4eq2vd9MUL7hhIyw
znyoiHbxh/fPxuCBE+2GQGKw6p5aNEyfBuI8d2HaJVxYEwhq5lsTbSIWe0MzA9hv
jxcU1yJjqoAu0kMaG9jj2w3K+h6bgqxfPvcEcrShi1o4M7g6gxWbpcFbLmc8MSis
GLVzjZPiPJgt36d920J9B2t/jupwA9P4mxs0SEyUypY2AY6btZmRFxe84MBs2EkI
ky8TcKftl8ao+Ch/nF/+j4Fz5KJjXGEARmZtQ4Kx/GY8+BTAwTSO90DKJOSuIW8H
/Q+u/VhLRhGJeRdMD8W8ApM8vj4CjaSqQduqJkKWfwWTcvn8uaTLNYWBj+AO5gQB
xiX2GQHeyH4qadL0dnMgJqc0cUj/79tOE6C1dcO0SlaIuvpfSxdbdWvvLDsRfTkD
Agx0DRbuc30+WZ97wKcqsOxCfjaGIGiUjkOHz5cBiwGBn6H9QyH50x6ne4J8LWna
NJNfOOHYk3waCS/TlYSmjipSbq36k24GS73xVgfkusVhwqgKtSedJEtZrvse+yyO
Ij969uozNvhejEy7LGhH+NvhfzM+gRiItGT05XPYYsMcZIpNZ1tR3hC5jiJ1T+I8
0kZPaRuGwkfGikPwxHi4cTu9QcE+ZV8/UmJqYVrTPOoTvsrQA68wWDxuS+Ps4QQq
xFcOkno90VoCmMxavkZAflzS0eyPFJ7ZYgEjax3HusW54zB7RRfiUMdOhN5/Kx5i
HpJrYJYMyftTjp//czM8Hb36KcVz9NwCii0JYES3j2nj5yexIFRSKmQUfaGmR8Qg
oKb84Fj8rjyoUCtq1Z0dzR4brk7t3OcLGcI4Wm47NIMYNYAm4YOvCL9y0B7Kzi7S
BJ9pPreRdo8gyP4IgK3QM/6wdb+NtpLhLjYNkngA1GLJxmwxwgAIcbprILxYrdae
sUsLavAI3gCKKBFXQwzT3IfNQgxlVvd9tX8732P3FHSXOG3IM1gYXy4fJwGtuuC1
jHen7B2jHdIJw+h+y8gy3WR2iRzZTbwBsXOBOD/YcbuOX7vZDV0A9Zs6VDw93f1a
DbGgzm59DdXI3vV6S6U8dU976YTqiMPfH+0f0dSLUnxXUuCC904SNi+pdTbE1bg8
/lpFmyRNVgKfFDu2B+0zFQQd6T6QMIU31d2rRkMwumEGVPI9WC3o0uBS4oTErUgV
vDU5S7qYUuAa6GVUKU+s1SC7yNoPg4dZ8lej3+FrBsJuHgY3jXmBHI5q24cyT1Ra
6o21So+Vo23dpjcmFD2cf7XBAKL2iKKUz06NeSCLZ9sGNyDmE2m/xOxc9wGpjdnL
G0MM3rxpVW2ooDG099g2nrzZ2EiX/TxusxWOxnw9lo7ZeduZYT4ONCM4AqvRtPa2
Je1pEwNs7Pr0jgELCV+nPXEAbFY7fiosv/zOO+GJvJwxFPeRK72lAAT4HpDfh5S0
3E/tVSbVlNJ5X7NAUFjOLym7udf72LrT75lOEVEzi8sjcF/e5J7Lf61psRo4XRax
aSPdS8TpEGdwzcPnBDC22fRzckuMsKCwCx1hLH/r0w2rqZ+OAqZSyW82bYevj6vd
+MVjfJ/TZGFUGwF8fxHRI6KdFv4CqMEYCIfdd1PIy4OWmrWHVJnhBUFfoAL/jXzt
CzfDqPVDZj1OlMuCahugrlFL66rV5Wc4i3Uk6UvR9gePPt2BTXtDXo15uLlRQfGE
Qc8+dyoP+wlLyyfrHD4LOwejPfjWM2KmlZEN3x3vX12GYb87ZkJ45nwlQstC5BLG
VAqI0KDf6HA3E/MCWcAotXOQxXTMV38B5fAWzIua/D6JVhjqzknitJ7S+q3IJuUb
Jf+qGPeoa3MLKDZWdQ8ef0ZFMRotuNdmnV1CLfDzWVgcg4P5R4Vq7P2SL/ewU5II
DbbEZFdNx6BWY9ra6iAo0YL999pgWkh8KXPC8PllzvecD+TFPT0PbbGVtIxF7Fm1
Zhodp5SjuBIpbYJCJpmIVbn0YOHxwZO87Lwf4KfNX2MgBuUi2ULvWv3A350vIdSD
1u98E6+FiCC8lRODOHjZRQT/tOXxWThMZJUR+d6f139Z+jPLoTjI+AkslsOz2Oip
MaArEuYjnkuRoVo4zAfWw2rTg8rZiT+xXUfYHv+FpUDMvWDyibBVU+XL54RuLMP3
bdxT/oaO4Eh/BL2ywbjlA2qfU1Kgz9qU0JtoywNJP7aYJ6zuCrq51wL9d2BmczyT
jg8rckdlzHt80deOQqp3gI5F6z9kmufFXrBMCRfkJnzEe/sXzza9Yz8+Krs4YZjp
cuF/yMdGBBcDunRteDDPFWgzWNw84FB3Xun31JIjeRdcJ/ocp7Iu/lUxGHX2BQnN
G2KLFHk5b/Dg6yiGGAHZn3toPMp88RXiXXmJcmFSBleMBuPQ7z14uqgqXMcVBx8I
lyHwT0gLKz6ALPtiUFtoIm01PamJxYMSvdKopOkDsmcxEtdExYyb/9cpM7QieGO+
yxRZRW0vN9YkhiGJ5Vy/yEWYz8mlfK18s5JtYFmjWaLhcs1pp50Hq9N/3T1DEZZH
mCY3N3hzsJyR6Mdo9LZ0+w1qSQq4w68Mz39akbFCHTxs4+zZTTWGzfRmh3umf3WP
i3H5p6qAWXJ0Dshzol3rkchidlhkhQXKipijSXQlZzjBrHzXqPYI2Tgi9NL2+rsN
Qh4ukl59uwlvNl3BwxMWEXZmGlf+S5iK5cx6ftkxW02k2mALNUflRaJG/mkMdvmU
GLx1dyni4IdMSgU3wkF684UAcqZUAcqDz4HLhyVB4sleSddrLwxCvEKTpQdN1vZF
7ek9PLkZX0u0eUjgWCKPBARPAlTRcUsdknMZW9GOI7MKqTXQFcqWkC7ZlRWF1Du/
EYz5bXTt0PKIWyLu7lEO8vrhCLd3of8S3eVwMbKQQSEgteYPh4eZngNgKUNlEKSY
bv0oZQnhnWeIMYEyyaF4smHcrxQ3K/C/xZM6aPbHtm9DyBXXAK1E2GcqPzbGk/mY
aN3ebADffwv6D3mrgHuOc2AL1ygBM+vDvzF6KbS9s2VkM3XR/v8aMUXZuYz0mC4c
ENFt1UiQomX15BvFfKC93yeqAISQOjDLyBlqSUpAKMlc+tPBKh+Cv2dEYept6256
qU62DTDF3nAMhdf114NDHO8ndXYx7PCNFUoew0s0Gb07F2er06ENOcOPg3IMPoSM
Wkmvhc0oxk9U7GdX6D5c5OwBj5J13JpjZUxaMVb0YrS6pBEKzCNN+sPEnZ6piS6n
Yd5VdRI6qHFTbZJLxbPqmLpM5Wn0SOMQCw6n8+/lJEuejJaeg83QaCC8oUzM7zIq
pTFLsX6iN2mB40m/JxbqwNBPQh66N6ZK/FAdJyn+pqY3rcc6N9mFKqHHPuaL1YZC
i0a1fxgGol7nE0VsYrzfjK5ObJLKR+I31A/RF4JsES+LJv+yZAAv+uzEUeBBJOrh
rfmzcdzxlsGqv+OUHwzrDZx30UQATLfEBvUcYYMaQDeyXqWSetJ3dzZHhEtkyChL
eMbLgcPvSWPNNA3M8f3jZY3QrmJCUW4zNdwZG+JlwbkHYnMK/MI/fWJq7Ry9eN04
5VNEwCEg9t/09uCpFy/GZcyyWgJxXn3o8/q0dI0gvQbMmtDw2V5Y8APPT/MF2rh9
ARAu/gdwYg91373fGbvdc3aT+JEORVElWHQ5UBVeczEzniwj3SKOiWnEOpD2wZW0
irogq+0uCfpvaqESRi7N/fxNf8kEE61kM1NXxihQ/u/7fsfVUI68Erg9mjH9bmeq
s9n4O97isCejM3jMhdDQcT/1pPZh3kMe9CBrRtAMy684VEm0VS2JNYvLcf+mk/dJ
JpZk8ATgAXbJ7+Ql2NuMZwwpfrf95ovZULdKh3QQubfj0UNdizJkbuLtqF5ezofe
eiaKIeUULkQbFEm/D8Gd2lAH3/ezQfFrtWk9/qRHiNojemTLvqNC2aZKJIfUGdoz
l71ea5RZdd5MyvZdb73yEG8ZbcO58Tgub0OFPzeVSLoAZyh+qtkqlP9TE1hzC0PC
BBoPal3K0KhQw86GRhJCPQD697vDM7t3SzEag757KJy/T2ML14Qi5kNheWliM/Oi
yP5V7aw0bqN82KJbdMGEl/FJRVXfRnRllwj+zGMlXPExhkWOU/dVdsnPTU02CglU
c/K43tSOR3xR3QSFjucvwDurEi7oSxP5oboP86/BYDh2Rrp2Xa8oEuRuZG6SAYx7
STwbNpGqsmRKWdLmZrndyHgJCkz+qlMC1NslSl3iycZ1foxUlycPONrdZhU3Su2d
1V2a9RSMdNl8Lmb+U9h8+HR6O0vDR1YQ59/55klykq241WN19+ovV6HTFTejW6uH
mmYyx/TVN1xVYm2PmVrIAmzeMftgLx03adBfiVFPsqUSyIYUYigUdtgUR1HjTaR+
PKx3C9Y5mXx5ng+iaIQV+jTtpUddef+QaL0WFOhFAY99yGmI1Fy7lAOmOn7Ut12o
dkF8YSeIUE2rZmATyGX9yGoWqKY2IjcG9KrLn9NNyn8Qnm/fDf4DY0kHqY4qvptQ
fVBNLktc+LcdH+3Lpz411nC3bFIIoYflFZnVO2jQuaXAsZ12hse1C/p8jr+6xNu4
ujSgWPcxfayRtRLBI4rs71GUWjBMWzy2Yw6utOLfJlU5tvu59hfmSKLlRzdzoqTS
4kj7dnikEy3XKrdqq/38t4LdkYUCQCpPKhalrcpmPX98vl2Bpe/Y1Ay7pjJsshzC
bOFeXeuwdwRd1oncDGP/sXhYVgG9Xmn5B6sATN/j94SjA4MEl9xvtoJL3KU0Ts+L
q7us+yTXKWs8M2k28SNd/TefkcLv9ZIDuPZkZBAWYUnOa8FI9fg4rVybItCevmQh
EZqWQVqIFWUIkUXOls+vrNer3W/yf9c3RKNU0B9chNKquoPqMKkTYfer54T3xSV/
0Es8Zz6mVrRtL+CFtAuHyaVtAfC5s02bi3FQPpRYGsWlTB5CBgTnmPrOUrlcnnBo
yfigsZNIIjpd2Z1PkdkRuIykboSVhWtfB7d6FE8rVyN3m0snr1BhOwlCDRLzAP2x
ievmhnyuHLluisRb6ytlbrA1Yh2wzNML5bCDtPdUXKojpXRnpS4i8HYn842QYjqi
jq4+rC/MfwZBEbZrMLhUgu9Ebb8vmnVPVDB+dSDfR8xoCLKWqEzR8kJnYuvyjgBf
8aruiSZG0hVLBTiaV56234i4lAJ+QbaktBfaKaRSkaO3AVjL2WzCwn0qgr3yG4DG
tvTQIZbOX08jMYaY1FbBah/0GXX5+m1KC1fnxxeRXYvdkOir1wpzd4m9xgiIWn+T
8i59qJ+ZAeyrJWASUdygMMPfeq5dY6H+fHiSh2THfR0SJlUjO3xTDo2rY3TeG9jI
qn66s55uA5m54O9hKUegA5a77mLDjjpVklG84mwkS/6WBZ4kc9ELwk779LJOFLys
xe32XUrV+DQMc9V1Vl+ZUWgCtSWGwD2WvZNRcBtpQlPKCraDpZMRF5FadTqpXXXZ
aMhO+55/XFxFtD7qEBVoYY0+uDDJ6jGyw8IuLm5RzY5VI+RAfLt3CSVuaj5nW6z8
YsvNZ7YTMWUpKPBc+hDhl7oORKw69XMyifWMIYDZp8p7xF/i9a+Y0mOb0uhkUdDC
3i9WAJZJW1YXfg6BVirxji+EqHR6BUacGVy0hHtb8US+5kyVv4erI0KivXtJgbpi
tIkRpPpN4Exc0eRPxrOUy6VRNnTv3kysd/S7PHASIGH+sBwgJ1foQDMSG7IIC2x+
0aoywcrnpzZcVhXG5nia1oUxgaJZQRsrtNJ3kZhI8rsBB4+16oe02WF07SfGQx4G
iGfUC48MazZOlRTggfHItoEViqUcclWmNysNPAOJlT2PaphjeMk83ovC22tVmE2w
8/zeu79pPWqqIgxUg6YO+HDEodTxq3z1nnYmAvxIhiVGkyGpUZzaeZUed4R0IX5p
ZFyjZWkCiCqxZrRhJGeUaeX6cmTBjd8NIlqzFaYk7mQHVAMa3rPWl1DZCMCE8sov
VnTR4vNYXc/pfqHcX10ueb8HLljmLUNmGCGpxNJ7EZRa8JbhzDNEsQImGd0KYXaK
sL2pYnhrj8c5s2q9PpCSlI5HxM9HXihuYDHq+E386rFKpq/KEYpx9Oz7CV6Ssy+6
5LG3onqwG9Op0F3qLDHdEI0dmK4Rn+3p4UB1oXFTxOv5KXXOprdwqG703OY/q0TM
jZZhYViaUxLoj9s/ivk9u9glRnab8irRc0mRLt98OCexQ83iO+4WKd0f2+35Dijw
8NQ8J3ZPkRRd18JGlQbXBVeFwjM+2G3vDQn95TQNKaf+gqgQs2c8I8hba3OsepGk
OueH2W5nNdK/bT0efkSufK9LdGD1wVnYV1Zq4NhixoPMd/i4rPFz3/sV3GpD6hCX
SsXDJNriUoF/VIcH6ckvnRHENqIx9U0Xn3xLa7MASC+qChtR0R+KtyEKkPd2Hm4+
+XxjLrfFNZD8rL8o8Q7TA7vLTSIZ7dF+77lAfHcxJFb54LKpeJkh6ZdsxSHx3YRQ
n7qz+uFRgg/r9VDTMnWitIkGNLoi4ZS/fMxjeqgrnAjv/9blXhVfx45f5Hyq8N8A
XxbCQhaX7l7SDsWiUVxOvjzl50I7vAcYc2IhugFYvL/ewNQ35uoWUQvmSLrmcCHY
RLbjpqsHZ4I28xDA8lppQj4FI4qM5anv5kQtMBdk7pFRL4Ge2jdeeTUURnSSn9fw
bwu1eoEUSC2Oz8osUlBNwkVXP0Ms/L3ShN35tAO2bgv2wIdMjW8j3ljmZC0WTWlx
XovITAS7voA9xLxil/0z6hUQ2EpLlPZDwKKJI9lg/B/p67FVmFSPrc/HLsYet71L
pBlDGZsw2VePTzRdvFC6usTy5Tr1uS4M+7x+JersMkaV11pyFK3kdo8Xsw6Y/Tcv
yRGBl4AUJR3hyhNyirKv4XuKyyY65k6rrDx/2J2Q7HXPxq7LWlKhlUfvLzzmp2I1
pkfbDBeofH6D4PAeQHt/IaTTl9b+2Y1jvzpuynmzbf/W/Rgc9VHfDz86vET5ND5+
WDm6MKG1IWy3DNcn9VH4fGB/LlFa14K9ClAcGzdB6WXBvGq0FYbXPruY+w5WWIEu
sbVjsZj0qbOBEo7SJDohsY2fsicmf+K81fC2jkKNSS0b7B8OUn+Pz7Jzayn+pt/G
nomGJhFNc28dXMg3lrwdw3sYGRwC5TN2vW24ax5Lu0zOa7RqLQMOeEF4DQdgZN/+
zjK7xa4Kva2mrh+86YtNCFl56DqP/0eM6arPRX/vqYPP8z+W4zjB4tVRAMIOBEyi
PTGWYzihzgsP6kG64DBwLzTBK/3Uo1IR5703oUaIMYT2+sIGDd55ANd1JUrBnqvp
rvaGjNw2hDUKvP31ZcrHyumrrIZSyIkyNvz1U8n+dC1cPQeK0flChxiSviFiIocW
RYej6SMHdEPEoE2hDzOG8to0GHllHlZmm8HJ3ycKKIIZcu/VFP81FppqrGn/YHyI
aPncX9KNR/+xPhEgQiU5Bp03VUPP4uGVHv+qR2bohRXg/z3zkB6o5uAHdWE1H6bW
akqrn0JPxD21ovisGKO5GGspvO6g5FdiW24z3ogiQweZWGkPdaUZGDargo//M3Fj
K+x6b811AVJc90MB6QXjxB+c5kAzvd3K56cwKkFD13hOsMyc7V8skfdgyCLTF+eH
CGazkNsxrBbvlt3+eIZWeSfynjR+3YEl0uWywdEIxjtu6cKndvoN0DljA6S1GjJG
oesY5EhWlGuBtEzlVceaQV13h1WhzC2tejbOSGjSzdKnyIkYsZoWuL2M20xRJ25/
2CvmJkVhJmuKdp8ZRyLU5ytvWEA8mdhMBslY7bLPxfLkM7UA0R/mMmeGk7pqvst1
r8RFfeayiHtZ8cb3PMJOcvnL5BiP24Im6nGnVcmTp8D91+uVsGXYlFjUPzGciaAv
0pGm3tjI6KgPttkwK8zA4EgISXjb6YyQPZ9e3TyfDAb2WmNlLKD5ghlWs6Vbt3jg
1kk3zC9uO46QEQD1cDsmD/J5xvKDd7XMKEecGaB5Ed0mjVqZxzEOJWhIXI7IpB0s
DxMkgi2VcwpTVcLVermopEg2cxGu7xLSdCJfGYh5RQWzDCTvUdiaO8Atu/2CmLc0
9KVXdfmC5GhVI72Rqi2Rg0ZtuWGVLu1IJ31kvoKfT971u/daubM16uPyBQ2d2DqQ
RQTJZmmC/qke1VruKSA9gh/RORoJBrRCu06ehNkeToM5AlMG1We5khN5GKVqVz3Y
XuOYxTCYtTO4CD1Z3txpmTY/8mAliY5Fx49lqfySGMaqCbix449ND3wuR+bGB83E
BTo+V02HMO3DxKXv/ZxPEpang0WKn0knve0yIKZFx5nv+hvpXbLmUbvUWVkJezF9
cEfBCMrkMAxhV4upincU4CCc4OUL6KGRgCYA/VBVFeGGmEuNAm1dJIs/t43cWnLm
/5U/YPwdAZ1mxfY8s1NpjtEYINNxhlLjTVa57gB/ZFKjhlck5fXEhkxMvwBi1jz6
LeM2SU70yrLgYFq5KP0MYdCvP36lNDlnCqnjlWRanJHHGMl8cX6MDKk8C/JbqkDq
8roQc7QHnqEoDrO48092jHa6O8d36dbqyushx35NGpiZQVjJEeFmS/VnsI2Zox/7
WmFG9pN83bLReWKzpHfUzSY0x3cqS5Qyou+bPpnLV1SjIVvePYVcugj56vRV7dNB
leBVZTxnY3V+Ly4aBn6uzwNWUworsNmyNCjlfNxr4PEpl3vn9TFvinLUy9CQV03J
vj85vl2+xftqSxRaea/9GvEByokz6NwEJo97KwjoUw+0DxbuqddhWQKaiwYvfc8U
ThDbLdl08TbKt9k3hmlr2DrcFJyQ/VamaIj/Y0Yt6FVXMyD0FmiQEVtJ5Ga6bfLp
oCufQKqTMIJWcxE+XSIHgKmAvDIBJ8fFbHmEG/Cr7ltDnbmbUPvUkdX9lS2HDTyU
XxcuTq9PSc3iX3UKj9p38/qWHlhr4XyLSUR2OcpN48RXGWo4AX0Xs9TBjmdTOH2Y
vRYiBvoE7GsxXmemLqNP1jyCkSreAWcfH8vsHwvg2JffVkTTjOv9wdJyAD/FqU0n
wHCNd/S4BMGtaZV9ofm96glnS2sYu6EPdpoYnKgKn2bX6RAhvCcTPVPPkJBabdjL
rvnyyNaKSUwfN0nJ3hMPuWQ6qEoHKf3fTiMVMAXNTIswBJF8ayaAL2qgD+CWgvgi
GsSb/DI3Oi0jZLwjOmuXJBo5YRPrV+w6vJ3I2U4QAE6vLYE/DsAXgkIA6HUdBbuy
xGBmm9v47uwNbBGOvu2EvBk1oO85HXAYu7S8UaSTBqW7lnuNPperBqiiu9X8DUHs
MtMN0aZubQHfaXizo+yhRiuvFCRTgaYQLmvRZHFgjyG2+ID+eig/9kshqX3bduSt
CcZfaYHX+ZIX4+BitqFZJOLJI+dGaSiUSj9K1aRbr1YgxVNzY9263fw5hlcWC9qg
8Diua1YqylBdcvKG59r+mMZAgSqSt3757USn9D6Q1ggR3jar/bDFVEpcYPAOlGfR
t79LAJK3H4cIV64ySeTr1Zvknq9HO9AfApKU94GhCbknZKrPteKU0cTOvaXvUGUb
Q6FxNZ2V4DCyCF6WDWJLZGfGyZaqGFPOpAf1O4wMTuhJzffd5LYbanBr6NV1L/Al
NVejMT0+aXoqrBPBCgDzOpn4NxbgeD6AuQeJt/JhAiMV4UIHexn5BuhTxwqa9NVU
6WTqEzCyUnZrrHzIxaTldFzCasE9wJuBZWXQsAhvXvtNoUyX88WHnTEsr2/FKTRv
bP16jL4JMg3SvBeiPWKcqNez2Ir7JeO1V5ohn+95WPlOclp/kdF9yMSYHZUoNBKW
5MjoeqNDmJ3yUM8B52XI60UBkeSaTBkESJvQDe9PamfyXNpDt+FzJtsLcJ0Q+Hv+
mKSjLV3ow5SDnM4hiPVaeuw0ycKcKRHAfjowudbEjXvpMamhk9XXo0Z3KvO725UA
lcMemJ5a3eqeXK4TbmY88WOhOVALtQJKpIo7PKRfbWgPe6Unp6IRPWCGWvEJJMr2
LPqm6fRBFX+ZDfmYJ4be0YLZgBCyYl5NwYwc8oj+AMgipbTG6U1jk8EonnMS/6pR
Wa3DWH5/xXLjcwNiFNU6ffvA3sYGiLhNzYfbut4wbJam6yiFWT3hAbomXQtdYDP1
xpzArgXIBd5BoECt5f9bIAc+ZCCNL5KDwSFacLelCX1Ip7p5+YTh0Of8C1dqUbBn
ykOAOb5senE0W1hDdRTmntxjZbfWPe1ZGLoSfNjuYhKOTTzCF58rqXmWRBM34lGk
o7gOWYVDGyzdpvy7kIwtfLq9WVOhShdub9zRvZ566NcDHHyI0pkkBA/KMXjaCxAE
BfdKwS+derW+yzvkiufsy3acxs4zWt8wd5dZp6Ac1uUK2birDvWqWaLTbzDwxuJc
Klm+Qo8B32/F/aWWlnz1F61dHsWc6nXVYZtm1GGObo6tHvWxg87XtaI+RWmbqe/a
3vTSQN9kflxPXU6XzK2SJKnYry1Lh/67emTfk/17igmKbzzGIC0nw5VPm5jb+z7l
JbcqyWO4VEv+i+JurmDGU+yhwAn3k5TVwqCmlGeR4iNizRre2DKTsBBFTqTyIUQT
XLsTq0t50z4IHqsjCV2Y/7qdJYep5KG8AxufbK/5B7Y7rs/vUDN3ArQ9bfuVXbyo
JXUAGGtEViPTSLZyeQ7t+dixhpn329Ll+4cJrnFk9bvaoA1CU9aBIcelTGrRAkyP
FsJp6rb4UCvke4XRJs6iesHJf94IZZnyljiAT43W0yZghwHeIs3TJSk3aEdE1EFZ
//k46KPTy4+sMX2l83rrQmEub3lDjGYQ6guna+QutiEshHA3mZfuMYeQ+oIiG+dX
OJMFbx0b5GUZiv5RpYTEMGhFVEq1bD/TNVGYBIJXjmoKO/XxmrWkYlvn86Z/+IQ1
VITWt2PN4/ABdwkVwDloBwFNVb0C/00lt0r8VUnpOrZE8J2E59VhbE3ElpK6m4DH
zJb8TobYMbevTkQzLARDZECwFzq6N4zk65unYKPDPSnFQd/JR6gcRfyBXsptAUYN
oI1A7cePfl4eGIj/4RoIqDlptlhz7BIl0gCzuKFcyrk2ReTP2lijoU83qzDYeh2A
g8aVS3TyosBahBUZLuMNzxLyyny8l/A+L/tm2a2vUVHdC4aSiyEIOQ1S/vHV8947
4XZRAPsF/9LUOqLXJ97UqvuBqP5fFAO0F/5Qe8NnjT34BD6SLDiMuPT3Zj1eXPEu
pZSHxnowNOD1P0uqrT01psTwJV79sx6YDaQO0+uz1pw62CuPPYfZ+TnrmWegKMga
M3KCBVBowdXTLRYFeUZ2TkJ8lP11ANBhC011sVZXWJFxLheJkN2HAlAjIh77Rlbu
CW6abnQgTjyns8Xdn915Av0F/SoogZCNDHt3a/UhutqpP8Y9V7rGkv3jZTzQ5doc
tWzNcjcbv/+YmXkWS+q25YwEwTkLBceGeBeFKZg/6hP+E95yvbM01I/8G7+5nGZh
lA8Y/N90cBJiy0wWV7Q52IGMTS/p5Mib3nuqzC065WTh4DusGGPDQtAgjseVDPaO
LjUe1GiuEfqzNHTyvNy+NZyFmOIFKpgnaNv+IvakRKZBOHNlHS0adlFwsRrinNfD
05BwwDZlfL5Rt6y/Yp4HSGPZSeuTydptRexUu7sH0kwcldRAX6u3hrpJM7qYFEkm
LUnEhe9sibmI0AAujz+YBaY7IZqVjHrnm8c0DP4zzrrQZBoE6Ipvs87CU8ReDtMC
90dvf1MfpGJGuy9x1syL2aQZbmOBEdVAOBbrM5dZpGEinhxiPVZaKE5z8+Z5w0Yb
RXbaYauLAU7R007HP5fsNALvcifFgG+1VT67JYMKwp8RXhQUpjoLcSKmA6nJIf+O
HseoGkQsr96+kpalEBaXBtG+iWHVQMn/kGpjmd6meoKBAnJsIffUBj0hCAHDF8SZ
OkuHmCwmFQzFLBL0meSCaHtLPMzkiaP/FWddqVKrn3EBFUnTIBLrRjep7IteUx3J
HUl1cbgsX6jzmj3PR+LGjnai46L6AoFfL0AmYYzQm51WimkcxAW460ZP6pZVM7LJ
wrEspfqHef1YeewvwskW/5DX1jb1dfU/oc2AqH2GYJGmhcWYHmZkRwmInhKxUY58
wFIIaSq0dz43hs3eVhixAa+B/QydFewtmu+xTEySQWDK9dU0vv0QZR5wKGz0nSz/
W9SZJdCJDnmOE2P4/IjeBjP7hbT1ZlKqvKZ8tAFlcSMRb0wNFTfldSU1xYgyXUWS
H+jVOQSaaqgf3J2ZG6FdOK6QYjVVF40XWR5RAaHaV4+yFmYSUZcTvi9s+r65LpK4
W0I/adtfSSiiJtJDJXIHKMlqZs7UG5P5UCFGEZRTE1+BLSQGWV9pFuwA2eEJj5sS
ey9p6WasiKFmEiG2/cxWwn5YH2jIA5QAhzhNyQ9ZnvRQC00P/j/iRDroIOuATyty
9tbpkseT5TQT2BM9W4e8nHbXSbs/KeCQE9Ir8nqjBlHpG9LPC02pCQiogPo3aw7m
lmDLWQ9BvSDuhqsMZGazQhgMRaH7FD85n3hNxMcMNXkVkAXYyhEnptEoj3kQegXQ
9HNHQ8hiVBdcWd+r/7VP/RdIdu9hXZ4ExjTB+NuvpxYWlryIHCOMvjOLrcoSP12l
iYHQMDx5phBboH6KWlCfkAQBeh7rNTM0S7zBcXer6H/IoJAn3d0FLN6Zbz2AxPMI
3PqmsBXq2s1wdylkdcZ4w5KOkDlLp29SI74dX2PV3j/Z8gMPwexruVB9lvhMF+Em
LnwVKBcvrlXEUaaT1r0TF+7gU3cwD9jrsnwXT1g/CYAfh9mfx0toteXXFAXaE8cP
pFYZB2XWjRAiSRn83jbeMn+2LIdCiXRCAldb4rfHq8PnhDZtfRJOSMrKNTqDjg6F
6sCzNeB/F/ulcZJCVLGudlqLdCDw5wKklEiqZ2EyAufI3LvpzGi3T1/PxH7nTkZr
E91V/e8BEZdeOng5icWb2g19FQKYXLmqAXVo/pEUMBB/KHxpjw5HtjOb+KZtBWD3
0SJcpXNm3P9we53v2JBnK1GO8M1cDelUTrxbfqIbEQwDa8mD7MAxwjascLMw2Gt9
fAoeahRTxM62BnLQpCaKL0gtKVDqrLkfoK8ChOc2nV2uiyPJuNFk+NnfH1VzbvQX
bwjHUNV+zevVerQsPKV+TA/fu86OSvOOOzi1BcwmltEVyr/BdW0g+AoCxoe3PcF4
3HYuqsBpZ993OLAAFXA6AO5HhtnjkZQNYdZcW3d5a82NARxdk2jJ5IsB8cwWd1bF
oKKQUB6WHpX1MSfK5B55SqALW+boh8929+Ze8N4ErWvCmEmRWF3WN+n6mi6SMcwG
VD+/tNRrlPDt/LcmCkXzo1OOaZN09/QUv564fYfcxMazSdb81l7GEPemURTPubP1
PZWfP2UvJSwYf0aAaiANWL6glgnrmj2mtWCJKdKTVV6rI+iyh7y0mwlSoVf+tVTB
9Xt4cWK0KXDiixxA5uSQUZ6LMHbaIyADblrG6VGn55WxiwjUwljeZTGOc2ITXgW/
yfsQTHRH97bF0P66F3gBNic2nMCs+ax+5Wg6HZsBIhIwC2uneDudkvA9QIu/+U/s
GO9lE4adoWgl1D0tA21SAVLz3WnSXJEhZ8Pgkv9A1fqRzTIDyDJUGUx4OI8XEAyB
p6yMw1BMIEAkQcfEpdXvx9Zr268Z98emENUlFstv9+tDXaVzAWgdeQHwOia8dGix
BjjMLeYY00CF84hcn6Dte24rFASaiOS4I67AhLEMaw/rx4l5lg81X0L2BlMdYp7r
xtsLaZgTOop7lg184SZcPGoWyDbiHG3hjqob066NIF28nH37ARTSZ0i91p0DnvHy
Ocp+4b/9LCizMvZwe4TL7R6iojQZBdjaCyTGOWanwbXrBKxV0LFltFG4i8St8kR/
Pab22le78k3U443G6Zm44oJCCBryf9FF1nCnd39SYuZw34Bo9LCidNsT9PYu/WJF
phNlyMZxVOEkJBhSYnpEcoZJZlHHDshufYRtcbXhuw1gAchtqgfj4SBN7JqSYRLl
Xa1RWSSj6RLtjNAUqUOrUNyH/1tFktrZBRpiUq4dRNMDREKu7SR26TG2M/8yD6ML
RopCIpYX3+0hFazV6JCCMmrzuwefgq1dJflD0EngrNL/4ic0kWKzYRixQnJQvbRa
nbhkUax7xpJQaoVCfzyagw5OfkqbxCSVb7jpG1CAdo57Kh08BxcaA5eq+FsuQYk7
n0QnGSRS7mHow7JDkHnC5vOk/8Kh+Kc2z5PaY9xqre303JVlo6imcBUxqrS5f09B
0GukLvyq6AfXnKtAYtytfgNXXVXZmaMO01FQNMiiddp9pv7CzzabQaZhiT+wMxy8
gEXF9jBmMbrUwcwDwZXZLH9dvR3sFJU65E/dzPVu6X7GK6OBvHcogpv0HdSrBF0B
s+T9JDxah4kwm8HLezABg+t4XwZPBGoUVTyJw7aY7N+rTMSPfxUc9KPVtwZ0kwVe
j1iaTVaAa3bdgpG+H1Sow6svpcEMN5C3xquM3qxLJ4fiDsoqfEWF9fn1BzhhTahk
3Ojo7O9kuPYYheVl8/YTjMMUcPsnEEGGIJmPCxqu/C1Jil9lbnwWVVFkEa70naTP
lBOY+SpY9YWrm96mkpkXdJo2cwX6dXbIJzDq8GiEElGX81OC+rh7S8xKx18ioHTm
LMHErx5fkzCABBILvJI/kB3Mqgvilhc7VxGJkHSehZu6TGf7bnxSocz9OVTbl2Hm
LfZhIpAqd4skK71aePEgISagDDKSlLCbTr+o+8pXpk8GjMMOO/bvZ6hVuYFnSLbK
wmG4rWL0cOkHlVEn2MmjYwwOHFRSTPBPaz/0MhGxnnzDeegj7ykgYP/X+lUpRH33
nEIcCZmMrEt2x4Ewwu7GctPCUtZs8pG1H1ptol1V4dLbObZc41YV3yVCoXvSKJY2
4/fyiSLTvQPfcSBCWoZeMxewEhmcPyy2gp5y3BPkX2tzNxqwKRIbi9xNW61GhQql
sl+DhT9wODMNfg5r9FcmA5tMgKGAVt+rXRKUwoi0PcOLDfTTtz8/4bfoJ5l9/V77
B2zWylJhaLyxu8JA35J3x2/gOQzmLZ08fw/Oh6R672hkapDV91Kvgpc/epKbGZwf
vq/IVb64CemmxXTPr/LJeWjNTCFvNFWlrgsJVrQv5MHx+RQ3yxq+sWeZrgQD585H
kdbWVhxJDVT/hE6quFEPKLF0tNCq+/csl/1Oow+n+pcJk883pZsgEIPfW2/m7tfI
f85TogAASIMxuj3fdhvb8sMG/oNYBjAPUBeSHHnEThG05rrvw1IQAvDv0xxqAgCt
XOue8rz3z+XDViwKvnwq8+HG1SIGvjixGVrXu43XqHX2JjJsaVk5cNjRoGwDCxiN
3JUFnYexiXBLxY3MOUqWEWGiYiZDx9dGGI5mE15UOSlK+FZoyy+5UQ0RNFLGu84f
6jB1Z/vlZGMhR3kVlH/TNVrjMJKt95OlnasKekvmdlM78FxUnFstmFVvMzXkDWfe
s5ztBZVTsmJzrDps5x0XxrFVrlu9dM80DcihEtlEj+J/kIWdJSB+ZQFB0TG5021R
WPJw95beGlkhciEDPS4ubw9nf2i2DjROtnbfBVO4cKRyagfzsNQkp1NsRnirUspl
vtw3Eve7lwnP1Kh4JayHAApDoK+ombEJfExtBttIvicfT2YaiSEfSfXx6sS9Hh5u
hZFpFO/8wJxM/LKzDzmedDZkX6x8IoyigQ4UIjOQdlwIrM4RmdIeKBPAAWT6gcY5
K0uXvnZZ6XkGEfEPcnPTONBcsDiY+r+th4qzhfhlCsGbO3W8bdi0wAshkZZ5zLVL
XG4G27KQZGp4Bag4+Apu8p5VjYmW7nh8t2noZgENDtiUTonLUHi6QgS/N4AtQr2B
YjRrGqTMPKKyvfD+5AURHobcJttb5/uIPIrmaQIaFLljg/AUQq1KM/eBFhGE/BSx
Kx2umEtqaldDD09/2+Yg/wLs+vJjgZBJSo/7/IQgAh72NArPDHI+iMcCnN2Ui7+3
21GaVT5YPJo9PF6H+0mIS4EIjfAxw5obcpwzH8o7mSKunW9jiz1fk5t0AwqXsmxf
txkOCeDUhBbCAnHiRidXge9cfQTKGEa3N3VLkTXmrvLEQHmhd4wxCEwHH6QdURO5
MkmuFXv0Y9FVqlBuGcRfzZmlq4xQcV0Xq4fbXn5jlo+pvwM6zPtx4a9AdykMGGa1
qLJkPCOqV9nZdv5ar0xGPK1sPFuyeAU7YiAgfyXTEIH426lSu2+gc/ls3S2hgQL9
3HLhxfVOfBm9lCIX0wBvHqGtevN8k+eLJsMuYM9LIyQqZQarO7uW7YkDsPnRiVEH
qA7HbWm1mNL8Wcx9VITQVc4LTZVm5ulQNP1cQFfg4SIw8UvXtBXUxXB67Ik3UxC0
BcYQOJtqTO14+zUKj04PYDSl1mmdh8Dy8pQdSD8HLz1/xcHtxWgZLJnqozIGPxQe
5+6FswPW2k0LiEPjsMZhaySMHKAyDBhwLZvA2DadwIFGOpaN6mHazUXrg2TmKh6t
2rIf2bziO3BdDtPbe+2G3XnJHuDGSviTVxZYElGrz/exjGN3WI/wA7du/Wf/Kzyj
5bIe2y57E4WT6rgitvNDFQtyAVwGgUmCyrR6ClAS/kacOpdeMTuWZQcjL5UPbca/
oPh0PwAZO5ZgypItob6HLXcvENNcSgRnIJirmYZxBMf9QgELNSS8AWornZngzl9F
WYRFVUsnKj/HEbkbVAlrqt1NI9OI8Eawb4hHWyVMlbKTWRDjW3OxA/AibIFxtDBv
EKoLlhm6wHyRMaz3Ra2oEJJN94AxUAejWvWv7cRkylfEicu9TKdRNVdecleH/N9/
IVJDVwBpLiSLhND19QbTzT2g5RwCPvOHJlz/YjZJ420c74i2q6LfFUl+/ZbS9LAI
1bO7U38OtsON81VKBKKYfpotykkGqmOz8IK3+0SEOa9BPoJzY2uiQSLoF4fEm5yo
uJO+KyMrc8Bp7+SnJWQXYhF2PpDAAjH9FBlIZjUKrQahmTUTFkefixsmQmmYW+ej
chJaHTd7vRrf6jgueKBHYCVeAsHtCpv4Ry/7+zM3HBPCtgXsGmzVY7vzv6JGrPQi
r4fxqMwMlfmwbwwsUVd3sVWp1Z4PkqYuQibuU79EFCz5do8qYdYTrVgp3AmtNvZA
LOuusSwICbcDFBh33JUNjJU2kQPZ/DnMdQDrQCm58NYFfBVEZK+j5xBQP6fthmbt
JaTE68RkmrnH0T/mTyH7hLMjcGvS/G1k0ELEKXhkReWdP8box5zI9RiW0MgNFT4D
dCW3VAE/KvHm/c/0s56DBZ+lc2N1O6qycw/+gZpUMcIA2TEhzp60MyK1JyV2rzdA
hwnDi1MHXOMHRwD9xSb2RRpSxPpLMFfeJQ4w0HR2luhD2nUCkrkjeGyhOfPN97fS
raZb7ScrwAOyc/eKr5taLmpJjMvyWWkQiUQvG8JZ3jkr+sMIXcGtzOTHufIxaLTu
Jb/HgcWehBy5wC7mqGc6S3hCIws8AXsjYHWNL3PKWqY4oirq3CkOvTptqQ+8VYV8
OL8y7rx3LLVMofanapq3cOlWDGHeAGUu1z/dyhC9RE9RN8vQabUqzAtGe5EI6AR5
DgxpgcNGKbWf005oVnnNrJRBh1ZeaXMwjCkfcbhsjJpn/ppThjeA3aDhPDDdvNqJ
bFLfAjKzQT5elWz56/QhMbf6V3vP8Qp5wHu/dzWgEdUEaC3JF1zvdTeE3LYcO76x
5i8dE26ZHG52huxnN06C+fha5lEwv69nk1fqhH0Qpt0dGQuyPHVfBzwhhHRDT+Wq
ILT7uSTCT3R7JLw2EgX+VFaQ4vLjpLf8lDEi7Toa5/+1pckwg1kRJYMcRbIr2B23
b2uIc+/4qS2D5lbnlsQy78l7Bki+8/OnkhGcouOHI9Ygct9OyvXabNgbfUpRbPUs
sJN4gTnwOp/HCAIuoELsyyoQ5zY5GkwbvgQZGhIKbBzIkUnLAkSCI4jROtWHFf8S
d9isuYCeUlBO0pbgjJ3vtTuWKUwTCFhdmGAc/0mjZk/Ej/fJrhfR3A5HRM1lPPHu
gL5eLnQjPGqw3XgtpJLF+adUkxhPdfQrqXs7rUusGZoCd0VPcZBDKxXF/z81273j
kPRHiKUd1u7rauCn+6a9Jnx89xNTxAf64ZaNM6J20V45ERL4M78Sif0PtNmwxwfB
DHt2BY/u/HXuISdLv/Lm7HWXzd+fMr7DhUfQiqSkUw1JzT8026Ec6raf30KaIDgA
oEaUdu3iuiYOZkOeWXMcoYVQ27KpZvADb9ZbdHZ8DesYPX834heWBdElsBm16H0c
76rYkzex0NjyLlnd8gx+DnphEK0vhZT56HOP+ZuYjtlqBzJzC3DtNsNtGTJtasZw
nFqBxJmJBVTL4XUkovpnv147fGyfnwgZ4V7T5EMXzxMWtLcSIdWG/K1R24y1wBsZ
YL+E/EmNo70coXdTahcF6yRLK0o7jNuQVsscWHbZUsVBsGsE7ryvLK57my2aV78r
TDNHgvut51ygG3fjV0Y+u73dJzX6R7/IrWjrqoYi5wF+2lDM7l35zGmiGO6WUb+Z
kx7bXkl4w3f6VggEO8IFZY2iCFUaGv3h5Bt8CtUlJ9lc32I1k6//BygmKXVVjdAM
wcy7FHBzsXi+KSKq5410ZHoPngbewl6yOp2ZpC6x2mSaXnW+itVQlOb8P9QWJfud
mK0Amo0po7pdD5sgWuADTsJ22kSojnxlnnnrrhogyxMRaVjfmNEeMBrueDUcd7Sc
IvBjchTtQHM09Ih5fVwNG1q+76+QCTLQvjPQIuMxhELMFpPW/850X8xVXamMc60J
/gDgFyecnQEO0gtn2XvpkvEQYLMdxQBuDl2Ly3dFG9fRz5wrV7uE0ByOMajTd3rB
iLnoFen/Sb4dYYJdMQfCCpXBPBVkOVnawUOasTYJu062fVSya1HoRtPq6nVz8MTL
5uIVE8Dbr/krf2iK3xH8LcqXYIXs4ErgeSK0RXxc3bbhLzfwqQt7TRTzEAqSjU12
13w1lZ2feizyQEm+fr3dHh4W+JmocmpwvrS6gldqBbbJv802OPc5Y7TfvY7ea5q2
SR7To2H/XnQmUOhd2Ti9uRA1nHAIdBVUIII1zFyqq1jxtHW5bR7OR/UDnATkTzmV
jryHiBz58ymX3psTeXirYkVkxcFK1+bUN2kDFKHmDiQNy00sAphdEUokjC3V6A5r
llo1DeZgiv8fM/8c3bh6PYSOEaRMIx5swj6six78+3uAZTkcCSs23rhCyXaJbMOy
b/dKt89Ni+WIxEts//56btCs4QPIhRRiJNm3Z9XSY3WjUIWu4SVDY9xvIN07BTJW
eOh79vkghQe/fEVWnyxOZ5VENDFl9lYEuH/nWcOKBprf9KYWlHQmekRKCXAvNS6J
WKNk8c+32nMnkMqW+lo2FDVtKrEcUCbZy6glqgL9sLsR41bpxSJaoQ5CjuHZT7bY
dCSbd7AOWbFYfe4lNZ0q0MejozF4dH1RGBU6bSn7o1icXQw1eXJEDQnEbmf46ORY
ld1K9r55IYJoTeIvu0Ym3c5zBXRmcG4d0mgoHMOr7pb2W9lOIFRDWz11FzO9GEvK
Ki75zhipUZ3TYxE3Ci84l05j99xhkBaaaWCfbYMPmsx5HINP85WuK2xhB68PFXDi
1IPtj8h8gARIlltw8G0PoqswBrN/WsEBhaFuljfRqkyAD21yhshs7jTtAizVBSof
+AepW375I3VXoEzaPyANODCncazGmfQoK/0n+A7KtdIRSkcMnl81uaniuqqXrnNE
i47Unfcj1hxq/3WRStjB5bMBU41YINtIFO2CFh5jB+ndB4kmvN8Hn93AupAdzd20
XLUgNjsh8IjJMzedYl2riSLL3AptGBrfWU9pJHqgFv1Z7TWfFFivMFljpZz7tiM/
h/ayiDpYt0XKQpyNbHWiMu5MD3tDV4ACh/KGuBMA9fkVRyb0NnMvpet664vJH1Fz
jSYF7bEcGRriU01xCxdPsDWHALiIZjvrZW95M99x1/zyWL/MwCJEnU0CdR2I/dVB
SzAlO13N2Za6gNjawSzMlwshWJKs5lKPph7d2hX7ofDk3vlNvANwCayx/6xXxXZj
Kw+0ToJg7SPNWnkNfCE2hTRSAE62Bp8oELyCeWZFCKjAGuAqdUyxxyOXghzFSohz
6Z41M+15/zZuDroqoSlq80YepgzTu489ABn6Q+WpRb9R3873wUp2vBFL8sy81x2A
oYggoMHbVOGfHPDH0q5OysAmjSD4X22fm5QKz3l7LcgyUjJsM1I9ijRcYJquQAUQ
tGulSctPUQlnVl59ySPp8C6k4r3u1p5tmXBi5rLILtWEyYPwFnlCeTAvEsNJOJJR
m3UYeYksKytwdz67ctPHPbkFmm7PkU3h2pmgsbWYkh3enVs7PsSoYbolG1ivdYRy
ZdS/MjNg6QjKv1yyUT4+K+0k19qXucvbOJMCxJIDRKrHsXaNcgd6gK2qof5Mt+Yt
1crCJeo5OH3sUgYBd88AX01rZjfMHWlSQzQ97rh6TAR4QORIEHYNNfhn0+cX8LpK
tg+BHiB25ojF0CqQtnrX96Wy384gm8E9WUe4CzmUHzIPYInuRXe2D/cC/L68HGDt
nw2fkghxG3UXOaxaojuzLMXBSzAqMYlIa0oHcjYl9bM4yXlLqpZBlH2sZQTPeHWD
8pNGtkdN3jqq30JoPWexgxqIoHhBYeMpIBHUgJ6gIt1gI8fch+z5gJjtUsww5zpU
9EchdvXWhlXmYLz7lhICl724aN1oFI6IevNJA5kHef0OEDYeH6lRi+fzbc1doDUv
yV197/X779MTPQDUbU0ucLTkJJ0c1BX4Z4OwMAljTEa9uB0DnKOr9ywRrpbN47AS
dmVRX5h93hPrdm00MV8POkzHEzC7b9splok0AiOcxT5aB8MpwI6Wlvnc8GTll/RG
EROM96imQruxrIowBuhnE9pZVTk+GNVkiRsYmXnjurf9jThkUr/SEfoh4p6ZSd2M
3ypc4eLG23RU3vTEXBtwgrg+ZPCwVjL3n76hCBrM6kPSAq4B8CYO3L81l8janVAE
sC+QAxtqMMlxMoRqzgZKkIUbv9lb+8tzfKlwXziIJElAFRUitHFP6VhEiSN7nm0S
9jEVt4ERWLGkqHsgw9zHBcSBiuAGr14vKH10lkq7B1/Vt97dCuKeOzuZTcbYEt33
R3ZfOGLl2ksJABMCQQT6eTQ2I6wRle7nZGITTS7ejtVWBzq3SEdoMrLArG4EbGqF
U5bIrt6g7VH0ekJSAdjVLqmbMoa28MoYKByz6gOpj/k8OQbrC47qjv6Gw5VRHl3C
tMcgjI+UghYrTWZS5bGeaakDmwNqfeXey9rvA/fr+SmpLIePXEFd6O67cym5dU1R
9SA5orp4cznVWNvRzHRCyIOjwPNV3Z8BGs8zRTRTTazz53Iaq7xKa8L9TL8lJCzl
dMDlD9/MQfGjVLo3ghzOpK9NU7XEkH8LfNwBBl33UuOJdFgpaK7rE+mXpxHpgIC8
fdjZOgMzVWMSwqbdNw4aFILYuHQcBPUSdToxAbDUv2B7A4LhnRwipuhLa95ZxfFk
m+vJ5JpQjISe+Nya6GXVukFvtvDdX4VZwqpmiTm5C6tSYyNmWOAgeUFTrBpMQPIo
lJh0LyorebA/drnGTqMYKGQhvUfYn931V33e8eASqqs7tKg+yrT1vGQ/wItUWD3f
NjKJ0WrO2kdAXoHWfp9tDEKhPReCsUo6iuvf/ljyI2XYBBLaMSZMDAVQmTNxeloI
v6anwOupI8sHF/BnybRUIi0Dmp5HHKyjW5mVrmY9PQn7enm1KkNL37+7mKy4mi8x
jLffMDnmDJsh7omDDeDGkxQOVHeaUkp+I6Qh+VMEyhLFDHVA9Zdz2h8WFPFRFCCX
M9ig3EaWImj9AyxTGNeB8SpzhYyiDQDQ2tqcAZEhiFII37eRsGbJxi0iQXnpqRj9
7Fg8TMsmrIWMUsb+PC8XcA+Zm5Bb88u1Wiedfv0us+qw1MugDGDSEv1j0LLeURaJ
jq6QAdLkAI1B203ZWfXpKtHOth72KWyQfrqeUKziXfh4n2N7FW89fh7db7goGHEf
ZN4oDFZeK6QzQeRz6rt/lqOtjyZFPfVtBb8LP59UTXcf8hGbDLkG5MT4vFjhzwQ7
Ul/eIgVBNS3yUnp+Vxn58JSYfClkV4HQOmGbfsyq3WKbCloyuxwTBlD8+HvJY09v
zVoFIc5nJI9FHw29bMZFreje/5EgT6SaEgZnGl5jiHKmfvOaszg5l1pZFskxo7SR
GlB9sKw6XFTPDC7gwUSRZrZf5nReSi5iQl+2Mfw13zJ+IYIqROFjpdr0e8OCjUvm
ERzn6YQiQBmF/yd+sSAN0aHfmNnrmU+lMSrotLZTQrPZr3Q++OxiRZ3AjojZuZaX
HdAKe1iV7Rzkzkw4PHSzG35nWKOBCJNM32/LNmChF2jiEbPJcyYBwEPcY9CooCc1
8N0hJMoQ0zC72Ye+vJMIJyNFM4ji6Ta/7OKiJ3XPc+woyINtW1ftI4HCjgtfPgWP
vp3ahovwiQEdHfCpOBNji7dvsggCGACHuwKfXwP9nSen0bRdim98sgp/3vZPKP7I
o7E7Bg/x2RI2aG7C10Yd61ZxjaCkOMAjW80qyI1mj48d6uLUKha3sJpGzHWehGGP
xD4uY9rSl6YwB0U4GN2rvyYmCmvKK32q93Be7PPV185gnQEEpMKW9UtnBOBC69XK
DbtIoFrT0E8fXupNpbj9Ddj5WGcNC7ER6dFhwP99Khm0VataZg/zhcYWG8orvuPl
bYr4YrXUXX+//uJqb9UHOSLS1C0gg4E6I5gb7M4lPqojDCsxXbt0tYygwZbxN4Cv
K7g//lWz/a6N/n9lD/KXgNVfONP207hRnu/WWZFaK/W7svVEjw5MKIsPDTjJKKJd
alO73BB+u26UyXHJaXFz50Cwc8gDDIsgT8OWlDiumK3JW3yvrfO2wCTI7kricNNb
3vcF/8bGmYVjAwkVlK1Etb3HlbTMdIJ3x9C30f4A7wN+di7XWsXYrw3doCM32OQk
0gCQA6XnPQ6F3UE6MxOHlVBQPrIpmnWdIBZSlPugpeP2IEVv6KP0pDtqsuupD1zo
g0U9B2PMK31pMgfeOgFB0+Ma6rtq9ly9gzBZgDru/uD6FyvTchKMtV5AvDbSQahs
85Tg/j5Y+bhFsrPwWFYt/15eCoT396RUpj8Oj2OQ6EVmlgy6850v8buEo24XHIjF
D5Iv8B57F1L0ccxEa2s3fnteeiWz9yR44FVGk7J0Nlu4m7WvaRLhg2gXCl3KdzBR
M/XktPM4lc7r+RIS6e80n1TQDlG/8WB9Ntg5U+2rAGdwphZE0G1Xb03nvG5Y8Lul
AikOwFfMobJ/s6e1V84WCr4YwusrWnyLe0kUDkCPQ5TMUQ3wFWf68aw4OB08Iadw
jdXnguGafCeHmxYz7EGFsVX/QWtgG+BOhgJ8j6QWWQXOdilffJk5gIIHa4dcslJ9
izddwcDfZMI1WIT5599HhxL4zYoMobXK6UVxhj+HEvGPZ0V77L+X33I28+xARj1+
Vvk0kOyglmEkK4rkwlmT3c5VCd5pydrb0MIFKqjxVGg1gQmTlzp8r484/8paiJSG
00UwjaiTDE7dbumUMD64fpZO9zbNWA6I8+Na6z2e3wD0Mky1t4FYDTMH3g5xoRm4
xzoDW0rqny08PJLrOl3B7fuLISZ7CN5gcMG2yUqCyHivY55+pA8zjEY9ajdWt9mY
J0Z5F0CM4kLi4LuvUG9WkiV/r2YzL6ijt1nEQYNFCcussMCKFB28WMEp/2b/lWUv
EJE77j4DyuTx5o6Ze7x3E68b2jQwE7KWLN01+ImTWiObCVK1Vr0FULGvsBTudiCE
CiqcDne/Vg+HPdSAvMD++4c0tKFkbYt+peIN3zOD4vKaeB76aQ70tfnNuHKHtvf3
hdedloGXoY7NqTxNqDVQb5kIs8ZFcUeIW8yCFrrsSFKyH3yprjv/gTZiq/RnIlzG
pP8HPQ/kEfINOjC1YXx8pxYR9ACRZfy+zEX9yBos4I/sKKv3c40iCE9gXTYxKurm
Gaqg3aJ/yp1EWBvc5MEUZzzY4dajPiLOwig4miRNqRo1xzbClXgYXlaKM7QUPBlM
W1vUSKR0kNeN+exMwoJ6WeJ7QrO2Q9Ek0l36ZPbO4MdLFDeGahzU7ldqADu+2za+
y8qxy+2fnOBF2w5vxYi99N3ZYNKcRgmdps0KvlOBwcV0U0UIhWlgMmVkxIYdXyzt
W+6GnTNzlh2kCQN18K2DEFatZdY91TNAyuOmx6uumlqodVf5yAKDXFkwgKTKfEVK
0wY2hdkV7m1v6BhUbYfo3dVPq6YYrNfnn/VtB5/hHlFilFd7t7iE0LL90XzvzQVH
3+jDfKRzkW/DALsPgtlmECZlqLhXKZlyiK/KithplhP9/OTZX3okIGUUVdR2Nv4z
jD5jkaJLw2Ok25KRjt65l+GZPEoNc8DGWRtJfREWLO/n8LF/rvgnCPNyEeY08Rqv
K10I3d6d/Vw4L4unAIj9WjHu3g81nzP/GIbAuA2RBY+WTtgIPmvxgAuNg8RAuEE2
qXjJPV+O+/ndFuIqP/rGXXTFBJYvyB8mIC1ascg1fDQGzzbVLhQrBT0fNHEvrgev
1aGHv1gM3muM406KcfkQ1/hLAVq6Rq2x283oaIRk9Klu45ocOeDOt3HpcPTvrb9m
awQ0xh3HhFm/XSal8ab4eFEpnR+zAfDPjA/17OtjYCAqqzI9fnHw3POV0Pbw9elt
2Qx70YrkTCgnLn/WfXh7tZa9ca8PdbLjv4SO148XpI3rIHs4PVhQMnRDj7VBAnfP
wIPHg7xeF7BOPWMYoGaNqh3bBaqtuw2YeMCAmCjna4FKhKJPUHucDrnGBHf2h2Wn
adKcAC94pfUSsTW9kxl73BkJD0SqTeQAk+j/atfN+yItbb/G19c484L0/xn5sxxo
b2TSKmuFLsjFxENryLZ3U+it7jD+pcsjRFAMqKQCyMRfdQC9Y6IsfqkKNtc3Kcag
8tpztUPthn69Xxf3rm6ur6Lsu4gllnpAmN0sKoyLfgBQIokXfpnybQEToPbY0zDJ
uLLUCCkmyDbtljnpavulfcoVBShRKUekLOXStbM3Aju+bU5UXGaTJh/i0cWblxwg
LYLnSq4iNdm1hnjiIza0EG1I6ytfv4r2xCEgyOQvs1MItLD13Ut3J66leGpROgwj
F4gZj+ery1Xc70kmHrO2KjuPSH8scOOx9fR1r32GTe9PhkjDwwdAW2LBukG/LnzE
cxDYt1VKum60Y+gengwK/IagN/iZBy1xvaAbo1Xabyk+grwNHNJE9UZy7beEF8//
z5SjrrN3onBNzyD/4PR+S//C/zly9aDMVJ2IXsBnH1v3PkcgoOV0cCa4xvX3qzRZ
PGF+SDLdbRTD/Qu0f1wKIGy+XRmx6cbuzJ1OK8HxdWHR+dYQsP7O6yhr6LipKWuE
FQHLdgKODLF4RHYeZez64SQfrvUUUluKBRqTeRKUB/14TDyxzspL1kaFHBchNe8m
uQrnxWuHe8w7FS4K6g+xQx+dH3gTCmr+JjYad+079wTXcmobo3957OF3GOtES3Ff
E9+8mTTDNRiSs+E+L+p4+CcuieBCAPOGqO9iz7jgpA3+Hsajn2Gj10WAskRW+qHo
/bAVPy5XeZF564ZaklU/ZpXPlvLB+93TbT8eoPUVquleCKu6NAz6mTTT+npnCqZp
18iY49Myz5lkoXQ+Qdzey59QNQf4R+yFdkA7ZNY/2u2FTvUqgvSlkoEWKa/GQ5iE
yDdSV4d9/nRWLqAO/JdDKpywGy5dmFchmFRDLM1Q9AuVomH6toD2w1E88juAqr0Y
cOZVL20vAQbqAxtg265Uir+9iSB1UxQVP3ZuUe9/HnEVMjy8RSoWUb9ufv/K+eL+
YrxaiokakV1z0iLEmoYcQTsaMWEwwu+9YCxrr5S6QrUitcjgONaS2ng6nuoMSCdo
PluPXB/8kMjZ/O3wJgE/jdjdJHPoT2yqSw7PJXq3vveOe4WTEr2CEFhnoE3GHQv/
VcU7EXbWMSHdPyTdyY2pX78wL7GAklXGmhgEC+FOvVNUjlwbRHSzxKPqridA9i7T
i10qTtugU4nWCPt/63EiACwkSwNS2A346U2JrBVBa2U/mKVDfZAoNqyk4WgMFnEB
MIDhXzlglCr8ijngiNa+xcVRafEWMaWb8zfUVa2hZnLK2BG85jST8IJUNNVBNfQr
36w8Dq2r4V2WxH7ZceFWGDBV+9A4DLifespVFq6IYGwh+cmE0f1rdbUI4Kdyp94d
6ew70p/SQDaTynvMx/KdHllQ3Qjx2DkcX0bqttx4R+6WC0jWB/Ip45Lr8lCkZn32
z9wuzP+3BYr0VeDsT1UsX+17rDVfpRhrHBLbl6m5QR2slXRjNkj+nPFXDgvQrM5P
Isn07a3jt52cqZi0jmnJzypZbpCmF4JZVcqW1e6wVOM67FzceAn/ltfa9Ulr879D
RTQSLjiWMHCuINj8/cndvMjHPgV+VYb5BoEceW+rNDSv33zd7PSmZGk1v673STrn
KVdGdeC71bw5fUtuWQjljFndHWdpqtLeN6WKsfmtxrY4PMOglVWg0Q3YeMqf2qgD
SqqK4uIMtF41/NnOEZoPl1lfRqqH7BNXU/2GSthpqisyXJTM3I410vZYBdV1a/cW
r9+yhB7fcgrm/Ah6Kl0hmPSjfT6kXPDTVFbwzx/BbPn/gJZBzzbWvC3ISitFp+j1
AXK8L/4LFrHV7lRHs9e/iLS1c/f0Qq4JrbAC+p/Chp9hoEFE1Sv6AUmd5WimTvCS
nT8PPyUlz4nxkH15ANLTgV8CT8VM09+1/+ZPRnbCTcmXjes1unpC4FeKK0Uhfo7i
NLPCK8faDCGuHA/DyDHHESWkSa1Qp3O+AN/tmYPboU/rZWwGYJcp4UXzz4nt8Oa0
hehKt3DVT8faEWi2k0TF9033PoOL0aVkQ1ENXL1f2V1zKK7xgQVw2Zb1DSx2HoFm
HBpq/vH3YqFrRANj4/cpGvmqF7HLJmN3HW4jLVVU3YEoyOzz6+O5IXnNUBaukWfx
G5gkRWgMxgLvM/JbfY3M9KzTXmRyZyNymd+sHFPa0OhFSIkEGlIF5+4QNNcg1u8A
KpcWA+zrsX9rnCXaaBfGRyu3PxnPdy9UMArleM609ZO9t3Fb57L4vr2DHjPnAvCU
VU4frSjY4ZG43dW/vy6sMoxl1d6KUnvbuK+xlZApqMRT8L58abisqKbgBZeiqpZe
9zUzTggUAc0/StMY9viaWQ8M3Z4KlEE7I8z9fOaCoDUT6RscCHyflgjILhtdgpUj
T5wPp+A6krqK7Cg8XG+wvhQmmKeIadCsTqX2ka6UHl9Gx/rhOkg0oQZ4kRobyKrh
W7uRPUMP1l3YoXaHwTZBBl61o2C6g+ap72VLpaO+Cuv9T/x9ErQQ2mEB66Bls0HH
9IMll/A3oaK1C6sPTSVCsH7BpM71qlAepnkksp5/zGeLezqCUA8WIJz36t7ORy28
HPfqkM8C+/uNQUh+W9MP4n6phF56PUAjyNpC14pQlmYAT9IzbNcckKfqZrnsnbmh
5YhyJ17XZJEGqC/GVc7VpW6jd6EgXI4/cijM6mxBNwfYrDA/klLPLmoWGWy5ImU4
ltY5RkQW1nW62QC4kcqSmQOitXSveBbwoRTievIwU3NFYUfq0AD6qu6pmGAytnQD
exj6OALPzgSHhzrq91rrXRyPtb5My7iICifPX70PiZarE5Uen/0Nk7WhT9wIimvU
mok8UnBtPipeYtOeKMbTqpWyObjCgT9YBqb2qR+ooIitsYfnW0wi6FaFdfZuusrL
go1V0iebjlGVIzMOLQcOjXpezGz2PaUsIPbEBQAk9ROCobF6pIn86MyMJULZsktQ
s7Bw5Ucv2Nv1CgT3vOEfbMHg9PQYs+K6XKMJoJk3KQKrbidD71yts87Jt9OHWckZ
r1xkwPxuI+wjxq/A8ymadcbyTW+Z5pG2gButO/+eTT6HXJgHf1hOUrL3XABQEjfo
zrQvZTcGIDfzkHxUwPhg6DN33QbpIQ0Z4zg9VXbN9QX/oei6ay/SV+B58Lnx1SgC
+4NXogEZeLuGouDXBTS5Cz5CXyt75FXdf/AJTfYixMPADK+uO7hyoGhvp6rlFaVZ
EycoCgipjNAQwElROCRJEIEy39zCs+It6hMQEH/bT4c6z6MinQOninCnEh1EVg9U
pgTWYALibB+WiIUnE21+ZSB/bgvTaqbNz1/QHKB9FdtM7bM6tWZe+aI+R/OZsNdC
MIs8p3BUaFVhbeNZRqIlpA5AG+7mu018t1cmrO+0/MLNDfuYwTfMxjzagZvkeglC
p7e86P0oJNh+GZIp2t3SySdFJmeptNoLMJxEVHweH3+63Tmu3n02VOU/CHVDC1JM
zkc4Zl3OQekflp+XwJuFCMSIQIDizqQ9keUWKjC8XYxByel6xs8lhqO9wdKHa2SR
2idZFV5XYwCZ+W5Au8N67Lh5e0GeoUZDsNSBlFZOez5B972UA912MJTS07O8zmid
StH7wZNkxrSnfMuGFg/+q0ZwYJh3vVnfr8R7GfYs+ctWAB/ByZdJnj/p0jW0kvY8
117xLF3/GVpKSIaPPXh4rbZcp0Vdk02/O1ZrplIG4+AuWcKgxXQhtxceS2YGXdyt
XQlqfp/zzBfQS4Bg4RYxaYk2Y1K52+hl3OETMmCACwrltYv7tKgHms1zgFT6N+/H
8xAyLMiMoEEeM7DpaqIqgijiJIYdBivKwvHx2d7YP2gGODgEldCysYk6Bj6BU3QT
NJUjpuLZ0CxwyETCuLqCS2ZcprF48ysxgXjCVIyyjOJo7Hlod8tElpz5mJGiVRJj
RkxhaYbSfIvXskaCyWB2T9iZmo6rpQDGcOyu9pVUeVTnog4Ectkyn1PgcajqFwzE
jrzV9/4GwtBRR1T+ZMFAo+ABRNv5oklxrnpKbx3pGo/A9HjaVEPCL9Hzrmjn38qn
LxRP6MuLu38Hws/pkPNsD8hRzu0upHHePP8HieujUZOQErN/cMFppYYjXbABYf/M
jOP7IDF4cfBIYnAoU0tIuYtemC1EIVoHa6SZdjc7RYP2rjSSmYCTG9KKxsr3nBkC
r/8WHJ+nDm4g/kJHUrJYMML43SE4fWKbYrgSSxC32KAXG2s7Ym0Vc4yHK11bGmyz
KJjg65w2f+RMWeIXM8/o7zIOYqaGqxhSdXhSklgvur+o6J4thihlkET2zYzVFFgR
UObm3FKzb0LCveQRCHEhMQgJc7yaSRFIQ/C8MO6Ge9Imol/Y0ZIWpEb6Vtjs2seJ
JYPx7ZSSOLbVBkrrvqVSjOJZp7PyQwglDYy9Z4QdKB/qalRkCNuPpRGjydfbZAcv
CAbcb5SsJ9OjxVhP1xH9E2gmspjzVMF+A1Y8Z8twGQxtiRAcilgxLWEP4ym7iPHb
g5k79CYWs45E0l0d80k44v02nAnzjC+j18bv7TUd6SRrVl48oUTMUVttGsNyuI0k
6IREEgGV10iJRBwvwBocZAXeUzM0m9MKo0EXtYHW2kdM8tmg3d6I7nlI3jLH/Ue3
2Q3yDe0tdoe6GYWMVSmkljZzZ3HRM31cMpQtumHihegarqYhGABSIiurdTDt3eav
X76PXd02dqDqE5mnE1nnFdJxMdjH5XxCfdJ6LhezDi4=
`protect END_PROTECTED
