`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQCMeoPrvnzZPPpU/t0uc7rYOufgxT3DlaOOkvCqHxN06sZ8fKAFytT63lM57I+X
FOYDhosXfQcgf68qNmzEfz178PFgEO9OgtGa9LkENeGC8oYBopvrN+VkGg1n/Mn9
rBJP1RW9xqm6M0KcUxkUYpVGdg9CkVjLuGcgWyiE7XvlR4Yr1wm520D0QVaI7Nbd
KsEMp3NCF4C9QaB035fV62yNefC3AfztekDJKAjP5zZNTkqH4kcKWTP6A9O+iJbt
MI7VWhkKXsquo+61D1OYsUgADnKEHzhJarRjcPPBVBMyQZWlkZnCrMbt8f51JYe4
UDLWoFg27SP45lwStJ9AGye/Bg9DlY58olDDaW1ieT4NtGOQOzKBxceV8q6b6Dqf
0beV3N0/yPHpkayled3wdsXa5v6TChDz2OA2Fm4EqFCIbbEnlv/VtkZ/i/9gMAmF
gVhWvyucmpAO19aD/4SkqSE2gYxu1IiyZpAk1nZBMhuyKItbh9sqETVQVCx4VysT
ZNhhHx7NEtgKJPmVbJaDAjJO89zgbdk4ipMYBvzqiB+gjKRotq5ImnKG6zEsTLQs
3zO6oWjDdi89D7qCUipwzIe7xNrdDWT/2uwywSmz8obxzYhxqe56ZOrqWGaRuNLi
cffDGP67oJyCQqVrv2c8PBbtobdmX5oLd3Tos/9EA1U5rFIdli99KTL3C8l11Tbw
lc+vNQ1ytsKV7E3B4cHoJWFhWkzOU5xjZbneQ/57I32IqW8UO0HsGshDPsJWlN2W
l+WrGCrQBgTFQ41DY9+I07XXOUVbcSVeUxjJ0+A6jwqfoe2skiGUEsYXLNuZgc7z
5BW06J19tQeYbTzv2O4VtxT9FXlft/QPCe81AngvoZ9OZwb/PjtAjphgD+JcmD3i
MnaYYdOfXiszz/QiOTDWwvcENpb7kJ/FerHMy6dXHMazNARCXMCEelttYSEml3Yd
pMVbIkIPrxKWyRVmMH1GFqabY8ji8UZsV2g6jGGL4SZneJQPF8RMaWTGqhuBRsOU
CQag3qMnqYCKE7XBdX3sMQFM2b8vO79hrHDhNMxRQnJCCVEQrvbLu0ZhpYpNSiYw
YsyLDZu41PwSuFWPa9Tm9+6dBwJ1uqwTRngEZHNbk+utOXuIh5CDdrtlJJxbxmHU
q3TUIkEHXZ86yTVSEK3YDYiUjJrTIQj+knyuTNKmfDxAfGc6yfGwlwiNuu8M068C
BM68qdFXzlwvqHjPEy6b/hbbut9ZANFmce12kyVkW69C9zL68OpzqLlUaaUDWYs5
t/lf8ACyGurtHis37VibWo3fQnzEJUMkzig5ymB2QvZs9RHJIZrzpfKLVElfZEnk
kjFvi4Y7B3yO7ciLimCVAHsDBS9GqjJ79DiJ4xD7Birza989MvO1nmt2LTvmEcse
TyAZLf32RmS3EjqHuQeIjaLLhS+n2wHl8pewtdzsQDJbdAo6nGvJTGrpRvFkQ+hL
Ut3scbNVQTpDzXBdyEDh2i9/jURxywZIaqMb43ox5R8QctAIUPqtXhNbIXNEQmoQ
u/dG6yBS/op1DFo1Po9HpYP8waqhaUJ+3pyiQAdrZ0NnWUB810rRIfsVnBK3n83C
ovAgdv5upL4nbVxX5z8U2rFSbJAY6U2UVOmk6jiEKwyyol58nHhcntFmsGBKyqrf
k+5xFUxWlCh+HC0WGQjpROb/EtYDz/cyxnE0E7Ya/kGsNXwVGaP/bTXHsjR1k4D2
NLkldciBnnFX9nxoH2TuNp+fd5f98e2ux1gtd/fiv5lyrnvveeFw9nA/0LbcgauB
48g7n56LwSIW8hgpMWzc4ecsS9zPDWumHplELYHgT0kietyBajfZSQoN1B2vk/9C
JjFcesdHO8WhpaIddC4zMVQmfKBNKcZ8JvetXWUaHX0UDazW12dJi7ipdSbWzevh
7jh3JaRashE5nxJHMq2K2yU36Pdsqm3kwzIvz7VC4BDRpr7UsDn/MF60pRKLDl9/
TLC2bdFmNFt1NLdVz8bTRg156sRe7kDqZ7/fGDCgfyoymy0msMsZQ0sJj0euivNy
3t/9XgyhaaUZR25V4vL7f2OjolrjnKCVFSmO4DsupHlZKyitNo5jA2Pi9i3AVhon
Z5yuKiJGQILe1E6kydiwSDKqfjihDKddsROUxb+F1aJuK4nGrqhkpyCPhECt4PWY
o/uxZPBmfmBBpu20/ZXKkUCWTI51GwQ82VYLgL9AEqo=
`protect END_PROTECTED
