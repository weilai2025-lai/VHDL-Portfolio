`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZRFJvDLffdrA4tKBSWJFd16XfQfSvaMWatc2TlM7VjwhhY5Zfv7WYqVzDe8yNGx
VEmUK9Go9uhyXiiex+kH1IJZiK6idQqUEx4hn0GYGNoJvSAtoabJjUipvqxQgTIl
mMUfueOtTXmC6Xh7tV4jOSbVqw0pR712wooN3t/VtvpFtmi1IenebJwskEWMl26I
xmGiMakKd3jiE946gaiDUN10w07ph7KUfbgLyxlS890MpmGIQwRJsd828AXAk7oU
JDq3vIKSnaqYh6MxmUZJRwGH4a8YWmLDwYfi7rzJEzqOH/tlY4jDFoOxKKJdqiHM
CsBCqXK10HIgxcHYzHpPXxSOI3uG2ApjsidHKcTe7g7yk7r1PTkD2c3DxxnXqbaJ
Ip6S1c9yI18LwwBiJvJm+GSshAnT73n5sUN07aYICJS0ova1MxueF3FZO77XFFvj
q4s4ubokVAX07L6gprG5rK6lH7QlaaATGYinC3osjLu0tJhFkesT2Yqid6oev50H
f1pJ+p8hhBu7n6C+S+zTwNRk0pSVQAGpa35VfM+11qoYMdkTny1e7CnoGi/ZKW3w
o91HtwCKGuhuydNHgwCaV+ngGjzXWCdEP3Ns9iUacIpzkI+pyzBW0Edp0JCw7AXP
B/TzmrCAWy4mHaqmBJn1sF5jTR/X6D43AvFVYS/LFc9B+s6QWOWSl4Jghm+fZr0E
WzQjU4EZKlwx7AlgPMeo4NKpwugOWDdWDCYQyduH/abtohM892lcRfd2WLNQ0bqV
nMfR6gzJsRmLUTVJf4F0KsQ4wD7GyPEwz1zxOMX4KY6Sn+bRzhbB39FAiXj41EqO
jnbwMjyuLYSGwlvFZgycQfb4TAvxJ77oHVRvDhhZvgXE/qz++JkxrBRa691HhKqf
DiLVpevpI80N5M0NMYm/EpEVgACJog4WHhkokCspmxxjiUxsHWjytg/sIDf9a838
BTxDKdFcfkPxhjBHkPCcBABjCLZR2shH/jdx0muV8YVuIAmjU6WreGY+keI5PBnA
V+qinJ2l9+RPYECOACjHroHiHrElbndShXlH8UJ0Uz2G7YH/NCJAxTgqZ6/ACq72
VQV9woKg2NMfX00RUgKbHI7554XXK+rXtfQXKbSv43DQAwZtn6Ylg2YG0BXsQ8iz
U5bepG0i6RukJScxbkzoiOno/v+DWxpKi1HzxAB7jmnYk1psRlKiIl27cZMBYz6o
VDzg3c1cZJBMORGVUPeTSDT/Sos5cW49P2YVTDboSCHFIDSO74syMQtleA6mcZzb
WalKSC3s65GrWA6fPmRV7UyEW/SBwpe929tv6NJPpYYd2ilQQkCCwqn9Urn+L+II
3N4Rb0K7WwjVWX8esfC03T+BG9djJGuS1eyyDZiljBV5unYB507LeC3Ie5AofzzH
AiRQq1bkGysF8AGjt3vKbEPVgGlAkdKIsihvWInbaCCSQiONopwzpenbKaHsZ18t
kYENidB2d1UxYPFZVxPcoVGJUM8DtOy0opg+1A2kaZdnFsVkHnDLkOYhGFC3yCKE
qcx/VFUL350wdm+/lTTbzOnK5pA82UvoEKpTTz039zIMa3T04OCl3lwrEMNne71m
l5QBbTlQVs000oX1Nrxt+mlvi72bVhBUXP12C0FIfCMg4XFVfN7weF5/7jXhlySQ
jUuit9zwb25KKRRTKFJbf/L1fHZw3I3ofsoKEUfIHhdcaZtvSh4NjcFVyBe+fLal
q7H9mXXrP/fs2Ide5XfBebdKqniaOc6SqKrGJsH/wXlAWOfsO1Dl5JxvDU8/GE0M
P7Lx4TwwGZjJdkgb17wffSThJOyQHb9uup1t0iUNqDFXt0fxKBvF71ydUt7T+aWB
Xqu5b3eVhXEYNDQa6pbDngt57S5bRgZ9l0cusg4NN81p8HJNGGn8k2OH7/H5YuCS
IVid36U8N1Wx2vlBpsD6dg==
`protect END_PROTECTED
