`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CViodQ0AS0GmEnlbTQmSKu+I62eUBneBxzkr5D/Bdbn9SFSBXy1jzJtvVyqRXAL
1TnPjn0vd6l7wCKuWZ+nWgs83ypjHHRsZ9ctYdWSYb4getHlozKfN51SLINHX2G7
7NnWd7oW7RIBHGxoUs+GQtJUmDhaMVMPgl2qQV7J5B3zxn6bydUOFTIUq0mJ1kmD
g7afNib3DsAlVo4PPorpNyTwzyVT5X4y0Kx+lGI+BCwgxonJ8jzaKcs3yuJlWLCU
bZXDqEZsti8bTFaszlxA94tWwvUGgJfpsWglohAo23zmcJG4wvvlm6xX3o5FyrVk
nE8ulcsGpEfq6SMjp+9lL9v9AdHRgLZLpJJyLVtpF/Xo/wArgeCPgQ2PSu+P9Moz
uPLyGvW9nmsBEBhb/0xvS6gHiLKTU5whr5jquPqZnqdAIqOJhuY+EhLPUwqwN026
3BHvokwrtf+xSBa3H6G6PAT7LUH2yTHMPR1igE3ujfWE0hmtQRPIXXg5b2ipYH5m
xKuEbHGDkg0MLyN2MaJKGjlN5i9mudyCIPKBmIhXBqBD+6MccQlIllkTwedOoMH4
moffdHr3stOR3DGgQ251QkzgolEo8JifLE6EY80heW1do/eV4BCdZcvg0z1YvvXy
2ioptO6ivSYOlaET6bRiSdSG+WCT6eUA2MZggMKx4l+Q1hN2yYnxSY9GnsZD7qcb
Cn9WIfslFpo+PKrKyHy90GyLcXT/wNrBiM8wZm0Qytac+Pnjy49C8LXcZgsua9/a
78A5jMbU2dYau+nOfd5BX1WK1tVKyEGUIQsfj9V30CYaHu24mBSgYwwEkuPxbWiF
FKEBuHXej5VM6FfBeUiMEB3syp+F6eCtvKEvp1/aCljgUJu9tEkPiEK4Hun6ifBT
sAkke9hipMzBnZOJqSgNHCbeonQcXP+/FKFjbv8YsGssIKrB1063sgmkMHnhSKnH
7MP+jq3qkkbywdfMQSzt5UyM8TUlVb2UcyMXBX6vMj+zCVVQoTG0fnqTv4WkyOqo
GIW2R2sfT7gWnGog3SCUcD7PV5lPN4mHFlNiGQWHvzm1lmF2fFxby+j3rLXJlKEo
mebKVbWYUsGyjMGyfOzzHro2eT6fD55hIq+qTvBOi7xcmqnRlGwZS2mUhEtzAcQE
5OxL5oByDTuQrsKe6dwfhTv09OTmLMkiFBTDdFAWQqPjdUxxg1R55zQuvTujk49H
XM49V2BbtnSShG+6UWbjS760f0o6N214TxhrqDW98eccqhuAEq5nORAPXRYdI75n
31O+BdJC13O1EEexXY0k+6i1C1JZ0IE8OGwVUHc1Ac3MhcYNlNPm9rEEYCZg5Rlt
5dCD0ChiOSgYkqMZ828bq1OY1FIb9/y1ij20sirkL4mMclPLMK3HVC/TysmGhV6X
kvigHDqBDxm3tkvz/kjLKP/60gsHsaIvwSOL2/wQ4uNJJ11hIDbz5HNvtb6DxCBV
YDj/X8L34NRwvp/KX7GR/Jqv7vx3A3S9hcoZuehn4Gp73vehQrldr9xQ34qxls9G
Tv1fNBUz3fV/M+3FJzO7duIiufG9JVRVfuiPVkXlmpRJSPGJf4grqNRYh7ul9xWf
Z4lBQQtOEsiD0jgBoNuRQAuk47rf8K36N/vXyr2MGfjUsJ9571dyxb98m6zIg+/8
msHIvvMxPw4s7lvMGg9wN0KYb2Bn8jIx9EoEs4UtqYmEo8It08rYYthGIVRv9Hyy
Cce68r+QijCqKju6W7bx4uM6Df3lWuljGYomeCgUeWaMy5Zp8T5F/0C8P39fRXcZ
1CmaVAUKjuU/kg91V8S8EKwy5++Au8Q1DAlV/dS3JTEm7cCX3F8oxOfQ58shmof4
aciCN34UEKUSaJS2B540/Vpyl/wmm5wUE7lEMskgb3+KI8RbrIt58Q3NwwlUDNF5
hOcnlKYEWdEfp5T5qI5s+1PPj7BFjhusw7ZcwAqEzzWy5Vv7tOS8xHEs7i68Z2u5
AQGuD0EQ2QwUASseE/aFbQOqis+yDGSUlILOsIkkO3UWnT3my+Lz9zXLQfhQRljP
S6fqjhmlBf9ofdu4YMp2JJOfHdGbqsFY7fZZifSIyS5RzkBl3uLSsD39e4+HeV5j
dJuP8MlLKfFWkynpbbOjhZM0dobO/lc63+UI9Ent/oHR/n2ouEsG2gJv+duFT7Ag
467vrAFJespt1xK6ZM5iaCfltDwletVZBQK/OMrsxgwxJ4/QSRe5dnWozj5XqZrV
Liu+u5rJvEuKW/YsQSDgeKtrp7zm90MX0AlegUr6i5YAjU6/kltQPzay2qRmsOTV
udS58gtL1RldQKYj2+093A==
`protect END_PROTECTED
