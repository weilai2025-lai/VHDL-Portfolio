`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvObYUTurJ4c2VjC9CHdHsiEwUAiWe/aT2Nl+s19ePd3EMWQmoESPouXbXeBxn1I
iNxrI77gZ5id9Ig/RQ6Jyu0+SfxCCdev1RuevYoCZyi4XSDXnzBAa/fhoWqub0yi
5jHIIRHI1IgDYknDJonpI4OLnroZq6ZsfgoPMaK2YoG7LkoVs1JvWFH0mdCrzveP
mYcaior9/cRofFd7Uvd5EuHTBw8CeQYDcz5rIsR6U97Ss64APIBP5ICgjC83xrhJ
W1bcRLCe3erhUsPbsPArf/QEGplGnafKSfzfreenfBT1bImy/HGQ4XWf4AvxXvqB
jN1nrYHU/Akx1F1VLRaTtmQqZkYYPLa09BpYq70NpPry/KeDjsmwUbfw8ObkR64x
PTFsE4RGnibHs4Zr9hmhYxz5D6U+cqpFniz9ZLur2er9aHl0w/cdl3NI9A4E0sK6
QfETYvx/3zCoSqPfCnoACPvJxbSBFUZUMT5z/jwUFwgeVGmjQ3vLauFJlfYL+ohd
1qtWR67peMcP0kAPv9U0+mjUNc0IL53fHcvXbFmmRWiz0/m3j1i6Q1EdMFLQArzA
8QuX9B7rM9kACPRDpshpeAowI00EIPx/z0vXqea0WZAH+VwDlQtxBjxPGnZN/lL3
DpviEKUHYanE59oSsSJB9AW7IZETN9wZ40xso/MShYttsuus/Ab7oqFaRDRiayUn
otx68aUsb5XvbnnBzSXxpOMPIhatHebZC88O1W2IdxKfD9K1dxfN8uL7YRcg0JM5
46Zwmny/HCkOW7uBECy65vMHT5oQGOm2p45ZZwYbgqjZnz32LwSCeseYlUEX4Uor
0JL3so1MoinlC4KUBFhS8u+s23DmUL1+Er2UzEc2OULSEIyFEaUvtyBwwAxYpfwm
Xc1o9FH579AKzaEcQMzfXMQYNJo7XHYXOpU+Bp/gh/ztAVT87tPlJ2gcTHXi1+UD
F/Ld6gccAuys2xvjnYa7tgsUEH+xZCCOd2h/j9LmpQOCQuLiY2H5uXzqq99zDXX+
+d/BLgNqVVkQec8Tm/P7zTMwZ3BO3uDUfkSAQXTBlxdZIofIa2u0CrW+MKSoXmca
Hi1K2NlgS9/Umgjhs2BE/Iswf6rkpJIViVvrW53+Xqw/UoDpcjk3lIc8wgtK1acp
jQyzy6XExHglOCtcP6pZXYDz3wx/rdWzKJeGUKGD49DWJ90brxKvrgmv8uWomgEe
/SW50+Aw2GSOfZE3C+Nm6w==
`protect END_PROTECTED
