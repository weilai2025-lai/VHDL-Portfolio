`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WCD48D0IR/XDRvcwGNfVTR/SocDs0xIZb8E5ESmA3L2XwgU7pcFY/f9FCStNenu
3ngF5wa1QjK/Z9pBPCdH6mo+8r76q/ok8nZh5MAJjiHPwXfGkjgRvXoN/arjaVO9
0lIJB+EbbL+v2XTcke6uYV+XbGpek7RRTK+7XMQwKCGCjtzsJWIu+3bVv3ULQjPf
kGA02lMQAydswDnu7kH4mj5JgCaHokwBVcFafO4IJSQHqRYP8PUhkznJIhBbkQuZ
KOiIjW4vbO7/SP1w7yKtUjTR2za1raS3kV7bGJB17rPGCVL9G5PDg9mt+/kIb+ri
mBhQ582+qfwt/WMYYxLyuzIQF4l5S/Eexnx8N7UfOgz+OQqJkX4kqwHvbN/lwscX
Gb/kRn4Hc4HZ3TWAtxl9UeDFj24XkMx5kZdZzRThqxpWhobPjP5RBZUfGJYFP1al
RmbNExZKMbLj1LfUatcoI7xe6plRXvPcBvpZ9BRnuwzvbMyBiE2w5e4Qi5FrYHgH
1kToQOEY2K6NEgFy8a0i7q8jOTDI+ioU1TnB1RKCnyLbn0zcYA77i3Isgg8ywaqU
JW5HvoTWDIQuKhN4HWZiqWv4VXZK9G1RWtobvsCBhKl3VA81fFRSZ/3W94j1R4yd
/GOA6Yss17V2VBw4hEUbkEfRmt77uJbbKFxYtwLEfDXSdWLWgFHNuzz4C+PNcSIu
PUveDGuqv/LSvWt2RsYdORbu5PDO7dypCFP6kxEqUhy6mn+9oRX8nAtkBszxkHTw
IuiSt2wU63d0WnZbZq3u5CgqRM6+J0kAYuXEgaxmMIkgVSv2xAN6W926XsKW/G5G
iUL5Rz0SHo5dIqSIFQPj4kSJ98eLCwyKG+sk3W7wRBuJ8sxRGlFjmq9nMySnpNkS
LiHuL7KNktqmnZ1XTUGbkfGjPg7pRIhR9cgQgpuDUVIwUDIZTsEqZBdKu3Iv/iMK
qlyW8cqtzZk+88pna/ZUVhwOU4/E3n8DBXcsb/Kds30ePnv3V+KHG+1P3ObEmdbf
gVdFCiaOWvv0coaRzKxxKl5CxaYdHpfoeIf8SILw6f3j3K3YWqiuEU0l6GfzKXWR
/C/QVD+e1Rdi05ZQLQCtC2GoPRtA3u9SRTg75TPg14uSspkC+rTwHA4hnv8ivTqe
cJ9Cp2wk2MsOtWMAOIg0FAPYC5g+n3BzJZS8IVecMHffsN1D2oHf8AgvrEe3BcI1
k1pvbubFUYbK3rIeL7F1XtuLNr4XAxqFF9Yb2cBRD9ZpNaab7rsZ0YGTR9tkQZLw
iwWDWrJvn6Ilo1DpwE6RnwbOVp9gqzK7nl1vYKYDFJDtPO9j6e/13gqd/CNg1+O6
C6JlgqmafU56DW6JbXDkplpv+GJ6aL/bH9bj88twjXHHrJ7HyX1oIRF5AescNGBw
xHPQTQr3uIE3yoMTLcKv1Kyxj1ad79sjPdHbmehPGc7mshK0hs71gjt4EUVyhuRO
A+aaASQn1Vcbv1fk5pKy+Lh0Fag/bXZYu6SiEuQt48NqvWPSfOuLSbBOzlsYdxkq
OfxeNIZ8hw1oMfpan0e5DP5HrlJKKtMZ6IN6XQJ1zDZIt5TgAvmK/y3qs7OYCWqC
1j3FGQJE5aXavok6x7v+ZXSolJFeqG9E2YdsErplhgqxRnJNGRgwHcFkAAdHfus2
WiX004Ndf1GefB9Bb+xjYFs09e7hERIpwdVS7g+Cw/i9sR8hS29kEYWIJqeHhd8s
KbS+B6a1B1r6rzbbAxw0/vDRKwNePqjly+37RQQA64knUrztHXY2gid4+hzmv/vi
tK4M4p2ztmt0l/QxXcSe233AYN9EUNXO68YOyl6L1NvaTOBZLq+QRgM5FEBENHsW
eRucLpKEwZiW2Kj/nbrpo3ocVGvsTyzaVv0PyuVx2EyAUgYZSit2gP2cNaQGDahv
0ZLq7nDMHd7UJJmN+t9/Cvq278a0vXmTzpoElZnhvbAWyMVBAxkthupqoal7R9O8
e+HlhPvzaYMI0+VQYmJRoIhKb70aXZ5WefJHvDbWWHB3vZTW79mYeTQOq2KcMl/t
`protect END_PROTECTED
