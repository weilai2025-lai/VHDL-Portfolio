`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8eMUCijGTSAWwfF+OieTTTsQMMvF0WPe3RDYLV7RpeEIkO9QgM7ig+X8wb6MrFZ
62TrTsuH3Na+NvrTG/f7mk8JulE9NSXmwB4TnHs5of4QSIfaQ3Zu0MtyLwtktRig
ZiNHd5vR3rr6x0cG9oSJ6Z1X7czVhDvcsk+zdJBxcVDroywXO7luFJ09qfp7+gE5
g7M0nRW8CZoPqFGsShSooAoRRbZb3dqE1UG/1GwagdW/W1JjZ6SSdH8CROCix+L3
+0LGRRmBFOnV6tblzc/CthVsrSXoA7SF+NCITIDOME9FBmFZb+r2k6YgyrL/ozJe
EpjzYxLW8LJl14fuh7XgxAvFu51yXdDech/B8XywOYS0bhqerbZL5aoxnMSryC4D
NNgnWt0C3TzFqGp8lopwnBHvd1mPQbHo8jV8+8HMIMxxmjm1Qu3s8xJSOpZoKzMa
dB8NXR4uHmD9t5HBTF/xGuj54kRvRJYhaXBmY3PV9MH++Mo0/CTV4zUx5kl2opZV
QvAwZuvyUrqevSDfbpXo0kNxsFraxpczyMm19VQUCA1pY3qJHKpgTu2eV0PJUmwn
4yb9G2lpP6icwuv+ZP3CSSyGi/kGdSO4eMr5Kpw1uvPWRFCdhhBRCiR44Exhs6Tj
lCSYqeY92jTqsYDHAZW4VHfnz/CqgMn/RLEv/dqDnFwIkRGOJSgOTs4xR0BWbs21
o+D3DYmzTvbvPkDcbx/4oWUKppTkfGqU4KeKaYawcsv3rKhhvPP6FuTR3W6kb3W7
0a57HsF3gz5R6RFMQxPboKlPjFbMLq7lPQWVNLraMCoJT+GnZMK8ThS/ulH9Zq6D
azha3jB6HCSr5LakdiCZuKlMVy5taTS5Q24p+SsJyasxtfa3QmzTfNdNR1KhvXCY
70Kcjrrob6l+c1HuU2Yku/bv9K3iT4s8GJPnqbvX3QJo8PShXTReakRqQFx8lKBW
vpgbrroTPHhnyG+VqsQDFhux3xi/w9PecLQRUSFqSkDS63IHN3g7KoCpFaGIAfzr
bEENx8NWd4cR/Hp8pLw+cQFfyql35bO2i3c2pV3bUYda7PCvLQvPyk2Rwe4lL8RI
rBgECkUWMn3l17kEYWN2PnBbhZ5eHYoULyh3I3YILM0d3Vhdp5i+bwE4HHMKOqAT
SjAnAEkjdahho384K1RNm1FBYaqNn5sJ49Yg4lcwfZdRd+VAGdPOzNB19XTqc2p3
cBaOjQxC3SSvdsxvYdZlWY2En/k3NRxjMTZaD9afXIuKSKxcE8k0zHNZvYQ3EPEt
OECpnN7dlBUTTbbdgKYtHD31/qn3mR331qmBwPRHLcqCxvKZgSEYXkKwgegktjl2
afFWBNzfl6Gg2H6VJf7ELJpEhF2f2zjbCZyPWJyOiX8AP1liIjEaNg89h8D6HIts
B0HXhNULOFxYANsIFqNwgRpwIEujkS6MmiaFYgaaU9CMRQLZabLmPY/9ASONIujV
fs+ufl+ohGjDLurweTdP5FBRqDrlC97mTv9OaKC2xLrFYzZ3438qe8vl2A3QqGxf
e8j9hxRQQxIklDX9DaaOAgELgojPjX7J4Rf9VciuRBvsFDCOckY+KVzcw37N+cnN
JrOpQ2vM2730ODPynjPBwchYhX6I6ugbsGzdUbtT3vGei7bXqxUzbyBHZcS/o5Tt
ri91WYFTNNKoKTD5k0qiOftINUw6JLCNj7rNKvm9aF12/tJUjTEyW6lW/u1loYm8
XIY7nOCMMsK/s4SOM6D5mqaxht1lttbBoD9mmu2kZvMJeb3L7vpp0tT4iADvHZTC
45IOEJweGlhyvdDlfnw8IZP6m4q1JLw2WAdiP9d0PX7uUsF26gauphQyONEKJSk1
BklnhUbD2kbpFxPP0tCsBsjy/SMFOcy0V1yfaW1yfmeSLbY1ibsPjnZaBzewc2Vo
ELRoXAQyiZxWE5DyZw518Ek9R/eYyfsXwxl0NwBBlexowerQfUSw06lWQprrjRhk
VNTevUsHHKk8cldQinlFxxkeJMbc8ET2v8QwVGbBU9/2PxW7bjzlMxgfPWsVt6kv
bXfu/cmNIGllOUFslX6DGpp5qIKjHPmGzjg/aG0EH3pDF+CAFk/seW1MMHMgBVUD
2kCNl619K1vnTv7z6kELmGio5tGZ1ejc6ceZY8RHaP7zWf5oVeNRhwbjCkJyCHfv
SNHKao0UTvD2/FK9W/ZyXhKYWKaoS2N0Mpzu1yikPKd+JMBqYw2C7mHtIS/auDg1
wvSlunINtH+CfAWVeqChl7PUpwwnAjuz1OYVieAngd3MMwPkUXPJJw0P+dZIn6Mo
5UQmgpH+v2DQBOeWqKrsApOs8/TL3YjgZh7GbRwKuhD4g3sHZICQN0cfhjN0q/zd
d0V7RheLOdQJDLVg4zw3+LV5CuRbSONBYvNe42Y9+3nQCYgRzQiwoZlkvUN9v9AT
DFlFMxzj4FOK8UbNQi2JzR+45iZ7Jegkf+3dvX46pXR4VR4z8e97e9bobvRKQWU3
uIV2VvKM9D3ud0fig8WgryxdwPJcOobz1+vr5bdUayhfwudB7q4ntZipU9QdMj4V
qXvnByxQulCg6SDG58se9eghH8dZPKsZ35jg8eEpubFXkTH0L5psq3EI6oiMDZUO
5U7wMcMi9onP72gk7qz9N4r4in8/d4waUkeyJpLSs0DqX1ltrF0cXULksOQd81V4
t4F4+gdeKxbh4AJsGFscP54DjjZm2mLCA7ncM0wo38ho+9eKkhL7UGhVu73KwHtQ
pua5yi9Apn7op7nkbhHs+F0zRbIRvwocqsWab0kaQU9P0tNO8/xKPFb6jKY2Xbhm
TY8/0088qR9IEhFf57j7e8OY94t3OMnTmmvbUSQTDX14tylxszPc1qozqHz0ou43
BTSEmw70e+X+E6GPDk8isFIaomDztgBnZdujNea9coCmkeYFtEkc+ADWZ5UREfxv
AY23Sa671wy4oNPEXAHi0m8QK9COB9XWsdrbuVBFL4Oh82bJlcpHu8EM5+sOK7zu
1QwrnCflOnz9nLkhQlMYQUOSOI64A33tKjXIZBFBT4TgcyXOVsBEmse8o6a4M9R1
0UA7tvHzfruviDC8imGfWSKb37DYc7/8x2Z3pvRXpvJ9Z8ZVytztHNkYvsXPGhI9
7amDCQIF0FT+CV7KO336bAHtrgq2yJhZyy4V2LSa6pSTk9hqY3JhjAgYlwPR7XCS
xjAtghDNPQT58Ye6tuSCEB6RgLh3EmulURYVs4iYfk+JocXWwCDygAEjmy4asXLK
6Vv7QqLGy8ywyf+A0GiA3dPD3kC0xghXTHkobdhYGm0X62aWvyp2n6RT/1KBJLcb
ADMKMtaMlrXiVOc04DJobm9rAhSO/NQ4XXRtfC3Q9U/b02h1Hmavjc1so7om0TIg
Bd9KbNCRSkUI18eh3vPeZdFj3oaim4/v6vlxEB1oC4v7eV0Mvoe4/32hFcoJHQs1
Qdg4bFTf3CQsHhjF3aSf1d9ZEtMQDQa4vK4FTFJemQO4mZeLdm410Sd8PCit4b0g
XLa3AePpzoA3tXlr6WsKNsJADo5Y0jNFlEvV3PjMgt/hDRY4/IQBe1UrAYP2Z0VR
ysTmqGFbvX2zhITvzV93KT71Tm4MjkSIur5cRmLO/YORI7HF4xVoa/7ZE/iEkDu3
VGzIRaLM/1gzp0gFKi67OArGBWcaGx7D9Wm2qlW2U+oP+Si0UHRCtTP/edv7t3FY
Mcm718LyUttlKUNAgAz4JJf1UDsXgst7aHkNFhdfNjPner5nCu6EHW1eH8fMEdgY
9sEbfokP5r7/F6O0m9h2QblCbiW5bMz8PNSDukEqSg03wXmoZcWypveZdxEzVo8u
lAoOTBs+QgoEqzgFUlFlc+IWnWwcpsh7DLAGJp+W7hXKvN5+iX5hZFZOWqQPFHy4
7ZGZWKT9xEyDptPlxlEFH2c++rs7E9ncgDM2XEaiFlsdz1ZTVjWGjPv9wftN5n3k
XZhwW81bChe9y93jwGzKbixH5n+joHuDQucRSenAfYTcZS3N1VhCCgC28EMyMXPe
a3S2IyLoOihsx+hNmeYv0XNuZbYVULPJ/VLgqymaAASTRDrgsgrZ2rsBX3h0qmkL
gaDIn9jiHgCumEL0FH701S/QxZ3HYs75BXeL0mEiWr+U5zDqrsL0tD9YWPbhQE0K
BtD8cS00tBU/O398Nwa60ENeQ06lJ3L3Ewsy4ygpsP33KJSJ8C90Jg9wZT0AY5mw
V/VaqUCCWdlHfJSfPdImis362aowKQbiu6zjL5Jpu7FQ1zxOg50oqZKBO/f0prA/
VsEvvnEHs9q0AF3PnvCEfQFt2m8Fi4apd4Subqr8FNaXu2odutnjqUMAED+e8RGv
2s6yjAc41459mGMsUqiF+/eEV506V8cquZOC9Oehnl83wywkF3Gr7aqpUhuUFOdv
CFNcN2ghs7CcaEuKeQBi3kxN/epR6xbH1CHxNDLKQaCxtbh5Fzn9TUXcVf+pcseL
Fpv4gcR+gGUhqs1ytJYMaX2gZeA+b+5JQBGYJcHYw3XdBK1Gk/1tEoVzNPL01Qsk
Wnbns9CqaZ8XReFiceQBE7B6AkbJwp0dXFYU338zITVwUdz72A/nR3MqcVKLaLTW
jBuPVJWPHOj8LYyxLm2DHDPxGqUWm/LS6WYMhOLP6Bz3xm7QvyYHRzeCRkLCgGCH
1u9RaF4S6JSANoap4xhz0tKfloUxdCHYJKYRUeLKgf8W6dHa4mRJ7sYOidEE6pl3
fI8se8TZ0dxkjA9bj4Zk58VEMpdendI/TTXIXQI8jvS8PMvMX5ZW+63u6XN3hLpt
vBlk13Aue2cWDb/HyJMWsOwj4v7LPldo56i8S9OvNtYwbsls0CC/V5QSB40fy35k
8MZmZWnHV/qkszUNeW2ecxIzed8AGUBzX3w1dL2am5tCuYWWtgjqwlmEo5sqtdlV
ccZXWkjh2Lhr16KPcA9zPB42FNJw503cm1dW9nCdxlRiGFquGA7GSpitRl6Yquro
q4feLP106mruGvNZGACV/tiFqyKqfHWRrQKv62Gq+gBNQ/ro4mOzf1JPepUaLE3e
6df9lKCN38lh2g9EWfxCKUsyBIawRE3JAKDHStG8oYFLMVswvwRqx3W+pgV8wgYi
M9ZEo/921VXSJkPAJJulleeVjpm3bgQso6pE7dujFjorSVMNPQMP9REAjRJVGiU1
b/j99lQ2bsTZRKhEtQGy2/7yXjKB5p4skfDb498RVllrcPxgL4UayD+RBWfL2Efe
ImcC7hWrS0aAd9ZMZFTFqRDGOvu5MBl9ZzCsM50eEIWmL9kKbzvD3LVg/7o5o+GE
6gAq5I1QxCj10J6UKzlvR7zw12rwdhzAn+sDve2vj+vPx5+baa2z8yNXb2K+xgig
Opb9uH9+RCyalLyleilcjmdpALFnD1lxPf9Uk1YkNfdlrsySNasM/AyqzpJ+W/pG
Qq1JM+nYO4yAjoS9WWutTf8FPdHMjTvorqEWUlS0GrfPgS2aIWwk1b9yToYwiTIs
Wp0eFDvWBCHRrVJ3zOncDGfKM3v/vM3qSW5NZlG2DnwqkLlFigw27lC4pa6H9CE3
NkhR/z8+xx4krCh38el1eMMfMc+R9diZ/VoCX6df2JCECWNxbnoUAgewhNNK3GRr
H/D2ErxiO1bfnpOs80qQ+IwZ3R94LIejpIp5bjXHV3aMpH4SYM6lXKjUP2MMXOrF
US4hLgmSbD2U6Ng0JzHTRuBzm0WlPUOMQ+uYD/N2KbFsDv1IOqS8B7aguWZ9qxAd
dJaMjGRGRBDmiLZ6Bdy3HVDhOErhouiERRwALipUufCUNomvAUNVlO1oSAxTmfVQ
9KqPMEnpp33MWETHecUikh4yN4INZFDHCBRwYzRuOZZzo12TO4HKqWlYNf5hgMOS
J2btef7+keH15myLZcoXf0SGiKFInq+eeZ8I/bluMgPRVsRX8eVYPU7bsUCaMF4y
mF1ATRVJMhUVEHvQnzVBU76P9Pt4riYDvG6NphX4hoLES60OsOwbYbvalGwUuavU
M/rmz+0XhbzFZYxpEEKV0RHkL7QEeuYxPzFZTCD7IxoMvwqmriuixhknepYFUqdA
ODkRDB3z2Q4eQ2oly9mvC2fLlPvget2OaSYJhmuELCq1DCTCK+WvTSJVJQVxAwIc
tP8LVdWPK7GYZb9QN2FFcgjRYvzkcttSu0ZxKSIA6YxJ6OewVSNUJMnE8kfVAIIf
42jVOTSTc/Rs401kyY3BvmYJS3Oc4pmg1GFnPahBzBgPqwnL5NGDBtPOsV8FGoD7
xPRNHFCd61xwkJ0i3UAMvRbWcxd856zqi4YpDUlkta+WQJQr/IfUz7YUEtQHgdDh
XY+e8Ih1Zts2XI7inpK+WIwoSq4FpiMfC9ImXCrSfUO6PY2fFvC5n+WV7Q58He8/
uolAZ2Aqgx/+NcsfUzcT3SvjcelLLsN4ynWsVLeHxThWZ4V04IQkLbdPAUL0L9Cu
gsmc10gI8gdOaMc/COsI+/TTEaLWW7snn0AzhA5UtGb7JCSDo8/IPm5xLVpkBtRs
cRHKc6G/K13c+rv99aqum97lpEa0LfvOrAcIl5AbMIXwbeXM0yn/yvbfFxkUds5b
YTmfIFyBgRVku+iv4nU6qfs4+/vO+Uruwj0mvzg9nPSwn68N18BL2JotytiWvLHX
ZMShVtXfWmKGnpBF7SxejOFadGKrA/UWvHbQ0BUeVhGBvwdlCekJN/qOK6WIAAiT
BO4ps+4RwxJcN68orG42AiEWwq/+WU0eFITb/VAzFAXWL8rHRsBx105wnuA1K9Tx
hSEzJObzlo6b7+bU0ySKMcEdn+B/q1ZarUzsAsXsWHAegTVjplBLvl2hap5lms86
X4Oi9tU1OiVFeP3LyOhJjzoSW23VGz1Rve3tDljVYJWC9YaGhEbggau3IF55XFYK
jvnvajXwPZPckxPv2+zj0eIAuu4AP3wMkKeWDTb6mfBuX2AXIXmqWt/Gkzat7eh/
4aqnZEFANeY/JUjYUxLg6lzu2D8pkWEmHCJ/YxmR8efhTxJj6K5tt0fVPk6b8HS/
i8OJmXoMDDgxe8aAAAnzRCt4Hx3cQPLSAK86drfIx0xtUl/p+PFVwNJ7hjvEPbgu
cVRkUMwFBvBazSuTQpVdQ5q6eXb/OYSxDLvztmlSmX8jAdZZ8498s/VcLl5wEqhs
nrRRYVvEm81NNNsqf1ok6SHLQI1F1u//7vyFIdlBceWG383EFU5CFg/jboGoVd64
sGbgpqi3L4/5GGjy4Kr7ez9HC0q1/DZWEfWsdb06H8lgIkKskaZbOKDDOyBH0RB6
aAGFGICig5bdOCBDskL0h2JLW9zHH2YWhHtSoKloeo62fi9hwpIb9XYZpdmjLRiV
wG6NX86X1AaY5kgGRKy2FycfREBEZvknXnrVjn+DAdaCj8740KoB5q971Ki8NaJK
ihrob50+fxy5XdvFMJQvrl/4Ye0Q1/QN4HuiCZKDKTuarQZwtyeuMuatWRAbgeJp
RPPv1uafczGZgEB7BCPRgfptHj3GQJ57g4WeUQg5EEWmiFoGJuw7J2bY/5WW3aQS
pmHNzrV8BX9WacAOM1pgcwMP77uXutyxmv5/JoCnx5vFAFZ0HLbDTTWXik8Tdg7f
wRjvxYBf49DKCKJaZSwAQaP2UzXmcO4AcgVGFVsXqRkLbrKzm8Tu9pzePIf4QAOO
krqvBZciPnxMeeaTwM4YVuuHEGsHXcNOkldmHbbfGCGXM4DtKGEz28zxxFMp41uO
6wfSN7EgJF3yfAF9FbzHzcgAbQgrWh1IYWkAG8C1yUeMiHGyygTuPJBqv97U8fDd
v2h9n4n/qq8T9wDBeCb07Yd7BGEfJP3wOK1IYdVnVUBq7D3BtMkkJ51qKtHBOBJZ
t+Y4nCO68UcJ45z6vAg/yWDwZnCfXSSHENjn4jSyAAf9+Ct6isPLwTk5XFJeAyOQ
TQHGmNdVF7awVfLdxOHzH1JAM7lbeiebb4gPgD4g4MiYpyJQI3BVjTxbat8kqwFE
yfdc7avWZOlx+VAzRbLCdyK00HCOU96uS/FHknw1LacSXhE+KZguNPhVa+PbIcPF
Ma2FOBWTTQgAeBlrXNqBbO8AeC7mO047tP+nL87c5Ne/5kRP/jjAE//+TkApol8k
eM5qik6cbNJ6yEUto0QrxLKGZKv7akZX4mto1LWTDtY6gyEqgnlXSD1MhrbCktgy
7REFrsyYOQzpuhcrXFp7yge6FLODyHmOps9sctJcGrhdSFbdGPdmMQ3qLwhJr55L
O+RDSxzwvtGJz5UF9ixTjU5SBy0TKOr/m34cRgd4BYJiusOu7FyxuR7CqfFHvqPx
I6rOG8IDy0Arz/8x9nE+/U5xHkuWt8nMacg+CJw9JWnGju/3D585d34DecLRcour
4ZXHJWxAoA8mEPTV5ywLQZIbx+qUu85gTw7NIsFbkuoOsFkX3cYkZCxOUWRrp6cO
5QpCsGkc/l2rzBBt9hPLuNmg1FrD6oIHZYxv2q+2V17Ybowp9glMjvmBURGfYfaD
+FyyS4SsUgl3wNaKjBZt56ImOtDd0LbUgP5bns+E3kbZa1DPUyokJFIv16m/6deq
Tnpixra0NikvLgCYGBS1EtJlzv+5R/h8vx5a26Bjyr8V3H1rk1C8w6p4PagsXRQm
cKNK9Jfvg871IMOIvfQW7HqAtdFOk4VvveWLuTQXHuE+Y8JvKpdm5U7iOujzZcCY
kX9JGFCpFs35vu4DGxqdB4plOBLQpubEUVHaD+/kd8gMirvNwz7zxU89AjV0N83m
VDLI8ZUStJxMCCLTHHPy8Meey5hv5Jx125zdUy9QwCf6Y60aT5P1oa4pxO36/EQO
0SjGFP9yQPUQuIoWC0xSSmzm5fh8UjS4CFG/tMCNthuv6wDyOMvKzzVIryhgaDnr
8HKv8wqvpB0aN3LlMZMauDmamBxfZ59QmEsg8JFBlelJlx9Envn0aX+Lq2fZ8d1h
VWfPfWb6EeV8Ls+pr29Q0hady2tXSDra8wiw92s0BMkCCO5WOJYM583jd2HNDdJ5
t56Vg/xe/CXj9SynbVTa7JWxvAoe5gNyzZNjP0EmjHvhULbXeu3AyWeZHtxr1nY/
XlBA9NDnAmPvUET2WF5zZUnRrCfij+2DsRr7ccxcKcZTxEaKd22sc5TSIWhYiw98
aYN5ywhx/NaEZhxe/FBp0y3Sgw7Q6RVU8XwGvq1kietLEY54eCakgouQBEuRVqjB
hYKmHsjW5HWtLEKdlhnb8N8La3g4mfFuDJDh6G0i6KgBKBK+KMoMduXyORMV1zVN
L4A0YZMvM3IhBgHzxSFCJA5bhULbHKatggR7CPXRDyiLYI50smmVD+Qp9QiBLe1n
73TBCu1HsIPqbI8iUpg2NUS3o1O3hnw3F3TlkXZF+xOCeFn4tlVVjqa0B2K9w57I
MrxXlK+QRHd+CwMYjGuqbUpmUcJfEtzcuHFfdyTYcMv/pc8N1omMzDWy4T6s1ztq
W1mYheTuoxgK57HUaPNyGre/uPMYQMS/FEglFA4dXMfdAWHaCGCLnkq92VoIzg+w
KTlLs3Rru9lXnmGDGsdwAS1uYdpF1eyHKwViEMa+nwnkRZQFo9x1G8jebW0PDE8/
yiW1NoRh7uPVVoor4H1T2Vt88Ap0lzdlqaVh1x76x2fLds984WeDZ5LgOaI742pr
gJLbyK/3shevj4gmjJoE2LLIKdnnsNWrRrkKcuYeQ6lR4057/iJBzFiXeTsoDcFL
Vq8eHoRA4Pp3PGG0vFfK8oN8riNUAZjGiXLCX6EzSac/YCE1HCjK8S0ywycDipXJ
H/CNbjHrG645Z6iXYjH96OSo90jJgfQbfq9cPWzoWsmDNnRSVI9V6Qgi3OfpTbYs
ZgTj/vqlLKJmcx2+p/9cKMRDJfneoTA6KX41D9FilFpJhitmE+ipyeNybZIvkM3T
WFIDrnscwyM/GXuyx63IGSdakeDWtcUmF9vY4VzlYic1FReOeluoiXQEl/ukLIJD
skqvvenUk4C2oYQnfGwSRJtxwTiLENVB89w/bcAUbV5RPn/MQZ2asZ/aoPpU1+Ua
RC000RjN1zf6e4/YckWpOqce6lVys22NbuZ2aShO1X+OXLeClQgXlCCR1cxyFmUT
j/7FLuFEVRIqDDstxDFLw7DWPFzeutVDYGO81zQ+6gu6hNTCa5bblcxURbvHEhLG
8gebdlz35tyAvQdjCvWPlfoLY5TfSL5uEq+wdkjDPOy4BhvnW9lEdvbAhD2BmUR8
dDMQ62CvZZq1l4KXjUBrFxr7JSdZe4AyIahHwvpNiYV2GH85Fq5A4PkLI3pKhfeq
Y8Xa55abivYBU/QF8HEYQGRcbTWWzwYP8rePX4iiLO104iqva/5kvTWzLDq+VcPW
FLvOUK796isgiLBUrjMmA17mzy7y+Jyqc9DAbt3cBVv6dFF2lhvlsDZKUj6h3B5x
Mq89DUMM1QlpMNSXn5cqVuTvry0B625JFvZaGxvl3XpZnIpL3wEOVqJrRIoq0vlg
KkcNJ+Uv27u2Ii8dtFc3IuT4N7VkpBpR7GUZ5cUvqnr1HeqJf68PP9XGnU1zbSzH
QS+Z0eNI3Qic3oiXfOHeJ6Ik9nianH4LNKIZgNGwlIrreGh1PIvS1C1jUsx5f0Ez
wE4eeTTwvcC97AVlbJ3VAMTwSWJzMjU32rWwtM5IIgybas7O9R8xY3EVci2mpVZ8
nWReyIMDHAQY/Mgt1hKF5zupHoeN+PtxDnD4He6WU3jQ27SQ/S93HijXTalVydZu
PwelXGG2xD/myGmpPYBYEpDX0wlnLVq0PRLuUMH3D9w7/ZbNWZxQ5ADh9wENqSVM
QbMVuFCTvF2Kn7SP9essQDt5vDBzOBq1VOrz0Q3mQa77QG9gz/R4VeMasTZb24ey
bsXYXtUivcccFptkHdbz5mhbt8+jILGhUl7zsVBeifFX1QGmXxb5eLDNy4Dus0Jb
PJjYybHG3UgKpOkreEVdq2wlo9EYM+pC7pHXsc9+hhB9DO1LwPXQY3K3z3ayqI1c
ri+UBtGRfYeWDmPkpn2IK4K8ZC6uc/JGhdGkHfzKnKW+eLch8Q6KSKOEAJL8jWnf
5fTZXqQKcU8K2PNJES0VxhmopZnapjVvpuCtQF9Sa1VtKPqS+a7H36YDW9An7rT+
aHjn3hR0CHa6cKRa+5o/yGdyooprK/BBNQKA1MC/lMCoGBxibz4de21UYNExEHg1
NyM4iFkOqaAwExj4pfjfsk2oVa9UW0DjDMFvkDqL+Qq0vkSUHffXPS31KzUn1YH1
0E7ss7dzOfJM3UH/UXw3gpRztZ2WZrqT5pe6T7oRtfbHbC0RYNwU2xf8HODKsE9P
E4lPMJPoqxElicyvO+O25tM5rbpC8vJIb8XybzZWo85n0rTBjeJcE0uGEoLnjetT
4w38xdqFnWClAy8FxnLSrhZQ+oSWKBpAl1Li9fZ4m2LTeuomakuwM22cPQeog9Am
an3iiogZWu5kaXHNjGCMdkG4TaVJGkvPfPlhFJo63czysFEe3eYPYqxeIVHhJ2aK
qCfqYC8lTzUVx++rqQhqF6gecyj/NdfP3oPWDtmS24ktO+AiKLmoJVbnEz7UMfSm
rCdAFRA/Qjef39gWT1DgbjN0ihp/zR+zk2n5m+F/9v3e8ftewkl/FZ6YesRQdw16
QXydyxCLBT5BB4Iywhm/gHB0tO1vZoH8ti5pd4eq4H/pQe/w7iKegJ6KlPv6ZS6b
gJfFeejrBCfdIt7PeaMdeQvkq74Re9TO2z8rvLaPiuc8MYp0bpBy+OuP4arZoowj
TpPABQKDUunqC7JSjUObDbSDNKYOi8Rfhn+lt2dJ5Dxl0N+ag51Xem7g9qGZmYZK
SRvvdsJjhuLnzFNCkVHMKA/dY3VlDrpOy8RrZKNpzG7PngJhhjENMCUbXbrhR8x2
QPk9ETewD7MJXSLsizUrlmup0M6/pRB7/WvRb/vBRcN4NpnvRv+en1Fx+rKJrn9w
VVxPuQCy5vSIhhaIGQaqWgC0uW763UuHa6sAf8vgGi2mrvXN9x7DKjGEwgZD9hEe
s5yLOzar5/wdvwT/P/wOcOdlNBfI71Tn9JUW4hYCCbauzTDSmhK8WpDFED8uITWy
YAxHQdljtjMfHLNVK3R83idKQY8s0W9HeTaQMOtgmvmVhRVjSCzfUvfp3CbqcXg6
EVer8gHJNZin3/ymHjX3r2FWvUiqB6ruxKVYFT0dEaIAxDzikCGpfXjMM7mxRc63
ZfLBIA33PO5aBghL9n/59qJQdxDSfxSTUIpAXlW6S7egUiPVWp8ynCk2+qP29JmF
9GMF2zrC0wAwqcHWf8XzzQ8z4q0jLCYEVHgcu1zjg0zXNZ2idIxOm6ipThUY43md
DwKIkkEohAtOH3Zr5e4Bg88MqwqaVwnLtqSbB/PZC01xGH6DJXrNO3a9MYNzUKaB
wSs1EiAWgx029LkUSaGrTPerNoPQNdo0Lxu3qocW7jsQeCIRM9Ag1i28vmw24fa1
cSUGN7Lsla6IltNHly5tLnOxkNd7PpP/ssH106a1ykpF/HvKqTODE451XxkK+bnk
JshH/gDDr4QDPs6pIlyQQjO0+5rjOtnRZbKVXkZb2HCavkMOuFoCHPyBD80IbeZo
f2su2CJxtBq9+fHuZnOetXeb2VFT8vcKYhtiHCv1feI/2ZH5JsaF6LRB5uJ40+GT
dnhGkynOzM1ijDJD8Is0zM1djSwNzE3+5gyBEjMAK+m8BAYVkmobUt+LNT0SnYPG
MPU4jlyOBT+dE9nP3J2ReHFfd/7hcVvsCynfvz7sQ+XhAS4NlIuyM2P1IXK4TOtQ
8HTgvTmfP1b5T+/vhN4VBSSVrAL/7LJpsnZmQep9Vr7S/t1FG/7BFioQwhT8wpzj
1yky6/TOqqBDYDOXTdhBG0K79C56MwYkA2hhCaKoFu66IGkzNu67C6tjQIpijeDr
tv2HPkKWsQE7G55jRa+Zxibo1QiDV6xUZ9/LjfPvszwzJ8qAjh+gDsYPTbtDNa4e
FXnwRdtKMVdiBZMeC+jwSFDqxAOz7QG3uzhia8b6mqPb3fSw2sGwG8BZ7Z/+ZOFW
8YA+QYcMCH3Ln8kkV2n+jffenbl65tZjjNJGMVV6ixgTkZSRtTDxofvokMXxX2UV
wi3lqe4u8fa6PjlgzSAPQRgVgxIZFe4Sa5MZtxHZYDEO1nO2EBvv2rhRA7+/cw3j
sljNyIYz8VJNf38OHd4YcaNHaZ/t29MLExbQQsD1iA6jlJL3LTfT/VsZc1IbuEW+
/m5THkqXhA8NtZgLUtFLFOc++M0C2LWUSREfi3IgG05O54IMF/+YfWg/r2symfG0
p28xZ1Y3QajDzL945/4vFT6Mn0lom2liJy3SNLJibw/10gkXidz0xjZUmyAsqf5D
5E1eJ2t0DGR0gHvSDHKIzLWHt9egL3OqHRfUuUWEbzb8x5h2obDXYVwkOEp5TZ4F
lGaaAazTcgw7d0n/QxZdDcynk0KkfpQqRkIXJUlksbukANgtTaBjdOiPSvMCLtBm
0cy73DvzFNkI4gorGSkkOcXEWj8zINp6XfSvfPacEt5w4lyNZZauYfhMR0sjoJWs
221uLYWsaWc88YyDNCM8SzVkV1+klfJeO04QmJg+w36vF3D3R5VbtyNbvRN6ZeQ8
5dtj01vMb1Cj3npr1kJpDdXaDGADIVxTWDJAtVyJyvxvYZvSRtJbe3ZBsb5O8d3A
yR629hoa7KoVzpFSYrGTldsYJ7jxkUDjdzVS4cV7Gn5Ir1tpBoNa49SDib+nw4/s
JUiQOCU4vp3FCFJzvW4HGKQ3GEkY3D2JF5opXaMVTXhv0LWAy3F9Q1boLaO4wr9m
d+GN5B4GmBConVXlICZM5swyQmf2LRG7fGBu2F8D+P1g8v7UOfFU9vQv6GNzmoGJ
pP1T8WhUuFK3LKe92LgxiEKMxJpKK7qc6EVnbi5gT17iNRj0fzmmSl66iCl2sJa0
Dlsu1E8cVR2HgnmZyBZcxCt+nZNJeGZvp7PiPu/FKpjojKtwGkiPfdno1wShtHVS
ZAjjeDmG50YIQ0qaZL+ypTJyduM9Z1VjNf3hS4QmiXO5KhQfb5a/h28tMEvsysFW
nYW0jPYVAcuG86CAyFSzTJceDCKiX9rmMW7TwEIo1OsFrXinSH8cDI8hJ3PmMX5B
+tV9Bs0+v99rYVajg2ZFbN4wnOkbCpl7OIoAcIGdAL+enXCvVkRSIGqoSP0kYcpy
zIhUxSv3lulybKy2p4xyeiuVh9lBDTkM4SZjWqtbbDWs2YykNhoAyAZmBAtVAG1E
`protect END_PROTECTED
