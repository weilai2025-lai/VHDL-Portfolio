`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQ0WVasQTD9h0rMtIIkTOmwrUQuJYgQW0a13Ffb2l1adTOUGeqMq5o0gGeYyTFxR
zkiIrD6ZMYu7CNrOJNjRLTN8Sj/KTVed500JcSPFyXNeNZlZ5LwjXvzJTkGNvSyP
Zs8Qtl44728apvFpCFyOg2wAlkQu4P5HNTgvDK8Dm4diLhocQ4AewKzgK2HqZWwu
XYAV0KYcTbSPGwn8kOUaPiajOJnsbPOmBRYSDfINTjVvmPvHl7kyXxt566edzsKD
WGZtA7qZujT0r5+Mh7CTWuWV5v+SVgL3y1lRSvfsmQjQkhkA5q13dRJuJG5R44f/
BQtDNRxhxVHQIFH7HtYWiFctF1uIL31Gw+4GreS8QEPOe9pXmT31P+KKCmSJALuH
XFVXI4dQ27bjUI+VjqXJ2vrdB3Yfh9pBP/cpMoaQTvK0DyL8x3J2Of7BheszWJHF
/11EdMTBcYRb+zdB6Kxsbv8cLfrpXWr6vhEjbo6aJdt/DSNBEY3750+7+bYpJzhT
r9bRM8HYqNfki4DKZdLDS6ZhkC9jmQAd6pasTTVFXL8B4BBnGRkOsjAX/RpWsGBY
ldhSbzvRlUSw/9sWIgy0g8hdOiLc7UZUWgtDZAt+AywUNauhlUtcmc92vkT/wsMw
cF0bn8YzDtAQdmbq4xRQCYiuN6kDl7XUR4cQWTwe/l+xqxTkVlxphx6MuYh+rsf4
0Sywg5DtZKy+GMuL0MALhysgq9sXqFTFXOk9idW/ACAHzd/rXQgM6LigEQQgLGIp
Iscd83nXcHcRMyHRwfuoFRL6AbVwza0BKFolob/uMrjqFtSmtNuMuKKgVMTaqDqW
Tbh86Pbm/aUir34v//UUxQ==
`protect END_PROTECTED
