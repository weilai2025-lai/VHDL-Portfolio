`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dw7OWqX2DoAkZH433X8oxKFL+Ze83gpNBskp2eHphElqokw/yzdCSPvjZbHpIIL2
uyRQ9X1++8nMNHSB6v3viI/i/uVDM3caapxW9EU/5VMb9LBJUJH7mQ4nn8KlQii8
tZ467YCXuGiW0YwDRZDImfs3PazATR3XjeDIisbrAPxH8eplLiVqk+oLABDhwrh7
DqNwppn8yWGzgGIn9sw5bDGPDVkKEDBdOFqudOar+t7GOqUTYK8Mx5EWW5unftUX
HwTW57j7zEaxDsc2Av0Y0dPjR1U6RG+FT5pTC7Vwjw/RF25oSuAqsfJ9zuZX05OP
ZyxFzGjmQ5Yj7iqa5EnUvIPnXsxCw2YWugi5fT7Dm0cO9RlPmX6hQS2iyUowp8Fq
Y9Oa86NQEbcw+FOk4ClOD2/DZDttPC+KyWcEedfjNaxtN56+XkP08RPbLA5QoAnO
oq7sdm8NlaxVPUvpKdxxZko3k2VvAxIWMvOqZK52hM2c9BdFLuKlLMPLKJZK05q9
eaCuMyORQajvhG2ubUi4/SieQsRPdoWSETPXk2fP0Sv1dtlkLjH07Vm2xwXeRKdN
6OUISDCMotvptMZuWda1UmI1pSJcxA2Woed8Jw9/Lq0oHovggyidYa+Ht9epOyZ9
11OpeNG528W1eEp8RGlMO2+Vbe47yy1nZYRpaA8UlkR1P8QpYRHYyMzbSuT6zGvR
hIbNmVLPaaU8Q5NoIysb3KNmK12Av2CrrTLRHED1rqA3ajHxn0tNz8hBLW9HG6Xv
nGRrdjOajhJHkgcytSg40EDzBAOGibxvOj+TgUCQXpHkX1jWnO4QF1SXYi6O4NFT
z9SizCbwIuHozR4Spe0i4OaqNshPgvbEbW/BG/CaAKm7ABJvWfsVVx5e+1erMAnP
+tCCq5WL0yq0TApzYmAdJAAn7+It+XOO2BnVNAD1Y1olWJrduwAfBCVqyl4laifT
1honDTL71lASnVhb/yd3GI1JKEjYWJ4Eyj1QRZZjrhY4aqGv80KMfS7w/rvcd4t0
Z1DmpYvl8rF0rQkMDGNsAjwrbAipP7rOzM67pbGRbDhYrfqxwSKcZ8XKJrkU1GYI
ZB8pnA5rUtasJHRL26pfKJx5K7Y+PFnM4LXBYytDADU=
`protect END_PROTECTED
