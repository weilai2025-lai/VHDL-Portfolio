`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAHvvzgmHEp8bKnc5PjWyEsQN8WZVupjN1kGUmOk/iJzN7knspuHkz/iU8Wu4cwU
8nYajKyjPEsgS2Iqk/6Qo8tkVHGFOyef0NRAftME+VJ+WCcXhZtuPvmHmFG+WISR
TtNxn42KFSPFDk1eFoiM2Ony2m2zTqcUjvQmyLcee9i8pQcA1DJfNf7ywN5NAyCW
wmQZpQC7+v3aLjPtx8Gnl0kD9OI2x2kaT7PMxGUkq8q2Tgl9H/Y18uwmc8aYIBeB
SYDimR/P5mXs7qzrpXpkly14DyReZlo9AzBq39RDMtUlw3BrUnuxuf13P0DfK0kV
K/AdUuf1l0mLAwc/5Xb4O2PhoPp0U81vbYWyEopmRNdxTp35ZdQAlF4Dpw4iL3iQ
UOBJkDk/6IvBLRaYOGu5VeypfIe4KxJ5DDth/Kz6JvWyD+Dljsq/cEBBxlEEKe10
xeM777dhcu1uAxJQFoVEHhaL73XhnZ2qTKD3/J/E0TlTS6nPlXI5oBdQIGXOEpHH
vigvilZgqdcq2hZCPz9tTrNx7XVMV0K8OO909GCWvHcz2U6QbgDj1gp/kgVaD4uR
8BcKmOyi1mFfArB0uktAgK1NXqWrTrv/x0eUhMYvvSQOVVHmkJmfi6M424EtuMGq
tvOVw/4Ml4vsS0c6kX8drFFjI96eLOrB4x/Pm5SiUzKOVWs2YuJNtibpZZ9BGovi
M87BtnPS4s7XpUo+JD6/rZX/PLFNYkWS2rEnYiaC3iLDM3i45ctTVmArPc0An+2o
21tc0hoZNyeqLGM2/eDvkbSuUpMD06K9Es2grtSunPX2q1il5AftErZW+SOsEVES
aR6RsARY04qWGQ3Fp/WFfM2nv/6lUkRZ7uCg4HM8LWxGgHkIxAF0rfhmiYRFDGBh
JxBi3G0BWDZTClUz4/0PmfWhbFORZzjvmN4FNcQLtUHg2WSTFE51zFPik6tyolLU
QjLj2pNE5eftT3myw/yr9oYAz+qcB8VZoPjMckQHx4Uv24ehtzIfbINkKFmW8Pf+
nzlNH3u+2UAks/tnYYQBJEmX6gVf4Qbcbat1epVqrYUMVNpmtLc1UXmiLwwdYGj2
XXZahgnhypouJFolZtuqEHQB4wfyIBnIJPQqFoBuMhdmnQH2K/ALDn/Pjpt1RRmk
BIi1Q7z+uW04Tfgao+GzabV6BbV5N+j0hAofsO9orNCIfO1qHkHDFpUG+Ln5qy1B
qy1DTbB7NeAZQJQSFKMcCByl+qQGJZjnwQJrtj7BPN4ayrSiKAPfSCaGqazWZ8v4
baRSkhrMEUHlkFWtWfYj3SK0+emJm5EEg8jSigK6Z7teUIMn245ollYDvjO2lpZq
VvY/fF0A4OHbqEEkGOgg1OOhivw5gHsYKnJbIWDQue8=
`protect END_PROTECTED
