`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7jI4qv+Lq/bJaPn+f/E56C+Em5cuXC604TiSNN1D/lnq74zUn4v0HdAxpGdCU1Pn
GAWnerVYk3AAdASQU2hJsjjnUFduSWnHSbEcUjZz5jD5+QlfwXh7VquMstpPVElB
LrB3KatzOfzV16E7WVGx9wRsdvu92YGL0pRz2fCiLEGH7O/8NaHuB/y2r8VPJ7qP
plAPMKzSLIZD1z4w4MSocDg/X4lVSxjUjT7t08XHUqPhXbHjswUdICW/MmPqHIBB
XcCR70jjS2sEU27mOXfg+and3rLS+6f2O/7yPUNXQwzo/BzdSlo4KJT7iqy11ccK
y547LpRambIq82U0aVB4l2g2SCoTw3EnGzL34VR0Gh4QCQe8SUU6+o7MWWf/cjzx
mV1RoTUnPisPCD2m0et4gcZ7Lh7m2DnjbP9IBJKqvFuqpASrlJAy5W04BLIGjWF3
w9Hdf9maYQg0bYkco5ORAk5pWp9kEotp/LegoVnqIhxFn2MmcxgFh/MpJxvHNfvN
leFJRkScIJemqdZlMABUZgZFGipRa7kfjMgLJinZqm1lBvOyeMnZwBIsjYt15vI2
y1Q+2ep4eLqjgjk40GoNb7V8qi+703S4VLuR/8h1XwAA4pItVE0RuW2ZM8D8vy7/
oc8kta0z8h1HUXz1VhXSRE9lDpJ7AP6KbkBy0M1jzObIwHi1T2C/Uekcc9gcx3Q0
H5uthJodNDlF0nNN8pVJyP9BwbmDMG7wCsvFA756xsGNM+IAN/7de+JKpPq/mb/M
MMKe4+mOAg+CxoVU6iCzvkwFuPPEuU/UfqP1GkEDZB0YL2aA2cV+6rW83hB4754U
/G5BhAwzejAm9O3a3qSLsaK8tSCKBtEFUyp3h6LpFz1l8/meU/p7nCAcNh56gLA6
YQOJF2nuDOTLC+l3KO7EZ1GRraok7qh/QxZD6GOFzmztdx0L+pm6lNxO9MV9eJMW
nopcZayhQhlLks9bZ8Tdc1iGAB59XeE3tXuQMTPLYaYcSjvgSorbugxYo5rHvGms
DbSc2aiBe40pTq4eIZ9PdioJI8e/PKqk4seSC6OxLKOAAhMaBodyYpuKhdB0ymhq
zbKFvG5QAfaoKxdw5NTXPpbZWun3kftR1DwbsJnVACP8oV29GhY4ac84ees8bbx/
FrHRt35lN/0L//ijJ19G0JRKaNKt18sJHzl4KuZQXIf+3aYCqk7YCS/r89XOzHJH
olGdKzSmjxxaMaDQdPy69/UMVbx8qsU0vRu4VUbUn/PJX19ROFB71PV0dlAQwVlg
0basZiUGCGeSyXiZcWcB483hvio8o44Eqcsrku5jUQaHANdBUgkdjgAKCHwliD4W
qRWzvCca7alHP5ZsN46CUAZA5UNh2nWH2BdDXMRmWDr1FcatsVXiDXGIx2HC2Lcw
HOqrYIGFZg+Fr7Zed7oSy1XsPyZ/9JbzLYOVnY7PZ/C0Z8jqtSVdN1eFGUbt+yxe
SII2HvIXHnMrh82grL26TrYLKenFSPU3u7492wjlGDjU5bnVNfAH+/AgqQedwgUL
t94V+bQvSldKHXLtmj2uUYQu+zoyJ2f5Hd7bUSbUxARIv1mURVB4pGeebiJUD5s4
ODmOHtRN7CLjdo3m67Ww/N7jiKnDoeIIHy8QN4TP/CQaAT+UKo6PfAjv+4oRGccF
6ccFIWjfOgv/4qz7RqEW2VXbFqSx8iBR4PW11HkfsWdE6mfYpR2cfPJD3ajGd9KK
LaG1WwoGJ2/3K7jkuqHhzocXmKd09GuoradPYiakAGOSOhqHAmCJEKUjfTI5cSmF
J131YLz3RiJ8MXdX+tBhOA==
`protect END_PROTECTED
