`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yIZvYGuzwTzByZZXbghxSXrVV+X5P9lST6s5ooDbKjUdNJkgn7tTyE+VBbbhOOsJ
wQLeHPAiyhHnVZWh5LtOaGNUO0rIvsqQvJHIu8ZxGQQJzTgrhYJQUbB2pwLC/O/y
FPNVUFycCR1wImZdDFb6iSybNQZe3HFu0wttdzV9oy0U2FMTUsDRkvDXbrFT9asA
VhEtaRDU5dggI+y4RiBVaa3Hcjb3DMe6o1ipVmDFfVkB4dVL/SgxEaOyq+djMZqZ
+zjm2hTXLihcAuoUaqfjJLdqlgvmJ/qaKilZ9Yd5qI0HzC5a9dBS6TJ0rw6JFRyQ
shmgNMPo7AzTO6xKwDBIhtifebV8l+TK0RWlTOZ+D8tcSn8rbWN+Y1OWhOvIZMKi
M2UrsUD1KKwZ0WwkLPzGRE4kbK27NHqUrs8l4jncIac7ynyF44C1hhxWHuRiZmpL
fWlmNQxSqS0Y/mB395XXFvd76aDhdIGu7bjo0hJKeNl0nCcaVyaf/4LZ+uLnKv3v
lPv39UMCNNfMW9GRm0dkyOQDVsaSoia21QV2XlhGtXragmv0+pb93c4AeceWA+fw
gJ/i8Y6tsCL7rjB7A8QUwH2sKNUDE5Am0QDDLJjTbXWU2xjpaUX9+I6bfZ/Pfhah
I0E1ZTH6V67bD4ipSymTGr/DWjWKnHv/jbsJk6n2eK3B8pCus+JgZCWH9apsy7CQ
BcAxcZMif+jR8KiDnKbJAfrwVf5gHdKTVQQMJ6aIWIGQiRvub/KPm+uCKbVOK0il
QOdu8T9Gj+K+YMjHW2TuwGvX5bHSt71VQR4SIVoy5YGbrk9gPsEf6we3rpil7lWg
iiRiMfav8XhAV/jO5tmSQY4aUe1MY5GBnf/fv5p39Ie/Puk7i5TsbSnhu6rtUpTp
vpnY6l1ijlxC9C9DE8k6poUX9SuX+cdC3CYg/lyhxMYi5qwvE/1zJNi+cDY5jU1L
B9BLOmfQdgDwB+DNpeJprC7VaJHXJ4G7tIAPcbnbik7iur5Z6K9qKKl8J0OZX/+/
CJGuwR8Mn/hbnDmOcHYjcXiLMbrdzoB3A9u6aRqyaCLybYXBx9wFiCu8rzXomnt0
6paZ6G5STC6VDsPR5k7st1w/w4SPV5h0yGkRGCYhS8coErlafLZt/MPTPjnS7J58
+vYow/4L2oGDOvry4g/a2yQ7krQjzF/Eq6Fc4mtloCz1Hz8Cb/cbqN6mEQ0rOSsZ
+jqYrgA7QzV91O2UDDLIR96XvIieoGaQ3vmGDTJLBJkxmaXDIn453KBJt1n+6oNd
BBsvhqmSOgt/LkcZJvvzDTHYI8rpXg4gp9KqEFPh6kMsWALAYB1NhfcmndQVheRe
H4vcSiejA6fmJuhS4sc+ZBoyikv3D3JLwZMkzLuk7Xxn+7KNao+MXq7QBeDl5T+a
3bPm/kbT3Re0Mzf+WmCo8FpgYhIAVM7gLZoroX27E4kZnLUgxCC9G4qaPW+JepsE
g6HPBDlVgmyB2FRIZEbwHmAUqUJgr8rxDA7UxqkeoHjhGUsOgpn7Uqhub6pwD6Og
p7GXzXRhy0jnAhZDNegfZw==
`protect END_PROTECTED
