`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IZ7yr2i7M0OdmRVHvnnIQgdAnDDxok20xco+ReF56Qa1S2zDmxddqaWqx6pIIpb
fgDgWishjWUvrGlakPntU9HnJ2h8BmZyn/jjgNb5gjrN1gR34KH/4k/NLkK5ogEQ
LzMW0c6a+OdQ7+A9rKWmlUfChtmA1lK+QDNTIPMG+XQuidQUQk+ICfYvgMp1eBPQ
6GmOx6T+GaQkd2gL7wCfzhqLUs8HDbJjNkh4KsjizrDcaFfwJLw1+bLKkeC6CBDm
lRac014kqRpkMgsy9ulnwQBo+rS9jjthFdhSorKCukM3eXwM3030CjjnzmM1Vp3v
kWqQUBk6MqniOSJjvrqOolecFJjNdv0r51gdtEeByYsEh7OdBClW5vL/mHAygxSc
KFD0lUGJh5OLHunTKLN8Saoq+WaM5aveZMQeom/gWRW52pct1IzW6ubOvfPLwMAb
u/Yx9zKBEbv8CfDNsiZD/QpR2VmxuwzdYl/0H7Jr64xrL+IB4rsgCD1sW9qykWjg
wiIuKvP/iZk19sPeLKFeD+tkoS9fQsVnXtJ34zB8JttEzVuK5yq1RYL5x7JvJDHs
xwPJZ7tWNe1RJ4I0brnBEYeHVUfDbcxMpdWmr3C/OblooryFYaM5JVH6UX62y+6o
Gsj2tgrCHr9QZ1pre6JxhACwJG1C881w3uoBB3tsN11ju3tUvNXDjUsPShJD49Ok
vz1F4Udd9/qZQ05F+59JGLZrGih51vYsy2t8P2pRPCqCvSyurpFDkZmR3i39JVf+
tViqiPGNIB5PVCZNayPRAA0Gk4quplZ5aHLnfAqpLdAEGFtxteCi0smKbuvfOW+j
10gwILkAMu2anUl65Td1YS9+OWMXuV8Ksg/sDhVdMEqtNYmwjNKcsjiwwAprT24O
C9NygfxdyrTOnvM8/ARnBIDiOc14n/xmZEyxWZuYs43SPfXQLkdEmSVruHnhFi90
wjfji1yPj2E8mm+bSj6JbLFqAEQcWqrDWc98H8y1gYSp+xTZEZZoASZTRD9J89D6
VelYkpUY0yUeAh0LvaiP5r38CEAa+SRUyOn/6Hf6GdImKpGDTFeKCQfXAMw3bVpK
10UFpJWG+unlqagmNhPSfJyvrhJ0X0i5LPRZS6gbK/M6la1QvfYJ1a+hNM8QOKPB
D/Pw/g3JozRjXiNm7/+adKgnqNkEa4m2Zr81TMuf6Ct7g2WiEKr99EPCF/QbcRpm
YD/516HkvNZwIAx6l1/OtmG9Li6KHoOA+mlLaymOoGltGvTKjcg4CoAwWSCLcwZ6
/5SeoK3ysVUDcOlCk7qfcVk8v0WUpkKMa7cCdVb58WaZxdcWeGDCtnMlEtlk783T
KJuaN49VEz90P+KUlP6BZ+SihxOg5gTKEkLfUKteuEfhz6ukVgQietyyGLITgNpq
6IX78hf/IyReoVrMjA+BcGzHNjVTNVrixsdSZWp5IofpczFlBvM7lRrfjJj7Fylq
4iasF6BE1y0hX+XDVgXV6fQWX//bjtlLfTHavIt/2FOTqt1GmMaiIIFi8ECqjdVu
eIn+ByxoKoUWuJlG1DoiDbQh/wZrnD6LH+iYnsK4s92BT51YBnEHodEjw0lsz5Zc
paAvhAWxCks/TQ1EVrLeBOXl4SL/ZFcUX38+rjQc+sWXjVhW+K5C447NzsczX88J
8o7HelMQ8Fe/5Ka2hIEJFw==
`protect END_PROTECTED
