`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JhY8XkkKL/FPr04J1qOeW6HoNqpVN51ylOeZPQ9gDLvl7lVBo1Moc8sEwn+Z3qBY
xjEim1d8+KVI4S5Q9L14D1jgDkTbhSqlr3O0DxL2ym8hUJ2GIEZt3pjqbTJ6hEtR
6AY0GkBNn2CGkWBaVRzGpLXIStUcs710k1nGYejlkBO3/xq0AzUBhywcEgyncS02
hzxRrV0t/Si/KkFiwqIYU1kJRVKv7zjjExfu3lMHfnON5S8nzwZ+8zfVv31Zkuzm
J7wRn7NLyswayAYf3FXkIpE04I5jPWBmBhBmjKmHHqeVSigF8UtMiPe66+RPDJyq
4uLmaHXzV53tsX/XXF9Gi44yHOSRS+5k0vhZILazxq69gOlYQlkHWNswJnJ3/VW0
/OkrelX+LzTUSd64BMW95d+vfar1g3g/jU2BHZyR7n884W1cfoEBZ9NYMIboOmjD
zUX4cbhIGp7QeX4HeMYABY6MmRFqX+j918vNZYx0mNlbtoIkPhHDimHSwO2mVhsV
bCRyvTry+z+El/C4WSc468PyTpnPbwFWcgWudLHoN95d/y/lg6kIvLVTphWK9aB8
ELiiW7GzbJfW56aTak7l9X92a4iAPa2LrtWWqRr8DT7qh6z++TZheXKGtfqyhUiv
8LBAxlsjl/y8FNR6NqlAaSx2kSYADKCOhX1zh3aPjbZgpVpRrChvSb92gTYVs3LL
mZ0tFEdtdiTywcPfjcV2XBxrMTuxRPd3CGmqzdCOeVVReYVU+ug+5bib9gtKY4ku
APP+2MyKRZjlNwVUBZKelJ3oTdxQ8EXf/jndirsVv16qzgddzjs4Fsh2DQWn3Om7
EvKXfL2jqN6FJgWSt2t0wWRpy6mPGDGRQWi3UUi1ziKsxmnfBec7Oq7ycTCS9FaD
vDgARMBy0GfLGMxhARODzqTA5+b0WEt/Wq+EEytEo/8jhCr7bwqGnyDtEqf96X6F
uFsGDlUYLbYbp4QzIxkiUsZjHV4sjCT3ErnzRYbvWu4gUFmW2I/msKWco7ARaPys
g7kHNSa1NviAVxFn8NGtiT87eAvNKB+fWewh6PG6iqgXScF5STTO9xIn5SBU10/0
`protect END_PROTECTED
