`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NquECtaFSsHZw+4rntdx96WDCwGOJ8gzGFcndxYjlf6oa+ynxn2TRHLgE/Gj+Ds5
mCvWU+RiQuelb2LKwQIKxAsXBJd55rY+4I1+iwJOxM7S/ElcVKiILZe7NUIwGW1L
gVZn5+qpoiQU4Jt7UjF1cpNPRAsmtsu6IgA6sxbqFTV6s3ABp5f0eOWDux99yw/i
AYGd4quuYTjCmmiyEdBSe0GJwwIbSr5QXAlFxXg04jiUhjQ1ybO0rDgsqgi5JMx5
t8+tyF6wOgGsT+ae8hGotNUrz8/4eddD/+m0fOBPVLQ6MrPQyWMtYQ/+ZkT5Aymy
iBKvH1vp5lrC4NyAfn/oT1E7ZgfOX/yLw/95qMa439j61Oh9/yCWanJcrHD3+k9U
kfXHnG+g1k4T9htZT3nrlqqmQrZIv84whZzOM34ijHk8vW2jOXGdc/QpdPpVpdFH
fp9uKwAUE/FqIBN3T/WsMt13W9Yt4uncgoFyBzKaSU/XW9MNkl2kMoypBShedWVV
w9eco+w9wfU4HX7xzTlVc8dSLXmBAWAz6mfVnPpMOwCKVneiSn4NoRMm9jVE9Q/z
xfYzEtDkUUF0f9Ko+kWugm5Wey+DjmBrPIZMXZqLbZIJT3wOgsyZIviYFIo8Dp3W
KP5EBcm0YswmpqciYlSi2s/lkw2y5EAYwL5iZThJj8K5CkgeOUEcK84ewSKg2HIv
161LNLKobw3L3uvJIsFF6g==
`protect END_PROTECTED
