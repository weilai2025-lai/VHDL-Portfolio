`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gf0UQEUzMIvgXUGaxLwnhLF7zg23BI/F6cBGWZQmsJXr7zVVxtyMA/1P6yQMla5h
agADE9G6FEzsgsgyarx7k13MXGXPOcqZEYai84N+nVFpXcgLwUOlExIDd4ifffR2
s1s63sfNg8UY8l8vUo5rUBCZRFwx6KsoJL3EcSkLhHOQrPtlK3R1gEOyJI1dw+rX
jjYvMciM74U4gjMXP3jnLnOt3cFYcKIgb83It9NF4pLBHSlOW2nEEpyH/VKTT3CG
B+pAwlB0CG6qJTKBUGlIXd3N+FP/DEbHHoiDTNQHbRTKlq9qNmBwlMpkFty7H54k
HDnWEatvRdFDggBNAVoiGAq+Z6zlXhM2FDJcLe8iQXIYRjsv1WslTCe2OVqtVkb3
7fZr16lXy72btQHOziSBDemN/+PNYhVpuNjYZ6OIebqdN/rQr5r44QWLAuMT4LoV
mi1ofEKguSEP/9JPDZrWgqUYrqEPz2/a2ps/eZGU317oD41wY6XT1HY8j9foj7gN
FCtCydOsNQgbPKSweu1vpw/BEaUQM7tnpysjBODuyn7jTpGQH/cbBet7lKopjwdy
TolH7PjoKVe4TzM8I4UuX9OBgBpOy3SVfBABuwY7Kza44hbM32IWfNAYBxMcz0Bm
Klk+vglytYVEfwUrcfiWp2u1keU0Jhi+At1DMZVLa0fhYpcQtUgXQ7a3BAfZUVlv
Au2bLaMoI94MZywTDqwwElZOO/FCtqfkxErti/mruOej2bcRlbZ/eLtdwLYzu78c
tGNcMMH7V46QIgSIB0C6LjI02h3QhwJyhR8USqz1e/HSQLKnwdvxGAuGjiLR+YgV
7/EwjnuNTKC4zyCrM/0YxKvfN08S8gpu3bY7T5LUhZ/iLTKMOgTY7Lmowykl1M8k
4YucJWFW0zFN8zXmr4l9TWccx0LmeTSJSkhRfkqGQ2KoNwnA7hUh2U/UAaG6VnFl
caSEAe4ib30KPg1XkcWswIk4+qcwbldW4qnPhKue9ttrRfvIdS4MEYgyRmsZ7Js6
zCaLy0g/0Y9+12ocEmhhBfcOWrlfLdpR0kmQSIpclhu3WEgnrLhyz/xjZ4uXTA2Q
skqd2iRWP5zG/HUSV+Gz2wj+BSAHpumAtSMrEbmrCucyoDRAvFpIh6oGZe76nB9Y
8ESqPUR0LC/uiupl0IjETZkqi7WP/W7AfgD8ylSHPpG3RdMBZxElcWwvR0gO9y/Q
GSZR5oLS8NLvmvJy1vsFde7BX2SZtGsZHQT8jTJRiLI=
`protect END_PROTECTED
