`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLxA4B0cLQzx8bg4THP7b54P383erOfb26VdaKQ/jJDDtvblwsBX0pq3pFxyBnHL
voa9ixPxH6siir54TizstN0Oj3ND5GSGjC43xhFSIPDS5/BfNZONHDLOidWhsA+N
m4SNxTt7lAygZx0RA2oFgNwad3qDAnJ2X/uU4HKsMfHuZP5a+DWc0ALGXjbdNDg+
IjLH7p6PJ/KeEa4Uxf9PNf9PqA6M6ap2tXrwqDeGtsRSNR3heJyNhvDlzOaaDYdS
SL+FH3pvmCIrgJXu0g5QlFpPg6tO72PVTAmwV31Oe5U9BjFQB4ja8mKkUx5t462v
eWHCWFKZPhW/7lICvivG+8Qrx1zVNTNFAR1uJxBHU7evcbzMWnc+qaDfNmzaVXoM
P5H4gRBoCcg/xUgVO6ZIlTjQLfgyTMxevT5xwZ/hLF6ObFu6sMDYkSp388KuAVp7
VuQ54LFgGd7WAVSmSIulH579J9xZHjFeFjxlDBf6WVfuVafp9WfqOq683lcwBgZk
bEtYod6ZGblWPEdv1SXOJ8E4GZtR82aHMsTDHa7K/VppxkMJ5WSFaKe79i+8yVan
7aE5Cv5UR10cl1/d/mPgc1+WZkG/RL0u3MdQbvn/sJPdf7F95oS4/5GEy87Rz+cb
66RKJhIopRFY2psWED3jsx9JFl2r2ipn7dOMvniQzYN3M6GHJcxkF/ibmYMMTvUd
XqizwG4q/X1Qgrnup9ip9Nt9YMPjzs1s8+3eze8A4UEXJ6e0YF5qUE8UQ6oMeo9e
gx9soBNp7VMcz0L24afaetpQxZUca33iom8TT3odpYfHkmtKg8anEb7BIfLrPSuu
/oNhbNSuuyHJ5PiyyuHc7/PPBWKXrPv7MT6WoLiqE2OLFjNwV3pBfYgYOQeU+DAu
xB72heKyQaN6d4PDaDL3YENoTJn3myVR3XoG96aCFsDjRBBsLByio5Dt+R6LoqXW
9quQruQs9AOzinmRQ4d26xax+GoHfCVMvu841/x58EuWS9aETpv6J5KEaDVSdPZy
/nqTHHq6ghIES6GjNcWuKMHIzYV0n9j5KYMXB8jxORHpFiw4p48brSRPBaLvfWnp
2uJ1gQpTFJT47UczLbzzUwbLTVRf+HhINwUAAMbNK5T7LkAzN++BoGrByAdcDDdX
2VohodPBVq/K88s0IvPLuRO9qod+x7/TIZIWnDWUOW6907ZegalZDPrmUNS8q0Et
FCbzUDvcuyacb5L7UQTK//5GMG0XN4b2VTi6FoBdAXBAUWYsdRoWkieAYnMxfKce
o/Ar93doBuGG7kLqD8B/kEYVk83sbZ6FLZlb/YXFZzhHawcIaDrI1CzNcKqQHnjN
4y05IbgUthIjBsBACdd3deyCwE9McrdO42cVwxAxEoYVbIDSnUG7TvvmxpPiO/yW
qmKVbwKkUAkd+ztiEXxXfy+L3nyE25HLwNA71FoKFcWPyjwUaSZ06qHnujN//nUm
CEuhrvVXctTTst1inw5twYVeAuZv795aLhYb2QhnA03VKLqptGkTTviJioEF+0UG
Uo+l8ZYISpyw/Vhown1rmH6s0/S27pCrw1Ou4Th5FzwnkWKuF4lxHU0LrPKCpa/n
ZKralige0eXvyUhFXeRaYys2NhySkal6XdEd5Zh82jxJPefVr0cFEDc6oAgimzh/
5weN5e7jodhpp02BswCwXa562JXYTCWBItVuai5Ch6PDLHdryNplzW3FHM33yVW2
Ajp+w8D5RJGG/fANlKKVh/A5KQ+cw7femzIFenORfUmF1dqOZBL0blJtNvj2tYNq
sJqc6hDQkIXbRz0r8FmbSGx2HOhJ8Spe8ACLpMChpZmDYADpsZEpn/3KJ8NdHBgh
/B3O0kmjc/NZKwEks/+UhxBNy6oo/Her9rk8y8P/FgTNfsUlgF2CBHCotMAc9oTx
2a5PjeGHwnR8CtU49YQH06NiIQ4XyDKH87obdbePCOmOCPPJzgqh8KmtHI4yPMNj
C6HH1b7YXEUbYDPzdTgWMcI5IMundg5N/yqvJs5nPKEIJQwfvgtGCeJi6TRyooIc
2Nolb0qvUaoMGsUnUyqh9pon6WN3vTpnawaFh6SuwIYsfyIpnUNw4Bzyy2MPZhVT
UPJnVylCubyTiGxnpHLllBoVez5MwtmlvbNYJphixNSFdD0myVqRHVsQJKznLDZN
BWFXQHZ4hmc3vaeLkDKq4GYWUhH4VafMFiXpZ9bDV4MG9j4TSgxT8M3j0VXMJbUd
fIB6RB2AssxoiE4HZ7zdOT1y1x2/5Oxz4hZmWT5PeHPiX45RfMfbnNZAQto/yf1a
TXlLC9Dlx61kOirCacC8VDss3w/2sv/CivNPxKbn/DtDgXRIx6ku1Pnp/ww5t5sM
6vX65dBpUl1p9u/mK4c5uol7LWPww9xCEU1/EU9JgmIz10qMY6w/HT+CZaD0f5vu
tbknpbzWwa+pvBEZc2zucHMj0gEMDJZ99D8wB0K8WethpQUb/DryeokfIMChNPF4
amVc678cWV+t6oL1JLPEPUCT0+otsj80j+ltT0j4etdQbZazWXQH/yKySM+KZ/tj
W9s1Bv8Dzjc0ocznbXGth79LCUtznbK02nzpT3CHnBWOWqXHdXLlYUVw53HOF992
NrWJtAwXeaaixyNeNryXuQ==
`protect END_PROTECTED
