`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sE67BEbTmmlB8MnPAWfj7qmX2fU2M64hW1RyiSVICVJlXyYMp4LTbwU16hsJIxNQ
rhfzCoK3hqJ1FHBVgzSSeZIhFEKr0TfSiYT30vXkNyu44bCW8sMHOPHl81eleRKo
nCQI6cVMN2z7wUQiDgVJrGOIGYNhv+reA6mkaSHRv5DpCYp6fHIm8lf5xV5hPF0d
WeacMXfJrUaseTTf7wZcXK2ohfYU9cjHQAPU3p5ZgOfd72T46TshCSm+sm5igxrN
pG5Mej7cB54rCx1zISFX7x5wO1Cr0zIN/zVfSyKxVZbiVlykEN33m5LV4u6fbUm8
6m1ku3vflPh/pR1u3kYqzHDb3die1IwIaJegpC393JuRh6pt6PuF0NrsyqfkPb0C
RMnftOCwo3J+BPOg7nqUQVIO/nJZJhE6cFJXzwwNRpwgya8EWxpRyAWbHuEHv4ag
k7kxHIsJI4WUSn6EME7Dx12+yqg6jApy0/la5x0QUrPJyl+F/O5tOH4Bh5Lt67hY
J7BySj8xpgTPUSy0gEgCjVq9jFEwHD1YI6dXcHI6eHOyrrUYfhPkelgiMwPr1I3d
xUpsNp/UORXbNBRSKhL1LAeAsSmr29YzcYGZQUuIcno/fIKnSsBxxpQ+3dfiyrLH
lAI+9ikrMl2Y+ymEKLCNgCbcZlr5xVA79/lwpfNca0oGkFgazIzpLJK0LZBRp2fo
yXARVlBAlPKiNOf3M3s1rP1Uq+NSecTBJWINpPZq+1eMP5K/AA8ZGH/UUVTKFJVB
tdK05EyIBnTSBZowSdXJcVun4ysjJoZDuidx/zZo3qR+rnTJmKeiVUv0zQAL1EgE
VjMORCSx1P625FFCjsa0YskQzQbr/i1bTXQAugQ9J7PJ4eiGo5PXDn0Ks/c7z6c5
DYaiupJh2JufWsIQNerct1nWIFSJrvuhgA3xAfBTYB4=
`protect END_PROTECTED
