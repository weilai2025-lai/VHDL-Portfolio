`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tT5iGXl2UK4p0bKZLkFgeqtU0Vi791A4Hjs44a2Qa0dQFAd6HZurfw/WgTRPHiJ
kzJVvV2MfEUJYbjwZHWR00e7h37wZduOwWOJhL/Tz3JvR5QtPDfUdRNXxMicUi5j
DLfmLIh/kOjkBoxlhz8eZV+Zxr+XRIrY8Hc+Ezuq2UY21FtIkJYNdMBwP9HgkDAS
xHhWVWs/S1TovZsBV1at2KVOUZVtsCgxHbLgEUJreoAI0Y7CHNTN8X24g8SkaDA9
VyBY/2/o1tGURtEn7Arq/+Zi/wsjNJLxOOpbzN+LVRSoZBREqI3Buc3G0guvNehg
3aMj+F8+nUkz40mM6Xj7TaJ9jpffJVFF7xn3++ZS74p+c5d+Wcswyk0sGjRF/Vrq
MW4sfBHwWNnksoWQu7zwh2KLM4dR1fiMuMEukv416zC09jRO+MJ8tkfLuRWwdSbp
XYgupYrE1wppPyAt4Bx9j0VBqT+y8o8loPMkTm/+Wll16E7/CTcKM3XvHzN5QiRy
NURXmYjSSHub8N54XYEO60ODjKBzx8n62DICZIrdtMjV+YgSBxLkAFQeE7Q5sH3M
WpqEw91NZ46mUGTPInsnK68Ofi946Dr1/QuNlQ5t0TAOtQ6VOlGySDXAekGZhuVT
RARLxRmUbRHvR8GYSZrDWx4qmENMEZLO0xpRepeAe9UbX89oZbxorwLRVdcuLI++
6GNU5CeOHrUD9Kuwj4UBED80hvhiMJTBCoqz0kfDU7J5TFapm2X+M/0BLfH9Tjen
f9XTaaHY8TjddZmKi2PfOfpUyjcyNAtpZXxs4hz0RUcVyEctALZsPW8vNkSk7y/O
+eeweubj5X5QsQf64Ry+giykGxTlwiDSZCpl2ivBWZWAI6ikFnbKK8kJotA89wn4
yBqiOLm9uxCKZJQ8sA/RTgBBwb29KqDf4LmgKWd2uLm9RKaieArLWJlc0Lad+Ki2
2CQojiS7iqBeFOlLs35UVVky4uZ45XTTeIxs9JfpG1oO0wuVnSEQ+SADQ5FGkGov
2bibd4yBd0rDSpkPVf6f9k5CdTRz4wIadQZGD/C2qMuxC0Df1lejeU7up2E25hGU
Vjf+WAmXueeR/r7+Dh2KSCtLE2y/mgEnfJ9vxy2sK65MzTeV6MdGa/RZe0Ox1azX
7knkfv7u6vqqamYxAQX7lrRj/SR0BqCieKq73aa6QFN16JfbkfkxGGOg0CMYCbLu
DcV9YcX547X9O4zZtzkrrrDu8W8RroBVPgHk8u5VbBD+IGZ2BV7rxHhOWFESk2lJ
+laykZxNDkMLP7ZsPT57p82oE2deM3TRFFf7Zr8z9Ltu9I+ma4YfVfJK2QWNAqBS
sOj/erxA5qIyWJLMCLqjgd43B7GLVjS2zgUkZLe0Mx4kdZDnGJZFE2hdAznrXX/U
wvEKDUIwc8jiuydP73iunGHYsbUuDa948CydMBQpADaK0y7dVnNDB29oDE7WyRET
2feod/oWyEBHE/ZArWyQGa3931EQoNUDxE13JQbas+J1RU8ge1NT00Er/wUfgTi1
ZItnRHrwaynkmvYwF0IyObhjps4g4DKMFtaf77STdEDVH1o6I3I+/7QZJoa1Wtm9
ybNBaKeNdjMBbjnI3YdBT/PDxLNkA7jkNRS6Vs0DzXv7rWuwip7CvQGsdG2H+MIC
heLHg//NeHWVdFQ4nDRLYaEhXs+ToQG2qXDo1hhWmXMJsx/xhQnuxfQeATHtyDYS
rPEDuutW2cEDOSw2bN7drplRMh08Uza7udRVXnccuZIlF3PJPiNP5GTO8w/5CgPH
CrBa9WN0Fh3heDj2vDs0ike6wQZyIaKzrJAEsbUqv8HLAThg+CNrVvNEFuVVdjtw
DTgeAZIyEtON3FOO/Y0amM/hvDJFa6Nf5Qf4JdMvVeOyuCQylVdzKQb42Ka/IjFw
LO/C1x8n6NJ01wI6NBjYdOQ9+DabBwXsRfl7roFKA7Xr1BrXIohTssUc0VkM8YTz
HkjImwNuKg5CrqHnmbMLwZamTMiyjKG4DbbgQAInmQX8zO/sfLDTbVgFSQFhdFej
pYYxaYX3hNGTITm9ok+vtcww6mEd5VEOZNRiRL8Jdu4IEuhfZ0rg/l4lIUDBB4lc
N5CeCV6LJD+Ip0O7up2JrtNUMswyagJwXm6jI4xLTMNkDa5qYoWzd0YuVeQ/HzyU
bVtJsod6lplrkkWH6txBPNivoLaVOPaTGoAlNcDnLwx+b2GuNebXFeXU313mElyS
RSQoawnJ33oph3l2QcllMDzmtrAm/7m4TsfQn7/Thob6F+yROjEQxqP+rLE3r/NK
I6SssKUMSFP8ocxMhaV1W2eCz811q93D3ork7ZC8KBX82vriKWuj3Y/00KMzdjJd
/j9ggYf8PQVczDqEoPsiWOulAvaV6j0oc03e7mzHmrsSjHdM5k3jkvO+mlMucuWO
fdDMeyQXg42fjhNEaLkcdZmZ0nL8Hwgz17mWmamTFjIv3tNe600StQzq7Li3AamA
jBI+Be82SkC9bz50LVAXDBqruIZ+KorFSZ9kOFX0V3lHkZuVgE5pwsQaoIaBfL2N
msvFQEhdkBQ7ETeXAPIToqlWNUsxHnqa7roLu/soSU4KbUsVjRdgT8MUaThhWNNA
C+qyGQUVu77TeTZrghJq3wS0TrKZ9lKpGLO1ZWErT2Uq5r0ahWk9Shl/sBtK9uVm
HinJ6/4XB6Qhop76b8rvCC91reZCorWnfxK2vLLxybgWEe7+2uoqDv2u7LLQMhlK
wz4nqgAHkzgolOeq8eUpjdKDGuPIin/f0k7j1VpZiBK1eoa2VtF3xtyBUjGue1kC
F6mg/snk4KYhd0eKkBEYyteEV2najliflNYFcUY0SXcXcC98ndWgeHLl6VnDsr6B
JH87T8wAhuhaFlrUK//iEgBbQ1hZN6lGBfT7nBMPQVbr7tc6THzKMNoXow1tdWT0
KJr6ZqKjY65m8MGHrtO7wsFKwh1F9C3NmNyDffzi3v/fKsypETpu2EI9iD9VIym5
ewd2IFUpDbkXP5UlS88QvlBN3x+iqqSqNf897bMGvR9I1gH//uiRuxlwuAlRGDEJ
CEBycc4FTdoez9XPj36UvU2/TJ72jJ4o/BLGnvcyh8zEV/DlZ7B71d8e4iaGlWBd
fS13IBNKtYNpaSiK8EUtLRp069QElyv/HocqBQP6K0bmRwU0topSlQMLkjPCdIFm
cTPJ9WjyXR3JIlPyLZRQHBZQBgCJYuJ8kDU4UIWR9umJqdZBNP5uVtciXQWbjfZj
B0HHOOCuaTrKNCf0kY6eCHy1zXbTmJpis2/g/VZUsy8nVVIuYVWApHJk2nKL2q4d
TCDsyJ5NXBp8F5blYkZ9pa8BaHr2Y4Dxujv8C0Qq0hhQxdzBRMblybwKrzNaX5dr
Zh2dN7h0GK07FM0IynncKZ6v3PQwPkAoSQnyWYTtSOfYsO/wrFgaBNlaXnaFhP4L
5QKB6j4xCEYpjUC3fd/BVfo5M5w5+Rjz+7tiUKIUEsHBOTbo4PW0AR6ye6JYLV+5
7iJNyicYlBRVp6huccEkVQ136Qjk2HNOHrYkppPoFjnqsNXotm5kfNz5pg/DGEm0
PJCOCOBBld+jVeEmRLiDOw1awivpbk8MH3j6siMpyOUwQSm8Ic8VCBHZURsT1iCI
uFXzCmJpJ7DaC+jhiqtzCd39TvBU/Ka8BJyq0eYiXH2RAbZVqU2VlLjEYElRI7NS
Cc1xFORiL9ijW85YNd4J7glymfcsSA/88KMCnXr5yLqhLfqm+IA5IbeuZDclnD5L
dyPQGcphCamI2jUFF5a5WiS60bVYMCuul+iiIrdCVc4VYf0BC+XDcWmawSYYU3hw
GeSFATs2NsJTcOi1tnJwP0gowg0taJjhEHLKx/2NimFYmT/gSiMRByAxKXU2j1Ql
m0C66TN4AUmVWdT3ZCFiKtITCGuwCBq7gmYZLRGnlGFyLUHu1KIPhlinyBQQhG9v
Wt7AiIZ8+76Y4b4n+eD3+HxfcBXjZz/8aL56jwR4NJlGzFyxtqYy7NO/Ipj8ieiz
PsYD9aDq24KEOD94lTAEd5sBLTzL7lDQkLhdSwSnGgqPZ9M5kGKmX+V0tJBpwm1K
0p7NVBSX6LVNdRjhmvoOk8LjvBkzoXnYT1ANPGv8h2wCgpOn9jTcMOBOn/iVqcRS
sUPvlGAITziOL54IHOVPWLHtz7hD1x97+R/tBR67j6i0/nruQMoxJPjhbqrKG6fr
0U3HecCOtIGKLWr4NZOW9RfUV86MkSv5COuk76na/lCUIXSCzYYHgVr7Pa+o6+U6
ewBeVQRoBYZIkxEE2co/WKrBr+6zuuMLIG1bL5ZjKSjIPrr72+2Na+PyVkPAM5UA
HPtWMrscNH16A5ogD7Rv0IBfKLMhc9uQ6DQxOQZno7PZ5FvSVfjqz/qR+rngV6HW
bpEgweb+KNg+WVkzeUmoMrSg8XH/2kcXKg/DAnYLD3VX0XFM9eFgLtZgQ1+vu6sB
NjfddslWVKpOW1BAD2ZmSbkmWmbtz8tfbTF3zqYOgB/IBf9fccwivme83N8TTxBB
Pars0QkCep3SiojIuBOk6G3xy7Z4/Tm+jBMA5HvNXZZq2LfvOcqk1RzkMGf1nlec
9CLUnixOes63qj2I1jaJJySsRe1wD66dtiJ7TqBgLbWArr5Lnup6fiGQxDw02VJ1
4iwI3Ht90ZnqtNsy6AzPrZlvi+4DG6VuMllT32Ue7ht8pvwVk+x83jIRNYLlvQnr
ZPPl8slJEStCoeZ6+9jUV/u0u3gIbjreSAIYzmu3h45RJ/5kmPKu3qEfyPzjYSYj
OBWuqzFzHTGcd9HDxdpC8Kf5xkRgQ1Akd3jzFJiEy6I+mIVFbWORYPqRgBmKd5Qy
87wap3dL5+EXW5lAb/NYf7RHakcPyOuThlsOUx+jGXp0tjafAAWXgcue+49pvkOH
6PruWUZpIl9/h964/F399Nsv87ZK8QsRJTjYWf+w7aH7pLJaSgKfXQ4pst56rBlA
fxWrgFMQ/gel50sPEanMDrUDzafVm3xMxSsRWqH25/hNZaL3+4rkcAuRDv23RB+r
0EkbIagQAFM7hPcr6yfLD+b+CXNRkrmTgXigUdK6OUnleI6sxhf1Oh+t+1i2QLvt
usaOouBgiQ58HU7brBjEdcbrqSE8e2r9+7BrshKJqGuOa1bX29pFTlznY1KxmK08
TqZuXmze42PGNt8ZTjq7j+uEjDmGRyJaZZVvjAuJXKGm1yEKWSWrs+TKENWLL99E
64xIUXciPdR0eKoLW/xyfXTOfoFyP4MNLoy64tBJIR6UJkjr17wpYKpAbcjv+eG7
+BE0owcvSMuxJkYc54ML0ZRLhzSyhMf6UipnCBS49rKEHMU5ULznMeKk/KvOl4jp
nYGNuKe1ToM4VK8pWzm4LJZx7LZg6Cim/JSwwm51ClG1Q3UU1gH7PqXVNO6duEBH
CYqNuWuAWxUS+QmRJOjkRNPmqdkzo7i40vgrm3gOQuH1PaH6ksC5kjihRY5FJtMF
TGTx3dgQKrQvS1mynFSYUUWNvpAZNJVxls2VVn+KFB23vXkmPdiLegWl42ny1568
9+AuyXf2r4KIrThytNbTlIr+oXJgd2OF5EWB5vWirqvbbaGmZgLyWeFNXcR1Gws+
NHrkBi0WNvlE0fXTMc1nCWvcPflALLl/t+I6X48YS7QERCYrj7V9p+vAGul4xldc
3uf48Mile2WPqcKfvGVA+4/PyhisW+j/+/C07JovazsTHDx/DQCWuWa0s08vgTs/
4d6rWdnKOxYuAmREkj/kFwiLsBbk3S6n9r9d4ImlqPEErzktqsf0urjzvJjMmhcV
PRg7v2ak32gflfU54E+xtwTFBK+EMMqlcYGp7B8xRX80Zxrh2IWDN35JqGXtTUoU
Q+vIZ5CELGWm25U9OtZJz+8s1mAWnjk4M7/RM7gVi+oN89eTcnZfaLkj3fq6+/9T
l04UVFFkAYA0yxW2JFqHM9U2KcMGBRH4RAdGVg2W1mzH+M/zVr4o4msNBKYEqDri
YwZpccRWdQcCKUk4aX6fRHhcvs/GY7kLKUtvcS5vucqNbr3jRmEjCt/Y9rZAjMpa
5cMYLsftrqcZvvYavZO3MB/R679kfv+jQvgdjaibFkfGRuwQdkvDgt+5rhM5Y/bW
nI7Wvne+CaWVNmTKtDEZzTnVS+BLF1o2H1Ew9VH6050t/703StWbT+ycjdpsUhhc
3pGWkV574JlrDrzMFcfbh0Kq1YThz+2Z0AumSdqWW2QHAv+Yz11rWhSQ+tlzdxjP
MkQ/9Ny7UmuDIvO60bKO16EJsPW7hRTPUAMbqMpn+LNhxAJRFgXI5pCaWfFXJOrC
GrOR8Fk6BuZYDW3+jQ+pk4kDCVIxzzVizZMYyuo7/O4PJdVP8k8LrJj46aU2E1EP
zvo0vCOiob6wectt3gocwIM5ZZR4NHiqQWP0LcJ9peDqP8d6ySSi9aAR2/Kq1L7B
r/dlChJoW4k6MQECx/8J6zd3BHi5yd/Sw3Md/U8RoRY+bgfSXnx8bK41pDhbA0qJ
Tfxra4wYNdUaBs1NzUDA+KNz8o7vzP08AuY8G4z17giMh/hfHoFt8A7Q4f10juOk
EuX7UJybQ7RuDgYhgCYBp1XXzQmZ9qxPI0PgQGAa/X6xq73J2i4v2kTR8FnxMQF0
mpgcg/UP78MLWc6cfLdS1rpYl3oWQLtd3+cBrvJ3mZAAlSRbU9o7fAM4OkqQdDe8
Pm2ziHjq122yHSEkXD8LAg==
`protect END_PROTECTED
