`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJFQKcHxS5NZvR5V8OAFE8ejgcrJhEVleaQzBMI+c0ZbiwpFZzidiYsZ1K0Wg4mu
HwlstxzEPvXz4+BuiAU76s2m9Tw5gW2YZFyQIqyAN8jmxvHrIMi60BZNQupUQj78
zojQaOKvALWyye8tTkktuN/NknIdXO1BBpf25+IVt8k5FXtr/jb963C+Liytmk4A
2YvIDU2XGwo3xk0M/edaTE8v6VFRyir+tH8RNbzwWCwl3K2iIPvWfb/ecvOHzSA1
KadFk8cZHAl6GGl+ahDeW8KU3D3cxG4RwFP2F612dzqHtqqhCqIYINwsYUnOkzyd
yCoRYzlSMuH9/vtPpn6gdMaKBPPJuUi3UB6f3VKej96X6dJq0tv/ZZzlldip+G1q
O2OFeF0+nQPQjEvpZEmpXn2wqEUEzzBLvU2X5Byl4yA=
`protect END_PROTECTED
