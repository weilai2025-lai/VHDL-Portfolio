`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MUp+SPu9bhpz6fBKN3Z+jcVjL/EVf9zxGqiX975IznvTmNjyaelfPM2BXDRJadBb
o8fQtuuuuQ2umcppkoHdZfng1srd4GT++LynUaK4ta2Ng259jVBMVxptvhO2NoJI
Hhl3Gxn47hQ/nwMK35BkA1Xn1xEcDvfQ3Nzepl7bmQS1LVs1e0El6Ctdx4T6J39e
8oCtvmAM6xN4SucxZ+GxSvskoYi+qDnqDcV2JsPOCmGaZ6+Yb6ae3xOljBuWBX7g
vWKpypcx0nfeAszqte/a7+ogq0yOouGWq/v3Zbd7Q37FHrRmH1hMP0E5FRWIiZqV
RbAyxIZTtu9GLskrO/pq2V4c61dSOR0JdZW6Gs8uQKM42WrtLsm8D2EvANmGh+qO
vTiMDdEQL4s2P2NjpyyhI6hPpTp0jbLU4DhyE67M3r8q5aHr5YFcA4SZlXWrXr17
Zm0EhdhfZ8w0+nmYdCG2Ew+2uO7i6H0lK1pD7G2IjkQGdI5WFvsvruALYNKB8qAu
ZQiw78YTCeyACmxzwEPbq49G5sjnQMN5PzJmn7icRu+/kfEmOBKG9UjOZM2ueuFn
FxkVlD3pIhmSSkz5lyv7iAbpxkyKzmU0CkfZ/bR3uQvgNReD0ftrx8Zu6zBpJDTP
KDM/trGhN/ZFO0PyjoPqWYeyzrRcsMgpfhe90//k/woU1SoECaEfQI4Dn0rVI0lQ
on/hub9EKhmvatWywQr6DjXdOJZlxD3fqq02/VIfe9/A2soznM2GrrQvZqDaNlS9
sj+X3U1e5wdKrVnuFoeZBxihaSIPQW9NyqEMwZIA01b8fzynGsIQYUojAbEFdnyG
CfCU/dNPUY/sgjVww+Ktdw7DdVbL67qeGChrB7XpTRWyJqjvBmijJcQC7rPUyZkW
dtg0+R/4GvWle3MRcYpIImWw8A9VNos9DpPlXsFffZKoYgCKjz3CjSBELSjZkt0u
Q1chDpHuJkReTULDXOknfK5//Pnwvia6WB+/xR+/yWBQTh6WexJOyrxFhxURuBdS
YIKsKzx+/g+u2myiWBDjUs8wGGJm+NGrBIe8csUCl1hClm6ypD0UsMfzOW5lwX7c
`protect END_PROTECTED
