`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ImmkthiVQDeyWLqVbQudoF/jxmDuCM54Tjbn57tllTGJI3Aa64ASvIOwmi+vT2aF
nyATkcpTIlmCkTJj1Lh6iwPeKAy4xxrdNJFFJgYAG9F43Q6EhKipR2VteKtM12W7
lhbMHZZhlH9cxU0cQmRhxvYIqT/8KY9D8WpmTJ1+gkPdmIgeTZ8Oz2kf+BwAJYBE
+7TrpKvg6fE6rfkfCs5GdH3IMiwGfjL3Ghrt+QFQJWWWZWuVtufxPJ2tiWdmBdYy
KcYXjTEjRgpKbA1VpLXAYIuqpaGYTm1CwbNjc32hAgQxE4dXqBVZtdcr/p+7obzp
x6DSRCJSlY9ty+zXqOaPSZRCQEMT9J491VcVoOtrrSNSITFOKNjXRH9qIFepoYcW
b+sMrfNnerNwwJfu9Yh23hCsjU55tFTPQRfevkUaM03aXzAnZtcQJ+V759Cx0xcu
e95tQvBqLg4WuKPkKcmCjq/Lwps/B4iR7Ewa3OD7WsuUEY6X6kCZmyatW/M1NH+q
VR8PSE7aqCMXj7tkDqAhsfC/SwswuVlXtr7Gvcr+rlIkJ7cnewdxLxCVkGTo5zrG
wNxW78OoO9Yaud45mPlEWeeJXgkFI0ciSeA0j7lQNva2RVOLjReJWeXkaediVIhL
s8IuMZgOBHFBMgmrEfMD+GiIl+f6F2h9HpjFb/A0XXaRQdegZEZnaxI5KMI5lX2g
uvHukovFUU/5xoQ6Ooc4n+pCHLlatnCrNZfowZ1+Hh+Fk3+3BkUFsgPvZo8gMjis
dHq3ocUpnaIca3kMzqbAgvsyxwe123AnOqS6Q2WD4KTJqPQGPsglF82uDCTm1ump
6mrLxYoMyzlq1xXBI8G7aZQtAP7aA0wH7hOue18rH2hfAQaTwq+f/WHIvKXFcHxx
wzyfUvGVM4YN5SJjr71GjpgAUUqQbxYbcSI2cvcjjl8AvYamaFcaeeF/0cB4Jo80
tLuTRawfe4Kv1x4PKookRqB0OIuIP89Wx+eWVc5LoJebWzfeUM8U1lvFzmWlqRNJ
ZFwpV0lyxP3Aqa8qhyHL8Jyjd3xn9CkQ8o7K293AvUlFKRpZEqOPk2QOfYtZmAFF
OttubflzH82OvdQhshddCAgcMp3HnT8X2mdVnmLFd7scWQH5BO19VTtItZQ/y+PY
UxVxdod9cYb+Wc2tfeWCZJCssYo7Si5ldD1Fy7BkF9vfrBkJnp2QUpPn9+grI8fi
sONgR35eaJhaLe6vB7aGIYs3u+BtJrg85zocxvnT2YYW7odQ3nwLQNbQryuzfOi4
E7MRvTz39odacZb2yrS1QjhuMoXr1UhgjlNBW+5NhJRIXP+FwjRGDNaIndwn4S/H
kTdeeT69dOWNMbXJb1sjwT0BseMn3RQHdKjssdiFAUJqTAnJ7xcQwlnDEx3rwVio
CUXBP1L+++tgb6w2MUl9zXrfJKwGBV4oyJwt+LhSKBsEZV9j0NMebxedaPHeXZNY
GQ6SV/3iVJ0OF5PR6s+3mGU59JWO8jhVaDHMcM1gTfUcaGkZADLYgN7ogoJHZVkt
u+vOvAEizOLc1vBv3iH/+/6OKvKhVcjm4TbuaDCJnE2QFjkuGkE3PWcmEEn6689Q
6ZhlYg4U4iWJ8IgU9q9Fy/gaa/JVpQ1ztGZL+8QA3Kxs5LOKplGzOn7gw9cK4K06
ZzHnk5lV2qWJxIeBR7OFSCudEVwFZiJq3cvnoPBV7oVhLGSEIDttDp2kFkiYznBQ
oc5K1vKUuNDr0vOR/8n3+hhQjqzjpB0BZUm260QQ/KH+y4McpXro8E3dyyfT5c5h
439FaDIFFrO5qSedTyG+vY3JKifCn6sZPcZZ7rDLI0sitWDFAq94wwYGJ4F3sGD/
b7aECdkHseRP7Uc89SoejCUrAUeFDjQdoRkIWDQ1bLXotHDR4pVav7zio99xPghX
lEDIDLvzEARfhxhtu+ZkCruF3IAJ3qW1eZTNfUTZupb/CoQPIRHWqVtgZ6Qfh4ii
9ODi8IHfhV9jtNAV/72rLx+U30O5gaXAY7b6lJKdp0dMi3JWz6F2n5QXyt1j0/YI
q1PqD8Kv5OA7ttDyvFodVMkqopvCQsWDag7lgRRqJOacyZy7SAU4J5mP8lf9YZu9
6IneJU9jGTCmSp6u5EKOmEc9+/DdBvg2v1B1PS8+crQgY8AVyLLZWJBTCYvQ49Ob
dFrobUwNCD0acGnUVZFauQIk/HGJ8oDzay/gB/h5WIb0SPXJsFx0lDQn4N/gjlSD
FnrkxRfAMcAlh48GvkBQJTB/LnzNTKciFx1ER9nsvZq74cJ89WZLF1M/IX//TtWH
G+nY5VVemiLznz2ny3TM6KzikZI+MkP4FwG2SY0X1mtjThTxs9O0uavuOXUv0yKI
VnqEDCCqdDDEpi6xn/zz5YjTlHkg6x9WNpeeMFU6MD+uAXDZBUfzr/n58peh6kBY
`protect END_PROTECTED
