`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nIkmuXZ6N8xrR6ZuWJQJXDlRGTQM0x9BqOUBPs7x7BVs+myP6xUbnqLji7vboiIj
ObmlPbU6vrh9e77OTukvYck2wPQpCL7p/Rv5+0FMPGmFiaklw525c1/mYdIJMp+h
xbHZ+NSkT3+idrnbEgZ6FdXDMfeh8g/EAfSK/crpW6qG6dQNGys2pEe2VxiEqnoW
cqEYqIj4hBjMKwlbxTxmk7mU8vCCbWtXat7YTzewDTbvbpTRrtWfahPk8RlpE5Fe
N47ZsDWXAAxfvCQrB7v+Wo3P7fVIacj2/JPBaw5BDqndnaVB4P7pZFFhbaafMpeI
DIwZQXmbxQZfX7x6Gk28d/9SIysANOPEiakdNbJuuGpQAKtarRPuNkPVd2G5EALv
+4tAvG+XCpAkMduBn0PB8pGXeMzhvF6KFtii98atiOFFfpk8pdhEIDk/DJ/L987p
+NZ5mmlQcOKUq09wReEY2+85yGrJdkrswf0nVWh4tLgKrb5y/LbyFm7M561ZBkm8
kKGfrIbSFJr/5tjyF+o3dRBEwZozbmYd/LWnN9zcIwR/jWs5OlnHcdL9tHxoGv2p
etaHBfEoty/P+3+8MVzd4LvK65CladvPpTRiv9JfQxe251kbwhIcu0Z+Cpa9Iu0m
W3fhkf2OGo8QjZ3Xo4nDT0fVG9W302H/7lEhMbGXNfZ7QH7fzVnQ1t1D8Cx7PAR1
vSWli6UNEqMo06F2tA9b21OquW7pqy1afIzl9mPVGFt5UbESWzhsTVO3O8IcDvDE
tN5w/rUIVHB/K1+gAJiPsOG+7M1LeU6Ha7ApUcuIw1HwkdgUnfJ8V1EAskQbezEO
UBTIyM5zebz82b5PA1vIue8TZnR3q6w44Dch0naNt816v9/DDd4niHxcRWwr87gJ
cnFLwxZmxvVF6fiHVhZEY0oi0e7kpGqGo+fdsZmMiguXgqlhcqGZ500fooKKrMkv
AeUjCBbsXzUeWKSVousXs/sZ84n5ArEw46n1M1NDRrCjDi8M4oqv4Omb5vf4wDpB
kFWz4ldCQOvbzTXodlQBm4S6rFCNFE+RpVgoKUr50L/ULcmarQ05CNA7imiIeXNp
+7q4bjyFUJB3Ld4IpW3cJuv/aYcddD9KrYsJEJ6f7hMWpE++nQ0Pr4vxjH2d/CVI
sqFa/D7n+CCqq9puLeFTpOdwrfLW8VKS5BOq+og2+wGQerxaPM7ayg5dEdZOh+fL
dZJ4RIXk6hFLQRgqAoujyYF5jYB3AktXv5UqzG1eM3gpdRlDIleOn7WhNVtt7BIY
wQTrTg1lyR/pra/TM89Zv5qYFLSC7DD897XpmHAc4Fp3++YGlSmr+fEWGZk3IvH2
ljO1d5z6XcJCNpS5KW4C/q0lmNSmhKvNS4eQhjN4xuYvh6yLghWDQoGViivfyin2
`protect END_PROTECTED
