`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/YotsOe8VQiCvfv8AKVHnZguh7Vxbo93hk8A8TIUcg0EuJ5VejLhrw30oYpAu6y
eLgPdeVxecnu2/M7UjEw0aYC28Zeg1LvHaLwvGV6Tsl/tl5e/gA1Ic0PXrBEI+WA
fgdwjrCutVmrBnQKfJazwLrZsT+7T6EEKcVEX274srIRacOWyk7161KH6qBX1dHf
PsY6qM8Zc0BUQMqO7JB4OCPXTxqKOkfdqyRlloCksIm1xXHMy4UmoyA24t5x48b8
KXTLChoWgCAjH5aLHACCQjpKxFtYiVCbXkZ4QVlBBRDYqhrbrM2+CjjVP7MLwqNv
W2v2cx15enJfA/N/cd5VYDiJtIafuVAzdppHikNBlGDiCnbAyBXFYlSVF9N8aWMN
uTPelV7XDU4lqJ74kSBqKGQipTpwEnK14xrg7AtNrj4W4weS4t4n+KapG+xPogNR
SYGHB01E14I5enZcp+qr1rVcxRvswbHybmY6kNoBTtLJ4NuiJaSPRIX+ca9OKujs
cbRnLP0h9LQ7kpc+UmYFOGsR8Eqt6Uftfj9J27D4z0IjOWNKxQ5+SFn8Ldw4I8u3
XQGgSUWnlOWckOeHsBfS8Ci74K15rz9Ep6F+BLd+ojaM2WrptLIv2vIiGZaXbJdz
79PPEr55WU5+WPUqPcWSWv/CYpDWHCGPmtUga2T4iji/pI/WgxI3RpLblpDdK6Nl
oc3N5/sCbdkSHnVXRCY8kN+pFyAvAZ4CiGd/5LR1Mp7EsOKKdk+OIOsMAvGrHFCW
ENdZWekbojx0gLVBeO+uFjtMR0eoOSBzvbQVKBSRg94Duf0QzvUvQ9oQS6s1b0dr
SrPdUpH2Y5UfkXwN5sGnyWHQGuJyMoYI/RKzD8MXNJdHAvSU0L5zE373kpZzVyEH
0rrFrg62YmMcf4TqBiZfbfQgeTaXqiPoS4CV3x0YcMdPEfWriyNQ5F5tGwzqn6nO
02GZ4QZnMXQGRJt3eOuS8ra/ea6VggkKRcahOnnjLa84Pj51qfnqpJiXT65E5D8G
zFoUH0acyXPPUfmgQ7wYGyXCCYAzoADtULPrmiRb0OrRFs6NyIcQTNdCZQ1mxQdI
rbY93qgs8CReCei7LyKRpI9GenOAyq5nE+go7KFGetq7opTEOkGLXnMrpFUZ4cuw
ueUsKwgjiwe5zV+VeCHVCuKWX1gd/8pV4lIO0T19R5v7ErAox8esrnxu8mvrbOS4
2SAhDbaTc+viJ7p4HtC9J8yKp6Fhobtsl0IrLH74BJoArE5ZjQp88vfjMj3QUVIA
0sqWt096C8BoBhNWJouTLC6Hg5p7dt2+RQm/+xLAX0Px1gSv0S/y2R9TFGd7Q3FL
qRuDZQSsYIOHTaLCxqCjJbWMWfS4uiRPIWgXvKDOy+s0uTDGOixSfOlIwzpfH9eP
4RQc5wM3N6E7O4KoSK9bXjfI+dtFfgLYp0xsM3UnajOw32QNfFbDCZH3V6SNJV/r
X7RLFKaFwsVyFnS5J1bl7WfSWBYPmpppJpK40/v8J/CHFw80PQlckVvVQKDSGBwb
6TOlZT6JyMffxFVp+vWFWQ09+eWnRmLhB5s1jy5NrmwruPqgXh86jEJ/oeOG2Bqz
LxRyqOQFu7+ZCLEjJCS3FIXs1MujIdffVJpswdeqcJEwTNcS9rSVDuNYqZ7Mrlmd
B7OyX+nrsk0D78LfKKWXUG8gyvtZbvVlr3CXX+llgILo/KMKLnHPSaIEPOp4r0G3
pGe+aRhEU88xISyDCbl5uCn/soVcV2AbDTENzYg4g8LQ3LEixlIteNaH/HcNhlH4
hAe28nvLIqODQWsmgja3EAV6EK395DJCP+AS9rdCQi6fN3XBWtoTOY5VH6cdJHH2
MbXj2eyHQJA4qyKRGmb9ifI1dWSjYA8Ex4BqvR8xFXg51AqaXyThwoXgDzChczSI
m4B5HAzby2jl3acK7Tn2n5fF5BzKiuNp/4QZG5JRQTmgo4V7y4iovxRDKvSD59sN
7zAF0aedAFUmmr/DZ46r2ozqty6Ju6PENp5jrkwecyHx23ihgE/Hq2IzuH2xIht4
4rOXm+6kgk5J+uqpEkWIza2vqZXRo6OlssdRkmi1MYeuAkqSXp8WLRc5AgSg74Nt
FOMlCDGwxXacg8RkiK44BJ9hGuZP4T0U3PuYBOx9re2pynPnXBaiNKh4h9RvYo1b
fn0R8+8ftx1a/GL7xWs9nJBDjiS7paNTxEyCzPggpG7SDRUsYXGjCD18nm8YYRTU
NDskqULIEUIa0JtrVNqXTpV0fMJmjvAduJAY4ML7E5HaYQppGNxFwqS4gHFMaIFr
KRnQpDR+sa8/xIXDZTsSofniDuNWW41TpDH2QZ+Ldo1FGmkILsjxiZi5+DxblYJm
/X2NgbFQ2mCdImq4cyU26ME+p4mnN3UboD9vdREatGLcZoqUySaeNbFvze94Wco1
A7UPOqD1u07luhng2Cvmu5UkMz2naumPpd20NzRd9de7J83Riw2bMWnbH/iTTEVK
3UbBsy6aNxTLIW4qfvd3MXaZigKLNaoPzdwuKX951noEV0hyjFUlmrWg0TnBpeAm
VfqAjOm4MAtvFINYdBM9RxVPyTL7gYG+Q/mrYvBehSTG99fYRe0kdhynkx0yYa0x
vD9HUUy8ZviOd1x/a7o2J+RFcpSLTXs6aPoPtZ96tf2YzjMuPYbP4ara0LozCcZC
R18dKPcGFK4vqsoK42fZdUBVMXZYDoFLDI7F/8FeFs6+nBH2/7si99CdyTyQ+wWR
sByxsNRMrAE2HfEYWpOsYLPfKdDW/0eTc3XWJ/YkWjphmrUBXiKRroEvIvkUrEbI
KP7I061GJysfBB86AV7i9POAt60Xqf/y9S+kIP4mfTW4SEAlmx2m0flcSGEeM6MU
jHQANJCyTVI19zPBe87YtijFX5vjS/EgU8jc9vpELpjbocB7j65clzLJJHHMZve3
0BnE8UJCoo5ANkAhas2CV9ZCOabodC3n20d4EvNXQ0jjsFHuEkKvauYwDciBWb/p
G+Pk5dbmtFUi8l6OQmAgKUVHn+T/uUOVEwEOKCuQKZ2agKIPicNZ1oKQ9UnYQMg3
3f7URKIAVhOMsjG/Dds7AO9CDmLlB0Vzib4sKMLnFwY2giwKPmJo9Rfyx46dRuVW
3pxoQPNbJFtPoyDCPONQoYTzGxUUH00ojpWaOHmwnIKUZWPfpk7OkovAqerD0xdE
s19O66jDw4hOovdqReu/kMu4A9H+3sZgYhrO6ws9UByD36dyyANuPqj+QR5RtqBq
wuMqKmp33xFQDERXCwFLZtvI6KaLjBzzJFTzLCHAeXnqkEK4PCj2SEPxOhqnGrHX
hu8EC2wznYBsrQJzm6CYfkcDTi9vluaanZ/uGr+Iugo/culsRpt5TwzKM47h3cDE
N/HA59RW20hc8HcLQvM2xL9KfeiDJojdH5ncDAjLgd+fkUU0olBBgnyPjkC9UvKF
w5gCbAh8cVOZFJihrZt7Ltlvy2yrG0j+vQeVMpgbkc5dfw2OI4dfKCymS1PwGUnb
2utks0K3DpO1QuBJVz94tLgGkK5STe9JFz3EofAuPP9LyreOcurgAKdw4ZtFWpmH
hTgKqzCIMJcONbdYRmtSNdEen01f9RX/m3686G1iqJsaSR9kRW58qbxD2U2nV9i3
RVRrmb8mUYRXi5AS/TyKBl4vFczOGyfw7/gCkqhzO1ulK+3oSRBlYTXvuCJIXoNB
qiOE/jPQLqTBWS0wMQxi0PYZ98K5UkF4/hLkAX8hhirysMRZujXiRBirsD/4lH6V
Yg8pZCquzRfhmqXhfMpf86Q9DUk0rR+ax+xW0hDiAMM2Ix7hL5NuCGySMO5fohYX
sgZiFFgWUctQ9FqiELWLMe+o0Fg4Y4+IWTL8CaB0fB0wuEMs8vExsZMD5BADgFxl
r+AUfT7i2hZaVgctCEwcnhPEEOJ8yBcx98thRQiho0rlyms8jeZQ/voB+BbqDX0k
2LrdIYEYDR1A5i9S4r761URRWv5KEdZJIfl/1A1mb3VkeouyFq6T15AM/kboLdCD
yexGn7pu70d0C+jW2JhAkBg+UlgmBbO/iLfSExPeKYS31NxYjxnzIHe1tU1WwNh9
jpc9SeQjPCKxHyWCa1fUMbJC3GnBzr/1LzJeNjQ8Put9z2HVZ3YZHBXjTZnjgbh3
78P1rQadrDz9V3KHprNyVgAetzefV0sJwUOcZAT45NlFlGSuW6R2y1YobyDq+XeT
DunOWkpeqvw94zoLdGcQM44fmeWy+QJF6jeqXoErnEsJLr/+7l8+sL68Hy1XUDOQ
VvjCwKkYkcemIoL75Ih7cE/sMCsJCS91XvCYf24hC9GDghKnGA+LAXcUvAmrRERG
Bimb3ZFPo5RUNeR/5pe59VfLcIGr27tAm4P+k7t2GH7bpJPebFdSzhsyqVfXbMsN
Goi0yp4foy8xwakVmlQoYMpTS/VDjVxHcQXhLOlhcRrn62di1Zi7uw82kXr2ocqS
wlrgSFy3cGwlWQxW2xz7GmS7F7qUIy2wA9u3mYnlEympn2P6lhfflXrfwXNzoRYs
UpsM1TDY7rV+0rgLU7C2lMtfn+lxGXdp7nlWJohY6P5M97xrh7u3KxlF0Dl8oU/8
zM5SKEalBgOF4Hj/DpzVA4jASq/mBBZ7y2PcKOG6Cy3rlxxt0men7QPSxispSjk+
DLkim1xh3VL9fP/IM9s7GGPrjjXV6/qIDaoPycX09WbMOxgeeqRZNaeRFmvkOZIJ
Z/nGhCvyrV86KuhM6q/+MLSY/CQmV1hKDzkQPM2gYDLb/j2SKPg7ZUJKXGbHRiQO
Tdk1jbB+FO5cCoKUNUMqmAydYFhiCRznRoajxL8c/cvS+CZhGccZmvFvODjyyKjk
fs8RDMNQNG8UQEIYJqarix5UO0KQsUGKyx5AcqRk/altCU1B+CrJ+UV5hi8e6Q28
s1tAVrySm4AJH5KoUDaV25QLaBXX/UDZGaLcosJ1ZkXOyjtHoQc9dvKfbGYm2IB8
IkIi54W7DLF6vJxplF57hFnjSMY6EpUFF+vv7uLURcq+mYcimsejTJVoIAjaqhXT
hyw3cyfTBN1Hy1SLI4HWiLc6TekMXnPPfn69dx4F3TnytmFCsaCWgPgk5m/ia50D
kSAi9gxFwVlVdo8Vnh6PF8TyhHbFAB9LUkl87qaj7hoxGhGyFIBTtUMM1VVNTS+K
0HiQQKhB4zmewZgo/rN7ts7v+MfPglstqzJUiAM3Hvkwy2wuNOMvRPKZLfdsHdlP
gilt3sDDifuGnJ5DcVcdGJkPRh7DbsZ4twnvYNdnyMAkq2975PJxkL5zcqFRLaS9
aK050Gp325gD+XOnkEZpMnXTmxHD81NqEt92BrDTGF1LFz1440xcPCYbOdZ+bx5Q
j27W2Xw5u+MLbQnk3kk/OwhHNtuXe3TaBY30EOlJbKyRwHkDt0j1JVkNO7XlR/Nv
rX8Wn+8J5fFDqvvM4ArYQqfBmMpk+wuq/Fjgqn4Q7m1cT2YEj6e0P2TiEHOo4wGU
+rEpDxtvbHX02RFiCiI1fJAzQJQDcGlQ9ueX2d4o/HvgX7AcokW0zsZREKghO1rS
urUDhC+jUH5IBnSiVS+X75whSP1FDZz28/14TE8PiGV7PI8u3vcESpvH6h+t8ule
5ztE5vGDL042zsNL0ddcKSjhVH5HIe+lvTqWdoQjtUzk/1KZuE7RN0TJMXiRFC5M
cpiXllMQ8EbBIAD38M5hfE1nuTRZjyFXW5MSV6AnBT8Ev1NVfxKrzsmVErQVVV1E
d2vCFBcMZTMoU5wklTohAPJxGXGfdQjl8aS0dghjOcPBNGoZ+mjcTwh59omFmN2J
rG95e+Da6NFo4XyHH/tPaa5flqBRosa8c4Nn56P99g2MTJpPzUWsqLJDJaBVKZ9S
nIjjdosX+z8M1/v5vpWbNy0LW6GbaiIRhAaOXdlTYKX6z2uGiZVbL4mb7saWTHJT
QuIuH9A7o2GSXi+pv85UTLhUIbtVvyAldMc/Hrd0Mz6iitGZFBZNc0IHBIakHTXw
egUpzAQmDOByDSiVVI8jc/iy1r1wSDSOASG4dqNy5GO2wcg7B/CTTnZRtBR6p5cp
ATaPS8AtCMg0er4X/8ac5SGRnSaQNnpEmRA0q4Y6QLr1kcsu9/KpegC8tkjGVI2F
GSmC8H+CBgY0dXxPsJQGU+PFAcLjj5uUsMKbGrZJk+Y7hlnWPDZF9m+/E45XbrSW
1vY7or6FCTB82hUhJ6S8qgd+2l0nNWVMRCqwlxhDY9nVIumgP4iJzSYHMlpFzrbx
OMSS3SAXBBWDbGMakys+uT8ZzZZ/Y1TF0uOJZoyd2mGJFmPj25k/en95Pz/jtQWU
aCq7/nBOeqVQFF3PYw9sRCKRCvbAbyL2II6LuvNVFENc1kMAMz8vsB+bSrG5HcJs
IyylfXNfsyPtcPWgXxXf9bsHen3k3U2LuNs9c2I9lHxGdkf3K2ze0WQTXHVDDbu0
IOON2rboOapTne+pqOOOGfI1JVHg/+FBi5wvv5gxATqr/U5QdCGq8LfuX9D/xHpw
b2ya/bHxVg0Tj9n2SpnpZgUPIuJydg//MkT7uyPMzbX08bks618zm/mWXsIxrMja
W6PwSqCvNfaqe97NYs/GrrqFpoF0Z6/+ulSPLBlZgYt+BUCXQ7JadYQktnSO9A5R
G1tP0XzqS0wH99vP6Nhvjs3uO2D/VqSObqqUrFibXBbpCR/5bh+jZS5SBdAzg4+O
aaOmjOfvFlx49DeP3DdxC9QBvnHLRMs/4ClbAb2hzghRkLl5RrAJy2JExyNUNuI0
YAjv+URVadfWGdfNVjsSe3owIDcMddvmjGEhT/IN2CljtmLWcD2Y6SO0SAJ5O164
`protect END_PROTECTED
