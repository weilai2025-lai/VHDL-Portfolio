`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukS0mBgiaHc82irvxhRHknlx247uX5DpdfZsMLbHvnHp/BXW4mgbk8A1db/9w9mK
I4fq9KApaotHT1cI9omwhs9/yPYnbwVBAQ/dgMFfRXpyahGNX+Tm9Z8BNi4zApCA
t9ZRZ0lxsp9CUtpVbw2Q/WItkO2VW7XUJD9DYAQSBBaiusnC2f2Q2PpBoza7yf6R
y7NqOVU3bOn0bgnR1rsIoxu490NBvQcyICVGCf3FYdIgseoTWNrx7qA1ik4V526o
rUl1TV2yfbgRlHoCGxG1aT1mFpPGUX9Ivk5+wNv675wNM1BYqnEpzGtAWTFh4JQu
6Rfbv1silxtVSANC1KpfLGU4cxr8UT2X0iDIbooB4pSAf4+Blu3Ph60pWUsGZQRP
ysz0ZBU89oaAN/x5jK38z5wSbR1Im3JNe9gZ2lerpyiWgJR5T6XNHc1o35beSwgB
n8pBVekaCaIli3h6Wc8MY8XCgim5Hx7XFQcsgoIx5g0aYB13qGf0LYNqLIialKMQ
Y8G0yCoc+RWWHTN8V4XLrwdO7HiNYPauBUJHh7t+D4ozFP1VzmVx9N3PhaIynbMH
wk8Vh6826ZrTcnff4wxXE14KpsfEx8moTWJTxu6TV1raJ0QrMVl7KiTiHLHybv2I
yO6QeqQZmMZ58RD9unrEiV16hNHpZZ18sH8FYi2QDd051G6wMfX12Wa+1++Xv1Z1
joirtN9qTvxJzSVH8iZpE/b3XOrH3iBSxtBAboJstMm9PXB8/J96A9gpLw4UVA32
6cF+pK7CmIzQAQjFn5tiKspvizKf+R4SqAlt2TR8mnjomd3kSVt6Ro6LCi1NXPQ3
hGRQJ6M1/LgY3nTucyi/Rb9azqyRS749Repu+hoKBTR7SPC7tBU1o5nLes73ZJ/P
wwNE6Hnh29tEI8mtmbORxoMe01oN85gLrwRhVkvBC3268DpHZxp5qBJUzGteU/Hr
xAZRZDIWLkEDLKw3OuwIw57nuWrC2mahlp+2kSnFeqZ9j/F/zqoY15EjgnYRtzAd
ghPIbCyio/knLFuB5iEtvh4dpJ1cdfdK5H/VTXtqsW6pIol3WmiFW5z8w6XtMWbc
B6UmOpT9UDLIU2SDWPUWjb2MbSkzy3UQA7k2ZdVIt8Q9ju+efqm6aiBGT3XIQWS2
c4gLc/QiI01I8wrQhgpjv5L0ewswTqoBADXI6eTNPV9VxovZVgmaLyktnAhL1U6h
wlGrzJVbBP96Uvow/fWTnXchxrzEj4nEAPxA2aLFMaFFlSr7PP+5kPIx7Dayv1Ib
WlcBJ1WR9U3RNqIpjFoZspzJWL8+3rnHIj0RH/N5e2kwWI9Pa1MimUnVrEVGqw7g
aWGrIxvYkoanJmkNPYXFvtD3a/dFQyG6K0B/vK9w/0X/Fb932ilsWjP+rUZDBsnq
tD1hE3gr+KthiehJnNVf+YUUXELx5q4HkWexFkp9EjdqM/vBCs243Vx9qQqWWAmg
rGM2nZuWGlTpePqfhG2tlh8EOYe1CDES19RMQT/Qx2pAfH5Igkb9sFPkXClAFASA
tLKlm5jHM6nnQuqy1aGJl8uu+fOa+b/hgQfv0jV67DV1Z4tk7JR/z4wmLBMNp6UJ
m6h2QJ7FEDKhikucvDj2K9mXBGKkSu55cYVhHtwLcuuddE5LmGmLenXnyfhRkAPV
S3NyfZaHq6pP6t1NnMYdJ229lg2+oI7JcvHghnRhTSdOelFG8VG3SAIh9j6jMuv9
DIf2yRPYLnglB/MhTwGPPxOzwTfY39MbAaynpiWIzESmIJYzyfvt0n8+3Kday8Fq
dmWTjjtdD85vsevby/1ih20Y8hdrMtmPqq464K/1hnY4ywewNKjVz7R8lPTktrP4
W99eKlUMX18K+o1miS66aoCNkaRP9YQEDOp2ZVpRcC51vhzGs9/cr1nwAhsEt7AP
PVS8XONZacS4sGzYmqsRExGdlRqhBEIlH8VewApL/Kz64hgezUa1n+8tbRGmRJVQ
9q/vOzx1s39nkBB0SqQ1puK69n6IFDXZW/unK+0IQbRUaGbRNdyMT4wNs4spFlTH
Nv9nSHCu73aFbKMFbHCU6Ll8pwoQafQlYjZnz5qvP58Ly0LuKz1EbYaKrMo9XtL6
BGC0BhW0QOnHEkoeOGz5uhKzkIHLjuKBv6ANqZzKf503usZ1MJw9AWsDKg27RWnz
dMmIA2Zvm9zHxgPOovr0ojqp/Q2gZ1E+lCq6zo1vIcT71h0U9+HVi+J5nQG+PgnG
VPk/vt/D5XLjxGVMaxeCDMHNzatPReZXlap8Uq1j/QDk04ElSkn8JRWC6Ho6tAq3
31/onTrkJD+RcOUArpAXZlDY4lu7CbThZ06duomVVQeJEUqCkbpVbqa7xiCMioB6
jPCx8PrGqtjAWbhVkyxMt9uTHTgmO8se9iR64/+50FE8zi2n/tf7TvToSvXgSYOO
rThhgsCbYMUp88eGgZdKA9YgbNCIKxuzZnA0pPxC1++lsuocRkS+RCoV44HOczMq
Wa1h0+uf8s22BFtNoJ5Y00nxFzCcuQNtxOblG3zSnNRNsf3gWWlH4TVmdd759Czm
S29m/kMfI+yWtMVpINa0ITkZPWEFxXgfxEXm6t5XcfY9H+YxETTR9x3n0CBubc2j
Tr14jd5ahh0+kNynXpjwt1fRUqinkHyj0cAjXa3rl+2T8yusSHUvm54FuVyBwksD
0w+tWL8UkFFgj+rqwGRVNarXyxkHRyXmjzl96Sab1cGU66e6kro7WIHxqzKkxfB/
aEU2ORy3y7HsfK/HuwCHE/scKVZ6B85Qch2SfZXDZ3IjBbt4m2TP6t3lfgeoEp71
J+1+msJWiE3goWRfDyPBOBobUlVghVeVfnNEOklF5L8UTYCg1auh//y8huzJqO8+
OtIm43Zpt01Zrvb89CeS/aqNGCh13cxV0HBKTu+VHxv1pqixAyzWzeoTo8u29/8Z
NmexGoFddl4oc6jPwNRY/J4Y1rtg6d2S2b7D94jPbsuwn1KV7CM+rtOQHIyuOTQX
U1TkNJ/Ob34am6eb7JhmyyrNcI2Zj40korTM1M/JR5fA3Eik8Q9UtzaUahSat/CC
CDbs8Hz21C25Q75Ln2VYs3A5QonVZPquqJzYBKrZFkGZQ/czxsr5hT02n6jpZaTL
xtZWLc5FCLuKMX3hPkJjyvQTlrfyq+1/T+rbM1yKIrIb0xZdPDE2TmoSZ2wVuvDb
M6pmy8iLycPhWwSlyFj+hD6v+kIS7Ixtz5JxdcQUDmnbBCAYlkkFMnY7Ikh/wi4N
SEd3P6TlVVkaDATz/8sY9JoL/T5AP1vFM8OSvoupNc6akoH/wH/c8lzqxD1T50WT
2EOlM1f4bJ1uahxAT0IBQCJDcWpfZgHGdQT/ew7eMG3Lcu8sFx1sKX24eotBM5ab
+H/aY2XDjqPOSRk9FxRMUNAJfAaXauGfgRkjTBnqKTEsrON8dQf9Oei/Ynn2cEh/
s51xOikmhYqJL+dYv/BetZnAPGGmf5c0ulpHBMyE67yET8OBaVrR54loqwa9PqhH
cLSTXZ6GukSwoumQnm1lk+Xxaadjije/6dlUrNU1JEHsokp2mA56NoaYKHXoUWbh
Q7m0t6i7l6Asc47Pf0c3ne15bpp2cnpKT5N0tXjoeCHZ0L3/R+94JI5O7yImwsgL
SVBsecoTAD2hxoykzfMsTPbe1mdoc7Xi0GLnkAIV5z9K+CuB1DeSzR0S/oBAlIjo
Du5ZNyI0gzB9neQcj8waWBu0Eicr7rb8cR8PO9UX6idUm62sYFmlKXokGQxoAZlF
XJFpu+/m+2Cq4r/XWKFicMKiFEIJPthzNLtXIIurwfLOsvKiKdsnY3GCZ4Lkhibk
daw0UVsiih//UB/yE2kwOObD8ES9QhmYe1YA6/2armagCXUCzaWTAEeJSn/our1h
Bs+gj6I8+4LVsnPRUiEvUb+QxDFTdnOqJWWo3Oayfr1Xijgcll1wir5Z8coe9l80
FRazRbcUrWnJHARzE1YJd88e/VbuY/7cz4J1E0ZybNo6lq6fP2yFGzdyEleBEXph
Eh+oFgILPwlQuWHdjpA9JZ9k2Y5DmR+ceikhxH7K+9pDuoi0N3dqu0RM1XoBZ3IL
qOzt82sjPTXj2B2UPbNNTDysno3kqtJaiWmrvotNCF1lU77yKvpUw3vzokj3b8dC
9ZKL/GZYQKnoQhJS3I0gy/jsAg/qNsUzZUcVwXqIT9IcsHLKcjaEm4HVg4O/JFgm
fVhPmmntvIu1yvkX2iWYg8OWGgCt9qekgGJsp5h/RD0EzNBLczVLPHhhm/Fxus98
LUkpm+80Rat7VJxGGsJnJm8dwKjlBWUrMweUdesU01IH48pd+I/K+x2DiJ5K/nfB
9tyme00Vh8mYGmf/87MTm5FGE9bR19aW1PfVIRvb3iPr0N6unR5YobRBPFUBmBq4
la4b3H+fYDSF6qJ4FDfh0y3i5K+d0p6AHtVwQTLSmdOCPHFR6Fzk56rK68ZUlFCG
HL/AYOTfMtorEpvwyp1DZp/992KDXBabiM4GjYMgGnj+0pBw69k0BvEm7KV+hd9+
2DfK9HLJkM0NAuO7Pt2e8T4+jAsS5OLicWiiWip1QRWMUG2why7BudUPVB5dT2J2
KRBx289YgfXmAjt4I0lsePPVg0/Xzjn1dQM+nW4LfAS69fa+k/Zk9VOw0e0R4FI4
JO35r5wDdZNuZVmKRC79r4nEkMaVlYwinirxJpJ+yWxMroIpYU/0D2bFPl8QjrRf
Wdn/nsTAU454ENr2Me+HlTq/qkqRqc8HaUv5cWPfN4xucJHuhv58n+MSO2M7ezj7
N15T6cr8FB5BA60OBjUjj7u4w2u5MLEiVpeBiD77Q8LjcXOtpr2grX9u4/KokT1L
Bkv+yckKVO05vEmXwVhcC6eacFZVuaaPSK/ywYLTUo/PA5FAZHdm7RjLwQBvwdPv
Y+zW0dnbdH2zJzyN7Bj61jCFebOHurQfhJJQmOwbF6ioFaR31/VbKTR77rd/tIzG
yfKUJAWn+MXnAvbxCI8i1R2MIWeRZ3lWUA4gr3FmsIVTCjvWC9VPzrYPDrt+NGYp
Iu0iMQpzg5UbJDFcprBPOTzl1F74xPgQ0pH+PhF7B/Dtx4+l0DbOSRAT9xAKJeiZ
QAMNYhLumLdBvmpk1XtKuzKibLUVaJLcYxE1lsCLXV/i/sV1oW+i4Tw6Pr0D5xDY
M3oLKOlMCSg7qN9P2jyYt72/LGNR3CUps59BaDnkaNb1XdPiNTt68O+57XYHJWT0
st+zLOZFVC9tuR7h2o+88tbsiLaJYZzZk4AsGy/DVugBY4iiQ/lU8LzbeQnxSB6q
gZwhHbhARMsjiV2KbTMvahbFIV4eX/v3DGv8m75YS5mbD2jOK6y+UFOHwUWUCV7L
ffBJ2iXKvP9h1vehMfoSY1a6BIoUyG/lph60A7op98yI1NGE8oVSg5iF+niT4/Bo
NZn0IE6ss/LfbOEZjTWQE1zfOxSaMq2A5qso0nBGiXFK6iz6bU+uQJCXW2hTis0T
rgt236Pht6e8ex22RLwqvVTekAC3+yWHQz65Zf3onN+u9X1USOnNpZDcgOodgyJ5
7x1+RSIHWTJ9Wz7caC0RKIT8DRygaI36+n7ihUPxvHDBz+KKQ0jtC5/DkjJ0eQjx
UwPJe4YwMeefjVlNW/cBRWoO4wWdd8vKNMXF/SnJAyrKxldzycyMAKV5kPJF7SwX
Pt490hmpxFcpygIBdkhOw0/SxFjECDbEmZA6BGYpM9L1/uwQVKWLCTH9b3FuZ97s
zgW2XP1fqsvGD6O8WPsLCdOte0qhT2lHYogwEghhFgF7awHf6Ktyf4oHQH2q+B3s
tpXsn59jJXbdEuehEGiXfgmcPQ5LtuT5dK+Qeslxqg8=
`protect END_PROTECTED
