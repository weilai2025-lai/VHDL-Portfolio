`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJTKpOzljuKKvjSps+B+dQ5CVKNx8r7TcIZIAzhYuVelOsKZJMk7Kw4rECD8cdCd
AekhhsjK8FUKEEdaTcOGAiSFZ5hA0/AWrBaRVrhNXIAdMRHZz/+9Yi1LNJ1gBFcZ
2NVDG251eHjG2ZRslTgUcrpcla8ifMza5HQCupaBEEU0tXo5wmKZDaxlieC9SqNH
JNWJwJdSip+v10s8LvwvkeOGFwYdaRgxhxJyeylqqGCK72lBLqaeHjGsIqKvOX4E
1E+OLdcAoP6kMgjRmjCDlC6pBMLaujxkhU5lBSNzwQFwEk/ojOLjFjETw1utfxA4
QDxE1SbAYibIjTn7yrf+Nj75n/TQMnV8naZ97GUMCMdv+OAMw5bz8AYZi/1olVzC
skGJQ/HiBbk8k0w4tTmRI7AVt3jX0twDy8kjBmjOkr003tqoINhs2JhdrndDHY3N
Sf5XLW8rDXTWuyUQLGmbbFW9/XlQEjA/gAAC670pAhxqfxOkt8lStHMnsEEdeLex
JZS3NzhneOTGqw7gR0r37MVceBOKs0uw3+QPnl5Xsfls1WsOpMmRDv4zsbQDNJVh
K3svnd5hHsdOXUwUCzQaDsXzQlBvC4tqGcnesV2Tfi5NHGMmWG28pSZE7ITgUrmg
5vMCNRbUnSEQWDFraebrZ32flnlbfd1/NQRxDGUNFRdxmGD0+n/k+tMw+CXDWlH/
xpbnmwmc/y1oKRBYfSKfoPmBoEv7pa9nESMT9D6+wYFnXXnKBaixks6Qd8o9sP75
r0BDrpFaekmqVbRsLYUuTpIPPvFoylwjX9iAT3BBQOHEdIRMY1wqc3wqm5YTKYFO
w+yIB3xDAjFOS0O2WSzu7yeh7pBo4OSmRE0I0jpHdYMpzXGJt0MzPvSBDGFRaEOT
O+hD8m6unGNVc74DJgUlu3DpdharhYoLcGX2yqDOf+ry1Y0QeLAfCvVlJNS/VqWV
J2b0IZnu3VJ6QVbgjoCE3BTFFmZTAVLKOlT3tYxE+vGRIJoda/4TWxbv5Vnek82t
3IMZxqZfBDNOJvsGg7jYJr8ocb5XeHLpivsjle5w8N3opJkN52lB1siRr3zKYm+3
V+zkIdBAwvHF81UFofZeNU6Ke0q8LggfOGHg/ml2x7hpvBa1WPagpW0ZK6sdvUPa
p3LlQvgdO3Y5jOrkn+V3563mEZL+kDfxIxLfvIONAwkd0L3EYitM8rUdK1c4Y6Cv
SLpPBLPe+dQLeug2tfwso8vGfFziz8hUEbbhOLK91KYc6td3fyQpzY33rYwNNBjX
`protect END_PROTECTED
