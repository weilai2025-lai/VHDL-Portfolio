`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyy4o8ti6qWeqKP76o35z1mlF/iyXF23ieLv5cXHWHCa5bo7j5fnf5FtDL3dMW7J
TvSsewjTSLrK2kb6R15DCrOKwMQ9TOYc3isOX6siNM3vWfAO97c2FFK+Ks9+iLQ/
q+SYPt1I5ooKaaXiDF1OYMLmnovNSCzx7oUI96ujSZw6nzVkrWEXNCI4y9pX/D3t
Iq/ct319i+z/8a26Z/BChcFdKIfRWe/qGprZbY0L80/4Rd2fghG5bEHsnL/bQ7YN
18Pxr2QZ4ruUUm9Snt7lzc2JYePLJc7GpWdfVCLpI9GAupl6k7EiY+7oGEYiCmt7
y4brBCSHZk43SvR9zxBcmHHsuPjiSDZxbYOLSkS4e+QjixdpHGZEb0x4tOrQuNiC
d/rEp9C+XIym5y+B2BJ3FCBm4O0aKtEUmC9A0QbKcLb90VoO/bN13a42A//ngFcw
NlWHNqJ3qqLf/tKK0cXgJ9ivFmr/LvTdLqkK8jBF+e9aCR+06eRdht6rHSYVbabj
pWxmU3w1b2KjjkS4360WbuINv8bWni9bO9lfsHK5SU1FFuz1mn34xF5J6KULkRgo
8hJk2g0uEDgUhYH7YH8zD2LrX0A+UTFwx25LEodyA/QqaCa4xJR4nhA/lUmvk0Vd
5MB032bIhodE3liKTA94XCNNw5DCFNiaVshv+CXETyBuZwnPHFCV+0/dQGV5DqY6
rQOn0P+hKzGnnJrN6cYxdMlbGNz/SrvhwXWz757GRu5DpIrHzmDrSsJpxH+H61qd
Gie+PWvYbfnoszVREBJVbB+LJEw50KvVoAERzHo1IiIxu/cW8xVYNwj0M9trb1lc
C7Py8Tv+7lAlEgaZH1+wpMKx6MAqwaEWg10Oek6H7qhAP6EBtOiQ7b4drd/ova18
bGTcVADSFeSZVhSrW0+7723wVc4tyDSKRE6bUBZrMxeC4Qj+imk6FNiFYnMCbz0H
KAntoKeEdFDaO9g1FWheGGoAolOVoDjbezlvOR7vbLCF1d+WG1b7V9xkxXPRwfD6
nldVF5Bgk696DNUjzCG3WEaYEWJ9dkAACrsrvwOpjwLP0+Twk9DR/n4uETqQLTPj
n0Ypw1cK8vSsEcu2t/57ZUTDaRH8ojrXvS2LxmqgSVLUpA3zgvjb17qzViyy9hTq
GzP8bgqjwAGhjtgyNt4PxTmQPZDk8Xf2rWlz7Pv1Pib14DLvZThTgr/P1IxN2hQr
jC70dNlIPr4Ev0jCL5+UxHe0uyrfe1/z9sgMBKJ7gC27y+hLMD7Y9HaEaNEnbv+n
0FDyZ4YLnzCRhm+I8Ehkf/UOdRFleGtZMzayf5sowkUMbYoGMFrM01WFMNGkIFnZ
0+DwE5ml18UCKx4J41Sw3SIfTcqkydAnCiCfgAaje73+Jwo5oEXfHKlPpLICCdV8
Kf9S69kBjv6pWNLkkQA+K88dDynCduqKcGl/nkYPYk7JSi30lbLmaIL4v/jR5tVX
4uQVUDE8n4q/YydwFWBJvtNVgNqxspp2mL7xZkn3ABvWKsrpFcxUBLPiV3SBezTT
ob86j7nHmeZntOq0pTXkpxthKoJQ/sEfjEdtjQqEIcmyPE4Mi4+ZMNkp3GF8ijHV
bL5pNT8pTnHnM84WMj7N3YQny7ESKi/JL5+Zw781aA8=
`protect END_PROTECTED
