`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/HqyhyVzfE3WrPOxYnUZ95hzMu8hQJwBsF82TTgZLx1htliYOqaRC/aGRCoTnzlc
JhedQQLQjeBD4nI2JTDezbG4ntjsG2YPgcQx7vlCwGCbsg+s0n4dxx/7aVgmfjrh
JN69ZBZL7ZK1ymLcFQbt5Odtf/V1CA/Bvsh7xmpiImzHeDWomlVL61B+J7tV2Qgb
/nXliOhY/HxAOjqbi/CygeCcl5oBGvTDyTPYH4L7bx9OVx6ksNgiW5Bk3ESgDDaQ
3jhlXxbZT2vQ4+nUQ6l6y7H7bTGaG+9+RTM6E0oYLdMApnWuH7LwAbPEiZcifdMa
+G8p0scxSIbGJiKchv4wIxVRbxMiJCSiFDWSGMqjfU7qjfA8bPiUaGIA9t6lYMrh
y1/0/0ppJY6SZQI4Vr8sjy+5cnny1SKYSUmgdtU2f6ogy9NmzQEtKm7TKH22Vmex
e5YP6Yf3aoeF7nEOT/J9t26MknJ9PEWf3J//391EyoSH9QoYTH0kfb6H/1BBgPlU
JBXGxJNJBDwRTed5g2torWpszILWYbCf9gtVxYdJzj9vFJKXLWggpi0aoX4GWyWI
Q//Q4t0jHQmFsArCgit8yW14MLs16rxpJwEFq29b2cyxWvOz3ycklIDBo53zEbRM
k+5cpZLguA7VaygqbdFd6hHQYF7pM9mP/xi/Ry6Ln7cSkjCRM4tUMKu7dZSBxoR6
8xYe97NKOjGfKn1OGuqD+EFmiJnGauUxta0ALrt5OQ63yhwKEO6HJuHB6+v1JNx7
MMIjr2vYiwICZ7B/i297pB9aaml8wgVJa/qWTs0If2BLwUIq4Tvr/LWPIvx0vOis
yoxW8hngEK+kIY5ssmi+myeCwrehnB/vUX71t+b6LAqqxp+3JVUWCyafteJkM8cz
FR7FXUbtB2a8gNFOTEca1OsirLn2xQFyHAsNtgPoXp31LnBGgud85f2ZpWCYYx6n
h4EUaIooRkev13ni2QIrjVv1LeKpvtMPbM/2pk9gnTQZ0IX1CRIMRJJ529yOnTCe
OwPIs+AIgAHvTAIUnTLEZUuOg45PFxiLVki0OqJKvNiT2HJywggZv7vxY8jilkvF
9XI6J18xhYAzvgLOLa2FcAxZ3unbpKpYiDHYzex96GtTOVXFcyL8iBp8wpixApts
NFKB+FjUJ3RNB1rrMjAIb5XyjLFgFbg8iBTG7ClgH0J5MSfNd054yVvYY1FzsmUv
R7wj7fCTa3MZMSEeRRTe82/YSDAoDeooQBm3kUeNyFWyeLf+6IIorY89JSMP5/MZ
nbhzvLJCv1LjXpSwThSEOg==
`protect END_PROTECTED
