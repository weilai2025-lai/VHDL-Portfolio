`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYudQ/+wJ1zlXV0zbSHupDtkq+G9ZweQA9Y8ltWX56XrxqFI+qmwAi1djtZOKIB7
VIjE6IU+w1H1XEzf9wrxiCqvF5eNY2wrg6/eDAiGZVquDRAsLdtjXVPdzxHCnPEc
tjXwxExG5JIzIea/uDphyxOzlxyy2Kc69gKn8FikICSmegGCtXVjGh0gpgNenG5r
fgoeiWu9GUARqH0kDTQSG6qLpvj8xdb1FqEtrE7qhy3J/GzYj/Mp2nQE3LrfI4iY
IFrcexLkOWOZEYBdw5aqrldqlXNhG3jcLcXzSdSu3zVwRxQWrY9xcJ/ufHxow4KC
QqKWcmxbmq/+ZTS4ce+xtcFk7qaQT/b4yVI5aKx/VyW5R0HbtbnwRTRS/i97uFFI
qXDivJCsg2t60thg3dHCRN2Z/sd+GKjABB/e+mtipuA=
`protect END_PROTECTED
