`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gb29VfYaSLVq4ZDqh9Vjk7ZDl0Q3kXcNkf6SflDoVMQSSbpTdz8LJBp80t+FudBA
BPSE1JnI1wqk3l7TyPGfkVuNheFPsD0w1swU6KU3Qoz13p2ckQ9/4PHVr4vF3cOa
gbgBkRHaKAZk84pLM3kpKXWzsTiy2SzYvMy6lGboNPTltN/LXeyvrR8t+iHoMHHP
694Q5OWXqoCBguFfCyCmZujM6ITYTEnFR0TMMhyGTNTgzmGEyOWb8KZry0PSu83b
4bIBMk8Ut3bAyoyLIwqAA80NV3cEKEYSe9NNK6VSqljZyGYTDC3c6vilhjEHEr6q
MO2ePiMTDfzRPXqq7STp48i139eAQeZLFH1YJtR0S1RNFzd4Rus4UkaIgNeYrUR9
+fE5C7nCPQOuk1dFUC8kMrALGJUecxZ9atXsYRE88LxbEH0FHsKie4xCT09yUX7x
xayaDxwGR+fgh/q9hbdq8LfwDzkq76T3x3rooqgDjj3mOdaLLJJunVLB4hUn9aRQ
5qloM086fBVIzHwxmVvvr8/nQSSnMSCnnRBNhHhKHF28mV44aIEoSGbjfuZ8vxMP
8Vfi8huyqBNAvOAhzxPvX7cPXRY7DO1907Bgwq4EaNe40w9mdQTFZ4I/mC98//pw
7FUAlhi4O7SBxQMS3o5FfARmcj90dVMcgNufxxE0TK3wTyy3gxyxTTVvuniOPcZ3
tdn67JvNQ43yRZxsqRN26A27L0TNrquABav+hwpr3bfVWF36CVCpPKosXRGQv6U7
h2dbynM8mJhuIoYxDAN0ac/Qpt0xJHgKUdic7gr+t2f6ErWOh1lnC9e4aPZ1aAOr
YWf7SLPo3UK8sV2FaTidEEAUIoWBSyHW764QnLXnHq7rxk/1I1JNdd9w3KokN99D
gTZXpWZM/9c4JY22jyQUbmcHFfpyR0/6RJ2R6mhMYElMXsNy7SNmpnQHFUsLU5S/
+JCi2iG5Ytgwpo083HZw3sgVQv1T8M5D+PlVoyAZ/64pMfEx5E/jSKmUb1eEZ/pj
OTcaH7oxbGP21eM7TIio9dnFr0feLXYWFgzd3KdMnRvkaurItgk0Er4qklpLbTHo
F8RLyYtWmpFpCBaigYOBz2DAy+wWpfTnCCL7IKDnjXU0thq8fJH1aELbU9KDJMZU
7wUKa+dbGKboJMJ37sQGOLuaQWSlER3ia9eFDQFXk71yaJTh8X6SxyVGDeTrGxQR
EjCvyzy9uKXNrPmjECts9pRTmG1qYfndue2A9rItnjxKnrRkaxiL+npip6yA0fnZ
t8bjr6jJpmI8iXLAe7s7pCJuwyFX2ujMDFfNlfa8aSYzq3AzsgoddMCTQ9Xz2Ov1
bXdadTbCRREjh2Jo9CM6poEwmFcCANyFxXPDXUJqkvfo0L8ALDR3GoUgOVKykGeT
ocKVlHdYiN9D3ZeqGJ8eepL9z1bcczxcgovwLp+Dl0F4Xmz6yQbDE0hVadT23jnR
qQLWLbdXJTXCfsr2PoAHgdw7I0DQz7gYvhHRyhySFWC0fuAUVj9kPqN4W+atbCGr
/kNpnGgJKj0qe38NKcwNYyXPe97xRDxEZIrTNBLDhhZRvHEEF4OYwpseiHt1XkvD
I9u+pwggeMO5ixvWm6/gU53Y5oEb4pYSgYp+ZvBRp/PpcQbKl4L58dPIeXHmI09r
F7ecGXzqpPUpZmD6lYZYaYSdTQum5T1ZATRfB97FVpI8cgLYLqmNbTTx4uLM12WX
c1BIktPHuKTMxn2i6YfF1EqG7BctQpcZWSkETqWG39mKjOfE4k0lyhMikuN9JASq
E6LQYpk33fu+wd0FdyeMuZqEnvp7eMzAzU0kGH15kGxw4rR4aijsiLypfJKIz1vO
AFwc9JoqZIP6g7EUXGaQxiz+5Waq9eNYxZKODH2wfzSvZionh9ey+j9ExNMggCwS
UaJa2kOlcKlT/6fW4R5sNXcwr3ljPnm/aIUnJbcGic34qo+6FIo1Yi5nqGwsLZGu
svFBpLTljLb/SDI1G0SDeypux2zHEHXLHADEMUXy+BnxTBcE3Cd7QF/sfEz3qgtf
FJeACdSgPNcP/JMQCnym2hBJaQHVChbPAAG1rGcZOj2J7tyIEcBIr57cjROKUNea
o10SyI7yybgvEpykzYbM5KlF55TP/MqMmtsSRCY1tLrNjmkXhQyDZkTclbZ25FvC
HUdEfnnx4D+wCFVI+uIgW13QGyLQHiq33dmK047fPqV+OT4+eD0i0qtduNWjaVXZ
SvuoIzOCyKGnYcFKxu4yFmATsTn0IHh26RpM1K8eKSjGLlSc2BcBPIVH8y4kE4Il
UAKB8enUXd8/0Fv5gBsemHAo2f8AdVEvkOacUJd7sUa4n9d6fj+Yizdf5/FKl0uy
ydhvU+JcRwqbjcduc67lgA4liNTPCmkMfmUoDkn+v+sbOIvPPvxOTz97DiUKqiER
lQ79rBb+h30Y5CyAg7lna532QldxEWwRh65SuyIenOs54b+/xpODUC+X/eOO4/zS
HQVmMTT7A60oisciWOcSZAaoqu3hQdrj6bjvPkQqatjV181+WoWwVC90mT8TCkq2
5U4jbuTZ5ViiXH1Jtt5FCuHAkDjMs3K+hqs1gHq5ea9gFj1Qpqu4mUBZvg38oZGF
nmKXz52y2iTDjP+yOmO40mauOHJ7yTvqxJzlpDniCsaCAEYJBUDjFZOrWhTNASGz
QVLP9l2K0f2KAEjlUzcYWdtEtdFfSUGAoZRCh3gfu5qes/YtyZXdaDl6KRXYPo6M
/Jb5hlIqpGHw3kHDWEKHGsm8erDkLR11Y1Q2LN+5K21Ge0a0UpqAlm1MtofaOhuX
4u7Ig8rkVwvyxa2DuLz+X6aXH5uehxfrcknkpNK3xZDgtXERL005mb55IEZwqkpi
+lakKhoV4P8eQTshvtUkH6h6gkhfWliwac5V6ttDSwuncs+crDD5Ule3hz2PSqIs
yjRzfIV7C6r+wsI4fmjvmZk0TODgonubUSqpOsjL8fyrGvQLw2pGeEA4b6lwgpO4
fFcjhVccQtDwjaB93lvPgp56UFJEfkvt71gzOXPRXisRNuZNjCm6KqhJdzMjrorK
ymAJ4LIPnnVKRdyhUBoIIvPwD5GwRhQgMa+DGCvSza2ut3raZEer/Bv+A77x5LXu
lJGBgLa6+SKiZTSVUgr0ErFZPJB3wAW0cyPD6JoUxQOeUmxfxoNkjI3lP8Nmnmi/
7uqbr18b/m3i8jh+wSoB8Tmj+0xUNylUjx2Xx4pMeWhewnm7ifkVOo8UEe5WrjlY
2U/RAkd6JtoKxyF4j6mYBsY4HNlHGIawMPMp35JVsJU5RO2rswU8wypz2peOJDRO
RZ9zhFXA+mXjQJ/ay10QVqw+Hux2VzrsJbQAe+7Lyr2NcuT8Gi5CSPxdLOnM0Tbx
Osw5UxAWrh3votSZ54heLzucvOCWYou8aeM5fgzZNFvX59/ZUuMmB5YEKzJrQDIr
H2Lv/MX34x+s62FDTFzYDeKvf2to0mXPIzm5+RLTR+2N4dwXDcIQXAoMxlTgFSnf
HQUDKpIaUIrZ5/tT80DZvNQeNpPeFjjwUayAZ9WuEemIODGc+cVxQa37+ndy7XBo
cVOO0SyTuiSLpvf5a3k182Wj+LUZfscCE50i5lpArSuv9oRRgg+Op66LtU45bgah
TYg4vrgmHU5523HL0XXr+45ughOOm8ZDbgDRlY5pL9Hk8RaZITAk4n2+dwdAdXKo
b1GR5qmymzRl5bVTJjm+aIUw4SSNXjRKywzx9+v4MPLoZuxjr5deRdQnSTyOjrbe
SHWspIzINnfoMOUlpsvGmE0KdW3cKDpANkztBcV4/RUHiGtMgi3dao9UKZ1tBrdi
1KNKo9cTRygdlWSvhDZmHsb5Q0eLSjYU4vfjKOTBWaJ8qqFt78ne672/+JmwvGYF
+VePctVXSaO2CIypwXucrZ59HmZ7UhYZ0BFxHcgdLDhNzpuFumRhkZe4iwfQSeVS
hHloMYWq9fuhHjM/5mZFFNeDchY8FS72PyRdEaCVkuWpjP5NCn4CoWS5F6m2BpKy
7i98wgOz5Jter07fg6K5cNtsDq1CrQI50hcAelUNEJOBHHlWTzpt4uDZ+6MhjU1A
tPDb9sDuyz4+DakxIaMw7Aq9lWG14nNiSYxd8btFlOBp6JTjL/wbYprE1Eat8o4D
EJrpymgFe87oLks+x7Lih3N4MDB1ucY/BIxj+/oAFhLVmeGQZEHT2pTr1DvLt0gI
HmiPp7jSfOzPdJacEf81bZVkkjEcnhGta8qkOTul/I4kgZUukRa/+KPg3tjBcEP1
rloUnk4xg5SeIDnGaEAocEnWt9YiGk/CAdbee1eA6pagszUti50vPxiRQebtzkDK
R+XezLz96p4jPpdm0f+G8NJwRzHklQCioyAym5cyeFWGA9f3hUERWAmXhoWTD+vd
6Xb9DSHYri2or40A8Cmx1hsALRmBtIWZLJY/rbM1QXE2iBzkUCww/MfDoJv9baNn
OSnOfB3QdHsOoPSluApsTJW3XYY+o8bxAtTOkjjHZ1i5qVzANeUGUM7MldsRSjIb
RrB2hLQClkZ2cwQxR/pmIgaQnMORwDOrLB9RcpmECPX4EkG+QaxmE8yiDC7ll3g5
6WvMeUqwj0cQ7BR6EXlPTEfojtcushL0a/FxxZfEe5wxlzJv5RK3Ac0B7ACg1sDY
OjF2aCsiktvkUfGh595HpS9MAEI3nxeKJsDtyF0u24DKrN9KKVmuZ/pJlA1vZNGC
igSf16qdS4nBv95SNK9tjqbxXp6mUViYoOY+HPsP1pvJKieIE3Pheb1UJjT3FBFk
9VuKZl1rLAtVxWS/V1LCGuSoRatiApKHAitx5Jy9SHgTMGfUZhR1Yd5zSA1oMSJa
o2NIGueczCNRl5oDxM5ITyo8QR4EsRTSkcwh3fDtqkK1Gl9A455VOf+ePQtO9X/3
ISsk/k3bT1T+jaFW99wt11OsQuN0AUBkVeoMOs+RskK/lUI2XnAqu0xenlkHSh1t
Avy9cBB8xEvboM07tXszJyqVMesrFu7OINbVtzCofxYj18lP/FL46LSExp+d6OcE
ksTJHa06/lr23Ype/8zoVXp8jPHfKuJ+usrvbo+YWKGaj7N8EGO3bgnk8a9u0Qp+
hKGEftTHpLFr53HnBFdAE4dZA3l659lLfmJbYcfX+MZUPv2WNsfBCWJ9THmFBdOe
YMRYz1Uauy6sj6xCVkh7cdkNqbKOu8tjgwhx3Wfb+i9hqXwwHYWYWRz/yG+dZNK4
mg7j+LZ1pfhjSE4n99VVnWaQaoGAKHODFImBNuEF5H7oSVCEFWh9V/D2FtdZWsvV
a6j9HIU6Ua1YwnsbijYL+OsuPz38bnCkdsBcs2yhbbPvALxzlkqRa7IXWSSiC8qj
S3Yn1HvB6a950uFHqSY7Oofrpfq/3Ui01oTZhOLANFtqpHXQWUWr6R3+1EZ0EqN4
Vg0H3kUrthyfV5hL0ghKgeUOuBpkuQvGv+oYJJ8aP5GjKGDb2sMgqOeBsgj9mR4R
FApg8sv+vh8A4CkoEbmta2v8Kqvqa5N8pGgltJP5rCH36L788X4oPL+2DAn5NBqR
1QSY14T/hYV9rubBC5HNjTZOWbuVvNgBbVECsSRa1O+h1Eke+SXpY1TiMGXBsa83
luYSLSRM32aCza7Hewh1zQ==
`protect END_PROTECTED
