`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDnJRpnjtRXXbKWqMcn+/Ms3GuQVsfFqr4d9vn6vw2Zaad+IUN7YImohrSVMUjOq
ZGrJeXKQBobWTCxWYTa3mARJzL74nOzaGqu+v6ilSlsWK7ov/+gvkOUBnDIiBD48
8F/iWL08/N6qG9iZbfcrVLJJLl+QdYCfwRdmIcAfm0nQGbLH8obv5rwW7KDXH0M5
GoHjOd60bn7tI1SGKrK3LHQ0APBAOcN5DWD5oP0aKR+EBu79C5VcLzWlX6e+YE3G
izm2vb/7z4psLvjMGdu3239f/7tW5n9ydHWoVcXGHdZHaQBF6fkYoNG6QK6ivQiE
KH/cmORCogZfq8BnyyQQvC2a5f7Ef6gIqECXEcdoFqIqLDvc/tL3z4h3HRVy6keA
JKAZsoIVbNqTDy79e5E0k62V5xg3/Gf2H8lJj9GARknMbkfUD7TLBCugDdimZRhQ
g/PSV1c1RqJIxSCIwCZf0A==
`protect END_PROTECTED
