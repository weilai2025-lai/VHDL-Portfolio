`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rZeMkXmGndca3L89DWrjvH9k/LXPJBTOOhXIumrdc1X/wwzPlgUssMxjtmq5LlJi
+vfLwvElU7jaL1lgj+bhtn2F0YOTAYlSclyFN82Rj1Pc3RFyIVNuSXLnoA9NbHuq
NnGPZl9rLLPNr93hM4O7duLoHx4kxNMAO9CSHpyLFQUR6cO+VflbzpCfpiuSI1tA
pBvc0OJ9X5sAHrmEAwDGw4kz4jO9SpXH8jg321mygMoEyin43UuRht4YT4ntPwgz
N9m5dreEqCuU0Iqjik6ZRtPm+FDE/rWAoFv58uwshmc1DlCdgTBeciJifEA0TS6H
TMkeavFUgMZURBeLN7Eyg+5PpOV5Gw1/4YLA6cZhhqzP+qpvhh5c/x0iDETMA8ge
SkQ/46UFXUYSOBY5DFW7fw/uhUzAxE56tQlOdDozIN9zne1G/c6WZ4BVghWDKtqE
nPYwqtdVXTAohzqyDLB+BqNZQo/gxOHqzOfSEUn3+VwlkHAAUciLIH7+sJZPNKco
Ye/Rr1PQkF6aj5m+vrsKAtUyaYLXWfGyhmG2rWmPqh0wvHszulydP7RSILbJn44b
kT2zzv1O+ltLgmRc5Bu6cJ7cm65OT/waHjtfuMItleFcqREeroQ3fsMUmih3H7HX
91EAKdVIwFeVfq7IgUbL47ONXC1+5PO5MGIG9uy5bYoK2skvXkF4ZcscGf9fLYfc
Xy5omRWuQ8i9USJ+HnHDSAg37gH30oqW3dDNKdM+nxS1plf3sbcQK/z0+7FC17+E
P9G9AfeGNGP9UCtETvUOb5SnTJNQu6Zxzkh66qPjsW8jsh9qoqmjUW1zR6HLAy5M
EwgY/vfMFtj4Ci/hw7/y6siX0Hfe9AHV2PqbEuxu5/9eW2AKLABk5iR89ycHvfoc
cZx/yT6cpyui8Xqf0yV4z05Vp9b6G7eciWIgiXc7wB8defd0q5/uuZcZM/QcVIem
ZJfNNjnOsRqZq0koMuKTyxfXUxVGppkfUl5/TPa7atuDbjFVtZSNLIEA2v8buitN
54Azfm0lO1E8MbEITGNUT+O8kEoCzWN0WWeLA3I39p6zOM73c3j7m6VNJXj0M8Pc
dYgb5B6jHda/B9AvI/zGC4ogUfO/HWWEhYXP68y9T1kEaeub2BN8MlMp1GUuH7sz
FscZCWFwRs3hdQN9sqqNT09itDpNyJyqD3ZFP0Ld+eAGeWNKOx4na7Gj7muPB5P/
vvbhJTHqTyVANZspWdOdrIx9MtElq5hTamGOoMh1WfDp0FRhwSGQz3eLl0j8450F
NgnV7mkbnotcAAreESRdf7iLFGjKfw/uzuPs0fyqfKaaG60V8RxnPnn+qMlvwAQQ
5ZbZh+BlQQpREPV4vYVE6nnGi9Vr+Cr1nKeoww2ZwnGyjrf4tPKhAqG+blOBimLD
DT2oUIIo903Pla9gy7geSbksO5AZc6LZ6CmzXWl2eTQ4OZdZyjF4ymIKyWBziBT0
uRzK6CFhdx7733CKmOw4bie4cLcCV3iBagtUvHez0v77MdP3Gd0EOnEbllVtaRt8
0KZ4gmImR6Y5NDNFpM57+O6jUm9O4ALd7hlEOmAfq6qqvXqYKuoXSTO+mpEL9kIW
69sZhIZWvJyYL/Khhv/UEYXMdPePAreHJtdlkbPre04CGtcRc+VAgM88EW1JVQYj
ki8EHt5OaOBX3THC8zr/c+AspxfMFRUHAk6JhFbCXj8ESPhURwnxn50+G8JZQ8Yc
jS9BuDM0PiPIKy6NCGr+rAwLhSkuma4WYSwURzsgkOTWh2JYtRI/jgPgatIEU2SL
zvzXcWqN/Pw+lnq+JgxgA0qLy9QtLdOZhishP2zuIg0ddk68ympn6oD+1BUvVIor
s9k4D2ybKgXpagTuDJ8N/PqgNBIpCNSv0S1MuJMwRrdHegx0dnEkRUFGhzc1JB/Z
Bwx5/8zgcbsyyPqkhIkPAwH0Ny4Tigs+b89gPU+zEqRJeDzK8zKLDuwKFEbZOe8Q
h9F9oDD+L0E2ba/BYRUguvibg2ujMv4n54rZZrir2QK0xwYnqqESeFDh57sLUAo3
PJA65oDrNFFjUD0qHjtDMxXtQPUHAah1aMmv+9LY85ifqBOhe9axr/c5rLHqrWlG
xQGgs1WqEadAFi3eQhJ+aXPpiqYRmcb7VIYQmS7vQvUeG3ilWXMogt/FTIpszOZ2
IsAdvKV/7ncpXC6hi+JTwGHvC5A1q75EArQfLStdOQvhQ7iU6eAggx4gXjROj1DD
oiP3xu943B3f1LNRNiEsGRhKC97666whJQh3O63kcBHbOOAfdPZSe/du1xHyAek5
kTZK2kSfB3BlBjOwfwl5nUj2xeXiVSqoiwXBAhf+VwWLdydRoCq0uAJEPpoBJ8wT
dCoaM2WEoxdX4E3KXPt+sovXrUg1OE9cc2/Vpba5FpIrFwRJkc27Wm698VmrN4WJ
69O/VkMgAfyxduVLJRU/7Z7up2hFHWj4s1yb0baqAV1IyjI68vumYJLPNw3PDjvz
4klLjpN6gjcq+CeGHPvp84WZgYZtq5EZAfXWQycoOvfHjEpssJHcKwppwTs6Yjkk
pwoW//Uc9AxTESsTg59A0rEeMqZ54h7Slb+mQtXPvyv8Z3ds/coMXEEHW428oypp
Fan1YiOzSrF9mra+g9w/wDA2BeD90P+g0gAyuOZ50ViRTypN7HJmklUCfU1SnKGv
llgBRIW/AtZQXqQmkBWeyIjJEk5U0/mi+LB60NNMZAt+03KxKMKxGTWxFFyJ498a
FypKE3m93r3xGwjHnZTVWqHn/+p66oEKa9SSbFtcqv0q0EwQ3JOtuY6SgHez/NnM
6GVGW//pGemeV+IiItiSDsmKOyXRgd0y5HR6qQVt2h3X1uACI4lq3MO0ooivOnH4
b1RXRWa9Quc7Y1noJPc1ss32oqs//qzgp526OYQri0csWa+VHRSvYoa2XHVCmWYI
tNrKhx0is/rgqAGbVmpy3THWRm2LTGN/8HUG6Pj23h0eTEXsbXgjheHRpr7g+Llh
yzsE+HJIerIauIBnkllGb3MSaf+3UZLbaw1fbaxf62Q9gb4SMx8IzxJU8TW/gqLM
RwrGbh5QdbRcZ8vuR7BGgs/qGlujdDYIBWMQ9Q3veC3CuAR/LCkycWw39+GrS/yO
fJ2o69wA4VvhoY6EDFGzj71c+auesoA1c9Nls7OagQfXi7UovzxBL2GqGaPCCEcx
NQBhLOtNMOW7KfZpXH8vnzCfYgVB01yYK81nRBhMFF1YI9U9Bo6kS0Yn1WohzcnB
sLcymk4CLnW+bTjLLvMjxPmoyKIMgHzPk1aoUCf+FYwwNOE92iMLhvOKY1Yip8MR
KtK5C88Z3k5C6IM9xLEmqIezPvR9nVJIQbk+5Kpi/vBGIeNOu61FRU70nIMZHSry
LofYPP4jZ2RKclVhI5NR2BpSm3CZi2J8RnIeKWWRJd3fNfODZ47VnZsP15vVogZs
GQNzMoIWMrD8a+LexTj1vb4Xlms2TGbmT00pGQmHHdvHkRwQcki4mjBBjWptSzJ3
Jnvpu9YDSTsfAbn7ntsbqtgOdAuM9Um3rWkpj9KY+ZAYeB0f//EyYKOYYrXKneGt
nMVKuO/qrndDE1eflKxhEndUTJOIXkdEo3FB5BkrnK7n64tUWv60LoY5qgkpnTfs
VOF7aiPnjUISrujWfIYyUrwEFJwBLTsStF/ArR+ca5FgqtPVNCqmwbwR+B4knJZt
lAtmYU0Lkzz9LqA9HZJgezGhP4ohG2RQVdk+x9DY1Ux5T25j6KaYppDQuDfOQOAU
bKV3g4HxRdMH1k6SlgXZ/tb9ICIblVeUxOZFazaXNPfg7DmjoD+f6Kmr8aMpB0Nb
prHeZFJZvxqStAKUxdW/BrZ5Cbi4DgONqEus6IFxnv7yaVM6TotCwqT/KHXR5Nkj
ONokikJHrOfohTwXUKnmrLw+o/oeb3m69siBBgHyDNzlCcOWaD8gbTXv2LTfwRIL
23J3ecGFfY1NF41YFyOipVXfs9mTS8I6NmCjS4z4fEAaHcZed5JdSIA0qQRZ5pAV
sLytqJIb9LBTAfI9+5oKAxsFog420pqXi0HhrZX62vqmg3qdMGX5Asw3rZwS0+UW
vjEMK+dpRkhMnxcyY8qiLq4wm8bPsW8D47bes7zN8aJJYwI5usoZalRfFGMhiWOA
uzp+2T13ExTx5uNcDKVLJnDb+CU/ee+QB+lx6+7c7n8nMxZ4sI+igzQNflRDSr4B
OcEVIxJ2imdA5oximaA1v/OHFxKb3EDAQHWcKReA5HibiF2K1WHinKsX8NG1LiNi
BXA2Cu4vWZ8A1kInoy29JHYigA1ScQsSPYmfKuihqSCL5mX75JZYDW/B0OqPw24v
IdBrjUvCMxCQi3DoOrNsc3b0rKbKlO47q+dRgDr3woVXmmnEj05jmq7QMKbnWSfr
vi1qbWtJEbF9pw5MSJmFDgI123cwyEEbPRL2v2BBsLdjMdfqg9fNIPiVerb+eTu9
wyOIFWnpgnUDDjgIP3Cw/JFA3JrceCOpI9cun+QIzuD3XB9JezQY+bAJIiktTFe8
FqwlGdijK+Qtc8+yGFA58wF1GTZ+7XM3Sgf9NXEI8yzNyeiC666qS7N4c3Ix9ech
JBiy20hgUiyh7nUhgsVc73FX/5ycA82aNDozFZDiMLtKKXrtyrkyQl2VRAJnzLzO
vvRw+g0hMgxJF82TkTOzJ8csQlpi8G6nzEbgETvdA8aseE7TNq9Om9tRJaXh73Rc
M9TNwfmB1D6oAd8hkniLTkqyWRnOX/sGjTDgtK728ulxlLSB3XM2oOWNLku14Wzc
eMuQ++DtgrvZLChdOMHNzs4goywzWerNRGFBdT+0lXi5JHLEsjlFGqwKkMAd4G9D
TeZfFOKla13oQZLT3/Z5qJFCBVkcjM6gTrtCBJD3giewJHB+3gXLXO4GvnOx6keg
wnafKZ5domQ9ilCBlNEGb9NHrVDel4DU9NnNjMPPQTwecxwirSy+2n2ZGnF0Wkis
uAkYqxbiK5622PKGgn8u6LnKDLd0YtBd+cUqGsMt1MUhFgLay5/DFLl2vleetSEL
PCPZfwq4hyHJMKXsczf3r+sGK1iWVVqr/pUDnjccTbpjCQqwHVadggTHZiYjCgfW
DG3+okc6xlHrlSWNidzTIfxbpMJ+ZAJb7q7nNnvj97EplOdvyU8kEt8V0s/oIhq4
DfK/U0zpyH74PEb4XLvoxTkj9euYCNPA6zBD1qFpECaYvHSWjRiwcbYUfKDm6N+q
fS24NjlZj1NYzePZRYg6e8jR8sUkat/feje2cGEg9tHMWiZkdJ3Jp39ynkLGZIvN
Xpv1goiAFeosJ8YK4/TY0FuiS7apWfiknXjl0goAoGT07Jo7Mo0zBKvLIefzk0Ot
YB305X9841BbTylv2guYOZiwu+x3DvTkf4B+ed9Y/i/cejX7wPi1TauiSiHlThe3
izUEGupvAE7ypdV0OjeHYptClPmT1xFXnz3EADJIOI6uA+dsPwh14Uj0vXcJwGZH
ra8sw+NpjsWbRpgnxo9I2+b73/L/aB5tl+6mmbDejiJF1GFkc7mOIvlEblkexY0u
mOmnVbr4FtQ/lqb0q0mTvZufZIuONJVw33BT0XiPXTlC6V27OzB+1WZXkguatDLe
xCzaKmgCyf9HgmTVGZiCQx5WQXXrGhPu/3lvAcmYVqdSMRODWT/IP1UqAewiArsh
Aa2G1imq+UnwMeLxuIBys1fWKNhrsxO1v0LoHCOjMOEpgcAiJOcN7vFuS3qFVfkp
g4JnPI2mLwaWZyN/yRJUJ7s4cu7JwEsqy0lX4p2xNBGHi68iiguARiTQPylxDOu1
mlPSOvrZRY4/JyAeMnh1wfbmnnmFnIaNL58vO1oZzAnZuirvT4rGXhqWObL9g5vg
++c9HmJOb5yuDecaUSKBVGjmGnST9eEqJYDIkaJzRXPi4XKMBdZ+CPlfdmLXwDQg
ezTYv2CFK1taRUziKuqn5O+i/u8tVcYwIlJZGIQ7VexybAU9rJB3UQUU07mf1GyB
EbNdaQk1rJh+0WtJxh4JMdCKDcwHsrtBJ4P8qwVCAY/i5v3Ol1/OEEOx2ookQKUo
xJcyzQxYqSYtzZvoo1ApZYBkQf92lyDASYN+XdKbWRZQzERtjnMF7PcwpGLXiGX7
aSPlglrKjCXVHI8XZP0sMmVzdeEg5nO82OELWXD8fLmADRwmp2c04Wdmp+LNS7W7
BjuFUrQaurDB3S4UaLuAxNKWSpAruz0onv2XVhgG8Rgb0VTmDZ1kOd0GpxvIhike
s+mnGJknCNarjNdL0uIaxnihrF+vGXiXLVOk8GdOl5yG+4fnumAbVj5vfkbktbbx
Ctfe62V1zePiNMbR/y78R+oCDR0nwaxFciu+rOR97XgjzExhV1DM9eDRaWOn/FOR
LAVVa+6ppb7zI9lSQR+lFmqRDWaalJH5p5IfVodlNc1a3e42S3nyaorHC5HXzKjR
F/wtiE9lrKQw0uODmGpacb87bM1tjfgjQczADDk76o1Wlr+zvAQ29UENTdOpeIRQ
T3z+5JkQbBfMBKO9eJNC5Fukk/URwvAJSJ8GGcbH9rjas3/At0kllqRyLsUSFPdQ
aC3CzRoFUww5N+gyRkdSszhXmMQfjiUpkQjz4lGP04+peuSdRzlRCQVTstSUhNO2
Pc1nzmkbPnJHT07XbyCWe/fWRM5yWJdUHr2BR65KRwBYLa+FWxjo/jOgcngjZS3P
cd9fM+ntobqElSsONiNfa3HcuoceX0URLUF6OIe9rZCiLUvxOPebrkWuNoT0SqKY
6CPVaL409xd7PJ/xojQX6ex9XdXit2Ft9ODyQJC5j22FUiwO3NMjqpbYgotIcVG5
dRxaBkzpKDO1fA/QxvWwigSPL/HXrqRGgkmKzX1yzd4xLNOMXX7euN+vsPdlFGUh
dhsFWwsbqtIjCXRxKmsoo4SH0yUQWTZI3RiDaIE6f2rj6VDDO8/xXhxm8kq9SvvN
N/763H8oHrMSLX99BE2rdkptsUX6vDBx3acwoOUIke6Rvh4BmnDY/5KsPBX3c7LT
YjZrYY6OE0r7l66mbqZJEwCMwXi9EqyjYAmRkLM8kstGNA+XYF+pHLb6Jhr1h0XG
gXrcww4P/tr81i9tnx7AdpRTJJ9YxK8xQdnIbFVr/mgtdbysZDvEYM5suZ3w4UCl
a/AHyPQ8SasSmDaUgpEbdtkUB6PtIs/1BYeicDuFUY+Py5dMNhykltNhxUZQUd4T
MVN6Cuv/QaK44kkNic9WgOPjMMHmeopVNt0DKQqFNzWQBHtHgz/xFB+3iOY9dh8/
an64WbixFTwrQXI14jZmF7YISRMwuGNQw2mOVWNQwIuxXMH3L/8jz+OPCCVaE2rl
0rmwEusJrTdkgnQm8VRkC+oWbG4tbVW7WuHJYgVbJvsaAv4YxCUwT6HY5nyRsPMl
y8cOorUI1D+3VV0FUUwEs/S5kjb99airbW0cwiydJczbSvNLVb2q+N86Wi4zyQZO
qGEFOL7PWDFtyhWPD+tiKvp0DDZLItK43vTXkeD+BKtZIIHBno1e6v+6/RCuiuMn
foFi7ZmtreR5CZamirTvObHlwmFqxREfYPtK/7shcHpR7lDqakdOD8nEvYUD5/zv
nIVawaDMnlcLJAvo3uV7OiETEQGtsu7rp2xg4+AjqEkq55AEVkaMTh5SkCi/mQoQ
bk17ygMfdMGgbQzHsNb3fpcx5tuEUCY1HjY3jv65TkJ8fDMj5kzezTo4EL+W4f0e
MBYnI6IwLLcsG1a6i3c6f5qf0+KisEf5cDre43yTtMIdzYgZjBQ8OXTj39espzLq
XO4+iqg0EULGM+Pk1cgsp0Sh/xGX5nHdIvVesW5nhJVUa1YKOlWAsWDvlugSnlxJ
m7LEf5uQ87JyPobn7xEfcb+FKdirvuE58Sw5mY7P8ysHgsVYJZEOZMKmOR3gD9P3
L/2eJ3CIcbHj4JAQJE7rSJHZUBPuDAvaWN6YhRR7nOfZW/uz3BLQeYhvfhtC/v6t
5c3rhVJ4wPIuB1QCJ9nzgGhDphVbvU83UmjoDgvC4Gj2bgdEOUWsYE/iJAC846gf
X+cEysYD2nlPXip2BDXMSfVkqC6Dho4BFGNk04cntvQGKwpzm1Egwo3RkFFOFHFK
auPQ1Osm80oGK186v1yrc/2GcanaNsPAg/7v0VEFBZltbLgVYyi5Io3mFIhwQ1WS
R+dCPZ9WSf5TsUd1Z/F28pM1iy/g4WB/vLIvWGNtSBFHoX49pxJLBwoAhEe8EpHh
S+LgihjrU6h8uRbb6SEeFf3ecjJ1t+/w/FM4YlMoD4H3zUvr+kmrhketFLqw3CZQ
Pd5Ehfy9fYzwyljuIrvZBrQeBqzDEghCRv3+UKhfTuO1BAjeElYTLx/kjwXlAJMW
5hqJNjReaf+Oe5QvANWUyro+oMyiWf9yMnSB1HCg369wgQq1NlSqKJKpuTdZrU76
jIG6WdBA0sVrIHxHJdVngwu6YwEkOCtAvZpYpAOgz2mgMeIMxP99o8zeKryp6lyq
MnYPvnt2ExmY7oiiIvl3lyrchZeEanyLv2Hkz3sI5rHB2xExI6OrhibGqnK9tviU
ftas7MMAzzc6FIWMXEWo1UIbbAj+g3i7EqqmZfopabBICDLbVEsqB4Y9UGfU/aVM
UsJHNpGwF0T+ygx6UQx5TUAbBb4vGfp1mxNEyb/o7vStRXkFfSHSC0m15ZsojiRj
nFp5OtC/OVfizeUD7/mEKUpt5BbpNnOK7rvfl6H1SMoZo3r84jkIpMGe/Q0tpxwv
mEwsQiD49qggb7tXPA2J+pb4vvDhsftVvpIQCxFm8291UEBEDl2fl4hdkaT9Xe0s
Mv53N7vHAbutEpi82sEIuvLQWYXVoYyaZcsz4YYoXnErNJaBTsmVex4dwhcJ9iuU
7YVHx1zVgQ42JGH/GvcNuiDcoZ17ERtHXCDca4iACKpaBmRwwiRoPHf+I+09l6Me
AJ/SBCE9OuFqbn/sgHEGdZjX90Mw+xtIj9rjPEIpBYyzkD94upOjomkHAjwVlaNI
s/hEGfVmDxSsmSjunQcDktRJ+2cILOhahfrdWhE8mF/PJjjavfrt1daKTvYfKu/o
rUI2/aBAG9TcU4lww34zzh2zzxT7PRPOTNBEF5UBPuSIRvtnJt0i0d8vr2sLOs7H
v3zbcB21qV64/hYOxOXbjoxJhE1QIdm8cM08r5/6eLx0oS/4JlHzX7RcVSkKYCv0
T+het5PUqK2PchjjCyg2wo+qTg9b5PhLzhkESP+F6WqmOZStT3KZ7FSc9UZJRf+Q
i+7lxRr66NFcdb6rj1E4BUrmPxOPK53BjTfeS3Gezlh3HVyd2HHiPtWkyDsvr2fY
yaOl0RYI1nsb7QsLcoh3hVNiu0OaMjThDN6jU7AWEIdoeMgJQUP5MmiO9m/8V6B+
sK6Cf+QAM3NY+jT946aSfbGm5tuVAm0nbVSxtqdDWdcPzVBH63yOF/wQ0j/1IyGB
na799m5SIzNQ2TIkz+AnQr014xseO/3DDewvK0whUrvdedGAkBZw/zY0l0CXUW/z
2HJazBIS0MwqYw6Gn7R0lsEUhdtdeeXrmjZSXbgD2yfgZNdqcLG0RQ+kg3gZnZlC
B459a6J4XgcDNYaYAaPJ057+ZA3dcJ5XBO8I4hT4WTNvTQUmk3GD5flQRVqV6hS8
CvdCUV25AYv5uTDZ+TZ9/O60CHxgj3oeJzZS1PEQGw7bQqUUaL1iACEqEpaamJRT
AozfO3u85SVMvD9DIQpbiBR1WoG0ay5vZWrfq4ze0+J2IKDMmMjLuyh7ndxvoXgZ
oeVFd1ZiUrL4wZ3Ah4CfuiKri4Vhe9jvGdzrYiPuBthkYzIeRBpefbzWBNgyetbE
TkRXEEFlq/R0y5DPCUfe0A2FN7mqkgINYugQ2KQ81IvU+P5KFfv55EagGLgz2h5Z
B2CyAeEZCV0MbtnIRCPWeOms+a43yXNH3APAIp0HMEh/ou6h981jj5Qq4C6yObY6
XCZW4gjOpgM5IHMlkz6gHjLgJFKgPDlwjbyP8TBakwcKqUiBF5EFLA5McS3NI2sd
MeoMq8Vz9KB6Ngeeglwze3URzPp9XpqZHBOCxJ7wK6yb1LCJbxnzJURgDBIhQXc8
RR6tIiERBtN6dkyP2onJWp/2A4eHWBVO5W2y227NfwTMYRkkUZrM5djdJmK8Ogwd
HrZlQxZZAMjERAGJhMQ6h1AFsh/RmpVXKtYNyhlUGuY7penKJ1QOsq1HzP3L2nVF
FhsCqjVNtxZAv+KrWGgyF29sWN0wuGPZxmT5SUOnTuHhKF9UN5PCSJWnkm3sC5oZ
iQGEn+6ORXUQ7hXasIJrIsEsaBz0zvvHBYRiGjXpBzl7a2nKyMr//6EiecRA/218
yCUHJPROkJK8PMVzjcH4nrwkn+F1RS1u3EU6wNPV2WLpRLgsy5PgnipxPaWZFt2W
4iLDoR7kG3nQwBch0EeFlvOXjmArxlfAMvbHpmkk8qMDT8VZQ03a0lpwz8ForyBa
p0Kdsl+xEAiD5e583IeIEpi2LahvC+TuAo0wuvfBD01iFn1EGY+65smpCiwwoEZQ
GJ2ugmmaqU96xY5v7IF6nO+5NSQ4dig9I2HPjiihj+AHAPc7JHrhWys015OJ590y
hBcwQCPdemkjA9A1DmK69U7UXNEBFKE9qRHIyr5w52nwoX+ptLaAlhc0q10B7sTX
u86sZSuzZVfvuK2BUfLabbf75Z4xyWya+h2b9cYZM5fbGnRPGI4KfHAfZ4iOhU44
hxvAnEf1tXlne+Kh40eRLe2NkBBk5mV8+PiZ+XbW/k4r2NzUFH705IW8Ww0w4IVU
hATkJsgW5cSbR4fXsVFzIor3lIb4bgo5Fd43Q6CfvXZU+AStNmkbUldvEqgoUsLx
CupJKUIiylYEHWhDez+KljQl80p7QO8grNZROkXsBMbuy3Fq/kPZtJ/edgJa/ssU
4M6xW1M73i6hCxG2JuKyvNRO4Puc07aVtSYNBedGVTA1W5rCImjJmc9O2BB3ddyJ
Y3cF5ibA+SkvXcDj0j9svMQMYLxZgky/kzJLVpiECaE+1HemucDF/GxEw7eN4BIz
rlGIA3G7iYKygaFB17TOyqwieWZr+pbugFiymMMYzVg48gyQUKBBDMEWhfgokIKC
zzY5PR5aldrSPHw4TywtkOSSMhnF7wj5/LBxsthYwJhTy4jY/AEMTuW2LEGIHy/o
dol0pnwKX6oqkawNVQshoZR8/KOTniipemoa6I8SUfGWIzgtt8Wp1sEjtkmwiiek
hkbXWbXbwWkrufDZtCwHiS3BFBD2u8KNf0ZXRuTGNI4/7pcyvch8yrVEgPb5JKr+
+m9XdhqIbY6/FNhh03TB7BxKmLEdwCKLPOlIzkobs7qnEMQakE9UJOHZDYpYNfxb
fJfFfBfj3qr1WnLVFRze+dmDflQrdoQ/FtbmBahAj6dLE/kYhq4bBHjqobKMmSPN
qwyPhcXxach8V7/SX4GRjlctgbKwIuL8T2iDfKp1/QVQF5hNYmuRSjC1PC0DJTWu
UV7js8ZZUWmF8LA3KGLjR2Lg4fk2jjbf5bW4l2zHj2Ph3FDNakAMT6U/tkoaRC/4
hAc1SxKiT/Y9OpuW+I2pxpn6TbQdQ2aGvx882MAHczQJM6qC2oYWcemaG1sMnU01
QwjYGkv0YdTxJSZPMtsIVPNdivyu4DnIueYkLVbJjeJCyYENZPP4v7xyhpWCwIRm
/ubBmD22/LOZ6BitjmGpaGFLdZZJLl4pAdvHTEFzjPUiN5JLm6pHu0mOcTaAuuGv
QESzxujnHBClbQo73hDxInU2fgQ3c9luAbxucKf7FTrYdVsXCmFaQloDWBoDlH4Y
6uwwaYIOjOcaGNdvWc0bOT9PpN/JHhurj1N6wfo01cnF2BbqHaFBPx9nopl3NnhV
Sg0ZfnddPFvDeYdXp513KTepfp93QeqniZe+dh2Dp99cti5tPWdGjnLwFveAB4tz
HRCtEanYdS9pk18aA95fGVoLJmwCJMOSr8zi10Sx7e2m5U8dj4bSEjWwgoWM74eY
L7BR+ry2tb2ZcZDj5S2ccFiahqdMl7Nyf65kzVw04QzlQ3j0S6XbPcAvXS5To5Ie
tFtv7XxRDGaF8WEOZZEf1Xx2W3aS8Z0sBaEU0lAREKCjf8Fgkl8i3tupW9Hdrq43
sev1Hx0UNQDf65R3ii7zCZQbYf1PqY7uZYiNOIjTkcgGflM+9s7lBW+5mMzdx/Nw
3qQgxsz7m/j2bu2trnBRfGNX19OPJR8UJCh6xwN12EzuyMB/hDMbz74MJ5zlPkMu
PliTMe7rt+d2hd8Bz/93qETroqDmvTnv+LyCAuLotK9tS/3TKbASdtuetggSzDrt
fa9bU4DHUkfHszRRb7j9jOVrUPhdVCjwjN3WWuTz/wmW3BacSQTpyS8MwWyiSw1m
SxTI/zkZPXl6hB3oAW/s1m+rmo3Kxh8pQS/fyNutYmcQAKdO2/xnCqx+nO7Bxd0r
V88p1kxOiLNgc66+tuvDCrO9f371r4ab0qPxuHTMm0mFVyNuvCkhzQcVMd8xNvUG
IhcnXOqpqN1R06IY06QT4eLhOeHU6PTYQq0ps+/gyCIPT8VgNU+dyZo1aUBMJ/oA
jb075HGLOd2B2zAgSPcE9Plf4uaQ138DLsXapx3NnNY1f33AcxEbgzcX+cbIgjkg
z9AJJbWILx9wPrUAkBMaaDUj4JUFETScJXZOg0yDn6WpJEeiZ3FxsF+1KHh6TMpl
QMQMxNgSH8GfbY5c1dJXc2qH+Rn6YJRVfUk569Q5QyStARBj2eiITiTACLqnWWA7
G7JlVrV+Weui3mEPHDwI48YFsLRjSm1AKViaIYUqtiLrbhVG5rVRRCsE/9xxqqhm
S0FrX1SAAnlATQDAUxGol7O0xGrAOh1w4cepXRBazl0yYrk/wzGd2GwMIhMkj10/
cPBdzosb6AQDNF6PLqHW/fyMb/S1m/bg6I2SGe8BKBNndtJ/NDTwuIZGaYyNmM5d
B854QVnu8XFsnhv7LANsGwnSW4uZ5d6rcSMVLKcQvrZiX9LDqI0wmCSZJEFbEkm6
5anBX5Q+Y7A0M2mSd96odriRTqfv5b6zZa7FOpzrsG2Tu49M/t+SajtgTzLd4ALy
xakqML0Hgabktox9JAbwMuroI6foiRDrbhc+ubH068odKW/uMfMz1kEaUKORBIdf
ntLhuEyTcNtwn1plYUjEBHxCwzUWQ0ytQEUaHtR3QLAAiydqvV4m7B1MAGUOG+rI
buT0oNUDYaK3Sosnbk26wUK4Upguvt2HHq3uTy3afeU7lDE8uiKd14XjJ78+B53+
zjLNdkVgriwZs66Id3Fmr8gCxmAazfDpnxMqjl33Tu0ZcLXcISdqX5khcx9xCMFL
aaz88vPW6Fs5mHXCfGrXhnxqf43xHWIMm9sPqVJ/VimQVY+pJ2EumdbKgPtAeoVO
26OLuR+zCYi9mtQ2+Ae61nqes4aJ8DkQo/v11BkRoK1jLOmFpm3l6yXBGTfElLjX
9ThxDD05Pr56iIwosQj/vgKDJZMcXMpJVcLe6kpRo5WuAcQLvgu9gVXe8BMjlV2s
UI5YuuXfbixxdi9uHk9EMoLBgJLSObBUbxRPruea2B18KikQiigPeuGp20nTBAFi
DfcT4ZeAt8k6bXq4/cS9lZ25IOtW4wZY+b8v/7CntEnsx7x6MeP343rWzhaNecT0
OoMZekjohQvdGaD+6n/YxiaNkEgf5laoYU4yRso+6BUy3a9WXeH3Udemy0CRKylg
BvVFPyb2eOSF6pF2dVvBS3rN6prFrjXX/qkcJX+hJWSYe4Qth70WAOiOsCewm4wu
K0ISZbqac0otlBqimp0UlqSaqQ75khzonInygEBOhwgZIz1zOORSI1QH5R9EZdeM
ULkNejKCEwLfb4hvad3MAQH/vUoHpNCxc0fD8tNtioXGVQwn0zGaAXIqqMOISTIZ
zIwAx4MvygFBwmk/KXsbzWBR4i/KM0GF/TaJCmpebwJuPGEBC80iVcEtVrp6qbbZ
141DWMZ7z0N+/9FDxSptERrwzEacMLQ5ZlCSc1jijfiKyLCrr2gwFumlL8ULwP71
q17tmtMqxVppQAkWO9WZwBQ5yzcLcXM7jIsb/Ly2LKolMApc5C/P1eqHrO/bV9WZ
e1RdaHlGZZO7FwDeI6tE8VmYgGVt3jjZiW8wgP5mSw3QMJZmuGp81j4Z4mUGo7yL
PRWJ5ZO74mJbGXeTUOoGtwbfE2R+Q187L/iokcsbuZQ5s4fmt8XGgPCOJzQdfmv0
QxXL37GByY1z9YXmA+vSoHhuJrTJAI6wbIF+0f2jMgye3m6y4BBxomaPCQe+abvR
QoEkiDUwBBlK4vLg7vOzhNvQgtYBaXPDM6OKuktVusQFAXPkORnXI68iLoXnScbj
TFOvsm/nq7WnYrs4OEuQmKsG3YyG73iwdfeweKNwUOsNXip0T/vgmX+kWvSEpcz3
fv0XotV6g9ugbsMG3Zuz4oxEj87RKNpFTnC3Jckt6QDhimd0+UKDenaupx6c5O4Z
H4yW/9rLpb2MtsMYbGUrm6aBY5vcew6zHFJzBznm2sPgEMStyOHjsHSDh+ipWp/J
tkF6o61JVca2UkGCwjkq5sHzDisn0yIykC755Ha8k/Vm0qcOHt3v+u41jBnOxTgn
VMWzKXSnFrHDsKoYAqrmKH4JyJMhhJgFtyJc8it6Sg8vqnebYx2CcRrWN2/yPZO9
U7exSARlRkXIxY53cZd2HcjvK36p5qFni9mzqsxZMuMf9jN94vjtWOgVrvvKuV/N
SGZFBFNg9n51r3sGtn1fGqFq1RW3Jvz2XJZOh/xwppdoSFDMXVTPHq59/Ce7D1xU
G+47dBrcryXabyOpvHacycB5BGiDnc2r8Wnr+jFZ+a3/xoEL2Y296snD7r0wtR66
cHGFJqWdsKCOghQAQrK0mvnT5npZuLGQXFpRwBpj+j0i+R/9fBGjnJbZEbpjGMVu
fIAVyivwfVxjk6ni6R1ssAsBIcnRcvvXFlRTgJhsrWvcMmVuZechnYsny4GxT6zO
b1zbhvsBMINDCcvwVGie4lJHgCDDLBDcDsc+cS8QaYBN2o0K+v+jeXf5dF9SY86m
9cw+qDeyilzJROYxbU+cAygBqK32HJImk6hGo/FNdG4Rnx+65GAwZ1nJA21OXJRH
yJ0dg1aP3xqwpDT8M7Pq2f0Ioz6OBkBst5oXuoLZiFcxqs5wcbGZcmV8ucYYEaOP
qCS059nIB2GrNYUEcRtX9+jFpMqdOrPTaF3pieSy8lJZpI0rqF4KLrz1Z4x2QKnB
WblZBLnzl/LkQbGhoPT+Ce2Ml+DXucZbItaNPdOhPTjy0hbi/LkSEiGBxPo7M2S3
F/NYVOKURUyaPYkh8PsFLb0pD3mA1nKphk3UmE/KwryQRxa4YDAy3w7Hea8nPfdM
JmNcJTe/LIAfzBN3rFga4lfz2wIYA+jQayJRsEN617osqfw3NXkXzLXVTQb1sCmG
j2vT37BXlMTpDwBLT01QhADnIB+3yrL5m837u2FTJfbj1eXhb20l3W6Uxp+/Iaxk
Ieyx+CIVXn6cLbcqdjPxY5dClU73IYD14svX3nzXGNv5CYEsGiCwD/vlyMBvTaMR
axhnEZ7cSm3vOpqUNIdWppnSBO/lU/N7zytwGdLcems3jQMGoLSteeicnj1OC6OP
DsUCC/3nAAbAIwrF9sS4dOdbbq74TiPJJmOtHuE3h86aw8PNijcrSjJURnHEqurx
d3oD2t6jCA0SaJhmKLZMrh7URB5z29nEPy246LPXbQ3OMGryj11H/LrCqv6CmW5P
UpmvsMCaEMeLBrL2kWvvrF66pBlimoSHpH/O2V4GcdggBGRfQHf7lODwa0hVYKp2
jwAhWAPZHFWE1s4Z3K9gLgLoNGBNrJtvtGl6RfiKdU1nY99z/ab7jgQUOSdm80aa
8AOX+YxoSuBBnYiAsN6DA7MqRSskO7VLLC4CHYj8Hlr0zFd+jhOk6fa2+H8MNBZr
oaHrNf8TZ1sHUYcDD1T8vYFvRU274AoMwWhERz0mZ6yGDujyZXM/TRilkiuUOvO4
v9dcCF4wD1l8L0L03b9zw0qQE/gl0koIl5nKdykFuLn7iiMaQbH85uYRipXgWyYC
7h1ZYqHBPnZSoaT47xxbda15J3pBH1wlYVTWOQPtll6yc8eGPCPFSwAuruA9OmOM
82sF+t5yIJ6DfwWcvrK4RFN6dM7IWlW+Rgvh7aZ2PhMNVT9u5MFFqqGoj0uaptfS
uqYyKKUWtdnM+1L9qOqNG31GYgeX6j8kg32Wc6us+yT4dTT/NuZe8JTQXzHYG109
g+4KT8AU/iJxCdwOBJWAp3y52Yqh2WXBZXcovwipYnYZGiGFvSDtZTqXTt3pL2pf
4HuSR2zf/aCHGVx81FksOKJMLE+bz1ewXlYWWmsw5Aa1+UMxS2Sik6EFxhOj8/FI
PS/7x6tSk7uej2fKLHlQxLUS3LCtvDk+wUveKfoMdef8xorMTx/GqCEDRvx0Mwo3
VvFL7HWrf0VbQMpe3zt9C+PfEVM7p6CizofiLHJ0xNKuv2XxL1DAwzy2SjWVBxY9
Uty2fxgYIkiWg8qzuRebzstkQpkp95tyyNBhFRlrpfCFldvWfenspMyHS/BbEqW+
zc1pfWahoiAnsjlLiTJpaPwl2mh7GCzr3E3K6+zWWWOQ7Jet0ckiJ25ZOiP5eLy6
zfZ2bpYPSuXCgPpvX0/j3vlDYed3UFDLccfiOQfKc06RSZTrglK78JtnIfFfFKYQ
5Ay/osKEnDQoi4zuVSn5Trd+Ms6u7I6yfZqP839WEkEbXJucqMuFUZkBWAI+v0sQ
Yyy2ZbSc2INGnBID54G8pOC9tIAajzJ3pFnaDfGU3chh+y806dScbGvkdmxsJokn
axCcmTbZEyseAXdyVNAYJQRm8YtnOkVCWobneeKh3sovrhnal8K1HSBh3JGlCz2m
CrvMNQECQ+q+7l6D7Eg0TGabVM4+Zil+MWRGpkuDT9n/cJrCmjEexgQIWpEKQ4Ro
IjuyFgvgFnOlFOEZb8+D36Qol1ctGNnGuJGiYbgVXEBRT7YtoeX9tfkt0MTq1CZe
fK2UcsYup5q7w3fNPwx84q6LkLTPOCT0NB/Fq6T3SECrrhx7H+stlOLGfHRvKJeF
fby5kxPl7yb2dwYOT28z1SM07KNQ/TOVJEcL8tM0PST9XuPrwgBTpAsRdhtvReyZ
JuHA+7b4y8QDSdn7tMr9qYje0ITsSQGJNxO9r44PXOYcfD/9fHDWDM1uovIz3OPL
On70ucc5yUCpDuXVOO2dx/hRjDngm26mzimRR3sc/jKCO2N9yj1KZKKxtrJ7IYLu
EzyRIOxmsAZr8dVVdKHRGZxPqizY44AVgYIFczLW/Jbbp1tLcwZegMWiVC7N7nNn
1QhBa+WOlY7WsOaVnpc1ikBG13NdIdwAezXzI9Oqre/1q+EF+cCYvBfuufzNPoUY
Pg0toE0qzth7PUi3ZHv+RYiovbMW/mpi7SLTWUW9XWKS/CHcNf31HHfd1KKZKkPk
tZXAnTkkk0z0iKqhvB63q3Ol/3Hl2rEHHcBgIIa+HnciJZt2krwEGyZ+OMAHFg/I
u2JDZcht//1pd1r1eI2Y1W4+lEJIti2Uc+SKYx5k/CcOLt3yQPmWZEs2ugdV1z5S
BB2FIZvkbCmbhSsLaWBDBKiNbweVoHhcz57xD6mUyCUh1idXflCBJZd5kU9c3zmX
W7El/Plc3A0RJQzU+9Vepu4vWclv2fXl7yCor95mWzoamIG3Z/xoTaMU92bY61UE
jjrmJPBRNXp8D6tlv+HOPxq7nLnxGAFm7i54EPf4my4NhqXOZIztHZNEEfcqJw8v
BH/RE9z1ePVvudA3CdUTWQFRXFNQoM+bKQ5HK9ypl15+i/SiUE2ZCvelDWvlsasx
IvdB8PSnAdu3AJPlixEY7SFaKDeCyp4kJs50O+NpR0W3tXPbpUQXFwdUmZDTDtye
c6veEQbFCWH9JN/IvX51cpxqEWTooOXp5J1cpl2vdN7gn/Hg5OtOoazlKpa/VZ6g
v4m9Vd+8XiEU/cRh+7D2tG1hk2g7C3EUyW2Et8MENHNhC3m6YUy7UXekY0uP8Br8
/cAjNo/jl5nr5sQnuVXO4i3XGmx5AEgfjB0tC1QGUk2gUvqZYREKAwt6FSUm0ZG+
3nmns+qWM1vd2gsXwEiZ1hFVes2mzHxJ9XAPTNGkIp2a3a0TSmqTq1uZnniHxHlU
y0D+qpKZlbbjdfHQ9RIDPRzVOzw+Ez8eXBzMeOeQ2xoDpDZVFpY95p3/K3fh672t
aK8G7K4VTInSPYDNIsaUa7JYq13ZW51NGuN26qfINKMqCrCTAxDAN2XZkhqqOOk6
YCDVZ5l0YdjHwpWCdmHpGEmMsimMDSmp9DvYBaNDlauAgnMGt6+IbGscMJN6qMUz
eYV6gQuBFRDLXGipfGIqsDFgPEZ0ljaOH+urm1aFr5i6WGZFwbrr1rxreqFtw8eo
zQcL1O9TJweWBFEZyF3256JLHasZLIDpGHxC61tKSKh0SUEyXGLECryXobBdX4dz
gbIv04eZMy0OkClwo/jf547ipb4n2FC2xPEqzJbUjEJGwhbYxDgajAsCwonYI/9L
e/2FKDdAG/lV931BTfC3kOuquk+RNUerdP7SLOeFNMRRvmduL5mq91w0vOw2Uy8R
58dZoEpDctfwCllhA/10B5CwpEtoIzXeya74B2is13IWs5wKVqdFduQApyE4niWM
OunN5LW5vLL5Dy+MoAelbWnIOTxy9SSihlr2Xuf/YmdgO2sk6cWeEmVRI8hORSE5
Fj9XVmjFVZj2Msq1GTMavP+odh3ASOXTAal6AHLw8gPZCnT9hw2C8yKAMWdlPvqA
BTpDbERUjTKELHu6j5hpjQmzqxyJmR+H5p1IQLFpdxOEd9zdY03PaKPgUYEOLNm8
AcfN0tpt5Zzl1rQOemI1j3VKBhOmQ8/3p3Ie3iNcPICr60lM77XbXG1Ar6zR4vHD
ICCYP13dhL4e9poyeI1cb7tyJCjRk2f6b5C7JxGU4XYWy355YJzrzzoogowRXQIp
blsUUxCrR8wQfZk139XVg7FOISVTjFmbXYdz+qvEXL1hFPSYtf6Axl3NGP1mqIIz
iB84Xqi3ApZ0iI630W+nhPe+oImhWVbe4GVKjIc6J1TgTPGcXbBvd/7NWA168zxx
xcmIm6oVn4uWt4Rhlerju3Zq9UR+Tn74E9SMybSx3QlG5SRllkjQ8yMyqBi6JSw4
M39cixqmvnpJeeGYM3XLGlYFY5jIQ3TiXfft8j3n8DtA4ej2i5cnT29XTY+8MgcX
ZzXhmV/rMCRHS7mUvhSfvZVFUd+WZXVveV1UHHrQxTlq4nCSbiJCYJxej0KTUZq+
yzADIgsWrXSb//BOgf209QqCzBWe0brDh8HQs+9dIJFqTKijdVjET5ahzdWUTrG/
hYlc38uq6to3/AohsQjjPnDkDIxCJBt3wS0p1dhGgFaVins3yD6kgG3iDMLhLmNJ
SgaEA0XDL2E3f6ZBp4GjnVyeL9kHhNSmEEbftGPCSRWL3NtjQTqiE0TPzxxTwv1+
FjMZ9JMm1Ss/+bF4ybnZPquPcoTkZmJOhIWUMoxQBUYh+VTpiIW8Wlndj2MrQ08W
jPASA/E3aTgVdsuLhXmv+HFROHD9AIf+9wNyDg4JTT6p4ZYuFR9xZXT5rAtHtJlY
hgbCupRNa4vZG0Fb9ReacbcakY9JJted6bJ2KaWZG/z9jBIBSijiHXRe37gkc+Y6
tJULxyMwd8Jv9aSEdE7FQaOFyd9HEQISCUyJl3MVRqk/mjTMjpMJd5Xx1hgIWyRB
tqqC9cQW0jhUaS4tYnQCpWAt0CeAgNPlREJWebpe/3wEXdBilscii6oU8/+ASoWf
LU+NCpZIddB87Z1y4au8P2SEbBqvaEca9CSWEkMTMBLUZC0AOvXMISu04XKk6Hl3
TKd2/plyVHqRcbkU9TEAJx8TynUwk8qGlv1VS66EC9+uCPHdyn9SSe/PGPJXBXBt
aH8zfLUXjUBqiJDSl78rCrdy44RZltZ+1Nyzuwd8nJRiGgAtOd1FMWbAvyXJ7D+1
17KH5ixzTgyd91audt5nG3Hx3660mhGoaC/4Fpa3TrG1cZmabxUK3+/53eWJKNqK
1hCQfl55llydyhs8mZhLfFU/SDs1dfsMxI0NCXAnXMWDgbllz3Am3oAzaenM5gAX
2+OEmbImCnp1lQX/9Nf+YnWldKrp7VeTkd5IAntcc3HIxX/pAcjWigxt5ciwbeOi
mreh8/GfDd31S9FRJwc9MViUYx6sobpanM7Lxb9kvpUyi6lNqnwKh0ZYO05frgoM
ia5yAUtO5tOsTQtsJzTe02Q8hlq4ZnvIv+AzI4gO2qDGsj7sqUzqwaSs2GlGlgZT
B9UF0tPbXsaI7yoYT/RNvJW5xdQzTwafq0gvfXspevWCR4wj3eKICjKkVowJJ/1a
J+ryU6VzxoJ4QmwLrUL35no6uphEyScHKwvJy+dAJ5DWAVgQDVITYQ8nOdVUTcrG
3zOtOtIGDPSXP5IuJMUIwgp/qK7LmELo/Zxv6OXCCpxw4qyDWf8CRnJjqsHkWFya
9UL8DjYxqlBwz5X5yt/CzWuREDei3fwcd8tmkZDa7fRufy1NZBIRpO2hbrru2TZQ
RHqwjm2knBG8OmbV1VCUqcAG6THPcy8gLf0+JAmtrwayDGdjpNVqxpWxbSlzp/ds
BfM/uLHfO3nLXIBhdwMdudav0SQifJEp+KhRkBgwNdSExm6FLz8pvj+8LRvIfx46
wLHDbzkCbAQZRAnh5bR8YrNcM3P+CqyAqt6pyMIuQOF9GtcaiboGb107vYfIp76V
Pqm/Isz6BRIbkwRxU5fr8muIqh4k+UeMufikAKLOdy2RVY6giFWF6k3yIY9/Kvxz
ws/m/76vyyIKVyhIkOWC6lI9nPDlBe0W+mn7i7Q9KJpee055zDVgZ3xq/6Q+wDKn
k5DzHC150wG5RKKwjSTpTP/frMycMbW5ENhSNjptqnPpvVRxLkXxZ1wTKdUEVGo5
f95Cq0MZy2Q0YI2K3pbAaY/w8mQ+yU5fdfwm4znp4DDHtuhf26d2m/QiUUIo29OJ
QEEnCXlF0z8//hGtHliMLP22fAxPTbcVnkTBG9grdTom9ygHqUPSI9Y/xqi1Uz/E
tLWoNFJXarDLUKAtdXraSczVVdhHkG15uLNGZdsmpO3g3QnU08HBlMFwB8bM9nRJ
IaEW/Bfcl2rZmMYguWb3L6L9tTLDHfh26GpBF1HxzmvgeQzbEPwQ3lt1ylleSDVm
aah6Pwh7jXnmOEn+mfvcB0ztzTazZg6yPn+FGjEdDwR1icN0+ujIhXOqZmtRsx/V
RaKsVsd3G0imXgYQtAI9h6h3d6NiA7zDCfIYJlUbZpjEzvbYr62ZY61aMmyOvif0
C157JWXnmJIA5Qkz4/Wl6Pni0sJJpHAIRw5Of1OyiEjbIOvcgE/puQxHkRfT88Ro
44Uk56RhB28uu+2yQe+4uPTgrFHxL6Y9esJUgBMQKL9HrSO38W9IOnZOStagLodp
DTmLDah6+K9MEyNpAzK0Pb7oj55qAyeLe0W3lw+5QgA85Iku0wYz3HXe6r07O/7Q
x3Vb6QJ1sWwy0329lwD/d61MMHYLxBJGXuxA6AftgL6vLKg7rOiZ3R/PzcYff4kS
kIjxiCWmA2rQVEVs3sofixPzPU7aZ2K6VA+U8sdy3FesxzAFJv2RrVEsib/WGHV5
s843sZ1L9/BpZEoZ2IAucGwmrjE82mod9PuwAcFpNgNOOj8EGIOadT3XzUJUFubh
ynIQ675gy5bNLzVHZWeUL9n5tIJYdJTWCSOrIwn64IaXJCZf8XyQlqzkAcOw2Onk
iO6QxjEQ//uRcf2e3BpONkFIMbVIKZK9INMzaUHkTQ4l8xwh1BKd7vCcA3K928Wq
2ZAWqXIIfKhzR5u5qFvO/FyuyB9i9iuKOu02B8bVVonRIkASpferLQut3+6QOSWu
HV0Yk6r+htKofOkb8JjOARckhHu2sjTRp5DtOquzE04eoUJLMNZVw3rOXmXcNIoJ
+UAr9QcY0Lkl0ZBG0RXuY91d1jT6xGTrpAsIdqfTHnOAd/OYiRhWYLQSoHA+V688
HMZREC+8scsKgPgBmqWSUtqR7R/WfLrPHNIu+sDb6uR+strRr0T9GYLEc8PnyJ4g
uacxL6lsHoXIh+7pa8zGP9n+6ILcV9SKSrKrh9Lj+j7shjzKUj4EV8dAwKT6EZ43
Vj90L/doZda9Z9Ncgo2+8tmte+LFixIZ1FwwU2gF5mj3JFlKV7V/qFrbhIb0MBUe
/lJpzCtIKJ032mBp1GSblS3n5pVVnehRoi4/43OO5RDB8giZf47lbr+ZExX1tpuS
y+jB1c6Ecom+KebPI+ZiNQY8pnOKOk7pQvprjD8C7i6oZYJOeEfJpc1ncqse2YS8
jrCFm+wc91sxW/pm4cLHQNLAD7sun/h2NAaJTjeOrPN18bOwjqtWcPwFkPx5Cudn
ZZ0uLbwjU/MEld2qNcfqHKTi+DGSxxZk8WARQ2qT53KjVK1yrSsCkYnwf5JYsSPk
KcnDrXcZPocOhR4fMKoIFFOK7mp4BOvhxj1YmPdhfJoeqDksASAb4WOXYY1iJL1A
Wjt4gHJhVrn4Bg8GPn2gnpouxTrYi9wQJeYhZXZKbFYZOEObew2/Cpn0g5OTS6Ze
eTJCbRpttfpC0JgQz47OIjGbmhpIxG0hU/4uZ/c4LZu1c6XUmcjGpVzlvV2gLxEc
hZ3e4JCXNUnYIQZwx9CQ/PmROorL1ziVajGPdLmJCThSa6MYvjb9YlPavpu4M/hf
WXxAjS6eSgnTs/0mmAJ7BaQ4M0jpc7dhRYBce8rh+9xjJbFqPzgE4Sanx3prHGWY
GNlGerE+5+DAwHPs6i78/DMlvhO3UxwDrMrlzCnobBHXEWnJ4/JleTVHqhexkMf3
R10211xOHW7RRhpTLVzGeoQuAIO9bOsXSUCgRKkxiyx7ESOqng/n1YtuyRtUYiJ1
nPR+Rmnc/8naJQr/le1ski4657mI3lc6KWti+3CchEVMx+tRCzl6A9Tpai0PvK5x
cOfHeQ0Adbzt10FoXMHpYFq/zE80MBpp81eCMB5oTUiYQ/fi/E+X/idsLwTbE6+W
9waxCyzwD76fnHuIk71Ue7QwM28R7jH6fPQ7uGxPzmumzB4ioG887nOB6TSXdoKm
jEV5k6QH49zPYeibI4GcOQdIyBqkWtM9NhbCIXQ/HYJKjuFt8UKAZQ7vUkHLxMp0
Kd2SjTh7349ksXraAgXp0fEmdnbAqynFUh/S8oS3o5CuAn/bmonIhgMtRJhy264V
eYJWBqoSWFYumbfpd5no/WCZvAwGghFVnv4x+x4IHjgpNEtfTHqeNbhpR7r8Q9+1
EclGcVDOeqapUIK9usq8oDP54H2C8cIkL6AiFxBShqSeZS62hzMkzuYrrmSeLJnW
YAXShLJRqdO7OpRhWQimCq4pjymmBjLJKzvHqY5lEx9fVygcNIluUBylcA9RsHRr
JytZvj9GGw+Y1y3rLgMcaZUM7xykNz21thBPb5Dh8mtxlrTXUPQAK+N/JvDR0iAK
bRT303sg2z2WGcJi2Y5Nk2VYEc7UwgTtqNYSOZ2O/WI/eMqj4sbWUWuyD/amJrTd
YnjK+fjSQuI+km4dujdgtrK6r2LVFxddOdVO45+zUr+G62eVqQoQOTZFo1chKDOO
Rx5oGrLEHSX6KMAz69MdTcTXS+etL5XA8RL9XSCJlWhepxlKEEL7VY0cAqswZnyE
wkv/F9EafMAh0KwVKjbXRiVcXYpNtyQ++PMhCgTLhokesS7XGWgRYsS+CLwydqip
n3eq7Ub+bWi6zUa2WpDWaCumjlhAuMFu9Wu7fDX4YhA/sdVkNiBTlpVU8lX/Dbol
+QA0yjsuWDSwu7iNSeYSfUb+tnGGXVKQUzJBEQyAHA6pWRySpXnSOmc2hpykt4MK
geMLY6z6KfLxVv+2+jd1yKYA/W+YBPDsOmTZnrUre40=
`protect END_PROTECTED
