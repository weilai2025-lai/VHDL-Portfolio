`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMvh+b9Mz2awPQJyNcQvra8lf+I46II/9oIVzQuTZklphbjtHRCqd9qZeDnf9pCF
HzvxGg+psy3vrDY8uUqKPdwG8zxjzKJ8RrnSTFyTfOwP0CjwcPqOh8/lHdkLeVot
YclswwbBG78Ta20LX7gccgLSdt5yFFtNfsN0Grmo+0iKZLDYh6Mzxd0hZcUh8pKR
hoxWuHe7R7TyhKqJXw0F3to5jW/1y46jiGhJLTz78eu5ak0hPWoLGlJ7JND1xrf4
0fkq7GIcHZK+q2MqQPKJvBqTI77bf9hnFiQUYJqRmh2t86t+4Ml3ghM6sDqfr0Ms
p3zTL8wrjHRfK60ghHDPQ9GEL8fRaRGvNTBJsQ1bm6YETwSlim/ZDBYP0hHaTenx
VG+H27tm6XyAz/5bT4Pxvg01mKq75H5TPL3kZgzETO0zOY9ZkqKzi8oM1rznAFLO
I9E0FuyzHWNJMIE9R/pGh84vdqxgcMDaAeDhKB3WI//gnqkBFGoLTeFMhcj7j9No
n7AXXDOGLPEHXeDmxk5eJkmtDTLuy3lqjdRp/h/IZXzH5CXRbwW060te2t7sLfXx
o12lBxbQkK2ucJwKGzCLcojKfXyEzrxpQJvGYfxIZvqIxwyMuiq/DZE80PlrC6Gj
8J+31k+jleglSQLDq+wYBym9Y8qnCB70niSvac8+FwTgRzsj2vuwPzTo1T7F/sk2
LNbRZTTJ795NAse0ubjnBk05y02myIQJEwYBL9iN6/bsQLzTfPSvd8fI6gvWd3RF
uJZ+3iR3xCv+ExZiq+cQCwtrcDscGsJCsq6vz5P3/W+YY9ZoDHBIvxdz7DGLWvIN
D/jdFxsfMLwDYzEDK1ja/DR/HCUZ2LdemZJ/TkI3kjO3LZZ8HAS0PJwCzrEk/hdR
3vdoqDHuZxFHTqJwCFRIHcUA85dJCUSP393ONer5SrxWOFrlgtHynQXQSJVsBTrZ
Qsc3zJX39V2eyUPCR78bB4OfjxvZ+uQGnxAbRVmJE8klXWjpJ0S9fIr1lrh5hZFV
rqmmHnGejbsYrJc77CHwgxHFqyakopopksFD2eZ9iEb2/kD3mifkkQdbBV0zpYtX
i/KtzOyPpZmMoerS4e/T3QxGUtLScQ9ARj4dJ5AAyWZX5y23eNG91EXP+2i4CXyX
oI4nN0PJIVmkx/pRS6UAI1vQUprmcnmewPuJBZLp+sjkOVE7M5xvOV7vybPaYaHq
OBXmBOYM5RB2/gGZB83P0/LK6R1JRgJEhGs4+oeD1Ac7/6Zae60UXSok9t6IFCQW
4/S6DXLJUpxIRzSOmZnLvQsLnu2a6+6yPbEtluWzBUAJBCZPnze3VUI/mUTmqVZK
JEK3488j+VCN8L/RtA3P6KJK8LH41+41jSfb6DK6XmPN6DS3DuewjxrgVhKeRDI0
jD1su0xvzbqsZoVG5/guazKsGM3FI+I1UvA4Daj/eGlrKiJfOUpipf7rsq7aBoNE
2xM9kpn4TZmJxcGX61HyghA/y60zlhijJeqKJY/jXKawztMWYlopFxdKDZgXo2iy
ynoJVZzCFYPrUeCHfwPjWiV/8QytJMBU0DVd+OGh7+CvGPrqXJ4pgaizUQ5imvZX
2XOQ+toZEThwSLnp0Q/npKvygpS/6znKZRKIyd73TvC+WFaxIa0r9aCTgKqyYOr7
Jw4VGaEks73ukNJ7lkPK0fur9dPI6An5eXLPA1kX141MOGSwPgZ1RqcVEflB8VRK
0xckpcUhzorrujxFnYFFz/CdpYKDI0PGzmqgA5UtZKf6ZxkslLq347bX/C7gxvUL
V7164rAiFdt2SXAINwi1Eb4W3ZKNckeHsiSJcvf3cQRrD5SX7A8qkKZNMcBOYkSc
xFYreDX4AmKTCP56Y4zzZ08rGapSp724tO4SCdeEK9T6Ts1jHSK6pN4vKErpMnxM
THNJcaiYEbnh68QPMdVo/yK3flG2xRlTYeEyyb3rSlEqdau73zMzyYR6R8fCd35g
mksKsxi2ajEYFh6LOiIaQvFcBxJe583V2Qk8J42A87Zydyn+v6nx3RsvvgIQfd9/
TiBkpaFpNCt6reAQzgB0gubo5VA8wxxH6xYTo1MQsG4iQFTSVbMzK3viyCIv+P9R
K95IoBEutD958ddT9ojJXEWjXW/+C9ZudMYgCcHKLxF8VXVphcyywYYpEf4DxMbw
rVszQdPALuhlqc/OVWwihwwWMFLsa6GyJ4Q3vHOGhR275UBaEG3yoicYyqQaKcHZ
PaUIIMfYIG8eZY4qsICU6lnUjInMmuoi8Prd7/cAZQPWfFLOOpd0UQzB2RTNenwf
juKN4ijQWO5GWhjFl/Ugrg5LixvCmgy8zCaX12bxakO1t/hpOYhoRQqDLN556NGL
qxupZN+TNrx6zdGoPsevWj7IwADDUA4wjOMly2vCudcav3tBy5rv2yZ/J+gOeee9
GplrLBoTmHb63O77hc2062WfQJt6tHpYtnbUdMlwnz30NFv5qYr8bkhzZEvLa11Q
ajb6QIzWCGJ92OsspRW+YXtD+ZMcyY+chvv80R01Yc+dKzNEXGMNjQSWUBmfBuHc
+wMlo1sSiyGbRuWDmD9aeT2d0sMLtVkymG7mDBj4vZ4AJW+BeCvYLepiJd9OW+ub
1pZH4bQUQn7JREPvrNEEwQSaS9yevgeO/pluCkFfMEp3VyT0MscDxA8RiywX0tHE
MGcLjwUoMyGOVxRg80JkkglzmTIpURnH4CT2frBAUa8O/aN9mJmuZLQLoh8B/Bw8
Vb9NmJJB/VzC07cwDK1aylAtxT3bcXFD2DVbdFsKgpbTGF/3pVBv7zDsaG0IzWtZ
6q/tu8MpCSlGUqU1JbD0QvVe7nkYV4NQbHulzOmhzc89EzIUbsdFsCMu4/89x0NN
xlYYVSZn8KANMilhJMZ7oI7j6x24nylX6vKrbWzsuuQDhqZCHRVx/jefiF2zJDCW
vtszWAashDMnnQA/3F4QCxRUPdex0yFcQjR0LlloJ38pq0EcC9gTc/EwSvWDoN2T
z8yjhoSFqn30YflOtMwVq8fW5MxIsm6/RpFgXWRxEMYkc/+4W/T1y4EEuO4fDn3/
LYIxgFYnNEN3s8Gy1hRoBkQLC1GMh4rBXnrkVNNgRSbgS7Uapff/0hwQKElc2p6T
hdGnHwlGJw0leFO5P5qJkavBEBSNJTHNjklTf+dj8V5OMKxVfOOyNzT1byF4sfPp
XTFIobInI6mZgkomuoR1j725mIlp1qhRCvZU8fKoKpOu4pMx2GLQ4+wp54aDrShV
+td9cw8d5kDVUe8XZ1rjbEhrOpAAKtr4CdDvo9nAGCs2OzOWwhX7piztEXvFg3aV
`protect END_PROTECTED
