`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqNvWWAI3OfkmbHlHS8nLwH3wAMBKv3fRjRLrZWw1c3kNdIStXVabPALAci45qnz
oOUKeVizZFD5M2kIGJgzwAF06+LP1GDgJvx/KaklMpgFUpNTDVdW9bRC+RJpg5YZ
+kb6p2oRsgz+h2uUL5qRO7R1xh9tnOVyYE2OFqtTzstyJheafvKkNbCQozyuCm34
SYU6IiKvevxIBkMTaPg/tADlZfkDbRp1dDptZnN98TtYTFNruHgW6Kf/8kurndyS
zKLu/EW6ravlwLraXg7Uq5eey2otceFCyckuo++aBlqV04pct2YGbx3rt3SX1as8
jJqK+hcoGmnaNhIsD3ofRW88X7oPxJsCWX5OfHXAyw6CkVaD3bApvn8QP3Xdqrh7
NkW4EOIRIqhiuHd3RCZ3cm01eJ7i2Jp7zHB6ztXvtY3WqhltcE26cwx+A1DmRHXJ
uxZHWGshX7ZpRyHZQSAeG9b8YRqmkQnVl0ZWlurkiEcQDRmujHf4agelO/WOp0tv
7OFCCLTJFEYxP/ky1GpsG27fl1Az4BLjfESnrKHExp0LH7QfCfXn/uXEApJlJcwL
o31lHM3hUfcXcN/ArWSyww8j+lGCABFfo99mtCVUhazZEEdIKvre7IYCRBCYgbhU
jYfjHaqTY4jE+zsmr04NOM4BfY/jnYw+ZZS5zNXxVvBNBzEq4HX5niQFPno3frgT
bg366o9QLrO620lhcayP+WZkVxUoCSw6aKJcUbr1Oe1uOlWK9uoRlV9XImgWO9jJ
7N2lAtlgzlD5dYo9mnmnF5n4giDBuQXDiD8G8U5BRyQaW6Uh8efasY8I2o6crJaA
5lbPrbNnc6ZKx8AmPWlBKL3oBeGpAFWFmJYfxzYg5X/QdAUWF31LHW4PXh/mCm9o
4X8yAvN7YWrq2Ab7BeodamHuU9+3TuOsP+yOVqU6fp0UuuLDf4oZG8GtwY9pSnl1
7EwZ/6gP+mj1P4J7OYqpLkmzsAsBue87tjPvzcnmzOa8L/BOwuRy20SprSEbEK/7
svYDiiuHPzNCFymANuivK5vVEz8E1LRMJm2TmLRbnWnN/q6BsEdnZC8LmRWtCK1Y
CJbR1KKtTyG6X+EbvCrpz4ZrRMyijtG9pO/x0P58R5kIr3PtNhNo8YDq0uShVuc3
SiZrVdmsSZyCo3C0whAY/uZr6E6mXoiZ1dKZQXaUep//Yqhl+Hn9tL0TH6chOZFW
/5M5pmREZ9nfusqzJKyOJJYy8W6sX9yuErbA9+hoyzQhu03tDKeybptv2k6XzHqP
7wI39xORytYouLYbbtnwzxsovVhWBIOBdT8cr490CyEPTOkiMLdejkF4VWw2LnsZ
eHh/VJu1hZYHhSprVDFUlDV1b4GP03vX3OZ+DraVAedSwNmn8IQlEE8R2sKiBNfL
Qxw/WjvG1E7BRVbx6P87WaLQ7w+XV+6mVwZ4EYyxfSGBJDaPxqJ0q2BkEdtV6dCw
5oXMPi42GAnEkRyHyty+A7oA5O4RBAtgkslWgnJ6m9Aq6LQHP6MDEVWq5lOXa5K7
mUQ2AJZSlB2aDBB2/GPA349KVsL2BNd8oKPjoz5jC8FEYm958plHiTHbymhqiAic
Lj68LM27cgmPBpBBNw4UAntc+H40m2EzHIwexhBroXytx/7sMaRnHvkvpH/Zt/tc
mYhAOTCPErKy6gfoLYbToDvpChmJl4VKy+vhtOj5yN3iouxzJorWcTWwLW3h9ftQ
FGAk0yIp7JnolbEZ4NKlTcIJLqChS4Nsawbpjt4OZSjRrfAR3mLjQSsZSpBfh+y9
GEPtk9jdrp64d5r06eLVyuJMz7HO4sB7KJwGDdQOBUpmOqclBU0SMRKKGpyV/ZSW
2BlQVLZeCXQ4rn5XLroSH2DcSSIxyK0ttlWI40tcrFNTUt4yhi8X5Q6Mt49HwPUv
2dIEPymGty/vo9ypxWhbQiZY3f3r/FmTuNBH50TEgA/zj8+FETeOY/YlTCidmDF/
OlrR7iLoFjJ0CQH/IZ7naGytE89bpdWhPytKMgIMsTZkunaa5JUmjybxA0n6pTCx
F2LowlwNjOp+YSqFoA1EejSJrNmwh//kt0CCbEuywqS2OYxOKsJ/25okkhBDZxTN
k3QOVbVA9g/OixW/ShnDdNAfcIw/lG9h+EyoGNkDWEmcZ8W8gyAOi8mmy0m0s8Jw
jinF0k3uZxkSUDrHNv0ujG4K/6mcyZBq5+zaW/3jynkyfhhSQf+opy7cJ2b+m1EA
Pc/wxdoZrs4VW+19k9O5oPZeyaRDukqwtJ8A8se52qjQgUiJ7LHs9shc785ZWxpP
gKGSs0pUKMYhjqjjjYIUA0Q1T6xqs/Y3Xw+qt2SV4XzjEj30JWGAQXZybhNazioB
`protect END_PROTECTED
