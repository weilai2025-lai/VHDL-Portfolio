`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raeBItPqT9lEUyw9T5QXteeAHoet3AAvuKkTCwEg5FdYmfSvedWniqRRhZv+MivV
MMfNJPoMOPVSCkRjlOV9ynTmrVr8iSBtZ8NsFxPPSms8NeYhVQsp1Xk8FE+LlUmU
09bx/lDjam/XQSeJ7cHdXDNUOw4TqOomQnnChK2C012oKgBjWZZgtJsUls7JHQGg
WwS6IJKjy0P91bXaQIP4sHf7g/hzXMPThl8rPqjl+AeJffpLcshFtJSy/Sz9oUXY
auF6giXeTwNnob/ozSDuvEG9t47vxo3/ARGHKYfz/LQ5DVcn9WRckc3JiITmsjdB
TcCu2FIl6BEZgIIq2dtuSh3aqaHGtqd9NNSQQaw6XV/8gj7iFmWn4M+8F3JYU/U7
yE6q92pRhPKUzZvBiKpTN1RG+IyXo/OFRkMaXGqJIKsrjhLfrENDFLAhY4YISdLZ
j80az4qxWQJb5dOfDFbu8wg/g8d7aRPxKzNrD0yLT8UGymrZaPlHFOBVwpBTxH9m
c5/vK3+oYQWGrlrS4iSNC6Kr2qZOAA7H3iB7dUdPdqe9VQdyB5cswsOQx+xUimHy
ipNr5a/DNmEUobe/VvvAlGuoKXddOEYZ2xCBhlqtinOD/qw86uVTmSTBFTzsvBYH
e7NMoZdX5+t4zviwmI5RZiLUAEMFN1588wfQnjMVi7vubHEgdszoHcvUs4xysgAL
mGLikpxcVFMqKznEKoZuftaDmId2Fh6jWHg5aIg6BiQ=
`protect END_PROTECTED
