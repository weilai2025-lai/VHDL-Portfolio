`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldcWcG2iZnnuH1cemA4+NiEhDyy+Poqd10SUiiq2aUnlhUj6n0YyJE3yVoZBt8Dn
EXFmbOXPcWx4MXqB+V7fj1YJmXwyzorLxzZtoYBJBEaJlIi87n6T09AefiL3uGcB
PSf7Ek2wt58Noq0sS9L//w5aUBNKSBgWZX+qfy0DiQ+B2vewKdMbNYs3I6vEqTEs
RSDBM3xun1Uat8md0OuKc7deffl6mmEoFTu96Cy3b/cX7Gto4vuOXK3D5Toias4/
zKBxiZ9q/Yl8YGx9Vpw5VZijxsKtPVxEC/pD/1zfPplxRhYOJPWapvPZ+kd15H2L
dpEwlfVEx3QnwmKgxrKetxwZknHo5VcCvMxEIOyf47yleFwdGnjqVodHQ8ch8ATr
XlHV+KDYseUtVBTA6KiZ/Yo9x0NYsLUef8XYiPD9y0RQpBXSVkfjgiwwh9Ce3sEf
mqXS+j1kO8bxuZw3frIKIf67xL6Q+M0gcWi4oqNReOIyVB+hkABsPuLqs/GaGKXJ
JOCD7O2pREiTV4mbhul0leQxC5f/Km74d9N4bFgLH3yX60YFlzouUUGxtm3LOg3/
84p6j3r0olNUx3nYXeVsE+SfGsmYxK+yDEjdLPyZnlpajEw+E8TY2eSIvBGsbol/
1ZxhGA08BTGcXXa1Op0GOfSuFqYfCRsCuFqeIc4bY0gd3eBgP5+O7Ha7osRaWBAg
OtuxeC9fkeir74wEr0MJYTALh4+w48Vx9UHlNMADiMmvZJK3U9S5Ke0r8i75l7Sp
YWQUBVd01sjSg0xVUyFvbqBjOn91MGuQ8N0rcHE3nlawtdyFATlQ8zInZ+9CG7j1
6QLY4c5noGsW/guHYgBY329+4YF7Ls067kgTlUtMkJLi8+6mRbrCED5XKqO5Hzwi
4BQR2mxHfSgsW7K4PU+BPcJIZMxnsbg1z4WorW0BKcyDmQ3aZiqqckahtwIV1VgE
TLIaXeQjxzrcn7knthQiQ+xL1ysQWZ2q4YodtpLemRM9cNIXC8d0+6WBTncI/aTz
7zCtOYafSaP8LuSD4uXh4wkCQVdUu2pK8by0gQl0PgPkT97Ve8OapXCWPvY8qja4
+ErSaL+BuUnsfMoEx034c3ZV+id6AWk02kYoQjETCvYwigFCNwKrr8tpok4RBqNg
GK1CrLf97uZ/cQQaqm3AxPTe1x07JErjT7hwnSbNNTDVhJ5vqSVBO58VPw4S1nv4
QCw3DEXQ2kArqGur6pXbwcj1oiGVAILTLB0HKRm3rM3yhNBgFjUcBnIZnUgn94vl
LvH+qZwNsUKRXF89b/Z6K8ckQeO6pikQNkg1MImm0LcwejbzcqCvuVYJ0TV24nof
GMLI1Iqqvn1esX7KIT33O9n5+sWPC9eOKEROgtx7vsUum0wNNlGu/pNmbT/kjx8w
6Oa/qn1m+jLwybOlrsy9wod69IJuuTLyk5UdC6qNlODPIJjeFCUkQRlN/LuDl8f4
CNduRL/m5oLU7lGofVecReltcPTy0f34ZyQBSo7W6sPwGDFieK5obth2ijn7mS5J
WRrOMlfdoEeTyQ8wq9jq7JT/zEQHsep7uKeXs6aXszi+iIfL33jauZ8iCnqavRPv
GfKAXv+igytijE7jjE5ec8NKBSXjx6YkV//3SeRV2IcuK55F3BpqmwMsCC5HTu7u
8moDgSfrFOHeu064MfLwBheniNUvtMp07YvAfTf2BOP+d94vj3HxAzRpY6dXnsbm
JRq/Uw3d+OMqgVZtNUZqOYTMpXK63VHbwKLaHAVyqc+f7ubWbsaW9y+W9/XxeKk7
C8gXqcn1BZp0p51r4CQkkL+BKQzRej4lc7O4MjEprlrcZMXuwYedBvOVn9JgDQvG
UhJkLx4kQ5EN2K7du3Q/jAPRdN1JOIvMt9V7K6Yvjz6KhcsMzsXqzpeLjMpvfkXG
3/qHzZreYcjY+Sa+O4sDjxkEMoYsLsNe1DpoJ8uMS4TGvkYZR9vsJx9XDlMhJcaq
9RWjI1McztgYlEjRuEoRr4l7NUf/46gn2XbVZU8bKMM7eBLDZXYvk313k7BxvAOV
tNoNfwQ+o+8pT1YOjlePn1ZQzYmy5TQHDs2T+/UEEBcTbCaZ/aWz/Q2cCP/XVM1M
A/eBZgkw5Ekd1AHrpARdq1fMrAVBE0UPeHcOMsqDE2iOQjzgrKqWNRgdAVRvowej
Jn+4Sj+xtNyDcf/q+d1t5LKURXoC2minepdI0wYeVlqImwLNu29WgegeKNRaDUQ3
rMM+B0SlTwD/rPqPorSBAUVX4Uqdx2+8bNcCAPNulns8WtQkvNp2Qz5L7oEeXh82
4+t3Imw1ObfgpmB2QNWi9/kJgTKxaIQM2cEZfaHMK2wPFMWJORwq/VhELdhkk1jl
x6UgcU2f0ID8qouTzPTM7C1M3e+3Tq1KSgiwFSI069GEIJXBvh3C4EiQuOGXVGgq
TkQv8G0BPFgCwXxGC/ohLCTzXYeRhu+WKKS7+pth1dvYbfE3ljKxwkHW3hBY4L/m
P/lYBlkU1OUYFkFiYxZaieIXMRDxwB3F++2lIHQO/L1dCbGetR6AJVvGWo/BlCe5
J8EQhTRiuhtu5X2mogC8q0o7d5tqGcee+FNcrK5ds/kGkETFkOAV1LBMclBlRh5i
qHgcDehPnIvpq68axvYcmkWQrwY6OTqBaG/S79jjU4De+YsypOU0Me6/wrByHlGi
WaxuH10QW+P1+gdaeIIE1rZRBd0mx8yHDUfWJZiQQCS9TeTSCiFzsYQV4fEcEG2w
JenWocqqVpAudsTVKFgUfpuMkV8iuyRR54HN8nAY9b2Y0vXrjOGZKWfvHPjvTYGC
A6X2t7bICdFme4X3pvwiecCO1dNRBEaXbMomvdXTsfpgBYijqJHh9XlYo6zZq72/
qFWxnsvp1llJdCehyCqnKiV1JtAoAkhhHvW3j6aTdsJdDPSSXt+i4WOK/ZUos4/0
nk8eim4YR7xhFgrd58W4qVCed39w7wZe4VTn9sAlAABjQnbUo8BJ2ba70UetxrrD
j5bLXx+mARTY3EQk9VA4EDcoduPthb9/WwaJ+i5d68DpsB9XNezYg/HtvB5G3JUv
9uVXb84J60EO1Be/rzHrKL62Np5jNkyOqxH5ORFokwgTBztGqfGf6AJIHgo4HcUS
1v7kBhL4bQjVm6gOMvGJvZZUHlXYvpiZAOEKKH86+UhZKAr888bpesnjno37oqhO
srPB9+H9BIB41MvUv2ZFi39BhxGmssTYtJQwU1HE9BewhSy3b/zeQgUlkgWey7zi
WMxewe3ui2pnrqPRjCmVe5D9hsejfrri1foPzqMAsKDN7zDAYPiH8AEQVbi21fj9
D045yi0RoABCJ0/lSfKNpIblOKoW3aJk5raNthpDXkKVp5o0x5LImBEVT5bLrVvg
IaF/uTa4jukkT/tPCRzm/DN6zm8BiTaPDmtwc+4D4tTLV2T+DDOBnJld764YMhCu
1D1B+yvQS586oHZLmcrfa3SRrWRaavqVbMVpsXE2fJvq45BxdpICZJjO85sndLGC
GHE6sXDzOxKmDgIogytLQe91kqBia7qkv8ZsLdcAAlwiZHD7a1DN5plHH72caIX6
cOYJV0wk/UmCZuTvdgVVvSJASJEBmRkzpt5yHsl3v33XN5H8qIuPg2Zs41uh/fAu
NSg69k8TxcKyWsJu4lSWipAXYhLt1Rc6j98gKTaz54ShlIgK5iDqd1JD/DzKtcPk
oIGNTRMjkrgBZzAQrqs6ZMNL3832Q3q/wB3rHiNo4lda+cO9XkNNbqERmCiJ1PNi
0xNBHj15eBtLG+q7lhyT9wDukW+45vvaKRJAzESq4GFxteIBZ49RQEFCNX5X7KTD
7wxF971K72mFHY6NkrOr8OARVIxeu5VgX0qTyc7wjJTIbJ4vBlXaxIbrEE+YXfol
Cfqk0ofH5qMHFyDAD9AFpfBm4GezrjWF8T/9nS8wFVCk/fAOKE9dLE0Bl40N8QR3
sqvvI+syFTOLUy/78H/2yFoDBRGXUSfyf74N7F68BppSLFizFsrm6gbkBd4TcKVG
GPQWINZDGqMKpiW8DAJEzqmx0SdnJvgCnTl10ORF5AvM62Q8AlpxLix2TwUySyQH
ebcYYeekZRsm+O7XG6FqqgQtgbfzi7DPoVbRUjBzqAcea4U2CRc8GpOR0zlj8auM
63ZA4+ew5WFMh0I4zSzoPBqENdDOCZP1m4bOTCOe3CqfxVNzq9oIECA08TySDUQ5
O7N0pdhh/A9NpScJCycNO23U50eKWQjzytgQCr4dIk3QBAktuTi51v3axzH8H/pm
ppgyIxKbkB4m+zGB4Z3gcCbuRJ8AukOtQATpxQcV2LgAFGagRVgzYpmm9e422Ibj
Na89AXBdPS7yHA1Qs6bXcPujCFylWczs8HnEgw6jbKwWoUS5j6472kRSXch0JijQ
G66J/PD5LDwSBfAv/lOfg+B9neqz6WE/S6KE72Pz4ipj5Wou76qLq+mbULR/YbKL
VzIKdHom58fSQdwLWuoGP6xLiZNJCLCmvmQlmcHhmZm+vEb5S1AZwbKgk53FeY/S
gHgthePiXetAQ8HZ0+ZOpUj1lUVWh17vgqaZlnVW3PXobmOPm+xlfShnH7ZsWtTE
T9U0ICrQB5lZDo6vjfGujlY1h6NpI4Agjaph5I9EecHtQAPhljRkecEbwsvV0XEd
9ZQGz5h1Vh3EFsnBj04zK1o+ke5roI15BJLeVv+eek8NHovy05pqtO7ZWXKxQg/c
RkDwBOMa9U5nOV5weqM0Pc/zsXq6yqRNb5UhXnBUDQX21wKLuOKiYy/jVYMGBu4N
hlvcGeh/pXFDxk8YjE1zIQvK1u2aE6bzkr+l/P5MTgV1NBAc1rE+r8LvqtvtpBCZ
Gda+WzuvHpvYREiNAOGGJ1A93fkFT+PttEUFHDEDg5batbYT/+ktkitW8uDkjcDo
7BC16ZJKvvOa8reCTat6Xy0Glhtbfi5ie3rt32bRJj767iDL/jADcEcUpKmtxEzi
CimmITv9OUZf/nsuX1ybHyds8WF00Kry4ZIvKNEdHkBXCAzTVq/t/CgH9xhiTwTi
5/6sPuUP9z1aM9bnZvtLtIfEu+hg5dpqegRyVKBXmzWfsSX3piqaTYj0qrI0rLW9
0lrm9lZZ8xvpTTRNHSggFOdlSqW4BAFYxD+4i/55v+sBa55yNi8wt2/j2gTObz/E
g5Gq5LdjbpkNFcNFHAGjC88PFuN94YPJAQwE1qBndplavs6/pH8WejMLHELgGQHq
fmDRBv4j3yNp4qeYLtVdO1oZtnh64irz3CRdBMcAkPTGu3SeN7IRf6TdSDkSikFs
i3WOELrZm3V4BkLTiQE5tuvBgY1FN11GfpyyRDu6fW//Oa8n4E180VQyTSwaksH9
p9Lss7J+/1hJcU+LSKG4Z5Lm+wUnEWCgRnGF9cvBynvH3UIRJd0Uf3Y2a6nHRZ7c
ipmPkf/j1tFyIir1AI/x+pf11ObQz5ggc6/wvtWySlvTDAOr6TzaDB2IS8D+FSLl
htlrZ/XxwzWBupXuLpHAId42rG798R7PEknAv2ncT88y9mP+ZVccErRIMEvm7l5F
tJz+w2bt9pe4v0Yl99O4hjNwun5EhzJUsG/+LOoYeeYwflRwu0t9GppVOxQvh7gZ
C4IRPMXYMJqIQQswp7epOxLsBD8J2idMmRGyLvwoRRmy8vhX4XO4Xmp88y5pjPj9
Ts0x2XAQFq6Y9ovhInBYjwsFbYoOcapwppu5I6MdsxrFS02uPV2mBdwT6umCZ1iL
hwA/xf81VTpGfcy28naezPDD6gPOAA9IpBFIOKPOevkNE8NKpcXwlKqmjSUuu06c
arjRs9ZdAZ2gSBxDtZB2xzyicLlDNbKMjwsfgZyqjxQ1rmlcPiV3R6PoqmBzFy0L
qVsApRGaFxaPqIQN8P0Gry208jcp4XGO8Wfk1iuPhyEZl3P4d7xHXHFIkD48ldLe
XlquxfQV4feLgf55iSGd3wM9m7uhKbM9KwIpJ3Skrv1r5o4e9VOZSY11OXE+Mvj3
3C/+/twYjQoEL3wWtwM/TVXwYOA1UW1U2T9edZvP8XvE6sGjkSHBnANnMbJYSMzg
5+pNQ73oWeBEyo4xtMcaMZKx30LL8mCqbaSQllJjZ5GpMHeILFU87a/64ap0CWz+
Jfj9K88+TVJ7j9zW8ipteXKXfWgPrQkPa2Cm/bWDJqLriuAndnNHRF7AP0n6Scdx
vIftHfq8+riJMjICpk8Jzght5oRZCmsFl9En+Cj0agHb2kpFIQapJreer/ta7v55
t/gg1KJ9iWyDNaXIowRvwcZ16vdxLUNY3xTJC+6o0OdUXJxtPz4y9BNnMrF/HOSE
x+Vzwp+F8C7BsfE6BnJelTWCYbxRuefmn7yfemFShtoqEUzMKn4/Lc3I5z8kdAy3
e3+nfKXVJBeo/kh0C+ye5S+SXpHjdnbARBVrHkPyI9d/Xm9+OLdwLE39mM1dg/k3
jnTr91R4rkJf9Z1xU04Spt00anj2PabOX1316L9/z89qjbxOky/Tt1Bh9Sb+nxbu
Xow1r4Ut9DgGbCt+IWtC+EnpVjunrcCIQzwOmUb8GYnOS0IpGeLTxJwRED2eqYUo
tlqr5dTBuIuCsdi6tjcLf8Y4XPDUb+U1jnCmNr6LHSFbiVw3krtJoHYvbmo2OzKn
Flwp/M/BaoYU1+E+m3gTogVZ/oVUcNbStnluBPNJT8Vbpv5gzjoMH3bzGT+Z4mZ6
q0WdFVQoD4UH0vnSLOCmNSj1tUxLRQ6Cc+bsF64mu5+sodrPri3H7wW6BItxWJ+U
df175nM84+Rc5UZAOgFtB4hRHkUEq+PsWVMHCFK7X2h3/EqcEfO/jiGDifpuC/Iz
n00XUYCpOyjYqOprQHjZ9+4c1yFv7gAieYVTCAbEfSeh3xW4rWpO5U3YboAvRYMS
xB2ud+RPeF3AIYxATvtllzfiK386UDf5W5MguKVxYB0jAu+kQvT9GXqLOYtlvg+5
NIh0MQeP5c5GSYhRBlLQ6+PiL4ofhlmP1gAtXmh2nIUMNVK82yj999y8g6CWBRWG
Eoo3owQ3rywOzkRUnSB+LXs4mmoWU5sN/tVBJO2WHq/3P+k6D1/ZPhxhoNixVEmI
+ULQI4PUqbBjYU22vvc2LLYl2REVqWwjdLr4pa8NhzMflCKQoVXS5HPFHNJzQzFQ
LqIShqSyAn9H3tWrO+DvOxYyiTw48fHyKJYqVSlwoXPS/WIaRB4WBO1JBCFuo9fc
xgB0MUewQFYKT3jgdon+1cQ0JbWBPY0aDoKZaJ+1HdAcX/yixRKVEQr75O7p/dDE
VZU5ZEcS2zNLfpLY3MWbaiOIGkfmeHwta3D1j7ryf/OWTKRXdjZUJ4MQLo1+Jl7p
3zUtq8aQMrSqgZ0UQmP2Be8B+L73YWR4EIPPVXCTgUP1Z1todxeXHvT+95SD0ckh
detPeIMIhfh0Fj1dYOFL/zWwE3PQnHsmYHcBFScnX8rLb2W4WC2K+n+4+HH2f+xX
ZvsHhifj24U6HDgW8uObJsY+M7w1oPoQF1dHwarqpUai/J3wKbaTyLSJPdySEwx2
pXPGkfvzFAYxnKniu8JUf1f11wLYwuYv3JapYTZmoKYQjTAhlAFtdkcSxpaIeIrP
amNJm5jA4zWQZ17c+uFLNmgkJwbDfmhMgIVoMSmaJqX+i7xrCx9W9ojD8MQPJw5O
GaMyAKVikQKUq4uGKRTNe2p1Xt9w+dlqr8SXX37hxJ1D8ni5pu0TG4Y8CvgdH2gh
oIxC02Gt9gKhBgzVNqIdT8/YBfLgB/A8HVt5itA/RmB3u5cwaZgd9fM7MTxnay93
Z78+x6fQjSYurqg6DuBCtHsH/wg8kxNV9MJFKPMsd6sydTiRL/Vy77BoCaHDeNxQ
JTBT/B+tEkuCZw+Q0q12QA6ezwuxbLggcMUrl/Ed1n0qNvSwan1thRRNx8Q+koY9
1BXGKimcextS+AoV89+3lK/TRNAf3uWHrb5GDVPY4Fti9D/LFjtsgdolAD2dcg6N
PqgrvSh+3EsPFRLA38qnd3SBBTlRUGkK/BPFJDzKnFileqcJZ0aqeG0jUxwnFZh8
nQHVw324QJKXfagvllxpQazt0ZYktQLqJroKyWzixR4Om37Ljmer5YHC3I+XhS+p
q+F9mQaXmhNEWwTZ8yTTT1yN7owshjoB959N/pdGVjaqwnKoMLT3B291yTu1AXZe
cnsIXPvuWhcIW7DoJbbkiCLYESfdE1HPPFeVolBxxH3U3QUOgr1QwcJNhTih30tx
9Joah5cO63Gd0McNA7wk9XNx0+SsCJHzBx/VKK40WDiQEf250iw19i+frQ+egZa3
A0NQ7ca9bWl1av+kqi2fLYB4n4sIGNNhEm4f2sMkPPb/pfV6ELgwxdDam9H7qu3F
UF4M6WYhagpC9GG2It0Tnyl6BwUpbeNLJaYn6M3dBCmzgytFSsJMJC/uLp06zC2l
0gVSkbrBKZUj6rCp7Qk7h412E7FGg9QyZhok5/Yz+vtSI5+hSc8OoSs+EKM97yEW
5GmaanAyoql+NDk2lawQIOwM3TJ5imVCxFdNEm/xkV42aJEVJ4+2Jsib1hFv3Ulj
Pc5E2ln0OXUnOLvosseSkFC/yeNS0p2B0ZPNblhZz4URfvpy3GrzDhgAAEV701De
KweWe3kUcj0BdkEUT5bGaXI8dKfHPZa/URNmVIXfuoBAacBU3a9xHoVkAGhHvbN9
Y+8CFvqYVwmM4khLwNJHSoMxa3IymfXuZzLh0e5SCg6G5Iq6MgyhWe4tEJ+TwsyZ
SUCGdE67vF1zK5cUPJ/HLWTQeUCh/PrK3FCnYk9ruXqyQb2vjgnPUzYR9QpwR6WK
UgMXtf3DDi+59wEc9OasNwRd/ehuu2xJepwUVV8QqUOFYHJIsh8BSXSgG1aMCIaE
4IEI0qXrHMQpdr3jRxr3VzsSWHI8T8JuDFHrTWGun9cwRKyrMb88lxDpM+HiaxBM
6ywRnBHZ/TJWvucRcoN7ZGklCgUuVSU8ni7QOOkGlFfL2ZPO7X8gDEpbwIk/c/SQ
ZW7PSro9QgP0b1sJg4IZY5owcqMmzpfeHE2iZBAmT8d5z5g91DSDfxQS7E22R/sG
Zis2XQlxdvUoRYxjcmtsMgJMp7feIG0FjSywitjLqeVJvrO4ShLup2v80tNK5a2E
Sj+xPCj4xZ/BHAAF8p+Z6jWROoBeARIH9D4WtrdnYQMGS0kdlXnaYLCqWQjpTPmw
s+fmwjM6G6rQN8QrtbhWf/GzePUbgWrP16vbTwKQh8OLQQzWWoYmfR9Wnybkq31R
al08r9+ngPgYbmx+e3CkO0d5vE8bwkekdzcB12cAKPGjma6clt+OvR1BGpr5PrSD
IPn/dPjENpyh+MEL2utL/+PSR1c0Y0VwAmq4afgALKyPQTnE4VuNwPbG71BEHCrF
xJSWUHnJxnkxxB8VvGKIfuJBLrZIb7Ek9O/K3/Hq5HIBkmvSSapsCJmXKtZnRiVt
f5VtqKQsAcGvfM4kbN3qxyPO2niNpc/9W7ky7sZM11HTAc9NxCnNsfj1MKJz/rAG
7vHbDFyrfcKWkq60bJeHYI7xwL5bVVO0q7Wru7Z7AB62oc2X5KLbd0c8O0kbCy1Z
lRS5P92+AIv0x7e0mivGSIckab4OPQMNycPx4kVp67CJlYekQeuS/6IRY76uh4tM
b/1RfZMscBtrdaNtYitmMDTSwk4WX22yE6EVoIPG5wpoTUnmqlz4yPCQDo2fROW+
WTNtmmdskzJMuIwczvXWFH5v2jFVGWewTI+gD3j4lZvRi7MwGj6raE3xYQb0mYdb
U+5XfnSx5im6/2EeUWI7LNHp46e2wa+h+o0jKUW1YpIqb1IZhzK1MmIXJB4SHuNl
4pma+3c89bDrWaIE56/W2EHJrlws/Z5CxwDhlzXtQ0LmPdAkI8PAnhCGyTkSbfmX
gEYabaLsg4FPgr/yujFUb4MhLJ4BN/dUp8BLlIBCl63NlyNsqIeQ4EbnfJsfF6rk
MNnCytNIZCKQDHZqobyPTTjeDSkllUODbIPARpOKefgoCGs/rwFEJahe0DV6RbQ9
RqmYYk/2H+yMoRjrkjULGYpkQHZNE/TWENWBRp8jCOMWrrSrhKwySvW3mofY8qJP
Onap2oy95TYU/V1v8mJHl+Izu2TRtwLGy83DLl0Z59AisTdC85uLUkZejj1k+E02
GBSOV+RqCMlCJlfcZhffPJnNRa2T7S1m9NzLz4yWV/DUS3hyVdLsHedelyjCeO3I
5xBLRM5HR9Ofk9tc72G1/QJXjV1tOvxOOHBuvi3afw4B8HofxRmhKGdxGAxTcSMB
dNOE98LWEkVvcwiQJevlxgRwZN+LnV35b45wbChqSVkVQ4ADlNiKNhETTN6JAgTq
QGrZl8HM6ZxqUZaengCgqve7Z22Y1YA5USv+tNF372Rq2FykdT6UqIKqYOn1FNg7
PIVNkrCK1WTbMZQdAEVuzZLxtp60Y8ic/Jlg4KvGox8TnS7g5W37e1VbEwcBizfA
Fr8hDDkEGurpgm4LpYQO9bquKISPX6N87sR7EGMRvQYECSGjMq2n8a9o1pIgkexR
N9CLgbAAd9jc/pxSu6is9TiepxfMCmqqNKNlhQ3V/DimddL8UYM+cNpAId+GZd8n
LWXU6chHlcZ/AnMDpQHzRFxaGXgJjq4426eigdGkYhFmbTCSy4X73OcHc3o04iMn
YnPH32d/BIoXsPbXNDv/PpGCKKu3y0leoaJ0m/6rhIj0gk/SEHqBJz1A6G25hqRl
PAXavs5f/rTAyFtYHku1Ny6+nMnz827Lckt0yV4dXFuB+l+hHRONgaYFVVwSs6CS
GBLTflla+AY+7nIFKMdTV4NeH7JRD9IJirf9YpZ3fo0=
`protect END_PROTECTED
