`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFBIuYr8jt+KU1zoRJxhTKk0h9zCwsu6CfUcp/L5CIJ8GKu30cZJ1FFHBLgwVci4
q5cSN1eqMRDKXh8GhLUTuCpufOqSk9XmuRsGzcyUhv/sj1uLpB1Oad8mSP/kpQuk
hC9c4T7EnGVe9PMHcV7eiLR2bHlZixD8yH4q1wjjg4HvDXdgQ/f2fYR16C4eWdqj
AfQQUHh7zLNjkO1caImHnS3zajUDqn4ugER5lwTJW7EMZwGjy77NNKz/7UFpO6li
1QdXlBfhzmYbvFJDBrOi310RxfGSTH7O77/wecJ1/OIXxMJ/jJrIJjRiWfrTbq9p
V6cUxkONAuKDZ+ovSsor6pgjHMR49d5VaQ5rg2DVUfvTujtGnyehLNMEb0bzAcQ7
kAZcRASL2PyOR1i5C7ApnlB2rg7QqxqKdk6KLRDGIJNE6hcOCoRHmIEdsQ1SlqmO
/wN30sE+5QYuFbpVGVa/5dUK7r2vZnWZ8l/mX3K3tK+ORKL0z9zW6LFymUaXAedf
VOTNeWzjFwZhGkoPwCKkQ8/o08xuxtk6bhKmQmfqSWb+Ui02pSvprH2AjR4Ob1On
CrCeC3z49tgxW0fliB3ROG5xmUWukZhaahVWruCjB68=
`protect END_PROTECTED
