`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R/5lyMuRFzQXSxKwI3H/rFSUqZck2/blV0ictMQjxaDvrc3ICiH31jw+Q/rZkeDf
cVb2GE7U2gFzkqqrXo6vN8cDNEEAphbDfvdGMOx2Prf5+oE1IfkC04bzPShJaYY3
RzbAUw15yA2lDuonJ4F7K5YOGO53diahWHCpSig0+FRp7bTL8QnsUqpefeFww154
KkjqPh0Tj4XWEuaUUIDR1nc7CUEFNKCziJ0lDEvgjGc/3MPOO90fp4p11FaBtYjB
oAgp13mswzJfHEdQTRlhi8tKJY8/C5ORce076K5AvZ7CKh4lDgqhUotT4/O35OGk
XHPdE+RjCzn5u0UGiabi+i8a32YXriMrJ9j+ihntAzMCrPGl4Xvf3+wpWbfW1wk5
ufnR2q52IWNOIk52uFXiCb0wwcChsTR63eQdIwzZvs05r6hNn63e4fCbdn/NZsdX
Iziw0UBchWur6caDt3rG929KEwdWnSebRYhPta/0aGeydhFmWTLikfN+TlwX7YdY
2yi3SqSxde+71vOFmERMkxNJ5JFpYrnXx4ZP5nYqabIl2SOFwdwYpL2f1+WYCYB5
hGmdU0MVfHhMkLiwSj45ySL/Q5hzHV33y1ACqGWXVhZyOi+Q4HGZRAUN6xI4+lZk
57qWSc/foRKRzzLoXUqxhtYXFJv3IdGUBqJMCRp1JizdynKWdqRe7NnvmEGtgvE2
dWpt3d2wJSZRbdVz7i/zpWKZmWwZFHtgsrbRcMATKs20WqbA6fSHlfYqSuGfePHi
3ZMfvJr3efAmzv+0M8c4FTH3mPJ7V8pJU0tfdDc9QQQ9dln1bOCTpgQ1Odnnlk92
fcaYUz3XcsnVf1Xah9D1EgMPShTevNZ987ABf7FCAwZRFRUlJIg3JnqNUgHgWxC6
tUmr+Qnzmd+9dVOdXInqkYf1YotppItCoaAlfPmCErC1xX2GejeBHJMond/yt2NS
W13EcVVhXajX/ZMKpXR1uJ7oeEqAVVfmiawkj0SioULDHRtGe4BzZllqOX7X4Qs2
0MwsZHzASlynY6nDtxw5gs5QPITgPGl5iQbKMRi0c1mFrilSW28YxZ16A0JF1MhP
ng+hu5aieScTehtG4ocuoXvTHT7BZ6Xnlp29dRJ07PXROjMsybe82DnaHQ9A+frM
iqrjFUL2UDE3u0po0BfLgIpyIGoaY1Kh8qJW5+5SQVEOKh4zoQw4vWIvRdu8FfYG
gmKxgLue6JZHmzNMfJ5mxMEE87dgFSGlKJmzWTH7/wlWjgBGXm9yugrQcGwXgtuN
T+kF1Nvst8S1hd5iyRr8k8mD1Pa/RijSQWjeE8WJI4FC8jsadAbtTq0UCWhJpaqU
xIc08YApATzOOddWx/3RLuWEDeB6GUnnJP7kzzVudx0V+vv+RhXmHwU/bhLTM5Kr
TKUMWpjTfIgTMWRYsZoKgGbooq4h+Nd3nZSu/tEdBTqg6NMsOh/hLOhn0y67A/Mu
XnYG3tbvlAb0AgSEmKSO/kBoYWndexCyBWG+aTdTNc3K1bNgpl+Zs2Wx/SASjiwH
x7py9YWONsdTjNs+TBZfaErj8dGc8OjzPdtZA2px5WcKv7yQ8z5oFI5wsOFrzrwL
oMHNIaEJ6hi6sInhE5mNJWJ3hoOyQ4EpwIr59l2snAY97fk84v9G+pgVfvpAuQpP
+SRnabP1De8Hnej7Elr8XyRiargpBDYxqnlIhNEgewX1Prhx/RDFYO6YJLh51iVX
b6HF4YBsqwjgge8DnIql9kBfNONegpRFGF5vCJ2xdCmOMp3rr8T6/XcxNBVtRFZh
VpfjGej82bzQiuCo3vauUUSv/v/QDWzSn/Gquiakff/dXwebmzd5qm/wpYcHTcW/
OBt/gv03Hoy2XBZw0EIl++qJyV/CkR8kvwqGKieacEuZ/sY1rsMQm07K4/O0xR9W
/YBOG2IDN95vak3p/AeOF4mp1s+kCqv0TlHsjWeVmF3t1mxm+CW+acOeAn4sg7z6
99haBtiiNSg5RaMWc4WgCMQItyEdC5IThosELHHzBuJwupeNMJB5cgSHeC1u666h
7gQ6GFxLfCxuYmE9XwYK8Eu0Q+GDoTJru1EFy4S8SEDTtWJ/wXAIfQpzHPhWuBnC
W/EqnZN2D3uqR7Fh1IgcIOFU0nxKQ7gRMS9Yc02+svJu0sxZGjGlrHiIgCMVLb73
aTZP6FWf5PSJyaaUaqWXT+p7JS2Hmy6Y+5qLmNKXDHeadF+nj2otc6OkZcEbzDTk
UX2khpVpCkGwjkvi5wmsVEaKTWFo9npysHbOcdki0D7IdgEDH9BKCE6JHvYg1f19
PfxlZrzYHIlszUd43FhdNbM4UHgKSjRNEXFUVR17FSbK9iD0nTQSnu+d2AU1yaKF
Q8mnnMyuuQEfDuquxwnMV+bmQBxZj3wlaDawvjgA7rwqL4aFSkEy25mGbW0FEGGm
FvDKU/F9Z90QwQCADYMefwjzPTOG93NN8hOMtCuazFcjmxJUOeqAc+aFDFREc6c0
j50+8JgZxoXcXByLhhIHyUPCtqZXT4L7w+2EWmgGdaWG+KS/sMfqwJaePnGMZka3
OG/dbVLTSdlLmq5U2sQi6BmU7meImZlJs/uqc8pR5f5ko7vqtQAtBNpkdfBjRIfA
O2HqS7HkgDpajiWR9X2h+6fG5ICurxSXmyX4UkfX09H0tyKOoacMVJqr/FIcOxeA
TqsmLgMtU1JZsMT+T/rul8RlG/9oaE8LacuEBanG1i+tmOO8Y7iBqLypVeJbkx7i
/WNTk5/XBbsvzFu70tmigoH5CfXUCm3yrdyrTkYKmr0nqL3X+uJuQtXD40OtG61D
EV4vEdtOluIfl3xykXajyviNd59tzkyySbpuK+SDEuxRH6MxPypahUpN4QH9bYWx
Jkri05oktQqaHsmTqeVkyNO8trQnUaRoEF+TUsuRL1kBuhYoA3YxrlWLwM3l2WTJ
ISGbUo3XqHUDnEPsI8dfpD3JMlCczYN3BZKUw2WndN/3HGIlcxaRcOKjRuWLoM4/
0xuKadWQ85W/onHFJ+oR8w81CZLNsUAq2AW99ZS5uqFcEZrci3MVJFKKOuWzDMeK
W160a/9JLKISOvDVkpiIf4Ofc8Gwgt2o9dhM+gN/BfmBlS3i8KMGWlV3wOPouPth
iT7oUQEJdTt7aF664DGQ5Pjfh4saILvAPl7Hr4MuezWWa3J1jQBYU8inBSbQqDu6
IBVRevS54n7oXYuZ7a92K/A0+whwP3npicih0Ddb4HbyTlzpb3IFTYiakS3w9t48
XiJQMrRCvynF3N6XAzANsw==
`protect END_PROTECTED
