`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTBnzurOc4xNmxSMGNdEwPxIgPKNHRbXxvtpKtQDM+qLMGU40XVXLDQ+a749sb4Y
CCm2w3vAA+5fnNXQhAEcb0ZCAs64BbioBAaRrCnmaogPAqFMvmoZylpcGoss8CeS
RGNVd1E2+m3sh9VsBhqZzxZAS/HsbaJUb2tR70tgqzUC1eO9zv9WvRZDvWh85BU3
IqT1jXVYbo+Ld4EKMVsq2jf7rNvj3CRAAmgh2VFRluoSNaBdrYVcDLtrIAnl9Mjx
ntxrb139r2aHs4EHk3Ol/4ffPayngWw9ZLYMxsi7gcVeE29piklegoEAkRQu0QSf
B4I1tPSsy/J9dHxr/zLsgUMf7lcEVsd1L+FgIVP5sibiJ+CEUkaGKfqQ4sZjuR4a
BJUeHZwcygA0xgBQeSub4XsifK3fT8ipY7Ub7mSh/EP2XiPXZASxn9u+9HK7LOgN
aEurKUocS34+dJMovY+bUgXbPI4afGyeEueouK834mpvqbDggpKiNYNi5LlB/LM7
OWXP+y7Qbu/FgnJBEUj8ZR/6hFQWlFBbIlqwjHWX+mbgTtP8aNugfuY7SgYAQQ8C
F80ZY3WwX3uvgpvV3Sq769OsfSesSoZnSn1MYthJtmppksXaCVuQWczEUYDje8ok
ufY7TcL7eqmu8sHcaOD592+wYFoE4N4N5L5qwY7FO0wSAI26o/yhyd/UYI8WYKLC
QQrytOTYNd/pyA40kNpb0Ok4l982W0YG71Zu1OOJzYGUjz4wxcg7MiKLJ/6jVeJK
H6mMzPFUEz5ntrTHgUX3bI2uz6keFMUt2XrdqsAguLm84HFC3jwYCP8bH4kXkfvI
TWHDtvR/ZwegKDjuzTc0DWKK1O/z4YysyYCKA6ZcwwFRcAzXK1RliXnZbfa/+SIr
7XLs8gduWWe8YxKpAFFVSJVTUDQCIPYl8Fotl3krxWIOp6o2GjMzJ19aRsx9suHg
t81QVXC45yOSfYw3wLtTFE7xf9UlMjwYJyt5XKbYX1U7vqE6nag7c2Y3tWDXOi4+
Eh1PZB4N1gA2N2YkbxgkBRdQiC79O49ARMq1CTWwFh5AQLHJeJ4i/QTJTrZMMQE0
KtmB+T/yFVMgBvn9gQePY1Uck9CkUIhBVNHWwpB7hDGiXAfuDHdcRAaNJKeByxMP
R8ZGBVMK7Q8tzURcrCdqi8Dlk9Uk/ELfQKI1//JmoElS8xdLuMn5uQM3pMxiNfke
EVLxPO7ql4T0U6nHcV6GkYnKvyAZkWBnvshroj1MKdHIUqRfRJUpNHzN1kVW2Hup
rOYMF/88vskg9Z7eVhd0yA7xaZ+au2UrHvfzjVvpP94RgV2qqL3bR1BjEpyeCE/j
TYDrL8QDsMYF2PKSOc/S49CpUjFYukWVycLCeRsbH9eCAldKxz4v3THtwcagIKjG
pG9HjnpSK9y9+VrFMkIvddlGteBJHvYZ64uAlNDRyxx85cJloS5TmdLl0HE6+p2G
fDAtkWb8qwJttltTp4Fk39eiLw1Mt/f/9UsPZzNIeM+z9y0QbukaZ6HNI+bxa14n
joeuIBkxF2HKKmXJKauM4pcleejPUXDv6byOPhmGApadEPqB98A8izwSdeng9jKS
mw85mtIy4SdZQ6fD0qb3YUVUDGaV9ZkElQYeMdIFQsrRylOAL7OTMSKZe1T8f+pL
nsGHerBBkaT4eqLvTQVvziONNh7gZHTJfKkn0bNkRK1ZsazXf4BPjdUzwOEFxP5r
GX57ptdlJ1foZCIw/LC7EzfCWNODUkm+qfUvVieqttk/VcqEYTAK1XdA3G7Wo/9T
`protect END_PROTECTED
