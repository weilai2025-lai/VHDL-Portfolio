`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVQK/DNfA1sbx3wDN2jFEb2/t4fY+TDDmafn8PvPDRG4XZwthW/kSPAsWAmqCifH
KuGldv8YhMFZTFQ7ar05eE3T7A/hNOWj5p8H+/TbGQTRbYiAe3td9/VnV7NKhdhZ
0G9eKGiVaTvjwgVfYbdCaHLeo0i5459xCCtRuhsrhyPAl1c/uRWBv1+p63DYnxQK
wzPefhCS2CIV6c9oQyvTSZXKkV5cq4yjimLH/kZy7PY1zoQ8Ul5OpR84V9bp9xXf
NQ/VBECF3pKtVPDbu44evrmfzf3Fp5PDgfGCNocrhrODvV2mBGgKdwemrNKGYaBk
KUIoq9fL/MqOvuY66wMidwnUWtEPZubHsHKuB21/jsOtLPcB6YUl3yJMAPcdPHTc
KJLPhT5epqDOjMMwXY1J93X2YVA0pDm9SAY9HYzgyBCZLsf16Ealm4UI9IumjEaQ
FRD7P5yzF5BsJOE7agGgCUmHSOkG9rBZ5WIZcVUpVS0sUfc1sdT+uNx2XjNxmZqx
UWP/RN9WOxUAm+mUPR3g6dtUq9U20/uPIBsBre5CWfcLXnB6TgcEzZNp9Bn/Frri
NH+VRJuXE6RM4whEu368AHVIhIFJyGpCOEf6IaeVP46z91ufa6QGVBgi5uzC1Rhx
BKmeu0osWGzcbV9BWQUtKdjJH1EPmRtNxW8yzOHMlvmLN9hxD8NKxav544OVxAch
LHy8ad+647HuPL4kXF+WomTxObDsKagIhufUkmTxFx8bSmpUP1v1i3Q6ju8mherU
0rK6iY7RrE1Hz22pBPloj/bqplkIp/NdQa52qbt2RNgZhQfpBUOQRfBhX/CocMtx
liXu4tYMMkffSDtK1+aq7toNprWFC6Ij8McJlSte9lS5VQN/u3Okp/sUeRKr4Rkx
tn/JINcfNJUcryQdCjlE5kaWulQwbBKJx6q7SkZAvySoKrJhbgo9YiJolTGYDsfD
sk3g+WhOQ9s5mp+5Q8czyCjLbwhFQPxIbtC7r5VVIFyzzeF4BIjo0mxmvVPBo2AW
W60WnqOzI1VDw+SXSQejBU/JUdd032qn4P87z5GyIBtVoAadMQEl0/aB7Pz8Ta7f
eGwwBDFH4pYkBdYWaGsfsJHIangPEwtBUKf5rgjzyfERfUK33p2sVdoBqSOKewFG
WsAvR4B6jXrVkax5JDHTTWtOj+dSxAGhwx24wBTgymCPnH/q7NesgS1MPTiw9BFu
Yd3tK7aRumv9LRs+R6UJMaeBPcLRCyvPXKGjD2k9AHYZdntQhYmtsj53cjDMgtNn
m+x50oRzFB2+pcs9EJu9Tu+B0vEFm7reaoclmu9H43uV+QGUptPkCaACTNLtY5mQ
LrO1bVyzVmASLM9SoYWIGs6ndfDHntZrmbZdKs25mUEsHfPzTT4XbgxfsM/H+iw/
a7idUjeDz6lr0RoWMCbokesTtFdSJ7klmjoxR/PP3ZHHJVlPU3TWYX5fmi/omh/8
UcDHPnl2apuNXrvxmvFVXXNk0m/9J5USPSxXZzw1KodwMkoUlwt5uc61yWMGOnSV
CEuU8wiubFaRW5yeGgafIL7cIKSOnxeIzv804rLiA9W+ZLORzt7A/FrH6QR+urto
/Qdu+HyQ0SbSxuYynYa68Bckr8ZOBCa5pg+kmyZFA5ODb3zxk4caM3bTtD21UB5r
zm3eF2k9R4qGk04NVn6plu+VGMvKi/PejCSfdSVOhLxIFcX2NurLkEH9VKwQk1vD
Z1qAtmK0IqtFmaNNTnm6l3p3l3hRkp3+CLAnzZe8aJXp5w5FdCWqq185D1TKJveM
rR/s9LaS8LRGRCNO7K3PWuAsAgr969Ja8G7YxP/f36vvcEKfYgmrcHJD7JcAPDAO
CYJT/PKBwv6YdyWMWd9yfA==
`protect END_PROTECTED
