`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0w9YNmhAfw4MouT2gHzGwd0hErBh47xMvYxJMu7ej6o7yjYqFXdE9h9+T/Pb/7kE
MgTDHgcfpVTvBZeJl+rCiqPq9nvoscr8jjTpbVAQiJoCIUZx40apOBpiGSODZj2Q
f88h4PZ3OUmNuCgPJ+Bewl5G1M61taOKkGxYoDo7EYldw6y9bB2+5qH/7E4SdDQU
mcvc1D80VvtdlksF9+WGRGS7iWvUsx28x7JCSSGxKSJbUoLMWxh/FQVB/XaqXWzD
TfSri3XyObcj2TCmiTvvZD2o0z6pKDXd32IrsyNAvMuSAcSjNY0OSXXsdRJ4EbdP
nNOHRdPxoNXCqH9QkcV2Eo4bDE/h5UupQaXoo6xzsyfWsE0ZcdvnRvrhaYjSF3fQ
Ai2OUGZvVl6Vv0xcsLUabhnNMmxPno82dEzL2Am+rYAv1qRTAocKdg2t9jG0K1/9
aYSy8lrBqOkOffFcyUwsMjfeRLdz23Gi87l7EiXVoFWQSl6uLt6tuCqV5uSxos0p
xfe10wBwT6t4T3TN0+a+vZiFf7LJL40E0ijfqhYJZWS9p1I/G9rR+2IPMyS0Jm7g
kvm4/2ZbRPoX1I1Xld/1I71IOBCWDz9/bByvXZQ9V1lVFP4CsrRlSWRXE2tWsiZe
FLslexwj/vVYau3MEpcm8pVc+P+UdxJdwCoqP9v+GN1BtCPBK0JjcbIkbpmSURsQ
vgrv2ECi/UqEoZs5Lejl+sWnVI1OiDkKzPTx65ge1CmXkj4sk3AWjoCpobJwwKA0
L2g/V+1K2LUi4+58HMhfJb3cKJoMt9b8Gd4R9vZ3SNvxy7xR0tq8UA1Kti/JMPtW
gUD+WwHDBI2yQ0yjiofFxsXir0OCh0/v3k0aI4Sr5JiI1QsyKlI4cByouIdg7iWp
jZytXpS3pvwio38VuahcttN1uGmT1bCd6Vr9zXt6jlb50rfAm6I4X/tM2qmBNDHP
4rFCIC86mcQbsPSE5yNfR4D0luLfX0m2noY4zlbh6frCDu1CTU0kQ1/4v7uabwoc
bvldBuTEhvWwuaWY9ci0eiA4qNBAlgsxzpZMEcnY5HKIXHCyI2xG7Ecd9cL56pps
Bz1YcWBINGp4VnAU07SxNigTuMTGObR6qC+cN+5ADCCTwaiM38n2fWTDJWnaDpn/
BL9bjMpfIIU0UPObMSrF5XaBwZVRSHrgFdLeb0EoFGLi5BKgl4iX1n1tAcePUgwW
YLyogCeCSTn2fEoM1I00VjsVOEowzK33n1lbVHDPxZaua1Ra2LQ1AQAjcjeykZQQ
1yuVVaJvzUTmJaqZwnYzz766EM+hfkuQhq7Vfswfv/S2y6o6aG9Rt88KzgBa3+Zz
pCU1OjRhejPmbIjX60tvYG/F4GIlzvRAf9mMojCfiwNs+wZRd9R04njYffU9ea75
NNNvXwh2DL9HpwNGVq5AAo9yCg5Ko28LG1/8VseeaUug22sShHzISBkb4swQaFBb
WGklNkVpxdevq1LQVoqh3DrNNR6JJGFgkJyoPN6mjK++hwWoXX+LrMxDyfsF28tG
Xq2nVz+1CJ5lx5+lqr70XoD91YoJbLBPu7VPIAC8o5c9YmtTOhreUAzSY7r5r2cP
90xfC4W4D+Wq6z4l/kn7RlsdeHSxTwKTLxiC6P2otKI2oF/PX7I7ye5ZTi/0N1Qp
Xll2DIxhOHZUnVlzvPWPZAtHsIPxFcJia2cQ7i7Pfo4jhVvw40aWY5P6fJcHwZPR
ji02yoGzok8DYKNVneTsxEVYtA3GsJ6PXXEBeC9y2DqFONOkWx4H0C3AArgAOXLR
kLNnanVSk6PT8hMK/xAX3cAiMEoarFpKIHL5R8FqPXvtmq9Ons1BZI51JyAjth4S
L3aAZUp/iNGS4lnmGjvzcy+Y2yVZTfJmgBTJcJM0w+DawhZLpKC+oVHb5i68PQh/
LRHWrkBCK7gTkvz/8k5mpJjeu7PGRUe+6HX4W/teOwiV0Sj3xQFpufM7D75rqUBh
tkCUHsuoi5UduU92QZNu7zqBwE8S/nNrWyFPEKVUKXtAC/dFXgApzvTmDNpNTBCo
FvpaNfd7Mir+gRLxPKXMGUbwHT4Zev9AYERFbAQBpfCtLPDNb2MNmrdHtveGHfZ4
TJ4LlbUcy7ZS8Fr/UfK5WaHApw+TmYCBNp4bEcDPw9uyWrHbvci7k0TG9j/aSn9o
Hy2Wv5VwfhT5eq0xxnHm2Kiqlvfg8tUq+5kAAZyj4JIhpA8ORL8F+n97iSicgoMM
ZIBpTIfpnk0mM0LlKraQYHk4+lL9YsNrWXyCUGTgJrDVO3pniha2N4FxAL1cWM6o
ZnrWqbmLpedvfrfsk6cnrItF42c5W/R7Si5yxAW9MnzTmsZ0jOMRJaXIJUQM4kjQ
0155l4hWlUdduAf8uk/1pA90kqH4uklCSHQiK/soUlVptfiynXJ1cjJ3yB6KLVYV
hYz2TZl0qlqpcFtmnOAtQOA58YB/zPvBZ5HTmYg8dyDaClIIoyBktsOLd/cX34ru
C1O7vVX3dz9MGXyTpgV/QZuLdZUMRI/5OEyLaFeEohTeCeUdX3KFo6ieCwP1o7Ss
yaJRXY/6uP1X48doSggk9NStNgNrBm56GXlcZAszBbpGGMmymkvlB3Nd055KzK8P
aj+4esLdTsaortvfcqMfjpbokNm9T4Dt2B630Wf9cfh8fpsNt1R5cVbKcuGIVO9x
9O8IXnbWQ4FV3qoBAxyvCosSS5J8jTtblAM4Aqxxd+FaJgmRQ1BaOIrK2px0/dM1
Z+hivFf9sXTunoWoweTj8KOKKx1ok3Kt+kjIu4t4NcLX2O1X536mHmBZC9hrsfxJ
H87lw+pOCp2kvJabPzafA9p2RJuMCwvmcSgOxXBIWdDXM/udPojwYaQqQ+XM3Y0v
2sFmCXwriPK/5MlDBCkg1dsm+ok7udD3DIX+J2bKj2WSj1ErnzNdfaWZprqva0Xo
jdrvrIOY2JMvg+Lc6TCOTTbePDqaItdErVnPycIBwIFUFLYAzVejiMUlpq/VEIYG
/xp/0JL2iTFwfLJH3NOw+XYfNGpywB1qegYACVlihxuzZlDUsZxTSHERRtTaiRk2
CB5VgjcK+eZ0Rj7i1PMzcUkwGhjwKHMq7LEuiOra0D1BCeq9uMbTHnLfl9LFlzop
jmClKWvqfUtVGZ3rn1bSFHiNyOBxxTvJ4XyZKHACY8CdS2+xcanRBRh4EjvKQwoE
XzM2y6DXC/wHeTXmD+qqW7v9++2G+TOpn2B6mo4C8nQ4tQlrBroWUtklHdR3l/G3
BW3E/hNTW4/nPoRJy76OcllDanrCaHuyIJwg4ZtQhNzwd21MqP82u9ovYrpMvHPw
0c24TkL8dosoTeRgwxHqHjdtPqGP9hwFgsEeIKgVl4Efab3QSwg34mmkqo42JQYb
KWtEQUmFSdlo/yS0RgLZUFyj1X41deLnNkO+tDgemZ7bSI0PCFUCvFyuLvUgKPFV
0sJTf1AMTanCUoScXKaaSB7nOZHdGj+ibjUZVvCz/eDoHwCvZIXwt5Wb6u+rjmO/
vdoQf9DpSMyeLcsgFY34Sh9oeLlw+Cl7GUUxyxPjlmfQqazL2kd1fBznfDN2mlpA
0wA39O2yWxDb+hbK5FAsyrKhekHgPIgJvQZjbvcH/CtersR5Jcv9fmzN2QOrwGZl
GK51jAw7VXAJnAwlJo3m8Zl8+LtY1f6v2+osCHxjdw4J71S9C0wXQmelSttbHT0u
anpVBiUp0nnHhJ7rclsWhjf8WZujHbeQhAPIMrrtXbaOIPvfmofxuj5dTHeBk4zr
it0NZRm4FYrcIgdwC+C8N80UK8A+6/oRLSc4dluhPr9Pu/9aZobXX07vrC9/4a7t
lYDwKZ7qxDdqWWlzheKMwkbQ4yvnNr+SHq4UfyAbbvRdj1hYHwUGN5argC4YoCVV
YwR15nePJFLr9+T8vSQt4BKoBqJSf1Hk4r3HiSRmo7dotivC8u7KZfZ1bP71jCBx
vteqZvXrIzB/LC1Ss0OeEpSKM7G4JAI7ptoaiAF4i5wLrfTeHzrutzaLp//Jy8Qe
8Z63f6YR72o7I+iCgitvw+zScuvHDfeZfqB2LJdohKyL8vGJkl4I6OaO5XTK9bMe
IdvIInZvSXvzseKZeCpLq6cC6Aotex7VPLklzqAD5eUJkvRQC3Ha2EWWUBLiONwO
QYbIe7l+aj5kp+OFD8ykHg5hSoK8ALLQN2TjjuIX2zwRixd67sEkkUzQ/B0fLxFU
FxebFmqYWQ4oTn+89pWr9Kc0ro2IgyK5cwjfHYBEoWq8RAUknkUPCq+V8UiPblG6
DxY5VnWaOlM+jQZ3I70CS0mwcB0pb9a9GqWV/j3/R8vtos72NHVDgI3wWTxtoHDD
D3m4VOdsAe2WIyDnHKZGCHDDHqWBVU/io9Gn0f45XIKEtMEUzv6oD5pKTkNoDYlM
jSK/glafluNwNpInL5QGd3tEnj03bEckJGzOSlKXPN3TerggXNOYNyoaaUpk2bqP
OvY1WJZMDY+2v3vtG0B7GlqqxMoCHzv4+SWnZYqJn66G64og35JJVI0kFcOplOnt
GfIaYRoiwE5hg3iQfkNA7ut3TJoq2rrL2qLLtRn2o5SL/papLYR66RGXNW75c60l
VRkrcjh45LnAf33PQuBK7KIoS6lmHz3yyaVLns+MU82xVq0hTkxrt95SZ5fohFCQ
pfMT9YzEgUPSYE1G2djsAAyI6YcX9bOn6qrQf9aT7tk6E1UeJTay/QJsg7hALco3
+Y3N4LSQ7j+hpVwaNRgfJkn9TB6jMs648G3E9JwHG6aej2wlHKRWRY8Lhob5Vkvi
7qIbXeB4HhFgHu2wJ1OeTCytASXAHApRwFoT0kDr/Ym9LMCGVT8uuLJP4KFkVH8z
QHeBEwYC0rIE63IUWlM+3ilQSDAeVUDXWhM7lesNSwax6CIXDxtSCnOS+/i3uQXK
/tlDcW2f42EMBfzyLmDJ/UGAfcbymBiZ0UU8nipcVgtiOlto6sjqPE5gtAaxXcg6
dpq2sXRtlYEXy2eJX42QdwUv5PyNX9Wh42kNLSOHLXWT2aV7eKy+SRMTVtdrvhJw
5/mp/o3hmp5QsmW6JcJSTqWoaltpL2eDigM6fAkgEnAt6GCk4+RwWwh+zm4I1t3M
vc9RAB78ui25U6Iy0PIsTHc++H08xBWALGF0CrKk80mC9aQockiveyiTi5GNDK0o
uSeT16GBDOA4PHk49mza6frSWvUDjuiYHRVGE9jempru3YEx1089KkEA8mrG8GIs
9bYZo00kzxk61Ytk+H2xNAOVCCq5BDZAmc7Ew8PUSQ9fk/UiH4fKBsslMP1DKhUt
hzGAf2HWB1pejaO17LpHLQ3rNflVKd6L4llhmCWMQsK6wcOciUJElNZfYTi1EfWv
PRqAql6lrEtI5I6sywQPbt2vmNbb/zAI3iKPBJeHjP3eS+ga9TvvOpUY/apCI20r
StEqITcjEOULu6+0L83F2HtX+wqgqKiAvuDBxVjSFDWu0wHmYx9lSg3SA1R5oKyu
Ck0WEdxiXLn1LjwX2tIZmq5RWWWNqKv2CfM7SdtB1Z6UI1UljFPlRtvIxyyFt2kx
xBjP1ocuwa94ZqVftVnmExQScrCGA0HclHO0iZx/sd5PAMAFrcNxglNFOMuOnOuV
oVPcD9p+hnvkN96B4FCsmyGjS0E7SpbsIKCYuGL24rP0AL1VSt1O6kEMxUQF1SRQ
+ja57j5O7X1miBWZvoCTdIClhfUWyyKgbeSMLoTB/I4hCw9FoQMo3ahQQMUyqXYE
LsoWNvld6RCQsQkHAEg7rweruBcviKjHwLxyjIeQBjVWDp2uGHgsp9VLdgPUL99I
7s/7rLpf4ttB/AzzWNPTalNgAu2Z5hRMeWpUxMHh3q8CgluFmLwTURF7bK7oEPCl
y7Le8b51dm/ProwTOBZbBIZn9TaEjwDZLMl/NCibeIAhaVZN1cdZebatLDDhwylJ
BkaNnL67NeIMDC2w2u3r/Ru/AAasO0H4WWQkXoKBJWWgNs0+OuSgUN44A/R6LPUN
Wgy0OB3VgNOi45i+vaCBXhmRREsxSxGA8bDFSu7TeTG7zc58UwU83fiFwincwfPt
fNTXDsEAoRBvWW/FRQS2k4KkzqSVuNsWGKr77/Zo8Qasw/ZklPmvBkjR/xS2MaMN
yFy78jZjgc79hLFM7PN1RM69p76jm0Gsr/+j7PNo9Cd3ztvfxj5OYWfmx1kKqvKH
+rFbOoZfICX/Uxh94myrsTVSi4ByVoio58iGLkF91mhZEgafYV4/+2z2uws0QNus
AWy8fx1+mSPJpPMIRDb78N1Qe8qv4qSdCG1DXdjiMl2bBOd46+yRobZ732mDE319
GmXtPGIcActa31MGR1BvxwTASkUvYcQCz4Wbv4bw53TFYdwMGRLUgVXEagg83Z+D
8gXOINmNS9okBWq917H5jFbQOyWRl1UEWXCrBZwjpEReFUzOSBmAlWaBKstAyw2Z
EE5IOJ8Fjl/Pkh19VRGEHBd4ocGw+AKCm+8qoa/OF6eRzGncD0y0cf3LFdlfHCtI
PXsk12JZgrPeKzaHZaodyn733EUiAN5+3vgJT6TYPIY8i2ou+VnCISVe1Zp+bvCP
hUUVSv9drzhpebJ9uSVOxVkIYri1eOXIoLEnFLAFTLtSl7atk7lDNT2b4XMVtesH
eokp2dp7YqGIk25gfTWlomEAaHl49buKQ45KwXa5ntrN24bkmvjH91wZRvpFPAw7
eD6QAbOmZtg2LZ0i9NsnOm09DCJfz3/b5/Vos9obUPKruPpP0Du9e/ps2nCEb/l9
fHK3iT/8hIivsUOc9FO5gqVDegI6rb+plSHPS7u+XPuGaqxDSbx/FUhAa02EVEqO
ohgTM2ateRgbzM3s4imdv+b65g66TSanhXnhV8WPAG+9Lc1z+EGQfmQdhVkRbwar
i8abpUCf5t6lNz8w0B8T4CIhjQoC4W1rVXGOqNO8Or4KQ3PNj3RZ8ZlmIx2jLWij
S/1Dvaw7a3cd2uHgTHYJXS0EFxAV/U72SF8gHT/u3gjvo8KfaedL8sabKP/zsaDn
4TbLSm+3FWuf1n9VAnvvjSlxqCVh6COQc/YR7pOnPGOCAzMBct2Y79muUww8kdle
DBwDNAdkIo7lPEc/Ws71KNN4WB4YYDJeSr4qPpArn7quCdpD+OL5PB9zruJC3I6i
Vcu8/XPJB8dnymQcae2YhCiZjugWb8Jrp0DaNWaCHNt0OQVpQTUQzU3qAyVW+Qxp
r46OvsQBwmP7hG9lA6gCs7ttnPCeRpD9BlOeNmfFO1K/kkhw8XbU2O1b3UBrYTZS
kwDMEFoRtJWCR/yZKd4beQIsFQWI/byeyjkX4fz2U5IYr/gWZLMAaSssc0Itdoxz
fvqjPdtG76wrY1ean6gDQBYDkGVTZ8yE6gKP5qziEQ+fUOEt6IKMYpnZu8mXqy3w
+LJIpV1VCooirUEWwGgFsf21A8yz4xQmuHSf8oj95FpDZiRBpuI2ljpd593eiCR7
zFF2iwIRqPylybrkulghIapFOKkRxHNotK80q68xRl0K3Zse7FWoNPnVlelvbicW
AVDPkWAiIoucVXz77zo1uxvuK49Yoo7HZ4SHjFYmcAIe6nSjZ2Siup6oh6oXX6v7
G+swqB1VuKhgE6gQpy73Eh1wjw7GV3wINrdBDccWUkGbbZyGglWjgZ9wG7+wnuTR
/KP/AfX6ndkE0YPj8W+DtErRGfUjsoY8QLIxZR8rNoLSVG3JurXlT0GeKG6NyLpX
cWySI9xlPw0eqPZ2u+dZ+XQbnFrPWYosIHA1TIzxUW9ePtZdm/LflGNqHiU/yJDl
HbHBIpMvOiRHcecD8xF5FfxilyzdKZruwvXRghh8hwMoaYXRIbtQhziMMDzepAUp
kTpz9RaU5nynUnL/RqgwlSK4fTILDzqL++O7ZxYg03sBiv76peVfPt+M/19bR85P
wPyB9fxXywhihgdcn1uUHgBuetOIby3zwfs4eqtCGFYKjp0tH5GW1r4NUNJSyUrm
NESr/jCO4GcdHmHp072fkjNHrSxmkbSc9nAcOyBn64/s8gsFa1ldy7ynX8W3boUr
LI5W/C1OUsYX5lMgvwdia007LmOpl8elYX2zy+MWvwiXbDoXceblDQigcBTkQ7Bd
VUsj7staUUrUSxZV871ypxGLgzJhVsVg/EiAfyPboXleoTXMfLKVAVrMPcPwiHA0
8DeT9D4BCEzGmWQE8FgFtZi3e3EXsHgliGHQalQiIGpFd5tERoZuO7ZwJuFk09fF
ZdLQT7PMlCucmyKmmFBch4Uvgoqxd3oe1kUTsPlS0YYQUSX8sjxNOJ1mbY6vmw2d
GTqNZrzDWGa+DuOm9Vca0NWAIz+oE6cH/IU8VzWSGzUC5HzL5C5dsWPYp5A4cGrO
4CiKNcOxAkYPTZaMpaVbLLC/FZBTWoJIg423VdGSu91sJydX35oZh8xtLQ//CFFE
fxNiq/EKN1Gmap3gzv80Fk61fUNAS/RM3ObE8WOiaR15ftHYbPYIDuczgMm8Bbmz
JUCjdL4YcZXaVn1X8C/PhkS/jDhcoHwnbrQJdgQ3HG7c1JvehKjNiw4zdxBPotUL
FeUbHwVGvd1Z6u0qsNIV37b2yiz4KlUguoCkl4NddI4qXnjJro+wSrGDLtKgY8cc
LZRXDYil8O7reLE33zhE0wnWGh7si2Fjvvt7Qly083XD4H899pO/e0HG2Wmzx3/R
2DlHiLaTaw+at2X0X4QzNogKdhp6Q3rLnbco2LU/8Ap6YNbSsPdzI84VddikNjbE
/P3zq88GGu37H4pc7DCpUWUeU7lbwlhbbqg7xLfhLjq7vAsUEEnj/bTAq7ZXQFTT
u1KgY7dXbnOn5/iIDYevKY1UZN4apC5C8oFoP1vnKFSYPE5BfR1ZrSXtTuou2Rhn
vucpbzKNEX86cwdEb2pOf7R/H3rPTUU9jn5u5bQ8xy2iWJd5r47Sg6Er7+8POSaA
26jiEdBtHl7mFFedrVjljOz98wicsm5Xn76fDBQutSKbbCowlC8RH539MlGfhA8M
6cmUH/eewwFYub3RvUn4UTiMFSLvy82BbT5TOJFI+A+fHuNGjE7GSWs6nokIwWSf
vsshveryhknteP1dblfAnZfDbfZIyoD5+DzyAmDTRLPNQMC72Dr6JqeNW0dgaqAT
wDpdbLvoeOUxNq5HeekVsZ5XF5Elh9O8kIc8pKbQgGbXWtMk8n1RqBUF0H5E3Zdy
Or5P9aHhEZE6q7hD8dvf1no5eP0JvTdOdR/k4dry8vdy4mHLxnREPuwTT0xUtx8e
oh34qJFfjhzU8x5wknxAyJFFIfRFhlVk3vKxnjlylNZx7te3Q5gHGIq+oO6iVQSO
IluLY7xNFvRhbelTAILMJt7+l/pHScWd5Rphll5X883DZyIeqwKTA75Z/TSAbnfX
5VECO42QqNXsNeCOEx3GTXA0HUvWElmcOvKHQxyuZBNPsIaJrGAfFcwu2OhV/TiF
EISEkle9RD6ztXbvGvcDwO3SKBzROG4TE8adpZEdLrqcGGOsJAhT/gTVxIWF7NGQ
TuHzfC9Fzqapx0A+2U4N3Zc5GqFkJ6Z1/dBmQBjGD5WAQfeNkvf8wVKDNFs2apcg
0OJvxpX1o0AXmWVAj9IOAEGNJuFk99TGWowyRtxJJXUJ4ba3kWr3IuDopwFiI2OX
wziL1oTl5jtEWj8Gk8KxtE6s1V0EQGQFXps2SLCi7kK520KQRwVS4UQGeAfwc/XE
uPVNsTUPA1s3zCpXzsnj53PYmw/m7hQDJHyDwhobYY2qCVKrLJyzfrhLCiEmsG1e
mI2fbfkLclY0r090LeqpKyf9Y1ZlJaDr5q0DnZ81aFWstX4nMDxT4XCdazwgKHC8
Q0Qfvs33QeuIWmYS9xhn7bamH44Mojfya90Py/mLxx+K+5D+CNBBBJEzPgZG1LSg
CL2yFj7YHPloFTjmBWCtkyL/UiNUCqZPZH21GNrRNZGFOk2HvakFA5j3IjU40faI
RZN3CvKlxOonRWu/XZ/U0l8FZFZ+5pHDV9anp8m/fBPbb+ybuWSNgZnBhJt79joE
r2Y4ifvD9WzpvySvwAhaVPi6ad8FsytiAX92BdhiZ1aEwl1aBxQdcDoL1njDuOJ9
MyZG91lC0+7IiJlENkpZRt3cKwbqh5LBA48gNJ2fWaAc6UYcjIrSnnjA1gG9QppV
RR4YKDCYRa2tMCJGP9OxmxtikhMvnJj7lgF7EgFhdS+sKrFDPe4cKsobFHbB+1fG
dR1wFOyzxEr1gxUeXRriUhxFTHGU22+2eoKpe3ZAzdrMdS33T9PGawW39P0TzFX6
R9/Sp0/8fkbI0zsleDEv8WRgd+KtckoM2MQFrpjo77XBWpqH7VVMk6p66U377tj8
AfI2VoDlhlRJC0ogs8lb80kKixglvpyrzik0w6XD1SAT2mU0FDOeHsMVR93wJu1L
Flxnrypiy7OiAQdo3Xn5jrh/0oW58QTAQSymSP1b39dn149mXb0patR16jDnf7NM
xqm739leg8R5ejqJwwP+6aBE5XgzaM2B3VnT/jT+1OVQVFirLiFZk8Qy+/Kodv6a
L2H4/a9HjfCmTCfjnF5fOoE0QRevEAKBc6W+Z0dWiVC2OhQ8YdwEqlsiaO90PBmk
xtoi4J2bDvLMzYMoCOaFARTV/s5dSOU6OqDsLe8tePpeKnVI64HcTLl8l3WuYqvV
JUXk40NQ0Dogdpssbwo/JxhcwGhStoUqVEr15dbNVHl//eyfodrLtwYCY2KMn69Y
UbyKFS14WjuOPTPQwCVfzjJSN6m+cHydLOk77PJy/DVs7orMNYTvxnzU9qkkVSdN
e4h0OOD73hHxgBkQV6XIF5CaceLlTtEm9/yar5PEDjFZV2wa7gBgDqo2CNSzYO/0
DJPNevYquGdq7wDrK/7piEtChr2hDItN/tCL/6fHJ+TKHU+nTcmeJ78bXSDSeQA1
8r04Mx7sZDRzIyRJeBvjmKqmHp148FRkSzdg5Wv2E/WB0nMECVKnFE1rIZJeawxZ
YAppZxTp6OUAq1Gi0bnoFlYu3DzZg1uCvaEfgLyNp4fs4sHeLslj20sA8D84bMlg
hLxMY6NNL5COASGIGdCtAlrT3urlQSq2d1W4/1ohb3+NJwrGIdVO7H0GHK0htNpY
HiiDrZ3o51yHcLz3MtEoE+NmNwavFxB5qwy3y7b8hBodH/fAh47unrQO9uJD1rN+
a1wUq/RGHawf8YOGm8TtCQVMNHDHip1TbymQsqn9hRIoGiuBaEjqVffhhSzktX8k
1b6zWgY9Yfs3DVYGb0YLi4taAVzuaLfSATDdCgFazYocEk6keQ4br8V+IJP9cp98
V/HmYZtgOkU5s+pVTpRqRm3w+HyFUIUAD/BB7OMpp4j9Bh7y+Cuw3mNrWUBltOdv
MX5QSxfG7SqCFDhY0vVe3+FAegkhT00vbnj2xTfk6jk7i6jzIMk/Nw2D6goZyeBk
ugjCyvNb4WzvAu9j9GWG/F5/3smAYdeBjaSqmvBJAXlGSz6XqUtLoSTF3Maj/0Eo
hsi7sFUxGS4aWtxDDTUpykZEeTzAjaD/MqpBw3pj1808GuH59s604VEGprDH+fO0
uM33XK5nHu3QOTq8+r9Xh1tqOCUqhcxiZymYIsVrdXb0Yb96VE1VnhY+MYbhIXO0
g4AreKk7lXYqjC92QH3rH2rxFjtYH5PcwcmjxWcb2n1Cmi+B1h4zMGPyyWCFSws8
QSjz3GlLQ0k9HFttOxbho8CRDn9J5767TZAh4kCRogQBGxw5QU08uRHuT9K9/tZU
XYG7nyo2osQMYmUXOecQ49COlQNoQg1x6BaieIpBm6RHf8Xby0YdHRLjFtXU6cNq
9qjd8WpTyTs8KCeF+tkVRO03k9shZgSNAK9NNk4oXOIKjEVkkH7Jzs2XEN/iDeMR
W+VR/N8is4M51LbHLm933/ozjm2hQmNYu8cHwz5qPImPcEX99+lHxloy8SjLuViV
C2wrJL3E2D/nQzDxh2vAnuaE8hrVntEdv9yIlKiNu0iK3ojFJP6d9P5bAnz7KbSb
Zb3fAX40KuIzNxRoXHF2SJS6En8OYUD6TaQkK4TMujcw20XofwmCY5a94Yl8kydf
ccqSdn+UR1Lf06nyc2b6nbROMUaXAOv3HRpNBeOL5E3CAtrcfPlro1iHty/07oB0
nZSkrXumzWCbFs/nohgOWifQYNYIdX2RCZQlKOo9b2Aa/noIQWxPO0xvKgtW0xsS
dap1brSHNSUQPZ4IB41VH+wE5/Dj4b5apz+Bk199tslAMAk8ueKqO3y4N4gux9Or
V7FVvodqsAOlc9t/ypCKLL55XJ/zWP2SOwiQveyqs2JO4NZ9bBp3YKx7Qodsf0S8
wp4IzX63cWcAuCNoFTj/0M5AUgAeqAXBqCF6z+Tni6ADFx+BgU9MGe+4Ix+XRFsJ
vEENA3e7ecM9S1ulOTDSZI2hACBxCJyJ4SArIENP0vTDOPdCemiLoraGxyHZrVnS
8bmuVH0xFVfgXL/cnk1YjTvp5KOwRpfK83aE7UiZ9gPCuBgVRUskeZkq4fhA6TqF
3DWo36ipyTQHNfnaLff90VjVNh+5gETl648T7qZmDy20Fz9+idXow4+NGeO46+5H
g4P8ukhli+rQSE7z31Qh6rDBwnpo9jyOUeEVUYxWOUIeS9Fyj1FbHOPr+CfWaMUn
x32UvR8f8+5UTBwojS0WvdHMQUTBnq/TueKfcogCR5y3prSZp+wnu72iK/PGXbfB
bAybiqAImcFqRED2WwgXndtiCKzf1hkIlwRbDiZ5Qd8eIrPCSfCZspaT2oKzMjmw
9zefr1SgLgmvKXstl7z/oxxfgL3rmPaeI/P7I8TP7eGlfylDGSk7FaJj+CvIV4b5
fiiwtwY6OgT2cnpV/AjiKhQ++qkP6RPFZi7zhbWcCJH8gOCldhQj0M53jfQC2Ddm
f9HQfD5xEQBELuAqR9jbJevLU1l66g1Z5SyzyaOJnNftazPp7d+llPV2LVqNx1lE
DifEvvEHt07PfQzIqvtztNolX53+cJ4ga/H6Vmx/FmZxN4jsER82pxiL85z6nxgC
u22aMRTev7ckORye92pBcE0wWCgnNpsmc/yYctMZ67kKLV3oc0BiY3OFT3BY3Y3B
26feius5SiDJ4TGQhmJNnaes45mX+r79JhWcqLdmopG3FUeK416E0NugAO9LsNCl
wdhMeV3Uq+QBwSv+nu64XmjwoZ69ikTSXP/T6IFZ0d52USBt1ufsGl575mbHYCZN
Scl0kbKUnpulAHw0iFnMQ9ROO/UJ1MC27czEy0K+umdQMyR3gqLxxX1xoy/BwJ/2
tNEfjyMImnmihEvEwpcngVVZVb9YUhBPm6RiADFanKn3YOzv06eqdfGy7OHJiq6H
kwFxMTpu2e8YBCVFfhrX9d12wWdmevlZa9SUPkeqDet6O5HzkGl/CG+HPEg4DsfT
kZ/8yLB8d7LzdQ4r9KoWvXJ+CtSYpwDCodxCl7MOPEFxbVRFIq1wSK0CKZpDMxuR
2S8BLjW/zG3AjwQuS8Pntize9nmzaaXrwlJcmQZOXOsqvfuffPY/v0d2e2UmOuNu
+AanF5bIqepamoH4LHWTHt9/Fy2dbbE4Jy6eH2wNP5Ni+yiuXDUpLiXN8eIQxJzn
znyjMsZ9T313VIxSQ3xYHyp8Ll+x73BAK1n9ZYlX2GVMogqwN7NQUxqPaz7BNjiB
Kgn+Of4DpVUj1yrtq+gPv7Rpu8CLMMzNaINXQ6GIXl+30MhMRBS3NtcQapQfD5qZ
wgmzzUl+04wNOCKWzEtYyurAwbyjCjQf6RXCOOb00WRymW6G5T8Jq0GKIpebxlK/
QyTrhYKi5Q80ulqcC/t2+KUQtPlxGV/9RaBbDIBRlEjTTY7+WEwQhl6OOn5P91nn
oBkzjCITr/ZvHBxE8/llDpmw/3E0STzSMYQOO4iGewkkTmGM0BrPFSBjDeOIRLxo
o2K2T2C8IyCZl3EPvvThS9zfjPjEhuRSXo9UPCg4hh0rJjN1fPvKpHjH1AiCYdjK
zYeu+6S3WFSbGyNK8nDDXaxJgEx5FGS8wZapHk07AfO6nupTC5ov3VB1SWU+swUR
b0+mPngl1n7Mrq5THJAuskX4TzvPvOSw2C3vxxytiHkW/ubaCCS1ABMrgO0YD5lV
G8Ut+wr1rrikz6iy91tjFq6skD70WYgS7iyVshvtc3vmfdoU+dEk4n7IGqbYh6hx
JBTIKRoraOxtxfiknzBoxJHwWZsdBvhmncLfYMTq53N6AsrEKQyBQFnd3TTFLXU8
VPGoH5J34a7GVBlA2QOocWLW1EUkVWmm1brzOvsKpqZVrNWjGHhRDjo11LbqwlNq
yI4kRqGpDs+s6K2VyxLg+AOiNE6LQSbycW38sOMkt8Cwk1yjF8qQjwLgs7r5zjg5
/LK90i2POzB5+I+kMNiK8Lc5p439WQhuejNHKaq66angS3K7+jMN4T4NH6/DhuZu
xwb27DcAblwZ0ZhFIQAiKTgBHe4AzjIW0QnMg/0mHhx0N1PFtgr07ElmY5rlm6Tl
UFlxiiGQz8QTXQfPRFo+GibZR2168l3inMp57QsRN0Yw9exr7zcg2yqRQsZvCNtu
AlJDkOsYyUj1UI7lh9/1b7iQWQt+vlHooCFITeYZCOO3V9uSUpk69oqTWT8JsJXr
s5CKt7JhSKapdp+j/MitsmE8m9wZWbi1bclVNmvbWP41ElmU/iGYCla2mwNTVbW2
HUz7CCG17fQfKqocGNbB3bKI0QSdszD3ZzgvB3aubyVb5wZiZpsAAQDKdvJO9plf
KA1qC1MKjqG6q3n8qf+TmbJ+LXOfkRI0jQjdQYzrKM0uhKDsGHVtPtFcf0F6gFXs
vDOo7hkNEGWdBD8voCrKG6XPdD+42hrRFHQRrjsmlRlkDYLesmNnHeNnsRqFmDo8
yfBZueKGVcyHb2x4TPIlymXlLaj4VzOOcJga5npKz0kOf9R4zHJxw13/3PIwCgfc
keKxgLfU8hVVO3ws66aUkYIgxM0Wci78kAh/VnVEgahi/zkFn5oPo0GuB7aHxpvP
Z+kMQvLq6nIjIfa20NBIPDzc9SmWXjA5R3s9of/MxYv+9fTK2nvr5AXrChb8P4dP
sIiHffMfErvLkpjaIS7JY3QepGyKjslO0PZ+FRQpMs/r4fGXfBj+AFGChzhHVlTB
yfKv3zU5SPtgDKL74K3TXAnGQoTS4Ua/VEEl1C1FTiNaCVUu3j9nrgs3TMnlFhby
CKKWcW/iLPZqghu4k/p0TM91WeTXO7LpaE3KpGqLtgcFihSAK2k7EGuS0S4lIfBf
uCOlnXC4YWNYSpi20ukec3hPGs/27OUkbo/1iZQetnc0nIl49yiEtnwO7TSotrEJ
q5Ky64Jn9LeL0fFqq2jT/i9gm9TZCl76owQ1yzCUIH0ey5SiIHj7JR5ruGb0OpBi
WdZnyrrb7X4aX+ni9ag7RAiuonGnJT/JzOp860z+5jqmZqIBYkrSkSJVaVHyHMgt
DMjh2mQVijHLQJbQXE1d5aBXwcv4G+esYnhlnxnvT24=
`protect END_PROTECTED
