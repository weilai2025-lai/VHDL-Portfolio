`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAEqID8ZHY0WK0LMcQNougDeyXhA5EeW+ewYJ9ZSlf4V4tElNW+z8CgjxQvT91U2
T/XUEeEO86s8KuT4C5KEzsICj8VbT8UqH9TwuiDEgKFnvfJNW9lGav9x0m5lcchJ
ke/FQGRId5tH80o7ocgZQ+GeMw2RQK72hyruabAk9rXg8+DWnMFVhfi1W9NF3obg
ec44/z1DIuqouVbMIiCo9xUIXvHOcqS77qDvx3q53y/M7RI9HpxfCl/g+yq7ibSz
pqvoGo/q68Z21bExSeRK0W5moBKg9fZNVpHFzG8Jp7WeXEp7CCoF6OEeKjsuaKYo
gTWv00XFTJSGHqeKebhxXA==
`protect END_PROTECTED
