`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Tx9LHcppS8qXgMka3hDuixr7syUAD2AAxMDbhsEfiAip9w0ObN/3uxnA8n4BpQ0
tl72ONyl8xV5guOilzhU6oZeXfrOH7WQShARUhjoqVrjlldHsEOd71K/DQuLJbTq
9HBpTjhy9n5rzjT/GirYdd0lRxTDgFtTr0bkVUieio2SRPyeiVEL/4u3kInoy4rn
W4uiD7WcL6l6H1n5hS5tpSC3d2b4ew3TBd/U1kxcQcKNr8NaUsCbw0TNY3ZfyMaK
HCG9FCGIv9sElIQpFuV7sy0AyeZ4uyYs/2M2O5xKj80G28oQQrTrnxxGaohSfLQg
H5aimHyQBjNNCZK1Rl0hM/1smYO1lnAD2+XGrU3zgv9GpeSzCGTburVmAtMU74JL
r9kLjoBvAXMshG1ICDOFAkB0NQucW9LQ0xKtAgNdA0WApDPZcMjTLhyrihVh7++V
OVemmihbLgVLxLoTlovbzJUB74JF/GtRfCFf0p4bE+UFCFhk90yMbjyYKrehr06+
sh5RQi7lSv3B+KZ0uFqBezJJjcFSvfN2rCGqdFvww2B58QWGT0KhmdPh85QiegwK
VqkWQuVS0kiBTHKDdJa6VacoX9lJczzM6t7clZ6cZOBVeiDGAQpoHlf1abyTWg3K
jHFK0bQYeuIWCOKgenYqG6Oooaet49D/DvD1nPHvdHdMvq4xbBspTH938ZRIrGU7
DulBs4MJo5zAdEH8caOLTMUNZrqrKp4wiveMdfqKm/GG8zEQyUDV6ksA1Qy9n9Rz
mS8y6rRkcFKrl+yvcMnKPhCRvzVcmg2Jr49p3ZZCIbl59vqHddo0PNXD0tfhVOgM
69Jls4MKtxF2k7A8FPSzTaATyGPNHPF+uYPv4KwXYwSU9fAngoB+n5yo7Qcs7Vmz
fEgyd6YKARG9L2jIYtdBTFFMpPYmiNbcZ1tejyiLh84iyr90CujFAGr4aiPHJ/zW
gfzWWvn9AC/Yo5dZU4/LnHKRGmJmVm+sKKRMimufALv0iu+p0ClC6dkK1Cjlo6HQ
4vAgPw2bo0UKQvu8WdYByL5/53kc8pK2Uq7GrpcINqqqYH78K0wMhLDp3m1yUvdn
v21TxG3LKWv+Ma040wbcQU79XJBrxcWAORiBxNC3JbFpgBh7H0O++9Y49v5byY4s
oLHzovDb+o2TryHBhFN/cBD8Z9u4OjjD0CiTs2O8Y2+mFNayVT7rXNpvVrzwn/NI
PVTFSE4fsAPzB2EmnmePPswo4qKsWusVNC+6wn0ljrAZqH0Pt/EgIz/z611zPZk8
9zrXQaXkuXEkh5xXlurzONCvIG3dlTvPwL0Jkza+9jP7gQSWYRDlAo/Sxl9UxcMi
PzY4L4LxM4CpEDkPvs9DIFSBQprWjWh/o6tdmRTNVRbkaqmwUCGs+iCMUvyrbcBv
aA2vfBzcz/es9ZmAzTJgOUplMA545nQ9oKg404nyngnPKjId7fKfQ1pXI87U3B1U
8A7o1SXvOnXWZgGLf9bwEw2/KmLq/2S6uc/rEefdnzjYMrw7Be1ieWLbM06IFHKo
zHlbbIDIPRHNtdCsCpYjTPMw21F+RZO2oDLn+9dw9O5CjB94DwQjcpA4Jn+2X5Np
uHHXKtsno19NGBxiHwTMvati2G1a2loSfkjciQD2KYWb+KACmXfvSpOjCGA8eIEL
VGUjrbjXA/LKcgYyVzGZvk7rfam4OUe1KSXTP6MBx+AGm+VIEXIb53AGc5qxCAi/
mvF+r4XNk/1B+NhsDSvpded3DnRmdYjyDvZPVSyi+/KMmg3aOQUhNcOOsqcBXU7F
7LGRDwGZ0O7ZVODdj1mxSfOR6XZEgYEndUJ8au04Ju9m1xr8m+VNNiH/Y/vzDAQc
2APT7YNShkyredPjXQMrKOWd1GYXsQ+VmE4TuYxgHyKulZphYeE+IB8mcb/Dz3sr
tIyytUrV5dhXG/D+ga77Yly8ZAqvEoNnws6o9702G+oVekO44SMM4qxOcFt3LL+L
3nfFh0S4yKBnZPnxGsAOqpUOinnQyXLUI72VEkfCAxyHsz/DbST8g3wNoZ4kC7jf
CjZmdzVO5tP8nzQrTrwgHiufhQtsMKlSROZRZkd03kwYVjwTA6O8yKPQ01VmGAOe
5jq4x7GcPCpeMrVPB43r84AiAQvoEHKsE4/yNixDXXtwfYcAcPRL8Y3oHzhaMsnV
WnnNfyzZfoyZ2ytGUKTre9jt1Y92ZW3e7/L8c5oFIT3HvDvxwL23pNuqrTj03esS
yk0Q3RS73a4P2wMN9Etg+lSog+4H139F//kDxK0DdB4rMu4Cge9farNmpMi7XAWT
uXocgf/UHK+TbyrwX2cdNQ7I5OXribMm+r3okwCt93XvJv4XXKeqVkBFy4YrumQA
m2HnnqFiHY1fy8GSIj7vH6ulXFUaFpg675xTFF8dWXNH3auHowd7i7A0MBvV4L9P
9mwuvbwBh3bR5M1cYVg88XFxt+60Z51Z73h5rVmU2eaLOEVT1JTTQuCN5NLY/KVk
R7WhmZGfTPpqgU5AGhVLAXMh1mf3isHf438VLMl0vt18+CKmSp5gMqMZHCDe9L3A
UBu32AFS8T4AxZGGGfRaDy+NwJp9WaWbEDXWo7G86MfklQMbJ9GojI1OQ+AyceTp
MvTouk8ktATPKnI9vE4oxi23m6cLeaFGORZ7JAYS9GbmI4WnGj8bzEnqXBP6H3V6
eiNzOlKjH7i9+JDNMM12J4MdcSGWVTM6LWm3Rzq9koKlzrL6xj77hrxNPec1BAmF
l0gxKKoE2/oVYEmLtfvs6Y+0hEo7jAeW/G62jKRoxb/GaGurVABsivu1ZdZvpJ2Q
2Ozzf/LSM8pOW5GiGmG1Md2R4f0mtn1tocY3ijDBNDZi9eyVUX6PhS7x8YW2wWvc
9A0WfluJkp4qoBF2ufjGprHioFW8zxRgF42ecCiOonMg5TTpvAIO+sLk5ukK63jv
jXu/Fc9J3Njrve/IIJ870Cyf7Kg1EYF2b3atGu29qWHGsq2L2NYooaT11ic+EVNg
mpWcd/NYttBvOP1VQz1mtvX3Vn1kNzzgPc4lM5C9gdzScpDpqlAHdnqrN3ZkJe4x
NXh7m84kKZ7wY8MTKElFPe3r8g5B1Yz/23tstZwXn+acImgi4vC2nrlpKPT3olGN
sHG/uYvhITR6T1xN/n6YW/eL8IC2G1VFb+a32Lvf4sf3XHQWrSsMGzNHIXCNoBUu
wJ8mwA8gVqgGGSZWD6UjuOIiz746wbw1WxRrzxffoT1LZPQO/GL2QKVQgfK7hfNm
Z0PeYdkWUtM25rmy6WxiGSS1+TcNLqJd9VNWuEOuYkw4WgqG4/yU7tsijjxmWVmS
1yNngWIDhE/Y9wdMQJQ8DjFRQVVz8jGuTD3G3oF7GIve+v6G2TR56b0EbDRXPMqp
HKzyYbLRgytEGo/vghFn7o0/STLKMhsk8I0ZOfXmXvdm3xYjsB0FVAXI2WgyUhTM
QFQanNVl5i14t3nu2QXkxuLUFgrUVDU+SHKAMC0aTt8OC8CUbeBcJTHUkkWVS7xc
LE5n8m94UJJA9/aWEON9NmBSz8MgiPOgvdG4nZTGmXrWh8sV+CpO+BzReugYu2w8
jE2Cn7PKtRD1hqkVJIU2xFgnbxd793vJ0rQU1Us0uN/7l6uCIb9g1+ILowep2kvP
YyQ+NJNF9EdCduze/wjRftkUrb8SrgN7JGsA9WYalM63fmFnTrINZYwTlxTSjYLY
b/VErTkVwBW2C1ghEu7QJHG3q1A5jQHFhMwhGRkrBRghHm9IbBHTziS4fEpuXIaa
5fjsUyXWiEZc+3WWkZT07AHqTXh/WtZI2Qd61KxmusnlAe3JZaXM9vBtE1+Jxg/c
gmaHYXLWxmJo8w5ObPscvYk//Ha8hZ1qMJS4SkcOd6sf5hwK/wY71sjbWQ0pvy9A
eOGmTd3OW3iv6I7rmXu+bh6fljf0chyXZWAD50l0Dau3pb+eytJmEXZE7Gvb3wp4
9USsxAQROwzVTOxxeruEbydPpgepYq8h6K72hky1MEub24lj6LwQ/5nSMOmFCRXR
ZwF17gtk95HDwfvqw+HyKdWET9S64ytzFupZTw9Hf2UvNZOB5zFRO4fXkoFi+uDd
9a/oygfGUzmPouWRX5/HL4GrcpRGTDtfIlmksnm9CI4151IrLK1qy/sH6vLy6aZs
ZVHvOGRHyxkFSsUnl8PmDYpW3h1YlXqg0mYKqqz9tKCMTxiJyU79IEvR1dPyVOPO
Hd36ogoS6tDgUKa1cWrBE0KGw5AZipk6qcXF3hSQk8OppPAKfIoiazMA8YCyPpD8
3bkNizn4407pX+/Fh0hYy+IXroCi1UWDOgnAKPIMYYPmDU7yH724ZCQtO2eciiZB
V7KzF9qQ/NDxYljn2uLt3HPqrY65+CqR/JWMdYZ1u9GgJiJ+nGxrZKRVHlRs/9HG
XvVTKLW1S6Z9eHQbhzd/QOJuERxo4qWFJdtYL7iXb8VC5kt25LE3ZummH5gjqnh8
sptEHLuB4jWlIrhFOVrTJEfgsaRJo4lf9U2XQA1m3qAp/y9pfAN16qxgw8lHVoWj
Qh3xXp3I7Qve8XAWM1MyCHuN7CUSSlMSk4fh9+3sECljCry5t4UwPiaD8knKb6JZ
1MSGTyxCeoTNDRIaW8O7CgaB5ZQFrWNnDc10cxMnTN7X8x5BnO97H1iDRiorg262
t7p4cMQN7auvQfVaYNi/nFA0s1SBu+VGQjIE65xFR+RFn6fHsFnAaebpyMApjjVO
sNDsEqxoEZdSpixhJC4qZnC7DwhXK6oJqfw9nmcptGZbD2eMjgXnutYlbDaMDLGI
ABV+Q6A4kxDcwQ4GdZxVaw/InEEA3q0QxiiHA3C7Hjr8Po8zVhSLr0uqjc47ODn/
rBDF4GcJ4IgGEOLPwvmRQ/os3+1YcScj8iFtAqhw9lDPn3//R+12tQZcfce7Hf+S
q3mVCNqbQQDeuqGWo26XUAdn7H4gEzazUhujXmJqwmRiIsZIR1fSc6VeAxmmtImh
QJlUf9eQ6zMw3TWLi7j0xOyrlbuf4bn3MypbbqcbCkgeC8gdgRMeDAAetxWP970r
JCJ+rGjFANYuGbGR73Uf33XmfCO+L/kWblN351Q4gzZtChTUOr223KJH4+Q2OP5/
/6wiI7FpOoqn8sPFW0P6gt0oDLtfGjy39pnvlbMmJlLwrFe6T1TTelKooTYd0AT7
1My38bGsfe8yydujf9JfdJahte0Y9qgCxhQSsL/hdd2BwAfKdaa7z018PAoQIKDv
08h8/CmEjuBQGNzuCXSEcLgWKtSAO5qWBkV10cj1lb3XDOL8OPZ+EmZXXDf3AIgv
sOI13uy0qmZVxaF3zoPSzA2Bsz7PxJa0bl6q7rkDKB5W1+0YX4gK4dHJJKDs9O3b
g0ucDvuon8BxfixcIlwE8QOBEH6oFKQpBTd4ARK7gaoj9Mh83V9MiKwvqiUzwq4S
1ZNA9j2VLvGmHoK6yestjw==
`protect END_PROTECTED
