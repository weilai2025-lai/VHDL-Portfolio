library verilog;
use verilog.vl_types.all;
entity fulladd_4bit_generate_vlg_vec_tst is
end fulladd_4bit_generate_vlg_vec_tst;
