`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoQwTuH8S77N0dKuNeniMwuloGynURP3gJnmsxM6k/WZfw6sX1dKlnnfhE65KoJC
Wml8GeNg4wiOS+vjbRfYrqi3uoAhdCfu05TTjpRdy+9up7WUC5uwW/17myhrYH64
MhxzWFayVXUPRhKl9a6wdxfPxU7pim2OXhHWZz+LflFHJryVcnK9O8p6117ZfFRi
Kc6MXc/D62npgXniyHDb00uTRT+mIiVfaqWiMtX9UkflmjGxIvDnZqAh89tbXVw4
TgkGvNi/uWTM0UEHmZJ+00c5e+qI7SSVT16V0wnsZFdD2s5RNPadu5yqbIGiIah9
WmRZVxv+1ofiOmVRErpMyXAPYp+ITDE00TqJ8N4pXDQH5n6He7cKUcR7gpB8afZY
mV9tWtTC1TPscn1GaJuezkaYLRrydyjcNfENQpd7rtpSbfIGuB17SA7foii1DUJc
sP6o8xzcGwIGTIx/iEeUqGnYJ9DGgLz7KFzf3bWM7YnsU81z/WF/uxrPhVSPj0mV
YbTf+w96aoebGtFZbe5warvxK4yNAhEyhwXRfP1rbINfQmIAxSTIQUD/divkz8Vl
lO1E9nTgN3ijULrrtjEJj5qUQGZrlBI+daWuzJ6Jj/PlJEckzZajsiJHfFQFPigx
5cxN0czkP7qtFGUYOaDJufk+pSqj4jv/o5FF116t1dPR2HidLcxs9AJor5WEjKzv
D5jURjWPc4LTIgpmeWT6WJeOn+/tjTcn9cxV9lRNdeTbFRFPcHd98zb2k7ScpbQx
kfUWKa52HJTpQ0UFe/oL/w==
`protect END_PROTECTED
