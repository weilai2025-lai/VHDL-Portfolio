`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcuOsCzO8j7DwoVzUx9VfGXXaAXssT+aTlFZGueBlEi/TG+2ygndw7TA6mRMAL3Y
/PvnnVFgh8mi1QJuNqEPRcsPFoanykGQKqCqnYnbBIoFNgisrhWsVNIhT972jq0o
VGYRdDarxgWD9yyLHubOUAFF4JIQ8Tye/YRmMOaYvuLOWausvdP4vZQ8gTx0xPRj
yU/tQwJE6QUy2hDYHBqUuaW0djCA4gVVYvy/6zUeUUm9n+KndV5SSPq63AuZ14Dr
axvzZnOkMqed44nWTTtTvAR//haJlhkV/NOC/hw76L3bR7RKXCZwVnZRqsZS0uzd
ULoNGmsmzjKPE1q8IsbyVnJeeIA9iTZrBrHLu1IlVmO+FExFICSDBNNqmRPXfLQV
+BIK2mNxjeVTygQPNVf1PhZXJskNqxFFMSitjszIWXbNg/hc8MRU89eslESNPBKg
vCqV90XYJG0u14RUiYnoybf6FoFJvlCFW1OZbNqq0ytzC/DG1/TKERD2Z2P+QQbB
ZDhsty57jXo7lymtx4U18kdfZTEdr+ieVYRNMF6o5rgFDyRRWEdO3Z1kpXr3J7Dr
K0HrOLLcPuxfNxTgZ4kRocnSP7dqiiHhxPTPtZ1U3VWreNUfvQjbiwRjj2jf1YpR
sRUv2RllFBJYF9c+5CSaWyTZ4fb2RpIyNv9+pwxEIbb7CZphHoMjHDtMDKascoVd
vEmm8RDHtEqfnkHN10xvFRvicm91zS/PWf6YN68b0NeLSaKyjIBoG6WDmvWT6Xsu
2Z2G4XwKnWlEgJolbkvF6KTtfNig2A2UQ9dTFfH+WpY=
`protect END_PROTECTED
