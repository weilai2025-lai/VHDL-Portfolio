`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMkynZa4L8nHp9Gkf/B1dQMIZCI4ahJ+Hk4lGdJ4h3rAhiXznjuW2AUwnzO+l3SZ
UCNwm/RxProPVSpalEwCe3WGir8QAS5YfuhBJYr290RHqg6F1dRYQa5FY2qaakdP
4k12QMcAkwaBumH4Pa7p/Ko06vN2SpCJGb5vfQMfUnHPv9F1+lsNhhhKQ3S4dNsh
nLt5dQBfg3RLkPet+JNsBkkF0uic5ko0hti7BZ+DTk7RUEP/ugHPqeBN+JVHwExL
fJV0E6mKmJKrt7v5Ll4X1qIilZbzjbb7k+OEEsjsQbZVnbw22pSPWd8rrx2agSU9
/dHDKp5rU763xD6C4XC5QT0Lan32WG1b0fdWjcV73cS7ZF8JwLfjX+EvTfYd6g7r
cRaMHJW1ltbF/Zs611CAf3jOpo0WKyqBCv03hhZILri8lOBqfHul5qoUu8YBSNfA
5PYhFBjldS8MswxYXZt+rsbsh+DOi7t3mabZa+hkpiy5EqFlWYdPR7NQI7DcpMUi
ztLjjZIy1V2DnKYxGn0COo/Xh44E70+VoXIwMQrkZ5DmA4qcCxkqjykoubSzvCek
J4rYcDEFItQxxuUysk7hDGABLMXgyT5JDBBkYA8bEbRrRLUUDnhy2PEIX5filMFy
TUMbgBlgplZcofZsfKms5lSi4axvoK7AB38EuBHQG/AgiLdODwUeDYBWSiVhfVNJ
uvg1sHEPDjppDaVBXrVVlUV+EpZ+h+NGm1BiJHjy9+Al1zBnZvWVV5mNAPucnw6A
4fkCWzn5gXOXVBNMlJC1+C49VP6DTNHtheAuS7Z98kZfEy1vVI8phBgBBPnajBDE
sbQ6i+4osEMRCBY2Vxd7gOl87s4yDOj1r7+U1fF4Icq81f7UE8qJB4v94/HQsnWN
LBRGElWOEl5Ebz8O/2+q0ltpLst9pcewHvCLfHEp6/knk94rNV89SJnjYlxMuZHi
hYqhjQz9jSJiB69jYQfRPvGHHTDqRQIPoGAMF+9UKsQuJF5kP0FLLoc2pWLOBK9j
Tm536347F4c6YOyTDSYzDS5S+NVpN6H4thsgBHynqXSF/p2X0/f8aJtChne6QzYO
cTyXOW3olBJViYHKpxfWPylcihTfKem+IQoujNABIkWHfegTn7WTrjz76geN1mo6
da5DGTIx8qNxDMVl8LiwD+PEX8wrp0xas+hmOaqf5zhzTLtyEmDWQ2Xhk4T3iOno
vOyQheNpu11oCu6mO8vyAZ+vIU7UJ2xVm+WAedPsQMkdFEZnANd3cu6/sStU8aHb
ZZ0TVOfGtE4zwtx/xNjRyApfFXLyMHa6lju7QhashcpTcy2YXqz94M+3qSXcm24k
Ea37w8ZqMLQ+60AlQzzOTg==
`protect END_PROTECTED
