`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2WqR9TyidJg59CzoU3QxwFF8t8m6o0OZm1Px8/z9CH1X576cqowUlQznNyuX9o9
RHSDfFBeKGn7UP+ATWBLLr5kOMqMihKuK+0p6nTX6m8DDt+Fi3yJU+gpYlvqNZz4
AQ7VX3QkEe+korEWF2GzPpKad+KqqhmiXf+mFnL9E+o8zmHO1HcHJsETOReOeJ5g
cuM/3ysa59r//MvDwbaYmtDqWKlUsGrVfGutdPBIyQNxyrFwGWr3Rm4vtVejHzQc
S0izsD7PAX+Zkfn/UAw/Q85ZRV2yBz5vtqoVS4uNTAxbJVnvnUTPtz8EM1WY+EFU
1IALAJ/0ml4/iJRrqtJkOHjCN8h6b+36cZ2HI3zjiWA78m0tpyRaU11xDt+McqBI
bLlv40r1IktWylrb7hPQuyNedz+A+sXDjQi2i3rYU/YQWFLeRRbRTItouHJCtCOs
n4e38XsJ+FKdm8nRguOrA+wykluUIGo3Dlj+28NzKODGN9J5QRwLWymXrcSFa6DI
9eAc5LM7YbuA7nwLuKuvmHzUW+DkcvkWEZ1czSO/LtnneSRjh6voEDBxm3mbPvGi
LWhjQawT9+sVKRypUDKfUfOn5orm5yCnxdOcjA/ZLXgTB60An4ZQo61LxEW/uZn6
`protect END_PROTECTED
