`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjIgwho1MnoB910TdL7oI8Hb2z0vioKf9T5G/2wUSbBOpiJVzllTHd3LUZ66iQux
ZWApSn1x0Wx+XQV4Pim1gicNuUGFNu2tH/DcV/czZRYFYaBokoT2PKCEa71K0Sqm
36y1ablwiaEbJ62Fn3MhJnKMPtFRtlxVX0TE9uNdzWdjcBLkhF8X2HQZEm/xISB/
Zro7S/URd0QCuuCn1ccwDs/sP22ANhcrK6dElsHMfrdKjd7aoQdQbKMfNyWtnMw7
RNWc+nRMdALR0PU/8iqAvWLK48OroSEdXYAFn+sAg9X+9g3iXOYDAMfkQQdLUv4f
Pz5gGM9j0aWhJXLgtUlKjzjxAiOmEhvm/qnFxcJWVwDnOmszJ0Zz09B2HiitYsTc
jqV6Vupe6tu1mBVGIZNfO7mbm5Zl5Io5RurdOXKAtB7PTIJkqLRmjktWXz0ARnad
yo+3gp+4JneRuorYvFftQlZvlGk++ReBkFSQY7xeUEtHQQh8V5Qmj9zjSI+lbJVk
ejUP+Q4TAWRLGZ6zUSei6oRZjRmQCyI8OZk4zWWe2MmYfwM43fsWbPIoywaJAmpC
tQ2FGumd8/e5J+3JUh6k/FASpDWVfjWWo0NTF0sqqAAH2lLEdKcSc4+NCiuOoaYg
dxfbiFRB9wYSKiYFV5JLaCbYJfEuWrJBy2ItctBZgvGwO0DSwHmaRjX0hFelvJw0
w/OH/SGyfQctSgRFxqClOP6w7kWmSgIJS1x5znS0QaqB9XsMjonalUcGi2BMmmxx
BkAEEmbJX2lAN/jzv4NBcDFqXfrgqLjkfLono5mP707aqYR/KptJOdwdDpdjlIXT
5hA2KMkJfjZfg4/3N6PhQj5+rxVOJ7SXKX9WWdQxo3CLMAweHaj9s1LVbbfNDHtV
Evqg9AaH9+KkTDEFZXD1wZ3xn2ChdQnXmj8Cl/4j+C2ElmazmQDoQKm7r395Cpqu
+XLCs74/n6CDWjo1tT9isXSVaQDqaZ9uAfNgtZI24RqaaP2SYZdb8VDfxwjP3SB6
buK786bnLg0P9z9SrrOcOnaXS3a0niOQyiM+G06GVzhkuWHJ4HmJlBwElA3ZHLpr
OeY9GfOB9+KKabJTYToxyMaG18Di+5IhTXNN0MM0Ino8xeT439GGCBYOL4ZZKjXa
oDlKiv2sSsy8cSMrZJscUNsw65Db6pEjxxNJ0Av0vxT2YpCEsFce9++9SRSJm/WN
kVEPr0CjkWvXWGh/8yn9NlTQ86LqJ/rG8qoU0//cbUtVBYDcV9QIdmN4xbStY86X
Q9ZDqSNem7zhIEp6bFmTfkNyzLFNr4JrVzAazKeqohl6USXAXuqZB3j8TFJON6VL
N4KVhjsSN4OQgow9C9YtVGJZWD84nreCIXd/jDXzMpap2oniTrEb1YfmAdvHgY4T
F3Z4XGFamuX9nA9nbEKjIkE/3FSIS7xkfADuHZvKC1A=
`protect END_PROTECTED
