`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOvc8uVSSAcipUFYb6xlEZwwZcuN4tr7Ug1pFBXYq1pgnq1uvMT4c79c7N5rkyEy
pQQIfFN73h7NWkxtUuv7kO3uRziLRBjqjxH42neuj60iamSWBAnUIdi5FSzRQ4aw
2l3SSGOdTm7sKdqOt+oVwNgx8yQ8+3AWJ98qSzgij4O47Lx7cTXgzAzLRBA8sJrD
1OJgWWauYzs3icMaHkLswPp3k3l36Cny7mB+ADcXbFGnDkOXnm5oDaPaf2ORZuKT
Lbix/WIY+HnRCLLBq2djyBUIDkO+4BGn+qhc3bc/wnP6YIBnT9XA76WTbRsbb0XD
3G3nC77fgPom5jQbaFJ/L3dy+HUMVvzl+vexgEl3IepMMmLIfgmhgpzU2CaKICHz
jzVyoFWzpP03BrWYZVuiGdayPaZIHOJlvDti7+42i/43WmP0a3eCVFoi13u4w3De
J9MyGtLpYtJNG8EzWDa03CGcPRiHCKkEGyAXPtdqXxKcWuCg2RihYUK1BgueyV2T
vo8tZojnrHa/ZiB28Ko4yebTdYhKLzp4GyFmuzOTBRvYYhLwes0x8j3FsKS8Z63J
Je+zkZOy8KhQpql1ZJSTUNQacxifXILO0VNFeSjab6oMx0n4VWSb7f8iSaVCCIWC
BszDTKUEDLF71APJHXrzyzM/D0XQy1WQOUHed0PtXBfwoCIet2ASz7ayvRK3BU8j
duLssCgcDKlN7SNxTnc9e4gjvLosixw298jICLp5qYzM/dM3DHFxCuZYOwNXECfQ
EwOTV+t+o0quEe+BH6o3lCv0msGzZRi1xvrL3ndBLLxTnugiPMRbWTj4AL+J3xF9
wY00TLxwpKvgocaLPMiQUbS2asAhMadh7BqLEJ4i+lmkXdoaS0pxP5V9P9mqFxM1
tPL/zbnXJMOKdPnXB4f34NzKOMBX+Fjjirb2ysYi93h9N7Rm/gpPf2QhwXBKvq9C
Rml7V6T0XXuEo931oKimeoFHukYspNk9KdNGnAfAi+hiRjTE9NjdfCN+UAkRcXOr
w+x2281iqsJy48PYR1vUMFmNx3lkyXpx8aB7EqbteIxy49mZAEpZjSeJhqSLLfY2
EEGrOAJ0j0KQfewl84aOokWR1CTLcP/cFipAyYN8TUSrlyHKuNubkSHmU0f7Pr/v
LLcHRmmwkxkXBOmbLGC7WJXYwu0gnVQLufqMZVtH8hQXPGUmwY11/8/89GPl59Fd
P4dovji6ynRLT33Cx9wX7BZyfX+DfXuw/DYVAgv8B1PZkPT2G5QMavjBtMGuvw3/
r34wUELK/zYo/EekZEjzK/ojrZhy8TnF4mHPZ1Jo5bi5JyIh0a5+Jz93GZqAwbcz
0BiGK4OzGqHmcIssKhIua+5U4FjTHXOWlwIU0L6T1vJ30rCsNDlhGatGVptP4R7e
OwuXcZtrNVmJ4hakZdp9L0rZBQ3BWP3O/oJrugrAgawMutQL9cgzOOCI8NDQVLZ4
U8X/Sp1XXg0FgakWX0/R6HdYnG926415vb6YR0OKraXmJnFLFfkKuYGHPziFBMct
ZXyuMrjbUOmRHgCagiEMH1rBVE2xcprGt30tgXgpVy+6T+YuQc40+KH2t/QNnFqT
9ORHQt9th4iuwn5yopKKSNaoYDE+fAImUkxmMn+jnzSEqGfhlyh/muzVHFxb1fTV
ZMy6F2QAKP2G9jAE2qr6buCkrNeFhjmsEKX4VhQ7m/jQULxfEqmPzcTJHa1WhqxF
inGmqHf75P5dlswS0VUPyo9CPkCpq8jF+jdalFmpNEWYkUSWIPttZiwZKN9H+fch
tlK5vj8cuwHemd/o6R+PMoK5mi50GH/q3ixoOP5dOv/u7r6JVUo0JQhrBIazbxhu
nwFmFRK96ZRet29fxIT1CxFV/dI+SxOuef3u+TpR3SuODvqdGrrwQforBSRSyhqn
NGXIsxho7F9vuTtuU+9ecNxRyddOaPKYeutvq9CgmQPHzh0h8Y1hMpe12PGDYzz6
VLEBnMTsK1USOouxP4sPzXDC1t36MlsJxGyFiXk7idWtt2q4nWPV/D2Gjp/ZuBPN
Md/2YlNyTJKGruA+02IrHk0LKc3g8x+/K8jR55zt5MwX7EeM7A7aB/vCzdIJyhss
BZp+jM/f5pjFfN3WXSZEmH3D5dhwcIL3s4pwCM7vw0wichnJcNaz769ZzcRCbfRq
tztxOQbJaC+Pxl0CoDDnmVu40eC1/IZbdUl/J4t6XPY6Tr2Ikr9rbMhhHLzRPSem
KjO9FysHdj/tFwX4lY1WuzOCYVjR28GEVIcs/GFTeEgqipcU1FxfAK6m7GDcaZ80
rCLTC5vemEST2UMjBFNuml06R5yk+ITby8qvacQGsg1k3SjwR9qSAM4BgxGyruvl
MPnmEMewBUmta95vnjM2ERk2dIY9BfTO3R1ZlKzyVvcWiAwTJ+1XG9oXj9g1qzdi
wFc3OP4FWqw2bgSFEmjLGRghGXg6zXTzn/JIK4TvCSNbYDADxJ8mR3HO8eLZqMtq
qi1wgnvASwS5f7WAVk+OnOFbAjXRovtcIsEt+UHhb/4FhKxORpIPccllaudziGUv
eYefXUcgd7F60Y40SoHvSVlONGGNAYrfQ386u/a+q/sbm9cHiRlCks+I95dSXHyx
Ao0ZTHmLpruIhy3nD57vwDVPFXWYkSf1TalFbxEju1z2D1AnTU+Fmr6fis2jU4n9
7wjEnDhVtLL6mc/1GSYTHFI35lJRt3jUW9eh5dFqUBagtQt7BJluVH6Ku97OeIbF
sPfRtr6lHMWOUSj8H4ifZ2PJbYpM0EbCApHSrVxv24mf6W2sZir63DVTjjPHI1xi
DfFrBAdfH+tq7/8r6o+lSIqM8cKD9LDHiEgBeqp1STUDV7dRGS/1mFTKasYLp49w
E4FKB+i1evrS6C3eWvHoahw686YokaLmB+UY44sgaWZoD6zO/GRWKkqbcgSNEfDc
0y6EO75PAHqys1aAAd9WCle82eXCV0hZgRU2liod982pOiO2d3md9ucO+OXQt/Px
VppbbKffGcZYziERDN4jHZObTcwGLco2XA6z1/sHLQrONaEUfsnJxgLsB8Geejsj
9qztbznj8XoeTWdiGWgbvlm7U6f5JVPZcXT0HVPoSOJ3MqQ08CspGGWeziPqcCIG
K2Qn+znsvfw7KoEUNaut6+8AnvdntQM03jW9bhPqk8t4qAZaQUyf+0R5Q1/PJgqu
qLWCXwRz8kU0o7x5pGWPBi2YliTHCwlHwphGUMDJOCO6j+RZ7pow2O7aezB0cg50
LmxTl2Ng5aPnaCGZbvOcMMMyOE8UFP+Z1yinxBlkQLA9P9Xraw3+c6+nkVjyy+sw
YznlPDW+6ggf7VzZxKm58uiqLjCLWYWegHbYoAShdb2DJO9k2fciM7vDzVBMu6Bf
YkfXwxUO3zLYXMkriJS2HpVQKJ6Ifl1UXZYix4N09vtT9S57F9OjAd34tcYI7ku9
H6+6bgO1JTABOadCtdlKm12WI8WKXkuPuUh255xyaTFmbHv+YZettnQoS+nrflYp
dgjZlVmA324mGLsjr181YnByokMJwycTE0412+Ywfyip7arqPkoe/JO5endWVQx6
+IKeAYbImjgP5Wyo2H27ZjYM3ThwdW0M0lUSCDd52IbHyBSz+GhbR8Rl8/rC+NGO
q98wrDGm8rgK2iRi8u1f4bt19f77vbC+r/4H51VIcXWHdMLwx75EOf8vsB1VMCEN
nVZ1Pfg1iZTpnDKnTzf0k8CWgMY0UY2NX1P8j/RNmLh/W6mV7Z82yEAer0nNr1z1
gSneCAsmDIExkFCjYOssEcz8pv1BEtm2w0oUwpanTmVllhLwH4Ry+a1b9pyl4K+/
fDRTSh9VXZsYeOxlNopJI6kEcR5eA4XnMZffVMA6FkL8k2kYwgsYdVU2uk/g7nJs
360basHQ7yMZCBVn7UJL7qwPM8KTFP1z+i2Jhvu8N0cLAyCG4ElgouexpNrGcr4i
33GnvyPstT3ts8ay0O2KSOj1jx4xUDZiaJZ9zHLzlTQratkcu+kGmBxPl//R0Sln
Atseki8W39vLg5HDfxZd/L+yUezurHhq5n8XWfupfllWZvuRIGVTrPkMZnR52S2n
wD2IBCVIOm1MhsJPsooEaLP80UMrm8kzgl9lzB73JBw6L95KoUIsSFb9siHFa83/
qtHAOnsLXCvXEDWVDHkbtRqvgXRyQw1gHaua1eDLJgOdVBe5eduJjLnmYbt5OfW9
uJqzthEmCBQv88nU7bhFN4v/pDVvnmGt+4Q04EeNLr5W8wR99Gr11M5LCxkav2cP
QDWxvMA6kLaEh27GAt4hnbkhhRk5p4MYgrGthyn9tUjieDgV3s1qGSTYSClM0Aj2
XI3NQpyDOxjCf7UqXQbPhbIWzxm1/3t1Z0z+3bRLOZnCdhSU0inEuxujHgfz1uoI
f0ZCuqXEV3zyjV00O0GIoBiMYnKvbEQmyo3lDf76muEHh4q0xrlQ9SPV0t6uDefq
F+LKJaIP82CMkGhMZHYV0nq3Zr9NxpcUP4okf0RCPgbY9Upk6meQclNsx546ZtKp
WDVCq5l766Mi3DtoDpHuVWJKFIhMw3P61+PuPZTrMRtGyjAVZb1h+2Znu78xeVdp
Xj2fj/DGzKcgWvq6tqMIzOTFzcUWkItXaoVi0HpPwm7cLWr2TWA+Acbrown3Wto9
j6seOLZlW+4hfJ4xBmvkeFid2Juo/SNvClHleCWbgnYY3Ea/IL48yDc5uPoQvWfU
CzqeeihyVTzzEavnKvEIqe6pTDrZTA474K7UGeI9ln3WZ7junI0uK0EA157AuNYR
TkXg8ZGAGj2clOPWhAYS4cYys1ZbuErMXAgRW7aV2Ucn7JS0NNKyzNswADK/9kO1
k3QQ5fTjDFfPU9t28VeIkHEGYz4uKLW46POgMSNytQMb/Ya9kOOPcY9ZmlQVvvRw
gzbG3hr/l9VKWR4fXWC26JwXBmawC6JCrKyk5zilekb6irkjgUj/HUBQeDLRFgZe
6kQBNnQoRllnp4UCip2MSYj1j5hAe4Xzgl1rMl5KcwYOMliPKHdH1DR5NROhozSW
8T2RpyA9Yl942KNZdmz/LBxZ6A9SlmZPh6FJkipI7Bn38UtV1DNXhD7Xw1Oaqm6o
pDaBJr43f/A9WvWLTl0l2E/wWMjk5rWvHawJqLDR17lWBj/fUfMp2gqiu08zd5vm
fNVpIm5OWHspcryuKy3G18MN1w+SErrxb10v51wNbbtocsvcNoh99fjX2/NIJNbr
Qnq+//X/4gmxO02A7vgjBHUGmXddNpQrcJZPr1q1lLi7yghr00Y1q+UY0BCaRE9D
QSdlRC339CzpRmzjBcu/YG8GlwTYdd+yVPXUuE4tlvFFOLKce1weCdsr1DPOZyDr
IRxH+vzlSRcvW5pkJM1o5PLov4+lbhLQQbE2QYHw0r5Pv2ZStlsXnNQ01wHcnkhe
0tJTpqUhGbIO0Yz2Nw17k3+AFsU1XnjL/7gQzsb4OjFZZhLIwsehaXyMuEnUAGIw
HSa+axkreW5NJwHxNUtguU13ZtIOOHzG59Jq4T/4TY9HfZXfG+3hCua18LlQhuZg
nNAj46cncqjmtkU59aLLVtglKXahpUdDYXffuAYpGUJPisi95hVrZFE/BQGnwUng
ovO4DwiMRh6jCpq1sbsMP6gEUDfhT4tS7Wfb7R4+Fa1EPgnqsciGQ2t8Gdu1SPXG
OVbuE6e7HZTl9/JvrRg7rQB3lLGXRKaegoDdj+O60XImKhahFNZ5t4zuV6Vv8M9b
W4JlbH9kW0kQ171MDVCSlV0HyLPmb5KYS6MunhzpMdAcB1JjA/7IHx6EdDZ9r0pW
agc/gYuzHg04t1tgMMjstw0/G9SEgjTUJM/ThsQdThbeNspfa818alfvaq30gylj
iXuvuSa6Y/HqSl9FUbOQq5Aoy8jLOIRRpKChPI2xq9ShB3FgQNHe1cMZcjQQs2Gb
kbDjuFMKqqweNtTIWBiPdIkdyYJnOrG+PdrBpbf3mQiQuNbS6m0HmMcYqOIzYy3s
cdLSTh/Rz9vM7UG1hnMwfR5dDKr5qre5ZA1a/YmeG3c=
`protect END_PROTECTED
