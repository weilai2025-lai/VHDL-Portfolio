`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+F+ifDYOn26bXHXmS1HTjTYlAqspAw2pDMXaesbAVBWs8rjwdTAkTlDyVGFRXqr
IVLEcvPQHOlNOIM7R/NKWpFElqGlgg7y7GgZkyLjeJLrsulclp6xxhF36dqjkaJn
qLqVHtUHB5K+kDb5d+VfShJXE5VpBIJQjGnnNbO1Rh9aYqVAd1+MICaQO+Bar11A
v/aUxasjan66GtV2G+tOmus8eSaG/pU6GscN5ojDE5OJhmZXlzpE3CRTT2aJCe97
DUvcHPGxUrHhNDV+LxqTSArD3ozNfDt7VERV96K/0Lw52Dx0ZWT1Q8EZ2cSz/hYa
LdirwXODkl9hD9em1CbjKx1zrqf/PmvjeW346aI2gh350pEQxuqgMij9jasAxI55
NinIEpL5rMRqE1MmN0/U9AYB638ZWeiPZSW4qx+s0hBMyQZMQgKrkr9okqwLtVQs
els4lxozz64F6YbZwSExeHbOE7+huIv8hY87Sxz6qKZwAV47dbdh/dA6b4xPXau8
P9WQLvjo/eR7ar2+mm1qlttbwflIMApNFA4gH7+foPZ2AciBAOCzKUxX/R7/hqAG
RtwUx+MyjCrdAd/J+wJCOIJ85DgzcTUXMcSjWo9m7tT58ZWj2i9DWFobfIgbfjr+
8Aey1rpVU+KziN/y48gx+J1f2xbsKljt8j1F7zYqY7M=
`protect END_PROTECTED
