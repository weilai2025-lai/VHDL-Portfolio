`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8TNPWTsWDS6Cvq4je8Tc9Nf2QRNetzxRHdwdOM0RYmTjv2RtZ9DtzApGhFTqHbO
kqg4m3zrpUPPldjBAypmwGVI192MXucf1kljCqD9kFXBOoSQWCU85fPqAqzI3vqN
ibqFienb75eTzNqUWPztBghc2AnyUubiVW92kzAatNgtHSAiFf7RydYdQPY5gEGp
kkNJi9SmH/ZaO/ni+8B86BgFzYWNSti/SstDnij0TeA78aLxBNyDuPSGDOdWlRQD
ku96IesRw+5whZYhuan1PZXFkU5Ne9XIJxMJ3TCjeHggACCLR/Rp+GYGLg2hSS2B
CbbFjP0hy2Nbj9DJKNt91dUm9SkqNiwOEOCJjrx4A/HM9muvkCEe/wpmGp6cZSaN
yJ56zYF54BwRD5PwjFU5qLz4yJ3RxSVwBPdQFcZp9BzbM8YxhcMEivKXxa6ao5dw
jwWf7dB42N9fqN36f34AhkqixykPn51cfIVqiRVPlHa4LdBYFnprayEB6seWBoGN
LYP0RMVrCn/Y7dBwaR9B538eZT0yQTviWWfEfwT1e39+0y/94rE3guBv8tL9Ndk3
CHf/WGf0uppdzQzusV1OsYsultgNfLj+660Y4acRtGch0/1EGsxPF8eAI9WCLVgP
qxpL4Jsr2AUrRNGL64XSvUeJLobQYbzMlwLlOjTQ2ghEO9FUXbYj92ezBn8fo5MM
AIMbaDztyEdOba8xYywfZhqHYUOG7KAh0DDLAOHEnW4h8ytZgvPRWKXWUE9CyPUg
fGToxABQ8OFfdQ7UF4j6P327qeOe+pNL1el5kbiqEeusYtiJKjToNh3rP2ACXEkv
UypxDfbWxWi5g9vS6ll1kiMfziiY8uhriZAXR2xDxt2O4Xqxt3JKgN6UF5SL7JmF
RXvP/9DMEq/uuGJg9VH8WvjMiHyY99dqdbpNz9fKmHyH6e7YM/sdBUmToSonvOBE
J9doIYnfzS33g7ulVWybVmdk8slBUxXOUjjJROOOuBa1o8iIOFb8SZNkpKeTEnNA
S8gWvR3STWKvvTZr0gNH5XdMMxoCKC/MngfmTT4VVJVb0zSSd8Ru5O54zeXwdE/z
w8a2KTPgR9wt/5vPRLGeEEvw4vkWDg4yjKkE6BU/UqHwR27aX7qPlYgFX7q3n4aE
GwHe48l1UXV5B7IsUnVa5i6lyiFhbiachqzaxbhTPqAvUTltZslBwdOy2++WI7Se
oRDsApFQRfMj5s3m3tntr9oPyeNUNbB4fUTOhL4tKYzga5zSsKaZQW0CScfdZLCs
`protect END_PROTECTED
