`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFm6Eew+ass2ddO0cT8bWMPPzaheSXnz4kCXwx9hS+Y6BUtKh/q0jIoqOFYdd9J+
flSsQaHVSDho41+xorFH+MXEL3w/SVFrCD91F6esEZx239IuzbEvQESG5GWxbBJ8
R9rnCJgwTd8HFoeQmVSoStjSfwZ7E76GQssg0EcJsmMy1PlNrnTwFjJD0bYMb1Lx
tLrJYtDp3bD8I5/9/5EOzkvpuvyeoX3+73T7Y+7gQDZAbzWxtnuXo1bQ9OrZC94X
74hbRQDqzl+ClYMTzjGfOORwWy4wEcT+xfpHvlXJieKDkAfj0EDpL3IEIeU0CZ6T
cJfWZpUxceBZBiGbEu73GPQct4AhQLmUOuJztFlX1PvbuORUXVFZFRqqx/uaWChA
cabVDukgEsgwmcecOW4ryG2s5Qt3P+Zp0aPMkPd9FTnBsE09KYQ4AuEfLzKD0dZv
9xAldqocW0BOOCiRU9xdQvWUUEDoMNUerYvnQR8QgdC+WnhuVLkiyNXJ7vbv7YWx
TXTP17dG2ch1T59y+ipKmbyj08Qb4aq6uwO1EFcTP5Y=
`protect END_PROTECTED
