`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmNRwjakASNGVNZm34hpW6apN+ZJm7j8HdZhxevto4rRzrfCSzNKaK+GZkfA5mgL
/0bkiC8ff2hifgXQiwwHD7ZpKD6YX9tJ35fBgnP9NZw5iz38cy+aVcwEvehIZKuz
sq6UeCSfuNOf+DH22aEkdvwZZc+kNjNz9GcbzYJeb+9yx+cqxlLGNk13LLOet9Yn
HaQ32GL+jxTyxHHo5S8kAwbu+sxB3VuCfqKRc1qWRl18zKX1+1KwUFzeRBDZBe23
UlVMw8mAmC/6V0PuOZTFf0Xfa/KnTtE27Cq6k7KAcICCQ1gPr7lXbsapDhANzOQ1
1e0t3FztA9cXW/nwBWfcz5gei7ShqR3336H+xGd6HEJci0meRrwMw66E/dWCSkEp
+PZirNvKW9YLDe696s+GSDRmXK35i/3oL0zrfU9c+AJohBZUtJL07N5lbY8J4D3D
gW2mnJ6l4b8v9eN/vAyYRhMkD4cQ3XGXzstaRcIe/jL99P1peNA8vHLqM4/cnDN2
t4uKtQsbWwRcxP3+aFP/aqqf6ZrC+Wy22iL+zAthKia2BvlWGH82v4M/jkrbqSK9
SihkeQP/FXMh6eZjazLmh6jMnO7mkuXzybSSN+qiiLRXPNNDIORadHOsxB1eQ0U9
9I5QZoPZvN8zdVssTROVYX+6xqtLrhIw3drm3RyP1oAngKFQ/UyMo/l2xsFWNCUC
hypiNXvMnPy5F1qyoGpEED80PvmDWx+NfjGTLvk5NEV/ZNTvUyBYlBo9aZfsBSUZ
N+tww/GTWstAzZJjB2sSz0vF3ntTdjoALzGEw9OuIwn1PxaNSSC33/BeTzIOfZ6H
BZPaTb/A3QVPFM60eVPYslv54GcA6gFOneqU99ZEtHbflDbKQpiZ6XJ7jzLrOkry
J2EgAXQSYWLk8Watdk3WIQh2am57/1T7NGHMF08pmegXCAn5gXOv37bpiYi4jXPy
FnyQ0WN3bdtNNjkXZRZVbx1/L1XXsRjnPPYWuyF3hkIlOeZ1xlOdlxSgIWNHghYN
PyZ+H0pyHAHhjF3eW/YBctllYn5lM1jrdxPUc+gzTNtsaAUX5RnmF5jhDd3LI3GK
0fCoC7sxKqdCoHZgMxQelXRW7GgE7PX6S5ZgfHGIQZUClPxlOQWsRQ3jl21VHcjA
a4JZQXi1fvUWnTFV4zVzyE5bEmIQxFGlzCUhgoIU5Z7wzqiPK1KmipX+v32wDFmA
ZZlIrPn9/x5poO5nIMUaGtx6cX12ke5i9gSnUalAAwv7OChBeuUn9Yu7NTBlIqG3
MvOC7xq75gvThIGklFkCfiEmvMYgjVzAHZAQzUNZEuHsKPsJRet0Y+gW8QCuIa7u
VvYRkCLAAjsdR50tvjpFnm8t+zYGKTahJ5qPOYRm955gZGmQS0akd64oDPrdHuPD
M9XpyP6njIyl5yHOTGl1fsKEsgr4PbPxpsBVRBl5z8iDlgGwrucMNTizlWGFFzzh
JEErMHHRIOMX1g4Z1J26c4w9KE9gF2d/85bITzQ/uIEPHHPa0VO9xf6FTkNs0pGV
OVmREwD0xH2lmDCORRVYKY/qT3wMLMY1RQgesP/coSCppVSKh7bf3m4+L3r0g13e
mvB7NipYwvWKchPc8Cr/qPXrsCeTrTqEUyEkemm7XcOxmGSyAkSV6BORs+GH/Oy7
cJnj2FpxilJ2FLHwyp4b7Ym0hNNw1EcFH0DX/WR1REgFQsUgLe7S6LCrGpkQvtyn
Cagk8fHi8aMHwDXvxd/9wTrQ/hrLMCmGSJwJLkErD2DEbAXfycsD412pJjEVRrO4
8RiOCNVhVROkVAXyc/vIds7fdZUThZiR/6GkpNWl2KPYod1WWJwuGU2CqWagBPLp
zdzz0OyignF1rqmZuJU2BcR1Rkrtr4J+ed3U+xnlQ8sHc/Hsb4rUc+BpvUUpzTpa
Cu3W+UX56tgJo0fg985i82fE91peYIxt/IZrAPWGPEkEGCKvgYl4AHQJsoMETFew
ZJ0dqizueQ9iwBGofw48PUqySD6QxfrSqcZqqlT6mVEcX+bWDjB1grDYl1x6D14V
uTVzQ3YYpfjXwo2e91DRn9TpwBpDHdjyyMgvHh/ubEsxyklPtmyv+bEL7gC4iT+Z
oi3hGfZE6EV+s8BuOAf8P2wdwnSmtHVDZP740ltZ6jUDHE4CaDLJHF45/kpwwUlM
QH7hZDfK8RVzwKOzuY0jEeU77jZa2FIsE9bk76cIYrCcvmjCUiiyDyrnoP30kJ96
V+nKtifLt8rPDEH200SqG3OnyE7XHiZMFWKrfBUVkECJ8qXSH41j2DgWtgEBXuE7
aonhkVzI3H494w3kEhGn7ydeYdt/Gy3f00fuXmsut4Ep1MlAIM2zuy4NxKZhDbhO
C4+FK0TTPunE6t7X5NuhI7YsDd2SgW+2AuOgSsBxSUqKu8Z6XKhUZRcYHsaYvagl
w8G33B8AR0YGZ+/LBFEkVi3JM7vkSvMkRF3dkw7hkOy32lCJ9a6Xs2+q+qQDPsZd
YsyhhfWrj2vcbQhJOLF/W5iiDUXo+tC4XA0Z/yWWdqytMnwEkzT+cwADeYkml4sE
r/zSUBW6qTsrEe7/qHEZP64ZuJB0WSBfxZrZFipvhCUqNOEM6m1ywEBXNPxtssDs
QGFkvVoKGHGSQvykOCaAs2o7IdpGcfC1xim73xO8jxc72RQX16/8UnQqyuxEkVhu
nAYaARYuC0oeCkB+DD2Y2H4NvkG1ApMgNKT7L5KhVXeFLPjYfG44G0Uk1VZ8dJ54
QPbBsPWjng+TLYLHscR3mjYd9g9/55brKMRRwAHJCZZvlWqti6tGoh/1h2gH7UVT
etzKiCg7wNFSroUDumM7saBKOf9FRmcLMi9MqdmVjKmDgQuSqnundy6/5AqpHSaE
HAL9l7nn7wrY+FeYFNvjqIc0egi4fite1t6pgU/s+GvdgyHbP91MeZUbFgixDQhG
P/RgUklI3jnDXiGDHrfKA5/xWdPRQHEXRnFycurPDGCfLa9xA1szU0xIAfgAHOiG
OcXa4zih4xKGEybAuKXyuVcT2p+1nNjaA9FWVnoJEyUNzQtV3q05QsuUTYrLvo9e
oaUcviCyAayHspnMx1/f/kQ6RVETEsC5Y0gq4bvXrsAHoZrZJOtZSJ47Q1ZZX4e9
o7BXQSZbgys0IQRojVPYappFVID2x/qdLPMK4lK7AkATYZnj6g2N+eDVRP006FH4
GnK+7M4kl5i7JTFYl5EtcT9sNTq7un0ZoUAdkGETqaK9+e+nylQ/joKhN37QT9Ze
ubcEoTZHZUrg1UT7Ifato9pGBvgZi4EdGYr29/1c9EibBgWuGrB/JFYU8k0RTfqT
nQ2otfTiqq1otjDzMCytjhyVR2nYvg9Pn2ceDNvf8LnnQEMxm2qg3JcBB8U1hajC
IUkRevDzKGqSpOvysG1i47yKiE/aYbRL53ohrTna46RrUQqDTLrRwZb63t/1GWr7
gRw9uXOShULPB7kp2+o42TrZS8JgKg9H2V3n9N0Z+LBPadcP4THg/gQ9tBoqK3em
qRrczJjJAJyCS6iTZk2OLIjgFe+XpwMCXqRjfL6BuSqtm6srEF49I9yXJbYhBSy8
bC3FgDpagLGR/mseyrmGNKqURtgnDamZqI8Qm1sFZWrTQcXO/jFXMVTGQGObGQhw
sLa8td9erEv7ajphuNzHActhH5f1ZkXbs+BFzLBSn+zOnlGjhGx6vr8FLp6las8C
++tfB29QGxW+eo8HcAEzf53i+sG02VMByjtWiwTXB6lOCj2kGyG1BARGN6dEqtqv
38d2v+3GEU+HwnsGjF3jaRIg1ZGDR+fkSkGvyFGovqzrfU86DM8js92SHgLtZuLB
GetTlgUfe9DlAYDQao7M9ClMFGfYitmw9Bm94SZVLognZrpC7kUQJybEaQX7Y7Ql
c8OsBMlK/ByMcsKhakPqJmFj5Bl7MxeBgsgBtaoPwAeL7e21medMwtZ6IBVkLBZo
BIaaODHNS3BP73U7YkfEXTGAbqVzPs35E2ENJLOrohuKkBCjm2MwtgUaLSZxkzW5
3kSbXKwTGIwEs+8VtAWRo5Cn8dZuPSKZt0w9nz9JMX4wDQuwUmqy7hGK3jS3/cy/
HCWXTijJqzWjSZJmReF2qyPnaJzNPoeFyeHr84+XDFzCGiHWKPSoG3zi5qwuG2j3
D139b3VKPnEEUvsBjhG/n5Xjxia25+wRT80khZq6JH7r+scmKPnuOFwwX9WZogb4
tts+UFrxL4QJJMwqSeP7lNmViso0/eJJfDbSzYT1ihQkdi9Mf0N+oMc8s2UJwYs7
vxZyh31a3l/2cTi0rqHiHCdFdYsTU+cA27AcmBuZAe+GuZ4uegVXBf7XwBb/JCCF
jEd8A9619wb4LErcPsTL9nlLPuqWcpqXsx7tLUATHv2lwVuQtaBg+PR4QNov+cdT
bGje6Tc7fCHFrMLyhUGgjUpg64fN1mQ8egaVg1PQIOItYu6HhpgOa+M7PgLybDQB
BVVLuHJ1csvd1p2xFTDjpyms1ITMXIg6Hrjj3QEWBBNQRWxfOaVctSJ9yM/GysX3
2JD56zQ1wHU+ytfhSEl5NV94Tc3TuSNs3Laydq4GzSxKW9QJtXS/xUBRhyyxdaxb
ibqFIjhMY1pDRWAPc7ber+R31l+TI26jMZ0d/EeQKJP//ExvsJAjAAT+V9nK2j+D
NDLiK6frTePOtYHzPCjbUBaFW+wzyKf1epANom8QWnuZhsWYUAKiwM0oUxyKdbqO
DsnmMos8QbGqOk1b4DPFDOy+dbv2IzMvzRbX+sYyEF+wx0bX/2p9BwG6xduJc0nb
AQPBCYFpnSxzzFig7quwOzNBTD0yb9zbxPDrHKCATn0NdHIoqr5jVd+v/qVErZmL
u0OB0z6hFQM5Z8IbUasLyp0E45eKAkXQ/DSrEv8YvNougNx2ZK60tJeNRpH2wSq5
VLKL+JmrQeUbJaCkqH4oHsbsfinwuBl5732N82pynsC1kqXZSFYZ7eE4B17HAt9p
4fUlsZ5bo6ktVoigz9gXwXx3tpIpkQXdrMqQNUsPtDLm2bN8Jq4E3iUYToIRcwVd
pheM5HDF1jTqUyxajLNZTwWfamutdKSGZRNCjdomBfAJUsC5RyYkpdc8eWSJ7on4
keO6Ryhx9wnef9dOQOmI/+GHRV9HQHo7wt6dmN5/RtbI8QFoMIcFr1fC/AWTXYUY
V0+F9m7zpBRE+yPIs8vVkVHDSu8PrKwsgxML60eb1H50uekUH1O+oveGKwwwHDH5
R/MN2uhaGv4u/7HxQsLBlu0+nBlOwppwviIQO9u5Sh/GJ/hYQilYGkiMPzcBSMCg
0H3+RKVyiVtmrAjXKPFbpy3/lVnoP/Lw5vRVD98jEs9IUs4pAqP9PqWubex8i7qK
siO4Z5YsJUALkKKdKjANRLdfeth+5ReZZENMBkL0CLOLogAaqRfFfsOjcB5/wTCR
29qnfCETuMFmrRdFaXEyCWJxEWxjlviTvNjusOWHBPXJKarux6Vj15vj5yqgr3AH
U2xIP2AYnd6Jteozsfe/jM3fecJJs/KOZBuzSti+ReiUFuRSo0kxywxzRzx2yiBB
WKqIZFb6xHBvyqBHTUK7Td6iJ7DUUj9JeTeVLp1/FQpo6e0R7ucwtP1Owtse16j2
6H5Vdgv6KKFERN25ToKFrBqP860BbgvilVi7hS20vCppTTWwN/ZLmWj8JmTpo8bA
DXy7cNpWfBF69N6nBrANj6vfityQIrDS2zdRfNxyhjElp7Y+oMihe/OVAJ8OCgp8
a2trYjYnGt++AsS9pq+E8Eij1D0O2mCTOzq2rk43DxrDV0mipldHuBc17KLH8/Ta
cvdoqyp4dreYSEIm45Y3qcdtXV/dXLDQ3R7BeI1bKEVsmygiDaExrWYnupyNMwBl
s1gonCtkMuEwqN3Ci8+iJdYViW7969WYxGK6bBLQBxRlnWp+zzCiZtTX8MpSlyVN
3E8zHASwAMdT8BFf9S5DeNOFOPVVY9Wrz1AHfK6AvuZCGibKorz8skTiVa6fVlmV
AiHI0j27TsL6h4NlxfP8uGcV362mYyDMOBAhCH3BJKhuC4KG9UTnoTVpfKYFt66o
cOHe8yWZ3KlgNaDwPHGK5gsC4RIE1JM9rDK6WDMr2pktPmdSAH59F4XJNdJAn6/g
SsSCy/BctTYHm9D8r+G+bDFjXm9avF5mCPz6JRD/CkY4L0aDVz3nhn+RTGy4gXjv
ZNse6//Ix7WF/WO3SSUnQGY5l/+7h82zWJpbIjlqZ9tZrDVDT8qDrJUaIrnhTLnv
2Rmi7LdgR7zzkEkJ7QhU4SIqtjl5RwBDVKGxvyQFy9lXRgr7P6QxZWUc/Ds7Ydzl
AqAQMjnO/F6mT7rT6P8cKayxbpncbz8Rx9z2YV+55R3f3Mw285l4yVIDgGh3XZIo
vjLIWugkAKhdfugYEmEA+PhOVQrGatGXvQ/x1znBsTB6WbboPuYMJTknoafsacrk
IBVosYvcllViwuT96I0zWNYsDokwHmpl3ISh2u/ruoSJT4CyQXeGFucFk6STYdIT
26DoSlcq6/skg5j8cVhzF/agUu6060Qs0tugQ+iQ+5drpuxQQKHU2Iwf85bdkoGa
saMYRG8MXDs1EK/h3bR+hiqRSWXi6laCUBQ++lpdT4sHOXusHxM20lqRnVS6BLyn
ruDaVxhH0jxIEhoRevHSg8Gqz6uivbdH98EE2uhEeAAq+6L+RKAxa1mUj7SADyRr
gJTg/rfQxmjvywZAyV1+fiDej2Mo/ur2bxJo52WDnGOCkmNVxyiaXRhH52gAHzJ0
kA4Q8cOlzzxZAg3F7T54xjq6+Kr8BySu3/8/V1sl/SrLLnPuracKHLYGyLuoQJeH
9rXOFaBpATCpBD0gG6mWghBXSh4x7porsbqaN99lKDdPj+768QgqV5uH1IiGEt2L
C672cdVbheK+eNsMfdh/+QCtBPQ0/0HlUrke8IuoAM4IzEAbA49GYg3fsKfBIamA
BeWEfbomc2NdPpnktO83RUmO6stm5mbpgBewuaRSaEGGuGX88Z/D3hD5ZD6ZLNIz
GCyihttKHk212t8I8zDnl0J1Hze17qQAOafH4yrewA6tu04WCtaSZXUuC9dV8m9/
xHNe/dIeNAChfdb3CXDblg/8L0o6jKOWsqDEI9523LxCPR1v4HwSV41DWA3hZgsQ
UXWC3tXEpyK5Tuwtbn5YRT7uZYMinvjpGOjwFRDU5bXDPkje3p4WhNZtsxXr5APr
sguXDkNHphW723pSRaegjUqQbdLIhpxF58iqsM2FtQUbYIBOdTdJz0ZATP4TPUvs
YWBblZ7wZumVB353pUc2mA1Cd+2vKB7UYGhQID9n09akoptOIn+5qu1mN8mWlion
4bWJHvIEo0zSJaEom94tqOor/Ym5ekjYyafc/EeA7pTc53ALg7nrFAoGqS/EYPSz
afEuEVipzn1bUb8q78feaizWKwTzlsPJ7I18ktAFDLvVqd5ebt13zg+WtKhGew3O
OtooFPIaONV0tVFO9vU1j/877E14CV/nClqPLZ1gLk+pTW5oTjdt36WfQ2CDrIaG
NTkCAAX4rXlCCFNhMUGN1rgeYmQEWsXQqEL3IUxJfn2iEmBUxe0Q+EEhLnzEYjWk
VyyBTIOecOqdir+6IFXL1Jj+eZNjnXowU8f6/xulok+HL9a7JhfdJ3bK4f5vQ1B5
SWaAXwKfxPRi9VVf9gL80rHRYYiOhl6Yhb54t2KAJuAdxtmveHSPD/obhbjGeYem
jtBHibnyRCWWHcVcuPS/MrL2KCfauMGOd0JU8tLQYIDCArFFyQTnMZycb6mNWt2c
c+VlyMiebIImFTs0MNDZIWmvNicQjGbOnkDPYjuVpT0PZmm6k2ume+lS22edoEsm
jgyuQ1f9zGwfnSSZYFLUL38oxxb3IjN42BOcpfsGVF7NqmlWLsBzCwTNQLz5lEs7
UUcVzlQHwwiMiwpjtlt3zpTOcF1ZlL08AYc2pSsH0AKkwil5GkWhYHILtZ9xUVS5
dID3bo20g//9p45cifBfx+F7QdtSa9QGEFuMi1xsEZmACUSgaXGFBxoEkUi5t8ur
dHAI5E7JgFjXi9cOnbueqGwpM7RgAmqPA/X2Mfb1HV7grXiIugApH1OkscM8nhSW
GTrc/eKCMRt6gXFXsKtnQKAkEIUvhuxPgfdX0JYsLFndZMffT09HRVHGfHpj0MQK
iiBskBE/LaDKyGuqdOW7d7N8pf9EBRlODoqOemx2v+0dcL7eHM0iNfco83NKKtOS
1jAc8OANAlA/wDFK265kkaddhD5CEXJf5/NgbeHBeIzcAfdddXp+mTqpUiJSbVQf
dZGFPBzLVFMkkTt0Wu9ug7+Sr0gKJ5sdHzZBw4jBD/r1TIEVKUUNZtSyOEWp3108
eUD0UELxXDY6nT+x6nf6jsJsPJ6h9w7Wb8u3Y0lbeLRXuEYb0gojtzeY2k/06Tn+
I7VniBEC1i0M/Bbr7F6CcPjjVxacYcxtKOW2ewz7rI3/+z+vee/zosVnIahBn3Pb
LyCON6BTzamIybkkf5243OkjbYbMOXAwvld2jdRMI1/wa5nYjGPfgNWQbRp3pxn1
aHgi6YXZGWv5coogb7/sg1w2teHsNeTSJI9/DFiiGmDkPj6dWL394bla4tafQDOM
pmzZQRXOMMv+7cj6tgpZEglVpGhGe1AObKKnXcSbagHbmNKQ67bS0qaZ1Sdh2VXQ
3NF9dndnoNUCmFZd9Z6zsg3Nof2RBpBOoP5WyTIDOMoeiSdM8lOPo9gKg+oZBhXs
TSSGSLK3a/RaQfqvpX8m+OIMZFQofHKSC+8ITgDmxaLYSlvGngHAPTgPgD/CGvmU
fHdbeBSuDjJRijxHum1P5q1VaQ5MP8V7k0NSXCb+0G6wLew7KfCdIFRuATjmb71X
sjxJDs1OwPA0DPTz5mI0KAtHYmYX0t+URh16Ri0AT3ex4SFO8zI8zlbkPeYYs1y6
7WQWh4jnTCWeoDRBrT6a4m62aYlp1PspbkUVgjE0MYxQ27po4uEy5Oi8BXsGZAl0
9ZPeakRRY23gNHf6tmHA/bY98yGWdbpAO4iIvinOVzdfr8k0L7bL46CfLqFk8m5N
SYN9fNP2lDqMZkdtDqkQvc7MKORGlyveHl6zB59CLhLr59sZZ66WEd28sXxmQ+Zv
g4j3l4qm+IFn15b6IQT29vmHcGCwBoeApfqJ5H/T9Che4uX8mrWQlKfJ7QFhSNAE
2PZ+t0UjYYSeqGLNwPyGmn408dmNxNEabeZySV5gsd4tJwf7dacN8si9kf69/gEa
vRhRNNfv9YgOTXtda7mdBxUQch4ZY5sv5RQIHopnpwM6x1dsp48iYB1qBKqUmskx
m+kWb5IKfFRJlrd3Fp0gmqKwCRjCLsIgEy10KyHwfA3ipUJpn3cWrdSY7i7RpFIF
8SRAUJUlb8YJ1+mHfa5TEIZIo2rWfe+p6K88IsResDC4huw1sxDE695s/JRYXkba
VLK6f3f7BAyRLnisDcvCKshHRLgGla9NpYL/4k7BsDX+xIIuHhVx6yzuovWY0uXq
gQ3SxEvWyMOlJTMwn/SB3BTuGnj+CFRulauy51hitvt32+W0a6eAhwvZyPgwe5Gn
KJhVuSqBLI5D7Wh/5VL14yjjaMmhiRkNnW0apB3nGutz1KbVyL0Y92O8iBb8oL24
Rw4nnFumI7gm3U1ZM6HIfapHWD04AVDRTOw4ZnKTeLqXLZ/NRQEtAsjpbWjtXyzk
p+DINNZe9UqwR0L2AngR2y1ZdbtrquqmBAXw+P+V5KQBTRyK3m1+XqINZ1ctkboi
Xqn8FHQkRGn78MYx3ACRrvTkEE7yjQ4NbsI7G1yG28u2WH195BXpM9clanOUdAZw
v9ttcVfd5ClEbmkpw4Cztntzq3vXnGJ5ciH2JBwr97w7XhP2rMvMcr17AgvQqj/F
BzPTDR3MwvSfCFPvbXAzrmUHgI5YfdiVkZ/KTkGc4gfKztahX+fzxkpaOOIyC4Z3
XCMV0baGv8AhC5lapjYVXS7EiM8gecsEqfTEgX0/obDq2Z7gUfkP+TOhw1KuJdp+
GUTgURgFIpk3ZEr+wEhCHNtcnwe4rUcrXMGYy+v0NM/26gKXVmzUIBCU7DhFPqZL
Pa8sX51UWY4RpvuknryF1Msz0sEeNEBwlucl1z3YI3jdLIK6VkgNzqbMu8kERyQk
btW/U0ID24LErZXcxfSpNUcUlOrSiQYt/vvNC/8d6JAh1rnrK5Xl49X+pO2j1c3+
u/oi+yxtEvJNDc+eUV+CXsmUtib45mIdCGt1hA4VSuwyxfFmqpO5ke8vrkOaZzDA
aS8yhmbf0t37StUnkZK0MKFchJGjyqUHujvMTVvnlvE5MtsgbI31xyimq+X2HmId
tVzXfVVXEEuMYzsbiT2199mBZaFf+5/TwokPszp3sXw0tm7rNExt2waRAw8UOMRe
74VNDiymTkIgtWkInHGZj+HApiACunmYqBFavkXpsoY8EowLl26/Y10FUCelXNjA
ElZnuAD5HFzwq1xjdHoA2SYruxyoJYwCNoom46nAZ2aBMAwYhd0gGL/l0xQ1TEFu
ajApKrbpY3C8dujpT23TaRvGxssUYbrDUpj/fy48YEKdkp6s+a6TE42gd+DMA1g3
OifwWm1n0fUyi+HeFbrjgCezXrpNuq89p+JxWCnwIJhWLZp5srk79uQA/Li7umz7
YD+PA0AfBMl3Jhhxv1p1FHn380TPWmOE9p8j4lFI7tXvwy6KbyQRv41CgFRw9iNI
NJ9pzwchOX+9lIFjrdTocTG3vGsERZtmlhKcFx+TqiCNBMtyZut9ydIb14LcHQYm
oVaM7sPtA2DVuHgHmaiIXvTehJOyJpAIKqjeOEFjze65b3MajXogU8/qrks2cBj5
Fuk97jnGyGEH98pHOS+0oz0XgNppgUclA7/3hh63jBFVzgjAvDLXyyQsAbArQt05
5wd4CFLcvam33DPba/lJV3x/pnux9KDiCQcLAgACo71oOu1UKGpGlr/cqVvjVCvo
yN4x/R1jQxLu514kuPYIH9QZYVkN5rlhAi/56xgyvxhRcQ15SDaDTetDb5Pte9CZ
rqHKOMpcJcpNLPcdbrQ9RJXl0saEk5mLS6xShDkDhuih4eRPmoetb10BHvW2rVeS
p46pYFAC2FN6UFYkLZcP1xoV5CK9IJI/viuwb1+zFtbYUqIvjEcWmWue1gX3mYB1
RI5w6lJUr+3TL/NAwAcIPQblxRav7R+3KYNGLUpunpdkNrRkXcPWJIwjvKP7+Dbw
LoyuFsD/UmnCImICuXxkn83e520Ojk4mvXaoCYB3abgBmtKuXHIz1+IcdnlHO/14
ug4N3c9Z7uZ2igliGgclbFD0i6defHz6q5jt/3JFpZDdKTf0+nJ9uvVSL8ZTAy/I
kv+G8DfGwHUDWFWMuzTAnWWBKBuC0ZlPcyFHII6oIlJtDIHvuGJmAzy9zkd39oF8
Tc1JVhFlk8SpAEKnHk7Jf0qaILKuZUEkEM6SK6AlMnDiCJOYLLgJkZKcwndajfFY
oIOgxtHEL+vHEbLcpifvIK64JNzp3dKxmtMhryN75vwr/uMB3Jnld1np47IjmVLc
Lnr21ccAV4de0JLsenUABfCwJipsdkYFnbg+SkHtWOXdfj+Dz4QBWQgNlldRT3Q9
SfPwVaJ2jyp+o5zAFiImy9NNXj3QuOO62VuNfy1yZGcM4QlwXU4AqHVusOoPzFEi
yKrs7Nk/OkaqJKNDUI099BhJzFT5W7G5hR2NX9ZGH4/Y/XTE3hLq1P9uTnSWUtiG
+9r4/44C2IvOw+H3xIPHFKXhld1tZtpZOPbFTNN9uaQWDvqBg/aW24ypScrXrpkf
vKARtFdsFM1RMdAL+Wpncs/y7gMs3HVk/9qrvNUH7envaMtZd6CKQzx9OeKIojAp
PBcGbvSsFOXQaLU3SYRaSElxfJr7+0tvmA3hbUJdzdIbeE7Qzto5/bjzwjF/j+vi
5l2sM3ACq15dTZ8dG1VSXuP2M0JzAsw5rIZsmxgQMZI3XYVRIKNqLuCf9rfRXssk
3F0w0Bu/N850ig3FCqRai53bOXWJocX4pSESc9BcvMBE4d7cssms/pqbvrGAQLNO
oM4YeFO0Th14KKgoUxDlg22TiAfcog880rzPdpfaM0IJFbgvmymGcLn+QrU2sbwp
/SlHDggMDcauLUF20f+TMhKvXczKtwGFMhOh2YIttGqb5Wjy8baWrCajKBuqhSLs
8os4HE7CN5crHDKfJKCBKqV9UMmiebm4Qrlh315kFNwesS4beS1gHRMQJ2cU4AJ5
ohnrELeVc1pYzf17jzFbw1d/PTlmzr3GoFGD1lBXvIRxtt4NsmL1hNKYFpdylb80
hz6SBWbOFKs+3EFsOm8Bw6ueq9QkIEYbH/S9aEd/vm5ZbImXDKYKfKFxtAlE35aL
Vjr0i+ICZoO7C8syv/4TbNTYtjv6loPa4EbAHjaodc5/9VVWtqrgGRj2rPluY1IZ
N5bziKOqJs8d2OQAsbQlEaFOrJQABJvDgtzNOEV4f9Itrn6lVjbNgcWnAfjiGDt2
nYZ5bg+qEAvAFTYH2jFl92H+vXZwZUTLpMwo8NUFAc3B7Pb6XkBeD4rHI8E3odvT
3MQELKDnwWUwxZRRWgegHO2l8QL9NbZmPWkZRFp6p9P69a1ZCZMbljp1C2ohH06R
HhAxdL4jKqJdg4azNMO+qOaQwyRmqFEFwdcMgs1A1+HQNQvmA02DbMk4CtRNV8HQ
oe+BknO8WUD7ps3puSc9wSZ2a+8CmGwyFi8CfVN6Xds5P9krVLQyA2Bo7b+YJWai
DCAV6Ow21FATwp/+5btL9eV7B1+LJzWHnEAL/vYVuTXuZ3lG9b/90EGRrfhiXYhn
W1wpDl6dkUQxvIpmBxlVlwFgpzLNx7gSCg3hrstjGOermwrsxpEBl8f+FxticxLH
vDQm71BVRSSIgcKRlTPRkXIRVehBAmWrj4pcwPXNyK5IiNAZG/bpg/ySsPGYDYR4
Fl6IGnQwEp7Cp5QodnAqO5kZu+oY68Pr+dRkIS2dmy7zeID9nsZ9e/SW+00rkjB7
eHgZZt5zbkD3CJZ7sGeaMI9TZbL8TVwmfnFAqfBJdv5uaJ3310yBo6ki7MspxLX0
oQX0D1vsfxvbbiopHVruVV5stwLqtQYGnvVSxVy23LS9j6F7/HQaTYDjWrc5a0XH
Sl46W+1hgAPMi+d/qf4mIyZweinjxZuhOWgvN27+s1Ar+XzkAY9gMvi3n5EixryO
RYgic4zyG9/YpA5D4dSzxOvSP4DTG3NqA3DllMQcQd61AIc6xAPH79Ekk9HuokvS
657lVCV+eOk8PQEr0NZsz6zhoJ7TMuBLKWt9KymDvcnDE4Ef+CqnLSNQ18qi+q0L
R4IlNjZLumz42V/Yq7/C5qtEc9MB+VUegdby0YhdXZI7EycYdcA+50c43KhQf6wl
yG3g7y+oCSVwB58DIqwusyPga0GzRLjY5S2nwn1Ct3D1gCrQCpns9gqyWmJhUnVd
PmtTPdx3Ojcwq179Bk9XCAkEcaoP84T2UbyyU1YGN0kduzGcgWLTO0PYRZ0GmN7s
4Rhe+VIa5ejyvZvbLueO7k+/3yeOV4Cj16yxBAy0N+6S6/ptUJfKddl3dErnLlQQ
rt7P4ORobcTJ/gqLCpT5nUZdJ49BOqmUYaJEswP7YWkl4L7jOKUNNKNytdwIWUGl
qt7WaMR4RBSnhfbA3le1g5dR/9XaR0fks6B2eWTvLqcTdrsMYDjb+TNVcs7kqnfd
l6Ep9kP2RkCrFfXTw0OG/Jr2Ce5rda/Nc65sbpj4p2xqzmt2JhXT6dvoZce6C+ut
vcRNxCzr8vLg16hZNJ41rKfTkm//vJw17eU6AIBTF6KdFdqKBkwdgrootlWJFDwA
tBhRUSWgSjYD9W29x7VAwZrXw77X0IOPRCebYL+hmLhht8nDsmR5QmZi6BjKe37s
yfxC0glm93M81r0eEHlWjCL0+ZZMud6DtATCRWXehlukrnXPar0DspCj8HGVG4Kg
pY+K4ejsg7gzunpqEq8T6vuD05ubi4j7krCmKMnr3vOvmuyE+wZDnH1O+zoL7yGF
gTd+0sDqLiM0AWqAu/mEKFW09DPRwC9isY01rKgUo9XPH7dvg9BB4P93YO6u0Leg
xjUS4fRwItxYuinsDlk7TXl3G57pZtzRqxZ5wzjiXaIfj2RIEqTnUR85f6rzUoyX
GLdlOATi4PvlOEOLIMYIQYL8nN5zwTq754guBVmF89e5vE+Co5q0+xRib/UclsOp
mbie8pwzqsUNfMkPQ0+yVvj/07A6H0T+n3PBQlTuppG5kfrNrRBTsScOPI+jVKnQ
FDPPPgrlCOPqN/so5GBicVnO7wQwZ9Wrqs8JBDBz086N0/0/G+ad8uNLEBPKZl5j
op6GnTeaJqF6ZU6QqXfjPsPj69rCp/FH/m6erppKaJQq5b629KQL5g+XjtS2SBm4
g+2CiNcJhrBIaiGWOdxlotGj06yzrf9KVd8dhpQCbX+OdX5BRLzValmCEBPxWjRD
dplI+EnyZwLYF9N7j5Jqvr3QYwO2dXkbLCs4omHfpV1fEIRKVp0/6SmKqf6Lacc/
Cz28qYfaqWMLbaz0D2vRXGF/H8SuX7L9ZSa8GLeS1W6ATyiKnu4YC4veLHKBSU/2
G0b6d+KLB4PnkYl2iesv1mqH+L5lYB4jSn8a1lEPcxf2zavQPCfRvejKb0mv6frI
JBDL6O+GCdd8B01lo8/bZU9/+hSK0tXRoDXMycvpZCCmL+GNYs4CLJuuUgxa7Lit
p1p+7PPvao7tcciuYAl39kvCat7v7Qd2Awz8d6Iz82Rh3tQqP+tW98ymNbKnOimn
84ld4ca0JDPtvu6U7hf5MGYdHSuthIXeSXYR5Q70Xo1VncKxfifRmr372qFRfL6A
twLZNSg7o8IglQcEfGfgT7/2U0NpZk8r/WYcLu8y3WBTdvZAyhKG9g//5wI7uBTh
JoytjbZcHVCFFFjkkPgFE4JVmCFwaW8oCe1B68k+Vw3d91kSm97E2o1FvgLt2y6q
+4B8K+ddnUUuef+3XFbiatKNfuaNyTAd3s7mcpqU84/jfHY0604SBW8kySy6ADgV
a1DOVveQbMdbzoCEueZiTOIA/IocLhG6mOu5sP40OSwNlNxvF9fUluCR+LoW/PeQ
eu83C1PY2dKErrAImxvw7vGTzQ0J5Qu9zq01/G2Xu9Y9K9RgGVfhF3lXl0N35EMt
uPsogzji7BekEOO5KBeNZGnfjAxXTWYl12Jlg2VfXTgiL+TPmzYmXnxVtNme5O6S
+9nM/hUn11tUE5HO+bVjr6Qz6LDzuewDSZLM7tyj9w34bb+sAW0g5CciLEk1JX/V
jsBlTRZ4DQVvupKiojQhu6vWkVxHzhMhs6UWfZSmunOI9SPGhLuJJ7awyFoT0qTv
m2gPDQEOKDwShVfW1S1OlHmhNZ6/MR2ywuqvprbDwuP4cXhHzv7Om4zVDf5Gjc2j
Q+Da8iL31vk6md+ep5InpShALZp3M+RP1WA8uekj/aZ1W0TH+BMqGz49QLaAjl4J
PuTzgzv79y4TKplTBdM9ihOT0m2dPp7lKlR7DbdikSIRfNz9cZ03hmiCPnYz6Y8m
E5BX7S7z9my8gjhf22R7JrMFLDe1k7EWxbDdiFi7cHW0NHtbuvst/FFzRe8mIdIM
IkVHmcBZTqWQywck5W16IqljkIcgIyE5feoOHXaI8gxBY0cGq9IXNyu+0F87Qd7C
vBgpZYcIUWWyV4Ip/+tHGLGGYqN2Mt5v9ZKK3ZahEgIY+UGJ7eDzKgXMy8u7GFWf
cv8pCF2xzuenG3g9Dy4kLVGZrcfKr3+NPu+8NqvHdWbKc+YB5rvUa+KQuFniShiN
FMqIweoikHCZTIII5eLBWkF+5dKXap2LvQ9BZrpn5sGdvD4wSLT7CiEhdkMl4i+1
xCjU6cYmdCVjRLMm4cwUfPjzhritDxwxxK2vKCDqWT2mHB7IPnjN1WD21jlq7MB5
dQix9c7XnKxmLbHzWbDhIL4N7O4eJg02HuAAZIk4bj4JEOjMHxM7grs+2MledDBM
I1bGAnajCT6vzmT/fk588L1BVD/pcRgIlqm2F/LhMfvdxfnT19BkNgnx4ZtaoHKd
x1LTXD8Z+2KJiqO36PffmOJeDYw/zhiqfVvDTPLaSJD8suxswflkd+SK38jJhd8L
UYYyL9W2GEOm0e8YKQLFnrA3+xAJbH68rRNn1HmJwtLbnDIWlgG19jyqF9mZeImr
MxKCqbO9g2nxi42060c2vUZKfTl0bRY8g/7rWDchIYZDLLsyJi3T9TX86mVA7qNe
iAJSQByG/aYArjnb9MixXEtoVZsZyTKugTJoGhsSlb/KRZhbLkaYPaNIbd8Z5OQc
QIrykQNm3+RHBHTaxeCvIeDcpYSDzmuSiA9rGB7U6eAiyZRreEgKtYtZO9SPUC0m
BULVafwiXJTYnwwy66XCllJIdR+xDLxGhjqmDf/lhPu+L9G0ADe6Rd4iPeyQJG1D
2Bo+HSXgxgJTAmk+jEuFpSwl5VghfNqocrhEjmb6X868McqNk+Aftw1raF5sR47d
uo5+qu+dC5dVhLw9NLoz/wNMdVY0sryXkH4xpfd8CqEnNbtoysJTVS++r/9ce2oV
rInaB3hR1tvnf4mST/iIWXSBq9erUT+kP5QdblT2fTA9qMrpVCegAoeeHL3vFIzl
BmtUAknVcJYqXpgFkY03XRTDIh10h/EEDHAz4nDLRZHy32u+QvmfkLc1YM8YjPWC
X/Oy2JWsw/MTUQ3V16XOwMeonp8JV6WEHcT/B7M6rsIH0VgMrW429Vt5BRPGYlh4
7LcHlUubOAVPf57nHcB0KiI+sKZN9P4L5CKgMT6LE38z3YhY/wRxmUxJJQumDvqF
tax6PSVnxk6u3HqY5ZFIFfQky1XPqEbYHVwNjf7BhCTGgRqznAuoXS/LFM41FuaG
M1E9LMHiAy8FU4X0AFdpk1xiHwnIA5ZjFjQd5BZeEsET8EaluyBxBTPnmf1IT0aP
ZmEjz8V/iXeui0e1vuhkwvijbGt/SiHkfSw9gQnXxI66m05iHkPrlbG3/T8G+oS5
anakuK+hYMuKzS/0+pWIGwCrzXHOHSnu6d5wG2i6ys33ecBGYjOxpuQby3SQuCis
1PVbBwPXFvKnfVz5yaQBuylDLq0GKK/OriU3P7QoYEwE443+7GjINV7f8sPnlwU6
3GDbGf0kUryy2GfWqCamzPqmaA3o73gPDqYpln9BYMKgXYqH5ubhjUhsahk+/66Y
m34JaI36k2L8jdjcig4OI1MIbkyiAeJcgIonnpCEaRffMOwNH4w2IhYjbJ3X94qN
R/vKK2S10MO8BpF+D+ImqcZwHEDY6UZttbAvZJzzqI2IbdKohpnZdHyaVJYq2FXE
Af4WTGSnVL3scPX+nfb09PlvBoAUYxiAFvoTXHnARwz3YENJG1ZIbOBGtO9uUUzR
Tw3aOLzNojmMPF0lNhC6FmbzOBCp5nTPDs1X+x3X+tcj0/i2h3rPpBfbHPYR6+T7
TJ+jQExPK8gVqiSnZd62BuXYMZYrePApyGphExXMkCtR5348RFFnzkSkw42SQWCJ
Jl7LpLFcmcNATpF3NO0FqUo3ymMZvGj3cJEGoqUjxlfFqrRKSj8jT/MIrealxh9z
lpGrXYlOVLBYCDQ2XswpbAlFOThxUbymruwt/tKwi2mo5zQGuuEQe+ZQvs+yOJWO
8NLitFDehLZpaJ7fLRLNksNAlyOM/bC2sPE9yaj42S/Glo2N0S8wt/BIRxTWv9Ru
hVTGyi3aVCse3dQm6X3Nx44jMzY6n2rXLUUf6I+DYNxPX1VippGcUp944SSOhtAo
iUqwx2GQxw1GMwngfE2e7XWLcGAE0GoNQNd/zENbp0oEzURs2NNRb+evqxww/6QL
f8DnZ61VRLu8P54tAvMzDy7A6QI+enQoZRgEeaJeof/qx8+XdsjMLVE3EkcTfZEW
e/5zWBzAhADAXUKOFhRl+4fpVcNsltXkjRiuiSFKj8HXpYwUJsu3gBIhJVE+1JIh
KonPGCgw+F5bcWrGMXGwPpkCuGFwhZNNPlrQ64eZOY2zDFGnOzilHISSK8srGkZz
SvxNdkzNiC1FsXfC2IyxhF0m8A9KGchXnZ6iG/C9ocpD53TMIO2B4ftZ1IQ0+BXp
ozEXZ2TZr1p9Y2disj7nmb9lRfkGrHzoj+PC7htyczsgPSU8iVoKwPUUQPKpHDsL
AePgTyZcwpNf4AVAAfV/FFNMupJahSj/tPksE/aT3kzpqc6ugDnVVfKCGp0/QZMn
0BmSnU62p5UHDvHsEnwBs8Txeoy07Ot74nHC8I2+pzjUq5KiONc6W+UsQpAojzq7
w7F+AetHkGoRGWfDFrZ/qvcfuHkrHbtSwIXsZ6m5q6rO8A+ykZ0XFG2n7mB9YNuj
EqvUCbgC15JUhzfeJ16Fm0NRT+DqDVnp7n1dhGFgfmOmequJB8rudJS1kBKcxeFG
h2o7w9WZJ58Gui41njuZFrjpp+boByQK+hMEz5BhZqH88FbxZgeKwFTBWIPQwdPn
zKAfrkRX5qGNp/Aw1klDG6Q5liSHm6L1IYRmnclBsOjd3soBl8xywM6lBn1mo8vY
mATj8nKTOhLDYFpxnPUveeXkwVLSGNiYH+6UxtwEaLhpodIeUAvZImgLRB2pWzQg
h8+EBgLMDDrxz0tZNxyn2psezAuEvW+DPAOjeexshsxy/xEvHFuAu6sQZSP0jqyX
6ax4TzDo2Ov/J0yPnDNaJFO+zPQvkLl35tSNJdaVew6ZMe5vfGYAmwh+H+SA26Qt
fWZWFbxkQoBL9HW1xHOc8CtSMInq/jyjrhOgtI6J6LX6PtN/dzKHfGSbakmxtkma
JYOfNZBwWY79MfNBEeue64FTqpac0njbtBU0JsA6Z0/by9vfPV3CT2qtFWtajSIY
mR1nbWpGl9MgAbqAegKlvpL59DRZbDUVg68Mg3w+lY7FQEyvWw+Z6A01nTJSZyMh
iD81Pb0bkOgjLqCWNrH3ifSKIuKzDvhPLA+zH/wWbjofRThPUKBzDTwocwv5VPBx
qtJwAqRJPbJ8HYrz6kG9vG2ViKegmUKRzZXSbNz6sYArOFPJCJrjvSlG+ye5DQmG
QoEcvJ4nrKjmAslwiJ04DIu4IppE+1nzBJd6Fx1PHP93UmMuepxvXnTcHuyMiOaR
aIbUp629y/WsggqRYzr3guX1978SVEGDNyO90V8btn+a3NA3dqP73e6M6/NkaH0F
eQ0hcv1Yl68UoNZiGBVaS21FLyY4f92c1+o90RdFOGj4BOg0xBdQV8wkxByqCWlQ
84T05m9dBcyZTZEjjk+e4V9BJEJ9suaDAWbOyRaTh1IamXMbeRKKXTzIVgCAD8Vs
2ZHvOnAJ2J2g6s+TnOlBfUyNy/7Qu0x0SgGwYYV8fKjeo+Ik90ggTGOFzlDCS57b
LNLUhssz1e4iXaXVO2bRHoHTeFaQO7cSCfqBR49nWuylo0UAd0Lcv1iRCkVC14Fy
7ovYtvJ4cvz0Mosrq9FmNRlPTrq+wu0Dv+CSsr+2ReBOfuXu3pnkB8hAfHeymog6
AYZHRHBpo2Tf9RlRmBPFwmR6JsOewQXd8sb0zbeokrhaxaI0Lh/upR3M/wAbbHON
oc9sf+7VfN0mPHggtUrXBMjB6jfqr+0KUYHnBmWIt7giwcClp9swCYP0FUwcQkzX
Sg+M0/0jD7ZrlxGR2z749J6DHPGwgmNczYU/L1xPuUCBi+FLqZMEUkdDsiMPaC82
9Us3dGdzMygIyf8wfs7WqI4p7CtOX/GGokw7Lrxe4DuqVxD53Vv5LV590PYjUTU0
VmqJ2cm+PDCMuV7f3S5CWxnRvqNAzjnta4iDgJCjWjnKCvG2N50fWelDDBl7Nwod
Jau7S1Av/GmWEw7BnEQxdvHTYgyU5qerIU7UDje4QgS9uuavkTRHZ8o+xwesMH6f
UNtI5krgNoLMEzvjCpUPv+uul6HYVhtSMjbBeJpjaDuukwvbdCkQmnpL0fuJlrZU
JYu+BCzuCShDQPF/+ll+dmkYj6cNrH6T0MZsX89mp6s5dFIkOaJ5nJeUwZhZOCyl
AKMZM114wLXpJponWQ70+NqD948s3Ys43rDMnJzMhV5gvM4Q3WlEqlcRKQSsBM/t
tiIkthiVC61x28hzCXaC0ZbHxUyZGVDeitFIuD1NqMHp0aIHAftU/AFOgg/Eufad
UdYJpVuuOJnDObBXjPgi6Ql9JLZALHABUk9iQWoS1zt3aQok1pGWRtXrOspYU2DD
C5vlmytBw3HWhAh+lZWKjHJ5m5GDkQDc59JnqscWLtf8UvnW6j0XqOtCtuQt0+ld
uxO8lEcskZTrNSCUutZLwhX6PI5KcYSHYrB0gOwoIRcBvcpKn+92VbO2XX2AyV5E
JH5zFUPSpt/Xg+klQPxTu0LgXXHOopf4OX9LpRV6spqY4h3pNLp8/n6jJpL7ROVk
W0LbmN4MwpGLxea0w3+Bld11NYktukuN4zCIcc3Br5HHdQ0T6vkwe/r6R/myEObZ
+uNsEfkQM6HEiRlfyxxNivGLLKQiNnphvkEktkty14CKy2Egpo2vhqEl/iT5wF5E
YTbnSVr9BDS1KOtfgLWKxBUSCMfsegWxE+rnfd3Mtq1T/LyHAkysbx8ubOd16ICb
xZHTlaYNZLrG8M7/hYfzfFQ43usONw8HWroCMFF2f71lO4gffoQ8eyuvKFk/u7Re
0ijcr4lUdqAvGzblk7lBYIkYTUcutMRtKR2OdmBWVuQ44UZ78SXy4Qd/QuMZdO25
7inLUjL3vpi7lbKqlN7WXq+1Bb2rWxn9gP6JCw6C+PcAxZQIE3fpuvm3Z5mhfTGF
CGYjPNoebiHiVbDloaFEcnwk+CfFrmSX7mN8WlNrESsPLy2tcEeu5+fTk/l1jTGz
TxzMBNS/jcuOl8fXYrS/SqfawPRktWuf48HjqSyaAsaefM1JdXjv4pMvZLugYaTS
B1f/mzJ+POVwoDSocH0nsJ4XswKMoR2FKV4AGasboqM4A607VncJETbkYDkFiyoI
mydn4crTlND4UFe+1iFLdE3GQ4z2vPZeaY4IkwD9HrUmfsujoBL7IO7AHlfjggVU
bXO8yihJwIQy7spEq0185FnJn3YNJmSbYn3WVnUCY+wPFXV/PP1g6AXh92hE4/M5
2FeRYzb20jKcqypEGhzkgVBfgC3MWjvc0M08IfR+XjLqUSjJRITOYX4xPkhFm57I
77DT1DhfPyxMp1y75JBu0pbUzU6b8i0yDWEorZbvhSungeasROy755foILs7SykH
2eK0rMmJDEq+hAxMk08YzKzYz+KoWD52VwLGQm37Xl0cZsETW+ixvFRYZvGaUd2v
viQzs/UX0fsiComt4bOmtnb5q2S9h6aMYQexi4g7ERdnKCMU3AOiLKLIupdI8idj
TIFrCbrbQkpzOYHvKrQaumOkdbHN8iEMXRHgPWzo//RECMoAHMs3Vi9Ng5Dxlopw
TDpFOY0P/nmF01Bn9ppROjRA7S4UTrs+yPWa5/0m+3MNRgNWXG6Gix5OGH7o193C
tpz6AwLOMMUXPfpusv8rqkdA6UBpDsSQvt8DbvGb4zOP8nti+mq7weufkKQW6X3p
lr1BEJjtbn589RMEYNbCtAF8u7sV5g5z4W87g22rAOPEVMyRiQk0iSnbXLrNgA1j
tplritP6qZjCT3VO3p0J70UPz0zR3WbrZAzM1OjwnMakSOI1YhTbHwRSENxEr6dX
I9CgdtgiFl5api0DA38bsFAqwi3gpluy2N1BH9kkrOPFODMXhtAzF9GUjDT31F5z
Ns8m1kKUYXaGVIuuaFiJtt/iYfRDkJQYizW56SGa0bXfk2511hpP1cQ971qMbyM7
8EPwmJZs6KH4B9WRaKJMaW6LB7hfZQ6EQZw7SSNNr6DVy9OQc0FoakhofScAVGvW
5tPIqmyLoJYdUAqRm2ZOE9L/U4h34YUiA/PEMwTkmsnlImDw49/q0ulSCQuUJUS/
ZOT2UMRss4mfNoQs88AIoFAuTn3/JTE4SYhvMJ8FWVjlZkXwLZUy3TwqNZf40Nc7
s2Ops82q8JZkSsHzJ01DgT+qrAC1+Ya+jQwzqVRxFtVGejV316rQxrOZCF+8tKgZ
WPEG0zyufRX7vHhmJ3Yd5QRwEG05XxDwPd2u3JYcwJc/5Vo5X1SMKlpUxSGgyoP8
HdoH04tTbb2wmf9DfFCjykoq9reu+m5YaP2dawfr8gSKrgs+tWsZaSn9tKBidCP2
Y3x6dGbrcUWFSR8/yxKRTDKIqzEDPqIRX4c7cVKfdm+BepAfg0TGvdRMzExTCXK2
MUgmAk3BO9os8dmhdPutnYoN+g3Wv4Ws9IELjV0mkCMZohpkRMK6XpbbXZ01l1kr
DUxHptfLHM8ALiMCAfzrXeR7UoAqR4D7+YXyeEd1FVfrZyC3N2JTOKuKdAF8Tdlk
/rRMl4K2QQ6xo49x5WVPaqDgxmQ72VqZsCVgzJtImJVLZ8Xfx6K3oW5mfH67SEHp
TAl7SJaDs/OcW05a4ImtuePjlc5KP2ace6uWOhYhKWCSmvWumRbsEnsLpG2UbVI0
ocV8Sikp4geaULYGtYnCPpZjL0hIDE5TnKNu5fjCTPsK3B+rHZRmujPB3zzuGyeW
LzV6GMDYv/k2+YqBaVxKNqzZHU0U+Ksb9ihNhsZuVpFpLgloq/ZAQfDzsvKmbPwR
dFciHX8lQlla63+yzzn3tUiye5eott+JuJ55Q42kOfUdxohXk63xGWbIXkTGM0i3
tbl2xKXDnoMAIVWueqqYRmqgoz787BuvNg/eNi2gTGSSzmJBOiVU5HiKoHlu6EpL
QqMMNS28m/+y0D3UVzjfOLZ4yorW8JjYaXhNlpRifpg/tyKIdQH+TdWXAK+P5Qj2
yAEu/cG+w/dZwKkfaSCmAgSGkgcdzCZjDVFlpvODED/yPCFkcru03O5odml2I+lZ
KpRk29ZTQBD6budL8qJR2qnVPcAEqXAXz2lde4JOxJnZlfjVC/+mEo8Z8V3DK16L
32fKcvJyN6XU7m9daCHL4W9ERqsgYefsBz+J47jYQClcudLM/f1Z6VQz7ySPaxXe
PBebAuWsmiDoVHP2+4lSRCW/tX+Su2bhc5x1gQZjOmkPNwSyncfPHkqBK3IxetGU
uRrzmP50fxAwYacSsNgoFaQrIaKBcBwSzYR6trq9K26cCqm4xeipVsJ5DLuUeXsf
fNbw5wixI6FjieNSkcVTl2lYY5y4zZ2q6kX4dFTpvImpZG/9LP8mAA1tLOpbnYJ1
7u8FMZx8HPoftw/p206RRhEHsD7CXicdnfkhm9YQBxnXEP3GYGSgnny74seo1nNI
sMCRpTxXOGsFQALv3RwlPgOjcDXsW5PJo5bcV1q3Kc64fzEy05nOzc9NxlBdwMAZ
dJe9TQihEq6hUmPrVhrjrJHL4+1TTRn2t1hMIzIFyPIFdwxg7t7rMB8J7fsPhlUo
GMfl+KZN81JUlMHG4ADHK7uuK+tt9Hwy/O+Af48WmrtXeaWbesq43BD/eN1WG8vS
gJ4OqvvQISV/FtTSKzZA6mPlUxb/1hbZnGAn8eA11ZNvcJpR71jT5C+bgaBbnl4d
ldSRIxG21oH4raOoUf9B9k8i5Gq3TtfIKsuFRiedxpKdaR3ifw45VGL9idLBvmBo
yrmUQT829RBrVCVvPw4JdmO5Nm4stUeQjOPcULq3SaqhjuLENBb5rWuP7kcr3Saw
8011OYAdLLY3VOlRuUwLTSLYa2iyvNCDTug6TBdjXGAzdcKYyyx6N8+BF6Q9ZGfy
ZfKkEkotjBd0RMS9kVzMoXD89x/q37OAY1OqQXN+x+9reFDrbeTN84NoZaqnbvPu
2m3ZHs9r4VeA3FyBD623+Ex3W6giYAd45EiRZ5oqIi8Vxc8msxyXsiv/9UbtwHzg
4XQODpr3ddpXXWM1ADRXY27yDk+PCNBhCAChAVkLrdI13gMW3a5hZ3FGZshMuMws
3ZBD5rJpTh8QVGAUim6QJ7x0jJNG0K5jNAN7IQky0LlS2G2kR35ruY/3vH1+Opy3
7Iolf95F9UpN0x1F9X+Uv18uPYVg373Pqe0rV/EHxafml07zS056r/oslcTMaKdq
NBPcmZYOE3sK5EejDRpk6oEQIY5NCnxUEDSTRgfi5CiQkg5YpANxH+uxgNBFeFcM
QCDEPu9r2ww7JBmOoBoQMmVcQmz2iaQtc9Ju8X8/ZRGoEk5OPb3ORwiSdpgkYULp
c2PXKC0Oh1Nc3kemPB5KaJAVA+iRA0098Dj/7Th8bQpAEjra+7cCVL5uWYSbord8
/oePPs0GrB+wyEmahJe8d3QiIB51GPWrLuIV/jerh0orxduyz0ymPJ7QgUIe5s2/
0AEFI7+iUzOoYxuT+mxy2zgh8im5qKb7Mh2aophWH+CFy4tFiX5HL+OKrkh7Yb02
n238hj/HOSsEoH3evcoN7IZQdO70mjMA9NFVXsdpy4+rVSSqwFZm9Qe+Slnl7YmL
C8zMu1a1gdrsBUetCvj156/TZPoei44zugcsbbBQcna9QWgJgqhMVdX0llvO2CIY
p4nECqyAHI9szj5ZBncNUb6ss66X0ISH+Exn7CoulEqAaxk7IvUi3jF+uzj2RvAA
zKa80oOSZ98yi80Wmcfo52DyVU9jD6v6nE1J1HmrzZKc0lFVj8zWJv4xUNrL+KwM
/XH0DB+ISogN2sJHpB3SjM8v8T1smz7kKXZh4w9L7C+0FORnCWW625MBe39YaS0N
HS92A1FTcocMT2uILG2A7NZJQtXaZIKHNxqI8RJ4lDABPXKGOzyBTHpua09EL/xQ
JqFI7Gc3qcmIsHxnuoRjii5X9NCRLU1ZPaOkWA/0GBFySeIEFP5Q4sttrfFTjVRF
gWC/fhU4Oc0EDkxyI5s+QADoF/XUVZ76RidddpHPCojLkV8Hggk6e6pjJUdEr4cy
4Jw0JwDR5y0A5YOqfaaDM1i42V0oLjyYDEfWO3xvaTcQtpL4567aN1Qvr71n1ETU
XuG1+vXgXS65UH+fvtRW+0mUhBUNJDO+UxSmwo3Equ2XJpm7ozq8ibRaMxgdYyFe
iEiVrG6nyEY7N65Tr8n4HKc4rR9x0o7/WcA9Vr2/VLOmEsrJAeQ0kCqr6U/D2Ics
jZTZi6ZdvGUVc5KgiU4eUHinQTE7ezcdxy0mlskmlRM6jmBNhMZPwLOFCodLwQqY
Wgw9j0WWbLqGbzs0bM1zDLqEZqi7YNfFAO6RstihsUmdVGUYWTn7UNjSprg2DgEb
ytUR8f8mGjisXZjGr2zVmK9avbrfwJ9vHN0OS1HOu9wx/i2II3Oz5pqlbtUblvT2
ZhehsJ12+h3hYYrxVSPYuxH0aUuPP4L9W4hLhByBbJ2vXgqh5JGZr+x4cq2JCNXh
xSur409aq+g8vre1sMHSx+2S5FOjX583dCByPMqvCb6hvEKJSHAUeqRmiHmhyJZc
CZhpF8dhMc8+4x5rmIhxV9tY1WkM/9rCf4BM2d2kIExf7K8lT3J1vAlUnWgarxRt
zRIxKXhP/HEp3KPQ48YueuMxgt0trf8p40jg5pcNMxAYPruCHvV1lh6+EF+D1vB1
Lj5BGxLz8RxD1389eS25fG1hVCYq5Ydx5A9D3Qu8ckepu5hCAD7FCCb20UPE1DSl
XYjjNDkNVfdrs6fm4Cy+73XBLWrfzWuSSmvM4r/HSg+9o9OZTgHpANwzdLI1z8Wd
lc62fkVx1o41tB6CBtAj/Xtig42FZFedVMkot3S6i+jXmxiRL7Cxf36kknk9jAf2
r7GQ/4AUn1H/E64XP3p87IppLX6jQddewWYpdX7ApV/+oyRBtBPVj4lERrwreJlw
ucHp24z4QNClh/QTxpcuhKoY1wos1okiigFRMCqo8/uWewZSvO+vEOLu3/DiG5zb
24EBGGffySHxewLrvnHt9KAbM9wW4rG8YTXn7OuH2+yemdfU3PCx6oInOBzHjNEX
ie5xCiNos5lmsErQ7LqkREqlri08rX43iZqm/gmvAVGvj7TSy+oTQ9vQ2JHnKuF6
/uTaMyTZkvp99lFgDDUnILujVWtzbCbTueSPPPlOSCcC63FRRu2WgeQePCw1kQn0
rCw6XLpPCPbwmvyxFIVK4K6jr9M9oxXSAyoe06NV+jTRRWm+bKlZMq1Fbyph1tRp
fgr5yt9K9X+zQ1SZadxphAHLubNYf3UqwVSUVHp+HliXDfKAm4DcZ7uoesSEqACZ
CdGcfnopNLpy+Yt2Xj6uf7RSIsnskJojbaCTcGhgWiPxoU+anPzmLUreZ2A09Lmo
gjP9+/wL80SkxrJFEDU3BGAOXfhw3MwLMxr2F+poyRKEzfzuS9FN1P6Nbwwkjqln
9pvuQ0O6VbGCbCw0Bfg+jwu3HXQffGyOekbJKyiwUej2KlabFUUEWHu5y7rGRgpW
bcKQeB4/a3I9xr93e3bME7bzhKLaI9Eh0gJv9YqMLtWISYWPrkQYkoz2lEQ0TyIy
oSHS5yVKk8CkdWmD6Yv3JBwkPmtmPydzL9bOybC1Dqx8ErBVSTeQALD2udoQckI1
kWMszyv+ZvD75EA2G1fDfAcEWZOARkuit2mt+Jv4zeSmj3zu/0mXHYoAGvF7EvAt
Xkjr1xqFj5Aq0O/NAWFmrsIWwXaWQPF8/T4DjAX3KRodemwhDqbz/stYJPJWdkj2
Vtlt1sP17/KDacuUrfyk6Nl/PBQe7cTANe+UgYHN1Tr967SGwVHiJISGRVnFWXR1
zQuk6WD0sIgk4Qy026lIS1OQ87AwGjRaOSUSDEFUXTi7qTDFa3tIf4idhdwsmbqo
noX5DmWr/tjnoNaPEjIhS5n4bmRG0p/MKmb0LMs7P0sK5N5WQhVfdnAK1SNx4Fow
Y3rWsAuCV9zTPnY464QR6PMnPcZ1oJZL3Uzwbugs8lzJVCDpGagPOZgvBWAtg7Ay
slwliYO/dW0aonBaZm1IWhCLLd1VMWuQJlC89D/kBWmhq5u6fvnqtHfXOP7JBOyx
oAnj2Yz3mJD+ilkwD3sGW6o2nyWBwdEYDlTUnasPwj+8jDLae0x4wc1QShu7RsAs
YS9fU63sTDhTLsj7qBChh/n1xoxCD53qemNXgVXFrRsEnv4hbx8GSM1fGRCbhlj6
UmKjTzi3QUwVHtae1qVHETzkSyh0zb7zTRose7lvl4UiUDo2BMNEUs8AeoirNd3m
mzfc29r/IJz0mAEf8wH2KZHpyv6K+qo7FP7EQE3N5QHK6Mx0cF8E5QsmiHEqo9G1
3YZPe6G1f+yPMCANkTodOUIcAMS1H7ljX+i2xevw42jkN2Ob34XIzcvdTckzcARC
Xy7ZuF28dejZEzrPG2QYdCSEO5s+5KdxBRWmqWwt+6aF8zm3aOglmPf/Lf+ipoFn
6k5YTioGj/pGnTprHrbMXEHRcElqQEdGjrS70MWhJp5FwofgqabPEzYxfzRXXMyY
Ezwvx88chj7+c8NXkufX9ZsDpFJJUU4HJ0y1GAgD8kN93rRtKtJ+vtDCn1ZWMTRE
il0Q6kbxUvZvZaDRr9eMMMT+gY+OHzQuLqg33YbENhBrUCwArT2WAlIIF7zpScQ6
A7aiZBXIgEDsbTrQFtUfrkGBXmQ4frZzwfDj4W+wQZfRP1xrsTAuBn/en5m12IMN
d8Hku9XE6JEnALZzAPTQf8ZKCRghFgEP3alGsOLn/MhdfERkMCEFvlrh3mdpYOY0
B7TBqDHNX8D/3dneSQ8DufLvvQ6g8FoHCwqbTwlvsgfNosnhaURPnlVA3SaUNlO7
gYp4MARPJhgC0NDozUODhcITmyXnLx8rFN6QZP4UXfwLfoaKLhIiI+3XPP+nqQn4
yNnWvRtHe+yHWTNIjGDHRbjMAl7wF0druXWD7mdN4n9LrWCarX+R93RvOicwF3ec
k+p8+ni3G/ZDDG/4gGdpy9b4CAX3nxZT5iE9gZGvbhnuiSCZQL3QEGSjiiSpwM+h
ZREuD9VZjNTDUCv16udMJSGj5NqmkA1MP31RQ9k+l4PJ6yWEAYQ/swcY00b4E14e
2Ye2bp+n7h/jH8Q5UkX5qvTt6tvbdNi0fzkD8uwwCLYi6nt9D2eCzJ7LmmL8ONGO
bCoWxh41XwMZvZ5qbNmy0FUfKX4cY13hNhFtcL4UoGjbZJQNGGdcb95zmUkodCkX
fpexD204QG3Vh5dlWco+brdxcLTpucmzCxRxn6qhajj+juxLjxGoWCnb4XW9WM0w
/QAMuGC1P5T7tEljRc5V+ZpOe1GjVmQz+6IPVG8oaU4oLjqCd2d8AtshSlx84F4U
4ZSJiCRnN0fp1pZ4roHYa/dlrAUSM8qySOwXHH8N5UtdVcmUEDsXuuipPlhbPprN
phBwjfjkBUX/Dgot/5pWe/xK52kyOrZm7cFZ4ZqjlZpApyE5tsTQDY/0RyWtT4Ma
qvp5QrvywV+CFHbyuBOiBNi2PHSStMmtxtifZDM2mbOWxIgTpIHc40dsRphyt6G1
NZi3WyY7uKClRiifetywzRx/6tBv5DxxaUtt/H6leONm/aH9e8be6VvVCdxI3rOk
68zbyO0NMxzH6qKN0dSBe7asw1S7h63kUmJjWZ209998yNB6c2+zOlGdFdFCrPMb
JVsmJiYlYp7YFRbNQSTG0rE4rzVOR+LWyHLQS149aguMBl/AZeMwmz6zJ8Se/bGA
EzKALK78FdP+/MOpKOiWssauKrosgQCFknpbBwXSKXg800SJlqrxOsgqDb1i9WfZ
6yrNZxtbLiTu1vSrwoOAMizK0NRr6ipvxWFOCTKw+peI0MEec2+yQy2INVWxZZmZ
VgpLmNhyNIEgZcPcCv6kd5RbF3e9GwawAzwFf+CxaoeC9hh9pFcMOHqYbZQxiCa3
nTsGkmGXLgsz2BFNMawoR3DLq4eW9i9umk4qU0c5Od2WfZB0wnafHs3W0RaG+Vil
OLGiNXtY9HpAIgiHADpNfIyLaIG+cnfMt8sbQW49ljFLn+qGYHUGyW7hcegSxrib
hjtHU1s1OUWzvlqOALQ03wgFt17R7HwEQ6WC7ZDslkMA+X7H5HN4ycm7ay4Z1w2I
kzPQSwfACdUVomRGh8B0WMwYBTtdBx/Y/VJyr82Mi/a1opgAo6L+AfJKG8M/Bgo7
w+rzndLaNEsdyhC94egctFl/mcYB5AnTgeBdZvM5LN+Kgxi5CfFwUI5DsDmXcgCU
AGIgwCj1+XE4ocuOqrLF65qcOdUtXllCC3Xx7PLN6kK9kYW5OgwR174Xw7iKfru2
i5dxIbpaejF9ikVHWK2t27OuQ5bI0/Bm4ITJ18Kd4ncCt/0ssNmv28zFeJ0omd0Y
Buun01Zj3toFyOKWeRxROAdLVMbPDrTJGSLFiZ8O4Ufn5867m27AQRE55MgOwmPt
sUILoKQh8Lq1bYjLrNe6zvx8sUlbiS3i1epXV1pbVGlAQEoaeOtHd3EAxuDdTIdx
73LooyUon8vsmOfxDWqXTaNvw0OmffDEhTVLjdTadbwCHN2TRarD243moAfCnrRk
eDA0Ehh1dwATFBX9hO+bZXeWiILa2p3j2WtZyVIr9hg/J7OuPKen3wlHCZ20eUn5
sjvxeuaECWX0QF2bPiUrE9GAXI6DPKdhHgZgPYUi7ViIQmh1LJ/4Uu6E0LiPWj7r
SwiAWKDQdPp4IUlsXFbhp4fZ3KOVcQ9/ZRFF1Dkr4sRHUV4RykhJzyW+7UHv7mV4
h3xNEjgkKyGnP4LeqSOv0RSIF+QI4+DLPS09V8L5mthoVGq6/XeStrM+wIa91Hd5
1+toMiuqo72JdaSvBuEYN0DAz63aSK1WrzI0hqc9JkqTDMtvojD6qfxPnzdrG1JX
ZOga7plp2BcUoapQVd3x5/UDmcaDM04lKtF4UKSPwbHAeTF9mu7K67cVkFjRa41S
LPn5prfxTXrGxZ66aedwNokDLj76QSb7uXfsuBXVwrwxQdH25Pzrwj1E3mMwR+CB
kyaKU+Rqv1QwO4A9qdIf/3rGnFxm7bKmccpFi9aubnkmblIx9uIo232sovHlsTIT
Go9IFOJ6gsCjQp/tawwJYMuHhWkS37UXzcdHQ8BZZO2wuSHzQVYm+a6ii20sLAWj
KoZ8Z7dKvR8Z2J+I9ics50Ma+9bxxO7o7VBs1P9puqygaA5zF+pocXh+v9jupk/D
iUais0wRJm75efxrQ6N8vKKY8Qfp8aiv+eL7ODg5wPWvcvmuqA+Epk5LBOMMAiD5
9xie0PYgbCoE8FLgHoYPL9d0cUoTGJcHmzXu+mQOqfd7m5yBNL2y9GU9wjq69euV
LSkJt+iYj5v7y4M4V7/PtpvYS8zKZXt8sOZVxToZvo1jXtD2fjRYAcWwIItksWTN
gFYS72lUfIZLk9ATxitTY36bSxVfctupgRdYKx3UtZBvrJE7LYh/Qyt7+aGBYWZZ
dVL52YhekusmKNqgTyArRwgj0gON0SaxNRKa54zXB3FNY01HqTV35OJCtllfzuYy
IHPm/AIlZ6jNPfXHkqJJzw9KupDJ+5ENZxxzft5kP6WrqxOZdlgmS/ykiTCQeY8B
TsSUzlaXnQksJPcNShVM+B383vzJEO5GB+s+GgYKs8R2ogvhXtvvMQaOInxSNuld
9jrew/xNGm3xQhpNdVgg6e7ZIt0zjVJywSd2xgzKefaYFF8/Bj1fuMrsvSs7AoxN
PuT05WJ12u75By8Y8mctD6dv2BrYFXxX2t5NxQAPMvlJOa602RBcUfwI4brNibfA
+DNby8lmAgwXyQCV3FDRpGfwCJXMMXFRGypVyyvtbDXK4EJqhbd8ZJL/jY5rz18p
22QYVwJ9+EbtZPDmWSZQwFz22Y5TY6Nfx1SU7XDbgDK+espu5Gj9h+t+DbGvjz7o
+HQomNgwfCQ12E4J/p2po4RdAEIQ/TjMu1Y3cTe/1my4Rt8Qzbt41hCSC7/2Kim/
YZ7X9yr4GU1YiizSXdPF6PQg0WHD8qmwuzXW7sUEa+DQJEB+7Kr+W08BnNRysV8y
yw1MPB7AS7795p0IlC3n3rTZPIHHwGMdN01XRKsptdtc4GUUB5pJdnJq8iEzNomi
CzWyWfyJhAFUfPzxb5LereVNMb6j8yFbFfiKP6IVpwtUwjWR83+mPIGSe5bckklU
bGbaAPJq1wdT87KonjyNOT7CW9TCjGKFYxzrodLjg1zsFoMXDRRdU1hDqkn4ZfqL
uXQWwz8WDFbSH53iworoJUCvnGINiv0mPGtI8vigBCDhZ82GvniJOBRZ/I49Te+v
0CYa02++xibds31cJi2vANBpuQ+rfgF+Jancf5R14Cn1STKKM9u48UJ+ut6EroBu
VH0QlbTSm9ZWmeQhKHNY1PVJrbPtnaAnwegTi8RATG5wwkcFd30ozD7HHUNOUtnc
Feu1HUqUPTNmcySluiivmoO23UAORZEyqUceadAKH+VXsck//RHyR7REABYfrxdv
HH9PVhNa+DalWNjUgB22yoilmcQQB8jy1b9GwEwxOsTj3LDTLYzrGAo8tmhVQIBD
du2PxyA+Uh9VgzqPV9q8mVP2jHxp+YsvX8NzLsjAGhOGJBU2xSLn3+lie2mzzPCx
7ZrI+TfTzBypyiTOZl6L120974kXq/bYBxRKq9dZTfwCBUDd7FvhYSnpApnr5nz/
99A/SCFCchJonPiXeGRhEWJ3CcNOWKmloqkz2KxgJ/jFaCX1BvfwOVzFmbv3Aihc
Z8awrIe+lq2EzYXhoi9R6hSOFV+XqFG36j7ZQmaW0+dtAXKfKolhtj56zvwhMmDQ
vkqhNjyJD0iT9vBKLp8raHtOa5sFiXNP2JNgjJyAv/MhVlqZIVVaBuBkv8+J71Oq
p/1VAX7pU7ls7+9P9OA1PIWgsPr8Xi5aKMj1cl0vkhLhsIVfLWOI64+XSjdkbz0c
1PoYJp57vKWeam4XuIi+QYPUaf2Kt6GDkZwVOlKMmeFwOpDRly7smXxBd0VojakG
dh845riB7qsoYNkK+RxbgLGoeZ03CVaQUTv5E8G8WGGhoN0eyOfkkzME0sUEpQmS
x+Dy7fCaeX+Sin8JSkhUBp5d6IrSpzIJeEuAUu5hUGNMlTCsG97sjssb8Q6P+QTI
YaNiIoULghevFpBbm+2a8LsJPFhVI0ur9Zv3CJ3PTt6/MVQt6DHJM73faLDKx0hn
modMAUjE5ZlSnPVuZiY2+RYMS+KdELEYp3IoJQxsNcaEvn1ZU4AyIMoR5HeZwCBH
iNOTNJQgbw8II6lGwY09TiAIYiWwac4jsi8hm+jmggM1vZqIkVshjFEmD3FwhlV0
auXeHwZrVZTrePbJA0DyXIQvhOVApeYx5eL+p5bk40pVfFi67DysJOzWlJ6iC6RA
XMZeTNKN39bQz/X1VVt2gskNd+N/Xx8p9ol6kmpxo1K62XWI6qw9KLy7003KNsRa
zZNSCjLT5s/NrAxNKo2LMz6mqCFcMaCUxsw8RoNKLzR9esPAh66oHzYNPXfT7WZi
5mmCAcvWfjFwPlJ0qXxxbslpSryMdkv6Oa5B8O4BuYZtyvy8qXnUT6mPm2cVncd9
49X67zdDijFN8xAEZYux2DafzB1nbCqmOKsFIuwaNsMHpyBsaN2wplJZDTvo2JOY
VgHp+YuFscy8M2Nkj2OsYp9Sc86ZifU4Tjdwl0ovaCyBClV5Xx/aQyYnGVad+49f
odGzyFcIaCWvZUpzGq/vVppTsFHq84yZp82Tu8RgxAAaNLv9pRP5pdQNdw7zVdVN
cHSgdFe7sGBzBkHTBgToorwYi0rrxLQDu8YbvB3OWqqO3QRzQK8F2ihMVTvyOPaW
5J4CpJwzzVC+GrPmTLat8+VcRd/Z2hmq2xtSOnG8vkewfI2MiJ6j7uZf6YOgRRMV
NSfvdgfQ+fnVTK9o0Sy+oKIdGgZPMQYwC5Sbz1HVHkl4d7ScCtjTzHVoLBsWm6Nh
jjztq0lW6CcJ2wbeVDe77NPDdjyr711RAf7WoUSZKzqs0E2BwlM/2kw2GDkTT0vk
+R/2UATiu8k0ODzN7qXRsZ3v8fOr+eozJFnnk2r0azxMIjNLLS/GdaRI8ZPCr4tp
M7kSYLRSJhD1CI+cGZhp8n+Qiu5q781us9rUI94DhsTZbgeF5GiC12EHsP2+QR0Q
nF/aurUc4GB/7BtuVu6vBY0m/iOS4hozWBhc0SEV0SkkA6msxJbCavGijoYmx6Cn
7a4xlQnBUSUpV0svJtX36Yc9TFSpkl1ZLoJMP+pK2NmhL+m+quOACA08XtcLY46Q
MmB540/57l6gtFKScG87ZT8ZVdg1HRqDVVV2pRd17fc7CffhkxO6Hshsfo46QyYY
DEM2ls+Q0zDKObPgVnU9dTALroSvlfDV4GCH3vlsLQsiilZAzVoXgD5ki/lfQKsw
h8ABbHfx1rfP2MBUe4WxBy4oY+0nSVFHSjULfbLz8ZV5Z8+GZo5CY2M738P2J2ps
X+jGH6T/hOA/zbpgQOUB/oUZePADwcmCJKGe2yZTbppQyPpAC0nWn8+hIVLKxbJL
FDzPBsHuDCEfrxSBiykhfzp2Qy3IP48Xigao2W7lx2eweiJ0+mi1anNbB0w1fr8g
Fsy9xK+Qy2XPoR94kDlayhXzBoiqlmvp4bQbEJFZ1ZdD8xmw8XrumPQhJngXQrEw
2Ik99F12MhbQWJ/JP9TNzPfwdYV1MqGEpUoLVP2f/5t6c7J+PogGTFIHbyVsuu2n
3p63OEoMcMw1I9UjPvAIURUMYV5/sM/7DvcV0NFCZic2nzYgyE9+LCMZgSvb5kGQ
rBacAPfk3I2dHwt90RU9gibJ1sEIfRBXOoxIucF1VxOMB4SGSZDTdtScFxEwZjVg
AWxWc7bAGSCT/kPrDiKpeObd39fA/tJob27dVM/TkVQIdVCWdPcRBufkfu91QO5g
8yUxWZ6nlZ4D/2JtfaHDWi5exczm/JXEcUsuuKBGY5LJj0EBKoN3MGjIl9TaMfPk
0BhJ76w42JFaJ/6eg++l1y9V51/CXIJC5nrIUmOYkEGFYYTG1ChXMzkfK1vnUpAj
9E0ya6R+zps/myJI5DQb808m5KVSMlT4mEg6QxgkReVG1+je+HBFEas+iwFZQJVd
auMynC8N1aAzQvS86Tq4U4JC/FBhmomvqo3qKJKYffuWfOfHh1bUePlfmQZRSFIw
CFvqhoL9vKsC8hu8kv5CGx8RNNUBbaVFltqAApFiXV6gQzDHdpT6dbFrEtuPCDdZ
lrH+TUpXXgGLANK8OHMu5JXfAWsgF+cZK5/xjOiEL4aJxeiaN/hEvGZ/KLNhXqCy
bqRSa6i6a5wFT1Avd0/QP9mRLry7dqSSBoriuzuAyKjnsbn5uBX3iqcZ3Sw0g+cT
f0PFbATGUEk6gsu3SVy7GyaP1liYooBxtbZluNLUwBdfIzKstAePKrWRTYCRJ/u8
MOa77gBqlz1Xi1heHgyXa1QAZWJHIlQGeUE6N4Wd467rXaZJVzXDIms9O47teCyC
DwjMAVebk6SIccXQb8mHdSdLy+IPbV37fqzKWSDo4oh0EgWIEOoWFcvLSVekk3xs
P3/7/YbHGhuy715jHeAEMbmnapaevot4+5baPIS+z2NmhSxQv3VeBCsgBdgeY4CS
n+ouyR0l8rUG5ZlyQIztvoBpf/TlXQOCnH1FHlOSqA7jY5Dj/rZv/57pqY8w4XS9
fdnCO03QKurFGnNeCgI8FP1UX1dStlw7mEmRjrmqgYGe6zdiLq08B1Ey222X/+CL
/E+3GWrNPRukJWxqyGhd4wkX723Z3Yc88CKZUWIiabe9p1EFWwFfw5gUvnV74dp8
64n6rLHEuRaCrvp5pk6Y/GiX6aeC5NzOdgFimK2dyV7lwYRYga5Dpx3jYjW2SwaO
G9OdAGkbOfT6mtsV2BsIMbGj7FEin3MpVYMnmVI7ecb5CSWzq9Vv96XptOcImhJD
gM+HjWuuK7ezpAuXBjY5baSpqvQujjRSX3NcRb2p/2woKIONoyG1+ZG0bGtjJ2S3
VQU4muYg1kRzvAQ8r1wGq9c1YF+gMxMmZko3xessRrxUU85eXE1+H8/bKRupFl8V
g0nGVkx2nSpCQgBqI/piUJ6WVinBn9ECKs5bo1qVJ0LO3FKXxobfNCQXtFmhKFOq
pPPaCJPtWJTopas+wibr6NZlYSZA97Ccrt0Lg+eERngMGVl0XWfXTnV05X2gIGDa
b7JnEYAdihbVGoP9LiMyPBFRG1sXy9ENTzg+qFCo5c8yOlb4j6pfI7yCHuLFBV8Y
+oYW61DfYworGqh1MgAPtH1NLjW6xVs9DDmhrn8ku3SQHp0/r0Ics5DFLClrNZsl
kYUrQU9QC2K7OvPo0azuQ7rYq3IWuHF1x9vr7Jl1Aer8TnolRb0LjxQ6noIzxlmG
uxMSrv1YMutwv7VGc2olqnU1KiCC4J85WJUu+7x74EcKSbZ5KkiRq/mVr/lbotOg
DxShl5L6CLwrJKJyMNRqrG4rkUyvkztrkGuC4OeVZVqFXdlVD5Ckf5iGq4AUMuw1
i4zCre9VToBCYKZhn9duf2RRidxqC+2PbyL5s/+pBR9DXyAdbUcjG/IfI2gWiP72
GqWhWw7X6MJOkK8r9eiWj6L0KctS2EBYM9Z+Gl8OquJG7SpcNzZkp2KQ47ntMNrs
VxX3WnYHceL4Ms2sgICLaBGsrOrmozqbIbyKRXX7rGYfE2chzPt+lwpzHWJ+g3Ub
8Oi/oGHHnDyuyUZeFX21GS53NCl2xiwXFqLRlZ/BgpxAcUSXlREth4xwaaao70ki
C41hbwNyqD42/yBeAubVaaWc8qQ5NDV8Lt7+tTC9zQzERQW0VuMs96WLKWyn45B6
w/1BbrEghbl9TOy6YtPCTR8/gMiOWL+A4zMrYgI3hb9Uf8Nkbi5om+7s09c0TN+a
WOK6i54y5cHKD83OyK+yUcpq1uO+Jm/T2ET9w7JsS5Nlg473ZotocNgWbp+CDLtb
73QG/T5nS0r+Okb7tCnSTPVNerKqgvCWbefJkIA+323Om2xCMuf7L8jTYNMAT0aE
MxP4PRIXPSHyxWoXoq9k+rZma5IIeJ68px2V3eAFMpARW2H6PeYIlZoUHGDEV5V1
U9L+xKLCKuP8PAoZdMgcRPBEcaqUla4B2nGyVG1MtTCFWbum0NLfemau/t9eqSz+
p6RbGp7lUDk/zIDZnMZIMkgAHgEaXzlZ9LnxhHkRoYz8G2jBF85Zw2sk9RpabGJx
EAHkUC/DKy+7yAH+blRaPsXhe/VHudvgqNakgVU+gY8ph12tp4+89J8u/HvNLUd2
Z6PB1n9WWJIPlZVh19rkfvdUmhm79jsD/p7MDj7PhiUj4U6utTzdi1mmQpjzDmjj
l+mVbr8HkFYmTaMrxgQu9DXNeKhHEqAQyrMKMvOZEkh+ztYmTqLnIt5NH1Ieic7j
Fizq1PcOXoYEXnhOAJ95FP2P0F/YPUzJaUXwW3rMH4ieuBc7o8cH85rqN6otSnUf
Q6zbOliDcXR4ymACYk3i4gcTUmWk63IEV88fdIMsLqpPOLLL9qTWxCGDsuAD7wcf
Tm7tCWmmlQbMnFAc9YNzo9lbGn30jYxYubjRC11d7vvapAmQkbcUTZQGkf0pVN+j
3R53qRIXhRoFkW6gLAPTxp47Hhn+vuA3hWOFF6RpURLzaKAVycOHC+QTET8uipjk
t7FdLm96zVL0bIwpU+Q8xGBgV+CDwR3mu1S+Je3No5YJPLS4QAIZ3coLt8H4D/L5
HXANK14CipTN7X1tG2X08a7JYBeVrxSQSQ52JZYA3lG7bzTfQxNXNFXjHyXydKKh
/eF0gyBTFe2U5wj2ZDTn9d/OkNVchWEi9TYup6WxUL2c/1eqtWzBBzTfsr5jWBvw
O2NkLr21Tg+QYaF9M0nWTs3ktLXvpzWHzTMtL9vdVEGxdPruT1VdswORa8f56LUj
51jsBCxZAQRyxh+Hlm31pVahX5NtbNcdVpsk+ekuUMA7GP2/8b4xeLhh7hjjwD+Y
QMyPIbQ9s2o/ncoIKLHe/qih8CG7f2Y2QsCCcRHotH/Z1EF1vsImi6VKLQFXn3+H
QdYBIi3SAw8LQ3Cj4ssz+MweqLLYfZJ37CRPhroyKLS1pRLD+W6AE1dZ38BfBEp6
ezOwqBBcK0VuNkTkb8vcuUlXJDNlgbpvC9lz6lTah7oAMN3L1gmW9nLahM0dmvmt
klihHrPt/OFP1BGYBRnYeMLO9rPQI6hm/eQDiQBA4mLt9mkuzd+vIr8X6ZdJXfQn
vy9QTiUnSRfhik8EhqP0vgK/GQaVX40gOfTcT6TuDuxLr5XvsYcJ5Vriyk4xiZRj
krQHQkelFvIFfEl07HBihB1QY/U9IreVS+pbJvwvYjQvDUcxGc1C5OdLLW0rPEQq
3yrijDr0VlVWP4UQb+TqNbjLQRWYloQmIuC5CIZNepGrHVZo0dV3fi4uMTCAL1Ds
UPpTfgWFUnT+pKJPdnVGPn5/US0L4CWfr0MBDZ3hC7Ez0bfy72v2daF0HDia8htd
t7WGO7E9PWEse+jqKyXX7+1KsENFGmCdKn0r+yDpS+wSH7mtPkY4pmYVS9sypw6U
+aWa340ibVV/tTGwfU2NMj2rGe1kF5c2Moy+Qdo2TCu6uG8ZHH+410hjcpyOCyXM
rp3omubEDfoawFga2ZV3GMoYPJK/simLEMrdxQEPL+4/3RyhmY9/NrFrFoxnHfoi
vpeJLc4+ueMMJqiijDtTTUJYMva69hz6TaARnynC1/Tn8G0kPnzD8lQLHtrYvkpk
F2XqUOlvhQOrBn8Dkg7oCL65nqzai2uN57wAiyr5afBpfhoA1FexQ+oILcTaAcJp
dq/dof8oPS40sM5XLyrrUGhMqGmOZaw2jaeCjxpGc7hgDxIBrF9hct77HYz36x3Q
890MHLq8v/97gMyttkqqFvMLVCB0C32PH0AsZNqjrQrHNlMIOtpRjeF4Z+//Flnm
DVjFlai/V9ANiljYl5cWEUk0qoSAVwOB/+/RvOv1e0ft4cEiNb+5HnV5cDo0Kq9N
k1aJhkegK7h4ER/+X8GzlrEx/MSZVks2Pyvzhlupsi7u1873/9OI4GmGNlYu1ZbG
q3+Ti+RK+WALH+MeD31CiEOPYlkHOvGbn5FzxsQePSpI/3sS+OUVhGEwc9NMUtHo
3iCA1iGc8dIYrCAO4+J+dpJfC2oQ/P0EFAaiQo8N3rBtvUvHqBGDtulb5yGn3Xp1
2O1Xw0YIDqsSxDIuH07xZX8+0VSfcl1WQGhXERvuxvarDDrK6BEeVFbPUmWHUW3O
DshNBpFvQ5sucyhyjaWocQzQua6v8W3oYY+cd2byR9rvMAJGw6fLb4eW9L3vmK6S
plKk56eF4LozC3zsl6PQY4idS/MK/if6ZnoYmEO9Gt93ToGB69j72l44POWGmLqD
Yy50gfotFzItN7lnTDM+z6zPZ/mALy+MU9wnWMj4WHGekkaz5sk9GxjnsgQprXiz
wUeG/VnihzajNPp/POE5e6irKxSn1egD8hZ9LPTxL/g6AYn9NT9hCOsp+2VtVt8Q
IG1G1lwJ7pHoRYkHydkHZ2e6eZMENBOU4OjRbhXTNAaoxvKYaCmeWvsDJ4P+hXOC
YhFMc/PlDrgZNA1n229tJ4yum/2DRQTBxXcAV1BDuyLTkGcVlMfaCV6WpFx/ESiT
QG/1k8vAmXp9NhRmLpoKhLpYRGzFlbZv7+qlvo/zwXmG+PLZYC3PI06kvJwxUser
uRBujFFPepZ8d9rFVQzODJ6QuVKW/eMbHCnGMWklD2QdbMDbU4ABGtwMz1Xh6s97
iwmxgboBeW3JFddAjc18skR2RIWCgJtCiAsunpfz+OXjloFIRRRQhyHpqkRW6hJ6
fD5VB88el5D+Hq1WIsmhp4awfyUZ1vk3CWBkUehwg8ek8VfcBESBLoDCvHbvR+Ap
tIUEa4yUtrcbiZVhopaJia++wqi3vY2bbxqIFd8KsxnGomQcKMICoBAzd4N1DpBl
r5MGyKVEHm4Yhx+s/hh2P9nO/Wzr5LYCoh/gCK6BDJQ64FaT2zuIKB4thEJqYHwM
MgNHoD/SXxjjPu5KMZx86xSg3Qte6vigcmoGeLaNOI16DzhQSMuRpNV6YIyciWKH
0MIhC30rlNsLY2gPP7v/fpzDNwqFIxTVibiEHDXIsPfG24wj0anwwYbhlcr6Kkg/
/ppf9c3ykIw964sZaLLzb9u7I9IBemgnTqNT56eULHWoctBRuo4vRBJGDx9/F0yL
HXo6nDXfQOP83mG4oVsOKiz8WTwFN/0v2LuoTYsD8D6FCx4letxzmYMNoIjWE7il
SZYTzp2e07xTs7n9hvht5oTrwi3k/0z1g3HCQNeP3HAWh3hG6P6yWSw62lieFZxb
XPFBaJGEir2at6J2dhw5zq66NPwaA1xkw8AkgwP7wB2K4qQcE2DelFtrNlZvpRoK
8X88jnB7Z2dPhzUYvnMS2bsTFv4WYjbh4Lwkfn8HF/98PyXd2VXkoEGOWa+WSj25
zbEA1IenJDcFTUxbFUTVC78KS7/qdfegeGhcCG1k8v3LzCVpYxF+8j1KttStMHSC
aQaJm5hJ2gzmouFaSAhWXqT3Ya7HiuprWxLk//MGly8UE9p+aDbSeMdFd8WIbbbi
4pdnR2LJjutAkAZhWu6NCxrGhOaK37vI5wi/wp9ViNd3VX11/MKrpNwlugEKa7JV
4cJACC30ZInTq7uMFBmPwwP8+trXP8Vem9I61sI+R+BnuFoVEhKWmqu5l/HZmAki
7m8OFBk33gcdxqWbMNvKS00Of4rucSIW92qe6p1ojG7W08rrucmBsRQeRQB04IJi
qJ8T7UCGWnZNSbfK9BuVELjVyMGakOOon0nPI/QVKDd1pXLtPMZFYMlYh3UX6aLV
onbtCnaP2SVgvtL8MqXX3Je5Xz/j+VAuAS0lZdcaSuBjJ+M3m8JSTds14c+EzUBw
RESHngnJY87FMxlDyQBeUAvX9VqdKsESh2i55qxbEXLod0xVqovIkA1R0soXeR/2
rJMAZBtGTMp6txRs3DZZnUASVed++2nFz3I2efOmSI4ysMRhB5+JWGyyhqE/TzuE
7JyJ0GrZiO/6Y06bURsGe+jkTTrG8tmZMO1QCX3OOT4rsk4ILuypIWB14afRTrzX
2slWzBZ2v5/+/sR8HWsz6pr/cPOas1YDatJUUkxphJbuDg+g4At+CVYW0uy+I4mq
zf/DGREESF9qEGNsTX34OzvIsV+vAsHCpJBr3xiONRGAOi2vU23Jtij7waJIcGX7
35Vf+KVpuxxLyHwV2Khs7oRgKgrmfd6M0BMxYc+H2oGqWskEVDBB6eKFrbtHUS5U
nDFA7aE8ukqrGx+N+VleJnmjAlFtQhSUpL5MXpC5KNRTLd01oYlco8o0bTdCPlHF
Fqtb5Hn6f2LTzc17VZcKFB0RkDYjMzaQ59gMAy8YGuNTZ57AwtYEzl91Rq1QPl/j
XuQb2lCSBPyHX7h0eo7QyQDeDcMwTXrzxGX12FwFL/5nWWeqKIZvStIwjNi2iUQU
w6m57Z18d0L9vvFf0KcYzA/hpxZJqtY/dsMuxzadn7M0SVcidN3JWThjA8GJq3Qo
OUuvKZtJdfEKqU9UNw0qdfCPq7QkeoM1EZ5c4nxCOMg65yplHYgq+n/n4blfrYF0
HZ/JMf8geMHvKJut075rw6XzESRyJT7wLGoQTAhgs9mp3FQemsQgKqYiDFphVWZK
GZpKBycPcdGxiwEJTLPNjFeXqPauDLbibWTyiPoXsUYPg69bGJ3WcbYEaAJYg7+Y
olQKB3/IwOaSqbAk5miVLk/SERB7hL0Nu/87j6/VRIqCA5AjW94TGWbFr7RXjvUi
/iLy/V8fkRX6UCcEr4j7qGmdJroGLSJYaB7LwqC0+V69PTf9zqx1D6hIYsOMhcCk
Pq/0K0oTHMVZDubaBKAqK0jih2xeVaSVIO0ctFiFy0kyhlhIUXev8L6pIdbeJLK/
9OULi7PgzfJtW/XcLT84/2eRpyOoPgTCQGIz3dBxd/jOgka8lrL+A/IPUXT9bk7V
clQI4JrucuHqo1KvJ5RsfvBrB6UsVsI4Q4ByHrRP3IPEGUilweZV9lEErlTmuhW/
FLCciU6xtLhdq7GAJAUlp98mYVOYtSBq+toXCA0OBEV/smslEjwOQA8SA634VTpE
w6R6Cl7q8If3+CoICDT3yWHlvw48JqNsPqFpFp2JWVOUvLdS+XAHJYe1UiRAJKum
JmfcJ2v6RtCCfqQZBsH9UyzlYQCqYq0D011WlZ2MBllRB8SHF0IXakjqtfVpeMJk
MPI/yYDBzIVUQdhiEN+8CxaMrNB0iKmwqifl2GnwQUxLH7TZlXQ45FMM78XBqiXI
fV9+pebtFrqU3Bu1HrMFAIjo3gm9ZehaMV+w73P23EfUHd+TZimy5vsHLqabdZ+5
a+fZkYX52FnJLSncff2HmEH7lDx1DJvyy2cwKhtZWX7hlSn8uAeC7M4h6zRakoOD
Q52SBzN0/u4Nka9sIanojxJ8m3BD8VOJNPTpCz5VhagJQ4GaUF8/NxcYJUeP905m
qYMKhK2ePGmPNZ/65hlJuu+DdWc+Xx1gQJJUPYl8MNWK0/mIudxUtdtPICK1GJxk
a6EfurS4FqtBwmRluuvbJ7VgqHiaLwaD1gZEnyWOa8z3SVdvS6k509Ga1e1eyyu2
6ancWVNgp8jeF0ClZv6t1nNxmyFLHXnQbXdqk+UznCVpc8MuaQKqCmBZ09jyKbNA
Fa8z5iYGkYju3mSpNP8Cmh5Ykh6UdkEOO9Tz+/bQnwjAqXHgg5RMi/I5fY6hN/5z
vymA73edds5MmWCfdPO2KvdADb76kK+yVAzPWLVSEv3rU2DXS1GNaEUJnnRUnb6h
z4a3g+RTAOtkdm0oz3JrmauzXbRBMz15tXAZFbQIdKA87BIfKFZd3UwlwRpcAgX/
vf8Riu0bmzurOWnmwT+cLpA3IMGaB4IbtYz7SgMaqQQRUvgWmilqa/tOynrNStDT
CxhM7wuB0IieZtYcwA7k0yCiDVwnVbWMMwYRgmGEmPRlacbxlmt0SB7UKFKEMK9p
zzTM7fYamkwhsvxUFv6BiZ34QGmH9UPZ7bYzLbBNMDdVtkulcci6G/fftMRlFuXW
tJ9bBihUfgJGAMZjZjIX9unbgVWqKMBwAuAa5Swmnuf59E3bjsYUrm2/wEuxPGd4
vkzu8Ky7EAC9jLIiTs3DJMhwWWLSRpre8rgRPEve+p64XTfBehinzOz0etwoCkRc
yxfh/F3DyMpo/P3wi3N6eJCyMsJ5aGfiVnc9n7uy92evCdDCsRusvdC0HLtDqdB3
gHXefmMAdeH1LoLLwam1DuTDGNdjmTqR2CG5PXQItmtYfPZZhTCxk/oQg2y7ETZI
1okraJedsGQk5N7LprsnVtjVbfyWzzgjDUMIYRjVZAVVInsv9NtNjYltapiRBOY1
Q2f3Dl26nxC7gTBWpviYNbbf3Wfo4Yrf06LnB5g80Ba2+nRpjVOly3WLxoqhbbxh
mMmv92jD8YFjPiyOv79hxU8PC8FtawSVkZKVWct2GtlEEzSJo+Cndr/EmGQS+/SV
nNDJgUctdG5f3RiRtKtdy8fjk6tCbPBBgvnRu65LMSLs4NU2Boqd2fcHQsZsOKUv
MRDejF3o68ygGLuIUuOza4XZcs9znLQ5C5Ua3x49JOudClPv+ISV65CJiqHkLlMv
eRV4obsLvc6bZ0wMTf0qNc7YrIkuWmimWUc1hXU6C3CF7caALlVHK3jb67fxdVc/
oDjV2a2mDPJNsqW8h5fs4pW+OMUOOtls2eRAE72Q6XIwjj7LJHJuLuQ3pQNcRCrs
SxUz7QXIPYK/upR7RKXUee4L1Ijy+5jFVPVVV9yG0wlCTwbQTepSXm4QuIUOaHul
p9fNN94U6v7B5WOYfXMCkpO8HrYT9k97fo8EUhAyeCE/2+RGISsYdQQHVreofUQP
WyLLp89ILzf0MBCG/IAKFVG7OpePDv0KJP3EqDAGyJmU9zSJiYIXYgJoWiqfLav1
mppZdc5UEeG1kt7gCTqZAkO9Aqb4DYeG+A/36RQOvs08E1bEcOvnYjjg3O/kpotS
muDAjdTOF0yH7WNVHuVL/LwPey+FJX5xqxAQtq1Kh5rb23+3+kt+drH0TcKNWgff
DjyKSDWFFRzd8yLdYOk7CNZxSCG+BxoGz+DKduBOIQ9B7EZaqg/XfltCdJVPrpRI
h3T6T3knG738QhZbDocNPeiMKQoXUdM26FcybGNoYr8T5z4AFZ9A6/5HVSwNty5Y
gqFg253PJ0p7Tw0CoZJmepfP71SJoXjE+vkyppizX3HmnPNOOKiYjAjaEg+TRBPJ
DjqEIdoiBQBN19D63mOMPb87I9fAtcPgXzt+rUYMsv8HmEACgA/GVgANq9b4yLNz
eHzK44HIg+wIS+qguKIJxtpsPy4SrL85xCLFFytR5Xa+QOi7uhvWgFeiS5yg7YLO
PWFjfTVvrtLhUoq531hNLRq9AdpNeJHvpnfxUdIgYvZpFNefYhhh9CSn8HBXvkcY
PGvIp6T75DeHxgeU9IsjxKsWl0zVoqcgU7iouL4mauioUBdCgGZYyF4eCVyeo93H
GKMJYmHFBAbJcWCJH+m5qFpfDVWItJAbpKQwnW6pzZHcWpCBQjCL2UUEoLpEUO5o
PPm9YLF+I8BKBEeunO4d+iXN4o4m091Z5SKH2jkjAhyRi68OV7hrC7LwLeBGnp3b
6vBhz+/gQk8ASvu3a8aIt4ZVRQtSTgKQderlHMAgJ5h752R1+ts3EBsJwW/+SU5c
DNO26T7yGUNia4ItiAMbELtaDE9k/cvmc3xbY1Yb/14HSNxcHvQLCzMDTXQDZkyv
VdO6dvcemSC+uNNBPgMAoWy+YWcyL8tBcs+9shEoSybcx6k2ne0xqtul+Yan0eK0
W3p2xTvD0+9yERFyvbc1qBmByGDqTOebB5EaMv6ewHORPRj3MfOeUMasxo4X7ExQ
Shpvtla+qiZ2RyXd5SWSam9mfU9Zw+dwXg+qylKS0y7wCWNSHiK+zJeF1JUBV6o1
y+cjg9pa/62AKC8aLfpXK3VGhxMiNysy6LbSynGl92gXTGZPnkyHels1RfvutHJb
2QFa7fkUQTYjsyaE91oZkauuMcz1843r8eVT+eOE3zqBbyW9EJfhVVLFVEf4T+Kl
ujPwxIOjXw38rhnWrRjiUk+cPdxi4voq+DzX8WP/dnsB2cQOLivzsr3DyIN3GzQ4
1H81YEq97LNkRA0y0YmgZsp2JREl5WZSsAt29W08GTIkc4amQ1pu02maAcPwntdY
TBcqExg2AG2e7Z5gqxsjjFrCOpQp2Amg0MmDRbW4vxFUiwJB2vlZnwrx/h+sBLBT
PkZicCX4rCm6KJZnUds4SUwUJ4KYlTBAOpTmScovDvAuUtKRv7Ro8rRE1I8Psw2L
jBdU1tAPJ9DqHU/YNwYGcCCwLEU0wQ0SoDMbUAyaEpAVSeyvM1vv9VQnLY/mjJ5S
MmG1Z8upNasd8OUZxur+p0YKVGg7a6w4nez6S/VZz7QQAYLZlsx9K6CZnd1Vt60T
belSBbk6ZwXhD15Yq2gezdqiUXkAj5dOXWdQ1QTvdk8d23RSpRiPmWJ9y2/YlVnJ
467yoB5xEBNcRgGcEcrKNGjozsYhL3W3uLWzPqKgjsFR1BfFNYe9izkFr+9pWnTj
JJ9vm403Jg3U0m4cSqzSy77X51fqp97pZOhR37vZc3ZEDT1lVGQxAk1p7R6fLmgn
H20gL83uN4wGw1Cxicy+j1jXCZ4gr0ZuJET7UrWxIy8sV0PmSwflDOt0Pb84f3iW
Sw23YevxI8X12ySHD6ngeR9RvBrJiy9J/ihsgl+fnnh5fnWim1LakJJQWUV+m/pp
DBoK62m3E8EGMVGswyGCh79/2QWfm9RfKBGCheRJlt7n0k81tufLqUd94FJ7s3hm
+JQkgysRCQDfAje715NHRJB1GJUKc599nraGSqKFKpbrLAk4vOQdX6ALyH1I5mZQ
zPDjbb3raTrneTwd8TopfGnwb3ubOBC3soh5+CWa/dYT0ppTwio2+CJrihxfyZx/
5GMkphh4GOpfESFNvxX4GxxGGJASsBuOImpRAFI10l7aWgy0iHghhRrgX7c/FQsM
t7OTnVY4qU1O6dquKLNnawwx1o59OBJVj+pydyojq1kpa5wS74Ja1cvUeBC9umN/
h43sY/bdf+llaI9wDSgr8ixfGrkE8Yrap633J5921jFTDrT6RYlDu0JE22jJ5u4D
KBRbM4xFQYkIfvrSVP4bGInWf5tzVzVkzR+vZcZhyFTUrUXHlzvrHRGBAKOCc+KR
sJ5wv7Z44PQ8rC4YPunNmNzcM4WbtIXE2P8racXUzEM99pvatgRLVCBrUSjugiZ2
2+3LJK360cyrq8UIWi4GOcuWkTCGL5AJ0TNmNczRb6bQf5b8fwqH8GCFiqtL5KRV
ssuTsavylibOtWcPCy7tieH7EzUFML6e5HDRiazbLgu3J4/V0fcuBl21xyJ9TuqN
KcmoGjbT/QhR4mhn8b4mAizumYKovKIyRD8PY2LU2f62FQkWL8SGHtWYF6nWdTWN
VNUFM61VdFBabS5j0Togmhqi9tOwVdjTvqMHZ2iIGJyfZrdQv7TNhsAlAb/fpIkZ
8JiR1v+QoTJnI8NhsV7E8u3SBzkKEc8Gno4f4eM0Ca4Iw3CYV+eIvqX6v8cxstuq
rmGL5aUE4QSHWwpznY5hGrgVofjjbFROC27OGwNHuxhNxJlsd50O7Yca3NNZGQrB
G9D9SScY2EkjW1fRpkSoknfm8PZJ4vqxAipoUoF/e7RD481wN1VckX6njdgzxJUH
y3GAaQu2DuIUlsrHe9iWkYWlT+30R/bq2X87vcUwJGdOnHdA5s/f5AsWlma8LkpF
d7uDm20MckAuN+RMDUklxzql4RD73KzlJQV911xs2DVMtNK330bPsL7EUalqiMxp
zDWi8IQ/vPQbTTfbwX4TZVvdx4+yoWn1J9JAQbfLR9Pia0is7jY7fGDaw0VzIuBd
4bTCMPNne0tGlGm2Qu+h8qQoBbB7hDSIxPDYbPyKURFlic+1/NYwq3UMZdtYc73V
B1UOMsNSSUi/S9J2pQqkVJjiFLrytcZkcl9gbnPcw25r37Quqcp3LYmqS58nlmMp
2hiF38CIbwXsx0OiKvdex8Tpc5vFBI0Y1F2hrILW74vaMA+SgiK/z/DS+EtF81y8
gqAuCtZa5tRPR3EjH7pL0IuuvzH7NGrY6gTf885PxRm8D/dOkpXjjxp75feNXvUH
4ZRLrlkKVMV3tP0+SEX1ypmCqLUzFGqubxAi2lsEOan2oeimRR4pge0a+qjmrKmm
pDBoYxUmK/ZKj7KHoSgkgc/aEcf8K7cT9xUpTiBTDXMqgNnlwogUCnL8+NsxRJCE
VaZ/qlhuinGCf2RGtQpXkC1vZTJADK/nrbi/WNCoucosTLjS+Yj4CxqJv/P2Pec2
/IjvLSbPQ+QJaXVWs4ZkmuIpuApuRgO76Wl2tZ4KsgvZzzDfRfTNoAPgRVzLKcHh
rh/EzZZXrS2cM05U8QObEz53I/2RH2H3MYKX2jZmmeyTi3opeBRyDDZuhmzaQPFy
kxV+GNkKBX+pEyOTHvtunYzAQTg0RkK1t2BXAKylG0lSq3k8+WnyhNUWKFQUR4q/
dimpuMXeGfMxnrnPRyX4OkIBsfikMtckdm//GnYHXyaMe473KK5XCL5hY0LJTYhW
br9kedyy8uADXqDuHLX2W/WtkgdbpzrU4NaLAbyqvw/LYLjYa9Iq+p7ubXNAsUet
hiZcw66IveXVrwDhduiCWOh1gJ7FzmOEvp6WfLJ+Uhp3Ap/1YJrDu5FLjBkCLgKR
rmodkoRpvxJpwSkmXmK0BFU2mYekEymD/+yZunZ1z6S16Blt51Hoi1xF+cBg1JhA
GqPxCZkilRKcBpaVsoaT+so+Kmx9RlLK3SZSop0l6uVh2J7Dm3Ki9cYXI99lr8G1
BRS/AwN31epy40rZ9OKu2i67BsoFy3Oy601NJEQyb/WjAsh8OhtcYikCx/wSzNdl
GahZz8x2MULKB6GnJlgaHCkae9aRUX0yd7uIxUIKS9oQ8eDXjusl1DdBDDuppVye
NdXrXZZZfo0C2B+nfGmrOcSkPQG5Z7f9aViu9QRfYC1ByiMrHlDvLWga8eoELyBE
zl6l8SwsB02RTT9Py3IcPI62DtwE7SYrXtEWoMvNwMDHNzEk/ZAQpdftR699wjs4
WmMvYfrg631+SxMXBgNpb42uYhxhtzGUSp/W9q1WMpYqB/hOGmkD+paCsnpkOJVE
EZrApaSJcfi67Ksr3Rr7xNCsTW2nu0+PHgWaoACxw88sM2kYhmi65RKAz6taGKGP
ddQFA4w6nFC3ZAYm8VrpKKBbL4jH18seyqre7v5g/1rIa9P1vOfvQQj2I70+z48u
YR0hS0xEWCAtM/E2H+JWMcECgfHSVkTUAMsETtOQ+RBFYfDa5CjlVjKBpj8EeykE
x+cmrqF88Mb73sbeubqMMvQpTRgrU8ehebRXJib/R5gyhdyi5+MlSAVBgqhpodrN
DoqEsBM29GDUVqW/MrC8c6RDtwT2+woMw+ty3MRLKuGnvkQuGzq2srCLZHjZtHu/
tk11i56TVJFFkUYj0xPa48zDddEIkurLcbghBQYOgjJlXu4yXTSaYR1Q3SybJ8f/
UNYVqnY/il6xXV+tcsO7GE3zcXFvofBUSfm4zX1R7fplpgSUlChiI1hjdQ+VshOY
mDbQRe9fDAKVAA7S0XNQh7vlG0ozcLbIhQV3Bt8EWU9y58nb17dWkRuKqEiwQ059
02irio30ig5JmBrhwDrWEm4IJKF1cb6AXtsc7eVQ13+QZVF2DliC/zlCugfeSfKX
P8DEGxF+1xu1mb1bTqc3YHxC1dJD0ey7dOzuWCOsG0WizPfCvyxXaJtkkCtbB7aW
CokjtaGGXbdqCbSQk3iZw2RGfTtVPEpiXIv+d/9FyCzvmS3pLHhjhaFSxGwZ+qwI
zOPfZwa0MWfkpPq2/Xu2p+Ml6MVH0AedjuCHXY2V+kizddLACY2zBY5s9orUgWNi
2Tk7Yf5xJFyjdrSZDVlsG/giHK5zBwfGewV0ljowUmSOdcuS7SMU64yXQhwCu4sA
tGw95lNQrrqromxUUI5in+uTlLgVX1Kk9Wbo1pG26zJYvfCyMTkq7UnkgK7vDzm4
Xhpz7UwTQUVL3dWUHfCjMwp8qgMbqMduP5VqTKRwaYkbFdenI9XK91D1jpgCYL7K
DVvOcpPkrVWycPWpNuwnA7Ns4mV8wZ7tcP6nVtdt4TRZ1jLOafJXNyiieXQ3bJIi
zVOPCvoR3z08EliP98fxQhGgaNoI5p9QHrJ0TSdxtCsgSS2q0k5SDpxraWKhBHHA
fxyOhuGX2zEgQI4mTuLQMqwnimV/6IvZ8Cg2cQuIWxyK8D7hSNy2/jUlZf8nBWLO
gMe1FHZQimYHiHcfdyZWQUNPtWmUG/uwMFNTpWHnH3fJ0miH9ADqDMfzo2FsPLk3
SPfv9vCkNskcniwaH8PYDZWLVV0jlxly7mPVmtQ4d3ozD8pA2lAry50+lWjhCp5i
pUySnIhBiviM1/lMVFCIfCAYAl9FK8T4C1f1rSfgYBN5lNIUELZYcdYPhkvvLotn
GTeH6vZTauHQPQaDkQVcZLMAELbOHUyInMUCBSMpTbX9VZXW8ekmnvypw5Weq2LH
T66zXx2KOekZiUxh1+oVVl/E+PrIybUAQKgmmpHsrm2m/RAw8UOOi14iejwjNUG8
wqMEq3ZYiSeWgHTiqDg/6suoqV5MQiTna1mvyJthKnRxZe719m07ftqfM/4Bp6hY
cosrt1yGf0R9fwKyz+Sot/Ha8mri/ShT46Y3mcNvqOe2ejISqKObSeR4IC/d9e1g
+P5Rrcy3RJgjWmgGaNtTD5qT+s+sEhM7FtMipsfNmRKlDofwWR/ii+TQOYn2x++t
UDsNJPQQmgR1jgP6sUarm/iMmYfKCWgWUP+lX+PIqXf+B/S8dwEy7yK9qWN5QhcX
1+ddkqr444YsrKw7kRDcxbmAj4WcpRpNlKy+PtGn97PW94ACpwHDf7vBE9UmhpHz
vz+SAzt7nc9PXpR0UtPDmfvtR36VNjLwjfi0MQXrcxsQ2K3WrMCuEbvSIgVlkmTW
Pj3Bw0nD0OW/ND+SObdZ9ud0gztQc51QrOjBA/Tv+wTXaZ/aiZjKCxwJvH4qbFve
N6Y7F7ZjpnXjdOa68vvMZQpZonxSU2SbD0MSj0lB8WjAQD7WNLaEy6/hwZHzFy3V
OICnk116LiQbiFjQWYcq8FDb0vd3xq/LcU6IbW/NLdqYcnMhdkb9eXO8IxLC3DxX
spVVtYboeEDi5uV6pK9htqaQ58+jNZ2WfFkp+0aHO8e+5nd/8yBzh1vDr29mi3Br
RZpLsdI09XHthVWLdZFozGj6W6HoKnNHKzk5JRaualtueVfF/LTv96maNSWMyFEi
ajYmcB4VhdvKP82SDEPUnX+RjQNUHGCg8yeDH+Lx4zrC9VCgetcZi2vTjEqLndA2
4zEtq+zeV1/Uz71epUMhvtskQP+T73BN2fg29TbXl1k6H2S6i4qd37+uDzxYeNge
McZthk54KmQWepjA4GBbdnheWuytaMo1MwFGA4BPHGYwi4JLqbc1MOBtDvoxLZMh
EV08p2WCOqD5X3F2+buCieYfE4GJubvPM1gKEH37UNzxnDOwdEiIWisUZyMFjWPy
oiH7pktFPXGDjcab3IjmcxnJyEFVvShvRpBYmSnc8hqNg4oCdvmGtJhOToQT8o/+
wIXXePt+CknhIpMvGloqpR0ZzslF6caNi3R41dvVf1PjhdhQtzq67Wpt/hkj98xn
uD9Mk4diE46uPR5ldx8rHtyBniQKA0tPh/0RFUELWaoas1nxWHIK3U0KUFkP6mBH
E7uvD0yoW9Q4SvTNEuTe1NoMbhABhvkcBpalyjEsWlXvxmAJlQdbm8B/D5HJIv3h
tGSjexoq/beLqWFSYoXtmSecdZRIoVg9N4UpzO0LjuS0qAS/T3eBROpUkL1e9aPk
nqwesD7rYY11pLkqfWPv2Bi4pXKHgpaXWacrP/8xNGxeumoc3i3kCHBcSQ+ruwR0
Sszw+Fns2IkdCGpdCPFDc/eMLMPb6d5aAVSHxlx7FUmdpYIbvmD/pY9n37Xf/vqn
gIuo8r2KNJiwRS0RyInSITPFQennDn0JoSnoMaGqd6wQb+ncKE6Po2Adu/4AekFP
bMqBLSYBlYOYR9BA9gAcAYt/qrdGjhQdIUWXy9VsE/8N5gx9C8MPswt0InGQFDwd
8HfDqdGg6OkgLZM85Jj/BU0n2vWcXX/YL3cYI2udgNibKBatT/VJKL1Avq4vu2fM
eW9gWw+ydFu32G3RoOFXUNg8uqtSedBTuBNzIpQPbpeUjD9FvrBI36eRIrgWIfj1
u+Kgm8vHr+jfzJbcwDKj3C/nwwwgoN5KiDicjwK45GKtreuzCJYbUN0OcHDdGMbH
+LJ1+mJVt9C0kHM0zxGbct5z2Ytsdg7QKIDU/awWkX6vnmu7M/04AuxV8copN7yI
lRwkgvqVvAI2tCaCkrNCXhDPUoPGPKbyXXgwUicUvfsdQhQQXRnC9F2xEnA27HsQ
ebe+zhyOhxxeCxDmBETnnctvGhWt4k3K2BVjYNZDOpTx1SXG9KtFN8a3ZY1a+FdU
1IwnKAyxdmgsU8YuVaw5kauyY7IyHY3Dybr8R93Kd8dG4Rd3ZjgITuihO7UYnlqE
v85HDQAroLeBLHYn7dqFsmUackuMHhWHkKz8LiX1s6YaLl9z8+AI7mRT+TJxvcj3
Iuc/YmimIPGpKHrc/515DmDh7/PiofGtG8qCNIIkN2ghOxlHeanifZjZDm63zC/l
LUiD0vyLneV0Fm3vzwHzvKHzJLDa5acaTOtwW5EisKIW/n5KYxh9HL6mGLZ3wmHF
T2h7Q8nSRqXZ6rmv9cvxixu8Z7vu8zYDMlF+xDQ/Uu77TuXA0yFKK8vniTsAdDNI
aXlpYGMkwu3fKwEAT5WwfGnwGZLYjUmpnkjB+OmQJhVr4bQD0OWvJdzr3/qBXFRv
sGXWCogiXjpof5jnNMJnTf0wwCv7/U5MwSUJgP81T0xMigjXxi5/NHNInk+ypxok
/NH7qrPuEHLJO7ry2q/X2j3NwWO5rzgNnQmlkUJ9ieWU3jFP4iSmTRYJl0rktsKa
OmM5axrJsETNu6JGOJa2k/aPq1aAWv9/jeqG6bhWCmsRdmpkHXirUgKM7Y+b36Mb
8s8tl943yG4c6rJfP6Pq28YvmXvwiF05/79rgRz8uxNpF3EdJ10Q7NZLC5jS9TVT
p8R/d/qZlpLEUL/tsJo8nUwLavnhH6/OM0EWWf7DWaaLR9TEYewmsbA7oLMfXZaX
Wzf1+E7L2cHFfGFGltqlxHNY/koc7+33YHEfywREZt5zwM5UBFKE/jixInOnhgkr
LUuWkNGRJYsMdSR3a0G+Fcl+YniOQgZpo+J7zbwf+RnAYJI6OWsxy/anpwAY1QFv
APch+/yH7wzHf50/DkcafLUn0EphR0ua7DGNg1xp3jT2+aJvwD+kwK9XhaNPnfni
dOCWB0Cx99gFUYEJWyOy1SgT+hByIpweEU3Y+97JkhLQVNYhJzzHYRNAVL2WgENk
oSfhLplJ2EkXs63OUgDmiTZk2PZL4qQdPDSEsaanus3J5lY/DbKtblcVaxjRVfYA
OVIf4g/M5C3s86jfTqwdK6nH0DHaZq3Fn3eIa1Z/Na4KZq0SqI3htu85q/2WoRBs
JG8BRu9vuD/iycHbk8rIJhsME493X+2Oz+WrMJbcw9gVEn3fHtK/RzmPOlv0qKal
ipaH9WOQO8hOTXJqSaSeB84aQc9DXLECoRAXCmBK9mBnuV5vP43x+Q/p4gaUSyV7
8wUVafKJfSBC3InMvdzAgFkfGB5UItW2uiqryr9rISa245+OKwaqRp1tuG6OJS65
0HZBZmoGIU0BFIPTULHrrZy5Le7Hhpyhps7gMJyCKgH5a6VssjkUCf8i6LC+QJsL
vuiqjAA7hO7x9v/6Zjqre0BWyvBjt5V2blTxvB93QQTlNtv5kBFzDg1oo8HXbkkO
g/ZE+OkuNLDDnWHtZMOA9ByHSaQ7ffC2Cusb9Gnr2AUnvW+vGAillnhty6YGi3xj
C1zPJRkww+VMcrlkqU1Od2ag0K/RtpeOaoRUahtWt29FQw2WuQ9HUxm/SEBLkbTi
TzMN/CX1TA2dTiGHpD/1baxAFpo6E8ytuML9BNZYKN7m7CPNNeD1HQsfmduVjsgD
lVDn0MdGGOi+SDYzoGavuGM5p2BwLm/nn4bKZKwjt4WPaF8l4b/6BctuGZIjQTMG
cM3MkxKXda2eW+g/ZAJDxP+EhYHy3QiK/ye0LcjcWGjnwwXqNAol2I5UsD1TMI7Z
wy/Lb0zcy96VmMTNpTbabrWi9l7LL7hSlAHJYbi8mgsHZ38FWN9A6e/61gTmbm1u
SVgeRE2aa7W11UcwHbTdCsDUYRofno2MNGkr2POsGzb9wxoOzUuXhyqa5W6xRDUH
Kja9tflK1tFjvcgDR4aFElYRzIoqCEfqPFkuYbXDCiVZsEHJ+YNtBEZhUmamTRfT
KRq6tZRAzkyvVOsXOyJSLVnf2sLCLOOGuSAQD0GQMqTaMl4GFqFldoflQ6Oed4oy
D/t20BRwcNH7Km+PmS/rsJ8YvGYA0DHDvCQMNOwI0h8xW3SqHi8LxIFFZFPCh73b
R7/lzlcPvGNRpMlRvuvu5O3qBiOER81++WMkP9fc7J2e6OoBVgA9bdmy9f7ifDLZ
aRDfp6BnDWt/YVYo47CyGDCg6McbJ8f1Dbw8KzUUtk8R3faZhZfSUYQhLevQvN0G
kTQVy+TE7evPk9q77hPK6qINaSEO07zA77lQCLrJw10puttgoTyWb58CZokwkKAC
J0oWksjFFy045EHyoZqClULw7CsLfL9G6WgtVvpu4I5KTlQ2mIM1MwbFGhRpapnA
6IeH13B5m7TNWUAlAsUmz3zyPJhNRPBdQqj9uHfB4bVEX/sRQ9RCRv/dGtzJiZ5v
ott6TG/+wi7eBJgo5DHobH5ZK6ZSWi4hiuAs1aSCK2lu3+zOhN+fjCa7HkJ4YqYT
E7RcgDfaCkku91x9QoFm2reBVyFKS9vphFtad4C9fEdNo7sN6mB5ZZR4JkMZ6vGJ
UhVN7GiZmLBXs/CNNWIelYaKqyQemWfmMYIJBbI5yy23AadBaVP/yU3gyeod2eva
AgP6mdcRfga3INREkKBFF0VF0Wc/fQzoMaVpUkYgyU/uJfu5jaT3RlymO4DEfqHv
Ukf4C6ULD7bv/HY3i4t7bJfhhPZQnISAV4W4uLq3G8mNRmpn6Fb7aXPu++s8CLrA
jNDDKK/pEKpNPUmYoCLiMd2YU1fL2Q6r68dboIU5q1zxRDxWuz1qEn8RLLBSXLS3
/1rinJvygv4xx8psDZkGwmTffYqkk8Tty0H6OsaF0C6iw79arM0JE3xoAYLN5cu6
Ir3xxdowZvxRVjrVyn2mH7IVXDFVF1iDb1HaxBvcqMA0D8ztRYq2hv42Ad1qUXBr
QfVrFVM8ddX67K9idrEo/u5zoTNM7cp2Cisuc9zFQhFquOGSdYB+wH5AfrYNH1l/
HMda7Tz8VhdxxcooJHPKiO6XCwVRO5I38tPcfwwMq8Z/i4NZYQEiRnsMoJ5UmFYD
Z+zJPAgk8FEWUNrea1v1dld8pGFpXjp63tuyxUe01FeZg0Tyx+girBogIU/Ila7V
R2WBoK8HtfRTF+cDmYhPXV9/1RxMDWR8BDvAB4hSYVHlqLJA1d/ZvUqdsvYCCWkv
cb9Ldfx2MbWLMLia0v7pP1Jt8bE31jjy9q9lA2fnqbUtzalLWfyFS6uUgFT9GJ7p
hY/KvIFKguZghi5I7YHm7yAP9PsgDLAtpXAITYsfQzaWXlkQg3FUQ/sr13ijEuWl
OlmopyP+YQ5A+fUMEqs7X66xBsEFiuXeqXagDpZgKJFCZoRmgOa3HmgfXf6BV/l6
S5x7uyKJqAuFbnYgfMrluJ212w7y4ikicqZWvnjzlRCTzojhV0TX+juISOUeFvuu
yooWQJC4R2T+DtOdYeweiOQifCyoEyb6K4VIP51z9L9yd5fLlHjdcaH1Vtn7jg0N
xF0K7c9V75gJEwmAxl1Z0Q9eAb36PCdqU+86rg8AnXvklKOxo+ny95FWpvyxPynf
eIVnRY2F11cvKZ7rx1IuHJOvyLsVtjLX9DHlQceR4QbnTUOoK0CxxpgjtNEjntCC
Rnl/slWtnyzjcCpw8qAzHyWU0UZDlQP/noMrUhuWfJ12fTWiXzaJ4iZ2+/FAvJui
Nz4ofarGCrQS2ngHXi6vih59JDBub6lsWw8APrG8MAyNz7/ADjk+3Ve3ZGICXQyp
MRTXwO2G1GtfrdnK31WOFl+uA+rHcInfOPAgYSlibp5YQnxVOT/G0nn2GJZbYlwz
GvaUndBwrHzuByjpsL7f5hQVTqBdePIQzq7YHu6LYRQwCIjqKDqQUFB5rjiA8Z5X
EwFZ0SnkXxEqHVA6M+5ZpRuuIMtPdGDNtKlrR9zGYXcQY9OwstDRGQ4R6JOyhZLS
V948YPM1K8iTffN+6FnvtDk6fxC9g0u4ujZvW0LzPtlu1f9ZWbBcNEVar+cOrPYX
+1GmQtMh0iZAaQAWSzQ2T5MCgq5pNNozBY9xLAuXyRyf0jY/3KAL8UnQEui8DHWC
ODIXG7o9rRbXHfZs94Wvj9lkGZTvOPasKRoxpozCvWG5tzqQOEb9V6p6fl2uB74j
ug479A+FRSg9WUhAtRJlxEdhlI/fJEkL/BWADjmhQ+SIucGtZXgr+Z/UTMAuhA/5
hG9fSMrIxjGMGgBqYl2Dyl2RjnRTSir0wGC+kuSVcK3DGO+nsJdxsVmX6uidNxt5
82dMhdyA/IX+TOExbkjsoE1rKMbn7WC659fxkYFcW1fUxL2bdv2V5XyNHSmcWDSr
W3NPqtb0pAiWHF55YY9oQauWc/c7I7Owx1+cD4gt1AjY9Kij7xV7YGLRnlZ1rIrW
vrHWFRLqsHIJXXmHmpz2IB3QpW652O13CrjXvx4uHKDpCFTiKfZ+fZYCA1nYR6jJ
mcJGF52NY7ZfcwuQ+r7Im+5rlj5PfDjSFHjKkZv0nZpweD4m0iNtranuFcCz0/mS
2RDXjlHyX6lbIqo6aHOwjZtmcEXuXlcnSqvjP1v9Eo7yTIPUI/V7RTcYqS79y7zJ
JFv4toczQFQHQphloX2H3PiPr7oLSTeMixVYHb06XeGrkQmVcXcXBPuoniRVyd8i
+Vb+2UvMijxsBnuGdkzQCh7UoGicFbfHIH3wepqZksL2dVr4vLlCPmRDiuPbOuu+
PoHnLTnFeXvYCaEEnzWCRxIQbzjcZA+7qsCM7nHuiiRSoUMtzmZYPaOC/v/MLI/M
yn6+Y+RoWFtF5qslBZNPmuRnvch1mgJYmM8wRGahYRsWRPomOwFan2FLC903UdAb
9I0q2VvLRZpfDmOthmIWF5H1I8e7DyMSJRATcURw9l6Xj1b3NIc+w+O9yczdxeFL
ZESAZHzA8ieTY7W2kwjX+1GoLR/7LThA15FAvrldmkAK0c7x5o5h0ooZSWuKKXVB
Mas4ZB3FwbkT5rCRvt545ILKEkY0zLBcoXLbvn3O0O4W/E386zB+Yn8wWmFbKwg4
yTPTmGPNesQiYLP7j7hFMOuaSYCNaHT/PEGSDvGgBAx3HesKiSm3WxCuXVJ7CHTn
y1GOgy07hSO0iXzuJ7oFg4mphl63g1ZnOYHQ6YiLoY4qS6PIN21GdQ95ImTEF6Ne
+DgP7Fej//AHfFtdpi9lJAlaUkcC8p5hS1RLqEDO1/cZkEfkbgUx3zj9xpw66seO
1Eh2hItyXexGx/Mg/5KvxtPdvJcWcUQ/pvxXMxBvnZH9G1gwwM7gAjj1dUJzfbNh
iBpmzT2l0OIiZkv9y2veWf7TtMChHh6T/HE96+FCX50wG6o94DsoClJbMQ04sFQP
cEQk9h06seg1NziiOSnwrQ0r1RwgtQvwVER2dwyKsxXsR/+4Jq7yEfb27N6+SZWP
XkBtl1qKswURiqnKYwF5Guprh0001OufbHkINo5B+cV2A1e6ZwKp62YGyPEqfof7
RGwooY4XGtSm8LoACc3ENo/CazcIRkKy6tXMrmiluBTTH4+EUDLZOiceY2Jri28p
UtNNsi94kWqr55Fj9aCyFu4/r57yjXlxOlRlJT9GEIfVNEGBTapeT4DbsWhsyQ1/
1ad99yReAKKhgmWtWonVu7f6AmDcKJENfMA1/cSBAZKz19c/yW6NraRtEI779RMW
bC0O4vlzlC8wqtmiosQcOwzjKUcTTtjlFzTJWWvv3yAmqn3ppb5fGnkivuTd4jgA
Zs5fq2F0ILKfg9Szq6X47AW1XPQJId/Jakz2e3oNdtJdwAAMhCD2eDx22QKrixDd
EYr8jR5Ku4mMTM2vguGg3w5yi+tO75x/Mlkn4K1HN0RRkYhkOsKcdt6Dq3XeOW1B
9tPfmA4UDVW8CMQXBxnuTED4kPJghPSJnxwNireDWqhPzS2dS3JyryZkcCGzAQTc
MzINVYX5rxewXSDt2T58SDzVHkXlqULSbNisbOJlaOli+Faig7v+G/XfgKzVeJKC
vn0z3gd41FI/zvcep3ljjVp8X6s0xtYKNvLB3d342HEw+6Sy/eqYzp879BYhQzxQ
vbIKUcdvuKjNz6r3xrNLxKNlp4VEwTg+1X1CHA3KuICdx5LsR/6A4CZZdVV8bnWw
CVY7QESkD6HffVc+xiDjCiD4CNW1erhVnDPj1zGQzUA/xHSh0FSw/BmVZ6YgSbNe
9EMNGH0nL9SZ2GDtyUC/5uS3MHK96xPI5GzEeFLdCd5ApFt5J7Nb6ui4NrZL+RDo
WVuY5NH41b/ppCh7bHNoYuC7LDynFXpmlXBY3Z9ZarzDtgSHiTMKc2NeY1SSobA1
lI39jfidIXhE5PRx0U2+XNLRgiShiRc1Z+ahZK1R7ZgSGFN/DtNJjPtzzZQk16wR
BUpyRvcxWRcQa7XsfRSeiuOJ5yyoUwEzv6I+TybJr/Bb3+DOmZczBlXKC/DR/dew
fWfKNkuNxIA8L8rfKc2pyueQ+nKwrylmyTo122nHPZFoxzIpuVCZqGMPutrrysVM
xZU9ozgWF0ekbuaxSch/W06bjYj/gJssE69q2gvkD4VtZvldCOk8rNOTY6KtlcN6
jnCiysxeL9qgnuvo/H0yJOxhCNSJrb9OTo50VnUgNHPnuxa+F5o7TyOXAsS6NOL3
nXz+V1Alk2k3yy39xTcoSsU3SwrL/fLRLWhr6oGJN/wwEFla+K+CvbRmblu95kAh
eTl/J1jbpT1ropfCel5ACKzSb0bd1+F6T+boBc5tB/9/J983ysjRChZCv6EBWnmE
AsI7F2W+SwUVJO0+85Gy2ANQrWUe6WZ9xQgJl+T/suNhldOUo2qLEo3R1N5LaX7r
+BPLjCqhuW9hGnWLEGDRouQTkUzOrYgTUa+X4FmsOcXGeca7YraifAbE8hantASr
1NMifXUf/G9h7pyrq2K3DpMrxVhHJwKV4QWIlYoC+9KuVQpQutQigulg0ewBLrqQ
GFAncCH7LJsTLC0BTjc2UWodU4gTaY3SecV0WKbk26hqAQ1dU+cZ9H+u9ZslGtNB
CR9ntJ6bIhR2wyKbDcrWikjGE7qzEjeVzVHcNny643zowCz1cU5w6fv3VO1qRgDA
7X7uQQdWPBTDCrKk/tq/NjrCnhkenw6dhuFm/dAYSZyg9DrYTbaBC2ApWUDnAGaR
GQHfjXB3VnvdeFG6hJXq4NDgl/zw5XnRRXTiSy99McbRcn9i2LynEv69dOocyb6Z
6/AwGwguq6k5+G+9aAToxBj6UmTUSqyoqTzmAQSuJi4IiCq93Y2nF8db0/wRWT2V
ziLPJVfRS/+ZphsAa2N2j7MEQ30yv5hIzxvTn+g3K9/wAa0k+vRfW2sgI3/NLkq8
pkvI+Dqy28r+xyVe337ea0MusWHKowrVabgRIQrkvW+bG4vK5UU4PXmnbCJpOqZt
GKEKQQtd3hfYSdg8xLRKjXxhC3nwfvdGaYaZ4/7I1xQuD0Klhs+THao4/U+s0LgB
Bvwvq2/ap7KBGtfldkdAtSm6WVZlDx3/G+2/KwhblMUc+e7ZmFBzIB8E2Zvu9tDx
Pii39L+vJ4/v/LjcM25PGgWv+zCyZaMns25jkxredIQObH0NRZGplXVjYPlwTVg8
VN43vBH3S0wPLZcqg3Nc8Za1vsBui8fFAfKoZMYTYub4Pdspx1wHiNqZPsX5L9dm
CXfvc6BrnLZxNT8swkKKvuZOe09tuL0ipLudlAp4EdPSU+LJFlr4Y6YsPqJEpSVG
Sq1Dn4pof5r4GfHnIqBTkZ2OWA3kiRCQNxzwAg0+DJKxVbP9af4wJSN2eVZqyVXL
azbbuk4hNRhCnDETfCDtlSI/SOOm0OaZU64MWTdRCCUWPiug5c1OAjTCe8//F5iO
rZK2f0Z2b26R5S1fw0FyjS3wPIv44JP/UygZLZhywjduF6XuLYib2+tNpSl5YSko
cpwGtV+AkMn6zvjVKHzCJrPyuvvOY/E1kssiyO2MBrwVo38NIgA/nywVbolTGqDR
mRdLybV5pM7snGd7bVq+vOSkaqrmuNy+z5cpOMczjA1RTtAYi5UxpU/QQWtfJYfy
QOYY7cpMbp9l44wj2Azd+c4jNLiq9otNa7kOGkHrhwVwI2z+7okylonZFteCiiEH
nDL1Xzen/y/Myfu9ZpWviAWl8Q4qZ32JYtfzZrSvM7SwunsED0/cbbbjerJI7m1L
8kxb1GrDssUMv9LIentspxmk2KD1j5xXIUZAN9lLLek1RHgBzQNaBzyrp/U2+GJ1
GlMtolsPunZ3Ryh0Qj1s8bOW9pkd3cRAvaHLsF3raKrV6cUOPx1S9izabDL28CVz
cWx6tlUE042vzKvouoeBF4qfJEhjcvFLyvXeERWYubJAOLvbmMIGO6WM/NpcQEEk
T0Li27yjnjpXqee9XGBU+S29yz9Oi38mK309HniMdAUl16GA44MWKAeg9DluD2W4
oaiqx1IPSv31DNVzVKXLUgm1ouvX+usI35SP0OoTw2NQna/nz7guHONFfugdpCC5
RrH+TLDItj8rNm/twf7h9stF8StDAaQOqq9mGLNRubct0Guc4o920vUhkqXQ/kU5
XPNhaE7t/aENcYTpo+ZF/aipAYRtX7/GKxO0td37mtd65R/AYTfwMMId7DpVO4ur
6NXkJHj57aYNnVMl4KxfRTzObrqGP/XovlC9VgmzY9RFXV56u83QQJ4aWsIwYJc5
qryOT+f1ZAsLlAyCzoAhZb9HQMSa92yT7Sv038ugUq6rOOnlLgQ4DsSg0WdXtlPM
Gq/WK96glFftnG1i85P9jj9nh09IGXFScPNl6EKsB8jL5UZU+rL/32BOXAqtps3A
6WMGlqHQ2iozspWLfaJ32czWes1RyAs+P1geyj6Vr8S/wzqn4AcXeEHrAz+HxoQM
9rrIMavwIMxAkDTTmDONwdFexVp1+egYoV3fvrh8xrQE51PN6ad40euK1ocip9Xz
glvEbX5ZUjKdYdxsOCUOYfA38P/UTFj3B8c6shS1cbGrjzkDisOfQAP41mqXUvG3
Jr1TDljFSD3wjmJucXi5aCoc74Rv8QL++yRcl/g0MsvznhFxO2cC2Q3fZmkZtQIz
RweDG3fKCKRkvpv6KMTyELO0YTc3k/1kIWEofXQKDrH9qO9kRB/y6yGTromZvAxc
Vq+WflmHGmoEGSoEZ4RfVmwGbxPeJOvRuUHpupxeTo+KXKOTHhz6Ja/C0tORzD7l
QS5UBO79OlwtU0ZKkjJ1zFNmTkueiFO2rrQ4E/TKCxHjkigT6NM1gIwc2wXPObAU
SBMnp/1oiSGV8GuBL2M2FgrAv+Oma5DDFM0GZdExEaMoalL3yJJF+tfxPvHvXP/O
By0JWWVItO0Xy2x0AG4j6DruvLlZ2AQmZXKVQtyjw3Wd0IrEr4T/sx1bpBzgQeIg
BljtVqB5960CaKQ/tczCmn3EFPllExUrzvFQfiWh0TuG9aAvI8tLCPWDZ2Nnctk1
Bmw2i1S57L8lug+c1A9XSFxmT6z4+7vV21bjDX9zZbmKzezpoWgWmUYiWTn4Ez8d
xKSh3BsJ7qPuLnu8rXyERiENf6cLskiuxbam98HUCpLT55ZfYMw4DM5dNqeKcouB
UZFjzR1b4YB2GSeRZhHb4BFlH8EtjHA13VaBYAmxy4Lea4bfOQmSTEVbKjS2jh6P
SVv7hlwf0IssHM8uUzAGR5AsZTxIz4pTlM3Qpsla0SRRqiRhGXsyXVkHbGzq2Zx/
fa7yjyZxi4GOrZgDU62oBwzIeiNfo8acKLSBbVVYObY93+wZwNarLazJOwA71e/O
HulTvv/2FcKWIMqJxDNAMp6fnWf0OkSXPmBH5R/GmnAXqPNxs25rP6zL85FrfiEg
QkVmnAYa31wy1uN8Q+YY/gaUjtWdVUAIRDAp7PqUMlozsQ05gDRs7Tr23VG+8MCw
7TTWyUkchreLtgn+6OoXJhM84tGiWy67rFmYme/L9mljtzbdYXgIWpcmV3Bbqwr6
igYVVs64TlUu9Y0aOS2MFoijNmwOgvLDVQFVu/c59Cgr+QLPadZ0UvLV7/uJRzb4
VBB4ZXQAPCLuYH7WCy1HpNWW80XnoMxCq4387t1Ru/5rmITn6Uc60suvwNLIQokM
6fqMn4o2NxR9j0LLZMRyGCOPLZLCwkcOM8kYPxHah9GT0vm2AA3mx1r+g21+8PeJ
JQE4LhfJI/n2ejHfr0OqPG1IC4CzbArgKQI7LsODlLKM3DF/oV0ojgpXSNujJCOJ
+ii/+JzO7GTnGlp+CEo5YamHNeeZYMopK1NR2dCMkBNDp892NiNDsaEzgycK5NqX
DcCzPpyQPcl+ehxxEskO58YhhLAp1hAIO9yZrDraPDwu9/DjQ8PfMddTBfY4fs7f
o2Ve2Iqwh9FlcCE5xbhY5igwrAsWJ9c5kzea9/jeX5YsinfOPnMJD6tyFOh3uAYU
u8kTrotZQs/D3qgCBWxQxtC2pVSGxYdBvO1dWuemh4WkfSibrTEbiGydM8fqJFDZ
p7yfjUmdPxZvWqJXMQZTV7CrI3yj1mz08Ot4pKvVgPm33AIhOR9Xr6Q1k3UDwqc1
TWIvNo7M/4eIFU5U26Pq3ySUYAzr7Y5B0qdHtRxRJiWhkidFBK2eXTNYlfOS+YhO
AX6dWBMhcV1BFxQbHMvGhgGiNXvuptZWXk2Tj8EoY9BP1ZXVXHtCzEKBN2lQ1sti
T/EGpSjdqjnAHiZsrIAjVYh1UL0D3bGmPolnGy5cOl2NiGAZFhYwVHkeZ0tPwwvx
J/OG8qX2p8wiR7XYIY8kQLbhh35PdlQP3p+KHqVDqEyFN7zER2mE3fyz768HL8GK
dnZ53gJ/RaRGuOd1NnyUgSlC7lCoRC5QA6optrNvt9FdhzwPw8QCKDiP9BkNEE2E
u8IFNC4Wk5OqoQvohcG6sUltyY3jdkWZ8Gjme/ckzCdd2ITdJmFRh2MCBPSDX2eV
7j+IDmO9hupiXP8m2e/Gz9iovSitNRSCzYUdcBQEWAEo2iMpw+HEM6nHjYOCcSKb
Yb3eVIXi4VTe5wZTxzYZM1/JTePeVc5sWVzU7AMbrly2fQLUaEl8vO7oz9mt17QN
Gb9SCQJlk5gP9Mn7TPDBY7rxskVw4ST1i+oDy09DoOeHYj/VXtbYJeET0ilZD0ls
jnNfXIgqWwlR6Y6LinrB9ujE69qiwBh18qBiBjR1UX2brz/Yatb6OwPVzHO+q7B3
O37+v/McKLQe9XRLlRx0VO8/FC3aUW4TSRM0woAI8d4q0s/LO289ETy/awEi+uMD
gdak+7zGuIOcoh0tgXhG2t5iHP/r69RRkSa3x6TMbQYt+srjjTP6sgtDd+TKBjXP
X7JT34AfBjfyr58Lqug3zyIrSt3j2Fz3E9dTb5BXmQiArxDsEaUCGyvOiDK9iIzO
4bAaZVXDzSSGiqDJgpXZxNRfHIl0yvVOS6jojQ9DEKMoFPgV3c+sBKytvR3Jmdp7
vubT6i0r+4nvrQGwGtpvUZDqM1ut65JVpGoo4xD2foNulbqLzIOJPWxkEobJlJFb
dAc2n1GAWZfG9PVkWdnJJ7N6jI5Xxf07AMtpk8bL8CJedXSWVMb3LW+kzW+UqI/R
3HpCH8lMC4p7pertXos7GDmYne9rv59vv94BIjQQ4khm8ae2TfV1Mypcf2QWVl5y
6xYLeUXxDPuwD9mku8Sy1Tv/7GOilLuYuc5H55+GSDuuC6wVTXDi4H1cf7R5Xz7h
pYwqzLoEEGks7QyLqsCKsAskMCqo1HKlkiASc1cIn12FGT9hueero9UytxZYbjez
QskfueVo3mde+DcmMXntXP7fAolPHjS2Zl4mReVJsnfnQkfcDJnf1dh/wkxI61Hn
U11PpbC3f2XSe+N3+5oLhQ1PsNXwoUvHWY5yQxE9IpZNKu2usgZI6AihmKIsAvVC
CM2O8Sxtv/6jU06go2kUEcYyT3yFz94878yYGJkvXmAOGrO6F+Hav6ntogM5ecvy
L5cXxT6Xa2hNXn2jSnns7xtpf4rHINaZHLpxy/E00AEG72C4N7XRIr06Jt2q1+DY
SFC6R71VC3SQn97vFX1+7FAl5bwRe3UiJj3Lt12/6Zum/BhBP5AZbZ9marh1X5vU
vnKPbQuz/mfotr8gF07dYMnJLq0mCIzaPRTjaa8Axkmolol/NtEfAZGz4ivVnyXt
00WVEq5JDSHaeUFrUrRuEvPSCPRLe3+smkjijIO/MH2nNvV3YOiZq43PwPJnl107
7ImhpfpyCF3YeDf6AMzS+39IiOXRkdFWMYxhTLNpIBDvqY68YNunYQz5aug775P3
i8TinI2+faYYUePtSVEZvp5NyOhgLP+ixyrpPMSIvRp2ZPRm36rkB38H+fO3/T9z
0y9xRnadh4T6g7UtAUTgzyuQ/f0gBQ+2Nqfy8+toQirWmzqQ9QmqSPYq0/5TZ6ce
Xy8xUh3sKMgr6QqJbO89haQ6J8QFMk1XBHk43h19nnuo/rDKBdvbgyFqtgiKzVJC
om+c5XLfFjqP2ZReqpKNzIrBkkDecMzR3C8GsOJyWSS/SHrs+1GzY8NrfnBozGia
uRi2GMpBwPJ7evXsJ1tVJtHGZzPSXtDp7m53FOFwPTpxi4dyV8PLhrF1nsQGT6F6
NGCLkhlEcJBsTQfnOGt23XH27/sTh0WRIuf6vS7UI/EeT6kpdtEjENN+WMDvKmGB
ylgDdrtw2kxkm9lRV+Y6oMJ1kCASDISXrv+HFfdNEw3RnuiSPR/Syv/TqeYCLetk
YsmOpyuJMNgf45VmRuuTW8u0vSWDkWiYyNgmmyFcN09vZ2pgfYSgBfccOq9vtnB7
+Wo3zHc1B/rusivNwRckax36wP3DEpeP5Pi0eENpPFUaF+IxvRrNMwezFQP9KM6Y
ValMnv0rATwRPSt+w2V9hnRQowV6V0BppqiDJCX69lXeoNMpctJb2ygjkN4szSYq
6tvQPh8epZP66t5Ym2TN/BsMGvlLdUWxVfjvdVPSbYNhew+i+CmBF6ZMKaZDxyPU
YK/c9R8QXWZqzvKpRX+Dq2viQFF0aoh/cxGDT6Ae3qMvfxgIR/NbqaoYVGwfkM98
HNhf1eU4SKhK0LmjdAjGtDFyEfgMyR3Op2OMC5sZTFtv+Uc+0+Ts8rTQYT8LI2xA
VvP9D6UBvC0nrHoCboU0+ly95YYTQ38dd0ttxQb1ogJyo3raZbgcNoWf2u5dngwQ
ypCpAztpCkarAJE+p3JpOahHtNeH9Ofcr2174vWBtNe4Cxc6Ifk4HTTi4+lsOx51
6zwBJmWFdcS6E8GrioHCjWabfb86ALnUVZNhoShka/x7iu7hPEU+cJhPc0Ei2gNz
3y9lz2vUWMqUeNaPVzcjDKirdmZQjkN2rRZEf2R8ckHPQ1Z6fCYyLmTz90/6VwCI
RRLldqEn7jmSq0D6B7AyYVZ6AzjG7QUG8hF3YY92seUl68eorYjDpcr9hqGDL2Bg
8oCrXioA3Xp0+TNB2y2seBdEhzy8KSTcRs8fbNKjkwCdpE+dIVZY6UUsu0yKmT+H
KP1VurSnnjVhd7Kgvx1DL9vBPJ4rF5QBCf+q/SBjnUOj21nUw0tABNghSxIukWUe
h0ujXWuzokfI9HXoGnb6znrf0wOg6FNfIY0ygYLGqeCjRwuI1k5FVjAIZUtVpIxl
JDRaTPcBGjHGkgfvDIAR/EbhUO6qzhWbWpm/pTM+xMGC6+OFsSyALwKVdou2Rr+E
geU/f3pbH8xNI2HN8WGccQOGG5MdTkZN/WO+jUcOYgS0cvgQTGr3FfMSaMuka+Ct
qJ/97jp8xhw0gfF1iSqm9fczexPbnmXF55U4A/WnExeEG9U7aMvrSHgEQXzDepo3
yrK0+jnZXud0DzT16OGA9TuqfD0maRIrvOO/ue443rLIfVi8hSYjquGT7zs+ffIH
6v0/+F0VhFr9KtySVvW5EnQOK1YaAIGQMP5z1u5tw9LXvcMN/flAVJ0lYaf4OIPU
zRIpypTbBSceg+rR20+tNx76zs1AmwFRxpaSfujzTTg65mY3ezjZTaKrzHGIQ0PW
E68u61cnXSvNu2xQ4+vsmBzu4qTYa3H9fiGRvDm9FjOAH20FfkAvDKxBkJwec5tv
ux8rJuqCkG71RToT1wuIlkfVCPVkkQ3sx2Uk3iFodnvjIvBMQqf6BcwUwTkrk4yl
u+JJ2d7JtgjTZRL5ofdqClc+Ng//SIyYODuZveg4YtaqLFQFD6k42obimXxN7uYi
6mNrsaMMPoEhA5rdTwY7c8yVIVJFhfbS66BfbEO9YXug9kc91v63AeCQ31XbFXR9
Qu2/W2nPIJhvwHdzkdoqI3+Bawt7gOq40kHkPfzXl6hF3J0umWN9dgmBW3ziK+Xh
Q2BwtaWS9zAWDyuq3Jp5x7QhD7KGX5EAsnvKZgit5gUWz8KB1amWbsoqTdS4zlQH
Fj0k6DWAelszDrU263UGcyryqxTZ7Ip8krMSqt7mHXodkv9wR9g1I52e66A7y/FE
uHPiyCPFolcWvhQOZ+ztvkeN4MCdajP3PLX9oZqJpKFRG1EdGzO1y0fdWC42nIUv
k7w+G5Cv4FqQRSuEcSPcoeWimJ3jYeoScCqeoL6yHhrbReMC6Jj77mrNjUHjh4T2
vz4frYNQYbr0VgeIhRbxzJMfWourTer/82404Qm7x2/+HB2jjr6OkhyTOYPkaic9
mXx47SrRZiSy2dg7bEyJfLqOailFeFmUh95AyrUWn1C+JkTFSIPayseZGYEcXA75
rZ63r/gSmQqcGgpXBZuN16b3WxJaWp5U6rSMaXb8/0i4+SaJJTJ7wV/UwxXSN3L7
Z8drXdlHWdKzWxDFtEhNcq/u+0hSAWZv4iSQyn+EkOiNjo1RB/oohX9IXuNG20E/
y7BKhgoDpmllpVi2ytu9qf/VcjsjQnjJXtXGFfRkaLvVrS83OOOh1hsf4mN1C7QM
7uU+HIEJ0HUBrPaaWeRQJ8l8iojXh3nF80WWv60/pzsSqwwm4vATftjQlMkK3/B4
Sh9/Ba862FH54NrMEzad++4vXF3GJQowvrW/b73FBck/uhZE0vKy3ltcaehZaqiP
X6R9VuzqRaa1CzOzLu3FPN0xVd4X0HgqmN11xd6RCUZY80yB7nPMVeXoBbuzgDNL
qRSs9JHCkaYse246Ftl2qByt5qHnRyB0TJkr9wCYSRr32LxhN90DoSQOXNic0sxq
O8at9+oyX6BHMm/5wGwQ2i53USgzxsT/LX2Kzc+n9ZbVOY7r9ZA5FQUByfOk878Z
iuiDOv0KOk6XK2XgyjwQzDpaTvkhtJYwg7m0Ohp76grxWWCQQxLNiLfidYo7MG2w
NlnZqQzO4+iTJrT6WGlAHS9Ut3DbJSR7whkYQ/ZkfvBWfDVIXTrJ7MAE56WEyVF7
0pzmwcJOT6rz0I67/u9tHAlZJzC9kbIxY1dyTqTrSHBD4tgusBRGd2D59fdrsBJF
na9HlLgRYneQ5OCKq1Aik+4T9q+0dMMIU3BnK9FXse9XKwsJYVt0d+EBcisM2A/C
dgxC8oknFUimwI+mRhdCp60hF6xFBWsmp5S2I6TI8S3wwsATIA/gZJm3Ek++AfvH
K7b5hlyfAVmIeVzNyEp5W0ud5Kumf7OHMbyqNBNvemZ1d620fZjLz+rdEoi0UPi6
iAJYqTCj73LKjCKg9VNkNTCaPBzs1Hoq3HkjACQwV9U0neUVSWvJUX7a89Zjg55+
6KMMS36QySpXV5xlVvSBlvAF/SxsaPwU1gKQQjWvZGY6Zwm92qcjd1QkOfGCRlgs
HJ9XzrUSPaHBoFIQAiv7+nw4kYfcFm786WYnxrlffzKLlbIcUeL8qu87J+ZlG1Wh
UsRW0hDi9viC3Q4ghY7/a7809x65HhK6+K3ptopSyWx8QvBWpD1fX4P2r7FINl+9
bFnSnmmzl+75vkkPXtIFN3nSmxdB4pRVqwSYa+/rvDYtU+OSKgc5QSraxl1jgmHH
JX+vleaiwwyoR4KJAdzYb43d5N1WUwn8bbLxrLr/epech5inEuxELkzwJFjy7HUG
L6VVNjUrvy1ugj9Ccb6/AYWdYR3HtthVR/8eJ/rLvK+1COQSjxqnRCOitgm2lMDO
JKHiWT8127Jhpb3TqueLmCUdA0oKSTWulnEaTzAd4CH5zsdOrT4MnRrR+SUgo3+T
g+Yw056J5mKxauGBDWsiarEFJTILy3R4BXBqf9goi9gUquMPKheDiVEWfb12dwEi
Fy0X4o4py/xqZHnVhI5p5OIx2bLmB9+yc/WaR982Er3VxYUd/Lu/5vqPgyT8xtqj
iH8xmAQUF+p33rzw4/m7iYKBn3mwgnQ2xLvL/oXlqJyn5z/NWq7fMeHTIIxaWKnu
Wf4A+v7H98ljtATgByeEPL/UJ8/rlltyw3JLPSVkuORptGs67RuEi5EugpppMU8P
+f9CDF34fgPDQJyHerNDm1UihWtJmDq7EvGrXlsJRrKHsuVStC/WQegrhMTnImbh
T96UxXPHHy7PV59u8zhGy9NCEwNEXJXE2Z/iQs/7NDD/djDRbDdfdT9fZaBk/kUK
qZZLf7sQejX1sQbsy5T0CSw+T/nyH/2XOuBLFvr0jAduiUL2sDDdtrdxppvnnlCb
0HOF0qMRLfl8fPvGe3vN3YzO4H/+pUZy+Z8vq70SPTU5CnPTeNwvZ7dfju6UdO9N
7R+0S81piAsytAjGkI60ZIW6QmKgXwu9Id0tY/QFebnrGqwi/gCBDaEj1SBisZhv
OkW9Ca5vXNrHpccnS/jbTOgBcGyFxT3KSQpeCmw5j/wir0wAhJIuX5JivLTHkRwi
O3jZET/aadJ4FJr+OXV92sICEP8v4u45tgyIeA6CABqjwicrb6KPDXgcE44K8CHq
2m65OF2p7e+RUX3QAGzdXg+U8mxFroKQqMCaILp4JhidEA8FxbTYw8XhlIoJBmP7
PS4SfhgAwZUHSdE3gDghqcL+mRksc4E89MEQbxRXzI5dD7/SctiOFybgtJh4LpoP
TsJFmf/F3+gYf7gbdjCQrPn+s3HYpLBckdBJQMWldNGDdhIbCoAEtZlBQ7eU/xoC
n8O1z7GOm1a56tjarrJhX8Dp7B+57K5j10w+fQ6+kkZhUIWdl58YhJX1Rf24Bq+5
3cHl1FK4TPWJ655LxT61PSjRik8iIo6YZrsBJNEd9Q+vtb8YOEya+2e9fJ5v0pfQ
4Fy7Tk8h2OikS9mehvgZ2GCeg3vLXuBEGgPDlCioCJW+5WXV0md9yiyt3yvsxgs9
bzWh8POLhV8n70ct64FzWPQ6Ay2KaAsU3d2Kp4GffgUYDH8AVJ0QQfaH2Hu9a2RN
KmtVEsruy8JmtJmpyfkuapvv30hzrm592aGfxGTjBU/ks2Yi9QTels+Pm5uRZRpM
ALak2ZCKG7a89MBw6tl+u0/cut9yvddEs6j3jX5GcQsHHGH5tzaywnIvThaT3kTn
GsOY05B2AajA+GEgg8gsvr09aLnCQ9a4qkqn5YtYqhrqrbmIOWbrk/7+S1vnGiGh
1o6e6GJbBHQ2aEAxP3x1lAibsVjzuh/SQOH+qBxBzR/K7JMNc49BnGeliX7eRWO7
VC6NDrMPdDPlFkLZhPc7ZRiLffdFL552ztm/FqFazPHyzHA3MkVitE3vuLob+K0y
e4/9B44KrwyKppeopOKN9r1H41aOegQ02twAob0NwkIK8nnXm1XuRh6eeob8GuNX
wqMaE0r3NlL++Dss8NCsU0ApaHb1/8JHLTeKow8dEcYfn8UULRf7ISL6fCRq37nz
swP4tVzdn0o5cFIZyBPmo3oHZAc07O01NuWNeCOJSijtHyEIPC1WxCHXZh4usWqs
YcHVeaTZoWqWTrsiPYEAg/6BSRNwYtMNKVAx4JqrHYEuF0JkGH9fWtxQbvbDhBPK
0Gdk2V8oD5B0Ly3G4ueZwV2SxjI/Z1Z+yr8g7VtvoVSXRCkqFHGYDUCGxPgic0Gs
GTKd6pbHHGdiWc6KU3QLDED/vIE3R02fKQxzatibZ18EY/oArricHohIHueoJWi4
7p1pT9KiIYoa6fH30vX2BGsnQWykreaIKayCgoaFO6vPivQPwP2M/7f36iTyU6tu
XaXZzRWOTexWYjoKkKPCy8Ix726bNqs89QXcuD7QVzhU1ml9cakQCgGIoZVelErB
iCPMfsgc/wBW5OG+mLm/efxpzBgHONHGML6mWIKytBEtzgunlwCe/WGq2Jxw/VHK
oPV9zmBfZ+VuvVXBZhLra6PY+wSgzLxTDL+iEeCf2S3C/GKmF3RZ1PMk4QzDDPey
1ZdgIxslyo2gBlv+p9DqrSrAKQKuF0fv1/4oOuweaiW/bBU26QsUFhvHpVesIPKf
aKzA2qOkyft3Y3k8uTMQYnJ6H7/uvYiTYTJdrPx+1u5ISEkzHNnWd5/lRHj53BSF
MFi3GRsf4SsPlwB4ojNP9NB71Az8+CmJPZoro6idPSz4cnvRXbW1VMnzb1vTlkfH
QbpyHGjnIVtz77/yfvmix8jIGtzrmylsH6xehlntVHkhvKsKzal9EYsP7VJDCvwX
nozS9xLONwXftySCMl+pYLddvWx7HLxJD05xQRxw5a20OkmzlSZTnmYX6Yz86GKN
qmZs48AJVdH1To8q95mShCY/5EvGZM2IUwv5VPYFeokct2d4wsGbD23GkDd4Mv/B
oiqgidqxm7cBr1Fp2jkyx0eHFQjOVOUKo3silgTRPxy+q8tQi+hl79sNA5rBNF9V
BfVfQBIZMxIy4PSeLEL/4pSDRBKJHgKM4cvEA1ukiIp+bs5IxTF5ZBELDEESii7R
4q8552EedaXthdLxTuvwOWa8lWUes2FO09rRXutXvZgK997pL7JfIOfvIczVZuBh
kLTNm2uwNUzo/cYQeTZmyRtlvZ7hGB1+qeEJDJ5LRqo/9izWVbkg2dTIZrmrcLkq
Eh8I2F6SHjGC5z5ZjlQ3P9HdAx6mPhpN8wuc0vQZTUQ9/bV6qn8z/s5RLqf3vU1U
o7dEW3Hs71tO2Ka/vuOvhsqXrKfW2f4idfMeH1XjNaQQNBh7LG7FXPJQlr4n8pCd
J5u04wZhNDpR2OzGYoM19RJFPBugjhD7e1kQq3/Ae4Y5W7+Q445vZK7hXQyjWt91
nd/bkRPTTnetsqx8NWR+8+QaAR8SP/7aO/m1zr71vLZdI+dZRuIfe4/ouqb3S/hF
DQ4fK2Wof3EpdbHfP581cvrS/3DVuMSfVh4F3XR5YZQXR0pJCTytTdgnWHNe3Iac
c5Kh6k0Ripnwyx6hSkfjyMsDT5hNkm1xWaawcZJXx7i+b6iCV6Zl8E/CLLCnCF9w
rrNnFMd507xrsJjk/Ei+7osAjkkBadI2dQnpYV+c7qZhF9iD/wdaVNxqHTxeUx2v
AnLpi1a79VY5psffUBm6tZhiFwiZMbQOgfG/BqAjxer7pHq9UuRByZV4pmTCiMY+
Ro87lhxBNmDSC++C53BxYa743iziozaBDlZ+aNb4LoLCx8vPojl07UQn7M8s9diu
YkeawNHhZdqMaOUUm4ZCKlVbVpe4y97ifV6qH3LfhJJ7ok1K6O9weiOj2epFLX9e
ee5nnb00vsmNBJ08o/26lYk+3S3I8P22/SuW7ZAmiGymN8/LZB7x7zubevWQWmfU
F6D3AzMV00t6nqyVW6tcAruK3pmV79OOu0QpL5lMl08nFOnuEfEn8UA0vx/NOM5q
GdQFkAKaAKyT3FKj54Ob/ywEW2dvNq956W6XV6I3k88HkKJSkF3JRgJGZ6X+e/cg
+hOfhg+YP1RnecHExOGAYnUYqfjU88dH2VCLvBNberUv7Is30F+nB7+aKB0zRCAd
Aaqr3oumamp9GdKRxpDyjGdwh6OVTnyNIauyX+16xSoPaxJkD2doAW1M0aKQIFHW
yjgyfGl74IKXiwfG435Xlm0bKCUqO1aLXJenhEpI8ym5xPVhGnoHdXLDj6KKyHuy
S3+NF7r+EOIZzoG1PCwuaF8FYY45nmDp+AgNpvfFgWEbo7zS/Vjzjqd3s/NzKJjF
slm8v1EUinch0JmEBa4Dhxnc1nQN30gH0a3Zjna8hNyfRuWEe9HJBD6xnKwOeePS
pSUTiGWbX0m6SMK/znErATpifp7lqXRqwW4dQKthEEBdNRqaAVURcA03WtTel9ZS
uGBl/0QLt22mT9WA30CMT3nT1g0whw/F61Il12t0hnh7VVt9pgdlsX5+Vgw/ycDx
mSOgPGANdx3F7Ii1UABYy3diXtxCqjusSkE+MdIKSGoV/r2LM2+pcosSzLDhkrYj
t0PDJ3thq6hYoFVGvg560BJEpIrAYQsZUdqdTNdcMDXWrMKzrLaYV1oDfpefkHL+
w0neNgZ7v2jfsrUdQTUNr8m0MDXDiX8dL+ZkkAuaZ8KdaC5RoOl6zTDpzNC77/c4
pE4AQddqhB39IQBvC4qaMD+A1GcLnc2x30wtwyExRbY7+q4ByzpjVCbiIWbGRZHj
ufALyKQaSa2JZLQnw43trfIALLOOGmZuHya1I06AxFKowpX/INsFb24HW4j6EFYM
+v+9nG77bS/WL5ujOgqTCGHzzzzYffIAXQRjiNy1t5CXR5vkkx/y16svgeU/QdEL
cDK+rI6rcu/wxBo8rtltZ3ltWmXYXdPeEazc9WLeBGosQGWDAzxlWsNeecgv4CUs
gg0qBSBQuGheP6MRGqEz+g8HjPsHqNX6NuQuCuIUuh1/62ipNgtDY2+njT0V3iKJ
1jqZUo2U6+JVkpicSAQ9jyqrxuucN0wHzDqEBCepUYmdtVW1qZdX9h+1JplYmM2N
ks6KMVQcK02f2tWUhtvfPQvs+Ba7StQQRO6GibgoVzfWbISsgx5caqip8vU2W9iw
VafU2F7VZFZZQbIHy9AcCjlAwYlGIMQiPp2zNij9kCvQ++zW/ySEIo+mEoawaDbd
BAWZqZTXs42rSbAo0l1YDXueCMSJxJOJV8mV+7vqLvlM5ul7psx2GeDewI3tVvcd
8knnhjKsCm5Ak9a/7/2xEPJbC/5E2wUI8qQBs6hvdBR6UpuvSEYJF6uspNtDO6Tm
Pr0+42U1t0QiFQjh/jOsXpV3kgmCRbepfp99iwj/V/XmxFbzJ7xS32kFFbd7rlJL
HDy0Wq6vrJb/gprabhYKQO2mmsEdBuFqHSDmEOAMEmt0mfsWzrVnNEwtdxAnZd19
vG2+F58FWCE3Yf/BtKpezV3zXLoOTz95NWF6QFZOOoTxDc6tvxsPUg1pvDEkKhX0
oJyGt7ThR1C4R0iLda/KGGKeA6AZi5D0OtAu3/fbz5M7YY9fPJt5hK+vEI1NAzo7
RrKlIqj0rQINd8m1zpavVk8N1Re0zHT5MEeQp3/gYFFosIdLyuqd3HRf5ncB2Lk6
gWd3xbmzmswEhnu/2zLn/4X9vo9dSrzxXyYAmKv2w1hS6XpooutujuTERl++zEcF
DqmrbykPxRtQcEn53rEsDAcZr5W120S0TDzQdANMuBNflHTZYDZlYIsklKDqI+Aq
+eb+UQ+O6q3EFqKWA5jfRrbEQMCmaSSaSzqVaHErNxt4FXHpxftVgMt3UcyJSVsL
J8no4aYezdtpEXkEUAiw43sGY/KpejB/hx47P81+0ruYYrvgEDw0PDqClnzl+6Pm
RRhNwsA+5zt3f8S7KlRgNVuqTQIZfTGZzd7gY/GUq5gmB/p/NkZPWt8Va+5rYaaH
6OlVqXhFEijkMTfay7plrUweGFCsJOeFVM8+NabpXBcR7OMXqUT9rYqAnQ1YkLJ9
7mPuHwzEFQWiySthsCqAGgHPfOToSDzjvLTHMZz9Tddd9GQhlRPEV/Bmh0kfcBO6
8rTjvMTjArSV5oS1h42N1+QxuHqLYwUpizBIwlHb8LzuTgAgznEPnT1fObyitAYI
qO5yZjBGSD2X4R8v4QA3Mb760o/EW08x56Yr6Y/V4EoX7TCURNDRPYz1VcGGcO8+
4UbSmQFUyQuSaZ6BWybIDpYE67YCz+3/VNH2fZ9HKGmEZFZlTYTmzkDbywqFJHI0
CbypYIfSV4mBvN3PK/X/X576j8ylAesEuJmOAdQvnhkqYu6EOnCfVl/gUQZu4oc2
9/7eanfe0KUuOdnwUOqgX/bkFHwQfS2dAkpklATfplbn1JKheA3e3dkpMH/XmE/u
J9731gtMqohLhJGmGpTBK3hBmhSYdFnAebDQyFB0VNNBWQSIixqDhbm5PWhYgl9Q
tp6XJDjNEyDAXi+eMfQ799VU74ciJX0pRGAtICvGu54MFRQsJjaTXYv+hl4L2SgC
I4TkpGAYpeEExi1ijydbBR9Tq/kBUW7+JrxVIWBsQN4ML8jpUP1XnsAToGUc7J8c
pBmxmLGhI4n0tCKyv9gypMu+DX0GJ7eWZu1Qx4jRiIwZJsp53Bye0BAxzqFye3ch
4c/JHNw/IWlMXiCbFzQcbD99YAmgTOGJuhKyJgi6gX0b/PB9RR2b1XahQ0SNg/vc
e37zX2IO9uR/3cCKXSpD8Nu4HYqoXRbI+fPIqQExGLZV/8g53ebPf1lR3o+uEs4V
eGtNOZibv47SRf9iIqW5XXVUtjNcGv3zgY85wkTfr5btck0yCXb3zKiGfE490FqB
sqXNdDriBR6fxjGshn84BLafcWc+mlB4I43vxEH6EMlFV6VIjLFxvgoFy4bBFxoX
sPVfP9129JsBBL0HEjVnCyL2tGLcyVmj6mzUIxgxJldG28Tf+Xr7t8UA4VInyFDj
jOE5Itn7Q5dwDcKPacY+JnKmNC6nxRbws2vc6d/bF5nyyXyVUls/bEBCza2n5gUc
J3nTZUNVDXUCQs8KvYnhq+2vzjTQ++yeyN1vty+qb4Z4NnPpiFnaQUpAtTF/MFBL
N1k+DMLyvWMe9eXUv2spiyV0WWIEknGgFlpUV/2LTu5WACJpvp8rLRwTI5neiA6J
R+8ANar5iEqq+TYWdtF888qINuK6cZK2Ih0EUoIVL62JTBlTyPQmdkdSA7tzGKIW
GSUKdK5dEFeCoKw6zeb+WRYrC3uT6jqFQGpRbXQ6yhA1e69satJT0XR0ral/Leei
Q30UZF1tkW5E3S9pC8X+OFt6ucOgB/wKcIWwHy00QZAjM0uYJfx5udMELD3x2Q/F
/R60FV44Za6Tkna2PxXjTTyO1krecpqN/7ksCXVPbZ4K3CakHXoauYRXFjcr4X7J
4iTAD3k6muPl4RlJLA4scDiscXqeYVtcJ78f2mpRtQHX/8865NY78g3iD/fGgxsk
g0d3Iby9Fjo3CDcNYCc6FWiaN6t6Ue3h8JuBIUAZwqct/ONMkNvRC8HdDcIUvTyl
74oW5oAoQEOdJHBGI91yV/QrRPa+jJTdVVstTMi5evvvnwAA91RivAFqyD8Z1XzE
Nfkwm9rV2kmcIfxMQ/dm+fgk4nBSIeCjzTgZIfKY0fWrAwBz4g+5lNA7rJaNsKnb
t8ORuAASC7TnhQKRv4dJ3vQtR3u8a6FBvr31vJb//ypiyjVSSljsieSMI9Wn2ccH
S4ySqsBd0xeJRJvX5w5L/e7ubidTvHgT2NJtlP3mnLtjM1p9h+UNmC5kMb6cCS/v
k9sP9yTyGc9BqUw4bfs7iyNhMfYZXY3mwRGJ3673vBBzNHco1W/vyVFSuSrtcGoG
XYmyWD4YQ/kz5nevN3OfnoJICwo/r+NeESFGCsSIiwBd1jY7osZq+qSS143f5Tku
ysos6V1WAE2gchKejz6SUOP4w4nH5wrLr8AKmeZVI3Hd7fPJEC8x+n7ziMJqG/OW
1s6ddzKSfhMwi1SiaCEG2XhXemRidsXgdx2suOVOr3M1xbSR76cPKu0UFDxJ9SFq
gMKC/U37yJzHusO8bs7t+sJRfsyD5h/U4AZzh2Ho9ckxzkT1yL+F+TVFME1Ve3HX
vgrkRkVRxNAIu7wzXVEoq4u2uwC4JKb2H9CbCF77jH283pR+gRTCxv+Y092qxhKD
JhSXyAF4SCszBAFHOwMC4/VTOwY0yYA04H9IyBc+M1b7CrPE1ITgozcGtYIoXiY2
EBWRAAECX/q4VWng4HnwSH9evtLEFpahcGWK4zoWsQDZhYIHB9M8rjgiVQw6yxaE
ZyHV+NkTJ1OOnRLM+0q15E0NRXyevSxdYnNIO7af2XG+0Xt5SWvUQSj9yPpauKiU
nlYWJJN373+/9vilJjCuFfcBNxFKliE6gK3FKYn4FGtszak4iJJNRa4A+smgWs3Q
Hp16gPbjcjOpRMYZ9eaumLLgXfMQmwkr9mDpycCkFT+Gv3tfMkFCCwrk+g5rxQS8
spM018sMg7KyX6K/BZ/vrlMdAqtd6bXa/HY4fxK0Z0FTrqrckSnWfofXsiKRpDaC
UH4BSpVcx5ZK5oyxbfxT8VctxbM/tKoelFkjqcPfIIeA/j+GFR1AmrW2bg/dq1+U
34wp6zKKvFtsuJp3fVGooPn1TGZVGQB615N9YQc+9EfOWlU6zLsAhBdaB994HWIC
msev2E5+4JJs4XHIvQlmyOmv1xFYQwKgsq9iJnOBmB2zPU7PvR94uiwiykA8M5ZO
9MNYnUQ6QH97/GygkRoZF/WL1SdYAJdCUHwgUWhC+aoVvpgtik6sjsivzvJub1FR
sMxpHzCFY25Dc61IIDJtsnyzptDCroiprQ5a/U/SIpDRFMRWazERpaU1zimT8g+4
zQqut9M7rv6S52Dy24vSZRuinS2MZzkMCj3YydaBZlovTG/MgpVY2RTZKMh592+G
f+6g+l9XquyPM6rYr4DUO5B7EfSdeiyP/MHXXB96nZ7RcMGBb/AfbNSaDn8ZaQBK
MSkB7bmhyHMr7lmqJSGIjq+S3psTW2RxZNE3nvGpNreu2Aijp8O+vnf1877onbR+
ipOgXNlYdjOGm5ji4NuUwIV9g90NvNcsXAxm6JFbv7EIcSZUK+4IZFWsGl2YyD7m
G4d2Y58MT0Lgdblim46xz9pds2zHYAYAm7guxJygg4IG39kAAa24d1YBHSiNEek5
7oqRmpKFmvmhgoQi+93bAE2QCz74GYxBlETjyKMtSkbUIJkpxSYg7ANkRd0EZezV
V12aLTqjUJD4063kookDLljMgqo8/UgdUQy4Px7/Ni9tGBHWKk0v+Gi896/kNFJf
kw4GHEAMPGkbnKcrzoEBWlwNu2B6hXIaEzfSV8GVrxn9DPwYAMWzwGr9QSE/88S7
wAVLJwe6ooEukHyvHNsNQGk65+4rMtXG5jheLar8SB3ihrKKgg5ELymgacIwuoYT
7ByoWCcmc+axR/HFpdhKl47y09Ty+MzscLWYtrPy8UljIou+8xnk2GNOduHkCyPx
i/raHfNfv8XYIE00bfgQy/mtPOvqle0c4RDSpY7qosSTMJydiNxX9pTWqr1MV8OT
TcafPo8rIVh9LQhg5Gv/C86xY1BkY+n6tTKTnc0yY4MPmlDcDgYzEYTjG1cgmXAR
LsxEyRkg8/kXr/KYrpgd/oSOVrooSU6gqQHMfpMeadZbGPdxm4qzHhy+TV0e4ccW
mSPAR2VGRfBFm4wO0YPUM9/4WDQxs08jjzBu9bR0PQlePKwAVsC67sN77gV2b1PB
HO1MFvl5qaETv4BP2H4XkR1ev73VCYh5CEgk1GZwlxRBA54SnEDaptYEyCwfB69c
W74A/QvJJCGFoIfLvEsq21D4Qh2FWE4UiTvKFsa7uqTd9jaANxaPuLvlYhmTpUGq
Y/2gMNZFCn9CA0iK3DU2nhE4xPuHQkm1oAHapqyQi4Fl8Y96jp1+iWHyt6Brqsla
Q8rMEZz70SAbPv9NgzbDr0CxAGWSjpzjNft61Lz+DpxCBqvriGqeBB8avpekm5b2
Cn9F4JfJwuPbDU8X/wf7+dqyKtc3y/aQgKXuXrPIpbhaYDICtGeBTuUmEPyD/W5C
JYrSaYCFliUH+QpESZshyueOgOXu1aMl3oNjGn07huescoqoPQgCdhqTktiXoZCj
gLzmZrj88EFZWSlF4ulE2q/3hWFwIv+QdSAh9StiJLM=
`protect END_PROTECTED
