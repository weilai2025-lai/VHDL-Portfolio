`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wGNbiCihJ6U2eGpfRTE741wuNQoIlIEYAlgLfFmkETnImJnIwbU8Egc9fUU1vlOV
oulZCunjQa4jH2AMaJSJ1q57tC8XoXhpNFVCzsmF8PX/g852XzaXW/DjLzwVy8Ik
beAEybTI9zzd9p6eUvelUgzP51OxXkHTqH24/1nXKwRm8cxDuJcZFwmxlPHAfHdk
l2qwbc/NlSJhe0t0DEDXngjQLRDQx4pmvb/RiARQkMlbXjkmklJlEhmuo2wzjYds
VObRwIpAG3S66aZ/Gv45+eH9F85CSSH0LlurAR7GgYecHuCgvfdAjo+1pFxeUPhu
kWthikmSNQnx5VJfgyvFt4L3LaOQPG2CqdU2vcgAfombKkpWo++3B56ZUAnZYJJI
pnhtXBQUrt/AZ4MmG5F5eXWt0Mu4BH2VBt+5Hgp+JXb76CO/BDk2SXjDxFAdCiZM
j1BjPsIB/JwtjfhpeEnPW/ux0QQcleBrFhzrjQXat8ouXunKe51xklCjsxSUeI8d
gHgJcBnbVdNY9gY3XrgkDCxIPMHXtEeQAXYBWC5/YqLvgE+FJyrhX49XGUs1puiR
hdRLMsq+SPiJfjMGlw29JG7aAVDtP9qaySt0lSEs8Dv9RKdCpCiYHu/xTaCG8tLx
1UkqyoOaa4PgfS9ga6P3uM9xgbv2zfECcLbfAeivBntrl9MnQqLYSMLrZ/u3obvW
2AaXbSP8Rv87e+Ek0zCsYPCZMpruLKQwYfinAZsuJmjDxdsDr8OrT1XUV7Y30ACl
vcbb4GCloWnleB2BgEkOUUy5pW7M9LpPpesE+SdDjQNj15JeHuP9514PUWxrncNX
HBoXAmnBL1W5SXzRA859qY2WOnmt+PflOpf7goWJ+holATL2p8z57Ydeh+YWyVxF
QSQPXmcJs6xrS4/8NYQ8JnFAheVes8OqaoLiwG7lq867jdS+r1bAU8BXPuEqng3d
nnUWpu5hHOlrktIvFe6pdmqMtCWB+5CkblsXOCPQCAwiVf6szPqzhIwd0sF/wIyB
ftaiIxUeFtxFALBLWC5fUaoWRW9N4NjppJ1dSxSh8FGVtL9QBrvj0QWZLrUY+Mz3
W6GWpEzrNASQ1XYxQDo5dm+b8KBv9JJ2BYRKbB+OkM65lnC48fm07rPu+I3IPzYm
D2PgP9OnjxkvhRv//0GzSy6EM27Ow1E7dWgv5702m2xQ9Mto9Dy4ybI/IoIHcpqV
sG+7kx3XpcA1IyRlDNXaazfCPaSeneOwzARfXbsph8k9nxsKc6A90y5K+dbFAcPH
Xhy2CKsJK6zsD6Qf78IQPHkVvarQG4H8NlzyoLYcP9bt9pxcMHKRmaEOzeO3+lrS
f/NFQ4y3ihc7PUbzRH9NZqL+6Qr3rZSNNDht5ygRaUdNJSD7I6hy6BScagK5ls8d
t9JyNj71xWPMfyvw+9Fu0+u3yqawLot1c/i6RLTYxM8JC/WB0q29I6SM80Abv0z4
zT+7c+IGztmO0dAAg5oW8FGae2j/2RRYg1otfF6LA5u4FYuRPz9wTOSz4XFyastW
1YCsyBnc6vZ28avlT7fTztWkTJH2R36MBk4UQpIa0Ofp5+ljhcTT0nyGhQ5sKyOT
ntdJqe+xwVoZ3HKBBtP1AZHbD62UUHC7z9EhTy52IdhKWm+0JKha+xMX99JtTqQi
GSjfmrVfcK6d9Z7YHss2p7/hefcVg8F9yLf2Z60Wm5djyQZft2MeAB8hTTVe4G5Q
4FpPrXKSu6PWwIaJlZJT70piB3l8k8N/DtiVm5RDEaJq9wEplLnxyudOwUnHSDBO
+GnkkiWR+ZvJbYdj/rSb+q+TtA2ghlQ6lBKjUjI5fKWE8Zjs9X6CH4PmOpGEXLQ9
7t/TtAHoX+TioAJMXVa4L423RGVytJVfwrgcB83caCALyv+QlZ2LU8olID9agGOz
IBvSl7MIM360q8xvtNE2G9cX4ROANYj0rJmM39G6T7JKD/zhy/N9rSBStvf4UGma
DXM1qcloyDINHDn7c/2H0Cj2N3LSN5L5/4ddsb+1B8xMAXI8zBoTUpsN+I6hACgA
t6giS3TJNxK7+b85ssBn8kZv+BWSsM7h9TKp8Bq+aZd1+BHUkbwpw46vpP9O88lH
Fx+DrtwWgNtseLyYXTU5DhbOT5tB0aVGCC0dVAkOIMbAzDucPpCcIuKnY7LTpgpK
W12t25SqjxBN+vqbaAvobthXfC9OK9j6jXdz//j4PASWIIwCgTMAlme44/Dt3WXn
k1C+R51zTuRwOmFDgrMnCEZh+stzUt1TUohlTbQzU1xoKPR6Fj+7qOtuDpvFxluG
GXP74s4zUcTuOLHEv4lx9nngjJ2KOBUpmjBqUFqNqXNO/LgrAinYy/lLc22OFp+W
cb3gS9YolCXSAHeyo8QVUb/3jnaZaSwoBkzznMpy+uC0sSulOPwYT29inOa53aAY
8HMN/XHqKl+IlL/3Sj7kXmHfom6STKDcnd7Ge6L8ZNQ74cYznZd4Q579xJGjNwMr
ZgAzScA/08S40DpYzsYj6dPhX0H/TV/eikvIrj0JCd07TEKg3YlfUZOXv9TztuGT
NuDOqHioTdHe6XU9UG4fd1kw/fWWc9VaX4cX/JG2zAmCfm0xVpa+oRDr5jAq7fWS
emkg3TLAv/hqt2u7hIHe1fUHd7wIROBCvjyA+LGnJIO10o6EonsdfaSVD626lPgO
NI37cGp2Lgm1HI25g2b6sCULI1xK1OWvZGM/vcjJ25bNhlSL9507QOp4kAwQ+FND
6vmKWprr/N/ubM0vdtrga783/bCt9SKFR2FEz+rN99PUJHY/Zw48Io3UcP6RnM7k
SCL61esyWFCMLbRpwVzTfWK3BWtJgmhMNhgNIgZ9VXCrRtapyj8B/vJ75lrM56Bb
GNEqdjZN4Tt1mD72pFbg/5DmWwE9lQi8L1lBAWcaSS50BSksZx1EMLYZ1Ffq/U1X
NKWrXLjx1MLYV70+Su4RBBWrOb+PMDFtmBc5dvq5OTo8kOiW2YwGsc6dKxgIvUy0
PQz+ZoSAseP1bkN4Sq33xqsRT12KXRyZL1drwKGT6HHrCiHAtxBk2DyCg+6Z/kP0
u4+GKP7D3uAIdFRilErSIgSTd2zUjSNsuSsKCBeQOKXmGawitswVQZpYd0FobSYF
x9/iXe9qfjDWEsZTa6vYrwdu43qh+G6HxArUTOETZiKu56qjhN0SLF0jUASQobOM
JHWaCjbZQh5xYgiwNEY4tMw29iOVXxuMmFA8nQqF6ApQteoQzDFTxvVrZge7vf1h
rWMJtRUpmFyCJecz5R0JeoVx9JY37dYWRxWcvznVAjkPImsVT5ZERfKFCewzk3pI
D7dctJdTK99QzFebPbZu41Bl0HNsjtsMfhEM2fymyIGVabS0V5Rd+4S7l0nGQ0Nw
ldMTdGPIjpkSrU64PhcLbtPQzMQs7GGmgyKWKLH8bgvgiHrGV0QY6m5AfUX7qOJh
2yl8Smr/4Xxo4RJuqnXXDXg47MDLdQrABLoo/aQup3BZRg41gZ0gQKCEFRF98570
5LFBlT6LFMEIxvd/O1QJVwa2sYWT3G8bn4iD6QY3wxxGi4eovDDDCqIrOtQetQNh
GwhVdrTGPAHG7L17jrh1O7BoFIK8d0LE0jYhof8/Ah4Ae8jAf5v/dIpByOkUsV/E
WQapRstK0ezSM4nPlTZaQWskOH3vNEJbBWx8dBjTTG8NFecJOeS/U8GgODLxug64
pSF8Hjub+BT4fcr++/GaCfe5mPEVRVthBs2zAjHfGOPmchbBxRd93gDfit1TM9Kr
B4i6y5LPPvBJSlD1HI1kfhd1uVdjpo4pAhnJwP43Zbv1fetiv6O2Sls3ygQLY2/0
psdNawoVdx2ctgG0dBz9ssJ4SFQXnGCrMduFmfiRk/MWJK05/DiJKXKYTBuoSNcp
IagdjW8SnYHB4yXOCJlyyShkMwj2ez0zcCDeLzg/YnNU6pfqj9N0GJD0Jzzqg8/Z
m00vtdMLf+8xkgNqFeWkfI5xL6r4q7Y5l0+G56IorZMpsn5/2S1oMqjW73Lh7Ql7
/pmbIgTNlXTNIHyiyU8Qnjz+fZD4ZtRzJNdXyIKxM8aoAalaRFgNnR8wrhvWfdve
1e61L0//fLH1L+J4cX39SkAoc2h1jiw8bFHqwozDQcblycp2S2/4zwZTi3w0wDWM
u875AY4Gaqk6i6ppQ4Wp69Nai/8ISrhNQcWAvaylfMgW+1uGtuYJCmuQFIdgVnsI
y/Ua7QT28lt62uA1VDY24ApnOnIhDD7juLteiiEdjIAoze8TvtdUQVWYUAeQs78q
EY0Q8UPK2u5aXArbe30rg8QBeiZJYWVnAI5Iz4eASRDiAowe9/6ovYY6C5RjaeSd
39c+u8b1kqk9RaIBhlIXPKhdjzrIVh+7FkpZDGviIlsGMKmHZZm3DEe51JByhRDO
T8j4nkkCkTbk2+WONwwp9HgW+zmq7M5R2RkTXfdRaQR/ftxALanmRaIzohCgNjkA
4B9Xi6ukFQf05oQQ90hpW8WNkIQ/qrd1oY7IT5M9cJ77UnQG85v+JNiFMnkJ6JtG
4yt51273LAR7BGctjvFN2Yxwg0f2KsBurVG2FSKNVM5gNJvFulAsTu+l7VzDyrgC
`protect END_PROTECTED
