`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2KnqvFN1dGCT0MtM/Tvi2HFJ1P10DdFPeZJYpSHOob2Ymc8Eo9POpnfNgcdjyka
HGaglHksBQT/DljNQZMjkeeYwipXbSZfkhQtSIKTTzTEFuV365ai1/J6S76/tzKO
oPxzbOUwiIH4YpLoaEfTGDvqKMqD43wD+XB04QZv3YlvAQj4DIwTPaEQ3ajj12MV
rmPrJTfGCjhLxJ+zsBco+ZutARIFlEl6DPsdQUZq2CKiU+O7jEB5nYs4fHAPBKJU
Z/coOg082UvXP0shN0LGjHki1bcRPVY+Ac+D0crojDg/uqhAz/oLpy7keyWU6zw9
iTuJK0wwnngEToikR2UUehInpswHsofO9bc37JpqvVTu6RcsVeL+K+YnStIu12/L
54CiuSIV2lrmWSGKeVHQKkz0VU1a3P1GW5g+AVoDJ/YVm0LuqFXTUTvUAbb/R1Gs
Fm34jGc0XISpA+5exb8tIuNu72hs75+qMbGGUp9HkF0TLZMJJNZRHDXOcVEYdb2W
`protect END_PROTECTED
