`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZ/CI2bI/vSVz7GBCs2U8pPM8dTIXh6FTxIvLkIb2AfJ11DyWNefKJOI1A9Q4JBJ
sMiyrrixdw/YvZvgwO/I0FhOZGvwxC4u3CTSJkK3YHMeSnz1AHCPsgCHHOPxwuvJ
95kGlIHhsWfYUYgjrFYcnlfF3aXJs0/zAQPNiQ4Ynjxx0zvFO7nngWL0xJs90bsk
amqqUp2e0O8kVziPMhTYScT4C1zDZrz5AAjts8/wLKHjDz/ASHzIMH425BSVE92I
a6mH5ihSjerGPhMU7CCl/PdUNdkIPyE0ND4GthA23gbEOXO46TSWXIbF0dX0vb9C
d+yBOFnsDx1eqpOny08GI/wLUgUpM2FsOgysJW137jXFv3j86ycPeqwrpyC0P6Gr
6dTC8FxvfMNh8ZnZDqeMpYao/AsJnqk1ctNQ0wfFjpteDfuRuaD902lMGlI3SLyI
bhu7n1X/1ANp3Qs4gEOMyGrzhM1iJq8Q5pCvTw8gMQ9AdnbnunaJBGFSM1hUxAmd
7feZGJs/ek0wif6S9Y/xeMRuCGsUBPkOSalBtyfuGOy5dzYfWYhNetApC8xuSRvv
hbCWQB14tgIr9VZOjGLngUrKyQwH6fPTGa3kmN48XGGbBZvOiUDmUeiaLtXIQs0D
nUjwmL1aU4Q/yanJKgXTWVdo1RXt/++NvD5NDfuC6OMdpBm9gKQ0/+n45QMm7ZPK
HIcjxVAM4qL83fefy62i+QnJSMiM3WZ1UbSUS3VRlEkoT409PJqhXGA08wSkbao4
8JgmUVsP/uau5jts7ao/feFt38dyjSOraePYTOgagIMJdcWnRRZdsIEiy6gIMLQy
hL0t+inhOWmiegKX7JtvWI5wj/iS69OHow1Hg2odJvitpQbNpMekPdzogmupNqQ0
tIVGaVvl6S9UdXo3nUEimDhUaqpD89H4EOf/8o6dzNM7pETfTSRNak8Vp/za2vDo
h6Q/qpvaTSAdCOiwkyrtg4GT2aIpeRLLQFtP+IoMVYOlf/O9CBNLuNnBTeQ7uRPE
vkEXVe5PCtBU0fy2T2m9R3MW1GXIodBKaBx5Iv37VQu3/RCNse8qB35y1sZUlRut
i6Obbeyk2WI6As/3MBLoUv5wfP3eJdLYEil3fXo9Idgqk82I68j62jGhN1ydDS/C
0YQuAwrxLW4PPxBhtQH7eoEcEHsmb6PJX85aLmDOnr4dLOP0fdEIGZyPpUUMMIcK
hbS7y8MWWDhTnB2jPOqeA2zMmew11ojeVpUd5pboT6cMPFkqDWPgPuPmJUh28RKB
XF04lde6NMaeXvszrx5r5d+1hLLjebtB2Xx/4SHbSzL+P2zxEkYpSwuGJFPliCS5
J3+g1E3aUGWxL2vCNCEXIr5/mPlk2T3yfrfYxerhYrPJxO4SQabwti2kjb33YcEW
Ev4hvd8n946eX6u9FV891r52VB2cYDFlNLuDs3LXMduo7UyI1thPoHt7V+5tuq5j
CbluMLvNhFa+QiZ2mOINaT54cpwnFUn7kRRZxZ+CH4sl7NMhYyno+XXk76MOKy8i
yeIZf04n8cz8ZZwgtb2MYGYdZ8Dp5YlPhPMIUjnmg/uMTIFm05MbvaRw31IWN2pH
C7Kfrj2+D9N4tnSZRn5ziCumUWmFP7zoJdqgcC5/N23vNDG6bDG03ZhdEG7TCgR5
BSPnfSQYB7L5vY3WF7qHyBaWEXZKgUJX+ctTA0CwgS303nX2u5cuuxLRC2l28miK
px8WLG5yAtQHnHxbHxyTQMyJF544royFuvN5myz2zw1TXjeYWJv9NvpddYw5uq5p
U/e3hmqtyuKjuqrUspHqCdB0uC7Poba12lUiebl2QoNACYm65DoCxVs0keuLK4/T
6v0MuEPVCTOntj2YxzyCQdQIHMgOUCAs8ThuKWgxainQS6EDNo1kgppIr9sf3Ytb
gvM+K4GObfH1G7Fsx4RzfeVjMh2G4N2dYRmQbSyr3M8CSTDoqxWSht9NGEbcicEq
R9xxxA9zyvlguc9cHnJKKLWR+zvsSX0RvHJTTUn0xfMVOm2p5+ouu5uw0csz97nE
faioBz/9MzRuNN7TZOXj6tvJMtXUkhvEZiji+F4IP9H2rVXJRme+4u6qKn8DnP3j
zxf6aUZN5Uht/shY7alM+7LGraajl4YoxYV9+r6jDjDZU25tL/dXLULWD0CwX5aL
PaNm3lzSpVcT2i6Z90TsD6J6SVgsHmcOelD0SdW9BB9Qv+FqnVhC/5yTcwvvYTEZ
liHr1jbDy4tOxxaTOj2+UJ/3YVhKQsvcoW1Kop1yqdY99vpGE6L26YvRwFtQfdh9
geLguOco7+M30XF80G3d7mQmxbaoYYxIu/rrqPgNXtVaL/XK5uaI4EKRcdu4rS7e
wc/kv/5HQXBtZaERAGDj0+7akjJxVJRJ8ViD4rEzQXA4OjWMJTc2LJmpT/AynOZq
i2yszidYecigjGFi7QsNGvk0XEDRHmm6y8W6n0f8uaIP/JEd52UfvknvYFUDQKJn
cYSh3bU4nIOmbFzPr52WGOblS6W8GMrATEj8pNlAVXCWoUjysmaoBU7KoO+/hd2i
EtHGj6glpwYc+VPfMCrGKAXYTjgrdtVafbOz/IICHIElZBS0Jo34+Gk/bAgisgKG
um7CbkNbQZN3mgDG37vt4fAOVIBABz09DLeYUJdvlFZ18RPN1dT1mvMTChcwYu5V
YLDyO+hD2D7F56FchniW60BOyG4C0+RCc48zNErjEh3oFxZzkpqM2brT9/CLJJam
05BkocPs3Sqpc7s07dCb/eMJ1miwAsN3nxbYFTWPhuhZP/HahxXnxgEZNEyM1zMk
N05iwFiPoSpfGHdWSIaY4DnxUz+EM27juT6RLTSU/fBzR9+rYkPjAEJdarLrDqPv
W1Ld0HjqddLB68N3Zm9I3NrXm2lHMT04kGM+19OKmRudswSvA2UaXhhQRT2UIN2U
MZmN37zzGSbVRmBxOAmjG78yrFdbWLGOW9zGeq4YiWhGSzoyh774GzVUtnrmz4+6
26jTfBSLGrV0SuO7VC4/CSf/le+fxrqFd/zUbln9+2MTPjFNq9AP1A3ENWZCuXcJ
G4mz9OiAx3r0dfJaRuC3G355R+4G5GVxgIWa8rpzdl8Byrfspst2Mwsyqpp3UWA3
b0Tenw2ELiKqBNlkmDuJ+s5hSgH0fE1ugKkhRYRXMheyfLUL46Xtb3COD+VRGkCV
NbXPGeUQLdNVJp1yJiYyJz32TV1OPv5vzLV5grvw7kwQliJxXC6awW/bZJkAZ4lN
wp9ndHbNhdbBQhDg/qhXqM/pAxtxcS81w8P3bRQmWyVEsJB37CiqHNBK6VFqcQss
AWm1AgEOWHFqoVqP3ixqTe0Xt97FkGABpXH7WsFYLCwcD+PPTiPKL9e3WHEgSdj/
f0dqNCcEZCb9R3n32mQleMRIrHqWlnqMNhWoYeQ9XAetlfB2g3IYADA2kFMvKeqR
e3yYbXu9H2ZY1Lz28DubuXL3Hm3WwaY0LtVphQyMA/P9EwwtrhxrYEIXBM8L3XNI
3h1yfZ99ZETYK2IyFoNYe+XNhnVJePWEyme+QtbiZObJPQADSPnkGK9NhnD0CD1b
uwE3KxU6U/gpDnuf+QWPPL0Vpr2QmwOZu6cxxxZzQyIgAcRGjRcCO849AWA4Mw0t
XIJFXtYhsH4KnW3sXbLsUN9LW0vkGuRoV3HC+O63wADoQvC7yWgQShAPG53DzZls
`protect END_PROTECTED
