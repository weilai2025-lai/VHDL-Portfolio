`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z06mC7xXZ1P0iIpkPwianG4PNVZHzTLvoOtmJrIqKwuD0W15W6gOBDb99iYHR/qI
HHiu7xpJhgccgoH6S6d3//4XXclMkiahfE8/dJ+RRgEWL/jWQwxayW/vGdaNybR2
bFpmPp0n4beJicGYxCgkJrxuZ7RAxOvvw1n5Vkb/0wHjrCEV6ztxSgycilDmFwE1
f2Atu3CU81flt81ectXodEM6k3m06itgJVvC6x8cSNOipxdUIcMPMzXfqB3K7V0B
yePzfTMlLOe9QcOkFWz27rbNBiC6YNNomHhMe80yOC2P4cgbJm7XcQdeO1JQtbWh
pvAsH4+OZwwLLKlRzfvw1wlRyp+zjGZlHF4yNEtEjeC5ypRHae93ObjD1oYXi7bU
hfQkj8vHl69IIiFk256BfH+934mwAFT/dn7jhp1Fa5gF+DVCp43V0TNC+8Gfk9Dn
rzh6qIf4VirGKIpVIIhfWRWxLg/ltK/GWZWrEEW+66l60byjs51bdEOkbwh4yydF
FSNJomB35ZL8EVg6N1okcD2VY8ItSaIhFOWT/+wIgYwbD8Tqh3wnTQKa/LAydHJK
38Er1qMue7yksG2KGttuc730gcAiyIk6S1S6Kdfz5AFfunAt0dSMHGnKH6dfq0v5
Zh+wwlPjjrGJ35Nbk/kLBYvOeJOTlUBR6WbTxjU5jCvh+XOPkoQTdHpMFEO30wZm
tm/gFTNyLXYuY2VyXM9YdHDlT+I80cdNaWwtRMAflBun9Wws7x3SIBjmvxCJ+Kl7
/w1DURrrQXAa+tPqXpa0f8u6a6w1guy2098m5A+n/77SmRHvxZa6ihstSMNWChEc
N3Z7IgoW+zMmsgVesdTCbZI8lZWvLWPpbYBKGh6Wbfo9EWZEGn4PhlhQP1edtVg/
eohKhjbcbYwZM9APqUjKtBvF9OkWAjswgAdX7JJddi+M0ksbqbf5oCJjVLp8cUMx
DA3/KzanwUf74xxWx2LhKDEqJ8bpNEgt0PMYpOHuX9sx5Lj51NhuEUpgxLBY05A3
JqlPt+keZx76kAl4LVHajSiVJYdtNMPU1FAH4Ce5L0VEC0zifqQHM8+HZCPEIcTH
7qQhcfzrByOf3jsYaYailcXlQZHyo4yAUeEgKubeThbiEtTvgORyAeXNZ+OEqRlD
EwZ22d3nFITcg8XKPAVgXSMEU5dR/RkHUQs6HXxQLjkt1GgX1xRXS6R1/LmqAXer
bQCvYqeZ8meKv90NHL9TinYYqDLL1r3BcMGQyztmEIYCF3+wff3NJ9i0dUnxraI2
YOSUfjELqM/BzDNsv6JAGIAvYeNL4NCBx256xC+nKQS1znh7fHinf1r2sLRCWXSl
ut9wYuPCTSSxgz3WczFCM6a9DRBYfwyWXZRcJuq4aNbyoEUXZsNMWBiM4w0QJOXG
eWwGQs36pnPdzLdyj1qrUzUI/Yarvww3DqY5Pu1kQp4L2h9h2qJj+NGIlte1boxD
AydIIkqc51A1VGdVw9VTmWqpbSoFeV0qYn8YnZNfB5SR+tcZD+WH3Zk0ZvC7Sd5m
AFLkL7Odh+4IgTpaR8FChfHT+W47r8uNIPJ9g6vOMaPcCtBepY/zLJ05jVXMwHIp
fc6Hcu82vrlp0BkpUlGTeFZFFUZkCYWJEpE80Y5RTXh9oE7wrMO7HzhhNwMEJ/y9
Gb6ElcJfDggRepvtdr/anIEOaqaWi4U5tx9TuO6xn9S9629JlyGOyJvJoj2iqAkX
+JdN7WCc/oPNqOztWrIrCMpj/XNrhfG6U8qGtmIwH3VoFrQVQ2piKCAoImMubGGl
hZzgLrVDprQE/AMz1WNfTA0p3TbSGgXdNQku8tpIbDP5aBmHmF2OeEl5UXBZ+aVY
PLWiG+PvKmU7seXM/IgYyRlx+PYy7lCYEQnbnMkK8uFx/8VkCtjCFCYu9xlIjr0D
tdv7109gHf1iht04zaWlbzwCjE3SPfcgPAUTefgTwzITe2yXj8XD3lFpc94TYORK
BWdP54vtbuUi5juZkRIanz+8Y7BKkxwtjQ81R1NRls8RdApPf9mwqGXaziD51QGg
TAI/hdXJnjCl6vB9mPw8POlgzPD9kMUSjLbaSdgg/xbOIOjHBiwitdOz0jOyt0qf
Ly9VzqScv7GiedF6vQ9tmlCY9aX+tongnlERTcrlvQJjMpppTpIm3Sj4/5YntAkZ
XkMfCowL1bAqJMRB0JQGRrqLqTb7hOtkUy/47+AVPwXIa275y0WIFssnqNwNPs+f
QXCCGLuQ2Erpel9LuXFjtXhSxUC3Y45XE33bGXf7DBUPe7rvzVIXOzyvhFTj9LR0
JToVkhp2XqlKPfM6gymVjqSYQyjq46drtD3cI1qGRp+QRIXQJLBMRRCEH3jDbM6P
+6D4aNmP6Ouaysqot+Tw6ui1F98k5wq8b7nyfNsRKl1xyUo340EOrvqb3PT9rw++
YGL9YQ9hzWPhkwrpPM6R78IRsbxiFMs9v2DxZzRpSXzWFmqiPgnV04Bq0P0QvNn9
XMl3VdUUFOe3W7VFv6GRF+I28LyDxpFcpUjpcll6NnB4KasMalb2RMfb9zypuY4i
bsd0XgygfyE8Fs7PNA2xU8WB51rj3IJUhCvRDEZ4qMNqsYS1Uo1G7cflaXqje66L
Qn89mkwEFEfrRFVM3St77bnAiOX9RYE9iBuD/6EcrzVCQUEwaDHv9m2KROLxIBW4
SYA6zorSZEXIEZIxItb4puX4Sqrna/dpGSieF3IYzzsccZZAfMVOdMtUI68d05nd
joeZl43SjkKMolaGtfSHkrC2hsdvXun2CxofLKRtAXGDQMZvsi8bgb3+hmwk5trr
Z2RBXXl4pFKbXUA8zL+7ybeAtmDYodS4wv0ZEdhbB9IXRaRkX74E+dqtiraJ56vx
uZbxocnXwWr2s7vvW2uPyxcKWLicsaQc26gPKICZx+UJUEZtIgnVzOgr5B8rv/P+
nv5VoAd1AWMnlVPr/7AULkUqn6jxylhTeb7RsY9IHn4BkR4FE3B52MmNphcrN725
jviYuwunj7Qxo03bajHJqP6pS884YKnyfsFS/0Cm7amG9vxDSWy+w1bfZpWCoCTA
dmFiK22f5Fa8I86aH3C406qSyGVidUdi5wtpf0ovZSFwxXVC8kzueXk9DVVJH8+M
f5MRj3KoFKnJu6rlVIXxTGRGBpzzP6a3W6xchuEjQLNiV6yXjd3/LaItrhcH2e1R
+f2ry0pZaw/q/7rPYTcbOTY9onFHnRnrceLZFb9MWf4dfPdl19ybUw/nPzAxTfyr
Mu/5KJiK6Fy2JzfsW7Teq6FomzMS2gS/gxXdr4STf5dxyo/NDk5WnpRU/+C5LaUM
vEdkg8Z2DUbvBKk1tNF0Zc393u9mtMV556F1yTkMXHezb1huTe/EsK4b4TyPOPFc
wv3An0W4lwIfLAhT2iPWmGbvviv+x95UKPBT+fjmzutbGMsQGPbgEZvqrv/fiJhb
MmtXhZhhqRv9OSUMvQMiga+wGb9qRKqbeAywvUIpch2dcohHw1otsfTGpLg2Mf1c
7xAFWcG5+Cvs1Wu06/+DcC0D023HmkhyjFbP6cWjSouhwg1uuTwZPGs+aEWHPpQC
Url/RRC2cQareG8eGNs+4OBy9fe1ifBVM7W8tNyjloGF9LT4Bl7bzoXh6pEj2Fz/
dFikgN6gPryhPrs0Cjvh7Ki/s/H/UJOVre6W9yrA5BL+HJuaW4MkuHoN0KRQlb0+
A60/73H70sCzr2EI3RG9BFD8bUBs38xipf3zivnVzKk4oFTGIZPLvs0r10g7jLgS
lFGWaG+J2G6YRhJouekFbXNKr6IVrsXKyjwDhNZJh/YPMxhVAnJ2vgnl76geNSm5
2rMmjibnhIV21zvqc+IWBuA/CyclQvR72FfejC/3nmY3ncrRhDGHppaEmDOu3Gzk
aTUsaiwl0vJ/yDoiCLE1AejqR20DaRoq9zKpS+6tmpAYvoKCBJkaaBYW+3iAqOOv
a1tGbbBqWqEkFUV6TDmnoSS3+2XNg0HlVWqU7QjraqTcIcdsQfLcudU55pWf6jyl
hzpD5BsrXmKgD8BX45uhPmccukiir5N3TCIebEov7VTDKqb7Z2qbWW8HVfFjIbqK
eCHWgyIcc6r/KNKrtaqqv6EiGjJC4CxtiD2caz7pxnQ5W9raFCv4YpjkRRWSfdjK
WZLykR9n9C489xp4hBCD1EvcF8BbnChddGrgk+h1N68ut51Vv+WVrR6L5KcWjdDn
9DC4t1TzUsjZwaDW2J+FauiRgcN2qHYhiKWX4bRFPi0LcSurzWHf64cKJaWUaJ4n
qS/w3qmHDZUAJNDwUleLfOj1EC2kL0J6k4OTFVGNufNDeJfyWnLAcrQqInxtva/C
2MB9D+vSNKXfUJyVzSriMS17CrHJYy7LByVq8BYe66MT2mRv5hiOTWol9Yec/eZ7
mFBNMaJoExze0kI3RBYap77IKPynH1gcFXKy7z6+s2avTNwn6W6raQ0Wr6rKgWKa
UKo0PnmkkIPUs/SYZaDTlB0xHLH1QdiwrRBPLFqH0uV4f3eY15+ml/Q2apHs1c5O
B6J5lrgQOax8iitXbPzYXt2E5J695B1g6FmWuhyGKpF0MAT5h0SZHGAMUlRa6DpS
xrG+9rKzB0VeOTDOtEFwVAQi11qQJ7zkgxmr6aiLkM1IdetyM+SDfFGsuPzhA51Y
mmmUbWWR8YxgzyqnqObZWrPG0d4er5iwff7iuMD5xAQUixCCpAiXCsBuQVQv2gO3
UDtCnwQQqhlaeiDaCjb0BvBefacKBRhhmiktzuXuB7lfF5NVk04zhn5sBJd1xnkj
7mOK84wqui0CTXiUQENYYd8GOcznmXl2nn6HtOykzYk2qtZoizVGKP/XQijlVQY0
/CJmiw1VcMWjLUNwZ7cl2/tJwPdPnfTnwfTkaH+SiIebuhS9XpdrMdH0WYcUwJKR
ytOsE6VIJKNPYjzGB42KV7OrkaZgNvC0pdQ01iz+czW+4I7w+xdUaL5lMs4UX4PZ
qA9qMogUHFuLjhRrvkXxkDt0s0dCF33+ELAYswGMA/GvdPo+6YKv+gHoYcEJUEby
WlNk9AhhDamMIT0HJKmMl72yEd3P3psDRyguB6MmzxIE6tIfd60nWgdUrLuhKWE3
efiCI9PiqaUG2salzESHA/sxoPbw+G4k2RHmW+htxq+73bAyW91RnYWRzISeGqbB
WCef3sfDke4U6SA8v/lqJ5u22YSO20pM7oAfFZ6mDx/ATRBMjEe7PRAjLtd9R+DK
PiuraFA2qbqNBD6VnCBmoieTSrMSi4SqeAaCRy8FgkAMftVASI8yado4dwN/hO8O
sblq4cCkmKU3G3EkI0rwmWkjXvTWamjQ8iqwvxV+dtRL+PUtMxx2hgE6+MIg08+k
pYEuSnQL01hQiem+IWtDcRKIo7osU8kwHXJ650A3fgJ9v88iH9K/9PmIQwRpMvja
2Vfs1OH5hXyITEVilEytLRc2nI6hfTgtvdFSq8wJ8cyN9+A2McYZEysrppX7aFhW
3aXEvkX1Lu8q/QTe6/kGA5MbuEFJekDOGFUVUs+E379Oii253feOznpjxxXZrKfX
AF0RYSkHVQQ0j84uUVFWVk2auYMC+2lBMU5cXz0hUbLFBUPNIaIONunXlc/7d3Un
pwszpql64hEopMORIjkFrFVyf1z+Pr1mVFM3+tHAdW4LZy3Uxr5avw4GUN2advbt
Cgpk9p17gpfK4tAnlMue7wk7UcMSchGg9BZyKwXQOalC+bM1st5Lrc0ff5KI5dMk
PDShQcv1S1KqaqnMx2H7/CT8qjJjRsrNFe1gXPLphvamG+gCjr0L4IScyHpvMi8J
KnJGPd+2LUre2N0Jde1E28lctxy3hd+dWvQMP68A/KY0JxTO+2V6JOQODt1avy4G
albnt2wiSynt/HcFcNEquKaii0NLp4Cv+2NElcAgSW4XpU65SOKS2356pO50suo/
2ziMqwErYm634Ca+Vbo8H4HEqDHf9eyv4moB2txx8Sl47jtztaNolV26qe/ZcvWX
SxC8m6AuESP+gHQIh4Ep8Z9hlMAniF6FSNgEdvRJZUDgUf7uQd2OzsnljPbUpUzJ
Vf3TccpuZ2vxfldXEiUuKYUMjkqRNkq6dpmtvtluyYw/pWWavoK25w/ZIefqOMyl
l3dROmMO7x081u5wY+9sY3nZpX//AsgMkYijDm/oPZgObDxHsN2oHMO5jwjlq1uR
OZ312Bo/WbpxwPbpDbsBVvsFcxXUb/SMBfJueiogoIGzHcAivBRf5ZGlKNotL6lM
OZrhoIT7YkMMtOkbGTCaUEVlze7osJP0FZALsGsFdYMZtX7ZmkFnKutkMwSQrQ3O
VN5x4iCRFs7u2vp2ZIz0up1OE9Fli8C0wTT2KpAPDfBGO71R6hbUeq4UDdIr80rP
OayEvjN4TS7rZkwJbQoLI6rHjJH0sq48ZDyLCD615/7Ih9AW8rLTNn9UC9FtG+P5
Ht0w3aQOeqZftljAysp02E+bk+ToglzP/wxXxUvQbCOhHVnK/xKhn0FrPgvOwJRh
raKo1WEeBfx8MePDvR0U4hEoBIdb8FcXrwgxODqoZhV+5+z42BvxylqZC/aFOcj9
Oh5CEahK0XMpFVls6gQheWHks6YlthbHiEbLeiEduKv/Ak6E3+gRTRfa/gN8C/rb
SQEMcjZ2PwUvvGvCheFMW1j59WI2f2+ltlwib3G8U1NEpcaacfiTDdjSuz27RGLM
D11/sKaDv0WLgUmi4nHpbChXFgaxz2c02AoYKu9t2awDb6rmkNOqX7gWjCs1vzCt
koEXpPYMTJ+5v+TA/GvIDCegk0Lpu/q+8BYDQ5aYq2J6GynuZVR/QyCbdSmjtz13
4dpsAqeQpIJycjcZ55QHvCzmU9Q+LwVzd1hhQi2eNxzV0vZioAjvLVV89jxw3tmx
VQCM3Ys9oJHk57DdNH4b/aBrUifGCQ9FMH1CcmEgQezShYu19NDkn6PIV81Phw07
rxBtD1wbCntXVN+4Z1kTaQl6ttFYbRbsalH2ktkXZ9Byzt+kgWE80HLS6cAq3Qgj
hDNhEhWIVtspGaaaZPJa1ScmDvT8/WzbQmV/sAjOPkOTfr7cOKUeq6A1c7j6iAGa
PRjTGss5768fHra7cCa6Hf/8EJqdWU9D8B49Dop+nFWXKh/2RC06EKkGrpWp7v0i
qGxmFhhAcq4qiHH1Gbj4kLdPCU3bSCsw8uu+51YDkEZFpyofcMDSUYmFqbMBJBzx
dFsvsZS62pO9WRceTWeomf6ko3JkJ2TjSl/2k6vbSjmBn+/4DkxChFtntyBw3Iv1
2O0WGnr3ioKp/RXtxi5tDvLaKMjDOChduC9I2E8z3OrYpWleZWNlpzgiSgkOENCt
1ir7ccvUvx6cnN1Wre2GJuCOMGDoY//7S3WzEPjzkAHlQtK1WvcZJq30Uq00iZjB
+svq0XikbOhDTfERXJnwgpJQhkl22Zuarwld1lPe4N98STdGlDl9LrWd7q0971cp
8fUB/C/9npV0ULip5fq/w4xhk/yCXWNBZiZsyqaGB4Zgdshds6tkh+uGcmCBpH54
YN5najy+hh1POIhi4VPjPv50e/mVgCSq2xrB2WXBO1GvLy8buDPi031b3nEd4MUs
5PsuVAlOYizxlE1RiXIqOQSaczKap87FZFMfSJtqw2TdlLDZCHaA1HLnY323b64n
Z8CH3usD37TpaO88INp7xYSEkwvqpA1je9WuSqchlhcT9THssgE7FzhRbKDjlSpu
boEEMAeRuJ76nVxpvsOhDemoC8jquAE6scVabKII89TbIsg04XG7jK0cLkQSvuKB
hg20NtVGkMLPrnORqNSQQncyf8Af7joCWNkMWRRgEAdZgto2h7fcNt+UgN+g+/4O
eU/OGn5tFh3+OIs7LNpZEhnTuJvzFukRnhxsA8jSGayrF9xP4Q3U0lrzHk3iLBbF
Wl/TEOErv3UUtj3Qp0cgHEMS8zSrqP8wS0MR10bmZs4X3v8/QpAHAwOVyDOLc44Z
gAXdunDGTM7a9O6o10FOqN8N8a2FYUKaEj058wedbRa1oXT3BsRtCQ2uQP6XQoZI
65WZOHP5bL0W1klWjEfwRCCtpaAmgI+j01TSDWoR1k/vGIsNmJma/SLGnHwovOYi
5unIQNJwvgA22bZgMMVlvxRfmmoDV3ue1Az17tzdEGg+U9N57MkQUafD62xODojO
wuC+OeBwYLEHKYyQIt2PdTg5dMPLJAEkfBs/rIr9J0gF2qRp2moQj2fZBWC1+G+f
9/tNfIM5XD6Uk1ovUGahERfwvLnmmNUJ/nU6aldZfZEiatWGEydivssHEIAQg1ud
52TSrCzWFcVWClPM8LtccOEHyJQy/aq9m43dAq8YKUdAp4y86IBtxg/ElDZhfrEx
yHhsddyIqIyrGv38jbtoHWd6m3MxggM7LrSvH7/TnHPBacjpdvUZAfcgk5mX2sAD
/MJxPe2X0XRk5Otu6wmO68Fdc0bRZGDxeQVOjfVtP11/sYDZ99eoa2rfRrtqofAb
XYabkfe2N0e/moR3gsbsO9/OOVPxws0KJB6M7asMN5AraluHPYTscU1gOzcAA3OY
u3Trphen6aIpoLAFD9t9vfGmut9S6w9PThbNVD5VYzkKQoxzcOxgpDc/PqtZf71a
z+158WijsP7v7xL2jcHef7zlyHXq2xVDj4Lzitanbrj15gRuVXkDeYIIuBCm8dHE
Ayvi6BawTKSwvpdjz1VDx36+FTCzv72CYljH50uPEB0v80ML6voKY1nZ/Oq8fbb3
HGlTKpGpmXWkInqpO3V5Vc0AXiRenBIoggPEvkdKJtCyGHw9nyMVLLvpPqqXzc/N
+sk02ofb8FOT09tzhwF6SCKRAwvoUggpQiAPukJ6JqfvRtPQcTci+bVc/JcM9z/r
LM/VyJzCMvelJlMXwh8wYGHV53aOxEzQIMc+U1xtIUx/DXh9JURvIkKzM7bAiRXB
by9S2snyARbyneJIuo0tRTvdwDVAnl+FXz2NJ05oCEL/cvnWIqQKlQOeBO8J5FQa
d1ohLQ8x4ZUQZjkkk11sKouvuOa89L/HYCewXGhROTfajOLHTqBCEMdDxF/ebB4y
g5hCJA8TVSuy2VgbWL8lfvqccQmL3lewlGa5P2ChjfSOB8Ja+j//c7JQGnLZ01Qx
ZhFcFn/D+hLLQ0/ni3pAf3za+rCPSrYHbBzKvIvR68PErinxtg8ClDte4Nfthf+A
XVW9TwDrKZnaGU22S5Vzw07NEQ0CjEwr2X0U2DAGSrAQtE+ujFRlMY8qWFf4RQYX
WsL67jfg/cNY7tbq17EOqOw0sMFvUxoWj6vVcGkacMl2GB88phvgsDdDDT0VKw9p
sJEtiBHL4Grvog3Cf8HX2dgcwyyI3iS0YhavNQSIqPfpBepdkB/id133xFY3YMMv
qM2liFgbBdurJ/cXkkAa38XMlVYRpHcYJ1yt+s0ZNlmyW6l0XS9NmB+E1hS6hwmW
0mG+O0VgZLw62MmRKYHwGxaMLCssDP1efIaEfgGFRERC6FVeYVthC/dRwunec/cR
VdA8jMQoPbv7Pw9rQV2fVhrnsFN+EMtII7r1w1f8czRSPOUbnLTbRLLnGAWyqzNq
z2B+M1gU8z5jUnaRwov9RT6aotGtfrvXQFgxHLBE3LyGC7iqs2E5q9FySOnMSXvV
61T/iIYx29dT7gdKRn0JPAN5WHe1Yxm1V991OTEwNpu12Z5Ljgxn0HnO1HFwurrL
H4OXCykPx6WX+ExYbnXtkw5P451z5+Z6qaDD2uWDc2h8SENoXQRjolsNGsG3tc2s
Zp9IkqQRmMyWn0pnIKe6nkqVw+ts1J8dgoIMZz5a8vanLR+f6yJO1KQmAMp69Wi5
72s2kK7S6jY0dqwJXQVjrT3HkTvQUi8hzdzdbdLgUUEfr0Y/+tUa8qW3vIEgAz5O
+LiAOcj7vYNi2G1625Og/7gUppwJoAjxX9+eSb4ujInve28td1UGT7/TSANTrE/G
JZCm6BZvXV7hxGOiIeIbYOnOlBabFHrP6irn9ygHLDcKZzfGrWFfA66SNCbcrAxM
kPhNOlQhu3yHyfUfA52THX0VPfSkRD20n0/vhv187a+HvPJnCaEmJA9kvPkFnrg3
WV5ta8zOXa3p/REviDFHZ1BrWenYjpHbFbKRJjqduMfXksFecPWz3wsbMp4Xlf/G
nrP0JtK7clNryHUX79rgXWSbzlg21+v+eRxAE/8/acKARrLMgQ6twge8B04C7ait
mVCqg1WhfltxZM+uH2zNiEnBDeH9WuNSQUPB7VJOFPS/sGte3DwpMkbp1G3xa8B6
OyNRv6SxdFvh+uj8B5LJ+zJy/xE0PFx5EmrbB7bKHb6mS3fVlJZkLVBv6f+M9c1S
5rQIxIK1oXw7MD5mMsL1hmNorOHDCNJh85dCfCN83Wmv9siu/BjUyer84V4qfInY
cj1MCtrvtNxTXDAQPyMq40G8F7KRy2mfScTYy7c2heanFeUXT7fegmW/6bLmngMn
jB71dr39Esj9jN2TwGQiuy2frIDpoqsZgluqlBHI8/Mo53/LGo3OpC1h5ykJft3N
8qa3sWCwTf341MPITfof6XZXJ+p4/U4c1kPtFRe8nlO/COA6E9ZOd8qgqmyXLQDo
A7muHLW4kzjJiIg1frI2aXtotqYn/qYFnCvjCRJI+PFLE4CFtBfqpTNuNTWtMyf4
YzClugGcSOzJZiV73q0rlAZH0mI2smz8Lwcq9Nl3zLI9B4m78TEwbOqxCVTl1NwG
3U3W+xgmAepcDvmKnha915p2IdMYmJ+98yVE+bE/qy3YdcqOzvt3GwCV8vnLU6xp
WDSra1VOUKj8j1ooB4MAatSPciRtT76dbRARureaJuX2XdOm9RKKcUG/PXaYdliR
TduI2KAxD/pZTGbxn+JLGl/9R+yHu3ptn17H1Pvbmuxneynh6dnX9wThqgGR0ldp
HERcttJ4BaUxZkVVjsjS5PFNqt/agjiBNQTn3LWlEns90Wd8pHWzZQUHKGZnbyJV
4+x2rpwf4Ehv5zx9FEBqiMHsdnLmmgDNfZ+4FAshVCWu81svh18v9xkkUcTiwuJJ
99w+wjl3K6pUEZp/F2vS5hiUGkm+p2nFwXdjyGFqBmDlAIcfnwhSWGpXO2ba/sLE
U15WvkXA6146jTKhw6bQ0mpxV7y6NoRvmqT7oLwy+ODD24gs6snrlYddP9DcY4OB
mPssEe1LiImQ9i9E4C3RWCZCFSvW1qZpBS/iabvEGqgxxeXfiXm1B/vRXxI+tIiN
rCrTp5f3zcExqnIZX21CRgklFrL69aXOAs+++vlh9gv8pElNPwzmUhNhrq/3bxg1
kALMX21zfDSXJttRPlditsQsYswTKsCLzP+VRLpYjTgvvmVgqWsksUEvGsVNbJxI
8BAFme3kFwNqQ8WIRyzC6C+xug0tz9wcrRd29L7bCKy5+rK8mryy0KH98c/nzAWr
8M5OVN0uoOBDeodaKhm8yL2+nV/DLyyLBhpIl817tHlooY3T2HnwByK0JYhIpQYx
2hMfgMpjHQnQef+4rfMslsLZJ5CqfyXyzx27hO0IxcBE1Luk6owYlv1umpCUyDLF
MrSx2Tu8YVszQNPu8UoIczc0ZyAVyBhpHWDTFRpoNqO5Tft3ZVe6QC+u23Mw7mpX
ba9QvmpIKHRONw0RjnkzWuygUFFVJeqvPDmeitgdz1Tf0QFTwbLZ1fUSkqZQHg4C
VnLyMzrf0e9xhILjd4PPAdTcbKohaH2frGHe3Zbko523ak2CyNfgYYSxxndGly56
uBZYCLyCtXkK7ZUtHpdolEx1gnbrsqZ8PdjYURYmM6AX4+n/nOobE0MfF/uSgpFd
0PsZ/EaJwbVtO9CL2IVwI8oFtAOEPYMo51iDzS5vV0pldpY6TRql5uc6fvmzulaL
tl2hTUZw6wHencDPaUBVQTvhxa20/pmcYVFG5QCp0ogR2tkWEhQqtbAaSe0fbMZD
1hmTLBNpEtz0V72CyI6QpsVE9kxmL1vaC2vvH9u5ezoaJ4NQgb2bUR4p7GgnJf9o
/K+36IpWRiTcUlnY6TUM4EsF92sX5Gsf5HUkfo9l7Y7j+zCV+pWjmDbG07AV0jxp
jQW4EQKIMpcPLmhYF+w0r1Rmu1JmzWM3BDsMQ+43AKCCpyQ1D8+rDRzQOkov9DvV
TS6ZDJnoJqNHjIxJ0FVn1psErCg/gs5V1OprdSB8pqzNO40G/Ls/yS7H0k4QM0rd
15c/bERCT6YBk/OSOeBros3KLtVszEBxBJA6cGqVAj9C5hlTwAIkNoxuJnkMH9oZ
sExO6ROcIOaChnfIUInZSSq0imVbKztebVWEt9q+6RyoPMBvN8UrHaRVSl0V5dr2
mVJsiKSK5FRXWdNe+1c4elTHY4PySPJ+YTQDetg4j3qvOnC5bQAMKzg9QLIr4E/M
h6PwPPemuM6ndSD1BoJKf13/zbQ6rh0cfZgYxuAgcDpljjnlox+hT9oewSaO4Va2
mJdKQT5P1PhuqAaamAmQ7Qx64tGyqV0thUtZ6O1U0KU3fw+KRZ2wVUjVsegEu2sr
vH9PrEMlwzQCUajFCmZJBuHxMwCIJKbDei+SNTF41XA8ELqU2BRqttjz1GZPqsmY
xCrBzvo0Rpg53gpShGXi3EAKCwObegL/BcJdwfmst5y0nNtw++8jgNkutEzV79SI
/Saw/Y4JKqcGUZeYqi32ul6moKW6GqmKQX+byCnuN7e94d7xpwJ4SE4Y8ZGJbHGO
ezqvunSmOPhK26EzkF1oZMF9CdMcU6nj1bdaY6/nE7b3SjzInUKoAZ98U2uEmNt4
Ih6IaiHLfcDXkcY1yM6dTK3scjt6+MdI5ITCyz8eadh301SByvGo7D88zfK7AKmX
xFt95dkA3s8IUgQIbm+Om4OIvPOJuuPsN2XV+diwLsb+akfkExmhE0a2cD133mJ3
BlWMwb0KdNW0tRUHXnFZ7GNyGVPOAJJlFKbHm0t6X8jOts4Qt7FVR12HyDEiqpHC
PFKvB7Q0xwKELI4FJrQ2wdqQnRDimBtreVzP6Q7GJCMtgQY3tvFDFx7naD1rlh9c
9OsIIJ8WwmVcHpLSdzJmD7LwwEs7loDHE4hDXRvB0b0AAOLQJXxeZ7B5PwDqcU4d
4jicXP7/U1EQrvKAWZi2aMwE0Ibr7eDUM/BrUUzOytGCcdA6HYFMTTKaBCENcSg3
twNsEAM5pbFHkEaO37H4SxFQKBgcdC9pN9dY/v4NwEAklGFWcjk6msaUfZFl9qKY
bNEN6o24OzTQa5lCOuCo1vBivaj+QV9SNWXYo7G4VZodGTQ4egnpJlS5PtSd5NZH
38YJf1POxydzJ/m0IOQ6EkdUvfbbjrcDJ51E5m4umJ+GUvPw6ZEHCKBg3uzd2OkF
pr5b/NiwVZ4KHvh4oaQ45XYwUhinhf/2LSjpO1u7vaFWloGIVQnyU6ZbDLbgcbL0
3hXs8RDqtR4IlQMVjIiU+JWT6aknf3R0y5Vs4c8XnpII7QE/bCe3YdCVpgyHtdRY
5iMop3UXR1MM8TtRWdS2Whl3LWYpi3CKxvPl9uUSWWklQqAKegPF3aNSDp30UqQ7
2MjI0vaNZaC2Fhy8DfFBWZuJPrgVMPWLqNr0YirEkLE0ZUQagaqmm87DdGpp6KFS
JnhPIPgNY7LWyOJyrWOYbkCeTr4l5eP5G+XQqklGVkD57xHPBIhOFLoJPBPztf7c
48bAEX8+g6+qFcG9yy8JCA5Ntqn71BNtlgT7XuQ1SM5nhlEYE77kBGXmx0z+/+83
HRCxOtxbyOw+rOaBqbWJBLnX/WugFwOT7Vhl/J66Gl04Y4LOw93m7dggpza8BuJE
LfJWsKKfgDEo45Eje1JL0+vnbU13vnT1LSqkk61XUiLyj/iYeAPuZKJvzefT0WUg
Y2ICNS5Zpf5hjcq+FCwRUmRiq043zOrcMAgFAOSFnjDTq5q/XdXjgqyARTx+yLab
v0riHtFXKh8dFT2UqZJdQEdIIStCpxt+sxJR3tV6PjGCy558cp2C3HClW0w3m1Fd
fFQ/fa4eeJFjIvysLcywbjRIH4IQ/3h/+eA7+L9/sCq2ta167jOIa1ybsUKp4Kdm
E5nyKN9Jlixt3Is1cFvT5wSrOg8iFZkPAMt2fT5ik4g7bputwTGuoumwm31ZM6pu
uNTdDtU6TJust7lkJbKhHenARF/SCxuOjdMdQ9lxtHjdJTwobrC4TOSAAIxKWOgc
ePV03Xcx3ubt4AZCPCz/tgxvBI0PTRsuNoRL5dfsQTQpIRrRcI4swQofk7T/bBmm
SLMYI40pHXoe7jVXECqnjfnf1pa5lG0POU3Xp8GNgNCyZe+EGxvBakYwXzDshH38
TJnKc1iFA1NWm0hfVhQL0vZ2kZp7YU2gZo56GkYYb5UM53eorQodl0LwFByizhaW
MZJaaxSck4v6N/8QMZRngtjxBmk/r+2cQr9W5PG+a1re2sRnGTLNe7knXmlJIt1O
YoKiXrjB6lCBTg0F265KAhf37II/eOmdWVpGJTuU1EPCfEt8vcLllVLswXuLco8k
Sw/zUsHnC7rGXeTsFADGDAUFrwXh5yrjNdCMA6h1ecdrMZulpq3s5g9eITVcBCtq
FWIsqVmkJdOMMcfs7AfdtHspWEdkwa5td+Fi88LgiM6azMD2FPE4knEZVE0tGBRR
CjRhmzsh8dDVv0aS9F+vpSQupLKk0fAYD7KPxmQ4QXVTgL1TVYiA+fEG5DdAqJ91
yX13H30/odhMRkHrCbif9X16PoR7LK529dN3Gji6oYMRanSH4zX9ZHAwAVADIuUL
6GzXphEEDUxmHNpsJz/G7oVsT+E3wA8IBtlvtYY9ECakYNLY2B6/e32/qY/a7Eb1
2xo3hdvVzUAWTr6N9kbzryOVoQr9lBVPq3lP0VBco8C05KJ7tMB5F1sCWnv7G8XN
NHiSnK4LDTX4bTwQSlqg8XpP1DfYSo8WKO0fXoPZF09U9JvHuyjUXreNmJk5//1h
T4rGj1+wIGrlRXMGG2EX672GxKIOkzwsAce1QAAigUDzCxfW7vcHCppVRLGZ+JUX
3s5Uy20SmKan9r0rv/bepuo3koFk6zON2l/yfqjZGmJAAVZJr3VPWinpkPerE4T3
4HoCAPUFWy2dPKkSYVt9CTL0i9RzKmONXxVnQYhagz2aGYx0BhiMcbhtHyjZW+tp
hKGWAjezlTqla9n4qZAQNQv6kGbxwtRWmpLA741AnkElohdEjkaFQcFJpuKZzBWI
Dp0N4/LcrDSXN5RMfq4vrFY+1xA1cFfOVyvdUk9tPQ3f9kIdkEZTDUn9bcKfnvhN
FZklue5hxBjbpJsitXvjXVvjjEYNRiwzhocP23LlYeI5ytej7uJ2JkMDUybJfEsm
rVZQcQLHY+0J0jaB9KBTgV+/QWnuOSgOZ9xMJFOWNi6YMzpZkpWlI4vU/BEU1zuG
FeNeZF9vZr6acF3pWgE52Ys12Kt2++KAy5nH9vXqVEj1u9SZYgbrYgar7T2zo0jM
8aN+7iDwvV5jioskOHuYFZcQcKDQ57KBRAPf09DljxZNNMus2+ujsLwSMPW7FfWl
ChfV4BfHrbNAH5gGtooDDMPxVbaVDcbcklmz1TWrFSjkNyd4dbG3LFBdqXDE1uBu
Puv4EsfD2gWnES10RJO+u1udvU7Arsmp4bsjNCsYNXZ4Tt5/JNRkYzlrAGUh6ouu
v6ary5uSYJa/hVEqUOUMHmAbL7Mx1v62ulo0/knNl5g4lFKzpJCfQhGEIJ4FelXe
3hKCkelMagdNQIMO/duQM3uSeC0TKu7TFDVI74ul36O/6kDttYlAW7koyavLBWqb
lANWoGe9IqLae5ys5jSrjCgvIBvOvjNK5rK65ZHhKZR+jsGZcF0Ei2jQmTzVI3gy
GsT05sg0Tt9sr5eQHCUQ51Op42ShFIgoUz/yiNOKp946zDFgTcgPxdN0reqKl+B8
61w9vIeYObYuD9s3cCF1Vt6RfZuvZynLnWWgOGpjVl0+jG4KBxhGbPOx36uNSQQa
vKovr7ib2LM01UXyJD8fbUAhnK1Rfx3Y+InYIE0J5Ha00FlSh2DIvLHbrdJn1Lcm
Q8cgE8FjCJZaqNV5mXJ89bgVycnLDxUGYASaG44r989RuiC2x0vv2twUHOa9MNF3
nVaMHrmxJBBhwfDmg9bR0G0zDuR0B404VEBD0iZqyjMGHkWChve+4AZcm7d6YzIL
dXm8xNprM//ziqd28h8qHkvsW7P0hCXlOEu+CIn7OWc+vvPACM4SdoDtH9xe6Mt6
d2RVVz4REsPKUrdewlxYpZkzX1Ley3ylkUePZNVsJCVbbUivHkrY3tOtFzsyZdXv
niEdJ09IE9qUdPS77Z7s9hTin8Y1ouCLaQ2xBs/VGDONAjZaNQVB8crBPMASEiiV
4LvMwvsQfTG5ZUQqCi5mC1Iy9UGFz/vv1ODmoTMhxtAV4TNVfBH8hCcgXIFd6ofJ
owCUBGVYTOrtv/j6B8vLmwJQI7hiGwNmTrbkm+oRhz2a/jt8IXqsUwWp86VW82p8
5zHBM4fCDyPGIISBMzJ1zVzCLwFWIHJxfL80aUtcVNP/OqcDS1RjYN8s+PJjU06I
7cePHupufemLmYUvpFzkT1rzD0L0QRiiWfmDNCYAP2qvy3p2p34fBHGvM8K3N3u/
czhMiO+2jsGGPqUwhcc84XN1WJgpqlaxhkwYwJg1NNQTPuzVTlDViTJqCygM/v7I
qnMwomT2+5QfOPaT0kalSy+Jyd3/CNtmSR/hCN7nMwVxSmRnG/VfIJjEhzyDzLP2
nkkx05paL0yeZ665INfaoVOYojZxc8m9h+vIXA6beilURiSn+fSjBQJBoAS0m3gw
pFChK86x43VNLyC6pWmfU9do67REFvIk61WboJaWu9/mfdG100CoQJIJ0RijsuPu
hAYLAWPr5QCKBwY0CnU9JDnFp2xam1lqj4MPpihMSJ+xabtoRqI4PCp1z626fxX8
NQ/X3xVq2SX3E/KP9egAJ2V9t0iW4VUUhZ8JltzfGQTN13ZycGh0/R5AZ/JrPlM7
d9H+aR7a8rModwxy04eXszOKASS0lQyDwLWT/6Q3dq0X3fMT41nQGjsD6QKgT/B7
iZRwHDi6v+drqYpt385NjHhXotqRsgMlwseW5zXGxQzvVF92Qny7bX8AI9Ub7gtV
xWmnJ48/E+J1A8prCs9TVgq383dYNXp8nxu0OHWBIQiItpMZ4i439BiyJmF+KkQj
Y8sdzaT3jWiGbJ/dQrSzdAT8M/Tn/pFtwKMXtSofhRgwvejlMIthCohuFKrPX4Rw
gjX1SG2tVxJRHaeu1fe38RZSo8fJjPZZ58gBtWXrPRPjBgQHATkzfInh0siP5zds
H7+QcFbbIRtIy8AHdpYdhadGK5iMdIAUCKwyduC2hZnegdDsSU4je0BMILJLwopP
29IPEuvPYsXG+ieCgwZsSvQzWt3wppm4NYI7Ak1cQiNukV8WuxO+QfIf/z/RDfP/
xr6kJ32ger51VzO5MJ5Glr0IrMJkpv2TKbJ6UdEQ63671ZMi7aC9yn0dlPMhAay1
QV0C/lVLjnWLJ3QNbEiosqVVMNjIKGUebzbHjIGSSEGtlmm8cvjtxQqaQGNFHW6G
wyiP40uGS456buffQP0NhhW41anKjjbWN5fcYjTLNhA95XiPwVjf0n3GnAD1DWUB
Sfev4uIhdMBMfFoBT9oaBGlc0+EnxdqRjEyqUYDqpOcNIHA2HHQt3mDktQuFNPin
5G8YHDY3Q1+C677QZIjnQmjyONJgQZMLXaf1gHJDjNepywORdwGcnXe92GXRgy1h
YyUg3l8rca3HkfuWQgrVO45zgR6A2SQXvOzRGxvI8zDf2IRL6nG9nB87PTBCyEb7
9toz3hAeZaFfnhXuSVLuCOC1Nq3LxyF5pAQysBg4ZkURW5rKtqj35a+uH/kC2Y6l
U/Jj42pLhw1hgdInbeLRiIx8ZgciHfAU002Kj5ub43TOTkmI1n8G0IRMjKWIs4dp
OTNKoTCa47j90xUIYrpNicSTCIYXCGf9je+U3PBn9Ak+zTi8kb2GVoxguQzLYA2t
EydiHpZJ5FCzeXLQ5T0S4PSY0HAjP9tyGUsB3Y9U1hH7k0dLj4J1H+Edu/cqUf92
rL4oljmNPwoSA6TuhTGqyoGEeCSA3s9850gLHl2jEUxnrSmwuUH0NP5Gv66ta+gk
T7j6phGbsAYRrz+wYGX3SletVDlgA1+UT1O7HZJp1fX3wXISJJlRGW6wdoLiOkK2
sfvhrfrSIZd38EgOjHst07EKQ2dLVKOMDJ/aMbikKxrsEw/UVNi8oNlJpkaq/Dya
g/T2ERr9rf8uNTBMwCZvS8TDj+unBd3wrQbW4s/XWGbQDI56/eGwFA4tUIZgVOcx
62Ids8OtH0PFVIrpnDPXsuivIC2yTQiO8XNnyxZsILp5Jk1YfqUQaT9MRCslqEjZ
2WJ5itC2lf6UN2SqYVjo5R9KWlU+d3ItBvaxSf46GGrcllAdc2uWxkKV7xtdQhB3
cv618YSclaliGQe+UpzWts8X47+zQ5intYZ8K6EoUbXy74LEjiAwhidXwb5aI6u1
f1TZMQwOYDqzLd6r+88dE7YtMlQOqJJpsGHBElqzuN7pv9pws0xmuWEh9x1fYmHp
/J/IyyFrfIHDKyuXfFZRlrSyPg71EqH5ViIXIPgvEDNIZeA5BOXzJxdUpuVNz6+M
1kDhEJZ04/CWz3FnHw0FN2p1K0NJDYmwhtbrElLlxNR/xnb4Dk9VFBMyA9x28yix
2KSulLK3bztucILxo7ROH71eJYWrGUXeAN/hIc1EG1mI72Eyens91GWXApb3XeCn
VSDYKKIHaM5gtplOlSaILSLkW6fkcBh/CSJOyQSYS2SdaL5WHCrvlhXkDu77uJP0
rcjhrtwvzrUVQZFd9DOGrox4KJy9GwKGIiak/XKGuIU0HFB/8SZpVX/9oJdLgazQ
CbyNWXwAhYl2h969m7kbBXcCATn45PKCu1gpMAmJh8u2jHj910UvBzAihPT4cSU+
GYVpTkCsWP8owSc1zoZW3GmQ2r9hUttoZZw67dBioQVlXdRkydRran8dWip2QwuP
31TlvB8sT/NfVR/YlYm3Ftmg/d/jBv8JTMrOvR+VDN4UGWpJdQ4nmMLGhmr5J4RD
00akMJC9k9v6UnIK3yY2yYD7elTBWvEJ6aUntOteNT9fwit70lGAaBl044l3VOIL
uHiJQTsQ0bOmho9M/VlJhsrG/pqwUWq1OtIVfFrUVeCzOX8uMHzR0n+7mfctUGG6
xKAdQbpP0vIVEvotEj9gn8d1KCQXnVGU6XzTqt06o0NDLru9d7P8uZ8YJMmBDXXu
yl4NgkEi09ZxQsqvrQc3dxkgbKTPxf7FA/+T4tFYTcB1rz+TAjfBgXLILj3LFwse
B/Kgo4Asfm+XODIcvpSv1rDmObLX47rGyuuIYJrx9Ht943RoaRK1Bsr48qrK0t/B
Mzuk7Qaf3Df6wdyIPP8lL7ijszWyglFcm1kMjam2CL6s+nbNE8UMZ3nJNiZdBZtF
Rm19lXbpCGz4iFl2YTEGEW+prL5mrQIlJdtgj09JJhw816Fc6mCftHwMTHxE8oN3
aafBPw0ox/fLGBwT9qT8HFRvczizsxN7AszBzIoJh36AAIPV8WTPVhEV6H7xO/AR
E6RDXSudcqfCNYAF7/IZItQ+/bqTi4UN6O/UW7xigMSpRLvUaojcIonTwJ7XVcER
0f8lZUIX4jbtnyCiqW420QUM/FcF00IA6kaSFGoEovq7fbMazhhtoYTz4bOV97lY
KyADcSRAZHIIZKR/Ng8OXZN4IjHXA7MAi0wDer0OsSXNsZoJpVeL/ZHzo+p4+odC
tbqXfuZ4lD5/S+MWlfpblXybveDTZHQoh5JrYCSTQQDOZcctDVzcPlJsfhKYXIg2
hI0DNStXhvGbTrnEe/hqpNIj1CjsfjeSwgksQBa+OngFQWED7ETtq8pkXPHrOic9
AHMb5zzMdN/xRzd6TLQpM/q6EhQTLFXSZxgs0FLuldxEccWeSZSVBnRcViaTg+fk
1bpeSD33beU9sPQErCjTl6CvnfppkGNBBEYb0TWksSE5yhNhq6409hVxLzxnZtDB
XxuF92jkeW1vvFqR+NXjYhQ6EPi8MyonBl13BrV8bBno1F3IqWpHnAsVQN4o09aO
SKquqHdc3ROQoI9BWT4C5DyrWfKEZMXhSbu8Y/GFEas41HoFF1reDGBoTMsurT+9
z+H4zU4ilHPUKk1kAIPhkombxAYQoJSLaa31zDQLNvmgLTKRmxgmEMWoE+OFN4LX
0lgCfM+/76XnDFEGmyma6mHZc2fiSrLkQHwLuzmJTBfd3+Vf+kyGU1HIVuX6PbmY
0LC9Pb7LQubiBWSk4iEIvFuyhUaTo/JPWtFZZqLtPramL0Yw890OowMQ2k4hDeh+
obbFg9BzZe6ju1edVfjMpCCE6Urr50bJeDxB3IzdgbQR7AitwFEyMBXZBqqWhloQ
iKRrCWa13052DYzfjvzoOaBh0q0kGm2MMjcPQ8EUQnb4hITEqKTmfk2YNCjM1+O9
IbGSGB1qnAaRA7CP99/6NoLmxkceBG8HuZ1bKA57QlAaeMqx0lPJxXDvoMwxJy3d
gLdScjfXqA/GmoVlIHcBEfRqjc4+pEdXx3XSj2Ei3WM8usKZbSZJGNUg2OMsw+uN
ARWbF6gSdy8koT50kWOpUTCGAzi5vNAqfGGVjIX8aXlA8HLCSqTONkJrK2hxQZ0W
7AqdME1PZAWZZWgxZmrSyZTnOQDo9AnkNDp5vZxWzQHMNZV2skohin8fWWgRfsYK
OxdrLZeWu2yNyNCBqdHrbp9Lshoeko+/07YIbTDmSEXsTRUwGKYs3Wfm61cwW1no
Wk1HS96Unbs90Z/Isn5zdHYm3IMwW3rn6YYXhLQIXO6SDIhnutQjZ4alyCxm18A5
U1Ojii+gkxCMCDSUnAeMGxMBYHbE3cUCX8rOETCoZAILNqOFkuQfQk69kA0VvwPs
ycRMzNRoG9zUPlAExMLrGDIzjHIMsdBzua17Z4b6vsRNnZ6/S3TdJsib7me598EM
y2cucTZKTodiWnuFrjGig1G7TyW6+zcNrNI4FoYXnx/hZEDhhHblrXwLofpDxW4w
TR1OFk0oMX5Vivc5M8UjGMVyWhDTF9jV+A1asbz2kbsKdE9XZRrM/um/tbYm+uqN
K+Jxje6KdwR2wg197N2pmFeTA0NbHL0ZbPyvFbctvFKqtzhSjXHz/jPmP5b6WRPK
Z0n5NCBh5LHPDWZCZJbg3aaGskRW9QbpKJblkLjPtdu2HrOEWRn9+NiWjwtxOCGe
zc0dBAxtP2ovKnnHEQ04QYbtrVcYtbQKv0Tf8htqdx2b9Aan+q1mvanrbMBwdamm
twFNB4uYO7A9tJkRcAdO1ZLc3PMTVeNiRRvI82efFut95L7ulXDC7PuhEMrRVpIy
z13TkVrnFMXHfUS7DHIhf5iH+6cmJIF8kRY4YRY3bS0ZuK6W6+dRXoazFe5BKddu
wn20UVF/zfEPktvYGNExsFLEK0G6yQqEW3bF45URlhF4mv6/t0/SJ3I8WR8UH/XA
xe4YRneJ/2yYNQHXOkzTHODStGi/ZbpIbc5lUsqb6oEcqla9T7QAG1LpwErSAyg7
cEFapGeHq3f7A/YyYIZZ0+LJhnDJEALDWgIVvBx5ulRrqGCc5GE6kkapj5mVZlkU
JeIpshNST4lP0SBpHax00ZiVWFqk4xZNbcXBJxwbnm8iHDajFIuZOuKzSAX5+3cl
WiP7Kh3w5cRH+P3Dxf6WmTx+sDBN5bDXTGVGEXZxC/hlvcmpCbNtv2uegpvHZvyG
4nU33uvm8uY3DbYINXTsTj/UHHbMMFUhZ9Aofcrf8KzqPkF9yOb8e3IsOHaz5FZr
wBv57lhlTcG3LEEvIwHDRm+tYn2clAgrhhWemIUiyv82qj7Cru7/zItXgsCTc1lO
OUjy7XeVRIVY4nxY49UYAcSDKh9cc2Nz3YWHyx8McuD+4a/rTgxcFGy96GzwD6qC
dj1zZimB3h8notFw7m0QOKVSUsGOhwbWwcB6P9CVgRdSrlDK/ulJOdq9nRTBMSQA
Hiwvun8XsmH4eVHu/5S+Z7Ouaz0cJEoDI7llkVnobcEGoMdAsmV1aRrkDBVnIpPt
BLqH7TvLYYDKB4meLkWgGlz7duXBszGU3fWH5y++3gsM86wNv42RN1LUh2ZZp7Y7
vMfjp7x9VzxIXCQgvVa7cqe1Gu6MmBi/ynZWCusaGRX79WHA/A4K0l4f5x88ABfe
KfDfnA0TA14Thf0UdWsEpuifv6jZx95ibQKft9YDYLh4lyx/OomDgwmpj75SmKWM
eMmUa/ITrMZEqS3hrdgNCIo6k5CP9fyiEA7/1P7iqaVDU8STp2LNKnuOpmhJAig3
e8CdRCGuysNzOvuD3zwu8HGhsotsr6KsCH+SNWMzPswGN3kTStDTrnxYdLHklL7g
X3AWK+92YNssrIBRre15xUUnLS5qtm9YMWheeQuPiAZQG6TZNGdCDGNBDQHcnfsR
t7jwo8jSYevBDHqbA9xv3Tt4+feUEOXxuQSVF/nrUx8WenTCCgUB+4iUni4T90/K
bstOL+kxAQI49amsty7UtYYPi4Rvim76qkSM4Sl9ThwLETLdLnPIWCA/E4fSP+jH
ZTu+iz9AlhBNvWif0m7eQr0TvgUbElYM+9n1UQZjkwScGlyatoLs4CJe1I0dJcl+
QXDlqRpDmagQwcF+2E6NCTrCIRmG7Ozz2bTn+f0h6H9HbtYjcq/uMuNLysAZ9H1M
mE3ELKZdER2JUK8R6TJB1XFEMmp9ScPx5CAX1IxZmhiIO77Kg9Fb7NYxEsFzxai9
gNeND5+7IQ0OpXPCKWWyvhOFHJhA7hgOk65sUObvz9ZljkIojQyMdxnSiKAYWj4n
vkGLzPRzN6mkHUjxeXdmPaACbVmSu+abpU0TKg5bpDqjWZD2NwrVfAsOceNmDSOl
+7FesVIiLUrio5fFjJxcy5MHXXInq4OyZvlgPlil3bpTfcRa8sag6xcqRvE8N6eO
dvlX43+rQ4z9ev2/mMxllZISPwrMW7r2EiAHh0VW2b3Ih0c+6d3kB7MbNIkmNUhq
yXZGGP5scjYAyqDR9uPzhvMG2fv3DLJupqzZopFM/zYQ5INoHSvPQHLyR5z1mLRP
pnR/ltpo58lnkyzlm9Sv84clZMS+UuA/+SO4ApHLcJWm2yNHUIlNWJUpFqjR5587
QEjzCxkilqLv4Fp68Xc5RvME9azITSdNw5EXRtDk9zUtK90twM6gan1tw8SkjIeQ
8K8bXwcU0sqWSSIgcjO6kpdRgxRrb9KqlUkhs/xwEYXir94/dtxpdoE2Jz+aAGYh
nekKEN7V+R6SoiPukO/svMd85RMTfvpCfPyErRItd0whrx4+IK0KLNVj3x7zrDLh
7LCBsVJ1yL91V3Fgv1HpwiZElCRONECQ21FDuxnUTGLOfItvSEEWylxU4cyTDeqq
dp+bwqy0X3U1tPWcPMC5KRMy1TZ599KqWBvE/VB4W8os4Za7k4B516U3pneArUyV
/jzLYNcaS3T5QVgl3admPE0y6W0IfIag5gs0SQUrsRNj6exXQOfNfljbM+aVdvdV
j/SUm45LIrfxNaYwPvAy7qh7yja9a5g4xekGXV0sr4/S96G6pm3Zgu0JRo6GGWMA
xdN6Vck+ys0jwbMEuo3ehpNsYJA/SbFnK5GmSZVifYvsrI56NQ4lZf4OBW1aQArn
+0M2T6i6YKqqIrwgZYUiWBH+fR+nWcEJ2htda/0VWNYvbwf/qo0eHFxL4H9Iy/tn
FVnX8qGI9PhEtyWb0+AU1hSXx7D4iZT3Hkz8XpvIGI082VGK5GtJ08kflIr7oiKC
VCUG8g+kFSXKEma6sa7US6kbL6qk9YHMlhQ+Xg1EmHC4QszRYCbtF9V/PusSafUs
YYT+Aj77oE4f9NtbQMDoRAJC4u2AykhFp/iwCQsE/E/gDHU0upOfDlbM4xoUOVZR
YeN3i+mHqQIC6SSvroAcalHfOZ6esrN/u/RIjpsZECHxXkj0lfDxDRzz94hCDKR/
Q+g193cTKm1fm+K0DA1staItd3JXXXC2s6oCd4uB5SoY/6NZ09OqjddeWN+OjQQf
WVJaYhkgXD/d0N3cEEA9tKFk0oAfb6NYVjTVdP6FssWzqbGkIfn1KydWtsOoio/N
rR4BJvzx6csWnuCc8AqlkUIDeUppGadAZB2HYZsPxynthcEAMIdhnpGatEPNyqet
/2EgA45DC4cFawBbihuY7IlCWNCqIsr9dAfPz9m2Brz2Hfk4m7ZlCQ993M6y0BAI
ofR2M9L0P4CltY0xnMbu8QrQkZvePeD2DAUjcYsAj3fONukwMayZogy1GO4A3jte
WQW9CoRLbpE2MaV2KnY4A6hHv5PLDbRypZRExtr2gALEw/c851i2R1dS0ePbqvu/
xG5DnZkOhQ8Liz1OCoSBj/nXv37QGm+xr2kJvEJB/pYrd/TdIAAoGvGXeD2++by9
VsTUAp7kMoFC/+lcTQCdS9P3gKV0r8nmQzuM6SrLoVJz59iGMLHoNm9cazuWqFTy
j54fwB2qMA2xQGL19GzzSQCn3lfl/vDXCq7T6vfpSvBM7sVpj2xNnwNrJV1XFqL6
4zlPJM2kDRROdSH8EFY8WBJhRnB1tkmEEMeyf/ooBdBixm+j9UNTM+DIXBbky+kY
3F9z0MsNUobtnE0ZYMklX6caUZJTLemD5iY7KXs46LECIdGcvp5IQBY0rPik7c/5
aIA/a80HLXM+gH7KaGsLenjwSy5YPRRE8z2kPdPBXcmc5iMkqbKBFg08vb3+xBA9
TG+Uet49p2VnoxCGd8Cx0kHFhzgdJyirbEyooDZNjpxb0Iln4YznJEF/YgeM7tau
8PYkca4p0UdCUBNQ5/MigZGcWsM0LIrchV1Cr8ffvF+o56gMh5mMFPOPC/9XXVE2
/hEn0GI5FSpgN5CUC+i5vozJR/wxEMcnX7dzbh1GkLzWfrKmcshItw1i7cRgkpgp
Za+Rg3IEHnmw8JEHiMl613bN1rYwDGyfln7TD9l+Jv0XKTiQ0tO5NsJahYqc7rnn
S6ZFCLB9bx50GEAKY+3IZAnuloQ+t7SyyC+Lsq3PUmmynkfxCsuczxUNGZzSYW+P
wYhbdxfZc36ljHlF9cD2TnUcEBCuKov0AWYto+RN20C/1cMVumqodI8/uSN0CsQA
ElGQGLrBAZG59e7qMhazijOAAtjcOmyN9KxAGmEtGXq9UqsFhiln41Va+tLsrAVA
CX/TnH1NPeHqFKnrdkisQD2+DAf1IC8MU0k8xyfRbkiFOIhIOO4ugrIMrmHK7rFt
qb6QrZIWnv7rHMLLQA+CIi5jS7soT8tj2SICl4C3CFnvS8MnU5IMsEzdr+LRsPqp
BpltYvRLMnta8R7nmCuwIZeA/a5moRMscs70H1iak/Nsnpa6AeUSMH0LE1J5s1MV
TbSgmlSWcwj+Qu8iGbuXgv8TiT0mxLNFwvSVFY7uG2/+fs2TxlSvxROu7/L1uDzL
C3yvAXzVjt8hIhhXWb1aKuF7PRcTnOWtoyKKGujxR6CcRZxrbVAb2lCZXe0X9WFl
EGFTSMAoIQAD/ejH5Z1E7JGJjUwZ4ytG/V4X4XnK/6YNdPPHGuLC/1+B5F+5uETh
lz94Ae/O8/Chxs2YOYgDktMH3I2rfEkCONNEipnR7UsMBrsIlAaaE1r/5WkAeGz5
+aPNZOZHDHgZp/M6dAk+k9sDxll9mtuSfuZUDSD2eZhmuToAsiocKl2X0lJ5V6vu
JOE+PP2O328bJMGIa69m2ltei+L+ET+nPuHwl6dANf//l3MCpuGNdYLd4vv3d6mx
DSR7BpASx4kAWtsR6bYeX4ZiA0lBeC83DZBbnN+WizAx/sxhQD+HpA+HQfcRxWLX
ChNnm5GVXnaChCYV33TbYa2PjJwmPMfl35u6Glp3Yr1KBir70V+5svoTvWJnQkwb
gwR3S9OLA8wqgm/qt26Qs/cjzyUfbjIQDc36ZtyTEGoV8ckRLFmcezbfSZ1A6WFe
38o4AAPEXAXgqbWBkDeVfuHvcPe2WKFVI2dkxM1LrwExBK8Wt6dE2Of/5M6Yp4rg
AgAf+iDJPpRfLc2tf4fDu7hINKr7rHKTzskYpuEdNN9wMKykpZ31m6sXajwdZGdz
ukaIAVNahuEZB//n+fEqmHXl88IRcgHwSPyNKnZYzDxOtwen98+fKCTJkZvPQOsg
DI6BFbgzGKBKWrRoByGj1KMKx4r1qBHx3r2BsnItUqGPVmKtM23VOkgmsHaAkK+r
S/FJLotPApXkU96bJ/Ep0eG6st7DIqQwhc40X5Ha6BdO3lmAkpwVpGWzBKwRcy3t
IZpipK0Ybv7biTKwlwBhH5GaGx6xLskSHYkNtDV0FWJ6EHj5IZ3lqxbvfJA+P6Ul
+kRLl3DApua1pD2uEPemHYiqFRmnoNmWisLiF7c6JblyWLCp1W9cXNmaSMyYGVPO
tusdBwLlG/AKzNEOHF+MbX0fmxQzXBz91/kH5z1MrgRg/e/ge5ZadT71X6NO5Jci
gYAnx44n8FfRZ8gtcmkQCK/nGFN38hAx/jaRQF56Fmwq7H7k9pyboOcrEqT4vg89
7rtAnIXDqcRsVHurqDAlSukZAYKT08j9zujrS01yVgn7Ojb9YgsrhIQfscmu43GX
EzldFhANMzEvKN0uLvOTJb/V5kLDnAJg5+GktqPY6qKwXGYmPoB3c0wEKXRV/3dg
9iCYxEwbp+IjQJ+naTVuNfFQFR3QohpNCfOWCPoxaQ4owUJ5OrWduij3gVqXQK8r
Am67d+3UNvRUzOJOWrfkQEaV+dDVbnYHkOBJqDAFNQ/AjfVb/nvc3YijQK7sodTl
zQF2fOseP/xq5e5tl20w9hKtdSAeUdYdd3K/nOp5jnRCROtfWfzlWUnWcfgQYcaW
lPi7DegzHThL0iLglmM8d2iAk1cJ45q7H5OmzIdzxIgCHCzJeXOMNauLOrZmMTKw
PF8CiHbieudiilgvuEMYr37t8Hh6GDkJV8Jd/YEpk2kYRvZUL02jh0rokhsfGu1t
Lm+bYaKngk4KjTQV7R4Bs8YgrhKUU1wzu5ow+/9eh4HXl5ePdtoaxoLSURVqucci
rM/9/KpnLDVAGsY5i5Z1K/xuMi3eGmfvZ8nqHn1wIK3zgFKCuYm8hHQT5V0/ftae
L330dOeAJgT6zHdePfG8y+0uCb2XLaEJ0CDn21TyoS8NZ1vFW3RNaTL9nns8kwkI
dFaWiZkMcE41l8FHqzv3GMA+ypiuM1hKMnOEdYZF3Yhyhtzn0QixqRfkZMGU+sKV
3LdiAgBFjr80GFt4YJ0YGB5FLT03EAc3cjMFA07+HYpe0o6sUlKvGVuLXBf93JeB
jrhOEubGnRXeMW7s8u+/sk45vsThSPLvpGRpAAEZkO9wwGh77MLtWqdXjNFikibC
FpSnAyiD7KvAakiC8zOZTtuznzmjL68E6uoD/a2/mEzwb9gv3rcPo8PfY2ds6mqo
dCjwSt/EphdDsmNQRtUElNrWqaeDOPoD+NP+HBbuKfqWaaTpoJ5EOHTkv0Exfd5I
DB4mAcaprPfjWzxE+XNA9PxeRZYKuABvXTT0izBiNV+UcQXFQxksuvO+hW6Paeo1
+cV9XKeX1hvIWFojLNFUjaXzvb4sFzwvfCGZQeasEP6vsU0pdtexy/DKtKRawipU
G1j/Ro36qGPO0YHVkt0UcZX0yXVtqsTFia3YDTsLkezRaMo2VK0mZ/OurEBgUixZ
mqAdY1qsm0Uiy5F5wy+oTY2bY4sHCYoxMlaB7+1rRxGDaM33grLBZm3Y/LK79SiJ
uCD7mFsYdPN8X5BwoMMs6X04rcXgtLiAISB0eMwXagJqdJ2AKHlNH6+p9//ScjVs
hD/VpWFREI2gYYYKTUq3RxDOTad+BOSOETmKl/hhNQkqq7GKxzAsSV0KhyQ6tbJT
m9aBH3ic+8Ew9P5w6K1uG6HnvW9FKbZPiCheuu6uXcVSjmwy/nzTVm22kG5IDEhP
2WzT2mrdZ4ysLGPXwsGpiHN0F/M76ZB7SUOeo+Lm3mlekZ9qiKbpAd73AX4pKqkF
Rv02fN0c9BjBgbfhq/yOSwUzMt3PRdX7ha/22T3CTlsW3JNxlnWOSnWsRQUaP0Ft
zmpwP/fBRpvGYWW4FfbzycRa4RnEoRQlVWaoS0VJTfLvHI8KJPcw4QQHNtvWeFmd
+nO8g1pfCliqQ7tNNtnbaXgHg2SxM5vaD6pqbhu/pWU83JMGaqAK8FMH0SNy5LQu
28EZJPJl6FEjioLAQ/4JkCzvEysS4Wz+DPCwhTNB6PAIFfViObUwKGB4HJrx7zYq
ZtGKpHOPBozS34DvwQ3GR+gI0vcxVHGuV1ehrzzDisX37JFJGXYp2tq4/EZ4PZo8
Wm28bDPvXaDId7ozRqMJHghTkr7/fOPgF2aEzVPxp3kp8oolYEPgpuZuPp+3puS/
1EJaiip+V22Z0FGMgxrL3cXsP97V3y+ACX6Tm7O8pTcnh1YzJ3AGUa/0mfl29g83
NNV5cyiUmQpu0BAYi0x7nt4odrolQ/+FCi7/CIAc80q8fmvT/gx4OsxmiBXemITS
8Og8dlDfLozkFmwLr2FdLYJYkXCLf4jX0MJ6BaD9OBZYw8cxV05ZUX/XlDNZ5AG9
TrJf3OVDbh/yBe3WjNQOUVWebKsJ6XZ/CkWPL9D7UOSitCQjaZclL+nhXnTCRxYU
w1NCCe9luvdVRb8k3khp6vQqoMawRAIkTXRYNuJs1pnwax2rhTVS57M3ClKd+pAq
nydI8I5UuDnTZ8KuBRFPKkxRSE+aYUzEOJUO+BxCnQCoxVoYpJ/ouJhAKvgtDZWS
BEFOXupMrahxSrOb7iI/XlYwFXxoTjVLAPelRKzpqEsxwQmYpfWcm62XSZrrbwxO
Azg+Z0Pg8XfMuzEftDkXs11+l0giVMK0EfdiiVVy7dPCk6t/hMzwyD8wvyuQJbyW
Rzc5hlZYzfVT8Pq2wz1QEwCnrm2XfOdIJsQWpDXcrBCxcTte0szn4oxNpIlIgn89
5LqE2NwaUEx0KeDLDteVEB8RrVJo1rsWkm2noxHw9aAowxc2E0hL9khTvsopPZq7
IbJ7vGcyPNU1OgdT0egtmhISkF37TyklK7z9k7N92vtpyBU2tWnn22NMjmm8Nioa
oxhokI+Lf+kG1vgxpAH7TdHTSWb0XlpLpJHChF7XFciWCiPUoeu3EGPHvCy74sOO
Tlxo3zzyHYhmo71EwYOAzIoF+w+B0yuAU/h3pJWrVc4cJ5abcNhyCfmSZQGgxTEq
pJXVYaq9ZvdtGczjXpkW+BarZhdpzhn+JgCKBHJgTmFqoGZfXiVw3MBeu5kyLGtQ
2l8BCdp3O2j+T57ZwrwPkQC7TTLD2JrK7pp/IcCMd4l/S7BU8OhVmuJjsdB8M6f8
Q2HeukGTmqoSY44YkwKKIEd2Fg0mwmn51NN2jffGvQ7tX7Wv5rApfqYE0wsXsCjR
ZBF2bCnIno7fa9CIJFmmxcr6mwbXqGD/njT8uQI9jGmj2O4I4tNegzM68KUa2Vyq
H2LfOJew0Xx756q4JI+WVSg0yBrIM7uQ2Xt1lZ+QS2WnpcM6wjuzWWUY+vK6WUix
+QmYE3JZoQLoRqEljvXsja+OGbP3HGtOpYwunHGi9okRpM956OF/M5zuZuPqFsGP
uB/xLoVVcH3JpthqTh0jdWS1PhAI2Sm3zCTmz1+OiS976beQehND9P2bjPU4ijGb
NVwpbHj15nIPU4WXPjOtH6jLPaX8TSA52PGWcVHkInLIaXe/tzYz69zPQbte2M9g
R03Wum7ol3gYnwlGCC/eJJ7Ai30GH81qLTzlTMDTZOSebLjk13r3yGkV6A497EAL
hxrBorFIrX0pf7XrOqHWdbq9v46CkvGSfa81hhqUOsGTSUL13WdDJq9ApCiWRVrQ
OzR+92O/Zc8XguK+3E0A4DPzagAmQ04FrlWUEQxLc4Nv8NLmxRnQHbnm6mneXmC5
U4ugcAb/dg9vB2KOnBdbcgkTubzyukpOLV055UsjjUJ51ZR+/hyFy/NGed1jpPSj
0ToZvwjXnjSgTTclzcPEpO9HUhujhC+D8HftejrjbSX+xa9dirMg4XJYSHGw5G3Q
gD2fz9wpiizbsdbMPiShFzCwDqZFBO8ceZppkXH6Iap7Q+oxvftV4q26ec+ZODWF
0lXehoGntAkr78zvE9gtsemMhaLE911G2LHR3wwKWcZ3wS6kkA5P0jjBqV5lki4l
SzEoF9NCznU5GY1Atd33v464oaiXEKsPi+WPy1sqpFvTV2OIfJ1G1bRv0w2oWY9S
iHjdhy7PS7A+6hs07/sHqCwqL7soALZ3b6FZpzqPl+sjEfqf8T6MyoCRIsJ/yyKC
F/R2axX6XRX3LPEI1S6eSyH6Rbq5DfBRfVOw90dINWz8r39u4W81S6Ryo2Lc8fKm
fyJhhsr70n6SDpd7bCppKabsTACZH6bZ4eNlZ3lOfMsw95tpwEtYUgsyZjkTRkS0
zmhyPblwDeNV3w15stV23b7KjXFvkEVaPBMbdOyzxeS61vATr+zIJayeIRMoUOMv
0878yo866OS5nC3xc/JkTze4kC0jkM0RX9o89tueoWKOArqW57NyX7MFf2Z/Zzu/
op0Y60zmdXIoTdkxbJmCL522DfvNa6KovW1fTzF1jArAIf/tUIccu73yZlKRCctf
++ba1JYsCoNophqqJNDtYSNcXpmPEwI1xvMTdIKcdS7nSZtCO6WsNetQl1jyTmnC
0h7hs5NlrzlzvGgl6mIDPt1/IUxixYkgcMa1tJMK1I0Dn+0g1PRQQ2T6mQ6tJofQ
TXXAXXD5u3l6e5bFX6c/yzAbWlDmFbRIehmRqS5+rHuf5Se7ZEitqmdakEph5Pja
cybXpz9aBC79NK6rncH+UjphzHKXA7noh5CMM4zcjoyasgwbslnjv8nE9+8GJz/A
ADkqa5fk8BrNqB0VpJALAaws0UbmgQq2gjhYh0jaj46aLkAtVGz/75sdG+iGwZ17
JZ5EnL5+pRF0c+jNn206bAyPJMDIzQcxdupdJy557aEI0W+ULIo54vdkkbYWQeks
7hFey2ln4iOWUsnwXSo2D78YWj3W0IT2gH5M9L1gACP5sdelSZ1c43qOSdwY/g1o
PW04IzNhpmjiZ8omVAElra9gvgxCJt7MVABbHTUS9lOkFOtpPfLHkBXdpqQay+35
4vtVMU25AjRXHC/uNW3ShQ6Ab7oxkPay5wCBbk2h/BlronpKTy3f7f/13v3tIcIN
6MRojMxIjYADuDm730Ejo7Y9aCoD2UyeHY3hmxAtu1Xt8Imv1hY/+flEjolgy7ME
StUQtsnZSjpU3NxkDo/NEYsOn+UP1oNgtEPzTxKCbvmzkxCQ2uczt7+m2qljqw44
OFnK9qQbtxxxCZNic1b28cKsadEayvr+D1InnXh+Du738r1qDGYDZ5XRnuP9xkZy
8hSzraXCqv0XtfAEqB782HOSNjofa8fCLZzZShe8X2znfoS4Igkae64dfhjaeVO/
tBLqf3otHudyghIQvtOlrMd9tfqVcJQZpjUAwJ4MEKGnBi7L9JQ3BYd0Z2mzDk3v
hlOlAOen3UdtNqxsCI3gV9sP8+PVZoi1hcG0hiE+0qcn8cg7JVeubWXEhB6knuvO
Flw20HPsoSx1/BHUKYgGcvL+WwoQ82MZF4VtxdkGBDMIsI5nVr9as2748SMPhAfI
EuXABrhTdsdQHfqoVyhdifkzRMUDRFyoLbCOEJV6Y6mEWB9pyzU+6KrQ+RQ0Pv2w
IQn3kP5RKqHJyufM/nCwLJ6EiZJ9jNwzNcpA0+MsbWpx4U3P0GOZPp/BWaFRXA3r
jlAnXUh7rpTMNflVR5dWJOCCJ2Dp6wgg361oo2WE2MYV/MCiVgVhQOObmOcQG/Sf
bw4frn00pH9/YLOfKBiOOkEA3sactPgCtisrDlDWMfdPRIM2d5V2uBDRYBVNFsBr
rgnw3mxR6D7aOWxWJCxfMrSH7po7q/UYmvcfu63ESlBl8B9bedDf8Mu+MJ+o1+Lp
3Gnnqz8bZ3eyRfN60S4kzjEhepE3aJuIhm5qlWZAPlPQvCGB2G9lN6Ct0bo37bUf
zuHWCmEL7H/KnOoKqCDALLdwLeokywMQCxlE+c7V2r7zaGDt8gVSKL9/Nk5L9/lv
fPu9KnpwZBh/noNVasZb1gF8ZmApNSGrvh7ZwFpMK9qtkTGKlvhRVoMVa15a+Snb
7DztTxlumDVXIg1wEyIyLYqoZAGO5vz80svK/ByQSojUO2v+VmMV0sXReAqNKxM+
v9JXe5/4AZ5zglvyz7Vaz+E4meEYEiwmgsWCbB/mTNVRsDnC6ViIz1o8kfN+7tnJ
wjuFXcaECKOQjCxA/S+PpXePL6HuNoCGMjmJCMekQw964Gw5rErLYHRGHRMHmg7m
fMZdVWUoF0FIP6/7/KZIgYOdOpOX9dpiMArVasAASYCYepCtZ6IgX+/sOUFHVAca
lPN1H0KW5s0Jc/gMKu5i708VrFhrOBi8UhnbA3v7euHPAE4E7vwpjHGCTL+xSOMV
w+6ZnvbFntPpJxRKIXTRw9h1t8G5OmfyrKqMLXF/GFOdtcjGNUoCrrDOHAVcAIiU
vsPfs6C3lCTRIppq13EN0FgRDgW/Z8vg7AgbY+OHcE5fROD6oJmcOSCynnNyQtUD
k/EhT9+XFgBFkKfEwh3RGcntirVdiBZ5tM2ptgM6A6Ho17h7FcRKtGTpQG9vuC/N
assud/4zFKskZXkby5ys5cWjs1zXmK5jvOqaMWQ1/iZ4masI9wLjpAEyOLsyhOEp
oBT6ytIcDXkqnG1WmNJzrVJ1onbRhQVangT3Qs8XNI5F5ah7xUsz2SCxE6islbtM
Tb2POfkPsh7tZ0b59bQgCOB5gMl3wbKmVW+3CnjmNzJVn6HFJwwi2ZfLKWyED/nt
ti2bTTSF12oSRix86IzeKmBMH4fHBXw/YU4hRR4HLNaOUzjRBmvCsAx2ZAzt9xfY
uAdQ6PRjUumQwaLskMGUleumrJ+/nH4YlkzoCEHoaFlOxNG+qmq/q+5A19zNDBwS
AFvuo3xhfP6ZzVWwPstwNN6ZgaN19kNtVAOZHq7+1m4HBL1UQnU7knOmK2fWG1Xw
1feHDJY4AxZUnA0Y1xMeUunThrrErjDoj28J3n0fPHUpr2HKPVH7B51K13Ey4jHp
ZpRCGSvFbUHyQg8ItuWuQ4PSpkwRk+8U/zIZhc5EwmjEAESaBvrqdL+L+g8m+U4H
qq5yMd0hjWWyBIWfuarqHVPw9c+WTWbTAPMUeItHnfZShjNIeV2JkM5AVArJrwKi
BUjTheGO59GPvzlO4BFSa3E4tqtDsAxbIWqRJpyB7lF0DEJI27aTpMMoKKxiMb4X
Aj16A9qqEoCdApvx2LcjA7McmMq7D20NH/oLdc7LASfEhQGxZP7NUW0m9T5row3L
iThsOJA+wtofbU5SBxFfQoXXAB/5v/XgNN8cEgL85WxWZG+uO3nZlHjr10V/dZfs
IrbqF4ec4L1FixrHhHhYccAVq87qtUAoy3FRMxxLV+PrQU+Ou247gnkZ5d1hu5sX
aJ/jlku67yclGw7aYmAu5lrDL8qdzxgRuv1qsKgHGfv5fRW8z/TvxbeoNxltDwh2
xqokBehckc6zL/yirCbxomAskuMVbnGpHc520hKAm7+AZXSonRJ35Z+wcaeBUtYU
Sj4vSXYz/sIXmArp0XPsxPL5GLFafi8kubg9ItXkmIgmwiqaI+BG/10zUaax4uNp
B3wASFMnNJF+HMcCpbIUDm0IePnuttsKw7lCFuxwerQKJ6N4VhR+bH8h9/blll7a
vEwV6YK7FA/VPQigVYmF43rJcMUspaq+YH7dqa/bVdUE1tf4pFKiKNqUf2/bLcKp
EnbFhiWlXVeLG5V4SsNJCXxLuzTGO8+bOvVOX331FKf3mXUKTlFLIfUEGCGLOh/C
Ye+eESevxMl/wM8udHQ9yqYjj+QzAP4NERtEfAAfYSUsb52Ggg7BaR6HlPe23Hqx
X9B5p7zESZ87N3TwB3rpq5cL3/TwwvDhLd8yB0s1+Y17G8ItY0jI2bg9MIZ1SZpW
AxhJqA/Vv7M2aFD7VEBrPov46qAVg4dphdcfUezyK0YGAuiJY0+V9ag8MN8o13F2
3KiDvPrya6iiAfR+9abrLh2/FfLiMIGqVJg5QgSgKI/acEAQd3GXAc7cQNBqe5Os
rrr+9QlsUUwzaW/R+Ngm+3RvKffifSLCvxr/OfxSWm80erF+vMm1tV9S6Sgogpda
u+ljCBlYWaiN6cxWeuAuXEr3lkkWTfpSBn6yhxrG/vzjpCxkI13qlUqTsDKyjRHJ
jkNCV0+1ZUu1nhWwYuHaZFLWITEcggk8uznTeceobwScDclcUZ3+V8ckM9Jufm9d
qEy1w4IE/92rkvRiw8GnKtR200ZL8i2jQ3JLBZkq0XQx+JtbNGv0GDhBeUgGYsbW
KgXirIx5K2abEH/rq8wca/IZoeKRWmDs/ZG8asgUfHe1dqe0G82FM9Sz27HN9Djj
2sxW09rVuxMK+Bnv8gpGY2wsSSi/GuhIA/D/NX0+s36nMbsVcnLUBe+kYiOJTMHN
+v7ATvLVnOxcK49btlmL1eFFwtGmnKJkNMSqMdrKFt+xj7A6wVkPDkMKuiJqifZp
yfpVMtvy5FZa+WAr210T7oqVJo5/aVWpL7Dr3AIdWSYPlOd5eYzYqj6R2thZfm0O
zgSPAFLbSyPm7qupwWpkA/VAwor5NKXD/ttvaIX6BYJ4G2x+akWGtsg3oFWrP36M
7bs7NabQXC2qXwVPx8kOcx21lgERGN1Sia2+GDh7A4M7CjGqFZB9phh1sVoG3ggm
N6glZi2HICdbNuiQRgsMQbJo/Uhha0LDcwclVWpXNRu0Q56Uq4J9oVt1tNeaKjJi
f1kp6rphUjKT/bmrJqfdiIhtkrQbi3G3zl9iv9fCMRFDrbb3h5/JxSdlI2iQb7+d
zTa94qCDfOX6ET4mBDswY+jzOAWkbLOrUfUgc2+wT6bxwx5iS2qBkjr3dGIeLCal
4HlPhXygl6W++2fCYRaS7Mq6AB+TafFdSGDqDPTfFNDwz/Wm3lhxYl/xwyb3gMva
mt4juhmhJBxwOQiN8X58fFDs/RVUD3dWaJaoJD9VjPIgqZdXuHAygs0B5IuiA14V
WkHCaGg0Ai5dUbPXWy2Ktzk9EU8Qh6X2hCs7o4OY1Iy8azIswac5S3PDBxOYwZqJ
e4M8OprdZcBShn1AqIz4VD4ClJuYBqSQW8Eo2suOYdpHEYpmHWFtX5JhpHhALFLn
BVTxBY2mNyszqZVLV3qu+HtxYfDE5hGbg+G5XRzspaIyEseUT8JvkJu5iMeV1WgE
24itLHVNa3NSG5RNLJFOCML22I8iGimmTZIImR72yIKk+bOFeVu12jed8fKus8L/
2oMEP+CCu+k99oq+vlCnxLVq1Kky0uHB5TyFVAnxCzfQtvyUvQW2s8xqVxDuiNp0
U8+Bl4VEmOwEZjK2UQsoSqRTmGj4aFxvXVteoqLvF/Awx9Lt3QxDjjkmvYboF0FV
ViEt4RRDMRjQEQb0+RlEV+HVoV0/tL77D+fy7GZn73OdTTp0Pfji/IHIdCXZq0gn
ABd1mABcpHT4CUmjMbs8858QI+P0rnGYlM8tuKiG/iHNHtDa9AM3kuI/iAN/fPKU
Ms248eY4HFZa5+ZSdlkYcvQG+ehUXoraD4Y8lPbShBNTLVlrk1ikMITyTfEOVDqX
2iwafUwVg9o0pAv1hAZ69QKjbYSwIl8rlT97q5+lUigJIAyciFWvmdJsNBDdlGQf
ka46n6OdGQbEVuRMsT8n9dpabaPoiIf1VEeK8azoDoM/9xiyHvZpDbNoUcbLYWUY
DgMewUj3bPqzRVayG+kui4Z6Uda/tIdX+Q7pKZUHQwAZu0svdBcS8y+5vYpHdwh6
UPxc187B4t6qb73nuOZJh8Xu5DslGlQjjfRsSe2cA5IviNt1RdTEPwR2JCWhf9Bt
bajudxmAKATtxa5XzJJazNyjNji2h0gnIwft/keOKw72l0jHK8hDmy7ADGiIx7h8
8WAF3wiWj5xmGL5OiWx7wsEN3erTBAHHEFpsXRnvvcWmywT8N4H+dArawzJwwY+6
vaNjdA0GLQfzF9thCHf+i4NOyppkBdscHPcsGmbJMEQPdzKvoTVhskaisXmBkg1w
BMgpmc9Y7xPPXMpDE6mFefIoVq2ANJX8k3qFYvqqjDJF+ZeXbuNIU9ah/tzAnM0c
8hESRlQR8fClTfR90tYgIVC2BTm+NQWQiF8/mQhKd1KzmP4q3KnaoQhrVE424guk
1JeXODOdj4SRRsVmpopwDwsXmvZHgUvUvZFVscojnPEog+yeuX7bRX7C+Xaqv7JH
4D2xqvVa3+qx5jiTSpuGQJEC4eJK5dr/NeTEwK9RVBgqvMD1g6AR2TQ/kGcXGzMP
NTbXIlfsiR5GvZlYFcKH+/gSRQKC2xytykt3PIJoY6elAGvr/u3ODVx216ytqbNL
EvqQ2vP0h1nkJcIWWoEaiuXi9KoWQMo7ZYU57rwh1Vl+z1Vs4Zq1HxYb3XKTm3j7
wk+wTBRXyey8HdkgSByZvJuoWLwFtDsedRiq4BSBMULdkKhnJGijXqpUZheqAkyE
Sn3PsLxKMp+EfG2coPLBMdnVvD16CnTfV5oYwAfNEqmleHrs9KPEmXnp+msd3JYJ
74J/JnGPxzKJxhSez9LjBtjwt5SmOb70XsbcM0BKhRk0751VPnpqrXhi4VRwQ2s3
zangiYE/nCmy1dXathQEgORtpnfoLmxy05zgxO5K80CRo+awpMZ8s2nFWkZVDHlH
ml8yIZwqz/foVQiD5uskr2oXd8E1J1FeFlecu4K7IPCmWK/Itn6c2bM3G2JbkyIG
c3aNQc/LpVIpqTH1c9O1Jyr0APG78Qb0GymsJp2Jd8CxgeUCvpiSZ3htuvE9X2hu
fR4D/1wMhtS6TsTXDxTAk1xnmYUFUXOf3DJhWTI/89OejFRdfbvEw3TF+EG5bX4J
BYnUThDmUvUDNyYyMjPkC5G9e2gTO4pYEpn8e0Bn9KTDIDBb9JyZe3eHIXgcrv8V
zCdbcLYioGhCVrMvz9p5q4p/WQ1kKu5ASEeNE4Vtq+ilC1sPO29OKjNxzDMuJioq
l0by1VwIO3UNjZBQxmxuHbphhc/J1Qh4xLxZpAsvgsWlA8kThw8xYcU1lNOkaLJ8
VqrigofQTIZkZD4KL77pcdbuvjWmK0uMBDUjuv7vOYyV/X44y4tCZpidgvOusPub
zTYgyIo+CKE0j6DZ+fztwKtPlK3bLQDzWQ++KObty+z1MGdC6tvBrQLZVDyC+AO/
gg7w37M1ISPlr3mmEs4v7fZDfWmd3Rj4oXkCApY1ajhFtN67ddPO5W4br3NkjZ4j
eZuNdCHHvoDs0agpQnECN4u3NM0w+fPFsM4TmwM5A+v3R8J3xuEafXYnilGzIZEL
AvnKPlUWugGE/B6HuDDFBA6T2OgMvfCoF3GhnRBnR3g2yFdAWyQQH4x3BB8LMo3g
S6cpUiOADlDydBwO7sZwIRu6LdWQOVlZpiGREvCXjOdG3ZfBCdgUHPRuD1vnHtrt
3RTQ1dmFKDiKT5TbP+bpyUgeAwRGSiuFpsL1C1sJZqQ32Wbb/P0WRjg6CXeunv1a
9KvGuT4beYt4pKosTnmu2j4vC6+fwjUm4KU5/+ApVEAmctob40ZVnORFqJDq/Khw
4+iFRuBkVJLIi/Zy/cDyfCl5n5/YZocbSodaxskRcdO5Zl8Cg3juZTy3jyNutPR+
pCL5kOaHFe6vxsT9Z3ea+QI5IIGL4b7491Qu5Pm1Nhmsd9cX/rRCdvEHQiU1UvbC
m7y+aoAmRybZMH8k22eYdfMDWU1I3tDdhYo2KlMWzlADYL/qVyimhDG8aDmX0qFG
tpZnC2ow0FGSzBkk1uPNFucNYs4gNFOjAUKHL/5vYACsYLw7MyciZt61Sbk6+IcD
F3WeL94o+3S7Zgcur8FHb/1ME18MrNWujyWjuyUyQcJYjVaft+D9+wTGZRgyNVTL
YNMcR3MA7xNruRSb+0RYQgf0bLmqZjFcJnBmJKgUjWhPK9hR13HEWsda1hgoTfGr
IcytoL+T7scuEV2ZFoRTP53tkfNSzfKREMNoCdevb1W7nvn4D3/HQGdP+QfXwCCO
iMJ8Mp1clruZblMm50Bc+mu9J7av7oEp0T6ZGWaqsH/yy7KGONKZDC6bnYR/C6yQ
r1Oy5zXPzYxkZw+X9JqBuEL3nrPvC6cTmHTzjYJq0jDHx1JP8hYyRHL/N9H+qTUc
54f7+pt9D6s9u63JDHm7wY7x6P/ZyfzZ6i728CDK4PUOc9SqFhMvcAijbeSsYQaQ
OYXjQqLzet0QXLW1vbg35da+U2fSHZh7WV5AUyqXoE/OFtbMTbh6MytbQSeyp/Yc
3G4f/ua5lac8VZ2KZEhwukdEX+lgp0frrKNtwLBEUNgz3K99AgBxjQyJteBIa0yT
eN9hARk0LKKmCblWvI9eWCqPqAakLlpPXLERkKhF0bDw93D3LZoAj+HsdRUNPMat
3L1oLL1btzp4h1nm6N2smbJOPTeLudeGuShbjjDIt1g5s1lhSjvZiKJ/hWL+8dC4
1nydblwoxtV7maM9J5nrzNZBnAPKoLh8uXv7KXCR87RfHCaVDA5Lzr4TvFV7A7X9
stxHA6fWwOG+XoS6joTK/ZP+9ZhKucr76T805mGmA0JxGkXrqrKoaZt7PZ74hg+v
lyuAbEN/k9JceJ+P0FgAijsR6Uoa8HngXk3B/b498+JmKqDNBwwy5F+GMVh82zLX
rI5lqQ/VYxfnlt7CXiS7Nzm7otMN3GmnqxxXfhMNVBrW4AcdXKkvlP9wrUtBesqO
DY1k9YlKSJZ9RaClh7weFnmR4Xjox8KO10WRMKtQywQ2fwvTCncYQnrTENVgt8Nr
rBliuHcdYdgDPVdzglizPRE89RfF7tTM5qAa2eESI+1ISMKwN5KLujI9UDxTXsSl
JWkkDZKNyFB+XOea6JTPGRsqAOKUPOHmHDwvVtlvsx6b8qUQzh/9I86h0ml/VS17
hCAZK7FqT21Rls7f2V/b1drEMGzU/AhOJci/NMVFB2iHXZyV1dJVLdlQ8BdrOGKw
o/rl1NjjN7fW57c0I9QHcaHCrWcj71SYwLQi8rizCJUSd9U03xw02qvrQYBpqH4Q
bteptNEqGxv+OW02dbHarwv+UTMp3DqSP2XIL5EE9g21i9d9k5snKNObUtMdPMQ1
ElublBMSbJ5bIYhsdcnESFoXqCGS0d6AjwMZJSILHDyQq7ebLWsyObAplh2e4G2z
toTLzAdLfM//7h7HgFq9PCw5Zi8nXhkHZhgbautNlFqT7b+Ngx2VpTp2nXZZfcOs
qSKxhA6DANPs2qmpyn6FNWoGme9gCUfoBLjKrtESMV7k6cIxwNxwe0bnkIurR65+
gP4I5Cwcs4LTDJnkrakdWIzOe6yYQ2+iUb2VFyfX5C9NBuVhWe2hLj9Dkech+xZK
iVM2ULZN8igiUNxUt+lRVvXxvpEF1S1Ji/LZ6BxKBleRCkTRuo7DKSRO0YP1t0Z/
BtHhd59nO/7QY60RwdMlVjxDRShwx4kp/C4jDT6LoQLGHLAvafY1FKofrxra77dX
bqPPsrhLt0e0K34nW7yUsuuC0DzENWzBxOLxPX9JuXerS1RQspeMS+3fLZisQrGa
Wh4zMkz+0xGBN1fCehr1EZi0RuZ4gRmbz/3LTub5UXdcac0snzAFLgm4xV9cDElW
rShM8BKwQJ961blNWXIeNgakvsnFrtD1DkpfxPHLcEIsl+deIPGrPV2EtEbQlrUT
p7x1nZUeKylNGq2uggFjIm3LL/tfYRI2hiZCec3VKL4S5+X4glKBDtkWm5qJP9oU
rG7ou7qKsJ+hvEIJHwP6dZp0e+Tyn15DN/BF+t+8O+ExxUag4SmRDrAq7UC+xzqT
JqqzKT4/SkfpNx50T+M+wt1uAT60c6E/2LRVNYYIRnv8243x/kg2jMR7tW95tKYM
DS/4BSoudbBEO3Rr3zRBEKmG2DVv5cseUJ2mb7QvxJ8G/q/sjjkR0K0LCgH7t4+H
f5ipzjuVtHKZixyYtw8SPyQqPWnfn8shgNO/LOcGH20QnF/bjMRe6GUuljocWwI2
X3Sezq6UfWg07b92MPb0rum1YHDXC9dLo6JumEX3/mQlxwQo3QHw/BYOgqcVQY0O
cotiXKAbGxCsXD8fLjmqqmPn3q2UcmoeTgJLm/2mQzjogjqVWQurZnE7Qc+9JMPf
LZzE7tAUz/8n8MMAtvtQ/IH6MRT3sG8ealveLMuOUDwhlOFDwaSCGAwnrFMm9BtO
tjdkT6qvmJnngl2kzXS4JzoyoXRsEBUUbhHXb7H+HTenIWxYED14DmKw25XhmfjB
LmLbrqsRElJFo6QJmSog4ahgNRziy+WlgN2J1yT7YWyIAh3bA0P1SCVyUPgn27ZJ
6m8wcG2m42+w3+JqeIzG6lv3bBhMhGZ35n1AihUFZ2sVEj6tt0+u2GoKlPgZ8KmK
/XENIh5C0kWAdOHZmK/r4UvFnXqcACFA0ut5A+Y1A+88xj4k+zoEPRSkKSiNkhZ+
GXyUYVycFHM4RTlqjPAtM/rkvstshrKHxbMJvjgNX/bCSIaFJ8UEo1K7aYR6gI3g
R6pEQHP7Quxf8Sm8vqc/iHGhtBXAtsRTGWmKVf9OoMzWTPTqz+wOsnGl2ItDRjKI
T+0nugUibjW6RDKUg/k/uepVOQkjWKBe6JWDu5ni9qWauX98xUVO8NB1Vedqy8lG
5S8ADK3JZ+KdUDYdn4EVHlZgGaoqG383ehQTbAg7IUHP+ASdjlXaG5zqfBT0mHIE
Ypz25lb7oyWzFXp9aojEXwfBh+rLzofFfTyr7vWoOTH+ThkGV/A1Qpeu8eT2AW1G
M8GL+OIr5kL6lW+Tayf3FqCPXmvyhrGgg/CDTcWxUn+MRKVvHvUgOG+kXz8bqysn
oUeXffP/Q8Kgsdxw4x1RDthVMdXi00wN1VO6hoPkoWvrMgN1pf67TipPbnDDqfLn
s2ISYUEx1mDVCQBWwzDHtfrUoSfFK8Dqg+QK0AhpdYgDsQxCuluOcf2lmIwEoMEj
YdTznH3yuBmd6Cd7rKpSl3yJXgOrhfyUsKGGAxx6jm/BgyuvNBKuL1J4vhUVDH9d
ewpT53/d3O9T3x32n+XGnfCl2DlCoPEdBuUgtU5X2X7t+fU6IgKIXuwnZbNhVAsX
qd7cWVKO2bdH7LmXLLF0iJtEDfucw2DCdqQe0E9nk+CE4+VgnhufHZIiR5cbesA8
5d1TfnR0d5JJjmxwKuBIzFSbCLaP0RxFen1+EGEUsgDd7xLgo0A2lfXo9yqY/SRL
OH2dqqggfwnBepGrqhKmy/AtF0UMfwPTEX2UdWWl8ttTdNaD0OQt43kp5+9xpJLs
xP19RLYP7RP7jcQZowz9LVKEm7lw+rKacHnIV7ktQl9Rx9qp8Mju467bAG+XLTnO
9hEyYdrMUiA0fOgquva7KKJz/OXllXw68hwPT1cD5A3X1F7kGJ44zfSYw4Qx3wKW
jUmxVu+LS1Ws4I+bb8/XuqBt+RKJZ2hyrcNbj5/NtlJqlqZsPsbh+OK8ktK+RVrJ
fxCyQcthFStheseKpwgbOLbnHm2Nxf6IlSCQP0hUSYY4yR9EDusdFEoXhPOXdhFB
F+L/aW52HsHHogjJbiPrCEJ3wiiCC4qbj70BTZRVgTzE+71hi/6J/vwGxfLGDdeU
lacx0hxxV+jwIAXn6pZwOxZSIdgye+CaIndPpf6+BXlKoroLZyE2o90u8BoWyi30
oR8K6mE+eCwzlHCAgVQQ0QMm+J7667VuoVYntON8rsWrhAIeDfa9PnSafZf+Zj7K
Epm/ZNK9GzFrolVKlR044W8zuRzw5nXCqpXh7rrAyaOBNbhExKNM+KDMkGTO9PS8
MdDRLvG+g4VpuD06WlE+5QujdiwIeOLFvNnRYnxvnyjmCQgrzL7w4+aI/h78qkJ9
E/VzNim4wTFgGhv5dUtBAAw0oN48k7cphd/SQ5dAztbqIh2Vc/Nt7M3uQfSYTT02
cGdvPVDNtQnOGtnmEcVHwVWb2vpGd0gQSMQodIQH8VVSebwaVT+WmcCAzgyAFHNH
GWwj4S8vRbzkK2zc4WCHK/ZnZlFI62WtYyw0p/iUgR8jFlWrQxwHrHKS4nvj+EcW
aRcBtLhMd5pJaEbC/dvW06xCTf1JvXjHEV5Ovo2cJVw9dPYh2z7YEDaQssDqwyMl
bnUZWhD9L8xEKGQCNmN7u9aUITcABNBeG6eqNpZnQZ3VJGeqICr44oBeq/BUIvVu
9W9AOpBanBsx1YNwYevaZICRDJ4X+tIP3D3+Tz+N0v3pYb2LFHGBAutdRWNPWppy
oNNCnPFpge1ME3TRDHqg1ef9BKji33rr632mdwLAQkYCfOhgVy+plIsRhXALTs0E
3KXZnUDgvvYJfEv2eYE/5KkL1R+H+SXZXjeH0NOY0ELOMBp5cw//QYVuB4Nm9Ew2
HPTGeYLo7HhQ6XVjGMA74lqYbiaHyd6qvEVKs+i0BF3TBuNq6QvXZkYZ1fnBVgbN
cjQkyofFqr0+YXugMrIiYQa7RpPwwGiSJWIdbVflDkY+DwQQUMl1HBVt7d19Z7VN
d1Px9EIsIYJV0DLLgeUvob1Pz74V6Fv6AlC60VfTIrIXg/Woh86mEGuB8da5/iGQ
X83UJKSCI4S/Xa0dsFYNhjOXM2vs6yqvQ3MHGEJgSrIsY0VlW4I/a9bbmTxlbB4H
03Xd1s2fdDoIsZR6F2Wkwyz1uEwlGfyhX4KpaHD6A/ZPVCR2wTrEM0LysJmQV/eB
I6wGLJBmLZ44dJ8aX0XBqXnsxNsr9EtmCStfAMzSYZPSqs8o2+qQ8clA9KX540jT
CeGiogDrMa5GIG6PKkIJ1UjCaKUX1R0YetrJWZJ23AsyUACjrhgmNr9LcYsuUWiK
8F+Txr9fKCbrVe04K8rIGhFV/jmjPaX9G3SWEb7+kWzyzpeyFhhMZ7GJHf6LCqoy
dCrxx0b5c6/sgF/ngXiPrxmFsavs0jpk/tsWR+vS6VwJ6zy1gNBuEigfYvygrBrp
6hWJrFXzD/FE2Z7+3SvjePOaii+zPT9x/+vlW7T1ivmM74rDKR2FlDMUFodRd+Dc
STcgJXy72x5CbU6ukSSt0PlX20pS9arJe5cRcbQyWqm0Nxe+TXJ0s/9zMMf/v0pi
A+49Wla7QaUvlIFGQNuY4HQJnyi7/sHkxhOwhjo4tDvl01izaKNxRX4akDor9HsX
nsrUu+0R7qZQYGZmQhb/AeHvPqmYN+iomCiOCsNHSbdu5CR0ShM5MSB6AhPWxW6I
n3RaKQOtYCpzww6/1wpGPnzoRy/P7JhNJr5AutkeTdKtA0sKyz32YjRjftqVkdiD
6fbtI3AtPgv9qMM+QIpoAcfGYPOpjJPiqyPZE6LOHOWUzTb+4HVly6lMnpJvwaTM
nFJbXeP7dcwHF1oU88BXaP271WMOL7W2lBMJ9RWZeZ7PaBtoBBbagXfpZJ91cq9Y
QCuP5tdWokRZqFrBW8YfuZl69vM+QMsNR4Tqu3JPTpltKmM+rnjBInQyV1KjBMMg
kPJt9w+Dm1HQy+39pCzYubCpr3LJgqnIq0WkSksPvOG9OGo5ltYX51GPVuB038Ur
4H0HxWK+BNp9Wfz7F6sIAVWa2T7T4FMqkoNI6Yihn2nBd+Cdic89r8fEl0Ys4FZv
L2+JphMZVWblOW99VS4Y0p/X6kkWeB12eWB3bovnp4uL/IZrZ8Z9a0dJhlnvnMUf
e4Cx42CvLhbIskhr9kXePBq6SCmt1nlnw1ripS3VgPsnNnpxyXu3hNW2iYWsavMV
/4BYCJBdq+DGk1/gVWtoUF0b+k9C5JG1b6qtEcSJnow+2WhXd1DEIMWyqqxsAq6p
pY1Na68Y7IDgqoUHBJIgf20ZsagwJ2C4h7JTQz3tFeeKc/tub8RdI4ALxu3LbIeB
fTZ4hz0TRi4uQn9WmsielAz8G6KHhHnVET2dvRbF/4QAQef5KhmzXyoGxxyafgks
QK/9u4UM4Y7WZGeeF1+D45/0BFOzZXFR2uZjuGQa/kQzbl4E8xZg+FyU83xqSPtA
gZgIE/lV6yJZiYjhMlNKyTbAG6hx2VobvEzZ//L0krlUK3N1gPRrdqG1xmLYdwIe
czgkgihwY9aC0am/MSFItH3M5sgyt490Jg5Ukpb9vy92AqLch4XWgNJLtUsjAXoB
M9iYc1/L0gLGlmzu5ugDWFW462szIfoeXR66E/8n9T9lJ4W+bEHLz6KmRJ5q7Zwl
keCzTmJh1FAl6nnT6OrKsM75Sk158N8kEaw2FIeX2pUIMt/tRPcrEANPqu4C9847
YhytwTl6lw9kEqrGLHwXQV3n83MHv2KebzsOKN22ZxBthdFtgqO2/tl3HcDKYBQo
wAbZRmLWP7LXb4RKPZLAWUw0OBYelpdDm8o4D35+zekyJsraRWgqtRNPiig2B4H1
fcoAewD9DUhQpQps67IuavKoQC0NM5Rm5A2mlb4a8riOvLEtkQb3fuIzFt3yHkKX
RdCV4CwwRIUe8jmbtHlcG6k/x45Na941FbEE1BsgCbF8j2y8PVu92hasVlsyPxJk
7X3ULmNgLcNbt41LxfuG+QrvPI0EV/PC3IaZzg02UdyigepaV5+DVACtsaRE224E
toXwIoCA6gBInvdwSG9R67fPc2hIge1r2Hct7vydO/yusUxT708ES7G9btxt0A0R
7ZglJZlv7gxE1g4k8stPOhwdoiz8IjaziYsys9o6ZoKFeX9M6QkYRK/2latGalD1
0RC9m7GKQarIisWZb2vX7Grn44qNDXbryaUUIW8mpeT8zKrj2HFfeN0VjrAO1CEZ
D1llcOSYXAq2sEpnIxDTMEk69HLH1SDnwTX4u3J/g2+zwFR0taAoiQGNghH37cdI
ZllAkRj9N8I20TpK3bwxyt+L7LI4zq9qRAFtQ2m6NDb0dhaxUBEmAiNit38dOH8a
2vBzLiCTd2/CvFP51iOixrAad8rJ9hThrMqF3Q4YNjvRkJ0nsZWWkFBjnyKuREao
mvVxPgtT0TcyMFxQJ78JgtJjH0wGCB2QKoXeO04vUlt8ZXBjpGFiri6R6bfGp4sq
IJKqbfmlEnyORT/HyI33dDnj5Pfd9H0V/1tcE0pqgcw9Loq5EuBx8eQMQYAtwtRN
DyVsrLNRrZ5xJofirRbrI0R9D5nljQZZLCJikSeDUxgkkjzOuE92RVq9G3ueC6ko
2Rb/cG9zi3DK/KBraSoqFN3rIypq2A5Eshmac1WD+uajC4vHEN7DQmvFLCu5BFs+
LIUA5G9YO+FGwGxuZeyTSx4+aJieJdk0O48AdXzHajelR846Lszt7kqE8eG0/XYP
1TWXTdzWvaKPXWeXS9SUp8r2bO7+28gYRuUFKkFfaVkMn/RFn7PREX4CGzw8DI6C
vYsh2iK6wKirHwSJsTyECMF9znjXx/i/P88HvGpd6XBCmgbnMuCR27lSHeDbOFtL
J9MUb6LTY8yl0QtC4Gtqt/kCM/ophePqWn8vVrsrBxw5b/VZaX7CFHh4LQDEjKrS
rzTJWAiPM5otyMrf0iA9Qq5JZz1iGKFiNSBjVSldAhqkTGF5O0D9cRkLz3nBfRud
P0UdrO3ZmcBXFzJ3LPwP+oKv2MaEm6dbeYC51UqPojl29Yj7lnU+cqMKAMSxhSI+
vH8e5wEs6iT508e8hkFDC49digtnLpARu6ne4JexHAhCRiv1Ykz81+9l4GTm0BbU
JXKIFD8QUh+ER9XD3XQE+ATs3UeNpWMh/78hh7zRvBQv/3qIpmPk2fiNpgVfFoNr
hFJxYYrEfw4Kg8AZQWaUmb7wSC9OGmoGfu+wzEeEDu7WCtWj0sfbzxGx/pcv/aya
O2tTmKwlUYZ0uWcJiXu3nAC6u1I/nhtEwca8vvCfLu1uCXpQR/3SzQWJWEknxOn9
L9LwgEZFDl8rJ0pFTkUt54h7fVLmjRcSAEApMLpSsBIei/N9W+bHNqWIMnwd2F7t
LRMkJ9mGiFIRf2oktNvIi5tFRou1E5lrGz+prW2xd1WpzumVhers9Z/iXpmizTIa
Ufw9XnKLFba1bS8P6LDKYp81FZWM+4lgjWRRxy9N3Ciy7Z/zeEPQs3lzNMGkN3fh
ANU2XFvqb41Nrjo4RIBpRT6u/mKeYZXsP775DE6MqUxeN1gbpUL+bGE7yRXt+SS+
cA1arW6HTHGQzP8fImdPSy/bKjA+OW60Ryv5RJwwJccP4bCMJnYqCldHdI8qPpDJ
6epFSUMJ1j03s96F83YsE1zg9E6+B60NyjWDrtsBXz+bW948RYTqeCq8D4UoSz/Y
gSo0gumTxwyEuAJZlshIWFGMgAlLD5ealEs2V4I/ToTaqLOWxL5mflJf+CQX1pb6
82Zj3xgx84RCx/2B/vw33UD+E4/fxH4E4+lux2ei/kEHatWjBakFPLw0L5YVeXNL
4GLHcpfd5Xz86KePHVLjXMz2qe60HWJz+YgF1nwYM6Pe+tvaUBGx0LdSWq67lyGI
pdpr/k1hn8YS863vAMr6NIiaUqofhfbTvKULLE7rNjo7Hdb1rlJ0qzT3Yt6ID65F
tpdoqeKz7c0hbwxqjO29p7LdPmRJ1MmNdrtmbU6qVFl9yNUlIyYoknrvLvcwNzPv
ZKdyHLPi5E1vIm1wutFJ0fZvLgT6pPsvnUBQKWfULC3jPxWEWmS63yAQR+FiWCAX
VpRCqlaBKazt43UcVJkhOIXOXDpoTLhsaBzAXApsrtIGyyWousTvJyYN+Ix7E9Zi
QAfECQ39E910KyNgIhlwP7+FJDNZ4jqTkVwDaZr1lKGb6+P4SnddAGSy3jwf8XXo
m1G8i3jsID0igNiT1BRlgz1cOgoqUd13tMCLC7tai0xUM4cHW7MFFa/TOEBYD8KG
HriWE8oh0uVwcuAJvCN1JyzdG34Gxkq7O2ieS6P/B15IWp5eNAUFnPC17Blrg1N1
b+5n9MfOpwM9bvbMRh1dUO+BMQ+E2YK9HmXhg7eY1vnOGKuxzWZBwJdvFhTvbeYO
PcBXmYEnGIA2KUqzcE/I2nkCzJfI/gMf3H3CiFXFPr/KIGoCDwAq1vl/v+zOKUWo
GNBgvnoDIScJZBTHMXVKpgcUv5sZC44Zd/J6uylWWDNU5m1R8KmXG63ADJlpi6XI
GhWcaB1Hu54QJVw063t9dBjLZKiuTGW89RQx8EV6jNMS39rBQHPR+0EbNhtLxNUF
ANpZpsmuNi+djaIJNyshHfuh+bkPZNyUb3J2V6yIUAUjIl7YWzoQvcneWV0oRSVf
kCjtBcvp+cG0mlnrli7Wd3SZfUW++eJpa+hJSWhH2c55OuM1JOSSnPCHdxj/Whra
i1Zb0AYm+GBrXxvD/C1jcZJz19PdPPNJGgExg4JcKmYYqClgM2n3d35eG/CaTFr4
0EeO0ceCr8MvJxptuXTfNODwJ/Z8PhzyU/XHMb1awPlP2+RGRnx4nl1WPodxLBMT
K51ErWGH1VGbDKHdPInnHzmIu+nATSftKnBSbXEIUdEsNtwR3/Vp+rdsKgYW7463
ghZxXvY6w+xBeWogf2km5xK9V+RutgRN6tglcdnql/NETxjD/0Ccl0KFXZPR7GM/
dyQctjkK7a7I323WIy0P8RrY2inlwuwfUsyBsuj8hm3sxuspqX3PS/kAXVQ4jqzC
0KkqmNG2nxF5DikoH7j58aeyeYKpqsHNtswk+2ySWAUZEA/G265aaJRKstqj7FU3
NxrWljaIwFhQ2d7aMipMWO7DXUqvX6A8GgSun2Glwt9yb4SZHdg2vBG5PtfQhWBA
6ENBVPG8XErRmeUP/u2L/B3w/MrmugGgbFW3BjqHv7C1FKzkQbyY/1oveQ8mxUwH
Zu5b65jtnkFcCmaC8AQlf/CAklNl7bkD36EZErXbfPANpKABNMoxC9rd2f2VRuA3
DN+7tWQ2kWOeFmx+pIZAwK6Mpova1SMtlcqdC6PmkilhiFJ8ovfwuU6ZttA0ilWH
4CIZE9VO0RRR8030W2p+L/STVZ7adweHbxApn9yOT9N+JZCOXOIEG96uVvQwx8Tr
0M85ahhnjG8Ze0HZlwG9AeCI1atmJtYqsT4H+SWL4LZb6krtmLBKhRsyi863aQlE
KVsWxH5AWYVgqHYTIrrrsoaUeYudfw9U9cla9m1OT9CMbGKLq6yRIvIXx2NNvf4F
ndQVmXKAzNmR7ViPaIf3qQwc4n4c6uTMiSg9UdVYFNkzuQ9YNThVk/jpiCnPmbAR
TraukYfUjmpLIISHT2ZkWkdbzfy+6FiRN8/2Cki38qYDDbQez9aYcc5vOYwZ0iPB
wENyHG1k3DTAWmRU7OJ2g3fJIVKG7lIuLWsosztCgozZD1Jq5KUC7muhuPonoNoO
6Zczz9hY5Ponn850d3U8hEdQJmcejMVAbwVs4NVQ+Y+Sy5TdSjeW20CLgJ1bU+bj
C4vVzPGRwdAu5/3af8cep29LOsQjtruYpj/LneCDnF/mLtMplh+MWjSLR8cfo7lP
OLYaqYIdjEwJrov0TWvkoBfeUoG3BfcJ5zLw6ludXvAudwypBNP1QU8FyINspJng
4zDucuCaiVkAMLw6g9rlWpGoW5KHSbMLhhItJ+vuI3BmhAC3I/pfk5FLM1GGXqUB
3IYXb3O2zVhJ3QDQ2NLptdThEU4MwsNB3tpcEFH8q4zl464lFWTvnD99qUP9HObO
4YZq8pmHsZQcSqnhhzBNF1USnYASeaWNPPNgDoPFHA6Kfq0l43Vln3LAaArwEE5I
WMvVnVVIa9M1zKpJxfLaOwL/R+F7SP/B5QOjbksZVCJa7QhevIjLc01zaXxZcxE5
Fda7/hi0FLANYu40CA/+x81kiFUKC4JQxBsbd8ySoaGPCILynIAdRdPmNnMqbO/S
fZQqQRQ6Fe3YxrSAu2fSU521AwSM+AnSHVXEixNDM5tTWcJjJq1d8Nsm9R5QHNYN
Urm54WYQWzwegD63PHEE6GUDfGoNturv+Vky6Idib9aBCLboHYb3gHFryhEJnHo1
Es17+eWOsnJ88j+EjS/kyN28C0iK1UhaIc9MOe1iTwXc51E2jea7QDhzb6vQOD4s
vn7T2dFVNDXZ9PLJNfFXAqZrZ1HbpDVGmBCKF0cSnuU3Y5A5jHW83PYWkNllKR3j
8rTUfv34hKFQPctVLUD6kPtnq/B6u+BM8oHevOdAWtZ9PytQx+HT8VMgTMNiriMF
asoTH2x4+VsK9ZU8mQ4S4dcGdK6L0tWkSEv+fA0Yxfcx6O+wybj4Dmd9V6E5sKLO
YF6d48PyNxN6U8Uk2SobIwagP4H7lS7PtkLpUQad3PeE2+I3jDkhcmJII6MicVob
ln8p1EKO6vl5RqclAVER7wer3W//FJNk37stiM/xzYF2Y2ZKFEFRlhIRbZimis1V
unY9UH3hPo0ZJHPG4EdqmV99bnZqXc/f2UpbxeqN5xzSVQJID8Hch2unqkN3aSVu
DxGFfpIIhyRUmvqwp8bA6GpZesvsGE0dUUyCicuvNlBZwaH9wP5Yqbt3uApLExI+
Q6E4CXtIErcPGP8hq5rii/GeLCaEuvP4SoyVmLKCEomfLvwlK0WnP31TB8qx/3wf
tYsQliTSSUw0iA3lSOThLkIOIDWDl1gRMi87Z4IgtF+mmo88EC2yWBDf2TKlB58S
D88wMWDTgWV4x+KaMYLxknxR/2IdXccVnFuhZKAAFX5/W62c9iFhg9dys5Dc/rwd
NvD2tFTNPqPwghIwQpzhlKeEmtu6XaDsPeGEr5zJEEO5bgJVbsVqG7oj3s5dLIcI
H1Avfre5uvK2nHHsMpNvos63D8ajbgBmwluKnBQ98WrGgM7CzwlaDLqx1FKeppsZ
B9+x8Epf3qqinazWfyAa14Ddyxt4YCvfGY311tRAfwln699Jsj6o2Bf6bmer8eCW
HjMLumaw3Ru6Xn3urg4nbMvTF3kCqKpAMx7AqCHVr29GfadSnU2vvsYTfmn4RmUq
tgzkbDkcrtZ3vVe30gJBcm7QVUNdXyrcB9FAfgppyJx4XV2TAwHVoUrtgFAtYH+T
nQIrUSgW9DYsLrY6N474pCnoeeAIJDuvKK+goeHnWTpSsrKLXRzgajK9WTZ/XqYi
LrCXzmGKCWQNPtIwDmofSMwCwKYIsRcbSjAUGt+urmDPwE6dmPPc3DpoXdV5kkhk
d+cpYoc2zcKi67T0drYG8ei4wXasAs3s2iNmP6W9upWIzO+hSoA1kr8+g2hNAxnp
OLz/0NWCiJ49Ez41Qh3wEhDnaoDw4fd9jmwp5lSAwt26ejfMtKYtiqCwebfIr8YC
tZSbFCh2BurUyGFu8oCKYUJJxJkeCVn+/QNQNRjdrIPSt58uVNkNrB1UXijnfQx+
knwVUvvHeaw9bGTmkc5dMBrD8pTck3Wmw3r8+ier5TXAMODcuyHTdHlBUHmr9oug
5CM2aqR/OvArkQXil9XPcw3eFynwmOs2SMPIotlS9zItMmiqouGPFVijNByiggz6
NPRZYN559yiw8krSJ2KcACAvKygFtL4jFFQDexu3bUAHRy6PQi9d4VL9gdX0Goir
OSlwgNCE9utMikbjtv4wWPZ+Iy/oBF1hdKqHUGsKSV5Idw8naubkTqNcGW6DYqzG
1jsR/YIz4xnsRK/D/n6LT1VK80vutDClBBYRDORnycQCkn1XAQ8JDPG+qErT407s
qS5SLn1L9RHKdm8WTTUDe9BrcPhtp6zWh+gMtsGCswskeJGw2r/pSLFx6M827sSA
6xnxXjrNU1UJvLNgKTslDkjCDNO/sk1+VKy32YqfLRUhqdSff/onOArdwQsziy2C
B9n/q1Fl1Vzqirl1Ex3pXh0aP1WZN+vV1xC1yFoHMw3vRcnzDO+340+bm1WLlDd3
MdD5f7Me3Owuw+iKwsh2QtYNBhRcCkpae1xKkqCPbjr1AuXCcVW0MWsUh+IoLUjF
lUMmgn/4TmI220Pbz+QyUy/KPHFQ0NEDh1zHbDw3wpaNfiYTbuyE4ZEke77VraEO
FlM673CQi8xVHM4EQrWjOessEzr0xDjq0ahLGPB/OYuMR2d0BYKaVDgMBZXiW+nk
O5EPxxDLKEXjF4JrkVxgrEp9+i2nsLr1lFc42Vd0SJ3cVuUE3MxtM0mvROWd+xHY
CwMiEAHtSGL5xHA102k/FpeIb4rE5QYwMlL2y0EAay7Q/81G/0gUIebewS3MfRPd
uvj1b2ne78cVNXjpH3pFkSP1BJ07anwKsLCs0gbYKDUJ2Gt0eyPaPcMFFIDV/5C7
o2DlrY27nCFeJvpWMcS6o70prZWZm95SoxEKhHTC3m1iNVu1Usj0P/l3bS+Skyy/
CydQh+yEFwzbOV4g4UCA2DtCxTra5TgXOPpG0yBEJ8m2HiSxic5gbm4pT9mIc5Ic
KMG5IdvCKn1n/4C+TOlDmSvRUyMLCNHBHm8Np06zaf6t4aScd2CfP3AcCNdPmObh
yoveDOcQx6qodZ5/UD+AbJGHDGciNSX9TtQbtpX2kTNHhTGoYr/nnoRJ7Hd5g1kZ
/MtjoAs6dJumD9z6lcwogkUB9FwJonQlVyMtQYIlFOWDdgwtF6L3MuTRy5ZCChR2
vqO63huIiHILP/gJKbTGQp0ZU0d3A8QdF8NhwEfF4WB6C+vkoG9KkVa5DLgRLWN/
ZxjTH+T5AIAM0ZIysqfMwJ5+sxs79f23qstp5B/RbKvytqnqWtT7RW72QI29vs5I
86uhx1BAKFGZGj0U9pRFwldnrizMYaPr7WCeuXAMXzhlIIU/XW3i/WAp8NaxayFo
GjRJi+OAjz2EHfXrREk82Mx73RC5Pia9ESlkT84EMjGk+M1VZa4MpE6q80tIZj3c
VPXwLbhXYDHMxHdgfYqzCKqc5IrPwntYg4GC9uOkrH/WQuDELTVkTpVMCouJLJvv
kWizwXhibNjCRPhLkjIog6XAqHwrSvnBdfeZWCqBMUadm/g0OX0EIoMkeEugy4k0
HQX0Pws/yqe4FaR9Si2rvKJdLzS5HFKsnYkQMCg56A5A4z4feevymuRCOIrWf7th
T1ZDYO84t7G1qIgxikxP7ZN7x2g7dPqaTqVETtsNuaTvd+QAs9hNvQkF0LjGKzie
AcM0X49HQ653xtXlNwPH4aCJd6MPFmXqxobPCGds2iyIQxzOjFevFj2YUz6xxHzL
ZHYeegvx1lihMcCzpe8kTV8bUvWHDJ1L3+Sk5xLSFJzOX4fo3gRnhQgiUf0Rjlms
oq4xvqzxCZm/EBL2rZ/HXb+aYVBLplQ+e6Q/jN/rEONY0bvwE1qx9JP+K4ME4xmh
TE6KcMBMgVx1dZj6W1Ni3Sx0abxyQWlb2TCVGUfQFDcr2NnnaR5UyJzUTGcXZpew
uG54M0oCwCsduTSdBAI9Yb1lzkTbXP3j8B9nfGgSOLOMNeuqRwyKDVl3/AtmNfSB
qikcJXOV6TOkT4ZibZxsYu4vzC9ph1wtaYhkvHdjJWnVX33SX9Rao/UrJvRln/E6
5KDtaYZuAhTs64uAJQPliCRxUMNy7FTxVHhaq+OFCgQV49R6O2hwdA7O3+qdza/f
VM2uVLS2aWMtSZk7SyXbi+/FJX89b+OpbD+BBm+VsO6E0de+wPzHDVsbYXSSU113
upAd/WCjWHhX3Ei82kKGKDmbDeWYVlQnRPHaCEAtATBfOUWSJ1hlM66xlENfr5xx
Vb0JyS+s7ghijZ5rmhMl7i+wzsTlpjVc8OHWJuW53/wotOoX1ya6G74PzRPRsOeH
Ac7RlYARUiMpxTgeKOUreyBrkX7sJgfKimjsFr2HUawCWRk8AlnrlmXsLraJnQ8F
LIFrTKPXcozJOLdYEFZc1HNbOOK8eLytv8Jp06uQgF4wT6Hg+VTQ3m0h7uwXI938
FZNRiFzkKCjP6ADjm7X/PlaSQfYWX21yuKlgs8c4Q7JzDUMKSPsOmiMaeNgTyzMa
TxMDNSKYmteFFgQUeMnlLNo/5IY65Ur8HcAWeW7o++R07mnG9luRK3dqdvoPfhU7
6tdQOc8j57uKHgUXZLfpXbx6FKNpo4R1KrhFjTwVt4wJIaNwvDBgxpSgxm8vytVf
JHqJnMAU+F9dMvE9ep+H5OGHbXzYRAgxgfrLp+4Ce5LYTgnkCd7jjtwOix9oIQj+
eY5bHhFaFNOq/l5m3O4Pfh6j+4ELU1qNUJh6vWQeM4I5Smljbm14GA9/rCw+d33Q
DASNIRGSvW8/S7VOmF7ZzxNJEd97f/+J5upSAYs5xC6sMyEDLHSgwDgO3dJdOadl
5RwMSXpTNRDzJtd5BKquLmo+DgIharrd8pD+sA1kiCx/KbykxWZwCbdpTQs+YGJF
/9lix6mKxYfuxoF3ieLu1jxr0j+xV8WOi/q1mPbIGw8Cch3eOjg9heMI+q2yB6W9
V4BMHZ9NN1I4uT1VByjOkuynQSOsBS/LnEfyu6uWaJs9t5dT33f7si+oD3LbQZyO
ypWk2sm4OvvXQrbx+TpnLvKJ3OPXa2G1PQlA4Fy1+0h3qc4OI99hNN9pGzbJXPVv
XrU4rve6+S20sI9FQZy35MO7OTpr8mDjOz4WyU9+9FrOOTLCADklyP6OJh0wHf5Y
Gib3SK6Lym3AkvG9Yhx5O+zJ8DkaE3uK1xHCqQ2m6jGvhy5XfG+6HQ7hCMlsSpHR
biWs9ysWXUWoV/SQrzDaq9nx64XZ+ZhCZdQQLfQcaQpVVeh2E+abdp3CTpfvmxHT
qkj4gLVIW8qGmjrQAcVI4nhDf6l24XQijsddYRBRPDCGGbEUndR2kWDN8RQ7j3h4
jYYPpxuJIip7EikNoWk6av6z+DtiAGAm+sJDKvMSMInXRvC5rUHrysdXGM3jMMa/
//7yTgawLyKicx7PZhto6BVQwyrb+Ot0yQ4i0KzbNcPGDHRWfhv/3jsOrTB3fojh
mxdR6q/CvknUs+XfZsMQQCZFekTr5C/xKlqrzWZZ0xCL/34LzFGd2TxQaAoakmRN
CI5Oi6VO3D0tPfy3tXJ0kjODu9dTgapu5nHcguMVsGhIw1JljvGfYegIdpIwYyp1
C4Qq+F8T7pjnbTjOFCkc8RxsJwM5hClzgW3+Ai8tXSw3/uEdtZfbIurvu4xxMy+1
AT4M1mInscBteR33rRer32E8W5LwfLHfJziW2wFX6YQMVFrbUNpMQMM/cr4js0qu
0y2669sXmpoY1KCCT/TKs6hf9ToLOgNCPk6QUWzsSn2Kh1Q++EPMxyfDO301D9Lc
kbWNMvyduxclY0SQMeaNV3Be0dFjgBi75DOrz6KxcNqnc1I4FtHMbyNFPHKueEUN
N0UwlBffq/XUCiz5ce6OfGl8wn8wSEdaSDvldl7my3MQ+x1C2S6UJcFzGrQ5X64p
QFz91i+klxYqmyctr/kTLj9cL+S1eaI8+vPlUrZ/xtopcTVbP6lRXHzGUB0KqzPn
tLCWYTpVkZhNopAG415YZuBLaADcuZ87W7fJpo52whSsVQOYUpnVCeN06ZS6VtH0
EZ2xM97WONOHghLEsUO0MqSQVQhfwTE9bq2L6UBMJOa3UFbl99LOahKzS7FVMNm7
MmnKkAaPpsYB44wHw7zbzdvo6r4Nncn/oNCumuVu9t5spJstyhzP29JrTiMo1LQX
vNl8yBPu+o6ZG8F+4PptQreV08Jhk6ophteJNfXvilbjzqmnXopUDyXSEqsWfp5n
H3ecIu4pfnf+LDhvJeMVZksxoOtjfDXyDpgbUU7rwYIdBAhhDOlIJ9/msJfSL85m
9YSN9Ob0sFP7yxPyGcNJvr5xhI2EfiNkQf2c8M2TivIYTNiEuitzhmDwnQhKqWPE
T61LGCBDbf9Bq6ojqlNSSL4e4rQSRVhKtHGRqGpElKrDYAxNYhBXepDoTzTlshkM
6Fmc5DiY2Rziwu20m0qtX4hmWbPOZNIEZditUK3deVTvnx0VNycYDNsqNv7x5GGJ
BGZ0ubvZelLXzmntJMwi9qLdXLCN+POfcgYwFlshOvBhpoiSAfgtspXT5a3zBX3E
K1cvJis0zBQeMM8u5SGaE1TJtF1FUQhHsqLk7b8VjeyONO3L+OFAuKFp7P8KYWcf
RKnGlJkRtLptpHPdkXaHDqcMMouVgQ8uIBcgbYn3QDsr8jyqgDALCFZv9sj/or8c
dYPAxcpvcRDz+g08iHi48CEslPjRLDgs5VvedlQdK3rs//fTX6MG/SvwJnSNUTF+
yJofp4GFRbBdcFg0UXt9mau6RE8inw9nmwEGYDjnXHEKu5wcKhsEpb2QeSX3KEYe
pPMZo8BUW8g2BziK3hx2rrCO2KXkG1eBiO9ufvqSQwB3GAFjxfL17Dq/lUKgpgNA
2ukNBLxDEYpLuy1MPkAsROLcu08keeOeAbLKrBz5vBevjLpx3qwXCjxHeumu7rcD
4uSUgFxvvUPfsQhThNt+0r1CcRZNw7qc88OHPNJTSFdk3Xs/khWi1XgXRGKZAqou
Tnsgpa4XxZVR0cdQQNTR/SxkS7pcK62BfTL6q5L/ZVBntues6Im2W51yodmD60iu
nNkoTTA7bU9u0k5ujHyRimGJqlCqKPwcHv/tWGMLZYyEnYUYvCwYFBRPyvSQkMf/
aL1l+hBfSBABbQDLjjXd8mRv+3nWWvgWUit5r8zqDpBD7xlUROqKG0XmXxFvhCGE
DTzzwkPP0vBr1Ek7DArL0AEXm2n+qvkFwvtb/EBcmQDjEuT0vinxklerGMolHhhP
uG2iC4LYyqzsCDU0eczJQTq8njydR4G5f7PoNmVsUeGvDR8nhAu+OPFFjAwt2Spd
diRh7Q1cryzQf57OCe+0/4C9CsoZi0oOdtnDvQR2mdz1zD4/K1fjHNXXPrUByyV/
Sz8CGRBc3MjsqiJ4qlWLvrOfMgzr/RlSLOFZ/i1hqQyc/tyxhNtQqMDnE8puNNII
R+qrgSBfcskSXzGQvWUy18Qus4UWnMwly1cO/W6oh905DjytcXQnhMXxjXlPXIMH
JpGY1+JgBFhEANbrdLMRJcfwj0aGZf7dX9Nq3wiacSE+6rHyWqC75s2KnNmbb0rQ
DieUgk55wvHsMblW7cy3cWn/If0DLcWHZKK9MExCiVJJlx+7ULJ4BXR195yWnWEW
9eKjEkS3fnJiA3nrsefQS2A1w03zzEeDhlwEmDa3XzpqyF6lFshOi2l8dbfXXQSR
kgYJskiBxGudMO1sw8zFCoHiAxkBohliqTu1wVmW8F7XEU6DGKdq3RksMpfGj0Z1
5qXtOEJhdALaQYSAooY7mXK9eMFRcdnfLOel0b6VLDIfJUyY0TLF7Rd5yxUnnbc8
Ya1S/J0ljYy6rIq+LfOoLLBLQnCTZfSji94UtBRaCYb/hk5ytfNQ2n5pMj7rJ+4Q
2hdywdBS9QgEwr4jBCD/65NkK3gyM4zKONRrOx3BS5R7U3oD7W6WFdJdW+HSfSrv
LPK1pZ7POeT4XgPMT8sQXqayWl4e/hUpn3qyA/gbqY11J5874eJGo2n3fNzFYbn+
ww7GiqJcDK9jjBwsek1gHmHTe2tG5KBCrkEO+qYRZYdwAZ33MbCEieM7Zzozax2h
pXcX98zATjO4D6dZ/Y8OR1cmc/xgr5GpO5L6yRUtlcfu2ALpZpvSKoCFHZATPPiO
kXLW4j/kYnxg5R3vYJWxrcedfowuwLzGixuDTTCAgd6xmw5nTUG5k3G+z+x/3dNF
ZTL/9H2BomLh4IakWadpEOWO5ATZbnkKozzJQFso9pzuMKmMMIXsT2D5iMqIhhqj
bu/qprFDtagenAkIyQZ0mO0Ps1P+htqLZYHoJXuGh+S/I3txbwXIvaFJ+alu4PNL
MapCiQLFQSrSB5YgrSSukJ5IPOwtAmG1rbaesSLVfuCI6sIrvatTJ7LgBGo7AyXZ
3IgZQcFStobbkw7Ua0qqGa3Siejl3bceAEyo9qKQO6lYE4oznmJQzLq2UdJFeWXC
344BnTAcm1haC7Gi0hbuh7mmccABAs7Iunwu5zisBsY9uGk9w0hKsBtveHm3RaxE
/Y/IXv/N00K0cRmWMI9a1XoraqprIK8jA2JqxDEkFNpngiWjorROwYQY4pvCb6yz
0g/DUqmaQh7SWyZEG1hAJuuK81mow9khbKQX7q1rpCt92tabU7OH2TaEwNF6yNoH
+vbGFhvY9vWTPDKWnj4dYEbEPBeQMERZVemJzFGm93T+lSct+IOHDMN3IwF0x9W1
YUfH3HFGOAcRyWcrQY5w7g99McNOR1xN6OwpEe7hzVuioejuTRLgvbjyTwyqy3cZ
vjyA95qn8DOorCDhEwh3TW/PJyhnQJAVKUiH0Qq5M9ul141e550fYet1I31ZXZgA
zP6ykWNVnGuV6mbXk6b2AuQwVL5vNHjlBp0ZTAmvycNFy1QQHjbkPyrtg+XtGs5g
9g+KKr9eKQQjQS7DpzBNlu3GRAyQiKcoVNArkAr+S2pHxb2DORxNCFP+U8sVJ+bM
HHPxRGMy3ooztjWbpe/y3B1zF28zXHzb0tOI1Ujajvn/rW8jAr7tlY/N1oyqiTtJ
H9sX6ZVZzDTt6bZbrrU6+RUQJMWQl617nW1YjFW9oT00Qtw0kuFJ+zdHpHHlPIsk
uV9WVdsw/dkopWB36xGvZtjfiOAbtn2lB1NCbyDOiYRNjGLm+ii1X9RLay7MZmaG
Gj0IAyoL1TWD3iWWNN1u+rENoKldGeoSid22dnZa73s3w0uEFbcwI8IY9/ZZgcvn
wyECNkZs1eMKiejbEwx+wcnNeoprD2LneiSCxOvpoTFM7xHeqJZIf/khXBdXcb4u
mf957ZxeCcIYWp7WiI/calAyKuzPR5ipA0q8f8HwLrgDJ5htim3lIlUxd+aEd0JF
OdJ5SC2JPJbCa/bbpFCT8QKnO4SUThpP62KK2dLYIWqJ60qBXH8/ILmSlwgulaND
S9ETAu0r7nyJJ4eNN7/brhZ1ufCHrDgn2Hn1q3g56SwfICQY/pvbTBuZxyoCFB6p
gz5ALfhpeAZ3FGRZ6T0XfqM5mZFtFEPyvDXb+QxLKWSPMVnBYJcE+U2MAPbq6dLN
OqzrYQ/zIM35/TGScPPPPZNOZkvGghOUqVjTFtDa2UCRD9IMJuNNGtH3eHaDmBWW
viPwDOlvjt9yPMn20ZrM3oLrKYrTCotOKSkwOuo9kEGR3Z7+iXi4njrwlPmaG3/L
zp2V72Z8x1t/26UuAAzMbmD2000TUM6gXYIkGs+roUkRh3ObOqTfccrkIhcPnai7
xG4kPNCp/EujLt/12KOaTO+/AWmcdPzJ8VofiITXY43Z896Okuga/QbJpkxwAOjt
nw+8EleF6boTjGXOzQBoOn5J7BdOGD7/ad88cdkDX1Hu4snC0GM53tx2XRxma9C0
8G2JmFs2S0BOqvizbXAXRFHpxjfE6hxInWAjETqNdg3lbyxKv856botDHhcQprl4
Y27rBQ5j0IQDh/j6bpQUSQNvFtK+ElFTxs8r7sP36m5zg+y0QwuOp40R3xqBN/kY
EH1rpG5H943kf0GD2pwagKpIiGnb4rn/ZqEJQayIWwkC6Lm2M+P1o4RXj75bX8uD
wMpVGJIrvgfJ9JfWcKEefEcrf2vnzKifuhXEggwT+WTuVMYmFNDlNlvI4r3XlJbQ
cZ2Vr/BYdvau3Neu+Q4VFTdtN8uAfCZfjMS8CH0xbhoh7VuSFn0QTDAMN+v5FOC2
4Lx1Kp7fSiwuGRT/KJht8/g5VAyqXStM6gC2OQhJojf/FB6hFXRvjMehMqYHkJZn
/grYgl7OrNzCIKXCk/VZWCzfRiUL9glqy6XVo27OPg3pjDtrfLQVOk42D7s7YqP1
5YwRaf3tE/rZcl82FWqWlAaYi+q+Z6T0Wp9bHzjFIF/peSV9KOcLeQaEhEAMN1d9
QhuqgmMe3qlT0Rn9kVCeCgJjVVkQf2W5yCAEqy+AqLzzxXXNpqw1pJep6EIdNkUW
6BNgTvRUGijXelx7Lke62eZsq738pvlk1m6neEfRvwzZuWaQTRtyunZnixHp1X70
Y25y3y29Lavjl7b6lkYWyDLJK+X6t9ZHJP28KJLfaTf4+zbW32o/v+FsGI3uPRDi
N0i1wjXuzh7bFJm3sr2kwxzp9a+g31sN8Pik9MebTHyKL8gxsjzescqUkX5F/veI
l7226BCuu2A35FGcBHR11NtqZxooNKfG058kbY0b0V0Hstt/P+WQQeuMJ8ByH5hH
c6bij+xGT3V/03tbxdlnrY05AZd8azEHI1lNID6wCRz25LGL4OJWVAKMEInG6sQ6
6+F9bzj5a8InwUBLjHfCAKcYH+1Ch2JCmwHtGWFJs5hPb0VYagjp/X1HjuNfBloe
O/IC+UskVqnKdWUff+1MmLkGETjy5D5siMz+0oWmRdi+Wnp+tes3tdCvH/bs2A62
sLS376vxkPMU7ElufF+B4/viK7Ssgjoze1cbpvZwvTDZy30C5+/uvVR7DRkFt730
tH0Y+Qv0yD+R/No+HALb54zi+uGzmtRArvOFyTP2afWDLIwYksCpVqe6TuDaOcxk
Nl7ouzdrvjsbuz4ZF4sQsc4CqgxgjtRWXGqtMyv2cpj/uhp8sfAkv8Ym4PVDxqn0
VA7KTpJLnvD3pUS/RT3+NHQMnFn6BYM2UEmkpsx6N3wwCgzgpS12lgnY1/GNnzhu
h2+p5Oz96vZaIQIxRZIVdCxG+goJa/4LsFyDwi0ZZiUpHHGJ3iiA9IaeJmBPeN2V
D7BVgufDmx0ow9cyJbVHad8u6b7dVTBOwPUcHNsH+jZEPqIaKYWioD1jsQ772tgr
Y7m/D93dE5epvfonxi3BQ4CbNntVmD5vA+q8xUnyDZMAFisyZSQjY0ecCbxn+lu2
xPnL3TNecRy5tJduqe0xcIIhtwhUV+1up3dAy0llSEoKpIdHBPx3C1wwzqydEoUe
WS82hRvf3aQbuKe+7DuiRALZMLmq9tGz09FkBPpRBtf4yFn0/5HNYCLTzwG4keWu
2stq0YcKH9nATTyWQEG+0StkfHvD9jsi2wJilrhwNodWjC5SKMSJGEOhL4Ojqcrg
1SzlB3eMwz4Q/mIn9Y5EG+Vw2W0s7szLyiwaSxFPcJjtPBSrQs/mG7N0mIFnaLwR
TCT444rBUhnAHqyZdRDHsx20SUriBq2ZRy7rBTjSLyhyjYeSL4XvSdMOQFJ0GX8F
2BE6rbJ9rDkV/pIHHvaGGFt+iYDP/Lcv21zz5yQPytgg05hT9/iaO79ksH8BV2dL
A6JyGW34fJOjjZvdpwgpplgccJMpyaihW1nb1BpTaCrBkh31MKCWyknFNcw+wGWm
8DzDD4c3SGi5w1SEKvg1eAVjYbXvJLFl9j9wDM9oRnEyXx81Z/YtxYV15FZCEgqo
41DDd/5PAYTLOE3LMpua5ZUInCOAyHgCkkZ5OtYS9lzXilIpvPMIxLA6eLpO3a0c
3uWFcC96hI4HKsajJvkLyFSfFHAF49/yBX1XMSiQT/KFlmetry18yTHNpU+ABbNM
fb3JZ4oRLgXSdkXeM735SO8rDsovdo7WzHKev1cadj3HysKP6J1lLJAVzd2wz3Wb
jK+yt31MXzlFZ3T5JG9kdHlNYCRSNE2z1JMWCscmHaX/p71c2mE7xKJnks5Q+oIS
sFoK6QyGyc6dDBmHTWFUVfGUrbe+3gXH5n86LsoNcdOQCwY1266S1kCfovB5IyWk
06aW009GjByjDVJIc6qUj6OAZYKgE7z+duDBcyujRwV0xlsa1Das+ZLohVsdVmS+
18bpdEnZa7tIvy0LF/Q3vCNT5IjpEYkZVgEKD11xO9XlxT7oSaHZsAhgWnufIEAn
nLAyuu3BzihNBGs8dgGqGGcP/WLwsUCL3hgCbguc2EUWx7L/4u3GQZy0UhR/HqKL
6rUeIUBMUdza362VWnZoZ79hLBIGmfTkwO8EWTo2YBmf8+IaN10kOSomqWSsfWPM
VXhTyLQb59mxHhYGEf5LBeOUhOO48p3Fl9CIMadgXzDYtSeEtF6cTPGqN53VYm6Y
/Wnbx4IwfFXSVtTmgXb06QGXlAuy7X1R2LksHd9l/kp/PgxZ93RtI+c26wSiUbUp
2GiEQ2bSKgqsNiY5z/OxGbHd9TIzjA2JSFXMPQiWAZn5nwZjxcT/5gufN730gOLt
Sj1u8GWr/g1U0bp1avs6utBZtE3hrEwOdRUYW+31fJwZPmiU+0h6B7aqbE4+lJSM
DMvsGa84c5WN9+JPy4be8b5qDWqIRmLuO3ZjsCTTUXtCIoDpqTL8kQJbz304tA2f
6az9eMEbJO45GabupAN4zR40s7yVIxHHi49o5Xx9quTirvxZkUb5js/NDsn2ZhNW
vQHGd4QAqQGjwM0c0mK9BAbH/z1WG/cSWAwkpmQmUZbV3AxTXViWyOS0QY2FfFYs
BxAhI+TVTdg4/La/X/OVFYyStZ+6ydl19cqArooY+79kiqzxxBgRXCADv30u81f/
NfpqfllwB/kUQrA6SVqAjcX0V+G/ZtBYctyKgOWDWdiYW3+UIdiT2lf0JLeAZYTT
bALKUzsNIZ//057WB0P14KRF7CxuuY/aq/YyBkWXNj2wwCIuSZ7tx1SXl/3p5M1e
aMHIoHlLcVCjWlR7zjY9Tdt9yHdH4zU0m6QbbAUnZVAvY869kyBJIcZQTCrBQlqS
FvkVCXnWZ9CaQeyPAnXhJiBlIL0PoOJCNdOMNYVQ7XCjhLuORwpTgx7s5oJL2X6i
uyM86PERBx4yN+b+TJWHFDfcYxdX+4VRoycLxaF6Xt8Rvb9ONai/qF4yYV4zZKG0
1Wh/BHxL2HRNisBeynjVbwRHbBY5qkROws992dlgTG+4wziJoTEKvLrtEVszpq3m
DwDQnxA/fmPAbmFXFAn5Vq4ZQeKcX27LH8Gm+8uEmVGVmCPMDIiE2SeDYwKoOT75
zR/1Sm03MlOYq2bNk/5IiDYK0O9XzIEn7FvWqunOTrmJmfsOsgTvOBzfZbLtwWjk
BzSEtRl/j+v1SulHAYPOGTv3TJEFj2uPWbco8NvI/j1TfgIaDmuoKmeFyuPYp6QU
34vJfoYlqntQW058Scp7cPcxYPa25hMibZ2zmHLTnKTsp0/hvdjnqkA5i/Wx15Kl
I1a4ceys4yoCTVi8+ruxcwLNOBicg8UYO0lIy5cMAJFrmUkgrJEFFHAQPn/m02wT
92RdqlRpVQcGZScy3bBW6KB4wXAvfbJuxSMvtpgjvy8GIXEIJqYXfex68PV5KVY8
1zbhrz7xiUKUq1rSg87N2HP9bgbrgPRTPTqrDlPbV38DCUYeF1HP32bvqnvV5DCt
UFoUmqNRboHT+5VQqI/BjwB3owHdUNWiiqER7G6zMjCXjrLBbUzu2I+0FkzZeCkv
gKFylYVwUjwRPkFtlVGJ6QaYodkz9OvfSAeo3e+7SpbSSBXzMkOyPUAvbowVQfej
ZhbbJ1M+9+J+cIi5vC7FdbNEvCKfETkbfpE1TBqkdaiRBS7N3ZVxXMoEsfrVa1Tw
opfN9Pb0St2on4dgNjYC5A8kRZO094DbOiUA+R83EFerjjR43QfuS1oxRQbwuFjh
mmHggG1QQJC1GOAQ3f5FhGVWRhM5bXsiiyRk53BBmS2VF3D/frMmnNAfn0CAAuTw
VfjzN9LR5JUp0QmwL2LxdH3XQvy9K233kA2ofKC3+Qpxo1WCAocHYHXRya9qC2UW
UnD7FQwC/ma3pq68lQItmDHLMOCgwvW0jLXVFtMPRdZoEGeGZn7gv0J7UxzNLlNV
27tT5+2ps5M4qtYWmceeajGt/JzrVHxqui2NuFfuqQFf9ZZmV2d7KatX4Yc8M6wf
k6w5atBIgSNdQcMMUCIT+T/XwC+jGc8OBOM7XXwENf8VS94WqZDKnflPbwE2ms9M
RqDQmd1/34Emr26xQEAAqcXUX1fc4xQU71nCUVf+KGwW4+8RLEPjNZxn1BvdaaNR
X4pqMhmgbb1zCDQMFr5eOl09ZkY1LkXU1XT+15C+y9hJdpyw843AGJqAku5pBvy6
d6E9/NGzmYJe/WkxoG3TY6UkFNToQHz32sRpgAUN+3RxYcZFzN7frgqF4N0yecPc
Fh3VlravsUojP1oSL2F08Cm7woDG2CAqGlyhv4yHb8KiwrqU+n8+WH4mBsAwbC9f
m8/XjG44ujZ/RjNs4n8h44ApJ9e+6SR0gPmb7m9AD9LS5pJ9jj2ZL9k/JS0pQtOu
zSczDVTWyjv7/48zbNEF5++FvBvvm8PwdtaHiyRWIcZ43iAiY+/tDUC7UpD86WJn
v8ccdWVBkHx+cYkq4+QmYBionGLs0sGb+rccUf/7BGIzzudW62qHW88EHsFKb6ka
Wp42ISz4BZE8ORvZUbRGye3mkdx9LTtBCPNEYL/09SNzWo6SysY9CUzjI94/d/Wp
NUm1WHHwOx4XBhGtfsZT45Mz4FU2v4+6UIvkocVQP+o3urCfRsZyV/q0xyZo5HfI
4hlqDhr+02U+HD40kFuW3OBWnwoOiHwI51fqGAemWcRXLC16NRbegfQfZ9Ly//MP
292VaLGDPH1G0FE2+JgJPiyfwtPzoC6Eydqdh+VpABeTj0UTsJO/JVgKXQuGwlu1
BMAZr47yYguCPPNRnpcCd4YUqzycW8L4iWSoR8i9qvye5wTpj7DvfckCeQ0xgX6s
PLZel03ARBP4Cr2lh7iyftbOoGB/fSCD6jIDqC2ItYLQi9yVGXzX8tny3vW9ohPv
rAIQRJmKNNyKDRU9ljW+fXDt70mpaKQLYKe0ltjoygsHIuKJoNpQPa4po/zxXJpo
Nb6ZZ2qYyTv2cQ0sjxH8x5jU2ycDFaHuMCiwEWfshz+MsrArLd1pd+FjI0mriztA
an7odW9hlHnVZQQKeEruDn6pLCy6/H89JiQtZRuyue7oD/VpqtkjWWHSGnlGxq9f
lmBMR3wPaeDyEWiM3WpwjsHiti2A2ZDEjHd+O4DRDwDsugKId2w8ohmGdgsdsCUB
joBnyuE+jLZqWnBfHUTs+hUNObF2XRULFBgMyU6Kovo82Iixnntk2Nz4K/dm0G24
D6RPKV7tmcB1gedgEMXYbG1Cm+6/50tYAhe08TGga1ZhHIf5wWFW0QqS9iGciWeO
/60SX20ttUkNrFQxX1fq4F62UFM3lNAhWEg+nEDI46pmlQ+dKVnlhL48cvRvWnu6
6MjdQg6Tpc6hurfignzy1fAw2N0LeqCIMB1RDKT9E88KVxPHMbz3lF4N0oGnBxim
fn4V1A8XyOZ3lh/P7E07MaBLWCXzz2LJmn3I3mooKZwgjOy2rZWeHdmuJAerybPe
KtXjjGccDcHJHErekjCmx7BT192VkDxGguASpLvkNYQbi7B+fvlmUFtMAPukLyCP
Ke2+gSDRJ34K9i4dI4waOpeBoHztjY7c9xMALoMK66pPMKRtD2sRt4Kg+uXXLdmG
KmUeYgzNJCs8BfAJfq0C8IW1jp+yfshxjhdBDEyI6KgSxo9gRY56oyjWoGZdQBsQ
LaMHL7DsflXK6SvcF7CQPEXHFOO9xbB0RioMUSlZKJymSWvCpISrMrqO9UAHEwUw
Av0Dzi+wT0jYpg83DJFeed2jOoVGdxoJL+wIdjGOvQZ1/znM2B63k/1L14IlmHh1
10k14E6cUygFHEdS8pWpAQOoaK+TJD66mvFRUcXx7jOdQJrMziShaTUPNEFuaqoK
wrRaebf+rWt1QgOgm+YolJQYMtdtYY2B4BbnsEYpvBmKLjyJIEEfl1zOojpTarwY
rUW6FU91KDIG8DnvJxztkt7Uj5QJYHVqGOV5RGMQe5WEsuFjfLZgsvXfWbidwaZo
5w35wXHj0xcLuKShGeIptPb8FHhobisLQ8dALxTBWNI4WIsE3Bb3Mmw7zfWphbsk
IKXHbqYyTfUJwTrdH0zXqloOxdRe5bIRMvjBpoWtcQ3M37MZRUqiHUSYEaqt4o3t
wLoQBVbcH6TpT4+eIGyKXfhenNHdCKB+8k130DjSZSrJ1Tauyf9V8fD/WmFhUois
urUlJA/83Iiy7ZfL3cBzDcItAuo+WwPj8f8g3DKq/NKoZ3xBntg6/m0KJz+nImHe
2XNheTashNXmzT1m+rnEJij9S946BcDa8ZKbhlpST1jaqqevXkeNPUEAmUtnx1X3
PdQkzFbet6PrTm05ldUIB6HALeklCg7SLPZPAJ2tqBlmRfXuA/tAg7OtxfQfoCth
YIOkfYL9ntr4mgVQewyZEpB3b1OWyLPm8Wijlq91Ie7BOx1Q3opRXkJ2o1uNbOPS
4wCUPvB/sKwUeYOldEXfer8cmf7UibfK/jUbbZeGfdaTd1sRYqGlxI1x23Sz0zlN
niZiOf2FiIIHbqCTDYezYykmLrre370KOz8lGw7EM22mfQc4jueBfUABzSy4SBES
azYmNjkUUx+wsfzjMTGhpJzt3UqQyiEBcV4yvJDvEXo+Wd2DOOMhgIzTH93rBBr+
CNBbmIe3fVSaofBHBJaR/WylwEAQ740DLGRA5PWKfAKOmhjK5Hy1SJlsEol4y3Wv
QLik3XCmeofrimTFS5KP2I1XSkmj8tfTbV5InXQQ1oh6z68qB8wO6fZ/xMvUA75L
U7DsPoaCCrTzW2ddza3GeJKYBLLOcsmBraUBld2cS9RtZtg+qIM6zrfgbiSobSW3
HA8Le76yUP6Qv/E3mcdtv67Pk/DChCRHYHlYDB6KWMxM6sEefL+GlnAS68JufnD+
qxUrqZvPUA5og5U/RLP/WpG6+ZermYYK1/XOPa0yl3YqcG08RdeCo74W6RRLYaEW
orVCta2drYUsAYSFqpUL6OL3rv3MMevb1RcQGKbMQ0VqVMi0jNha6Vb5nxD+4O1h
dHvaN6GkJghp7E81DtA1UUQcuEGERcZAc9FHZ0en5XgU7a8ygrZIEJUUrJq5jqZO
5N5BWgFVa2Q3p3AQKkthmw85jOVCMccHy/Qw4ic5ppCZE+xAUmgpzrLXLE04O98u
jdevicHnXEFjeOZC8XZAtn4lOy9GG3izP0H37uOchHPVil/FAbLh4dnmDUWjLdFP
KMarCenms/lRrMRNZeULwCe1Z1LJfYcmzFtomIHy7ShjVKnuLbefCFmd0HTUEUF/
YJQoRq+feqkNZfZ6NKuFuvI+WOiA2GWmmQXMBAmX5oDGxY6zdj+xGQKL67RYnr3E
27CUwHxXNJeM2QpDLUr4JQ/tyb7PDf7bYUlrNkk6cd+C0KP8cUJr/2zcmSxjXEv9
zxu6oQjahb+yyFoNn3SKVLGybiD2ltlmRDkPgTJYRbT81c0uQSZLaew4ahrNsZwV
/AM+r+wmDf+ziVWgt8KV4CYDEm+BCZNMF44eMXgBncEklyvExKJ1w5TWSIv9WV2q
IXxktx6euFLgYfU/rB+W0Gw/d/XUUCgLuXRdxGHS3zVAnYYspelTKYrbpTMgayEP
z+xCW073caoV2QzFb1dZdUtpA/pacCIdvDZ9eab7F2uYya0O14Eh1/DuIoQWLLpi
5uNv9j1NNH3YhtkviACdFP9i/DkhHRpWKyeLHVjsVAYxZ97NpMSMZue9QU2s8tww
ONA5JLGlM1RBX6TL1PyXqFh1trv1bqLfJ6Y3Rl89DY6NNcsfh6zM85k5r3Aj976O
uqcUtS7GKtLoQzRsMHbhPlsYM5Fq6DRrzBdPutSxcwMDYKaDkDc0qyAycj/9W3XX
x89V+Pi2uP6u8gF5L9tbvr9f4PaKQKRuJEEoDOe8kv+yM1KlQDhgjUjDjMPhsLtp
OGgKxDn8R/JJFn9/ByqO5lAY42LSCLoslsnDe7F4gO1kkIH3A07qmxds0vLNzbWp
+2sG2oaObxdSnC229howZpC5eu2uP2h+90dcobu5f+5sYQy1hFsymh5CIhRE0RCb
kv7fLQIizbOuOsfPylHbH2DoL0TzfsJqe1+qjjUrOYC4XBw9/WwElvUtBI2+gHhn
v7CYwrisMqIW4eHzWt0pvaX0ge+dTdxU7iCpq+18/T2jZ/7VJZ6YcDVCw/ntTNYC
jHkk56GKoKOcFkBfi/zaFPvP/Kh8BIa8zI9WtZyoaKWWxrCfikI0wuZV0OB/dpJ+
qHOEtIdgS5feIHpGqDZ4LSi5Oc9T8ESI21uqXTK0TYSjeLnytuAS2d7LTzT7nCvr
n28W/JXY6rAPGqz+D6nRrkn8Ll8ZlP7/ewOIz9s1DnoN7j7vq9zyzSpf9rkG5Ylf
oEDkLognbneEcqI4QsENjFccqO4jYsPhTy8sNW4nZyoYvEq1e/oahpNjhjZ267l6
GhRLXhYshULzMaQg6WtsRFqWIlIV1AbKJ3WC1umO9gPvWncUYaxXuGEeu5SIaZuM
q6HLpwZIlU+TiJoy9Aq7i7uJWeCUavMhBUC5TcobON47S2b0P9pX5+r+960XVk1H
AZLiyoY9ySft1VAnn9LBRZMTDANeu+Rtla+wa8AHpw/8cL45gvFxFN1RAHXY2Nz6
rr1XZDdjoKPEkjBNxpbxQ9IS+XMEudNHhfUrdwcR6Wwln9Z+5XsnY7EmPkpKjMgJ
q5+nUC9FdTh9TASkcM57nlq3Sw6Yu1HY5rDENkwnkh1+OQOf8HF55uLSvnNaJati
fjw8C37A2NelRySmUBM3aicZ6rc8DQFqgj9XmyL1q57ptNV1AjiAaS8YTd8I79W2
1GmRjyLBNvsOiGa0gU6nMWDPnIcJ1GXQeuTGFGSAqdukOr3dtB5qHy7VT8/Wp7yq
DmWIWBElH0YkurcCpXE8YqHkUkcfHpKRfmfAyyjSGXJt3IZNlQnZK1/pjl0PNSmj
YU6sN7LBNRkE62V/EOv56fTphWaRTX2slktafJemEQcBpvufE9X2eIACKRi+XPU5
aCCJoHuY/9KG4+J0gFI/bIZc1qcsQDXbowdYDZYG2NqpMgvTq0rcI/h0x7BBxcBp
JZHxnhBaZqSTn6mQzlW3NSSVrUQlWIG5x6nkeVe1uwZQCrv1XnHMPs4w6phWoUbU
poieTzVVlSLYaFW0tavz3vuFpxPP8qZcYe++uzRN4CSMIFKgiSKO8Gw+sGumoC45
OPH6I9vpooGi/friIPf/6uLuqZono6uW9v8qlbbc2M2ZjbffgGLXmh6UFaiJzN7e
UfSv5O4njMOCs0aNKeeopGuqw4vBnWN0vShOj2V+2tMruxhzUpZkM72iSXHYadp9
jVYAT21iRj92Jx7egWS6bwc+fleVd8mgqysGVZ8U4baFMyvtkI0pS+AIiXw8/ucE
9tU6S3DrAqrRdZKqt71euv8WMY6mWt08++p9GHElWdZezW3gCjmALd5eEv9t1XeP
D+tFMx119i340YK/TqY7Q3VEKOlFTXzYCHQToXKSyCq2VCXwcPNmZWpicOb6zPrO
bdW9IgaN+2VWpoDnq2mGNFtrvgw0t91vMRGqpAdlGyXNRLxqhqUm6Yr+bksBL1wX
BFOYRmH+jTOiL+2BnB9ddtR86c3JRJYJagDDWlGHlA/WtJRSlQnUjzCZ3q7YmnBF
Zsk2qrx0SvF18yJnh7WdxJc5yzYSrAb2IxtTDjGPvojLviABBmH/3oGTr66k0ffb
9Z13w2sUiznmfZHTBmlhqfupvKwr1+Ws/iwFrPMls6ZZ2ptpbLHiQgyQIU+hOakq
EHpNJ+X70DNhSBvsFMYgUqAW5lCSXxjJR8xGtpFiJPq46HD9rz6SWdqKsZMWJS2b
x/BkaWCztaYkDL1MjJom7UkPTuPDq0lnP6b/41aKaPA5hdsUU5MfBuOBBbMYS8Jg
i/YNxQJC4v3Ivr8kC3e+YGICZRYs1Q6Fu8sXhQfR42f3MNp+WQBpkTDLxvTf/5QC
y5CujOclEucxx1EMpFw+vJDfamGy8Tz+mW+k6Mqv3wFf0XwSUAt6W6Z26ZoGBDYp
vASvHA2MgopYhziScUND1lurJpL02nL6pfzXYovjYCxRv2t6r+8p//Z7hIxOb4Tv
7vhlPiqlEHc/Gss/Y4nUzkGBhposIkBMA27hYfuJA8EbVtih88yCTfB9KxauNpUP
T5TZiEf2zzoEG1yrKVqX1sFReZX6XxzIpzQ6p7NFCIwX3RW7+DLlTv/syz6dz116
0laOWT07sH+VF6i8DKz7F0szuU34iBcGkXd6WPiLFse7xW3wFgrYmlzQanrY7AQg
yjx8Z+Q/u3B/cszC28+xJr2GHZ6XEZYiq8Li9bC6ANeMtJlq9ZAFZJAK8hGJoO2O
P5gHx0QtmyjFqpTsYygqeIm/k4/RF4xAnrFLs4QQVxmdd22XVQrKZyzSF5+fXDwS
pKij6QXp7PV3WLnA7ba1Wvx7jqFAF24/PpcJMEO7RzBW6g4fRWOufZnLW9YRJU6n
X4ZYssHw7Ccf7ai7YBbyByhQR/ewEDmaNEv/CQuYNk0Pm7CAd4ADpNv1oUxdv0d0
xpliygKeuz9ssREMmKVhDGI8MMtgmhtn52S8II9xmRr3jP8Ww5Paot820iQ7a+Lf
FHZowWYuX7qhpE9Q8YArbHC0qjIuVfkn39hbyHApP1Z9f3hx5DAjKiFUFjEqo8Uq
AXQm1a3Hatl2CoHM/0S5hx54mYeHSEgr8mDqgpcV0PYLmqsQLqKXLeo61DVyOrZO
aopK7rSW1qhESRGehy2OFSs4v2SkIo9pLzcgkcV8jYf9d3J0s2sXMU7qzoDYnJdP
2l57nYvhczTFUXe1mvpA5ePVmch4HXfXr1K8jWgAQ7UEaGzHegQSRXrU0DHStDNX
7S2dnOTwm/oFrQOwq3YJGNo4pbxfW5+BUNN1wV00B6re5qc020ju5lHZc5Inqpl5
Fty1rjpL3iYdEGk+D75vJDCd2c3f23IV4JO3hjPiRVDD5IqNHpmoN5Ammku3yKDb
iGUhj0pWXHp1IsTxb5RpmyHpQu6C6S/oEsQGy0riL1qeMGldlkzX+jWtFSOfZOCY
LRRUPr9JfwzK2luIZC6XuoDI1IKgiwDCCsF7TDGPxQGrJQxbU3lFPADbnBl9a9FU
vgVCBRouTKqUVNhIyWAWdv+HBThcIduD1Wf+Kftj/+zbXE6U6mKW0wjKgmIZ4Mz9
nT/brqUo3Gl9/Z72JgRULPlMaNfIvISz7JW+Aho5xIJ2HMjN3ossJ6HI46gOOt28
ZiCgdLL4iN6ZSjuFay3TFUKscYWFiQbuSJOQ5P6/Gr2uSfAE2ZaTTr2KUGylYmSK
O1YqiNa4Mz02dZPDWPGLynEoURvSGeM9NfRJTd1qz0x3y9G4XrrvkqZQ+aAOYIhg
EAqoKgeql9TBlEqRg4yNNc6pTmrZFIcJkIn6H7aI0B4izK7k8AK6OJFZpjr99kdp
3ne20OVcKvIAwJOqB7uzg6yc3uBLv/4zNV4QwhGUJurr6K2Cy9I52G3LXd4pepMw
w8d1Rsn/53PTxarHWKZBm+Cz3Zf2n8lBLVceHyRHxP6jsxnVSteANz/P1ZG4LZbX
+eViV/s8jVxdRsXUQcfru75WqH6Yr8dz72Gbcw9myv4M3UMdd3wduCCqoHbl+HoO
UOhakPciNBNzzf76VrqAqrKu2Wt1KkmPWCWAnZ5AgAwXQt0nA5tIhyRT9/OqHl98
g7UvA0eqTzVGc8Tk8d54qHzb/0XXBqERM5nk1iFBbrvG0zgxLxsPd8nCPtSif9A7
L7jm2fShZj22AvBPyfXqbGVcdRBcC5Z4YJHMhG+hhNQ5Zt1GCtl4abW1KwqZ7KSd
dVBQ8tljAd4cBpdxYUtjfqecVtM4l3nOMft/A7kmGU/F/gOfm76QWXqpoL8Bxho5
LO5Ond0GWrCUfbBlWR/n73b4LCDBNbvzhQA1sQGqfMA4zwQJyRdUlMVu8dVO7/Ig
j3WHB9RjUh46EM2eD5gcxr+GYc3bFR1ZkDP9zQ/5ldXKJSjm57ZiBeXcM0BU308+
HApzKZxERHL8WexazGBTAQ76fr7hvm/MrjKYrXFE2jNlVi7wyV9QToLisFxLQx8a
g4QWZHBWqF0Jectk4+fbMRRWVqmAYj28lqBujui/vE0SY/rt5ssSNqSJD+cU7Wyx
aZFubU0IlZUkK8E3hwKwQIfSIYZGhdvVDo1PP7pWX0gx62ibu6sbrUik0bsiuaq1
Kn9t3sp1N6J19JpO/ELv7//LKt5W/26LFCFy1lv3M2KdTdXzDP+elnz/YkS/DR4i
2Dogo1RpFspsiygs0QCT/fQ3IA/aXLdKaErDwi+DMXgGWEy46Nqh3stwCf73V3pe
6/c22Td6icOimMRbH6KMkKjs/t0IM83MfywqMTAHbFOw1YypCRTXL2gW+/xODHjD
4UkeOC8SGQeiDZ7VABdVlrBgJ0oauru0LNxM2VCit63jWDvhX/qNgWNz1oUK8f74
cFxxyvi8itUtiZDajx7P6lh99dn9CZX7omIGR84X/n7+wfSSXf/xNgkiepjdVdPq
5Wf7m5pY81dJ1iTfrxly2dR2rwmndXlp8mkdK2hjWtDoYGif0jJ9tg7Lr5Heu7O1
Lq7+pXuCLRhTa+P15/gjihzfFzdabVXFKjaT0WclWF59d3XjdG3euX6h0r6jmGMs
1sXo0tQlYMxWT2hogjtfpeJqKaZmQPslCL4DmQsnrwb06Us5qfsqssLgrBJNp5GH
ptfyPjCCDOQdo/O1aWkg8PolP/U4t2sY8ICApAs5ojdmrcSG4Y4QIerndvn7jWjw
tOFWE9E1J3SN4oUNF9aH0hGZ1PDhxTuNIk6zA61yosCCM9HxQeLfBmaYrmIyzOB2
h42LQXyo0idHyzUOvcgpodmLY26ZevMnmI0K4IR63ghF1FGAvABU81VjCaWRuoDa
ft3mIQglCtd+x0hyi+I89NR+A1m1/wY8XtgOpXae4fl8c8N02HdI2mD0B9xrcO5E
EHAqkrlJOnAHrfTS94BjiONFHShLV+IXqAcycMTcU+2juM/C5zEYfQcBKwtFrtAC
4H5WPA0QOuMtHffk6W6zg5T4uvG50ITsfsLOQUZ5VcvM/eWPZkMb+lVRvN/9iGKM
B1UNJoChyjQBQvWo+YNebquUP7IX/V+LmZ0TSmWE4mCJ2l3oNkPcBl8D4sN06nZv
jdtWMEtZaYoHlmApc/7/UK7EFKla2dFSffqz40kx5JcY+zKaZlrb5zILsBwSSMRc
+3qGqRAJ8RA35FaFH37Cg73cccOSHcp/Yh5Ad/ofOp8Uk38tE7NmM7waqsXD/sRZ
NcMC2cEVEMX97yqMXj6sY2IzwN0LEzkmIQfV/JUFTtSfApM6HoKqxdK2WawKs+eZ
TZKEvRZuHQkWe2SyntxXWbIclhl2Gg+IE/i2uO5WNxzqeybT98bpOKj5H468pLeG
tKSWE1bJF1kxCIGh4kPZBoElnv79A9wjWu1YAfvE8vDMePMqfBiXqv2HUe6zYhC8
nJCcMNS83A+d6JH1vrBI2rVK5i8F6gNZvq8oXOX9GS9C1H9VzZa3+kL6ahGOakx3
KR3RBhijwn75W0iwvkGmWoZWEFTeh/BlSmz2IFV3l0FNlf5pWAmxKkalMBqsGQqZ
9KMgOuzba1oRN3Zip3NSd/57cEv7CiNVsOGb8/4kCpX+PAJ15yuxInPEOjvfh+SQ
BINowtFaF0rwGclWyS6N9c8/pIr79pFAKAbmg3jC0kjKvm94RWawcAxVQM4ptJ+/
TKAKLrqX86GO+agSBclO5QOPeJwq/XU0DL7a5tJ1AlzvwD+i4Wuf0F/25RNpzgpA
T49rmDxJ/NfnfgSXiZyVrZ5yCHpJTb52uaCVYnTo99LtHQtcfRADgDG4rZU+NIOX
Cf3UTPWbodYdRLO47N9wIj0/gECCB+GgncoBK48ugE0mpnizJhPX+W42uXVX5zXQ
4myr+zI+r1lc+xY3zW4KIg1hveAJbb7zj1deobqC2qO7mdEBZY6FwZlvWJz6mYG5
ZskbHjaVmNT2pT6xQ86xd68fKvMDrLieCrbVD4VUybO4mPjaZBWPdIoyXNsf3jqH
A7gFUYK6TiHlIMKyQzUyamgJmf/yv1c4JPsTpSPJlo+ESXEuw6Yww63C0DGmDfD7
O7deYBcTo7HW59OIBHG+M8iJlpzJnWb4DY6TwwwZ/fBYV/vLpQ0jFfqeP0aOIUTX
PCLXiOFHOeCtp9HuxfmxOPF0D4M/wd+8LCQiyGE1HyJpIzr4vzkMWu9vB/QAoYiO
kHXnpUUacuktxMIw4ARstxyyk032I9OR0+dTcSSLrtTcMeJww3+UgkbXYSVjqZ5d
AGOdFZXlpniZGzubH+md0kBS0XrIdqu/m5L7Q8Cv62VocBz0hhNsX8lpxKCJaI6c
enBxXR1mx3jiOezGMDODmGL/Md/qrzPne5lDu5KrC+slVqg03oBwf1bDwcYJag+E
SkLD2Qz5UTApXFfx883Ezp9Z/viaumiT5eIfwFTGxVsggffnuAzXjS4tDtfqlJ4X
+BPXU8IpixYBRvO1eLM4G8PY2OocNFFQgR8XKdI/F22n2GjwzLAP5mNS3eslYsLS
MuTiXGdkRWrntoH4BTmKiB6czuX3hf00JMDzNvYct/yLeXJ8aQpbmd4spdNUmiI9
0oPYiWbc8v7aW+tb/0HhH7gXzAntWoCweADogEcigoqf8kRMy9DZbak655WrY73p
i5WZqHZ8lg1q+HBO5zEYcnwhmWZssaCei8Nm8pZLcXsVtWrRxsVdXBdAjIZigrmr
J8FCVDIEYQPpVakfoOvcfm6qPgaBfBwTAd1bFwcgK8K1mMBaa03uGHhPvZ+dmdYS
bLQ3rGdS5cMeHSvL586IAuqGjmL8Xeep05AAzImrBQtG6wSMP/jNrLKlLHFG2Uew
LP5/RPPRxUUg2bCU+yNHeM7kx6H9wMIeFzRg/EpeIOimioDJkgazA/eYxpp2M/It
GpoqsbcB6trySXmQCJZhlkq7qjqoD+InmL3OxNvW68AvXtiuSK5jAuKLQX1hMb62
VKmT+iqKtnOTx7ijsAI8Gx2ydm4O0zbyE2cUrkGmnJUiqvDaCwRtrTePaONe2f+r
kfEEsxnLtXltZeIaRufvYHeEbUoGcrVeEkBgVWqYywKLkY7ogyRSPvtVlJ6MPvcd
ngJYXnhtzoZL1uGlOgzhuI2T+P/LExIfs+XlKPhBESXOIwbmzo4yAPEsniDfydX+
A6j1Wh1LMj9k6KjVgCBwz0V5qLLspHRJWlHl/4f+1o+QNzny/23yULKqYUxVBJma
BNAEpCpWsKwqAaNbPmTR1AzKDuy1g4J35X9kTyEUen3wMoczWuovc129YThnovci
3oXQHaeuOuX42pRpvE5hzTxNjxELLogvivH+w7kYOE3240caGKGD9FkxeCwmDdEv
gAtkEPFs7CElPfXmEGvcESs3mZjfooqzX9qVe9KFJb0l7E8wj9f4McyT73w1WyU9
097N9SFqwoDixA/782czkQew/J1hcjG/QcucBAG4Mo/1HBs6C0viGrWcIT0sTRk/
psYAKyKMMvbPlIwUhEUr2X0t6cF19oI1Al7hIv2mPGUPOmlxFXns7sWXSKNiKLAk
eycqeeIkLw3WjYBRONDWSWp3nSBkk7NV75qoTI/xzy9VH4XHVYGrAsXdV/u0+QG3
7mIZ0eGISIhZ+p8C6DyZm+MfIG4jjNjz9/DZIGsaQb34gY/ElFYU8PcsSFtf08A5
0gg4+NqRbVJvaYvUutTyg4fZvWRkPYqf0bDHpQR14xPy8BwePgBQuwCg5Q9o2BY9
hJrIF9GJ165Xurd0FMi94W041Vv+4FI99khuHiOAAg39z47Mo+kocHhXhicURlw1
Tm2oXpriQsn9lDJyEQI1Xg+bi1rDm3KaCHNFA5BV8y58rJqk8iDIefFIj7BiVD6s
qCo75gIuN8xDr8yCeg/ACTcqUhZSnSwphEqLNkj532xvqnFVAUZ2PkgIYh7r8pWy
syoUzb2v6c1+Z7ogJrGA0u+7p370L8NPhQSpRbiSFq4arHelMGHsBkhWHZmBVJ1b
g4Z+XT2t8+vjdG5TtlmiQcM+0pi2KWzTwyUyJqQg7CwjVPRHjIqsaJJKjf4BP74y
YmATMBr0v8nXNxQjb4X8TSRYo1TE7tSLn/bji+7eMNz2rb0HTLlAXHcuB5ApofH7
wvwntngO3ervRCD5ajGUIm+cpCbrgseomUzS6h4if3cPs7QK7xpewofywC/8vDqk
W3Z9MfuMwk5KZlTP8y+8v4GIEPZsgXFpe4qrpGmf7wYUgNaYzfQB9madYiWtqjmN
wC4/4ClYO7KrwE/StiuMu2OwhM8DK9H3Zg9wv7g7YiiEwvac1TVKjwh1BK4dwW+r
nMduWB17UMQorvMOtKQKw+QmqgTUrGGlNgojotwY6oj6c/WcHJAcQLjQ1WWVwTy0
7CS3MxbsW99r2gswRIQ7GXtuooL1uY0YgPBTCcPJT9e6cjUaSnP3G4Iib3/znt7f
0AulRzYCXjmicEznQAIpv3PKutfk/n6sdIHeYP4JHL3FDCWToMxFNodEEo3C93M/
B859ROwJlSpcBNAWHfBV79ziwq7Sd971tpyg1rwqtQZG63IJ/1ziB1Sj3+k/KJaR
id2OCfc2vN0/476/V6Sys73C3jtsYlYjlDADN7ojWEBj7ASN320q9Z3IOOjRH7It
lLHdO2qEth5aGxCaqcEysN05A9Py2x9EgOm57A+wRJuAlLEICvwoX6wsOOzM/nJf
kx89h2TlyvFs0hfJ+FkNGprT6F1Zsbn/OTgNxvliezpv3exReidkMtRpDlTu5h/i
uvIJImohWACqmvY+L7mEMTzSik8PvWNRhUZAf0GU+CtLcLIQYZfiuSM+qFQZuJpz
KyqULODSdZE4dnk/BzrujYs8We3lQzGwd58D9pFYojrY9JtakbzIMc7pBMjmSttC
J9f7nJRqIRbZ4AygtJuDxiwTrJ/5yZ1yi22h2hDC0F3NxGLcz2VorZOoaqM8Kjqo
FgvhX1V04op/QcQl8r/hLnpb0wgiMO/MeN2XOvw+e9FSd/XIC1+oQe9o+Lu98st3
gs1MM/vZdB2zsuHb8uqYmD2ZBms0Bn/9HB9tqTuJerTO5LTCUyccstecW9HQrzO3
Eghk5d+XqdyMY0SGJ9pccvxAN9OltxaLrGfjg+B8LHqog1nzvmyNmxA/H1jTl3yJ
4bTUEC7xgt++1HPfoNIGC9C+hqHccUU4qPKbkL0emCv/Jmqqc0WSwQ6gSibm/p4p
ZqgFo+yTIYvCNSI5DZ3QFWB5BxRz+oF7MEVkOlU66idoWNgZolGDCpwuTwfnx6/i
fSmC/l3HzctUuS0D5sFVx3xEmaX5leEyYX1XSlGqRrQR6ZFF/e/Fcf6ZIqzSf+wR
HCyEyrLfpjN8zKaZBDGAiDiaUnjsOq9jcj7XQcJuEw/LV6bAofbKVhEoFJ5vCVT7
KiAJQ3S1LJbwVpjOdWP/KflX2BxsbyK0ojoUqBAgEbJLuE6QI8MHB5Dq7Ne3aixE
YAf4ICP+WWX/4VLqwy0CFoknXZPTR3gV/ddz0bJejgL0P4oDcitU5D/4GIxHf3Gm
Jp0RzQZJvmesO5rhGMVdaqVrb6My1Tjtk/d6T1GWajNtf+Ji3o+ZdXqITG/r7DlM
0nKRLQVupc/aUeVHuAgmtog9vD3LvUySPQa9/kKqfEzl3thwL+4sKo+I82nA+ryB
EQUI2a1+M6ObGEb6YapiVei1fJe939agMKuFN1nOanJCn0wWiGjxl3JCcf3B8BfK
ereFlH5JofGMKa6NSVJFYniTK4s5qockZcaP6Tn9LJQe9cWsUg6g1OBWcwVFiIGp
8i38cQhOVXYQblwf2wIAAKYm8/8f7dUapM4aQfGA2HTF9FsxSEJIg1MuM0LzkJC4
kEggbNbrrZyN/NP4OLOiRA1sbk/T7l/gFGmyKdgakh2uQ8ZqwNbs79HRQKEvVgFG
jfyLeyIhOc6aXjjm6dN7RBtIbtwh8eqs8jVfhiB7hb2zo8gJ5Y6YfbbQhk6dQ5oh
w5LZt22flvUh5STR9HygcravysS7LhGQE/cDq8XkHOK9peolZO5WiStK6tENmfQn
ziJFd3O3aCshtTxsjvzcee2snsFJDTBWVYpycX9yh2B/zo0PZxsSA9ifEPLP02zL
NROyLHznvjpIJnmgvSREfRBFRm1pqOAiJYN71jtn9gksy2T185cdBGEufjkyyQ60
U+c76LG70SnWpZ5Na2xRQOgKgM1vGH2XtsToSneTY9eXg748oNMzj1GDlrFxbTwm
hoKeOGAYj6mdXe/GpRpr4f5rfbM7q/OFip4eIYcTpJE6N/ceub/U5JtHSILFhBch
WlVsFSxitELGXOtShPLaqd8FRRP1iiSLlBWlXqF6/5WUnBt+H15kREsuHSUcFwBp
tv1c766ka9x5UCtsIlhmZW3usgUpGiNcfiGQH8JeMb2O5rUvbjWG1XHyfrlul/4I
Ln4R4DYD95iSYGaqn13E00siXfJn/DIwZjuvOtlOLvYfhytEjubOVynqWkPktmHh
6Qzl9k4odCLTE9a884xaMfYsDSHLhopjVqgEUq6k/iYYTx6DDSt3cZxjCmLaHiwE
JiFn1WXqVAdfmfoCkGajPO8Ne3uau/AACzTGHf+UhzeieeNh+vginGZ+LfNbv5cX
44uyo6ZcwO9lpyQXGC3o1u8GjYxTdUEqaBpnhjeH4i8S/Nx+8IC+5+V05mM0Ysk6
nKltNz5+QZ2DIGbOWDNUCJ7TCiPGFk6shaix4Yl466sShGcGPLQBtYZFdL2JbQJx
t6qUE4Pimwx/nPIp6Diqs9KEchB81SOG5pxvU7YybZE1LMXyDypZ9UHn0Ew2cYmx
ihBY/l2N2yUGMTEGi2SBZ+HoxTAW/Mr8SUke/FnAb+L7visXKTIhiEC/GNPEhavZ
SykXz4Elq/h12/qKwHcS4hw1gSb3MKsqrsxK4lR/9+CGIJF9x3W/oHJ3BNe3Nj3T
dUyhsycAWDnlbKyJzZGO/WNv2+Ga6lz926jG+dt1d4ZuNODJReVAoR+rjrF9UVK/
WoAWy2IEEPTA6K4HKDSm3wmzjU1MoqptAJdpo99sbYJAVlOckAwMSGpl4bHCmK3U
xbxIISzhbcaOKd/Gu6kaCVCMiEneBf+NREs75m4EwvZ9id3xA+tjD7kCkrtvkKI1
cXefYAOnT11MuAP64+aIbOn5U1wDaOaFdhK0WOt0aCrQhYYauyfbuD87JpOWGcvb
EBfSWxtG258WNBIPHZC0eGOQexCZTQTBLHLr/IEFjeOAqMyK1kNqSGB05m6IdZ7d
FDOkOLSBw+5x9tF+YTKqyJvUsc3b7AwO0I1VPOn6tioBskEWaN98MLcO5JO54xyW
Q9xJLDt/txR+VJEeV8CCU1bVs0CVHRvxZw4QBplQKJeCBByGSFt9Tjd/7PVfCq/m
4LvbY7tQ67AN1RuV3c/RLsnCjRiEWcEBhBjBH3R+CWI2kB6Nh37eUue3bdtjEazP
zXLxKCMLkuipmeBd/xKzZo5rdJ23oFR3QXNwo6X1UFEW/sbCNCbehnTl+6FbEMFN
sMs0+lfjIWfzOzGVzBMHLOaUNm3Dd/e7poS5TVsSizpQMEA8AUeIdS9YnMnWoa1f
qINSMxGDJlkh8dTgxYCKKdZISAf02OaKt0+SyKwXonXqaPwbXJKXczvBtaZ5qlXm
nMCRHw4K2Ld8yrfIRUh1JYrlzhNpwxunyy07rwkKarU38/DJfMzb5jQpjalWas1V
1ZzITSRpQJr5cFUJjYI5If3NHsWhCNSaezYWB8bexM616c2LuRnV2QsBEUPx5qIg
V/+76wRdEFv65/C2kvS6TaKzBi/XnAnilBUxZOdB2l7pr/k72tUn9vtQvBGaeg/q
swQk4m8mE/6QywQA0ZeQxDzIdF8n5HfQgmOs7wZHVl3VlUOjzTEnBFDc8XiSdbLb
NscsL0ug9DE/neTfPSMWihe035FFfyo2u0THj5vAxasfiiTVFgNOSsMgqSXbzwLU
43Qcg9ht336Vwo4M4k2V8w67O9SfGQQejpeCr5RdvXse/NkjnT/b2Z2z7Rc+vnl4
3sQtNlGLsY6N9ysej9JFTmxlFJnjLQ1eKYOzhtFjgY+Cqr8ATBvxTnL9z3AbgGtD
yGp6Y/s6qDPiSYsafUrZ5NiY3IUFlnoH9rZe2Qj88Ep8iXUxQ0r+jl3e8QdbTjZB
GiaAg3z5EHpOwODQitcf303ybs4FfiWfeRoyNwTy5tpWWjruk0QR+v70LBuind2A
nJxSN9y6bgRfBJ2q5uLo04FEI12rLPagqLfqVTBQaiWzbSx/OsgwsdxELBS9c1sc
ABbZM27fk6KWC3r0dNhJOmhj0hOFZq9HAXuZBQNQGydmypNG5+4DcDlx1ibvBn4L
nds4gZzxhmsBwKCSl1r2pVsk2w5X6N8qH/KOWh5wReCAldT9ysoeEPfewxAbwjeA
Uf4su2QUlE7Ch4MBNVOTIosZ2rYzs1JI0mw/pnOgrY6IW4++qGUwJRq21wHmfKLf
HCft+UiVPVYYbEhaPq9Y8lr14PxwpsMPupcP59HIobqqKii8zL/3aSKtbqltPQXV
6k86EQnolLytkKCONhcv6nAgA2sJhbkm5a745LnyxMU0B9amMUkphGM+tGVaBSNN
gpQkC5bJGRiIF/HzsLfJ7StY00EuIKOrkHS+tU7tloTvRhQ2C+jbSHZ8fjbNEI/H
w/4F508DuHwf1ZLOgtjBkSO8hZ+KNK9j/iOnJfUs2GY38dWFPdydvCSz35J9QPTE
6KBbOUwpECcxho+3L63aDlpB2FsZ0/ep14p1lcXFhCJrxYXWJxYVlGUTEz1yHPqk
1kRG6/BQhZpVB8zMsCJDvg9ijeykFbHt9HEwmXG+yEdX2xZHac18cof5y8YZXyq+
eYyUMXkRJ3e3ZiPv3jswwtJXy7dvCQFMmVH0G77yogWPV2A7Tof9CHPxMjsI4g2v
uRlhZGXy2CtCHkNxuMzMZ9gC9rjmQyteRIamDNnXetxLG6exKstziesmksNYDm5J
0Cy5f1E2v2ArT3ZFJ7wBDd3o8AKoWlwCMetOHVND0byINVvGYmAgpdqMrk51Mw3X
p6px0zGRNIcP5ajvA2PWH6M1BUG6ELUpv0FLtJc57xUux380E4tCzxd47fZ5czsa
793Pmifo5qgcfJEHCC4E33g7p1TbVlI08rCVSYbTAN+jK7awkrwN1WSFQ82an7yi
OirpwIe8zZr5OBEH8Eba+SCxR7xE7W3nQb33EK1cbqxZVkohZ+MClM3oXvtYa6dp
1PANxMpAgq9GnILYJK2gyQy4I8YhC3JEMjFM47L5Lu9Rut/ZqoAkPMeswda23e0W
OIy8o1fOJDjF4OHHKHUK01Ed07kFbF7qje4KE/6xhyK7OgOINXsc1UD9rmrxmXgR
u1AKr2NvMHJ+qEMuApyXlnpPXfG0jemVRTmueSh7MjAEX3SpRXClHxmU70dYVHff
2Y2xEIawKZwK5ihInxZqOF65sX0mSoYE+7Dj7JQ2+a6u1SAqkzAP5s1twuFTSvVr
cuQIuaT56ooJKcxFd3Q7Cef8JILglbFpNpyZn/phDdHwCPsrOotDG8oFdQDPqwlN
NFYLY/ZT/CT3v/GzajfsRGgiHjJ46ffTBCLaB3VRrhm08U7I+0DD0RIIGiHH+uwY
DJ5VNa5Fax8SCUEcKCZZGQsyDzmFmOl2XH8THmzquBmUCdQyFICCw50Laakkm/sR
iSgWxPJSMzhHnWcb7OhAskk4YELrEqrR8QLy4ZWTqyfF0xUMAw0Eg8z/7tUlXAwW
Hpxs2wgognKQaabRPaffC4FEUME0it3AJnltuBWWXU/IM1zNI1SPMe0CclsqYpkF
/mk5i6DQtZUG5fD0lgN3FF1rLWpEnK0tA3QU9eKLGzkXryqQO97Ar5ssf+Unce+v
zOSgVqHepoJiHztNZiIM6wtmGfES6AO3qsGD/2nX+qVQ5bbxf2leLjwD03gctJzT
RZ/ZMhSSC8/Qy7/vr1FRDTC+YTJFNl4h8n6TTw9m7UkclAwro7J0G0LqugZa5jXj
VYJEohEVz9YI915bJqVJ6G5KSBbczSuSLCHIQ6I3PyYCoXw50EehLWkkf09aykTg
9Rq8/YY1fPEI2ceOMNGXXPjU1c8wGKArygzlCUqNcMrVbrXjixRWeozXfJi/bRVv
Z4ntv+F5y6xAvBJEHMm24WgFkDFTGmtCXfXtsNZHOunt4c+X4J2lpakmGTbGT5nP
kPeScR98ipOcBQ6NPjTQMw+fpoytUIn5QlkkX8bWzTTEJpfXqR8WOYYpr5yaql9g
3dPXoHpcuuhbPgs0TwWGAcvALpMoD3F3zGAjmfYEKAahNx4lZp372Ahl033EyAq+
x9EVNmnowTO2HI5m/ROIIU4lf2N/5IQh3qWG4hrhZy/T784iuPC7yBSHS8nVoob9
1DK2FuEmjNecQfWexcM7woQ0k5wbdkJYAKDRvFzrTPefPVS3luTXEUdmP92053EV
UsAxdLMTP4YUCwfUGnlvmRgU5eky6vbm62+fDfhesMXinuNxxwxPPD+NvbB9UIKW
SmYNvIb7rUh7OMRQaiF0q7Dd8y+/5jQMDfTjLRzBtlX63HvPbJ7gZKSIbELv86v+
WcZjV79Z+z88TyDdWEmNQ60544lyw5tfu9ow9vPSECA9nDal2FteZ6V7Kny+NPn9
hzavqgScJ/1cGr2wqOAzvGjHvVjWTW4o6pU9Zpg7LeY++IWXTEGL7tO7ol+RrdT9
II5aJW17YG2B0q38rBdnuaS+bGm/beFjc72uoY+lawGQ2Uhru2UblWNwWzo0u6y5
SwdSCzCorE+UMMUzqkN05GOjW3tp4NecePfTRy56Wv3DD8inhTP4T7zy4HbHK8fR
/yu9MA63cZu6GCGS1UvPbHSzA6XW+Fx4p1arLh29hkdbFomrIOZ6OsdCwrSYKYRo
IBJIJ1N9jB3rScdhb4FO6BJrEsLTXkEqHU722rp7tZXwFaI2U38gOO9ioue7l+Lv
hwUZZO2YlTdcMyBpk8e0O2nMfszCCMi0LSdaGIJvSymkVxboBsnDfN2BqlIuFSjz
ToTAyzWfPWQBbn2A4SyeDnORumIZtj3TaXK5Am6zOrN/L993b02+ITH/R3mgtE3p
6uLsVhUrP5491McPN+YM6wi2FmDA/Fv27PdfYCauYicShftJNjvrpxxBgpbfXy+h
RB8Strn4dbzdYB9DAOb3rZHxV1U+RQFH96J/ghk27ScE4Gcy19Y0LQxw8k9QZxye
Eg6X+kEAY8hypXeQK3ua2t+vhEQeUNwwxjm4rpIT0dBiZ1GAZym7HunumjKaM6Hj
2a9uXh+HItafRk6iv1xIX9cI0lxsyVxbctOwJSPHkwQuDf+BEB7PoOz0oB9qWJXh
mnW5cnEe18VlV4Axhc9f84d2SjH3CkDX1H8AWQnwppNtp3PLG10F9I+IS1rUweEl
zkQXazMrL9FICvD2Q90z8caR4yObKXUR+syLFK/6lOypB3grHSnicndGvwV2BhZj
vVlRb726qyd2WjPyJg/HKpNuhPQQDpCfGGGF30BKMTRGiTCv/8vz9HItDp4a7qiV
aXux3kHcqZ/Ce+DD9+9+hozWrYTgrGDrJ3b42v31GAfIofrJeMP8N3dXdxBZy9F0
p+dQScaO/X3YTfY1JHdgS370zEm7SSsJ9Y1D0KweKijCMABOCGaDkU5X1gXXhSbl
FHjwiNgTHZZLolZa9/igmxX8LMH0te3K24JyP/9jCzXKdBygX52k9uxZDbOmeZDf
OlVcnAb6Tr1sJxPQREE6TGlWsHMrgisBwLzYyOXZN2HXKRxIekPjjIIYNAYpq+TT
VJUHex2wp7G8wmI6kf9hUxHIUQCXwgpOOCd8ys2Lhr4jYK9Oe+7e5IVxYcL8yxSq
YVoD5RbdWcMYrT4s+TN+76ZOo/7jo3T/8PSpfoa5ruGH3Rf3axqPfaWmZkVkhSOY
meEgL30AUj6FOoxbt5i+AiUfNXFIs+rlbD+rVL/2ShOt4NVoNAXVYQSH3sWEoa4z
eDLE1ZwhtO7FjvLtdhkOfA6ZTeVM5+c2kjr9WV11pAnpIYZB2dvUv3sF+jDDEYq/
xYG+ct2duqsg6xFT+o5BZiBE/HakzTXX/yWnBRtE3D0duEAPxi+alFs9Hi7ObJDr
S7I3UaiMxhz+yoHV6ocLW4bqNcVjgfOGjMQJn4qrAXhnZjsTAW2w1GXxbUPw8G+j
2QGBLa/dceZri+LE9y62nKIZf6ZbybWR3PqB4EUouVJMEo4guqgHy///34GOSknk
1sa3CHaouXlQYoONUzIhqtfWD1M4VCGDbCSiVG1vqeScqSBzc2BeRBpJ32pGcfVx
WdOfUjX941PPcd+OglbrzqIfsFfbfeYyOfVGo/vxinjuLl+TbuGp6z+PqRLwM7N1
IUwftZjtngtxDF4AqnPQhwCri1j8VZZUW5k0ZvDCk/lJHEs5GRTv41P7e5PHG/C2
wu+DvY4e9ueBI2uTPOdDUOC7jAN/po7e3/Y6a2Wn7qw/IVY9gRDrflJbcu50dWv4
FQaAPt/FnJb4OLhxKDYwVw6tUvvO6TgaDYeeYAhbkteML+Fnrz/wh4pDa2RYgfRw
KBGIVjho15GEh24ya+laBG8AMVl1xIZMM0WVbAslsXqXZw8EV8PuTlsE1YXmWPC7
OnijP6H+mcvbQi4uPItA/NCptUMMFWpVJN6g86kmR+1CKAKYCokMmNeuDdnFROL9
mecpaSATCw8iXiiTDYgZIcgGxW+ONB1Y80D1PwRb6On7X78YlQjEl8ArA4dmBTi/
Ha26TNV+6m8Ez1Q5eIn3cx9KhzYSGz/rEAwYiWr9jlbD7qvtpC8d6Wfqa77cwDTm
p+4WMJ4pGXq96sWBI/wK/oOOVQxHZSyWHemIAS0PWp0Kb6R+nTST2h/V6BgxhPi6
5Cim27Za19STa84zP1+ipcb+9AD4dh+3cpWEWEW+UDijYT+DGW7FZscOZgLHFtvJ
nnW/n7j8YgZguucG3LsEZLxPYpZxOdpMBR3HpvhhUASRcdD5G1pxYxZ6KN77eTB6
PglfrUxCeQVfLdY6F2AX9Jy+RMe5OqIu8fc9PpoeJa3m4DTUn56Nv0ywSgNp+plP
x1ALRdFTN+amFYA/uWaIzWM3BWPi1zRZrJ+JfNHz/1ZWCoDPy47hNbMteTudEw4r
ncAJasMZNjJpkB8vEESlUsIKrcTKNUL6EeDiSmhVtxwHXMFKwBcBJvCHEHJR1YDT
v3i2s2rx5WywCeLsIGIQk8AAEP1vXteD2T/3cRIM+ZthrWTyLyoqlHJzLGNHD2Nr
yyRbjC7cj/CB3bTYTkqUbpEOE7ZLW+uIKr21uUhEjvzj7T0C1K+L1E5avSkAAuBH
FGsgwoVtJZWrkKRiZCUs5J+ZRrYOlBvtBI80s2a4sB9AQObP02T9ooq3WxV3VVXj
VaHkosBuAkngHLGiYNyYzplcnqHN36OTDNGZHBpOMVCB2zYv1p3riyrDBvgyeKHt
PUGsMcm8eIy079IDlXEhgGigXrGChShkr/9rlZ7N8qBQC9E5sc+Lfbszl69VQK0I
Yp0BPgwTcWkg6SO2vmf5HfnwQZMowmHxwtJHOVnSJ0Jqkr///xQ5J3BxOw7ESC7N
XkQZjooK06YT8CNpeTtnihCzO1saAwUaSy7YxoXemcMpe3LZ7huIoKKSuWRMwmvx
qx1RDv83u61rP3utR3QYyFbrZfzgm2J4mlS4zOHh5120eXb+gIWyJPrmLESRLJEq
DlVgC7qq5nqQxZ73r2EqUCFPgExCZ0TaQjdwnLRvk0RemBLZ61e7BpO36vVI64bM
/x3lW6B1fCSy8BdaJpd8XK3s+UqSFBapn6spuwISxyMlXjYGEgxkv2lP62iRK/qe
5eU3K0bAZUmzJkVyxS4DCXMxmX8029ztcoLUcMVX1j8hslXd1BfHCi6KeMHeKscP
IjSsH65m5IRCAYvnC3sT4sUP0Sl2pxrqqazENYoySzl98Wlh2fNMZ5YQuXRMwEyF
anbc2EAkYhCZWX2zSj+Z4hdQAvhpBcZAAeTz3FVDDt4cBIwL+dGKjtVD3/u/MOKs
Tfk7/5+K+3XR/wMSH6gwWVuAUJwWGJrTmWMqi7/2AdFIaQYmyAlwQK6U2B844rVM
W83dn8AAVz/CLLRoGxnqbAV+wcf3s4z0yBmMhHLUuE2mXUDiMRoXoXO+vMO4EuFh
jZNcgzMCeZsUj2uYZtqeQWe7NhTrhRdE1SGK33Tp5Cc4IYDsYaY0tYT0+EY3lhFP
iWf3v1sEZutGj8pj/7wFiauJ15NDIG6OwWqqDLjeWm9ww2rUCTrigGQfjCq5qIoG
Mf88hl2godoL2D0Mtu4OUOPsTS0qRORCcy8NvK+yEB2MjV6NObtQCf4C72RQ38fv
1jl1adOo0mHkq8pz0BXHAEO2LbidgHJDC95fYX88BJU8WTdi5v21HltOV9gtr3EB
BsxJHJfgWDTSu7s6xHJR+8vgQApjtkBSoNzjF9cM/bo6UYrwufnavTisL80qx/vX
TKidgoxn5DuwI9/e77A8qGNIYRkTLFouYQhuCqhaY+NpTmaY4F7Es+A5IRoze/2Z
KmaIElT2TAvfRLJQ+ynG7PtATFKtOATyMBu/GVTXa1NQY1/rDV5BXXDk1nr0v6q5
pp+BpEIbAzU5qVbfwTdN1Xr7ncZslTUebhpHe6zi8MziLc3ncUbvkLDT0zvZ3aKk
6BFPxTRfvGSOZUIHD8W0bb+pkPYrVUxTAqHlIvMl1ouUFXj7r9Vk/UxxAYThdgZg
db9qF7DsvfpbFsEJ2ZgskyQLtnHLWzHwNkr30URStkilnyFZDEfPUihBz1cQsCot
Ds2BZ1YSwle+dOA25/ipbuZ3oYXu5fUEdZOrV/2AHdATFXct8sN9MAreuMIwAlN1
AIoDBqSbcU0ZF1wFhh3oBUPhzb0SWItQ8OY8wFjPLURCRgenJI1A0AypbqdYe/GG
ciNZDT4H3VNuSFbQyDltD68wQXN+la2li9rhZwId2UmcfKzZ55faBDOSdoU8IzkJ
NrETwV/xTDQWphTkbslkb583H49RhHSKZ4MMhIJYW3QJth8JOHQwgoEjIFDrBOFB
0T7vIEShZY4YkybMVltTLqSHAivzemnzyELFH8VuQglyxtoJMo39LafaM8sXlg7C
v0R4+JxL9ZcWTpHQ5gVOmn7FJeF+yvJsgVElXLP/MQr5kiGz7ZADrDtcfd4e9th9
R+pDDezwTRS8PKD8hdFVklq8GnfNnJ5QV+MclQyVXUS9DClG7PQBlwFLiSMem0Gm
MeROvivNdsE5sK9mDoyuew7VahZvGq+L8bsR5vesUXWGh2ePhVPEViCthh5pokSs
AbaeZ3wfUOlgZmKlO4cj9Q/64FN6ckxWESD0xBRCX5YEJJxqYiJHCmAPWnX1hyD9
7yiFZm8FqywfkT9shH5Ja2x2skCqznD9+ECagjOx2ixD7qi5BKMpBxrcl9O6YnL1
8ZjR/sCnJwqCYfclBNefGCSI0UuN1X0x2wx+k5e4K9ypYB8UmttqjjIDu82X/WUe
qQ8jOJyC7lil7W4djAhuWI7Q2TcTS0Qwn4J3y03CQrsbo9vNEo2HZSBN43ABNppy
tSwYNQo6T9qnW0XIwYBVSWIk/USLWCmwyOE9bK5LjLgU5IxIotBQYWFb48UBTgpO
M+EdEm7BY1f2mdOXBDYqjKTn2s5ifgqPVflu8OJ+hldJhu8og8nXLrtdBzTiB46c
DjDw+medMYXpRPsf6WIs0X4j6RRTDM3ZE+BX3//iwYtS1lhVC8eKwXOE3TowWdZx
phGEQSmnNbkY4t963Uk56hFZpryr48b/8XfKVkuVzHSdZ5COm4LZvj+ptSPm9psr
VC0i0yeCNvBGsVdRyeAvolAVbSfi5ot4XDR2uR6vif6JwGgDVQHbHGf/q8LIMgkd
ckKeqHFWpY6DLVXKZSp1THlrm9kepgpSVfx/NkrQJfIpZtedAc4EGhOzVYfsKP7M
f0cGN11zv7cLpy6Wh1mnVWgMWAZAmByyjsBwyjUC2OHRa8u2MiQvzVP41k2eHgQM
saoU+2k4whogBs8FGZUdthMG1dvH/0Nz0GVA1WZd1fpckFB1TkSHe0w3eacESGvH
1i6Nd9f74jSoS0sJJvLqCqRM/HYzNl2Ai86IxKrnxAA7aOIaOYUwF6Dw/PqDcqaW
7q1TBY9Aat+2cSDpUcQbbO92GFEpkolr3d2dnIThD1YfPctznNDLmwwP5dME8krt
HtqqbHUo9R7N47FYgA8hx8SNB0wIUHTW5UOyZ2AsJjYaKvZvU13cY24YhpISWgdt
1R454LHbR3PZh4eqcXTrF6ZLDCIhPW8yYxVblt8aby8phU1vSq+nEOc4ENTd+Hft
MnuIgLKpXu3ufSIVY35lXF4Dq8KWr7IexybCVxBlceZZhYPYEfcYPig1nWOwa1MQ
Salw7N5PHIfGIjtGCWRGcCFjcfrFc54c33k3XGKBDkLrghyjC1J10dwvirHK/6jK
6Zt/Ce961IF2QgXbQofvPU8QhxxBLaaGfiln6gcVKYKXOsxuVcJjZ0sSI4ShyF00
uGfTF16h9dYFmqA+mFlKch1xV42ZxdWm1q4k3iRYlXZNzk86kMBvojcP9M4/7+NO
8r+rbwXNw+1wbrZfiSylwbZF0Xnw3GowKGroBjAyBV4643jm0oZy7QGtoMCi34W1
KNOLz1uWvz1yO+GW6iWDWpe5qynXouLh3tBjZ0RNinadrBXgxvVb3c0I29ciqFk7
u/l4/1NBXQifQYLpwQWasm0gW7MZ3MaFYIN3OF7npt5kT5b9az2Ljo394ZhqoxAL
F1uqqy4OZKsqZIkPZf+0PV5SVQjfW8/eDAq8Q3JssFn4pjtp5IgLE5gYlOhloEzC
a9xPnT+56e4USWi/AwAY355397Aa0oy3NzR+O4Ig8zHicJyl5E2p6NnbUEjcneVn
O6/5PAaFlzOe3fc7O4LMT5GcxUzW04PGfZFfvS1OmhKXF5F43q4mhkrQDgURQonY
drvNZp5cNizCQd/nVfozT8nACJugFnVQZxDhThXra5I8F0wTk0q7ZtN6g6HF8HAK
rjxhJwfSstfPuJQvHJofABGDohMxHYEKNA4QRDxxMTq9WRxxNQy/qmtJIl+tN1py
Jvy/HSjl1k/PUhaJStEkuldx9IslFOecx2iS3VWLUliXhpVTZNwr8GWKw1Fdc+ha
bxb2CgtnKVYK/BvKTxDHCwc/9QKbsoe52a3BJMrrvDVZLhQK66lkzqgoEBSryT5s
jC86hPkNB3H3jyarrkk9YVmOCTQl27X4tksYthz3a14Ir+5vMMQOAmtxNG0tQSPA
BqKKbeAaI7ZHI7fGZvv5v+3LuLoAI0JdgU+gE8PhP+wZj8aExDFiTk8JNxXoX0QN
9g9gerHVAqVQGdYCjKe7vvQZsaqmh15Fnw+nW3q2WNswVGO522YkKEdDy2DTNzBM
dknD+AXCl5xN2hRWPa0lAARKbwMxwPFJ69uP13D5CBNQ87op+oKpMxlvGdavEIqA
xiaIJXecoZPRANCvgTZYaZwFw1lOotvYiK+D9mWIRy3euoOqDXAn7bHqGIVTo4Cp
u3+jTCJUs5jdbyEuzWNWyb4+gwuEytiUVxTrzyvZTGOMwIyDZiKmu9Zs+tSZe8eh
KYxILBYvhTDyGaYoXbwkfTosc0C1q4eHMDp+THw16kSwNMbsQMmVrggYhk07enqe
IlrLVIAeAGzgSqTNke/O5W50qb3w/tXxc1ChNtB6khi1FHPHHE4HyhrdKdSaMUnP
H5vGFRMV6OJ7ou/ot/ZMX9caJ+0WF6Ot8TpHlcV+z8CTn0d1iSMnPI4WJvSgsEB3
NIcD8CtHaxHKfFxCJGz29f7m5/y0SpVM/cnp9Yh3ehxfOwva3POsJWBf9xXM+J9o
y0rr0ydz+ppXyWT+IGN4T8q7xZvdNfBr1JV4JMLSRzZg81qQPHrLNkea4Hk8lWqI
ozEmeEcek0c+TGX62mOG2FVbGrI0Q0jGd0+Zrjmshe/vTQJqclfBpAUPL1e3JzeS
13NExBixD6rgwQ6inf6XdDKCHS/ENGwk+Zfqax8NTdAKTWChUSR5cOWeZCmVayRs
YUGV8BMtXdBYxpmPsITp438cswAE4E2W+kWM/nQLVKE4UxmVW/78hN+SGP0q9gMO
iRjiBL8cx+Y9UcnM/QERdPUZETDSnuSV3mXUshUBi7i9iNBuQU1MwIXwGLqI7bJI
zTp88r6gNzq0HfSCZxEQkyRu6Puok4tyLZFq9AMaYd8clsJTNM9JCLTvBSBpPmQN
V61r7pn8O+p9KdPmEXlDNCMh0MMZexbdt/Wa7E1NwpGXUkPq0u7YEeZEcLv6cdcp
qijNJ0kyZUeh+4aC+dkmaCpWjv/smseOf9KlwiZCSJRxYPZmVO0LHOH4PWshQhU2
07Mbr9pKtu9MizQyD4juR407wWqYvvIyuL+jg/mUq5LTVunlVe1GVp2z0Ox2Pww5
B0A/QzfYtKOy7beAbrfmOASAIBGainfUmm98P2eMScKE7Hgv8GY+5HC5+0KFi69G
NwayVOJV7dinQTmNwTwT1TFDSRvzaURP9HXyoTMstovH9146T2XPKis6tkjtZRnt
os+5mh0nmclG0Aa9/OV1l99KfRzr1Z3eFT5apPCwsFgqt//GqYIZJZrhoG4vpxeP
RGv7VyawgBy63mhQxS3AAScg+nzTPrVdLmdY0GFyDzIiLx3GPkyxQ/zY790vsrwD
33lJBQOM1G8SUqLkfVW788H7S0dJIqC8qFDxP9AqHOc3PDv5ETTfq0O9EvpAFzXu
q9av9GMuRRiatypL5z341zKBgEZX+RREdJCDTtklhz+Ww0d9p9ft7GqJeut4/n4+
PMHQn7ObQbwynCgZJ0bVd5QVoyI7tZruPyExUD/Y8qJDV0obOEYIZztYFavrPPsR
yRS6rbwBdTaHFQPtj+6p2WWhXru6HwJInbxD04x9i9WeAfzL8TRJGO1JaD61yhGR
ThARoc8xdoB5mGlwacbtPqWpbaYyETSujWKw960XP4Z1AE9oDjmN7m8v7ev+N+f1
zPyQUjK5zNikxtWifwokxNrTb1Amhtf6tGPswJ2CipHb/rDLZ3TVayulgarAkqDI
XNxEVN1RYRtJ8mv8GMPCY37R6o7P2kVCz8d/favfpGG88+rwf+NXeP+/gdbOS+/W
5QvdFG9FIB0+rqs8fD7d9IpqEKXAe6ncB37AY/Xc4XPxjPl/W8FQAsSeaUNQCkVS
l0VjPDuAikaMqKrFMOWVr/i0TYuKt0i73v2YBLg6KGKaKmCJKT9PTn+WoQdiGASI
Fq7LY3FNpScuR+UdLIoYM02gNXRUlTJf3NGLPpbRPGZX5+Ss+RuJf1WZ0+a4Aw0g
/L/8XCi/+vG2AMSCHpc4WII1HbQ7DyymxykYryPLmE7ta7URt54HJYDLfCcWa82i
LxHAHMtguHFWklzbq/p9A3ouf46GAXBDWPUh8ri02yGAWc0HQROdE54yvzrzSlMN
fcXYEE4ONyi0ek4aNZmdUjAt+Xyf74YoFgrq3pJvumd6kr1xlya2gH9Ye11tIVVG
wXANNXHf5ojo+8Trl73f7gCvdZUyjcLp9KVImPLMnMeXw0JLARjAX9NFkaddVBD2
FyKWT0FR2xiKQt0sfU/0CQBFfEvx6gI8dW63MaplVMWuEzYUElCz/k1mDo25QzB6
SHteMqvxMlQ+iy9lWLILqYHTLKNGaFWJfh81a5gUJ8LjkmHdGPijVecr7NHmdCCQ
H6ScP6pFJX5G1L34oOYybQ5q0+4ENEiMZOx8KnX7Q4dU0351a6quLCKC4NGrbh82
Hva5wJbtjZ6rz16ObPlgXP4TrvrpaFKd7xcjIIIAmBRiuMDcOtsn1vAyflHKaeT9
/Zk1qJW+wvMT7Zk8VRCNj3lBKRXXDz/kypevZAwQAT3wQi9s6G5QAJGz6SOyFfl0
oeIxlqA4Bpa/UqA3eijRS8LN7q2GPISZw/84xJfywX/6f9cKlpdnF72t4bCCCamd
Y4fBrWERJdYL3iOGFpVAYtAh6tx03lq5n/7eggiEH8x9ScRySGuqOUeDT440P7Ay
8BRqXlj126YhXFSXMlxltIlol/t/PbfqqNjbGXGe5ydGT/ns8Ztmx6B125/XjWYj
Es9c7ZnltKQ70Nuhvce4+A8pdP3naolR+mZKCaPxlDOOE+cCydDyrkYZwFH99MhT
aef3bsFLVER19FQPibJTno/1QjzR8UG6hC14GSSWLP57n2LPcga5l/8DoFLi6T36
N3XS1a76NU8jHB3ceV1kPwJreD0DMwWiKFl2N9WUcw30FTLFHosP9cZV/CdeQ1oQ
sSgH/u0zfV3wSZwgM1qbbrVlNxn9yHeiwKSPbnf4+lJcETVE0RfseuBjidvj1Ncb
em67mH6+jUJs5xaEYqeO2ORSIS+VoKNBUHzGX5klPf2baBDrKKsoJUYAUKCaaMUh
mycIZiK7crXOxkAaluXrqeKrXb7bXjkG8x4V879RDruvoy88ehUb+jy86DAx1nIM
ixqtn9/S24lOcqehGQ4E7PRJT+c0qX6zqUE+vGWeXsNX/T8OdSfDP2mPkIJU4xru
EU+pKdxFgTVYaZKzjxwesi4GxPcbPE70HuzeEwSAq9EWK9NM6NTBVLZBf5hqFTS6
09QAoUN5tobLxbYAGJk62JS0cBBBA1w+dHt4yF0TnmpCActK8W1gWcPAP503bpzP
a3oiWiIqu0hNUH7OE9bFOZD/SbZDEoZCqxCoqAnJ0VyVxLkUoJo4e/eo1Uq0W4Gr
MXM3YIF5SkxIeoTpWA/5twKnnnukZdDpT6dAbWh4Yqq8VA5R9Mn4IAPDR97riYwx
go+ndnOx5AUenB947KZfr/88aqXSMBupaSaKgWQTILjyutUFPF8mglWDkANUTpaw
EJMvTUP2T+S1g5whBYBBy8Z5ZqW3oqy7F7+1RpoW4+ueyRFc+LZeG/D4ehC2skfj
tNvHKCzBDW8xOQt/dGkyt1OW2jZw01D5qD7ZP98SnY9VBRbr2Go97L4/VV6Sopjr
nVoy1LEgLV2CR3Hpjrj/NZ/LzJ5fV47J7lvc10f+x6enewLDapkJIa7Az3SSgGzJ
1sg0Q+SpjOlMkG8Gi6+bieUXcMiIlDiHJXo7YQj4JT1/yJd/ssTf6vpV/NfmbHDp
Tk1nklmowWVhU8mDQJkxuV/LyHVA+IULZn0ToAnF+PscUysQG4X4bMmSo1GLZeOX
jF7LkvwGfFtxIsE36rkHHftKSjV/DQWkRxdKgxZ23yzLGJWf9hlzl4NwwQuyMU9M
SVKMOQK9cGoTuI2zFRTy4cNjPvr0wntI1o8mM9fv8elbDm6gPdquZT3sQlCm7B/0
ADJihY4ZU7eEOzzR2woA6EUZ9py+ApkgN9oTePfOiL62ZkJW1o/4lvS7jh+TWiKh
CRbMWpKlm6uUXAIni3A3fAcYMzR/GRJq90ms+nBMSPehzowx+5TqkBltrdkg1RQ5
uu6J3cm/CcWDDbaeXGAhjpJDJt2rRl58UvU+gtswYYJoJI4VYGSKRgpr/p3NpnaS
UZHpqfS5A0T9VFZSfzbUY3vzHIJ8J8LCmj3rFvUv7dnbstcGGjJFuMSIqLARmEO6
CwmwxRtU0DehNjn9VFNn2JQOZFMSHXgor4YTiPIZ2ljDgQ0Wr8sOX2WqezGTf7X2
u44Lwj6lEK/JXSwIGou9rsLaaDlV1WHQce43DzqK7v9kIfdO7v+I56Dcwjkscc1G
8rsUHu8c9+RI6ozRcTYKBGPmJc5vwc3pzRwRxYnV/IyN6kqiKoyJ/NziqxhKCJfh
olcjooQK5xAp7ynKxljctpjqCZ7PiFbRnLR9s1maK1cawba4oMC0twyjeck3NrJW
0ceXRcKIqkJl8F2gJ/NOXFsvImu7vEppte7yFguAv+3CMbx/46Lf5GUBrDiP80k1
1WYy09UO/n8kWSWPuZflv3hUcbm7PMeCyFAIa4IBN8Tjbi2cCKrV3j++xNi/iL2q
4RWi6FSGTnzNX7mGL07hOkZt9ogNH44qjvtJd5E4rQ3TWxkaqW/KQGb8Lgr4vrqM
+3fhGb3truyBYny+LtOniPueDs13uxGcwuqUozAXyYPLD0HMwdHLj4n1JAmmR5gF
s7OkYk1TyybjqT9ahMwO4jKXjRTnlsgY9BSu110LfZ8felT2CZ8S1gpwcApaDfQm
9m6cBq74s6j6p0twVXiBTsP6tIJ/LSxp3E6Eg0UxDjqLiYskMvcS0d0Ebdjj9fgh
nbvf200BYYDxK/OPgELrBu7f4zmEU+pIGWhDDGCFBvl5OWdTXtxmJg+4DKpskQrr
8u5ummZM0xyWVPuR3P64hMh2XRBIajLB3c0fUpl2UFXpvgo0B0AZJafieoWynP+i
N0IJyDhZVuD1Lrv9q0/expNVdLT5LUXiWyMp09/m/uyPCCGEueP8PPNJi6V73xGs
Hjhqp/a+szTT1ZaJHaqv0RF/pUp0YWTRTlvzhwLRjSCIjbaZSfmkfJ8zNeD2CjKz
fGOndu706mu2kvxeTm+L3FcSyDOKIEjmtazqFaUqmUzEgtGd+5IF1vrRMD7HXtOC
IDEyElZfnVPXb/Rhf3g8aohJIpMsrqr5FE0G/SS7skM7Scm3wAiloSF1WwYl8ay+
yLq5h5NXowmNRpEPMlMsvHimm5oPLwtbeq6dkoICL3a89lvkwtjAsjK80azp21ht
h4z5x2ZgGp9oEtovEMubPS8mcOojOu4Et9wL9/exauNng9x91JRCnGMW07kd0DiT
cQxBz/mVaJ8tmD4uOMIMjb+SekjURxSqK29be0pbRDygFS7SA9br8LMPq6D79ev5
0C08NHQhoZ93HZMlZEXEBhqvB0jsd4TjHDG4983OyuhXp3B8m5KpXzoxF++j9lnz
0bMGN4ax6gnURpaVrJgWXiTHR8iExq6UuXTjhCN7EXhMvqPvhv9IDXGTz634rd05
6lVctE+Z0OqLaM2+pwjFR9Ps8i0jwDVme5bMa+prunLxlJSwSa+sQoqX0dzwE4Ta
3aMySdcBA/l5tOskG8yHCqiiISGiUrfgO06BsaY+otibHSTNOwCeldkGQwtmvPb/
8by6CZGvAYuSNVh4/rycD1a91ZhRY12xbQwauXXC0U6JFKTtWrj3fKWIktmOxOaC
7dWTKKhVPjOdKFRH3rHTXUbpa9YhSs59UKZBMt9QYqaioNFHPNmq+/bD0/NeQSg+
8/DDPygkVpllQuZyL9MMjE7OiyuA/IScwQXi6TGkGWSvunZkDzzViaLLu1Z29GCz
vU8DCaRwY1+cQMP5rUvqCZMlfD9x/xHYo83tghyYCAM0zBTb7sCVRLUaDiYHpGQR
hJ15MkDiYQ1U1IOA9el0Djk2gl6rRLREdV2d2a9FBfVJmh2EnCgQRmFLp0OQcacp
U8z7ynOnQqb56jfuAw+O3AlEI96fZAUZ4tL/XwKzpyc2PjSLRnqNgyRYZV9fJ/QX
RpX5rEK4wf2IbsdICQUkG72nbReZQEkH7vfCpccq8rx0B7oqx/a5hO9SD9Iup1xE
k/ltZ3d2LepuwOU9pVWPKhfkCPKu8dYL6TDK2ff36eCdrBw4kNXP08MQmJ9KBS05
Zj/MErid/8+vp8f7PnUq67WRPY1PUoYVUcV+kA5KV7xWXfFVoCi1LPZKOWa9LlOG
577+F4LH/IRPgvPtdVU2raC77C55m/ad1vkUIBgxuIYVGG9eU6susxx1dLj6d2H/
iNDDa6iXEW8kSR9ekKTZWg7QQs3qpSC/EHDoU5EhFOlxmbw/JBXxtHKryuO0yJkh
4xFWPG2spGkfVjdjlp5AXi0+2nKRRbOc/hyGVbtHtDIkpI8nsuCAezgJU5KV02gK
0na70NBBvc7//TwksTwJcgwnfSWsTwyLCvnPYAn0PqDahTL+i+Luo1u8gWAhOb3e
oisTOMqvAmupXeEL8jJfY9FHVJ67XQn62ibVmrrjEeOSMfoPB2vQ8mxbUoYbLL1e
tw2rExcy7S3USDXm4ZqDNzk3vtTMATtwCMKnrk3WmRUTUu5BHVV1EEbPk+NnMW36
CwVYzWKWgdtXa2t6hQ15orS+2LVJC3EbrfjnnpF8UoM4rLfmlZLSx6e7o4zceQVb
BM8gw3hC+jDL5T6yvboC6L0gDOP2CEniV4R+NiuuLDzVJQCeFojCtB4jeZojGsNn
V5Zk42gnfTRIsykod/jlcs5vprPdz05iUVeOrr1HhxYwOfO253aEH/vselh623LP
1nRlaED4b0AV20Koj9PixvCWgsrIkdQVLHBiLlzMiYAcy7VD4pfYF4F9JVaCWTne
x46mI8HLy4lj/eAbrNcTXVowgeQS6LSAr/D/A5A00CA6t64XRVuuzZedc3VRhqPY
jlK2HspCdnBrju6CV7mkeu6iRwfxvlqypAPO1006dS16VVebv00YrV6T70SvJzE9
kd7zuCrzEvZzN0tNm0VX3h+UBQTBSirtmrqIQezxGjcZg0Y+CZIpAqwYDx9sidUk
4p0hSVMbBlfzhbBuSTiBgZkMdOazwKY04vbUpi0kgBnRDHZH+dPZhs0uiUVmUzcK
nbWkV2bFGh5rGQnOc9Bv0DzXQkZ4Nyaex2OBuKqlXoDYm4t8dFqpjkhT3NbKMCwI
MXcWxDv65E7DWUNC7nr/3VpiNwiUgoHgA9By/5EbadRYAjR7d8JubnV6MgLoqDxO
38K4iapow1cA1jK99jLpGQF+jFSaaNgYkgsT7F88wmGjAndah7RjrFLUY+OUwzlJ
NwUJZLhBXJZJIR2nINbz8ThLN6eUQ9TGInx8LRgNx0GCsFTnzPFSrYhuPVMMYVog
ymUpv7T4sooyJus6G2Rm3GTo/Scf7YzRR6Sm2l/klBNuy/eBOgYAKr4TTeq4aTNh
Q7cZ0HaWv8HvHQwJcv+EdIhjJZ5um+FMEtPNIIZmSt3SryzrdSODyLzifQ3IfRkk
tvlN6WfPzri5E3FKKR21Zb9TrToTMSOkqHLq3exXrpCU6Z6JhV0UuRC7ZLRqFpML
MAr4y49YPcesTEBzxzpRFbKJKjpesMEtF3PWIXwmFbPNSUUVxrSIwepq8Ao/T0oy
2Wq+in3TEst3suQCeEBuDR0I1XXfIe+KQvRevb/tIoaU/gIg0r6NTtXdxpXga/rm
9ownz1I1z4U2D5fiupOtMZ+PSdWEiwRtgznlWvCVbGBQyd24pITPENdizO/bOkCF
juJ/ZeERYove36tYtERdKi2bmf22stcaeBax9hnJLNuFiDaeOGtyBT8nDAfBR0wL
7Kwbi+64naARzvuXHSVl+Q4WTnKFQ+qxbj4W7O3YVt6b3E3zvhrXDtSxij5AMsps
owpLvqpQ3P7jmVFYhrqDY3ZmmKOmwVnY4na8Ue/9a++C8p/gZEtV6+YvSCwfEaPh
R+c1oeZjqBzsr+6xU1xvG1e8aM+OWtFPEZeVDZMVASbJ5MDcPPzJBtD/N0k8j/02
40R7lB/tZ8lgbZaBHd2V4bJnaD8ycA/pA1uwFSKMiJ/7sfFo4d8H9OFcJ6h4N+8B
FABl7ovIC5uWHyBDrk3d7/UZgZhMCITZJUlblfB1YKnvbnCBukMo9yo1bkG9LAEo
i+AGE2xyr6SxowqN42ASrB4r+tAWtp5KsTqpJADRhWq/gNMOJMxO5TRV2f6+RVku
QXWC8aKX+vWrR/0nn0zB7ngQSWYrmQXvm4OFVWphjnoMXsMlCsl2cbOAGs/2CrsQ
fPEfpQpClhHanc+Kdvy47R4kikc7JZNbnIyS970rtIqByO3i2ch/v60+8QhyfsZJ
/BhoFZbDo1FAeUZakB0bqoiprgCVABRmUXTBgZ5e2ZWY5Lqd0yJShMPuymJyvmJk
uZUEqLj/alySMi3tHLBI6GKVcU0T4du4X0dITcl+fowl/1rQVYvx6bsvpuOc72Nw
SgKOi+lfLJWbp98oyHWlJjw1UhLBEJ+Vi6b47gvxaXlQdGm1IpWSEi0M+Fi0kD+w
fqF0dRdUGvESkiuLCZHy6HgpMGqx7/wUIhpuV/rdUVRkx/nKTHFvWMAvPJEjE46r
I42QPJA2Xk41HPQNi4F3wThbzCIeG3GAdISZFfLlfQeUGRISBrAH+3fF+3/dBI+T
JJvzgFSqYK+r/rPwYH4cCE2uzFlc4K9Uy9TQPFEHznx5ys7wfmsVH6QaAPgHUuVx
yNuu6VJ+6QeXfD55a3b/Ozv8z4Cu18ccSRrzj32ezwzCeaU88kLGxGG3Ky7+CbcM
l1RLTfm8kYsxbVeuebQiQ9gMgPuG3Azc2hvf96IH7hlHFVgXfuxh4WZZyaJwgvsm
Jd6awp4M6BGGfpGPPAHQWvfGwd4QB5J/BrgkOCVdoI79xeKEtglb23KKRAgHrvsx
l7UrxnL1UEm4+MtUZxNSWTihaMvaCjZas463w3VnPkgPOTAp2S+e+H0tQnk2nCSN
mu72EdTZw/EZwfmjkl0tLCiXJlpUooR0AhuzVcBmaDbiX0KbMLm6ypu3bP9oxtY2
InFWZuDzw+zZvyIiNSRW4Cz1makak8cc4MOjIQhQb2Ci3SyzxT7NbWdTk0WbJpnS
6Eu4gx2U8lVWNHYIGxuo4kq6nu04O3V05qNoF4kodF17/dSzefsdtWrlAj2EqkLI
pRp/uHqpmiZPx3yny687SpDbj8jvZUQ7tTO2DY75DmPiN8J4Vxa3GWSGvDuJLiOS
hndXlvzk9Hwa8GAeT2faOuEaWZujEEgQijOnRtskN7Wasu53lE+ChajM5KxYjksl
UuR/k/06qdRCgtFsNgzsP2I9EeM4LkqUdx8bFrWVfsTVUE3AqC8zPeIR85yW+aAc
Zfw8oMEbdAMYrTB46N8lqUOl1ywtgwz7YTHtNigvqvcjJQGCj1WZ/aRaqHGYQWuI
mBWpNt0u2x/CijUl4gSswUkUVfy71a9YkkWyD2atkG3QchE2eQGk6NR0X2DXAUYv
1uh6C+KRmMvMRlUrQswRDHuGZF4DT/y/+03oFzoLt/0Y6Fp3hjlPSHRShZ+zOhIz
igAksGo8EWxcLsC1dp1PXinJM4S3gKc+WZxwOlxmyPG/pmehp9ZiUbbszLTy6D2X
oiOQzSHlp+2oaLwe7LSUjgDNeKXbSxkw2Kkhj6mvhGjgp9/kXDrJFDDYZH8t3e3a
MJ+hGNCGQ4LBbUpIhemRXIuKNdW/UbJSr+21NbUZpqNLuBscNmLO0I2V6O0fAE2/
sA+wiWuyXzvVEiOXACV7GIeDMBQV6ynYPAKXFMzntFOFhqBadVvkGLiiiIRiD8Fp
7rc7mvs1guTxspuomM8BVEb+miV9ooTtKVnA8PR7W8WVJypJ2Ah8RX47pSl9DO80
GYKf1eY6PmOj3hePSVbmKQ/ot+rWhJNUw9kBzxPxWy9jx1J0dO1GJpycl0fgM5Sr
uGiLYOELkr16Hag0+TMjWXavaGvb6iaYq1FSKKxxPIc8xQ8CzoUJduf2lIx784Po
eN0Bmv2sTDROadjM7v1LYpCk4Imo7eaIy1JJOFZ0gva/Jo0qTX65hDG3OhPmyiU4
BI1ou408H/FrxcFA1olpIpxzGl9GLldE4x1XPhdFraRgOpZJT87hnMV1fRzCa/1e
1SfRUnFMTdxnhck2o2KI3AhPReuAZES2aGuGFTMBhzScG6e1DvqzQmmIJVw9HveN
LlSvza+LnsAfWMXhD3udqshBEZu7059QGOXkkDkJSoLfJiYz0LY6cpIw3YsE7bnN
3qAUrT10lCewps++Su276m2Zjvh6nQc2TEsYEo/aFqspo6piFfhS3L5rVYNfG2Eg
NGU2IuT0wDG2Nvel6/MlFk4Vvt7wn3eAsUm04+55ldts0pSupRPvEgGHxLtQ8SFS
omdSCeK5wzcA0YRCLiexxFBWb59N1X4E84w1fZtk+KlKUKj0QoB2hFUyD4ps6vm7
AMpCy2jcV6srf5vHvJEzHMjbgTWItD/sz3QrAblOj06gZghjB2Icbacninc04Dxx
52inGi/zGxCuv1xt+qu/sGEjAKFZ0bGEbuswvaKsxTRP7Zzh4G/ew+148pMT2tSL
4G93daBUlgOvYwwIm6szbLQJvOjmsWKdA0ZCXpeBNP88V1hTcCpAuQnD68ZpILbe
hfw4btMh/RL7oaAAOsmqTRnA7z5F/AFqSoPt2UFirKlnt8w8RcXh9EXFncA7orgl
lQrmq0QruYjj0D/voi0sgcoGwkvOq15ovoQpJYuSLHWl0jYT92EJrRaH0d2z25nd
NjRrbGDWPGNtoak/rhLb1DcdkHubcU9dgwl1BswIvbH68hL9ktwHHCfXZPNhCYNz
AOGR45WUOTWNF6NvKn7Wber1T8Jhb/hceX/wcVdEJMYJD9SUk9mEajMfh2u66vTD
9NwHd1/G83kIT+Mx/GyFGv+ZML5u5yz1trUYpaoOt9F3qos4dKijPb/Y9iGQ72H+
inUSitz0d8s7DR/wKWlZ3vGdKcLJcF1CyVCQFSdtHc6ceFAS+GmjnCfbhtQY/tSK
ShT9XR19WxgplU29hMIWznd0ryNEju8qAAQ1iJnGeAZ4C5mI3nZ4CWtZoO8eb5nr
ruQDua/NbFGD4jyVKqKTJrLBZqcleSK5D1+l3DfO+p+9mDpREVv5kyh9Y9FyfwXT
/5tB0YgKxZjQbUMSxxm+rGENQiA7iZxVTcn8fMa8odaW/mXSHfk+NI1ndEZgntbG
40IMIsOSiFE2ZVOTTJnPaJUMkdF3YrFSObF8rvQ1PILNnp/DJ3jrTRlllpJWNFeN
pUhMyl6tZLf1ycDG67fqqw2v8NCQs1B1lqfwb8jW/CR25+amW6xyvEyUHlQCdLOk
5c64HBjdxCUYDagiT5DUgNFqCHK1wevD8jgt8BOZ2W7j94xeHEz6MTKuQD+HvA9o
0Ygezt8bBf3U310SAjdtFdRFYPpEww4w30eZ/g6Loy/BhLcMxMA0ooov8e121Nd5
aws+9ao6Bt5iP+xxx1n5zYt3s5C9mlL1+JHLn3Pciu6zV9t0wKo7WS8o97K/tAof
pYjZU7dJ82DzcCa4r7X02xBP2CjPez1n4qmkXzOlxrdqPTHJzGlu2zY5KpWyl9O2
OenIP9QkoLBAKdPSLDfV/IeU2QHnL7QwbuajojKyUTZ1dVu/XhqZBxHrSDFnRAc9
gJeFNuyCUYepZl2d2zzeY9FDfeL4clMup9x+PZS+Z6+Bbb/HMEaWjsivH1kiwrVA
ezYQW5+7wEW9pkehhiXEH+fjWhNzZryGkWy0b3CWR+tUO3+q0FOiLUI3MlPREa1n
dbDRTxmxxkvhLRjZdTD70dRETSyeN9xeA+FN5cOHQgHEP7YGjGPY79KonCdRVQmV
qyk6YjQs+bSQJWil+EtFpA9xLRKSrzAKLfIvVM40rI0L/iSLq2TfjPl4yrb/NLt4
0r8g9FAwKfFX9MDx80uBHpxqOmHuKNN0kZCDexuC5xfaCDEtm6pS5YOFPcq8KgpV
49BCMyDJ/HSP6HEw7ZjcqBgoOQecKLYF1WM2Fhh6YAYrpYkrFUvnH+1NfPfgHwJk
EuUKtcIqkp2kUySRg+bj4RHUtlk0i8Fk+4iMAfSVlzxsAYnoFkp1Xo1UpDI0qzCG
V+54m4fM589DhhymBjs6v3TbGX/EAnav8I+1f4gaJkA+iC9tGiT63fgpg5hTPB/N
murUNcpaAit86kh2zM5dHV6OibBd7G2RcExeFuCjrc0ElsB8JwcL/FL4lgBa3lZ0
ie8LWkRK8CW/qn+aO0WJouRiHg/khSCxeBCuRiImIh0zm7EsTPU6DZSoZmuE9LXo
jZsbYk/FRPoBKP92fM29z1gsU9kTAAWOUEwWsKXfYdDwV1ISLU9KoWHt2sJ0ZERN
vLNeYWjzXp93WKfNe2gOzEIHBmeAn8LA2uH9JlPp2kK9prblAqasSYDvoFp64beD
iE2lZSDkG8AGJmUPpL53n9md7A2a7Z24ld/SP/CVcw+7b9WOLIMtxs5ckBNxIp51
X3R4gzmHh+UyMmw7gQa6DL4LxyMPRSy3q0QgJ++y9c0SdyBYktMWbVJTTlfUtPYa
OE6QZxN53ZLH7HbgvPr362NqDW1XqLeFHpPoZb15QTpNNT1nbbCUJC/8eD7vKJbZ
WJ0mAem37JXrj6o24qfEaC4TJ6SytNUGX8NLaaX00FlAbS8EASO3MzRoqub8Wfqn
J2dILg6rqGs8sriYoxVsGW8/ZrfvA0nMs4GUoCYIcGiwMkj2fK19XLiQJjr4fNdB
dk9rNd5EQpWBMFmkFsovaDV42gY41d+sAU/TdeSXZSdm/IPpSYy1vgbF9gxueB8u
4EaDmFTa1ncw3VRQyXdaWUsDqLUYZfELT0grTP7FLJF985WmE3VhisrV0c60DKZB
dPmgJRLFakJhlEOGf0LbzuzuEyhj3gDk8E4T804Jfp1glQ0Tg7vcvzjHyLYmgkk0
0c9zIJ2nXGiexsry2txsyFbwC4nFuc0hM8RQwbVrv3/MkqPn0wROUgG3I7nh9+Qv
7PFBvNt7zHt5zuqQpVnoWy6qD1Da1ETG0qDeSaCvB6jlMQWhxJ+oGRCHuzQg0H+P
Xd1Lg3s2HNmzkz0WYvfSi36uLz5UPSHzJ9obQB7P/AwabEpgwrN67Pwq00B68vUU
VFP+5Qt1wcEBbjEAc25Oun1wKqfb3KMyL4tRe8f2jL+3bj1/GeLQW9BaJooB9PSo
Bs1nKg8lh9f0AxozI9b/gj92Mswu8uPGd1tCAkjxhpsCLDmtoI9R9c/Hr3ddMBdi
Z5wXSUCB/hmv+ItVZ7QaMq//d9MWhfGyDEfpQ3mvk5Gs83tO9v5RYcZqBg+bS2gt
eCWoWlu9M8dkioa/iPpNiWXUVaayu/teCvMBPsy2cbW9dvkrU3l6W7IrDYPxo276
kITV1anvhLLlbOlEYx0hVIcQKCcmrHKrbiOVy30KwjkwCeNlRfiTDSf3B0+sOCMr
lxmFfyHmgKuQGuGJXtB1mSR8Qg9XK9UFEChSWx3z6eQssLVonRF3aCIv4s1zN10c
KPu0q0X+sGOrxNSPix4dvF/fAoVXqDE0CROS3WrxG+KGW0qh2M+v2q545fuTiorp
PtIDSGvDCN8yqBjQD4o6m/G+s1zyhUzMCDaoQg5dymk/wUe+ePihgeSilWBKvaYZ
gTuj81MSkZwstV9GbMh8MC4aUBKJYAIYNtebS7OTKxf0pV3XrPlbdnvUJI0nfFoR
OyYHmUeHQiJ+Wp+lyL/meXLrSSDsMrxeGeIPi0ldoKpr2aDT3qbuXzGgVv5g6VM4
0QW3TQRSL//9ibvML2gg2MGL1176zoCABn/xSgSwyEah0QJ5CNYP20kB9+Ixk6pK
9QVxtG4blYtIMXz7SqZeFRbA3JY790StS0Oy2g2igRFeyb+8LUGMGFt2KuJS3TpR
A2oPQ+CM5h3vzdMkNsX2RjK08u31gjzvaZgqzXmh+jhRoae81mLjrsv46PvMYnTq
BA0EeT+fTSzTjWCyWtMMMvSk2aTTi5yovNFEoZ8XNixo/aSM/tu47BQW6Yvpvc4i
/p9TYwF5/dR3oCQob4XbAIMKwzCrbCBoapnf3azddye5BBWVty0vdZ/JYO+jXXu+
mypzOb9yAAJ8uER5CCfBkGyNp8j9h9NTlTmnWEElbjljzXsBNw8WSJg+SJ59qf1I
JEDgNmFtyRxJEJCE3hr3B65Ow+DnuoZ+mGRKJhJAArGB1vhDtJQPpTHKzFKhkJPs
svMQTd0y5gMhI0QlNbcqmwCCfTce5x2XZAmwlCpmsEyYYSuv96OQaslw6dZmJ2jH
3v/oz13pm/732nOAOuUvvtG8DxRoEWJwZQwwTQmq6QR+hG9qWKo0GgnTZNvzLfn8
XLot7Ihl6ESpcFQO3e6uVoNqOQ1f68WTQTn1UwBcr7kcUeH6PrfO4TI2UB46o7XF
Ru/cqrtKjezL1uD607yuMDeSx1/Jki2o4yiYZTL7+GetA/XzufY10hu/PYehTcQn
j6glEOjfRTcjVggiEYomlD2kfUo7lD3YgQa/W0GlI/s9ehTY8pw+6SBtvW2KFF+F
J+eSQxLvp5mXWjPFGaUzK22bQa7+hsNaHXHp9bjty6mSjOYscScOONDbWzAjTDUr
5WlugyNCNuZiATtL0NGtrOpfr6yLt2PFW45W4Phc6HqfEIvR6azwPY5Hn8hAlh2w
FTFDkLa+ZBDxlFLhiYbhKv3WyNyFZvFpRE8hMcSpX177l5kk8TsE9Cy6Zy7xouq5
h9ItkVrlVYXldrk60jeeyDgVbPU4/RRapYz1wTh2GF4Lcwq7g0lGl/Lk+R+ToMYf
NYs9ordY7/uMhW87vlcBdGXjEE+I1f5tvFh0y13Mww3O09FErqDvUViZSgYlzPBt
w/TMfm1uzububuYEDtfoQ8kb6TbEbDhoI5krwrobu0BYJjoQNvyiwOJb4Ym+PWs7
Xc1IMq3A9Zc3mvkHc8IPqDGGnQxz4kg1u0n8S1/N3EMqOD3k+CSj5k0MQBQgHXBd
8Yb+NSCqmXwirwU4C2uSDmfGAz7RxtWeSXBmblp27RaBh4jHo8obv/RM0vCQCMR1
33XFytGGtOFUGnTHc83/pCnJCXN3eDtjRuXLUqH6XcwIi0EBI2CpCouPq1HA5C2d
A7MUmYJIp+wB3pLt1K5lt9WqmcUsHW8C3uNECilzj6Ajqcd2g4F5EQ+4rwEBpRoX
YduDRoNvKgHgPBxY0H5JMWkts/vTSsU/yBQcuGdCN7azW2vymnPNbzEKWi/eM2Pe
N/bqSKCSD9ttSpZxPNdgQSxwqMRxb7W4EwPXEut7FAS+xusJ8XDYXVtseG2aCdJI
aXZbx1Ja8rJTp/p+8QrdsGI6Uww1khpsT99yM4krp7l8WvTUn7PDFQDa8lN3/kb9
F53KL7bcqDd8Ngpd7PRsE7vewCE+m0EzTdh5OL3M+Gb1yJXRxeyfa0YH3A1j7B9M
5YQ4r5Y2HSO79M2LqhG83FOvRSBGTJXbyX2OyiuL46YdMGaYh+5bZBNJ1mKszV54
2WQZlKGrC9XJ5esNMMuedQ6DnzWGY+JtslGDTapi+GK/LiS258EwcGNCXr3fLZ5I
N+/avsAGgpufRxz/3fzl78xPRoy52dtRuYKgNmNF1cZqrNLzd7iu//humTnrq8sF
6jybkp/6jaq8h08G1U6pWwk06qNa1NdmB4hw5mowfpIX04rKc3cLtcy6p697dUEX
krfH38t2pi6TFodGHzavIbSTegAGv0tFJxd7mF3P0i1U0E75x7peS706zNfAk7c5
SVQdJv6K12rc0S4Qe0fWOUdrQhENd+glqKB2ig0BKZjvoIWrZxAmbTFY9ao5Ibw5
SJ3Y+PxE5jnpBjNL+x5XS5KeQG5QJrR4ql1zMgvJef3VkNUfQ/o3/GLYYKNG7T6p
1SMm9ESN/jcWjhKSJjKr8PJ5hbJqJw6cyjoHoQvi7xuibYZMUyOVxD06FI3s14rO
v/hWpFD8GzaoYgY55hLjb8bSmNvjqiMcvf1jLPnSI5U3YafmjsHiuEa4ND92OXE7
ZCUl0MVNZo3mWXCW0Gi9YOj+Mi1yb4SGn3ohyf54Z1H+/Kg0G0X3wzdLMbtoFn09
v/ZHSQKZmHtxIM7+uMwp/qv/+C2abLtdOCKYZdHuy0NpmIWSnutGFEHdyaVp4yd8
dB8/APMk9FbR2rnrlGITDRKiV0sZxietA1/WB5sBsKx4Q0MpxF0t0TW3IsFwlK9q
V1PuzwquxcdnBnVZfVJiqG7ZEEoX/1130cbCtwO2ZIK1ScZgLaZ7jQCWuSsu6ktW
CLveCL8BN4+YpsdOjZiJkgR+wozLaiD4Z0PFx39vTAvUF+5Vs/gdXfL6oXb8gFng
Xk5k6rYE5Soq+pmtQ6sKXtYPPMLPXwlo97evw1bu+NLLAeKJuKzUJyN3kVeMpYwt
YGO8cKl8iN/V/ak+AbeMpV4gSMr8ulI6thyFXkCtaHDV/NdpnUb1RNqJNIY0oUgz
qBQbmKWZXNHKOtgkeEiKieszmYRAXvbKcotnbN/IVKqB7pimf6yyyNAoNs1c5P+E
5nKV7d2WxDck46+keJOeAnlPij3Yv04EzK+WUnIe8LqBUl/rVRWIBYECOF4J0OJX
NmRknLE/mf2RU5ozthszjLVSDfzFSedYkev6IO/oQK/Ebfegwat3BhrCyiiZ0QX/
6zqbc9l95tWo1sPQTp8eCD+UX+Q7983jJom4rWehxMxCDWhH1jyfyz6Xx7/c91TR
DLD7upBj7E3jSG7Q7lm6Ds43lxuQiVn1P4KsHGsaEttRqehskwuL4ktaVsf5y8FK
v+0wi5kcmwQqV2MNs6FuuqQXUGxAwOgCdkqH1oYWm/wqESeaL0TOwQTykbpJvj51
DXa0OeSaEemx4slbmr7BHN2VPk9xLDsqSSIx7L7T73cSI3/Q2Zt0taeMCXHv8fNW
huSzZsy9bMuFEBhnZUMaUmBjDYvm9Q1NyaaEtI+3RYR49IY2jLr423vtvUL5qZxO
atCt///q78pBLWhSOgbP98wHJC8ZcvUz2H+uZkkWcR8BlJsBbDdbU/g8my4FQ7wi
YvdpBOgE2AlQAHvGW/U2Z6OCn9da76Lf1UvEn764M0F5Qs+rVGbfqntJIxaNhb3c
sRusxcnnxWIk5EUb5XP5w+rNq0he3UCKIsPFGJ8WHjYAJtXRflNeOZFNP/rcQBwR
dSCfFTmXyVWaNTsuMHwdeUFnahqIP43QEb73x6xRYJS2JbGB0ETpPtdLOswHyL4P
3mEoKwPbnwVMNQVuaP9aifPgtxOtmdI4K9ayRBFB5N5pJ0iFbWY2AvSORFBSrRz7
Y4/4TfLwuWsn8FyhQFLhTJCN+f5r0pXPWYuOMddttukgAEZc0zvFgRj3fgSJSLK+
JF1wYniO+dJMeL7pH7PtOWlwUzu/IFZTcFY3rzP96kzbahI/ul5r+MjgcgFo0NcH
zLC+2GiI2wMff+jg6lCyo/06g0QTdFOEFn4pdwipSjRXHqNx9Wy2KZEeIOjoF0WW
82RwYvkpfuHKAVsxzTH/qEkKTrFZiSNEQN81lAkHbkk4R2OeNOx5cYNxTikotCBs
EBbR+pZKi01r0HniaWPy4yAbZgFkd8TSrTRzRo+QXJkwKd+zzkDgmVSX+ozfScGA
5lj0bmDgypEnPGlZhsFsoVBdCE58EUvc6ZM5p7yug8m31e3hT4l9aE92RYejcaLf
aOhn1kyqoLE8bFYqPuc8c/OtBJrVjw1flXNtXtZPcAp/sTLZJHmHMu7pr5UwIqhU
Nf0bXkz+VFAWB0Is98Gwn8VUX896tH3q1xL13YsoaG5PCPLJBZFGSW/Eby7N32Yl
XKyXSrjvXwmZHQ9LReSrsOOVaK4CbJ6NACzM4RpucUuaCw51TPs7XD5xNFDpD6oS
0gQwN+nkIhzXCBa3MH/nDMBLX0k6R7QA2xvnbdZu0wD3PhkOMm1PFjuHAc8FXRN9
oTGyif3KFFLjH+IVwU4jiqYRjbTY0i/QPiHrzwaIlcm8GNIInEW0sSV36Ts0NsO3
9BiYuruILF8SJC+4eeRIgyaUSKHRihs1f7YLIppfMjBS8pPdXesrheBCGOCLqIdJ
OgKXqGghdNEttGJ8Okw/CTxWsKmv592C7/SQbaeTOtgfE995rhZ/FJGoZ49rjW1r
2MPqHEoigVAKC52qe9zcW8Y5MUwzjLmVcj+mhb+wY7puL6o5Y55ZSZP8SEGm5NVd
6Yadgz1MKcE/bQcBEvXuF2W7ei2sK+B4aSca8Ls9QIpzwWTVn9fmRUuJmECnH1d7
H2SE/HahKrvzDzxwNpZ4B5wm0xRi4ctBBp09J5qTRNrAl6+M0tA85e7S2CZQdi13
ko64uWWQBwRIWq0t1bMJhxpivRYZXTdI0ruaKwzVaa+uTG13JBDPpK2v3jz5lMwh
59zWUTjBHyJnFt6mMkUvTjPJm77CwBq+o6OTwWPl+Z9942Ug32YzfahMyP/dAx5m
tzAcccTnAWVY/05OEc39l+RUkMpi5lx3iuuoofCBn8B1L5k1Q5MsgdaeC5WHwqvG
P+6rNsdxY1rMN4a8zVkHgENz4WQ2E9EilXF3MkKM/XI0QhwDg1R4xiUOUJBhK3+X
XB9qM5/1CD/MXPxOrg6Rk8rffB+mfpPPkYFjFs+s1VMUAmXWVWENpRBQIw33Q2fa
8szWc7yv3nhRJRMrGBpZbGXkiPqrSoRMAaLo5xUBEyilo8nBgoESP23yakxW6zBg
q9+VVMJ0DIcw7IO46GM2osh764MCBGM1V8w/6uwKPEcA/V/jkMzBS50wkx9zhXM4
W8C8SLpFaMETfNLAP3QZBgDimGFb/YEFR/gmP07bZqG/+f13EVKCyCeUmxW7XRu6
Tw/jh94KGUGpGo8WcrUB3F2a3lBV+0ArDXAX5d1P/DxANh4CpbaXJYpwua5ZQEWp
cGh3FQR/U2MysFG9qFYWfFQ72ZEuB4HuT08rc0vVJpX8aSNUbQ+N9CKGW0Fc+nTU
FNY9GZx5UHDcxmM3p1i+iyrTGbCqUV2umKf1Y52oM40AN6ETZlaGajohn48REOSZ
dJYydGVqoGoG/27uYdX+hieKRputMATmKOblYrzPjmY4SUsB5TfsFXY2F6LMjY18
19ZcPvljS6MCD56/lTfixL/EOPRdv/5LMIekLkdpfYmWLzHU83FVTLrSzok773f/
ZOR31iI0E5rXCshT6zEiPoK/e12YrW1Q3ki+xumtgKSLBQBj4i8jvkGwB0M0FCRA
q1f7lPTj+fMdJW3kHkZEQHvPxGP0M2zm4E0W4pChOzMqUWxgjYjulNCpCzUWklq+
K4kegACHqFEzFuIwox9TQSj5OzGL7+uq7d/Nj/QgFOFZntzHFkhl4Q8tnZPvcEw4
aPATH+y//DX+dO8hOu/SomNOe09oIOorkggq4G62YcRvzbvvHYG3q6u1mk7EzhjF
zm0G0C4Cw8lc94aJFwEi22WlCaI1ZC1edt1ijDroptXHlTc4yh/iXZRB27GM9hia
MV3zs3GFFL+7sBfxWTseKJIU70+B8elGIaO1CmYgB/cG5La5xwwCrML/W0iuggt7
QZltwIRzctn43Jn0RWPAJ5EvvZLisofGUQkgk5HJ6/rsTheAQf9uPgPsJyfBS59C
xTy2vk01LN5QsbPVvi8CYkojQRM2KJbDtgwObICHsOJFoGhycJBfHYZ2AZe9NJLy
yJZ0h+rjCX/uVtU0AYHKLSIbYRBzqMLHQpolv6b7tHAOYuGRL8q4iJXHR+3HgjAG
uvdf8ovRiIOwa6hY5lXGPlyoCk+paLsHJMX8qejAySWApifvBsu5aqXXXlq0iH0q
z5RIve3D1E0qGE2IKGpKDCsOhLne3FUiBOTFV0SJm7NXek6vjjt1Yh65g5J2wUxe
92ATr38uJnBb1K6GAbcmSPKjqZ/vClen8QwJQidSBKeeUff7ukgw73z4bgbvh7Wc
OSnjR/bKO+NlQkhp45vgSVoLF3XfJKI1AaEX1pI3r2TFDVDx3OHecSguWRo9wxi2
WHq+0QD0JQyPno944YjiJgxl9cp6WGfqe5XRVzsdQV4UFpzaWJuH1APw0B6FGgmu
bs7MUS2ry3lsvv8SvIdhML7TqGyNMmCG9e0IP3XR12DfLRc+S2w3FpwLyk00DR2X
ZeElLxoBsb8hhohtXdWBsZBMdA2vrJKi7Y3hwF0qgyEAQs6SXe86jz01kYD4Ow+I
j3Y//Xar5BrgRVsxQysQEMfZyMUxQQbilEeU+aqd3hosPSC35Lk2U85WDsRiUxjr
B0ZyhaTe2QQsBsjbiE4AYdzp+i2AB6FWsUn2WQBaA2QPr0Sdt5vHzHdoSLZ1lG3h
C9sBJeiAizDKBYX06KX5qn2DuWQ0qM/I6o75PEBMiWnSzLH66CNRStVNk0AyyUKc
qTQJoaSAGpshp/JPJrt/KD+GsNxd2GaoB9y1SERfTAlM68UeI2p8ICjzuZlvLjrj
mKNj4KWaIG0mVw17w9AUcf2CsyqDq0AfoGHfH+OF9X8/ZnsCUcMeq8FaRD2y3lJY
EBBHTTuChSG/2LYXMHpJoJO+379+C1umSx55WXWVVfbZCE/bQEvO8rBXla5uCkHe
YnoesbHOgfYkhIQPecqNSnqL2958xB2NlvFoeHJVR9Sqf0Z8liFXlaAOQQpDf6CY
+MlImYc8uanL40SPBoVaDtBV50ACYksDXXv5QN5CLDNgR0tPGaT36fIc8ci2HFn+
avqf65dhO7gkfgfv5e4UUtkbU4AiA1r8EuVmORYZxzofoPq1enXv4donjp8U0ohg
01N7IsgGVtvDwpgzqT4oLlktRocRrIn7CUwnYLSpDMvBuoL1v7TlpLg32bjwkbkP
lcCXMJhhh+HRsEUKBgq1VejIzp4WMDmzurx9kqUwgslRPk8h/S8zRnY4wrXZB36x
QlSL4lOq7bVy4yuqZxhKJI22Dum5do+rD6xTb4/+iNj1TZjnStcKrhEbWo7Sfygm
7lvB3N9wxn3Q96OQRNbD69dr0pJMaY1VRBCMI4X2JdjMWuaYfQEE4GOi203lvsWQ
Dy/LaykbVJk2wKTDz5Zr2w2BswyeFwjPieGfOWVl9NPEdqOE4DVzDRP+oN6b70Qm
KFwEioTBmEnCYm05BeuJAjMb+fy0MphlgdmEGGAl8LQ7erP6kJCANjXEgxdh0+xY
ST4lpTXlqbz7dYqNMWCVuUVz09O9VWS3XbjPUSuUMAev3NHSHb3AsSWy8nuQbqN5
DMewSAbd1PXHjD78D5S7tZ2GyDVwaL72nlYmZMZsCSE=
`protect END_PROTECTED
