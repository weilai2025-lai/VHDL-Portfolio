`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Z2lxoyY8pBM+Y0M17054LVGqMMW8bimSSePoavRQhpi+ywoghbN2lCepyqLXZL2
NVcJuU5kDrcB3IjSeMedVAQJ+DpZtx67ZRbXMIevavmPEO0iHYmf+HyU9sApIwQ2
7k7odUvB6YuEvd3jBRUN/n74LPJMVFJ5mjkK1UwIs+IpTLQHisBh5V82zaclrZFc
ZArWywassKApUG18rOJBNdZu3NDfEvYga49jwk6a/h0aWt6RW0VmjUb8Su4FOpoz
ebMs2jEFtVDMfuMsZPS0b/3rUlYYk1uiZrATiLvdKqhqVEzFsAhKkFT5nlKa73Dg
FvJNsDsYcD3X0Mh+9dp7xNr72w5mxUxPpTmTCfaWGhcBwycDOco96ybaFMuXULpe
`protect END_PROTECTED
