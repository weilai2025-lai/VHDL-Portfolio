`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3f/UUL4OvBQJOGXxAznZgqMYRiqBO3eRVwjpOLX/oSHIJg0GwgH6tFOK95XCoUKz
N/rpjVyGSD9fq15lSd7ob0x0J2P/UOcTJvY0v1NB7cZzb+Reyok8Tl+DF2mh48NT
kL2wRWRX6P0MzNowAsSLq3YgSJplZVE/MV/TpOTGZamGpRQPdZeiKYwymCpxjnZ1
WASyFo6HlBCtfaBurWeApOQaZ/HYnHNUo2TZR4nPUNP3v/ZSIRToed5dHLAI1mfI
mXALMYY/q5dBZHtKk3c2YF0aTfHfUk9nz1feHeIwuzfYzOZ19SBAHD1eJ+wctMZU
6mEYDNv2JeU0lRx83QxdwGOT2dGfmKta/OOJTIi7U6l0pDcrNpdxHtd7SUZdmApa
KBJpZxPt7UkrMNL+xuAMy82PgbWC3v2iIE1/QubRnARk/Eaq+eCpw4xwjywvIxuT
lFaXm2b858LBdRPd9SyZXokb3qCV3rXsI1wuIm5dH1D0NzusB0aS+Yn7QdO9dqnB
km1sk3pkTto0ElaYAEvIQ9tIhs9RkOTkl1wWYUijKo0UUKuLqf+NR6NtWjYqjV+1
9WXTDhWOAIWzDS/Ljp+xJo/zVZogidSGxJJq7WwIt/5WEHwSV6Wv/hPJL5nn/PVB
ljuyJzOTjyGGVKejtMbNBU/x4e440o/+GswYRAacC7su0oYlPzuSRFoqjU2PRPPa
UEJTeblteK2tuDq8nvpp4APQnoUrWoVVHpMDSi9Ew+BSBZoXKvC1Pqfx60/t7bjp
JLW71pp2nmMsGAqY35NiDMw4o7PkXZiBVliKOk3+ydGHoN9P/dup97PcclQSYCke
fxX1MGHVPXNI0QphOVzF5c4mhYjDI+bwZev1FBSIucc3EWuaKeV9RODTq4SJAj/g
hQyBLksQhDv6NxxgAp33ofLP0py/kMejjDeg1gCELQ0=
`protect END_PROTECTED
