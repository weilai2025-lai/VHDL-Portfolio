`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvAU+wKuseLAYqVEmczAEPBFcv2WcJpt8WnfPXTopr4/7xBahwC2MV/VljDH6H/o
LP9A1YLVmbm333DTI5g12cOlIpGicGd0MqIvztt1fsAOXn6cob+CCoDqLM9rRDxv
/IhvLn6GtTtWFLDiynJYCE3+efppv1vmqCKG5nclJrNEtTWuzTUvg7WCLp3Kkwq7
YkSUMsQFHoq3BEpx7SwuvRw66Ola4+Kuze2EbHph3ZaPkmPUehzjS6JlqSmLJgw4
K3yRd8cVdVRE7R0duwCp/2gAlzhdTuDjX5xRh59EnBWhLm5nk6QUVvrD4HtiVhS3
WuiUG8Z06Ci8O5mWUPPY5S1ck6MF95vNuyjGlyfy2tZlrThTzIq1kuYw5P1UARpO
pPiJEEAWDr0uRY0e52aL+aBq0ez5GZrg8b9lAa1YVKy4xOeE+7oc+6PZl4t4Q3EK
2yQFT6ukylaZNyCrdQLoUXPZNt5oIyhBCae0RtTYhmnJjBmPTeGtn3QSl1BsWAWM
YPZH3THBl34gxQhX2sEYC6kTXSvVrWsIwgNDyRo3av5TpJQaYhVV2HjKDd/EzogT
/g/1ousMnVrAzR9vkkD1ujKuvze26hB5nBXEOfp5p5R/gsp/XK8rV3hQWAko+OGp
Y56O9Po2rP7rZGlKSGEVI6egM6ZRjTlxusA8s9HecS+S6x5YDr6rzFkfpILOIbjJ
laPtIwzHRRwFECG7NT1/A9RjYmiJhUxW4308Xs1+pCjUVK8vcWrFclhkZpIPY9kU
HdBZ12H+dS52xk/RzvFgj8fdeL5wS0K8EktC2jRn58tbUOC8woFbCg+QM5EqL0Ex
Ddbwjn8Q+IWHCrJYiCI1q897sRBLksGDEy8RSTBMqqRWSgCd184GNVxO7/QzZujZ
68SiR8xnfIprI2ywQtcSra9N3MFFLXthHoK+uEqNavdc3mVnWBpMGb+K529ZDx5N
ij0J2BnhuT0wM4YHK3Kn4nd4riHwK0R8cKuozrGvhoiewdD1fZyAy3Cqy2bue3do
aCcoPvVROjfOfWisxIU1QQOlaBIeThU1N4RxrwYijBLopj9L3iWyFbFgmc6NMAaB
`protect END_PROTECTED
