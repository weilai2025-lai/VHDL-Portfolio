`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLkTAFHyygj+3np59MmN36o56fddK2DSWn/oxULxiWMKUahU0riS750MLG+6FusZ
6oqBvInRY6nYS8k5VeNjGZr0UnRR8RpSNmKvcth0Vq6UFosX79fXP3OX4WyZ8dSz
ybIfzy/xkFtyqipz5h7zZumkmrj+Q6tYiC2EZIE8rinaqSjJAhi8koF3jujXvTBp
Om/SYswZDUXcyL2sEtf5emuBqB00DPreyZh0DZ+N2VMb9OrkOQXBSSt9tgnp1tpA
ZBYREoB0l4EHn1KCjtPqZrns1qfNf1nMyWIXiwEvCFU5wp6jswgZR0JOTWvqGMf7
WjXUt8jpdFE8/+FhIMD3VlcGlZjCk7FP9TfRItclZ6ItvomYV2CAJ9V8OQ0CrAcd
Vu4bNLxaulXwKpGE+yN4yRZKcNb3IIUpdNR3gBrOn5sLjV3gOuRM1TWebi9gjLZJ
Ebw5PMX4QOzEQMLnICtfHi4ltlTWVqVaQCVQlRwNDPe6EJBgNrp9njYjiVtNG+nT
Iy9lZzpdVnq6jAUpFnC17pI8iKBFQpm1XzCLnSincGGaTzfuupv8h6fcfaH4COHZ
mg6tYqMIhVT4CFxQ5SP/gEDc7smXZBHl44szcy3ZREbL1CGrJ7zlQNHPOOTYo4Ec
yqz7mjdzHK6qFAe7tYsZT/jTO50BtaLzkXsQvHy1W9UW3gmVZPKea0d3CHsFvw0h
0FLDrFoVVAW8n7euf1B+Y7TodbYZGcSsjAy9Rdp9ImA4QmM2WkK9mJVrYs+fzcRS
K8+8/j/26trZ6K5fkpqx6P+EOJorkFkL6V7rjoTTqAFq2ju7mmJKHRVh10D3eISg
LzCxDMAogYMW9V+1F72KWwPzO3/LVLC2BNZdrMw70SCZhgvQw5sK/k2iVWB7xVCB
gqgx6ovB2V96yKZh8gRGC3vNZuxFFRyLti/O+KS8lywttcHyqCl6KGrDOtiyjvqK
ZH9bUo1WpsCzY0B7k1TsskrZ4GwaQVSSj5iJ3OH8qVWNIhd96TTtWql6RFJWCeeY
BqjqxdGxFMW1n2HMJ+H0zXyyK+oTMnR/87wV0d8VhglhbUXQDc6cKnuLCK+nLN5+
KwLu+04RTNU96rx+5DlcRmHvttfvcrpbE86DoRz4efT/WtbBSBlGrIDRaf7OcIuk
KgAPkT/KR9Fgqg48+RuzKcUgC4VcaqgQOtMP7ZqyCsKXaRUp3lR0Ys0wu51oy+r5
DIN4aZzsK3OvImZaTj9KIIeR8LP0HbbX2K6QLtwlrd62u1UlK7iSmagHRP85KOmn
NArRBGLwYkAvueS2/SYHrYksDfstHc7uJ5KGLQkfdJY=
`protect END_PROTECTED
