`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIV/+b3qYOE6ub5FxDpF6cP5xVb0ughMGjiLjYxFOudIcR0RSCaHnUuMwkSaxRcj
nlrlTCAdf/2+escBPwrTzomxkTcUc2POEAFbMNHKW/gBwCi3IvnoIqcTVROugg/w
PYQBOXZRMkztiegPQub9rFolrHuCfEC42yiO7TuO5c3GBsSDn114fe6YAWImO5Za
cEa7j5x6/BFXnvxfON+Y6E7ZorQuHIROtFjlnt2uPjPVKDcYp11Uo51hu1b9yBoT
y4xeQAMA52FpFQaEko21Yvvzdpsct0mEZq9+AYBOEqJ5omyhmEX8Z3zM9ZssyBUu
nIIZtSqH9W83nJhnle7eOZE7ctNY/UjvyPG+H5Twt9Y3bdez2sjLHgUs/4LUl07Q
T60QngWusWWqKF/TGhFN9kW3q7PWLPXXLfJTUzI3vIodYtK7lrgJA6B03Sp5iZDc
Uu1himSahRSGHiQzn/XGslXAzU+px7mdZ5f4sV1GwxpYQD/j+y8sqpk7gKQGkAon
7ioArmg6E+hkpJkkrmo9ujeL2TasPqdzg0vF/uEs/yY1Gc2Qr+3oBSyGXAfycTHb
gtsP7r2oV1lpnnp2qpINq2ACxhrRbUqlyvzR9YEeTFZiWMDEbJjJtzzTzqPkBWdJ
T56NJSIPzihYsISvUq+ZLIHuxluwsbLdAzE1fqnBOQy3KzeW0ORaepA2pQqLfuhn
OEUwnMZ0jFSmvVPj+eZdUqi5qMZmXY0zSCYvza0p+0xEG/F5mEdvHwwVNvseO9tU
VGD5jNwiHw86lCERGhFU8KDaNDYZxZLZxrq8sy3O255Rx/J2H0YWLvm696o2jAFp
IOkFGh2vxmXEZMRvCjHe9vRqCbXAmDv5ROAo1Q5WxkseFF3Zj8ahJWmJ5XowQ46v
S8CjLumj+6+tOBtJK8SuC5aEMGQKgllLu2W4TyHuQly3SHmOFVmeK2ZxJVcLlGUo
qrtt7H0A3eHwPtw855tmL6Sn/5zN3zwRn6q9CydAmbeZ+Al2+Ij4wMQ+npnuNzzC
LvPn1a/9zZyfGhzKoegxpdeAh66fc6thsEiIq46OLVE7SX5/FkOoCmXX6/Y8nvjX
jqieo3FXsY/h6MwbcBSXEi/7xjpl29pyTDTtr56UXD0q2cZ9KrrLowXHPKDyk6lD
OPlLp3jhsU9KvJl26fNG8UkWglaNAMa5pBHR8v5qYUMvekgERw7XnybAwkUG4Kta
Tt8D5a2W6PehS5k4SNl3i0PQSogBgRlyHgrYBgRDKY+qQfyQ7/Nl4k03j0R1e9SQ
odqaw1f8GhjVkbkri1DDjDmn9iAa6DesrM7BPLNsUWEOQCh2TYV+IkTHx7+on89i
ZYs57/FZdWrVWakZvwnj6FOi8IukmUtgh9Qcsho50DyiGSirTFeWbTo5K4oknekE
wxHH9kkYhN2NNIUeM+cXXeb3kc50Jz5+h/jqlrkQXig46tGdei4pjj+562jlX3c+
/gqPFGEySQnTtCrYqhf2lvLVV2E8JC8VmkXE5rFsreyH9Hy9+o1h87f0mrgeYAN4
4XegKImtwp0q1PDRRvnLzmIBSV1XS5fTJuX7zcz2oprXgnIldDDqlc31Kh6/I+J5
aFJ3LPcb5EftDgl1eNJg4laaIG4BvGdjmJQ/cNW2QLvZMnfhXt5H2hks3fs1eMUV
GXLPONAR5DbGxFLG4CFFeRnu7gPBsPEuOMs96CP7wIMXVyVyWP9NZmR3FTf/r+GH
ngAA0PKbQYigJ9kygNHxkvDy0E/Lu1/pNdS24wdx3kpmqSbO76/MBKl6jo2MA4We
5z0tOmXsflEnpk7R2NosX52zkwdOHWFFtF4+m+JhCfCRkNG1osKM3GCnMhbyN+u6
QPSiPNwcVEq5N97qmft8OM7ssZVx8+OB6Dem3enOJMLsv6rp/TfbcYhWGINOBU33
DmTAAC3+lYoTMQwcjMEWaW6W/ApDWEOAoU7ji7uFsVuAzdGLrFCEyusEGSV6Uect
/xQVkSyQaD8nZOCKEgWm7uzlHInidUwdQNVjCLeUN2V3ZM/ArmDbe2GgsD+upAFb
GaMATVJNeplR6e0Xsqiapi0K0cS60Zdbjp1wQ0DvRLfQ4Vip4tmDr2WGflEgrLY0
aQmSmhY6MHOxNmFpz08bj5NgH0ZvnDzEn1thN06uzDEfgMh5mNl9uPUDgSQS6b56
IGr3f+tJZlOnuORm3z3E9FINXMLkX1XuweC6sETaig5aBFSfEeZcdal5gCtKQP9I
jDR/h0HN+zvPK+eXT0/cV7uvnhS469rZBLPxOMuxHCRjOwWzh3V/W9JgloUBIC/4
fhRyy1kBiQFZ3lw580WsI8+5VOgdgq0bMUOBvuHwqGNbeX+1WmsLVig5eHtlxeay
nY7BPYtXhfd33diT8YcucGgJUu0F6zM7G0qskQppnQ7lhzP7vMSU9nJEW7FY0p+v
sMmm0jAuw0DfVhPwn8SaT9cEH6S8t87vr50G7FIJgrBtZ20qO6DS4jgCGNtyvTNq
B5nhEK6hc4Xh4r2ERYFBz81azKpMI04Ea7urPnTIdmTH9fqrXisOFk5Cnz8+hUHg
G6nBmyhxVadUfkSN8ynSZgarguseis9/1vnzWMAiSQRb9nB7cGUE1opEZ1qblgmj
5IQ9PNTjJn7jp0AkUvrk7nCWcBYCm3Y/6j3cj8MGhwEvEKgtLc62pCm8Qb1q1fnX
wACHEhyorpdYJXqZjBAiS7bIW0ObSng60G/ZyksArk5VF6ks0hfd/SPUUUxQlMvV
DYdhz65B1GJldl2rLfiDsb8keRTGaQvosPUS5XLJfxIXOqQDHLk2kd8iWHxx7mU1
mGpKA+dNXf6kVf21H/ygJJlTWn136Il+xbxwOr2K9WqeyQhONh8aJF+k83/x4fTL
QGHxN3m0A6gmJjapvW2RCejAqtKaoxkowLPrUQBXB7a+14qEmW4w56wwiNN5We3B
B+D22XtpvEzH97c4IJ9R7mQcoXs+TMGIjXYSpTnYi5Rd5qNPzVoS4/c1o5s9Pqeh
XJA/PsOpRlYl7aEodtkphT7wruqnBGeJnwoRRR0+9aMj2LtV2zGZSyjXxlho0xsE
0VlGvm78E+nl8GTcJ9zpn1BPYMNLsh8YhiAd5kVqu5LWavRj8e4rALED3qiWi6E7
vrBJuorjpMJCjmdQBhJCJ8P7odg0tf2NI8hgGKqR94gY10iY0CCMInLwz/nVo/hZ
lbt84JkoX8PjkBykS+UOh6FkotXK1HZMWv+sm9FcFryhkzlBzi9p0eJp7+iRDGpq
4kfoTsUVOZ32PoIwmzGSvNg5UuDtDHzhlmWnm6ioBOuq0A7iLUT8JrXgRM6i2Mdy
x6cupWxoTNVztfGcq/1vDqVjXC4u5nq/2AyaBw1nfWNAJD/9A+Jvi+AQY6j9QGMq
sl96j0T8DcNRYjy3ZhqhQ7yDH6mbrLHqgOxmyOptlU+NpKnDiyFtOy2Njk2fTIYo
9MHTk1McrI2fSHClaJFDvAPb6DbwyvETVIAC24uJq61tuPGJYHpwj6TYhbTLzWkE
oHlSy7mE/JXUR1S3atWq5ig1P28LDK+lfXfWu4T7dQ+YNUzr/V8N8mmhC2ujdnzD
ZaIGD0FUjDbSN43dbqa1aRnbnUYOtxs7gNUhyYG/THW7heBU3wD0arEEQE5kCF/j
r8wWV1NZTfsskBT79Vwsz4iow3uCa/yTk5NHwwcpMBW5aGadaxt6gwaDWMW87GdE
hzo+QYt1kIvDVF7rtBE35dzguYgq+1uyIcem6MRf3Pv5ffg6YmE6ZJgNOWhADMzd
YWbGXG4/lFhyqIS2qR9X1NgMeIWjZ98YivdjLQbCkT9dpQHnLuVECTbD5FOXcD0l
FBP5259FKbytKmwuF4ZTyD1xTBmedy7HPin/uxCSZtJ2HXEUmis/QKNDNKgV/JqY
NPk1l+FJTnM717dnQbKQdnzkeX3svLsltmveH2vaMWJgj/PtJQp9hEWDLFaKnnjS
WoQ91yytvQKvDjv+ozFhO3PBoU7TcK/Z4UxCC7a48ZgWaEiYfXC2NK2Zd7h+9o+8
9c/vasq7AKS21jSj7alXiOEQNIGAztUPoq8PvYMRC9QcGNZJBiI351mMHcd8/MuG
Z2KnujtmGbpHVFmlGUx3sMqPVEZ0VFkZ+mYXqlIT7+HRVL9z2ui/6BBHlf84fDZj
V8pT0e3PKMJz2R/JSOUyye6i9bNdP0KVYxjLCr55nV6SSThIsWFNiJIM/mxE1gQF
sYpsGux3fdsQk2c95hljkIsQ1Qjr7s/8hu6SkunODeQAYUpNogacqQN4o+t9FWs4
ryx8Huvsh/Ik93wc7+xAQsrT/e7iYx2SYseisWlldnEwgOsNSUv7Nf5TKPyM/IZw
oaMy0ThWcPcIxafMvsnJ+VuYytBBciUy4ltqtlPS787E9q4c5zbsIxDCho8mcZkv
xvs5FDBlHNFoRcborNRGQpqPzbwWxzWbDlEeyOhy7fYgjt+UwAg0ex6pElhHjpQl
xy1lFzjCLSWiMoesMP8oEN+cIvm70MPcj6o18msrim3Mx5wv5lM/VCJenGT7e4pX
S9Z/YP2GAvpcN4GFdk912rmiSgR7vnKrd/JPKO1yHuvG5LH+RjsiG40GJwEDn7Bv
ee0nZ28vo2Dr9lFLIL5GciE+H4HXM+ODAdgtMd+cGM+QGRiHwuvhJp3wCsginP1G
2h+R8iOwjDzs309TnkFkCTQ3AowC0veW2dQ39fCrnzcquwClMu+uLP/3vTPcYG0d
n3KGnCpGCW1Iy0qi8zHmoq6Zs2AVPwPkUSIWD159yMwFBebVR+sULtNcVJ6BXy8B
oiEZy37BmWTp7KDFQgPCVZ6fSlMGwA9xoUWQ5UraLy+7Xu8lum2U35ucoAXkzKjG
Nb9qadvb7BTxJv7dKqrPt6bt8e6uBnsga/bjeQcc6wdouxFOGFB4jXJCWV3vXMQ3
5AthvyG635H9x2cHwR2ePx0Go0u3hemQQFZgNIMmPf4ei8nlI7+G2v3WHFroTyqe
m4UkFmwP2NkprzrjtvR1Gn30NONYsrizGtru7X7L5MrkLobt8CcGL3uB6EKqr5Nh
coS1doEKsYZLc1qz37L0yjDC/7RFhbVKgc2xphFboHzITgsJFe/Is9HWOUTFAGeQ
4Nk3GvC0Dv3wRTJlw7eL3lbmZv5cW4ck7y2IWYodE81klQ6YIXAkAWCTTEpbWkGB
y9W3jiQc3D+hsAyj2lvWeW4uVpSyn/sPh3zyqwUF/SqsbOckbjxLfsEXpsxhtRiN
DO9Z4573iGJ74lLToUdKe4gg2mfZ88A73A7dwCmoc7vZA3IPKOknIU9+2O4RFVAI
`protect END_PROTECTED
