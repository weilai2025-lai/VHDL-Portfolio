`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qR7nKvFKFobah+R05OWFSA9vf/zQU8i4xRyIdaR5GpbG+PUg8rKhgirUwfpOw3Z
zyqK8urC33/VmzF0o8owK5OJCnZ2J1CbxfJ7TDKR42kcUJQOClN6lcOeWxdoODkq
KUkLDFxpVPQzCfwA2FRRANXPn+uHAuDJ3I2kl+ijQd2GMY/OAzJwQkbdZfZ/n9bq
5gG+J1lPrT058ET1zgu+xgHVdfdXCUEue5zbZsVrnXjQBvg/HFw9kM227bL5CMdy
qe3sroL3+8stWG2/01nZ9HgcecWBhg2ii0Rsp8fql9TYSiEGtG6VtzqdSz5GVDRx
B2wCQlrh9F8TAfG5bYa40ipGfdYWfBjZyHuVwWCfdE34HX8rastHyi0aV2RoRgFG
U/hJDlM7Gg4n/krwHWI2KLAky1K/9ObORh+V7L34m8jPWFkvla5HmsPvdmQacOhQ
l2wXFySN1+MX9bAXOgwjc3HC4sQ9656fm/PDEYhu6y1pQ8dFaItbfq0qxOdFlHUY
rgm0PWSFflMp/dGDlytarElTpII5SLsKFGBSfbHrxnxVfLNHtbWhrmfDHuxi7yoC
+iUn+Qxw2kTesz01iQpidekx2+fcdBfugvs9TvMV8vL3IubNRWC0hUo5B5XyKR1Y
q5l06xp2OeV6LmzWTSjAF2R5LES/RmLA88TWg9icB3mbcgYJg9lfRhNvwsLYYkGO
oQtzmbe6a1J+/+HaH4wArtY3LUiZ0BtWOJmagpgH1bjvwxV6EoJ0/1xDhIUzeIy4
SWpoP7MdjlD+Bh9iP/tbzxTOKv5RNFWvzzJL45+oNhISdtsP5IYdtg043P8KyIGL
tbMf4e6eUHmwGi8H7Ud53VNcqJefroDnvI50e8GbBREZ2bkA0TLOPtp2U3r/yFjq
6iTKkpo52HHU4ZKsNs4OtD2YuRm5zTdY2KU5Ve8a+FyBa52/dLEgooBBt4ieq8/W
UhMB5fSh6EzucNewRpCnPDuJWRzzXSEPeU7Pg7zhPhqVkQXj9KxjG/KOB+VITOsx
BeV7e1dkKmQH8EpvPYBURldYWgpsCNOwt/1suCLM3s0N2/mODXba52W7GAuRmNjw
YUkbgA7ftC6QJEJeZVi0C93vKsUcLVNDGdT/1d88BqqyOQKogK4VVft7M2ThI6/n
jD3A2s5VcUmdOQteBl0miVhPLc+rF1/b90LTTTHZJAZwPLTWr6nuKFTmCjhNlQqE
zaKq/EmZj7EQnVV6l0peAo0b7Ni1h8XS8gLN/Y/8wDAJD2uyBkZmDcwxRSutFiD2
DE8E0SM4wWJAanD+CI19/qDFlpdcPOFITY1RT4CqypQm2qNnWh5WRWEPFwwpeIIb
trs5j9Q9m6F99RLPHsNZoUYLnx22MB79Z2m7655C+xyIozE6HvPEfb+ADsyw3iKN
4nR8CEUwVgpChP3Nj8/WYftget6whg+1IfjjWVwv8hiLueWE20GgijD+fAEOxH8f
xgIvSb+OFN5uKN4N0PykIpZpEBGTFGgEkEp9WvOMiGGcy91Ccb0rrFViQjczwNIx
wrNqR71qn7zEgi4homFv52WRfP2oZq+Q/AI4LsAW/bzAys2M1mz6KkBwV5pUSg+X
YXDP0LSbJUcAUIlB7EAiwIvzL1yOoHiEhE4wNW5n2XCprpel3m6GsMeOXxv9J0Jr
qOtqfRYVUi547t7ANXEsFx1yLTHKBFCbkZiohM2UEGl9SXVNp9lgSdxCKYW4/xRO
BlMbf6wuQcBY3giTgrzu88A50Z9UNjV1VDJAgOwl4y0x18VL+HtKcY3c969CqvXB
Ovr1nrZ57KmGQ68HLbSQRgu768XKvZS8/TiBWQzpr8qJ8WTiTjsoBDXpqMl/Xt+h
nTsOdlkrpQ/i3o3+/sdVqcFwfSh+HuZAOFYZIefzcVdZH32dZPCEQngVD7C8Uqlm
6ng+IAYE/peTxU1X5Gd3SUSjTCAyJ2lEkJQBtlbRu0TsYf9cF4fmWX0GILLGlCfC
MfurSUYTzkAFL3JCep1Oqp/H95HO724hylBrvZTRqH72ekEhZGqrJ0+Edhkgsim4
BCwWrbwmeb0nmG9E78zfwWmFHtG9WlBO1FXtWH9CBnn++/C2GXCEPg7ek214vslx
gEkHjlKBcRt6WHS4aIDL1zArvgg4s3lBW+indbegrAAITXfC3pxZdKHNjl75AoZr
m6f0197CGZTq7IZr3njAaWspgLvjJ5dbltJtwtTze7eujlFMQvDIYiBYcXoCBZd4
Idne2LOYEbOF9V2Vfv6Q71irH59dj8Q4l8PkxvRbv1X6HMALcxQQK5Vp16uh0+8c
OQala/KbPinDxj80yzRKEBRwzDea30MYlME43xcuXpfn/H4/8o6G7gFuRIMWvJmV
RPzzdwmK22EonKi9gzOOBNqa3tMCTVDwHHasDkVsdBpJSZA+A613ifH7emr/id3b
PlXTeHagmT3oJzVIYGV0nI0mKE68ef9ZwCNvZrqdruZescv/QCxICXesrAI+g0mb
8s7ZZyuLPWUXnLOGmeLH3kJhleEURW8EZ2MuZn7r+zRjNSBN5gSlrzrc3obATqRb
yLCUWKidRFZmpvr+RAdakULHs+UNzvRTWEVYoGbclTkncw3hYtRAaO9R/yEWN9HO
Vu7JuCS09ZCJPdPGUvoWFBZt7peCTnbMlvMe/vKyrw60WVIu9azw2DcniIqbPUKs
W0/AMTl5G12cwU9Ojwot64DLzumBkD6Jlz2BAwDFJK9dqVxYZAq8JCuxazytgmC1
NBvc5e8jeKHswhsl7uYgqRdn2oy0NW42PabYstyPKlLHl3F/i4CX5FlKqAScgpzr
c1c4FlTW0gSsJ0tNATPvVqCIiX36bxlg1jc4xnngkcguind2A/U92oc4m9iJajiQ
ybf/5iUosJn1EYsXWv5VK5H3JiUmj7/eb0t8ETsZKQkLEJVKIC5+9pgZHrYI6D0c
ZQF7cYiRLupF03M/1mg1PwBt7EZl+w0YqJgRQdzc9liAMaNy4zpfZSbStlwXzoFk
P8NYlJ4O37SksTX5r354ep5j7IfXW2wX5k3EsNvnh/a6l/rPgH3nuVGVhLZ3p0k2
zqMsvHGWDm01SCfdaF4MAESImjEeY10jxS+T5LYV/PvDM7EBwKXuCZ4u/Okp3IPy
rumZDNAQLzCd8KPoF+dWSGWvH7xngEzN/4NbTfo1AmYB0yOYpjyGX8/FVOVIZj+W
qtLVG6KVDU84qSewYaVYNfy8cw5jyT+HTSU6RaR25FqdnGl2kwyiCy42eiQykv4H
1nNCZktFM/glkK4hk3soRAMLMOODmRowQHnsmkxCNFiQKWiOaTKxEfUFaXMsBE7G
qMrGYKmgKWblDrXCK111y0054HgB0bbWcjDJ7HmbxtuXVQkyJjV8um1FlwFbh9MQ
b4Vgbu8R6CwaAIPTvxZcFv/BiuD9zbyS9FLUqmX06WqyBsVuyAokavcQMjRwaBKl
dXtgygcRrlDTWwAXTxwf5XWD+mOekB4d903kcNe98qJQZ/WRZ6VdIuzf47glcqoT
tfaolwPVZhu1JFBjUvY8CCHMfGUxB3kVYYdUm9Delz/CwLc2Omd6+uzJdN24EoFc
9yUUwwFUsuF4MmxhrZnXelXTQRkfehPEcV73u+/kkyecbfXEzUcz4P4ih02Zupl0
cIDAZlxTh5KFhGxMgR77lYuVomJPu994mxrGenXvdPcdrRoLpqDGPEmu6Mt00jGx
B7R6LeCRp3BgVlW0mLCTnM0WmNdUMYmtT6ueG+NYWzAyjNqhazx36VaDW6sxL/DQ
dIj2+VPmI60KWlpCpqUCXidxz1LFKZvIYmQkmGegYDB+oa/t8IkYIiSMNb8c886B
Qu4eQfe4SvNQNXP0mvJk5B3lHO1aKEMsRRQgcNpZh8shzPwjiE5X12wR/sTkquuO
Qi5z31Dh65J8yUzwitXYCTaB3n5xyFyIMp1r+SuzeH1+yTgny75ibfF+ByCZmanA
o6Bp2mVhciLuF6IgyO+ZPz2FCn/TBHxPMCqbmC5QkoiilFCbPjaL6lCz9197OdNZ
JFpmEnXNgK3CWvY0tCnrgYn71oE3JXYJ4a3C6gSogbT7VhiDHyKw1QXfs30X3R8T
hPwebyH5uZD33pSJNDF9JBMFU4QXxobZAnFw6Dy32XRXVBFYnoBGSfydMzLyKksg
eSFPnHzebKcCiMbpUTJ00MAVv60BfmJQk2WYEZ3DmWTlABGfjvvesZzwMyCJ3MSr
CDEk7Z49h6o7Q4lt7LqcGtLcuMRrNL+FqAzOnrdUARKR76csm519qPxPdCysxWkN
+hlS7oRtPCWDe5UshbWu/+tjEcDibsjONpmWQFAZtHDuciu+ybHOoR8zIh5nnLlG
7I/tNtSqlbch7eyCTsN32HKK4tUb1hWKj9uQyPlTWqMmXYPD8gJjQ168JXcShAlr
k1vacByGp4+eC9TVoAJx7thcWqZ23Ync5EITdQ62ipAz5Y368IBPDTBxcyrialEB
hhWZbo5Lm+jNv0KDyjRr/Cch3mUBzpUXFjd3EoFl1mQQREHs00LO4v4YyCrJ9WY9
AH7L4I/boRc8td2Eq1RaxGeMKKFlr8McqM5Yl79hiUr5b80SHJHYxm8mtOg5tcNr
dg2DLc0i7YvWfMxAO+JiJkEuGDB/9yh7NgMQzlQd+4O2NpG8Rr5eOXWIVGWfVSef
whrUTVNMZJmjndUpWptebk2KwGl3rX3Id33MyI2FGypJi3/kfqGqZeoqydhBej79
CAZ22dZA8gdy6jbRFoSsO6C4xC9O6BioQSL3CLMxcomqpdKyzD9CBt25GHyyORCj
eH1EvafQsy4OzKOVLm+FXItQx9+6IOyW/cVL7FQ9SnlLDlnCrnNcnieKEChTsMVx
V5n1CystGz8rl3kYUOUzWo2rGgnK13G6TWbvrsZjEXwLxKrSIfNSetgmfZp/5gCt
sZKzdgDevb3GZAezMy2xnU4oegdsAnpvzh8AEaXhiyM=
`protect END_PROTECTED
