`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gqj6nVvoSMyYapcjB9nJEYTaTN5QEqOUXELx73TNb4VGjSmPjRAgedxfESjptFgP
RBb9O4ZL0jJI8nqo/zoOVAf7C7+fRxaJQ6wXx+2/P/YK4jsEHUYL/sGkxRR+jdiu
BYqLD0b54OL/3xnImRfJDie2CyNRHwEynF0SgTOPb9DYoAmG5uSvCMeH2WDs4V5l
KFjxeVVutRSyXtzxOih51+Cdmgkl6O4LRljEuK4TSkYY3apV8dQFKycJZ/5qM8qq
KXP7XK0WR9jQ2T2HS7Rw2hVlvlru/Be4Bc9JLH4GuNy9S+I+44lpE21xLOiOqTk2
OftkJv2I2l1rE+9y7grlJZO365WP9KnYbxAnpCpjT6BSu5hgCB5qBCdxspgnTwag
903kJOeplUwfCLaMctzXEBR1cONCoIVT/VVO6rSrSDPYZdJEEa2VUUSnZ4fqAH3Q
BzO2vMw9SUSsULVsr4GfpIR9AzGlblyDuVnA6Bq7vD/wOvMcI2VrXySZvNxFlceO
vi5dgT2mHy0ER1TsdcJFUc8TbU4oLSZ4ZJSnywEM7N54KC9pYBKGWTFwx/Ab4icw
D24pIcRZdNyEuCMTmQRxzMnxmN8TVyywCkpUUKZFNpqJiPZZuO3gZFwO7VqAu3dh
0St6LD2BAgD7AkuxDW+Ney+FdIz08teu1nxbpPyeuVxmR8jlxFTu4ambQAm+sZzS
OffFHBqfH555gpBHv6pD2I6/0zwbXhMLwYkJzIT5CqxJx6P0TUm6zHEjKsFTFaTf
fq/fU7DmeVnFUJlLBXwdbqJbZJxoI49PwBQS6M5OeaCzTPya21c7GW+bDjeaZU25
9L06tkO5HGjsmktkPo5JTQ==
`protect END_PROTECTED
