`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNvAjL0u05XoqgpCn3Ahkk3yOAnhoMDTPvlfW9JtJq2LDu5NzizSlvLoPi0j0aLy
3RWk5UTIgs9PHx91UWw6xxe1m0K7YrBFYDLq6WPsY1zHI8LJnoN9Pmi+fC3KcOBl
PEN6CZD4XpqGSrmVkQyKTtlwznDm76zSlMKW7EM2iQsuBhqEhi9eBDXUXd1Oz0BI
ZgvaihPxOFyo8HMfzBJFj0ahmHOezQbgSxpQw/133GeCA6RmAxQIZyAGAPvC0sRy
eAM4MMQImlVZ7ehJtxMc2/QcJgzFTFe99FeIoZ48ITOp63M3RS7Vyle81bnafFOX
MtpRFLO43LywFVcgcwPBU2PXp2O7fkKtSE3IZgUflSyVLQ9AgOIlu8Svul9+Z073
ZUzlXJDpF51muBE9AlPK+Rh/Ar8DvufdTjXmgZHp3U9rn2xrsyFiblqdRI28QvMY
ovgVEBu+Jh7SP5TnIo6LhBsL7WU15Pcf5E2utPGK5Yv7/adHOhi/Uw4qEFoPk9UB
mTgzeG90JLFN8YdyOSxpvMY5M3sFtUvweJ2iAxHhZNwBU1mdS9VeoLdNfQmdb+Vm
xf2A3i01VtCWqbhFAS3nxFUddd8zPBad1kTSksHzD1sdLRPx4Ymgea2pYwtVjUWH
02Qj1TEQ516GsjmXavj8xYBNXRiDpwcR5hf0DXuQqKDyf0ETatXVgja7cNA1jAuV
9x6HbG1JcpAW6gdePZdb82mVheG2HHV49lX2hCxrBogbo4ujhHLTRN6M/dzrzvzF
EalGbNj08flsuAfufME34ISab93TgI340zG3nj6vVA/aHldy1e53e3QcVE14yDOL
Kria48t4sqZxkjVYbDg1v1LCi2KedTgDN5tZaP2AdLCIWTqRpqBK5nSRYcaP1QwA
HMQOg0gj4dOh5EFi2FSFYPg58lEdlD8h7jNst/7PQ/Dt10KgyUG76fae3x4GqjP7
W1sTxCQbRUTaX5U4y7U5DF8AxZcYpSbNcS96P6kkOPB/ruWycW1D3JONvmacSuIe
8Vk9k27AcDhf1Qth4tAIRIOKAxaeazPgPy0Skyvh5HljOLO+zQVFyCjzGbeGFUUz
JLZEJhRH+SrPx6IEdrDeCi6eewIQvUTTCBU1fC5Di9rQsZK7+6MEqdc5HL+5BgjM
RHwFoJsthoK1Xp+npmXziJLXLDAdTto9CetNQiLWtkn+j6Qpxf+Qn8B0Jn5wHrNy
6hVRKRLBdt5mVpQcGkSyKqHz+dgZw1rfjg5hGHQbD5cGJPahy+iHPXYqKwgJqkB+
KFNzRrzVuM2CU70QB0gOGpIVXj8p9oovl8rwlRK5ykNuVLGwmwS83xs6jhiWgNz0
oHma+FdzYskPnn8+84tdC+QeRmEmUD2KOdfE3Gnf2A3XpKZfzDMXeLFzH8h15cZq
A0odM+4glRl9EW6VPAitXKtmZE3Yh18Lqbs+tIYapoXPdMztaKawhEa08B+J/gDj
xq0Heh5vUt55CMb3mje5wyshh3Wn/O1QE7mgDZJUk26wU4lthwS2rP+xjllf7imW
9+RtKFm75/dhtS/JDNpk52fRF4RWTQykVAqAxpe4s+sF9yFrHfPA2fzsh1tA+gj0
g7yZ/cS31GysHbqEeT71xBT96Y8ehGXcbVGM2zdUEcobsvfKe0XURFYGS1B2SOiZ
WHfvORktU1Y0jPx8Ijm3vAZYHhC0ja5T8S27hu9pdpYuPoOXvJ6s/fbCaEjaR6GR
cLXANDOKppg42zBuVPnc//WcNqy0SP3Ac/2dZShHr3zWiAVhdgTGcZT5tymIgv4O
ckROC9Z3JS1L/qU+lek0zERdRww88kKz9X2CPC1v/Lg=
`protect END_PROTECTED
