`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
95myEPVAh3EDryFYX2LRAR3OAQaQuMhWqv6O3qNEKPbLqdLtCsPWAVm4MSBEnD1n
leyXeQRGne13aTqGnlxHu6di1gD4Af4QyztKmRzIFQtgz00c7efPVYmaOEJnJ+w/
6tgcrP4Q9B4XCP8L0Ee6xlTILXwuscjeNF3BmfUjUkejIYYHEZfqP8HzvNpFvNhw
bCu/k9BY6yZpqW2Z62FhpwKI1CWqpO0vaMbNV5xDeG6GfqMQsxRBbLLDMQznx4fC
bb1Ndpr329KN5ksZaVwFycmDDk70B+R9b3HarYPV0wJy/XGA+qQ/qQVAnw2czOUl
TuiBBoVuty0AZI+3DqrNOWYy12XDqnNWnLZ6kVv2I5EoUEwRvR+GI8NYfEvgk2FF
VeI1UDHYnHYGGpUxJtF4nB6gsv9K+ZAdQpFfE+GHTMkFP1+EAmrNheOZy3A4Du5D
Vo+lBCYHwWbk15sD415TWwXWt87FBqUY3A/YKx55rvQ/6xNEm0xXHOKH3vVHgHzd
687oyIIWnkFdbSqunr4QngGuM6iydtyfALB4Pxb9kRswZZNS0aPmCQoBNGaXafJA
gRsAlwTznwpOcyzHeZru59OrKnT/RHvLUOBoTDGw8SCyy2Uy0gdpfuTz5X9of9mX
1s8axLLSEpjxtWv8Oql8aN0hxGQamdrz6JKl/Bh/mSW1mIkBfEnhdekVebZRuDk2
CIHnBrDzTkeRFn0jzHSZYSpM3qcQTB4n0ZZuUa8HbnB0r8+sPCMkBwlRUOJrh4Vp
b+3Tb59GkkeT6XISTNswbVggkdZ0KmzMqn8/ucgnl3Nfxv0F7ZsOvc/z7XlIHet2
GfMut+5sY2GRODKIllpn3QqPXxlkGKDcnNJr/S12MvQ3DAW8mu5cUEGWeg5V4s+D
Tm/hnPTlsg3scVr+zhqSQEE1C5sn85ETkvzNRbY+DxtcaVz2F4sFm1fHIYPwq6M4
72eq96zdkNCAO2JK6Ek//PtTEXGz1NPzkGiGRR09H5QAnwQMUa7x1aQZjfHaoMEc
keDeyL7ZxLaVeT6RqQgns0vOKcOj51C9LoB45XwXTH1aFD5mwWrYlk1d3pS+b9n0
+vXXmhCQxKfUkkWnxk4OiH7QMit8k9n7AhgNyTFfzZ+LoZcB6ymh8OjLxTLQ8Pdm
TIrWkAeIIdLPKEmtWUhCGfnZLrVNvf+xisZFKyqvo1Cl1vG4dHIlJkQr5+1S4tRF
O0bVpp6vleDK0OI2EdtX6lccHgc5KQoR3KDfjY3TB6utj+qOhY/zx/SWQ7eyCbz2
owQ2qlQGqbVONn/49YiEBlPJfI6Iei5DWo4bzQTfEQ1+OxRKSH9OYghF53wq5g65
hQO9DA7xRqtBtPS+JLBg/806lR9JGxN+rXnuhDifAzGzIWayeiNGCvHFzPOlh0Do
HmdaJDMJIdAHo/qoBAx4RrfZc9Gj7c5qnE6bRxiVl/5kNHbtvtXJANrL7+ZgCrha
0hiCjbvoXwancrZ0F+DuaawdUwvFTLA4WPyr0M3FduIAt6fZlBrkABiVffFSGVN9
5Kg6IwXPG9jryWXLdzpqM3xDoyd4HlG8I+hL567fuaqPnceFUaEjqWFy+9lCATry
z/He9lceFqLk9HzsgPE5d15YbqLkfcYQ8akz4wtmqsUqchB+k5pvE+Djyi9QUFhm
tUAeVA/0fPB9ixDL4DiUBewNeCuSTpjvXXqZg2JdXzawlVY67+ueoIUUxETKSb6m
lhts1w9lW4aJOYfX//FCfHTghAUNO9CDFrGgfj8nhvs5B5ELBPGQCfWJ6fJJTV0w
LTf2tNICRrXW/FjOhxs9NK9xneRrRZyFR08cdHMWjsUkK3J7zCFyCdzRe4iEU5jd
VwYjAeXzB6YSzARRPEFD1LzyEtonYcHDNX7b71hGQaQmVSDZZKAopQpeNPi0vHiY
Fuf/r/fiio/GN58jB8OP6yby+mqmarslg/RVeNuEmt7DAXmQKLaszUG3tLN8Bzip
pPlhEwOuIxOscrKorE94FTqy32DqUZf5l9KY1NLEUn8uehMd1FStjlrZUggR8jcW
ssegQLjiMn6HrvB3cNZM/P6H4w6rHsrH0U1VSH481CJz3RaartH/XPCAsL9XUqVA
ge3Aq7PEfI9Fxgfo+R451OkwqVgzvGhIk5Bj2wYsmp66N4R1xAdwSNwaS98nPUfa
SXf0xQJ69dBDp1WE5Gt0b3VqkmM4HdrwjuT5NLxw3o6JIm8d/j+SyjVKmYpk1kO9
Slne2YA0byK+RJWMQMXkvENaEMTt0AtEnfZfSSk3DP4GPjjKp2eMCbTWnE1jRSs1
n185B0qm87oC00KAJG79lj09zUytlzTWtYz9b7vzVoSwTVJclMmR2uMEi/1HheL9
hgfbMKjzuJWy30d3P5hdOp5QP+ehn5RvVu5t95nsS8L/jJRlgobFemE2rVbkDXI5
lCV9y5QKJNkMWrH4uIEfueI8CAoBXKjTUvKru2v24rwaKnK8i3ry7cYW/3fdPYpi
Q+EMO6sgq5kQPwBTikyQ5ixlgm41+0VgtHj8BDH0TIRfC7+ykHf7ggJlgP2e7kM+
QxWeY+iRl/nImwegztZLdDt1Kboht87WbttPMGiKLy1WG5AMdk9ozK/QKu55H0tv
pO6Ws/rwB5RCUc31a6T2XRrFNIN7J7TMD7UYSYrrSCwY9JHm/iba346A48GlZQ1t
xcTiz6/cr3T0olkWOf8mkJp4qi44gFDeIQGmwhThR1hNlSmKGaLoXTAUBZbVttXx
0hwdjS2cnvspwrmK0uUgQE0xoVVtRxOmm2c0vpJshdnUaeH6FQefJBfflP3aakla
KYgo5J9SeDvQNsEPVbHz4JB2UepLRKvOpFx8MVToijrOp+J2vXadIUbjH5JYeVYh
t8cRGamKAcGFGQVTUS2IWU0zaH6sVgPZGC0O8PP6mg7yzVwCgEzV6fq80f5+xWMA
FcVfOwfn3P3+sDP+Ga7dXwlGMyWkppsYRmUPQL4s0Dd0+aRnZ4kxmMHdHK/9Buzj
uZ4+9D3GcujS5XQ7u14azUX0Bgn69L6BK5nMr6/5d9jO8OiRN7Li0mux9WYgIybv
HXdo6Q5FDBvczU28NKlaK9Y4k2UdU1CBal6BglA//anYBExMotIZMgNeuOvs+n6T
8+jvt2NPejXkdopnnVsAtQPKuSyvrDqJMFsu+Gh8NBMBsKJpRi/ec4j1bWPpriR1
zJ8UJr5UqfcIizZsGgR+3woGgSFTjqHbnnJbNEZ5/OcjIfhHez1hP8kkY+de7CIV
ICoFshjcUMsvSwRpoSe/1zl6D783DPgBQMwCERr7Eyqz5qYHxjx2Wmjj+3U8ljTO
T0UmN0SSaOvoG7+wKCDadnDlPX9ffodcYUgAY3iIb4NAQrNYeOxJC+m8HhzwSvma
baXIzDG/JBLQ0sRBvBQImHllgRBRESXhc7VysArWwux59g0aD5e9Rs2VAbPkh43u
V0GGo/4+A4TVsAAbjZoIzwSMCiyywj/5pPry6mI7zsMLG8rBp09zwPdkwjpLUxm7
gcDEgvw8Mu0hXiCtiCXyUq9mJXJZ/3dmp5phnxcgDF3bGiHUtL6USf/K6/c8fAKN
UstQ57VPqq5U3K9hF4yZKW/1dpURfI23gm35zn6BAMylg4hXICUfKmAC7ae7HtM/
LAEJddc/gpOf7QquoYmfhbJF5WU4Pnfcfxton7WtE6eum2DFTHZ9WMlYTNcf51n0
a4+x2gK24jbG2fWK437+Tduza7v3ZCKmFLiWVscM1uXk1Aw619EF0ooalFcBT39Z
BA+xdgHAhrIsKEr1Ty2mlkM6prFukE/8QisT0xvVz3TumKLkioOIvylo803uFqPA
wBXbyFpTP1i8NPKh4C+PRy+DH1yEY5Gc5hBTAk/07HeiT7X3wjbQwbyyOxK0kmcn
ZkNT0ykl0D/1CXjb30VkcdFFjKXIaxB2P+XHCJTplDxfbLXwrYiX7IgNgCVDl9z9
4bT9RYoOJ0gbErWOepLmfIFyVTxXYIFbAO76UrIU3JB3D9fmsAy7ADWQQ/H9uEJp
500fkzDLnikmTQ0RakB3ObTA5DIe98JVhhHdF9y0FzLtQc/26/CV+ZXheQ/q0arF
+t8QKTkmZMGm831cy0e8Yj9IWVBwhxMWqjloMeyMlx3DpNLZUxR2sUdpjqgWamyy
SjLaBKwHZYH+Ab+dBFuYwWxo8ltpWKvPlALqlafqFE6ulclw2koLD/e/wu5KN8bV
Q7sMTNqoYnIV+ux8M30PnkU8GRoexSSuDxaeFf0LAtyl+GWZFUoFmpB+Bgs5t98e
NIR0yao21kzKLBMGAHzk+dXzH7gzMMWnWTNwP3Qro0EY2ko8OH9NuLh/Gd4l8niT
XLFpv8tPixLVhZR/g5vyh7dttR87kXVD4E7X3xznL2ln8uUWZJnBV0ZJUNr7Ve2J
rQDVBvRM/zK0mLBqEQ41+DyaU0+vYafXffXPXAYmEgPo1ccswKe9mXy+g1U3sxQT
qYQSMII4vcgeqOKhfjfdpgWNcHd1MgGzg2KvW6Oru6RXddCjvqZAE4p0iHvBqGDu
xDEg5D9ub+xXiNDoqKlMRWe8k+NrdaLPSxht6hTyy84sFSlQHoy1azFP9RtPWCMp
vXvWmr/drHGfRocoQ8P6jj7/twZ0R9VMI71DyQFe+jFKjUC/gXyS/9Zfkjcgi6fA
tFpCksy4GUoFygVHqk5OHj2OxxvVJYIT5NvdZfa2rlEW2ms9jrQZ6dCieEeSkyke
mW5FVqNWe/VRd3MAbvkyheXAmYhXrnkH0vZ5Ehwrw86WdJNrCfB+klLALYBeflpK
zWWxAbUdCliYbCc03lYBVNeQXDqYchB7f19imKHxX4uZfmbBw+N80Ws/MB9HDKyz
V2DyVce6iCgqYJuybmFQJtnyhSIeW+iXIeCLuWl+aUTeDb3cB0CLE0rYgRC50uoP
L/5oG6Lz4uChajcyjx4+OoEqBlSWKcDylP83uq8fQ9P7X8dibgZniviijjzGN2vY
PUudzxzPZ0w9CTHrAa+AVcGdb2MRHOsUJxxyI1JLhP4t8LhYZb4sxsvX0aWVQHXB
wAMu0BWgmFrjAsXawW1ZBQjCz41DIBcK1SZew6omJHB6Lw3zz7kcFRZoTsqmYoj2
fVTVyyBbmzxD2otwSNfwpce3Q5fU1rB7woDWTYTn+TWqTBqQWBPqBEYG/9ePicRd
BanIe94AtxNQCVeSu1XeYNneLq8lj3IR6odZygz2lgiiKwSWMR0I9/mDfvoTMmJM
Pisf9kJpXx/qu5FFXvxF7tEBRy8AGmFDNhIovzxwixB1uNDNIP9THa5moy0TFLs2
u1itFCSJTm7/a4bRev3dx9m0UtOP6bH7hzkkicwgFeTOQ57n79GB0p6amSGIO8PA
W/0CgYlCRvpT0oQMjxBsCtNKEHChhoaukSKCD7yuEjEjExfHFIOeNoYDtDLJEeFE
XNMJKzo7y6WAj6jfkWA4yaUD7l0fQryoods4CF8+IwVoGsrKozu8kebKgPiHjxj+
8p0wu45FFhGVUj62f02oBOgdUnw5EB/dbZSFLEgXqKU0KYiXhglYJuyOnKbHQb4F
hVTSK16d7UYR9d7loyGzYk+UYKXjL/9BCry13Vk7s1LgXOLDK6JYDQl5pEmUrUU1
+Tw3oCj2VKsogwp8YlgjV7IFVv0ChCxovD9kCi5czfwDFORAPSJCzTqG69L2wyyB
O4HBxPIUU2xK+MLUjsQv0318ZLm7TFNVhEQyk3v6JTHBKUqEaZlyoe4djv7N/8P3
3e7Aq0IAnzTJZLU/0pQwJNJYNQOBjOxq0143RSaITsioLzAWLLLRF/+TdHl9TrFi
fyWztZwSpCWW7k3bT+ybcp3zBZUnr3SEmMesrDEKQz8E65d61SJukQ0FVHWu+6dh
REMOrEN2CZUBGuf56xu0dqlERsloh52f+edSOZINxFFoUrUd33zDGS5ozTIPRkSW
6f+DLIgcC7P4/bGzQUNVbwykIJCIYJzLTSPcz2UGW1jfQ6dnv6Nk1uB9WXHMq1ks
0qivf83wcXc7KMk3zx78Sxv4AkfOKtZOrqcqMRfb/r1ffQjeVnjlu1gf/oKfakuJ
MwDrikXau7u2uozT96eS1/8i/iYrN6XHOkhH0NBtRFb6cmt6VT0ZNGE9ch/Lr+Yn
OaEylYwC4jVUy2uLaZpodGs7/LaEOw6M4QUvv5uTNhce/e7IdE8GBmilsllhePWh
py7sUoMaIfyCiAQghf9L1TlFoAg82bASICw8OMoSpqJypb2RoUnrEM/reNJ2LiMT
ez7zDz2c1GZvJRC0tl9re6Tg2KvMVvdUNCraPf7D6pxbx5Ij8Hn/FDXR1wCbii4m
kY0JXeLyDYNQxg8s+9yXTgbqwtz9Te9GemorVIytbk0rTL7/N6DhSvSXO7yGjAT8
FFek4P2/yUP4vJkj/qsf28Vb2KY4VRitYhl4uzTIkWWkLWtxI9DmqqRqBPti8Cf8
2JcGODiZViXfYUVuHEQgNag9hLQ9Vo9Dv9xPk7gd5FYl/1TNxtVlNOjE1/Qac1fo
eKSSX0fmQ3JJTT9mof39PpomEY3F9CMPD7bKBD/Kx1pl0dhFcGnp7geTARtLGtIu
4cJh2nJRBa9LQwvNkzOPyk8OEX0OJjbfc/XEA3SX1U1r+QySiY75+0zdq0mg1s9x
3cEJI7Y4M9CybcOGygK79bOj16hS8hQTvrAKpdyritx1fEpy8QFbDohDY1T5A33P
UO2BRHHtnAPoHF02176SwKTJNek0Tu3MEF5PyCVgjBXiSD9SjFe//i0pNI3Iqqe+
fQaKNtGxIrcSn7scCZ0kjAX/D/b6/lY+i14Vyw++JDTZAkmrkTFEmwmbxtIdnq8j
Pw77AvsX404WGPXD0rsrhEj7fAWSQ44wJtKZkiDufhiHXWMxsnD3gjIApk6aP3NJ
HqptoD7HZJswKzLB0pwyIy6GJA1gXxzvUjP8uLZGaIg2cqa5hThFumplx8Tr7kIH
IlFIYOreH32jgT8vLFQCFLnFxy3NXo01myzjdIQYsvK7aclI/E+TjHg/8kP2Jh5a
vO+PrzjYR9Wkl3dB0Um+YHMZikCRAmr5TbitrPXS3VsbegXp/2PVmisIoPS0kLVi
Lc64+VXlla8kdU1pYw/MaP0oDz0I99T42tnLk6HjII77GdweZ2GduK0jPzrtFv/h
EbHxnPhKE3m5zCsfdVCP6mQaZReJOYGBD6UMEhgsICtXtUFBUpDU0BSDLaNyjpCg
xzuh3YMRMtEgLjQR28qJ/tbgUlnQOlj0VLj28eoXyMWvibXDo7C2yF/ClTDunRYZ
Wel5p41PzCgJFFaYtiRLc590eT6t6VCHyFAuKjLRhV1jL/vK70+cfGt33z8tENLY
w2CmbkS10wDt9N77mto2oTL1wq6fvezhMFZFkjEnFTwdjdJsbBY7DhsLh0xbaLjg
N0MNGbvTiOqWVXsoC1nPkrB3A0hTbcwuUHAgr8IWqbAH4ldoIeqHsS9eqFxg87iQ
1wsSbV4mwAmGwsyNDd3LtuCro//cbMLuSDioB67LHyAl1SQS8kdcmECwm1fIzpK1
RLjyNzFYi2fuv/4ySebvgE59MY3Pd+f+6GfwEweUWfnEtHo2onZfPIL7u3YvMb+q
1B8RtYAzVSjKSnNCsq3KrFtSb2sEE15UGhu8/0gRA0j5f/9LAp7sbW1hRy27408y
hnIUB5zINwuqjHELUNf/VEJQHeo7NpQmX2LZuB5gpVd76R+U37hJBZ91ZkTQWKVa
Wdv5/6mjK+siDfL4AFSUXbu4976rScvZbNJVV+LpdiQAfCPgTyqkSapAk/bQeXfa
K0V5C4LfWd1zLcSIXbhDfk6B0M012DdodAbZlDlsnKIXC7FCJ3Qbqj6le9ed0g+c
sgmqVAXIfJ0I+/nwS0i6ru82ZN/0wP3iwrYpq1MuxeIs0DgUulNqUK9ph4VkiNPv
lS4zxM5rG0AkokggDFTwLm2MDBD+Mbow6yFna4nSyrgF/v0yDNTfVq41i6J/Jjo2
fBNKmdzsj6c53AYNKSPpQpiQDZAUrtzWt3DhrsJ29zhDMgMmROQmdnp07/ZgmUPr
3Zv5aEXXiW4VJxpTFTOiJJ9KdfWiV7be9RaYUSfM+SVy7MAQPr/w1Jkknm/K33Ey
2pWCyew49emVTC9MrQTqbFZJBKhwRG10tYAU4GU3uyFGUHsOCL3iryLOcp1yXYzJ
o0PG+tBDOLaMzw3Hcbi6wdcooOPYHQsIm4MICvwKQgze0+VVjV7l2CanD5SP0BYu
dYfKRj/GQDvEtPanPyeR6/RbxdSt8lQC7UG1o+f0PkMx8GRYhbkYpvupnFGJdHli
XQxqAL/KXZp5wm5faT2ee49hQrCBjf/CN1erK0kmgJdunG++bNUrjCV+6UyZNu30
R4uMOSBmS1jzJdxaG7b2noSi5cHbRvIEXYr5SMbb/H6pzl6rssUeTBEgeJiwAK6X
zXOqjcQhOEYktQXYVE4BIp//ckXgpuv38c9cU6O9LmwHnby+MDD6WNdrXgX3mCFw
lHAOZCAhB7GQTXhNTOA4+8QTMYV56HaZbNVcsVzP/wtaB4jr/xF4gYEZt2+FExTv
+HFPkGi4xo19SUFx1UZFiTaw3mmCTJ8dgVaplQwHzoFGCo6A7ndWXSHBIn4PRSQw
AfC2cvyKTsEGgE7F+rrXZz249x9inIHXFxo8zrLJUwA9SwvC7yDnrJBgdfsLr+7h
aZa+fXtvBjTOngZawC+3+bEobsEKNwDBDz93iL9/DFdX7LFYLJcu//RDi1AsqTP1
Xm3HJk37nB972sirHEvb85sZ0Khl1dlUEqrQQTMc4g15MtvbWkIp+WqI/YTBEIC3
e2G50xCZm3AbltLHW1w526gvcLjkrAuGTsPqqPmhUHEvyJcAH62Tah1vpvNzNp69
+Q8SbwN0tbibpiLeS00ARt4FNQd6gZTjNi8v2l7pDURuckfi252E8zF3X77fsW5y
Ftq21KhSEmG927++gPq1MqjL35UllX/ds82AlVhBAFy4tXxF8M8avIIOHOf11LfB
RjLiWMY4fA71xTpzyHwVCDfO0YiszsIGOseW3JgzB78xl+KfeqznXRAtWg4yBgVJ
UOgdQ4Iy9Z32f0OpUCX8BWPx9gaZHd3sOiQ3JA+z7CPT4NvkBuuTXfPhUcYrPXuZ
cV2a/9THJfKNSrxX3JT8Kb3mDdhrZ+U1UB+iu2Il9bGknWwLZg6T6wblUnFbvsjs
E0NJmcRLVdbHEdaQkPAWcx8YndJ+OfbOnfCmtMBg3NFXl4jI9D9nqZbjYsOPkxg9
zA7TocZl7pRhxR/QngfFutWCVhxG1UbmnaxKM15I1iz3tNZmRMW2/IDfejmTyLdA
wRNj7eKpkcZ5w/LyVACNFlrjdFDmBdj7lmNe3LNg3Zkip+bXpVr0SOu2E2gGJQ3C
B6zW1JfuX2P7eLX2Z1CWa9OFVgf9YxszovPB98raJiUn6pf4DnkNBZTSU4yuPKP1
qoEKKnsRW9hF90wwv1DN+HXbyqUfsqMAX+5GTDRURvxM8CN23Q0IDzH9Qt1SMQAt
AWG2CmqK/+ZXBEsDy3uAq6fu7+/1o9nwc0YzKfGDfL4juCWm0lIwyBncTR918/EE
VWse+xZGvxfpqxmteZRxcRMxXnYdn1e5QYryhDqA1lESRfJUUn5fCUKiPNHVJkBB
bSaG7O8fzmOsFmx1k0VWVd6jDO2wMIO6ZJEThAcKCPNqoCUDdNVmdIiNqHdKYa5c
g8Z1Q4QynDtFyBnUksMld8DAtd2+ekzxf0Aq9F+xPYEs2TIQoJOuQSFucahfcp3F
pHZG+dUjelxlU3o6dAgiTO+to0n06fVPZ+9n/rbhhoEEaSybj2KPaEr4HvZjGWGK
wzMJX0DeVId0yWA6hNrKwS+TIEcbPilIjPdsADNIJpjPi36WSVRn5yPzHL3KsoMy
2jOkSQLxqHdlQw49IrqwS2unJNRU0JavlmROP6pJQwXaoAZyFkphiPREXY6QGYjY
/XeiTqgz/2ierJltBzxyAL/89+octZAbVZxqm+oWPmTjEwEWyUQ6y1R4IIh5C4E1
OKLIr7/+blPu4dc0yWP7+YBFPrv9NM3rmksvWk1ezesGQwkeFzb2GdmvCXN3EbFj
iYGX1UHJnJTzE2ghC/1w4VW7iNjgvLE4VwJrtCxK0BkqscRtTjetqminxYxO0k9n
YpyJMxs9oI6EPnvtkeiax0ztDftcA3qFb24LWdwexqKiiHod74yE4eoTsE3j9nDu
O4n+QeeHyCMbg8dkjnXM+6a3IN0p583b0pxkzkQeIBlIJmFy7PPIljQZDzbtfHhN
WwMZFSfmKeCe3jFVM96qLq3zi5VnOLhju+dtPm7ci/gTPlBdD1ej0PRkZGCzKYir
c+hRS6R/611wKAwuFuZZ6hoosDxgUP8iruMkEd4IIhIlECoQ+HD9smUelMncURA1
LNjWMgG5wJpdk5Z8Rvlvx5TcfZndybxUTJjIBzyiW8TdBIEu9CSjk3O//82/2/DY
Ri8eZq2h2dzWIxuKIqVnkQLSPrEtx+Ukv1NY5VJX5/8M1tkrq7q2eWgZi6CfSscf
Ah+c/r3gWT1nbe+D7VqYn4/MfqBfP4LbcIY5ifIpYPkCmE7Wjm54Hc8GUFA1wJE/
LH8w6p7jh+jS0akFdc3iItLpyscYaPPkkkb0RnJani058hhPnrYseOxaSAVHdFLK
/MWqSpIyXK55wxEPUgXl34EnsoEL/huxn64H+jAIPhJr0PTsnnXLPs2wkQ7+4gWW
ZJzVAFgiLZP5ycb3dJaSfqxAiohVY57zZv/UvFZZqewUqOhsZn1xekKY4WU7iH8B
/VZqPHw4ymldHzninjbXRPhNl1eHU7wTRe0jNoK+YU0XeVKD3eOQ/sacb4UoqGQB
hdA2elOs4U1oXrZbNTtO21WbF42cmCptfJBEB4RQlI93qrTwddYAAPEnF4Cx6fDx
lg4QmdHg6NpLjA9JD8+ukugLYHtsI+sQn/dlWAJQeYKmKofr/e8oBPesQWpRFQyC
JS2lwZF/QBq+ug15HDTkd1ZqsIxPLow3t9vjx3ilJOiFzCxRi33J+wPJrTk7ln3r
+C6/34LBLboT+7AviQXTboe0FjAUSxQUaKPiHpP9nFk4toiHKfG5if372GDG57B8
A/Ac5nuBVwq690R+p1HSTJ0TiotHSUN0D0hhDuHy4KW9El6Ty5q/Ym71kzOD2Ybe
AJplqEJPwhGOuhSS031kXdCFidAOS3Aylgx1r+23E0h7mNC3cAPPpsEJ4FzrmuBS
wwhCOagQkJuFwgWgqTuvsavGoA01rSDSoEzr08Mwhm48ho6879XEJoB1zqIDP432
jcwESmlPKFa35sqQ0CZxHw6xRKgblrjLDnD/zIf79o6TAZ4j4DRGJBBpvVbY3SdQ
z1KeN3M4JPXsBCI8k2yBqL26BQsfREGzLuTj5ZZdW4zLYD89iUhUHgpDC82JAlAl
ncEGOrjVfhBF3zO/c0XvrkrjBHF5IOKkzYsdbCXNkCFE/Pk4s+solpW/fJR7zehU
JKYHHVwDBWRKGoM8yhtWPl/2APjE7h14hV1X14kzNXMbpgEmYMXFWLglhl+ysiOm
Or4gnWVRQPy167cizZyDplydKRgFyqVR3g+g74Q0+Lq/EC5jLkDcRdq2XlkJXQLn
/viFqdYP4kdXB6XYZdtdR8VUb3o5nxP4ED787LqGaEV4hj9+djAAYojP3f7BalJn
ygowubJjyNQjV7VSfr+KUmO6PIWaqtH6n43VMUbpCgYAAC4iSIhfd0kaJKFyYrHT
POp82TdpJMTtSVz1iIqV0wLNnlV9XjaN+NhNp/dT58zYXyjczKJcbcDqYS9kvldi
dCW0zkWQ846wCZY1j1xHuG8M/1LQaJb4eVwfeRkHujo0HQEYoStTpYVwBf7KmW9q
ZMwaPsAbezhbdcAjwrMlUV4he10GdR2e28Ph49FiniBFwCwp0GSfso4krdbgjb7C
f9hK/QVr4qhzC+bZ1r6i6fpIWXAxjOzOaU87VPVZ8xc/7mHEZie1HJB6Qeg/Ma3U
tFGGwRVessuVGo0XqQ+nl3PCOwD4Mb1sxv/cpYk9EFVIiPgYoQeHCXMTrLSxzbMU
oJQEE6ZJtgsC410nWjJ5i49RUkEFdflP2HfckoKUrbEJEf1lX7LHqt4F7qxoHFzl
0xbUlnel/Ks80FNmeS1xhQ0Ic2p6Uv0WX2MjQLyOibWiddSWZ3X/lPXgcM5FhH4U
BgQoM6sO7IgWNnLjDWhfqyC5O7MfmetNiARhdFLNeK3pB97OgXaO1YERFCvagZVT
2tQ1HAequPpGFtAWO9XfBkD2or5Wb3k80WZGqKETRpwvpr4u/UGt3YPi6paL0xJg
Jt6mptdfgoCCYIQ6/hWtrRxyR9wmFipCifZ+9GkmINWk2223HPCiiU+oK0wBl1Hd
+Dc91CO3H/loH6bQ39sESlAA74NOoW0hzVDYdAWdxKED3MpxWn6ZDZZCcI+XRoz9
x3RHTe2m/z8vC6HBMlCWdw0IP8doyGLArQB/tJ7QPC+kv5ohk7xYsrGFBlSKGxD4
hzYdHLIhnnJ57Q216TGWug3qVyd6AUHNjeKHRoVIRM2w4Vxu/DkAt6iBw9cuDnzM
og1WfE839GacQ/5kRYe6HBQh2zNbKbgKpcsUTPVgbDHlnuDtfNw1D7/SSTGLIDfL
bUmlJ0NNhqUX/94pitjDV+Bi32c9bEMOysWAh9EQ5IM5z2wGQ+Wr3P7s0g4l01a5
MhVmvfmXRtfeMPPHAtPgb835wIrrvjQtItlvaKispHV/FChXHntU7cvhAifQblse
ExBYNreqVz9trZghIGwiemtBkHb7o7lxDZaGyy95JmYPm+TInwB/KbG6JGu1t11c
OQZnPSfHK4A6TrtmX2PO72BhJ20jp6Qhq+7KfBg9WQ26yvuIpiVhH9w7Xi+pobXU
WjAGAuQW7DrwcgSzluo8kPPUsbmtdVfR+fG5iDLgSRkj+XklhuAPxtJJyHu2d0ZQ
z5exPvbXBQHK43B153ogu03uBSJhvyIj/1nrksdKv9R5vbeRvmhMrCLwDrPEbEc9
CCyehWwqL75CeJeyUGaCzGTxF+UCYG879xukoHnv/gQr4/YLCnIjtR7JGC7eHT8c
Dx5GLsHmtKHOZTilBVygdE9ePM8sqPIS5XSPpSQ07xbHNRHgVFoawPqk8bwBtZcK
qbVRlGB+8K4KNiDzc1OIQj7PoomnGa9+GxsIrqus7HYdyxDw001wS7TXrmeRNBBa
CcLdMu5sOffVR+KISYOMrIUdOpkiEOCWcNos6x39VeeNwvG2WajbkcxtMEfUuY5c
CtaFS2svf+gfqkSIIVC8gL6jSORvMncMYs0bmZ+N9gVztLfdxH9k4muLdHxyBFC+
pNivt5DWZQWBVUwJwQ0xcFAYV8pqjjzLf4jq48fiMmFHg8iYLhWCFSrbXIx4IQXS
4h4yvWbUHt1+hHnJgX76AG9dq5KvyblOAtSjcD2FCmN3RjgqHcK3fiuPavr4PJ30
YgSn+SbeZBdQkJwM/j5GDQv8rFNoClYZDzF5lUSVqwihq1/8qvVk6ao1Zny/uqTh
TNVc7ejYQ6/zFbGIvkzvMerWPlmJ/gZmNLjWxBYrHeqjwloTbO3MrfR2iHwTX8tP
wDvKla/rbgSukMUiyVtlD0giTOU8Sp8MdNfrfh9BHYCND5JA+cleR/Uv0vWSZQxA
Y580RpdNpbQnFP9QO7FeGXH1YKkCLC2T1aWrFG919/ghSZ0ylU4QmORau5cD7hOJ
KkwpLL6YtOQhqpGGrcvmvo5qEcHmvzV+3SdqXGmJ8NH1T2QlJ1Zx8vF8W8d3022/
XVpZcEQhvxvW8ZrsVgbHAt3zV+Fh/PrSGMS0o6cW7A5ZSYp7+zXHuFb8sbPNceqV
0SXJs1wM6QXLOBeeNSiW650apdVTZos/WrhYcSpEUZbVw5OhBVSu8SOH2CNxdjp+
2g3aZuizvzmLOECYsPfRF0vrBu5uGLHFhm5OObC7jIynpIEZj8cG6WJ50SCKAbyr
gPy5IO6SXCnm0WxEKzH1ONTAYiCExCyZsK9sYG28WwXrFZGCFmQuDw3Dj7j/2nt7
AHWp5S4cmItouHtAIk57c2aFtZ89J0sFd07wRZ02RlVKGt/zJma4T2PIuG6gHid2
Or9qkSAc95HUUv5PM1yP+gmuScBMKIQgB2dCzOU4wFdwI67yI524vl13lXfHhTtW
ACYKPUunTOgsauIXd+eySDz/Rl9H0xEL+xL8dqEZe8H6IaFXxlVYVwb4g8jiIFJP
R8VPTnDGYMgdBNk4YtEzPjGtamMILHHTEfpLEynvEc5ZltI9Nm+XPmLthYCUy39K
Oixg5Sah6p1tkfDV7HLFSyOZv7YxX5msEixdRBdNiSgwgGiMIytp2Y8AXWuUmCs+
qiso/EWC/g8Wwm+gew2ufQx1vgNCbU/+pous+ter9EwlxkeH9p2482ywRov/xvbq
E5tQB20EhkUzkWsVXD9KOWfDDJfTwm+eQMr1fWTs4iteDooT1flW3FOq15O930VG
xO7ZqY9B05qm50YIS0n52BCa/B2v9nHMGbiZ4DMLsADNv60026YzB0pFFq2XfwDi
laLGi/2qGobgPDmFXVA5wvcUYoF2ZOVH1ZasRJu235dIwolv6PQxIooWsezsnUU1
/WRUWVsGTbHwz4zJZE2BNvfoIMFhNGzI7vYUu1DQNkelGqotjpPDmapkFthceTwa
pxjOANoFDk7DLNnNGXjJ21k0Khl+K58VW5e3jhlyub/Ju8SIlpRef9sAdz5tJjlv
d9dxzbvBkLvkPDkBDcp0H0/LH7v+StG9HuWkvgJKbhp4UFA7jXHU2j45Azk4VuUf
LH6GHsX0Dueuym/oQ9Xhg9tk6akrB8T6UJ5S3Ss2o0xk+sgyBS5IcqRXbPO4WCJ6
mDe+PaKHKUib4Pi0SyADxeBRgfbWo23946QI2c6udOJk6XRX6eEnWovRoTLb2IaQ
WoqGN9oZxZAo+3hsPc0fo89+WeyS3tApHbEas2mzvKQM4TwJzZDbaqiqAJXq1AUD
yL37EFA4WVPF66BBI7XrO47j7LPSzqnC7povMzU2kzKx30dLUAnNI3e4CFFeaYP8
HittKc56tICJstyQNPH3+S4rNL0FI4RQnyKn1RDSgNsFZNY+HzQiA2EnKRwUAp6I
BX0L0pxorzeJ1BCL1IhjaZfk/n3oeQxAGGyWEb3mrH7ildoTyd1SeswNjObH1OsV
v9bUNn8PzI2Oc39bhgh7Ea4lUORzf3y5pAtGOx3X3ZUonCY8Fk/WKhJAiFyDJ487
LyuOiAQdvaYn0U2WhOWV2EQ8fLc/zy1xDBJmDWqpTe/LCMVIZLwZmXxVoMTF8GaJ
G8sm4GckZBLHsqzO1OxQJ1jMNby1lrFOsP4956zbj+rsReR7Py3qB9E99Rq5Jnrr
YYHfQR+qSGm1W5Lx5sszcTkOTCFFEdwjU6z4PhWqe8W2XswdFNbz9vZBqlAnGJoS
JxkSlAU0XN29Ka/itBUd9+z6rkRLtVP+f9dC84e43qclLM2lJJ4nUkqNmFKYy8j/
GTwd8irtc74EuWgvn0QafSvcKT5/TEUUhTGRgrjrKMZz6Su11PQjeql5TiTO+BcW
Xne0tuPXyTmuIll/5NdGK3s//xQlQrDoDklWg9oSnkf8fjTvTex7jsIt1dZ1jUEq
0sd0NkDlmQoLNT8f4T4VHk4yTPQwrigu3e49TmRaux49E+vRDT2dvwETRbo7s+rm
6JDy4IUM6SxIFlbljwzI2MmvKljqu7fmdJWz1ERfcZXo4sykz+Ah3l3GXMhyI9ik
s3TZkcNkB97pVadBOTMqXlE7qwSq3nroyvxSXv9TNdYmpeDKY1rBmhPeeP9LDoHh
pYMblNyRQ5IUGQ8y4HQAlOFP/RD1pCfEPTgE2C2q1Q7ZBTI0cpSOq2tkzNdaV14U
mAZvpJ10rzV76WlpSoTqUn4Ypl9m3u1vA+7BD97cYFsOvXbgWNGygg6rwH7XQkFO
JOiIgeOw/aNlodO+J6ZdwXh/M/asssFM4it1TidnnNjpTU0JhVX810FPb3uP0RG5
3E82hxVZIMyqP2k7IOjw69AJhtrswDGaosOjyUq0yTQh7J+lltH93zWZvRMrtqd0
9WM4OseTNP6/ok6W5nC+q1xid++iRikQh56asrRkSqtDxznQsKAHqXBdy/beUpUz
CyKs4oh2AXlf0JuSQiwf4fOKafay5C1aoQrZVDs1c56YVYvCcbdrCafUYqG6chab
s+AodlyhzkYTTT1QBIWrNXfmf6Wr3Tm7CMjT+XWyrrVdGJKm+0jNtwzF7Ua3ThEe
P7jhcjc+46xA/Ee4qqPasjPS0Ybj110rhE3qGFKXHdvZO93/FVf1O/93mqmKzBM4
S1a//7fonyWWZBu1DbuyeXWBftGlEeUwhYW8B0OIpDeXHxM+EXjFKA80pSiV92xQ
l07M1ykVJFSEnda7UFyIHWuYOk+akY0OfQ55jqCspFRNFTLvSVAlNZgwdBFRzeza
BAe9PGp/EkRk5SUbSqZxDIhc4R9mxkGeRlSRVJE5yDepAWzORFI4S+iiop/F8Vk8
mUNoTZa+JccBq392vNAVJOlmuBMBEx89DGhmUxn9hfbyZis4qgr0X+wuCe0j1iPF
OdD/GvwzmP1DUO1rHk7rdo+6f9Eskkg7n7m2SzcI8YhwiZhvOjFfTuAQdhyq9BPf
cxCPKrHYgqOqB+dAFoY+ngLL+j0fHaNWHjCc7O+8jzhJgQTTe5Dcsi6l0awfeUAz
F35k0cQD3prU4Gmyt8vHZezV64ENtAiqeqZUq9gr/mOB05iKyyCgNWNTEr4o1zgv
pJo93F9dUM6T/Wv16uzhrN6w7Q2G6wRUvgIU5xpXskUafo9C98Y8ekGD97+vX0mH
o95ICbb631mkFjtKDtt7r+QnmjM6//w4re12KmzMczVyeyJYGk3GtlDnZY9nKfFA
mCC/XAUm3LiP9Az/tZyB3NoinJP3weOZLmzbLyr6+QyscdiCQm/4OWHP/2EsDY8B
WqURYdPJVZkCd2AGC7TFzocPJ4DBWAEFqA/zrlR4ICnypP7/714I3hKWpyx2Jq1y
s5rYGYjGx1Fy3ib9Cztykcs8ZjeXB4v0PLBJK0xHiZyVWLnZ2N7fZu999v7/PT+0
x+FN1F7vtU+wMm+axlNE1eEqUgS5CEjsaLgge7PnNp0BdhJckqccL7AtcOqga1Ix
Gav9Yzn7zU7fUr6whSeJc5Qrxk7t+IWYrrkiEYJWAYBU+0k1xGOZ9D3kK2pEsm0k
XsNNE0ubjy7idOZBOLOoJ16UxpeZRt2uqQflrtWuRGWrufJzZCiByS135eyz0aJh
Ya5a3KqkejGAWD1uy4QKiOUErV6EV4+mi73c+84Vnxssw5rNfqRccbXsnv0AS9St
2PsfAWVb/7qjh49BE/HzxWdXsdfSRf2QiOprHB2ZZb12vlFYcGZIyOzb1sFiCRgV
BaHX1MzBOQYR7sZDqZfnBaUK/4Lzgwdnx497efd255YBbERUB/qEbi1jFDINuPN2
pzJjm1gscwkBs0reK9Qra3WhRlokLxTZngmYQlFNvaWrNyFrgSJ6TRWVykM+Pqnp
lBIr2oxYv/KlhNqJG1Q8GMzca0xRzh9JyXAIJqz0hK4GdMO1Q5WVXBUoOlSXDOw0
VlOUpXYeUetVnXTs6tS1HEtu0q+io6Fb8peQKUJNZpe9Ig376SISS89lhengMYKE
+WUHpyIdzdgQmYFFO2DlXk8ur0Y2iy8oCGwoVQm0691J5ozU6VpnmLcka0AYLXRG
lJ3S2apKPBjouUFHhmI7qlj5foeWyOobIud9Nhs7oLsewTjY9RnCshVmrG0GymEV
KyPhJPR0HmtOrvvGWkGhBJ9w11Md3QfbamZap/ZE3oilMxcB8JLYSq93ErOMWOJA
atTV8WXHq6IBeDnYRhOaAcXx/wrWL8qCtb6aepJyVapFMqlf8uepHmbSLf4tTiql
HznXBWR7QMsPy5xVjmyYeAX0goRu13A38qow9o4dOR1LATjYXlKmDoiwWGmSpNeF
CHrSEyIDtRvNRA0OK7mbLrlQr/aXrGYe21ai472eGPDQCEP2z/hiPvNiQ8mYznrt
EkzAELGt61s/JheQ3K95MMOiQD+qOhO/4ijcOgoHnJoOFatkkhCAYFZsLhwiALxt
+Ay3l+vwC8eJYxAXBAK0cJThv8OcJkbwRhxVFFsYq/TgSj3ICkXRotakVuz1Eu4/
tiSYNLKnyyVXT4D2ZRW4wT4Ft8pfj1TA4y+rHzfoKSSqFn63j0K+5qcCXDrWvMVh
ix6kUNN/uolFTH5CwEf4jZXEFsgzSRS5SO2i/kjljTU8G/P4lEIkABvSlXig+TlD
BswxsfryAx/BRnIU+SwRAjf66L6TaN0d6tfuzTRS3jZ9/8y7rpFf43WTvPK3wY2g
2/EF6TFfxUeEmEn9PpmkiFea0dRnxwjLkSWFwdxx9XT8VjZ8cmJHE2Jbwb3kv2rz
236mHmmS2xBaaCol7yo0EXcQP4VuwmR5M9QSnSA2Vzg63FSwgUkfywb/O00QRgrx
MOULOOMDd1JAIle7LHWZmQPyarumVAuptJJKp40DEMpFmWr5zIZXSGU39kqX11VO
eLte7Hx5f6on4Ac8dZA8OrVTUrMbHdtj84g0GyuRTSjjYd852Fa/WZoXWvyvflyh
yDnlhDrldTuuBmvX15lK/7BxkdpRXuRHtGwJHNlCAZkXdbqGNN4kMDBZrJIQup2F
SbpQBx4xYxO/YBe4iWJ1p3gWr501LqRp0XNl8HVZ7zMHp/qdNaCndgxTKrf3nkU4
V2anCCXThNWt64Y2J+j5/1j5fdl3F+k3n07qqiRuf8sSlHNETaimv/aAK1L3EDOU
UEEbCK3a33gyvj+jd4xzcnkKIVC03chEuEo/XoYIOGNa8OSZzUZlNd/GbkgxLJb3
9t/d+7sroLDHGuEIGzHgWCjdFnaoO3DpUQGs+AsUn9qo2FD+66pnz8y9QayQiMlx
L2C5PygNeWVo9SXsfTLQk2EjHiibzGL3MTJwXQErSP94tz5Bt5COmbast/qzLMTw
RxByomWbIpmtS6q7UCc/OgdJePQuKl2Gi8AZ7aHw4MTeKZjXxvg2HNL5wTAkJCC8
AAdIGfrZZNsmjGa8QX6WiXmABJmtydwJULZlkp2hhfnj5fDaOnfAs0owdh0OUarV
8jVjWNTi+mLw1lDWXa09cjmeO0uZ1o238P+Fqw2SK0DiOJSuYgFeHqFy2exn7z2E
Qfk6hiSu667jPR/kkaouacCXB9kslCv4zraHbMfXVkNwFSpvE8F2cYstj8VQchNr
H767+G56oTFi3fltV5L1o5zTWLZVfI+4OPoRJJrbzhaEM+FoZJLtZH0jIXuLjl5T
G6LGsDAB9BbESco+uh0gMdUy33bUEkGzyaxuDowpA6PSCRfw1GqV+YVosksDClUf
k0TEDTt5fEAeHGt0PAYfCX5sLFfzJ26B/pHX28t1us6MUVshs+dX9zYfS0oz9iPT
TMZrvXhfL4s/CdHiaypMBpkEP2NRCaLNVQBqjDArQ/YkS4SYw67kC4Y9EVEDyGSH
4V2ZKurC32XLI9NqfjE6BnJ+bm+i6GCjqj6LwgamUl/EV+J4Auz2lNKLlhxaXYFo
TmgUHHK/4sGA8yvk5UCU0m0jyGLBKkvPG0UO3+so+uWPcmN3ryAVXkac9r67DGBw
CpNf7eYxlKYF71Ozx1/wGEuirTchDl6sMUsQxNDldSPoYLdcnKnwev7c+XFWOdX7
Q2Cyv4P9PcLZdZgOhSrvlHwfoYBQD0x9ORDxMSGish4FpIMZ5pt6NorW519DOvFQ
K7fYHAVFTYvnCujw1+hRN3I2fgOxke2BfVV2f0PXM0LIRfFQNqBmpGFIa1AJBh+K
c9ualVwiu0zZYE6f4J+RUWDww8mFQ8xmK71b7YHbP7kmlt387181Db30cpGEJ6jg
3+sAof5B2kOMlLlCkg5HHL8C+oSAdzSi2krMsdKtRG/H179Ni4dSF1J8Jk5Z2v6Y
f3X/zmgu7uiaW5j6+Z8jei0Z82RdE8guy63gfZdm+hf7KMOE+K5R3N3oEhYEc16n
6J20CzGhwHuv8Wr1YG/WP3RubKl4fwwRMaUYHWO88ekQgLkC9iZqT8jZjWEfHXJ6
p3OIZGwmNPVcfUDbqkJ1uAqoCTBFbd4UxHyINKVIHOevPPLZlm0pLOjdNKCQwXPM
tDKKywubj+6zGFyqL0Hp4pHX0n1U/PJIdUocl3pEhwYUY9ccVAfrsQIORwwOgaky
ZvCAHnW7b/uaMZ+iQxLlAiuJANVN4jitwRI5xYIGYVZIvQSLJJbnmxBPdL05pi6c
ccKdE38r6ubgd6X6f06hgVfYJgdeNXtHHHvCyItzgfp/5gpnzwrLmxwSL1tD8a6d
NXAzbU8p5Hf3VpwMjeP87qm7F4jxZD72AbPqbJQUqEQU3n8GE4v7Wy3Ax1Rew0mr
YVWM996RJ2n7/y0bsaBovJ6CZCDOVmGEpynV+S3flLpXrbCUYNXOqUqC22W+DwZb
34//tUwo62nABiiyGKT+9nReZs2S9mkNBY++D9akhl1ybjKtwoZgUkFLiD1109Ke
opeYJSnZTxkfnuiKzr+MK7tPAKPMNyXyBHTlbjz4Hlto1d6AHdMGEHXdQnpLzP/G
xmublMismVYaXskk+NHZwcQ+/GEd8VAdKS7A0TL8eixF5/hTJ4ouvDz1I4IsKvOq
wZdQltaL9Jd1E5Qe2/m+njzegXK/KbBXZQk1DCWpGa95nA87kqwqB4Nbnjj4pBoI
hIdDs8v33RISe0LgKQi8OgqySlL5WcDu3HB6GfIQyUkfTD72BGA0lx36bnhu5yKO
/W5cj8eQ69nNiY9w/ngqD+I+x3i9yyX/6GuXetZT36FvQO1rwxL9O6IEqINooFgT
jEy6W+p3lfVcQnkZZUFNAsv+3RESYx/lZy5fbEItcwHcSj3R2aBgA+GnZYEDjT2E
3xQ49JylCH6vRu0uTvOAEZ+wGT4ISpMsHSVnM1s+5LjSwCjTqkzJwUiGgei2HbND
jYt+iXhVS4LBsMT73bZyzFPMs5/hCrQvE+WaBghISGHrF4e9rIG7YycbdAILkPjG
3Qi74ZR+SvX9c+7mV+Gu9MoADIkbpN3cv8pwROmynnEUxFsi37K3MDHCXFlWg8le
6djDJGXLUq1gy9p4puTKgTdFi2oooiAKfL9IIMJYP6PyYN+RqSeonlZWk2SsmGOy
ZCMLZPnuifNT2RaT8+HZvgBFHPtsSVVQFRsG5WXEFp4=
`protect END_PROTECTED
