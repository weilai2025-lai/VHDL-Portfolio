`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qk/kvhAzO/fG6B7S3XhIZl800JltWWKB69AxXxcErxOIySSPiHnK1M6OsUx2OJk
xgo28uheG3PzRo3dXa44hMlMGDcm2+BTBX54NfWs5TFtDKR7+F2jsI3c78eTKA1N
AssGg+5o/EueZfIkmBUl/MvVNUb05yPnBOICv4vouSeHDubO2uGeIy3gLCmyJYi/
Be5VjNoO6RdAoYm4KCI7cUWxWMkop5K9wtePyvz41OTRzhlrY38YPU8bXbUh/yAr
u6DgUzWB9tM1oqdjB8D5uRGM+86DSWikltHGWHC/F2/ygC3CYx0LySzuWXbCSPVh
d7AJEUGO6Fhr56V28/UehOKsAqL0YDIlzS9NjFrktxwxJ7xUDsDCS5j8Lj/zmlyS
e3NJi1yH+9et5Xf5EGvICeggRvtKnavhEoFDE9at+rE9j6iGOLytN1NmOb5S6ERR
xu9Fjs1su7FeH1GnBYndgyY4UWH7u8z0M1mJQ1JVqUp5V/SjViY+h5XncXkLMtf6
AkrNfS1HIY9mqXxVCVCWRgoWCYjZppPBP/0huPWhoMQflMowaDTlxwr68z2cJC+K
PU5WXFMkxkczZbpw24cQ4bO4KOapTj/ddYleRqQ05/2Z7qy84rR737yFV4Td5qlv
INI9ClFk6pDkq4PgaEvTnbb4vhxbI8RnekQj3hZ5pi63TmTZntlcPQ63iHEDpO9h
j5IfNqHSwOLjZHk5FXMulfbeUK2No1MBKBhZ7sjYHFaNGur66jecZZYx9f0jYjyo
mCmpXn3wYCzbRRDDPdNhdDi+kMrnyd47r5mBTpaNeHvw9u0mCfLeUrb+matrKW9R
gUDmzjrDV7LDmTdM+Y8mgmVaf3BYIcYO3bnV3lNY3QVe+Gmb6srsIxcEVxsuDGKk
/F5VYtNQ71voDGFFQD571WWa5AcS3SQM5ud7BwMJ3GbBOrANEMsH5wjgbPa/tIVk
RSZEwU/Jsr9jK7IiTk8k0EYlcXfp1gHkEjrjzGQ30u8osg0EwtM3T1g+JTJBIVkE
pC/j65aW8I2pPJnxmqIVmEti58Lurfci4DumJmWO/QGsnHTaUNCOGzrLaRqGL1SU
AiG+pz1Nw/GIRQdML1p2h16BWrEIpxrlwqUhf3tpuZxGKk4M5/cWWUArTFcMj0Ni
3AQndgttOI2JsQqKxYHZMFJV3aPeldiDXeK9qmaEnhgTdnh+PVBgOrI+6c41IQCz
CPb9jONIrX0fSXTTOmOIZUcmi0TCZdld0j8LGFwARgVa1D8FpwKbIKeQ/aHforaE
hCCk8KeEJBOzSGqI0MrzZJ3OSzrx3S7mTKL+r4E4ipRjscRIq3ta/QLlzWgkoCUb
s82f3UUb1i/CgrWK2cd+NI/0KNJkzsHiPGuLBTJlodIuki9BMYwrZZ0mqD5YxjId
lb+73jJwu9rr9TiThBrk7jdYZNOeavgQPRCxPVX4kNyFXdR5OQi3k4oiwgVWM9v8
kvsfPKI1BOPDjN4zxoUut7xCfEMQ2cUBR2domoFLd7ZhS/xFT1Y3s85RFefe4PPg
/OjMD5Ueh3ESLP2pVo4YLruxTkTnZePI5vOMCDQl/2HYy6qJd5miWf9QBLCsaMkv
TPA6G+cGGWzVwX/1qhk7yODAP2car7YqAiihqxnk/WJ6sP+hiPByEFYjq48PHtVg
df+u007ex8Gnbw4RpAku9oHvUkDCfcP0FKvTI01KtQRn5xD1rueYBgL5ECj8Qw5M
jU09WIcnGmX0OtXNEbiDXlUZJcKI4jgPOv3lzNtRA6rmQ5Cxfp7WCZVNuY+fu6VB
mhkoZuaON6A5q/Vnu1gt/AB8X4RZp4bJ4BT7kFmNWGrfogR8JyFOxkwaMjHzlGEP
6fmpTVTqwz+kytg4wfoetjzRhA9zDiy6QlsECYo7DeGLa67z+0jevFhfSfE8dOHe
XDtBJ1GTJNswmO2HVPzLi8zgUplei69i7F6t5SaJZ+NkhgFDPe0UtOZZKoQyZgIw
BXHXalkUSa7CiF0SZJAN8scGVcINpTYcxD1V3dRWKofLVVFZONfAENiEHCt7tYIi
5YBOjhshKFMiZR7KNccj0BM6UO3M9qzErJES1HU7cehLKTVGmpDzM+oG21mHRS8H
PsD8gLNiNkOeV3CFo+JM3CPAK5fUeYkD6/fC0OkRpgOpktdQ0d7sFRrKYStg1WqA
iHjj1gCalcsS1j3zHves3qVB3BWn/WiC/x0QFUVDW3gf9tokB3vXEymrNRS5MvkM
wb2C5eEtxFqOjA2a75hW1jj7u1wgdcIpD/2N9gPvxWBnCCYP9DU0vwXi3lVvgKGx
gkpn9lsPOlJX7tBIjwuqau0m8ZPMUx7TuOG1ColgbWO6+VmPVABH98bTPEMqHI/u
HrKst4qv9LwyUlemXQV/x7+B6i8pWODewPCgNpfN7sD6u8yb23nKOpU8Xkq3TpvZ
AH7gGcFJZ+ub87gKaTI/CxNNpdPw8swyA3SVc/LdGurqZuxzZvrRnF8WEN5a+maT
QKRbZYHy+jfIMtkNjGS+5GE3tjhu0sjqe5tyZyDXsaC552Lt0qCWUSxQuQonKoJ3
WcULI8Fd9ol3JdaLfoYImgE6m2LtclieUfFwWRtXXoCCvloS/MO4OJr0H3Ruva1R
JoWGvlfLI1GO/obuIAi1yocO/ikpLjqOQDXxXKxr82m7WQLHs733RLNr7KOH0/CH
xpKfizWCu4XIPfK7vu4zdFuJsDm+wuku++sYpUMClDn2YJpm9TN61JYONCY2dwBf
/rz3nmhS+wyoa1m6oPqCDzvmXhHYmBJ5tC1IYtNj5fk4sHW399OOyHW/nR4jo19S
iakdH82q6BSBr+o5iCgJHufAQvomFQHAwwpz7QnM0pN5VX+LSrBJU08ERhh7drgt
B5uCvy3BVqF4O9M4DRB/u0NJgZIWG+p8k13QZl89yOF40EMp/K5lqy1cpkFQsLVl
b6GE5uJu/Zb0twXTLuEyxiBnOx1W3Se6CnmyymKZguc7xqn7Ex2h7jCYjHRcequd
QOxS1SMYhagXmSurlDtDIJn3dzJrl0Hv9djn4M9P0yoxhz8HnsOmCtLJNMeoJTuo
GLpOKm6UMevaM1l6J/u+FZJu6pNE2AFgakCg0NC7uidq5W1VLAyISCUvjDVXb1Ar
WsHyf24Qg/LU8QOloxajRbXSOUWLODO2aFKNiTd9RDtn0jsheJ3Td8VlhKYYyBrf
v5xTn8/DmNZGTLXi/e2IVmDwMKcib6ZfLQL2HMnRvHlkpn6bDYM/+83my0tvg1Yh
bUDAuXilpZsL4ly5MDitt+ktG3VEM80sWeIqahKF4N1rLaeOoPmnilc23r51Lz35
l8wZ2UR7zZLYJIEy0nNbZ08DDBmn+uMfQFWX0m9QeFcW0tfUGVASyidCy55FDwQP
dvZIjbrfdQGOjtbW62GasUx08JbJgJTiBXOffBCR+SXaiuXFoIdE+gFAmL2kUvvt
ukGtnKaTJREKAxQNUqWTbmarXtEDEF2h//dOGQhtlw9JEvvYE0e//JiDEcqthm2W
Na21G5D8bGVmZdKoTeuZmdY6Za4A9LS7Zh+RKaZnjQSkbCavzwNfXXPZQF1stZhi
k/rOSIcno4W9TT57zR76skJLCzR6030wc1axRI3steDwHGSoPBgBSwZNmmMwtttV
gDqBXy/nuinOxvXTBusSLRa4/dwpZIuXLKc+YLMAZEz9ygpWBrTqxMI4UC0fgbvW
Rr4T9d9kN7OAQ4NJ3vzr3qphJ15dMVeyDVyYzXRXRJ96S/lB3J43P60A297McvHj
vnflTbXgzD5DUL6TKAxN0EQGu18TW95Tm6OLThuIr/zpvyCLlnVohOLByBCycx6S
gbduiu4hAZF+uUUCzGJ4Dp6iIGbnc7Tet+CXwwlBGAOi8f/9GUxrq5ksDjrlIkYN
IN+yxDfcTDukX4zixiVvvN6U2fDmHaQ6n4LdsyZwSNqkPFtFqUxqtJoZ7bcGn+0R
/KBtaE3BBLWMtGWEMkPVOJKsL5+nd02zebWV/fdw90tKtigjH8myvskn1O0ZNDSd
jyqqTafn2s4JJ5M+l5cs9hAMOJf85ViwXqFlfUZ1h3VkwjdInw49J1JIugyrjy3N
Mx6M6KXFB272TTy6YNA69+lW7uG7wFlWwrYUZGL/kAuLlx1oOHyi2CCHFlezFBxi
xryhUxI6hqrLiUHDD1Spg53Uy6EG4AHfxKTShTvgwIexqAse3FS12e51ZPgoTKWh
I2n50LqBC38u5A8ASZCrC8Y0+IJqX2pArv6kxnFawGZxRJbUUJBO9qhe6iNPilr6
o+QlwUhJd8vTS2GdbLUCmJ1q1Lk8r/Zt6w1VbAOjQdDKsI3uEGAlFLkGtEQEXGNF
o8b+05pie8hqECh9wrlnOpYuco9RVcKNxeQngvI7SJx1NCrW2+hSIeiaTve/oIAE
Mn18VgqX5712kjnttTnSNacURVmwntzD9U1Wx9RqoaU0FYnDePYbmZoICBYghuan
p5gNk2UWMY3B4z3FUt+37XwxH9E045weE7Duw6AP9hNpGXu+MpAjeqQMhtXjS2qE
M1FqryuqJL5gkIhJXg1OOKdM4PYYrA4bXpxaqmTIyt24l+uuZkX8+Lt5D1uRPrmp
eRoYwVaUi//LasAvnTVdk0tAAU/rKxkm+LO/xQrQ186QFpJnFT274bLM7TIVBhF0
DBCj7bza5z6ZEhvn+w+JvMFiVgUwVy8acXejFXmvxYAXi7mQggdCCZdTirVAc1pd
FfNxLPVOLO4BZGz19hACSUttlq3BEHLb8c5mWdnZJDshf95Avj+YhpQc3eGuqZIG
EAzT2prBvnwcOhe7Mkj1kBv+EGWuRknoZpiDZgTJqfG/23QxWt+K+VJj7D7BNad8
8c8IcbttWFCRQJjzoBhuEwkDQoW9v3BZaPwmL4gTl/bdEjBFiCdRP+DD31+8r3mv
K+MWg7ekDuDaUJEQ2uFUNUKzAj7AkWcnb78XBVMzvKR6mYJgzqKVMvrsZvmz9VrP
nfzfybEq8o99LSs6iM5gzXon/3/BRcH/NvoKTZJb5p2TQnMbSd3iTvFYNfW8PTIG
TFaiuRXG7d4ZIewiHbCbEW7a2dKCLO/ZT0q7shqv7UnOUCjde0hvtPMfvIFS6oFu
rNgz6sbly2ftbbXCTmiE4AMghFvd4HyvnMoMyZLB8Cok7Ll4FZhnqI/3AXrh5lgR
nHLwC9oaP0J2sZ95IR6RIpEzd83I81S+NEwtCq/FUBPMn6/aWSt9NAIClWuQ23wk
47BqNOehnzXZD/q69tVQLVhIcrZ3hoLA5Typb+B+V7GSoCecSdoXZjS2t3QpMTbu
M9O8WupssGXu33BDixlwSmw/YQbxSxeoyWJetXj661AzbA7PTyJAbKsIfT3vQ3U0
eXOfy6R7iF7nHrZHdTq9oVQoxR0E2ZxqtcXjz+y7cJz4iwVlsz5Qn1q0PKO98P5w
l97cBd+ukLtxJIRjDqqgvkyloXuG8VSvjxEEUSDL5CbquiPui8oxiHcIynVPqVb+
amIekfyQKcUPwLW4g9sALepiMp4jgH7SUpnQMD01+O6h3BN3g6mkPeo1ucKM65/4
51R5gEiA0tgeV5mV+f/ZINDqVBOrkOXMbrcdIbKq+wktwNxWBLe3bKqShyRI3ANN
lKK2WH5/7KCVWXIk5Vn0o73y0EvV8Gymya17EHVqjdtfTNlC4p2bH2mVqsVMtUcs
8/TiKRmw2OriWNRfPdLeMiT0dYlqgByAZCqQnJMFF7CF+CE4M3pUrezbmh5ywOBH
xV7KKSM3HYrupMCXjfoDMmGT35LtqsDEb2IFqrR1inSbza77S11BUX/+RNO4Plyy
cXc3sMWlftFndouGK92ZUWjNsLLUbJ7er+1gDgEXo1hKZn1LDJv+lfHeAEgsCNMy
kMEkoUX9w6Dj2XCp0nMZ2KUPqb0uWP781iN52rNCPbinJOhcRZtw5vJt5GalpLiL
u+ss/oSOCyn302I9e6hrspS9jMOgAvoH1qjwGdYvQe+tNElv/lXkxdMtJ74/W3zy
b1JwsXhyZcY3LDpQqwhk/iJVJt8U5e3rpVnUsVap/yVDEjl+segWJvP8VkHqCTHj
graCp8ZtguKDU7QOs6spsgbF+Lu+noayh2krk+00IATGoAsPLKFkDIkWQQ7SFeIj
F+dGcSCYC5BR9fx/uYYcFHb6qdZkGV9Gi0yedl/XNcUrCrPbqeFd1le2+yg6DyD9
kizDUVPr3ReifqsoCb6L78FXmvu2MgQTGwgLQafDmKmlz8ZFwsQPCDWTk+HAso2A
f1pKfXJVcxeqHON5GQsAeODQrgBT4B2WzZrPSgJFFfOzAHGRGxFq1Plm6h2W2GVg
ub+ouAPSGe9Vle4kVwtBf6SpMtAD/4dE9KsFuoqiHLlKTLLRXz7HkyGwqBu0QahU
ZshMp+xifPSEGxt3JJNgOzxbN/E8LnPrGhtZuDDJHCso0Bvuxk80cP2lEPoe1NNV
nf0weLYNc5m9oWQjbKTNG/IS6fXM0sqilluiuIHMmqabi6ABicSqv0MSoU0cMTUa
jMMqEPMrWc2r6tetVIktuXcqBmMdRWaPBqEa/+80wZUmCTNhCumBH14cK3Ti4weu
Wl10b0Ae8oczlRN65YKRhFAAjopBQOlnnmfl0ewxidc8lGZPDVTXCTfkmy6Wv+4B
sVK0dfSWhDrrzPdINubBaYajNzkICML1Fgwjq9YPAYUR0yURuytRLNoBmHH+tSIj
plwEy9TDoiDGggQvblkV459g1cG+kXjKbDARFR+rbC0+KWkvqPo/HLIYQJmMuz9q
6gUA7vWS4HtWO4naO0F8Mg1LM9Kh35Tgrthi+d3W2bBB+iAEv9xVBdKiHviBuiYF
eCMXQqMrGS0PJabWFXlKu83OUt/OMRD1eNuS9mHyZjF0Vfx2FwArP22kAytU8C2y
fIgOINBZ9sWKU75oCWXT3awPAYnaJClS7t6/ZoCXnp79/aBqbr0Q3VxFMrRuPME6
vLsA4MbWxX0R4MT0fLKHLDEt9m3+igdn4ghOarjYEGvO7G16GNpO3D2+MB8wZS++
Ef5EgR1AKK6QrEEA4mB7wAARXYXfl+uUV0C1vlFH3NWGr3Dml8ga8hjBKp1O4I6M
7CURNh3EdzuaknenL4ZxCcpIM18RavQz1dxBxUEEwt/vX4354tD5Rby58azdzwHQ
dlzmo1tCmE64ErvWUYCNdrAb+c7eihpUYQYKT81k/I60UCm3iFwuJtnBF/KZP0ab
zjH9G8l/aMi1MDmRfwBAkC6/dXueS50hIPxrkEtzn5dw8mJjADJSzkLIcoCRivK/
ZjmknvJXR5NAvVlA+mEP0w==
`protect END_PROTECTED
