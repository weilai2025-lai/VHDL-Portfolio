`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qbblzz6ddk+4wvIMaosfDng3ZMwyeFLgClEMIjrDiLbd7rScr8XGxxj2KgAWcFB
5hGz0dWPR/SdjgvdU/OCKO76l9/ndgvHImdjdZb6q8JwkUqtP3jYo14aQYLjZATh
uOT1dtUp/On0DOSygteHrXkbUFdS4/VKRjirM5+4WzAaFCi1BvqzhQILF3RW87RS
SzDxyBDsKPzFxCXaG5DjruUIp2T6LDLSWJSpBzoYnNgmjvDHynMzSjN9Lej02hdv
jnNlrIYvTcSsRCwqBwYbvWFw9w/BR5hXIola16ZBIvwLYRWJe3VUXQDG8cIiXR+5
LVTbGGNm8Xyt18WxEio5X+uvPg4rhfy6yFQhfAYPLnxUO3WmI5PL9gpQwu4vs9pv
OULc5Uov4a4AjksBYrv8uQRFe3yNHZTC2JMOUyZ3JnSiOt/s9cP6mpDu2W1MzVPL
8H09XGteJh1vJ082tNOCYG8rGqQj0Qfc9S173hYk5UNeY9UgzhJZsaUOFAa3U/N7
VPBdryM818kLHn3BkS6tuzKLVFEJpiqLPwDKcyauvVK6/6SoBm03EQDMxX93ZaH5
e9PJV3q+TbBmyqJLyXfStr4SPoKElJz0nSX3BrG1Px/RmYCD9Wc4fwRY/OkFR7/u
yBMurMuenDerf93xAme+d3NMQARIilbXbcrbZcmngkwfWLv+XTHm/nOUsLeTa9Td
UaV/58RjkEh7eOwzdqBvq6sexfQo+NMjziT+FqmsnZaer1xkYSwQmaHdeLDrbjfV
/uQPPWJQUF6KlFkJffCDaWe3/qM7VWInm35qolRpn9lD6DNliHrlPO2eg4VgeD9Q
m9JeykmZdoJYUAJOhAg8HnV+6YImugXvnkH9AIQ8zA8dbSqlMTQ30qIlt7HYYeva
QV91bTlWNlMt43iqihvmqM0xc+mkHD/XKpGdHc1xTlF6loL93mIvUtb/E/zzy997
F5mZDNRZ9n6tui4VxO7HXOF5z6JMR6q1pF+xtN1xHWDMOVAULjtwiyj83IqjrGaP
ssN4/QFXlS4HCEE1iiBsErZ2y8UsWBH/U0tE1xLzB7h6n3BGvFGvJKk91Cb2WSRR
hVHSaMhHihEJeGp8rodVKrqscaAWGdfzy4En1o7mSLfQkQJ6VeBmPahPxwMLB0F3
BI3P6BqTq1GJLsbyjihLRtZ+T5a4CyaTOCvaewY7HV+yBesZrpQTMAWt/CWVm2hr
6PbBCQf4DRZL0843QEygK56Vw+Zv1qO+RpTMkaqEvaK18BEJw+wFrwQyMsN05E4t
+43H26pUPAWH3SZaqzxRaZrLEAjHOzJCP9oJ8v4KLX5QATv3nq5Yx5/zZpY2UpIg
CYkuzo4ZqpUOeakHbAocNNzHEYWqkkvH3yvNILG80Zn70A72Vg9hQ+VqUw3mTtmz
HoFpeeVp4ThqBeqF9pJGpxorAfFGjQ9qI8WwVhl2ImmoSMwZ0D8DbYjMU8nNNBFG
XX298/Jf43t9JTRrXiMKteKC0CL5fq4tJxO9owg+WqvuuOYWA03YG1t5ZKZtUknw
TGZ5nlxNy8palbbAufGhpPIuyiYZKbBXaDh/01Imy28atqt4k9xSJMCQ98iNcDkq
PhrrTAHCkDw4p7lb3HZ8h2TCErl51zDdknLvSz3yYRrcUbxeKOfLTu5srkHdp4Nz
MBvtANqesg8x1pnitJmQjnWEvu7f7llESRQ2gTXdqUQCkrklYzGiccLOp8JWN6/p
8GDnYyPpJYiSk+CwbhnmCvRH/pRWVtP6OaKOCGq16b9HXI4a0wMGRem3GotZb8op
A9vhdJflwGwMpKAP0vWqq4Q/5GZeee90N21mH+BPeoifAJbZ0Myqy47ln8ADs34I
Hy8mlG6RfFMGd/jr1WaLXGveamV3vhoqq6pnS1OCDVhNtB1tsFRW+Wvcm4yKzCUW
fb4w1s5TrsHOrVYBXdgXhOvlqW9po05Sja5GuqS3iRSoLB51l+0dgS76CtljzQs5
Dr8qwaJIxIRK0TOkBOU6xbRphYzPXbnTWYFozIyMQclr51IPAnCD/gJ58hl9t0eO
5c6rnjrJe2M6UEvnlPfOsE1vZSchaG6m94m4Ikh//K5bt2tw2njmcymyAMyBj27P
GsI8W+gPRMnbmVUOJoqL0lQKdHiAEB9mO5lgXfhJLLYU1jtInrn6AJ1vXCssirp8
iNtU+bi/Vkcb2Jpc4objGG4zotwdf66WVa8NUaXr3/hJmjy/aVSOlCmZoWKOFXxV
SpzRXC4APhOY9Y6UmH1hf6Q6XO7hh2YAisSRxDpnuWt4JbZIzUDnhr1pc0Tw9TZ0
Idns+f6vogexWj+S0/WBx1ChoPOFpa29yKMpEKXez6NhF5sn+DbtRv08dmFKko6S
mQ36uASS6zJMCJfPF/Nu0TSrVQGoP/NTL/jhlYBRPA3C/I7wbLpuLUy36PSa20NG
KOYn3GFEuAb/n5D4bnSCsGI4L7YlUgPg9g68j/cWfAGFmy0Fyr8g+d+qHyS8mzC8
/xy4nn+kcvoTgaycbhWmqOVTdFL+P/+InHkw58HLXczb+gs7pjgULASpF5cxtHlN
srFrUuZmSaMjbK4DFoxoZFyRG8p6Z3kUoIcShXYqnaAO3KqAIle73545oS4MD/1y
J4ZgufWA7zKxUtVwnUrVMqG9QO3+GANrtAPronaKVh/05h41xpVAhqYVfp3hbggc
huOaCVmsZJ0sM0DWd/90enQC3qJCERz4az9AqYFAbkGMFmaHEh2wWzr53qzkbENQ
afTAoHWQQhd4nJ8xDqI4uNmeCDTYr03wlTpBg+MZoJyKGBffknLxBmv9qyoymzkh
7OYDh09HA992tGSzBmvxpqXG3RhYF6XB34DFkR2z9QOM2TD9rDuQG53KCW4tU9Hz
ULKuhfR6Mdn1s8uaW/yRQ9BVTXYxE8xT4fApeEm6oMWFY74lDtiU2yw5mdetEAbZ
K3SWXQsVgQ828uKxeYCQ0KrL63kUByajlnQAp4jIqqY2sKnjJ/yM4E0PdB5NkmGz
YX/HUcDWialWHTxh0TBvAIKFEG8r54FEeF6OAMgxWbBi7NxqJBgkSp9PYiFiOPA+
JsgjoRFP9/XNfHm1h9ANRwEFqjxpQxGssG0+IpT53NgovABpZmBl1FlGD2XMcUuW
eS9aqZE30p1RJBUoknae5mi5d1lQ8ECj2qC7DLxHj2Lri/eOHI6rMxT3H2k5Reyo
9ps19zCHJ99GnEtikYv/YCZGPseGGBquhfFLF+Ku3bZDfIxfkCaBFvPi7+vZL6hW
kr87vzTEdgTPL6JrR2RqfeHHST/9Dn0VVnv0wSX7Yr16WwlwAeKxEUONwhKUJ1FD
ksRAIjD2ncsBkOcJ5cYbuvWA0GyaWEr55zgOkxwyMlHjOiWYMXKg30Twceu5Po85
bljlpeGEFHEx3qW8TbirJdOdS1SmNJoBTgeIMgtYhTqF0/PLYGmIu947v5hNElM3
ty1dEChHCie9P+PD/EcgCQu3ps+FihooyDbcIPiR8WcAkZR/yHNlu11ktOpnV3Pz
/GhPaiiKB7rONuEvCRlrzA7i8AOZjSYWaw3yEeBkxoHsR26t4NWSJQMjUP2I70bL
QfniXB2ofiTlYb7mjWI1rxEOFY5AR5JDECRLe5CzvB98TDNLn7Oxp66bZ2IU1H0P
eZHhgvcIPcQFPns22MRVC69L1OSlWQFTaEsm592/gxFVaJFlxxhda26Q/PoGcafz
yYoyg+iYFUd9yvGXiv+BQ1Eh/Ncqa8+TrNKmcifW39TSpWSxT2hmnY1nQmsK6gx1
ZAcwqkgA83MRO9VOcktxxIzLAtU767BQhgvf48DAeJObrBARCTmeynSyiP1hpBVT
KocP3qvJrIdds9rT2UCIHjEVwo64VMSY+h1ZOO4Cro7Xeq9LPCKBPFuf8hsxqd47
soNgDhifQjRbJYJFyqtw73Sq8ZvEL0q1o1781L6immTIqZ9JpeglY/Ab6y5+/t48
eOlw2hdZSn+3e+X1ggVU4fIJyfmIx9Wtz1XjpYBRYGI5/a5c6NZHhgXZBx4w0joj
5vkJEJJqGV/Pbohd6v1fvfqvJDNGUNZXkR88YvOKmmyllrXq6XOKsNzDf2VlzJye
LBemkF+92PVtqjXK7Xs+Uxt3zUX+TLhhi4lRqvXOcX4Lo8j/G+neILlzpv/Sdug4
H9hO1/Oyq4TFdwgL//6zrpMRe6dQ4AMhYjtYnt1sJRsiwLQMx0HvFIwGex8xDb45
bMRkR3TpQLhismJ0QAZalfxTbOurb6C0ZfOD0r0LVqUQtoyJtyIxYCfd4B9Pyb6C
+SmuDfduT6HdhTq0SR44E0Mde3SCR4oomf3FaQxUR8mO+U4GXI/bcrbfX4WCav/G
gvN2DHYvju1/QFEXBilTWv5h+tLjmu8wM1ORRBL3TsYqrmoHUDdwegHzEnMUYVWh
u+rE4Bx4QNyUFpETaHFqwWe2P9saLCgmaBQfGTV4bRNGrfzgwbce4807pyavhrDB
wcCEhnP3ZmnnG5OFj2dyRr+rYdIdaCEPG4lex69vh+PxLbp1bMBl/Ooef2ohe8RP
V8IkhdEhg43Chf30vIK2oHGVfc6AekXxiVBF/HFFAEDeGRGgPIbn8F4EYaG9xkZz
iVMtkrEyy4TEAQwNUbiPLxiyuy8epGCnxs2855wr98jg+2lgSp12cV5hsFpaTOih
Hy4X8XtMAOY2RcRCf5hf4lDlIKvc/2ClkuqnmTcLrH+Qt2Q+K6RUlFPav/EP2pEo
InJqi0Y9s5iOJm/UPYfIv0xka6ZVYNaiX7fcDrwObY7yiIWuSgnBdVoyeIC1uRbp
4bNYbDSEni7DWMgWKQalokmdApYxEEI5rIjlyqy3lMxw/2upd5lZZvJPHzDybD3C
x+xmeKqJ7nvKjfb7TjImco/uSlSw8Q2wyCr6AXnVHHZnUlRlbhzy82xtzrNXJ8gr
ib9HmWtp9jOSBb5tT5hTTv+a5GnZV2krr4vvqwvDBx8x31MofE3DDe056/asDa14
PEJlsiDzfaaJ+iKMQuHqrL1F1SX933ZzE1ruua5GGh4ybKFrT5N6SMbw8OxV/dhm
ZofVTzM47lgotKDiDhvuyjXN8ToRY97WpWsQZp7sqfmHROma2VPdB+HlymX6fY5i
1UFn/WhCPJLbPUCrW6trQVDdlAo4R7L91r/MaNC0mlEQfXHqMYjStWkvfZqewlHl
F28aQLtW5lIYPXzF925LfY0DrHd0URIP/3dpEBMWcaRXXsz3NP3gysbuNoXKQ/9E
wOqqQ1V1UplsJZ1XMyqCWJFRiC/SEEg3/5giCinuAha+Mf889iXBZljDjitKWZUp
mjlR+42fhHRMc8/LRAWI6u+6vFcU9rddgnBXubhRDNNDdIJx7X2Dkn2edIG0T/PE
C2h/TsPqlPvkGjBFWpA8S2I6Iyg/eRUu984fGHEJhQJrCjaYssfCy5Diy8MQWuhd
bSreO6p+78XJrTToRxaMEzg20ebBfBhqxHIq8k6CxXnm5V97Gj6jSTyiJHLW9KvQ
LCcwMCoBbYupZiAYJsoFklDMBMamI3DAChS68wceTbGua0UlFd2RSZEmEPnDBUmN
etx+pi9WLCLtcGwL1btAyB04Kuv+ETzdFe4kZ3qydpY+q8Guis4uNuCQujP70yLw
UutLx6s5GFIH7CsHrcwmtI32ZoY4JV/Pr6bqYG7lh0M8/84Ge4vEfqJqVpP9+5QU
1AT85NA91JjjeTfk2j7U9aTZ0gfLGxBlDxXrCRfBsPI1eDbf02nbq/c33aDXs54c
UFltM73YTm/KJRLKl0nfUm968vo9HtZaryTbPy/9SZfR2O76VABjiMvR6tuZ+9Vd
eWMnEX1NqPNxk/y4mq6UvIKqbPQnTbfqptgo9/MzIaRUQdUBt/KK426J6H9gR018
Vu5vlzDMgSqS1K+mWD9Aw13UX850zTjoygNLNW0TBc8fn8RimaHUeA8HRl2DF/lK
Fq2xnxw95Yb5wfu64LzNLM33czVos5qqKmcFjLSHWF/t3TMTJff7zsDeQ0KgBNGg
Lp5Vk3FvwEipnBU3/LS6tRfmALl+AtPEcT+E/maIb7NgaZeZxqjhjZcElI85Jk1E
8WVPcDvcN/rU7gZa1UFnSwcfCnrbicwdKvv1IxAS1KpeIAu8Y1bC1SBwu1LhUMQC
iXa9mE0KhNpCu76r16QDETc342pGYEkG45AOYFUwZhLSdQavmAS38ZrCIdnHwLnr
x0UL/arXRoTXCDeF54h/b7GxKQst0pM6gOBFh6oqsYqIJOpVtEfeRqej8y4X8ae0
cTsudoXnigKv3QOLLnRN2z7Sls+Wwq9+v9AFHJKfpRLZWkMillQXvzIHuU/1zFCM
Dt5Z03o88rHYIpl4MO3ZbF1ts7cOLyF/9eXtUnC3FcKDpIYa5zqZj1bkw9QPRDb/
1zDk7vXNjDIYaTXdWeZ7vm+0dPdp5CZJIIwJJic/WNiYYSNcMfuCoAbd0KsxT9CO
ARLn6mIq66BXSZGksL9+3xq80TbtAySVLyi302R28Y6DCkeMDHNnAmCmBWBHmwf6
IL9DtBnDK0CNEc5DybnOlBKj6BfKjdhzkzyeR/uHm4l/detLJisV2e7zlzzghDJq
JiENRctqOwjvUHhgK1eEUOV14GGfo014LT1avuMWZ3JjhrJJRdIfcaNrnQGsjpgW
`protect END_PROTECTED
