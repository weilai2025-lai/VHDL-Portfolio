`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
popFQKvQFglqzFtvGSG7SSK+EFFdLWt/qGszqikH5enPvG877E8ei01cbZn2Ragv
pK9JhClkifESWQfsLtsc+EeZ2RoISn0GWC0jwtDnxaaT/+Ds2maxWwzdDR7UWFLP
QKjp8qB+x4WELRUqOKGe6iJWI0aqE0PYfa429LFUbETS9tTOtvIHMZG69yA5dfBQ
cFTMi/wGlNaaf7KpXUmPh39AS+D3LIrVv9OH5cjUEWd0BwdvahesGSnAxGNUw4VN
tEWjBvF2Kdp0vciwRje0pHi1z/+x8VLFYt9CVWYrEl1BiS2Xy5N/N1mEcQ+dN1zH
LZNGAHvfgd3j4iumiFssfSbT47nz9qw68/+MipldHuqzVIaC+HqirAPzwci+EfyL
Y3bHy+rlty/wj0g/m4SkIuFB+ebssXrRILTdmLcAI1j4+XRBWWeg2u9oWJ6P7IBI
El9MF+GTIF0e3oPcRNAFeDmfxM6MbNzVccE45RmROhnfNDcSao0BOJAWELx/L+p6
J6kUhfpy2+8vG0J/+NHQUxIMbTImI/4HgGoywpoBk7oSC3O2ktgwo873KXzSR2FO
pAuSsFZWJeN8cVGc8nQzMOd5yxsdXWyxsRKwr82pC3rGsZkOdqVQf1hF8MXMKBO8
i8PqWlZanRlRGGdH0qcZXKqyUbz35odTPJSC9eDWA+Tp+2rq3Nl4bMa41AqXKsIN
BjQyBIbgtaPl5rOS0YDSM6Y/WZcvzW/s2Nh77Ag2u+RmEdNgmzdGXcLALAxnrgO/
5UpRN0i5/AcCDoyV9AKU9/SXFRVt05d0pDUUQUN/hjnZD7JgWOXdAiSIdyoiB8qx
wDj0pyLiQ6vNoP2y0doX2XafmAmK4gTUfQvolPe6qhGd7YK7Hp/7QMWIwliXHaGM
cT+mILIQmj2C7U6jZe+41o9Yx+jwdwjOVqQKDlZRYKoH12Pbqe7MkYcd/gPR9yvV
LjAgqWEn1tHjQm5jc4XTy0CvurKkBmzd51auKvs+J30lflx5AwxwRhGyxrf4MVLl
DOyH5pffhnZlkhUonUF+cC+I0WDzIPGQCM+MjbIn3MLbd1YRWni1AwKELFha1Dfm
asYhH33uVndRQjoxAbNbkVNzjFk5Pj0S0zOY6stF6hVZRINfD8O9eo7jRdEOF8sR
QDOLR661D1ic5XJSo22BdIVYNbc5pPUfiih0q3QoGfSkXbSzZuL8HwagX4yO04my
BS983haS9lsDI50RTlQs3hoXJW8NRy31P8mGgq/vL2kPS0HeYBtS6Y9jFB+oZj+U
I5V1oXqoi0BjwSwfUN6el6lRNTj/1TgHVyhclBNRV1T0k36p+5hszu8JxMTF0fH/
49HChjaw2tW9hyyUqNO+RveKSsJMkz7ItdLD1hUiq0Dpn6Bkoo3fdLGzvAJpyPpj
HJKYGTOJswmhkZTkpcg8GE3ltkPakgAvi2E3kAsvOQKi47dlHPAky1idt85R2c8T
M74Zphw0otmDIybgfunl+gY1METh9NnoNYHYSsBXnptMsLlc7mUx3o4Et5q4gZ2J
vw/7+dlyjhiXfM96aRWuZxf6piHqrmjvACutfeMj3hq5nAo1yvsrW3At+gH9XNpJ
XIrFOXzPQuI0ISWcW8HhVwGzx05lka4vDe1L/PIdZjd0d/+12+gvHum5eXqb8Fc9
mxGZjr1VBCmQtuJ6j5j1TweCqpQ/86A/GToVPEYNk7bUcYWDwPIUkiIrNGhLER2M
N7flq9WFcnAsTtaktCFmXIaQIaryVyqMXTcJW+0OncNJ3BQEaUOQLkNoK1kOlMKt
AksRPXt34XlfxRRkn21jhumjdzzXJFhsI7NqPXp7+4/Ja3YUf/0/xF60UBbtxKGz
U8QdwgtgKjDPngpVJaxRehpxFjA4Y2G3A3C/nvUoGcO+MrOTwPoL5uAS6/MRuLwN
tTJ0Iy0MSy7vik0XsxfATTd2XhXYzxPEIdNTUx5/Qw7fla0ZRNRrddN8ZkvvZk9L
NjDZT/sFNVirpaIT1qp1ncA3Mb9obShGqIrmBhxfC6CMgxf1p0r38xp8rnGcyQaw
xH4hD5ZrUIR3IFXJIPPbHK12sE4t1PpN4Wf8cgy8AuQh2SnZlsVzjqXUA8IyZhuK
7+aClAMoXv5Xrz0l4dvrksMApbkDOcQZHMQ7J9Nz4Q7SKMuB/nKmzWrpNgZcnXex
k4oW3zTVapfJtVRDjF80NIV5oFKxquYwOgmV+UC0KxvY4UnXeMgmStwD6gvnpr1w
iV2kj2AebKx4c7P+xgmHKAeU67DDfDP6OSpor4k0rmRIyA0Ykvi5DaKcSqy3ZPwo
53D4fOjNn2iwMGx45pTKtk1TEiy5BOHGzeBDhzkRwckAheM+kwRJox7HZquthhPz
oSJ5KlqcG2cH7xAPxnt6RQ19QFTlpYYMlkzZYUBcRqg+HgZJ5N/yxGT2fGEMPHuB
D1yG+LZdT4xr3HOrKJQysNnNNb595tSBjSCvEvhzDM3xQ1HImYeDRxctHj8aXqrW
DOfA4j34KmstSqBu10pj3q72uMgLTUQkZ2TLPZzzdX6DgISOydAM33a0Vp18PN5+
IFy1onHJkmlTk0VEb0R6IihKHgewCLiITniQKKLVp2r+8FNdwcoDhvyyH6NI/20R
vJcmDK6YDcXcktlW6WExKvy6kh77lQAwC2xPr7c5NbifS1QJ/ke9EeOL2dRFLs4C
OB1+dT3nmRJHwmhZaHQnJo1stfYEXEq9W10zsb55nF5FEVrnuX4E0KoTclbedbqT
19FddL5EZdn26IPrHYquCroXLwsTrm2TpdQtaBgkRxg1itqp0/XlKZxX1FvP72/E
3RbWF5ra6ybu2bJCL/j/48Y5p2nsWHG1wuFYlcvMU/kSCCUAIewUftXtSBzRN4IF
JWi6n053N48D5PZJmTojKrlcl+6O2FIdrW9BbHOX7UbBR2NuZO8lWdyv6O9wPzqM
08siNhEMeHKxSVJSdtcHNYXCjcCW921cw/yF296rB91GNDbC29m3FUOaWGkwFw/P
h3vvnTadCzIr1Ur9U7/i2Y0GNccG4bAZE+uutD/Pae5SZevLyqurvi3id4vcNJh7
GMpEIgRfGY5mf6G7uBoY489m6kPSpQ2hxwIxOmbqFZF5hRC7d4P9Af9VntzrzBK8
tMi1U1eLDmsNwRuf4R0k1MaxouF1LiN6WUhNFfVlvilvh/v9IPYdKYgIpgegqK9R
Fp5TQJIqXxi9FNUpPR1746BCQaVkr7W1WQ2Gl8zRJ2lzm3TdsGjRipMmb/R2ZgXS
caqXWCRgJ252e8tPYWPLi6KCAZVqnWq9SMyPLifL4ZqIAMt5hskl9JyJn+0Uas/z
2vrC77H9fBUq8LbrXLiV9RDYDOODQWaWY5WQQO3McAHognJ3201nrzdV407ihfH+
/v9V18VhrFB9yBS2ULdbkBO7BZ5EsT+UJ3Ljn5+5z7ST/QWh4Dc63Nb3o0sJi9bp
`protect END_PROTECTED
