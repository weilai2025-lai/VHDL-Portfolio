`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjgGu00BkAW22mZVNUz6PbOkoEFt5dA+xr+/nKDU2OZyzG6Z/zAaB4P46u9VxNbI
goCNebKF2CP1Il9hIqwGwueAreOHGftBCXriGiyRg9txGWcg9xSTAQDjirdLTJnc
EpVyEVPp2u0o+T0zqJwXgs5dIuosCWjf6m5SQk9Co8R/wbVISl4IiHlqwdXSpzEE
g405TXsIS0rUogke7hNya1NwboqyBkpclw2UfTE5eM6wykul1YPXWsERugF1898i
p20vJx1Z6NI+IrdgyCCBfPcON8pEQKM/eYGfX/nyEEechOH3UHdJ0o7QOW2a0R0V
aEkZctFWZuIm7eftwNNme1ZDiTZdq6IkSjK3TvQXyjYR4v61USJYIsn9Go9lHMYp
kQYHS4FpX5j8nT4TEj83asU24ei5gpx3lCjofnEmFopiE4rPwnbkCrkGgTggqEE2
8H0NMdqynqFF3Sn51AUQUDhqJqNZ/FV6SpzKaiytKanX8p1w3t3BngxeDHB70DpU
vnK8wcCiki36P7ZNUVpRReb97B87Y8PX5XUblfOHUA7vG38wBkWJGTiNNCs9pBDG
BpY/rnvcXrpCJ/mMgw5ErjA5j3NQ/ZEEgKsIR/XWfkpahLc5pYI1XvB6QiWl1wqE
7WeSRxumwzBdYi+kP6WIi2EHNddz/kpCv78yi1TppdgwM3JyObUz/Sbw2+YwRD9T
otIRihuv8Ac73tdB2RMTgNWJ+Uh3LNS5mILMx4HiwOEA51SDHQ3DtNWalVit17nQ
2qbaiq6RLKCIdUcYI5HxGaYrNQSlUsVj29RqcpI7HJmjFH+dB1uhnyzM1vNQFe0X
KlKR2crPNCoY9tekfuoz8W6RFsvmKIo1JDQT15vzBvzKi3HpJUY5aZsVykWanixE
UsqbYVPmgSUaap+5SsyKcTn3mqawdVZlicknsI0YjXI+lsY0xNMgVXA3zEYdNpp5
rM685NaxkHg9KV80wKze6LGPD4L5XFD6B03IoeUz9HgrauAWREQkBDRXOYGh6I1E
lGSazry0JN05dr/03Zj3PI8XdGVdT3yiH5qZMw+y1Nf8eW0O+L2GPVE3I2j57Aa6
YDjzJSWC/xG9A8F9fflBYHclZgyQta0iCKfSIAJbcMIpdZ0cactw4rKM8K6hbzVb
Wy+adEdZ/5anqC/3p50lMSnXGKT3PXu14N2gQTBPsmydT8VArnu7SRntXt6VTPOz
qcdczTNSO5rRrJRIKCQu/oz9I7e+33OqX0tkQpDyJw5kFApuJ0g55qQHgPzWkHHJ
PhwVRgMVBbAq8uVNm6hbRM44XZ4IJYU/MMtLdLC/lcd2I0IdAUreA/zHcaNaEsep
AKkEf270EkncdGtMCosoyXB09u1wospJU7i2S2zmTpeMMFJGBN9BjRktQQw/Eqde
58OHShzRWnC0uogIuNd0euMvQ9WWrch0mVRQB+Sj4JP9Gs/gqCeWFTqvdjURt3Hd
RWWKgWlgRac5melll0i/e5BPCrhrl2Lg2TtAnIj7pHJ6epYsqxm+KasIr6IosoQ3
K4z3SCQXeQH9YZlIYWenSmAppEYusoW3EGFrZkzDmCZxjbofTdxTNJ9No9uWSvzq
fpZxr4wOeqpWm277iCmul1VtZ2Q9sse45v8Lpcnsxl7ik333vCfQDGryC5nDGAc/
oFBxA7zcELcA6oM3cmCfzGingFcSJNgniM75PisWk++IQVtQKAdTshKnnejPKTJS
hgZw/wH18nZYXEZmHQ7+8f8x3wIa+qlTbxzFz6GP847ume1QpbhqW39VNPnuuflA
2L7dTIXKmrcdu/mYt3/7ybyAacapuYpWj8xZJozJ07nIZlUrjgKzWh2fAHc7l60b
+0nQcJyvigKU9o1F7NC+1w==
`protect END_PROTECTED
