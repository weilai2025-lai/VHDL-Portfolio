`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zu4foGbc2V5RQr1LE5DfaX6Cu4Mj6L+5VMbenRvLjstJtsX/YOu0GJabw/lwwQF/
Bw8Vwlm0lv9UY27LoWfp+YL/7/3I6CMzXBaJTAWwWGSIuFj0gZjY40xkzFVz6Sti
7HeNROyA3S1+uZseDiaKBRvW4/sCeMM6gvTti0Mj0G3O+GaG0nJeccoEpmt/eoKN
CanuKan7JYns2vaWcsWwzu6dbRtymjul/iktYa8nmQDBfMv770nTwBLd2Jl/Sl63
T95WGTv4sN1PRfvmgZrkEXF4tqf2sgF1oJMZ7Q/3fBVyOwERT+79CZ3Cdvoc5KxS
cZ6lQ1LPOlLldNOpgnrXcxb85T7Swr6fRrFC7+SMF1gKWYOynA8sjWv/GQeEQqt0
H4jwn6VSi9+MdGiH0b7J5+A3VREedZ4AwYsmdQzzg+KXMgVFGOXa9bczKUpMrJPp
1/J7yxfN37O8hekvF6/WGpglxrEjZY8DaB4XnJghTZm3glIkqFkL4g2JmWvUvI3P
nPos6fCArsodopjX6SlsiAfOnAmFqz2Sk7nawEbp/8/5BfbJzsySe2DPu4sic4bx
QjtBxVqljeN1gCeB6GWzFyeDvNv67XipA1ysrHEmPHe+7smt/qKjhd7tBDCqr5en
dRfHe2nEWtOUUISY2e8E6/ZVVzYwJ0DuFe9RS82GRBqlxBvZJoZk7FLzdtyzwf0z
QXYKGvrQ8AHAlUkd8ke3QpoTtx1BYYHCEXXX0na0o9/+TmOrbP2yj1e3zb499zoK
N5hoER/vB95auzxIDIKveum9eFmyy+Ht8oYTYRuOwdAE8e7sjcihfytCwg50k4jY
V4Yyh+kBrMe4glnU/uIevz2JMwgZr6V7Mr8yxkxiya7ZqAyfBMS6x52uMDQEVMh9
TUr7GwPCA3pnMt51CPMLGM5VETAwLTPg7Au1RnYSffYMmhshwPuQgiqowJr/wqka
DNgehgcbdsVCUsUb1PQc9mwbxAjWBukYvNx8NILetsEMP4DkYhqNPyqTTr/BB0Kk
2bZQQCJkwkR9ZYDujda/tKjI16wm3xXmA/0+DKoul0gCAFVw+a3t4IHM1CNY5UEt
D9Ng2O1sgjptanfRL9NQznZdMN+CFBrJmo02LKxv8lZhou8D4+CkHrp3sCx0FjZR
cmrwP9QBFqcdgzX15Y6GnfThsHmZ9pN71EG+/d1D77F07gqmqzQ92BiHlQJmlrRM
26mKeWG2XJFjjr2tJGO+ACWS4h+ipAUM+B05pD7/4ZbUeKlM+eM1zFtqhcAREwuF
778SWKnQz8gTBUu4jwb9aiDwemAonDs3Xsic8RQDqZGSprQ8kqVTlLiR0iZKgyZK
SM1oqJy2JG8r32c0dNDZeEASDQJJnnw71nJ8TP6SQL0ZLHwob4T2BtGWH28VL6yH
2KPjc9gbvdE7EasW0uSqPQ==
`protect END_PROTECTED
