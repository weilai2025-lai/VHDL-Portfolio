`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcmGj5isr3yf41n52hxRbOPcG2sAuqdUSCQacdFlUFNepFPUpicwPxvFtszDnaVT
NN0fyusYhryWE2n+vF+8bcGdI6RHKHtGSASyGD0EAkaBEQfFvHjAiE+5iLfC13Ng
INEAZ6RqOpc1EKbi3Uibeg7+uNHbmebKejS5Gh0OJwSj/+r8CH5FaE4V+vZWdZ3+
YnWWtmOBoAWvIWT5POxpX92BJeWZh4gR/aW2zWKvqzHZHVjX23bECtS/8eZV0GQG
ZsIAXVeCAJs+P8/68hb3yo+czrZsMwRUS3TKr63oRyuFMR9mnQLQFQSAmcAxbIbA
ZpYNYIL/sx+NhKYrrUnRX3MD+Is1BNZ0lo9HpxkAaHFE/Eb6mdtzfjfxN2NC2e2m
tqrtefW4c9G8jXXxGE5yBw+pQcFrpcUd56RYouiJfbUGGdUlagJE1wAUSOsYWv5D
lfAdOsqOpD6lK6rHgUnii0T/NsivS+pqcRTa9aK+Xjc4rxMZI7uvG0jmqiCdmkVt
moRzwUzGHZoGRME058PxDyqAzvfo0C+3HPAiKEqAN8EjPTXG4+XkLciSZK7jYPTh
Y+xo+2hCDiAxP2KiNwNK7+RNlS3Al7yOg450C3COwrlDzfsSkZ+1zWFgiNy/55Va
+vwPBNMXUniBt/0JDc0oERr914DxBA0PL5icr3IgDWo8+Cj8eCyHkL2gkQ6IndOY
897+IWPLx6MFqUVar6R60aQcJw/XJm81DyEIyiYBSjQEbrWCJOr/tc3r9TEe4EaF
r8sLOCGBwToxEGEEX3ueHBR9f5QhdvyF/Bbxtit6HW5kaHbCQ435nvMaSfV0XS2K
eQoYl9NRoZZY8IrfDQNpigFMlj3q1x5TYqhgQLLvqvxXOTzAwp+LoPNsfQOeETTc
8UZwLk1nKhjOhWWtk3w3W2oZhFTpQPDYz36VDT2sWmA+VhcNoYIwtJW6vpVsmZho
V8jyyYUeh2W4N7ObGYifIxxvytvY9ww7lnzOhMsqFXbpXF5uDwF264ZVP6aM8Hxp
C8bWfKzuU0yDIPsFJ/YIwkNjMPh86H6+0zhimXfp70Mbiw/apwt+fZICpwzroEUo
oxqs5cP+v+Rh3vmJrJUo4YNNO43hoKufGqbg3K+5Z20=
`protect END_PROTECTED
