`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rzn5ZylHo+XPrXxAWEI4dybu2DylZgE5po1hgX7oQBEstoBgL/+l+eLesWNFLwVw
2vfyVTv67ytbUcMR2Ua9Hr77rxPklJPfAC1QtlduPh5pmBxAf8NBSGKGi8Vyu4qV
6hjBXrSkAV9VJB9GHexsNL+2k7xa9fGI71+ddLToquGnh3oSSsoZjxcIqb2ucgsh
UCk7SkNW/gcDV71ox19BXAWMpYVYYwjjunBa8bOvQXAK8UozN3uZyfj5NMUGRUhz
jKYIiCX0VtEUqIZl7c9dQCYblVyLctkJpckzyvklQ4/C1Nd04quR6yu7sAvGqAy+
ftWQs/QBl2k3zr6M0J9o9zRgn79vl7+2fJPrgJZ1JJM54M2sNOBD1BHsq8CKfV5C
/beOVHWMZtIKaO0TvF0YQSpsTKn5ln+AsMRyZ/XLqpOefrCrlX6pKAeyzgRNp70G
mBU1/fKq0eLWasCUhrBbM82sJY65+otZbv/imKx9sUBIO5UjSN6rf4CZnx4tV7EB
tXBfndf/X2CpzMQ6roPOfr2ZD/Pl3BSo5GBZrIx6ajYq03gsGxIpnvGTWBotBIvN
xVFuQ+Gz+yPgHyMLxCM/lxzW2FgGYYzz2uSXRpmdQ9oVDG1JD4nSHhpeC1uiNrDM
Fd2w0DYvlscU9E/KOwY2EoQc3GTLopoh3AygZLNPTfQkWsYPxM+6Ki3RveidM/Mh
S6Nfn/Rpna1SsA4Hf2VE5+DSxD2yYXRmIXkAZM/+ip9bRPICYy18hJqIkz9q3oaX
vh7u0PES6oxWUvZ0MGTa7o/Lx8ApiWF8IS++77AQPPHVC5BAAyBiEWBkAoQO5kI0
GYrc9ydh8bodoenw51KsR3Z9DjEgVZJeycbI+4RrOYpOIHgyJBD6aITY4dsDBuDR
9hTsZ+QHzCaAL2y4yqe7CecRffvFj4NxHSjlL0TJiWSCyZy7QOX4uLPDVNUFlP77
Zoo67OjPEoNgaUMV3BoEupV3ScrhN25SBwArnNT0836KRrXxlc7mFQbwND2A+4AS
64c12M4d8SWDT38nUrSalbGTWfJJbh05w+04HDyOS/PIv9hDdLGeMFoKwRmtawKw
RorpbYeHZ2kCE4sgtt6G6iy9lUDvTN+hy/olqpzYDrTenMOG94PoFmWs4JQVieJb
akfE8qVdVXrUG9EKTlvfgZOE/paE6kxTG7e4y7CMdFg7pWTs+4RKjzzBgSf6lImi
ovpW+RfNCOPHjoRUXhKyDZ2KKJWmLsVg1JxciZ2FyLBtxQ8gzE6dUtKx9OXRUhHW
0jChZhJmNx1rmQkFW8Et7gO6ulr1pBio5pmCiKq+XOGNqvXdYAaJEt+rUusIG72C
U0gKH7AnE+4DKW1VMsQdLZRzEbQQpGLVjrqsA6ntDnxUwBl9JLYkAbgGLrUoh31F
`protect END_PROTECTED
