`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZCtlgr4fUnu3BAIZhR39hyqM5x4x0dVSUlKqm4QOdHHqF2HW5aL2o6L1AKfnS6X
tzdeZISGJ4eF+k0owjxi7yS/ibgbFJ0y5Bu9aVAYi52K2wcePFYyQGk7bElgcQeP
gWYZv7Cof5hKsltg2H2faS75dCG7skhh4sklzVwSLM12cv+HvVsJcYK4EMnbJRaX
4hmlCqSh1rZH/Uno4GZ6kaIdtzBGSsJRStCL31e/gGofErkuETFe9P9U+1qp7fkf
7yiMDPP/mapr9WiXovDVOV2PtW3Nsxn2gaGavx7b8nHRahbRluxC4vgoddU0haAE
zgGi1eeuFgSTyLhM09ZDcPPmvqILf5kOtDWhhhpFANfqLxvTNT0+SYNCfCQc2klw
k3VtlDH8zN8hV6qqqVUg4XFx8H8Sz8nTHL5rkVaA6OLE5uFVso/owD/Nqe8HlXxA
VnF1cbd+wIb9/MCVoyUxtDXiAVzRprNy3eFNmZnexjbTEqiWo0SuqkEQpIcXBvJ+
IovD7DJugOXVZXGTOX5YTVvLM9FVItNfL8F165K7DiUghGfML4jSySGNyHfQmqUc
N5qyaebzQnBZaArvuBOsB8litbeCrwll15VoQMq5/0b5/Ac4ZiwCvuvlJNQ5IfZQ
vuw0nwVpJNjZj76wrM+qo61hjjrxGlh8hpkh2N1w3hkffzVx/7a/qJMrebBOqMWG
6SZq8KGBmbNmyG0QTXPIqccDHKaDlrnsyLQIQb2Z+3RBZG9thHY767KvhZktmYrF
Mb3yjS9A8a1CVTMoj0MRitHB0IxK1049phGetHurza8HZRujCRsPo1nUiJ2p8wVf
HD9R4yRGBz85PI2apw9Zr2xVLvcF4W+Q7qo4DT1EjBcJnLk0BbmV/e1dA89uFXej
3EIUhb4YVXxXZzAXOHqko9naoiSR09u19X+lGpvzkdALCJ+plnWcOfELnDYKuddZ
LERgAKjmzyHQyGjul6H6OjnzuBSbVjLmnOHRG5C5JUzPQgp3lwnV8LeI7s+MURdy
S0fZiuUu7HmFJFMT17oD8W3Z8UFC44OwJUwaC8Q7SWFhrblLVDx0t64K2TaPfCzH
O946ZCXlHvFy+tMlMbTsF3iAGtIDGwT3nfPkYBbJHUcoA7ZuNtmqFPGnnPtztifK
GD3Z1yt6Ey400GOMqMg6jcXb26H8L4/Slinuo6Orsv+hIij8dVl1ff2qASY49ojM
1AJuPdgnPjB1QGmY4DsTlaKEgxcjhyImGNsbV9qIySZw0JGBVD85ojNgSEQAdJ62
zZuvtcGJKietgp4wu0kwbEwHf0/0oLFJAMQGW1JsIb8zLeSg+VVOYn/j5zbGXJk/
MsnWkEJfuszafNq3gBQpguz0XV5BhPBaSNMbPlbxEQSRkZGfUAn57YjbhraAGOxj
VWo8TvP+9JZreTUgnclaCri+fbh4RkO8KuzujKZTXa/iIrUikr8WOAygVAs4xcWm
ON0JSro99KRxFnCaHdOykSqPcCIDoDUijBMQME57Oz8cW7pEIjyNnBSjrp+X8F5e
zzescU22FrOvIxOepq4jz8X1QLfobUpJNF0lWztKvOFLL37mtilS2ORibbLyZng+
5edarix0arg/+RHVlhGatPGS6QYo4H94BRgReZiuE45isDfTiaQWxfrhICIXunUF
miyLr2pdtBIj2FJVoRrjuiUCwyK7hEq9ZX6kyWvah4D74F/M9hOd+3X8rRBj1lz8
FL6riVU7PkILCsE9oMhVzx8AjdKz1U5RykiHL2L+vg5+S86VMGKVeqph3LvZXSAB
aVFGrbJ0mNTtzI4hV9eLhLzN/X5dWnC+xR4asEjTLQsL7MeqJcfwv3hEGm52sKZO
CBSBCGJRvziGDXziv63JaMN4/4bU1a67Pm8/KQFzeW/XLwPSy6aDWDipAG2NhnE+
rXZO73KQzFMBqpvQ2pMtiC/ckEmu6xhHEu0AEE/dUIiXLyliWixwvDQ5w5YnvHVt
/D5NHMgk+52dU3WylxXyX6F3RY6qJ08lUPE0jcr03nKkLRLWxexUzcuEj+NhJD0H
V6Nysr2o65wIoymo3yXrQFAaDS858BmDYY1r2zpfss6DHdk9c+H80YgLRBJNQeTq
78UD4IFVX7ChM4Zlz+XBXh1rCjYpvhufh5L7fR+cf7EYkxY4lgyFR7ihYUjDAJ/8
YcpHKXKOcZnD9tuDcsvHoxUVQPT5cMANbR5//oV8rCBiSn9wK5Fi+mgT1BJ5kqwB
uZ51M+Iixz36372SHqcCqaMlbrHdEsDnX4U8iIaIEfy6gG0suPppV7vTA5CB0Yvv
5Bp951kg/Yl/qonkjtNg37hxLF3mU6yvR/fPWXARHArV0gmqHHcKmgTNhDXgZkI9
6jFwiCygpssyvkdp9Jaesgz3rOZZg+R6QgMKfMHaBCHxWZkQH4nteit1kvXMeKQV
c8kO3qJC07acj6X/av6dFeyms7p6yhRpNlYfRxoJJpunVjcQchKL34NINfMkylMA
7QodkudJlGT3rxa3b0zrhgNOfcIjO9B3nfM085TJjRq8MpLiLM6glKbNFvc/XIxd
LIcV6tic/QvZ4gWWSnVUjQxlsuJbCtlCtNRxM5Qvs4feTDFSOxa37sVA5d3Pl1wg
q84aRMxK/xvaYIMi1sadhOW6u8f7VtLN/7Kh9NL+kQBrIfTI4B9eOlJlZkrvvMSV
5+ZX+5Ml16rNze77N2YLIljuo2PKio3D35yISuLg2pldiWvnWHQ/GRLfXLs6t5AE
s39a9bizJ/fkD4OQEJDrSZSHBSC6JElnq41O/NjOihDmtcBjAcsh/w7grJvkbglt
Us5cKjKQusiH65MQ2+wsIC7VzkQR2OYppo6I7kAOZJo=
`protect END_PROTECTED
