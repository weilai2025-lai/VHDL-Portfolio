`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rz6YXOu6MG6xH6+ZAxXJqLJU2tzJIV+pziSytw2LN1Ap9H7w9xj1uWTWcIThlAg2
+GrU4z1WyOijZFk94tMKx5p9KPz9AYAZ2nfQ3I3bRdER7jhlgh6mnJm/4mfQ6DZi
zqrf+cuiloXVJjvXKgB85gxGSQYvbDBz46CRRCiw1Q94+gzpeUr0VsmyKGAWkVvt
m+qrZQ3Ch7ktiAbdCn/K3h1BtG+sHzF3JFOiJ4xO3RpdhssA/7qnqIFOfoFfnsyS
ID98vP6+nx0IDT4FK4HgcBzORBq9FxU4amBid036sadPC5zoR3Ej+BxZf2y/Xvgz
DnuqXhAMFaXTE7RNJkKc9DqsCiGUsgJs2xQMff50ToxBiw6hqoflk/FYyQyzKdqa
xqj2xyzfgV3CIyfYJyN6quMLEJMzcQW+TBq5Fy8TlEqovgzdTygoe+8elUW/sRwG
gq1iB5/sjy942tsAbsdctEvF0kDnSbRklg7O8hzLAbohvv7yEnsiVoenmZyYfbF5
nMirnppoq3dOZ9L0ZyeHUNAsbiKpz71sTbsUOTIZzIiJOAikopolB0wgtxyQ2uKa
9RJCVSXAYJuGBT5Na+T6PdbhzBmsjX7DOg32hWPSYj9yAV4Mq9WwgXRfUVgqZbPa
zb/t6PChi94ojmJIQLb1xw2zjRTbrzL+sDn3otyZ0HdaYGJqe2CPfTooh+NRx7dI
friV+M2lxFK7QbBHhG6sUOjW4/VmRs+X0ItL3TCaYkprXX3/qEPlUqn/nlMDltUr
i8p8Ot3PNhz338MkawB/IUGlWyvGhfOSr+7NlLfsP3ZKxhfNqFvJbENY9B/sjfVG
LNAfROl3wyjWoztg996T6ZjXB+tkgyvkGX75sC4AdZUTXRa4O+qjtzFP3D4iapYD
tt3JihMV3pAlsu15WXPH70u9DlzxQQcO8iRaMZr7RWBMzQqzXKY0tZSHQSTNgXXD
R/1lLKbF/qmoqDh+5NnUdBzALbOSa5oXJ53/npKkqo4JiLDE9mbvW9/G3rxmh0QP
fnTzihWiyikcCOcub15we9TB5GbLRAc0N+92Y6U8Sw9rcPw9CM8aRGLX5tXIZcwb
0YaxeB//gwv6fy8KDhw9gkDSsPCai1f+4PbIQKafOKhRZ+t0rgqBYoin8lXr0eHW
f30kZkTVWiIXSaUUYcAt7luru9uNTti+4za6WY91U8NP4gqCJ0J30O5fqrP7gz/z
mKu6Z/miHqvj7IqLz9+mNkOS5j9udaFn7QiumZP4S2uBzUlbLjwq60Vrs4qisNQv
27537CWOiA3yXYUAYBP2U4EQpJmeakFb3RASrrhT7PkmoS4zOY9o8R56G5nmmeAG
v4wAjhamolVv7ciPtNWZ7tftYZsK8NmvuLBDjeH5B0mi+xHogusa6ejf0wRC9fSy
PyIuwLQS3qDg/JzfOGE+BvSrFh/XOb29T4j2R072qyoZEavOqqXGw+VzRYAlSdIa
yMUol9nsj7LpGpWWu9JfW0EzOtPl86NLHfjlKcWdj7g4tDyibQyqLOrJy/T9C7/a
fRjAlMlyiiOlvGjJNCbQDs68x9egGY7sHNozlwnTxJ9sTJRlkUUkyxFFr10sz7yQ
ue03D3/+096MZd0gEAYVRwBV8FokS39AYhFSrM+yS5enzdh9Z952w+KRDbm0c0mu
sXmxiwQYxaJsMUpSZfQ4uRi/a5j/2UuB03ZP/mnm0w1tcAZiTRzHjNkeXBVVux2l
6ASmmiwkzIjV0Uge1UyzEGvOjZcJrKTxvbFusvqGPsTc85nhrBptnLlYDBE8iSWD
HQ/Yh3bMK+uyZMDnlDYo9vlfTtIATgssJhbVsem/86MzUF5vYSrKa1e+3Edb0ssf
OgdJ9RThsC7cd/v8J1G/e9NZ56Q9+UG01QxF4C+soYoYX1+nim+bZF/WVg0mRkCa
l0WXmIR7WD6uFBiJqglhyvBRFt4PCbVHJhKh4JQZ/17gnp2bjSYfdwF4aJIUntzj
dYXHh/WLEO0JOQXdk4QnZo6U+S/LtpyTegPhQu49bzP/rrNzGC297iDHgeIkzZIc
/QLsLfNHpXJp+zoFzQ6dOIB7DZI5eAOv+DRc6F82oz0PZJIofpXhMLV8vogFVdkm
2UOs8Ws8mIEBArFZ6LVig8LKg4HtEkHUUJA0bXYGxPGKUR3f0EDRq8d/Cp4S+luT
4rPl/H5NVc+88L+4UZQivvK2GLDZATubSiAxovHrvstrEv1JUn0hpcZM0lSBQV87
5wWRH3a2bhxevv3jlY+e+L5aLccfIgeAOu8Glv7nCA7LS8RDPd43QsCzQflyoJfK
GFLmxPzNySX7gSDyqrY3iVwp3M+f6+DUTERu3SpDpT3XKmnl9na+M2CQvx6PWVGQ
2itPdigiyC+qt8hrTa0IJcStq29JMqDUGZ48cFyTZStTnKjesA1W/i2f6xIO6qcf
YCtjQf8khppVNsM6V997Fk7GiXoBnfi/nehObt3v5L6kf9gXb18F4OCmfkNXyO7J
XSsdOoLj83QgYBq8h6hfQaBh0sNu6co2BBR+Zka7pKwUtZJOW1Sx6RCTvXh/zNsD
cFm0mL3lq7oL0yjlZNBZDv05lBp/oqlZbIUHW+bDGDRPODm5oKRAlPzcRDzvuybJ
VtbPdZiKxj2VOMKFzGwEtJePNb9Pvz5fOFnYqCpJi0SH6KnxR5vgl0lvfstMMfdC
7FBwc4ydwpZ8r8icxHnykhHM1wwh+s9d3TiyGne0JvjqlzkZ5/nMqvYQwnbfH1K6
jyp9aFimjoNb0UTlKQeVqKXDPkplvovoUy0JFsdRDpbTQXV/obfY5bKA4tmdeHFt
TASZbeD4M/aHxnNmShKOS/k9I23ZcYcdGQGKy3uIBybqLYqySpX4w+SXild7YNDb
ZqodfNHtkBThSyuDEpD9pE69H0UtPFfqFjLayyZYcn3SxBaFdtBjaaJ9JcGCsSWv
LftJ1VAv+BZiD9gzUOWjVhHg4xSIuyRM0R9xIapHcDSX8yp3rfmvJrfl8sr7Vw0T
/dGAeeiWrHPcpMfo2dZH/Th2Njz4HvPO7NBSOLkcV//3I9m4oAKl6mpwWvz8O9bx
sQGP9giGW7YCGx3kdnCNzKxkZPotpu7n/hwK2xIjwOftNbhtam+KjODfP/vfbFhl
tABsZqYeoNXb3HHYP8HCvLSWUff5Ap0us3Nv4iiNPsZPEYtbPNizUxwg+6OmdIhk
actiFDRJt9KgSkFZc4KnHU44UsCpV4cymy7/xNiBe+Gd8Q1QwVcEhwtUdc023l9S
GCmUbwLl4oCRz78yFer9QaKkSth+9hrHXv1RZ9RWfpzrKiclc6yX70K/HeTF0wlq
NGpUzDCB97ZuZ0An8+mF3gMQmNSMwwC3YuVi5DuBPzO4L1i63P8baV7hLYyavyKJ
BNDTY4ZV1993Ch+nya90vhfcpaVXE3PEyQsz4TwdNdSiEiIQftUjM9ssnxfbxmMU
KgoHppVJSz+V/GRVm+q/TAQimL7elw7oiZ7WTRvQeVuQQxKw527Ma8LhcHD2RI5i
L5J0FpI3LBxMzV00wXkk7tEpiLzU0qYKNXZI+GLGG8AzW9cakZxPw81zJeWXzu9L
7j7F/BVZy6j2B+yZ4LZonUQkoDlMX70s8o0TIYfOm5wnd9UcZ8kOVUg+JaPwyQcw
S2C6pQGB0sVlKxe65XNH2hS87qKjuFF2YIfc3asRa3nBBhPmM498ecLjIDQYdP7+
rRf2TWjxi/G3BHoOumJAlhKeCDisCBmkC1vbbwoTKnH0ngvyceVlxK6wy5sFvz+D
WlZrvarqqyn3OlYAFthr4+5WCdG+NKwLl/Rvcjjcp+gtkclEc+eRyJq+GXUCPibz
2vIvqvbqbZm/D13Lq5fjDTNEJ8/7a8Sk/kBw30s9pOpL2XEDbPRmI5P38kE7Cxci
DIFzMOON+XZqOqIfjbfqpvwFazrTLx3O6LEit+F2t5wUsszqyu/DJD3hbjXpgh7z
q8dCDRK+9rc/FcJxu24FSIxKhfAot0JwBDZwNn7pi+4GyRH/H1EUNaaRU3K986/j
Z2QSSXgG0M+sFdPoHjmP7lAg9XYZOIeuvKmGCRS5QMra0fQrJuRu/4We/rmbWhF2
4Vg2e+aDfQq/Zg2iGHZA9yNJ5BGi6wl8JPMjS0PtRonlgdwOQs2TA3BWrhjEn0Ed
QxtuPRiI4gs4QXPMo6/mRzGNch/8dO8/MMSsYYuz5fuRF2so6fwqt8kXmEAkXAK5
tgewTMFLGFnzoC/H7ibix9wLgERhyWSmySH0paf15qW4jg1lNGVR6YW8hq28KtZ0
1tpIquwxcj1egSNRr7DV/fVYK/WcjgmSTRmLOoYPksTLruvEapYXEdQ6GMDw5Ubs
Ej9vPm5O4f6egen6PYo7zyqyds/cqSmg0v8OUuTIfQ/CUGOhTA+UH5sfq4VGWmes
lgjOoX3c2oJPcrPwu0uT2gCNHb80xcQ6V9FBvoQ0CnIAUUsqe3HA+mYxo3w2VRi5
ziBYNcY+bKPU1lYqiA8MBxVdPjgv5p7/lIAGUEq1+03sOnUKbFl0ZX+nR+vOoPvY
Td78927JgF0MiM3nBp6kDzfJxk3+ZaSYIUmwv8/4eWEFu/de47zXG3K9bTFpXQ1s
rs9xCsoQ19I/BZaHDJkhU5Gwt/+dwJ6dVf2u1QgOS5OTp5hUgwvqTymDogJ3HA43
KhKXBDgbS/wiMqWJS5YIn0BLE3vxDHHFS/nQrL9seYahXcFDIXZQnzZUFTGTA+Pb
7BQCnl0Fw2DdJ+Wg4417O0y0HNdLRUmGFIY4/2coJt13QrNIbbUyvFqx7ulRlnXz
71oYihADKaHvGVCoIU/jasTQWps49IhYz3cmt+b9L8ltZOUEJg+6zR3Go5paAIfZ
Bbs/F5W5nLE1pIRZyofFMXcHc5/kVuTbubuNBL9+tr07cJcPTbfbYwt+ElTdZbRh
qEfvLUwg0kUWpeOhlOLsZgGWosqgucMDhFgy7QJuCPvneVPKMOX0OYU2/Gvs6HJq
hGeuhNgpunzWMIdVKzqp7lQj1eaUU25hK2+GiZreoinlovO7AywA1Iq2/c/0niR8
AOa9T+5SpPpdAsvVfN+q+y7MkdvTApH4olKRTTbbPFNjVz2uihSG4Xyj4TOJ9bpx
85pjSdopSHc0STlKE5sH7VjmPsKeE/ytV7nEnw4r2iSXbq1BViJCQ9qtlGjuvpQ7
rPnZysuJuAzpN8Ma9qQHl2PUdqPR6ItVZzvqtOcMHpTvR5axxuMn3ECOr6J7ZVJF
3rRYjtOyq+Vu2oElIShQS9i8tQUr5qdAHZV8bW5YBOU+HapK9RbQprrlG7WVR6xm
AigZgckNSP00ShlHlZ0iQAkNEu2gBy1qiv/NqCOfxB8+eBJg/Lnnklu91SOYuqi0
gqibMuJosjTHV7l6HOWSyMgIZWSG9gBbiPQt8gmieqUCWwWiaYswHKaCHXW/SUpQ
HbDlmzggw1IIohMTxRWQHxgcsdSoAq+OKq0xypBwiQc/8BQGxlDasTAHz9H8C/v4
X8YlUJzbjprm8jYdL7QhkQd/0jPrxePrQkN7r6Co1gA4NPNob9xPPTnmq8HJpQk5
BkgHluNySPM1acZW2ElDWsPOEO6uIjtt04RRRsFjr3EBOHyRLD1N9oY2ISJJ9N9b
wB3Fa76SJNw/N/55IkQmjImwwECoBQrGQruQPxhTBMr2A6p1VYOGbwQyUN/o/3lZ
4FHx/EFB5TdBUmHZsRHzz+klQTBqwl3i/Vn77fkFSRm5mVMWKxm58jZaKUL+6YXR
VyDyUYNzC6TDPc1IxPW3t7LkLPN0ndi2TP3Zdz9JhrZFiRjZoC9lmR2sJ4j63tVf
xMQWLIgakwpY9nUzIEzzDy0eOXrWW/18tT4fMbD/zUjXCZPwEdtS5UgHvvFZvhny
KM8r+ymz61m0PJ7KD5rsRX2Gk8xorMdTGhrjzSjKCdmSZ0LWowEHOp1bJGqxAkG2
0LGbUAFNzYcRWvtFnXVMIgCaTbGUooPtaf7iMXb0SsTxksrSg4TV6qXKV6Ho9N5K
eJoAs1F8NVlYNTf4ocSxLWdR+94ejvljhWI5MJHY4znz09nFJIs5WArceyLICjsw
3WGD1ZSiwLI3ffANCJWOAjBnJO6r2mJum9o4cPjZgK0oK0w6rZfLGyru0HY9G4mt
Ip8S9zme8UDgva3L1dQAB/bkex9NiLcDmUwHG9zQ1gI3yFFPydw/LSNzrEX6+cPs
ZKVhyXqY81LBjOxrHX2AaXUEQ6Pi7tygUui8UWCGgg/KBPiroWYIZqa/G7nLbCOX
CUf412vWM85uZQrt2CxE6EuWR9GMiHagjPu2OGQMh7k96j2RJR4Oycmkh3ld+YvF
52WfiN4S05dxruyfdN04N3v6/3B+dEAb2hTHwlNObzNShKaqE+C/RPMFn7CF1CK+
WvmlLPetAGiXIOaw/beQKQYzYoLLJTRPRTjUTl+qLt/e1EYjX1EZY175mC/Wpu6p
SLth+LlB36XmIKDOX6pZov4Fc1TZMVlm4QPRUr8FLq3Kmq/NF7O70JoyvLQ8thrJ
jpUGxN0rKjBLiecxqnblN4PQdmWhr+2z4VpAu5nscAOwQNj3FeUDzokQ2o0CGdse
4eDwzoFPR+l4LLiB9Va3b8aY7ixJmzPJEVTSl43u4x0JKgL9LZml1QTDWVEs7V9w
f4wFpr+wGMMKrgSOFJOdgHGE5xyEjGAwQ4VZGg737oGx3JUQCaa/RhiaXi8bhA+Q
aRMdnZ2kpSzaGwzVqVH/2XxIwrQ/E3YZDqxZISy9GkjzJvy8Qpn5bRIrK0o6YTFG
q0ar7xgRQmrjqNYGrw0ZsZ3Gq2QNpAD7KbAsc8yE0n93rsLNCbdXEq1ojtzqs+/l
6myzhHVbd/zLIC7I+BenSHfmmCK0KrTgh1iQAD2PikxeJScRLS9B+iuMtPUqHlyv
xaJR+W65Gw4GdNv73FXm8HkUxhi9HyGb+NGDZpzwrIpbqUKy+XTDPn+lja0dd/nb
`protect END_PROTECTED
