`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cv8a2eEmJrVZp7NNdxy9XcU4wFjhYKXwhPQCzFcLTgtiro8W593TwaqE+XZztNHy
ikv1Pw66xZP32FL0eQuviynU2EHNJQ6tJ7Ujjea1MsKggZv5pvZ7rTXAQfEUJqJg
TeR4rCIqADr7ZzTu9uiC42cyiKpocHbVRCm2TalBL89xpN8CSqEqvREMxk33TgNX
RHnE9BbAthwrT2XcYTqOTDsSD/w0uIUvAUhy4YgFTCdsLbYsKPPBreiRf8UnKtj4
+PVtoIvp81MHP6Q8JeibYLSAKWYLXgPe3/6cG5peZLhQYdJTDi2YHjj4ybfJX10S
xRZQ+gAj4tpD41KWRsNUISGp4j3jjLwCf/1gz9nd24vpwC5dkuyU6N2tjfcmTvMI
8iP7jgAN0hvomLiF+BrWYQeEtMQHLbAPiZJgoZM3VBnQ5TSWlEFmAXIZ22nW4Ksc
M2TmV+MW9d2+Cn6oc6+3k1OoZ552xr92LYSwWT3gD5HlVvZ0cCPnbg0z1AsnqAtN
0aPZDHnkL6mxC1C2f0vH8C5l8aHiHovtIjEJXTuR2JZmN7/vfqWAIQ4J9kWbYLnW
3nJ2i/ZNZTPNbJg4Zht5QpQzFfVlrybdsff+hdBJwfgv066RPNWJZ1PZb6lo7Paz
FxhJzMiWhNZ+/x2XNVLmU3tGKsrTDhpvqmwyU1JApd2L58HgFgRQOAXiehRWppZh
eWg5E3A/IRjAw3T4ayBWKevabZJLxfhgMQ3lx/FLhrK5LznyKnS1j4BSOtK1SxpG
21uDk/WAr231ZffGluJm7S8sgGcFB0kvFyfysS53GSNVc3RUA2Vn9/N2EgAGl4Rd
W37GUQvl4SxL+uqiOqGFich/GQMetL7au9vpW681XPIYZpyw+SnrKqG6LeKIXH2g
SGCuiQDX1Q6c70ulGiO9nl2eUMebBRm+f+cedrESMuVUiqLL7inPbd3uizQOZFsY
ZGF/5x4gz1+NIlWDUdcBFoXUeoolkkMhgk4kqgmTUpUQ3E69yttM+Vv3C3nOfHxf
3Tt6WQCrD4wvZrzo6UFDDQqSZ1DHmT1gSO7JUgCzq9fh0+Ct9abOZp5oXYzwIHP5
L28t8WWYfg1jieK4mYSV6xrHIG6enT2bY25/t9PNVluiGIYS0UuAtWZGwppjBX/F
ahonQXlWW6gcTw+5TNHdBPru8614gE9vnU3HToLmxWbJDufSzPUunglJ+19Ysz7j
B3jw8IQ5Rza1qkZEYY0EU/VNpJZVCIGmFctAvzxbhVIabviOmiBJeN7F0ivLhpfB
c4Pobv605RVt0UDXzzKcedaY6BvpuUV4QzyQDTC08DPRaQNAmAA587vXfPmlIdPG
ECs0rxry8XKyUQxl+VZu/zXODzGsrNVCdGcyeP/57lpvg1GOjNrmu4/HkdlYqMuX
BtK5w5cxekX4WHXrOyB5LGWu2BkVXYfrgKtMLKwqQOoNOpA4wUCpZXfHcT74zmPH
tZnky/xWu+jqoaln4GsnHMBlrnvMtJTZTUuLNhAknfMSRG8gYlcAMg17ZrDFzfJt
lPcynzOIs2KF5QC6/BaSEOlIp7ReiGXupJ5+q/MFc0tuhW+KLuqwOBwr4WXXIYHJ
XcnhSuUg5IWcQOfRj2XlZiQAcc0wHkp68Okcm5gOHDg3Qp7S0cKRyQ9kyYRKCSeq
4/O+6G7fkeQHWra5TboqVuedv05mxNJaYRTvd91NdSzU+3FTGncJjPuFTB90RoeK
zYLSKFyP50SVhWOPFhweDasNYDYrqYKNajCJ1qDM21cwGowPAt4dKL7od7o5gZHk
D+VacCoduui8y4zE1VXuJQkBJWF7II1pnrZUk2UK2p1yqmiy7hzSr4MP8RXWXVt4
da7AkCSN5hTK6OFG5v92lK5w33yJ3nS6RtQNn1H/f1Rr9y9Zg6qnYlCmUUDwJVwA
hVuq/ZEu7QkFR2UmYU+OsCd5ssmBHZnrFoBM4bCscUeRidLeKTfujB8Kbg9Gc5bx
4C6zW+/uMoObEOYcY8t0CSKmxPfSWyRVRy3zqPsDXjKYsMVHam6YWO18pjBp/4Yu
hWL5+za11dSuXpIt3u8Ep/iLkbHydgBLhTLARiIQMisotEBjogk6tvHplnmeZq0X
0Imu0g5JVA6SbbQEkmFhzttgpCvD/OmWV2Aqe8u66q+7l/RytJ6c4JMTzd7KUC/P
REFGvmE1J7fzfTaTu2uxn1M5U+vQFfxvZhcLzGqcM5gsxq4w5Ui3qDQoC1CmJJYJ
n65iz/98HoIxvnDg23ZqzDzRavX/6U0iEw1hQB5A9PetgQMTfnDojCsR2+R/XGiK
sY8HFnpXN9NM7CKwrssS42+Kp5VuUIB3DRLh5PSZu52dIa6tndTbkS78hjeWbhsP
Uofr6dwyCBC7lnaxRkBnYwYOmrNg8bayAbb2G6kJq1Dxcyf6Y/s9ms2QQSpwnAcF
v68+xeqhKGPWMjzCo+0cOkOMze8+r6rZVUpU1EeONgbo69B8xz0yZ5WvAF0ARV39
pEcidtYv/ka7E8GPcYVS3rHCD8qGRvANTdo/vCgtkBF1ff7gQLXcmXMj9vsaMzyI
0U82dBTdIYcNJXpdtbsjIGn8kxrXMDtAZyzUl6DTETPMfOjoAuyGuvGHrx2od2Oz
5VPohcB5rYoYLJDzJEdeLxkCClOXtO3sP6uT+26xRpi0KYWJ+upj/pvd1G9GC5Gw
+xYsqdtiJWLP0j8s4kI8HXEYHueHUqV/uGH6a+HpbE52bNWI6M8dqLuuY+tHX/I9
YmmGYsjLMxU2GZeRNtgF9ga+DqFGv46qb/VUrHy+XvZ43fCEHHE2N5UjiYwX71db
6vpEZ9YL0kumbo3UkhRnwkixEritFqY7/MawRSWT8Xypyg9zRGdiFDfCxc6Q5Ph7
3MrTM7aKFpngGwSzjrjnZ3G2z9CscFImVgtMzYLvNs4+QSrG7rCNdvRGGe5XbH8w
aiOaqU1aS2PYZHO/8ZCiOo96kzyj6yhhch0sOmarcvFVwwhVVFVKGT8tFFP66ZqA
8X1wh0ikY47JCLSjDuSDLGBr6GC9NbACd7Wn98nlnybEuH6W5GxYtLZaJJNd4dya
VcHR47jlKf4CDzfj/W+SNJ6q5x1R6R9ezNd0kAo/hW82JU9IKODertCDmyOosO/p
BHmBl/Mx6/WeIH3rTIE3g1pmhXXB1IJVQbkpIYEEpfCM/4MFDOkK9UcUyoBLYwPW
mc1l5rxBZ1TUc9swXOWD19r2OnG+Fw46wgo7hhgPoumgq/ttirML9lKhQFNEvLi/
hAq9/KlIXiGPyQAr9dsSSGVA7JFu7sBBQNiiRELZzhvoda0r+pFAjpS3zQOvS3Hi
JOaWDFu0iwPZEU1qSUzvx5aDCFELAWxiM1/OuPaxLM7G1lnYzkXfX2fyjRWueBGY
4EAsMMSfgqxy+pyJdBAUV3n8hqMxZJ2jzWvkt3tACeHQ7bhJ+0QqggefuF2J74VQ
DFwL78XwoY1qNJht8B+YkVcB3UazNUvSSmhjQsbGq7TB7KpqxtCgPmjgjIv4ucPM
UL0EnW5AxouI8qLi9JJ7PkTfyxctqWT4S3CMzwjJA9r2SFVFuBElx/3gge1IK2Z8
DTl2tr9cE/eDIzwwTvdgguAnGGhnkJ8JLbtESW+HAIuQWokjc3GaKRn1LDVxyF4J
QIHIvY26CDPAlZizHXfkCiD2NLYZB0fNZd5TuUBKY0yyOiwxXHBLs9t7HejUGVBn
hE5w1kGSNQAnStx9u6Kd9mWIM5vaW0EVwWBlvHOncDzmgu4Z9K9aqwzwWVjOIhPd
BoexiZHyfeRqBvzsgsEf1dVNjPa2jqWQBexbEI9VKZ8x3T//IW5+w5zMEERbzMjc
1pEBWI/NE3JLzH0/9llDh35kJFHhgG8cARmdyD2+OMl43In6U5ln5wFTGA6LhS8s
PtTfC1JU5ZSR3OG/03QXneayVLb+0m1OzbEdapeHix9S/b1a8CIN1xINl4B8fKAR
ADNgNm4QVGJb9TgT1Y9ex2bMCMaPr10E0YW5s8P+w01B5EekP17slDpQ4Q4xhLiB
EpjqlWt+zEVHD9StnWFzFf2nelBVCbVp+lH7tx01c1auaQ3d2RD4Nff4PyXXWZA9
nrsvlabcDIFojCb1F5Hovw2/EnM6JATPpAThggk4DvImrcNkksptJYoiyP9p8GaX
Fe4PQMvUhbacdGtPQj/wMURj4i5QUHFlSsls9latERfS74w2nkiako/KyF29SFzj
RGQzkVQ/0gbMyWs/+uPwr57K17uw7dfXk9b1r0lF68tHMMOid0UdAoiFJF2V/Ify
HqvnI0uTtJbpupRXYcGwYKQaP4o32qwhYO8Ra351XIT2HFsctv96fVsf7F7hSw+4
hqFr+d6qCf8iGI9irG/q/YEiLfFefbcX14u7aUoFCOSuzVZYWkQ8yPk5wNWGGHnQ
FkCLKxxQ+2WPkY2tGFQx5crmqCUaPdG2GBOD2m3WaVTdyTT+AZSAgbQSjLxrKkze
ko955dXNHWvdW77c821zt5WtHPaPPTQamexZ7W1pc/HKcd7C4tZymSPSgFAUpyCO
LxnfekIf+0YVbgshdUMNHI9Jld8ivEIlR8O6DR2/GLLfloD648PA9SQwlXfsOqVm
9E80qmLaz4B1aYEpiX95IzG5QHDg0LCv6PypssOKa4bBRK6KqbLAu/jPDVD7hRJ/
jVuGvNwHVlBl+2sudn6AtO3lcba/55dhv5ql97dqwUUCJdY07Xv3UQt0ktZnJJKA
+ugPCGD7uqBTftj47amjWUnMywS2EOfGTig7Nf1TazIhRMGkaGKBQCs4ScsXhHBb
B8sQOEE327BJdSjkBXpo9mF9DYKyDtORiDwrq1dDrzjN1ybT/Iyp/9gcQeZ9nQJL
41QRzD2VCzi5EvQtJk/8lzakj+F9JtsaWuXofaAaUBNnPJjTasVYP8YEhTYWJn84
Uj/HvHCgm3UmFEWfYWB2cUUkbk2CrtEDSpZOLf5cE/vWIHsAYNfFsBGJfL62L4TX
2cRdmE0Xv31lCXPP6tXIl2RUZg+00Burl0gZ/8sM14d5Mg5Q2aiU+2pX5Z7sKVHE
KSPtPhg+RPus3YybNerYwQ5Kj4DecnMq9k6PFBsHm45zCeYE7b/WiDDu4R9N53ZH
4TNyVoObs1RNdFA+FPTyaIklfnxyrMCG2NfCbeJpIci1LSK8BS/ZFq0jTDkmrTI4
Vi57JJtzqQxbpv7N7VVJehBHBBXy4x/qUUASw2AFpWvA04yrIem2FCEFBvkwQb8/
YPXJmxN89ysR220VieIzLnjgi5PhnmNYN7Gz19acwKyA08bAwkkwI1/9drwv60KA
b3qskAsV8RnEcxJEEE0yYfSbWf2eQBY9/5oDmVHFNlEVnCD/gfEPm8PgrEIzItix
7xr261JIqfubN3KiCwDwHw27BiTC13nSH5QKJH+7wF8hV7IuE93TbvWHXyCuWrvj
sTiZTJB3V+LidCYn5aBSvmzEkWKiCkSTTnQNykWquR2CouGg6raIen2OXxRb+Ek0
yQmIo1GBbinTTK6OE+76PxA5bp3hdTHzN/Ov26H8pXTN1JS4SazbPkr/PV15D14P
r5QU3SEVJjOaolLUoNPufYbPYFwU8ut1pO97VrndwG234yChOVuUchfYvL9W6g32
1DruVAkHlSM2kWwiUjOBmPmHjM2ti4Nnv2Ns+EYu9liTNL0Mku5eMxY9U+yC+QSC
GTALHR1gltuaWRZMyo/Nei77mbP4QTvtTjVWgsoUAqoG4WEhivYuCEAm/BNysiZD
jD4VNK2CzR2O469qIq1R2S2oy9Xq/j4lOsslWTAXgUEGaWx8m+4QseVJszGt4JPX
XEQ01ndZbQ0iAJLDou8VuLteVOO7zDCw2UcEe+TRNUa51TNILnt94Oo+kXLjlcGu
DmSKsygjTM88g/0IninVXPnxEUTAFt9hMBM1jP/zkrkzYT/Mm+AJ+C8o2smQwir+
dxOcNaVOC/10vfUd1uUeLfGrE+syIewjkwW1LekcTpSJ5mn3HrRmTIsXDhwKtZHK
zaD8RWHSF/MwEWcm8+gbQdEgu4X91FzaD6fkp/0vfQCEsO8hn2uBoquO8A+iT1A+
M8EZ4a5DS2T5jo3Yq4djngu64hCNwMbEZsaJue4kfbGDkAYvY2UxmZ8+LaizmQw/
sk/3aARvrezMwd6cyxMumDizbj4kDayofJzI+45Qt+adq9xyGbuQ1QE4wb4wxHOA
O86AF50YVki+fp5uy29nrfjiyKTMPgofIkwYRdjIt3VpMzzNCdy0hy5D9NkE17Qi
h3fS2UjVTapu7e3627BXFdFXoqKT2hRdXdRlrmhTdIKh0OSXemNLctICDCo8iuqA
l18Jt2E98sOOJNFf0CNpM/ALoC8Cih77uLPpJ6wwRolkGSalh+bS9wkvRPiwPewX
e8Is/G3DMj3pxLnZFvExOJ03WiwY++kjIefkFWhKQ8pRWI3nitNrJBbC9NPSgJe4
4Q9fUwMJO4Th8FhkISuPY2IBe8awN5ar7DAc8Tk/CZNRetlFQKyH01bIfLCGvfSO
xpkcc9JBnFTj2L/WOO1vuoWE3kUKKyJ4x2+nqBkotdXbrS+BBgv4vwVHgqyBCJXf
cRx9+QnvK6Km8nRDThYOBBsKVDzNP+WTw2NJVXx96YzB4+Hdc1rsGs1YOC5bE9GK
K7rSD+qUih+D4APH/aa72MJlceqKsfHQfIf1vi0mpLfl00ugp17wF+hJAw/iPGgm
r+Z87SrP9UUYfPhwoaEyiFORGgrUpv76x+hFTdx6IrNZH6wPIU2oO2WUMj6WxrPV
rn0qxUZV1c0WejolkBxbkuMqfWT61orWSExWLfQ9l2u3OGygMXTd182IVpjmgzC0
SaF9UlrmObe6R4RMQs/5vG+HmFKR/QgctIJ28flHvH77nsmKREHZ2LVZLvOHincz
zlyiR/iuKiLHWpVF/PteZJwqChmeWkwcYRK+gBgREl+4nCqLU+W5YGfMJvIh8rnD
kNLjClBZmrKwMaeKVFUPIjw4hp9vdS8wCA9smQbt0Cvo5wLskEOreS4BKHEZ1wEQ
SjbCSm1z629o1mrDnmIVZB2M7JsKaf1UU5SMhXTKvQMm8s3eLApyqp223fi1P68e
fOLvHS5u2FSDEVfFicbyicaR0cOvO7Wz6YZlgp68tp3AlvzebanGOjgLjvMYBYBX
bg2JMF57gnzg+DMY2nC5GEpa2uR9HXRsrLVPEaa1Yn82ADvykB4E+3qpMDTaw6tg
7ySgtVHMy+ftMRGyQ5sgD1WvcajkNXw6knACML4yt8tHXhZFcyiVB4iDCfBfCO4d
d+0/sgDFyqg+qcX8HyNjmrBqFmffl7VKJbiSCmK/1tfrx3XJijj56JhOOXRY9dU5
RIQMCW3WnHchV5leLogdAtiECHgcmiihKVpeSEbqrw2ekx3oI1NT19YYPJwaPwfD
rnBEZ7P33OjYDdQ/B6GjOa+pyJy6+8IxXBzXyk7vlf12Z6Xo3BSWEuKzZcFFkEGi
F0PBtj5zcGOty2Xjv45k2VT4DyTWD0SzDfyNnVJdut25XSgZgPhKyLjItnAeoJ6F
Fu050HNTUxV/bX7NW3IxNXgAb2Z2Q0Tun1R5rMr1CoeouwG8ooV8AUcipa4iY9cK
z/YcZ0d64+1nZhh15lhtszEPlq/AutQRTdTlGag/5gRmVfukXrTIsdmnEy9Xt2F2
Oy67gSrm3xaj3w00OANcXENz6iSec1detKb4SQUoFqpueIMngd9LL6ZpyGF50Zi/
6ws26WwizzucdP7kQNHjd/I5NBRkAMLxy14jwiXcLt+JRuPu3Qs7+SzkQnS5F5Il
ztpkREVZBuJKgy1H0SOvM/DyW57isKjl+9EvIYzk49whqQ3jYDEStcA2xDX301sO
tjBpA78CK0dTOUb3tRBTW9fxTVWl9tsqC4X2YT5/FzVClKZrBGHl2n73U9OGJwwU
30vCfG/8nnkAosFjFDa0iIBnFATifU91w4adWfbzX3oMN+EsbMOsKUS6IhaBpcU1
Z29aW5/v3CqG/q3+aOpLvErOkKD8sNVSUo5BMCFpmdqdbXc7NCrV3N5nvVEzyIQn
N9uskS7jPml2T2Kz36eGb829c5/yr76JYBMvZ2Hm9OafR6Yor/0OgoFbfXLKinlU
K4/RE6PBDDyl7Qj74u6CTcY/A5lOr4F/ASRPwoHXCs1W6x5p5WKuQAzYLwblniM9
r3RVUjbbYlWO2c2uuLMOghCbFfKEcF+dwwGaeAT+F4J++GXx+DaZMd1LtUhZL/Iy
JVzao05sBJJU7Bf9M1whQ52vqsnma1N4cQlXYqUb+Pgy4HPKP6xaoaqA5ed+snkc
m21u9AC1K2nSFfjuHV4ZrIrXlXvCnxaTnMcRB3Jp/ntH3t5EnJD+L+4LfoxHwQpH
cz6NZTQKkb49WGG8RtRGBZiQrl36NOO3e/5hgrNtVoYUQ/E42fWtDCJEB51rBmFe
pF9fJ5FRfXPl6GZvd1oBqEhcJ4aiPPgAYvn852LaIGaJcTUtSqW+Pz8Pm3BceoYw
507Vtt4oi2z8uoESXw2dlc1KuMBg/jEWCyqlUeKz05wgCx8vIhVy3CDIhP1/CAUZ
E1gZ5UNhr59YlmMmwnIif+nPhqZTsdI+mhxieD3NxZcO9YiF9GxDzUwDioNutKhn
NmkWAMi1nYZCAATEwJxfu4ItvjxdAI3zhvbSCsqwYRp7mMFbmxX7kni1fM+3Noid
L491y9kh/PVLHGEne775cOJ6mWkvw1sWGnNlfduR1QFJu3W0Z7ouw74C9k/8Ibc7
L1glAo6Mk5wI/FVpaZD8nzKMQRVIWI9GJMiNrMNp8h3lghEWyGY6OgcU7W5qvM0I
aACBvT/Zh3LjpQDfNxTCB8oM4NvQEwcvQV0BSX94NHUuZaHfVo5BwHQkXxGV8knY
S0uJEaI4KnfVilz4qtslQxVvhUlcuXosbGPC10Y1ntwivDNeEIeH6oY5nPy2VdNx
mGPBM4osx+wnksHQvLcIJ7T/lzU0fbwyMtR9kkNHROr6UoFm7s35EiuDKsubZbnw
ahkYz9KhlKGdvWAXl/Q4HP/xck/iM7lxiEGs16IuvoFaT7U+0V8E5hidQbEYmVcl
nuQSBlWNZBl9JVDtU5eHlV8aKyJI2tnhi6791qI5ywc93J86BMfCtygxJGc79qZI
tMjsjhj2V69X/OS2uS+LGM5Nu1LhFL3wg+uyOMhu8nUwJXkKJ3dpYER9CPMl+iJW
XSlqSIan3zOwLdnEvGQ7+CFWlxt639wwNf7g3/COYTY6OLTZo5LzBhocQSg9ABax
Bt8l3ILiHsnKVbVrC5cB+djP8Gu+W1uWBvHqxVlRtRNxTOhk4oQ+XAGtSmOsLkCw
95iuDtv4srsN7es3Ch6vqk/H5K1cwekHQH0vMmGwYNk0Cjr1iYEGHeg+PKBj5L6J
XiswniDhW77P1+XydaE/vS121ovrMTZ/hKqf/GzoYJCZxmDVQC13WfnoLiyjq95k
2GNUT/ZLeeyLByO+dYQrLktwAZ8QPfGFBjn/eXmZ7Bp9yIXmklYBrPHscuuZ4bx1
2LqR17nr7iyilyTWZtJhrShS97TtTJgxGE4Au1VJCYETj+KvbfI+ZnG0GN8mCbbd
WJfBtAWT9qJHtZlRk3H2fpY66Eh0AUGAq6+lDoi5JuG8UeJD6FRmrv+ZZvnxdd//
GFerbInBqEfy1FO36RGjcyzyEQV5AFpY7mNt8WDOlz1ge4hD27tLwJwb87+0fXNh
lcXjeLJTgibVfWv2bccBJB+S+kTLtEvhLwdCzCl2Oh7QpEwjC/63ZlEP+8oFAhyT
EylJ0AayCjNykoIOqaOBBFdmS0W2IMukZwxH2AleWW3cK8Z505g2AfHjemAb/g51
PcE6UTsBoy6UpL+J3tQOdiUxGtymuF7pIsDL6My9jhZIP71IPousKM3YgNe4WekI
ZqLQkxxyxo5XhJ2pRuT4yrn5qjtGh0ltivBOdUYE+uitzy3/xP2X/kiOzxbS8Dfv
IfUYbwYB6+an170OvkCY5+IBuFPKPbpHFu96Ca+BvggYw8nnpe1oDvhwsNySg967
ub86r7GxOMh/gYa61s3Vvbm/wlWAXEAYmLiM2mXuaJ48/79zAgif3xm3vYCNQ8fi
AqTjjCrE/gWNvUcw0jCVsgA9/J4P34GWloz8CWIIiPQmgaSOEYNL6v6TJfYhsr1j
WyW0B3eZXT8jJPX5BzSS03pI1XWI0Oux7JfrdHxnm5jZfO8SyetiHukVY7DYxTwy
WMnMb+8KKuucAE3QQx7kZDW904P8EPnfiqlDjFXOERgZqH86dhhrl34/+8cNkNwX
ZDGUTLSHpwPzOzlRRXhbNlKpMcTzEq4ZfQj+KnaDX5L4bYsv7DUVdJPFEaRo4dlE
/K5U6JdFdx9WGjAHQ4EdICMpdaRGqbwZ9ur8mAhmNcpNLFIwoVs+w3WJEywcjq4T
7H0gvbpH6ABr4GRczJT+BBK1QRjWYXFXcuIZM5LgvGVMH2qdFEOEb+OhEOYlIcSw
4bkm66aLv8LGyBwf95/CEYR1e4MUD5bOtmqE37wZ8zcAKoPsiOFE4hu8BGhZyAdi
IJsrsxGAPImnTDdCDSf9Cexxb040KK/CI0g63YjyK5WpVk7Ozw6u0YzdLslOUcvx
WEjpEG4W6yKfQHeDS6ZicLHpSEoTlXMGRuXIo8L8OhjUXZpaAbUYxpZIaqgAD3S0
ZyTri5SQpEDbZKxU5X2GMPKaZazEyd5t0gMDaV35BKcJBzdSXNkIgAXU68JrZJlX
O8bQH3D/I9KI2d9zOicou2sHsw2AsIrvQJPGwvK90xBaZfzEhxlIQ0mfSTmrQXj5
L+I43Yk6M5CdtjLzPgUcd1Pi05MwwRbVNGh6kIrpR8la6oSL0oAS1LYVOsOtx1RO
4shbcTXbrjkg2cXJ1GiQDZhXcmADLQHISWv0idTk0hhNAbne5eyOoeiNpOwOIpJ2
js1SZrTmgTgswAuBewgNogg9Lcxz6VvmIYJveGAk67rY+Y/QwY5kKMdoU1t7yR2N
H2kaHOKlVOOK2B513/7xup8yCWW36BWrG9zMBr7EPorUorBkH7URD05fLJKVE/rv
De2vlD067dpMAVSCFy+3imyH1i6Oey2WNfw3k8PPstOKbg5fp11BAPcLB/YZiYW8
vaGm3a5TNbXBkttHye8YbQ3dacZt+cMcF5/QsZvvM1Us6kx/KYfjrJiWfDmF2OXa
Pw3rqezTxu4g/UzNkJ3CsYmQFMuxZnJUSOwqhheErSXzV55W1S5aLq8TH8RW2bjf
+QFBXFOR0wTCRrCvSBpvip9ZV/XDxDpIfsUl3cohbSi/XKOh3/MOJFvd8bIhgrKx
P/IBl+iOk5jiNRbO5sA2C3RmdjMKRPMlk4Mo028N2UHNrNDmK47n8Zz/7VQgUk78
t1xeTVrr74HUlIy0msIyiuQP2coAbKv0wGwUIikf8LUbNS4LRrZ+k+XMZcOjyGeb
2o4ue2fnqzmA6g5b1VVJF0rPfkz2B+1K/Vv2/9YudV2H0Esa0K9nWQkXwfvshYQV
GPQ0vvKVm+TIVZ7aVEnNTcGCaOZwuixRi4WLQfh+/jqbE327q4qQLzgtQlAIgID9
MNjsAn8LrYuPHRzX1vbbNPdnjSbrdjumY+L0PcGdMfqUsZuCaodsfW/mv/g5iIt7
0TEB1gFMMpLvEJ9CqcYrRjrGBNxziQS8Cq7KZzmnt8ZEPnG/7n1hPq3HwZRAP1wG
oZcWM8oboyuJ5GaNqVPNEIdgaS3ijxYg7KTd8uFzHLwhup0jzBJmT0m/PgZkfp8W
DWl1RmGKhW/ZMeByL4FLq16mWqY0gqRXIG+0u74Jewt9LVqHctrKC/BAHBaaY5Vj
xPVa2uWe+dZSRItKaP+75NsEoHKwHiStREZ5TlQaH1A/GVDGUIa5H/HZ8Kd0pYFK
z5l5HfmU7BaERApPzfMbcZ9tlgAAMWvpelAm2L/62q7wULP1+SPMkHNGPW7Mscp5
ltQSd3l8i9czUPk/4IVzn2JnK8ASgaZrIP/16aloDmT1P4PNkzXocS9OjU5XNZRX
MBWBJD6pXDDq4FxGZuJV/3m5J2Vel/0mZihCzKoxMw5NJoAykOHAarlXJbOTfmSt
rNruuJ+cIvb7rlr50ku7qQTCiL75abYKnXm6/1Y5U0h8BAje8sUq4Rl0VTQKjpt4
HiPOrmfYg7MG6nazaj5p4nhFQ27k3GUmlQx7IRs4Ra1FVNuOWoqdOsMPJ6H2AT4H
W+BEeDvBmujyrJKAQlv2vyjz/unTpq+D6Y3ALr684ANwY45DgvjWu6jL2iV+JViH
Sn6Uvnzhev6Tb+2oG0cSibk9DpMkItmJmxgTgPCQ1aChYlgM5zYuW6s4Uwt6YGAi
D3yQ0xVbaiWQVtgnyJ/507z/aqr7MzM6YUDo2n94Ak0e9H+I+BZKQMX/9Xi9t6Qs
5xWbiHrLxZei7M462Nr0MfWIk/1Fp5mFjfv02YhaYuy8+GbmaKRazaGguQXZG/1E
bB00w7nNp7BTOffkkMvyj4s0zJ/AnvjmQWe8XpPyG1PVmtOS1KGtaHUz2+DHR86z
c4/pbBXCcPt0hSspqJa2yShbdgEbGUrISL7HddG3FK1j4d44g2E/trPs87UVc/uo
r7l+JHTHYUaRJj9w5cuCROnzeORfhWgIjvqYV9mBgb8WMGbNdP5vuCq7DoRfWV5g
lImkswlkOVXvwwe1E3Mns8+fsXvX/XEGkme5kkZH9R3EetnT02WT4JFaSiTerzfl
DJViXqNTEo5Cskf3QwL9w0L5cDCWqkpfZCNfPUBkUXwH7hql4LZGaJxqsi6ii1g+
vs36fjrJ/vuQfEjWIdXjZcrl0YY4nlgqw7L9vlxcUMgmkXv17GZx3duh4wd1xVbl
Dd8eQy21ptmL6lhTIpGtcQbdXF0hMirwlrnRb+oEik0zui72r1LQ5zvk041/H0KX
HVBjtPxhwHWfNgJk6OejQ/nLyQeLb0dgUfJ102A599P6DJQgGnTIevCStu4mqUs9
jQRyjqPdV07k2it5qYTHu3eAhT2cUsd3uPDZtHNL9ZgJetv2dGpEDwP/MuVrKzFx
ECcR9L1edr/M7ctwpsrCVjlYukiuQMMORRpQ2xE7iulOLev+m48Phh8vEFHGuOpm
Uj3J+RXKKARlF4DkFw03xqcrAL73d7yFrg8gVsD6/ek48IX2e26H2j2frvTUMSJx
AOGXLdeCzVCP1aNzLAI6IUhqi4F4qmWnrupJkE1nJm9t9uHa1fIex3QeOOUdkpN1
GBrKWVptcIECciVOJ9BYLVzc6On2rIKA8sKC9QuJdR67aYRX834rOGjlGedbchfw
7BIvcZqXp6/XHhLFszVr1zU5kitxLXI5uODBpwrW6jakz4FaUF3VNTTp5T9pjqGy
RMqYXRuILs2s4ZYl2SQXSZGiipxnWoMIr8ZTdReySKFhNDWAD4hmubOHdtPt4ZrX
4xRLVHo+QdeNltHcWyPp7YWCWdm96gpMsFkKd+UDb9YXB2Zw7B19vU7AnaIwjg2q
lP9huhsqVKUDpwnsTysbHbB/ArVcHBdcfXTgFx55YEyvESmK/tdZXNehEUMgAGB1
TA8kg8Dwk9jMsVxVuLT2SVZuP8SK64SZ/JyF4b7q7uiU2yLfRVNMyN06kV9v5q4Z
hpG7oypDffd7CZY55Wxe0hg9lBrRaiZOAzuZPS2SnD4AFzBneEXY9wZylmFGyN2n
nYjakjaMU9r9c7DtItvY3V17X6qgao2Rs9QLl9hzreVpad8ixRNJI/q/B3M+vYm9
zF2N/GMVsGSH/Z8bR/z+CLK9Wmfr6Hu4tTzp3UKRTkLahzxjMSBpUStAQEH2sThu
VcT1u5yA3iXTe535rFfr4Jdq4Z+Yebb+YTBMWvWPvTgiGNeZbBOGN4a/8iCtYeJd
KqlY7w+GGr8N7IyLf+fM8MbsOc87jF4GiC7gMFyemj8PNeQVvfTxVphPdPoYqC6Z
B5WT0aFhD8q9El5NF7UHWQdGGDQRt+R8OPiqIVdi2XcVyolPAdjhbO6IgeIO5wUy
+JAKtmwN6dIopZJnSV1P2z3kz2GQ6jG3M7lZ9N8Jy4N9JEUJXRCFA3phTCA5B5uo
79fXlvnBNCRXdV12j6gESFiCVScfJYkYCRBKWVvxh5W9BGcSHwVRNj04Md+yLd/M
PYW17VmT0MMor+H+LxcGmWTNB7Y7os8VtIVkpihafailRacrp9HAlMzh55ZIUqub
UaRQp3GZnZgBaz3/d2YhAvYwpnNxSYmQaq2S8br7b7iR56uo/1NSVaXCkv3Kh1Vf
cdcKsbh0/26fj1v137LddsLX+lRttjPvqWwF/G4xw+sRdoQU2YYoSW02djyKmHS7
jYAOy/hk6qZ36OHB2WpKnwFOBAJ/GsZ6+IW7+kHbXxw/95vQaDM+sKKcSICBmCeF
G3YFvYW1a/a/kRmfozFLJlpMP1u2QtIn2MK1HafJYtpSxc4mWabSBElhDJOIhkoE
ieipp93t289giy+1DU/9TINFuqauxt1I9uMczUjavlxd2g6hQkVNITJ+yKaGaWbj
CRP8svxov2CTAebK1mRqas2tb3gX8Z51Fr7NBye8aEDGIbbh2UZOKY7aymv2t1c9
Ck2pJAQGyzvLmQZtfpNiy8es7x3KG3ggguJQtjg39bFYQnOM26k6bxpiZQL6PWVI
xU9yugLrcMCrC1n4TwOZr3fZfu8SB5zkwRBZsngzjw28HCJudzM8Z74qRDzRLM5e
5GVCELw+lbwSJ2zKal+w2RIWTigYM0eSnXakcfoGxSNvV1DlsQ4FwAP4vLYDImgW
hR5rHQAXdIqn7wMQNJEpbDTkjKWcizNR+gh8K7iQH9/+qCAaX6g/ybfvYMWRbPVq
B7JeO8sZyLR5g0hyjggWQuLNtCgMb4TFtQ+sJljuV0iupt6K9Zb0jpbJKobGpV4I
r3ekcWnbjdYtEQKVawByYkoM0qmcMMXkSRqUYnclXBIDC6UWyAaXF7S7tju2+t/y
7nlZ8Zkq8FCzlGshyROgS7P+t4hG4xM4LhS/FrM/HVn3s6p8yYnoop8/d57UlzT0
z4XTU9KxDcNBbRF8x8bKoLjECD4Vm2QNwvjuGs25zSLzY/qCzsccBIOCa9u+ec9G
q2ts8kzg3+6R+6lymm8KLfvagVrc+IX9tcddBc3iwVa1akn/gsV7ZyS7GN8kdlYd
U58AhutzHs1ncD+XnqxJnMGVsbvIPpwcIRHh9trtkxNF4IPjkdvQle8BaYEuJIE2
PhAMO1jPJigKh4waFnTEx6SRrBSNDVntDc1tZypGWA/kpD19BIT6qolVHYjoa75q
r9Jr7w7tK6La8K/GrWBdl6PbwQCJ9xkgpEuj9B0r4tHwiOCTL1d7Lv7z4ITk1OVT
CCIPQNAab5fu0KRFaGYB6NiE9rEiMNtJvZqfD+V2yUeDKWzmF+wVtqMpBQI2PYJi
JKRYyqnD73ZNhl5KhUhZcQeW7ebmhOAhXw8psdsX5HzZAF+njsCqi/JhyvrvLxRa
My7f1yvDO1NYkgRmMUZCHa8z30oW5ci5Sm9+a2bCnUP8ryyn4GvD6OLbPwug0qUg
AkdoCI1FD/5UXDe+nnamBGRFQ/hX+BoKQct0YPZ4qw5JvSgsXX6OVMuQkXVhNwao
I0ewX/ICXjOdh+90PwYuDpfCRNq9lo+Q1JkaGRuIZ7SxCP7FIaewgywv0v7LWuy2
jTPupLpN6ybWSs3HBIjbnDhlonmeJEq3IdjKjrV/lMcMdQHm3OvJvhqLwCfI5yzw
c+P7RbjIcZUOaV4FZ1u2W9vyG6rMPLBb9GTX2ZTaaleSoc5QZp2wvoea3js2vzXi
anrI7WhErDf8xK2ZniXVC28/lYT+hNWCJVGTX4lIjAaCqJ1RPHU4rxz6Bx9zZrwt
6GOQD2wGe2H/YTMwLsmhgPSKwn6h22jXHgHJGp9YDffVWMt2/2AN6vEAt9patoLn
r31xRCpTYYTw3r1m5XM1Yx90X9LCyzLxoEzbQ4KuMjIdmErbHL/wZHPNBQPZb3mC
aTApqF3jtq0cxL8p/Ejn68bfrkRjswXkVH9yTLY9eqL64WVOgAaBOYA/zP9aCNpE
dAHnZyXwGIku2B6SdZ0mcok/GETVg9WxFdVqjHK6haPMmfixlvxQzV/ElvWnqEUI
63d8TzUEe9r4mvEtM2X0qNWn5jGrlD+V0bjBz3tgNm/LGuL7PW9c0F4Kwzzm4u/g
yyMsWU+e12fBwz+jlW6Lw2bT4p9937ie5r79tDFuoV6itaeXIfG7leSp4XTHoMxh
LpVaH0gP3bsc4SEPtYtUH4DNnCve1nWtsI9TO6r1YfSAIuJ1hvFZ2uFwCrP5f1WA
6aUPouVyKFLOV3VDyDSDHt5AZS6nZD+WD7wB6iAvX78as/Df4stmET9I1wMq1p30
mii43iBHmqGIArvqteWXd2tt9G20RjdLQZ7nVHkP0WwjVz6NEZzltUCm/S4rQ22b
sV+FuoLiNaKzKwx1SiuY0GbsE8ZPPxuesJc+3FGDRq5IaE0QwMzQGtr3giruabNu
RMJU0Dzv0XO5sEVgbi7H+HqaoVKd0mN2VJYzfVE9vCYTMg8sWI/tcF7/GTcBJY6V
qh3GoSr3RM4elBTUlwXCPWKpWcuBJ5SjtHznFhy+dbBe8iqqorQf8bLkvkRxKtB4
vwY0YEtxZdqjUMO3rS67NcFOcij3SqG6HooYSOHvygOgxdhNMMMfQC1mheGVk+SQ
BHqe60/jyCDR9/Kaa//uNkUATw746TTgAMVN9apPU1WowMnD1cNSD5PuUUx5SvCs
2KJXR0MYE1bxVNexFPvHN3qZUe29wgGk9J3W1vW1BJgUTcBzLMUYZgzy0rmgQXSl
Zh2mwlbaGyldzllBkrbYOUruNdymjhF2b5J8KKeO2Vg6alWLqPvmOGId3RgEBbfP
sQoH3cdRmdFP9N+s/xgCkifOQL4N2FIkZPKPPz7XjnB9BRYzM2EzZFi353bkbrQG
GXHNOmY8uxMiIbHgRSmbi3g2mOfxCociHW1jXXGs8pjwgPIrfgy3kyZ296UdUPyY
icw1AWtoZwO9mt/Fh6fFP5VeGt3F++qtr3eKfMsZPVToJy8c1mI8iKOb6uobSwiU
gYL5Ph62U3+doqN4k2lfxoKebuTFd8h99XMXTiu3/oNmzfP0zgntidm01E7Mp7oZ
txdYBBP5ncFQ1Ud2drkw2OaZy4AQ2wwYk0rJT6wd/JKUYrdIV37EUA34vHwnt6Dk
F9lWVZmtJPBKj93t0OfcCPy4IRjH+Yz0ZZRelgx0rirWRwxnSR9dhA3qMyiy6bkp
VtDGXHlyPO/Gw5VaCz4Zusqnzr4hILC5rsNjd1f/MNpwu2E0pzMYkBz13DcMM/g+
uUlfXUbPwRyZC8fFwoJfQyF9vNFzx2C4YTpiQA9NCOuaIBdN8BpDX6bltO97QT/e
igXnRaHwypRI8UICz+0RFX3o7z6Ra0PBeYqfvDVXHG92X6VHc3AfaypcwC3h/Gn+
s5aZX1qlfkP4vsqd1Ac/mauabPD/VumZkQqlJogEH3Xmv8iCSg4TGkykgKEDPkrO
P9qC3ANLfRcg/QHjQxZeRaZ0dDFWVsjG8bDAbPVhqofZ150AUViPu3YI2TnNc5CJ
1nSFaHrocII4ZQXXxbUIjh+kV9Llf99lDqYjXDFFiinr7ylGiBbFTk+5I8aod6Ne
G0GTtuUCoMhOULKtMYsR0/7tQVB7qLNQqVEzaMdpsRCjidvgM35wBUELXCU1DBsa
UlTrYH+gPh6SFjjqiTjV072Q7slkxDO2OjZJXHe0xzBCIgiVpBcDnbQP8zDaRvNd
jy9Hq6QDSNj5rJrx/3Gsed7XolpGACFvsDY79JcQLBrBJ1VT1DYrzPqJRGVgfiva
HIMKueqmWVpxUexpDdEf4j2TjiW652OLKokS+Aok487MgA5iqe6DGcSDKBV8cKv0
V4mafKpi9Yp0gdqHJdi+DW8IvvIGoE4wzhYJEUK1qFJc4PMG4NSLqFMg2lTKmPJY
L05SHlzt6M7py/PxSP62eD6fqoWxIRtYZrItlKMRERDMxnm86Ng/tfoOgFgFFzTk
mLd+TgSYol0DSDOCTAEVhxBQBsexEHDjjtx0fjx30qtJqtxW9M3Gg+teWxlF0ksf
FOR5XFVm3ETDUZJ/XZ+TmPbWLK2iHqBp0DVMFvVE9AOaG5mmWu71SgM1AF4R4XF3
IzJvCneVs2uVmjih8oV7eYIgOu7pmjRhR8+MRIsrDWSOX2ec+XMyNZGP6MWeUL9/
Hms8SJVQk2QD3mcexKc/kKQWI9oVA78f/GtGJp7Edl+O16i90Cf0MoLHHD90S6gz
hqXVcK96QGi3tQKzPlCXQUuzi3sZjjMvnAxj2h8nRyb24ldofVK+EL4k+oHAKYCf
oOx3/P+3heh59C5/XrYTcDR5ddRiwVq9A4I+KJRwI/yt2bidUTBjWvsY0JkZtV/e
vcJQLAnFQgHopqw9Wq6kn6J+PBsdJxW9T50x85R5VapgTQm3Y+rQf1kB07c4264v
Eel2O2QngZso/Ma5aDWIxQDx+H6IapwwM7HzuoHVEawKHOZ/13qmGXMo/f3zApq9
VhXgGoLiDd0pOCaYm0HUTdOTPCRwYI5OVKiXhvfWrepJh+HERI0zKmCZBsooLJlE
787dJCnIwFyC82IiDr+NrzmEZX0yJKJHWl45or23aVTxgcUX1lDJXk0v4kvNy5R/
M+u6hkudLRTJyKXeuAkNtIG+l5FxR/JmY7NZ5xabfrNj98E4mqCsmJSJGSnz3IA9
Q3kxDXDJVImG1TFpOWVanjqKFNcaIbsT7iDcJuVE+33VErKY73KMmfuibm5rkw55
vHYz7S+CO8tiz1PfudEcMrKxiD2dIqxfjNF7yFDKY/ngm3QTcc1Jjt1ljMN4vi1U
eqSjpBehJi5UaC5k8Wn6cPKavMWtk7Vtl5fPTh0VH8LPa0MGFWYLGPkh9e+g8PDQ
RyHLzvGJ92EThTtm92nDh2cwivscVAEyqLripR7prPjiRq+8TbyTobhr3rLJA6oe
PRZjjOdperoWgxMPUndlPQ4IbTsob3iebv6pfdnt687S8CB7Q/6+fj2wtN9ZX5ST
tV2dQZX0Ip6dFdBaOw1II9WDC2dCzZBbgInJSfkp7XUrRJ+B1YsXMCy47SFv9ast
fTxySIQEdGJmgHi06+wiwebBrittloj091HoluMrF68qZFuu5l8FSB5CgSkvJqQH
Rml6NddGr/CV3pvoJQ/pnZHBtzJLOhRyEOeu8O+4IWiESdbPJkb2/ixVq75Zl/g5
wfNCDL0KaLiaedNomICzYgDK0oL73GTIOxAFIfq8QDai6YZx5bKD6BVxGeEhGE9F
ZXpaZp95U8xMt/I4ZirxdHpdpYi826MtUjwizVBScrCKj4LR6zj0Dwan14faEVaS
5uGgWsU7Fq4DWv0a51MzzzZ2+k8lFqgJc7xhTCxlS/0f2nG1Y1PZm1jNrXJIk1nT
pzrPXyRwlJGP7+IYQMptmITIKuoX2T0AEft5YThQR+TlFMKKyAQSLwNNIsm+GxTL
EuK/u+4hikIP4X9VXYi5lChAMhI08L/Fn9+vN/b/QYKXTDTbs1xLy0WURb3sxmi7
D5wsNWYbt+Tn9Ls1EivEGQsIkXRw/FEm0bpxss+W+aL8a9cHXK1RuEGBJbYoGmDK
oaTO2E7oEeMxQ52aKeyaTjooDAqqmtFXvxeRXoD7eB3l/BSFGQIF6PGrmb+FUqB+
Oi3LPXKlxLZ2+grPb9op1gxQRXQLiDXWRLN+IQc6tqYOPzkl/lbv8kG4foZldDE0
XGc8J+hq0Wfci/AAJrhXENKljuNadQHDX3j4Jg1J848xJOT71EOFcLV27pqHvCe8
9RPXmDQ55ifcB/rj6QIQ7rNsdc/1vXloqhUVEghb7IuObfRnL0to8P1WkxThSvrH
bv7yu24q/W8be0yngoni5jvKOZ5NKCKvtgHGohcgCQK6vIOPsRTMerOcpWk/Bg9+
dPngIMzGZFxmYu/k7eLgava4H3k1+6BLXbrqiyi5SZUqind0Xi6dwpRh/BaVcsQ9
pI/SV5aqX/1xmhWSxRFpTP8AC5blsR2RcHsnL4kK/7yc+Vh3krlmizS3feCqGxHW
Qvw204Vt6tEKVwAPneRbqthH8nPYWmwBkqauLBQAeoOBYG5obmvMmfCg3aNXDwO+
kXTps/k0hpn70GZfdpkXwvHXVIEUkqHFx+F4TfWXctBDOnqdyEUvU5HPtGwlJP2p
AsSn1+IKwzCqpnwxcoKO6Qc/w9j4u7i4egNeDkQ/iaSNmVgsObsi/rvamlm2pStn
5wgoT6KaUiXofWhL/MpFvCIBhmjQaHPr873TV/qrZhuhXRPk3cS0OYHvQuHc2fdT
YCQ5wiURiqTj5HQuyKXeShYcBitbCGTYkgRbqMSTho8Vy80Dy5WRg0wBaVojKUzM
x/LMuLstHPok2Mhdcy2UvYt/Pjczz0bOxKlpWpIsHIoghuddu9pEyBTEpcSyUG74
Ye848KsrWBKoGufPLrc8hacFdGxM3cN45ZErsXYFEVfY+mjgCI80lQ1qErT6Jw5v
xN4Sua9xCjSdIjpYQ0y5uohuTBQNocUWIegzTfh4WCdx7PYG+nThvELrTJyJov+6
Yh0bAc0UupTv2NVdS6UD4kn1Fmk0drsl2gZEpUCnGDGVhRAvdGlG/4uzetEd33Eq
wFqr/ckLcCM+6Jj5mGNiAVgC4MRdjKFMZJCwfeDLcgcXVo4ybopZdC4jC6PyHBYa
MZfg6RL2P/XFKB02w2SorYGFEnMIq+2TkAWnAfnTjq4QKqWbAKbHuhBbm8iVi6RH
qAdenh2DdpTTaG1PRiRxMkjiQ+d0YMuocXAHxdxhx4jd6IjzYQ4gI4ZG6tu1WYa7
HntnG0iey7eYToCVqO7SK4hb5vFwocPJlLuKnD0c18Tj/ww3HkE8VkhAfdu5mDpa
QRwrNgDoUyp5RkmxCFLvzd94VrSB27Cm+9KIs63NL3YovSpLEmsR6acYmohNuW9M
p4HPi6S9/sbOOnUMqaBbbdsZmi2u0cWXU3jyvfWW+OhaQTNka2uAV/yvATflHPNH
aXL3iYjW07zOA7HuUFH3qA2Wb5EvNDf4TJArHT3SlS7fjgXRqQAYJsfBjL8tuwpU
sqsOlUHbsZayLyYYvMrbonQooV1rea5nvlrh/I4h/YO+rDgFtb777Y6c699Pmnn4
SWnwgj/YGMDqpe9onzb/i5fUky2/s9psWS+gaH12ccFWq8Y/Xs827XPmksn2MjEW
aubMhh0h9DnvII/tEX9U3UTclvB09ZHkocxqUGfFRu+bzm61+Ht48aq9r3GAdc1t
u8odv/s1SYymxZyauTSNyfXnHdvhZ0Hd3ZVylOzDDpca69r+tk9PQIDu/XQH0OBo
+Ezx3AS9JNqeGG2jBVGc9FDZJ3FBIMdV4qJGudnPk6mW16vZrbT2NRQdLfg6UK0s
MjRMKl+dSfnlkeClb3lOaovGQH5gAjZDVs2QHx6I8K18pMS6cC4GWrjXkWb+0Kdp
o4JxRp3htBxtJDAEeF72E1zRiODKJY6NEYqJv67tPF8pmgYa1MuS4nGCkRcflt4O
FNk3k5WnXneJ8CXewmHlJCSXEepVNVLsPxq1NDa78Hx8AEI6QhPnQhb9c+FjHLTA
4O3n+bnoY+Hbh4yhJ2yNqDYETXM+RFnTFevyPBdNn+SHu6hRVi5zY79sGltOw6xp
MQXUjiQpi7hN3egSQBLVwCmNpfNGGhK/YWqRS/iI1Dfx4LDKxZ22/2cNsnivi4DT
ZZDvUk3dRUWvF1KRLQQNg/pUNCvN8RuYqn5NEl0FsnXt1V3QSsYpLIliqiBA1gg4
AGfGTLh38ue4XwRRK1QJV8XiVnXObZsIE86/i7HSourp/AlUad4vdZpegl0kv2/f
0pyu8J4UJWQuuHdo0mo4hKZZkPRPLhj4GiyTiypKVeIe8dIpTUXytNd3eKR/VEnF
gslAqmHNjZrOjyYaReWo52J3finxvS8qT1Zl3QIIGn3WLWLhjPeK4ri1ZhpQicJv
YZEhuZj77BDgg2JvSJuK+ZUkVVoIPxATvs32c5/iLZqFL8dQfRUsdrBUkv8iujUV
NPeMZXRMGFrIzi87sntSWb/giLHjqGlemaaLRrIjONnszlQLxMrZdF/PsWFaNVu+
8kiDY1BxSK1px3euLunmuZFxFHklNFhOaCU0TGUsZmVuAp/jNhV9ULHUiMMcl+yS
hRdhZDwLynKsOxYAfisIwqIatBgGGsBFsf0Tu7qkA9L0iEhDhLf+M3V3Ua0w8C1U
qqP5rXSMZQSOXKUrVauAPBwSnuBJ+rPjssc1w55gSmwaPrGeDB8DS577y24ws+jX
CrKQSkC5YVTDQ2qt2MdNe+CniA2WmuK7gBEZZMeGn4YHscyv+lrlTn8qoderAfP3
WnpzCkdr/SN6oX3XKPH+CVjoyTof31JxlLz4DpTQ8YFeyWzIxNozD0bNFLOeGmLp
Ky74rE/3xI+O9feZU+q7BRK/w5VTQAt2pHoPvTcge2k7+AbGLweiticzw63vmZ+3
KeyIIDSvl1Lu7bdvmoAntrQVYrABj3GoJuoAzKvr4WO9oqtOJ0At7ti8doP5vrRB
LXxDkZteKiR0SiCOyG4bbd6JJlnI8WHv1UGVz4JzOukRXh6hFq1OOq/mLYlpwI/m
SeE03buW7EKem+FOKZQPmQDXy52qf1X2Lvclnybo+IYVYEUwn6wGO17sIPLDAxgW
et7C4O+qW5Om/WSy48rq2QBSXSUibpYQJ4Inly8Y+WfMdHvjZA5xslxkFI6J0Sh5
oVT9+QQ8srkCJQz6kaQBIZZXCbGm+puYuj57Ve7sSQcAP2LmJczu/ML2HLKZ9+t3
4QpdyRCc+RPncCXGjDyQIGZlLoxqR6g89AtAgWDwixxgib1uekzbgZlZk93vKL62
9V9HGXBlC0jJc2QwpnC8E2vV6dyMyUC8Hx2Q0LI7sTHw6OafdfVo18/ifMFewxJT
IMO3dakIGo562hCQPaJJkqL7EZ+O7ndUllvTK9WrjqRAZ98S/MUhGvCc9eXa/v5N
OFRhJGd0mH6LKRcvjIdlFoBQbwEOC+Hbij51JJT5VTld4JvPu3ft85EH4INw1hc7
Lx8pn3/hB3vkgSrku+Rtdr02Gs7YsXvLMqrqL8mefXklqR4gWyxFuDcyacQtq8NT
sIWsowreN7RfSuL1Mx1hdxRBOknPk82mQj/scX+nHb1gtuIt+YIMkO1Nu+Sf/sm2
YeQyGCoqeTsFJJ9mmRCBZAgx3thPsCsopWeDyM7TDfcZuPFvMZanDq4F4QDG1+yS
eHrYufTtCvL2XZ/xt3cFYSSZNUEg1+GJh/nQlrE7158DKS2Pbkr82OhQMWIFQ1CU
g635zYobvZtGaRX/tN3EP8vPFrMNWURr6LfrUMujPYcl8socuVz6vHk9ocFRJ4p7
BBE0veKF+hWEuKF7rWzo2MdQRjblWPzQ955ASpliCthYthAokBchGLlrOCmcdixX
g72WUtlOSC5sh4MdjG3djlpRe4K327BDdl9ApyWkVkcIsUAXAIqAM7+8zHE4pLsH
UugXg2ekXMD9HCfRpZXjO7wlMo/2JlwyW/erIbX+sRz+/eJzprkg1zkOc7QEtqYO
dgW1Zu+gEVGprQujhwEMzixhM8axXtJguF2T5OTmPdxXH8oV9qWL8y2p6SidFpl2
/ztagYlgPL1aZwKjf/B15pq+OehmMdP/CdqIUIEMzQYgw5+q/mmpUPI/NlnYfm9H
MGjj97yBRhcfOyisYDN+YxTejUwiXILd5ESIXPZggAvRrJebpl/MylwL/Q+8Wwel
vWh/asPJrZWfsZ7l1+STEDjTP0zACj+WlOHCPWDld7jQTf3wcGvgsdAERm5wnOd8
oBpIBB1ya71JTWpCBWqNFtQw2qjd3y1glJUgVwFO49kGsHtYXHUPhFc/jwRC9gLG
jxsNPiBMWjlKLuPtJjSyZDHGsiSbSCLHEBXW5B+aamiUWRoqoCVgPqeyZZFxUAvx
BBrp4WhAKbRhicclCIg+dXNZ1+O1sdgysEIzrXXWo2MvHo/rDwCBFChu/fBetsFZ
o4oFf6EM4U7okTW6xSN2DH9KFY4Fx18LC9I3V7fEXB4B894kLGZtg9EdiDAav//x
pg0WTbmYXhMEIsFGSRaIct/oliBzQHTh3TlYQ77n3onI2drz3AbQvcxJGtKj86us
tgkn3AXLvqoIFc4aeaS7Ng3qk+BRINujQuclplJPJmG/m6zNNLkxFt7Kl7GTOO+q
1hq1KYwIVLoOThktxx7JxcDdaD+6n688yOqut0JbbcW2JcVSp4M38vIHBLGSH0qM
5atFmnDZK3ZxbOecglv/QONukKQt8bXR63stkBFhPaihP9p4Aqkf9AHlPFJT1o/M
W956972Z4EfAOy045mYhXEIFBfmF9zIOX3a16ropVLr2fsJOviDhf1B5gyxRzcOY
Cy/hsL6ViStz4CzLB6CPoc7aA9AKBHWeqWLHA5lX7qKG4CLm2WXB1jCPKUlaeYId
rnShxnT1UjnRqashB8Mz7riCDG+anZBQS+LRsREVQpXh5GVoU7d3qp+CYKil8LY9
VbvBtwWv8BQbluMYj/iZXjWnvCyhgiHgjj2DOVmA0e2aK1a3xb0hG9FN6Xwhe1qy
r7kZrdlnA2wZnGQRBz+X9r9/FAL5Og/L6Zijy6dHDPx8yjxabVGMqGRB6xCf34cd
0s3tntAa/TKn+l7OyurfayE0xrQY8usYAiCgBEHePNscpjYFpsuwBdeFc59jt2JR
BGdrmPMpcfqQEnZSz1ddRth8nx1Oy8+pEOh+xXDTl+tghuHx5GVUhWwUdYRV+ncX
qf7HHgx21rHRsCZbFGgXVbCbHNqH+bXbqz+bcO9ol1P2Ojy7BomvYbY8AHPpWtm2
mng0AzA3Gu06zHh5WaiCG/YySKPq3B53yZtRLDng3OMMIAQ2gu+Lc8ERGNguj4wN
wuqHzIO3gZ5vd6qIQMxSylPO4bVsrUTm1NdkMCOrhvsacCqR9DcNRhqLuTo3OTaq
oRsOeguzNka2LZ5HVQnReNAjkD9rX2M7eHRjfOTALcji/8Vr39Re4Zmyu1lg9rbW
aFWHhttdq0vuGyHXvy8PBeUtcIrJgxkH5jogTd+3tSRBn/fJbu5eWm6MZaT2rKn4
C53rpOhoFHUFDz2LjtIMiPHyBc5y8UdOB3BtPTntFBtqEuVUTcGRXZhyPHfurfuq
SUbnziTj1abU1Zm1yVCkq8ei2CBVIXxNBA4BvFmLBwbzyKX4mZHzGYlXwnh19OyJ
3i0SFkRHQClCmjU0s9bLUEPDmZAh5Jwezu5bzT9aqjEcLSeKxOaeJOQSeKLiVU4W
PGB4CYtLtjgOt1du4bDYwFr8XzIPqvd0QHgFkBnOW+x/oGcuphRa+PEq4dCtMh2W
oQXzD9UcRgExb2NfJ9TX4RZmTsqPyDaEZ9L3AJNdo5/4p4fy/7l1PQeube+5qjo9
zLiN90R012ZaN+3u+apqFRjL87URdorQMmRu8oT3hAYHhkVSjTfl+VPHdOt9lkhi
8qUBRj6PIfAQfIlZ5vgF5nmJM7EekLLKy0XCDAH1FFBjYJAz3yNAAX7vlOOTGzLv
t663AOiFTzG/QsGYpOul9bRtkAWHPsLQP62JSAG8ZEsRY9jo2P6SdzTa+z2NrBd7
ygqNPw9GnKYjc7O7a1aMUEYHA+EfkGaIhvdRgHNxrVawz7NWWVa671AUFwVuzSgY
muqgtvP2mHV9IdaPeDeASi0OhKqSKAt7oaunisdfORVQLF+zVtspGBp0Qz2Fg6ay
hrB2+JjgtuD+KLv9SdhOBDlviMFDFF3pa4Xo6nokPXMCEFYqKvvM6HjzApp35bfD
NFbx4epeLG9K8JAxgr/SM5/1fzD7E+JqVPBi7aLstDr0QPkWKMOZMDiSXX6BC33L
/OdRdFyahW3A0FDeGot9srYt6UqbaQ6jQFR1aS8PxNFbeSXlIm5ZSAptYSqthwzZ
DDmhYpOFu572WiI8WbbuKB7pAqwfXAL5E/NsuMFlsizFIU6Y0Dl+Ticadbt92Ay3
uM4JARJ12F5FydW8ofaO8vh1gyHhRs+zRt78etASZB+99m0/YfDPe3ESTLp5UrkM
CJtFw+XVC+0WZi+afq/vh/au+pSNfby4viPyNIm/KwCbWug2DGHnbFuT194iNarv
xfr5zGGOX3oGcx8U/dpiqTsvstCEmiIfrMr32cgttg2nQCDjXUkxKjjHer04i/9c
gav7JsPvRltOvsYMUhO4SpTTHYtwMeGO+Bcsu3Zf9/CgmP/du4ecSyVOD/0YHE/T
kIzNvlenS6IYz3lXRGEypwADA6wBwtHAu2kE9uFCF7AQqL5OejqgCN4oJFD+W4vC
dtcIVVKR4Jx/3rhqnlqRHzjeB/cBqomNGGJtUkm0K3Skp0Vaz+dUrycx5MGa318z
Q94mBjc6DJI0lGDHfebucTxkeK2N07dJKlupCS+vQ6v7PR2l4GEDTBJ8Hf3lhINC
BedlvvbQex4C4lqiwHROvTRfV/N+GeeiuTBV/IAe3yvKBhzejvgZQR+k8WoactpZ
0izqGCH1OWvTs0iDDMNYOH/MD5Zgd9Rk7GaT4tbK6qQWARNyMVpUNNWQxvkCLL0e
R2pMjuBZUtjWIAcdbmPehFXk9RNjiOoWJUx+DGxHFjprNtui0dHKwvqnxYMVeov7
8uymUbcAd97nAkAwX33LD5VdzvmgEC9xpwQ4bLtR1Jx6tXPq4RDmi7bcbOD0iMnH
u+2pwJj3f8UoFhu4rfQQGlJjZYKETCNUAzWr01lj40vcWU1ct/BWhD+kbHZtesNj
KoYca2Bt2ALJbwuEPYjPyafz5E9NPwvS+oyr/CGe3PDG0j6Va9ZZZHVMskZcK3SA
BTPgp4p+YwgNusjPAtY73HjAp+iZDDzyAjcTattBzNZfK3cacUZMwwlmfz9Vzj0y
zH57Df6bWCytrRCvhgus4sRGLQIeSD5nBsroYPAB/Xuy2isBqqsffF6AiiPWU9Q5
nS67+7ibHfBy7yUnE4jrNZF8ENcQK/FQMDccu2VmozmdZqBDvNB19F5SaJLsQjIe
yphl8F+0agapVigKeD7dgF8jCqTZWE3Dl1HhE2aV8TMdIHyX2jlMvA7pbCBVxrOf
aeyYY+qyJU9RuC+qQLpLqaMh5wvE7pLH8kI8zSBUEu6aB8NmJQl5RYMJaxWj+FlM
ztWCiXLTcqVCa8mK0F9NisscUL53Xm+Ecz2FfhaWSgP5lztzckbXiwPZDSKMUvAG
MaL0tD8UwrCQIg24jZfgsj+lH5L2zPPaEg61StU3+3hPfBGwNH3bbnwTTbTC2OM+
Zd02IbkdYmCWgOSicB20KVP1aiiLh00OnxEqnmad1+VUZkzM4Lp2GiJaHwTZEvid
8csc06R2iYDvTU6iNGqAevKCaP2Yg5fAidvpgQK5c3HEf1j44uTix5r9ksYO09Vf
y2rzanxaxm9y+cqeTE0NjAfDuZzR+MeKkMKD5DkxYt2lDn9QaLFkhN0wUL15pGi3
36QLEh6WevfuYgosqp1McfHcNrPT/+0V5YNG5Im3H8sDdxkm/rXoj3BBEtm2HWBs
kOCU1M3iSyCEADrXNeWkGr3ymYRpyrNKAa7dp6EXlRb9tsrUMhncj+eMkJiwwtiW
T5MImff7kfhJZ5/ZrDz6+Lica3xxkH+SiAd56/SeGIRY8Qc3oeTSJ74cjjvjZnA9
QC9pLdaLBoVTKZTy2qpL9vhWKMAXGyAUFsUpN7kk79x6+x6mlfUzhXJLNKoF83Hf
r79YrlhWmdhzeuNyTlhOdsyK603yz9dFmOei+7VGIUXFCUAf77gSunqYEliB0XsO
J0ebcCpXDVX/47bg8iQHRgcLvk+gx2ftAI84TZ8DfaZzeUt+FeH2t/rqrrgLWA+3
vTUEcP9PBUxdhUYsRKLISsmCQ0ihSFutZXivfkp4b6yLVMusSROaci0VzojFO8Nq
0ROStMQRkNS2zbu08EBZjFutZB9YY6o/lSaDk1O+08U0mhtPLcRPwwIDPSb1AAk+
d3q++7+F2fawGmKvIOvqaqDzk25l82+zKttt0zseE5dwxAJdpmtRB5YNJoykVxFK
UGx7OsQbJDFM1NZ+TUwc0KJZnvKlP5QOBBWQdRkzInDse68lCtCJDSUM9nNWLsTQ
w3gh8ZcdPo9nCA7jPb6sap+rIUBNlaucI6D6PZUvGDzqXAFVi0sLxGSGOiYsEDSW
dBfkVxSq4Xryg5ssS7vp9IYMcibLIRLHyYnM//JFN7Q9ivTxkKCgPI6z5zaFXLUY
5YWgQ6apyfUmevKdYRqMpyok7qUjgLkcEBxohysWI8htBtDJ0QwRwrZgxChn63yy
Ipe34HWAsN1QMa8lV6BN03WlyLQ9BzGQ7wP2BMHar1xP1+38wzdapNQsx0HIdwcy
4mXJhjL8dg3x1XqLufJ+7sEHQedkxjqWaAjio4oDIpg2+nxhucAG7MhdaQoIVWfY
i0cMRIy+S81DfEmg8wTNq8OJywCb9/rywpC4FdGX88xsTAArv9vuw9Jgq74JOr+n
u7bf2E9SH5KuPs/luvyN5AE/oO2MyiPC52Uz/lVwXmY0T5esv5BomAdJ7L9Woymn
EZQh0c0Un9FERHS+iVGBVUf/7gN4b7kUXRcul2SZK3+3jyMT7GTIOSWn8RmKAp+9
OzgOs6s/XvvxyaXbGdrceI17yEVH6VuowS68IP2Wj1KtY52NJqkWJZF+JTyeehal
OY0BJ4+jI37MU/FqIPSkGJgQidisxtpkRbPHMdA4/x62X+C+zXFvYex060abvsJb
qlv/fKr90tF29ilHccEZjnAOZDRt9EhUHFgBwrxeLEFTp+W5TQVPKCQ/RXPH/X9v
WxLs8ACx9jhkDDk+Dwg0tvTJL4+gZL3g9BQy0FRzjWljVzRLcPinylZguMTjTTIC
a2IbIMmQ3i+6hRTLFy8BOZxzPXlu3f6tHFYnEqI8aiOB+BPDZMAXZILUuzJZwNrq
4CDp2Soj4jXI4Nd2wCbV1NRa0gTTs/43or7bFqk6Qzm58TRCA4Mpk7JHZULVbZHt
scF3L8jI+Sm5kZMpMwuWQkNosL+L8QHTI1S/Fk1CJenR5OnEVtDhtVdZabdxdii2
14nm3DiNRT4DougS/klR+AtFBQRH+LR4vGEozFUB49Q0EGtR5PEzSNM+Hv3Tdo/y
srNUjHVaV6ojkWqfcIRtcYpm0NDyal+Hk9NVg3UFVA3NZZUjdvyDQpNOGGuVKtOk
uQZQA9SWBeiOR3ImssBy8C31Kf1isqizvo150+/9/sg15UKFVSmyhGHIP7LOZM0e
Ah7s+OKS/VLjFOhgdDuX37aWbakOj+LrlL+D9XKIBjRdaxrutaGn73wHpb29NGUp
xVQRjEsyBYVLQg6gNOEAnJ1/gCNYwJaiQ1oksD77oqsG8o0VLBIJ/CyDcK7pJpqx
tQi33cIvTrQ2c7Yt0pUtEKdnDCiRModZ2RjIIuk8DmDqjQG6O2o3o7LJr99zjWRV
Is4Lb44B/yIv3MAd0O+9RW7oozalziVDqErxTkkOZVn3hzZz5x/bKaBoKqpUsP7m
sS1+V3/G8S/X36Ds4Vo+jktfXs7SQ7LQG3CpuhvITBqlsxzncY+hhPqZE03MO1NL
zmNvqVGK2Wj5ZnooiCNRkYCj+MCn68xTremAes664XwYUZmWVqx3wtutGqGz9CxA
VNDtqszsuzq8DZJ4Jynw6xjZYOwLhXpvI7O1HrS+31QmenglFbBHjUVUga38Cf+p
JFmty6X/Uo1AIhulxrdQcQZMmB6jlGfan+H5rBXyixFoGiMawFoPPBWeLSSew9VM
coE5glYwumXL9dllpGSeEz366f6PgShxh23IUfZkZJqcaV3xOUkNqRmpcyabXZA/
TF3h1RQoDbcrlck4lKZEJP0B/TWxl9uwP73ks4sLL9AC+3s7APjXYX2cfY1yLbGE
stOcpsLsJBx4k3cuw86sVXaPyT2PF8dNPbn5sUy7Gx5FsoJtEkZNNVNbaF6gCpdi
B39byMJc+HQgoQZ/MGs3Ib0WGdq4jpNDTnZK5iNhoLrUpg54D02yNN926jY4kG25
R7yr8dW5JAt+/Tu9JDrpbIJ+Va20LkIRhdLsZiQ2I5RPp36RAFuuQcLquvVAupTH
WxQKpIsZF6nyd81tx8mguSLtknhSl3hiPoefYRgC17su9UfuWvg8NszXvySMQT+6
1NbjPmLrmLtkurmuUA0khtrp2rVE9pykt8iibqmeoDnHhnpDXOTLaMb3TqY+MCzr
wEKw8kW1Lh9NZ5YIlRrz2Ba5yxqOTt+Uevu9V9ja+tCow2k4Mpc24W4k+gE8APGo
5KYRiggEV6/+ghXJcrTMJykk08fUso6muOwsbBnqBWEGVCdjpepSUbShyl9Ku/q8
uTyTCLMkZxlvXi9jyC3knsA/F6FpWJUTjo7VNKExE9jpZE2Njg8bR57axVW8/yIa
W+7KFLQeHnQD9MAoRQIpz/g+05ns1ILnlAI5RVuSvug//C0189suafBa2V2ragA9
F68Dedae/zBwhEytLwKhvTv2WMqW20+Uk9EOO720fo0NXwpX00bEbVJ2Fg3tZvWg
pwJdD/GnDyvPYkB0k/RX9KEu+c5V7//SphWSSTJjuzJmMEjU4X0QZcwZEK+jI6Vu
BOseKyy1CRypOiyrWEG3PgZXhifdheDprNuKkS151M7t7xxZLwnqAZ4oe8ZZ0Tdk
Wpcn0aPNA2GsmJ8nZZ0MTCckIAaiWE7mFVar8BqcJzNG5ssdB7pvx3IhEuC2i/Z7
fNjQ7ykVnxtNDAfyLl+bmdFK1hDAjoKKC5ClVSSLp5j4tXEWkTooG2uQoDBvEa/I
6cS+WY8Z9KdQP5WPCUM3ZgTlM11aLotiVzp2VnarDOjoRI67wFEQBOZq0TcOtjBv
WUcShWRaWfXVKHI+Wqkp+9ENYePH9VsYGmm04DKqBX9+hoR93gn2hM/HnU3ull8h
ITL49lEH9Qc82boHVMvAJKmoFBdb2pDu0bW6rmZeZ99k0225gwEDjLiyYDr+GxJt
MXFWWjP9FZV1H6WvSGkt//ao5xzgnpZ0gQFCAj1SH6PAQYAvY7oijByGUU8iNHQM
wzNi4Mtos9TkmU7oObgDcgBBEUbphCn1uubbriULKdAO2TjkgvBji4zzUPqReaH6
zOp0ngFDSNII9Xg/nl7QDuX/55DLQ2FDwQMU6CAZaSAUyigQX9qNmQfTqrvVAesm
riDs6QzLxsLdDBcTqLsd5Ok/VDLb2Zf4A4unGdB51jEXvcD4YB49EH1nSNobXcxi
Veuc54EitB14Yq4PtlbFnDkpQI7JlPtoJzXTAB3nGdL1BaIEmD225lL89UA/O9ij
MM4M1kVXJ3HSivZZYFd7IXE5X8e8HdaJ+AGNE5frFP2T5TpwbrY2ytQgFtnWEYgy
5FhNEdDZFxrleOqAy2Pn01kjXHYnCQZ2YXPHgvhyqp92JSWgzOSHZROGkYioaMdU
vf55H7tqqcU/NzvtNhKlwwQ3FHrBd4wJLEBzWpiTzedHEXo3kMF4EJSrnGcd9NDU
yRq9z4NZDWRYp0ec3zSWI2VY8aN4GM54beNLRIAWjWa6PfpPydmZbCWvXoLTPzny
ZxU5MYod1MA2Iv4nC/CorXiSHTXf/4PTscmFLsVbEMs7vSD7kHpkvUZ0sSiVEaEU
Q4PhN94d2u6UgARCT5rqr+LTDNGaa63S8tBd1STv2yC+njQSuwBnfbS1DeoferS/
bfjLeW3PQa4Ekq9cOOamDE/aJ7cOHp/+6P/G03htYxkKsjSKSTigdO8CHF5gfQSb
4bHvVj1t0t2ZTt0y8jaregDYflfHgUpI/R1oTaE90eCgq/6WKKreDYE+rbxGS8yn
BxAa526/KDmc0DaRooaVNLYbPJsHrg0M3i5V339RSUE366Ar+FgePcEKetF39v+H
ldIyHkxQOGY7e5ZpNOkLUBZ6mldj6Mn2LhIwEdNs0k59Kv4Cg78fyXhZGYJU8DEA
EMuMzd5/JtBCWZ4paR5GTXxkoOUg81QIIqLeLeMqfBOddHnrbESfBFfwlwA6F64/
ccgFqxBqnZpZmQbh7BNJMNAbtaJjvmxz01q1gCvWXHACGg0Ebp1kdRklAmja8cuE
R/wg9Xl1h6llTMQSvLwKk6XWTlp/PAMmU6El9aScst2tHg5X0lHHKnDVJxuk1nPd
S9ihClIEbGKtpgBy6Hai2J4cfg27HkdUAA2aJjeraHwl13EZ2t7vFTWx86v2Anxx
QMqomcWpxtiXhzFkwrBR+dJMlRRxQIN8vueaL6jh1OSXlWlGfTctCZXCH7YAlYZv
7GwzXZq1ncXbpKQLQpaJRwPFWJgSD5Hvr98Yw5HODj2yIFi3PY3J3N3oiW6/g5ga
1yabZ/3mVwk0o3FgLjmLuxJYAmnr8o998ZbbnFRXDvhkLGKRrxxv9hnNAGe5A8Rj
40dNb+BklKMSiQ+M5UFodQfmzMmq41EM4PADXjmAX62U8IddvmwbkR892qNn0CEO
JlJ4dgNGuobiskNQ/rRoFBl2HnfJW2xw/RMmwISoX3hRcu/QS76Odz8TEpf9t1Zu
KnpgruHPeLWn8BJ8Jq27B0aBXryOa45gSRGqwlBhLflBr65LkwMhUlPCWsKc3pP2
c0nMS0RC8YPZbiq2sy1xXAflnsqRYFj37nNIfyBNRNhlrz0UGukPy4uIhU9aN48m
3yXyXsDG7Y1a/b4f+5sEqLM0O78ZLbRPnVY1iqQfWij2vBgipxVYieHc67kd7rZF
e3TEsbHcw4eNFcOr4VzN0m4IHH1R/GscFfPQgyN8JCf7NCoQ46EYcYhlpKbnGiib
FluoU+ogPuo+cmECpd+rFdlk+/fBdi394lOtDBZ5RlJfpzq2oZ1esCC3qooscqE1
CD5fw9TDQ5wVnMuzLkxAF/1s4EKMqwd/6cBZK//Hj09kI39aY1G9kU9ZWkE2Nb+i
g1O+mVRWEfpu3WXygbMACiLsGwBL1xplD4ZbcKQorX9l28Tmk/EKWwo83hXe/Oiy
5teVQOgWg3nQWx8iPS1G1a20ZKWAPhNcKR1uw4Ar9PkCHTAcD+WOj9AA1VdMh1oT
SZxzC6qYuF0dt+Scc2JQ/MuaqEmVT37U4HmTuerbEYDe2hVk0v4YNXtZVqZ+uUmE
fZONU+E348jSzwYXYxApcaTKCp84tcAtFCN84c9e0cLLc3TVd+qQfAO0WlXHxXjM
RS5vN78Je26yowysSd2Y580kVJrmNFfCuDY/J1ajrn7MLtR8tLKhZ+DT/ISsjVg/
7v8fg7L8sWKEgtNs0fgpKBZp0w9xjJdCGB4TLPada81DZ4Ao2WsugEWhJa8rJRUk
o5lV5Sgj61SwbXEUJ6qj1hlddObz/2TN3nfQopKBF3qrlh64y0hiEeUZmaB9vWFW
BeXFqXUZXj3im5dqFFIQQzUFNJ/jKsWCfPlxOrok2ausRZoTA0LDoGfAU/nC2qd5
vdr+uqIJEL5hQcJ/IPXLZzQCOEO95YiVuHmKGPj11g11MlV2wOL8idnSQtdb6ABf
zzR3GDwnchZOGD70JHmqKP7pe/X9NYmVL6P1QcSUZeRiwWqaCrF4Tu0JKdVgc3R1
wu8puyStuz5tGhKA1b9xBZqbpeotZJ0CJCCkm8qVMm1eaww188dl3ciq1j39e4xj
xMOD5rAHIccPPwAoB3+NUFwmOcvQdv8R4j+6gZ4ZpvF+NvfNjmXMaNcUbSJNKFca
1eLKx+lVX9/tSe5Xx5N0dKRRO6wLMa8i9WHzZzX0BfAjLkrW1AzOSQOtmzebc1aa
g4nR7oK0chTQlg/Ws8boJHrrT7c1Q4zd5IxMGhM6/+Unb42RQnUcxPntS3xYoyFO
z4axhJLXwZSmwORziKkU2cuTwLz/o1SB28nrkPebw/MU+VhFj9JTYLEeGKb4lcDE
mkKoCv9iYsSdBICoh8C6BZ4uJLbD86knXN785d2TbE0xpYaLCdboQMB3aFr2nLSr
wN1UIhwe4eSAnHjCsuzIsbLhmGK9T5IQEzusFjlXCJvGLFSAHC0NR4dKuperV1KQ
Ejvr2DjCWTlpeJJWJEhLBY4p+qHsC8+J3fxe2HXVDmNXhrPGV7ef9FwtBJ9zGILb
LsRGmOD+dtpNP4brUsgqlBlkZ3LlAFLIjMRy7HztonqukuFSHu9pdhtP+XHBP5rq
g4UqhbNoFzhszVtawlxiXhSDQzLJG+XN7xwTVWUWf78fu9wf6DMQCFl6ja9OQTN7
e5R5jHh4VBUZokJYwtAxBYOTh1P4K2CnPYZ2G8RV/d0CEyTOxWpng2bafI9j/NOs
eekKLZUsJEAa4dAjhUP01yTLqQ2nA9ZMMOxi41WrLgrk6Lm+KjMtMkZhRbBHByjP
hIUpQqKdwJD98BGhDLUs5wKgglS1XPVOa1ZvYcEwDzYlJJ3dzihe/hBSojhI5YcO
zcI0jiTxQX6rGc02qkTSJrI5ocP8NiHW8QPlAxjTPC+YfuZk6RBu8rPuWdUUWdnq
pFit5O6ApzhNpkIk09qpfYzcI3JWpvQUTalsyrvGGJLoqFHWyo7RZXjU9pQAHjBi
ZJcCCTbZHvCsk44egb3YIRmFIO+pINHo9ASDFhIRulsvfka84anKE7vtSawP1vpq
aqEHCIWgey5VJTDAPKaZhaqCJZ7BrMRfOFkswdn2tCzlOlGVQoVjfuIwkiL2pHNB
8BwGCLirG6LgqLq8k2YZ0YAO4H5Mpnej17+laxQnfvD+CUwRbl/jOuaq8tu7X0nP
67RVu5iU2c9CADE4oDvj7askcrt/DJs/EyCmCfRlcm1eelLT7z8TVOFKiyOIG0yT
AbS1oZhPn3iHXnVQWyHnoBLLobjgyoGkoq5yJq5zYvS+/Ygbbj9O+k+J4Q16wurX
3UMxdwDL8OidT3dldEB7llTGGlQ6bSEZee2/sPsVr/IQvGQ1dmZB4vQ5h2Ij3Ce9
isVbASkxAcOKnPCBAORW3xScNBoCIZzadXi6AtUxJUPyn7nBwVLXaVaXGOqPDxvy
m+mXgC7dNW4ZaPu7e868ceynwm4abU+sc/yQSFoMCeundo12NbjDGhCzW7aLqvzR
0D2SkLLP+DnFqv2uDGOsN2ARhB6sIHDLMZz38B9edPU0eF/oq0yLcbWhyeij2Zpi
SEZwWdLVxhNpHHeJ4VLVSDPMbAsTTpqDgVfiTbRqlR1AIHHuFBVhiDas2IGk4Ll/
jUHEupyzZmtZMpdz63X0eRe3rzsp+y5DBCqE888Ivzcv7EOjnKe3abAwJcjCBihy
uazNn4+hjQK71bIihX7KYrLsbEbJXcHzd1gexw1O87fuimWrO6uRopnZ805ueF6q
NxeJdOnByIwgIlsAMRXuy0adJ1k2tOM5H6x6Kxy5LAIlE0Y+RpI8YQjrBNb2eN+w
MCpPxm9kRHBlVwRqLOv9x1n3lRENESSD99/tmHD3a3UnOOkL/jy8iigRpLHfgYpY
CE9dj4e+F92SsQX2KiX+NG23Lf8gnVUCJTVLT4R8bAihFTV1O2PhOWjU7mJh9aoh
kaAgnPn1+avFD783sCrGre9C5+bvJug7w3ZbmDNM8HHbxgpNEvSb3nuYND1q2ClO
Zd9Nc51P7SPCAi3E4cv6XLSzVchnPlcnGv/vZdqq5Ugxblpp50phCY/CjuXF8TCO
3r+Y3QqBOOVLmBTK1Uyzxxwqn8/p87HVs9AwKSx4a7x7+kTXPl+G7+Z4rTJSU9VQ
2LNBtMYcSsqadOeiiK5bh5ye9rjg07mRLZBaAEDdvitKTsX0fFhKobXAdLjfeaz4
2k+kuPsUddN7HJQkEl7pqzW4hpuFB2kXeZYNAXqhiInKj4hUPiMXMYvp06qp4ojd
EsMKeU4BnkQc0hzhzAffP3p6g9afnKO2q/m8o87sfiCs59T/38w1H7W5OdRW3Ip8
EkD2GR3VjIvPzoNWcXA/JYcrAjrxYF0KJw3dLPtel0YAixM7YaIIXrCvfZnsUIah
sk6QKrm8eUqY9VCpQgOGgwGNfoMJo+Fk02lJkK2O3pw69wk39qtVP6BPtIpBQFGd
IsO1WVCzIgjJNpnZLkzPWarZBO2+7zVMjHtm6WVLzeuf/PKANIf1s9CHgGigR5Ei
S2dlAUxX7vwdCwEIj5hvpKhk3wbz3dGMmuW9OGQWzTrUPWKvgx0P6bMw5gLur/ir
0WeC0R7SrM1LmwoxXHsI54VbMkPQ26AEC5zJLvajouWTzuY8jugn699Ah6zUiqVK
9joLsp0HbDEcvgnUrWt2qeS5eMRZfdYcv96QKRCKTh5JfBqKV723S6rf9yHxoW0H
W9VNBBrKBJfr4+y6kuPu7L5d0/T3SFObmP3uRN7eCWuOiA5M9PYvrrvILc7QmPEf
uzlg5OpaqmWeDueOkANRTt7rE71PlM6PEalM2PTSjfJ9jZAe6LYq5tdLVjkuSYSn
hoyOZF2k+tOHD6Cd4PLhW2oLHny2UKMT2zsJbmc+X56LaxiK5TWxcUdOXHa/udB7
c+zOUD3b/3kKCc72mutz5m70KWPmlJkVf8y3CWVbdpH2xHMzD0FgBMDHD7pX1Qm3
TeDKEA7shRFTttlCJjbrBcxMNNPW6IRMfP2jt/gt6dpK+Gf18vlWq/ME5366j/6I
aUVcxiIyjlsVrD6xBVezDsekKjdVNVWI1mZ0kQjsBfZImi1Dd+jRU8dkiMdHsFXb
4b0CFfnugmviKln3vJ9jhAFVGSVW7iFG3fRjhgJPblt4Bb9jHvvHULmopYKdFVmZ
2RDAUrZN0Yrpo0uCpls1qTgS04BnOxA/C/QwevIQS5kDfOkEKND8mideitdGmyt0
9UUdmS6seeURudZ62YE0S6Xp4U7A9j/RmkbJzJY2zHAISl4frV8CFgTc5g3QTMal
naqW0ZmoXFPUSaU1HiWjGJwuhZU1qK4y6MiJej8hsaiE+1t8G6JoAOCg6xXdeYi6
XybGDoX9hEb5Cphgw8fRiQCwCglLYf51WrAl2OE1XtCRn7F0O8iq4/A0wXprQWkk
KHQHKorSN3xumEvbQ32Mv5OFgKBaW/wr8/fQ+sZhg1QW77PHjgwUYp//v1V0md97
YVISBXJWuM9jzOUsJyj9zKhzZ2pdCXVNiNksCe8Ve+/0KGRGcnWDIrWIQHrply3u
smLnkeSQLcQcF6eWt1XBqB0oe5YAg5E72AbExQ+HaTkSxQ6hEjXBXpTDMlwihewd
62GzgHDDbRaXFx/eBTS8hLMSoXkHDtUMO2x5LN/gZB17bAMQboKYMB6Q8iYdq9sa
RXwc0cWa0f4mP1O9VaX0fTmXhTxbvY2t2BhrIprgy7B6qgpjoLvlrhlWffxiUFxJ
u+WHdBVuJM65rCO0rkQZh35NcC7iL4ndANKee/eP9fuKzTuYTzzW8Sxus8v/wzOk
Pgm093qGdeVUYeNOlEoXJLvtN5wa/DPk1u7v87dd3do913fgjFuF+Fn0oym0UyUf
Y85p9dgZ0NuAd8vRmgYDiT9CxPiXMXCP1/59Av13nQbTQuazLPFMx+5FeI6y258X
ldYNe9g8sBT6NDSap3NLZ0Aq9rESaaRlUkJ6KkWsllF0GoyH0WgDgtfADdJM6UUV
GpkAo/GZn94fuuOZoUJ9DoR8Zp5TOQToy1Jxn622MXkFgJ6k2onNcKqrBQsvFiP9
etcL3e8u4zIJNJQ02va58GnxdOBGwt3iVm+TN2gbiAG/tCEzcNbJ8skjDrJkisdp
6McvaX8OxxWNYv626Ksc/argtWJEG2BHSBdDdceZkJTzfxXIHgcVXXV+AJm/H9RK
44edvLIlXm1gzMEu1bEmRpM8gZ0d3adfzg+abH4sPtmCXixix9nfLrT0Bh4riF84
iqEoOiSQMds2FAKVRt704mlqrWXojvu6MAbp0ezk117EuSe7QLJeJ8j5TLffbOnb
YB2IFCzoysiCr3mLeaKY0Oji3JpaXpki/Lozs5ve5Qefj5z3M02/BfMaaJyVUB/u
nOIe927NVjCOSSYvEP4wyrcEDRzD9aUZrpIaCEYpEJPdzK4YVFj6u6amCHP9M5az
2UQti9XlyYhT/jQPSq5Z8jlD6kS2RBL2itX+WS9yNameDrlZHJn6XgeD8QMiCqx6
7MXmYIl08W4d0+0ADYmB1l+rvIK1yz0Klxyj6qfZCriZjIFr50Gxx2/JZ+oGh2Kb
+ghHnZWGaLMXkhXdbZEXR95QFYNr+k173dYNFkEP+Xew1wD1MxvTtYF5aeAHQcYG
cHIWyipJEuhm2YPaA6IqYxwYJMx+n+qFzmh/CGlu7oEEacraRjg/+fLLJC7A7Hj9
ahOq/Si8T2hBSizgkyPlcGWgyjuAQd5cZLzx9WdABdxbjadcsc+4oldCrMjaRxv0
EdE4lB8E+WBjXKYH7PTceH0L5hnQ4G1o2I54IUz7W8BxxbZsix86ZL1eD6ayzt7q
SJcO35TP/gVgs+BbVHSxnHOMXNTYN1CBKFW1WwaEOUqmk3Nbd9ABbjI0B+99i2lU
W0CsX29wN3pPJYj6uCm/weLsl6k/hTLPz+iYTLinojK48bATngD7D+Y4Lw7Zox0Z
Ktl3ZEHXht9xyIar788IAF0tvvQnbjD0MB6a08GKIHp6FFo8pZHeBp9l8FwMHrex
m9Da15yB2NKS/6xL2/XDdRorc9yCIFiKRQT7asO8g6RpDap3p+XfwBgLj1VK9UG6
mNWMx4fW7x5aIBJYyWh1lQq0Yqq7QYuY3+uLE4nKErxFoNDFdtpOL3vfCI8tlzp9
GATVdMoplcxW4QUPCtShc322bs5WMCxCQ1vWX2HrIANPr7efIRxVYMZmLNP6S1IV
Ft+RTUySQjkXd8AfVUByns12WlHqEVqIi6b5E6Auwo9pa7Li3VZFyb65QhQ9eGkk
ixkLfSM7HtYirQzWGrMczBdOMb0CP7yx5Uz+4+n4frUXO6GIvBrFndQs0T8xJbqZ
+eNDiVTFOouWHVdH5KaEuLC5h7kGCsJEkYpuLKo4bjP267xJgvzBmlcaJSsx0yHJ
3Qf9R9AYOvHZ4DvZgswzrDcslbVwYEwGz9rbeM70s1TPjMwWU6LOP+jXH0EKJu5x
nLu9fWG58XOwqU2yj/mMX47pJMYpYehop72qBCDYBSznDQTchmvZ18uFvanANT2+
oiolyubhXPMPUAB9dXa8NLaF15PFwt7TgQ0chsXfUTzsjna2jxUCIW7WE2qCM2lq
31nfXz7AcZ8qzJmYIthenz/9KHI2EJJpp0gNDbuVU0T+PqRoxEfsBRVA7XhadvRL
yTlZSWBniRLcDuz78IUh78RX3Wvvye7qGCYkkuUVEcvGnwdDvaj6JLAPuPqNQ3P7
E57pBMO8zZoElgTnvwf7x9MMziCAlxOKWJtS2XLw64x0O5bCCmz1ND7wr4OxPXHP
EjbUrfdWBh/Lqet2f6JRy7M+RdCHjqIqLA3pF5JysR4o714LsfEnFT9dFjVoSiQh
6Qt9qcS6yYMX14Z4wkUREPPJATXAAx12OurlfckjCngdEQKMnpNNwG9SKoL4iLRh
`protect END_PROTECTED
