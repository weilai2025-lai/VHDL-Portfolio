`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k4yA1O43WfNqoCogvbvLDQ5iekPzjvXncLSwuEzbYIve/3TfyUAShfJ56AqvVIHd
VG0vwMhIwERtt42k65xsWtz0Twxaj7zKKcf7bD62kAHGkuBWfh91VjmKecp8kjf+
Qmmme57dTp32JJjAEMYlV6SVTW6lIP9TfinjIIt3HLJCHbHHE7KSxlKAaP/l9AA9
0WVys/kBNCGaUOIB2KaYXpOKDdb/9DEd/qygQpXAIyie3JqiL12elMfMOBsB0yF6
2uw+i2inf/zBpR8RWlmzz7aFomgho+h4uSRH3spLaqv6PBEEz7Ygoxcnwp8pv13j
txtzxtwhmldHCyVu8Rub9kL0bVsKAcsoEYAL4CSEGn1pBqmvvjZddVV4cW647MWn
OqIK4UpQSeJo2W7D+SDMwUiYbo0cUtvMCgNBEjjeO4oIaZmYR+0VU4lCo4PH5EIv
FyzxYIoZpZ/qNKQiDgsL7SlPJpgkqZF21MGeSt6h3hFaTrar8xBx7oHmCM1lFFrn
9gFcFj8/Y4jeUY5gvkxV/5SbY0Z5+tHVFYElllkol8r7rlRr3BkXzjcfAv1hxHBb
ssc3Ikaa+MJSg+mk+FBFk4/9VERPkNbynnaNOTVEoqXljKZG77kK20e/AAa5hUWE
nekgohcLRoZ4+CGnuEHswCLlME7fXZrFEQRUVk5K9/Lu2HvFmeDoQPEiwjOZjzMW
gtrfmqB0t4Om4U0L3DbgshliLR/tkREK8vMaTQCIsDCYToCLPPYX8+vv+/QPu/pU
TNgEKwwzx9fZqGgNa7euMoAyqi4L5Bhfa0L3kLPOTbQ4pM/WdEcSOHTOCUrPNYHy
PumXrxlLpdTW9ouTAlhw7b255T5UmkiQ1lRrhnHst8J2USho9Ur1rrqidvCJvx+h
iLYlgQO5EiZtgwiZ2XNWXdv3JQGLWnz9ZNjIQqpQdaxNsm4in3tEGfvR83SNtlQp
OmAu40LGugqyRXYZ2ZY07du3t4Oc9XKzueZcBPMHzEVlyh7SCM26kVleAcP8Wc+Z
DZBE4rzqMkocBV77Z3S9bmrWO0XRI7Y/bucjtSoq6h+Z/J4oD4LbZJH6+QKes3jX
ceP0hOswfeP44+QsRmBZPKTRQIGDxKPJBz0UIjmTsoV8R41sMtbQIhDoR35o/7Pu
phTLGVhqElLFbMe3SQuzraEemTpefapIx661/c1C5AYPJdhn8Kwgjc0hA+H/L3ZE
HBcgupXaULRzPoWFkCLjOgcl1CDwq8I8bdJzlfOtkg3muYD38NKnb+sQ9R74uE8d
48p8bEu8/F3wRIuiB8zf4Iv3ee5pcUAXxm4e/lsb8Thzym/I1PdGBFs3C7ALZ/RU
2593Gl3wXt3Up2+TalGKAUJ8lf8HDHbLre8jn9U69uQAjyKLnLtoWszSQt59RENO
ruPXeJXlS8Ad+lijL1S2Q5TxQghiRk9c+3gmHiRCEYfFPw3NV7PmMfsvdPGGNp0J
C0MP80tEiYSWjHXeDuZTS6ul2gOTx/E5U1LTesxaE9sb32IkGIjgf6FL61g+1+Fu
vhO5enqBTW5Q5HajUQY5I2xJU8yhkrfabVBGwc7c6KUU5nvNg5HMoNeNrJIZB4aZ
0juq3a43EuxL1Bg1748kjROPJYnOym5L6NFVEtVHP94dkxKxbtx7RBuMF1JKZZXX
REEatTt1sAXDQoS7202MEr7lkhHRIxISxE2WV9iuqxv3eBj+jb05zSlrpeIX70jT
G6poSkfa2JCGNY3KezjGVLMBZKEYljrUHkseSHenc3PC78qr29gUHy5yuNf5jZ0T
BEtw/hvggT1qva0uA4LSHxPx1erZtJa355vV/4ulorJRP9reyoZ48SyaWzkbLpqZ
/sLqW3ri+kGwzg7vrJ7yGT8vBfnX0knWlAhrnRQw4Fkekc5OOHxCkz71sk+yt6k9
mScpq6TCX8qqCpAhWZVz3arCBCr5pEygJOJIuyBbPyt3noPjoDQ+A/NP9//zQVaU
TqhyRHBE934Z6dOew7apqItAc5ZX84wnbWknTf7ZoZtrKiRgP0xkCVIz54NkkdOU
B5Jwj9gE8WAMMCdtv8g4lFBtDzpXESOw6+rDRdcndUYuSdg3b4W1rmFtIQeFqo+r
6jlmMvUkglw9EayOjYlozkmiXpYYvf+f95ZfVFrDs7jPoYJfII1M/h1bF1jXuC9F
fqYDALBgmX9dMsxc5leyNxlDCvrwboY2EDKVCWMKu23xYs6Saz0FyN06ZvBZw1ay
m6bLOXE0BojOHtEAdDjTgsP06GXPCAvJ10aqVZhprWtjwBKlyVgB9AETfypD0xBL
NFXBi8PuKXl7QI/X/G+6PQH3C83uQWCJz0b3jqMDyHFEHWg5DIiUDGI8mO9mu3CA
OHOuI4D0vfLVZlkWKj+feMVdi159e2MFodUstz3Sac1/QaTl9D7ynjZfKL9ce1nf
AliqPDhaLkIFZyHUKc8iUJKUERexunJR/vWx4dBOrgpuO12GlYe4qg8ijbs55SXf
jvFP9WIry6CAethxWMXNjqNeeVViJaCLj5fLFXrhw5fT7a5uIiQI6C2/Lz8EdNGI
0MNW7YUTdjTRq8+jjoGS7BtlNdW7S0H3JO24AaO+DcKWKd/tTLy5XJyHHMi2j2st
9xDF/CE5dv5lR71uFH7oFtlDgIyZjfs83p92DWvq02Si+6BAGa0o47l5jzNxS1A8
dRjZDWLtPLfD06H/f3abzUmFIBJKGt9pNsztUR2NMssY7etvqZtdtTtoOZe2nvMr
8dwM5JYs5xEa/waombk63FbRO8sqRMJqiOnwRfYbU2mg4HbPXGWnu4pgjk+O+zX/
NUoXXlK2HsP9vJd7IGFwcgE5vsbEpr+SGw6eV8Uxo8Q5/82kiLJv/TN2+EktbXlD
PIVxYHzkLcBa8fJy6vAiXigx3Lr6KydoVSyio7LF1BD3ynJPH7IDoGAh2Pxrx7Zi
hyJ8gtGlmK39L8x21Mz/WUzhszAVLz6Lb8WccjBWTApp2j/jv5Tj2nRtsKK6FsBY
pNH4dp6xdExQ8ep1yA8uOGuZVbzdBMzMF6kym1rICft7arKVRnuAD1SusUbBHWiz
YrQt9sa0foD5NkmMN+ZzR9S6nu5vD2fjhryuiSZ1UxaFH97EQIS6CjEOsGcdc4id
LLP6K2l20PWma1QlpuSvjgXa8dEUJGC2w/UMUd+e0sU5sWsiRbkbE88mFFCdSj8S
XIlQ2rfRnA0pRsdPZjoLHIaxEj3BLcddEwiTxgg1ktQn7ZPLImgMYrqFtl2BwkEj
TTQL45KOUTJOccYX1kWUDnmJ7wI91Zp8KkfgfMR9TbrNVP8sSkU1d/HzHDTdbirp
mC5DTpg0xuddoKwE7WKK8J4drZ4o+a/Hb/hsrBpJ39Tn/kBptxqjph9slTZynSxn
SJx91IBnQ54N8SkqhoN/fv1dbJkCehwTNn81Fn88MOCLDoqZPrgAlkUTEAezOLW8
Q7ke5VS7P/J/yup2H58xFQyKlSVXYV7biJLHgPayDB/dCZVXUEtXDNstr7xgBGjG
4u/dcCmhL8zwWQjkV9VM0Sx40i2lw7t+zsgGj1K+AM1GGds9sQDdXJxf/QUSpnBj
C0lSgSU9WgG0llda66o0H1ofNa6zBCwNrgaVd4106hZmhEHfaIy6KZV+UTa3eFOK
eDAUngjV0zqV0GQaW/sy3K1IdkyKzt1rPK7ly/Cbo7YckqOYhudW0uraMbRD+yyE
b4jZMHI1EpYOK5xjyMl6mkxVnYFBoOjE3peEshoDmaS9EuVX1LvnwuZg/8UMlJRB
LRb+Z+nSB+ms1BFY/ge8HOo3TCSabvUb6tuEcwg3Przoso7pUJ7IjwNxUM5zrRHB
890lnVadeJJCDl4jQrLjaL0tNhjVuNGhHWNLdhlwusfoAgp7oN0rq4es12DlAh6T
0b7L3AKXFarzUvY/VEVLbMtqsDDzOWsIwoS3BODSJ4leVaLSm2hF256adPufkwgs
ghpIUa8UIits90w2QAEXDyyxWn6atGS9JC4Rk5kJf9Z/kTqGg5nRtvxIv6pe+co9
cTastdPPTsq5NXp36vU0IyppEPlbkv9P8Dy5y/A1rrzNoXYv2gKlgWXyU2Rh+2lj
YGqHUqJKAYDGPfshB72NZRLPeL4m2D2Ad/HiOBGr/Lp3JcLoibul5YmHaHaZ0Ii/
QKq7ZWLuuSMuU8VkyNsANVAGSyMjPrIoP8BtYv+JNC1/j/6dtcGTlmusvzevtz/h
eNHBehk3a35N9AUfvL6q2sAsl8l7ebmJSD+1ojQcPb1CGNSwTDI0TPqcQdhjlgDg
pJH8j7K9odAwn08gyylIvf9+elsX2QfPdaN9Cjm1DDiOBC46i9HD3t+njwpK+bR1
EL/tCjzTu4vmNL1eYzLVFupH+k+Lk9x3o7SOiZ6Z0FH2gQu2H7mIrX2z0ZE86UpH
bl/5KTWbQGWX2oOnPftPlXFQFDlMk4PG8t0whojVfGspPYfPVRoMgGvMIqlWcZDa
+HVdfK0BsrQVgDGaDiconJnKwh6RSlPOPRaHvd6QtcdWVUbLGf89MklbGLUUopOA
/xRWeV33oedYTmANFQyIQ2Ld/AaV5JhX2CwXVJwcbyzK4jpinAozHwRfrF3eV0O6
QZONuSh3MkQIZZmejTrk1x14mrVSlXVt0QlIjry+cyu+5rUBdZYD3Enlr4t7fpIt
VLOCYgmv/HffOur4lmZl9PDAnEwNXr6S2L9n7fIdI/Rkgv3FRvbXZwhevICs59Rq
1KSqoDnf0Z1s2WHHfUKVP6fWOOah2SwuzLl1DzHq1UgydUe7/YOHPPtj0Vnh2TH6
rpG5LLkfhFm+lCXwfoF1GFlqGDA5F9fPeqrebiYzpy3DU+3VUXusHCZgOLdgq6Ch
2/NXwGH1iYjvSbx4geWW7lb97Hit7oFP+KsmeaIw1ASytjLuhQb6NnyG5CEEY4n3
/zP1zgIX8XLNT8GrTqKXolMWwlvSuCMveJ6LB44LXcnlXsQIG1IC9fli9GQ9zccx
4s7Ok1YH3kJ7yd96B5VRRqACd8Xs4EzJxTkRpbcRp02P4+t+9yMiDY1Eqqpbrmv2
E2ljxV26L322gdYSWF6ZUbogOTzr2OXLWpawde0cdcvAEH74m7YE0YODuv7WR984
a+hs58R6O+3FJaL0hd2vo7Ayxd2w4rr84FYLoc6vXgn/v98WrGSl5h7x0leX2KvR
dspXAqqpQ+XvskgCQZENzeLheDWBOszvgJutSbXoa25bfnnFi/ZZ2VgD6Fuec9Hv
Q6dUbS0E3ESuTytx98V0xWPnFNXXr9ofgVTKKQ4hUmmPnhGe5LVRQ4P+LpG1bVR+
RAuFCZhDMcSBPR9mlkTtIQBreeYygiaiJ6cwsndIpSh6cjG0v3KMsQbzFzdtV6x2
N4dDI/7Xp0FVdtvT5s6Rx4/Addyt6nGj4d8UHe2lpUAy6a6DL0zkpvmBtSox/rHV
EwgltEaGFC8Sfgv8+3FSBn2RSpsmZdR3LLQsFXYvFkOnepfScimAUMaYwPVjKWmH
fM5HmxXwNLp+1hnY5Z6oEFYx0ev32uO/sSi9+I5+67IjZKvbWmXaj03DtXNVQ+E2
+yp8RrEwcRLgeR6ukh/rqEMGotwgZ2U+SIIxjUS1MnrSkibOMvQznxAbXT/27p7v
oBPl9jojgLlOBDpeuNSoMjPXoEbXiUFiFA6d51BtfJ2jPF4ah3GA2/vXtFatSB9h
jDBNG+/q5i9Hbl2cC8gUjQmabo/lM9x6qEaVrqDbtKnYFHiVmNNw2VlX2Z9297Q4
chHB3OlTVwXsrMoJvbKuF0b7XdzA2lu/CDf5lxjRtIMOG+nHSaBstLz3FPYLEHsw
0bHujvwZLK9RcBZWJ9AY+99ANDQFd0C1vr69sOYjsYI3BN5rRAhOsNtOgmAK+mdY
WpBzKnWogmOueKxl6OvPpu9uenG9VR9aeTZ1J5bCFI/dfy8ttJvXIednyPK5NgBK
JLjRNaNlbBUDSMyNQYAqhISXsOdpY1mpmnfGx+Q/AUaLSHRsWS/DBvejS3ggQcx1
CZJPEiMyuAK9idO0GasddNIv7DDLQYByhvJlH81RbU5NbxGnJew1WLDDhNmoJDc6
JXc4dUKsYvUuNdjBnhcqRKQlbLLmZMogvHmEgBYpwXi/hHeWZYrgG0IZjiKiotFe
a7Y6T/Ks28fs2so9QtG8kckCVS2DLJTdfYcoTXPyDW0hpPWXZPYbqypLUFPxnV/O
/JijZ9ISuLqL2HNa6qAV8XyyzPI1xHmXk3TFitd/uKbkj1AJalgXGdcisl0KKlix
1HS14M0SLzuyVHYk1vZBVnw9/EX6gscfEpj+43YaFrHYg8jKZ18gPiQ7yTbnlFnN
s7oqz44QlCII9fal5g1rrM+na0HMsabt44CgahwrdOGiabQkwqpRsVHarCwAQocI
veoH6pjlSdlEK6SDVcp1FNxxkOZBZmThhupv2G0o+MBAlgovSXUx27BYRyKxliw1
oqg42Qm1/vpP/O11O7ICJxeWkO5SvzvUQ5GXCeyvQzTFilB6AlwLDzfaXS6DkmDe
iLw+ZyGjAJQC1H6CebFBb84du/jqHBUJ9zzJTPEPxC0WzgcYkDAuSWZkYbp6gKYJ
b/9cYpaHzAq7lrqWcHpoJvjKmd+cWPExYZdE026PX/DTiDd6ULNzw7LnR89b1DJJ
BC4WaNThzHtxCTmGvXHK+IbClnWRTcsDPquiyZis2K1ju2DpjnI2I3k0UVXYyonp
8+NfX/R6CAE+B5xMy5wD2Q==
`protect END_PROTECTED
