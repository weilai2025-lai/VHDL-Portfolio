`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAEd4XarqiUEQwNdqROq2qaXka4X1Y0vW3wAzyWwsrnpmQsvL0X0zOJ36+MY2CgU
+oYpxM7U4L76M/NlhOS19nVHL1VohcDQcjI0eQT+MsZTAy4WJ37W2Sb+1ftrznYA
7d+NH1a3wShavtPN72vWY7PUopmjUnu34xZHALeKgXqm6LrgadZzI3F8xIzc/Q2h
85ZNDJsCbvV1L/UMGwnt1w3/xMs8MdeaJl5DcCsC7pect+LXZerWFdek0sbT0PMU
xzA1ltW9KKX2+gmy0NcWcrX57XbCpzlsrj1SMpFGzPevVP+QZRFXmSvj1lKzrQ3v
Dt2ZtMVdAIF/XPeeueUBvWBDHkeX2ZK381Sx0+xkH6PwNkQFN1hFjvo9BOke18hY
Gxfd9TXIg65jFyR5lWz+Zxss8u8Mvc45Y+tVLJycq+TLPJBsBa6RPwPL4IfLewK3
Ve7NFsUQOaDhEz2/9HmbFni/wKhKUA94LgFkgZAUmrmhFdHV3hym8toZYvGVFV7Q
KRcq470ZQYvruQ9/gcNgRn4dusYTYRbZJont6/8ucNuOGYwECCyEOAqiwTGpyOBD
iGpyTvYbQk1AR5teqjgpq+PdaXwVZzAP08cor2pmDppFaZ7ykSIOtHUjhP5jNnbm
vZZdXWh5BQQUmS/N59hNVd88FiaqwTSjQd1rjuz79psGWFG1LRUHpgd3Zo6WEc0M
Jt+N4M6q1rQIYdtIF83E15sfc7JIYhmn1obl5PZH0mU=
`protect END_PROTECTED
