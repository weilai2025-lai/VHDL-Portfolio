`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMTSdfG+rqR9rT4YajQi5dY+pVFhhm7rpSskok4eDAcR7E5MaQT5WR1EmGBJ5UEy
ebQ62NMSAEFW4DFxSjJ8caZ8zLRh42wL2qwAVu7ceIE2tbU4zbgm7ofRhvsN/3Kd
kzHaHEwzR9IkgdHz+zXcFVYvIRPSVgxRWyo8NPlNK8ZZA2xZvQpu0H+d4UwldRep
ZONJBf00YGjSTzgYcga9K2afMSQGtClt6SD/snd9xRaXfQpDbsuwPc7Yek6uIygR
tlCkp5kexZT7aKL6U3DcfBUCrKmSiedMYmpIqH9RzmuONPsQUCAsczQ+f3i0xFzi
jV8tbbYF9kgayBGMhMkXv6uGVgTiPITrR2nEutHUZ3K084jjXQVHx89YXtYCPsF8
IebyGSc/lZBrb2k0NpFgcBmsc8pB8ftjDSqjn9UWmApn99nOPobKZ2zQjMJ5Dr59
vb3JOqNJYHPoYNWhyM5yMIeUe6HzmIK1s7rWFZJZDUdtcrlY/tVVnIasXqZZEx48
tkWd0JhLW0uZ/eRPuRafoRNRy8CuKtBfZ68NGwDaCrHGjWdxaVEPVSkfNnZh0Dvx
34Yitp9tXpZVNdWdYmFzV29LGZLzc3ssRGcnvNayX8tRIS+m/SU2KGcI6Eq6VWgq
UkqI6ePZK/EdhJJFQOnCv99n4BMP66BqZ9jEtxL5qIF9IbgA+Vvz2MYvrWwz2wm9
ILMcWYFMHYzEHe/btt5U1dS79g8TbDxgNSrAGmqXULVdpl+6M6IrhkKq9UEMMM5o
aYSAyWNUXpivDznSD5tp7w==
`protect END_PROTECTED
