`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LY6KAbl2qVn/L8p90HQyelWKkhsjxwEQOjeWxH5/4bi9p4Sh9od/vxG/DnYAhwuZ
pbTRyNPgwb1Qu7VE8AIBajuXC7YVItA4W2E6mCRTnXofQSy+SoRE73FfXhhVBXrg
ZfaJI0osb043GYXxeQcjuEoT6p5CaHi3a+37N/168uEtjDAQV9ypcLUoypmAJEO0
sSV1xV6dkn04U5ClQV3YBkGT05O3KDNczHLXCsuBwzwPWhoY3GGqmKj4odtRJ0qr
CtBtUPB9WheDocw1wjt+BI630xCIAMvPAYm7dJKOvM9+tg9wrfCYau8FfIKnmkWM
PVVkPnUsl3vmRPmE0aaq3j2ITPJlSLFSF200WQ093czIskb6BZ8o8Fd2xipzggvq
euAmdBdkoHM34/lpvjJChq4wcz8g8/8G/t+jYvPyhG8G9cXX/5XYeHwAdx+ip5KW
jGlkh+gUrBQq/fxNOUZqx77Cbff0ugjNCBRgGbF31L5ZQVmpg7fpOQhAexNbkkhx
MFpaMn06Wef167vCdx63+ZC3/hlHPTiivPKhMsh2DUkmU1L0jaHQvXegT5t7f3Kb
RwcKVbmx0JiHmbhVYR3i3LlK7ICGJP/svNg3qKtvRo4+y7MqC9cLODKPKh5U8vzh
bBnvlToZQ3Alfj3YOaxH+Q2CCXw2TO1gz2udZz8RYgMYaj1NiK6Eg2yfHrTpsfGI
Vw1N2fkZfHj5zNS/ttsa6pgREsg3OE3ru57ysSLjif39RhL/bQw6toeQT+O1Fes6
aWFEcJlxRsgB40VL2Bp5C1rYwqXMkFHEwADgjHdmW7tMY1vJZRQ4PchO9aiy9876
/xMLNMbhFMkYiJ4EdfNKZX/+cea5K35b/ONfKchbxeZoQFLiPOXoPW+10YpQM0/W
UbTFNsNODZlWbkx9ykTtRZbo3UqEXa4vAoKe6/cF9HRWb96e/akOhq1seeSqeMYT
tPNMXPdW3rzagxPkAmDzc8yR9IiOw93jSBMN0WPLZMftMq+4IYQMzYwjn6+jFK5o
UyCupC8EMV2uaK2V+ZJBeMVJs0vxNS9zUNMy9edTubZj7Ak9IDRX2T4QEDDLc6Vj
v6A7uLGPrB1upjeXagxGwudtvRAMoFTbSeJ5dUa1FxUxShgwKexAsxkmSsJp5ZUf
BViNX90EEX8AY+kEj7LaVzlHCgMJG0myL/kn68yejy5l31z2SgAh7LchuCvg8uMe
m40WGCj3+ULSFWBf6jpvVkWgeQmIdlWTNhA/PDgJQLJxiecxkD6maOMCm/G5uWYi
1SkU56xERxcfZvlvr4GZnuWCQ0llcbGkhOm83fyu9eG2/vfyFDjIl/5LFh6scrMp
nBqajrN22eUHoMqImgFgt2nqR8LaWwtvDW9M4UdfXgRd1sw2/2zNsv/tNrrwjM2s
YqupriW5mKlRcqd6sKRnus8cD6arGk7Bh1D+yUgseIM62ol7iwfSUfBSbiytK16Y
UI9C3zA/s9eYfrqbvDt6EPSyAAS/Z2QeSPgFnNsgZ3wjZ0MLeLV8ffSG3uFs82vW
xy4ptOT9qeLvuJj5WQcfy38KCZDfrYm0xrP1p/Lw5zjW+rsVCWeS2paLBVxFGSPr
S0tutOeXbj0NebcM5aZ15LIHJCCj1qecnwoqwsS9V5AxVE/enH7mszt4RZ3+VhMw
LVI5xNo/Qx2ou+LmvmUma9pmE2BgB1TSUBmBiMNCEQvP1n/vm41S6DBebS/1AGWu
i1xMN+ZY2d9GpC8nntpNyspcELDP89WD3DmvnjvA3ulKoVgh52GpoVX+GD9iNhaF
isaOMflLmNnz/7+XgkrvoYuFdbUDAD4HzTiqj39FfEjn4CQBZ/ou5LmiRr3AGstW
0PAKnuxQh0t/M0tsJzok/ecc0Vb47Xc/R1c1Ti7dbzEGAMK183SbscvWpzCsbNcd
LqRCAwp7XdePufjGRmlrZAZC8g5kLKhGpcwGKt40UmxcdCsSGRYFYIZY24au1N0r
rCUdYXV7PQL9v4OLPU+A5Ti16NtknIUV7LlhQsgwbOibg/RAgRoh3aw9I4h3zPVo
KJyrzoBVdoOWmGZv75b/uYTfIXg/G1qMQaJzfWP+WTPOEasSQ/b4+fPXf+oEb6kj
I6rBNWe0KgoZbrpz7jMKohZfdOh0jMttIWSN+499Ke+nTeaOpjGgv98vYGBWzNiJ
Y72Kkd+xtcMSeyg5L3Yc7vBRLsXl2F02m7BKh+jPGDm2Ue4ZpOh0C7IBEGIw+0cn
oQhokHEWtNKKmv0njgyGuHQD32MkquZJBnhNZI6k3tIhLdbn75BD4q7rD3vaC4Mz
19LDVVPbRF9m8GKW49qJbVex73n12eOnuulV9Cq4lJflja3rEvIyGhSAkNnyAb38
bWmdLnynMYAPt/iwXW0jlgDy6dLDkRdZB9YMLjZXhsJPcPSZr4+DILHTOq1il4EX
ooXGnzFskB43RclLVBAhJoIQXrRBzqhLYb/8OgRcfKo7yMOS7HJk7JvgtlaExIRE
ZHHhCgOGOEtiR1dFhWDy9A6G9P1StQb4rUsNprAKpjTJdkHOwbUw3VFEGDNRp8yP
8KmEtrdRhkOMxSbfLqpp28y9X6K62W99tukDVT9Jyt+VAbam24H+wHJzUFUf4vJ0
l4q1cd+Yqt5vi6spKHoF9o2sHn8wD2KugWUx1RQZxQhWjWxu+VjAqLOciUCRBOmy
MMPbzmSXNCnOmHWTQUbVFcNJ6WqG2F1PeYQbpUl82ei7nGsGXrjloqzBxwXMWOjs
KHpzY0Py2WywkWDjXK6ZZazv1PzlwleygjKb0xlMSY80s5uxjmuIJjTgDkho+TDH
RFpbBSSdBVlzx10O+6GGRlQlumHUG9U6Hf2bGAfCImyLdKQ+yKWASp0h9/eELzUp
aRl/dEYG6Sn+iD90ekM1amZJIB77V8SH3XClpp3RV0gD1sTro5QQ0L4L0f+fXiBb
Ceh1PbZLJnOpZtp8RwyGSvNYtHLj0unABz9Exyj7rBrOQX4Dus6m9aIeJlOxH4GH
hCSD7yEkf7x2XQeVpDT9TCUCp4k1rgsqMHwRLBPPQ0evFXuX8O69RpCMFXedHxmu
Ii5VhnP9oXo4gW2Ma9bEzOkjsNkTElbdW+Qr/TNxhHMjO4ZmjsUd0F8kEEAcnEBW
C60nQbbFd9zGuoRz4nF1BJZKKWPAYGclX2/IEFxP6eKkb66S7mu1f5bTY8kodOOx
1z+XAInTwq7rc3CGBpLG7QvUz08LB7JgDDLSZ4HLdUP5CUtaNII03VGqIx9sFVsJ
2pULkLHRnX5LG3VKmOE65zL++v9/JrGVXv7O2gTBWgjD1JWq/UsT/2/5lG3ibVvq
F6mrLM/1rAgWvBQbbhklr6CNM11brusVJqtbA8xlAauOW4gVchGhBSUFbLAhUb9w
A14jhVjm7RJ8tAICWJdfoZyNPznRkJObEPj9dVN3VZmPWMjCjerSj6hRG0RZoMDh
zYYjknhs6lFFPGnNOQv1PsyWFv2klDOQZOh0/DoQsLQL9ApoX9OMstRwJB71AZR3
spB1S7nok1jRQKWzufjgfR1xrCIx81Udc8QZ66wF8X0WP/J5AU2cgGCK3ADi3nsr
6uQEp5nDqdj9bbk7KL6HI2vdBLe1S0a/8c0aaBecBHo4aqO1D3cBWSr4WPmUgGn9
ZiJUar3We6oVz0uREJIquZCk7R5X6QAzQOR8qep5Ry8V4CzUAjIBn204ml9v12hP
N+W5mt/KhKe1LU1TiZXg5S3mbbYP/SRACCMbmtp/n7gJsEaz0dVjmwTmg7cEF1nC
bD3N9cChlYQ1wKErcB0Rr3Zqzb96t9kexIxpylZ480i3WH2Xfw67opbxLdlJtUL7
fVCIyh3nl6BEraYZfuDUEKQLEIb52qYO4bq2Zko/tOMXd7OIf5Vh55+SV2G0LnR9
IWwjbpk22H3QhsoFafeTVbfT/Q5yLyKSekwj1GbsC/B52Gh1rG2HjQm2u1Xamx0x
Fy0Ucf90OqT1FbbBJA0WtlDb7GGrSB7Amb48NI0LCfXZUWQdsnxbAkTUWArm1YmN
YTPL7tZ9kdaXGVLpraCrTXssMTqwOwyyDulot7j8TYSPvbuCzgtnNdVQIv/ykEPG
6/OXM21aZakiHOPJVDiuPUfqwbN7K2wquj2Q4BpY9FCFswQOXLDeYMfDqx+925rP
jYyWf8MmsYXznt34SlgOC/s7w4s6F/eccssQyxgFfsCjVWU51uoJ98tKidQI90WK
2lnpunF78TudHCeYoJ+LfPo6F6yKOgawRKE214v9R3tVaPq4SYqLNg72j5X66jM5
YnDhY8AXTYoA9ERI5z+O0rxfgxbNtGEt4hqZegJyYzDBmLiJzkoh7o69uILi2+Ct
CpJba6jbCZdS8i4i7KK89RZm9mn976rThyM+79viKWGqYHaRb3V7XmrgD198TVHh
Dp60dBT5qIr4aeGTqhJaGwupAmMXR2P6DuZSxNuiHVnQ7u0fozfRZNAj1FNZYpcS
UCyCJTKvc5TIfgkOcG+kflCj2iIrjI8+RwL4e8jop3a/69+SZWdW4xqyyWCfu3QF
Ot5Q44f9BpVcKfyjg93opi8DnBy+bnOqCAWRzQmyjuMW4UAliRjsRuCVODM+pfMy
jggarMnZp1JmAW9ylKA9dx4umo9gVeroJaYRtXSgprXGaqGubQN3C3HuTCErvpPs
5e0YSIJxrHwnmYwxCyrcO0QRDZMIbxl/0he07xxXjdbchxtC23zwaAMH3EnkGTjo
1z2Owu44nY0LwBpIDAEiX7GAA+UBhPE6rpCOew9aQJEpoPwCK5AfWf2up1d+bJ0y
62MI8+fPsr1LFSQ7+lRbSOkk1T1vzeOILyhadcO+PgPmCJo5dxlH98MOwBzbpHMQ
GaFFXg3MwMTB/LJaxuJI5nALLLHxzOTYsBQmLsYlG6XRjU93Iv3UMMR6q7pJ3Hqq
ix/4II1ODBREVmRaaOPGZscz+buB0IfadSw3NtWQS51Vo7+wU0B2LfW8HoA82x7I
56ZIHAb4Qer8GhQND1ZB/ht5rpEwYmuLD/rZQIPodXz2mb1vkvnn26PU5aK2W7iT
Y3/ekAYhvWGWxjINNQ7Hwdlpx6A1UgKzY5cm0tUex70f/5pYhxwM7kqONKBQaiAb
GGPVKQkeUG/GGMH740Zno+/geqnusZgb554M6pS69ShCu0KKQFbD132uuRYKAiah
e4G8flHpFC5oaddZXW8gxcEsr9UXfEgicoJ4oteEP+AtI7XbOUlwo2Np4FlxT3hG
t3hiwUMW0TjHqZ36CFXOB2ACpU6DZ15hnc7vcIyhRgJwWNrD2BaVXYrGmmb/kcOd
+c+ax/kE3NavIJabBV/orskW6uAjsCukgClp3ma2m6nC4lPgS1M+B/GpJnzViff2
g3Oc4GVHkPThtbIcCOnrzsT1OASv9okCr0UxK094ZGp5lT+p0IJ9i3D9xwO0ozXP
DProwAae9vcFG+k657DMDPsSyOea8Pw5KrRMoiFgSKwCKRDzO3vcPmkylWP81Ncp
tsEHDM8QOm1Da3zPLsvOB6VJpoq2UJfbtDjI0QlMgwGeDJvs2EmY5CsoH20gUrLE
UNVHNCi904QM/BhmicTaV2tU0JLtLV6GXXn/dBIxVEsJgKg6+EMuy690NRnUytom
+HwRNppe6nem25QoS6ok7eG2E6Er8w9H7HtUoP6CyJa9J/AQLN/SPByDq/pML5GN
9jWC54RbfB0SJxy4b856AoeyQk++tLINnNBkgTGk9GYrXr8sp3eZG2UiEhYn7Ho2
s1MEl70+2au0NlR0W8/KYMR62fBg1OWjOAKTfchuPQlqHqdiHht0zZz5xggU2oGR
iTlbJDRu9RQ4Kian9lKUW0HF8PhpIi0n5LLWqndlEoibmkiwNspdGnvZlhpREPqW
P6+CDNLOl06YWoLVJTKo7r2VtPDSeZAcrsyBZNyYFpRpLdV1aAGGGU+xV+uQY/mQ
q5d0/y7u8szm84i/ao6mHwrkkrL2Yznn3hxafhKf5Xaa/w3SoFOtcXX9LjCoQdqI
DHU8Qo/j0xkya6mt64F1Wz6HCAGNb8pHMQhrQaxT/RejT1Akw9XIkgAds9Rpf7XL
m09OkOdgAwtpXtRawMuJBSj8ueTaE9x6EHdU9CjvzDDV2vEwBp9GB5lFBSXvpYpa
ay4c+LUnOBCaz7Aq51xjdNCzRYCXIAQYsUo/Lo1jA3ywenXaFdGdu3tt0sHdNeQ9
5syRqmIRt564fWvxMncVuF5m5NB9h288Ak55vmJJ5jr1NleiW5NPIn2PZy0HSEmx
03X+pqAoyhDFkU0K/WCtEC5WSihI+Ki7ke+xZHeG2YK361MuUpl6mSUhppDjAfXr
ffhdw3WdRUh+uA0ab2nCJoO78CAr07OKEu7Ca4RyI8kyf8DXohm1vOPtfoAF6suJ
sne/xZ9+5oMXfYiaYZcCXneo+8BOryX5ErDLszo7ljHMDyfffLsIHUpBRrhP1od9
tj24nJF38ZpFrVPc+I28kxUxdNV7hpknA1JkE8PPmZMX9Xumk16e2cxQmNan07Rw
1/JsJvuxbbnJfK09PMFlgrnr9a4BXFUrgzkCP1J0ZEiXkqyw8vMdIIw/zftU1oD7
jNt9uUomuLEixLjEc7KqSNoPbxQv0A0ADt5yiFLT1ve0Wrn2zSaWX+R793PgK6AF
kz0Bd+vsBJ+ycWCPeSVcy7O3nMURneFZ8fe0mTL3+LCJO6YmUyhchtrXtFdv2c4L
Z+L+o88MIyr19qfnrFn2iXJaLqkdBkyr5gfiNa1W9BqzACVp3zQ+PdErJCnoL7hS
VROMykzNIFZsVOstEDW6FpX4W2cqSTYzeeqo1JWb+oAyzyFyXcEwcwozTX0D2CeM
JblNDL+CDtKWX2L2nU8r2wZFBB/gBl/hXCYRbIyaOAyiukWCBEdnq35A1mVJ23tZ
oo4DZSaAjspj+SVgvCcekq10CSgbpuZL/EZXQQI/9uSu2caIJFV+borGLUj72Mbg
i6rtLnmOYSxbck06cgHBlImqXr3DQjF8Kv/bYZcZs1yzLlzuV2WHO6tgJL4kQqis
xrR7QQs90Qt0mdOMcySvoT//ajwmkjB2kq264v1lRU0wxLJO6hT30USvrE1rKGg4
S5XeI/lc7SztD9Vs8S0nLEotVvxDyerlYMnmC99sU8bKcPYDjUnp9NqRx7D7rrDZ
qgW6Bsebsipemi8Y6ROenuqgGJapWgbgqp1mPZJY3ZqNUbsEVMGMnkzDOSfY3src
ZEjLYAD/BZBRCNctngIlXKPACbINR2+VR6Tb5sVj6FZXwihhm6PGdsyuDrNGjXul
M3IbhP1gyZqGMfrcC06RmaqP0AkCUG7an64+xRhMnFP2waLb6Lm+aY791Fk1+Zdy
18Xbvyg3vpxnPb1Qd4jqAbp6bvqV/2/9GalRGOvnIWXDH54XBwacgXRyAJk75eOD
bxP6L9c6jYXkJNvCeIDsuDTYt4gu8PzTIjxL+UDDFisbhrVut1y5YI21rx1Sfnou
drBKEtDqfO3sei2BpYdaIbgg8XUzhk5nZZs2IFWBoMi0JaQqfbM2gTiiSR1zx7rF
4wva2kICt9N9Uks3GkDBA2C9eHqiQZjHWZxFwpOrlOF1dn9dC1lf6io3cA17KFYh
TtGAbpeK27Cg3tiqgbLZZvNmoFGDZjVbHMsHlV16VsFVab0uM1EEB0lzAM3eoSdI
12y/juy+Jm3vA2n25KTNSXOEPzUjBTXP8mGCurPR0Eqmo0LLbjD4xYS1lkIYzzQu
sePiX2Ic54J2+iUQvYUjrVOSU+nCO13xaewSdBb7E/zNZp+vNK4NeuTVOBAku0Fd
qtJ8PaxCufVUkGUGhMEeZu7Th/p1POBDzDP9/z2hOokGRCltPg64BITI87hElIFk
Nz460+ZKCGoquSZHpsCpH0C4hq3CHjYNiHXFld+6kb4gZbMzM+qtgjYNtSuqhX8r
AX9yCAml3m22YPD7UTzpgGw020bTjj7DH2e1ehHDvNBQ5940udzJROpw+0sUbWM+
n9JgbyQIJumCdjdlGPQBDyhDgh5rZFBZpqGHiy9kbYnEg58EgcUNViJQXu68TRDE
TLrYDWpcw2sJHDInmQurQ7jBCUSTc/0cPi9ks+Nme75bpZECaEBXh+YkpRc4LLiD
0RAq5chrpSpHivox2KGdQxHGO1wb6FNH9/QdWiFvLTyeQho3qGQvhR5Rl5+EXN/t
MNYatFNPaASIOkOqRESrccQ/JAujc66mfq4ZrsqdsWCDBjwpleZgfI6RK4F6ID27
+8obbVhSEiR1cvCOWEKJrzP1hdDNNKz07WTQvJvlmrzgzzUmoS26WjtD4M1ShCiW
FDpck+QXcol1goN7yw6paUealMvOyMB7wTbZuHiSfLhE0Z1dSA8dHkAqIkoKvaQj
ZyMytnWEZoLSJf8VpzwWs4i06PFKC3j1YcGoU3Vst0ZdRETEV3EIByEAEBWANq8a
onV1S27LToQF/yyH+WdVgg5kbJpc5bX+Q8Tmj3pxCTM7mCLZja33pr5VIMAh//w3
S+MHM7+wUfR1irF5OBhD5pLM4M5BKvSoI1sjafsI3hOjYxwBtwimfULeoK/iaauQ
kqmPouqMEEkDoMci8crteueP6pFt9MiE+M2F7WPluu8v8G21zT5xgozcMLXjoX4w
0ABIZPxXUJsEoPq2jRm/FiNOXhpC8v8GaYp6duGd64SXqqTPh69cB2W/8zbbaoiN
aJdgyDOWfgf3S9nErX8B0lgJxB/gEtV451GKixVj+ja9asuUHbkqOm9u5ASDHOaC
JbDM1/n7SaVqrq5KFQs0h/xIPBji18F+au43aQg/8lIduphx+NBbUqerQ/ZNrnN1
mfmwu/6nLGYKdBhgetjVSAFoUm3LhSF7kqZuhBDMYIup2BI64guEySHxpEj+2zle
tC08pBbH33owutQ7f6TKQhPS/aKSSWUATcJqtIkRwgvQrX7eyg+2SB1CYABXI+i8
IKZo9XogFhYpr0HyEa+7bPmuU1/e4tJ+e+yoBBYnBnoOGWmaVnp78cOxD3WoVGP2
8ExJ4k/LPAPL7W30qZFFVBdu3mxdeN6QyKpvsFgsP0w24+s/jBSLYYV9iFumOUbt
XWQnWM9yU7bvrX0Tow5+IAIETH6y4Wo0fnzCOgXjvnX4UzN396ddZYwF3yyPg0pS
IBU+Y8d9AmqGUC6XSUPeDgKU9IYikhDG56c/k2CYc//4u474I2v6SAjeutP16sXw
XNI3G52VjphzWqeTlE9EglzdEILStLPyR+CpEF1a/gXs88Y1oZsmQ/DaOVX+AIMH
WP5XPdubb5c2zRgbqb+kkrfW+xgvkYzNLLGzNvTJsMx0FDtXd6uqLDBSE/63lUxI
3MFTDohmKWxF03qKVwwbdO8pNIcePac07rIhH7raUsAS6HZLaT8pJveS0yNSy2YV
AA1yaMffv0/EH9Wl3UjMDCXb61nQqvzXCK9Elkw5B2GX7/URN/V1YW6xYKI8CuYV
fw3XOA/svShmodPr16zXRQChzHEFfXhWnf4S16cznSRXQLCQfsnvSz22UOQazOvf
o5UiEiJ38FBeDVNeF0yo4Axv+owxBITIi3XaHi4fbuENcdXvFuFmW/ywgUVt8uuu
7VTfzc+eb2YMbNVgmDU5f8IZqJ1Lzi4gaBZ+RQZQyXucx0cjFCRgV5NyAEyzhMtz
JO7Mpa9H3u9YABZKmNAQu3jorCclUjkSGNYH2dq/Q1mHaCFUOzwEwyG+j6VqbxVR
YnRc2KZSIggZxexaMFc6wYGea59M3I33b8CJHeqlqyEykd1boLO9fVvU7SgPOe7y
Je8+64BJoMok/eCawdtcFzyMyML4A8zaPW5OQagIPjFdO8FepbPcAlg7I91rsnHR
sjnLx1izqBG3QIgQvDERQlgJ9IyP1MdO0p3+UU8L9O0eZ67oOrOdaRTq4Hfwjl8b
WR8veazeqe8pesFtbBHwV0yMC0bvb9UbvfMoldctLx/M/K42erSdfpr4TfP4TDQF
bD18DEJ9Ebp9pTKx7wfsOI0DZEGCizcq1WcyediC6iEOz25AMk123OZ5bXl/b4wo
i3DuFgewuiL8Jxx1DF8IrmVLHxaUV/O56Osl501NBvZwZuALe0977I2qscbWhykx
qELK6K3yAxJcZa1IuMMY9A7tH2EspJRbti5jArBY5fRtEqF7nVXDOz+DWk/F2LTQ
kJPCLk5yMoFQNjNxBCyXdW2N7qAyTwCvntgpZRGVDAL8YFXbQKeqIORX3LPOwc/O
kukxEcV+bbty3yOaBymlqnn8+g4pYA0aTcidJJM2nhkOzXe43JPhQ9JE4b1f4Ury
gaeKTOgQteFV3t4Ttxi2q90HMhOovHPjbuPafgbHzPTdZq+xAUJNcbx5rSjb3FF5
ZcXLHHmD7QqZMs25eJQlAlocaiw+uzNSqZXyVWuk0Ori7z1SM97kID3H0ka69vyU
fzWePzCxE9R61sj7llIKeAqtf13+Q1wCfcOml2LO5hiUikRqyWVHpG0Nna16bt4w
0C9nx2+tOQoZScmfNuW9JH2k6pEghceuLdfX+Q8cYdbPiBVMN7UfNPuFgtrGby5K
lewSPKvf8/RrEfgkqB7AmFhW/riMCcu5InM0ghxjkF8ZYO0Oiz/lxaL8THnzcm/P
w7neM+l/0PZr76b0ySlAq/hMOlmgpQZJYDwy9t1ZEn3Pz/HZdBq2WUf99QmaLSg5
Mco3/SsMwFspakZvg0f+Jf5dIFcl6CMtgnjnskUADp1ZVLXO1nhSj/uKRWWvP9vI
fcjQj4IYX4prz0g2wK8fvL5grOoK0aYRTf3pFoh3hWRr1s92nZfFQ4UcFlsk/Uwx
ba3vgncF833EuUQFdNwZmAoJbNa5JuftT3VJkQPSbJp0BiSw8LKId8Ozx4mI0jun
Vk2afgadaDgUo+rPDz1yzFYUFlEooQGH89BOZJAu8/G0OI/GYZ/8Mu1C2iIg5exk
mw9lbOq8B3iRii3wqYeEOJM3Pi2RI3OiBJhSaJiYlHKht0zTx4FeCAsEVUTl94Dh
k+oEE6Z7FuCTS2x+DUZGNnc9tsVYkmT0NtzpjemHpu8hOuDHsctbyAiLB1V5sCAO
92eqe9Z2GxdEsoSOJ54ufzu6SZeu1CjAf6BSDkBKHbLumNlCsfh6BdZbkAcM5zYn
rIjn0C6zKbGG3LvOqpYFM20fJE+NSxzQmoYgG9y0nGsxlAWA1DFkOFmQm7rwApU2
gIr5gVgDdsKegaGRXYrfHL6kJ24kbMCBGz7Wq/Vr5n/SUUclT+nolMyskkfPyhFX
Gc+ug7ZPJpFnuWUcBP6ylnStmXvT91dijNmeyONFkE+WuSEC7aHrj83vnEV3hL75
JTF2QBP46OOoUZB06Sqlr+xb+ZUbJj9Mer0JZY8zyV2pbFZGOsm4c0lfm++qVpM3
mvG2zdKUPkxJ+is0eBmOUEBlOvmfe78MFm6soMsYRNEOPXl1vFrA5rxxw4jFKNZY
CaWTgoMLa3fvim8vKcIA169IUAPrqQyCATAvXhVCdsc495tBmhYvKx+6+X67+i+d
dv1e8ejDQUxdvX7fgdos6Wh2clG4ziv8xo3aRLscPyeOmT+StBCtw0DKSkoPdiQ7
SRikCyyk8p/fzJXMReoWnQ/sLgmYicKmgn9n35PmWyq5PuFvYxXb5vHNmHE63qvi
A/7h1UI6Uyds3V6Jjn1XkmIyhBId468y1Gu/lxTIS+NJ51c7QFBDihHq35IQJLEw
lnRZPySa1+faf532j28onhfZUzFO42Kof64rxCiW/6OiRmvMwoUSetmeI2cgbFPg
pX/Q1V2dME279UWcNx9rYbD3fl4e0jMasjrPqdCpxB8UsDaBrkQteALVHFohV5xR
tPD3/AMtO+/1srlkM+X6SGW+qI3FXx5cQY65AuT+4m1h4gcXoomIG6iArznRsz3a
hmcBZdU7rjxZ+gEd/QR2+N8yyuejfcgZjYis+GJ2IsHDKfB/krgH2id92P5iNgZa
Ckx6iQdirvSNGPaWsEiH8islsCS/63DFiKPgpNtVL43zEMIAHPuoNoMAcj9RAsG5
2tzjKKfC/LQUcBEsQ0lFjtLrbEwZV0tkC1H+DxvlzfSz9JE0ZLmbP+DVQgJVT/bQ
pLAIozyBWJ5uAR9LsFV6NW9gCkFwjWrjPnSyEX93EK7ZPIPgZGPN9v9oLQwaO9SY
HyfmJyPOwqXFCc5psk7giQsd2GifwBrHzuCB49aMPOOqDnID3G8PQCf49R0C7w1X
sGpxpSOnhc0+Z4H87EKJd6nZXqonLKmg/uHgW9JQ1vkDdRV5nTmqBkhG0zuRG5RW
jtHEg2A6Ryh3j5URVCDOZWx0diNk66TUjm1FNccqrJghe7x4LE8caycpovDb3A9N
NjgwDf8o5eu53q8oXLFcX8cYIhoxev5+2YwHoedSSafaCUp1orlmV/Qi2oIy89UY
uln4j43/51SW+poJ+nZP3LXQ9lwzsVHjsEGdbYuA5AzabZfFoM5R/9Ydsec7/hUN
coKFZ1AfZfkwNyrCqrJFvJXkdwRj9ytCM/Q54Y5rpxAQl5r0G5tnhkPv4uGntgPf
EwM69moQEbcr1w4JpJ0aygll4nEnnxqii+koP+8USHMA7uU7+RpD90kk0RnPcMVW
tr2EqtDXJFkC0Ua6c/tjyvUWZDsKVzK1B1jgNh8PcZXyzkO18LzGVN9eZ2v6I/Hi
fBQk48NR4XC5hCy2JQPQfoh3MPJQ08VweRVkHqX5D3PPZq16OhzyVqxXvms8mSzO
BRL20+RhiKSKx7cKhBE4duPR/B+I4/zIImkkmKAiDCQxlTTQPVyQ08BIoj7b3dtG
kqPzV0NcBzM1sQHigz7rRvc+Xg9bGe26hdOn03zEiT6raN/pWA+wCR1E71QTFXKm
sBXJ8hX824x95Dn9vrYKrPLZWzWNqQFH9MFTXQy8y8n1oJs/X/V8XgNctYgbkL2T
ZlVzDxBikqFS9OfgpcLryQJzUfLe1PfZAbQHG1lHGlFdiMvv3vIM1u+JSy7ovq+I
IdCKWtfKMzmUG4vI+LGFro61/mtgjI1YcW9gKYEUlWCy+tnrd6Ew7mwS+oI2uyZL
3VbefOEcuSAK2Qn6QOZ7ArnhBLT9sv2BtbeS43x0lLQV6Ew0uKAr+9I20RDLc110
SVjapE/VRrsc4fEyIihz/Wpe7OEf13ti4ezMjEN+W5kle15hU87qBekyDYomKTDG
DOHhZ1XNZY1YYnK+YEvMM07K9YD+V0N5ikwhKcE7BEJyAq5BLCKfP7hS5qUDX9QA
k3bXMsj7bpUjOPL+9XvmeFvqltr12CKMoP6yoKg2gLhEm1o45GliVI58GJ/BgNjk
RBMbYxtzVQJPp9WNIer5/SHVCuH/popoh/p4AMcMBKvk+XWZpaoZLPT/v1gZTuR4
orhB5mGMwwDjMT0ImYvIzOBCUhD4kcm5VslalZZfrolvJITqQNKfnhBbgBX5uDGj
hHhLzzds72XwmekaaGsvCoURl1asNg4zkK0+Dy3aULSDUpFDJH1ZQk6Y2Qf/B7RK
WNqIdyg23GprYGv77eNbqFxcpIha2K7xV4Wl+SLz8GKW5o/uJCx6Em0nW5gxQA0M
oPskzXW8ZzKik5oSu8YPZ4WmJSdMlXNMMSsKWI14KATi7/sDMq3jFjRGhu0BxEZ1
qD7kkQlG9ow6ZJogAGABL21j7yJpviXNl4LqgPyyVo94gmWcpAQAFlSWrVVqhDkm
4crQJprXPOWcG1+3H2CgNMVajkkw8J0xtTBzexnss2r8YAODd6zagj93YD4ZBMgG
kKlnNYWujApOPwizSR8hkEynzG8KnOenkfK01gDMHnd2faz5Y5cj8+3hvBG56S/w
ZHctEr54yo7tgTmrSJ16bPrh7D6l8+XvE/qnSgkp90559dYldLaoUbhlIkcduTlC
Ucpl2EvC+OCObEYqb4Bs4l0aghTT6xh2ph4kY9V2g+gA1hcKRdjNaw2rbRfxc02s
URgvJqOSp8cAHVuuvqBbnAVbDjL6GTvNPjneVmfSdWUOd2HIRD/FNtfWYCUUVHYx
mqyjA9gMMytLBVedZduf5mvWjnf2XKI6y5CwG8T8wI1zGJfdMxtg4/RrDhSqbCE6
JbZFxFs/WCwCaB7Xeoa5dZUkWK5mX0WKcALLLecFQNtvsKXrDXZZuQl/gcIkWUa3
DOtS8vEejY0npVzFX3ELO0huhANqK5f/F71wEz1vlQyCIujctGdjMf8jihmlb2bz
N+7Vdp0IdJt4EWtWl4jICejvqLNPpxjnxp1X87PTusPMFc8/OyPeddX+7pJ7RUgD
dRw+EU03Mle0IBZrREOCdxG2mxAzqVGQdfFPVM8HvuDOYC9QjPDTIdiJoFETu7Ye
lPvuC10T4mgyHHoKMszYVaVwmb7U7nFEiLuGe2mfFsLqGXGpt4cZcWttf1g8YxWK
DYYkbU1ghBFRl+BNhzcAsixnu67HmTBMWnHM0YYbASty0IaUVCqA4yCnZw5UMdQT
HoiF3rvAx4FGoR1BJhsECf/8PbOnQPS6oOAHz5m+dKJqU7WLnt4HFcHX5v6t8R3t
KZ1WD8UPCV1urVJm9zePCTEFd6mLmDZxrO7fgc+4KR25HPFyc6ijKaowfM4IWdUz
D/aee2j/chmajIJZLXzyHi4FF7ZorvdwqumNs4JbkUWECOrC1l1jrJtuepG/KGP7
l0/Wt2ldSQkmPCno7DHDz8iDo7Dy1YHtBx5+prBh00FTUf0lbaEEPleNlhOkTUlz
AHaOEIDxv428fT4LUSfuisT1zJK94MwwI/x+GlubPSj6MgcOAiTPZry2qkR0aT15
wlH6rxVQQBgMV63yXcs89I3KfT+/WZ2oVGRyxjeelu5nC9UPr/GIVC0iUI8c1s3a
i4rrBdUrpqQjo+Q7N6em27ekxaz53YMO99bbFQhiyRrLO/zXnkNCi6UnKzcGSKmr
A/D08WZd6UHEZlyqDgTDa2R2ZDk6k3ib3ayZMhyjXZC/FrQ0hpVZRE76/lSoC+im
XkbdZET9UpeR8yGSYRM/WMiV8iGmsLL0XxRg8/ExDoNd3VLqUTK3w2vei21Z+X6g
7HN3//RL1NAw9DE1bW+TuOpbFuapqj4xytWh9CL/Z50HsAJY1KZ3BznowHWdRsSm
k+yk7RZgrQDZ1cA+V+YRfebwaP6BJUiDBVZgDZS0DY98EKXD4/5EEdtTGDofaHQm
2lvT3OGV+uhKc9OFfoZ5ZEXZY7dY7AyPYkX0zIKmcEyn1yCU/UcQLdkmSQPDK+kj
KzBmZvjbBP+3CvJnO2vyE2Omhvs7rtExsR90f3SmbP969I5+xEPfpn9p76ak3upQ
h8JPYuFZNqXLEdsxLgWYEExRq7wOGASWalnMr9kfBdS70hkrey+y1a1m2wQ6Tn5+
dVvOHH07orc2KLxh+CU1iNtt5W/l7Sw3ZROHkH6ZZx+NAJxEO6i86FjBv0uoCuFr
UAt6qVqJ34n/l6onaQNPMhW1KzxqDeHDqGc06UtdrDVGcco5u2pr2AuxFchGe+2p
uqQtTXKnVyOibrFpHk7spWw7c7WCSIU4XIXI9l1z4KieSMrqRlOBFGhBEwfsMJIS
HSB5UgLbtqJBwEjMGBb5PGpUYCS/6ULisi1z3TrfnanaaQJN4SOxOdJ5IlKzn6GU
cX5wgdSE6+1aAJPcpjwPlnIBEdQl1i0POfOHJtL2H+dEtvxAMw1CVb15B7HodZdz
zT2l8ubhGVAWElAP9hTcc+IlEGBTOpeFnFS4JN2h2VSwuSce6dmKDshpVZB1rJn+
Pe+aLf+cESQ8tFQwn6Y/OxTbETTW/t2+sDqv80h3ckXJNRqs3hZr8PiiozfyC4+9
YBRiIBfJMjGDZCgI9qCAciO3J0Dc5sNfjire8SFGq7zOmyzJcNud75PiWfAW4E15
ftcPsglJ2/q/fxzWFpBBn6UsOucTqTWEqMCWTVJUevJ688huUG1WOv+ai9RKKjg7
WyLZ8+dH/CDtZj77DhTj53DZvwkEyD+HPtFTu9JbJDcI8dL55Nar4+uU2t0rE2qI
BcPQ4Sb6gkqi2xt3L9W52kJT6X2LnvPZd7JIfubUeCQykXVNEhqGtktArxcUJ9MF
zYVc+HHwzoBXpyE4oaze9JzJQGzEhWPOXJ3ay+Qe1ZP8oQCz4JMA+/vmqpg0rPER
yF8iVWwX3uP74YNuYa7Rh7qjvK7NnwEcrDd/SiL3zu84OF6xbx+6ACS8jlm9zJ9s
YyuBEfUE8O8yPgKLCFTM4YbvVhY9/ZXnruDwC2p4SqkvPIx1TAHf0o0KEzVNhkl+
7ugRlqdnf9/o5H+n9QZf3LsGgUowcNv71ebru0F1Erx1N/aCoU2BhS3BENV28wxv
RDMMhNImjj5Iori/ekEMQX/Aa2w+Z5x4PVd6AR7+hTyCDXVSO1h8DVAoG8cbtMdK
9kjqfmPOXvnlB5A71O/J5ki29MoW5319WIXBq4PyUCuUotAYcT3FaFgPgTM3nOgR
1bcEAMfeEg35BknSy+YaFbSR5/SVLH7PxWDdsVxULMJLdwyEDaHAyY8AoooYshyD
eu5INjpDEP1EiaCyh8MELRi3Bvw+0S/otctGaRCGqcGktEQyzoBLj9zmgOAqK5PA
PWbI2oQCXoLSYTtG8NjF0ZS6b50z7lnWuTeVYsYAn/VJEX5wzRgi3vXMM6fLUAAb
nlWlGa23X3kwdc2C6NkSHvfVEcKwXvdDllTa51fqpa3vNEcc9eXyKcG92lLXeH2y
bDcUV7QxaErb7ZL22CYxBLF9cgPYCCcVI5IZvmlNn7+4VIoeHlMFYF8nXkFOz01L
b4yjBJIecJVts5tPO51F6xt69e9ORYygN//lGuYkdWHASW4SRCMOX19kl2Y5IhEP
MxOmBNUrZa3fsnk/6fnttpm0+PCH4QKZhSq3/EqhnWpcnE9tKwXB/hkpc4zgBv2b
eSujWsnEM2xGC0vC8VDEghEVzsfNBdI/0RP+lH+THr9lh+X8YiBPj/lmOF5BafPa
ube1q2aMeLLcDO3pmCagVrV84eLmJzIIxBC71OIX3zH+J8xQYuZ0DL2O2zuiRoos
0Fk5rDVR6HC7ByM5ikyh0ABWcXaZ4P/xGVwTGErTKzti2luR+cCah9CWDPmYxrrM
tl0MKPgJiFpAjKpSgTL6q/o3AVCpeS9aMjp/DdVlRhNLf5IwKaFqyQHlulgWpVrX
crzaRUGqjSBCOgL6gJGNYLCE7PtJhrpS25HKJRXlpxbmdQDNGL3Lt4JpXDZ00yNy
WC5X00GlxwxW3mgOymYea6NLNgkQrydNMdrBpbpydi0bgs9wwau9phSPBT7ESBF7
J1k+3i3QfRSuV3s7bK1LqVtAphG13+o97CAiWvxl/tik07tANykoStbocF/6gONK
cCyQfz3qv50xJjtR+5PBdBR415FzMR67Qo5hx5VQkC+2WJGiWOWoyAm0sveitFPG
61NNaVoB6Y8JqD8nqARgi89kJo6hZH/HRYB/tEnEp7hDeabk+o2uG2ciwHKKH2iK
UL+oavY8dmxhVidf27XF+syfp2jeTXdiH9M+XYPD/0RQkr8dc2A6UFumhLDRmJI5
PCJmIPlxL1X3vFiZB1vq29hA400Hj7NkdTArwy3k5MtRdCSYrUAvA85TICP+yi4d
8BkTuKEmEy8CN2h+uJ8dmBBebhTzz+I2u/iXZWFP3JBghQsRIu3sGL35UegTaK1W
xqmX3kDpR9LfB6FnD+pOKVRGkwj7J+q/Xdza8lhzJubPHdP5bIGr/0/bGcGDEPIt
ZuVnQtELwEvdq3ACDkjEU/Mh4F1OtStvb0yqMzJtL4d7bs/uxg/kxoDW1Y8ypZRI
q0SFxx0AwFaV8PKkDNpaESiJjohIZ2oeC1pvPvzCxWPPDvzxJ2uLBF4Sd1t/dIAh
lP9Lnlu3yOd9IrtTehwQj3mhuCqdGC5uJBElWjbhP/R8RtWfEl6Rb0CoUtzB1OI2
yqNGE4wqjT+H29rqeXTsW8cP2q48NafmGv2t8VRAivczqd5Mhik3ZGrF6/V27Gmj
1wNZXNjtUvbmzsgo0o1wtJIZeAEOSpKIPjbYoST5kfV8vAUv3xmx+DsaOuK1gJ9I
GUeFbV0FybLzEHDhyFTHgDth6GWn3Ux05GJgQDXqlmMv9oCc+sLrndGWNcf/jniE
zJsW3qRbeVtCOtkyVGBrA9ERgQuJuLzVHlRNiIAu7pJnX+vCflGRaGC0RPPrCjeJ
JAWNBBGU+1R1jdMHQbfcCj3M6LNuuqJyiBqc6gm2OIFQXzAeVeltdnaepfaSWU5L
01xs42iIkYer/dca+W+svnUbJ+TJnzk3nLtvc2dUNqHdmgDttQolWdFiwi9Pamid
8+Kb116LMKEEeab3jBQHX5Um1MoFKEd/cfoGjTSEVkB1CHwvydGyOqW1L44mtRO7
ZXjsWOR9ipfaxIVlA50bR/RSQf8Rkv4SLnhmmCpo1n6K5UpmAobax7ZWB+zqPuVI
pujzqddXjBx+vZF3dA7oloic0t+8S2VmgBm149T8CsTJXEiK5d0xpvBYReBQeMyj
1cmQAYW71SI8FaupmGK7vfXAZBZ4cmdMLWar/n9fVukr307Zx6mqk7LZIOxwHcf8
UYOPzFu5/GGyuX8AhndAtBl1JZMj1PG1FYXDYxaS0MfX1AfRqDqN17Hj7pF4z124
AZP3mFbbzx+T3E1pK24JzkKjwbI/a9UNd96WE2cd+XyhkQe/TIzIgVkA+NrePQFE
n3EVR0AtOzaz8LAhurW2dPVSso9Xb16AgPPx1LetgO9nA18bOxe2xbz7Z2u+vOxL
kSrowEirDN0wBjBcnJsRpU5b5L3XjB+8eVqOK0HXhJFzWE9WSMnSwl5TF93LlGOA
mgqiJVAD3E/4e+zuwfVxznofVpeDvjjyyhBL6HmH3Z/2+7RrmAPNvO62JSMEYgE5
6zvH84oh+1HWF+JE4nohM0px+EOAZCZU0oDmBJkrBuMtvji9AMR8xW6obQpf7AZ0
qJ4ZYqBGY1KjvekVFiskSDgBOTZniHX6g8A+hdy/yQWC5sgRp7DAKPae84ZoVlwL
DsIfcvJjGZpYtlKap9dJEhnTsYYgVeRsvysiU54yW7oPO/oOtfeM8eeZpm5Y3Zwt
939ip03xa9wYtIJA3KOze6WsybOY2jhx0UqQPiEZmjMgQr8kF6Zqx95zeewhTI18
krg40gy3jkzE6mjXPo1vEoCyOChnZNmDeTNLfyUhyy7uLCehPHQSDAKz4yd1dGW/
GJBVzcLUBcPYNMDlxOsFQ43bfgcK0oBAA/JzgQM9o92pUxK7zwZg/BytVFobrpT3
E9bGMh94G0EHC8NvNVYIW51g0Iyo/uU8JfknmbJh5DCpKNxnIyN34m/0gCr8Xr/i
ZOQksTAosK+tmlmRgiFTqHx47VMzc0k5DCM4kyQr0/iRfD4taceTC2MG0MO8n2WC
0cLOQyBy5FX+c74kT33thXjpfOM/djhNBsu3qYVgkv1E/qCB4T2H7wx6ASWQAHql
6ttatKZ1qlZhHUpEFlKgjo1nIVFHZ88q37kWcUmov7vTOQQqGSncH85OKKSbsuCW
TYlvvxN1EUr1sho90UOEfWpYvaaQmiE7uyBD/Un2gXOI3O4spWlg+WZM4GQRbBAi
0NCvOat/vxUwAF3s4qxh5qGvq4/a0dS6xvvZ6eEXaAnW2YouGucdb1s3fP1hdVuX
LYD2orZT2gfwks2av1oyKkfLLIXzMz5m07hYLAVwJYKO7x1C0BIR1As77fYTVa8o
tfoh4bEPc0mDXfIRI49ku7aQY76o8bPhsw289bbyw5CI0nn+y+RHe6+WOoxA8JQj
wq2BZQMiyuZKO+eBwT/OjJ28Xrav6o+VJ/dFfY0NaNkbt7ioVMzYYR18rN6FldZr
PHslA0HlCWGlzHozSuVyAsH9wFkhD1dPH44+Cx1PHBGJ1FvTMp1xh5QN0gkq9TGU
CAxKW5gk63IEtOK24TKlI2V7xzu8EzeB41F5OBPSctw2C16fIsBOYr0AZOJdeAwZ
GeqPqYiSdiY1+xu1uI3LJLw8RqJGr5lIrsMeMXI1kpbxvZLw/UeTC/a4ynAD23Cg
A0Fi+0DqhXGYVZpRToXxPiF08OKak3BQnpKNx67JdJoyzcyXIgrfA9UzA8eAxG4h
zemjACdv42gLyKdutNNByXx0tVifoTHZTUmlelbX0S46qXtHn/Ut8GxsWO88Xmf9
Hh9JwKMKGlmTSBdMYHjv1AJmu2B90GEpLz7Ca+d1WPsKWVL/wx3KL0cvdvt46iS9
gYteNypw9XPxkZCFFnw2WvTno2aulTIm88kGGq9F+sOb3bqgwjirALiA7d0IyM/o
0meD2AvYKteqCTyJb2tMpglWs1iRu5zZy8jRtNBLliMyBLSfMIb1JdHlkPO0Pzdj
IzAr9cyPqSqiRmq9jUDGYKTgBmLKXRtCYU5xl2ytzEfHtCLKLZe4NQ6i4/i59z8b
GRlD0XRku5lR1n+LCQ756J0rjuZXo2vlmeixOKd7jV6KfEzgkhPfNGLtDfG2xY5Y
zKC/b1AT1i0JyIi4QDwTF6qSURn28JigePYj2TM9WM06uqf+f1UsuAZ2lyUC1Rrx
2JcY2SuVYHex5ll4By3ETgt6S1dOV/xwgaYJPuaMMCG+LLuxUkKOiRf++k2oeQK+
aZqaosoWLWNqujul/7Z1AdhUc/Gl2BBgVqG+TLgczMz+SMdra561Oi58zafCstTy
HlGYv2l4fhyHDDmJd0BoJ3Wp/GUBOAxAO6a5Ami56XMDMD6oGt89XPwAbnRRu1AT
51r9eLA6FEjn/x5HV6OPBdd6NEu5htsgjomogXzEosJ/QNj9QNCUbXB76oHmq30z
0OveORainu2TF9THwba0JJHyZ1GfQLGdreAb4mea6YlgAWASQTWtzIXOo9ejj7RR
mRc4CVdJf1Jv0Iy0Rj4JkAXDEj4QyQ5pNsMD23g9SdPNKtjc7YK/WD5U3eSXEt9A
ARcwr5zBtTS+OO46qzE5FWFzBn7OEUSd+22Mh8GodkytL9qWYeSi61VH9RV+NATt
CgtnQk+1SkjGcvncOKOvsjYAcLX58L+IjiP4GULxFP03F3wxUnS6hMXNLuSHb/7y
/VJdatWJidFXkUa3J81lIofy+XqttyiYqmxdsujtuTI6BXWDcqwXt1xfZGoHwCZQ
vrKHuVp0hKWovGLc/AaTO5FD72uN946ZcKJjM7/WW4tUFIWljuZEE7NTs1rrLIpf
bA4f8DZojfvTLuuanTcRSEDIvva5jUbrRqS64UwWdYAAYMWTLquRpPbOvIm4R31J
00CCoxKACXjmyNjVoyjfJQ9xljy/CCnNtQikpAaOkrlBpkW6NwknorUYB0M3iRz/
dSCRBJv7B/v6NPRm1OPUs3esxxRokkyDT4Kof4BRb21yEK4vkZF7SA0pg0wMd6gz
9BklicLnP9GIuTPOo1YKcldW+13TRbXeEThgwiQCnWl6mOzrZh5x9Yd0rjcl2dOO
NNUD/+HAve5hzg/M+p52ANmeGOphILBdfyMYR1xAr/3dlEjKe1jzp0DvQprVfJb9
xhUv8bRjH0o/k75TNLr44XDkp67SOUSdNOkPmDGc8aZqbER3J9Invjscnq/HsY2s
x3HaCCHdP6SGOLOUUOvmXlqNO8pkbNUV3wE3t8Egpmk9c8b0B38YSzccnhzZ4FlJ
G8S+K69IYJRAoq/JU8KO+XPfPE0hDwk6g/bu+QWzD9j/mktSTw3zXYH175GmXg/Z
eMIX4/ETIfrIVtlN607D3p5c3ikrhP3eNkXRRSKSjWtIG2UV3xp2SB5tHwCHoeAd
Y2vqWvzaEJxp05OTPzuo0ZbA2/qW1SkoyDqQNyLimZdjPnrauzcjCb0EQYMOiYSg
jHHnK7yOXvfmuh/4o43Dijndlk1A8UZe6T2FqYP1BWT7+oF/QmpNltGn+3UoW2Yq
WdxaJ/++8nCnOK/wI6kOvSUdyFP+ax844aQ1tjahmN14NTt+Jv7TefWb9DTZJgEI
UoUlB97baYLC+95EalZM1VqTStvomk7sX4NxUvkxQq1ljB82tAMyps7T9GBWDnDi
JkLhmhlSMQ3HLvILgj96DA/kyKvNVMqglKpdaSFUr+DKIUH0vvgtntdt9O/WVg9C
W/ld2C+82n/gXFX5WnMeJ6zaMvevspz4VeoisN3QMZYIE8vo15l7vvtRQRk9Del2
C7PzZMbEMWbTIZsN4lKSkDtFfnVXIz9qGSPxFwVaYloZ1gTvrWWPXxBRmFGl1Kf0
BdVK0ZHpFJiiD0Qbnm6KutT4bm+w4qBsPnxzkj6JRLf67RQxDMQRjULEdNOWkqaE
iJWzm2aqP10vVNPge7FPrWauZ11tZv7m0ciMus8KEmUxeDySVFHYYJ2NnMwUyd2e
ZdlBdjTgQJ0Vks1EsfkjaMRtDnH/5o0nosctERyEQubWwXjoliDEIBtJ7oYecQSc
nYMxDS43OhvyjbAbg4Nq5XGAWwtYY2b0MxMW5h0CPAiCJsEiORw7kC46M4DlrPMm
5fRLBUK85J4E08zGoX+3nTHe7vKyYE4mpcHzIChMJlrFLzSGeiTAIoheesPW4Dan
dNsU6gcNnUT8MtP3guaxv53UQ2PFYet8asypAvUe/IsZN95D4jaolM+W1zIVAtU4
k9WEYvLvRlfh26YWRtd5jwTGpvYc0Q2xAzBDTgsUCrHKDZgLdyfyI4frMR9t3aXj
i6HJFjR7XkiynkiceL0Gw65UXqIMBT6KR3u2fj0soi04hKuIBYZ1AnUBb90cop/X
GAqi0iV+trX5c18HV45BDWpZUlDI7lf89yT1A0ih9lYbfzQm36IkHHd1M6d9cfhN
nmBUzRUL8VK0AghRtHRo9XkYuMUU2j4K3HCg7h2ddozOKWQJ6hWd5w8iKgi7RB39
MWxGQfDnzDrWAOHyPIlFKi6Jr1uQ8LdxvU5Ki57rQ8dqwqGUdcadvxQo1BBRTSaS
Zlpc/z/qnST8xcz5y77DhK4FdsygbBoMetjMCwikU+kQDPmGEWLWIsHOpb4gjK3+
wGxYfXS+b+cmYejvqT9/+v4Kpq2UmclD10JDHAZFwwnNM+UFaSFmpypz16pCpxDB
xBB/mh9bZP6EwqKy1HVhCfrgFbvq7NkVg91mXFGIebSY76RQSNQyglsxyDw+ropv
hrwRP4V1r0VDit0Zq7Lu8lG4+jgkZ1BvHRBYd2z7CYjMIvPzj3o+D0C+YFnHPals
y8GFOymycGWVYKziR6gUDIYmOmYIYuOWnMZU1F/AvgjYUgt4G4Bs6UaaXA+fmvQE
yjDb0mnCRPaGaoW5RsqHIh464qMZvDaWtXN/Fzb8VJp8kiPXviCfytDLvjzekS7+
r/arss0n/SwHqwfagy2Mxulq1vDUWkOV9ee5dBVRzoQAhf/zp4Y+hYYrSAho+dfa
DvtFRJJuu6MM2bq4VAfQ+PsmH5+4l2n3ZEk/KNKDwCGEYBt1G9xOZlPKRZ9XOCtu
csDSjvOy6V4JETLifFs5TPdY+Z9pdTstcy2tvCdIb/XGBSeH0mOU72mRIWkweCtP
zm7ot3Sw+Eqcu/hfs9KwhErqmhtzBAVSJb153sNBbP4YcZlWz1RJa0XR6HnK4PBq
GdnD4Bn3PUvkrmAylYQfvhnJpc0Ov3DmGOrjZbUsvNszCVoldnHIKV9wvacKX6x+
2/j2ASMz5oSru6+4+pzYQN9xZSMS6C+inJSLTUFLRdmpPQ8/RQ/9VgoZuQsJNPAm
oFrE+bpmfE/591fcLL0eAMo27YRyrazx5qwj8CLz7gXJ5XAdCR5n0BpH5WcrRezE
PIZC3LN7s6JvWBL8temzNWNqKbGUJTFbWV76CI2J5gkqXO1k4cjEGaeU2ECvIRfG
RIPNxhN+j1fwZgCeL0ZezGgusnM1R8WxRc0mTSGbWrEVcqryIS3dz6x0Rq3fftRZ
pIyb8wzah6abn8mGz32vIytZIphC6kzoD17qnrkaCQBsRwUdj20sHIkxb0PXIXQP
AsU3PsEGc/l7WvpFoyzhnwkdeCixhxXFRZS/MVydvkGWhrpexqBdM3yGJC3XgJU6
Fz5d8QjERYkVII2YelT0Fk+Dss3DLSZwRRXO9064uemHBNvjTYxszgg03QWMq5LO
AHSenUZNxpCU+amy1VnpLQDhdU/ZInpJHs191ZaIgsqA7sEKaV6S/jHi3TaaQNEL
01KVl+XSr5dvYCLM1NX3utgRihznADrNYdbMBpsG7UUggGreLp0R5n4/Rsu/xLHG
dPr9aHj7Yid7tZ1UUsriaBjQ1fy1aGQ8JHE32147v6+/AuaupogExdFlTwfZrKoO
DlreGjG/YVUWIkGxzp4pb/cX/rjFbnGGDJfvP/CoUhgMWUsmSmH9zNbACEOrwLyS
/sdCIuLz51yOY0Qlkjafv9p9PFgnB77Tui9ov2Jdu7cxhEg7brrLsDoOP+8h8Use
kXdgHXWm4tUOcnc+vl17g467aFdioJMTMX7QZ2laVetNximJDKqWg/1qkcYP/89/
TXLfr4qgMN7UW3X+eoojCC3/TJYPXl4A4uVHxOiq7y6dtx4ttTJC/zbcHaeJ5ZIm
u2s+lrLVTJQzVCjOWvGTYb5Y2oldttsZy98m7dPBnFaP8oJCxXfVJiOuYcsD2Yo+
JTpvFz3Eg5O/ECR9I3CXxfJ20+U+N3TXIUt0c0C6PedvxUyYlQ4qG3s4KQv/aWfh
D1Gpr39VZNXDjQrLgXvd6EyqxRtQppc0wJmyH72MFta2synxxGTvYYPJe9L/xxTr
zJ1m0tV+VnbCDxoe06y30FdwB5QpridKjzzgQeBxkS2XKFRiAoRScPkWCUgqMSQc
GXm1OgATiy0CKdJZANZAXgi+n841kIQ8gXG2VDfGJuXIFMDCDOG9qq87BZoXpocw
YhouBfHjrppfel0QnHH8P/w6AlKf+1Uau7Vxu6jVnpWi5LUtL7g92txeIOW6fSsv
92D+kJOUSh1v02VUG5rkYMWiO00XK7YJkGR1ac9fvJM8Kqiybcyx2HLoWXfgqInv
zNnJjzw8xmPQcdWe/2UrNsnCJQVOXSS8U5kGpIAKEmBFi42DUId2uYSR409IB/ip
L5GRVGlh2CZi0DXpojNTh/77YEHSONOvrXTYoA2otIInvCWB/3uI+wiRr8twPDgT
mLwoyxffu92ccfGVlao9ZYuJ+AKMShoD4GwQJtxG7nypP1brzPbJogHO3MC6V5Jl
x1GSlbzCF7+rZdAfeS44X0uU3N1eabQIuccArz/oTgRugMgp31GAnVALSy/p67iv
eGWKddWtsHuAxvDemImbVE3tcUmP2KEqBqFXMeEEwtZUM4/mIeg1FEfV4kDWSrjh
+/ldUBjdYDlt6TTcXiOFE42eUodWTkFZIPEXMszlerK9YcfQLIdVNK+ziBxAUJFb
JNKvHpuTmwig4VnnnJpk5MAb6LYCMoizVfGcTjqk0tYLWmicSsdXzAqI/P9qNVc8
Yxt5eh+MCl+j9pvvl4WTnuhIgmV+Zzf5zfw+p6OjALtj5y8dQCcJMnfMTzW8Lstq
z+pGAAVL5QDQ+1JZHAoylOXxEdepRCAdQFWckB6aQGmRZvwBv42XbxogNDNQ8B/6
hQlQYWl5BOMp+7W/GhKYIZRzgaBFnR1bxQQajzHmriFJ6O0UyCSPlnNJqL/iTQ5R
KRwoHt9RJoZrEeH+ecNLzaG0QK/hlsdDeKClrOTtd1aUyJF9Ru2vA7uFm5l1yY9c
rmrCI6XtHEBHF0aSw7T6wKo9CrzynQ0Ta2/ajI0xJpHVV5+JptV7/vZdKueI/fjD
l17cCBKwC5j/kIi69wLNMsxc/LFsNi1I/wR63qZHMCQswn7BnPOqjkUGVirQpPlK
KuQC4PLzXBvXXyfpB/wlFAauV3bK1t/C5rj9vNtDEpXkIUDaPQAmv+9HYN+wGWdL
u21tmLQA0LQUstLM1ymVv1Tp+lxLHiBwQPKIpC1DiBIDJMZFzz0R0P1tTVvwHUQh
2Ae3t2vYGB0jBA1BCuYpcEoKHaFJsA77+ZlLG1/m0z47gflG2u/Pgtspsb0foIyp
wP1GYr7HafzUxcTuKmw2kWVQw7vw7hrfj5CHzlC50mANfcnSRxyvyz24r1E59Je7
c7WdFtkE4juKcSrQaHj+RzgpmrnnV4pV469NrYewksSsXor25e955Pj9GgxlYP9w
Bq1tZoVi28PEApfgFakxFlK5zSkaj1TsVIQyqAW+TuEHKZY9LdELah2sXFKh4fvU
KHIJRvTTi7KLGUTDQGZ8cilKfXG9BQZnuV81UveWTsMNzOrgs0MmFzMB1dzcZpW5
/FdqYwH8kp7dUX/Iljqo3q+J3Jc5TyP9tagcLO4ESCmB4/+VnqalHjk3tpqlAUi+
UiJhO5VyJd17KdHqr0OVwduO2AHchzt/pGytEFYSS5XlFevp6PtMMGINASxuxOZs
Z9TNxvLFxLZ6gV4e3o+LZvBQeJESHAcff1Z51nF99GbhRgzGnueMms6ruf7cwAiZ
vfpB6jCaKPemsYGqld3hZ9NOWNGiDTcUYDIWpdiwhJAVnV0PW0i3eFP77H6UpIDj
J4TiQ5YF9H2lWKHZswEYoNc/B5tGCob4kY2e1EPi4gM5ur+yASEkHjye0hKcKwNg
iqqwOBLz5jL4rTXHkJYU3qHH4Gq5O+Mv646JOWNDC72b9UvAcdNwTZ6mjdImo82b
x9FeY5x9kovdlcTlLGCUqxFq0mB7Ix8N+ujkCWCuQrI0lruYmZY+qVRxxtV8PaME
zhctp8O6A5lvugxw7RN4c8UhMPsZTJYZUtzkYNQ/ciX8bREc6DI07yzLa1Au+zVY
OCm1gpLfCk4mDXA3mLJOmjyZRmPXPJ97kNArEW/bziTJpP+Svf/7OC6nQFO1EChl
CPu6UkUixrKhIheVkLAPExKLJg1aRMEauKPVz0H/woF/QXBDoAzJXs8EQsU+AnmZ
OpuMP9N7iEQvPtzNgCG6su3WC2bwy38ae0WSrp1Hx5JqJt1v1a4ML7HOyY0k2/+R
eQrdVga6mv0V1xLXFPEPXxkOxwGeVlrUqXaoeJUY2eoJBlQ75JlGGXjFvjY9FPCb
2B0Drf5cqRBOvXVMr1dsvZA6wWTtGaR0n+TMVe1AvNOcpulT54HYQXghU3Ay7FJj
Xt2Gdva+OiDzy2eQx9admsMlEKn0ql6BBTyR90M1B/qHCo7A/e7u9UUYYY9jJ9k4
iZ7nS6UhPCz4NoJTx+5uxSmLMKgR6/n+CFsD5AN0HQxsR/ioQu7mqAyh6tt4SR1Y
+w9J7f4ET/QszOHYawj02lBG0SZRyr01B6nrEEJgxw1wsaDXJv8w9/MC03i2lIk0
iuCltyd/jhkszGSdcu+k3f1qrvcRlkSGAbXA2k3pLDwXPP0/e7gUvutGNI1QmwrV
QXi0mPHvX4LqhHZQCpUg8McC2jbexFqJEarEqcuzccI/yx6imSSQXB0dgOv/0eIj
axwVUDDPeyjyMyssuiMYVRKZGujnCpaVhplI3sAnDPgnGyOJIiBa/9zbvzOmH44n
zRCTs5hrD3blm47XG+38k7F8zbWnOjotEzMscsBR0xvaIf3HuHUvj3IoyyaXUFXW
84w0PwEzIaTTo0grH4lQLLJTM315+WuOe8FhOWLyZiL99ioDTI+vfnpMJCjlHPl6
ugAvpk1Mpz6ExBtB9fdfkAK8QAKTgedXla5biZ+2zWUZAT1h1ac/FMBGD9qFi1co
84td1NLENKHbsmYdmi6IKYT5IXHlg3dPyB86aObyHC75T4dDHoRvBrWh4ngdDDha
QCSHoC2AAtdJD2K2hSJx5qWgD4Mot6f036sw+uAXbDQd6ODlbg9dNlvxmJkKnAhg
/GcCmuW0bNaLpAXtRhy0sBStiFsNWWGnObaRB79QKu9uvZN4QzyzALFWNZMujGiX
dspGJmTCBveECztKwc8Dmj8kfHAZE8Ak8FnTZx5BDHPaknLXuy4/h2w6MNi7Di27
UU/V8JWpCaiGjPtcyMhS+qWuQ/8dD0BYSmG0x7bGbf2G/9/6rABZhCY6ELImBTF7
Zw07d9Fm/Tg+aOvjPq/vOjqSqIuXHK+wFeoUK4O2tJxjPpIFDBePZ7jEJYeKobHP
7mGgb9TppqB6h73C75pF82cIDDl+Uy9pbC3pEqNA+OenQkOUw/qn5XfcgMN5rP0q
2U88emy8VAKqH05YVf0+iTscdRtDJ8CN8RMV0ZM6bxbhnnA2smbZ2U/CMnmyanoS
Ua3gtJvphYctRzRcVeT0/ZhvUy31Mz7RdUpfm74P1I8VRqDX6rexb7n6unaO5J7f
L/NheUIClxUCQxONGlT/kVlWoOs8yaxP1wnZkyCIk/HnfNq3duT8eYUVIMmcsyD9
Sc0mDGlb0mzilhIzF689jyAXPbYPGPodVzok6pezCa8GoEeRmBUhTeB6UBb+Obkt
/ofIpu4NJw8U1+Ag6VaILoq1k3SbN9AlGsvyxs5SuIOl8Kqi98WrMHSuQkwE4ZEp
Qn/RGD25VQcEi6VNh+9ApfkIfvAJ1h31ipwjzrg1aoUgt86Yfp7Yyl18TMTibJqs
GeOiuezV56xdGiVmNKHRnuHvcRCLSfVvLcWA+W446XYx8US/B+SvwIF9TIF9fZlt
HbPUg53pF8ogC/U4f6iNkeO7nrBe7ss3eo5NzSJYsgCvJ7hS9av3cwf2SQM8+aoC
lOEZUKeJZo6oxRiPBPTPp7NzHcEIhtRVAK6U0FCUpoolRmImVNRRdk3o/s+ZPOT3
lRC9eqzU0xi8DT++jHQj5rHxnrWV5XBetqLdcOLp9L8ZXmaMK8JYsBejgLNlPYWe
vAsdV/ulePVFajaeq3aRJhquOF0a8VvHeMN1AopowFGbyluF6b/xVDx35I3nuJ3K
cxP0uxjYPwMkjgIwO+mTEQm60iwyULVcAHDUQPfcuNXITFxPq3grh9fg11ngd8Ev
NdqiC0yLpf3poBhjZ3U32bjbbemj9R8O3rpSgZfWAi+WQcAwJs0WMs/KuAGzhiPJ
ZgT7CG5ylUkX0kfS63aD+kaHnF1TWkjatmFR43rO28FVOY80luthA7MLedguNAZ7
5jrI9p0wjqgj+isvGSijfiZJHmjGG6qdrEkqUC74CamAEGBZ3+FIhnP6/yXCu4ox
X6mG9via8BmWUTD9dN5UdGrzYNdbWVbxo+bS1F99yVtvy+GwFEj0XPtSXk/aAs39
UJcCUR3j8fwm+sfmjS2u/ShuJ07MzkB002QFbcgzesyh+tU6+dqkx1u+k/A/USu6
4jRYyPkA3XlsWR52K4M3VSo6442g5vL4QuQ3M0XBZjvhRtADhqFZfW9Cs1R2eBuo
kIDUQ+5W/T9e9/W44TNS/KR+HlSm8b7Qn09ygzva92FDGjVJSP0Ns7mBDyQ2pr5F
Wn7BAR5lUHnvRrCytXqlHWhCgkA3vtxxCkMyGwnnbEc4HPjvSCb/1udrlbDzfXal
e5gHvkhVmbFej4ymYyY3pvBFUv1ByBuaVLS2wJtGrHCMfzXJpOnFQhBurC04hEWT
qyiCP0iGV6ttA2lBbXl99x02fwRgSDa/3krNEYDJOoKZeMSGHkbUSzgYp3mXrjOv
CHnYl/Ezd0gUsdKXY5ti5o7Ohgg/fGAFwK/Q2oPGUjXGa6MPXrBysvaBK43bxu8o
zRADFcyv95BNTHrwcawb6Dt0Sa33W1tKW9kT3VwR8m8GgmakXwmRoh3bv8Witxz3
jh83hNxXnXeDTE4qFHOMX7mulodfyjydB9FEmGQrMxZasXfYJb3E5ajwAc6akRHw
AhVksUiJZWCbNRi8SEIAcx+zvpvrqqPfJ2yU2bInhTmu/U2Ov7SDcT+S3Q9ok2mu
7Pch6VUhLr98S3I1NdtsqRakltFtojaeqLj6C3z0FM0eEOFipgSlWmLN3sf+c4js
ir3eaCRLVOi7dz5uPc4hT+oTQdL6jADVFBE4w7JxiH3NOXOfiWYiPgUHEfOSmAyu
aVUcGB4RsELf8RQa3jkwBgYIKMcTn7OLAX77hjmYiKB7n66FG3NA9MA5BqRZtXOw
RTaEgo8+Vw3mEcwxyxPIAQ44LBVwE6wzf315iyDKzEA4rEPhHgnL2Msx4T2y2hi8
Hl6v49T5QvoDBrExKt2chrjkkDkCywqVBVNUsPS7lXrsp3AlmrF0XTVdZ9CjBS+0
JVLhlU9v7qpOfIjl2JoZo0p0O8HUkJrdtsYoDbZspPq5Z+mv5/Lm6iZDp1w3C/vu
j3MkskBcihR/U8Lbc4oeD48H0iWzOAXYmmAJimKzm9OGepIL/uBPSv2C3lQ1ACxQ
oUAsBSQ386GqJNiiyehW8c4JoqpXy1jbygmcxSjRFZROPLK9svUaqTsygP/i63kG
HuT/FwqMbSAxVdBc6vTQUZt4rIvoMLZofe1zE3T7wAxixrkuefY3r3monGfWCG0r
YdRzFWcxwR6k6Byy6TWPsik8a1vwvdE0SdiHp4DO88o9pViaAEiXd5ZSLTjd2yGU
FHPgC4g+eqeu4S/oq8+ojGcwpDqQd22MC9R2mEznxnDIAcYBkFo1GjTxOBQjiLbC
G20I5vqe0sWvx9wCImzbYcdxvWs722CzihbWhMrZYNyVIm8IMVi6SCdNKvazPerp
JCDugHTN6aT/hG8jYk2con/zL92sMfTBqDgrHO4T7xlYTtYVQbYxr7OAzgOYlLhW
AoG1u991UMtVhgO5rfGdJlDywl0ezg0BXk/Cu325nDO2nDmwRju/6Pku3/zM2gae
O3mcfu6xj/ou0hQp6HYnN8Xbb7x3S1V9eW2qj6fVLLRHMgagpxRW8F+Y34m+7XgH
+j3wG5E8Vnz/BiOBKm4b6JhwktqsGq/MgzpMG+Xe4C5R4E3LQDYymPO9TB6SxaLo
s3H2lRfZsx7CjIr9A6Tu+0mZcGdN8yzh511sMYzK5EmtCbd2LRBJzo2+WbeW34f1
PtWbsxMkEju0/CgUM+aMHfcTVgvENqa6dSkreagxg3lEUgJFfz5fz0sFdns2cIG/
nuc5IFqexceSjOnpOyVPT8qzw6ggO0A1kWWx1QvlwXonFensTOlqsT//RCjWd6Zs
gS9kbJlKMKGNgFhUIu82iyWYuy+cIquGaYRdk+ec37ytVAXg47t3JbzkYXe4oYv/
//mbHx4gSs57N08YwjwD6qv9W/rP8umy6dqk4mwNBZU07Bgku8yCsF9U2/77J99e
yXds4FVqqhVzlH0MnZEJyfnHMc+RXggReIfHAxTqz74b0xHMEnECZZcqPCi7Na+S
kz6cX7tW2Ad5p1lkwE71oygLyKWDvpYmX12q6t9uowESue1JVtXae/1OG8FvxirG
HBEtDZvxDH6uGFUeyo8YggtjxG8tYCLq7uk+lYu6ZNHjVzU8Jh0QsM2HE7naeAZQ
dmJWs0XYbVBo1oRZZQyXQmIg3Ewqtz/XlN1MIFCv++mrZdn6BcJQJEh6VSMBJQ7D
LgDtzgaWYx8zl4dWfgfudIKGdwFWgpIPNwNVBgljkJxtm3hkN2w+JIoQPCNv6T1X
JvNS59C2oeTwUp5oZCXpwEPGjBZJ84hj7jJmJXhhb62upTzj5qQ2Ayj4lscapz4I
P90jJ5e6P9MINmGaYEt+zH42qkVGbiJKzkWA38Myn3jRWgOclHoVbvfsGUotwxSN
S4Lipo2KgdK/MhD20J5wn8r+xlWkI0T46WUuzBFxTUJq86JwUMtdlgxgUHHBnf0P
d33clRhDoiS0pEUfBGjTEfeu5ujDIQpDj+nzrafsxe4SOVpPIwxxwsfSvvz9k/zd
kPb7Qutf8FKxhnZSMXNekBcyJvQHtziT0Ljv1goVZkl2/RC5K64aXD59KrKSxxXn
CqWRLyz/NoboF/HRNrQ2mr+44G/MlvVZvq55WRAOBylgrJ4f0iON7TkYoD2mCSf3
AygZNbLuLpfo/mt2bPlafdyBljq4YEKKw60WmGTUOh5jTW/yp5WJMTtn1+nMlXoM
IyGKzCTCoBsHa2zqzD1GL4vJdE2+tzZfPkv4Z3O+Ijug9pONax2aB4YhkBzcsbxN
g3zmuT0zhljf8iuIUDUTsWczDJ162L4WaNVHBK5kohkVSKawUqLY7P38JMVnuRtk
b3HjeIWLfdnaZ48WTEcI0NSD02dBTSdGJB0NzAFd0N8A5wARHBw45foP0C9oq3HY
fq5QHzonaiPhP9OcqoKu3atKzpg8iJbinwzCEhIn+W43lm3Q8oC3bkSs5q4yoyeB
03u2i3x7sggXQpcY8ee6oixyrqpLoeapKWohXu2S+5zY/m8d6il+v7A+in9NzDAP
PtVleth4W3lIW2vMXoInJMSUXtg6PTE0mQAlBGNUEomVBN5GbB3ttm7rDzkHsrWZ
zHP5iFM9+OoCWnKOfBmKGHcQjxVj7w40ZLlEZjbgMAwJmWJDwESQ1oz1pmjYCVsm
GuK++UZspOnZequTjDxEQ6IBlFTWcAWH9kjQDN9lFIo8oSOxgdtaZwNMPfv4rGRc
pB2pFd8BBn3DGdbcFpNjoHjZWxLcSwRbyzCtRWERKNWsH+YEnVqj5DCyoMhOCTC2
B1NDq6nTYhodkh7tbv84S2E5tYLwi02OpDZQmVjdYUIV8d+ItQLJa4kj0l/MMf3B
hY8MYKCc7WXmCcnNFrqndF0OWML1fNwXiN7jzJqV/1Rl4RHjhuLaqWWqLqxGF4Bj
RxvLRMjhO15CoK2LQ9TQbV59OZRnzA+0nL+8jSXCYzt8/QGRfVhyWlCdjJ86tfS4
2ij5SPOlOcnjkiXu46H0YHlA5jHouof5DlnPFMIEKMxfAnt6Sf8XeE5h3zeUcqq1
6N5RxCMOaZZDS1hV6mkAaQEvZw6sut71n8kVKkVXp7yeZ/dR4hTLV6q9sV8b2P6C
ZmTW9wkorF9+XoX8RHIweOM2/qMvIomsiMPUTmIRhLmUdGZ9FtLVjeAX52JSHj6B
y7qyxKW7XGQS9ES+CvHf+dAsDS0LlTVRxKFBFvolLJO9KXwPorcb2F0W/Z+oNCLS
B+14fDYH/pnN5cMmizk+2iB1iiizfchXqJry1/DX+mAqrfHIg3RQRQWZ4RC9zN7q
UOmn+T3YCv3djZ6xOeSsw2zgn0YNAfV3gwMEmcg54ap0f3k94Il0O/21Kegwn72a
Z0T+pUal/GigQBUOpw837tau2EU6ExXZImqL2wnl8iq/8QV92/Of5lKE1uuunjfz
L4Vl+GHxV5auieLf/xifPvxd52mAzbByL3xaMMcQ0m8W9J+XG6PMmPJWdnbmICu1
ix5pxBtarU7wtOQjqzn63omZw38FG+dnCVXxvXo2Opts/r6sDQgTgLFyip3fheVW
TDOAv9cb8ltOZ2F7b9vcGrFVmEeY9xXhacth2hBU+wqOmWysTkcbWuPvbwLC6IzY
5iAcZjlK9EOpio5piwAg8Fky7/3syhWq6ldNoGiiav4A07eFIeOmTZI95Cf148cO
xUE5HiYOwKw9F0nLfBzBeAtMM/xTZP2Ozmxojyu9NOdDyw0V/FKotqnLWhZTsyDy
RqYjjmKbM5XoHw33Aw2AGvcJPPRXW7ts7V2R7LyZHCyPrudaIE6y1GI9n0N9nJfC
/tg48GUBON9ZignA+kjBJPteDXCZ/htU7f4mnLlUqu0aTOrUWkBGxO0cxuls2CkW
yAOH/G6IpxBPyti6BpyAHYTbUcs5sgqKhA/VVir7Ery8sPKpvlXHYyMMeVeVagMU
I4rYMLff+/LiVf2EH8ILYERZe/MbaQf1oNyrHDgATmYnHjlmS6bhV/aicGlNm5jr
7Wu74SNxAMH0TKSnLKp78Xeq3zlAi92N/B78CLrQaulBGw+LOKEi2ZMGGqEQOWbl
48JYZmTqm4eAFarYQjcuJFfgMzRuti2Q8IqZIOfR2qveJZZDpwk81swWPq0cY0Yi
6nKHioZrN1N7FJok9XPIk6yOjYbOqAhHIOYA3182YR61rfz8qn+g8xniS2SbEuV1
zU1wQF5s8g/uOjVrldIIaJwSZPs7SOg+M5INQq7+hLXDw3kmeu37WbYS1U2+cnfI
x5TTrXskHrQZXuXg8VXT7B4dRkhBLu2vxybObSA13uNBTJDuVVUFngDH+pYjerrU
bl9WV+1tV37/cr5884ZesoS9Ne7K3Q+pQcbLRBJQGjY2GUA6mVGUJwLJZtTiS3Iy
5q68tPVqN57nLb05+NdCn+5N6N5bpsyVcuglL0W1wAUAKhjRUH2Dh4+82BlDKHWS
Se6Hr6p2fI1e2IlqWrkCnnhcLv7S0chwAnL0QbUCG0EFyOCAAFkYY+EtQXOVx+zY
NTfiR7G12IBLQUYFSyP3vVvmRzIQbOvfXWs8nXYukRY5CbP7LK1nZqy78bI2z4zC
yTjHZaMuAUuSxrS7I+1UpXqW7STOfEKPpKgSBURrCFpiksai9Od6v7isN517h2yj
U3kLLn03eJZ7axWTZQJ2i0VFVD1lcuOEk5ignZmXautaQ+K0XRGN3w9RUnPIQZvY
BdeZLpOBi3/+VPVSDtcqkB9Kk5VKTA1XGKb0cA51+/8MyrHNsKbt5ynbamQnCFi/
O3X7C7V5B0R/XjKuqB2sHmQY/zIkXuSVqKvjUdWBYiVHHqRIldpNoDDvxjuK5NKS
6cZNOSVxWbRf1YgWpGDEfznKAjSxhdqq+jm2lnwrl/9c2PJHoY6vXzQRMnc9+K3S
jRYEARc5DtuosvXAwhNBuP2Itedc0CY3GJV26VQrzxYy2qqlCuTN5f37jnQw67qn
lV+IDodiLQrhtw9sb+jhpI6yERR0ehsU1y1sSDov8LZovtm9SB3xxO7cZtn8paXK
HiwqQFxzvokJadnJq8OIngG1j1ZtFYsNmmu3c6ihipmY9BFUCWf9PjvMB2d4IyiY
uOWK24oYfz2hWQQhyUkN0S2sDM3F/2BCNtnqCwlr6RaJ99B65IPar+gbeWn9grFV
7WHiX1xc1kLZ1X0yrdnYvCEuWjrUi53JUjhbZXEc9UczxgJsU8sY/q3WdXAoefXi
WNpSYH/xLLQ49Jsq7UbJ+ke66P95sFYMCra6Eqgz8sy4x+2hzgbSIUMHSPCPEKAi
fEO5s+MNtgCI3w6plBnBso90iUSE9C4TOw3+kLh97fNr4od571X7md96IehapzAa
nAMQJPuGkqxRtyXGlh1GZsPJwf5dfF5jl0xRbVmS86rUbGmx9m3GUKgv/dX2++8F
uTOYaa1G1sQpMKsbSeU+Hzq6rr3bmyNQ2Y9hdB88pP0UsWLbAi8kOAgFp7gGII2J
rLPyv0aCz7o+q2zvR+8n7izRjwKCqhddfLqUpL3eaO2O30eGub+idhwA4VdGAx7q
fc1GyTTPkYLzYY249zzF6H3fuOVDCu5i6m4yTj6nbYqEJMwxWeo/DjyU6X+9r+sL
zttUGZgXkbmnZql81PGXMprKOnI9Nt3ylx70kmcGhLYQNm6VpBrVcbJ9xdqJOo3N
7y3QCW+Juq8RMJo/SZgmc7RIVMIPhujHQsn5Fv7u2CK/SIjxH27Sju2XdIXFTDwA
qifanmoXWxBbN6ME5ptPThHenL7HIhnZOm/UeVCxI1m6l5KJ0mhBDy2nzyYld4hH
MPGqRvtX8cvxBt0Barou6/GRkxYNZ6ezt07A4Edf3nCina2o3B0CZVWOWl9y67wz
3qRZMbsKzVYASIkP+LuEJyUxC+7+uju+TgDYKdxD0ooW6donhDq6itYHUHYoWyXn
Z3Xx8NEYvFwKKywLf+T4JT96XTICUxQ654Wwk5JGFPd1UWHxaEY9TXds0JC0C5/h
jtS4KkwmxWjPE7FknZgdwok8vEczihdF3IpQlC2tJCAo5klUklk9RfAIqMSi4Us2
pWJWiTepqqfrYqGtFL48CAzNDT7oT1VoOwTRrdCspXYMNfr7vN+Adq94Ri7UJPLZ
SZMD0yxIL8mBLmUXLBIZZYZ0YoW96q3qla1G6zeU3oqn8qBB60/lq19wxuM5ElDR
eN9oYjo+VQSsl+S1PCDPYC9tyTdtmOnaknzihS35WdZiCE5/dDSPgbBI6GGNUOY8
KBV2mUy1WXCpR+hC5HPv4PRqoaBKypFooXLDZewE2JPyCjUZ9iOLmS2Vk/GTHpIQ
+6EvrOOSg6HoC+EWofbSKfaEi1dHxwai18v0jfJLiP6vl/1Ydlhs/AW+jNGwJC/I
IPemPtm9i5q1NOm7bFvZSGtl84zoSHwJUBcWAH0cy19yipGce98Nh54hKj2dLCIH
teZbdYAogoW3kSHolQ0HZhUeUfHtdC8nv+k5YEQe0u3DIsJOom9qDDZ1zur/bFzH
Bb4Q0LQgdoF1AtgT+emRymIqbqr7KdcvzBuk4IlrlHi6NrW6f2SkFtqyn+WtNzOW
PucuSRM6o1j3cwOlfj0OdiuExrMnbqPg4ddPOuyO8Ry3nVYSaLpPvLeeGD2K6OCm
NQvQyUYoQlKUP59EJOTJ6BqWCKKAW02LrBl7UBfHy87JdyLTsJ3ZRwfTdiXigd5I
hrCjvYpn07FFuppd8W4ME7xvAxzZeQV+7gvANri5DkC5c2ysAJn0OX/yBY5hkThg
zoWcOptVeRHA0TvQxd5+rfXRz7FHOgdtVx/1Gr75TaDvFsq8GH4pLTKn3C4zsY0E
L+3K406Hd0Bg3bp7oZpZ2JCsBX63lpejznLn2CnMBGA77zhHzyNMup19KLwyJ6py
sJNsCScFKQpX1K7QSO9+SgrsKN92q7YUau0bVXt+g10zbOvXEdssvhuJkNxXhcLm
jhsxhkhyLIp1sRHs5ykhaoCNaHtj0YuyY34SQobeO6hYEyBAK+klZN4/ew3HiVE0
9R3ghRhb3auSd50DhKvSUcoxxGisV5hgyaTZsnvDFE7D8gCmjmxE0wWcGOwdoxUe
fUwhiYQRTimFfdBBOk3qMKYwKWpr2ErzhCoySJhDp29l2dMGmqeWYgK7RO+SrcNu
21EwK5P9ADyfwuOLHJ+hYAJmnPJbEkGzKHtAGYLpbLlIR+gaOfY24FTktxNgJLDT
JdYEbm7+qmYvzeU9rICvRdWGk/tVzsDld2I5mmbflGJjxj2st1C0vtWJ3P0vfTxe
U0bdgT0jfNvmRFFrH+Aw6DjCwpbPM1qt0ha/TIcrxHuY5UEwPqm4iWP2VBBVbDns
zBwBVykdgXVGPJgsGmj3Hedci8awXIviFV6AosICy8KQOpWQYxohGIpoM29djKQH
hoEDYrwUmdhp26ctiQgi/pWXqe6zNcIz4fLX8W2Q66OmZj+gP1TXHI88KRa6/Xsi
4wstWRs1XJwvEHBgWwGEXiOVYZSFS5g3pk579h4LnDugyUVurxiNCzjAE1Q9Ttfd
FB8P6oHPHhJ5Jcgrw69FyqW5ziQPVPyyo7xlCsA10Ij2x20yp+OXzd2HCMKlhNI+
JMhAVel/CCgtushy3j+g8QAymWU/EkvoVcnJT9yfyTfXC0yNqr5uTI8WfNJm65S7
Qzxg2CZ8Q/Hc+SyXbJB5c1jxNt7v5g5q36KXg/yG2wBVZv0oMIyk/J0fGnFO+5cV
iwCXgpj2uKlC5TplzkcZL8J0jHHIJiAMjlubSOCp8rIp2sK7JAfkmHq5LDmaRd+a
BXQWkXStRU9+N1del/tQ/kfI0vSeGs8tgGbn30bNCzoBv3+zw+ckoB/gAWv71oYU
xzUvK14vFFPhnBVztDG4h0V+ejXA58e7Dri88TmGr19TnoiNcTb7J4/SAnTr3Ymm
NPr5bPBgWsjfSPgusBFvdtPcBAD4/a6Jwa0iPccqTiHjX49vQo3P+rONzjRQYBsZ
1vzcfWSir1il+9AOfoeYXd4yTfssJqW+2yyVLaVRNttZOoVp6MufBSjEtPqbaimw
`protect END_PROTECTED
