`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oi7ACIgdho1oxfGdaVrfqOYrM5uiW5A2DTcH7XqImEtVe7YBvY3epS/8a33dOsNx
UXEpIsvp00kL+pOu7mX9WCqpc2BFx3sY1I/VJZAOPXJXyW//NNzJenBq3kMglso+
q/AA32cKauiIXL9lY5gCdx6m/slDF8B1kLrSWRWkAJMqmIjEoaOEheE/EqyRvMQK
0fpjE4qXrXdxKKZLl1cMYeAANxrgQb3Cwq83PXsjQyE7kkbUak88U+MbWOEw6+q/
yawBqCyaJ8OFRFnWp/Qifn5aPl44Lrrla+VNGANQ+7/vpFC7wVlM+uDfAMna2VJL
Ll4Si9kGz50Z5mIXmwsLOpyEif9WSKeUv+9QEm7kt8JMVf8FDCO3x9KYen//99Cu
Cr7JVf/2hsrDj1oo/6IYka7P5Z41BOjEfW5iwAI29zKjAGfjUNBj+IfVcjkWqz+i
kxFoo6+Bf21pCkmyDq4rnFdyDxeccPd77jin/PMNoH05FDvjW9WdGKXkIzQHkkLO
J4Jmeiqv93SfjD9FKOt00ySSwpTZfHv2x44VibXyLPRCnJawiMnQXPD5HGdFDedI
egT4rI6Jt0708bDodlf1GgvJ5U3V8Lq/X2FFar3wp06D1PGeOxKa28ZzIE/a/yGd
07ScrEKf1hbyLl6lOlQjhWnJrvuOlTLCuWtrS5L1VBG3Ae+uOOCrXIAmNSaKHKfW
NgChjj7nLL4EiYSWwHz7xx/3Dck67GA+fy0OcJ0BRFi5qnUGQpSHORS7MmJtnE8b
XF6hgr1fcXJL/l2wxejafyX1nyV1TXnCRVcfgokn+SgkLrCPvU/J7nhb9Bl0W8tf
o0f4FjEwgszhDH0gb6kPdQdJUhg7o8tJRMnEeAGka5Pw8InGzzwQC7tiN/wYM0OV
Hu1HOaMZwMAZ73CJ+szDMYASrW5zX4oBAx3W8axuHp3p5FRGkkL0Pt9R37Z/APIx
lHkvdj0sYkE2d9BQs87BojO++JBwya1eXDJhalg+eDDDlIOv3tHeW96mUoOjyYSc
kK0l4u3Ob/Jl8CwMC0Siz4MKa9H0g29zNWodFqVgV7e97XwNJHlGCYMISBoppLn2
z8tjWCAgiFOZS+P0b1d7YPklmaucVjrjpQy5duHihCQGUaPG/gfVLbdmuJOgz2pg
OIb4Ix6IxaMyStB8tQSgbPN41xVHWidReeLeCho47P7MbeGVdatpKdvKc1VFl8uE
rk9Z1e4ZeJliSzk+W8JfPoKW6HhUoQgRSYxMDK1/cVon1lqw9qiDOnolunr0hzlj
e8SK1MxGcmwKgKyG/e45+Yepj131yNMI0jjy92vQ6a5sh8aq1Hftleaf18c87uQQ
SsLlzWu2HYWV3xdCLuyUgSeLtNhxX6IP4N16OVePpTGtklz9kh5wMbvVCtMx9Hh/
qUcesSaS4712Z5XQiUWsTRlFdzYLG3VIqxqFZgl0rXqAUjDP4QR06buB0GKvh0WD
cZ1otNIJTxJ/ROtm4OVjkqWHsDondafeErAgJLIcr9Hmm38HIMgShBex47kIvRxn
ytOc1mATYMFNm98Z2eqRLEF0bTwg1nyEXJfSWmuh+tZDqKDciRQwt6uamObk3jtr
cKtseJq4wzeR4QsmC/NQHGE/F/C7F62nscqXIBs7asmP1qViW4uywPrQxRAgtaQ+
3uQkcR5NcTRH0A0cse3k7tx74gUkkqV/hj3IOn+K5E9tt85scpE4n14JWsah2Y78
AiYTmJRQlGLsLcPKZKw1vB+RPP7io0ue19t6KGDgH+IZAC4dX9D5AtsBwF2nQI6B
sp9UzD8S1IZkakNcs+qpnMbsqAdCeouGroqaLstH9/KUUjeBgytUa7OMouayCn8l
9Lj5+JxXq4c48BUFCPRoqDrCchvsV888RCLJnSljTFdcQIMnFZGybvb3ncLPsoWC
mNOdLt+zQC5KcYTmXOtisb70klMk0tlPcbMv3o1WrQtRPr1431wu9wdJ9+89YN5K
Hjqeo41BKO/yzZAjJFaX9OvHVFOP5VnG6z1BjJ3+aMBgDTqUpspznx9ursA0IcBU
9ms8yM+ujCwgS5E5+4HeL5QoKBRdHC5rNV+o0GLz2G3XnyRA5QNJI+fG42sxgafe
hyYiajIL+jqBC7YWjRr28QcXcbL1gU+NQrFdX+TmKMpQJknVTDYeeM43dqbJBUh/
rO6AIxPQ8yxUT97AB0UldVMVVaEwa8wjBDDbWaHc+IWUmekNRvMUiICKz6AwTLkQ
ZfjAR8gx/8f24HYjKsUyuzLw6s2hhSK5LfYBv/mxTMFl2h3R8mQxQOEa3LxThyMA
6sFRN9IxjhZ6hV/RMA5j6sCktlkXI56lmIglx1NrTtFfYjLeIK1ogdT24e30modh
luiFM2NG0+DAyhibUHFbVPTugHu8ZbGvDdf2Ev4MetVAG3sRUOtcPwLhDjCf/5cg
TPHY/THRmzBhHObG7kzsAJO+KJsqjtMt5UZCmK6klnUvuEVdS80jKoBxYaQKefEP
ynFKoJa1HNZrzO8vW1Y+Rz97yqLOzsvdmRhhcYBDNngpB+KSPFrpTAQeB3/YdIRB
ego8ASJq6QfPs3sjk4SsyPZe45QuY8ZARSgTu0z2KtFI6pYTCzsENwgwXrvRJknA
n1znHKIPLmEPWN48fC6Es9DdGWkoF27Fdb29kTn5acA4DZGwtW1ptmBgCXQebOgd
JxYABgMyA8O91z3UCt4UMpNX1Dg9I60WEBkIcCMyTCZS3uZkVPnewYAGgEcezfuu
vo8lxTUrejnRMyvb2e3cIA4KI/bJ1faisTUXPWLwBipEcng8gJBtyQcwIJPJZb7r
s4uVmS0Vk/SScJrS27w1/OPsGHOEHbf5bfHc+dIjWF2mcCyRqmgptfTYbT2VDBDe
`protect END_PROTECTED
