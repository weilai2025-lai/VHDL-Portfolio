`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OuN02ItoT7By9KUK/s/SbRX+3fso4DDBnIxqV8cI4B7oHRWRzhYdfzFXqSUamxLj
53Juk5tu2oWIIS524JTSBWxFvBpNuSwdFSHb7+SsPgtOJppThSP41VszbnjFhme3
4iupJI1n+fUyi8/bOrmICEHIY/7m4iRs43lGZkkQR/SWwVSQBtvmvm9o14gg1tve
TC1qIAbDWL77nz0KYJfPpnkPA1a13NEJyZb2SxZkf/UlvtLudjjiVvfdQqO6yiKd
X5UIQSEL/Z6Dj24RN0SqKCDtuzbuzpqvmtC/yA7hlYGEqWkLAv0h0W3Ur43syDCp
1qY9RKdrZJP1/BV1hoMFuH3/yY8BrFT0oK1Nla49uoFsEAyMADy76++m10EwdxOx
nl0pU3gArjRl/m0YkglTlyuBIeP/UeEDHdRnaD7GqYg3LPI/4qRr3ZaHF+6pTp2p
E31VvGSQxDWx7so3h5PcHK6EkBcrKi+DkOZ79qwKKrgZQiwg0O/JKT2XUTuzwu+u
AhlhmQUBmTbPVP0McAponhcZU/3ZG9KBaQIFMLht+dezrrkqXsfP26MVjwAgGLOo
r2WAoTIA/QKOIljLiGNcQEM5RIr+R0JORmaOS/qspVYTTfsvnjBdDD5BnJaWGNJu
QAV4iHknCnCPIDmd9toRvok2wYL1P5nqJ9cjbbBL10XE6roCVtyF173cZtofW0Zj
8E3cxxJy2yY0SwPpN/d4BccxD3TAMHz5IeOMKIFl2I4xEUrFM9cCjMM5FXfSTpYs
I1bTEHyk8lS+6S72LuaeIJ//ymH8q3sr3CGHH8VtGnVv3ZMjWbX5ZkgU1wboJPqW
f/uwUQtZUFMEh19bDgCS/lwLRrEy5YnjN+yBXpoJjPIOFV1XKKobEwFBveTJQ7k6
Nxw29UYnvxHQzFUgn544sovXvlzWSa4s6/I+u0/XoT8PCn49A/okgPeDfla+GzOV
6rqS3dcfod5Drb+FSkPB2Ds6xhUKJ5PeIdZSZB6d8OgFR7sxgJFnmqZfOCkQHOia
8xwev2Y4zZ1hOfsL5BnWKgC5mVvWgZ+FcSsZeZ4iwhj1fFlRb71MTGej3Y6pRPLH
D241W/g4aoqfccvTr0Iuq7ahQCk14zDnm8fmf7BhtvcWS5dwsn2N0sxEglNnrEGY
mhob9xSqKH6PCwDyd7tNk0WrjjoVWxpy5fJVH9v78yYUyP8Dc0SCQLM3dAomxdBy
rjbHSXEY6MCrz45Vu2vpOd0w4bU5AmxoCweTf4jxrI2uXupWMX0QdhxJQbpBS7II
PTziL734OuEazR4UrH6gGJZjLNJrZ0UH+whbv/05lwwe0dgEuXX/7BMXp/MZrH+z
PwMj64qMVvi6twHXFf2Xg5NPMK/QAocOjtaVhTov3aOaNMwGZvFqtHTy5ep7HiIn
IGEUl+1BmsPCiPxbdSeNO5HKVNZ7U95FvaH6PQMLU5kUJyT7leIQ+ey34tWnZaWh
6tZUFUdFhjFmFVRJQPzHYqXSwfijWkwjEtoFtCOTJIBwxTx+vfd73d4bU3cRVd+3
fqcxDThrlTxXrL2MQ2rWpJYZMJYOhAZC/V5QKkDvomwqSgVDiCEJuHmUcDNslERF
mVNFmGuSf1OwiPsuainQ3nh/nQ7vqxFX52zBFl+yhyFTzp/Z32FweJZ+ndWu/xAT
XaczPnZS0QGpRC5mWGxwRmM9MbdBWPkGtSHlbQ+c4Jx8Zyooq8JPERb1/rChTT6C
JGkgdnyjtzGBd6WUOHsR7gGR0CUPdv/Vo04I+vNB5+BcFwSLAnOsS+FbGats88Tc
GEKj9ea+LauJTxsd+QUZoVmvn2VBFGBLnzneTYY2jH0a+3HyuHfmoAU67txkjd1x
G+FkvttVaDv6ItNd45FNUA==
`protect END_PROTECTED
