`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZ33FnqsaJ7oedTkSReYNuQEqq3OiJ3IIHHeWmDqmG8dug5eo9eAiL1r72O7SIAe
mRuaU2CzUAvs8RVpIs+vwOJ0Q8YDGtB9lU5zXNA7XZrVcLvO9ocz3w06xQaxk76r
xKapebLAfs4SrVV4axGPB+NXuywl549jcm9TKjSVy4Kpnu/bEoRPihF4B5yHGhwR
YtLqdp26hI9o0a6IPsoJ7N55wkZUE12CugykZh3VpqaK/W/2v2h/UhUs4Iifo5E7
02jOGqgHSII5sSYhFoFLdD0JGfapRLHLT5NCigrp7JvQjgjvjus2zDD4INCInGvY
fWcKxoMmS31kG3AeJnI2w2TMyVD51t2aAEOldWjvEhZRSJvzAM7IQXKZ4pbmKfAE
t90NUC8he7y5Na7dVwo6gO8yZoBKzixTCS3KDu7P5ZtbQ3eMhXUNMm5kQZgjpuer
h7sxAOwHyAka+B3oKBDqwhtXFM7uzM6t9mSdyXzbVuTqDWwdJKCUHRP4Mkbnemhb
X8q//W+NPYLyQm/1pvncz8MWA9/tVH+C6LIdbnYyK4lNPkTYhixD0FdVtNXKq0IZ
Xesz9NgNs9iwcy6fmGBqzudZqfU2w3aKO50GePzI2jgDq61prn7IyvRe6GVjWr8R
cE4fNGEDI2/JjJIq1eUah0u+P/1KXqiOStb2I7lAsHdgDBMYIDviYgxKjt8UcQqD
`protect END_PROTECTED
