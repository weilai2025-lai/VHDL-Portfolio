`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Yj7/vE/aZKgFDnuwaNXOw14r0cXULiBYuGmjkUEPAD0wr9zzcWYx4exszPW84Ak
/J85CaN0MpbGTJvUihy3jEJzXKXaYTps8yILWIO+LOUsMlx3jzZI2KBhrnQMw/7V
m+7M35fIezZwrN0L293w3dazuQPOaYiS4JNH225gWESt1xTZNMVjA/urTzlPv2/a
IyZoEBPb16KOxvSOjcJAlb3j4FYqv5Ooiv99tNMOJJy9bhjeiiCTJpgGDeUMLqQH
jtUFlum5TkrErofJt6kvdybDF68CxU3KUiP5/XKY15bWR7lsDmvSlxPsj4cR4cfH
+2SzzJ8YH6S2R2W0s47VZtX2h5y/hQBMAcrwqgUJC51rjB5qyXs2u9vs0I7+HkiB
8pnqDTuUjmjfIuiXjthchB33V5sj3TwPpCI79D2arXGlpVfDyuiBzLEYBjyHkbPV
p+gq4KPfoywn2G3/Jw0eYstVJPKhcplHjqGx7pt+2h0MeYRT5q1xpmVZxylbLJa6
F5Oei163T3OceQc4wPywG8S1WXQpKPN6Ss1tEWKgGmKG95SxtSmut/OxAQymprB3
4RsZO1gOWRyPgLBlg+xd/KbVtUS3aeoukJpi3zz6dQQrk30dNT0rrpoczeaAKeiY
HTIXZ1gHZRRbeWkMQELFMCfyLJSvbzrCifiDPfw4ERIIYZf0A1t4BrWsckuuZpyu
ywgYCKpSgwA160T8DRQte+IEWo2ZZmWXtGOtbA1euDHs12IrehHQ7YA89crUuZtD
TCaeT89koX5A71l5GazBE9hNE+tDHO+q5HxHZK++pnGA8W0D0YH9BaEiidOhCNqY
2xLP3k8RaGO/BAFsqD6v04/XtskoI2pGc2aWmP7Hyx0e7+TIvAOnNylp92+TdzMo
rs0+3uSsS8E9BOd23qlKk6yv8k8HXR8I6U/nhuH2yyri/y+ZaodLQ6NmpSS5R9+2
cLYOVsI6dFlt/mzE6I+pGjngg0IzxDyLjIegkbhVQo2hfSP5YdeDU7y0xkvePCU/
CGptPqjrn8rwuf0IyeCg7ELOtvn+4H0PAE7H/8WY+wj7TFI7gSXl+8wPaClrMJ9I
DjE5BmYA6Cfq892yti3ZbQXewROIK4CGMvtI2KOB3fmxgNpV49gnzEUrXE/Vr6nS
eZ6c3Y8PXTLIDtjJr4BKSUY4gWwHo5JYmWTgj7ibdQ8S+VDExvpMasJTl9VwtPj0
lhxA0QE6m1RgHLyZLpJJ13Ex0rAf9Nm2dE4rk1UGvQ3adJ8Jes7rQ/OAfByXxp+N
wlq6YHqy5/FsFRd41/6BAxY/RL7T1j6M8jlJ2eYpQF6wkpSrf7gd3t8gU4YGd7bF
Ql60Mn8LvG9EQX2MtFKdjOS6vVPZ9Pi5vczyC/FtkzMZYeXOgGs64jFtsRR1I22Y
zW+Rul77Xcey6SP29o7euE9+Htd3SdwuUxDakq4Gv3dDDZh/tVYipZSSEn/8FHNP
bcReLGgJyG8Exls0J9cWCF+cJHeMC5XL6YFIpQ879FajoUtIGpwaPe3aoFFIfMq4
K1R1p5FfmzpiWDM5gGskx/HycG8WtWwixH2l68vntRRWjahTKIxWLlovRgMzHpd2
8OJhPh8uriSDAsr8Ki20ctD66afDU5pKIB6jhNNUqUg/+2HCDlZadqYDyDCnntMb
LBacoJYcF8oCjPLKsXikNw==
`protect END_PROTECTED
