`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/WFb0JECsPDAtKwX3tzhDDFUCN5mpz3SM7Dt2BJIjveFlI5I+TWABAI/4/OKfea
x/8AJe2kqdOQ8MQ0qFYcaB+gcjz3OqunhIj044URecLOYZ03zpLj+IFHnOmaA0vK
6ra20P5fTfsXUO04yC0My2MWkb/nm0+CrsMBpU5suD46OQzoJQuOrqNFQGwpEYcx
cGdxmESmkYIHkbG+pa18hRdDwFYUnAbOHZcGan48SrRNZRSuYNOzU5VnM9+PeZRD
KhzPzDdof3iaN4rC5MQcV1Pn27+oyVdtI4gFGOkHmFetGOEmf5KfrKFrL8WFl42n
d53eKaFNDX6XiI+2PJ/CHzBgNlcrJUlCHAvZ+d+DyaLqb+2oTLKo8xBv162NMdmw
gkAp2m0q0e0xBm5yveH1Pmk2gv8OwW3AAYNneTVolUWpbfTLHkceBi8K1ySE6dku
BpW3g5ASNLje5p6UomJ/dwDTOJjqgC5zAbg0wAdvLkDgTBYwnEBHI5WCc7sKeQ6B
rVdnpwnHICLtoTNngYvJx0E44uAem8sRidy74Xk/CfNqdcKtE62GnU1TZ6IWwQ2O
w51yZht1hZVW7Aoum76Gl8Ca7Zjlk9NOrH3BzvIHpYeAsQ1Ry/IGA0NglaAbQCxK
syw6xu5G9swHZ8UVxobpMp8lShU1jphQtD+Cp43oPddQxhnp6tX0Pr8tVhoo4GBY
blUTnYjux2apjzaYoc54LNfLqIYvnnGXV+ZpN63VjT/6jp7+0jNsUK+FTaDWIZuo
gXUyema8TP+sU7vqxM3lnqrc/mlchQZFxIA2nS4AyLePNAUROnkYh8PDa49wCZq8
S2Bs0ws2VSqKHNGks0+3xCNmKgDhuw9xRLo2A0b8qX0FMdMluYUMyYc9NxD4JR+T
0uZd4PDlOpqCE/57Fg3evBLPnxMtY1exzHMUL0f1zYiU5eDTkApqFNv5cH8LQuwV
BEqu6lGMU8YJi6Dk4EgTusHBX46SEXHKx1PKBOCK6HkH4xCS4kdND80+5ALPCiUd
/IbhXnYRID62FQ5REMKhxh6TVE+RK5+I4dp+eYP/t2xKo/3PqxMr5jep3ga/fwVN
WP7aF8JbYjdMeKwc290WlutA93iBbra3gPxACAVvmPBhyT9bspRJ7ltqtkPH+8lR
Ci6V5yFFDEEfZFnEHk9lNZw42lLWdrt5jB5U6qTG2HlsdlUmFd7IY89JeT2sP8fI
resSQ6Ze9i7NQMRYdkQ4A0l3ooWgCvFkh/DdjFEqoCuGDIF+N1Y8lvl5HR/592ft
`protect END_PROTECTED
