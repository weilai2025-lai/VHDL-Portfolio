`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dBHUGXFmAF/rMvw60KazTya/xoClFAesDju4X/8tUQxcsNYpkI1NR/kDXEv5hYM
Yn+xrmSzLZu2nj5/u3lPA0831Vwn3HtGHoK9SzYYTs4wlt60H5hu74Qjbii7mPEX
Sbj9iS4Hlhl7b1Rw4grfKZDzPqZ3RkQMSXeN9KC/UcDJIoskRamGPFM3YVSoQLSR
kfZRxic3dQNcfpRmGhKU17BPuSfl/qqlmxeLhmnDzxLua44Fq/c4eoSZG4raYy+d
UU9B2SZuSIIaW0XkrckESsHMuoetB5nzA6Ybwh6GTweTxPfa23D+VqbDx9ux1bdH
9wsH2gEUmkeXgkdFmkVnhmZUW6I2zzMVRQq8x3yZKdz6GnjnSt4XlTImiBoGzQ+p
Kgi7YaQoc0vpMbte4xYZPff9P66bRp3F/LKI29h+3yPfLkOaEXr1zKnIgYYwdDH0
VfyKonV6EOW30z96XtkQSoKj1OIw+J+vmhrYmwsuwIdnwpqQ3tlmOzCvcV3H2Ncw
B0yl/pfpryLKpmaerf3/cxeha5DezegWBmCRzjvAF/P/c/OxpK31MtGRnbb/14zg
2c5JidTGvsnEuP/G6bePuUSaJS6fwbWg+9p0/PslwMwMifyeuEOLjdch42Qqjom3
sl2Zl8ZSUZhmO9RMbStig6WxKl6cVGyo9WA2yVxI3kkJZ5EkpXcZF3a6iqEPMAd8
oGx6lrRkIVw2rY7TqOKDUd14ftr0h4+65mAG3fEgQWm9LY/k5HmK1s2cEqT5l9i5
HcNcN/s9Pg9geWB4FRGwhIugjXsINS38xf392VL9VwWyxtUVqBB2UuzCQD2min+Q
JUqOdyDv/e4qMDUxXjqj+OyJbyKCZa5lVyQYHlDoKVsdvqeuZW2rH+IRecE+eDi9
um6iJYcoj/p/1V2zOx5/Uj9yPsLN3Ck9Hu9vw4P5+cdLbknxfX5ZZFa/ctwPY8Y4
qNruSX22TuoF/j2n6aZZ2DDksRKBqL2CkvolyzIrb04fYBPz97aYQ1E4OdAIn10s
fkN3T0vBNSZ5ZFcKlPJ6k20ZHS+cMH8Tr1x3xzVoJcM1BxJ0E1+ZWtJbwg/lePoi
QmBLvL40oKVoa9ASV3khb9nPxDtIloJcryXcdZL/JizJtL+CWz53XOOhesRZL3vG
jhTSw/r1SDPDa0tQ4cSb3c6bNODy1VVJ3uaXy9Zr0SrpgadzLoPecEU3Z1LbHVw3
VUaCGFjpAcfJ6RCEc/tsTg95ZqfhnX1NjZs0RbwRn3bfMHOZSYtHamHH9tsyH1ko
MzT1+PbKD0Rh92xLAu7DfU4TEJoZwZ+182YX1f3/vxbxKqfaNtjwohcQKZwLE5QZ
PBkSDIH/85/LeyMQOVQKaQR1llciLugENZAh2NMLcvCOf6GDf9SuYiboPt/LZIvr
8W4wmGGt1xMKauUTIjk4QyNRgnFujncIkRg+HbqDPbrcAybg+Osteyw+gTTRii4o
qPIUgAuBy/4c1UApzPcNgmGL5MtPqgyAyJiSBjsY3eebdH0DNDPac3n+PV7d7NHe
bQ7lOpsPtTtGOio/X6OJuoyCGaazJTL27KBXGS1MVK0AKLCK0LdcC1A1Yjt1y2A5
Nvux2WDmoQSvRso1TiRXGok3mjfWtIlTG09fx/6Ozr1XkO7LLDY1ldkb6CkvM9Ox
pFLRmPT989mJiEMY2Nwm6nNQix6y3wD1nE1bAIKFJPYRj1IHk9XXFpMKI8Ok53Ql
a4f+hCyqE4ScOugqGdV6Nz0QWr8VRQohFnGDoq/xUYAHHDJSYm50AB9Q7c0kwxBt
hVdMNNaybVfjC18qD8XGFrcRUa+80esQ7NO7KkgDT54puuFUotyrhRbiZR41wglh
4mGLtXDofo06E30GfO1TT0rS2d0p421f/PS/paIdvE8g34NeT0WTJReecDy46X10
jmfd3f/T4L6mfEKNFULlGH9E0pzmBxf+PoorbWwf1OJyFT7xHO9NE4i5sn4480KU
8MXkZh0RqSVlvUNdNhvf87fI0rmvbd8E76BpdCt7fmSrnI/xuudfVLXn1Tb/4Jjz
wpxWot8OPbigiB+VdjmIPTt7ujJErzJ4K89Z8EnywRYEN0LHHx5dmeypLlc9Y8A1
oiSZt7ukGjRprWMCiAumHPaOZsGVkTueArzMDXtyAiywVHKvv45zplcp5m8IZhTI
LaBBjc3mzV36yPPYQA4zEtAL6e2Dr7P1/5EzkaxlKZc13sd3qrxTDrzBIlDdkUXZ
8AZrOYH2ZLx4WB7iu4C4EapBG1r1njOKalI7XiPbFr3AGdds6I8s7VnqgQDL+0cg
PC1ktkTaKXgkh6IMtiQ/8hTrSGMQ01MdhPQe5KDFQz+mmAcz7m5yJfqR7TZy2y5O
M7b7uNZu74VZZgfkKz4FDKt+fIpppPm7Egvyv9QGChUN8j7EKnWOB4hpLNllQZzd
BxIERX3n9ZOxPnjXNw896oNyTE93V8rSe1Wtsc/P0FZAYcp2jogKgOfxNjd0DMMz
qS2RdrTTYCyi80RKBxG6RNksZAQHrzycfZNvysBsUa/MeB8XzMvstU0rrHlgW3Z5
Kb+1JLLr4lTXdhNCWTZNtFGfkGcB62tJb9CSQyuNea1HKxrjL+JE4PwMKxtCGl4D
VFhjJ4dV+w2L05E+9V3TM6Q62EINzTMfZuFU1uhmxUrz/hzQTSvnjViWtID9802O
jdXoVbpZLLviSVF0sNJpyMEh9pxzqI9Hd9y5MgU1VOK1tmVo2oK49i3O1nCDGSrq
1ma6FGUd+eh+SxeGJpkbnnuDVGdoF5CKLVdrfiXzR5BgoHe8sTW0zQFOFn9v0kVp
BGU6OteNOZ7AU0dnZZIivcSVg+8LueAqYNKFUSwW9kIMsqUv2UOzPsECYmCYkXLC
K0qVEtaVAGifoD9qsIv+Fkog+tBQJA9d0GnVkotz7Gaerph68H/w/gFJu823+HxH
e7MHu+vE9ySrhePIDwqg2mT2coIQQx8ANKc6QFbNTMAJLjb2IavXFEQ0NQ49TCcK
1bb5oDew/XVO1lTt4mV3le7C0mmgejxn/t0vd98NTCLsGYVVxsRJ5XUea1wX1Vg1
pn/2313tRIjGVYcGcAI9t7zOZK10C73nyLsFx3PBd4x0BS5MNspxIEVmq1odS7E1
vS5hXiPDoPvXU996maRKQNAMsDrZ/1UW3AXIcMZIupaJYNRtqdqJkIk0UL4SxZEH
D72wWCrz0Z3tjKnhAOqlRl3G36UaPqLpuahM5jw9/4f4fKfm1o2jQxR2m3L24FPv
lGzz99HJ1pCYpVcv4JB1tvnuU9KrSMRk0/CM0rJJYoeTLm/IrFMgVhNMQrhuXf0I
XwYjRzVPGncU5u55xDnq0gXJdu6YBE4SC2R8+MqIi0i7Zkj2CFXYeM3H1M8pxxCV
VgsTD5fja7W9QHLwrW1c+OC39Bgk4ainCl8XSHpyTdTTD4AA5km7IJvPgRrO24se
zp0Fi9dL02WbiSIsYEKTFS6Ef1DE6LiP5w/c+lc4dUmOG8vbHrZk6h37jTfrIwnC
AsDT2EvkgCfA6MTE0MKWyUdNLXdeHcEpyRjGQXGR/Eb/rk9rDeCmI+2uuqSZtn7b
WNO7ODB5wLfr4Uz1Ac2cf7crtNSY7+2cwgdUEoU8K8HQOe/u/3ews93vgUqg+0Dp
ATKfFdo0I8nxFH8MDhdkxskoVaCPU8LBPBuLOIkeIGqAZSOAHBZ5lv16Xz+lC4JJ
ffTaAV2PjDpUGNg8oV+u4eqg3sxWmRnGko/PyAkU+6ydyeTelYsGWuAmx345mGoQ
a4ksuMd37pmy8Gd360jdz0txCkISXakHoj4OhGwLlAI9sryn3z7hAAkUwHEgeC5X
PVPvBQkzQXVWTPTOaSg/HQ1QzjROsxmttqFHt8jgDdPNoG+87m7D6vU/Guogmsr8
QYM4EeWVaNEwd3SuXqd615qzoasbbwHEao7O+h+7xAUMHr3H9eMkZCV+vh//7RbN
zHn3vo0BCS8u/qZHzN3dMNKzz9osN1e9rgTKIxNQD/a628/l6qy4p0OowZZ6+j+h
rQDjS7CfUIq+zo7ffOGvq/KIKIZ2tjwF2Q7z+nf/DcYxIhsexLhXprVlIXb38BCy
BQXjt73/IqTkLBC/mRJMy2CJcjrF55Dq5BSkPOkfUr3f6+MJ/miWcv1FUKIribht
zPo7YsfZFZmGeIP2Vzq2aO/BuuT/pt/KvDm4wR7KuvMSILWNv03BTklaSgdElF3X
I5aaCNBY9/yY9oVSmfpUOC3eaF9V/yhVLu76KIxmCdCRtm2mgL2QhODbMgS9K1ov
8Lv81FxSc3MZPrqKeb0wZHyb8J/6ccRZfeA2dZYgOxYrEKizsyysFCqdz9UkEDiq
vVxGDj4EXb4HnKvpGzQyDT1kYjfWfnlMY9q2G6uOpw6sS1/rDv+UZsMcyzmSXBNO
S8m6jd4PCyB4bBv7F9fdW3704KKmjQYrgqaaWbKVNgTMUoM58vWNX+LmHF+wIOAR
j1GiB6+pbWuyRB1D4hL6gCfuzyOnE9MdE7WVotHwkNc5VONAORFBCmlVBOni4wMH
5fiCUEwK9pAzCI5GSYFOlb8hvQfPthLWDyEz+jaw/dDe41L+8d5V64h5tTJPq+E3
mlq5cxTiERp9nzpb38pxHbjVSht6tqSWnqQeodaHOYIID0TxO0PUR1TwXugKVIb+
OrDvdyxd8iPwktw6Q3nqiGlWIYCrxu8rAgIwuOLlrZdqv4Y0iHTblDYOcZNRNLbV
OtUHMfcBM8lkYhavwzzzj19cLjrn6fn3zMkr27gIGZaH3pHOEjpzvRMmaiDabDpM
6eqX+a9qL3fwnpAGfn+FnhMPX4sV4zNB2FW738D+aQoinDTtlyDo6HuEi6ICFp7Q
ydrNoeMAhJ2p1aromfw3NhXUiF8S21gSkKPKE+Yr4XKQvpAMg34obXjiQknCzYbF
50l9mkGsKmoiIt3CA9mT5+elsq9A4QvpYR8Utx4hljTbcfd37f1J/WqCTsAAogIU
v+74YZ5J9UsC34YV4H0fyHipZt2Gu4UNodtDLNFBFlvGt0LFf40iWmLKkY/f5We4
ESYXHEfqH0Jk1XxsjXloEfIxhzAKwo3nSN637Jlz0NECwSNiNreZrLuj2JTTKDNL
tI0GMPMb22kFU6uWz+FNaihBymlVzDe+3saQZ/JpNtLpdS+qIcVnHoan7v0Lf0Il
o4U4TXjSZlqh70fjOud1O87biAkvm2qMg0w9PhY5y0Lh/wK+Mq44PxFwzKfO6cy/
ju4h3Sd4TiWNvbfQGUXSwrioZ6ydt1p3oFHnRx3YtzvXip4ZVgYeC2BNlcs7PuXX
sFrPLvBcwquwSjRRMIRvraXnm9XNvBG6T5LIcjb1WLwbJA0ri+aB0IW+92M5UqPY
X1f8yc9EsGEPojbHn3dWZESDzdEitsW/ulq1MToZKskE0YUUOIfsiZDNzzkefar1
jR2/04+suMc0gje3vngy4O0LeDTu+wJkKjLpMpnwtRDh/gWtIxwKWZJFa6rRf2ZB
gX2qtJbuv50ZglGxFvswY5bdYT3jh6ENtsL1L+pNnA6cdDGVGJpR/2ac40P1damI
UFPXTVXTJKAVPnJZqsjVLyAO+UftlqX4rfjKYDNktDK/qmozcWrFmmIBrC33dpI2
oXx81MDVogeC3diMjpxqn0sNQEpQ4cfsgJ2aHV/YkAzp/HcUkxmovOYWctLRBaX2
PwlJopjJ9oWlqtKz1hznvy6Aq4U0eG6A3OV+U1/Ha+vizdqxRdkVevApEboWk5pT
WY3Ae6om0pYOcxExhfpygPjg++Y4eh39rSLjp+4NKk/D6OkxLSn8OgyMpc/alewk
5CBjwQ80rW+GXWwjOn4eltLISOVp1Zae9RPlHxlPz2p0fQ3fVDB3/31dNz9ECN4D
GyqUkpJmMlZN4f3+JpTL7Xf/PApBRij08e0zkF8YjEcT0yD/wuqL984vAuTjGpOs
/7jVLEHQm6WLBdKUTg8kwrz8PnRxTai5Ze4mFCvBE+C4ovLNTiCDHHbwbw0r1RE9
jvDMIfcjqDmqW8IREZQQslmqMyGUPOUOVmyMoNCpiNaZYnv4KWE36a8VqQGglk3b
3Ks+TbeRF2lM+O5yzpQDAYiBKYHCwecCr7n55PRHaiSnHLBp1wdfpwWEdxC6DYqM
aB+J6Q5Ib1u+ruohu9L828Detv9ji7MhqyObCAisWL26v8w++BUNoUTp8jkRWHWb
+qbvAgvBB7JK5g2AYnamMNd7hvDfgA7d/XXzZo+DzW/GX7Mitz+K3shYC2w8Ms1r
3/wZ8DdQKfvq2pA07i0mw1rvs9uAEMuPA9sXL9yEvgZU0jpitfOAXSj/IPyh1bWC
I/EpJrPafAaWYAOqy1EXxYfYi428AK20jyIiCxC84gIVt4pB1XkaoQbgqQrsrR3K
j61+m2T38006jna+S/ZB/sNY/BbiWKOqjvlhBdHklnBzF46+p3MYgojo+Mkq6vyR
N11bxZRez33O3TpH6T4UOL78CQMpworG0cDkaSf6YfARZXGDEGSJ7AMGDrF1E7Pa
skmAODEhlSrTicvpa0LQfoF10uQltIMI4SsxUHb909TwaqXpqVWN/o/kfC2XY16u
W+qlsnIig31eHkvt1KscZ94T6M8HAPKdmhYWIbBoAR6IiSqXRVScqrFK8+vW36yp
udHWgrc3JBDHa6uEJJ2YZ7RLw7UPgW00oc1MO5NnjnSqa6TsI8t8ODv5YJWNwWC/
sz0gUDZEBXTrbtlQl1irnZqhCRAMzENrIdQpCEu6dDNyLyEjSc/AjlvGnkhoK70d
jeDT75VeSw+fK9dGVjrYPVyYInGIAXO2q+ZUbv/Iagc5FrPLu4fvR94Fd0iQxYkI
99M9UpeFnWcOzLS4JcJGLfQpT6+h8bq+XkOhT+VlzDfptau+gdFSo1uTzRikMQQo
RNnTuvqBQGVt4o1gJey9sTJqvvPqiW7JtTFxzYaY6nGG+gz4QkxEhXWgDlse8bgZ
MsmzBsAS3NXQJgity781Fh1Rv/5itM6+N53o21vByP8g+ha0AVVcUGdPvEKSvRaB
S1PtMz/0nFXLYlwECf6e8vAB5LoPsqBU098rnVvNkLEdZeY7Kl7El3BSAWbPgVTR
o8uiJVKAytwRuhQEe2pH8DG09ZL3/b/sAcAyObgkoXZBYCKmmuMdY5tCtC7Wpo0j
SJjzWJG/Klh+Y+LYa0WD8RmW9imyPojUF+R3RoodaR0TnkF3JBi+oUOY8JD3W+5R
m3pCRCQ4KYMM8Zt1JSHqctM3bQGPmbf/qqNfvBliPGLMxHUR5nNH/4XCLwnvWEji
1GOFCVPIojqiiloCxNN3baa82qIS/b9vlTyXGpzuZ4e9J/fStC4sU8FXCWlUL24u
berhpSu1yp09pupDxQbVL1nxlRcFAJDyMWQONymVlho4AdXekDsmctFqSJ2udYyU
vFMgFVwP3EvoWlV5hAPuzVX9PwCLy7pcelJ3OfnmaJ3ikSknDDo++cmfcbjbnnOI
E1LBs4adtWDCzn/Aqe2T2ddqxXWU0gpl4QRMgjgkuxu4b2fEEnMqb2cTdS1j7jZu
ShQjm5khpLykm6lLzvRBsWmZr0MOngrgb7+2GXuImh1wAOG1JSdC7vnvbLRQdkvi
eW7YHq3s34oxleAHtAY3VuT5JnerkWVL+zmXAtk1WUYW5nxV5msQAliyxVaJTnDX
u2xwRlXf+B1g4WcsGQKzUaHcGDqbLzQqbOCkGNlVJNgesM9FxXg/lnF2e1nFrVaW
TjYeN21+esYjutEelX+EhJyx7H4nbjlFN78khyJPNCdZNkwG3563a1pUd8+ZTV/E
1JzxBi2ijquKKvLPJASAB6HMma3/Okde/HHiFwdU/MSCPgEo4tkFQuyTBR9H7Xzs
F6CkArMM+2PQOFcZyxLc9wdG9vOravBXinn50VVFfbujwvLn8egri96LvvWUNHVX
d01XSrNNWTbqRnVhLddPBC2a3HdMWa+B9TacrAnxPk70ql8gQDsZtq4MnVFuWzVh
0FTKCEmb20fL115itNwf2GFOntdubkEGP2OexKuuPQcSI8e5fpSDh7xEN045AdMx
kt2yOmTiPXlpfQhzdqJIYaZBUmb2E0qksIgHF3t67Bvj70BAX0z9bWaiCu1Axbx9
JXZhOOlRhCYoZutswYEohX9/IO57H6jqit7WUxxzcSf2aI/OZJ7flPgggafx4jYJ
KYcmk0KokGBLROPB/HUKOg8oNE7Cd6HhwbzKEyJgakBrKQHEDK7Sww4R6PKNu00W
XIbY5VPPRlIJxnDxp7X3dWMUeLApuqoy8+/xC7ldEOF/bScbRaMlatBIPMqGScNg
F/l0ctDcldqNX55iof1EPidlEm6V/W6ILWcJK+4/l1SAR9kBiIcg8SRWvl1rDRcd
7GHd14et7WlzwbS/qF5chMu91kRshwLFbziH1tJI50sKJSpbOvU94dEDeXrjQkmY
gewHjf8c1C2Sa70F20gAoC9cMmfHT6re7snIE0mnLmAhR6B85WfgfPmXLM3RlmzQ
9rhCRFKE8xa96tg8lp86OQpJqb4ypoE+4mscA8zjzwbijIiY2rnm1nMncb7rUmmo
JQmjjRNmm8EF94OJJLydNOYA36qYKVH12l4D35827kI0RgcR+w9DKzX8JNCDNw4n
r44YxdrEvVS/Hzb+68Cg/r424HVFQ6JScfFy8lNBY18MpD3UYHPO11TXGWpXs8Wj
Vp5ZNaVKQ31CL/6UegAgBNIf0N5tCNfhbA+79wnW9xju6I3lQ1WSt8jgeyhe51t9
nlVWsRos54mqSRnIhSnxjx+X3avMxBH0f1+ZUhMb0m7CBY52cSF3JJXfoIaaRs7F
0PXna9Z3kmlWlJLs4pRd+MLEZV0muvEsOOa/g1terx5Rb4jRLzey5C31XYHb1qxh
fcvELv2QNHFRCGJy6FV2sO8amT2FACTZxGSEfSLXWctw7pLXWWGndlT9W7ABqjRX
0JYOYnzsYMzgedIB8i9ldfKcnlF3zlNExhTu5prN7k/QHmY3artgV3E24drMnziB
VbI0DqMo1yqVVN/g+aMaT8lz3lz2fKqEZEOrINnyUFvIThGcY2zcEsIxFFhgMiZ9
rMRJ2cLvj+F1kkKSH+wY8jyOxohkUtpGtXm6BJLvthTB070m54cnPvV3FdgglJ8a
K2DL6Fel+/m3b1X7n36fNR8t4ZsuNcSu/muRmSHWZSe726NAqCjBWMJt/jd2T0PK
kypQHtmBgHUexkah/LwD3cBQZ07VLK/QJB4UTeXv6V6XBMItSB5fXTcFJDT6pEhc
u38y2Ew5JHuBVV27cssTY+MqxBm3XNGWFfltxTreeIUts+cThgK1YJUCOBaiyT2w
37KA+qpvsFWS0qiPy0KJdxT++o21dZ9394tHxGj5tBlACx1JSzzqr48p69ENZ60f
8p2roKWqNgjx/ZVDlUDlq+sIWK/mWFjNRvode60S1IGRMgBm3LXneK1+FLkkaNc1
CD59uWfWm1JSO+CG0EHQMBVLiYPOUbgg2V/R8IqbMWgvXCbCfQMzXNF8n71/AQSy
D838CuGBO4zGLmHEQxju1n3HbJXxtpFPlY8cUS1MamTV2PCiZGW4SPdVZAey24r6
ZbRyNvy13FzQO6vVpWtvRxbJ05RovkUsDL8azsxt24m/dpYhb1bMOwbmV++WZIXv
zu9gqUt5SRV4EOD2gNx823DnpYmwvwvPe/n/g3oKjxW63dxj7dbjOG76tRE+C+jO
NUFQjNVbGt00ddlWIh3oSmOedp7rALO+YvYNgVAPH+nboWRSrB4LTLfXCjmqWWcQ
DN8U6YVN7c2x2JxTSZozLvpVCsi+b2XII8Ct1lEpUj7nCbWprPKoFB55cStqqbEx
0epOtCN3nX0cZKpvbU/9uVu2fNW1ickoodmYINxAFO83DWlSGKhu/NMkrcxPE9xf
5ytU/oPhuQ3gLSgF2JJi/GoFAfxX2DrWeQZe8m7jP0SRB00dnrHfmEqQ66ymeunj
LB0fIgk7ATTc1SMQtQUHE8QB9VZYUtNvu4Le/ZCwub8tqs4dLttfdTm3opf0x71d
V8qKtQjpWfzQRih9iG6EOfXPxhwOVQbiDlCiR7xzTK9Ui0Wh8veBYQM5PenZmpoB
hNQoDuumtUCyg6COFhVGzqSjbcxLwQVew8x2aATdTjKtNmdGVqOnKQG1PcDepY99
zzFKObR/vqhQX+zHdVV2eQ+NOVGspFV80/SHDQreRzV1c4DktakrUS/Ko1yYXtto
wQOwm+ht3dWrIlJPpLox5jp2AwfyaXFgNK8EpmfkIKKbxCFnY26G/FxK9vaDgaBD
sn9R/5MYfHTWdRuTRN8C7XdWdZcFRAm4YKr4KFgtnmSRDhxix/iqo2VdAY5SRw5Y
kpZwtTFh8ov/+2cPEVNny+MrovFQ+XnCC3udZpx9lyW/f+hwBFe6jJix8IgNy4P5
kPkCuhg/cNEwqyqti+MP2dI+PWwrfERtDMm/i5THrrKX3eGowfNzUgIRTzUFrfmi
83uaFlg2wlP1+LEURXy9CkZM6klUgxncG1Jhmrpko1cWMkEYXCsHGIWdKqhxTk18
LR1D/c7KA0nmpJLAJpt+ZSqHGLWPvDYkYj7j9vE6YSdEkwCJ98gA3LaHn4/8zX/v
FHuJ44jagspgFGRm8IQK7Q7CfJCior+0xtQrZ+8/Ci4DPS4qJX0krEeQMM16IZAy
K9j/qr/COzLQmNuGehSPq4iEhOqw5EN4TbPTpghcPSbdPkrL2O3hZeiaeddZi8B0
2qKckZfDBZTovps79ra7FdGhfHa/uul6Ui4+C9I+TZ+BCrEvGWWRVFRpVK1AkSd6
V9TJyoPNfKS/tiigQUjW0EYMgL/LsDbh3VcJeSaqL4d8gv4Aa1suJaK/SslnA3oY
ntbZcO4PKAGUszw6SnLyNBnwOYby8l1NmjaZNsxhf2zDa/c1VE9aTusFMAb3b2Eb
DyI3dC2km9MOroyODyWpm97wUpM3vwUTzNwhJsA7lRelgTDrITclLKPEh5RXhw3j
yAcRVQ6qGjY9HzyQw1WQda3lRSf1b74Hipxpy7gHthIJi4HBF6JRph56otCg5ank
ZwqKgq2g2alY0zmYwbGd4dtzKykO5dseMvhcU/WgJ/zK8qtISi352cwHXmoI/MDe
TVZmVHlMNUjdX3QBMG0wz25aWW0XhkA+Bh1YO0WNpQRV4XdNWfOU3t1TCozPr2RK
aOx/6ZzdqCC1wDK1m69Pk96uDoZuKZf1kHmHvclaenZbT4bjmSd1MZZp7pLagVvG
kWlUQIa5r72G+jW6YjKt6/kYpcJGCyxudk1X5Bk+2r68y6PZ7RbCWVKGvi2+OpFN
DQd1Qr87GIpqRjlG4ygcmdqKy/9Cexmef12hKSvy0wWtVvhFnv88TnMBIUVk6Gqh
3p6X2snt4bXt7ln0JySeQ7qZz+fNsw12K0DhxvMA78yLxREKKVtkyebJJ98c9qUV
96fIiFA7Fh5+nCcnzGX3+lwZf4hac9drL4OmeRyXPZkLMpOs5wj8fxoEBMHMuE9z
qF0MSescykUFPNsqJSSxpSW/FM4sxoDVHzq8nKDPylSR0LjiBN6L0MxAdNDClPxA
EYeX3pXRSj3p2oYNWpPj0imnuxYlx4oqbJhXli4XnwPny/M3YnLZ01KkzVUTjgkz
7hWGu5wgILjS1kBrig9TreZPUDAQ6EntlGVdT98D+40pLfCHgh8DZMeteVWqwJtX
Pe/t7AHY/zzPsfB23+wnwFG2Y9hNeTZ/rDU7IE2bwVAsUyXNjGrUAR4A9zAoU2Kp
OntGa1A8ObqEDtiD/9EHJaF3etQxteELNsJJvjrytm4nm40jsGWpEnR8ZmVlVm+Q
m4XNx1UQarNUu05FogMYfVWdcol68W28Oar40ILskoufn+0Ir9KcBWu1/mrk/Mu/
appbhOsqclnFt+LmLgzfnTtxJyVEF0KiS8bdd5GeHFrzEmkuy/WYsGJJqPPlC0X4
1cnTI2+nL0Br0OXstbVRODBo9fJpgomtymu+W5okz9gsWkCjJKfkYCKvOzg7P4y5
HMTfeoAqbIliJJCIsIWmSRBtRTbSQQpbPveTe9piEzAmz3kWDlmJPo+tXMwL8epW
U955jngiW1ebhznOg/io0c+snl3ohQlN90KIb7aDUg0/asEmJgp5NDvdHe5hxMfD
0+w7RLtSJwPOhaX7rvcXTgQDujER/HxAY4A+g18MojHy/seHwMQZqQMk5/75m9R9
WqoTq7uDGBkas83dPaYShcP+jFubCSpYeZwynix0aiBKI5VDSuB47S1xubqbw7al
EgYAIG7INnjDq1O/3nEdSvWqyQwWBfX4hqtRL1bPFpTuZ8onobkpzS+2j1Ymbyj+
lDyTO6ct4mhFmrfQBeO6c/HToVExlRH29kQEstkNaw0l8KslVImMWWxqt9obxrt/
drWicrOYPqViWjeE9KVznxfBBlvh2vy1PxGQ8+WEJ25qBBJ6vLuMWpTMIhVZ80U8
qjaCxv5E9eUOAwmHCzJfaVOz0EOvY3g1xZ/986wcLV8nDyQHc3ezBftAoYrG7zIn
IYFBmDhNgHKkGyDpr/Nd6NYYehnPIdyUV0RiyCkTZPixLpbvkmK26tguKnKM4/0z
4rJjK5+Tdu/5iJnlQS+Eh3LWRSNCyZZEfXxL318pnRXgAvl9VguA9hSO4u4ye+Na
riWedf/euWB/r2uCdxQykpFBZg96/BHJlxt4V9huTBC48K7wQaOy58kCramsEueq
U6iQnUgT6SsQMeH14if/jRWi4FkmaRw4e+jEUXQxw+Kb5f1JOuyclXNlng33BGW5
45FCE2IORh6TEr/rFleR9dF3HrWfn/yqJj0HVLWS5hhJszDyxW20S2vO2dRE9kp3
ft8Q/TTr05mYPESviR8DhZQwnnKFJBmsdrQBFrbchBwWZjra8MLEYnYj408a1UYh
IDgyBCyY+An6BugW3QGxy+XUaZ1dxO9F8dWT/S6FoyBax6/OPgL92OP7EjW1l/Dk
EH8ksLrU/WJqD9mw/tnOVifDRzX7Emhi9Ev5KlwVvXRFUODKYdU3IfGozTungjcE
nx6MbBA5Zn1MYkURtloJsD9fDANabCX/ynFLwIp9cnvdxH/T3SeDqYZd3gopC8/K
inJEjk+TiGwf3AJkgkCn59rq57H85sXT+0qflDUEmAZH7/REAjqxO45YZntQSGxs
KQD1W6V+UeDR1hg9Ld5kvJEgLiDJUMTrG7VhwIpYFkY5G2lkdo+eL00nrWI6uFZn
krldrBcZa9b6DI1LS5K6sXsO2v19GhA2skwT8V9Aj3h7yzyrUMJWNBO6n0OKc5nt
MHNs+405/siGJYIqXeIytDA+lRmRW2JBoqqfQzo5GdtkZuO4kKv3T4neglet9fNX
3aVVAVYmlcKxZNWK71wGrMvERU/UXT1zQrcB17mtc7EIyXGKJheVpIK2gwHbPSwz
Stda7XS3ZqykRuSArR6Y3PSk64J1HPIKs4KxcFNkK7sPCmeCdIWDKXJkZiaBeGQi
hlaFjC6jQ6T/rhE5iCkwq/KaP9jO3SFXiq81qZSNP7x8jgN8o7MHjZT9oGlTocyL
ahFkoyFGc0fYi32CcEtpnRub9nUxbmtO/OWbSQ+M22ktniyPw+DnkjMyD3SE+ntI
1867/mxGOMMSgMsMejTj6jtmSonyeGVqxL4PJCe+YSuE43NJX67b7z3bW04T+lOp
btx9P6QP5v3ZIYOIq/F54FBBJgnyB7Hu9fFSUZxaHn44hPifmf4W5Gzw+Qfbpzh2
Aiel5H4X6w/ktPlB9wrnBXiGo4rXNuP436cBnS/KEOAaBU6jZTm0OCYq340Zc0w8
adYt001K5XTteK1QTYraBFGFnl7t5/k0505RLFWEFc26vFBvZkDa++8mjxRjQcFX
5UVA70VwNigeVxUQMR8BrTJVbPn2TxCARcppBMY4vkmx1nt0Ab0cOl8Pbf7qfJhM
V07BHqT0fmXp8c3U7uEKMWuHWGNkZ8iDraHyu+S9aaGjaYrW5lFvIXwgzanCTKUR
RfjqU4KGA7VvKGiQ1TK+7IwIxhe9kU86dDKz92atJdxC0QwQ4tOR2UQ381XhjsuG
GPK7av4gMlzkstTyacZdxdjkBuBwTUFc0qGByfp4dJETgqjRhegWN2nf8k57f41u
NNEoyQ8pMSu6vwP8FVZVSn8IsEFM9uBLPOgeVYdrwOPZXYGY7NT5zNW9coNwswxO
pRXHFaxFPcp4b0B2BbQqKWvvvzEflYc4kgJ43i05n3VtOLNvKJ+UVZnqymxuxKfb
bG4/eZ6Qs7faFaLH/Sz14mNN7fOCP0O4CACbKwcewMsc0wFNSIQuJS55Ek3L2anO
dfYWges8TbceMteFTbc5uMjESWGH8ieBD8G3OrrwpFDGLnvCth//BfMZpLXRRzBf
7UXgvEzcJo5GkPHx5qHinOiviSzqOI0Qh4uzYmGi2kLv+8WAoNNhl7iW3Ej8OBSb
UAx8edUO5FE+earjN70PkNwusLVng+5hqQsBGnxTbXQJsHuHNPuprGtQcUhSycx4
dejsf9vD5FK839ej8In3brUtNQqm3Y1rJPuad4RQpSfPdmTFxWpcLzjqEw8pmAPM
Md+yIVcQfAHOesOlJAAMm4hkaNXDNWjTMcDyz2WSg9lgnn+l7h/w4hglstD3qai6
Iiugr3b6NIUmw+LZcooyMltTH4qi8LVhqLfNd9jTRVSkZl45GUBG16AEOY1PxxkI
MbqHdDTvXT5aJpBtGpcj8qpAyfOpf+dSsr6fgkzD4CyjoDhOMNNbYnQXRSbPWJ8Y
TnmMtINZtZqTamWaYsMJKF3jSSeJh450gtTRigN01XX1P2MVK8KQIktOzf2KzPfg
bTMBdMIDo+gpOGJXUoSgLJZIMSt28CK/tQIT0jI4RM0kgr0iLwJCWud5Z2QAFHZk
XCEsi3vtuQ+7XPRuveFUllLqTzR9h0w/2WNUBe7OiOpQNy2YpcSTPPeYpP/lZ7Q1
WnmYqnxB1WFrLgyFpPqt9QsjejlE/JPwnYva2UK2eoUIWasMqZxsSKK3RfMKHkhu
/3+wTnSd2Ca9qed7oghemFYcOwsv/km2MpSZRZznvUHtdLYmF9pRkVnJ+PepWia9
msQd/raO6Sq02EWDe8hZzogLaSorR0H8/kA/GDzCYuSamVhtS5l6BupqR3FnbeDv
JZnzQ3CxcqNm7G1FuZcWUr/n9AZL0GaFtqD0VMwdmRUWoZErzlWTB1NJqsVGX+9f
vPzJXtfeYOqpuh+Uts5NEX9cd91vFuodXn3s8mKnr0iMNBm6S3e9UMmotI836gQJ
xD55k8BYOj5nkITROVFUF1gZKBJMhpPiF2XK+hFbl+HWAVlnc5fePNyLthRStVdw
ts7rceHBvunY5h7ijxbpSW1Aqio1Tm9LyXlZVfSmeQ4Ur3sgfDl7dTmpne9irvML
hLLqw1fA5VE1wQPA9rMazuEs6wCntgAQyBcrn23ecOJ2Qeunjk8v2kFLa5Ig3NKU
CetptsEY3haete06CMHCNiulainm3nUEbVLb1porkegT2XcSwuRZi+7uGvjtEOdB
vF7AmzatARGsSpJfHxIuwcMQWzCrh9jiMIU9qthj4dmALEpXS4NFx45rqF3OIsyZ
SnQQ/bzpva2sJ4V0nrKEq7evkOibX+Tlsp+XFlCLXMa3TN5AZyiOmopt0zU8R6rB
yZNS6/mLaicEn1XktDT4qT7wBZvZriDaua/kP48uCY0XibCNVTZdOcyY4VYQBaCp
IW6/Udkr+Sw+4/cBzdo7qSqS1dYnt6ZzE54df1nKwYg7efbZjdMw+MFUa7ce99En
/J/s2cig1CKjD32wAUZxZukxCI24jQ51dD1rvpoVIFAULj7bzKmDF95rJjtup4H9
exWMDtBrBRph/JtWnmhOYxZy5O3dGF+n5JVOy7i/1VNj8vojUjGzcQ7jnUQExfFq
8zG8VNXZlCa6JzPba1N7dB7s1OTMoy9ElrEvbuEExLs0vfQymRDyboXp8CBpK0Fd
KJt85oTYNA4i98hMUdk5EKJbzjtwj8DRLyex0zyzHPCptUIxm/sz6iSbx3vNau2/
DHX8CGO4+dU5p6dDWqgu590hAy88sniOl6HZB930ANV4E4y2mc6paDPBeGDp55pM
m5m/UjYRVzLDNMCmerE8/WYJ86VZMBpYdP72ECXCQGA8YHepOZroASqK2yztashf
R+zePL5qO5ISy67GYQmh5WRJr2IoIzfiK9O5JTUz4fiQ9dnb2pgwT6XqBjYQZDOf
MsNVIk0FZF49nJxGAOb6pubpskJ4w5LposU4PV3vnVQZfz5NMiLCUES2jUqdL4Zx
laK9oaRhgZBfM7Nlaxam/R5ECzUxXgfZ6WSeXPb4DeeJn09DQv41vLEu8W8/RATy
nK1+UK+bvcUM21jYxHJ2MVCof6v48a9YlbDpNdcdL4hOB8dFXBo8DgEimolchf3y
T2R7g7r53Wz3LYr9am97WuO/cEvoTGiGQ1o+CkR04ec49ClGPPIoIIf71ltk/Xz4
KmJZXmPy4KyA5hoNg9Y2V5KstRbQhmGYyIoo9Dt94/iPh/AJ3Lkm1KXKYZ3VMZ19
/5ufruv7302kVg1kex/oYCUKExT8kn+da9uHOd//OVa160P33nNoSmPiG6Io/c9+
OPgMGmE3LepIF7j5qDhexLGkedvOS44TWKatiNhJugY7SN1qGg+XgV1l6KZ1mIGJ
s+rwgRv4u2PdN/xwPxnXWDEovab7qa+2M6+LsM7QAziemyIFfnBrhj39noIUEeO4
gPWglOL3pXFL4vtymXDrbyC/60+q2z75xMeMUMa7n39eFxeTMJAU0yrx9mXP9h1D
8MxNo07GyoMovnY6cSzJ2qy6muiM1gCIzIC9duleW3nLmih+nyGO7CVJKef8Frd7
RABhFTpGaOtpQRKZWpqeo7tDUMRZi8ojcDQkCzho2uflQwHFCsk5kWclZDZGzVtl
HCZxTPlRZ3u30ST04bumXmSdmra3wAXDpqI9f6maRyXHoUn5owyE0eOnYXTX9Rlg
aEW2mAzbUOkaQLrrEFL2O802HnjOW5rMzzDYzXBJdrCL1pv3XOS5hu72/pVgsyAp
fK++hwQYSZKNL0RGtIy84w4aFjPY3t8S6+U+0XuVlOj9ehA9rNCZSTcLTJWQvl0i
bKefPihi9cdj6mKT+Le83xdol9J9Kh7ssqBV6XofJ0DRJsxpnf0kkXK6AnGeTCJg
jeovcgWbmbDfKUCKIifxgm+9zN/l6JWcITvZ3v94RfC2bBJxY9UH6/RfaqOL/fBp
oG8MZwqpjf+sUAMSXOiN31d3zRHGR0pHsUNYAi4t6d8+ErGrHGrT0BliFDaV31L/
upLhqhEWdCofd6+T/rRXcIuWUHCyZIBNP0u1Tc3aXs28wGgnXHQLwrs6PdX533Oc
/hKz4KGU5yoTAxUhCbxtrgWNvTJvMo6SrUvE+iT6cXbc2ierik2yXQcuB2lQV7RY
FnDFX3jARYsxjYghYk6yDY081VgxdYwztkB3QJtlLzOSdA+IIxo6+0Dsw3csfQd0
x9LqSWN+enJabOl49YmXJQQOGdHCxy0J9YeLjWhJE4+G+TzTzEJ5f8NUlnDOJxwT
MYdeWdspkEufmFy6SvMEWXXCBjWnIOdRjxuIaunk5pq1R2vsiAHUXIaW/LhVy31o
95IgyOBasrYRP2Kx1P7eHmdHRaTSSDucOndha6oiqdIX8TgTMDNew3TI1ckq19sl
HJx10sKLJDVB88nBXG+4sGvb38VPL/vrGKkPaV8ld4aCY4dBd1W3//vpaYU4rDmr
ISCpxtsyvctPJiuRoRsGxvWEVbQHgGWDqAZMrgvHzYAVSlM4wEjScS+Kd/3gp/qE
dlYC2TUn8i6tMXrb4PHXsIGUI7zOfSNlt+4pOh2I2XmiJ5CypwxApNpHZrhhqdP+
rnUv3MQ4Nwm+TaVFA4EgV9XMEpOCVVF0RxA/05dcMhEVivIlEztTly07qRo7WW6Y
L7VdkGrm/dkh7JuB4RmFqslHFRDu4/X7ts7C/JqNSnBZJnwrcvem6ogAk4GKi7Ff
8MgkJJ2j6cUIXMUuytjb2tiu9jADH2sL4q/Xhn3XIGj/fPdMHAt114RefPFVUf50
8e3a76RuQhSiBue6Z0MEmliQvJD8GbG40Bau6DTT7jCDJTxoCI63wxdJiBFl3+R6
l2cDdFwnzME3bOdnCZEOP+UO6zQbybgT5W59iD76uGYa12QgJ+Ovyrq0GoPtNzZ8
tlM4NxK/6fhRbCLeMVSrcFfjs/bsj0sFZ+33Bvt0jLa82+G2Ct0pA+vTG6zzPa/w
izuWKf+GUemqWVKh4i32Gjs21GpPaloCjNSMWqcfw1D4OtF6CUj7WE4XKYpgUozB
otlZ/92WyxqY3W/fxNIJcL/XUa0rQyN8dsscZZLfmsxzNXrnLdaGvgVxxgYVqWDc
k05yBbuU3fLeP115HgnlyuDS5B8Pv1E/5lAoHfAYobihXmTDUMCBLK0lUohDqA9E
QKAqEJ+hkwzLsrIODRXfGBiOqpbtz/5cnm/jSvoOm5m3xr2RMvCH1IJ4At40DngV
l8iMjMez+CvTkqxo+tLiEBuMk2a+thIkeAsEtlsvwDAUMbmsQqMRWxmxMnK5wm+E
/DWUXKwieBYayPrD2b9/uGpcVHYD731VBbmpzLERTAD12j1Qz5kt+XIInQktEErE
b53ZC1P4Z4/kCTRNnk1m2SohyPY11lsH2M/urczWjWPt74TUuaNDNY3cInl8MTf2
RvM2nwzEYdhVRdyt2x1w+YL790sqXKw3iqPyLPZTuUiL8RfJoGUiJSXAhTBjF2HN
AZBqBW5r4XqCmOYergPdP2TaqdCaH3M0XOaCeiqUca+qbV6Ik3VmCsGEdMA5UpS1
dLjUhL8CJd+H93vEG3Kx7XllMZNM4rnfco2b0Z1ASK4dZ0PhmDvTwbZyH0f7oKhX
zMOmKnZBvi7+wdvo00BCQcHmLiSWRZjsH2BdQOqRmIC/+jouDF9Mn66pof+dBapF
Elza+AZwzHGKMpaaKRfrJskUj/REqd4RYGbb0eM8asdGbfu6Fq7fpV3mz9d/TMRL
XPIRBA0ae+TOGIo/JpZFV3FIiJ0TMLzgUPLdPd+i8TLbgnfwglTjSBgs2L4xaM4e
g9NjW9ziw8FEeKGdO3oe91PyFtqpHXTRaiQc+DEaIZ0vt4rOBiWWUHGSfk93IWEv
ZzsFa7H8IcZf/HPRKo7ZCpEKILhOgsnJJAClLcTw3ILOuCZCX7DLNt2miRRz7vGT
84PivPQOGX+Jipdv9BKnILDdfrfaSys/SPiuC2OMETDpN1c1+saK/AtjJJ2fM53M
j2DzikY+Fe2Q+2VLsGActljXvX2H3ghAzjd0n69hkPAswqTzZ89Xb4aeyatAmGbB
p83944z0I0fw6VvyqiDIpCwh/gnweFabi5G7KB9AXDBJsiDAqQSe4fEG8T+3iCjm
fakO0Jv7RZfyymhu8H5xdWQFSQ86SKzEZa637/0FpncRWFpMvBRbfqiXKUVn2jOt
sRzPqdhnoPj2OTcGcYu4ySd3OfLutEGwc9eSaIAX4FUxNTHRfWIWFWUH9c6DRhwp
j5zc5JFnkaGQ4yEauyibzz2TZi8RjFg2pr7JxkSGJy4q2OBX1qYatN4Galk4JfEm
VtguTEwXcExFZnUr5jlNckA7CwdXrwgzA+moU7IGqdFfDyGVvYlyr49IJc7xEGO+
fKE96l8MH/cd37WYncQL5+8+Qo3m7w04rXlic0R9dml/vOsX8ETE9AtVqwLTH2kS
XBPFi+xAQqwTgP/Qrg76fP4ybVxwX2Jj53rEAMXr3SJYGKeJfTcKCYg0Bm5KLsep
BEttzgUseK7bX7OoUPIeaA8vNTg63yfLfJp/sFheRrs/XXJ6KpyH+Yu3JtS7zfyh
wF8Na1pgnZfRU3Mf1afILYySD10ZJcBcu+9SHUY1qm3SRY2EP2Gd1qymX9QBW2rr
vXfvpRauxq3Rvw/6HXvSk6HMTUmlcyDP74gURc8ksD44GufugEOUFE+2nBHNMV9X
A0njprBxJE4DzSV0/SirdMs+sgIRkSjrQkFa3nsRrh/8FnBWMfOmtmJkHUK2mEsq
1XVVGVaVu24hSngSWbiIEkJ6rEXKubM99caW99xKiGmYu+3zr3070glcEcRF6nF8
T0jR+4J1FLMMXDNfPQoisvJQxujtGTddifw75+2f6qA9442Foe5u67ZmmJCBcoMX
qX577ndgOJbl/Z9Uws+HN3WYVRtE/3WtIWcsvhAFclxHldXpho60mNXtB02yWYfE
S3wWlzEuTSD3VYKnwbknWdBj+m+54KihwC2y2xj5s8VDLfI24rk5WGcZUborXDWm
ga5LpqBYuIJHlHIg2JcaaMXVCIY8zcUQq8sSte6+aRuMJqJJuwywnv1wDmdqP0gH
jAfqPTfntTnblYNU5aoE+xxHFi1UfU21yw6cb1JfOctSjJDHOtXVUCTDFq1rewCK
5rby1eDXLw8sgLm7rERCurIKflKkgChYVnT3qWQAW9NpiEogofXCKjtwGetaoyYT
srj3o1CCGP7S5iTaVBUVJp5Jch0WBGdLlPUvD4svxj1+WMHT3LZ7Xsx9IW9kIV/3
nYttPuJ4BVc3AE7DsAWBzAXQdA9ctMYzlj9awSisZkhSuLzTJPYT0fQBSAAkVrMM
IGDEWw/2VucTc7WvNpfkJxQ9+diF0gMOCBNS37i54IofkkjuRrGUlHsHGkGAB2QD
v7HZfIZ7ai0XGf0M7ySBc9fBKkazh+8/Pe9ekug0mn+Jt7PXz39sa8N9BlMnZag5
uGtz4NUP/esR1SdCsXfOK3Vrrs/HxelZPmXkNTIKQ3LjqquJccPDhH2q/FFvCKxQ
sBQEwWYQTMFaritEnyzyNhne3y5XqweR9fXiSfULzacNUombfMo9+8cDviqtPGY2
TMi+TGLEbqMMViTq67ZKQBz6mrrj7JjTaT3kNw3yBi7x1HGF1K4tZuqoHj5+0l5V
tF0nvWVPjW6nktfDzzjOZpvHfBZ3Vwy0YQr7VnbRj5cFKOFWF0U+gqAGjFugVKNj
ltHYODm19Og2V6Mg5RpLox3EgRuQAndDQzLp/CtCUF0rfAmMpx3aSKHi9Dnd2U7s
0dCcS2NTd6SWue288Q/5z2zMMl3oUnR4+oXMj1LC1rXDlg5Sy/vI9VWRw1fCxdAT
Bl0K56PJa+emi96zEuvOZY9tCcG1dHZe6vdVzwO3pMD45NbO9209O8jg7k008yLP
B/BRRYdztEGOjc/So45gGDq1MoQJCX5t8svB2baoJiYMWNHJyztsJJffvSd+gvLh
LIK+TwwDPtGG1CKJECho73woO8vWQqn7/CGnd9VKStxAsH6SAAopdRrKD/lTSekn
wnnyxUQ4K4/jRZHQMLBc+FqJzboP6mmisgvAstfBLYeph78TyI2x0PkfHxfISCZR
Fh8CjDCvpKgyIIV7fbFhmxdPkI6YiZtQxGCUgd2dtdDvh1fz3yIe6gnwOeGDwt+y
9hKNzNpSoqh1Mriw93rkXaNj/oDmoWoyy3eIiPn2hCtZfhahyGcsroJ0BtSi1LAJ
0f1A3xuYmLkmzMoQb4T1B+3KqjMlD2ktLUQk/vxnHX2aNEDoNeQsP7maPDKmKxD2
kUwhMCz1zhk0pK1acTgGqSMRAe8VCWuVgYGFHn/pCyasKgn8qMsUuCRBAyiNwAbT
b7mcy2DMhRQJf6mWeVq0Li357SwLh3oP7sdU+cqxlOOFbr81B3o1Lkmb1rVpFOya
q0QPip6yo3GnuISWvrtXx0it0/I7yNCTmo1z/lW+sXnqpnXvocpE0KPeH+nmbzd+
1XtGYxOAViptf4VHzqTX6iFImfBVr61TCk8XWFxn0PiNq8ZDRqDsblBX+ReBSNwU
HbwxZgdWl/Lwl7POeNN0IQV1ILXx491wExjZRWFlGIMSM8HIwNLenXHJ1NCpziLg
L0qULgcfBWE9d3rzBXhglEVWjjdw73EBWx9zT9AY78EYY4l96oMcL6bZRtr07k9i
rMtngG0VQcBlyKWWhDsqGhiiYegMOP4CVZ3JCD9H/sH3G/X/I/YkKYX3cJLS2gPd
kAiMWLYzIZU2dVXsPR78TGl2QgDaRm6FFKEULwF27mxxUAI16u6LOs54oNBHjMjA
j7w0S72uIDoHW58coPVzyKUi9vXXxOAVOlM2aU7Vzh2EWBf1d0cVhELfqEjW+Kpm
8fulGWv11SlfFZBydCgZNsmNppY1+1tZNpjf8kbNqj04nLjH6CpT4SDOrbZ9m/2r
sxvMkT6RIbYmFT757DEVyK+3BNETtVo8GeaUgviKrhkU2jnM5iZMekLUXH1C8eyB
GMiN2q1o3x5x+Xxt+jPGERFhT1G2qIxmDR4r5kWRMoCukh4r6E79fDNOY01Q9Euo
GmTqj+CBpdry/43HbAP+/KlEMl8n0FYm27lvop/mjR0UWts7SV2I5BTN8suSyYCK
um6KtvXyCu22OZSXukwarig30tuKc3cIVTlVVyBnmlDu5o7x6qtebNBFSLWiscXW
1UfTvnBP3PnjoYWOAOSw06SrBegvM3CEwXF4If/2SAXwleZwuuijhcRLd1Ch2U/z
WfADen1c4FximsOigKI5ipNMqjkKCDuPbFEEZ/BBC2d/KvgrrAiiGuYYuU/ptHEe
cRv4Lh3pA0NwrOHXCTpQP2YMqNPXEmclQvpgMU13iOuXkGa5vpVBAnbCb+VItmAa
MStEwUL9VxgKB+iRdyo1/9/4cxwIotgK8+rPcgSwl6BfiXX7ccl0pRz6/TJd2r1V
rnPkr2dmEZkKj8ORGoX6X44hwRTCQxD05hDZgxj6LMiy+T7nTsAAUg3fmkoif25D
Isn4iOokAgzOYp0vaKmwH//1BddjdjB7A0f1krHqoq/VippOiD1sDa4ztfLVTNH7
mg3jmEUa2iw/SCfnPJ4/kzwCFHFroAYC17xgd73GuyXWDNL0mOGwBbeJdE1ler7e
9mHbHSrZachtzlhSaHHi7IWMwD/evSY0HA5gAtqvD2cuIPxDZW6VF7DOCPjQ/rrd
tWW9IyWJhpVPSi7JBM+ASs4SXo9k61IPyQlPX33T4JfH7oOct01+MhmA05iQ2z+P
yVhj56DuW0PimY+MmvcAChk++P2r/Dr6LJZ6nNB3FK80U/rZx8IMzTPwQXvWRL+b
Az1pdUVvAC51IoE878FMBcwnDj+fNEpVgFBDK0lrUZ2i1CWAjl62y0k0zshMB9Y+
EsaAvJIhhdfMfoOKulH47hCJZe2f+kVNptxgU8HKHD2Egp1rh3kc8+U2VTw0Dsy/
Okca1APkAe6nSnSxqVcSu3s9cwsV+X8y5dd6KFVF/+KZp1Kju9k+V4Df8qi1QV8I
7aOpkO36VTJN85OsfaL1EngabugdiYpJ5Watatvr+FFTSwkN0dTuQzVq7AKMHyG6
C2Gp67HqrmgPN7zNopmAILmTFePXxg/AkhqUSjQBzsnPXa1SsH5lLU2Ln8h8TPDz
R3VapAjOQVrsue4r2um94xlfNUA9xHTPR7L5CaEOJaYkAN04r73nq6T9me5QM/BU
2c2+OOp7I73ED6Sks8Zu5SXF1yL3A9auwCG+sNc53dUBm9r/revEa8vb+xamXWmN
9dEN3XUAsFLaE1roGFQhmowC2bFNh2rAT0yiwvQg3TRO+7pPWqCL2SLqJojKaIuY
dmPoL3JSKTCKA6XASJP1E85KfeO8WWN5pJMlmlLwybiMc4/zZ9nHcbYx1M2uxvOq
T14KTlMVVqPFAcy5utvrOAiRe0p1OOvFPzkKq3DgkN7vsd/BcBGkn3o5/nnGlXFv
Hu1pzD+zt4Xa9yUYXy4gwjFhB0BMzSdSVc+0nAKJqBLemflY3GblH3xtjS2Kx++a
7+lBT/KZ7Qqqq1c0+63Y+5JiaGkRdXhaMH7xqed4NDYX1VOiiZXKk8fYLD0RWAtK
cUjkve/GjDh3+Bgjkwc+ZAD4IenlFy517zbmExF4YS7MPeaRtRVkmQdVLWsmjsPM
a3vvcYcToef1IiEIi+0BbwgVluL2rw2GyoEJvMJ8jVGimXE38phcWc04nvNW/KKF
/2cuZty4fj5FhWeowxte3ABlAo0wRfZ/vzkULExcjj7EtNkGwF6K55Bmb3J+tLCW
eHN7Nmf3wQMd+izglhMWeQUzj7Pv9DuOLpxpXp+YWngwi2UT6XfYGwjEbBgjvLHM
fP3jQS1dei1tA79fuiKfw6AyhuE6roaONIugpb/mhSweD7sqqezuNS4fByBBI9+V
WWlopuSRAwBRwcVKTNy6SIXGg8iYb1YLyBbccXZAlrcm2WkaX1LcTzn5MfNla7el
DjVtnWg1t4n55LyH/HNlSx758GDqr+96/xzPxu7wjsR8EbVJZ31dGlxUQrgURvM2
HFfC89Iih6LEtvfdfCmNWtUXDe7C4dyjschVcOUU+eYa8qESYSADpAS/5VL6hCk2
otxeYvXqFffhdVYFf3050ssxVunEO6G6i+ZFhClQVVNOH6eEIZcPka+qS7gdum9a
CTvYEErf3dsgUb3ckjMUBlKCg9/h/mw1dUCRknS5kSH9phspPztknFgnV8AxtLW3
TcP0Eklc8WCrPL0BgaWNMbYlpLqmtdB0jAWLaZqRpkGiW6GkCCF/tS+hg0RIOoWn
LQjEU92CG3OONvewsDU771beNL+y6ZLOhU1b5x87oAtmyUyQuyIE5a+T1Tnk4Eea
fzJJqTcQwilqX9mx1aiuhQu/SWnqHQg7XriDxScazzA4w3kjvqC7FxVYdjXOPctF
YP+61n7rgPSlCisJAgZsJlQk7RXfHhb0GEJyqcRnlgJhchAdSqXITRj8ePsxzdh+
sqKd5nX+kMWrR46zOJjnYquMKboj2xpO92OnMPtuSVXAj+tKBVKJnMc3K0YHSvvd
q3fgnueHofp/8OxQbNn/gsSCuTz6fqzLI27iDpDszrn7ELJ8AQFxk8c1/EZfztd+
fGk1qLM6XaS4+IMnxNlJIGNKAToqd/pZnKwhd8LQ/UC436cVidxPNHCVYCm2sb0O
nGnjfybxJZ1U5yWASJG++BVvSlyEausU2AYeBGeyQvqopQez4TJB7qdlXW2974uy
rFp1bVpfIWSHTGd0OWoiRPCYIOSFcm2ksYZ6NjsEzF9CwAbUZpCon5aTm33Wih/h
E6bzFc2rt0XjxHJ4npek9k3P8sm5ma6a7K5pOeFzlLfY++6psWm9T9hLiVE13EaD
B0f9pXERxVU2a2WBOsc6yHe7BGawtc0y96fG1eg0PMcsyaYEvlN0dEQxp3iKf5Pn
SNQsqnmMTKA/p2GFy2HzNcj5prLl5+SnUMwZooqXvRb+Y8Uop3KqEEmTL4xpDCxu
M19BsI2NKaJnlo0+xQ250ZsEZ/68R9GMk38oZLUXajMTI9NGZGALXGpGhQZnugcK
1xLIpUlPyTE6oac1vBOIQp5KlXGuBOvIRAzzOBvpzvibuOzQx0i+FUvrHN5XLBcu
iccgLgkdY+a/3sk8ncUuroHPnV6Fli7ymnzUolAS17ARICjKRAHgCJfqhydMfy/q
NYZTHyhGjksfX/72TY0nDYRZxlAn12zCthF8qDzLfhrblLfDv8T4yawLOBEF11t4
HI1NAEch1dFlJgGPfHoTqJzX3ApUu1xzfYIRqZxiaLmoDvwKQcBRhQK7I0HZdtPZ
1vUmlRRkm3r9JMDgoUqQ6mjxJ5kmt9SS4HSb1VOm3IhEDpJM6HuXp2djpoO831BF
Dms56XWWN/S2epcJ9XUWs6rXb34WbI5kZkMxEdQPfazUCGminROERbOgqqeMOcbF
+Y8W10KYtFuL04ymI9kWA79WRPmhsMLcrjKX2T+VkS4WvgT4rWlJAhNzCWCMHbA3
zXbJjgMZl36yuecTbmoCOfehtciRAyN4tSLpbZ/JzinK1tdbQ+99x2GurRyM8lQ/
lJKsTULyQ7haVeEQUvCBskfW2oDUwY6lxYUnw2Le/oj9cG84bpoMf2g7BFC95DYQ
5kpJ4qsfH29LbHdaEJx2G0Q1rujKiLfdefbMkPO3jcqanWhg/Pk0NI9fqJ+6uZHB
3ZvOe5EuK3UlYSxO9KIxepbC9XgNJBdSg5ZWMf4vPgVpxyieB10CNTnkp9+6H/xB
8Ww0G5GjJa4cpNr1uEy4RXeZ0PUy8qlVYrG0/g6lXLmbe6NWTZ9NyS58lx6trC1a
sb7SIFPi4eIK+4wq+FnBkvDMKkEyHQ2CUt4xzSvPv+xtYST8f6C2dxO82pnTpkWn
0SIaYNBn1w4LbAMkI20qeID6Qt5s8p/CH4Xn37gu/+scwMhaqLOfDN3u7cI2N9w9
5z6560rm7mHfKQa+ENuv/5ojzY++rgh561iH6pF+q584KKAAx2Mg/sOboaNh3TmH
MU9Rjl4OeVrUeCmFSMaeARhlOveVbX+JKm5/z9ePKXhsgPDwz7ZlqIFfkw1TJRcL
m9zH0zOoUuREQflamV55JD4JA/YYJ4UXvCuX92eGU8uMFCt2K7jNpoiQK3rjnbZR
+MMNKn71dtYlagWIztV/S5p1Z/F6ZyIMovUpeQzQC4picbOtjrlqaJhJdvs9Vn7X
gjdikgRYjsO+DdUsApm43HU+O/dHEo/fToEA6Ys7IDdX1Z/t23kttnZNPgrx7wtI
hoh3Wu6eair7+eHqp/3WfKPiu+Z6NqnNaoG0VoL+czoks+Lm7KkMxEZnT+xoVwQN
3IHpIttI5LInbaZIEenuT/VGegfBSQWCfdEaDLXudY/qOBDFRnlAZfeF61+MTH1v
lJPcRRFcps4+t/OkgW5zqEuwXVWolParytcpe7RLyHYObhOSbs6x/Vw46zMYUYcb
cLq4u3H5SJDx6mwXaDgt2fyFjU7nbFhLWgZhbb4N+Faimxts9LW5/EvgBEBdvrtn
mHzLiK3Ql9359Bo5Vxf/vwXBa4EWDh7sJw3Q6JU4CF14sy0JOY9KKVpTRo7NHiFt
xvUDP3FqN/UIEH5YG53D3vEzR5S8Waqf6dGmzL9RtAyWvO78PxFyPylMrOOYZs5K
niOpcfVCY2va8FF/+aJ9kaaTJFfLg6pHYSOPKcwpmNAqPaIW2sH7SlAF3Qcbnybf
fSS8CjxLE5opeVMySOl5dYVc3GBWkfJJmirXZgrtggwaY2dFpS7ZolNYvG1Q2Qcz
Xh2oDHaRd6MUC/pY7aa3MsJd72OCNsqWfeSnM2fGMA63j8X1cBow9EvaI13nGdga
nWmgFwVR4VJRyQDcYDOmQ7ja6hCXrdkXC667d3Nnz+XvC+CxuX9bvX4m/7pBjYFD
GC0raEHnZuu7GoslwSvIOobALrEqMbbUog8v4lSugnF8muIacqUj8EPErl7NR5ar
eTGW5JLajoEeEnw8mkWZxKBaHFbfe+vh84SUNWKpkvxMxV5iDHCFLrh8i3en7sAY
OKeBJxJwqE5KByq9DJ0ZDHDf8wG4oUVSUHfJHRXM7H4uk4/iNW7+gD1W4iDf04dF
R6qM5bCGJPRRGGBsXNkCwMc8Rpuobn+wmbrGxlER8eLQHUkBPINCannDprvcxYzX
FMRBJLH94aPjF6vkghjlmEH5AebqwcPmRiP1OhGqOwus9ColBpcpS1/RimEE7koY
Qkca8rzQwLFsc9ZbtPU5TFA/TQLv2oZkiV2UPwBKYsjkAhbEc2/zJq6n9hxH3boB
jX/mAw+jTno/vQA/Oyq9Qg3EoIJOBSv4Us4Fimt8Ojs4Qr5SbKO5rTowvsBE7PHp
Q8Q1Mzo127jZPud0c1UJxRXxFzxYNcRADn7nn42TfDZJ4pmgY5nnp2DFm0CVa50B
6I4z7RjlCc/xyRCz4QFiHThqjv+QJkjvggeHkasxjHY9hoC47PGo86H3YUwlSqRk
BPaY5lYiegx5r8I/sMxyanZm1tCmjSkjzY3eZMOqnqemqpKztyH2gyQMLeuh2yqC
Wjy4SXcHi5Z8n9CbHDcrjcOKYjm+K2Tcm9jNiklvmXCac79xgND8on8Q8CKPS46U
G8RRMEIQTZJsjc4wQet7QcdfOkGXN+4c5cU/4VlRP+23dloYi4plcZTPlJv+/1TJ
VwaB0ox0xWzEqyT8fkr9Rbt1Ry1YdFhF7WjsbTr+V9OPdhn6RsKThNJXaWYxPwWP
fzBE3Ayf8klwdch27SWB52u0vLB2qHNZPD9CYqM9S7nBIbHjlOkSYxXdmE1AY5SV
Bag12WH1GVWdpK35+OZPNfOjR9to39kmKeIeLG4jqVbaePRLbCo2quaxQ81uTpzo
QmhNiIRuts6r73t2WeMcFOWTMWtFGBoFMVm3FV8v7DWqyHM9w5BO5zV9Fz9B6aGG
PXAVPRCBCH0zkCW2cEWpm7ifbd08PJsvRPq35PZVCAQUxYDJwY+oUrNnguCy21y1
Ir4G007G5ir/7X9lUoDjl87TS95RZ/nFMxQ9FdUWLSrWHgEOIf4FQVJ3r7knXf2c
4o7odKHZMNjhVg8tmUNIg8+A+oTrkY0JYB9JXgEGQ15y8v8DL7ovuKbSeZvEjEnU
ZhcCvsqEIRG/EQwSebiXipiCceOIFyxxpRBA3Gn8MZO5gHvGqmKZdzyieeOxx52L
jF1pEU8IKhDow9Y0qpFxTdNCFySR2pwzoY0h+/g4a5vl3e6kPdD3cG+Cnjx82p3T
dNJ3wC+QGFz5FqhEoPIqvxtCuSFMWtX21VFsoJ153JNALru7B8++Jsnll0BtONAR
HFBLhmkNl3q1D5NEQj5TwelThvroqRyc8SwipDReEbjjD7YEEfH1UdBKdQCqb0Xh
j6B8AFI0TcbHJ3BfdTxsug1rP5r6O3J8QFbrwMjzY4OSjWfR4ID3Lgew6GCJZ+71
Wtu3TcckuI10bWJjUCy1+ANzwjgeJIIk59AHdcdkKqkbGZhJyfvk3LYCPbogzZXL
Z6guLpgupntGvXRlcp/RwwHX3Yz8TUEcP5RvLk+Wrw8o0GnnpdFd47bjJpJ1709w
YrGTel5Tc1HCI85NnPF+RyV8eHiZ7D1jJZhdgQTaGzLy696mCwi6mwMe1jxwboDb
wHkJCIWn5pmTisg7yXYoAgBtrCuPMYdS7ZpSdONgIYZyOjnYzt2zAum4Ru+G74eL
wwkPCPrT1bIGomSIJwpALEXBvQjRMA1k1Nx9NjHaR83e9A+eknldc1dWr2MksqsJ
zH69DeDzz77OEKYmjMSlOH04YpGULudGJ2HqKv1UNTDqZomslH8gri0lMRVGE4tm
7otEvG3cjJm72ZjIt7i7jyFHW94ZVdRrfqxiclAhwa61pIxJcJ6MCqtHV8800/4j
bPSSprL8m8EYl4d5D3IG5wnEYpC8Lf0q8Tehlkveu8BrQUmdy9WDd5Mx11S9pVjA
sCn7w9E1Z1UN5sqCsMDghVW3EGXL23uUGYmY9+wlrIfHzQusofalozvvZXTz2mVn
st9GpDaNFiq5HR8cDpQs8wjdc4r4K/XDAuJTDS7qUhzZM5JV/ksSY/cz8Ewh7LBB
szY5qbnXEMA93+gNQEcfvkI8plolP3Tg+D0aknHGfmuTL03aqxRd/8kV2atciqon
l8vOsbOG0U9yb8ZQyI9D41q1WbIBJbOHZSjnwkW7VPE1okeEf0WR+Zb/rbZ99K1i
+Yu0WqkoMauRfZaReoKGrWz0aQq02sXGYdkVI53RMx0wNzOYrT4syZ4HBT38R2Cf
K3JJ9X0xDqxo3atErcHoxZFjw+tZKGlbk4j/RY3nD2+hitNhA4w453CD+ZspP2Pb
1w5krYcRbmIqyUFLK0mpcZJjhC3FUxf/SG+UPplzNaSWqgr13pdeKtzp6eJngIpx
3YitebtKwkVwPlUsm0rA7dY1CYzcZANBrFtrUEqGdsmCPHh9i3pBmrYKazKBtH4a
mVTQ2UuO6hjRYwuh9iy4lvsUKKG3pJHIdK9qxPIuSAuKVCHXqmDxUhFPxqWFYn/d
EljvqNHqwS7huqnu9qrDaAGcMcKthnKjfhtRbfd1cDENK8O9X2kTmXBtXlZS5bvj
N3wUBOgBfocHd0wiToiVfs17j3UKj8zvDudT4Y0Rjm06fhJQuUBaFf22ir3zAUQp
87y0gloZ3k4AflcMIebjePw9TC4mAGVrO3QVi0cgDOAFpDZF8KUJy4CJGFQqKX1w
fpRax+hI02GlXVc4eSE4r9gN37eEi4WEWOY3/4xIKgdqNwOhyyCQR7q53sRsvjw3
w19YbphnEKyhpqHTMwvoIj2oPrdKj9NDYWi/NRep00sBwMWzfRiInBtn2LZViCwZ
GV43U6LKYlEDKnGHfsFsnuBtwBnE4+uk0kWZfPoeF3wMZ/Gp6AKY1xH+Bob02bDv
d+3hBry8JPJCuvtpbtLQzlMN8Qi6j0CfD6qpGdAhu7f2e8gvSP+NyxO9R1AeAURX
B4YdBcUd3DSz5uylNe1ebMYB5wRxXVCKag/LgT+piBo6GJPVd/0+dBxxT47iILGq
TnKwmY3qz1qoZU0VxZ2SXA941cM0aCpogCgxB8yLvRk/QZKEpE5RIHkBitUb19vm
gWWZ0/PQfuYIyk+aVCO/wOZPGFfwQOCy+zrJP78EFZmkv5hF6dVPikg0qW1zWnBX
ujbfD7/GBmvTiQIhv/rEzNBqjsWOlTwJfNAOMPjdjSxkHbUVSVp+aXch9MVRIa8X
lZ1tB5XOJDdSlkwLiuqUkzC00jUO1RaE5S2T8UPALk+KvaM0CEaJc2WiyOKbluhe
VihLSfaPOa6C6//iDyUsP3OnXUcGQQWeefHPxiGs6npRbJdGn+MsYsflX3iplJWA
Imc5gSTf0K0/0beNTHiO19hd13REh5p/t5n9lgS6jnwZx5Cl+vqS42i5z9iTFYAc
9/cUXG2FvCVFaeJZ4dp5hOEO7j0peiygIImehFAI0gavJKOLvMavI33L3inFDmd/
e5/v0RuQMzKxUuyk9IoI13JqyL4GJ4HHwDxhV1hVpXE0Fl37sxwCjgPfnDuF+f15
IeBED0UHhj325Jn3zM7s3YFi9iJ5HUTGHNm7i1wpKh7W5ViGR6OkNJHSWr8lOGhX
x7r4G06axA5anb6VTpb8clesOySqxy+Yokhr683N5MM9NHxL7TvF9v3Il5D9njMx
z5YKNxi8kVddyWYvjYzjcJYTxVjihtz5cyTJBUs6PPNbraL2smCtJPKRUHmGTP/7
F5Y7k+BrbMVYz5XQaMJ5pUj919fFCn2HcRHm8xpscd3raacJaBkpK+5VT8+bNYj7
r1a1bfi4G4XcWawaylweo12wQhglNVLciMgMxfnUrYkBWg5Fc1M4t24PWwaYbGO/
Qk7aA/ligPES7Djz0KxEuCLtVUrPZs/UTYBiqwjA3EFhS8wTKnAEht7xoO3ZBqUR
o7cE8EAtbaqKgyipChI3Fyrfn8Uug+3gr1P8rGhKnpuavuEYfVg/uqSDlUEijTB7
/IJp4hlfPi1MY2pI31/83QgBTC+cgIKwDwXml8e3f9L30BFAy4iNj0UD+R5xN3Wb
cHgGD/h5hhkrpId4rPXWyaDcUtbc8xBKHHnVX9xjakjRoMT9hL5XEHK/mBv9iwiw
8yxh4MpNTBeTgG5XsMMbVdkSpUuqUANbtBXOn57EB2ZD5z3Uvy+z8gyBfip9meSv
XVEJB1ElxiW/zxnoDz7rRjwL9qCNlv3Q8HHSK5l/Z+P2xD/7fMzSgL/BBB8P/vc/
/lWrRkK4BTaSNQ5pSdBD6crLyPFugCgacpHuXdre359uLeOfo0I4BcsOOV6jg1ZI
UZ7WLZEBhuOdAgcfyrkNV7T0fidkVoCJbFGqVI1fwva0QPYB795/Co+5yFlgt3Qj
wZMx/mIWSTHXv4L4EiVCm9bUe+7JU02dcIqH85jWCYQNg1hw8g7/33sSNO7JriAK
tfGgK8dqj+bMS9my//X+MYvi557WE1jaBV2kisF5a3el6ixnfHahIJbAVtDMnBgD
CUvwjzzfS/BJeFOWey3Indr31RdiHCIivIwoAy/Np7Tl4Xh1ePuWpLvzmsuNW/TY
vtZpDdC0xIORetyaDUksN85dcxYwqjQpAYAVkJFHONnKznygVOtxPebmi5O3h6rO
zoJqDB0ZG2e/kIKT2q2r6HetZlctWQslxv7h7PWxSKSkS73GS2MFTGfJqs6KW2Ok
lcs7837OI7OWi1RxMOGeOx8BCprliNGLothcDYrTcpMHuqHqG+HWjjVIs49oAIBF
l/PkxGHDN8jOBAeqB7tbte+kpI7u3Jnar4JhEWybZVCiFQhQ6wRfpVFLHB7tMPHD
KXhbz4j5L6ig9iuA9rknvO8v5/m2ROw64nqj1ZfacBuVU90OMe0D5zYVmJ+/ohN+
rL58gKaP/fUHaGbBXV58IiX0KC9n/DP7aq6UpaCjpgT+lTy8cliunbYL9oV1/wj5
hvQKB2O9hvJXhGOHAKRq74kg4p0578a3SHBwanc6mAP1UPBIP3kIAAXLgB6YqYBO
DEB0zL6CwHRoZ2VZi2eoJQMDxyncnkIYfdhs3XAUOnzVszsAt7gL018JKS+Fw1qU
omeW1SFnduBwdd3it2wMwE4ohcQEaexMRn7b4nuIiOQa1v1x/7GKjqWM+PZoZL7h
C06sl6636phzI8HV25/fp0PfXm6ns6k22y3pCjbt9DUKtvMtAZ20lhuRppwa9aUF
lERqIjSmx92pRmvNDbaLgBIrGhhgrxDZZ9LGM5YJnn7JKc1tBUWPNjOmqg0jw3ci
UzPJ9ndz1xuMqxCXKTOCpnq1mpkoDu8EBiFHcOR3RvdbEthyWF+MPUR8+swE/7ix
e1fIXbqfHnnah7aqKMcwpLOoOfq97wnUKhzusNsOEvfRpe71roqKOrnx4bNvHcfm
46JQCF5+1uayUyqHg1nabp8MB2iZ9DTUfwiW/e/Od1xn9E9LSBqGvkxFuNfZ2YQu
eu3zJ6quh9iTvPDU1nXYCg7UbnFs0eZ+1qmuN39jv+rT+WAjpfpt+YIJXgt6XRUy
ah29z2VL5yGDQKfj38JKc/A6LIHhOI445qEu8lRDVfVbR3P6FjEhfpHGo6hW++9F
BVFY1+mxc1+9zZn2FTSmOdhUV+lTJ5x9T26sE6P1gIsV1zlmR2nvlgGiuDcvd2ht
LQxZeOtu/2jNIAKXiVW0b8lmlPc+H/L4waSOdtggsb86SU1EoluLSaSREUOKySD4
CZXCOGkk8DdfoVoDTkgjh7tX4PO6gYeijEIQCj4F6GHYHDwqry5Ws8lhbn8e10dw
Pqrk31XkkNdl8j/JJWPBwGHi/GzAb1NdqzNmFpz2Omfpu28vSIhGkwqFMh9ErDlP
Ynfbb93o0whGFj6DUINaIUsueTJDm8WlYWviGkSfZgk4s5QikToYRFz4ngVwhAqK
fk+WOddwhyAgKMaNqA6empFzym1j6n8EtFh0N9089FwhSiwh5jDasgIrXvaIhzWO
DF5RHWPCvC/XEeHs0730KwFgoiMKIt3MxqQira1eyHKD4JTvoPs6UUCCOFj7n10K
ju86pBpZTUm1f9IikasjqdUYuV2dioztqS4XAVtsiRBbflVMtN/++kGeGbk1WQto
wLd+ljEMKGaZkFDCwYtRVs/vcFsLXdHtLYHZEwYv5zHQ5AE0jog39rtRTn2UO6fe
uC9QdbUYv+46nnaummvJOZbJjkpLzTfVseLbcQXFZOTtt4d+xdzzQ7I6bNpYya1Y
3DazNbJJdkfG9DE8yXNhjQ9gmApbTAJT+1pC6ZGHE9w7XjBclN8C9DbKRNUMonrr
4r5se5Sk32YVQ6bPg5y3rjSZFk+fWRy74AhJ2LtG76/wLQ6/Jd0pecNCs1V7XfhL
oHC91PVF3TWx7/hHNG3s6PBwSwjdvP1fGxVWKdeNcceH+r1OdY4d290gaAsCvnxe
08yaT7uhw7RYmQou1rpMJ1txzjQx7fo31gLNBC82etwzEo153H5qyMSgVgM97tMs
YMP5AQoUK/kkZGlKa72eDUAedBltWCs4eb7s71WTW7Jp2NHPKeCWxIzoDcD1R6C4
NShMglrnem0ys9rPclZ3Ch19pMUw2d8GBx7Xl3DvebMCA1R4wTKQh7zzlon0IdhA
K8rC/dOXWsr8k+R1hFawiy8MToa5r24vcG/3R7z63sCkQ4u2s4WcxoXgGmNUmG8P
uj80S/3N8Z0YQJ/nvqYxcu7hgUjnmBLtotugovVuTRCaHjA/ZesqjF08z99l2hl+
7ghfQbsLwnKn6Rs6J22FxRFp3PgmLCWkv0wfjTzQFstPzyFrjaTkhmDKigsUgv+8
7hP0Zcqd48es2H9aQj9JR6hbRGjwbhT4g8QVtJkGqVN/09et4SQxRBmaGav4Q8z+
dD1VSIUesboClmyyKCqhTYwcnh98ypFCM0XnbYj/k7OlPe7zOOLse4E+iC5gAsAI
556lpC3PNis7zbMOkL/D9W3It2a9vVCk4PQ33ByqZRQwAhwhrMAphJ6aeAGs5NP6
kc7BId19AlH3j9V7S6uS9BPDz6KGtJt3fUQZ+CQQkVVk0qoJ1/mUFbGS0j615cgU
HSS71z9Tb9hjcmDBTYHHvmzRvU3L2Nt+PhRVFjkySyMjvPVtXuHd8FaLxUiGkBj+
9Z46EOHdoacRJrxty4nrdO57IR3gBsNlFtaXgeDjWJA7emSFJwz69TM427xRGy4Y
VV0x6DS4LP0bAVzFrGCERFbpyDWU8WY50C2RNNF5K8mWblAZSQMIZrD0wl+/IFGY
iW6CPVw0aRbjEJFzXA0+SFus07k7wTyKSEeVxmZI+hNj189b6YnP73OASrskD0JE
V9VSYipjL5pIRJ+yh7n5mGBgZQcly6b3uzeeP+BML4JlTxFI4Z6+BvoonWkLcnuG
2TlNjmCgiRA6OgtRN25C1LZUfxI1QwVwLm7Cw/IDSFqqeAp7LZAj3f2noqq0z4rc
lQmJmQ3tvVXy5xQLEHwbKCaUfmTjUx8hZjK5FQDEnJSvzRETqA+ZvZ3NvYHgPGIs
pRxqOwTPgk107WqRwMl0/sZ3n2MNt6wplR8A2o0AUdtZKqRUO6UL1M6vngpV/4yu
QM3Co+cRKJSIhZx8stfsBXtPUPlKqChVoNnCOWDaOl3BH/qeFLBm8+bSTDgbDZkS
0thtiNSYtvFswZd4/AYbibFUh/eLpS147klqsWoVeoaa+Dty8E9VngVhwxaFxj9g
hj4wyd9PyHDxftWKEaoIM9F42QcGcG1kheLqCTuMnX+PiKbWA5a7YB1lYKTkxVBN
pF/eu6EshI1q319raZgrRnlnt2zvkASSHb9aepe1qnaBs1HGnCv0T307gLwBUTzq
rNzcjuaLzCH1jbQC1pE9kAWsWdZT62UJfWHNpmY3lXnswg3GaRTAU7twy7PBsTmL
G2hRQw7ilTm906EF4glSWFINUvBJoK0PEDyyZ86SuaMEWuJgMZzKcqtb21qy+we/
+SGiB/K4gLG5UbgEhE+KQIKFboY/WNd+Iabl9+RJun7H8e+PLREQINfuc3SKrZxX
QB6fmWY706XeRiwe1yis6RYQ9387dn570NhmD5nc3ziNelj2YWYGoOKGaW7T4RkU
Ay6bM6x4LFdie2i5MihfatuVA32BD3IETK39MEqB8TGiyiVLFp3Ksfj39D6nQ3nJ
jdhM7tm/NUhwFSD68r2lCnw+1uaOC20Sxs7U2gOEZ+9AUIKnqxY5w5K/zlMBsHDf
19lbN8JesDmSBcAjjCfBnufmV9xSE6WCy8qBRrwNqoqa0fgeljl+gT/Gpiu8+w+y
akd7uj7FdDipgzCOMDjB2TGdKFoRLHm2Jb0QnJtXatqkMe7GHJeehhKxsGvsXx3A
Olka1Faj/MIpqGJxP3lRhomhzA06BYX9uynzUnoAtJ6D59LoLdTZY4/fFGAfkEBk
xBHTGKLWWBx3l0/WYzSy5/+BXn79Ry5In7gkF33AO4tLDtdCN3flhamZKKGsrS8V
7jTylUD7Y4xURTAckT1tAXf13dThs5P7M3/3A9gdAfhP+ThpZuf4J4WsJI5a0/uI
Trx8/YfXNRpz8G2ZakGPjXAMI2tleZnSqM8fX6PY9R20s8DUTAP58acrBdHI0x9t
SxQmKAdGT8zWZWqC9ZacukdEp87Mc5eK2AhBnjgbsS1H7GfZ6ahfu4HAzCev+yMs
e/eFzm7mOQjLTg2iVNHbefGsfDO8xLxX1qAfQmDksDUiBlA+563YQUpwoxc/nuty
Zr1lW1V2Lt1hpyB8Iy1eJBh+X1OxKswTuEmGaTqaWNQvuE+qtRMrBVUdosIb7gEd
hNz+pXC3OundCrjeKOX6PDYWzB7peXq1FPg28E5rQXXBGnI0XkqRrwwHKkfMO+3j
asKcHWy73xNgiXwWs+A5sziMUzf6FOQXKSdyFuyHNhQSzvuWeo8X953VboRW9deI
jqlajMefcov7x31iDjnRacxsTG0Rq5C7sELGYzlmNG8ISbRBW9/Mtht57Pw3pukW
yMebOQFQp9fftcUHMa6XPaEbWINKwVTMIlZi6iIRwA7I99htvZnZieTaRzrSOoPl
lXwWlMlX8xx9cP+nCRlHdJlGC28tv0xRst3vHiIfgOog2zDKcrxo1UYevNMvCzZ3
nfurm3PCfgqL51fzn4btQCN7Y1ehhInMlFZMkIU55RzcTLKanVq6/T162dZIO44I
q3WR0+FSpkbTJTqX0LHGV+/vwKGI2O1wT4JptpVQz4t0hXzc/y3+LpSDDf9M9zUI
UoM9MhiRqV/jndUulepARE12P0iPEbPoT6rcX0kFu8yim13lpTejAs/sSUewlIox
+fmL8Qdqf4t6fA/1sm+IcFgyDcvgyXkJtKS9FeM3rw2P2he20EgF3LbSzwsNfFCq
YNG19lXKCRHxHmD2ffSmjZnUhC/oGTrLc579/9bOVbmDClUOhS0aolmVqXBi1Nsd
lMqNKgy6cfAVMmAnH8NH8svMm88jAFFMjhVDoZJXT1Cx7nPBOODFf9zLCdG3A2s5
GiTernel9oq3dq855wvn9LLV/bMGVza7eIKxgzW2b8ectuAwjIzBqQKlpO2k01q+
nnLclIitcO/AtS+/C+ejUYylUlLzMVmf+GmcwieOwHqbH2kESiOe/Ab3er+g0wb5
MWi7f6RXd/t+/yzqPUv++NqGwwVyVgIDd1qYZMeIb/o6rFhd1IQq8aDMNc9EAT5p
w5EGKuhoGjCv3WfoW9qkNifKSxdqeADrsegaoKc2j3Na7EI3aC00oI0xh2F2tb3o
ua0gpwkwo/6UGoflajGbW18WQ0C7LDi8uDgsgntyWlDiTum5fJvVckxQ7SezARG7
+36FR7/QOedRiM+O+63ps8SvyQ8HdKkNvlfjayd9jMdnHfuHsUJdZ1oPicchyEdL
3XTY6XpnKHxa1TcZj1auIWh9nwtK+OFJoqUuuDJvCPdrk78WUjlH6fo9SWswWAUa
q/E04XQZdIwo1NnLUznDwmYcwm6Suk5NAZg3dCuehKOVvKPb0EulQ+4y7sIAQXfV
NZHYktQjo1jA4n2Z+7KajF0m0xF55iMthAJbiXW37X6pRnNLXccJRL+dzE4HmSsI
jbniF8EpfLevtMfNnKlWf9Sn6oY0XeCA+Q1qkO+vSw205tKU2HvmoEhWwTCAcCBj
PNDSd0CHypDEehRdtMPEqt+Ys0KXAhm66CN5oBCNXDqQoBwqysqw7QdgLoHthLh9
LEmAXk/oudbVGXXIdFd2IeGYxWWi1Nn30+rcytdxen5H7Vlx3TaoHFgeWTo/NAPh
JOXHFBH5HcVd+w/7Wdipc6QpX/VuN01Q+HfdhoKqbO0ReDanHTp4msclyJtbPzFw
OFxwAkBD9Kqluvw47XcBte6HOqP37T88H4PEUiah2Kqd/5mBGL1su7uAKFH7OMdg
59Qql+hG5Mr15142ovAcSZPAP6am95khpLZYOk0mTB2XEX25+pSI2y9gjFryDHUZ
1a8oUXpwgP+OiQBoxJnY0AvyTpNqo41WrnE/nGsm7N+AYbcZlXqbCN24QbVek6g1
p7DQHQiBIl5F+2UJohIyrGHtycbrTNoJa6SLaCCS6GlAjwAyhGSHjXYuZyQNmgkx
HyEPhCl2j7W+TKDIhJpCHArWGKGuwXs7VCJxvBmP5XiCu9SGVBaSM4TygSjnebso
hjQoId7LJX4OroZnZaYB0nN7lmd1tClju7NgVGTfWCQ+s9FrUYNVB++NZZT8hXRl
/v0bf9dRLlQvTcmu9De9SyKZdQuM0JZJHG/0y5ewoea/RB3l9hR371niuLzVGlYZ
J9Go3RIuQiWobdpcBj+UMM5s4PSF7RIkSpq0qAdXJh4OvsuTEfNiafVfG/wSbfCA
WYs7ldSji5b1O1TuGm4lsON/XcfHTvQqr69MrlYLCv/dA2GfX8jGZoMBRzjGNXtx
zFBAtnG5oMyT6q6K8FHUAPobMFlVlQGpNF4jHJA7be3FBeWVbgGA/2m0UWtlu4+f
44m/ePfRF9gkMWRiXfL2+iJR+lrcMQJii57zWmSH6NLA+LfteNsCe8t5p1Xgm75F
13uzfDu1miRLCwafj0N0NS7aIMQy03KKPu+et6IG511kfgGuIwnWJJ7VdKgW1xnY
8m2iAS6gDCycff/b56JaB3Vi57znS9eZzMhewwULDCFofql9NzduIxFThcvjcYAM
RFHcDu1YRkYHRrL4L7UolEeOdZxCo/r/QNddDRjP6HLmKUyS2AHAh1Lb3kAdpeSu
DiJRTy2K1A9LLEzveX0YprP0SD62ZkBLy5NnPDgndTkaKdSZO493dZkYke+KZYg/
vZb038ZNUIBn6teUm8aa44an9r4UwZQZArT/NBRLvn4Cl4gjhp6tJZVhOl2+e2bo
oV7T1M29Twkl3iwnvkEBbLVBeSMFGDKuKH7F9H+ibPbQGZlgBvx9J6lkyYehGR7d
Qtds+GsuW18AFFJqbsqetcHePJO8Zux+Z/1eVCVUX/2KCiM+aHyPOhXvgzmEHErS
q6jKAhnZIfggL8asUkoRm0PBxU+0aXeygzXuTEXvbqDu5IFw2s0+bCtVni54o46B
1FDqcRkJq8PaE7wk3VcMxaBOQ24T6gY1Mdra9fUBUVaKA+U+zckY7bE3EHMp1mg4
soJD4QiAqo1IDFX9cJob3qVYFA3uVWtcfs7l7Uu3XvqPGdnRJaZOgEYtehlBVXuF
wDyqKDlT5hb4AMe2D0iEd0jxb0eyskRhi8iiIx4Ye0sRCdcMS2K1WiUK5Rxti5Jw
Aym9JXHsgNwjouKh0OxvBiM91++/cVhXxlg81bbck3rqCTXES0BSSdHHnRcK2gUS
dO2oCtXlG6Mzq4tNLbAKvfHkHuCjdbZKRALVucCk7/E9sEj7d2UIavbF/ldm6g22
jAI/Eymk2swn7ia2QItAb2dxq1YhGT8EcmTyll4pggKM+B9h0koapqYDVGhKnN/F
hXjFKWJk/ZOI5IPLOpQ4+UaY7a8pZISTjpmFiQ0R3j3NRPdhidNmIL5yVe5b7vbO
lLkxidjFJehd1wLIsAVuaejFte8gAf+B2lI1cHKfal3PEa0XI1dA8mF8zPoHVZw6
ycqpaEylg3Kp13oAIMdHKW5BGvXFEzCRzW79ddoOz6SZpLOduVxGj7shLDE/YUqy
Kp7sb9UWQnj/txZ8Zt/8AwKOIYOFS1FAk9Ak1X3IiqK0A0Mi1JcHFgCGIYs9bVxq
qHlgdsGHFwCRZ80dlTBc93AZmbrx+ZR8FHYZM0OtQw4+8quFM4u3+gOtnJkcIFlf
UPk3+f1FXuhjTk4AjGpJe6f3igAQxfkP0gNlPx4eDy3YYFXMT2Vw3PU0Sh120Oti
310vtgXJjQVVhicu8w6qS2JZYLRXCSGsXYLtMpZU8JWaqwGvFwM6v4xK7QGNBuxG
HP6aSyYGaTXsqm2xN3RHbwUNosyau/YOZsjcXLu2s1ezFZw4ViEoEg7FJrtC6nOD
knNm0x87AnHeWiJAk5ZdDOjRU4Z1rPMqhfod4zrcqGeLbwnQXBiNAL2zvBdqMnZQ
m6YnqVl+MSONdcgGX6XkH4uSKzhYVGf9rSsY+R6M2IJS8FN2RNCiusMn36AktPCm
lg0ZvKgaVyJrfh7qXGu5Rif40mNXzRhGk7CA4Ml3NSCC6h/ymMLmK5Vm6L+mo3cx
IIMAFcOFiHX5EyQtgPVUDx9GIK0TtkWkiJhsT8H55ItDOj6Mr87WF/QUJphhpbXE
G22kRsRimLYhmz/W4Hgc/N44HxPV0SvUd96sizXuO1S3p7UU+OPUXXRKlPKYGASM
FqjmrhAMvImg4UU0ItAY4Y9bu3CB8VO4eRMKK+EkGBdHXQrN40Et2i4bX7GWh/f0
aBR4JtuoB9YPfNXBQ91+RquVQOd1FXf5/m7mdqTWAK7Ng3ae2jWRc/v2l9+RDWp0
zCXGspz2r5LxI8ffw4dhE+X4X5zwi3423NCVjLsZ8b9ch8OXO7dxBFmflk25/067
TygLlKZl5R1s5/M4CqUFHOBhTnHZH4lyQHXexCvOhQfbbs0nf2ea62bywp42p+O8
6rcoX3GT4l5B/jGSEo/htFwTneLOkuXhEKQrwsv55Y1rpPulToxNfm2s+Bx3dRaT
TSWQQ6FmtcKczxbdX2aToFCHsnTiVwtjOX/uiEVSdcZRGtuKFd80B7dpqP9wx6ov
3OvCYlKY/3qgRhNvH/Pc0a6rm8o6JTt0FVFGk/K20Do/43Ut2e82XwTY3uKt0LYf
bYV3nyBjZMIRvmEoSy6yz1SsBJ9TphB2d7SfREZkWTZlV3K6RMoVNU8HI7QbsJXM
kcThGBq9EmsNzYW2oTrvZpmOmhcBX2pleHvdUPxKcesJEo7C+4YDETZyyyb1oSii
NqizfHPXJUyG8z+rSVkCGj/5PIj+tIR5tuqlt/z/vwSmxRIxThp1KgPZAHyJTDGO
H9cjeMC0aL1Y3GxM+UCDfNQ5upHrbOjK8Tx6a3Sk6Myqz5tuymB8KOn7pacnaSJ2
rlSIVWo2Pt150d+lC9nafOEReAL9bUwkBf9MiLcV1RkU9ZOh8AxoUihd3NqNiEr4
8o9AztjCWltGGjl3Ro20jfX6WCmYA9sMCkzoPYtfxBWc+8dYozNW/Js2qXbcppmW
ItuRG1f7CgLRtgLLsanwuM1i6HUvFoOU7YaM3Px27+3JhToZa1TYgh3U+qE+kMnk
YxK27phJobfu15/kfzJuNyxHZgk4AbsDvHiyqarH9kCRFOBamOVjavybZFerAKm4
OwiWV1gq5HEgriTtuLeKuZbEgjsGysNTNb7yNXUr8uPvXj0yUgwNfQOug7fO/TCt
o8MjTuPvX2TTPjc+hGaZkoDxLuJ6jvOslSKR/eYuDfDNazN3Np26PVedna/kHVQb
ff4+IMa1IZCD755G/S1599X/+mx2hLbAhZaJgnM0CsTLkeQq2kCfLqFSU19U7wC+
056dTZPw+2QBAennIGU0kj+OejO+F2hx6ymYdihCMmkItDXZkSNl4lgZ5qY3p/qK
aQc+dbHjM3AexgIFPRY+5IYgP4m/QabV0xg1OMN9LnYtqOtku1fj+mnoBt4FlIAw
BGnSENAQYDZane0v5/XOAgEBh+wuluB5uuNGHdx8IJ/iC1QcgQMYMITPOAik9zGr
/wd+A1F9TrCuHii4N+Yt0telz5QaAnEl3VZihMb/sAjmQGANgH0Rf1b+z9iLCY/X
dDCDLXGsgOK311KnWzYVEFppasqxkzInNLdN8tOqTWtk8mcPki6spLxJNoKbQiTm
bhLWaaU2oYURg3sKjaEGwmgzRSloh3EnIJFIgVrxK0WQBLL32keugVeVGVRUHmfg
RW3RGluB5zBh139vnUnpLEaEwbEMSIwZkokA6k4pupTOLQZzAv7chNsMaWojUdFT
BVNiuy1denG9AJJZae/qlqw8GrTQ5HnUTTaKJU2TfStl4AbCK9u2pcq4tsa5mcTL
uWkVPLzxkE03m0OBXNMQPjir5Rx3KODXl2fq4319LTeTSH1FWDvZb/E2AbF/MGAm
4O+4ZwwmjMnI+FZKAdAdF8UwV2E1VuAbkBtNOxHYPhLQxbKr87e1VSh9t65shKzz
bY13vIBdTLJS1Qy94V15/PN+RyC3EC5tnkRQgDV3F39/Esh+FZtH8P1hvZ9M6tbQ
yQGoMCcW9QWyPnrgxP3NICBYwH0atDdcJqbAlPMlUpMkHVeXHT5xq11Ij8WWUR1x
ITSYw+v/FjLNchwMTTfF0sBGxVk2j0YP4BkJipFEs1wej/eWgo2ODMWzk8WkeBfa
pGvZkrB5OCdp/9ZjNztgkKrfHwCl1zM+ns65BRZuL/vCU6/4fn+G9zGXBNE0XkJY
jfZf0j8u0KinWL1I7vCBc8TK59ygpx9s2DAcwxmKVSu3H1M3XUkxZmy3y/yUzeL0
Jo3l0rWhTgtCyA+PN4+bVSCazHSz82ZTb0ZoqxiyZaPJ3M7pwDRF1zx/XXfhrdIW
pWNdzYRZSCgPdLY7zeot1wL1TbBHGF1WmsmMGuCiQaVXgW7HhSrO7BUWan8t8Y3J
9sOB8idauIcJxSozzW60nrHdflHKazxKmkSnK9URaSRlXX2Z1GtQcywi1q0PX4LZ
HwMJztQsdNQpWvwQtOovYCetH75Uq2vlTQXJTked2VEhye5mkEb1vEDL4AWTY2EJ
mjUCqq/O8IuqGdZ9mR3SQXMmbyKdpymSfViYKlPWJMjCPh49EfH2uoVnxHU5thP1
CARLZ1Yqz6TAmu3IUYxmXble4DpzyfYNq/oIGUNjKybyZ7RpMTQRYhiy06hz3+lf
m2pcRWU5OeLlKg9VQdVOEuHth8BGO5z1tXg2HmCwql5bgPkVVvFzdJT8oBE9udT5
rsE9RXI1j0NvpGFiWn2cc4QFP6tYCho3Z23sXiQ7bNg8DJIvSwzUfyDgNHCMrvy4
jMUd/PSkVAKtEGb5XshQ2ZdAfRWYxW5YGqa6/0GV1uxlq/F/lEg2PjcoFi70eyES
QYCUJXDAoRQft9AUxFL/jPrqgO7WeBvmze8PduL4bCtiFqenZYooeop6r8zr1WJ7
P6Zg4oA2HOwx3WwLzYTK3zGcxDNueErK05sy7Vktnk5tc/EL18Dg/3hh9oW5FS6+
BxY/DgMx+MXTthno7ZnRxuEMZ4acu0gFPvSRi+/7eBiRhmIxxSUYCBW+E1qfT5r3
uMfytMCnLHVMJC+aBrAkPrlbw5ZmJNB2QAtDyVEXY/AFVZtWtzIZPdUvUHBD5msx
aoFGVDbs55DP4YWnGjNGvK9P37257SlDz41TBx+joB96T8u99rCASqKbu81iy482
NTZ5Kp2Ek2OBOMfmpYQl3q5BTdE5ITM4ePesQw6Dzkaoae7bRhNmvw9DBNCvRTf1
Hi6DxzklgsNPEhcBc2HheNOkK+PUwvnA8ChtTy1c3Tr39U4bE37N9eLY+ozmml3W
bBWq7ZS4msogVJuNJdPqP5fP9g4fPrdr2zFzcUWIFhoTOOa+xtQF7X1AhSw0CWtR
DY3UfSJGCmSy8ln2FPzpN27sVzsAIG/xefytmGXN/d//xEZDQOunLynmzEc1aeo1
WnkfhQFNAk4l2ZMpQtfnmDooVhaHTYX/g+oEeSBaRAR/yHHj0IsCGOAKzyz1NQt/
7GdW2J0iO5DeG0SCvvgk0UMSkNWkgeiY1HBG1F0N7bCjeID/ka0eVUy4bIdikutz
TunCs2aIDPRsn3EHG4w9jMtxZaxCRCLKFukH7RHiQme/vMhSr3/O7UbYT5k55wVT
JA9KHTRqbur7rQCcIQV+97QREX5KNvrH+MZ1CLgG8848tiaiGqBTqej5Gq+nJSBX
xTJlzpXeJhqU5PpHX9jTq7LbWXTB4vcQBE5sodcVs0sVj0U9AlQsJqjCgvsC2J7G
ayxlXvq+1KYQ/pAM8NOm8uquJZ9T/4AQpkeQeI29GmXSfynPp/LPgWk/1z8PYEu1
LVSm1xbyD9G5uHTrvCEt4QTdGhNI3WkwaoHRNIB2vr/AoxYdT53rNrk0jJGAT/mK
VhcI9q+9WfmA8OwYxD6GkKL0X2atYJ2H6cE6wD0Lz700LVtvkNGbNV2WYUveA1Fv
h9drWTgf4CjsaPea7+EAXd0ImWXqqwqqe8EUKKJ4H4MIUOw9SaWwTwwYA/HrrZD6
h3GRSSbCS0UqfwD7e72k4XxI5JdYzbPUl5JDgtW9DcucANsEpe1fn3Ydy4UF61gz
h/26mx48UQ8tPCRS0aOsULA0B6W3gvyX2yOwzxuya8gu4EPTTrpLPE5UJMBXumxv
MMGhqtk0c0lof1oMFMb28f63hLqB5YWFSlitDrMHfNEV1B5IsLabe5L0DeMWr4xR
FxeSG5x38ZlNqdSSp/40o2jHmrWmBrGeE/IIlVP5dIYHnKZ+34KpDWPRXF0MC3w5
MQg6Mpdetq3lPpINtRnnHIxMTn7TUvVIFnD5KFhiG4NIF5ubIf6iMdbvD6fMq8GP
ZZz2YoxO3oWvlBNzbZn0TGwXyvBIDB1vaThVJswmnMcaB+Z5mymbfcqnqszTFUW9
IhcdBtdZHEbp1S1B42C5O7LoDmoCphFua1VLrJCZqzvT12Zv5AdGdxbPYvqOFpzG
9AJExCmyopsT0WmeMq0DfXJfZpSPLpW8y9m7xluDR4YPe040i5tmDdy2kJd5FQ2T
lwrqycjcV177BFyE9mUZM40gmF+0+OdvAMR4AQBLnw/EP/VJTS7btM7NyXitFkFD
U7fMPw9g8dN6YzAwWooHDPXiQZ1TVeObqxcXw6XWJdwSTgOHtBx6rr0asUI3v40S
dNf5XU1GNya5Ma++qtTyOTwhbxEiqg8P9m7jb75JEznavXPcJHDP5PTP+Fe5MBTN
iDsESCVDvFCV/FuWliHSg4YBTTnavvmuqO1T74DqC2keCckyhS05ufyJ0D3A2bUI
LZcW+m7WY6RvUR+XWrvSnWWR86mUJfhKdT9HI5Uyv9EvH2DeuArKh4FLllFAJXVs
IzYPV7eV/4S5SZJLsCk8qq1DftWMhj81vTNNAcWm4WOGCquY3NWxT+BhKF77tbWa
tIGIKjm/TIhO3LvfZVvuwVmZBlQA9VmLgJF25pESloHpOsllVNZkdVg3mmzPQ91m
2qZX9Pa5Rw403i2+UUFahfl/VDk2hwkcZVGicA2R4eJXJcn1dX7drDA6X5ijNCOh
tQ7W7rR8C8vP4Tm/jq/SWSdoNZzTHznGWGCiWp8JHVYgNh3nyez79g5zNlWXRvwi
4EnlrIMtagQmpnB5/dKjvQsJ7VDPcXQ7iI7gIG03L5oWjSJwkSRDWsUB8rcmg/u7
2mIBy38AySQaM/99NK+7XAenR2K2lfB7+JIcqkmpYjoYvp2Bxf2smOPaxsg19Cdc
mz3JriGw41HOg8Rp9lgMZMVdM1A3kecMcl5+KrLY7yHQ5W2qOh0B7iFECFL8rTmV
obxAcQUOoVW30UGPzY8FCyDD4EAgTZTh+YYotu905bm1/L0XSuOAbyn5xEH3d7A2
ob3+30vF8JVGtSYTsb2un5X4sfUfTmfjuuXpUSXmj66XDaGch2t12Sztu2jMCi/6
Ma2YqQTMSEcyjVfqmnsR/iOS2w3NdvaSXwdj8ssQC9PzjkW59zPh3YO2rcL96cHZ
VY2IWyNut0Gy4R6kb6SA7+7m0T0AzSuNhZLepMOBrtDxlL7+B4Y6EwUKn0yzh+si
bduBVeq+7Tyf2dCQBvm1Svyn7LHTcm6y383qb/nzbkYrAwVK/dazDrEGV1lWJi1D
ofw+HGQbVgrhDJTsPchXt2HrnJgnMR2VlU6X2KBipeLBYrWW927JCGabzFUzhrix
PykOyhiFfELaVEefZB5rYnvGzZyZgk4UoSd5g9juB4efR6w1AM8teX509xZ5Ba96
bCPjBMLtya0RZupooLmJLqT+T6z4vBtHaENRKn/Aked/UohvJwG2URpR/i4EFzcY
wKws7UPYnrgTprgNyBKJxIa1nw7dcgBGu1p7+nZNdPFB8AByjuf71PNfEJvdGtL5
z3uNI1nnVArSfZl5ObFHXdRSt8GNkjGla7+K6Qb5f//qh7Qt8/acyyPfgGmAjdOG
Fef9Q+9IdGO3jUzOSh4P57xgF+zpUQrLYCFiE02aM3ic+XlJuGX8IufA6W1s4tr9
cPcg5HIMdaBMvMiIQvYE8LwDAwjPvMU7reEHtAceBdKgSoHy8YbRH4BlzHyMZcp0
iJ3U8U5gnxUlNgijAzxBbfEXSpAiH8wRaw5VfqSvZiqzGVDD73Q7P379W8SM7fV+
DZegCRzaUM/ymok42EquY8bCdEMxkbOeIzb9+zmFzX2k5cY4dbhLpI92C31e0G8C
2Vf33E9V3M0IN6nYVBP1F8Of0OYSBzjqOvjLTR0WH4aIXbdZlQvj3K2Sh6/sKp9o
4vy2ogjD0GMhIdcwBPIzqr+vlbQUrzprMjTZgZMEg5/oOWxq+cKDBDRjq8uQ6vg1
FfgXqHwNb54NefbVDHcc4htplVOnqmhopf4vJS86y2nuZrH0VNqcey6VzZYYM4V5
pf/yOqF9x3VfxCB5FGErNBDSBKZlGYNcA1QP5MpVO/pjFn9NlLkIK23Dxz1Nq4CF
m4Krh9z4ppRaZhjgWPGL5JMoFKqIK3JJF/4+d6gCo6Fj68cc4iSgnXYDGAgKn6Ir
z/SrKbhAuxicRKUuxjcEfMVXw8K+axOs+auwxo1yU1Amhcv9CVN7DEZfHiXihrDO
uooZM1Q9Ep7/A/GnHfnqLmjRqwCdw8oYQfu2spKsp7sphk1zPzD5qocRwB3mrPUI
9R28W2KNHWPc4jv4yjdbjic5gG8VaMiV5b/slGuhqE7M6TKrWGCFFWOQRezHPLhl
ezH5vWuwqAwYX+iZkFAUJd95663ckWhcXrxUCh91DkKA0aGB63BmzftYP4d3NAPi
PaFcUWjx2Lh4K7gH/z7qyf1s9I6vq/4okov97gyiF9OXG+PvkNfEKZUGloMuuycN
MBOv2Hu5CbbAIxN6BPDgGspweLmVaAtYSou9VnY8NKXAWFdyHASAcjwrRrp1N9z6
+7x4cfNnmPYH7MbSo143bBIuBifuGTkXsDLIMJzgU1fFnBLrkBvZ97DMHfKtVPXF
eqrrCT3IAfRtumZm6tkGvTpN3jQPUh7UubAs197cVVgODQtbZHd7WPeMmyJA+4p6
5rDCcMX98CcuPAQ42EK3/PCaylJxbTpQJuAUFuCvQVUNzslullwViBlGNqjxdlsA
3QaF+FB0blL2pLP2B3vlwJgq6zdZtLpMGZ+9eWbFLqpxqZw/M8KPZtgMXHEnxFHP
qWN6E+/KGd7YqSB92BjEmGuf37q86JvKzElTy6vg4iQ+g+uzRi+xB1TD3fxelpVE
wWelSIV6kosw3ypEId7NtpgNaIplTFV0lDP1LUWbyzYyvThCQx4sasL/qD0E4cuK
FuJVkYt6dq4CcumZ0IZdetoiM9oQecgZF1TkkunAQZQijuSfZ1S6e59URn1TZVkl
wcDO6KsclP43OTUKRcrqvvxanIidJ9KOi4fsk3pJPNO0tqWGQsIONY+enwmRwdUT
64YuCAJ8w/jyfIgZMsi/EP6XRMwg9dUccBrAXMW818S7PkUEMgoex/XZ5vx+l8Zj
8koIC/GP/UOVqu5CvSUzOi70GJ7PMikR0Vd/7FjPOCepg8jKPleJfAUi6ayjEbAj
xXUEGe2Tt2L+3yeRWI8zsVEBPB0Qgps50i5r3M/OBcE3BuxDy09OpOHwXRiyb5VP
88qi6SG8YOAJ22aKDP7Yz4CdZMI5pCjZldvu5i1Vog95nuxXbaX3y3yNvB06iWi5
tVfxGGpnSfO2kvpFDIDBo5J39h0f/XFDA7ZvT9yt9GuYMax4UQpd4evPnWZ6mbRg
HARNrq1df6J8uZ1fXJ/j/YVgl+LxJWV9Y59oPYlwm+HsH9UjTwa+yHqAalppcZOe
CgAHWLljpJJvJy31prwAKVWWBHOBGdQinc/XKCxJsPGOi1W/aCTseepT7AYiMbUp
k4zfxabuzTNrIjUG42EX8UcRDIv0LgKaV2q6Iy9/Jy57Hysz9Mpu3WFiv6nsokKa
M9gJdUEgrUNhq2/K7VPKAxnDXYDZAujmV8fIkgv/t83yHMxHD5EOwrflokgabOOH
GzTHW26089WCDy4/vlz36cu9terC6nDHRy4+fPr4YuxFV5PnoG9xdCn2PX9WE1r6
ku3YLp+rfqGFyT5B2OHa7BIWxvpzSOUFDl0WhjQTwOQApMJ3bCC3cTLBbsxD4zqM
cqAmx0JWMwgZ0EivoBPZVxzGCnffI4/WUlXM5Ni6HDXqGelw3wCJwwbxWJBW6Mjp
yt0GtgbpHvJvm4tHyoyzG65lq5qsr3LnzJuP2XAmk5dBof2Y2kpNFKqF2pBjKYA1
RwFy486tVodjcb5zwdnHD4cgKnGh1olmkWwVr1WyvSuk3QRKahwm600danf8Siyy
lJ+h62mUTznPXrUozEUv7pX9xHK8SAmO4mtrmW1GnQsQT3hcDPn+k5v4kkOB7P+E
N0R0hrgAPv4JNpeqGyIrNaN+Lweaas+n/4Z2xK5pV5mkbQN0j64R8S3jI1tUW0Aj
2lhXPf0Ezc7kuMeNIliwsKmFmoih73iGbRPXK8JJggNDPrmoydn9wVR0Po5kDuBa
xUPlBR/WvO+zkjn5fmAmq1xkIgS1/fo4OWP4+DruCrbqUAT5D9f3jz7s7DYfO63t
dAy4z8xQEre6hIV6IMG044rXRmZBEEBAVWEItLwYrADiSHZEnKxCe3EZp0BI3FJR
8+B1sDMRqpjaK0XZtosDytna8Z4BfUoiULIlItlYwU33oMHr6QDe96YZ92q49XXG
Ekip6+0l8Lm2ptCu376LN+6sHhTZLAClzMNEVn+mO3NFp83uUn5X1BYPU7IiyT+Y
gPMC+E1UZ32IE3wl7zPnkpdt2qF7grETwXy1xxfWUxPFJVyi7mGOxrrXxI/dtuKb
F4F55SLdw4mU97Z8fapZmAne5ZWOZpv5krKP3lmWnr5mxGg+pqKNJ5WHlpKDn69R
Eap7aAKv+N6xhu5Az4iKYARIsfU96siUPQEq4JV0SgNU4UmC60ktuk+CyBYWlkzS
2B9t+PM9lsim1vXhR72DW9+bvuhWa972VIrLyn00t0R9Lf3tWcb5GbTu74Iy7wKX
1eZHtQ1OSL9JzjbWq2/j2nGeUuMpPy/7CApZF6ChGHPGkvuImiMliDQjSmHXIGYN
OKajxJy+fcMmYq4ZBuWJGUBPoJbZ07DT4J9Kpu5j0WgAjV+AAzV9uT946CMwU3EV
89K0qjjmNRkQlzfJ8wcItz7KdFdf2QUiaOp/izab9RDizbl7oCTZCkadFPZBkxRt
i5w/+WpMVReGvHEfKekMvNza4tISBBkoSfFgN0sYUdVdZgGcqhb+Xr8EFt02MCJq
O8o3c9K9LUyL1ZXw9m4SE0v1Yvi6Y7pmkL0S3abaqJ9UdtUJoAVPyEwAwTWfj+Td
D1yxzZuYv3tsibaZrMwhZ9xeySAOf/guFAifr7qiUKBmvVjr1TYw02WE9CnmNkiw
nwTiHrOrYLMztZps52nxksCqEuNB3UjO9skJvineDPumVAUcSLX2B24VoW4YNuVd
2fCthu44GQ4Dbs09evjpGFIuClmxgySpifn0FmRD+zfK6cjt9nKQQGpjElBwfNMs
QKxxLAWL7UiFuyPvESJczxH+VSpRmlFt629HcOyYQrLht5572I0dRvTt5aitPDZS
MGp59aie1ffQErHnI/SHQxPCEHpSBIRtvJPpbkia3ud3Aeuhk6IacZKoPiiHH1AC
oVJ+hhZ72PD3JEP6MLKdNzqt6XadS8+0BuWQJRiyQQz4r4RSVg4I2m8jJ9gr2cKi
WA3XDQ5shGwYQDBbYX5YEiL7P+bgBOnfFDgXcQM5gWLr3kQXrKSCO8KyNhgzirot
/cmgLp3C/esr8rPdCAjoTc9TDwWNfewsI3JgGMcKTEHtc3ZWjPQZHPiKEZWUKyCI
4BrsMq9PFGxenVbkUOIpFgkceTWfCQILFo/zTwNr7ImtaDf6AvLHbPA9UhJ5QCmf
VFAnQRjsIhRGnEJILwOwJZJ5WijkFVCF1shErD5p0UCKdr2pD8PPv2mlCOw0tyNc
OvV1LqfA0ccuEtAa9YX4AGVzyohJPEguBfn22lNSGs9AnK908DUHEzyVeqCm9JZ1
yqje3eGKaXjHzdC3mYHnZFbbKK3WbXm1nHqI9IlcL84MtqAoz5iMBMMsDTCAaRd3
IhIptE8PjHLV2ECcVTGOnxARdqA6cK6olfkm3Hz0Q9UDO8nzb58VsU9l/Ly1/woj
4wFnBlJLdnKwl8aACAxPAfO9W7vuCLFbEm6ghjYDovLaq/ge+jH87bLTgNqlqGpG
0VqEB9yuMjoJ4E5ZKuMxvwfblVquEKe3utr1pRQ2IaR1Tmf3Ws4cQ0qteOqgXqHB
jISBcoDVpHMl5hY28mcBnM4KmHxnbcyqFpSN8R6pxXr+iIf5T+dAnDvs6XHXYiuM
UUlsL71NOHqZBUawh/lZ6MiPqaEaqkVdk62KR4whWPQT+JAT+ctXUE7HzaxcxmWH
eDDeNobveMgTtuxMm2pUEiLUiEltr2hZASHoEoUoKjF3OPR/m3x7Q/TjSAdnsIXR
tQvaxafDgunGhtYfRYQvjXokcaeTuwB2I9WJSN2kVEUSL53rVQt2BDepBXdWh4MN
/3sTbnbdnY01y2Opyo2pFIDycXavBa1ymSiO53uLgUIIlv455DHa9y56TFaWXnb+
c0ePxxdutwshXn17BZYIdP/AoRUvW4DzQ2gG/I0VZaDlZflPyeRZhI8i7ElVqApN
4FVfOY9CcNq/0JU+YSZRLY9zV4GGo7u/qcbGoDUiVa7jo2+yfaG8lgQThkewBHfI
O/O/bJ84WhwkD7fgBcFSwyvRHsgCTxtzs/8bIfzWsrMGt3j69MPbAI22Z1q1mpTi
NlwFZXpARxDmI8OTrxbrPORwVxG9FcSMOIb+aNiOvpHUMOG2Y2VRCjvMHQWL1U08
AcAsLr1b+FsXBh2skL57CheKazDbBoIL0xjRvgH8EyPHvwyg+K+LTneT60U5rycU
i+qce93TgXIgwj+M1cEbubdwy/WRCvfdVqqrnth38VXjDpy78s9llPKIpv8FrAig
eFMsHIPjOy2mcEB85LCxkDkzqAISdYp7XMBnZuGTnIETfqHpLtOx+g036QfnGtvh
4WXHzjYP48Ou4N5IRNzU3wxZJt+XUkVnOZhMuoPUJqdDxK82wRUOgaSuJbExykmg
D2ScynG9hV2YspUJwVxxvA+XdlRYUR2O7MS3/QUz0RXNmtxPJ5R7Mqs3btTnOPQ7
E34scaSzj4p+S31/nf7BLpXIP6koS6Y3GcNmIu4jm8Ih6YMgxp9XRoo/9GFa/fLn
hXcNeS0xm4+4yifegFfIIaM7l6uOjgv4JyM5kdG4uvxFciV1DuSzvYWVAkqN5hAL
OTNohg51IlRRjDqGWzq1GL7lqCfGsoQzAnf7dUUhJwAPLsbJpy9h7sB02ydMVbzl
tKO1DpoA713i6HZ1tsxXX2Y2U/6/3M4W4peLCkPTNIZMlQw2XTaB3/XnAoeFFzWS
CbCpynDi493ON5u5wPBImVZXzzy1NUucvxwYDWqMAvA8eSyTFqi4irFaaP14ipLl
SH6sQmElwFJk3QDJ5sPFFf+/d3OmFVcUitYRdKWAX+dYtQSxNycqvFFG+Jz1wOvY
6V5J2ZzQwmqGy4pz+N7vSRsy+WtPW4hZtPd5aOYjAEuJpKp9D7ZvwMlu7UM9af5a
OYtgTqg2Wal7UgPjm3q1vvUwBGPSSIJp/32wxG6Gq1v1vshuNYtzjdcu+zCi4JyH
iN6DRRtLwAFaDKBhRlKhGR2hXmLOC4UmeriOZX4fOCOsUAOo1Xp2NyqMZ93/P/+x
1MGq8vV7spf4wurx8T5I2uAhv2PZJ3YTZSxRbpgncPsCgXIN1TBXEbTdb6gJzoxj
P1Y6d1jwFqGGyUotJcyuIjiwU9RxiquKn59y0UEmsr3Zwwd94wC86fk7S/gLrBdN
jBgX3Alxb8EclSICLUw2SMYGv6neStKCQQN8qJOlqP65IlFq5enQeGhKBKUUl+pE
xtEZOtxM82KIe5bQnzw+NeRjg9z0xgq2JGDPO14vLnDHXTOcT4/aSDs5NHV9fgbR
CmyXML7aWWC7D4UT3jZZPMgzLEjUIQdZD2gPi1lF03Ng9G8HNiptE9fFvFAnx6zK
sCjQSyZ1EO1u9j2jLVnSZN/36uxLc4fPxctrsaVX8BdPYrfN9vmzyeApXzx37uxO
ylU8LGjjMAFxXo6mXCxTMNqkRETsDdk0u49XL/njsL/bzLmEuB3ccNpDawBXtNz0
d6ITJ96/mcjVE+HZmrTa4iGmdq3XybLgcx1b5k8S3tgqJezswDwIS1qQ/6BYr5b7
1RBegMH5qs1B+FVJ744AuUHnqW1HwaKikvSwDNT8X6gaEwTyri+0FfXApBYw7lEn
6WBBVMoX0kthVAf4V7zBilWC9eh8l20pbD1sANMAbAOA8L6wTwY5yIRV5jHoCh8b
42au6tQ0EcxesxT7MDnkYGoB3woE72zpSca+nlnBUyQ8YgTN1Qe6eu2nYMEs0R36
72J70XpSc2OTuhmHi5GR9rBQFO4hVA3+Hh4wjE48rZTm93aGV5u2+Qd15BHm9btN
AUGJC/I1qlGoMapk50+Nl+LfwPIYBc9E757vm1vqULE47HlK6+jL7tKOOG5w6XdZ
ewdnArXwi8obAKU3L073OgK0AsgJXBr7Lzx3JtVIHeKeTtNjkgWPSxITfzXL0I/z
fnx5y1ehdyp/GMG4HoFQ4sPs6W5Z8O+593LWEoD5xCJaWrfVPNoOJ31+BgoDzAPU
QRBh5Sdf7FZH5ajDg6DT6DHh1zcFwNuyj8lJO+IkXmyuraeJ1aMVO56twOKrFDq5
/f+fq5atiGQX4Ii29/Pve7ZizaukDxy6sA12CqQNlPCW7TtLZ9Ndeczwg/O2PJ+/
Ff/Nv36RpFZ1uxsxqQDFj5P9onPmvgWctPJJJFZ73urigq3IvTxvEeAhKtahF9n6
1VanZK3pC0v6C1hyjUQd6l9G9w73GKDi+ozxr5u3Z66vXB8koCejiIlw3NCJjcMA
1Onya8MdBYAJm1nrBuux/saywZfz7GViZ/k4X8pyaJ8pCLoBk3qKu0dn4Vetwb2o
scsDOX9P0bvRCfwjCKlh9Sa5af2ATQB6VEM36eUxhls8iHjvkeM1YO11L/qb9bLE
r9pnvD73Sgbd0sH79iB789AVqJsRSQWygpDJX01AbY26T7NG135rJQUAtHS9M5Dc
i3jZ7NgNzO8Dqmt4eFsYyL/Bls69MTnKDA5UTktUavzvhoOx6sITqPp+7OZB/RWx
gODdeuxJvmqIVNV8hDT/yE+yjKcaK7pRqLBTz3flWmI3zuSVffKybUl10ic3u7OA
qT2BOvXORccBtDhBdmCfTdZp5bfmp1F0iDpXluUAIYdYjJ+XFEEdxz8Cm7UvHRut
zbEqQ2kr5k6+HxOfWhX7p6l5AL6+qnZucl+QjN4DYTQzltnEavYkwUoexbKWzV+e
7xOUEFsDwcypbFSN+B/Fhx1+eAQkDSKHB0DhujXMQGuWtVM4wWrQscqQ71hoL6uo
OUVG1gAAuAmP/ozi1F1TgtCbrwT9oXSxfiL3nH2AKEaGnvAlLPOVJlTUZAS5lw7I
qOwWHniEOXkpmcDgf5q8RxS5p+q6EGxNdapKwQAX7yi/DphxtMhdOEkYXjDg2ReR
0tvqBXcC0itckcMyXAxobBO63M3ESZ58M1EM2m3JZX8134w/GGy/9ivVM9sKxTQV
CWcPwrYjAFzCjPzdVsKWZuMayCRrfNb7oDl91cJVbmsAvYuqegg8KmHKqRZ2Yxxw
/k/3c+W8WCdVvnfqvRSRH2EUHh6s9sDOTA6l61AlzsmiBa4AIWshVlicYxRcrHq2
9sCRqGVEZQgJ8IJQYGlnLSybfl4hQ5F+ycZS/1WEvJ5E7zcXH0gnkN1B56H2SPBT
1BlfXNU16VRudWvNlOk2dEcr+Y45sdt0nMavqTiN+APBTGWXD0pJKwSEx7mZbul2
2Q8Hjdlj3xS8vAslp6Yq/79lw67DBGRJK+9MkhnPY7557JObeDOLBwsmfhh2Jx1T
WFmFFVUtIpgHwKmOLSy4vmOc4Kbn1m9iuJ+JIR7hS6NrmJ4upWjBHwfuc8p8A1eQ
NUquInyNKmqOLHw7lFJPAqrEqbpKMnxUPLOrKUb6VF+mnPW7Ib1ruPaU3Jbg32To
dFRXxkwUALgFJCbhLjXiQTdjvUNMl0zZfWQamoAZojzrnj6LSv0gWSTdRQNHf/n+
68zpvAp4u3ssAslmmPTjcsmw3xj9c31KlWBmaz09mAnWvPy0rEvdcpc8MprrcI4m
Us63IbH/FWYMJaUt7CGeabDvvnWjBnFAbvoXrLP4jokv1GpEX1ElBvUje2Bd5iko
ouY4v4VIkHKtjF4sO3zXitYOY4gTaetdbqiQ5GDVChjQe5ISVTtFwGzNYp6bjDgB
WIgsvcDrefnZpW82xfGZas3duzrNvVfD/JVG8F+TU6rnpSRtcCY19WwxlIeVaJzN
nl22EFiAYTXnKkEm0FwCDw0lkevcye0LL9RCWDDLRbkwddnnlyQTfZOiaDL18x4l
+Yu8AuKiXIShblEV1PKn1oZ+Uf1BV5AzbUAeQES6ulYX5aBSgBo2MF/Ey+skFoxp
OlW6pFr5HjcIpopfX8yxbF8twdwx/lKU1fyXa1i8o09zdhUyS8RgXxGqGAH9mXg9
8H0qJsaeDMlRw/8zGr4XbRiPzqaZ8IDmXhV6O37tYzrWuwtk+KhCu87cHsoP3VTZ
bE8l40wuOC0X/lZu+EaCJnH6Dy2G5QPo5949AGk7R8m4P5B39BZVIy8tECxdjsHz
i8O4EfQ9Qh1iBPFEx4SDdqLhZOlDhoJQf3wPQ47X5Cz/DWBWuDI2xp8u4tApkn+y
Mr/g65itou54Y8QPfw+Z5KVppIfdHT+ICSkRB7hukKuURRW9DED4c8Z3DsOL4BSv
92EcrvuG7qigtRRyZj7dNLRuWWEocGPehPETBWkQ+qbPw5x+v1aLQAkv/nKzZn9t
C/rsbAJfsmh3ehzPcAt7TBdSUZvCbjgzd8nW88foapZPOnMY0v5sniK1pYLiFDRW
2LbA4QDVbXZOvrBDaO6H3/qr6uuNlXp5bhKZ0nMAQpcoDyFOlIEGYW1Uf85WKmLH
d+GA7GMpgnjPcO70JQJ7TXiALkgQvf1AZYgB9NMuK/jYW5KyzPiLvuXRxEegJXS3
N1VyRlDKvGDVcl2pfDR9xVeAVFoyEPUGCG5ZyOTm7rZvbv/FMDXWMvmWZJsOv5HH
Pr3l8I4QkFxK2nIGoG2+Zxxo8RekOodwkzuehB02jN9UwoKJMTG3mb4ZOvR6V713
NP10u/12809VLRtjcQ/+DUxMVYiO5RloBwqq6eTp8dpbmamHqFjUfD1wWhe6H72s
NEx/zOjP0fSRD/u+uJkl1u3Xz2NsLp93ljiZTKrKsgoPNNIxoPdzTcATpC7qQEY0
bQec66if+qtutrQgE0GrTgWcHQUsk9OOPy8JKLqFvoGgv0Ac6HUJZoVdYbKhoPSK
QRhTZ4lbn3IyAk680YbzpJNm1PiqC/6Mzw+LFnMjJ9QbgdfsuTgbMamD959Zb/oJ
D9X4+D0VDqdJXEnxCdr4x8LQycpVm29WbKTVSUcPAq4411l+VSj93JzM3M31Sr8j
GkcMpx7oGyyFOnSksV/L/W0VAoFTt0d6AB20Jg8hlgpPS8iJqImZMHCvNQ51kGf+
IDaUIOrBv8FA2DVDwJYvbhXE+VkY4p4rBtVpN/+TeCpmFI1vdCDX00zuN9nUuCKE
5V91GGRdfLPEsYt+7S0Jdp4YfA2ns/domt/FbF4QT4rRVEbo2fBqObGMuh0Cj1Zm
d5e8ml1YDQxNRRFmqqzaCROGiwdKuZlbz3Ai/i7RVecK5e3fiTvi6+589luN6vVh
eT4mGbe+GQcx6BquDStMhHGsv/9jEqTEShDroF0t7Kj933snQQLbLiNhSNAtu34K
AbncB7va39S/JKLNwft2wk+nBVY5fK/o+tr+O7jQ5pnGg8JUqUFjeB3wyx9qiCBY
gvEzF52Au0ejmQg8cEVEzJiVSp7jG4zNlMq4xFXQsXT8g1hrHsRhFc/FWGeifpEm
8hSFrjBPmiWqJNTkyz0Nlm7WMZe5Gp+P0x80t4I8JX5rtBhWD1/mzZRX8xDB4nLH
vimbvSKr1DVfu1VMtMfSM6BFpAFmI0ixwxSeh4KNS4YcUApwz+gKixX/Cg/AQZ+3
c4SmxN0aMuKFzkBW3Xz40IF/CmkA0cFPmi7MLkSok+2QYS99wT0thgSimEzAoxOC
QRhIV/ijieOLVoD77+A/aVgQ+S8lHYNTcr9Cmr7QSjmZrTVMIIkPBVeedKzXrZgt
R3gDKNv9cGd3FMzChQTunCGH069F5Dod8t6L9GVa+isGV8lDDR+nFY4RHgMLcTsC
IJojhRDAX33mVt8osK0Dd9jvwLtRDx6PrpKH4OdVcpaiwQCztPkOEwdCfrbJ4fwc
m/lzwOyYAM6AJDEcgPF3aG64x+UfDV+1vNgME1Z7ZkpYlvFj0F7ya7gRG2ff4IKJ
hSoSusRsicHhzTNaG3qNw40h19j8Ag1Mt74vlQhn2DWao/WPMeDnjkQcKYfWBbq2
E4cZHpZMPGl0RgRkPZ+uwBZ2IygmI0tbFEoBzWZCaqoCmEwxGfN5hC90FVlDs4u1
vlJmlyJWLl/YKdxEBxOjQF73pygPZ6PibmXdvGWFe1QZ+IGEIxr4JmWju+FqqR3P
Ukw/pUsu0+Eha0mswi53Gl3bfyU8EeXoyn51p+60hnS+58YDRGPbXPgNOruwCsgn
H4NnMNYRbzrPpiYt/nePka6JGlWZdfid9giis2U6os6bPaSVU18zmb8xfPYYqs3y
Vj58VnwbMT+2Xmybdmu34sCuM2xAg3/dkXchzirf0QZCdLBSoYZTMh0vCVFWPtj5
rUuJ9nCNLlWg6hiXWi90Q3ucO8GjWuXQ1gGohRAFdSn+TYNgzFXWq3kGtdYSooMZ
ShSo8mOOaRXnEZrdE5f11f+vUEdWeYBaCX9SKO6gHPe/5pqiDbcZyPkInBMqt66p
45ZW3L2CIpnexWs6RCK3YuKKS12oR1gAvswP0yOD5CUq3ic0Oe1WKCtMOFpXOEmK
YtHUrLRrR0h81cFsjYNkG1UHmdPK7/QAcrq6o5+DZGDTJSM1Rx2WQsaPyw4rfFWc
onK4qv6m1g9mHbpZyneid8LgMX0f1VvA3UiOUz+iDbYfyKxfG1AnlqRa6OBz1UYd
/MmxKUsIWneqYf7EHTRjWQxIzR503EVmib7ruJrRP95zS7r/F2j2WTZ0x4znxwka
NbHsP/YD9ICzHL8sg5H73QqT6D3So0hjYA862lkdA6BDmWeCQwX2M3cHOc76aTs3
YPMBL7i9BkwqBR22shdbzp2EaBO/aogUuGZv7+OKOS7twPhajZ2AI9msy2VpGOwD
aNZBBid9h6178rG/yzw7gEZD6Mt70KX4lrpec2r6wW08XC1g/RvrImdTKB8s1BWw
5DTTHtTj/Oi5Nr2dWTW6o5kwmhiBIOlA8ShsBsJ3+RabVUl7ux7eaSrMoRVarSK5
KxG6X4O/6O0Wt53lvup/aVOmAlnHzt2flxZclW0Igcx8wug5GN1CqKKQL0YEj3RA
KCZHkPWiaHiySrIRdkTRKd03sOCRvifSrE6BeMaJ81goFXl7lAarerG23lb3z0at
19IHq2AgTxTRL7QaOSyukC7zNY5IlERin0UphWxfGYJfbp+p1RJAHMbqtW9Xrjvw
CY235mi2yjRe5PjLITD+iMUb5N6hedgpJIkkeJLZ9gyPorIYYFgDUYw8+HByRw+s
Tb9Xc8SnUvDwA0qLA2JCaBF5LHiQpJjVJiN6+n3eFPnA5hAENSmI+tXD5SvYyUj9
OdimlbE9R6C6kFNtdHq8HJ4uxNYofgVx5dOY7OfZG/R5DXEjc32CFns8tJs4dNbV
mupNPrB8DhygiBVdBAwG7JKown8/NQ/b2L41cCfDYNtlYsAhzlsiJOab1B2DTogY
qwWqj/6v5pXq32koNzpvRahpMJi+A7tll43Aq3r3QcyrANLvYPObmsnQvA1oJQup
L0RVvvRhiYARxYuwGOkdX+pFJdL1LzzBd/W1Qfa1XE+XDv+aCP0dv5sSo2zssGVl
vxQ1ZXAkuSLuypLg0ZiovAX0ZJqfHbOzZP759MqpQ96nAJ/cOgjheLZLi9zd12Yv
DxubQ6OoLBXX+qqzTsKBoZhh3BjUi2SkpWfEOp8cc5MGtnx1HekZJrHpzFJxThTV
nxuNobLJHeAOaeD6mOYQFi2SipoEKyBwXKNvz/P1k9VpYl4jwonwxWHGjOl1gD9L
AKE3Rp5oCUQNRerSWKdkfIeEJgPwYD/Xa90UDZqlwrtwr3Qi2ilerVlFkoSxmyv5
s1kmRErdiRmG5FAh+HDe/tur6oTLKgBR0731dqQS6rljR29p0w/cRN/LaLmOYOT6
WKZCvLkY+dJdQeXkbR+7ODYv/1YWUJidn1TcA8VkpPNtce2NdsUL9ejeXx5ok1dr
2OSstPXZZrGvsdCkTsVWwI0NGUdEVs0D+mUzvDcLwSGZcU9bGxIIinDG1vuAV3fR
IXrtIDGcTfRG2aXVcnsHJkMYhDMnkVcetHp8r8LOOD4ylEMyai28Xz1KbDxUeYbd
lvzIg+puAbH9MyQylCXZBsYTEq1gud1hf4UlLLL7PP0mI3U6k1MJuKypq3SDXpAM
e3wnvK0rmd5NUtcThVrWCCoGJXyA/tFcfJyEYUwH/0Z/a/kye3wyuP0v2XIO0m7c
WjSNNRGuwlkSC6FM+HTYY+n0X4wKeL0ut+UEehzT+V9Q4hMqxQwjAfuc7dV3vqBQ
Lhlp5wPEwHz2Hr0FMWz0PHNGF6STbVEbxK+r0uSd8/kNGnSFVpRiDHpwk0s2/IOa
634IODcNjV9/DjjRL2ocZS932/OqEWe1DFS8GnABx65z0tZE5kRdYbgNe5GkIh76
BaeaexSu9AlUQ8uEjW26EDcYRdIQhFzaWx/gIiNToV1BESv3NrnlZvpUCYC/0mq9
U7hVtzrkcZb7lUJY7w6bL8GyPmTCw6cxbATX434FtqocpmoDyHX2e7aji+rfDAVg
ZeDcsxkchmkgXE0vJRA8HiPKQStcS7jUhzSmx8jHETa/DQ57whwX5Aas7WAovsiL
uMk4S8TZ5Dr53kDRaaaYX4pF11F7EdHl3f6m6lYZ+dDnk7GGvj6EQr6zt4cE1EmK
BAtoIz5ynIr6t5XTZQ3mAkm1ivEdsxGERYyNIbcH80Ivuiq8IlPfuFw/OkdiFjz9
pqe/kfOe64WXhTw7YeqJKe2L0QCRHP9x4fGOnIhgpxLZ44SObDN/HLPsHKtIIWtt
rvoOWnOaEZUitLYm8NSd8IgD0TKMeEoUci/0giusDlJsTjhT47ZQ/fmvph9IcyL7
Cv2pJGgHrfyO+PlMoZLswhLpQ2Ye6mo5LrwSepAeyA3wGjrlDPjJw06oBhmVvy8k
AsVtfe8ZQOoZZPHYKK3KRnhvLbsVM1cHf2Lv5i/EbjXv09nE6MYetVPskx/wLSHn
xTBR/s7knWf1R0HWxpJlkRGT4Ka4zi2FRF58sQoFYtKKjGGYIvqrsnSz/Lxy+qL/
02hgJ1/2st2BULc6v2xwM6Da3/08FgFrhsGwveyQ+/4QtXfchEvbFw8P+lw+Home
R2OBmU1R4VI8M01SXgXMoFTfOipaUN07t45SMv9l4WCh4YL6trR+M/8srdcLX76n
xAmIklZxrlgKOSkyG1Kge674UbtM63dDGMa+Iwdux/WzjeJ4dd3kqZ7y8cT/SSSO
9oYN4TTdoi1nAeZTwItLSodpb6+Su3ch69Uh8OV/9Y5V0ujCPmmGOmKGkSm1x3lp
6lvOqwehRXQE1jU0SwOz7A3jAYjRqXSCV8cEQ9nbL3KUIIj6PI1SS/PPZNDYwt+o
lUi7nsUVMUWmng1UeOHvyiCv5zpipH17waZ94UtPn1sy+CX8g06MQv8Adu7uM7EJ
B59AmzOWjstAgDaaolWC8w0LRL85Cxl1/CLJ7l3i79wAszi8+ov8qaV9/ORcU9ux
QCmwKfn6+qA7xL4AWb+CVAsre68TssJZZv8e2W5xpuZyIe/uKD/a0vN5PgsUVM++
9OXDpHPYYraB3e1kKGILGO8hC2itnq9Jy+6Sl439TtcP/u9z4qyD6kPYHF6vyuEE
wdHa2/pfuefne/g7Dg0vbp8tT3xuExIVU0/mnmRH7szMjBs9tmg3UtQ5VD9WF2kp
KP5qyIC5TudQJu4l3Wvh7f6ElmirSuAi3EtXFDhLiAFdf/82e7iVVeFqMc+PphiL
+non3OGNbZZ0aLsHKBOOK3BKJYMSstnhnTlzeW0qRl17f81IH2zxluoHQnPVxcOQ
zIwU1a9YkHzFLvuAWxr202dDpgl9ePIxAVqjBmNN70bbHfkOIWKdsHk3k35rApZU
1q5WYWCrdY7klSOaVU85a1g+bkg1ZbZ5exWux3KKZOJAD8uhvHQNGIH+XiGcnI9Z
DM4/nXz9eSOlMNaj/7yZR9IWc54o7kzi+RmP7ZLfaxCrBfx31PH3kGgeksimB4UR
6WmOq4b69qUeT1PC/6mu4isI85pTOWzmCu5fcyuhyDzch0Mhy7AetHoqTLnp04D9
a+6ucyatEuavxQTkqzejh31p6iUofRcPkmSc6bTrGKwBeIa8pqE7xlyGp4lwmDtM
RTX+rgs2WVdnczp8tQaHJRXjOR4ha7gXPsOk3gKGJeRgiaYA6Q98kgLKf5G6Z4l7
soSqwtoGXW8e8h/Mw5Cq4r31VRMul2twi8kZG54XQAml6/6qg9fSXn81B538CHm1
4MrZ0WQp4DysnAaQ1FblU+a3eXqNiT+uAC11Obnae+/gzttbWgEeKHkQC2YIpHIY
K0eT9iENPGzC5cJ1xlXxu3GT/3rxbF3PpZwiNtv11BiYgMPDylkYknf4lIy5qL0R
NcAA6DhU8usdMQCRdBn4EhrMIXM7WqElPPrWMQY49bluF6W1+gVz5qw2uI6de07H
h9gA5Pqmq66lTR5Lc9qPmgHwRStdpYsL+hCiy3pmThxBpndMwDta65/kSSTsncru
GnkLy4JJzUgD+MYrX/pI6SRQyEMQVcPyG7eL+drimxguc4N83OudOZe8HlVwK042
XwY2ySmHs/h7ZvnMqXmRI4UchTfUY8ij0HygFUCYVXMQgju9gDA9bazG/wcsJ7B6
itAd1yTsdT9OQyL/p4JKzZIdDTj+42oRcT/bqH4YViYDlAqQ7nBEYqNWRSt4Tx5/
ZINj8Drmaf8GPaQxJiYwOh9o/aVt5E6aMS//pXYgRJ9Sm+9Hf3rn2+/KRaAx8J0P
3OcM2hCXlsBZYEyCuAEOPXr0u52WnLvEShnT/hv03j1eS7n8cQfcFGheaCgl1GGP
M+hf7nEarYsiq1hqa160C5ycbr3KCnA2F1lxhbsD5xKD+j44BjWcEvxvN+sL3F2d
mkIGDu1BaWu2odFWq4ocA9W788NxId9oOlCunLvc4ASOt8Ccx8DSCjELFmGGFWc5
y47ALU0aSXZwJL+7cr/IBvA+5eaOvz0kaYy9J+nzRRtYtSUTSM7HZfnND8HxlpYf
LdduFN8/ll3RDFk1OjRBgb/H2C1yFl8cmNdv5zyHZkZG3SOypZs1OQQPGpPCJbho
WcNEoudjOpEc9ncFsie+sX6Fi0Wdfq34roXEl+ZALMEDR5rFxoA2tFTU31eA1l4T
V3fAK5JTPnL1WbVhT4h9Rn5zYIm5fPcdQj4WP7r6UPV6K5K89Zgiq1cUwrmKxXAH
Xiw93eOuEyBECIIv8OAcYornF+qJaTJAUepFFjEwvWjARF/nZXoVxBBmi8zq2vXn
weQTB531xjej3A/3PlR71b0fZWPyeIGtCfZ+C6pCgKEVFGgPxPMQLT6qjYUh1Tyv
lGmAnIcwipA9C5ygk5/jR0NLsBMjYeE3sogycfHChdn3HU5LlhsewotMNxpj6wtj
d2M6TKZ1xNw2sqnIAcGKgeKLaj47Y/cCn4Fa2KwzIBjAed0ceHh6LrdYkNUvzJhA
/14+5D8Cjy+Bc3pSIHG3HvKfhMEx59UivgGSpC3mGLRuAoADPp4cFUYPHAg3UKr/
5bsiNnfw4ctnLhDriB5LVDmTyTXSgsFlagqhGwsdPDz3QK7q4qrh6KKAtaXgceeZ
7Ay5yW3YfynbWq/ZlaOatm+sdAhuVw1bR3YJQV4aq9UgNEhs0nvE55HmIpZZ6pWt
xPZOO/zGCvpYkMLSqgShHU8hJgPylOGY7DjI3OAoSIcOso/2iervCAa17IPnutUn
UiIR+ArDAGUhWxfsyIACfZ+zoJeCJWvUL4wxx9AM7+xKwNpTu79Z8jmTwLF7z0Qk
Az9vs06wqvsb7abBrRv6fHl2q0A9bnZLs6vMsTfuZsxV4DNgFzeUb5OCLEJTLQbH
oM8/qJIeh0rU7TzixdU5qpfvq6KC86TyZ+qCEAaNbrdNmRZRvKA/3PokE9zFQSDw
xsNswB3+GVLCH6fRJhILbKXn5suxr7r0cuqXRzvu+BmORxqssNY074+zqpBrV4Bk
IfQDlwtEr0Va5g+fXfDNwnomregFE7yIAjqpkeD4xnOiIJ6iT1uh6jeX6oMoIa/5
zNfW9sSTLJuxc+O8Ytej4Hr+QphLNAA+hDdIKlj5EJRKjKp2dk9cQHKh98C6fKJG
m45WspwD+jGCJ0sZh+doAw/DgIJvBlP4r/PK2Ydk5VU28rxoUkKj0+szrX9g37JV
WdfswUVZ+YhmonsL6A3Y3hjDGszO6sCZLwMOZyQRHiyahGEyrOasopyQfOX8enhv
EvwZpQRJNJQgjf/7BFtR3NX6+llFajsRKVXbDupPLJ7vIuWXJx837q0mbUKk2M7J
R8gaI4v/dbHQP1KZoyT+wfEkjXZAjLW6sOrLU1STXzzETFXgeZtGY7q+xyoOjcuH
y+SiZ2fiiKH7ylR21kp4I0E5yWGuWTnunbENM5WzvHqiFUv4xr0GyKNpG1D1TaVi
150b5AUCNCS0PKFBi5O6WdzSpYkix0qvWpn7Fdo5nx1kT3SQbI8KJtWj6aCcmGHe
x5imjxdI3oqjoigfe/q4EkS4sX67wHuIpMGxAIKMUEQB60I10PF+NGFfuS7tH+pI
G9HsBVl3cwspkolYNh7IBsZm1lFbepsWdTQAWZSZJPA1sQNrxJPyiv4EVV5IAPzz
Mv5C4FpzQVn9cEKC4wuroCgPELTzuQpNzK0HSFq7Xb7P4swsTlXLOYko3sB0BnvI
RZRPUOAvr85OEvCCUh1CbYnWTgtdZnFoQS54WKGh+XX7h71FR6nV62Wybc6bWoIR
a5nNkrnJfDPozREIlV6moEHbSiZlUY16tEk+WZZY6UQGVxVS8gc7Gd+aKj3GE0u2
wOyBrREpzU+USCySWV8hNCAmgZh9mXoB9E3ky/ghnIx5Zag+Je6uMaf+l1FIbJau
yA/hGvD0VfoMQTcAf1cLLdWSKBYdvb4CUkas5OwERQ4cjUcsadfbov7ZM41/lWSL
cfSsXyzrNBddcYTihBWTHY9plFuzaQejj4nSLvT5vIt5nuVmwox5t+xfobxlX+vG
LJc26yxwURPjltMaTpuXR/irRw76ievlRB6VGdKDsgfMxWiWva7RwA9btIqsZ02e
fYticCsK0960V0bSbd7F8EkcSWVAVvRsTpoX0bXeTAOwP3AF2OwlfxnutnXIp3pc
LLtL5IZRTPfX8jGlmqZqY0kuyD6Smy3FI8JlJxWDAt2GIJ+ChQf+WtNFbybdSKD0
3ye8QVxLwuo/fjKuIhTgxl4Xd11k4ZhO+9QN5v2N5XNzZlHPwpAfXBp9NqwpWL1C
usqOU/b4IL76LcLehtTn1AzQkIzvSUpC+vxjEG778GQoZLerNecGXWFSLdKMj7IL
RoX9lQXLfXeTX2HeySn/xG2aiEYEfEfacoDiKyClWkJD7Jr51spVbP/iP/bo1xnI
IKVNTjfY/0LqJr1zIRPiHi63IqVrg8J4BX1NxUSy3k0ChwazBmKKiSlJKPOhFfzu
wsn9xh+KFJIEmrwkYYa18CCOjzz0q5hzmImy/4DzYwxsI9fLGQmea3eE8gz2DJNz
/Qg89mZXlVB0DSJ3lFa1n26CKLhXo1ks6381qybswd11lhK+w8OqxNVKjQd/3wXZ
L+Znv5IyWTBuP0C9VqmbRXkTIDJ4pZkUDuF0zWkBzS9vDlPLdYo/8hLwBK3MeQlt
KXoCeoUFCbxNgoUtgkd1/zuOacGIOZa3ySr1f+cieA0eSIsTUL2u5yv32d9pfzzs
GRCkLhH0YGFWdYWsVXi0mpy4c2ID6XVU0qwNLQmNMNMkY5EB3bBXuS3BsHYFsuB2
/ummBnobllFd6g+6wpa1Ulz4vuVoeJU3NSsJgSJ4U2usUopRtsFmhvkhW7B/rI/3
YL6rJIH+EvIWAe0H603jlhz4893biF/Ss4mYMXvLvOBgdS0j60qrE0Vq3a8I2g0H
39T+v1/fiCGE99TI98DfGqbI+ecAPALozuPhdY+ZNuGBVkNcgn2C2563NcrMgn+6
xP5Gs71I0ddhx4nuhhXe0ZHLDGsfVZtYMZVuBtNDvBwx2al2/2zpFigFReZdQlG8
2NP5LiB0tB3hpXzhIq6pQQMi9D7mgct+HKFMdvYNt90ZCNYdw6U32d8MVTaO7ofG
wcv642gWbrwSRwQ5cytF2qTOgizyILTn9NPmZr8kVCmEwBopD3rI9A2LBz4zniFo
BnZ5AW2FCbXhX4I9iF7alQWjfOJWBZ/SqPsSg6hqmC+0OMbW3VbszfLReibDPXMD
A2mCTffKeH0qzyz3fQG1G5U27slSzgaoMDkjhpIURTG74SYBt8zYUu4UwMPPIVHf
koTus5eaaTARt8t1xcU2tMdXqj3Ex534jva/wXOrDAqhgq1N+Rxs0YEd9DZD/wg6
iNxnpImRCnbG+iCfTrPCv4IQFb+loRhWz0KAQZoz6p2VvTilkqRLqjbetP6UvsGq
cy8TofJ4tG+wNH0JIOoCdVS9bVOBHT2AJd6tYnjSv9vdLo8DjozIfBIvPLNt9VS1
vGxdEvG1Lit1LFmIQctTVZKuBLFPkUT0r6mWsAl/g/uUj7ySUWs2XVZnjTkdLoRd
kQh/5gWwG/GSR3j6Dwh3s85SnY/335+9HPoHpBfc87rsAoO3Y7OcscdN7q5sSPFw
VO1nKC9LJprDJJzSnN+ByaXVTMKwvhjGT7fx0ngmcr9VvxhrvUxWWB184DQ4bXiH
FC3QBm1/194VDaK55OfJdiliv7N8ct2sHgW6j7sqx6FpC/IzLBB2Rzh98Vxzv0Q+
ogQ/cVwcNzebgduzLYn23SpfqXFh/Gneqg4BrUBquxebOi8FnbFbzWFY+dgJCn5W
BhcwOVaDRMN1HwPWd17wHIHvZMlzJ7hWuoKVIplAQ7nfg/R+GFmO0f05saOuSZSJ
6EYx7X4iH2QKVpERI9CQh/tqUtpuBI/55wd+2Jxe58+FW718tgBIDUxpvkz0GOwT
wRiPQh202d7D4vtQl+DXiIdq8hyAxMDOUUv5pkM54hdpg7m0Eyrl5144tTIuQEwu
burclFV5n/hfSZBvuMFaMtAnoEq2phS82AD7eqzeE01jpsFU8LxFOjH0n9KzkVo1
4Lrya3WpuDoZSLlq238Lpew/C71EfTsPyKV9R45G0F8bQq4hmwbf4OqJFN3aeZyM
2cQrdGIjbhI/zQSDjJHishQMNnHmaeGb+GrZF2jLTk2BzC/N1S/kHt3fhvd1M/Ov
fyzYugtLy6O5kdoK854dBmuwrdOnPT8BcS9VPfwrFvUeTRkfJEf8ZLA8zeT2hgd6
qGAh78Wtas3ng/9YwAuoEqDeA+SP3cZf+n1sKCV4ODU2C5axd5VAelPktdFM/D22
Tcap4bmmVyAu6nqPuNpEV9tjA0o2Dig6d9fmy5De5LfdBeV+7S2cPhNMy3JwgpBm
b/xgOplupoxdJ2q9MzgueZA0XwYEtoc4O7mLhJ5ILM2hw3i9d8Qzztu9L7TN8079
nd3Qi0nrqofYfHgaR0YNM7lhEOpDmZ1cBY6+AmvFh+0xyuhjUkcPGgJv2QmkRcLQ
NUzf5VeSm74ffguBK0KyOHUpQltjmRPYLyeuAx8AOkthjptDp7Ukea+ks6ha/Io4
je8RObFlRYGwqW53sQRksUWOixk+2DaS0oYaViubLSplw5ZtQOisZ7XkVwn1m1QD
LjkK2bV/qwsv820kCoO5A3vaF/Z4BUm+LT0Iwj23Y2LSvfvLmn6yAtmhF2Q+k4ql
rCHQoOHqik61NZ2kA+c8u5dS1fesGSgqom3+Tc9pJ4RHSuitoUwJnViyr1zM+ZJ3
tiHPFm1kdBOBlPVJRi/XIxZg7+nQv7+mm2D1FOh5cG7NKdUHlUFhxAvvw/LtD4ON
9eGXus9qHpgb8Tp2sKLG4o6ZAt8693Z4pCsF5NLS8akKSzDXmX4IbN3fH+KP20mO
07x6mLFmZh3G9U6Zq1hTJWzX13lkrBbpaR5zI2oMlJ47c/XKldcRtSmIPOh6Gf8h
dUgCr8yLFfwfQtlfLEjI0lPhGsVllqBcpi8ecrDB0KXnJcQUziwzbUY9YJNPNh5m
AF1TeGXepfrLUwGsrC/KLm/h1cCz+i9QH3cEaLYc9d1SLZqzn5mS1FwLEhHDYucR
jqh+ubDPEfSB4rCg1WIumYb/zbD9pjbdsUe8nygYZzz/4dCx8YhEx7YbnAIj5han
YtsUnkfZeaDXItX0xfLgX/gFG+zQHL97MNLFj/+fZl7acRoKYi8FRs2fKjpT01iY
Dv+17r1huxqtqXJCy7KnM6nk8c9NK02GiVoAshvm+xQXRxy8rEn7gtVJN2C8Xmag
JHjbXletAb017ZX7r4HSJn5DYdQZezmv8dsNxEc50Q8If1RnjyORU/6pZL+Kth1I
2aaWmjweHQlkt2zbQnET5iZAzttRULuGe9Dq2skkEMjY+HNVPpX4eGGN6uFRkL+M
dfrIjIY3StgBp3DP18KjKGBuJA1X05g8MyO74QNAJDDOh0m5KglzHD+jYQjQWHBB
Xz87CY2XQ0N+c6sn1ygFCSVZgnoLwn7W+76ETPJRElzI5ArXGQFic3CfkAMAUM+f
sAeC8i2h5b+nmlrB7otmXYMqF5yYwZm5kOFAWtGz/RfBnHlPFLD6djlbR4u9Czk7
1s2wzn58eUKr/J4q1bwLH7KpfnBBXl1NuYrx0nUyvCeE2uXXa8j2OxrL5cdEvzwf
WC9cIo2/nnMRn9wZS/1Gs4+WK3wdDC0IFrtijXjm7QkQWfh41Vp08QiH+fOStdAX
nPk+h8zrbZKi0m72/sJ88kfhcgagxEalmR69XsptLXy0YXHFHq67lGSVfCwheUyV
dxPMJOaNRlqhSkIJaveq8xBVHa4VBPRPopOT3I8tKJGL49ERXwVM5m+841U2uh6K
xv5U/C10hyQX0u6L9XuBjhKVe/nT1h+D/d1yjC3u1B7qvNXgmWg0USj0K+5OY3fY
z+LLNwocl6TM3cUKkUeLmy3Qh+AGTQVOxPfW4wrsOKd/3i4RmMZvzqOTYuDbetLK
SBv1J/FRWxiwf/jSiU5RF4XvnSjQTPxtKGv0bMaggDdozgDuI87lgCV5oQBFDh3+
ycT3lVRAt6w4Jpmb6zEu/xNyS5s+2vU5Ys3EbCF1wcDjdkwYvci+CQJsVzT6KSLr
I3/AVn2l1heM1QSLz2/AlJvPpqlBTh6je9K+SOzObJz41tFN81J835AR9epXQFS/
UT1dfXGqcXhiubuNGuD0L934Fd0ijdVJOwhDa1XpdDuKbpqpL2P6tnJQ99g1k5ME
hapPeDDpgK01GyUNQGuAdXGcj1QzoLrH2NLFfq2GAsJq/kzk8eQo5f9eMoShd/QV
jjRybSeUT3lCx/eUfzkY0lfb1zqKApnegNoQuy4L1kE1O69/+PrUWPo2IeVDfkoh
Gdmh3Rs6k9+15XBcBMw7qW5UxwGPUXZD3AXQD1KfwG2i+lPNB4XRvqr3iSL94HC2
aAZp5M3qaDu439r8YWA8gbwtpjlrwkAqaTHR3wmNu4boDu1IJE5N+iLu7xxQ1xj7
EzJzatFbcDuUgMmsOIcEAiW9CiNDI8wN+GvOc9KnaVpOaYvwEQFLCczMyU2n7QRb
SvN6cJiejLsMvZYyYwrKvsYGRtvVNvl2l3dtTMTMwLkL6nYq1OY2INXpEDP+D2Q0
7TyV4pH5pxPSwXPcEbV5QhaKFVNK9b0LYuu9zxoNhojiVk70fd+lqlgEN/k+EpS6
pkXCVI5dKt5qmVAkwkf9Lt+4zwHI7s0KXRFKmIxlASVIC2XUR80K1zUk8RVtU9aR
DKxGRrmkL9yYFhMX/5mCzDEQRWc1Dy3no6TQOrzsttB75/0L2wyBmSGRFo7B6gpi
cnRJvGX2mgIBlbNWa1p2jSQgWQNNuXVualCvYDkcdirheEI9Mt+M43KqAC/J8y4m
0uBguOtbLA41Lg3vhLmpTgWEKeuzIx7MpRdRWoepD8VFDYg3YIztw3r0K3jzACXd
GS5umYXKB+/GTY8DjOGdbg9G43brKu8ioruI3R37mdQSFd5id4G4z15iAuC+WToU
KeoLBXCXBYFYRXx/xrwHFy/htVGNdaG2BdE41SiMbO/OTdtK/PwzpJq27gayUGBj
YfVu2tpIf+s0+RUrcgxoNXnIZHExwNlu/GQLXcvbvRNeUnp0cnFVuTk629IHwz2j
/CuOY3tRCHu+PwVzGw2I7Hh0pXMFUC3P5RmksHFIUv+VFKCtxU84uV3czl9qsnTt
JxVJkC3p4wdcs0Lx+L1J7Suo6fV/rgGFwuXMiqOuCkRIqsejSpSucXMPJbiPvaED
XZtYByMfK6Ou+2RZdvS3Fi51QRSGUvcPAe7/MTYjFmx6KiMn7NS7g28oE/NfVOCR
nL+pe/LGy3b111Tloh4iNZYlvNjtlbK3FDvCMy+r8l9Ia+98emN8tDf3WZCyfVyh
VcBWWhQbZ319H2RwgqXpxf8gqk102vpBu0y1hm8UqoMlR21RWSX/DFBJpILQET9p
eq/JLgLcGvhTKv0W63fj1fn3xL5RCn+BAKLP3chbcM2Rfd/WDVd5QR1Grqo7Bdcg
4h4GPdoD/iKvy8+n/ox3Ugezhj0Afnlxqj825k/+ORYoRgCO6TGvNa+1xHRmO/6/
yTxz790FjsfCFKlW1+r6wp3qzLJYJ/RfcCywxCupY/NwGrZvEAGlTNQc4TH690yC
uzHazyFDiJ+LEupk9gCSu+FxnDg5PBO9DKs4cxhkeqaih1IUE2fplNKMdA10/c/Y
omXtEDdhGXlevuaiTXtyxjAUA8mBGl10A81F39nFwGIQX1t9E0WqwP6u9zaKWHlV
+l15yCdJfclQyGGdxSRl/MnMA+RIYBKL7gEBkVZUk2TR/qGPH6NHRx35l57P2lO1
vJR02ZzBq5Z1NNaCYBD4+M7hH+Kqgsr27YmQ/ErjUOf/AHS73nx741pW7F1sK872
ljOqJRsx1QLvIdoLWPAlH2R3A6fnKT/efi8eelZya3K4DUOww5gTFNU9arrognxe
ruwjaBGKyuNNevg9X/dOe3IzJk/4Ne7JvI5xWZ+5soSOpEVJmJFIJot8kunidLho
RUJTqzg38/ibI2a5geZhV+pxiDNTgmVZvRoKVuASRWXdNNHGVlSWB9KINtFM295V
heWGmDLRTnajFs6Jj3UaXojrF1bdLi6O7vHtCdyPvrfSEY5H02DVkwc+0MB3fZZm
Fp0Lx8qEoa9JGw2nOim5rtyta7hmBXm5pUz1hYuVb8WvBh0CbhEZKwZ0T/4xYZKn
dS71s7f5frGWzQLlADJaCcrY1oPYypBHVI7tghUtMj8xLdRI21ai2KfG/UsRlBRy
eDrgD3P6UCE7KUibxiH5o7Xy8nCKZY0GDcNBZqf5i6aENotsPqMfBrR4YElUST7M
X9oFriwt0DhvlAYiHlQ5xFzqOJ5OsD6e0nnReUqYLK8n80ZtgYWumZS/TcOppGqF
PKF6Tl4PdUvV+qEv2X9tkDQAFojj5QVjj3Fv/JxANJ3f5uIL7OisoBhvYtgK/S47
UzZMxw45VUpw5/6y7Vtq1Mw6xcKausiCm/DccSM4za2XBNbt0x1r/KI5wCkhU7oi
GxiyLoYHTqciJSxIZsek1V3kP1RL1difbf5otu8TDzrKICINgMQnMeVcOvcyLg/n
SXSj6iiq550o+3wWO5O/bdroa0Efn5uPb98/tn9yRBAq8t43NgyxF5xduNFWpcwE
dmSQdkBejEaWbc768k7lSHvw5aD4t5HG3nkfCFrEY1MCqR8DHO9VkOFGFVayWbrA
Oi70JV5wetprTW+1+TwTniRlNqNZZlSqgzA/aCCGPpsy901+xZqNv3RrTZQqwgbk
9omll1x8OsIKXC/w2JEnG4FxxJpQyORuJ+0PtcQ7O1Hkk2SVt6CdSl0nIuyaqJD7
lsfJM+/MHWkfPSbiz9Kfb1F4H9ga/bT4XWFyIIlIloeug2IrNBdS3YqQlX/wVi1t
RpPRouTlG0e2G9S2tYRRhQLdRYuaTZ+qwlt+/fOhIaANKscTRljP1ZQeWU2XRW2H
55hPFcoPWPyXURdLbjBJlonoFsSUg4RT4xilOGcExgV//aSY1j65gwQ+qy/J33QR
4kWKkOIEHebk7nmER+uHt05AK3XNrhF/+As+sP+vlinKA9jO4hExoOp/Hbm/DtB9
yhh3lqd26b67o0I85JvFPkMMa53Rumi9MuUNsx8ZyCZ8Ucb6odzh3MBfxV2VasM6
qOidO+J4/tDYy8ZCTHcyx+uDAbc+HAOUSKVqAPWppcDv+zTbSuHYyUR1ICppu2NP
ulhHNW29GGPNjNaXjniU9JWQThM02i2S1/s+CHCIlU/xgX+OcMasDgWUwCpre2DZ
usxdgRbRJovO+13OcH28A+XInJ0K0GvWLrSFAEGJ7S2nbSF7gS0HPr2VWR9vHcbw
V2cF4Hbi8CSfAroydfhOYgDLCpP1aJ1LJ0IhD8ZxTYoZF9SsA6Pe9BOlizdjoY8p
resTvRrv/Pk/e6BE3DkhYXHji1FtyUSvBb47K/vh78E2Y+ekh9esObS1XWOiStwu
zCH4YX6ABmrju7+cQa61qkKhlpbnUzgPKAql55IfxVQheYn7FLB7EE2DP/Gp/7Gv
rVNi5ViBk43HN4CFK2KpAJjhZOAsD2JLPyxT5lRNg8Aqbh4rlHcGsBZTSv62GkPU
Qn2432MqVBSM1Nsv+XVMhqihEmYTYzcA60+PRLfpJdgbdgNz8Qak/q7u3I6YtY9p
zar1V4UgrNU5Lj3vmRUr+LEyV7xuWXUNullCc96Ro/WnhIYf+TgH4EN94tTO7lJn
rpkGuquI0XBwsj0vAvY0xVuwYpmPWdaG9+4o/FhfexgNMsPwsyzcjHv+SdwP1KHA
xGHvEMYEu9tZmeCoo1fRNegdpz79fP47sdm0dOX19Srv2WVrKbKiMbWxxX0dHo7L
73iUFQm4l2+76xhPDlNqVq3Blf/fgBHcQ+FLsbyoQojHVQIve841g4lZykJA7eXx
9g3Ek/jprjfxl+JJO+REniYYb9x48yFpby5XtlmjIdb6cO8fPJ+N7Eruy1exmLCM
yB2kFXHAwfkonOHfpP1uyyemVmh24lB17em4olUIupwHyRtVPk4wnWkCQEhwTQde
L+3qoHppsj7e1f8gq0GF0CVstEO55hG+hMcTFFLkBzs7PmbFgUoSQ1im82Y/ojE6
VwKtGHJyHJmZa9aJfmGbU7ZyplUNjNpMRsHkThmKNI6O4P2Q+YM2lsvxvcBMNthJ
okicYPJh0VqxAJurrob/oFjZxCMTnO7+kf00SD9cmwdVPPP6tkQ2vMKgs49riKwo
aGSza2fMNqtKpWqatlrLbIRpK4XwViNGeQrBGEezmWseXHQ5E0FlP2YqBPow7CEK
CW/I1bbrQUHlcGw1LK9oYLdcfZ0IgNymExRASAgDsHA8Ooj7azklKZ4GJG/+Bf5H
XTPz+Bfvyepn7AHj5AyVprf5NnW4BRh2UbPY0SPRjZinIdfS3PaMljUek8aW/yxf
e18vmzQR61H/vIRZ/1SIgS+NZkV62U3bz3NmL3jfmGFjYaitTnMUvkI1dYJXzhwE
4lUbaftQOJjbCHthCUzR6e5mMi8tj+F3MtBUDmj19WoJY5DEttvTlMK1Cdnbj6ya
r5vRS/L9635TLcvlFAL9JmIf1ze3l++ziZpnzTgu9iAO2ZrraXRW/vMZdaHHoYvd
INNMvE1CAhnjOGnJA06HJwhlMOfm5FgexVSzW0KaneGvgjo3hblYnZhhZ8wNvhzM
vhBHJ+3jFwhGYfEbLZk6EBzBoI6p9nplSa/amgBFGscwkwnRPlVzoUNPYNvZT9uZ
l2GX0wgCiYIrQ37o5Z8jMR9qDPiogCyYe/w9f8Qf/1D3372C8g1F5OoIjWx3xz7s
uD14/+3iiCBpSpRN0peZMjDvXK9Ll+Qh/k37li8ZYu2olLA/Ls4pGZvwHPCtgebz
zQeQz0MOBW/xLy5A3Oe6rPSMSTHNiewFY+dwvmqcM5AxlFgyFVe7+OBAlZD2V2zP
W/k1t/04smqyHzUz8hzZbrmMg9gz6+NaDMMoXDUnetGrhvdxABZ8IWJKgoVcD4cC
G//7kvMht5mCWTfisjzmWREe8NHyp+0LNRnIV7wsvOyJc/Dps7MnB9chR6jIyA9/
EaItaiJeyqZClKeUSthPA5+csXG2F3z9lDfoOVj5YpmQBfrnEdjzGOf0zed4ubvM
kbIKNp0nNQxSa3314cCULhgSS/gf5VjztfB0kRcB5Pd8MFOlBDPAtRCa/uT+qhtq
DcdRqqC4tfHKMdKJd6OJ5wTX0Z8nGsb1w/DuWVsyX9l+Llhvz0QJFG1H6PgNj2cL
gYddRaRwE0+C+1r6at3VPbPo5ZqZVbnCKyOchzNvdcLfemHXAG2wV44ntCnMTxFT
g8CSMqW73XESR514wxDUlo1OTlSTJorUjY6t3mFzb1JMPOUYda/FiCIp4uB+4gd5
kSPyl4p59pR5xcMfQlg/4Qd8UDLynFIL08g/WoTjTF5ltLSXqERq/ri3J4+44h5M
EK5Y1iWT2Gegk3zUpe1nnTnA18UEeAuTHaqKbrdyPEhuxsWur3917AzkjehON3C3
jXwl0q1jRGE1r7RO/dSXezRT7cRxVJ/VplohNOTh6+V3yzTSbBvI0fE1GGqAZio6
S74dh0MyRxJ0ICtQe2m1pY9Xsnbz+TRR4OFEDMo5xEJAc8BhnuRTA+Pl6DG9joR7
qjqwGYr1K0HT7Lxml9FOH8ts+veYgkz/tQMCOucEd6QCmAqdibSgjaDGgODpwTV9
X1/TF3YIxoQzUQN2bwETqYNEeBN6tH6kq/JgT4fcnY0yXr2fiC7xIT8+79J/O1ck
vWsJzs/ePPotRMA/sU42E2MxGta3fzE3M4cFBGuNSNWZCCebznOPRcE/G/PUwkM8
oo8ORoEJtT4KysGw/jO0pOB4xRHvZ/OUC6C5IS/0I5mjHxfMpIsOU7ComPJgds3i
0H0tm7jQGDuo6ISP3zO515Y7ADbTUdspT7F32AsvpPc9bNEE13DZvbYE5T7KWlhx
KcdKfAOQFSLwVVIoAl+MjDlPfD2dD+ZpoxgwB6gKGws=
`protect END_PROTECTED
