`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ChXF8N+oSSMzlVkMPqMS83uXDhvhxPGwKlVnDfcXbjGltvknS8Wk4URPBgG+L8nj
C2OboGVRClR8PJB2u/8nUEPQabx2X+ETbXEy7iPEyV6ith0p5n8ps19XKfKzBVFy
pWP79qSOfWSqjKGG/lL9E7uK9XSrSriHV1l0qcYaFQIuOzY1nek7a6qVUTcVPev+
kQjuSdhH/h59k867vsMEn7HuBpT+XQEMxeR3k1wQelHNTi3ZfH2FV4uiuCrT/dir
X/LpXp4lqq2nqk1DPZSrL2Eh4nLRVXXuDaY7TfqNK/WDqS8PELjd9Yk57GyWI8WC
xsIbkveQY/WpIGgpcjmIDLNqY1YVWGAUQu/Vx5R88d34zvc5TddaLQ0WKCnHeXYR
kVsOvMZ3o69qK3DLjDolehGVUsPjG48QGm+wWJ5QAcGSHLZiMuWnXF1H8wP79TJE
dKAFV5cK0+WND3VJxOJKkyWMRqAdZ3LjTfmAU4vTOLD6HdMpa7qZUL3Ptyp46Tdl
fe3KrGpU2jfLKZvlrM4IAM41bju4rTMby2Bo+o5c4wb03eEiHJqtC39FIHb4S+Fk
vlo+7Pmh8nvcVomoTU+0HbVoM2f08Gu+bYbPGnPnYlFWzl2saCEjGtKG7p8FFikG
d/YkIXcWJjQHJ+o5EiOAsPziNp03wZEojUhEyFQAESZnyoR33ZLEd3uD1n0WFPGN
x7PUKFN7RtOIctotfXLoL6E9ht1ZbsF+fpXOVDYYvI2wUxlk0LKw1DAdEE+qbU9t
AJMP98bKI950q5rq9FTlLyLL0s5x3hpLYLR1O93KReMfDsZ4r7dlYPavAMcG9K+C
E9hg4vpgL71iLs7R3BlnesZbutFjrUjvQknzgSW7Dtsqq5Zb5skf1Q3iPtdGAThr
627DKJciGBEfTmb8ghLEYqA5zGsqN3Rb2WuGwFI5V9MP+8jDwIZa+aANcpkw4F6T
hsiDINJc8WrSKswiMYZljXihO/YFDkRfdCeIAgJnwtI4ErVtO8T2TzeN2Fr+OPZe
Btemn3qyz6CVISDZ1zFGLYlxzoHrE+Gn2SwWVUqpD/M7lCXB2AWFY1b461DwJccw
xet1e6We9FFlhOndSCa67tf95qCriYln+EthLinH2Z6QKU+oy8hz1XynGvU7VkUd
MvBmZQUlZzZ9ejxcc2ouVMQtXbOM2ISG9Ge5X5UG0/tlb3YBGyNu4JGUAtT5YfTm
UUvJIKSXh2X8SgzmpxCXQg3UEFjxnpXjo61WJO9Y8oI18No13CUp+s5Gd9lg2D6B
pAR2U5MY8qqqAhDNyogCkZpP//zXhJZSYIQEZt9Pkvy0gI/THndPMoBozkuTUY+M
yT9AMjVsnZWetbKIX8VM/dFxiJ16AJaX6s7agzTaJus/AMFza4+UjKlkwg6YUVpH
LxByGaJzRXqPFEl2gnY1CWu5zYa0854s30n8uYm7QzrTWWiW1QI5cBZU4Oj/AgXM
754VtU6CUGl3gCpY9liEFDCs5/+8+riuLJ8IVA9cGz4+nm+Vq6V6JJvnqwmjA/wq
H8ZuXeTpYfCBFqV2B+l8pzy+jeiCWBnwDYK0W1F5Jy9+9xE2GsJiZU1Udb9buLcL
FNhIS4ABTt3gTAMbECWIGNn3lQ9yUVf0eyZ3Ucv6C03AGTjdIQJNorDfm4UBRpIP
Kn8lYTWAMVWLTXvKrdwDCmBNcUfTCiNlaspnV2x9Tuv8USMHNnO9LuD6ZEbGcBIE
eAYZbq2EQYrUG5wYlxgo5dFLHfGtgLsqsB3//KTvYHR+L15vsI0NrLCY2szZzLGJ
iBqgqDERMcw8TlsbrYRhxEeeCQz+rB2fig1/SZVso2v/y5nAEuC8mQXVxPTfK21o
rx/RHlHCd8Y0yHdqZrgHYGdEvt3/akxPdBGowKVeK5vJqlA6Xi6hUa/AvZUW42h3
l6GyukoWkru8pGepvPs0myH5xrgiF1CfIVjs4o/G7EOZgzmclpzor+lmRf2/YgZc
nVw1KWa9OZiESKBt+juo2vpPYLzXZeBqXRpFAinR4HdiiCtx7EKl5fsKKe3IAk6Y
PuBoOp6qSyLKM+vQ94Tq60Uox0007kC3FGN53lxqQrcUwptQmWc+q68EpyB2QfBC
p+qfrhr9lphQuEqhH1z3pEEMvP7tf3LPeoNOW4m1C8UCkR5TgPF/XW622ghu8Pkz
8txZXQweiv85Jng5EMOwGsp9AlQ4tSbFBNh4ybpQuNNxvok4VMUj0gkQMKJSIi4E
ZkrFc6BZCP5xSn61fQ/nAjXJOWBT8r3NPHTwSs8fuvM4TSKGujdDFETTWYz9pefx
u99AbD+81D87+nJomqUV1heJqj22o0hhmLkbDcZWgxSWK8Fa53u+aDH/xqFxcYy4
l5IGeT+M7URIhNmbVe4cBH9+XaPARrm8WvnP4p15PvitsYRoqE0PNtgYQxXuMox2
rsWVeq4i9XfFMrXloeXCVw85WIOFHrILpqxfRWIytS3MLRgrMcdqH3fnOhecufQG
inDNwFm9T8PSoki+NiTnwozAdd5Ke0yKsZxLrLcSaybi6Ao2uiiPLtzChwnq8bdK
+Md/3p/6kBAHIgoNAzS6e65IQnQ/56N2+P7e+l3hBvHvLMraKVucFpNHk6QsS/3+
z1SfvUkELy7aEhsA2Sa6FXDGBWFWwXF9tk1bRYk+b1/I/x6L/NGPaYMf2XCaqu/v
RruOUPJbe8wKX/BuG4HgdGiCiuKRjUEMg2nlWUTuoVyGxvQ89lZA2c91G00goqzP
A6FRInp7qUotcSnWYBNFkTJDTZD1V3G0BKOmoD54tySZ/upqGQSOQFAelcEJSYzE
rqeh8fehlmlaqY4A/Y4ij1PZ9frujltFWRnyMklX0QUrkYJpwO2wEWXA0GkguRV7
PyIbjG0sMekWggc7rMfXn5yjOHpkxmVKh9J6G1gf2mlftleh5OwmNIYg+jWYsi23
RJZ2wbUkPh6kvCHS6qA+Px8M1h2P6YPd3Jbf5L394EEpK1+OZ9Vslm/U6oHegyTH
cc/lrGhs6H4eBUhxQODqcGfxtRVKon+F9Jh+RP0ewNNrYwL/jEWNObdFpu75YRFm
9xCNZ+zFcQGAvuzgURL6oP4VVVHjy2FtgjVacvXqcXI9mhuRDVb6p3wYqXteIsBV
wADh0eJaEL45eaTawX80feVG6bUf7tm26vluBKLy7KNTJAnv9YTJdM7vUDo0THal
XyQjwRTlencmHpj8f+5l7iAbjmaO+bs8b5PcdujNHoWmMGOzKXWxKgBo/wD3kLZ2
DerZ40Qb6SoH2uVLY6CMA+AOSx3JGtFOsCG/VhMxSqshhNkVIdoT+1H7CAxwvT8c
Gcz7BvvaPfYK4CwRyeuOEuPWVZ9VlwpqzUuUpetIKZ+QLUeQVeCv1kQjFYl+MOmu
Reai85Hd50OLSZvfpouVeOKY/8vuT/Q8HjKCtjHEVrKeqBAM1L82ucTltyHStWrU
Xj6+fQ6k6mfqeUDVU3wOG83AycD8QOBb+pqy14x9h2bO54DZbgEJ/I5v+LVSzSHP
9qvW7pHSTlRlhAstWwDu11C7z3p+H3+e/DTwpn7d0SgOpmxGGxxm9yY0n/BEgjkA
+BiVBBof8slLCDTj+bNFF8fgSjQyPkSH3VgF5xDz/KmrkWjq90wOPHT7ZMAXISjE
mIMMWuKf9IF429MnwVpsMLmGIpPvgH5j7uwpGdnXqstYAS33+lPe1gQcbYuH7jFx
HoybeqXrAHqyNnUrOh/3LVxiyXUMqOugGJCnOf8+VT9BY8HhTdB6Q722exr9hiIY
czvQpohc28CjZfP29IZ8SoYerkmxzOgUsen4l8ujRlG3XucV0Fg9MvVGGbklS2Sn
wsYInrAXP8Pj3U/BIsaePnfefFwW/cleMzDur66w4hC7tN7vcegAZP0Yr+BozGbI
KdYSBUJQacZD9IM1WSkCjCpLegDD/YGkq9E29x38xee+92DWcwGzCkj9NIkg6WCa
/XKaofJuTiRWOk0hoZxq2k92yok2jkx7VGw756ciGd15dkrWicg5KVpWzT8t+olD
Gmmo63ZnhtzNL7NyngXLDIXVbg8m232WEura/64wn7q5L02o0eU1yJmjFB3Zj+dN
YBYkCnkTpqi0qeGk9Dnao6o1snKZz9m7rFrwBq6UX/DBahAl7C+mN8lmpOKUjNIG
eCTRZUwx0Cjpr6vJnagretHUphRs9SprryO9Mo7uOIRSJdx8vdYbvN3ElGCOswyt
BjOVbBCYpN3hhO/rt4s0DvlGAE7KXGhUtN41rBYmfd2IvT2BgknW92vDmWHav6rZ
+0okZrw9xe9VZ1DTl8u7Ko4V9HITiplS+UZUADCEp6uZuAyORsPlSOPIbfX6IosC
ooiRoAmjJAgDMAu4NIWSyJF3Dk/PMHHGRuFgMAz1Mn5r/pqyNroqerT22mpoxBk7
y60Hb3FCSiD1F0Vk8WX9jbtHHKJLJhyv1VDmpOdqsNR6fmKDv/z3BGTxory46LHK
ND2PBNnaH54Oede7qghnqaJho8fx1o1ZbCsOeUpTaBHk4ZmrF/YLP1183iEiJV3D
PRy55+rrjNseYHF+lb0vRmSZrrqbqZzj6zDIml0Yujf396fmGSXRt6yYRdDm+4l+
foYAS26tMl5vTnHFwS1RU18pyCWGmZmffSjRbkXKkP8cS8PMlUkJOfqX+GQeFNGe
lE5Gf8KEHOpXtUUl3Hsro6ndm7g3ViAp9oZOk6PJJxBFc6wUIhrFTBC+isoe0QYz
qdOhdNXuHVrYF0AY2igxZmVb4iFAcHJ9KKy+uFXSAKenpcgiZRWF6t4i5Silx0bH
x2GwXHAh29iX6zRw2sOl4H8l51BCJTlcwo0yh36Ygi8wuz815Ba436IIs0jCkK4p
2E8ZBnnthK24w0gdtHx4jiR0NTp5wVa62mOiCbvS0D16r1vXwtZdi5/3HQ0BAjeT
z8gsgOGn90PfeyLiGYoynsROB1e5R5zBAucBla/MKHNf9/+LIngw/kLKxJMrj7WJ
s/jhKIPwwmjBfHju9RHAay6dhVTpJ6NnThukpdily82DYz9dDSOwaOjW5tmoohuK
sNcODAk1yUzwK/NG1BrE8Ddi1Ay6IAoI8QsBDqBYK/jYI1Z1OumQvxvRQZOMgXGO
i3BQTwWXyYG6dl2m1n+QEn2TGJwKSsHeaB31mYI8GkRx5AaX7prgjnzdy5Tqzo1z
3f3GzJaogg7y6XRjpUvVk8pIhPn348Js1gaUQsijiGT6ejC8GtsUQqHZ8dIeEhRC
hoJbOdLU0EfYs65BSqdon/1lLpxB1Jt5gDZkCrqWCiXFThXenzLkvD3QLofDx6Mh
pVKpGUTituw7oSU0MSF3xMWAcAaauosaFM7Z9y7OZHByocPowmnPNbwLHg7x6MCj
Lp0t1TRQzx0OrcDukm5VPSJoC6H+8VSlv6AUhsrf3OcIvI/hyM1XO2Py+rj0hwOE
K/kqfh1RaoHE/sCmS1m/HqXk22BozPtm4sDzUvanBMb+dnB/eim8R5H0vyvUC/S4
cyQKinqSh68qywClZfM3ieUzznLdhux5uMbIjvrq7LQacixatWBOIdivbrvny3zf
9fD7B9tkfudkSx83WUl3jwi8GhEbCeGPM+J9oEGru8N7/gS1TYWEsaK49x8cTuVo
jpTeRhVvI0YLhYlCS4TjERwMxv5psJA64nf2Bj5svRQ6NDGCilLDRq/uwdH5DgVj
vGJ61R8VnChFP4AFzjKKKtgXPtfEZX5nBBtQA8solgozHqQuYtBjFY0HsARSQCmz
ipkHeYsXd0Ytks6ZZaCDtwEjbqSuPjbYJrPu+0P4mhFHoo54C8LlMmWZ3+LCI96h
F84+pZK3joe+OPNn7JoNzWzARXzIIB7EnjhIdx58d1USAXFi3jvPbdPDdl4ALUzQ
n+cQFDQXGHj/lnRLCU8qzyogycczvsF1uaIAb8dhXbWnUWaM4iV34Y691C64iFds
MesqKXSJe7Gm8hupZUgc1ifkg6U0slClWKDf9VbHO5QTg9UDraKypk2a9kKNb+J9
qpkPLiwzNj3zTXXIT95ZPeTdScihEaJ1nVjf8GsbeH1EN3G7FABFZS9VRRjzDeQV
y7kiSWiIH45SXlH/5BQzcicGvbv+hVkqZPSTVqUN+BDU4VEYrkDJiDf6aQRwZvwm
qzhGQHsxyRiTzqwkTKq7qCUyziWQNpsznLlLRRUcSD1UQPpDJKgA7i7V8cUbwylb
yclPBBp9Zwbh72SW7d/5HOoWGC7IUX00MrdWuEhvV47AfK5pkAwGETB5kITPRz84
ErOcBRfsqoiTYv/ARARtER6r8hCo00IpdqwcAqeoLbBQRpCz1XbUg+zDbYFTycBj
Wm5mM0f87enOs4A3YGIpgFHPNWFCuGVOyDNZbhTes75VXAixXH8ISShDyppF4vil
POEvmGClROuzjkqIXBiicdbbmwAeTRjcw2gnrkpns9I8QusO+ae001aof5wcs/XC
ZET/5xujL28Y0PkCd8yrd1KsX03UJi2VEebnSEqnCDH6baw6+K0/AuBc7d7vFxKt
cijETxEk+HxivPDyFrYg5J7fRz8zULPUCNB44XDIjFHbwgDzvgvxxmnaAvRq8oVm
dChAKgHUUwhepEvz1y+cmNYcv3NLxCkb6J4TbnvUWU3xN4kKNAR85d5YL6ipZZLB
ClUsK1aFcGqi+OKQRMPbKngaeTe3waZtNb626y6aSNnztqQErZnjXf2zcFAt7CfS
ZBk3FJ1su+7aL0HLE/vuxIDRZTL3cWSfsopBzOsKgFy794RKpaDJMl+HAkAa4yuN
gAJUPGmQcP8KJb0EVGAxWKvh0/Jydux0e522sNh1YWk8tn1FS/S9RTOyQQD+dsFT
jwTKuchw01RizeuclkPwlKiERgefSHN2lGOzFd2s1OapaKn5QntnY7C1tuHt2pyu
h4JSlqN9lfzSkyfRLUYEeeXsg0B1aeMpdPQzdJLCmY9pBP+dHAwfYPW9OHEuyFS1
dMByL6sFwaVyKGgCHS0/PG+iCqmH/RH2zDAaSn8aXgRXdRolCPvQ1bWq/WJB9bE6
hc2SeemddIqMhGRHtctvQyFBRIpKGzjOctaVglCiKeJcsOxGG/QAk0kLroTm8NMX
gryEsAAPMyD1wuRjsNkpGTXAvVzLjYa5ytO4lU9qhBnPt9Ek/8HyqvYh7pg7tEk+
fu3hnzuXUTCkkr1hiPoxXz7TrMKx/b2otZhdxbEqNaAx3YjGa3eBwRinAkpTJX+p
9sLvaLdOlQlt3j6BxDO0NGgRZl4HavY9zCl1Zu77GQqmtp5SraU9RHRDXhCyqYbc
6a3pvs6yt3tFMCunOJIxjnoXQhPRSmiPGr2czS/cgLYxgoxGJeyO4vxH7+Gv5bq5
ZAkP8OnGLfChA1F3b/jF1v2owAjT0iHPsVf8LdtM/2ittV76THgW7b/TS0kdqV5/
Z2pI2lrrFa51BHND7LBRc+Q32tmVTrJWWtCBCXt6gVDDhz2ALYTtoh2NDwLm/y3D
NdKg2zY1EnmesVjD+Ed/AZlQ1yuN9coyPDR8nWOYb+C66EuGsL/W116V274TJxnE
QEhBfqGY+UCJKZ5Q+3zHr6AznlMySc9idw3XEqqNQwjlKBSbQx+vO7MQnWMeMxEA
W5VDKGNVhtn2VACzFtVKEvNRsJAHMc9ZhjC3VOg7T8r+jZxuutM8tHkxHVmH+808
NxdrI6Kc95ZHwfrtl4z9LcNi+cnMqqOYUCKqacWT544dyEREIYyAR4GDZfONAkaf
zl4Gcdzf9cBzT7VZ69aewQ==
`protect END_PROTECTED
