`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DmYmJTzzdmVmRLpINfAqUzW7551hDMAAeNNFV0OYyr3yWa4hx6LDfIMC1A10b7Jz
d0VRcwlN8Afyn0ZI4hoqfHQfXpN4+TnP8ydlPpKOIqJS4KlPPgnDxkdw51N6TUPX
hrOeACrKg7C7ILhExTPBrgti+bwNK3vE1ITp9kpBj2U/XiBVBx4JRrAB1lSOrCTp
SuLs50/vlr2I8OMyd8qtj9fYX+nL030NNLll5/5Tv7cYc+eSTzyb82SMVHQJvXKk
BBCfvnbjtgCVWvWUN08AL5tZUg5qBfdbUvGp319T0fOLhiFXOkeHMHFLYxdTJB5R
xF4KJ6ER+jOXjP1iONV8BBjQG15BwuPvBTp8EhCY06I6iXTsHZkYvJTuanhhua2T
9LBlHClZdZAu1SLzNtw3AtPijQaGq9ysZA6NkqdI2LgtE2eTVdymgE7UJoVW3fnC
vtokjQeDSP+q1/wU7OPkUG7qhbdXOpuCn6YJ2B0LBcUotNM44We8roMT0puDZRex
1xMRaMz4tYdgF1iT6pdTU6bVZ6Mc/TW//REGPUK+u7wE26b2nOkpuEkTTb9Q7yHX
ZnNs1vhzpR952ZgdZXT9B7/QrKshmslifzTdVUK/s/8=
`protect END_PROTECTED
