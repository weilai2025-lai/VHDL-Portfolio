`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGVEUPdlH6NYnfVW6Cuh7z9gytoy6p3HRRjWXxs8dRsN61oKvt9h9THwSGXUxg5l
C8cdnVZg7FUKH7cY9inv46j/FF+lkTOcYWmD9+RQ50gsfxw2YQQwUyZ7lTY4BExH
jyLdu36hqtMFB6851XXy1IYwyzttVi6dqxTBox9E7WKnBfcgXK3S4AUF3COxEwW8
ue0Xi94Z9jt1qPQrgXiLAb0cD4lXn3E0T9neRt3YtMaJmJKpwIoz1tOvImOm+iG4
wT7pKhQsiD5NWbX7x2qqO4KP3ylFkxNFAOuKNlY2yME7fY5f/3MtCcBQYDNmqZC0
R6ZnR+EhIoCCwnaHfKcRer1qBpizPs7wxkkEdRGbSfv/y93yRSvy5M3lWc2Holjw
4aggL7sAWv2yegi3e3m1i5B+RW0fafGiMd7SQYL/GY9V/nmx+rSq63YyFIwRs0ON
84pDqmDyAnqFqnybHK7wJSv03IG4lsShsbIkdLjPpGs5YtXB+eHZnLq0PBnBCnQL
+b21kEvXKRfDPQUlUWgpeKLYu55p/O7rhgjLEIZj1bktSOl5eR0A9jEZT/ZUdAhf
w3THEvsa+cLDPP5LJ9XIRPeayTfV++2PPKGPkmi6rG5YzTbvTRCECqvSmZKMBOyR
pJ54Md9LoEpxkckvhU8ex3eID+TojBFJ3hp6SN1EwmYAtP6avyQZQ98zBLhafB5J
yHliYtXVhAu0ul8ZIiZ7jA2f3/UzzOqwFcJ3tlscB/Q3tojz0n++SYwhvHmFytoN
9qtqNd8R5MNGYFO1C4DvrPIh2+eIxfZM4v4rUvoVE4LbvH49JNMffccgFVItgYeU
LFIbNwhzvmdpqFZrFrTCztibhd/sI4UZRx1qI5amUYq6wc4AnV1ImI/xr6vmbq0/
vD+Z60fYvow9m/tdva0zHv2qzM/6cT7XWROnSdG7sxzBZ/WhJ0v+TLSHCSwxEw38
uhEQuMFNmGgFmAodrqTop1nPwJo8HQb0kGno0ir7kEl6zNxCTrxPtNKVgHFlUiYV
AepJNNwymVAjDV2awCaw9TRkJkBpeBwJTjLeb9fHa1+XZ19+jmtURjV0DKMeFvHt
W0CcVfAhsVgHwbCUSviA/A+uZ105srG9vHGPGDWESa4xFeAy17CahdkOCzMSaGG5
20ig0zwAicnhuSAxaeQVIOHWW+vxyXnKprSDVcMUDvF68mnj6xbxCeo+iL32Rcjb
pl8p0/RdnThi64ncU0Q3996Q3OtHX9G1Ey0z2LTpHU1/LxpKqpgmHyBIA7PzSpgI
rVLJ8koAdoo1l8npwppNDapc5MOVsKdLH8fEaqKKmeg8JOsELlH8vm3EUY9g7Kyu
bQRjA0mBoNUbbuTXZ83Fx09bGRcq3qy7ofSiNkYSjb7ScZ3AP8g6bFhySmHSxGs3
qhFtvlE0pdsW4h4G8VTRskg15n90NfU16H+Fuo9bL4cCbpO2hjW7217udgdS2Liu
SnbTgKJbjFZdaPkbkN2JRG/RmPpnOdik75qJSjpwW3jhPEpr6LQd0TdPrHaL30bP
OhI9q4HeUt/r7Rhqj34sfmRPZDuxIQbrZd6OdRpK23p7rpxzzJB4djLA49yN6SgG
Wxuy5Z2teYL/C12Fw/DknPfuIbUcAA0oiALyeUInck1vSNjHcafUqI385mvEGmyg
xsN2Dz6wuU75OjSM8dFox81OcJgwOqJ1j+fPFGrKO2gV/C34xpygrIqfKqUQVAOy
3jIlu1jyJO6+5KgKK2e1h5UFBUdrS8iJOdT3dcQazE06bDwUjnBjULJpJ8ejc/t6
1YR0D69H8fCcSv0SkPpC9pr0qb1AKFYPyUJl4+VYh3+kysdFQMNzoj9y++vPX7n7
4jhhRRRUTji40CjBRE4VgW1tFtQ8Ty4f+gYA/LyKa1GhbBMhkqw6mNtz2gIuJXba
nHbbCoyPuO7Ih/OHnje9omOt9BGkNZ9VcWW0a0LmdxcGIQfSz+8kHD0/agMbSNcj
NFLdgZsfZhamBY9zN/LiwUJAwrYu9EyQ7ZDwL4jtOmgIof1svej/T63X8eJIWB2h
kJN2RzIcB0uhFQ3ENG2lXfsqQ4jG8LwfgA1eyDA61+0l0Mr0Hebifbe4O+XnpHCz
W3xSTpPAvseawni0trgcHoXV7jwDxiKhV1r+vAzsQGOMjNs6C+zaxkXRBoixwsFS
/aScvMbxnARtxzVThiISkdu5/JtB2CObzHDHlFh7TXtmoV3L9UJRIzspyub2RtWU
CDkuh5rXpuNinn4R66j9G68bos/ivCUi6cYS/OupL0y4wF8J02o5BCiOBH6uv7Hz
eSxixs0xRRQDcVFfooYeVjdz65SGwIDhvLWq3kwfsPOVGX6ARKxSCvjhAwKFEHpq
oyFyQEabsFiNzX2wj/KRb7hVBRirKmiEMCEWQjU8OkO58EUFej96zLJIqeq+cBqe
C1E88GnXDhJzpOaGV6kaLigk1SGY1c8Oz4UKTnn9Ec5PuUV8EwAly1K/l/Guo+s2
wvBiscvX0jTFHxooQy1DGOfnlPl6y4zlrpC/tnWmC5UKOskhXoDYrjJ3WkhjSEHK
GMbOfdzPtVzHqMGb8eic3D3OiHAhErgU3cum2qNJrnDiNSA74MkwDQ1V3mA9+wpY
lWxjbvTDD2NLbaraByJyJlx9+5s/lm3LVdClAFBLzhw4f5cnxsURAQXbYnzicROW
iZRi7wHZOmVxHmaasG211YzG6izGf9d0gDVG4x7a4iFhyT2Vs6bXCwvy7IRXaZP6
noAcQn4j+SYqdpqBZkU+kbxq2hDntWBPKynR6FEs/0X+KmjwhjLZfI4tLvvLhQ2a
C+iz2lUETEOQDQlmYJj8elaMPq2M0u0ffGceY7W0sRugQkAjo0YCF6DvMDpRxacw
L+GRcL36A5Zq8Y9sQ18KnZ0q8ATZB7a8qMmDq87lpMhHAcdvYOe4RigsuvHOrnz9
8yJoo/tCdQcDTO9l4zoZrKHYdC49Mi3is7FBZNYfFsGtKlwy2MVWqHo6ydOlKmFX
K7PzXjPbFvYJJGzMi41frqPlroKjJTuYWHyDhRZ7mon3kfgAHrLAo+GspKWZRL8B
lwzuYQxdjv0n3HsxLv7vP0NMkaZ4I+7uFPNVSN6C+0XVo81lxgdDuig8AChDD9q8
/oCsdw8dZ6m3BYc0cB693WqJWiHAfSQRzQczxcjukQYwRuLcqnxHQTe5aNuTTjnV
yDJlw+HdvV1b0vSVX8Tou2EG0tfwY/8b5lUcF1puo4p5JIE+qfJLfWn6f0YUWKoq
fOcPep+qaxaSQu7r/m75S/CZHQzScbuB6WyJzB+W4tYUAEOyMGWU/ROslFRuZgCL
GWxLVOmKzIl5LAh+MhCZVdhO/5I5oKnJrXWioFhRMwLVfA/yUHxv+qmU/MCbtp7N
4tg4HYw6Dxe43D4ieyfO3I6uZSbSEhCTtQAQILOtdnYAqAMvzfUwFESSh028eWMU
bWZF4Fs0YO9BIW9BZXKuqLahiiOfJzATXlIUm10FsaZdAniNPq/yE0KsJGn5qZpB
t5EP6Q+qF8ZoHXnvrhwvCReoonzDXE19XfdpZemPs2QNTzRL5XTv1Ax1Gqo/d/4j
A1lsFLSCzlaSUIvKHVi2ahzBbPJP5kaULVtw5KBeo1qeEcvOgA8upaBopddqsfJ0
008vl41l0dkgCTgbkoxQTz2sHZ6Y7gzhFQkngTUw7FbMSym94UIXo9skAqEP1f/m
EYoJIHBLyUef68FYdUHXgp1Hz0Vv5AV1PxqckVnWtmxi2PIoWAjXQEfV5YLBWBYL
ylx21jQjtJpAuQkh9GE59NDv+2rPUYwvGmJa0d66dksU3qsOZvu89NWbyt+e3yBT
UmrGBWNZNVGasfo5rIe7UicoRgx4GBt8Bs9OMClLLm9ozLlI6NbXa9s3b24Sie5p
tiMh/BX0jJCaerIr88o3KmtCw9/malo+8/oKPpH2faxN2QltJA/BCfJOjOGpgZV/
sD/x5LBszM9CjAM8OTGnhIHtda3RcbSgpEOyj1aKocwhOXRuSOym/ECbd7Yl8roV
X+JEnusPC8AbY+sjRaKFSVJNukuJor9hSGfIkxsQ3EkTBIsI3t/HjRUFMaqmgBbC
khWzRBdbMubYZvQ+s69cLm+BqCoH3p2m01+y+itZBVTFkH0Pzt489301ylSixAJs
dhmFU48GRvHSj/nR75Nz5gfujdHFoRKW5DQKvhqMkdMB1ImjeB8taylJ+oLUv9Yv
Q/0MR2Gk23BHGPvuLxMt7UtWpMX2eV+k9SqqFEMbS/peXAuhoZullPr/xgYB8XSZ
V9rQj7qU6PlaWIhrlECN8P3GYV350L/m9xFDATP4voeaECV8z3Y7tlUlCpVLPlDS
G5U0wfyo21RKNrRKTgpyeY0RFhFZmZXqUtDhZfSbtQ723tns3frXH1556YkrSqrx
ONM3kYJHv4Pis7V7sU/zffja3h17dj5vQxfN1DL5cUvX62iuwNeZhkTGVW3lqdkZ
+W7tk7ssxvFRmiLLlD7xWgUEBmHuRT+3s4jA0kKjIodGrC+M0+3FbK6vmrwITHuN
X+nJuBh9YBnqdV+PZfXCZTIWfyXG9BeqJHEIa/vFvwYT7RStf1U+ODAx7DA63tqu
DxOqfPJbbWqmjqQAvoER15fvPPAauSCApW/frmIL4bJMdpGnu2tTjSyCaI2EmW1s
df1JeelAMnrI4OobzMa8RZnuXyAOg8yhOSAn438jd71Ujs0GaeyFhnoIeigt4kWB
83/HoGrnuoUttG52MxfbiaDzCi5erhYxj5XZSQ3HtsksNNqhHv30aZb75r4KF2fo
LFcTlnKKYb25t825Hy3+kcRc+N/DwoZhP8lwPc/INQ+edDjn/UsP1HpYaq/R0uEi
TvouFy1wV4ycXL0lAUqB4QC65hIzC7nlPcvyZI53qwPRRQAtuZnpY1V1HxWG10eV
G4EVme4W+mBW8SnPATYDWe3o/qQAU0vrwl9L/J2M0SipW39orWqSSl7ipyfHmdvb
ZindRQJ31ak81RUWKh7J964RcNUXvO5VNJCjm9+YAzziJe67PgZeW4IySJnZoYDI
T2H0Ai8vcKUZKuZV49Gjv3EEsywIh2E/D2crspZQuEocfJ4KptVeEwDSeq7xpTSv
Rpo7tLkPeeNvWZkntzPLHD+K9vdmbzjsRuklGGIyqK4i/2pAmAIITUHgLka8TKss
aXAe6z9O3XkLRidOCd2r2cJ5qGjbzumXh9cyP3O0OnF4YDvyxzSLTNY1UDBZmYm4
rpox1WvybOnirzRIo5bsZaxbTiUq2b8F7k+32eCNBpDIKzA5+6uO1k4RlAktNDsH
ypOAzCpxEYXjKVfgbpGr+bf7Kv0/sCsYR22M9Nl6IhjI4SY+a8mdM1Vw58uEGmd8
XvHCCD/oFh0nB+g9HXFEnX+eOmKwPwLJoru4KHwXX+b2+6aMIFnZc5fAH2mAfl20
/WDyDIfhcvQqZlKmK46fVmfkLztn0Ej7y28FaJh0mF4RwHSX8LqhYTKSW+C4Kd1X
+iBdHYHLADP8nLKM8IgwpKoaOjTDrq/GfAWWwpU9SBbOGlYx62r+PgZg0o+XJzl6
9POycChpmc5P9ZfJOLu7cXfmb8TKO4PDMEel/Cojm4lTGDCn+h6YXnPyYsH2Ap74
alJVW3DfjrCwZQ7+kVVlp1E8gqO/RAvKauogTb06AdrpSDXtyM+XdmWaRjmLYbYE
J8P5zCrtVD78cETgIQ5cUXv6SxRfpUTo77WYgYUi6wH5LHHFfQWEPKpVkSJb6NXn
c27eYrd87ueNPecmhl1aKVcMulGSkVtjFD2GjLlZOz6hyDAPycoS94JV5PSboVEt
Dli+qBXMp8HCbtJ9FB05aoDZHMGdiptp0qg2dE0tqz17lSep8OcD9Mgp2IG88Hgc
IFkPBp4l0eKKViWVUaorlK2rAkXqif+/esIxScSuJSNxJamNSI14AjRZnzsfUNCh
73uc0UC11AjmqNaSfw0sYVV94falDYZJ7d32v2/PGB8UdbVLvYcR8/R3aRBHmsxb
z8/hCrxIwQJsnDU92b5XbZPgVZCH1Ygef3tyui58ZG3kImabWUcVuWx82RQUJ5Jj
Ax4JyTF2Wk6CZUrRDd8bbATci9bM4BUM6Rq61zNpDU6PU5e7N1Bku9u5xzQ75/NG
l18imKa9BYWgDBj8ZDQXjlmv0eXjDtL6BhlyId/D4smiRy4UOfI8eNukQcvFbEfR
RqVP61JQfR1XJbwwjdDJ5Ef3RmFfrcwjtAct6rNeMQXJgCG0VmVJwBiLJqTUu/ss
tBPSq2EagfwpmONzcCeajOJxnnN9BHef60hzUhN5f549iuSwVPAoEDFYwvCsCFiO
PH+PBlp1/0HVsPcEg3/Sc/Gcj18dDlEhIdvXy9VhirP0N7a4pybbjiug22EIIN8d
sMlGK20Hi4Kg7IrSTu0CvmdooDia/627T/7FSXZeCMXHHtpGRQoG9QJ6Icgs1/Fh
8WDTS6u20v/Zd9u6GvQvVGL3zZUYnqmi1k9hbE6eDb9h4XiaaovXvKhA5kWhHP2a
6Fzo5kTeUTf0c56m60zIvK/+0kMA+L2ePE0vfG8lfOqg5JW9h+aXbNUizXpthyR4
ZUW/46MLd9lvI74OzHrHS+yuquRINVkn1oLscBb8QH5pjA/tNcAtxdX9UsTNWQi3
GEyNiZydysuLynCaiLEEruyRT6YTw0Nl03+uX8EAEQ5VHhuTp1XiejvEil97mQU1
gV0+aHEG3DUbNhZDJtmkvP6iN93IR/3NYAtXZP5RVTzhSfYw3xSR1L9NMrM8Hs8v
okEFQbOm6xQgxqVy1mEN1Cn1rJuafV84dE1XgVHRXkwbv2NCWp0y6/3WBwwxhJ7z
rn43A2Qb4t4w6sZWBEEZ+qZRNeWpKMZVC1YNLlMDwZxqBQmD+7hNl+430eg34ID3
LW4wR5Ds412/h5QmD3865h0JAKoj/UpedvqPT0HEdQVQNI2CgZNOT88YIE9dV5i6
SjiQBivY/iG4IO49vSxl8oCLbP3aOFRt6HS0v1e3fD7rs2XFYRVTfu2xNv2TwWEk
zpecZfWrQTZVZ427zs1aV9AL9IkwP5ZngtKtizpa9iQl4Ot0ajPgEYeWydXXujSx
tWcQXGuvLbRafZ7BzH+MqD9z3t/InPyYJc7SycpbJw4SM4FWtEXNl9ioP7+gE5Py
+EB60pwCGNN/QHesQ8V7JJi93MOWM8dINY0oXNQXytFl18nJEaeawvrrkpTHKnwO
3xYFc+b4qF/uxQHIjztq4VDavNV38CjE7zrX+xC35kai0r+Oe5zFNJuDK738+Cin
e3D+GXXjIc0PykBkyWriOmVMkTWoDk/hYm4cJF3QdJf0faHcawai4WooUbGLhxlC
kApO4zm6Xv77ebwjbIXlMOFaXTVjifIhHTK2+at9N/xdID2cJJPL8947T2vDMgv1
OuEpRO6XZ8Mlogl7BIqXwxwZbdByCDK5BJA+yMw3NYEwHOZxk9hBgNsdvjmFZMxU
rt5kWSrTgFi/8hWmDueut25joZfzFqUSr4UofZNSbkmjRIDUAoLPKfi/pgaJ/XUO
wBpFbH6frvwmAfDYLnWimZDOkOtIXKTL/871dBX4eqNhgLTFbJIeN0QbPTiNFx3x
F9UJBIgQCodWInkCcsILNU+B9IiWkCV2ZV9GbksUVT1lbOkukkEH61nkrF3htOFr
MGNhZA/qLmaaSIxE0dg3/KhR5a2+kkwSQOPwsnl5/7lZNk5Exq63JOYaazECs+4k
tLwyDHPrcM7nKNjvpR3Qsak2KF9J+GwmZ/Fo7MroHoKNLHYtdVW2JmpzDROHrH2b
QfN3EDehsHJRfj60EhxNTLwUCYkqFz5VPF7bXpJSuto8yZ2CMAMhtBrznaRxLCo2
YcwVzHF8UVGgAKSAZQ0LgqG79JT7MauRJaJ4YjHcPaUD2fDEH3ZjHY2/80b87i0g
ZFuwRJbWLE1v6io7evyxfUWhCNua6BBVDs8FOMtDucfGH7G7bmKDGrZQ+NNaiG+Q
D5xvb/vNbWmL41MWhwzWJfQi4gf5gIeOv0u13VCCEiLaNx2l65bbLUnhruR9geH2
v9e90sd0s/NVn93IpsWlYtgzTmHKrIMAzvxTyL2Nz6hKVqvau0iPnGfGvBjp5LxN
xFlvHIG4WEUg816+t9EkqZP6u0xRsqdJIC220/EZCf1KMKkhZF537+37DqpJYPb+
ff3zCEp4xQ/++M5M5Ikie2rDk8fYbBjlgXW85U3j7aGQEfFy2Si0h0bjXgcndwdP
t14dY+z1r/IaekenJVES1TnBPZovC4zLtiWscmHofb4xlXubUhC6UJf19L3y4O2o
5SzmulRODY13r6qaxGlyfo+C31ZwChWjHr1WEZltFB6o7o+9ynQfOSHJOQzuJY2H
X60bTi8dMlVE4FIen5H/zzXuIDlBFw4srFSzEZobllrIkavw8rWeuHGwl286ueth
5FTIEu9Gr/3nfICk7wXYcXLfmGKIgTpzdvMLmR3ocllZZkiecJAG9/4o0ArzFavm
gEUSiJqlL0a4txfbetAK/EATWY9dqEbIqa1U7zQZXWwaFcrQaURSt/GNlaeoY4yV
J5O0+9VpZardlwiypMUfOqyih8MlY5Z1A1JmDf/KmFZTMtDwimrCBH5c/kWfNEfv
13ray1rtJ46QybB39xtZ0nqIrWdHg5CmP0+Wql2o2LRRNJF3k6wCbch+B2wBd/9q
K/r2+X0vd0OuzOF1gF0fYP9ZsZfpKgH92+N4YDh0KZmJLvDrWAg9tBHuHKJNuRKn
CsLHNn65d0Ta+PilCjA/nI30KrIXHZdfCMfWDOKX6UOgtUl50zaX7LLiv1J4ZQTZ
wDLiIV2pVgH7oKmJ7qWU2UCwURsIN7MLnbrpJ+hxXwQBwQwn07whATVf7BUe9iAL
QE81jFKLFuVlTBKZG1W1oWV7CB/P/MftXiPctYVbpr0heCPQ3SnFfB0fL+J6QR0v
ewpIYtZ31YgEl+DPrr25TPq7nE/ku+HxaC5lRslulvQIDNXiRmxQii9cG7O2h72j
NLok4ZJ8KCgJsjH79t7TwG4jGDsQlJVMP40ikSlCJ/pt3BCHMv4SpfKE1mFIOZwH
8Gi8pnCLHT+6meFyTSoVSjV4hhHeciZR62xmxOO63QlzpVOSv/pVleUhhYnAO0Ke
JTWMG3TBvbmuIzOg2212mp7Q5fyqg9rJys7LJt0aHHUlY4WajwBRd9CkDmv/FSWi
21uzqMShjdMso0vGWKRgE9UVz7NDIer5s+UmiBBQ8JzCx2koTXxW/O8sB88cwB5E
FN5eRxqAiOEMHZmrywJX53CzpyrMm6N+BMo8EZmciLTdy6fdf1LVFEEbSrwzPgL0
UuOZ2lPVJoTbU2uGVCG+yaaAGzHG2sTJ+qyC6+GdJrsVJwblnne4uFLa9v+F5/ll
MCaz5sm3JCGyWt36iagaVUYY/hv6aJqsgKRRbj8mxMb2zlYYE69bIZ3J+ykdxNtZ
PUQ/JE3UpeRhGsSlWAkYazM5lt7Q6uSTP2T4BVCBpT1D6raC9iChNAQ/UuZGPJKJ
wJBkpfWqjD+kzC8gi2cCvXD0oVBXJLhF+7rPYMS/jNI78uXI3zwmJSTlI4D4zkLH
9tiWZpaA1OmTrypTdn60eRiJfBtMxSo92uP2k8jfzACt4mp+JkG2agXZnWWoqrJS
APWRX0oiIb3KzzVaSrMtU4H0+i4P5qZIirCUa47zG1fdEzZ4W8lvuyVV9NhXZ9Ml
mcBtzRklJRbbIwFvXK9ucU8r/futjxeXZyDF6MTQfS+S5VgJdc2RPcW87UUCmNFg
Ps7JTg4lW+Ml9yljnx6K9aDIXiahsiov1U0Kch4kfSb9vfHvAaLMJdY0V7Igu7hn
2nxoRnjr5dFxywP4Ed/prgxVx09WmqSFHOnUtLjzi4zOfFt+E60PFoWssF1pjaia
iKNGSpq/S7Awgo4beBmpQcD5p7Sf1uVPpIwYWXSZH3/+bu7ramdbMH3qc6GwmO1m
iZYwdlx53DaB/JA1EO/ojXxilhWgElJ/T2ZcI/FcqfVX4F4GzB2s4mmrBkUpc0SX
X/OkW8PHyv+nPu0+1ugi19DE6YjfG1OA3TqA0cWa30qF6mPE+5wIYNrx1IB0yTSg
2qoMStiB99KDxK8y7tBUheZV+43PkQSb1YvHd5KRicvCT5aUNA7EX0vEEFFpDlli
GfT36u7WpLBSZOwyres5cybyL00Daqxy4TnZBsg3UWwSD0cg5gU5OLFgcQ+5YOE7
hirHWyXCEk8VRD2J+QlC+d+Oh3uRf1mdFQJTbWkE3yX3c2QwaX+FovjTngIgwxNx
h45RKa2+d+51YE6jkVn6yJERYFFPN87Z7Hpad7doqJ4uOqs+A8kxar7FFMkXaJ5R
a5ue5n6h7Z6TlGk2VY/R0rzhsTKwb9PAfhTTV3XDckXRHJKBLX7YrJ+JtXhNR8cU
5nGVL6XI5gZTbbx53EcKqCZSeYKv7V1/NYZpl0xAflwKLtKDEiymFJHcd03BoWjH
kzKrEvNKtT8buxz7S4c4cv7cjs1h2ecwULCkHxoeEFJ4BG8yQiIrOg7A8rfcRSV8
GC4KgzS1WLu126u5bOhGHU3C7zwKoZQwiqyfgeRtqIs1Ff58XpVC5MZiCwnoa4IM
duyO1nPybXfgXqjxHeQwSyf1FDUarbeZlZb84YwWMJSrncrzoUNiWXB9cyJjdBXL
0WaBHezKsYTICci/btJeoEFz2LUG2yMh7/XzI8ahirL7+h1PxcNv1/dPRQCZyiGv
SmSaQIvbBX8eu9Pnp3Cpq9s2+HSnGBc/xjEE1xeRNi3ej2FmTcSkrCz/S52Odg5M
k8CRrcCCbNJ1nPFMVt4gQAT2lsUjz2Z8YUXJYTR9KP9F5u2FQXGa/PE8ckKh1ISY
w60kyj/BJvWz81Nzys8bgGUqzadMCuq19iq4rnf7vWC11X2zdnWJx9sYi1peZijM
f95FGveKcOLF78SBN2aB7oa5IJ4fzjur6Lm/+/qzGXoJjan49swXTCstbQtBpJhQ
tFksOMJaI7czKRCB1H9oTHR6HOe3uUpU4hGObKGwPxVK3UEkEUNNwtxxo6aOPNG0
+9ia/QWZFBsfSWU8FvujR5wWGduF0m+XH7RgQ+0ewqYrDSgqAbBg+dZXSdKnsk6U
JW/Ce/KOPATgxiCHoK2CA8L1tR5NNlf+W8x/vSxJA172Q3y//5L9CebVDBeKegG+
yrTLKNF7FSJCkVYGfqsur0pMMMv75wbKY8PA4c7x/q1sodbzycpw0MSPigdn4tMI
+E2uDyZtewH/3ndZxw5QhkVcHkFxfloozguxmvW6YTMPocfXBeaGo/wdc0yIPSP2
N/qqRnkhqadgBhYfAISRU9cuKcK/havJbD34refGGNwkiaiPct/AqSXHwYHQgKtf
nzJwa8ds8MHE5QHLF/nWs2niDqOdE1Cds+c0pJhOEMnWKjUkFQTDYIVQCC1FMZbB
pkseAw+ygVLaJ2f1BpW3HL1+veHQCduRxS67U9I7bThOlUDfo2g05fjwlT/o5+Rv
kTF1EvR8wC9+y1CXVqdNSv1CUwPXsK6nMV74BzRpPcnCH+B128r2iPg/W/9pPphy
alaMYyyWkmpm/Emj95lkZCLIMtMip7dJprFQHQHz8Rdl2DgEuFhgfts7BO7BGu7I
NRAYhYd6fn3gZpZv7wDXOOX21qrLH1rCGy19qKHMaskU6XKhbCosYjV5nd8hANgD
uZPCjtdw9auLRbfoGtjy2Tk8Kt5r/yPJZkzo+Q0yzbLtNfJk6L3Rgce+J1PaiGhj
Hz+Y0EVO39G9ahb01bx1uwahw2gOOvCR+Goa2DxavzjQnUTt+LAZC04BVYmksSpe
j4kpRm22e8fHei7kWwUTVtx3gasGhj07Pn578JBy82+Oc0Vf4pqzL+OyLHIGJTsW
/IbW+0inCk8ZiRaTE53d9t8gdfl8/rHAu8ilg9+wEYlWM04HDQeMeHElTNdN70yB
CbJK6fTh7uUFo2UwLN31GyOR0vQD/fMKfgKARynn8rx+XuNjDlMkfexdE9xGXe+3
CjLJMoGCgaHwJmikqjSSmLaH93P25HhjYZwrTTOVDK2UqAKXQHZWEoCpvnCvE/bH
PbtC2wEt96dLCwlNKVK3zm5/v6sODGwcFOwEzmLTUt6vRiUAmzSRjhNYht6AsiXc
hTlg8SwhUs+vezRR11bR+ncEhKEeI9nqDTMwSzhgXvQ1cfrm4wWWx6pyeWnG0ovX
GP8FJLNWtyNMTIZC5jDesnilogrYjmTnAg1h/iWkb7UTv2j3RJE8M556vBMHlgfC
5libCgM9NbgOHm6cizdNbZeQKO/aC8CxLErVCvXGIl+BWib1rQypw32nskQRXT61
ERZHEtOcTjwZCltk6rzZqwhj3QbZE8C2kJWkbuWg67PXBL9rMlNdaYB2NuoqyMIl
p0m2G+j6EhRA2azD+3JpAJQCAuXZD41vbDoCTZPeICaRDSiJFUAuH+HUAnpI0D9j
hUKEdNZV6JkiQHBb/qWiiH9ezix/3KDs6xPl3vLkACQv3Qkm4N93FOLqeQKkUrH0
OFFEWByBMvQ9Asr/xkUEVg3OBaeWSpFtapR+buWsLKTmCcgyV7FNAUwE6tFJ3Sqa
0rYJnLPZD4w+1awmZNDVeMHseYczt1r+M8yJtoVDZxeohcT3ZBfYod0fuJ2uWsvr
8aiIwlu6BZq/1xgs1JK4qiOig7sJTf4pFhr5imEYtxyFBW/vsM4gIAQ7venndkxr
rxcelt4Oef8hZ3Rcub+Dcz5DEnqGNi142Ns/muCD5o6PTSIDeEp/LKuI156B3jOH
2abkB7SSTXqvvmuS6+MJGujSF9j1lAY/9MJNV/3skt66mcSE7Q92wW1O3AAbPwco
WrPJe23lsurP20wwd938FcWo65qBAwhFhk/I0MAZmUHAciIMGIqkkQRRPZfDort+
jtrXfXMzlYN1hVuhod45Ir1+lUPJiNgKVDVoA6e44C4pdg94OLbPLb1XjCXFGjrE
6VtFyYOtk4xqcSSbU+tsVRUSJCcoNx0bx8/X+e+CuSXF2vnmNGf55fDNqlfo+6rZ
HGnAxGL9qEy7UB3i0yApUB7qEfQNtEv59v1ZGgQx3gpmyyzC1xG6U8lGQaH2/vlK
8U5Mz/aFuf1CeSW2PZ1iKj6AvBOCHOhNmI5f837PuArSIshs8cII0634hrQpXgFj
0AbVpsjSOUsEf0hl7w/KXBIwDcdvxuy/Ue6iiI6l7ojECfb8PZAayYBirmch7LXp
0Pks1HJFJLIIPY226EEXb3j+jj6sEd4IukFRf7q5XS6bLqwY7kPdwOvNCdceGTIO
tS/sxBcbQ3WgvZv6PORMdPDGX232lz4e0xrNjDx73xC7Uj8luDRbTXSK02/sCFr5
rnAIS09XyTFyufevn7Clsy91nu9e1q7GxwVy0EzZHp3ZlJxLn6BbctYCLkM+/8jb
Ky6d5LVGaQfM0y0HdwcP50WN+eqi6e7YzSniwuwdK6vUe/oRW/Q5ikPJkAZpcpL/
I2t3tSeNXHUFT8Qhe/VVoelJlIM9qqjWmvdA/1f25oGVK5ppamRNvSqXNRc3oO1k
0P4h9xnrUwvSKfsHx0SuzcOqGuAadK4V1WGJYLcYHn3wraMMTzOYcIHh2mvZBw45
CQLDL8F9UAbeBrJqwclf0sPKoQBlUHw4GHZISZhnaV1TuIc0dJO4KJ7dLLFTdwYD
7VDQwLOuOQdw9aLO897rnugdT7cNidTbQGN2rvxCwLuWHud9phZlh1zIGPgSFaKl
avnrLhAM8KRyHcaBDVw1YjigQii1i1JdDQRD9dlNUZ6jWr5ZJBo0/ctAflj1ntPU
bpaoO1sYyQX5gqkkp+SkQ1EwletxgXyTyV97Op5G9cGPe8fLMIGxcfPJIEPi+Mjs
KQSL8dOMsy5H2RX5SOLMYb6eWwS3ktUc8EoISUTIvKz99m0cfIANn/laxYXavG6L
x/PNI19eydQ/o7jp8deQ73yiix7WB+a++Wi9Q3m6AldXs6SFPROuga1vW65qDlLJ
l+eyjdLWSR1bmF+gxkVdJ0Uh5xHwx2OSkipGdZijzLGTPXhyVrDn1to5k3BFD6Dn
TM8exicIIcg7QY87KMeitqlPR3/YBCwbRGU+jKNoxs0B34U/nL9bzrWw5CCWMf5S
jpR3xpGbkCp+OTJ8qNzc8Zbv54+oKWnCVdHCIy+CYeKB5o4TfaJ6muzyK7rCNSJT
tjOFsNwm5kbTg9zX1LxYeLrc3isSMVuNylhvsGQjzumNiqpa/0Go+agaswC0jILd
h+RBAkOO08N6L5ajaDkOXhp/IebzupvzDN1a87ty2pUaLHFGQdluEAIp2W8Y1khm
0607zHyWHMdOFKh1oGZE303fE2ga90GaUXIC8iqJ4gjav5zT2d7ptFuB12OY2VnF
aro7+ECIlQA0hSRcLeC03D2Gz0daDehXu6VQ9hYNsAwS64KfHYPic8D7WlmIXn38
rXJxYGNSNZHQ0ob2D1H1y87ZCIbBSbhuPyhSqxcicLyuULmaC56z2rP9YchxstPz
SRHpGXS+I35+W2wE2j6gvUS1BBzsjcPrI9J288T+1sLMnAJvo8Ebd5dtuMN84WpH
jUMU4Lp6UMN8SDY6j+vBiM4vfxlaV4jazZykldcdAtZHwSzShth8Mssm9OXp0suK
jTbPIl7lVRyYCUkOxcLnuIg+kIB2haHASIESE9d2YyOZ+sdZGzRM3mkbX86UbtuL
cUtxASWTtgWUw7868mPpuKZR0gmx4WK5Uxoik3m0JtxLcWlctfPTv0wPmao8vDRd
eJ8XIEAtmQ/N3/WbuhmLPDN+BltmuQKW5zH2a8tgRgXfASrknrj5G5GPskhu1cxN
7LRJbVerxJEM+mclxQBq/ZU9eauB8G93yTK/kxLHrnhLl7l2mfcb61KCjVuqixpv
aljOXZt822mvYJi7uBqBIVI998HMenCsNXFea7SfT26uRM8g00Pi8JoGz74GR1hc
u0AeT/W6WPorfddJJTTl9Yd671UfAqwGkP6dbZrURuaSPdLyPi1FXB/DlAV6rdar
baTOC7C1L45Tnu3+LpfKKpH3uz/2LYgbz2F8bcKPkZfbCf+puG+BChZ2aAsdk5vr
TyRFyQ9eDH5g2VIezRl+vqA15EG3BvCdicjSoX9rfcoHrOSeVFiRUOtoRd2OHuxo
QZQrZ9q6dvW7RBnBpRkeUo7oJKJj91BWlS3X1BHkAE4Ehuz9LWJfytGHLLJL+SX5
q3tXE+OIVG5QzGu8wegT3TuORe4DzucxifvYJFWDu1Cd0q/xOLTjfm7w2lDaFawt
RiZh/Iz0gj2gZxo+IB93OLQXSR4glbGUK4h6+mE0TnmnY1st4eBB16DCLrQZM1Sc
2nHLGmUz37tyzwU7QPJhDSt9MBWhRNWMvXYKUEUvSSJjvRMrYltidtV7Bns+Hf/f
Ut8TeTjx875diW9kDSYQGSORGdCwxZFT38XrFxjeHzG7RAC7CAZpc0xglXbSCApQ
Na4no23eAv3x4LJcS/s4pcwQswOLDwHotDQnPgAtdXkFF0tJnqAJYyVhkYpFLFmx
tyfz6YZu2+543qNnyHHCVCnHDwzOoFSvDKWMVQ7qtSoZkfJPbWnqPdX/bO+uQfz7
jsF0DMR4q3R99/yh+L/403W1CiGsHkCxfUiUhpKTCOUGnEZk1VwBZLkYYIlpPxBq
lzIja2/pRplxbSmPTfeGUGnDtfzbUbbSI1YCVnkzc5VGXECwbAMO8c0TGWjzEpCj
LRWM3uq5WENk4GvReqnI5db4DFE03bTbP6JLDtG0yjumjmWsBQIM9C8rIDTqPEQ6
mdy7v8DWbr8hpWzx6+NwPVP6nyeRuZJum+Y2cN9+6ymmj+n/zHYO+lNsyjwXPtlz
xkXu99clZHs5EZYGXYEhk3+CxW1at0FxfeCwx3qoRIehhwqvQR5+h0HiRKnFAJcW
WT26DjwzWD/uaP6XR1/67EixOpqirzxpFGbMueBEm5Q4weQ4XPlLxQXg7IgCnfO0
jeqcpIRwjK7Jvpnd8GlNKbMekwLCtUREfsRhonUxOWCu+ONniLVSsWurnokDSh6C
qogJ/Lc/s4uCOU4q0ALTR62/DTB/HkqEIJjLrAoc0h135VpLiMFOXUn8HMLv9W6b
16KDJVWZVFLtX4TRD9IN16IF0wR1vu2vFHEKZ1wESZm8FgIaRa+z6G9d/RO8oxKm
2PjEjaBdirFoTRt7L9cE6XsW2/n04yh7oPR8RxrKTs+u9ZqLijco/8VcOq8IInG/
/EWCrkY8AsEZukWz1qqC9rl9WxTn6HdO1dbTE0C4F1bFDb45T5Y2B4uRdG6jCaE7
iXiPi9+hhney5POpIDM0psO6RZFsIRflw799abqplpQaKE+Iehu/MBvJFy0RUrG+
0OgY5WoaNvMmlpOP2JkMJ7L7GyWNKFrpy9zplAXyy/RNDMrNFnlosQ5F2cIIdDy1
ErLfuTl3oZeTH/dxj6UMU9wPydCkFoOmLv7Dbh5hmyZGKDUhnOa3Nsu2q6zte5aF
p6F3wNnY6KTXKaFc4u08omtd4nvIrxChLtdVsCy0HBwSjpY46+r/SCKFH4thYZj8
N3cMe0fpvAyQAYjcgdWO4+Eexjl/pqEh3rXVXPk9mk61NMOyVsXnaMsGklZNkNti
JKBCcIScTCidxYgVRDqtUs+9qBYYsO9Ep5jccknmWkhtnTIV823PoiUg7nulHgHf
NhY7QT4LcOAImN8KMlwDe74f57gKEwr2UsTYNNEFp7iU1Hqm/JlA+987TQ2vVcYT
LxayFRRKNGADjXHsJc7jTGK3F52Wox0rVxDEIgqlVGWtMrTL8xPVEIzKXSePXdi+
Z5bFY2IJ22i3iL8pICKI61djl/Ln2ygBSTRAqLHgtGjyTGPO5ctl0Ac0rf3HjPan
5BPMErujbi1FS8gPV/JzrVMBI0rUhH8Q3R2G7cRR2g9+RLxXqYEDcnETJFy56byi
4jLF2FmhesyRB5g/3ss/wDBrTZo9vhCELdC2Z5YY80pQTueHkpVQ6FfEwTXWyQuA
vGFXLCH3Nx25jqz9vAOzYcdN3Tp6d6TeYdQr7KTvJt4cdLMVOUiyFWDLMLXwceZJ
V0bxZkZJSA3hltri1/McoVDH5srl1Ni6tBmYInRJabgvy10ecwa9RXRj3zUrAfj5
v+lUAwUhxj18dI/38Zm2Pjf8NpVlxbQC3/1sIEn22meuWTxQEWMyeVJ2BylNFsAA
fZRZ/EblrmIq5F3xxoMXzdnccHfW/GpwLcCs4rDfNn3eMQ+6KtHkc25HliXTVdvs
lBBfuS60AT4cswITBTtE4FZK6c9QQjw+s1jYMpwZOth8DVlxrNG09O+mVPjy9EAs
c+w7+ZiPWCaHZLrUKsBD4q3G6M+4PF27acSzmjZD0e9J2Pm4khtrKU3PXTPdDEUS
IVw3iu7qNWrNUjirqernk+BJNEtjawwY/Nyjhrh8gWtA4iCdsBq+YNppoJ/CK1kX
A7dQajJummfw4t2BIk5vFzybo+fQpnCmvaoyeA0CgW1ztqkDxViuQFgQpaQyen/Z
S84+mET1Z63pkk3skS4uTJnxmM+jPF8VcthdMhVedzaNtEpPqr3VTfmUK+iT4QKZ
ItTzKDLQsqMaCKk9gvt+MCWoul47RebNwQk2IXogkBq78sWSs+gjEHKboSWdo6j2
M1F0OZ1B58mbJ17IFqEdJrjIFmZKzJTrBBVfpRdUFslUw4/PT3wpTOYwfAAgJGG2
3leQ1oHTuKhiWY05n4ifbERTcx82P6L+mQnn1LhKuI92PoIKIl4GQGqILyGO4VzS
KRGe5RqL9gWV6QUVyNluAyhdTLMj0Y0OXkH98HPdSMASCow7ix9Cfi8KZ61DprWg
PmBfSc3uTBiIGoTYVcZIiE5JSMaNj+vsO/ipstM8LcsTvDrshubYWCydo/9Mf39C
LpDsohq288J9Lxd3iODODlboteORMdk5c8DWK3HFhmqqFWI6rYIkQLwLmtoWOFyv
JzD2PWc3CWCjPa1ntvas2enyJtdtQRRoW7NY3qBN+zzygiP9CfnZp2ohNkPP0SlX
iYWLAnq2xtVCsEvipK6kYjmSG0Su4BLUitSnIZyJbVWY60cuRQYBdEdKDykHYdB5
J5+OhrnHCdNlWM/fxcwROoGGHFr7h+YixrkM2qzaoDc1E4yYX0HVq5hesML3QcO4
fEGYgxG6Wu5W1Xlau165Vn57bTJkNtNNzVx/4hoeI41iWmbbyC90irtLkrWoMSjv
UX1VnYlacHIj47GnqvgWCLlpnmSu/6Q+PePl5dOnv+/995cdNIVlS3rti6WYQwMH
tPOkDtmR86+pNgfjtsxxC/lgSnbDvypaUSytPM7ptAzL3FWofN6Ge+FiRvP4nYO7
nKbUU8tg52pqGEHamT3X/VGMreBbfzE+aPl25q2RMAzHrKYU64hL/w+jcff02t0w
WbEIvL5httfgB7zp1G1F92jy2sqlKQXNe0oX/6hYAmFOI6OGsnPDqgbMUKfcL+TT
5Yzgzg7Tal70qnIitqfzJrhM5k4W+UaAapvgnH2oKBrAKblz20The+Eh8Meq+sM+
4eGOA6Up2taZGWq1cZ7yvTbdmCmsb/fIx9nNGif6xA2jP/Fb6Z+VulpWSbe2RHft
iZ6o9Al3SUupCkOCe9cXxSSexKSifiIaWECZgiDSyyqQ9XXH8diMDjbUOeXX8353
p0FwewA7xOvHgIQJT6B0+j30LoOACJ7Ooie2Sj1jcVJzJebwMFGJpwiu8+1+xWWI
pqLLbtF7KhlOWb/EgqE6GuiDywZuMZ3ic98mChlq8ScAkVqNQ7GeIb9/4H3QV53l
y94pFYJvzqsdfP8C7oVl+J46bCWwHO5HIOeaImK1vS3ci8JebV6+MxT3rZ6oP1/i
cYYt+wTxGAB64+PTGwe6isWtDlhVc4VlaudozmKkoeMJe+TezbRkcVjNouzGDDMS
6b5S2oTqnXQa5l7BTs8pLs4hZjHSSXskhbNSK1LrbkuiOmSB5aN3MvezkEZxyYPM
Z8JL4duxNP16SyoAWviszskSFvwaYosUqskW5VNJxvGlQpHMiMsENQH4vJWoJfy7
Eb8aH8M/xUwQ3Vy/aNCHEJc2HGKI7SVS5duTFkj2LSIbqegcHZ/kfIWSwsYUS5IX
4brjI9tHzlkiPD1Fgwx/ls1dkvMabmmjiBXBFeTbnFOP/Dttt/Bh4wce/3Sb7zbc
TRFTiY56UiL2kQNxWSLuyhvNr4phAtVGuebEtxUefQLtunDUg7iHzpu/4vqjCfGO
CJRhI/NN9MxvZA4HJjRsUsBn+KC8JdE5PYBNXhd1SPlkn/mXk+x0Az8expf8u71U
80/wZLTQ1EEv/IH1HUIZdwoMarjblq688X0xWOO40OuOzGpdDs5N0JNXFSnBnNCC
37xd9d2FTBXtdGLof3XhjzEPEWpDSD2KigOjl2sPyMP247JdB3Yc33vNcmKipLj2
rFp+hqxbjWaq72T4IAzbZ9kEpnSJX/CPM/nSHD+BMFCiKnTbRQ/z/uXcOXNR1/5w
xY1ungY4JRa/0Z1uZeJZnoT+dpBV0l7RHSJLG+bwXbZqFrCjUbC0maCnyEN7KNz3
GVj8fS9C5IXLJfnIlZDcyU2t2WHLW4U8aaRMpPYcnot9lkFxyFmeAvN14RHfte1y
+I1tAQebMnjzPjiLfKEi9r86AWa6wFJwbpeau/pcnTpeCNp54mhva6TBAlu4Wa5p
xJSIk3YCQxLm0/oj2dPIn4/iDYYn845TWglYNu9ri+z7vTdVp4NQkW8yYEhMnHBR
AL+vgaQjFP7p+VdyEDf/cTscJOqKbN2NlXFrw1lHCuD4W9O80i/QlmjMcYOra4GD
Yes/j9HjMUc7VEDn5DKANytxjxnX1FyZ2GzQggfd7lZWTTLS5m6DUHExfO170m7H
BU0PWThKmps7wklu+84lFqdOOcBmV/LwcoYy6o3EjHYiZhj1Gufzgy1NreJhGqYy
tCDLhRULvY8zhEQBGbNbnuig82TSDEGIJdzttNg5GKP6MtTwr72hkSsM5cNvo8Xk
hB6ZI/xoD/Q64eCvV37pwTLq73+Nm28v7CkJpxFuIbtiLIbnqQIpmtXtlZXuweiB
HktpW2eNluwj8++GBfXFmlnzv0L8HaFa59xnRBtw8veaf1QGFkPnlX1i2srVB2rZ
vS7lBkKEnxBIFA7UPJjVtpyGVMxr1s3bJUKHDwvv/EwodL6+SpBBRdh+0p4Luq3T
TJHUzHwV4mmp8moyskVonvCciaQM6YPYNp3X5TzqRpimnYkrgLFeVPAVp+phRSqP
tgRT58sayzM6ca1ZNro7g2YeZiJzogZ1skWontBxn9rPCnTmMJc4YY5pbAypWIVX
5MIjIs6IYOe8riWzPKQcmYjA6sUl6OuyoMsTnV8pZNSPZWtJXYRuI598JFZ9T9qE
JqYZdUvHteVMyyIdpWYDrs3sFPKj4XvXNkBl56/LHsuieG04HVLykRS9vhZdR6/j
Yy/rW3VHebmjBCWAFf/vtsdMDo9J5ene5oxC3W7rHGwIMHx9tQgkFbBZ3zH7zdcS
NF1g3UxQAbsUQNA/mBOGxAWYjXuknQZLdwY2Sk30yOIEsDZY1fRpWCkXGONiD3H8
R4oqU3ECCzHs6YIviWdPB+aqjxtunf5SVVxiCGzDdnwSuBbHArM4tpCK5/B3alOh
ZF7ZwMdsGttY6UdT+uIHhIYqudBlSiZDYwTXkBxCl8sX5KKUzzu01LRzK7BQ9TQz
2w653x5Bck5o8fvY3VKhj2i3f1d3VyLyW7emPOOFzLAn/2nUHFxn9tHSAwa9R7KB
SmrEp+tSsv7FbT1dLyR/qiX9CHYU8UbAcycG5FLaAl2eQ5jfbMor37jQBlZeHLos
08ARd4FUWoUNeDSDjQc2GiOs7sh3RhzGMYIQXFW/Mjm5pK2JUSSgf2RZN4saKo5L
pOW0f1R7VHn61RSePIRak0r4XwDgyMjvQfR8sxpvt8jfqZeccSdQbb7NVYS1MOq9
XhsHwoctzUBWsROY7tHJhGFwOqN6drXd9QhDYyhskL+Cagrbjryujsi2f7ZIichJ
l1qgNbq1Q5Qpf0vdOviFKJUs2+wRKqcWsPv4Y/Mym2+kfd0z9KjrUg3oIPuX2Sck
Up8ur0kfvxNWq+l/I366XlPUTkmkxTmJY59GrEKCkxdCO0ejZqfKgG1d6AaliHbI
8j9Ket5dn2BvgSzcH97rKUSJp7Sb0l2g7BAspbMYbejySo4Tsv4JUt/3zOlz86K6
ThYLNEgozwkLO9u0FnEc7I4J2u1+oCKNcz4WVa++17CVZrilxe7QFiWI8Gh/FYqT
q+8fNTk1Rz8tM7mqCTm3Vcwgb8qItmyCYa5FSL17FrxYJ76d7RW64ps6Enihss16
xUZ05nCJoLmY3wzj1Nw+n3ZTRTvcJuPQKNEDottlaZbsam7CLXmJX7UtkvxkW8Fs
3fbAYTZXl6kwVqHllUTPoR4PQJyVTzDim4ssW6zuFnGl1MsUm3W1Ki/dKf2jzp5+
3q5hhgGjhmnCVG7pvRK/+uSb9ZTAo8g0QvZEs7aoTqOlDl9W8MMfAKBrYa2/JeO1
qGBKT9HiIrc6poqkiYknKjm5H8GsZIvlWaRKz66OUEXcGnyw7BMfI2I+C3MIH/X7
mbLYOi0Hw1Y2n9D7rYiPFMHsfx6YMREUL7ueIJGq1ujMeHlBUigFVJOWepNMXrg2
riZl7LW2A40vCAHtRTFg9xal/QeMhvXgTmEUFgVG+iZCbEF309PFrxv9L+tr0N4k
c2NAywUbzrXk1oeHFDDDTg582v+1WQQohaepKqGuIBOWoGiENAk6IWEb1dL5LUv9
TsZTjL14znnUhSelmDCzrYzil3o+sWM+1vZ33zQ6bRWxhLcpahXOes7XBlrUmlmX
p6DtCwttMoXp2YuXKYWRpnpVlYZVCoB57v3PTLdBq63xmclLxXDcaB3UQc0+J4zA
7ktN4kt10BQreckY+1g0/1RY1JF2AC/9awrOq45dFSe3quIt/rdl0V905a86zSCU
TvIZ4i5K7lo3sjepahGnIydxhzlPAv0polFXe6FEEQJHQ5fajuyB3E6b6P08DO6G
z5xIPGXclpx6TDGdrfHrPAxRKQZ/GV0QsXVt4FrXs/RtYQDUeb4V+OllcP/Itg+p
XADdjdRepkVv5pPw/kRGuohWf3CpltNPhprQvwpqNV3aYNXj2s/RojqrNSQ9wYQp
ZUgXobZz3TU6GEHylBRy9M9b+f4vKHpqMZrvGzlSFam4zfarN5yCMadzxqEIXxIP
XvjIRRLDwSZPGEBMHY3YK21C/xJEy6HJ3FrIgNpecUS1aaX9OXWgHk8k6GUvmBMS
VDzHIgCxBL78MwRzBjxDjmDA8oVaRLBEVQrIThLSC03jsj2kEZbudw/WP0Pc2i/Q
uXkLRB86OHGIVHW8j8UHlcEU88TT+eVxPMNTGMHGyxata8UN2F0ULBs32LEWnNZZ
4apyBOtolJ1nVAUHIewivaCBgMylWV88AzA51vl3NoOncb+5JmPjfuLIOFWcXt7/
v9m5+TPkdMW+LNLgbv5GcN1qNxr8RNzUaPCkbxWWHy4ytVaigvOM3SptA9eLU4i2
AP5sdTGTxyEMOcDZFr1qHk4iY/vdbTOfAZBmd+6wk4SqU+ecofXSbhlFaa9QS9vb
ZIna8GZ0vFF0gdVBoimXZskc95XuFA68xeBzC+JLw513Gy8IDF0p4ziH/jadEBap
4UiuoqSH02iZTQUXkTSnertZYJWMt/f3UnWyd2yUPtRhYEu8ibAgcdKr72SLlXWn
UK5puY7ej9s6/mA/eGazR0rjh4JTPwZmBRpK+qJtddD3za/P9r2IkxavLdyy6Hai
FGXgxY+uRY34Wx6jg7ZZ2V0iYaOK2p1d0dLVDzgeDytZ4qejpJXTABAolT7SCBXc
LNWP/N2mxkobg++/NtZpjHpb11DcHaGZfCRWtvZZXfsFVb+rU7SRVAeymFlkreIP
UR+rWOacsTYCXjYngSLyJnVSYSaL1pesm6/pnokZ2HNcMCWwBeCekaq2tpEycoBB
DajekwUwQvLOKU6bNwTeG69BJx0ixh3LgrF7mzgkS5/eSQL43KG+Qwqc5Xpp7IrA
jA11b/q3GeyqOPl2OXn28VQONR7DBcWI7xU4TO1PMGuVlVKurFaZM5JS1oadysbX
GZvuav6eyMimzEicLhBf7IVfqQd/UYazr9RITRpy39x17WBaHrSG0L3YSLlJKTAU
aDBtc1iikkTQyKwPcXL2nXOoQpJn5A1u1uZvzhOWqCjMIwkMfKaBzYhDLhtamhXA
TqBUGN8m3YVSO9geEO9Fk7bwFYlGHl0BeEOEZDpoXNR4DWseMDuJSRo13Wy1o3wK
+G4rnYlWy3A0q7LbxLxJfEUF8mnC0+uZwHsur9eO0e80bAtW9nOcjtmNQqntvbth
+gYJc9L47ZSnhGYw19pmUxhal1I9XoXdJIXNnLKRZqh5D+ObtJN60+4pOhUD4EZH
BA54HocT5eMAV/Dea7tB1DNNYI0ZIIK0RXIjDJ3DFX647+fkhGWh3im8rdyu9hoT
PMyeKcviqlsra2Y/K+8RP/q7ENd11kJieXC0eHOoiVWQaBuCHVliBFaogsfP6GlS
PKUYimA1AMXU4m/8aDEwsWXtUOH1h/dNPnHSO3+zbrsHlgK14WAJ/ChQASQQgJhP
n95R+fWZe2S8/6TvYglR5tBWLao6XC8i1LW4l2Vs2FlYOLYO8IHeDSpid33V1V/3
pMkxqvrladbijDFonr0xaEtFv2N+MbRHWhzMmEDnxGGQV8t1Gm1k1AH1TS7j5Q1h
0OejuClyUI5oMgBElpx8KAM8fGLVNgOttXCVewo5fZVdvbyduYcPznx/IGelaoaC
rSjz/2ISuj5brM7htdJfdfBMdw0w//tsvcn5BO+dtYWCfaiy89PvyskXJOLJviKj
doYOJMs2i6+ZaxH8w7hFfiOpjZSHZdmUj/Uw4UvvgrBfeiMXYyCw+gTBe7jgbPLW
IG87bcD8bu1EEXo324GTXufkjCEiN8E4ti/gIqhxIuOq+aTzKgYUgHd5jo68ruCr
HccnKtIBAWK8j85rFZ7fgmd6eXMy5LM2I8ni3wYcrdwKAlOLJOCaBioOPZNhgOYl
iNRKQ3ANUZw9eGDmcPf241vkzi9u2ji6+1+ctyncSjVhK0mJ5rveLqEfRfWGTdW8
rHtA/59LJDxegz8Hcu+L0glXsSzm3kboJMNzwDnrw0xc1zUSD06QSn+GoE5lGIsj
9dUhyv1MZla1Eskc5kp/x703GsVEuBe1oClNBf0jOtP0TSRCBk7Zk8IxioklvI8c
VUXNzKFacbrEgyGk48f67dNIX1yHMLC6Pagco7VYOKhCnh4rcs+4F42b+19wc3V5
L/hz3KKGVsW3Rc1lLLMZtDEClxbI0qG26aI5oXyfFZMgXRImK77cjfA8Y7QNjwfo
b47UmA4kGJEUdGRzuHaXurATEYe/onnMNgxGFe44zTtVkgh8y7b8G8TYrTFvw7ca
ZivTVvmODu8X6TiDY3lbl1ZWazVd4dupB57je9d5W9Y=
`protect END_PROTECTED
