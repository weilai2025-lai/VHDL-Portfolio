`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Edna7ArxmJeZQtUnzBG8BGPUxo0xTd2waCxweogfjoTdYrcYLKAA/Kmj44KynlGU
Nl1LagEvO/VDS6MQQhhjTF8gO6MZy7E2a/L4LT6NT8MG+CwKoPjvi0aGdDGBZ8Ib
GSWIlcYXaB9HUxVIyXPw6dB+TGzfaqy7L2ctQDMdXf0V39ZB/jVXi5H6Z+wyFmuM
uxRTN/2+QOokrwogtCZdHPXYvr2nbfC+uprt0LybRW6bPbwBBwDFERUDWdP+enPE
ebHFu9u0wNlWyfv1zgihkWGan5rLX76c9kuvApeWdERdRWQd3S5Qc+cds0dPS0yk
M1OcyOVkckFDskZ4hL+lUu60pWtipNO26Ai/b8Sp7wTru2E/68MEZBvf4dfKxDgG
xbmuxJOcl5kMlewA5KIatRIEf7znYlKgEuJlzhF/WQoJwhiQfVGvus+RnBvZpww1
C5OBPTpy/72tb5oeYXLMcs1CcovFZgql0p9BIh69Uj/ePFRc5tY75ADxrOulLgsI
DF6yDhh/Sll7MIH9niMd87jmUJwQPUlTSh1EcGMBUKBSSVGDaLCNrK2lFiXVzhPg
dqEeMOFZwmLQQEPV2KM7E6j1TtKEmA5+027HYNljKVviKiCfQOBsd+jaW0WX9EBu
t64UVJlnblzocx2dq/F9/O3N60xWiULzyZVhayQkHHbmNlY1Sr3wN7h1j3ZtL4Xa
Uh6KQm4uCLtLLnZM8iI6AISgxlO3BQK1KUut7APeybULobHcqouBHZoYbJh18dwY
LlD5ce9kNtTdM3KRn0KYQw==
`protect END_PROTECTED
