`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g94tMrewYyynPNlQGvGY5PVbdDDRDEb8LyjH8E6ssUnPiyAejfA4dBXL0KVYooFg
f5paaYoLGhdR9zbZrBPJtXsGPjxQhLSGWPtsMw9Kr4g3v6AAtblgSUf5Kn1qJM7v
USCHwdOeOqAY8Tj84ViOzAX1rSE7Ui823i90AiADvpDQN3rV9pnZv6zPr+i5afeB
n8a7OVVDapvmRk4b5AYrICZhzGq0qWxw+nAuaBDEl9xcs3TjiutUyfx0FFmwyFoW
QfBH0PrglMK0PT3DCRKyu0XpR4ZxsCcm06x1edD9MVMM9Gj9KSBYhjx1cBpgXJhH
vgV/ZtFa1x0SeWiHOfSQ+lGClOQcmBWRnjdfZ5xVvv2c51xw6fl2kcuXrja+r+HR
KLcrlX1te2mSg/41GkQ+atG6vbISqhV7HBUPkx5pMMFzykeUs2BNwCUWe9P5zdW/
`protect END_PROTECTED
