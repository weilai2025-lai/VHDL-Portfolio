`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oy/OaAN38gXqmL2de965HjgbPShrsT/CMYJXgFlMLW9grDDqa4LTxVnDwYG46Y+Y
DILUWxpZPh+O56KooXtz/YXAvJm6clhPqg4LnNoNQxWqvlC/LKDU65PXUKj4B5sz
xX0btzaiuIAgcaxSX3VlkIgQuLamSTiTJxoKUSyUUNTYTBCpiNa+ZTkuw8JJCpz/
z2WvoPrIIUUsKNqWXLZkMk6vRLEv/JLZJGS4kuKazysPzQvidIjKgDXtgzKhqUPr
9PGUtgqaT0ZB85QsBVXb+rleJPWe7A73wwLHoEN4cDPYcKoSKK1No0zfsyNpDZQY
0IL2ON3A6BZ7Hu2Ov932kx3goJg9uLwp7ytta7zM6un1un9e8N57G+fYiYLrxSgE
AIHixZ3waPMJGpQOv1jrpP5QXG2zn4DnCfOMGN6OsG+JFoTkyMLhWu8gvH7h07qe
g/emtCHPUwOPt/cFe/W3VdkENJBLOcMEiETwqmKpsPhQZishgJDx9rxFDoMzvbPD
TGMPvNl+ciQHHfom04kg+NSQhW8r6lGq+oB84pl4Zxt+0BOKhEWwPAfShss6XpPU
ECbPii/fXgAbOzIx1XOc7CgGT3WqgNfVj7nBg6s+5TmJx5aH/mJJsh6UttgYTLgR
doOXKyjfoV6tq4u6kHrcZ4Yx2q0wkY5RC0u6b0I8YLYEoqS52TLOXDmtHP01zb6s
4c3K6PXWFCGkMiHyiAbVe5KTsWA7+h8epx9MjtjCMic22I3Gn7fI6fsKT7CctHQn
x7mMpmTdRD/QnSBedhupEH79b/uFXmG/x91lOjaFiTyK2FdlBze0++QgW/StUj4A
bHAbt+NU+UhzKQ64S2WhM1EzRrl7MitAuYFl5al+jjCsIVzui6h4YV9jkgqoQT8R
zZZ6Wiatt7l180ne9HdeK1jpsbssAPwcLjhI0QUUimqVaFYjJJ3oF/tZ5s60TCPu
a4bx6YlcHkCtufe69o1K+2zswoelVu3M1DulunJv+uUIDeXmZ7d5gSAzN0hJs4Mt
OCZWRE4zMHXvF2DyOa4jcN+c5mVHZdnjwDdittpEBcny3teKia75qw6U9iXSkLgD
oDTtzmeUC6GYz8K2ok1LN/eCyeh4xP4tqqKCjROvFWGQMA8rRjpj2v7NmZ32VmzO
Q8MwJgRAPmzZUaTitLIcWZE0SNG2c2+0wKKBBdhnBRGILdg7qnf3lYbFOZQypaK3
oh9owUWguzku6oP5XD2tO3NKB2p1Vmwm8xX3jAB1u6tfSvRMPXog659y4pVJpT4m
FhjlSlYfgfc+zo+RKgmaTgrGvh/G2A7n3B+rRDvkoPzIUeS/R1MwRpEMQsjthsAj
qhcLLf7EKHq4LwSPmqzsaklMF3EA4Xv8MScIuQKoQvFyRCICWrvfAReqBwz+z5LU
/sg+iizugNu17VNbH/8e784+dH8I4eSxZYJ2a8bEMZ1cLuljApn31JX6TaIgUHIe
LkrXOKxc25N7VfVLx4m2pnFJKcs99vKLU/a7JZl7lpkP490SvwUdUw37MEl+e1ip
JDfhZvHF3YlPNHoP8copbzhRvbjC0JcTDK0UBMUhuBtqxSdujpe4tkZ0Fx7zOUg7
0g1NdrLF8kdvx+TrgYdoYqdOm2rg3XFBAGWc/TeQxwZ+X1b1kQr+48AOQ70upTKp
hWE0AMHp0PNvJ7n4lEHmBexAmx5nekdeNg5V5qOIJJ5h7xnQogY5P+nH+HEvsqhA
jFhVhGbem98/bbltJ/fL1iidkRMWLvmDUpQjDOdLN5ncFIvnEK15E92Jet8Gw9WT
ZkIXY1rf1gdkenUSB974UIZSHL0U/ukJKWRz2bSgQzVmhMuJ7ask26qpRx0k7MiN
WOL1VbkbZVfeAIjEYuPH54cyQ6m4WWsj6cwXHIYuISylRbGamBkS9G09Dd1uMO4F
5mojfxzILpKIo1uUHWPLkkDwkJZLfK5Y74OQQnkTJ82lhvQrhJ8i1282OmADEvjL
hN2NsvGrMJFehDOBbnPPMaPtLvdgKbovEsEypyZa3mmSBwe523wR+Lw+sS5hkzlU
O4Jxn04nk1LR1s1L8qOvH9A2dwV7WF+OgHNkoW0aTLg8NmPbmO10JjPGEB2W4Smn
6F7auBZnHmjLNZp1ueR3rolO57pvqU94J2qH/oOyAy47534VRTsm1Y9hQfnhpOaG
slPqeGG4JPz7pf13CDnE425+rAxRmI05mXc9exq1hbrGDHD/GGENZaiclM3xMTuI
5oJ9ndXANg1lS++wLxqipdSs+epEPIJ2li5fYv2c9RTInAVEyOszjLtDrW9f5e4p
80ZXWhw1j+oNy7XGlIIDByvX2SXpMgMcDadGFKe6iRaUfuXJRsdF+O7qyjrvv7Sq
EPl8E9prZtC4bfDgU0loiqItUppIJuV/LvDkRDxi75wAxy5o7SsuleBCIFxcIhGM
STfS3G0kTFhw7PyEzheBpJguR3ZLi2RdNX3OuKIj5StNKX32ACwRnlK+3Ewe/NXI
e2Fd0yEI5/yGSz5njJJnnw==
`protect END_PROTECTED
