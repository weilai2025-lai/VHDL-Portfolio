`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QFpGyci8iyqFrSxwZ0fRkzXcQJSpifqYvO41eiXb7QdkrXdytdD8Ai6cPxJS+gf
NPOLqZGYkdXp5OD8UYTcmYJl3DvNuizBJ7H3a65RWhh7LeXHzhJahEg47DPYBN4T
D2kP0IPHE9dkiqsi/gNTEoDJoYMTMCpBLeTiO4sVcawr/HTCLF2o3OJb88/ZvjNr
eNuCozpp8iYGOLlHnPKzv/+eSLHi2plscByKZuHskstC8yWc5vV/WnI8ExOnvnQs
m62XEHRshnSzWHx9QicegVHo4UR/QNUK4WrNxG2eoy9O+ExC76miVqaFQyeoSdkV
sTZl8yQIXJre7WbnVeBL4QcZttV5xj7OOmw2TIWM15ItTA1LLq8kjzEAlUJHfSAu
zH1KAu/ALwzgQaRgifwP9bg2JJfrLu67mBAPKSRfHUX3PXyEU4X0SySUS02j4gnG
VkUMMhdINk6WhbmC65oXWA5S8w6SjyUehHR7r7bPgU0qq2X1Hx53EeHUI7VAtdrv
TPWjHFrM2hDCV77rTEZeOlamJylVtMiVsskxhKDClpA08PB87p8STD8gnAjQ3gOB
AsDJJpBYlGXx9cNIMu/XKSAWJxg7dPOhGM5/dv9QctdDa5QTV80pgj6tsvGMjbaC
jN4ZjqRlvcoJyvjch9m7mCZI+wSEv9OdGaANVpiZrT4mzeBOUCbPb/07K9acYzeK
afIaRQ+it0zLLUWkuFsJaU5DQ06H+orZaE9Ea1Oj4LHKdEhQTBhLrEK//CwD0jis
7Ef4HITRoWK91HviVc+QiYhCy/rVrFi75MG/ZnRIYKZ9bDbYDYxGE6hoJfrWt712
chUiWFJYiiWIlvm5xK7Hjw==
`protect END_PROTECTED
