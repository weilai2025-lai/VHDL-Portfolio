`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6O0nCXyEHwwKiGC9rycCUrD/Rz/o4nxKlVcT8JcVx9uZCuIF2XDWYJucF3bW5EA
7NA1wc/9p+PVPNyn3Z1AOm/vrWHUdpW8OzTwOxfu/aH+cZYuhwFgYcuFRT2VFHE7
LVtv/K4CrDLPksPtvZGbeAd2VFYCpVm2Xzy8Yh8oc0a1qro7UqSWDvs9RmDNVJNV
LKXLeqVBYQrUL7Y7H3oxI8lyjWAEEwrQNQVBKmXzXiAINgC4mng1Ogiy3RYMIhWu
KwaMgLO9gtjLkMNOtOcwoBMs6lJSpP+8vSgOIObeEpZmLq5mNSQ2oK2VCEAj9ldT
wjDAcehBOguMBSqjp7DYIvBe5vZ9Y+7zCJXzXxRbpI+gYOM/3x9D+uJUMzXIssOI
4STT8xwx2fvMXfC4D0+02N8GbOYbXhSUOmjQeMK7BM0MHrGXvOe+F36ryl5tx38v
tiWy8xO/hVTYokB0uetcPWOykUpTZqBIayfEx3MaGoP5kAN3+L8IkpFL3pCqVzrM
YTxMm1dyXQXHFk5DDfYjw/OSgPI/sEzOB1hm5ljMQbiOIwA7mY6Sln6M8m7A7tDp
ZaQ7u0jU1j7IFJbdR0BsbOaTmVAckSLBZIO502mJuXwFmAd5HnwzDB1xmSC/5Apy
SDGQfPynGoxHj3xqzOtvwVpwy13su0Q86QRx/WWuUtrXsE9IJsUXlKkuPY8HBMfN
Qm3asStz97VnWWsTD70YiNCtvX9l/P4k0H1A6YrGeUbNQjZ6I4gV4EUUy0SQU5Mw
niL4XAd9yiQWQMMBpdOgSKEscdGUE38SKAOoFfSb08pBYomYETBQORHMInjSwfDV
m8/0HCgtBfnc9baOHscty5BrtB2DyxZxmD5xdKD9tVODrHXV7Itsr11nSHj9wjtx
wPksaJsdw5h2YCQjiZ6hDBtmq2Bv/tOg71RZhJ+XrZELZYv7uERe0mFTitjJCr/K
wv/YDDVUGcdKcYrb8f0MVPvzQyWJojJft5uLTHPFErgrqfLUHtKr2WvvhGCy2uIm
V65y96nvHcL2iIXov60f3/qnQgSr70XtscJJcZ8CRZ761Fnda8ExraIU/I9FfKfb
9GL9iruX48+tR+gcTWPqMItL5Ai8xWTg9LaqLCX0OXU=
`protect END_PROTECTED
