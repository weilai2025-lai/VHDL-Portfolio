`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkI/YDkYBXg0I3qesveUUo51eb+2xp1OfWC/YRtmNJz2p+vd9aXml7br4g3G1t3K
j1w9ZmfKzMqrj1ctg1hGibhI9zyrMYS7N5FmTkWz/WJIWH87yyRa18j1S3iIgeH2
4Fvmpt5zjlf6/qJsHAQdDg2zxQTNfucoJAP5vtVCBYc/c+RQmZO6BYyojXgwBx/j
LBocXSayIj6C9qlpfr/G6aus2T74WGLr6OGSpW9khJJz1uT3gOHaU/8t2nbvbXBM
We8ddDDjXVhCmLydSBU6YkrSVN6H1z8OgbfGBYwvAPDXb9HQymNWcLNQPMSWv4Iw
qQE0xN0v+rH24CwlDmRxbCxx3zACI87Szp1wC/eJ0Y5F0Og91Ljrm2CmrtiUFWrE
J5aVJquVOBH7arPi0b5M+p6eLCSo3qRpUwcx/dV6eVGsfcUxSoxDZQgNvww3MipG
qJhpPCM2nJbSJ1A2S8gRuV7gxhCQMXLxwbDcP6r4UbkO8lj4jUB9IyaYHAYpA3Q+
9liVciTgCsBhaqZaX0ynaJmDuYEaWYKOp5pgEVlbsbv1eZz53gADayM/fluGNCEn
ZsPyEqSjdoeTr1jSzZ8px9oMXC5D8aT1+9Wb6AQfeUhBg6ZtxBy/NvZvVqyzd/cT
3HzT+vNHkTPRMZ1JUi1k7gMBdunYht/PbGjL19GnywDTBwewMOA/41/75rYdWF7Y
29WE8Ic2wPZqwqXf+Qty5DdkMsskZkPSJFaRrjUt3ADDcmS4RLzIsfIceVOnuQbg
jPYvmOzJrS6sFc9XIxrpdVJYdyUAA/rmsC6Yd6ZEc3H6u7XvKR1E6JgRXjiAlHiH
4nQ6aQ+DkW5yXksMj7c6Ftq9FEmc8jTLnc7yX0eD6dPsNfzEeZwcG6b56/H1E/HG
CSpeBR6HmbkxPkuQ2nRZhHA7U/kVwoexmSAMruwdEIpfJmGjKSXPybsYAhwYvjEU
fby0BnPWCtRQ8VpW0NZN1AcDAXFSZ+/NJfI9nnYSGGf0i31Iol6c/PSuc3L4Wi56
P0j/064npcOHLcMIqxhVbvXkHhOR1V68quZiwW4HZBBvUeeRwpRgZ2hFnL+vcJA1
8zVGhYx0x194lcIKa8REaffbrZvl2V4RN2prlLNG6YaQz68rjjOms/xqid1+uz5Y
oVWogpVvMschp4HCuPWW7eWZqhc7H/5Q5D0BTzM3Jfr1Y4sDDUGNvgdwOuSEALFa
PFVfGamYLHa3fmVV6LkPe/ueYlFky+lVahwd+5M9bQFEXN3+dUH1VaCBOd2AA+S+
rIf4DfQ6dZlEw3wzmppviE6eGUFc771eHbXp7IBkUY3ThdpoCHqXsqsmWhR+wMJK
DAvEoiYipTfRzqcFudb16KbmXGaP57dRaNZrAY8vO1bpTtcvkyHGtLS6IqgiCSdz
TldoQdkSzYerLkos4Jal57RyeT+o7X5x2x9WmGCJMKPFkShIfHY0x9oRJhB8rJok
cRmBt8Wfw3hcF8Fsaoc8xfMTbTPmX6HpM9FfjDhhDzGlNzLEGoG/wbn9ZodgpWRd
RuCPS/F9e0/BZnqUA2HU3KGrU6LfSQgFz/M0T89yyiIpgZB8R61GQuFEbSLFLmsc
ghqnLv111zs/5FWJfXO/40SRf7ZnhH91QvE5zFmSCg/X/fPQlRm+oQ2H1sQBU6jx
Oh4AJE2I2hlsn5IdKKrdB3sYV1E2ySvPZ7cjZV2vnj15AijlrgR4hoAesR+XYkfw
IfOcy/OP3WJhLtdREaRvzf8eYSgPDYKOVu5CiF8ZTL1LvYb6i9LXjJuFRmDsDQHw
aJ9ZHsQYNw81JUlzCjt5lQKMJKIVL9dXqr2msj8/DWkNNWUvcLmJZNlulULanZ+H
/Gn9IDdONo9sbi3RodXBAgsAvgHcmyjC0dKCR1HN1wPz0XH8MuI7Ssn54ZpiTLv1
aiOFyyTCpUvK6j0ANJEAz/TqkLwoGPJEqgQr209XG8pvlFA2sGnEuOSSixHawto5
P+HdUVOHB1GlfZcwS23erRSZIk5bmrqMctNpavblOA2MiyZKOpd+RzAZB/qXwH/+
3ThEsL1K9QWpxOtccuL546E7SdYI2/LhrJpvX2x+4ajZXCvsPywgBUANPCuwcHMl
bRPvgd1etNOoBcaoGKlbRculJ01DWhyyZThAm5keLPv1OJztZ2eh1PsUgjsVomLO
xHFihPfRT7faTiLHj7qooP4zyLti1PC597hbM5qxBekhutNr/cQrSVyz5jV9muWH
D1A+ltvJPD430oza6zuUH//8nSiXwJ1pHcUnyTnPMiox24bnznxZThzrso/UITyz
VIO7BfMcfTm2vp34OT+453ptYlwwnhsiYMDbqJs3CsGTu9qJ6qYNrnis9bjEf0Zz
Pd1B7RXVasNda+40Jq+G+i5hZ6er4B1YZ71+DyPkLd4=
`protect END_PROTECTED
