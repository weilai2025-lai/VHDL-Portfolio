`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1maYXpKInpcNHjpzGX9W9uIL1vsJIxVrhpqmNo/7ZV9xjDUDE3RSoF78DwZHucay
S9VzEtHKwIIYVTq6gyp0us78RsHia7/+hKY5KLFpyXydfC0ddWLxwgRzXVTjsNbR
ca6AxobbPYAph4A2Kvi2P4pU7TzP/FqkmBAPIoF+evZpvtBErfTREmkF0vFA3yEK
YI5J39WLLGv54l/8KSQ6AJ303oVBsYvsQ3Zos8TH/F4ODNgS6Jr6xe9sUhtGqT2f
ZyJZ01BoYWwwo7UZnMD9Ufs3aA6AlkVyCXAB/t8y1IaQpuFkeTt0p+7ZWkf5Cmac
0HV9lSnQE474N0DCnuExIRdpExMSEMV3LTURM9/T8Phq9N+7b8GiG47DUvKrSFHQ
Fb26u+PETAXz4UadaHDP3zyQeTYsh0lqzrg8NEafNq+Nvgj6P+SZyb3AH5TIo0zY
iWD6pY1Im/VHMPpV62Lo3u4/ASWLM8XxsD/HV+xAFQmWrZvw2DhQHbjcr0pTeR1b
AXz/ogDHST696t5Jm5mysZLq5AUZkX1cQQMP3QOQ8R9n+jM3+gz2P6/2ZcgZLkha
CzhI1y1wgifj5rvd5y1DdDgQ2Hd7/tUDjYhJ9n9JwnkDXSF20iktiDadnBZE74Fq
Pgbyt9Bc5C1zdKrHACBm4rnGbB7REjJg1f9CMQZ2nYgsQIYhIAItFV5fhdIPGswv
eX4j1P09AV//asn9OMAee7V9NVvND5MFFwMK6CjnNOdApQXTa7L3aI5NGB23HIZw
ktf8ZvbB55v5eBA5NYy69jH3+N4lw9aiymozYsv3JxmI/31VJlARNHvV8HpLzjwM
0IXSCB9hmQFXR0AQkJRZuXu9qAXTY47Zo3xUaSq8MLlJaZCW/rLh14sS54l0PkWl
2GDQ23uLzo67CO8PCfRplZ55eNIYe75WACw+pdJc1UDfYVivCaxN+5SDlkVcGotS
7WuUNfrd1Ur/0DhYX9kj91MmAi7TGtqq2kAbUetrmjxDou+e5sQ46LmD41hHDfy9
OTqFhCWMy3ovZ6AhP+zB7yVnYm+dBglzqAJRW/t/XDNmsjQAeTJeQAnICk9/w+Ea
VdOb8vefQiKPY4Fcl4HETKbDwDtL6729EkUHQz2EKI73gstZmTAZZSIkT5HdVdvq
9pZPRSN52TIahsj+YQiMsdSyZYfLWCzGpDbtcGRAUa+r+uzrKvdVAnCpqJNXkDIh
UWa1/Q3Ix6ATy12uTuKm3sphHWG0vR7x499yimZOZUCUzp6vzDFMHQE+8lH2kyOM
Xh5VNQ58N1yR4n9bMKYx//MYvFVw3bwtwE+74W3gNysot8taL8/secVKO8jljcSk
Nx5NJqE8XKIENJgE6I1e5kdV2vgNi7WgGY69IHIhlq4/d8jnUGl8h1VIi+tTDcpT
14xp7hVS+z18mRwSTq0O2njH3R6J/EWkxvSdPcJi2512XXNfiISqGPC2zkwDjv2l
gkyN+yQ9hdogOM7iShjVUOITo1mZbf0iAF1hPgZ983eYdlQHHm9J7RPlDgFTRtPg
dUU5cnUqm+vDjZTBzeZssw==
`protect END_PROTECTED
