`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Yz7JwFGrksHQRLJVm0iKR+n9nzkJAIi3aiYLsXVhMlslCzRNKol8FFRwramibn6
aCSjl5dVifs248IR6qN4zfMclF839Q5wSO71DUBlUvO61kpwGOH9icZJ61rG3j8E
DfDzCpzYUSs00PyvE2Kba/8uZmY/Om+qNz49Cc73d7Ha6AbiGJX239Yxbk/GL4d0
bYD6ZCiRX/HsziNtpDShoVInSnIovYqXESg1PG4TSILPZo1/ZWKa4pVRi7OT1ZDZ
MEpks4OvtDa6z43ZhgpVWU5VBI2fPP5kvyHmJ/gF3biVkiNHJWXXZ/lQda910onz
0BwRCAl/zTqzBveauRM7zScEi1kw2avZf4qGA3y1DuW5Ai+uQC4B3dOBC2+cSJBi
qvaw3uTsVK/S366zlSDcMIcdVb2Z9+karc527j+45wguu8ExLP85NdvgCKu0wk1B
kRXO4k3q2nz1NyGNr9PCpGQQX/d/wIxMw5fAzW/vK8jOz/jscbZwI2U+S661yT1R
eSzJW27qB3p5PLmyiG20zjsmuIp8B8AdXlCZVgltEjRfjSJI5cmOZ9VRji9b6XXX
YXbTalZN/dXYAsvM3GbOB96zR9XlT1btk7S98d+QsBPQbs1rrFOxP8UWh1aVcguY
yVCli5CKEP6KTvVAw2lSFchWmUZ5VJQX+tXL7bp7qmBsQ7H7WEGYA7cj45OQPij1
JS+FA/aXmQlxGgh4Hujb9voRRaW89AD1isVweKKh7Dynt2d67FGFa6nz3+/atPuw
/ykXR22g29DFxA2hv4J2PK8f0LZcGuee5mOOHwe8+kCO6GR/rcRm78Rwp+yKF2Oj
lT9psFx9CUpz5ru40hzTQ/1XNEX1e2UQbVR7yGIy+InuGrjXzLqInZtHgx0gAC2c
+57Gw/kdzBVzzVPwaN9/n5r1SUbfumungTYkmPhA7AEkQgOjaZaA9ljM6YSlrZxr
Omlv84u8QdFi4oOCkfW9YA+pXYmr10w9s34jZmWCTvQq1rGY9vsOImRehke6hi82
HeLcnzInDqQEzmXYWNzvEogKdOgQFZJZF0O3C0ym+xzRowmT1Ni3CODevmEvy3MT
IYOO73wdMH6qybukT9rlDYj2dCuoM0p7DVN2JQlfZcVz1+tH0ahpQw+v9odkaifE
6szAz9OGsn9PyANqWDkoPyL3ZYUepDeIOdLW1aoQfQBd/U2yiGdgpY/p2C6+EuiL
pVGy1bQ3uakaTEVilRMYM1d/P+eHjWbHYTgiIhhtMd27hnYLoGXdOkwJxj/KKbDB
dRELUJaAWBhm4Kz7uUEnRkZF8CsUIx5rwclFln33upsQJROJuUe5irEi9ncTdTpC
4m4NjMgwM8wK/j5+l6gT9HTooFEZljW4jnq6GmYMoO8cAjbikpP9P2Bh7fdEK3i7
f8Mjeq+e/lHE2b/T8Wk19lzi2w7pmnwziVydnzRy59DYT+yhBpOXx/3zGkI29ML3
`protect END_PROTECTED
