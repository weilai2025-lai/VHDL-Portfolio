`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EdOi0BVLBNsw1XbyIsT5mGJU2f/3rYnI6MjYyeJgTdV60g5DuDhnfedk6x19/p0k
bn+dKK+tHoL0lbCa9V98uonibhR1MYyMJTbKZlKc+11hGOvvbEIlwKUDzMlSsxVu
4fBlAOTWXu2bJ8HqYDs6ObIJiC1OVihvqTJMzT9Kiaq8Fbt2+kZ5RT0J9sqxqqDe
sQeuvMdy5G7K+Hr4uayTsyr4cPAT2t2+dFdZKJTGXUuzjaS4IDD/0xEKUuBpX/Au
9RdcSxlRL8aEXsM2vBBnU30UFL/qYZ4Ul8Tpv1s4yFAegXqLL+Lctekg+sJ+mrDD
4Gng1KIOor6V+kUS1G/ZZtsNDYibo2JxOeY8IY7I0iiUVK+ckf3seGaTaG2TcxLB
Y8+1I3IO3mLGOWXa0Aq/QHQBw9Mkcreh67FaLHqxYXz/JGZo/QZT7U0MjTDg4ISY
4fBOwOlNUbu/3c/co58LV88K7VQlNsRogzI3s10bO1IMAhti0A6js6uPSuSo4y1a
uT932ZdR9+yvUACMyCTU6Gg3+hcclV4R1j5e6JkLEVxfyDI3HNwnF9T3JBKZolyL
pEchkJhIF94nOv3NX/ZxzzlZPVHKV8pWPJaPWFonpcY3tTs8g66QK88YWXXbGv/C
Hhegk98WNkM7sHsBG1H7KtjyBRJumqhaKWvsBbYI/J7ghb8iRdJgeBiIHD3uzwsk
92mTHVlZlUG/BO1hVKMGh7qXplaxao/CppmZyOM2cQoiu3jRE1ggrBdLOVme2afG
kfjC56AbKBSz5zEx8E+w6p3FgDs+diZgkyghqVzYp6IcV7Lw4KFE1MEP18OT8eAt
tfYgq68DUEF9bBSp3lyw8Io1/8fpSy0KusFUQQQIQfWBwsltDaFpdzp9NEVaS83N
SEWGsQKB2yQMr38//7Mi7AfCB2A4yiOYt7kBs9svS9dFQ//yMvjzBysZLkUPnz1Y
`protect END_PROTECTED
