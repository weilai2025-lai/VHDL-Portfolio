`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RB6rRSgG6X0GTtI80KuhSIbwzmVQBmtWBbM1PDx2OotvvkKlutOA4kaxo8g8sEd2
5B6Du5QCtIT7JMWpNGoMRqw4Mv3ZGMsWViJGqhPvgCfX0CCT6SRTek8sHw9a85Jw
6TZGeDjI9HLwHO2Mu1eBr8fP7WYi0UxYds2H3k0uNyhKR2BRGMFc8x5kqEBJi8zw
a4uae6vEn82CIiXnYxemsS32bm+jQRi1GE21r4rplBezUJXUlRFe6ZS/OTyHR0lI
0Qgr1P0yCz4hzsz5l/F7b8hmp/8BVsWCWGskBclrO4aB9godMT9KOGqBO0d2MZq+
ZqlbnuK40I+6xDuR5Nwx9IeryX8amLmD0pGxwLTgqdvUsLQVUk1tLcKkIq7xcgkd
RVG2Z0r7r6l2W2xHw9tQiVZ4GCFNOgm5GQj4menj9cNj46buegL25+XTzG6EO2qQ
XdJn2Bipm/35QLp45BpESzK3rHUClgHlaASm7pP1sNzkw1JAhYnKau1w+vdqJHpT
L8uC51tXsvpjRwcBNg4TL1fsun55HW0V0yrhdYs50l0zYBjRdfNislSndhaY9tQ5
a/DG2Q7bDJ2pK/sdZv04xzbuW+pCf9UXJNAsxTfTmaXDqZDBBQTOW4Bg/xkgdAK/
hk0sPhYJsYsHNlCYclLeC71IeN3tQ9k/x+bOcNMPyH5iVrfu1AkhKrzIY2Fpg18I
G/waRIFRSYXanHM7UKcy7og2iNaHtyj1SsNB4fbs6cYpa4fV8/GuXwhVSdPEvfNt
zDgTJKEqlgR07wUQEG1H1i6fBsOpgxRqzRHqws+czArwOcO8MXawo/Mj95yVQ5Ry
70gSvRJIwUFPrYfHqDqJ8sS/F+CQ0fwuyNYMUms6Cg9L+yTkalSvu0wSHEOZzcyo
Zhx4eeXk5VDK7RcgddsUipsTVive8kUPFzTynIvTOUGT/nn+qr4fzAEX9rLX6YBj
oXuGGgWbcsBbF2oxF/DB+DnArGVkotza5wM0/ko5sNm3KuSJpF2nmH9dyeRDdoJB
7U99TSeWVZrxBGhHr012Wu5ZQr3m7QgQRhRBXxoAjV+EIr301f27mPU0Cmkldw0u
rM95w4MoRyweSasEpKdM/cVsghcPs+y2wAiD6JFZwdNK7DGlOcD23DCAGa5lfIwb
ReGbuUanQN43KjRf0uqFAgjV6k7Z38agXbIgyDLlG/SPHigcDSNoLitGvtDB/GXP
/xlpvXuqiJIvJV5yKOT6j9TsoQ9Bo5057CTVWDdLB+RL7Ay4dxxdosH0n0Ykfx7Y
BOwkeg9mF6MxYjDLW0ir4xTvB+VemMs0VlN9+7F+rW1nl+lRQn5v0LYTfk5wT7i7
NldFjse3h/Pz2KFlw+wfAlAWkkMMT35zhKPMOO6/wjHHPMN8Wcw3nBCWuYnumviQ
9OvMCddQdUZknGIgpAwpR2oq0vvLbzYP+yzLuYRPLu9N80KVP/XyMKyUYWPg4DyM
zaRqNdR98mzlWnxBp1RpsbGglTpdySnOpvqdr910ioq1G/eSlvny0dXi9sZixid/
IlW817Gdn5y9cD1NvyeHpZqCLZSZEa+46k3t4RMQkYwopG+dHMAkB3aUTXJs9oUw
+zAt7SjofI5LM1d8UEOXFdak+TQGZzDo+aeVR8kJ+L16EJ+9CA63AIJ4f7+1Ce+h
1GZxmIyrBirB0TTmH0hWuuJnsluZ15YproMVz5126FAm6gnkpK816fWqFXQsARd0
GGwG3h2lKhwdtuY7pa+njWZjmDhdJPymymSSH9/dMGIDRqpRLYn8lJbwfJwpydtS
afk2hSY8ghkjZOo7EPiT/itTCC9/+kztlg8X7ftUPV+69fD7X0LbeD4DB/14HSD2
nn3K6uoYNlAFXD4AGqjc0C2AkXF2Hx/Y/K7is1NLyTIz1hvRQdtMy0E6Otz+3k7N
5whwWdgEum/WdUQDBcywsc3RQEQRpYJqNBj0Ypj20TRKtn/lAB4XGtpItJPWX/IV
P5kDiQ/EsB26tMbo0uMCAu6k/SdOe/ztpkJgHU36hbJp1JkI5gxRcneVUB0/T3yF
RfDt1lWGQVxMKjiOOtft9F8lJUKmgc/yOTJ9yh+Hhmh8Ob80ea+OCnJDDLKmoKaR
SUvh53xgzlaNiXtKe9Nxw4u6RhCLJvl9iSMbPYAyekq6IEVA4XCDderniLrmZroZ
p8KfTDtO2o69yEZLhLQ913tOfDxnbOViTfCfzNDtSf+DVsHH8Koj9QQFw+0mrho0
sG2Xby3HnJ9PjKR5l/U/OYNB4eGhurgwypthrNsQpg3tdhmWiB+xqpQZmzhdRXlD
vHoP4L8zMkYbnG1iqhXMcIADCNFhlXpyE2sABvwHVBzoikBE1TALiQHqmqFhmTHX
oUhJtaATLPri65EKFmZNQmallMn83eJDpYOyqned93n+7k+++ELTEeHlfC2EUsuU
Ni4xhMoS4yBK91IO+b19sY1vgLykio4d3upT0WeYunJWOVQ3jaCeX2/rCX9J6g6x
I3lX+wU5LX3lpyvUDhsOxRqHBdRPtxyVc+7wXY0NkXeMpOr2U70mgBQV5zjVVjWQ
QGpfsF12cAet2jugz8rp4JxvAv34ypuNa8SiiQb1VAb7M473LAFgPrPRiUf1xdMo
Il4ihwlozp4yipss//vGDRDN6bsgMq0+bPW0rvOnS1vcNv8aRoGp04lRk80Jx2wA
h023+d6rUQy/Db/hoocjOXG4BlSawSbDuwRw0WlxKn5wUf9lndMILcutb5mfJfLz
dQGda4gi0AbwByE0HIMzPODz3NMBkFRYKfOPw/YiFQ1muUWa1Qg5x5BUI0almOFD
1u3EPtXNS3bZjRYVnvz9+AKXRMWQuiXd9Elmfcg3aZNWaknQC7tvfzOxhn/nSeDo
q7gc71QsIB8TWaxEPRn8/HywXh6WbD9BQW7NRJPVdB/rgmYoMzBGs7KEEDbuZvxh
vVxRnXfVFV0FwXkmB6x2Zi4hDpftHTsdaOJEegBmHzDQ5eVJ7yAA7e3NWTkIGO6j
o5FnL6cxheK/NqeIelqHOa8hCVlphMm69DV029PDu6YpeEG3t8fSXQD/799RiSwh
hDEOFdFbB///r0VX5whCuYiCvg4cu4uapDvVoMAeT1J8mRC5Jk+MIGAq1ttC44iH
p8xwGnn0M76fAAY0X5Yjn96wknHWOt1FGL1wuHhMYwreR3EJoTpCQSkFIXlelbJ3
OJ8N0AOpVKku820G5jRCCSWvocxuA5vgyKGejeJ5a24K0uND59fhl/ExVJc2TMsL
/z+HU+pEWn/sc1Wlaqllk0EUIwCbGLxJ3yPgjYkBsFQuukhJjNjqWVv0Ah+HbwQd
XqDS05DptWygRHrqSuhVTn90YhNpI3RyphCd0qXXQ3qjUrxQiQn1g8ArnbKfmpEK
l9QI87SlZPFXPYmk9KR+klDfiHengnv/tCMLv/DrKBGAcJ079FxNw25qr3dhtd2g
jD25S6DPnh+j3fL3V9pgl6GQyEi38fqjZeLQsAcTXaWG8M9EJzv4cJ2pdzgvMECs
d1BJCWm9MBKPM6+FOCAaJeDTGc22YgGJzS+lDYZjGAPM8+zjkiQne9XxsI5/RHth
7Ie9qaaZxRRa7udcp9UvXupUpBy/4NK6JeRSGThu/zhz6/rKnO4yTgNb7pq/oYW4
CgqCHCHtk/urzLay5Kkx4MvugpCIi92SJ+QI4KAOPwt0MIY50OEU2/bEo06BTKDE
11Iz6gh1HRwzDnB6CMcFl0V863fI+lTEtmbo0pJBGM0CzNhHJ5PlnIloO3zqfV1D
WjbX4fHihSEicr7NRBInekp+vllg6RtGT2yw2PoNUpshVkc39i9ItlqNKhjuoGDC
WYlJggYcgM9XPGSGZwbzIdlkrWiL5K6sLibjMtF2UtzCmWd7KizSYcgfv0waEE9H
CnjEAF9Cfix89k/jJj0xdYMOLzLVlR7WLNbdm78yQja+aPhP06N4JqZLdfORsPvY
BxZbrG7KjNSr/MN4jTw8KYWo5XPwilqL39xKTVt7YlTGDmpBIah6uslfTt8Z3lEe
iGGUqIrrQWzabxEjWey75wkc3uW3YOSHllvFjkH+PPtFlMqT/bgHLV3U3ZT+fB1t
SzEONB8pwyHId58uU5HO7BeMgtEUQem9WaGkRtsE43tLBTZoH/Ic7JOWYP0lXjag
jxZB0WBqHgg5EAlwgn1ZPwKv79lcnavcQApI1Ho6XgSEcSfln2h4pAHXZZrs/BAB
REryD6L4cdA8IwiYTymEJGh2R5+HMO+Qvoeo2uipWNjT5DsobfuH8fwHQJe/65yD
OTayRb13U57fr5a4fh3hbTUi6KPGa+1UGVwpNADOzzcA1Juupxj7A7ozVWQ7SKMd
vU2jKCmKYJGOLR7pCKv0xuZJTm1tfyReG2IAlz5BKyA47e4mrW1nGfhoiDmQ1P8F
4504jXJDpFmPkrPj09F+Drd7jUittU3sQz643Y1gXKEHlcLqn7oa554N15zC0YY/
jMLA0AATiUc+C4+nbiBqnBhluFGundq5ATeVYWDw9WP8Qb1Po9kgVNQXqTWdfhx2
Su6oFxNPsEO8EQ+m9iVF/WefaAY+2shP+u6lgu6/Su0djBSBW9r0ahADYm2RUEhG
e5qv0xarx3WPGnrJS8CNwtWhxTEReNWLaHvMvZhDNyBtaeHw2UgSg3N68iryiVzX
DjdIjGOvihQAnr5LscDPVLRSVyreCe+HicseVlOghe8wFWNFEJl/XZwecCBM+st+
PyceNFQ0+APTdfw09XJfN0t3hU9s5CJmlemYaCRfC6tjdY+vC7olo7owUcJzY2YP
TB7tnGvFyKwC23Z1Y/+ehstaLhN13KvYElTYqp5a+BzOrgeAXi4UVeX4ald0KScj
p7JCCtYZWP7UUS930bc0zXJmaOyFHsoSwx8TBNAnIq9DcmB00CX4hYKlJ4D8Elvn
hayPYqQqq4aX9r+8AkdqOLaFeqkU87U9G9gcfoLUxU4M+OncVWyv3anIKrS/+sjz
ciFhHQ4Tp7EdFVF9TmF+B8eXDRP3x+kGNJmDVoEXn3MEEawGHmGnNYBRXB3xxsyW
Hu4FAHHUnWKfC7PU5JI8Vg==
`protect END_PROTECTED
