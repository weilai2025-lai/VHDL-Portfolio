`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTgEnQBtqW4WAYMK9XDT6JBkYZdQUUc1RNzmuetPnhsefi1JpiRxpNLCDGFJayZc
DGMCObIue6U1hupVFVfgF5DGt0YpWSWdLR32z5rrYjYKx6kIq/t0Nj6mgZGyb7QI
r4BrdQKK2V/aKlwpZcYqbtFOwnmRjg5alO40EdxuoTy5znaurlnpebIYqky32znG
6Kf8tXAo67MOL5Qli23bLzg+H9i28jLdsHMRyfr1JMzboGpougomCZFotELiHhi6
bcyPLhoO691Lgs6ltIuXWwvYHpZQFWuf294e3mD+u9XVBNwPN9iwUNHq4MNov/Qb
fHdwkR26IQ1HvVSAQ9XGjo/4qaCcpIEPGccHjWX7mNdl9xf75vywfKC2knC+EhFP
jCO/THBO5+Mudryfit3xDA==
`protect END_PROTECTED
