`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zT6m26PhjcKIa5BEA3UQOFCLjWA6H6LsN8XBQT6Gnd5kme9vLC8Cnk2xVT0yDHc+
FGen3dm3c224r7SJ4GWu6fxAQoADz1s2jrGbknNYyVBAJKpVk/3iXJFB2Kw/DgvE
Ay6wKPIiWmQ6/YNX8C9ny3lG6fmGZKydXqUNtf6uDdKZe/maU78/MpBVjcwI0RkY
d4o5BzHaICcH1Da96PXWzQ3JqBeE0S7YuvtZI/Eq83ZSiopJA6I4exRvW4D6aF09
gnty5XePDP5UCXOyLaQ8BZCv4RM+USunaZUTIJ7IRlurWTzIh7wV/P3Zf5Otaixp
HPZlAF+FYD9BeHltxGKZCSdPtMUKsY9qW3Ea/fgXO2LFphT7teSXJnSDAnsUqO/k
S4TSZBXkci9zunsWXR9F38esCskUSAyQusNuILhmLO8Twah5vb9+eawq4x/be+Qf
LjMFsAVzaRniijNqIjwCVv4DjtoTPoQFApUefLiD9MHp4OJIH8bSHaM4a7oZYam8
259s/TQ1eVJ/3FvRQgJjaxPjM1Ixc2UHcf9pII+bEIYF7anZ604UzOyyOQ91gXRP
EY71KwZ9fcU2vq7pTZFcJLcYlRawikFgq5XLduGmvJiSCQ2Fb530iz6e1P3WIItN
rdt9yiXDl4NQHNoIF3a2LRj46GzCH4T3VeRKi3pB469jSviKlWWFmbBSYHJBYa10
8efUxy/IKEUAkKhweqLxye0kZ+Qz9fufaoMTfYfORarFVi9lw2FYsYOvp174secR
HlmcK+rkHJs5yBSVSDgrGcsdbYJaHwwBbNTV8AlPtEsdU6ItHKGky6osq7WC5qUI
r/EEjqJRgGvIll7j/8eejdJqNRJsVQ2UiBZRIRTU2c+kBDU3co3lJdT4Jz28s5AW
w8gLxU/lqVniTB4bOpXQ44esnV3GAkKQ00V0/D+YQTdOctJ774ifcW3jlxrS0Cxo
`protect END_PROTECTED
