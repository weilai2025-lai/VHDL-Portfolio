`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhdXHSn8zSWVN8II/Vyws0gPgsfU8AQgnMbv5hqi3KesVgOrczESC8koz0DwiFGG
Q2cD5MDXeUuannPBX10WGbe5l0rNYDotz/4QZEUUqD5wIjY1Lo/icNtngx8PjVSL
1TcyrTdtTS1RHWDtv/AWBLWVo+pqgd2uS+YIX4/44hiT+spR8cf8NDO2XVIJ5w7J
5soAE0ehfZ9drZcSq4FCYgM5nn3S/3odGV8o6+McGkZmccJr/UvayWQw+XRYnCBG
nYHGGC0vcnWKlOeYCxe7l5Q5qMd4buKDIOViaYA1L8yq7AWESlluMTEcows0Pg5l
l+HCumBUwDOVaD2YYxRvR7BfoRAG5M3LmNw/fpMTk5IifiX6CKfaamXH/MU/9BKo
037z3MF3O1j+0+CEg6e6uQpdyCCG4kXLfCkD1LsZYhaEvNDQakWHR0dq4+c40EeQ
+cNBJ675lgJBvcAcKyxQkNMIqGFzoV4Zxaoa+7Lk3owlQPrkdrv/COHlKzll3rq/
lulduST8WEmucow73gcDgiLi3W0XvTd7rz9LtwAkVvr45qxtQbWgrMpIG0cKvDGB
Zh5a7XJjcU4rJElAsEPls8UTyevlpqU1ea2nj+0PAjTMHDgy7pRTDRj2Jt84YvgP
Fn3kHKb0OugDADdTYCHSq4Jl1RKqbKgBZ30Lqfg4w4Q=
`protect END_PROTECTED
