`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvd32Z/9xVjDxAKoEmlxmb5lqYQIRKtcj6sBg9gV+Fg8hyrcQlFOdzoEpMAkjVQV
Ef/EOxowuJLElgImlKHvQUNwutw/ngVIzzPnakL2EqqJGodIXeLNjBpKg6sLbfdw
fy1kBEbGjABJkLhMMg3y4TpwTtwT7n1LwnGAg15zwyspaIi0P53FTsYMnX9oc9Rv
MxjbCFR15xO4cVWMFfnk8/AwvO7j/We0Q90nN2typi7j+pKOCdYb3kcLLvW0CSms
KvwQUJ/wcemW/tlbWkjGBmM5wwksvdXk7m2VhuNlDrpXNbOADhBwAz+oRdk6YeU0
ddA8zg7KLrMe8tt8SPu2vYt1xW5vcW/BUTZYq3aN57dO0tOYACCatxacUPW2db3x
Yrm8jgj9vj0R2mGDgDEXdcJHUWz2ANwqHkzK66E/as16/f1Qov/28VVvJQ44F++H
GxWZqVlqGTBsFRr0WnW5KmUG+YHEHdzOylIu6+AyWHjmh6awWfJltNjsgWUu7NCS
i9SUDiLkZqbhZkATwaTvZzv8VStWVsCxFgK/Y+/88e0=
`protect END_PROTECTED
