`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spkcbcQag1iOeDRlI3usdyu3qRCYIM4v7bDbhTkgMnVEQWzZ+SvjEkuK7kAOPCgP
BgrSgbmNo1DamzuUzfngHroYps8xOpjOQWA+MKpyV/4Oa5oBVfol4+83cBp1FU7L
m85JEe7iPSdgl9ZoU88rtdne53qqWI7OuPRapCm6g10O++3pWEnjH1UaI5sgm8Ge
gH2Isyg5/m9Cqt0mMEOewzeGk10DMIW+cLZd/Lpk7jsRHZb7HrsUjmBj6PRqY3aL
ye8IFigh9wxfjv96x+rWJzL2XsmnPwqs8Ug10/dIg+Fr6+apGyiIbM1+L2w8o3J0
nFGtSSRRC43RCQo3mOXIyn1QoGANC37bvFYGTIfeW4+Uq4rldIdDY0++xAb1cFzv
SXpnZGNMPo1GhkZlPu6laKmb+kJd6qi11ZFFet5y6hu9kICz+AY8g/bJ+QgjNtuw
AqyemPvkER+Ld6ICJELVf6bysS2NgLOY4ce7ul/99dWhiYDZYUcncEL83Go/cUo+
1IybBxHKcmjguDXXC2qUtqEobYz1GjSdCvSD116/saucIdfgkiYbItEFKQowGEkH
Yc/XgL6faX8HowHFrR5t/kDGAyEsGH+ALdOWckcY7+92Zic59YiiaL5c8B/zjHBz
wunQ+NiCcIX+sGwHuzg+zZXXGqJ6RL31Lnwl/7w5ZUGpmZFWNhgNgHxKKsWUrxWa
XbOqvOd4AWRVrSEIT7Y5VPHMlvq028C83UNce9ODG7S6l2BAbjqj8ifDs35FpB2B
qQsX9q+1QLzdNKZ2CFOmRvr1IbZ9z4AE0o5LefIUBo+t9YzCd6PM8PnrxddQaGbA
nT6TmayxiI6anNOein4fI3mFEIGsW9MVFUtXKQBLf9ulb42UKe2+Y0DbriJJ1jNF
uuE2aUoqaoC4kiYQ5I+Lg9bFdo9vmi6wR4BlIpLD/uqX6ZYcb5XMzaxKoMlZB4zc
8EMVndKV6zDPMnIDbNKnE4keMS5VqIUjFo2gTEVDGgDiG0TiRplXYp8Q6NvRTcH7
F8JIy/shqMlfA9NmgF4lVmF+Su6xWY9vscyn8bkuflxqKwjcpcaXuRKrbHRe5TFW
I6U0QdXBhYHKmlU+DRbNxd9vwETN6IvoMv+RVSH2QRq2L6mQzzeVbB24TInOEbIb
4xzXaL6rvlE3tJyKXJk/9j5MM1FgGhZw4JN/0Kfw8kmsYj86TcPKZHyQrobIq3tM
6VMmgKYklsT2Y9QpqIv6SXIu+d34QfDAQkqQ7aTjy9omT2leLyTNaEwz4QjgscQU
V37tbEubBOvijgk7nnJfuARbAUqt3hgqIApa8WDj1v2D6zILt3hc4biIy0XFu2jG
gEbN28t4UFrmADQeGgJJaQXfmpyacPM86Nu8kfqdH/dgayiqeHvNZNpdIfvpHNRQ
dl7JGTZJe+0Psp1NsctnkGUI4AP9vE/hs3ruXzN4OsqlDazP1CGwN9dRgN+kO4X8
BSgpwri4kVwhWJFCTS1SOHKeJ8wvYhQwkSB/3Lg43u2K/dwD11zAyXEDcaNUDO0X
AXFDpBj/skOC/0bQMPu1HNp4xNv0QmE4t1CRRA1TQ4oAVJ/kxY4NyT8qfWUK0spJ
J1jZng0Sccpi4mvWVsZ/HePMZx1iZQMgg3aTNAqOrF6Upn5FfA/eu5iXMsnWMpxD
pcROAb9TUsZAZAMN4SFNQsGr+FVvzyd1VseWr9EgDS3009FHrWdSpE5aDxg9GO3s
FABfVo4xAGn/50z0Fl7kvennIGCduDigBXJhbUPK35mpIsUP4DIxCmow7Koct2PC
A1XWlptGYiUrofLJySqnxwpDFd6U1rBdop3A03Rtd1BHPtyBl8vJZtj73nZ16B4U
1ikJ1hDku5Tb3pKPNh91d/PrnDMZ6Yrizvlr+W1I1JX8v1P65n60rbZq/CDA28mS
z1wyKLazfoUhxJcVkpD5GIjcX8cDvv+rF747Gy3pqlg1M4GrKl3sNOuAmCX08B9g
eWXznHB4gav0A+kIoCfU36AT0ZJH4EZ5+lWU+gO56hUljUocLcNeIudck96GsbWV
Bb1vL45D6S3/TjStITaslHlv5T+b2/UZohO8kMQbuhsyNciykHJpTQnEHkwZjMW8
xZpqRLZ+RLoKc0667Nc8ZI1Hjw8CryQ8hwziO7qYulzWPmJTQRjWSyWTcmpse6Tj
gPkbSf039pIzXGKUWBLthvrUAEJveVl7BNbmFIdGso+YqZ/j6XPN1MorEiwuvz8i
DEr8R0hvn0+zqRLGUf+CTVy2UXkFI0QBcGQa476thJ3TMjQQydw07z5aAixBZ9RU
e0oSkXkJhC7FMM4jgpuaKJ63uNbLAmXttrRtwC+GNr/irrr2NZpz2s8HZNHIscxp
14FWU8iJYnhofxT851NwTdsQrRppt8mmjHKdHSiczrnB870+w6jahyU/bGckbI/w
ypHcVSYj7FBvThrEwZJvUSDj487T9FGAcJ/MAb4nRueznNfXVHp7Rp8WFau7v5vl
iS9p12AwLDvWMXj3sJRFre1WtdsPWpVS0rG9hNgMFymagt0EE3uTo6JRwcCOj6do
VMpJbx6AfDN7sHPp+RAZuS8EO9YuSSnW0xmNCJxRP2VEFvZDjLd+7uZ93YaK4ylx
HAbVkOgiVIe+9/phwBVVfO/Lgw0+UNqf09uNL5XD4+6eZz30al/pjv1i1tuKTfis
GlAHHtdsclFmoZyMEq7LIohbJ5TLdDi8eFUscUD7N1zhrCL+D6wyd6O7ff5/BLRu
3QWC/9IrZScwCkqs3XG9sKCbBq3WBdR62VxGidelm/yLA7HMDIg+445gJK3aeDQH
g+nIn3r0kPOmR44QEuMXJWuJWXL4OTbr4VPQRLNLfEAho0g6KKvHHqIEFnhzuzjj
uhR1t9ikB0FA1dn5PdAwfOju5QHHsXfhstOKo5sTtQbVt00s/HyHMCxrWsmzDr+4
/c/TpHahvOUi3qBIk/aOCIGwn1XGA6mDOaL6Qs46HGR+s1tXG6baBcohaije92En
giUoJvlu9TJq/GZzAAfeCuCbKBjU79nBYiJOGCPkULJ9yFDZ6CDSAXjEsUYp/yPC
U9KuyOSzk7rlckXEWDmyMWsyVYEdws39LbiqgHOGsy+aU0s5qKBEeS0NPL5qWwbZ
iRScQQ6kuehOdqiLfjHl4RF+00IcFO77wSINURdG5GOa3P8zu3VgMHwes7eVwg+n
5cNwfpHv3FNlNoxJAxA/vzfQOLLxNJyMdCOWbxclWSGLjkLGB/IDuY5BS1GECTEU
ThOt+iaMIeWiESUivPEM5ntXDsFxJz28JuGtshGFnISgbKRxBfNu/gqXcY+sRPqJ
4hBs3vuVu4pWe/nvu1m0i+3xKG992kigcSy+qf0AA5VeZBsvgvmC8ZY7oXlpDPl+
y997xwOVddeDpJw5eOjtINiBMJGp80kQU7MMFAmg1HBU9c/66//yeP9t+gJvTARS
D58whmAYtNLbk/8Rb9ifqmrhMWm7A+1iJwJdznKsMvyu9nTI/g9J+MP5yHY+xvuJ
fEKWN39idmwhbfo6h9LY2KrLb8DEOmLx4mubLlFPO1Hr1AvWSx23cK3G7Y5GTtC1
w0yF31v5mgqxg0qmlxshUEXnNFdyAOOo8b+S+4bjLy6pubbcRhPya5zMd58D+fln
c2uwJdmQ3m0gwYcwrjwswZht3vskGOFFeDYV4+1MgCtFOptDVuzE9fgsEEJTSbF/
+svxt77ssQNZXfyVSjTlsoaunKfzeuCVThZCdLEkOHeFUMQ/98Mgd0PB3O+jpZGT
KRrvu6Q83aLj/fcphc9aJCye1Izogv9gPmj7Mxy9okwGLcRBkgc3m1HMhiX9Nkre
2npjCCPtsyeCQvd0QFqX8Jh6j47YN0luiRAmX+qmcVh+zSmNB01yJ6kVKeBZhxqk
jqVTCqHdGQYe8Z5QydKoR7T2rPjvYY3+AMY7953ZrNz55FOItaLV+zrl+AOB+NKf
XblYAAqtPK/KYgb872QiPHdQPyAImHRzVB89sbfmqm6WBlPlcD7iJquXTZw1TEVf
dJRYFrPCU0LeFKxD1zgaUsYqb9ZfDEzXQbSlPcR7VmPkvJsvVcnKV65F5ei180v+
XW0kCPVaUFVs+vvUvDJJ3xQnv+DDJi3rMWX+P+ftQBXE8lzuNPmH63wBcYUVGCrm
`protect END_PROTECTED
