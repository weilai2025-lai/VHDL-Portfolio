`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiMTv1NHeSwfTG6HCGFOUYJLZw9N+I4cr5vfpLQIht9BU5iKoJ9R6F7wboHTXCeJ
KkXv+qzGFrwAvfzcJXQCxXDT1CX5YI4jxSWags7fp/YPANcojHdX8CylvSrEMV7+
msC4yscgOjKB+LxBCkPi0APXvtuaoqZtDJkk5LfWEYdemnBb56WiQptmcmFYVkiT
1RO9mE635Dn/EDeArssHpcumuiAk+yl4xAhqHYM2LwHG4o7YtvrrhITdDHVm8w07
Tlt7sHkwMeTcQisSvYaSQ8jivdstTRfWEt9HiFDseO/60ZG0RyfZHR++La7mfGQ2
0BoaJAnnIt9KwfObTarl+EstFCtybe+xm8HLp8iAJcIFgKNRQKZo7b/hg2Dc+sTC
WoPdQJ3iZq4K9EzgLkILc6woxc+5XLJuksaSPvGlZ3VEmFhDjDt8GK5XZGhRgfKv
Zv27n1/tVFFYO/TJxh99Te0EVYr1bb4Uh0fKkAMAvPvlYRAfxfgsX/ieoUHwZhqD
Pns8tQF7myOgtURxmpgzFJjxnfKIhwRk394VQJ1EhHdLZCHXWCi1gMJVs7ShTZ0B
jtOSWkth6MqGPa6AnpKsjVw5nOZpitgQ+ImY4XtiAV3jpElWnfoRu+pQ4dO9LA12
0N21gmCYt60hmpV9eFMfYs5hsgIP3wuAz0K4JRWIQ7rNL1TBAMl53auRrsTLSIJR
003cQpICPddPIEH9TjhDZKGjb18TNi8NZ+yb6rNJZG0Chh50MYEMD5AKnvsn8UFU
AxpcJlty6ikX+4PHtMLPm3DCCU/E3eWLXCn5JF+4Sq5/tQ8jv3PlW0Zrv0wc7Li7
dlSAz4nxfZXaQuA7IwTps+sm+dsWhY3gmndxGOhfeUvuNykNEd5H+7d33x44TyII
+qI4SZQGlSY3vm/JwjHskG+vG3DUZgfQ22sXtP2whiWkAVFsSvuQwA/4EdxqhP46
YtiUJOax4oKpuXws3n+CL84Hb36cKK8nUYPnzcxfit9QfiFvjomtxf81JdwRCP+h
TuPH6e11hCeXVkdU8sHshHsogpfUE4vL1XcaYNGdR1QiifxXk9+GUKHICo5H1+Q2
1H4aluqGW6wxFAz02rsR3MKHpVb0KkmWB+fabrt9cb5g2X1kdXLrpPIRN0pNLxvE
UjO2rQLaZ2ckcHwVVZ/ANHBXO7JmaHuQq6EnQCnvN43iwHZJ/oZqb/0f79GjgyBV
owonKsUV39RSDb+4HSiRJ4PqL5n2+9PJdNVjX3K9gcxSwDtec2BRCzHGI6nww8/e
fzXZph+srIXKB6TVsokU+prs/0qaDCB3UOB18EOWcoov4wyGoozl7zgq8RWVf8Xu
Y08MvVO9iTbzjcvId9xSJ5ZbdrNfICMh6VZEJlk6jmSE0WMXJh/DtHQMuObdEwsF
K6ylh7I5pi5RgNR47tE3sETgihb9bnCkKeiJ98gRMdRFj7SXasJi4HnmXgHr/Ra2
KDXzmBFgp1SZfmKK1c6v4FfveyKmaI7zdfPhgvNNCiAG5Pet+iw+uCRZ9K0+iOxu
/2HdX9MgdMWWqEBe5dN9oof3iSNGPtv2eZXz1SrelnpxHftgngdR6KY8xVB9v55/
s3Msv3xtF0FkuoJvFwo6V8bPkvb6nqCYVA9mb4vDdswJK6iNyMqt1o1GELjEGVZ8
14YPrOsHrRSd+R0JdcqGH9XjlW6DSBr/htpKfOVNVg2sP7o2VAq1NCfKueYjDRvw
k6hvevE0pzPZvbIDgqkaZ1uVe2L4fT7ljI0EUN3Aie92GDlRINGloZRIqIYGMtK4
tck2CbK9YvoKGsecAeBuBaA54SjixHNnfii7fjMc8sNFjAJtTc3+j1agAVwzxNZx
Xoom+oPWlKC0aAtAlU2ta1arLkMcl7yXwZWFXPZKIfFBvmZrf4ZIzoU2wYuPwpx4
niwcumcZwJ/E28iaZsZ0E8poStFXo9fgHMAnV/SJBgkc+29UzRb0DxFFugygdlOh
vPmIQ/TkvHJOtg28443yjMS+r1fGVaFz/5NAXee4u5xVpJ6JrYLwmQDxqC6gYYYs
fnXN5RxpCXni9Tt0Fzh8kAzVswJ3mP1JemSG8MmUAaSmxElnnz1JECXRUrCRp9lf
9YPG5Z1EQH3rB7cw8bpLP7e6bHpZ9rQMFaHvVkd2VpgrTdVrqmq0rJHOyjp1QdMv
VpYNEJ/WIt+gno6tw2dbPbtEUC6Dxwoi/4Ux0q503ViT3CIjtpAZ4znsIystpRJx
Jm2jobziiHRwCwc2WOV8FOJgUPM84dohzsz+hjGe6SYrrkAZDMnKRaFI1fxcbvCw
jAWhwksa/0J2ljylS4ZY/iWeYnyQDLoHBZA1Cvqwy0Sas1SmeFVSq9OcMnFDDe9t
1ovn+n5aeYLU5ntrnS55y6U1pVugTVVd+wAup1ayZVW1SiiyifI8+0e49UUk4yRl
WHDa74uMyNnGtkGTcPUJgIo0C3butAP02WvyI5GFHsGZMgK5nX6KJf6fxfTz9BV9
/meuuEURiMhymXjtK3zzV+8on6jVoS98ZDBUep2T/KjAgkGGtQk9/4ZdvDMSr5Ho
fQSd2IKzMvQ8KXZ4r3K0Xc68gZmLHU5G+asl5w0KD76DoQsr+oWZV1dY5ScfuiX9
xcmYWPCKC+zuzYDkksVULLmTBIQ5MgsUkitYWCfh9l0NfNgXkviFWXipG+lGkrc4
RFv1gkb5b7vvWSM4vEqaxmTngJx6zYpy9WMgDuT8IouTMzwWaenQnYyV5sfXhEK0
gNEn3uflzsR9PRNCCsxhrsCEcv494WmGWEeN23GuFMCZN+ZoHefKgswhgWIrIJA0
EfJV4kp7Uv9utnfisNyE0oYFXl9ljRd/DAo5c13J7+D/HL6/KZCI6tJkxexL6slK
3UTBZ/RWNJlocoRWsY/MVHGQq5PACkKiU4WIHf2MIiG9yFfbHSWHHfqRtIsK3iCy
ABml0chKfEUCGJr6p+TMMuEtCUh+7nKPk+4w/J9JlCBujgIlRF49YkSRb6iUqLyW
p70GnWJ1F2xGNjnIyqzEwYAFt/e+cTvDkwvAdDJ1mQ5jbG/EOK7MatsYwrKEU12I
bQsLbvFNk5fy4bXKeuCYn0/2EuhT9jJgaShTBtlJLcOC9MJs0qHrP8ZdM99Cgmfb
ELLEVCkkBFBJfV2VJhsV8Fjgg14i3Z4ukFGtmdjD6Aa/BFO2JXQUSTV4988QbVrm
v09wsBbxXwVK3WEExOP0fZUL5Y7C3k0oAl49LrbBSv+V31PvvMO0+TE1stnLSexP
sMl6WTN7jisp0pIexG/AfHm9o0vUgIwx1N75v5GufVQEQHJeBGVi7av+bROJtWFR
w8sB5bDOstN+OpSyPiHmosRwuEoGOBPI0nf0GTu/2ZAxDUuao7oz2lWdRpshJ1Qt
tNxiNUSGYrY8ejhnBbJ9Fw3167UxpzZOoUKZrUWGHiDXdPKoaOAqOG9+/pEdIXnr
x8IgewKzp3GJunTsh2N19P0zY8RsxUYBhTpozYhZYo8O2G9v+jR6oRfs1cNUlFgn
KS1kONlyMmOlyMzBUpGH3DNP+XLd5wFZlG+H5ajz83Iu7mDSoXg6FujhRPvB5Er+
qFXGa+X20K2GSPFQE2P/3yi3CizuQrOxagn0zsyfxf7GMoGyfoznSevZ/cIfEZqj
q++cewxUWxY1ZeOEOvkEhKTkRAWZbt9MV/7JtgCvyDnNTyWe2EJfKUN3oemazc1n
xwy4WyKtkcJYUd1bYBbWSM5M66L+0vl5rAzt5DvoYyicLOnxmisMfNd0+WaqbMn5
GE+PRvuM4rroIQ3+XPvuCm5Z2T9T5SkM23aeHsUtHQXp88WISHGPrfOoupMefO9q
5GwIvoc7uKpv31up3vGaP9WFb/CvSWpxOF/9UVUXJ3U=
`protect END_PROTECTED
