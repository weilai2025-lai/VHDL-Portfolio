`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K1JiImyt40QSaV7vqAj7p6PnuWwpWXHzGXho1LtIwJw81d1oyrz3EAa0+PoSDEU1
a1KczQJllBEsPDpefMF0iysTOgGb2IE4IKDbxSF6SA2JYlhpL26CgDnD/lidfVRv
SB8zrCXoAQO7fNfsPa2t1MhYYLx8Z9qV3A0sTjC466seC1UeCZvPorO2oQm5lr8S
sGTuPIknHRCTOr2CK0PuZLj8zukAg0IKpEbftH3V7tSQjShCfVBLJVZbFlGlQqv0
FlWDrWAHCDROLOf29Pp2FelYyxUdBeESuMfrLGkGsVpLofpCeWh68F44gJe7ojoy
USWoHKVb+BxZJMXOsHatE2LPlHoEID40jl/zcPU1MyHUusO8zBLooK1GxxRi79ED
XNfpwGErhlN4Nh51I5rgN8zRKiDRSYLyOYsOXZWPCQsErHWXxX6dTTHgds9rqflD
VoQu/qmFzQKG7A74r5HYcAxGOmmrP1tvOFAgjQH2hKQKD2REVcfGINGdHS3uCUe0
tJYn2D9h50Mre7QX7Q3OzKcx7Kcw8FoNiwHOgl5QlZOBes3o2Y2/MnyzbNe18IH/
vbCkIos+YpnEw+c7Clg6+8ei0SiHlmnyU6+RLkoz8gvEcqw+tZaJK8MKrGo7vvl8
rCrstA1VPXjrYoQqSOMPUr8pymrQJ5YlD7wMAbowK2RuKqDEnk6VIEZxDRgq6H+t
l5hpDHD/IouR3boKm9/fVfQefhycEP1/FYSOtrGwuUIWNHWKE6Fjh+dlVOQvY9FX
NR7LUxT4dsMqYkSOVRyHz5vrC+hHwiEEBcZnwnj6tH1FgbFol87Et5Gey4KDnc2f
yws3p7PUsUbd1LTO3NcTuwLhfoUkOY/6eFGppRpSTHo6ys6ejih3ckWNgC0d84XZ
EzoGamM8JkMeWrTpO3xwwSpq837w+o0tDgtu7hkvz+/fYM8HlToAI++n8dIfGVfK
gMzG3snG1y3oWxmXyybJvw4r1pNojWYZygs1ldbA2waaD942e1AblAzuqP5gY7V+
mXVKR/kk5soOAng57K27XPKnbEUJwVQ0M2saGWSc98/tmUSTBvcAMBHEbV6BJjq9
BqEQKhLlG6wJqSOthkxV60GdduNlN/UwQfXW+SzqdxvAFTLstpbCy2ULjvxE6pJg
yFQ90O3miuub0bd//6mYcFpgFkRPybMm5qmzqCByQnZotYIQx+85lKUKEzs8vbRd
1ZpyJo/e1NAM4FgSUX/k3OyAkbkAr7UExtO2EBs6HRbV156N8T0uCMlepy+28DKa
U/WQiyFewLewY5/DAMa5/8yEtosikabAt7J3NLT36MkJigihvBUeFTjE/J3fSRPn
GDBvsQZSPMzAGMVD3q4U3CE6JAS7sdiRNYFMEs+GhjwMwrCwzApofOADn77LpJT5
egxQlW0SsIKHUCsRwZtiWWnY9Ff9YcPPG/6Vb9cLZejHFNTz/+oE5iwIvWTjCNDR
3Ff/NsqrIbHMnwLTdAOTw/GG5xLsQJZrYm5MzZP9dggLKw3QU17d9vCdGDeCAT9F
yQUu1ieJRIWRPeFzoMDQZGwOeLcNHaGWO1m+VE3kWTcp/Egomj23IsddgPechyQ+
`protect END_PROTECTED
