`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ehff5inWOJb+eOkWjvh1fjbZGksFpUYPSu4p7eSp+Q6j/Syir1clDy6KHeDFzWC0
jFGCcOD1jJ3czgNPNzjY/wSRFEyvPuCrQwpVuV6EM+sNF1xpIAkorsjidRikBUM1
XoqG3fEkfTAy02umTySoqX1ofh8Y8jx7iCiivhdEyW2TuY6Yp8gbAtVuZl2oDhE2
lYZsC/AKrZy8V7SPef2t/aeKL8kqEXs/jWi0hDsrwXu6Ke/7SvInXCGa8NwDX0oV
L770JlQO3v1GC9/jThcR1sYMjqb3RqL/tO31vFxOlhnqUrN1HTJoyzdR4ih1dfHk
pNJ663SHP3TbXhcC5ZH0HkMF+WhWQbKfwUV1Cwmnpwhwz4XAhViCuRI2Cuw+X6uI
Xpv2omg9xmzjYtz1sgO/vnwtkuOyhzqET3s7prsq2jmyYaQFGyv2C27NnQ8dgqNi
WmmkcI+UZrml0WZUmSqG5a/VBO0N2HIJNOBubFxA1genc3GZmkQwi1lhA1zDqEEo
vxym2eLNqzLLHkk6Sv+szt2Ynvc+K4MVZLr3Cxoaft+pyrRVsQLwPelcCZlI8T5w
HaGmlkef910m4d1BGjb5uxf49Ou6qEJmxwKyqdUYvGMruFtQV+LyZSZ1kQIUwgb0
wucud7IO1tK9POutL5YPKOtRh/1SoBsVhKyjdK8BUbJAg+WQwtXQHH/C9hIgyMLM
ku+hBAhe9lGSdlzzKc55IFKe8wQa+xE/fTTaglHQZEJbpE+a5slb+6gzL/h9eL6/
SumNLPEIsQXqRcnuCmFkj+DhSzGcDMKaN+npxWNu/EqDXtK/wtoWYnbTqFPb4req
64BZ2Jx0VKYvFzPXECjxD5RMtGrP6B32U6E1q1aVLveaMh/VaJdrwF43ztif0JzO
e+98ZNxPRYpZTM1Saq3Dcee+l/U0v7D/Qop5RscnZ+rRmn/CFzvTvidyiC7e+wE6
BtbxVaFydmrbCI67Crwzb0VILQtgkStDLe52s7S8KLA=
`protect END_PROTECTED
