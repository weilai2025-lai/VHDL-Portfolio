`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwN/axNC965zCJ/lmAI3dglzII1a3pug5UeguBiRwX3v1QVppm9G5VuVsNcdqJ3H
zIzlwkXQUa8li1LamLR9DwJt7afoMSe59VkdsZl7PUm2vO45Fh+jKPZfA6+9b5/y
5DH5isfjsXU3GNaxNuYSD9lymABIVURynfkJrfZ9C/kUIU0ZFVlrn5KjQO/kA+Fl
KVn25CPxCayFijYCYb7W9LCXxQmpWhU8WZ5TYYPXta+uHXlDo23B30OOOAiEAzzx
zwvDYb+3jTbSzqw7eMsclsQjlSl1F+iFCOiaBA4cabq1LiY7fQWlzHWxaqU6ERqa
QpHrzl86ry39LZ+BBc47fs628lyTrAqJgJCC+pu9V9ieq/9BIRGDyu5axzuc/1dI
1UxrL5czMg1am9gLOVoi1zjHqUrPOVQPEYsRh00ZB+oNu7zSnWWuvyi1dB85zmo6
vaPqyiuFmN3xeqdS/13oLV46oOlZ3Nfiidwjqjac3MdcaIe0qTIxh9xCmSHF1KPQ
abelYASKHSY4qOqgRS3OuiGjOqM1iuUwbA3phNd9kxqEG6k0cqPy8uKsw/LHYtb4
z4msWdlEhMTAwvab/6w3Oj+OuqltkLFY9Cu18958vVcvVD8Jyc9K0YNqniZUpcng
1DcY4OsZZVqURK9fHjAiR1gYG5a9wzq5xWaRJu2tVKQWgTmp+ggikodv7IvyQGke
c2en/AfJWqW88rNUsa59K8wbGnpYEEqiKZEHalWx1nIU3BcVLB4iwG+5ha6LBnoq
CGNfKxawLgUXr861S0aNLzkePc3vRcPFe46+2u+iQhjQdDRYmzhLKW1pefOPG/oD
pn5ATYf9f0RNcwoAQM1gI8CG5jaDMht2hZHbedicXsSfof78sXWGrXoY15o+4Bux
L1qdT9r0s97Gni/v0RGE0a4EMJL9DlPKm+qqqKfGyT7tu58lPR4j8/Ze0wDZdJkJ
+3C9pH7TGuuUBHZL24n4k2tZX0UOMkpEd4CGGDHWQIBmCTPzYx7jZxdV88mVw2pj
EGR12a9A1HXlDYqAdB+50iwxOKactCOqX1ppXkSoUlADwFZ3aDq3lQ7uhyBQyhCS
9b4nrAQbpkn0GWbxKBeom7OZXD9botEBXSbf+T4vDoaLeoc5HUOkwA8f8LBcU6ih
xhI/JFDi85piWNSMAQYj+zFV8nBomI7HA3TzSEIVG26W3X3/EOSXEuJPcokpwXaN
M4ulAvAYTsGzeFGe7BHloVr0jvHZ2jgRXg7hdKLdfgAB0HbGrq3o86hEYEm4Hcw8
Rc/k25U2YGBUAz5DEjYI9AxuFOxU/eqqwrnLM8bn5p9H+84BpfEGyWJRiIXnonXl
NUtVIT1vVQxjSp7sIbStL5soOzHrJ7bM4oHFA4Mdvr/KLi1k4lp2bkhM8fPx37p2
+wJJarcfpSNTxnOTfIcZejG5i04qdX+fc+qPv9Cm4MmxeWaxiYDkFHTsEYWLrEyV
Mi/JvZJKteJwJbJhQtpT7etkr7KHal/UxTOV6g6cMeAMvuw/K553hId1ud15CBgl
gF4lQSSVWgSU+OH4p9QheVZaFSMu/J8i+MqYT6u5uBYfmTRcD0Qth8F923+t2HA5
v4Pb1S860ngrkHbyUjHitp9loxSud3guX8jGa2NMqCK2VB635A9V+iEEf1MoMEtH
FFR63guDFdtzJyNnNS78P+ylfXO0W6VlQR8/7dpWUQZNAnWrCbN/+Cg68z0LC0h0
axkwIToJ7HDho+q2xdrCXEhHmwxKyazBgVgfAqJLz4CKwh77vuoFblk7dRtb6mQI
vgGDfSy1keT6E+LHJNaxd4/XtLV7ElioXeLs/9ixGtxvkbn1daHAvsjlQHswibuc
u/q2gmuJr0XYmGjIXZsNC8l5vayK9NzJuqUykxxgWDQO0fcTt7PAaOJebDf6/IGI
`protect END_PROTECTED
