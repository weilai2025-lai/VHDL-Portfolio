`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BBu0391eQrNkiQZKoQbI8saXTrvGwoKAGaEzb/kJWDlWMGxbMMtjbkug1GbzznnW
waHX7wV7MiR+9Bgsd7iRh95uxdAhM0wiXek4HwwPo4smY4REb65RKoBV5bWrAXkT
GIeX9ur2RvgY8F71iVGTAqGQVWlUTNH0917eLu34QnJUGEsVpzWe4HT2LK5ntTmM
zCv8wijFHy45QD9xEFCmqXvAubL0eAnclHbyC8evoDTpW685ld/YicDYJjgcRw6I
SYhFqrOr3zGEUYsw0JudZjr25QA9JLieddbzVYQm8CW5Gq3TZs2EGgUby9QsUSxr
sghRqFYvdVoNQLyxyloMJ133UZPgpmYL7muLMH8ktaOvXqo+ONgLd4HXYsaV5/Uy
PRFPn4IQUD3N//XB2kNfwJCzK7SBGBXPKOYupn7de8hKjhxrYNLTOwkiEf7MyLYV
LTwhr4AapTn7dhZIFlXhtKVCgU8/mU7mGC7ozSlBcq88Vha9B8U2qWTuF20+JyjP
lj8gEiq+ZI+aRt6UihYkC3fgOyfFXayl+Bjwn82F8dhFOXEqaTZW2v0dUgFriJIV
u+zI6z0BqHWvsPO1cHza8+GJOndZhvCkZFRSn5qjO6vWxG6ko97XeFjVzxe5Ns+y
UJybweJgn6VU1hpQXmuG5HpqjD3k4lRSJbRfsLCcev0rLpEa/S3W+g7fbDqXQacF
FNN/oVSzcSjLZJZL8CnSER1QR2ZFp7HPBbjwXVP+jA4Lqldlv3mv4DnL+hRyHTt/
GcNiV7yO31UYMOABC1e9Cg==
`protect END_PROTECTED
