`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1CLd21RJ+w2/cTv1bx3PSXljS9k8sEudK4hyhxGw5WCTf5HatjMo1gNd9GpzxWj7
eIAjZAGVDuOMUsbFiKkeI//XvwslHILJc1dGYnjr9mEq+j2WCBCn+nGqtSvmZEcu
0kHxDXpcm0j2pTN9+SILfouk6DcHsu3Nt627A0oPb5kQ1xAi7Tc5pddlIAMIBMkx
AOx7YBjxyTIk2NUkr1/hQ/tQd5lSBLtLAojoPHCmHLJh07YRMDABTevOw5SOtgRA
cYwfAY03JKiSaKcCQURF/VfF8O5nWUd/NJmrMXv62w58SiXuCj/TKkhcl6stnrYf
q6ulPB81Fl2JGcIlUwcn8dP56Rml85DsEcC7Ot30fT0BfW5/cDAWYmBpgGs8qBXd
9q4sisoV4+cCKthG16+91nZR9x9C6fZK9QWG7Nnn9lJUneDCVUKXURnUBgxi+f7R
lF99Q1to9LQEZg7H5PAQjneui2y+tvqCfh3gGZojQJ+2juJeOS6lExeN+FWJ//lZ
YOvZr7YaPF1HgWHns9xEJgpAxZAJN3QXg1dk4Nz8bD7+NsHYWksyqqCejHsnpwsf
2FUaDwbwzyZr+xdCHx1FWcS6XLcXvzi/7FTCq7Z2dacjO2KBEBiAfVhjlW8cCjHT
EL+3DwRvy8iBhQLEBRbrSrvghAQzOYWDmDGHrz+r/pAN2oamxa14m32Gx8cSZ3dD
gwqAwGqx8lhJ/NPtYy/gn33ScKhhSf+GUU3fuZq/lKs75MjkXyF6EB95vxQn3eBS
3XEuywY8AnwUtxSbuVgMOErVwdBFxzozEiV12qkOYJQCiqVwWq0bIAsg3GqSjzqQ
OeOaDO8BnyxJw4BfiRK5Hw==
`protect END_PROTECTED
