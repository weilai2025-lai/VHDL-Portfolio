`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grKRva2vedxrl+8XFXeErZBVwEoprBCYO3OPmZSOiMngcmN4MAk3jsT3Fq/y8zru
MV4Pvu6/04CwuoLTR8cLpyVVxzIm9TxlylwxlkV2ZjbZah+9by3yMCFePaFpSbsD
na3dxU/CXKk9oI1oGRqv7727i3Z9OAuW2R3+T5XTatPW/md2JYcYN/nbmvLMuwKM
VxixAdqzAg8MzHZbAj4ZLiUKMu3GM394kA8Ph060kMWVE5uTlgNKHMwKn4hWjmo5
MwcxSe8bwiPi2ZEMJ9hf2KSLHLMNAuVrb8hlKIAPbhrLr+Mr5+PKr9pO39JOFKis
jdOBhTR5VcC38JZS4fn509GVIJNsoV797wiPbEe2sn4ua4tBTSyMVSuh6TIaCpA1
7EhDl1L0SWXL+PqSx5DJetji7EPrQpofBGbaIeViFL8tgtu8HcG6I48SDJso4HeV
wjqLfRoh09dF6Za8jXXgqUH1Lc/FiZll1A8ztvuD+081ww8E1+MYttvvPncCdAA+
TTTCvayiibaJT9idMH0r3Kn/kq3iNnawdFYUiVRB3NElLdQ2DQhAcjTK1OrGrsFC
Tv00LIgRGu0ML/3TQ7OfNr0L7NAuZ6x+INYSxKA+HWs+TZkL4djRVuStdtapVpL0
ad2UpRN8T49vYunQgig72A==
`protect END_PROTECTED
