`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gc/tquUHY8N5xuttBC53acK3WJHhj/d9obW0uKE95c/+WA90aHPXg97Iuaa8GB5E
F2dVN9dut2EMGwblipfa8Kmn4zYpL/u3tlbygeSxCoNwGPB9a5r80LX5k/96UBtH
sohSSorK0WlW3O7hf0WJZ2tS660EqjDEYIpY6cLLi8+vV5+ueuLxik6wVQ9YJRlF
cEwKebAnD9UG3+t0PxQZ4F6biIYuiPHzulc8401BpnMkexidXy/rjm2rnI/O4Uux
e6Y603bt2YitZ9aqDFNz+P5kDMjzX1MRZoQg3kgG1hz6bVIOZ2QJs6Cf0IBLhnT2
rujKdyjW7vePIth/UMxo+IBOnDw6iUzIZiUa9TB0MaA3IhPiVZkQUT32PFkhztAs
bAE5Etpft36OqCaNudosxuYcmXtVDUEbhuiANsi5t6Ob1fvf9EhcFfdKlaR2bmXy
JjSGXuMphWX97IXCP8EvxK6hXz+m1uysLBINtNak8OY=
`protect END_PROTECTED
