`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9Pi1B0EP6ezuwSxZFig5MYE7msYkzPOt8Q1amlhNcPZwApfqBit3Bnm2TPu2Iim
OdBscNSrOuSvrdn+gNW7PUiHUAZA2LD3/T5djSoHTqBqo+QBGGzYXtnDTfkCVeHG
M/redbum+J1gX2FKtZZbqwW8Qk2mgi+Hidvc+513/jsbicGp0K2CteKiFvj51VM5
gy+a1UonXQ3jMmXQaiLBzPsORZQKCQibwrAUKGjFTFIibQzayoA8V1i3lOkQpOYY
t6vhCmVfVLRD6jhQYD1+Shhs0uiRLSxh8WQ0+taZVCPu140rTtfHbxCzVXWE9u+c
zhb3DRSvVQtMWYPr1i/MhHBmPelny7zFZfjMnyZ8NDsogJ4P/x4hOwr9T0hZHVS6
C2GYpxg8g0IRZ56/aXlern7XbGI8ZKHt0rQzCQGSGGUzkcFbYZY6LERZh8uPgHWa
c5A+E/iR/rggzcj/idnrYWscAUKLUYYXhjPBcs16V3Y3crq65NomWFhTXwJ4ksCn
7jFNJFLn+P0SfYYQsHFLg6J5vYf6phuj3axpzEzY/W1d7pUAp4TKJjtMWh4Wsbzq
L8/0rEwxPOCBxJgIPKXA3KfOs3g0YytbvNxlA9NUdihNcGxFhYPPHK790Eei+fa2
hwV7cnYXW8JJEMESybrpECrJyw0w6CRVSCWHJWoezKvJCiupT7Ooof8eAteYJYaa
x5ujtt3Q90yagzuHRPRZBSZZtLj0rVVOBcSiUzgtkLQ=
`protect END_PROTECTED
