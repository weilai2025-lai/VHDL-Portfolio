`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPjhRmgpv6n2cg7cVJG2HKJ1LyVxh32LKmzuoUJIk6/ZlKDslflUroOYBV+21SNo
EBeihmcWENYG6izHbTLTBx9mr+yMMbwb8B8uT39ZUcdZxpkqTmSHzT04J1W2oV9Y
YK1UGBzlifTg9kZWffVMymt9q+OHSkIsIoU7FWWLyJ+x6v54AuPSuLkinYosbs14
0lSiaLVijo1cs3GZ3MVybnhtGZ/OyhIqh2da+3h0Q+sK96Prw4MvQIQfQghEjrfn
NMpO6Vf6IYbtgyBgajMxU8dC6La1Wrxt76eQKCTs/TwD3SyqbFhL4YTsZNkfjWbG
cgKpKAM4ywMl9WhG3DmUMWHcpY24V+fxR4dJeB02tYvkubB+iT+xVRmb0lyZP2gl
p5oohY4BV8kDEj8LYTPH3zqs49bBhFoilAosIykSVBaXvwo9hBWDlnvArWTJFfYy
X2OP1GwIiVWEOy/PMgP7b9ckNp0DTBr16owMSB+N1e1h0Zq5RacAUeAIVKjSoTHR
4T95m2eVkQO1rlepQzjIaApNvjv+h5lhyfLEGkCRwaE5XhlT6Mn29sr6V59nKMEM
QK4rP6btvHaD8xMsFYGLmRv1S5wRWN7YxwCkkbTHsFrFTYDb9cgXtDvstOUUb8sN
R1hhnixUGgBm7W7ZYorw72DnqFxkuLbPjpF28HE6L7QVamftsZjnjC1Qq9FIi3VN
ttkwDE+klN8J+p/XmpILHqdflXTb2UbuiESsgAVJXUZx088RJQBKbUnY4w9EPV+9
7zCXfz9GrlN1y5IJ1wXoxghHhkkAUmAdtqXZWpKalQPxHsyb5k2IrubrYd1Ixh5w
4dH5vz3OvR4nGOV4PTPUjq7xvYkyRbs+05SuXJltpZ6JfA9cJwmy0xV0HpdsSdH/
UPvH8lpu92Bid9ZgYWxdl5Oz5ZQWYTUwEJNyF0+LJuLbpqdwAZ1l9zb+Uf7+JjMz
g9m2+1MjjO0rL8T7bXTVuKUY7IA0PUKsDgTah2r0XZSXeL9ZLAsEMwmbFQjVhbD2
ImBWcz6JSYUWzHr4wMjKuy7hiaxjLhV+lQwn+Zg6msIP9zNLSRdqYt3S/4ZA//DZ
ocvEQBXgsPewCpZzjEL+DwyS9NBnLnfAjHJfHmzu9XPZ23jDrsTL04m6DKEmAbO+
jZviipg9WpL7Zt1dDAOf7H1r7UX189aIk3pPJiHbl4uZGMW2lTynwSbkLHb4aNG6
QxBDDRurhhnOsAVrBUw9Vi5A8sJcjgzVTa05pAa/YOWR4eb3K7FQ4sTRMDcnOiJ/
`protect END_PROTECTED
