`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bK6DT69f86aYbwjZSXNFItm0W8eRA8AyblzIPru9WBVaIfCeFaSkGvJnNSbT3gOB
bQw84fttYb7n4+iFlhXkwdgeGApHb31GbYTGFfttnaHINU0cgJPHlf26EYWp9dCM
qf5ysxraI17WAxixV09TORpZ5zB//hlLzpqveCPQTMb4j98OQlh26s+YodyKzQVn
qdLtZPA/rGfXS1LNHNO6+lzompfwYlvH5qNd13zPf9UxCbPa7uTYixvvSFD7PQ21
FLjtF/o+0BiuPRC5q9w+rQUggAgsqlEGBj2BmK7mS+JsoE18LRJuU6q+q9ECCmA5
j+i48P2u9UjYAyOWOHem82Y9Y9LlnaEAXVLK6lyb3nRhDQsQsj+DfApY6uI50jbg
lj2upTVBEep5b2gYTxU0trqU9mM0QzsG4MwK35rr9o9KzlXjHCBAAZ74fU5zjR+7
MXfcwLWkdVkW99jcW2633rFIBnMUfNvruR/VlNgTNRaAfViVv3RGv3awZ/U7M/qH
aQYfya3iDaK8bC9Y5L0aJFTB+Xo8cBXIEayCOk0rS3O4RVAyC5AIJdEw3eHJnqdE
ACj26Q6p3CAM1krNNbngLM3lkRLqOhDU2xJj/fDfX+MH580loHXFI+7ZJJ6fDc+i
jT9NN7mWuSg2ZfQ2dIa+ISrNF++cgirIxe4EaO1YiPPWcKW3ZcAIWwRIliLtc9IS
Z6P1SJe4aaxPoajovzCkEycWdBPhoJtX3WLB4U9PxK9DUdbSViAjjHxWSB+vboac
aE58ndAg6Nw85d4FG+R/1Gp4R0VQwihv7v2AaKP5k84i2Hh/0EffBnT/ElSMJwA6
PNj07moMzZOxJFmzMn3UoS7JBAMLIPBWayEmEu9HGzsAV7+Ev/KAkiHuYJOWwRrQ
5INc2ZfC8U/MR+QmTTyQTPgLR9NB4KyVQGCFM1EbvMnjzM0HHZzmRQG5tFZQ9wwH
R5jWgDdlgplVknRpaoSyJo3y9EeAcJiokY16OHQEp6/lKBbpbgTOW+wj39I/2OLB
5MZMXqjdgzjTvvUXd4BtmiSGVT0lNZT97aTS4fizwTOVLQgvw3Zsq+CvugzG/6aJ
r5Qg6R3O8Qp1amL9lirC1qgK56sIXTr9TTfyl81veKvpOci3TTX39Scz1+1MXWWY
aQKsqEq7k3902Ww6XZUEwAHGOuccC0ho/NuI7A9LFwFi8kol5EBWcn7jqf7b884z
BIWg0k46IRm416MToDf3Y6ttENleF4pX3S9/3uIuNsOeInEmYsKaoe50E1uILVFv
R2byKZcxUWhnh2yB+7R1ceypV8XC3zWkomS9bZVQe1X7w/bIJ9BsgeHC+atHjs2+
DpQS40W2WUO6diunXlJ1TZ5LgrgJxKJw8nrACyDPSy6IxuZmJIGhQ4bNBQ2nfyzg
UKxaq3SayyUK+RjuebQdETpbO/HKPpN9VRQjVF0+vRlrL+fh4HYfZfpGBozt6kG2
1hY7T8fvympcupGNv7LMHsNjPg4h2xe3oykDggUH9u1fX09G2Sd0QeGMUjAWrC5D
t0wlrQasA9tC2YL7agTJg56Qdm7a7HkCLPP6xWKZ5rZZePSHzwWyIaGSBRqCjg28
CYNaEqBGVbG6pFB1w0Sq3uAXDa10OE+d5n31+53i3rM=
`protect END_PROTECTED
