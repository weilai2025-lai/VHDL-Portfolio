`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nm1izl7S3P02DCUXRcxsAyaM/8ovUL9HecPc/LM1+wv75GFVzq9UbFSv2n1c5Z5
tk2kx2pyvS99hsJnWDCzs8K/A82hGWUdZC6oYcKkkJ9npI53ix8ow0uvOTzqRPUd
bjHdH04Xi+lDw7iSpUSp7LUx/tuBNJhxBIol79FFR+9c7KHUhXVQJOoT2YZO30I3
RO22ki+eTEhh7A0tRupf2aEkN43CN41ieyZwrdNFhnVoDUA35jva4mg/LWD2KYew
SpGeh4TrQXUWMoUHvMAdYPn+JS8r60bB1KR2gPzjcbUYBhFcqk2NUJkZr5kRiKm9
6KLuZu/XQau+d1DBycEEofz0MZXO3P+leXZaE22otmHMtn0DDk322JhClZhDylSs
Q/Ay7jmGJK29BwmUm5r5v05wL1Q9FtIxVqKlfWej8GTFxvn7R27o/rEuIV/gv6R7
uceHcVT7Agcs+ZbMtiWc3R7CQQ0/RtjXBre8c8NksFEZtoRHZIRAlJbGqhlqh1oK
CmL7DwkWl7TMuveQnx9oUzqzX5LKqHdlFajUPM0ztunF7nSFycjwR6cNLX8uFFTH
DFwx6za6kzgry0DHcSGcT1NM0zQXO1pNI/g1F3EWt5vyG2ZKRX9wiey9rI758uLV
PTt4Jh9xCqJ2qsH9OZsLjbYdAvlLH+zWTbxAxrNVBaYtVaICZpt4GXVGo0xJif47
0g1chwGVL11oTRtDSbtTkqbkT74ExGZU8MhmtFtAUoZkv6K5Kit33Zt221QTKsT5
RLtFa/z4TrDZPQ9Oxpp+c4Vd2h8LydRgAj3R/qFFNlR1KRYuqd9Jqfpvl3j4o8/H
aenDvwCs0O2FPRHGAz/fiFmjZw16M/BTqfhOmSrMpm7t9aQjO89veskKOMRk2UVs
qrlbcnQLIKtRQhHR6sUmMEnqAbTn1G8kE33KpWci02D/5yocNPR2Lg4FqT+T3hEZ
PPYjiJhGvWaR3Cu4HlyBsHoML7BfbVzqy0duFnQF7MDkQwF/r59/b4sf5LO0+2Sq
I9UYysKELywWPCDNUSUv+rIbiEPC8eblRQmqQfYw0uRdurHaM07tHpqEOG/EDfgR
3lSxLNym5x2TrTo61VAAISHAVS1U0Fq0fI0eGQc2sfDYFBt5m+Jhymm7fbKBltP+
7dqGSwXGrOYjdh1gUGbuHnUs/Rzu8vO2C1xhN/iGChVcZGc7cBR0rG6ugHmfxJ6m
Vu/y8vw52TJjj1AeUGyIUiny07flot1vhsDP6PAq4phuxi8sk7nWJfwRaURlYJMl
BRmO+XP0NrXLkxbUzIlA+yWBn+8Ez7YZV4BWr1D+TpnLX1qF12fFlwfYkA2XG35n
JZM2qmfm/iK1G43HY+vfM1rU5w+X7ZJoykWhJBPhz8xjy9bynLo3LVCkGHsLRs8I
qafHK86ex2mg94bXfrtGaaRo/7hjfOylks9EuQWM2uKd59h2Lu6CdaP2e9xKMivp
TDVIyqTBcRO+BGmE2NBvB9itANU3f+KdQcnLPrRpHTjnDeZo9qVMhdGKQlQ+Ero7
mDzHQp3+I/PiZ5ML2IGs4lWN7DVjE9jOqGwGkerYVj04XhBTNF0XIpRR61sSq0Kq
thoBL1mqTrQ9qkDeyquO0hVt0gvcgy68bCnZsbhG98KTFBRKcdTITxovdBoMZGvy
DJTWI+bgXnmMWs3rKLghlkrch+ecjyZFAsr4R4GUzKWQy8sIjy6epeU+AhvD7qQn
JWocrzQby8EVqfz3BM6rZIxjgXal+15vV2NfG4jR09L9+U489cYXDwizc2L+/DXX
DupvwNQARG+5Kv/E744C+nw2iZtENyKcoA1BjqM930vYVwwC82TcPDoi3Uk89PM/
Akfl2Le5y2dTBn5y4vqtfKJov2pqbXin8e0y0gcWkXmIjS6jiLIA1leeO4qruadS
8awlkHN8sC7jJGO/tgmaRVvuPVtgY1CGWGWAjw8D/TjbWXm57DBp/7MK03EAEAZE
tGVSaPhFvCPxt0QftSkldRggp6xGjZULcjPsrcIx8xiD4errdqSBu3zVfdyg8v+0
w1FGWEQlxTL7YF2U6p/eK99V/qXCbWXF1aWK0DcdFGzExdK+2mLY9Uvu9Ss+mqhG
Lmz0nB3WdrtoPuyTHyVfwZqm5DQeJPL6hB86gaaFQkdNSEkmz1du6ha3DcOCdcFQ
oS9HooMNZor5UOjnrzx6ZdvcdCsBi0QwJlhAf2+YkR3OXD7gy5Z6YECZzKUQ6kIz
zw4J07SCgs0c+kSfU5eH9caS/XTbWhNZIR7w5Qe5f60tsIWcJjzHpB84m2cWSV9n
TD2nJgx2pzKq7onLMIQdA6nPhVcu1xxplv9GMJ+OWhLr0qbNHA42EnxRI+qUzZpR
ULvnuKNRhMxIUk5iylqvwmLzCx1paPlunEE55Xmq3fL4r/7tTgUuDaf3pk7c1r9R
mqICUiYVDhx9t8GvvdlOYeN5lFQJ4lyJZ0dAtQpMSiE56gnH598f+uYSAetctdnp
JTiXi2q99c15Nbb6arLQr9u/VlBHM6SUytgYUOBhNToZFm9KtF1XNX2+Rlpx6RLX
F+ybDwPbbNv7IA9qZtD5D4gmeGtyDI0ylSNut5TzXaOd6/dLXo1iqXzvfsNXTlFW
0m8JMTuN3/g5rL4Q2f44a06tsHXBoB3hn726NDzoJ7vZ5QbNf2Va9S+JiQaHS3Jp
c/Cgvc3wRyKyt6HinWqUF2GVZ3oP/+9Y3LgRGpAwDCqOtsuK+XBYiJ8V6NbzRyc+
BOavVKIkRv31/ayjaGG7NNJJhwKaXNmB5+PwLFbw7titd/zYoD9rq1XF3XXURjHo
7NV7ePrVl0vPlJZeUbh6UNa+zGhNKC5SV5Z9/mgIaAR7fsySGz9/L76Mx/qmT3h8
rrNZew6E1k1mcE5Paw7WRBstRaEkdIC1uXD1FhaVdMXFsfH8vKSGfQvO0+A6ofGm
nQularweE04VD3tjFu1JVhOx9YCZPFGCVwZVg0yxjG/4shVNd9bEqaBir+FMIKRW
P/oBXJSNFfphR1PqMKKLrPVPo4fwIFMhVAclxWAKQT6+X6yFkmMLL0FK/xOCys62
JDA9iTSgBzV0BT7CpJI2/qT4LV2dV9x18OchqFlMwVTGNmU6xZRfV44Hn4FwIb4Z
0Zyhwr7nfnw09lq8CIWTKCBl/5JIo8wKPQx3e1bpM7LP3zcSs01aXxWmhpvG4Tak
f8YWPQ/xS3OZPNJF6j0iASCE4Km7eyPCIx75UTB3OXa4cvgiO8U/vZplgEq5d54H
An1r90VwV4EI8vz32vghkZjhUWyfA2nJGfhyylSXE2JmknEY/pjDxa6rQboiO/yL
+K2X4F/7/hEUik+2nUkBmDw/qwP1c0dvSmqEGzbQSECSUEmBsSFqgFK6jrOaztQi
W9qwv6Lp1mstEBupNFlfDwqQ+MzMkuSDudU6N8eT2o9jLc0FS7QXM9umD9xSC3J4
eHiWiDvqCx3QcmyGqvY4fGzGZp0DadvU5ooBqANXr1gAswR/ZzdD/lIIJAqCQSqK
ezwbYOMSTqSjCdQI1Pm+4K2ylBtSZYojtVBU3Jx7KRFS6STBpSW6EBgnHWvpfcZe
FRML57hIEBuU9WpDKWOikyQfyWQhDSthLhBoBOQeWpJc1qIiZphK/qAtOdFtp5nY
Gp/NSbSuE9Ku+8Po1gvNVyH7wb2uGCfXtAx3fkP1q+Oy2GzrKTa7N3YBUVI8gPJz
uTujr7QtPIc1XQGlChgsbxPIO7IGJOPTh4Glilwv82WXCI8v+RUZoRqKMvlOjd4B
DJM8KqxFX9ipbXxsN02chrapc2TyK84WAixF2P1g5ruZ+uJKFoM6y8lwUOFj7cIh
rxs6TPka/JnMovbg2O+JKFzZoq5WmlfELrXgD7Xi/MWsOrFbwFemWtCEW9Io9Gi/
xwaEtK2uuCIR3S3kSVz+JRUTU4AYRmECZFZdfgIZCzMEpfwipcO1ZtzxDGteNOBB
AWvnW+d1poNB8GW8ECp/lgxzTv/1M34aqUauTspQiQRKCe9FaMaNDJVGwLNl0YBO
AyFsFLxDXmGPCpQcGBUFOY73PN1quuM8b4uiZG+oaPJ+88uu8Gbt+OFWMv6agoZn
o0xDsuhEY9vy/yXFYhqEJgtaXCZlLY1m3Ux64Um/cH5iNLOE5sG1GEmmDN2395U9
gPqshfXiTZjVdTvkc8DLwDh9/tdLuK5Bb3KCijHkP0XoBNBFzz4TaowJcydWgrMe
G5qnULnK4Ue7rHiUVHt6GYQId4ztR/suT7m1075ZblEToEj1mjCnuArjwba4AG8e
gcKmsF9IbqE1FPS82nBp6Jiq2Fh/NESMdG4D1iUU/CFRzXsEHFr96A5UbHp5rcmk
3+jX4CT0A1hc/ViY1p951BkMUvk/SihpYbXwY59BUEVb0zfZUDKIter/NFPs9OoI
0CKHZ74MPVsEhzAcsEyPu+1C7hi3+vS6ZWpuLKzts8QH7iUvgzfl819o8fx4vxOG
duacfy8qc8KDbvjT06f8DU2rgRSxp6rJiMcfxzLoRIMNrAZfoLeOmgTG3JBdYW+V
XMRcl+J/TgU1mp565bZCnGf3chvbkT3KRY8gCOynFXfHuhMtwb2qlm1PzM32+NBz
DcWDJLstso1ozusfH7fZ/5XughtXRv3kDt0QmPbYNFrx7kfMPl2prEr1Xc7k0Ggp
YjXSnz0CBjiuTrOTGpHjCcdCD96CG7tuJO5kMt+zHXxnP1Ul6q8dHoJ0/hjUisEl
yT2eAOw3IRFUlAmi+ajXNXCNxkIqr4E5Z6CscX3d92KQNUOnqnwITvpGqYB0wo0O
QsnEzrPwJ4D5fnQvooUZrhknHA2GtrknYaY/oIr/C08Su0QLTgeAQovBAduvPWNy
/capCaFSsVl5uTq/XoeIFMq1KGlS0HgtTFGu4e5UWwuRDTBrQwLr3EPrjH5IKmGj
soXLpaJsMySYyyLlT0wdpD/zEdMCgiL1RoL71jSgPAE+BDElU+WlSxydjX8H4Enz
gS+DHdNFSuqEph6g1/GHRoKjioDHQYC3rfDT+qJ3vexJLqlVoQUqJt6G5czdFS9M
fKiRRvGqHKdyw0TnbeN3gA==
`protect END_PROTECTED
