`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SdQ4QlABZmJ1pNxbFyCvwkBXI7y/bt3JIR34D7u/ks7HJE4kIiEcB18m2WC+3fXs
7zJAIn3ZRyFTEkeWaFmHUQ5iWh4VukuTfU+4jFi3yGBMvElr6kqWbHOIVg26oG1I
F4NROPsSiOL32YzigVLxSv+EHyGpXwqComINqhbxVeyUvznQQ+2Rs3wiMSlmqQCM
rVjn9iJLrRcIVE5ybjDft49St3t9FUl/vh8SMEKlStxeua8jKnappsBBeD/mwi5P
9LgpVW2rGH9nGru6gUNeqAKATFxsl6abyXd+pwqX7fgniml02hcKioV02CfjHIAb
mYuVfjIfqV5cuC1ItE6bXeBFICSvcAY9ceK+/PJZMW3bzGp0Qo4HMaZWw7fJytf6
SHDP5WfI0m5q1roudz3ma3w+q3z5rVGNmmRT6nTZu7druCnFkcz85UrLL+8kA7rt
mjYA3Z3Vsmd3dLwd57aqkcjfocK/1jLxqtRQGTWsyUYnuV2gLBs5z72zxt1HJN85
RidMtUe37M7YOQ9RA1jRyZISlgAAVyaZKVKl17m2lkKdP4smiqB75MX2kwCiLGiO
8YA/ZJVq9ugUQLjUVQ18iD6+iugLdwVc1yTJ+Q1fSnWMeupT7PkkZQ2/3WnUM1Tt
mscD1K7BB4rOuoMIx87kIEPClgrU0G+u1uqM4LH6Z152BDdqXtJZzpvxZc3QTb+W
403WTxZmKmX8rL/114rNiXDed5v71s0B6uayJ5GZWJBJYU5V/hn5W8/9+4qL06x4
VeUuNyK4haNnEygNJRysKNPjhJd/9w/qdy93apOQBf+b8WsoNDTutBW2ZGtEGGsk
iOzySfeQQXXrDhC0DFcyQgrQ8hiuY9Z9NKeBU9eUkqaV+IRh6C+sm3HV7rwwBVp2
lUROA3tHcPvEgVg/z1BbYlhJsHWOPeUFpoqrWfvW858zjQqIPmfmJdvE0C6CyAS/
Fb0NL6n9cc+haK9dFmpWaMrx/VBBY1jYJXUFG2x3UqZpws6YiMrt7ZnJV06yu9Lw
px5V9XXrrahbVjHFeAf51H/I6PQEru2nq+Uax7dEM2t660Y5iTdB/vxIyySgOWm+
mJWS0TKVjQPY1Fpcs9xLi/C4S3CJcP+i0SPgxl9qcQtXKRODcTO8P8/8EslonoNq
xNyt+MvGQvTot0zhXAUai5Ck/6SRNk8c7VWJEOn7eoiS/keTgSm3pO2Kx4X6TUnw
92igd/TTczwh5K1I9zZheDchiMaM+pfdsXgca1Xke1iLGni78h06GvF55rjsR5ZS
5NgR/iN/HuryUrtuwu2jheiooM1V8tRyZs6L4PigOW6+yOyYJAQmOTNpiui3eA8C
AHHsBrkwD8XnYEizSv0lG1Obl+6LqPqK9zocBeacg1QlZ+rbJTT+rDY8Ax3lBixg
BHXrS1mIET/Amml/AZzMuqAD3ccap1B3UFdc/3MFssFo3o8tMYkQvmccfBZm9iLE
WbtjwWkJgC4EVij8c+jhJffUYbH1t1F3Hh/woGJpljh3pXDtsO7a2Y0aY1M/OWw+
ZOmKtRXjLU8IADGu4BislV67q17aLU9BGe1kVym+dwYRL991nVfjznBjxKnxOEUD
puiWHodWByNkTkQoJ7FDP+w4DPJEPBYt0kwE31I8l3otarj9+hNS72doJDJ8X27E
MQbMrxbaStdcIqqhaZaMsb9LfBb70Ky7EGUySAwcSQ3b48aAgEu2zeS8K27QR9Ku
7ivhVFX4YBfC8bXg47YUVs5FoRgywq0sH3oUnmXcWZFlW9iyI6+OqAC/sM0lBDaK
IzRXJAjROi4xrtNxMSuPA+bDVCJiIRFhvLlLkFDKHxk3US7LDsH3Qlps2Y6UxZJl
ItoAfFxLNjaCYk3wCFX0pj6YmRCtaZXOrvVKhT/LflzWZ69FndXErsHKlIc0XPa9
V+/NB5fVZJuUT26x+uTqRRvaQx5d3PEC+vdCDNbqt2C4vS5fRIfVHIx07nLRFHvf
wjIydu4eAxshvljhwTsbEKV1q5lYIwOSrNa0D9VDhcAleTzKSxSRFIuW1bMc/Zvx
eJtoBrWXf/vxCEDOVQ0d22qW4x9y/Q0yaXgyMRhYcYspYiB9CO7/6xFVm/vLP2AZ
HWxe7MEXQ/0c3CeHbY8UdXa4OL+IXysi6VPJqSxFIDY3TtJau22BBu62Y5r6bkeL
ImWK7k5fAzCE+rfLIdc0QmH7UHjKIe8cM4hXZTfNESocN5bLdsjoGRAocE7PELTG
fcdEQsZiGIS4RF9VSx+OptWwaLi/ggWkHx7MwYPhMNf/gO05jY60nlcLChUtG2Jy
ujjpfkPje04vng6oWgVKcVkbUYStCbI87d/PWcuHy/N/sB7plrzj6g5AYUWsK8zq
CSAENNqmXWjZ5yL4KwOzESmaFa9E/0TiRO8Nt8jAwxQ7waHpC/VPsDiGaWiAX3fX
Re04knLCIRyj6ywyDPOnNM8UPk+kTIdpx0LEsjewqmu3u3TT2Cd9yY3viEsBMDKK
L00IZNMilpOyhEkuA2bz25JlbU6B8jm8DhNkOutXZBkHKuNF0iDiPqquUXOpkDDM
go6YM+uFr+2ldR4KGg0Y1dgDTR2Vug17HUdl5FOPoy11h06gnZoeqc77U8eVL9tr
QwIhMG4Zd1aqvAOKpWWrcf6JHbGzdPwb9j/O/g5JJXPp2496rvWZBB2sGXogDrZd
YZLV59kTBE8HQHxxAclnF2KTuv4/E5zWfXWlKVvH7+DpUKLIoYlxZvW4jm8hI4at
L+t7BLNYGEp9tbwpDZTPKHqysfxvED+EKwiclaWeAIvYjrCOFIGB3IflfNIDOLlj
MxVlbhdBnC1SkbwF2HVl10VnvhrWr6IYUd8Kr0rJmooSzEWVL9pevp6x4MGza8P/
rE3Bwhuc9ZeZlUPSV9XehMXPqxaP4CuNNq7S7d88l3tLvEL14Xe9BxRtC2/PZqs6
sS4d2iWZwGD3n9fDnNa58yYPG8m4axKxfWAar7YtmL8e0ZjxeneFdFi4GRkz2Qt1
N1pDbqIbnK4qLxrC+6+cMBb5CtbFjAcPDSeu76a673gC2s2DOPlzaO6gpfy++DpL
rRi9ORDFbVt4UlN7fMOOhbxXlFrBcvZq4J8UKXtgI45zxPr4vBlvmVfd5kbXl0JQ
iPK0KjozLk1YL1762c7T4ox+oLQG/Wi61f6RBuwRlX3xYAoY30mwTMJS/q/uiBrW
b/d//V1qhpl4w7dYBRoI87AmqY/BmKuVMN5cVFi9J1qrsahZrlh4aWJzmRzVw0am
xtUC8j9TnJ+fAB7cwRz0R8VV/ktV1wakTT5rn6BQBiIjhh6GPrrUiVQiQHzr4Mz6
izkJ8Tl1vQJpLvFsGic5jjBSjv4B1GPZwyRY+SjpTJCMAcBQCLcGXhRR/+imIjby
g8CLK1WWxJKzMfJORlpsqcOcajjviJwOIUU+O+NxAZb7h/HPRNhcy3AiKi8Wmhl3
1rfEtCb8mdq2sddw9JIZ77ObuIy0pmFTZjtu1PaOGlS5cPlj7BratbOxTI6C9p1i
cmEe5urtbgM+g2YK686ujpfWU0FB6Yzu2YD3I+tNTI4nEsB0MbXizh0U5i0gzJBp
3iQ8HgzYqBBnooe3jtHz3Gvna7pObO9G82RJc5kLvZoEr1iRRMFFI1DNbWF9EPMD
7H91ygKqE5+OlB40a+yLEzA5cJKPPWMvaeAINx/uSd8iisHqgFI0KXKnz15Y3O14
pbG17zQeK1ll/Qi4nEJVwNsRt66YI8S09H0FUXCViiOPsDNFRPBvVzOn0r+mbsU0
PAz/JIP+CS4pWi5kwdfn1fueWZ+N1MfqFuHy9GxZJassTNUg9WYorBlwxWgAJHnN
qjat/qLc1Tox4OKoo9AqR9qgbun3pNgMPYxWyi3ItKx9C2E91seJdYc0KwngSBUt
dUTMf6tqpDYjkZf294XSEDHezZw+pMzio4qQhoNmXV+xJhOeQtfSftwl/teEAMn+
pQ8J7JtN05VrwXPfiuotapWoa2v3Qw5HsvV45fDCR0Y+gx8rL0q9DyrYp7KMdBcr
1uGvg6P1QiFOZGvkbz2E0NfbYNL8LmLMo7YuQ5f52CsLtaGSxLQIMWTCT36ISWkN
6Z0qoXVUeGHTRWE1NsthRNSUZd+WpbTPRgPlMCvNSStR5sf0akJ+YL9/3v2B55fY
jNdL7q1MkQDd7V1uaK2+QbvJeUG3RecXgx+tM65a5ZafMPi+6sbjemDfoCvTKxFA
BlntXK5X5rNW+L7epce8mKKY/Wr5Kt1yZ5yw7nvVber9PXwMPGxb9lslvpgt/U+X
rjEgAcqgJ3f6cLRur3Nx0ktd0yoDpagHG34/TqAwuGOVw2XUdaWfGy7cLNSeAIyJ
R6NO6hyeV+CbiybDpZqSoYzwkgIEUmdxVDWIBDq9PpLSHD8LAWYUWdmICgW5OnSU
u/Wmj8uVuQjxui3+WtBs5C3fbAM8h9J0hleQsV0/Mej7r5X2ubRGqn4S7kqqWzB4
CH/33p8Us8nGOEx/eP+BqFwnikzCxCRM1jzOggJ/RpFMtlYyHE26ic+Q5iw7d15k
YEppJV4fl0W7Z9JId3f2AAKQs2z3h8oPBHoNRJYgi2/gIFPl0iU4xxIa7Bg/LCNe
uPRXI6hhCxiH/azA9O1d+C1ZwWy/mjaRYuEY6Jdm4RurgZfWv7y92xJxWHjkQf6/
12m8rZ7E/FyhZkGgtEq/5B2O7kg3h5Op9KKxTrn5BgSQ7sypP5VQST4Hc0T0iEAW
7eCgzH4YtOMjgdMBbNOLp3dWDiHUKSNxr1ynZFWu3CncPz2s/vy/a4+ZSPILwk5x
dyqzmapk76GcJiVjMnqJcjYHUlfB5MSGujmJLRYeKqvecRPEhtbpr0k3kwbUdwaB
sU/uF3BgnZZzUw95Djqv535bZtmpiyUx10H7+ItF5tZLwJQp1vA4EcjIO2iUFj4l
5cRygKwCPAS19EBPC7+Ksj4CAFnIlljzObIe3+sPTR1wQ8JRq0McbIPhksQOVYBt
84+BU3jWK30PlXNt5S9LmeEpuIVo2M4pFhBGP42mLvHzAwFRntl3b/lBfnpkX8u9
n9BxupkuaOWzuaCJplYskG2FMgnTwbeHfiPB56WsbqdG6QfKiTA/OYaVsicaBiYM
ZXX81t1nLFZh0X0d/fP7IPz1eBVhdZkQ8Q2ChvUUu4/vVavn1MmrOKBus1QkML4o
veCMVI3iQe5V+E2zwDX4wg5wYGobM7Q0GsRESyUeHpKnwH1WOLKVJKPDnXGxeoQD
Zu6Qm9IV975d9GZTUyvTD3fzJw0UDQE7EBj26ozXMRk38PMWp5FIPLiQKP+OdQJs
YhCglA7ALiLST2B+WcAZNYJyrS/+nlw4UeTMK4VsS50zwJZfO0tKY0oekSH2SZwK
pgrAA8lxWftv76Q2t+S2u7KQZiVZGRpm63ojq1yyiiMYS0LjZw60mfoCbB5cOlUF
DhcgY5iJiPb7U1FYLpoRU7GdFcKtRYUM+tGoLUneMRe/or0eTkOP1oid5z/Nq1BX
4ty44mITVdJdQ3c8OwPNvqLLUdZDOOt7zrrFvDLtRYfu5lK9hkZslhQw8kK8ljGa
Sp6O2X+1b95iiv9qYDAKiupLYAJ/GYwp04vCkukUbBzPTqFEMkYxhoUQN2YxIbP0
p7upJN18OeFNkOxu9YPJL4JMQ3LvqUptjyfrocX/H4kT9IOq0KOirVrqbDEMWyVi
SPywWK74NCxPb5Hs3laGlevMUImLIcgX+i2WkSABBWGuB38cIDm4aOqyORxHMVIi
NSckAU22RuKR4Z2YeLc8pkWWH3uC2sd6zlhWG1t5LFJGMPPmyq4leaj4qGuhHySe
6R+Owu0drowTLrEswsnkhn3tsj7xKqemXXECS6hqN0sfF7fhHHUn5ikAEQPdikoR
jpY+PStUzWs2aRgQbZIkw9VvsB59PvQcDhfwDQDI4fXmSWXir8TjhUp9yliL3Wqk
IaRYLODQiYynOBbEgZ1lqasZ/qQm0fUO6G2XnbN0UncW5j3VSOnOpU27OMuDt2Pl
bF3rOTVOINE7Qo6TpuIDBlK1okwMEkpLkcVl+kRq4iFpNMJqccNVl7cIk544hrID
m4ww375rGS0I3QTCBkkD9+00CwAi5q4GMTJxRQC4+7GmTNnjyQ1JerSPHiJAuTcJ
9Ht7NW4gV4y5Qx8roJqSJKBsNw8IB0qKsr0x38hzy40dSwboYDVV9qw4NoVGNZJQ
iQGODgnOae1FOhYkC9vGh3g/cuSojSCj1qBAjiUpQHCQp6p4m9AO82BRsP5Ge/TZ
VAIdOG7sFBFAvMGDjnB2TWSZ1PEL8RJM1V/v2sBPzGW4hPWZkkZCwPAk9RKQM3Y4
bKsPyXMdj2HR/gV75X0NGQFHC6rIBnyGP+ZARY0KdoWbZa6eqm0d2oX6bsE8jVfn
+QSp4ApOjuDj27rO73Ridw1ly6jrv5z4+2bgiZwUMTPkfkQOl2ycFbojXkz62++t
rNsDJTaxOJB9w+N7gZtI0OcOMEXr3R0E1p4olmvHlthKoebYkNB9+DYua5xoXr2N
jqqZonEwLg9ULK8fCBc2EzSoOQlTzOosHKi4FpbuxOERWFwOYCf52PWX/KCjqpm0
zG9LDZem9g1BmlClScVRRPNWLPhR2qWY+gd2k32Lcx26n64x/IOLoNBfV/zXawUw
U2hpVc7KVNIrESZ99x8FtPE5VAEUeovQYvLlzNOUOxnB7NyTcB85lCwUdoovBGfA
QU/DsY1YmWgybEKUrwuDufHwJpsbQwYoRqxlo03TRPUyd291QR5zW07zxx7s3/3h
PP4H2tKufD+95hSY26mGS4aGXW6Ay8bqSuaKeJMh5ayl8aV9EdYBL8ecz2zoTUbl
6jm/R/9oauJGjo2YDrBqZCu3ymJKKbx5vYymDzAvgdLBmK5I9a4fBgc+jtDcIbBg
N6J3vkXj719N42U1FnKYB8bn0Q3DbA+Y+IRbi0Qw7e6+dr74BOksvWgfXQLrld7i
BxtM/dnmU5w9V9OiXHD/f/KDYc+BJ0PJVx29jupU65IwUkrG2Ut60I1+/LYLjv+K
QUwCSZT2l2bnbAIjGmA8IC3a84Fzu0UjVYUrXbRiNefLAiQfyJryWmEeIl0iQwfC
drkslGL9V5CsTAKp73Cw5i0MB+jyDzTj+qx+BmrrMNTTgHERbz26vuaFC3yaz0tG
0CHVd/eWuHWnt5z9j8NHIdczHGWnLepDtFTECvyVIcKRf96A7aPI9Gp5kvfp4rtv
LrOaNiCZB3gq8sEkcOU8x5ICw07BLIFcBeSEK8AkOYJPSJ7Q0hb0CpF1GF1mTunQ
BALcOKbRi3Kok0rJo5ky/lrqIYe5ysJusKvHrwYtnEOmkbUGQAU8HCKk+UGCfQ3x
wURgKmbtxYkkdd2xw/ama813qU8QxorVd7mKL4Ru8FRZ+q0tSWVhdOy6U/tZJmhj
WdHOSMXsJYBQvRaQdcgkIKMHHr+/4yokcPZBttAfrxZKRoTlzXg8gy1e813+bvWA
fQjUZZAhVMGRPGUR0a3hfeKJbF0eVXoAQle2G0bZIRwvPOOWu8GDRwQFcmDLsI3T
segyhpVTqJ+ipkhBjmATQJ5jKy3qvv46dzXmwf0A3DlGPL+uz/TjIAj38VF3yKVO
jDL+zbXp7esD0mDkWIBScsQ9apLbE5jAs0k37jM334pelUlriZCNWZy7/2sHiYE4
naPdkzyd+s0+WBQGkvOu+nmRu2z3MSVKmalTRRifFa7OdTyDPBrRVMFalbwUu7Gh
6ppLN0CGD/wXMILo9B03KxNNLX1Ap01bJ7Egz9qWI41Y2NX9MrOFRlpCvFxh03g4
Fp1LdX/g047SHaP0+aOckezaaVJKLRTzR1cSYhn1sLqIT3/gIHt976fDGyFtFaM4
0fUsFPT9N9eylKJHn20XqM+4j1ACwC5uv3C14v35n4vlm8BBPCA+MXlwB1JTLV32
Ylei7+IXyX8D37kJQBySCLb+LWccRxIcjbfb6zXAh00360yijSuCbgmK/uiGtzt0
d4pUjr6rXm6dWUZjZpKHxc5Pyjczt6yqV8bDxmzulo/7NFoj/MeGZpOW2fADLh0r
IQcj2LRZjMGfTeD6ZcdK0w73XDfWCUgkzlJ5CRCwqmj8/LRg4T0AeWAhfNaQHQNe
IiWyfgKvlJbweWH9kSBRhfXP7hTahMXGAClFerwFfu6ts3kQ+MW3MzhGa3m0zRBr
0v2QYpS0qD08mX+TG9BjhS1U4Ssuw6gioIqDGY1tJLh7gcQYQ0qpCDyqYnySYZRE
Xrpq8QHECMNe1XE/kfocJPX1EZf0IJ/udnoVdeaclO5A3ZT5tkpYqJpN5BSasvCI
pcsajRysnmIUcXmQzXG+Ph7/RXKbs7tvpmkku1Ru9jaiPn4vmlEePJyHN1HCp3nk
uG/Ddl/nw2vGWPBdJsnB9wnahE9TAS6OwF+IskOlwMRaE1U81w8X1fS1Wk/mhCcI
qZESBizBqcP90Vb+IomWy9BcLpCUOO2F8QDnHnYLd67iUgmY+4RuJnifO2l4iHSu
O8+l0poINnbFaTEDpMEpBBKjBtBbpQ4NChkvdEiub70QMZ0dRgIS7XUBzVXLnsjh
vwDv4XQqxfmPLq96cG+2vTmPS/7FAsvmRX0QwAIwgRUPgo2tCXffkpD2tLXeWxtk
jxmBhjVrCrfDyxONnwuoHnqBkdVe3jHt8roM4qbIASf1UnnO9j7eMJGyl5RUjjVq
5gkHjqDwTp1j/3Jf36Sbc6sKUcL2xpLiIOcltxhwc5NTe3q8h4bw+DQJ7QBIfsRb
BiiIGBypyFWoQUe2oVTqoxmUjlZJl0e0CZCnsHTrF6LW+V0jj89YgI11z3fDDkKZ
G6tavPuhcKijW+WFs/9TcqKGzqN0TFhxiKq7xLPiPw4RPGf/AqMHvQRJU732YGvA
sUGCN6jLlMSoRVyKEuUfbssViqmivAIu1sCCtMqxCr0eDMWp09js5Ug/MRfF140N
9YX8APuk83+UJQ/CLWf21PbFqOSHS4EfJa1sUyEippOfmkKqBIBhBlhG4QkNPd97
TfY/50YljDgwI16PEFbB3TC9JXaaHbiG1UlxMn/BW5rW/MuPcT4dnLaHQ3ZCxIIL
MC1WWgpb7m8b4UoNdz7I06ZaAnYWt+YFTHXQMjRJv2goHsu4UVLwplr0B3h4M0PP
i2egdptEX2m4koiZ2mIaPHz6onjdYOX+0TX0KOmIm9sPkoemRskXIlaS47fErqol
0+Hn8jQkweSdukWk9g8u0yWdhdg6+OTdMRT3z7rfsL/Oq9lLPQzf33w8jvjbyini
Y5VTjd1PEUFosx6TdvMNeGwbhQ3X8KYGBLzyBy+n4rS3dpMQ0a0RJiRIxAv28aYP
rWAlBlrZQQ87/jRkJ+mfOGavN/UnwMfHueijKgGf54UOCGmgNgEfsgAxmWJutx5I
RcJRM00OWbY5+vNzDtXklLFBWEHdZgG62m9D5S7FP6T8tK3/Vk3kAwHiSIwb3UWY
zV2PZZvfvjkXlIya8yFAztfePnQWXWhEpoLQIT11r+e3fkFi6iK66BXtDWpCMucl
WvlsfTvomQ+S+jxVctXERsxbafaMXE6kEIvorhIU+5OS+WFo47nQ+wedxV8kAlHy
n89xxNanlYXbV+OxTtYS43slXEj1Ljz6+HakKSrhtPBhlhgLxApm4tWho/HfwJfx
tp9WIWfijpborwvpIBsWtJ7Uf1P29tws9IKBL0uagYaHq5yHj2TJmiCdEWv526sd
quNsdm66ZKERu4O/FlY2qmUMtrbxd9ZYc1UhWn4Vl7jJAWQhKW/FvJpd/vR0OAim
FCn3mmeB/PFlUb5Gw92vFBmSXnN8wAwdzLvtJQTQeL8KGeVeYsnUu1SfkwbzVlow
l5DxKUUg51rqUIz2sGzNnPuP6kVw5i0bCgOFnBEzn5I8+r6vFDrYkE3wZmwlXrVe
8Zgv9pxsO/GLdz2KsA6xO4r8HkeB87e/wS/leJDW1+8ogKwSoqDITVSHPG+5zyyb
qQAZjCqqpMFgYAOc1Z8paUIg17eejtrshtCR5UAoHT+IrqIYgvhlR9E4tAlTC7Ro
zZjeszcnBxU1XbYRqK4tGxAzkaMkTEjHvYFOY44pd3tEQb3k/TVZTJYdDphdNkj1
Ei4ajk/Wrrx3/ODskhVqXxkuAYTAIHVT0IMfchWanJ4EjYbqI2R7RVj3+9G1P1BH
XgEJxbx6hOvVowsHNG5WwI/kkRaI9edIAj1NfII5hX3dVGpOSQQi4Qg8tnUTfnt/
At1v94lsX5oL0B1Nkwy6GQ+8OZmyNDLgNc7ebJmfo5KPb5beF50++uAlSEV8mom6
q0Wn1BuujLer6uVsIxnq9e35QCgXoL971o4yEZrbUIrF0nTGP+w+jDgKl1tGNc9g
dtgEXnFMf4YTol2dyZd4xC1p4+PE+CAWQ0GeytYddGKtGc0WxiSHcpL3S4HuJ5ss
1cwHa98x9+C4iorBoNYiIG04x7RBmdobzUSv8X4Dk4wshkjeLODhPmDHeHlr6e+n
5FAXzV3+1EoM5RWEeYoF0hoGqRRpfGCeNslJEGtjuRniInhbk5DjE0JMF2seoTbm
L1sPFl+guLdgev2CDqJQ+HvK8mXAhcodtjupg6ybKDptOOGF3FbXhr3BM4i8P12z
mR7T85afqiB74C4KnXAlMmwn3xdN+utSW/PmNiX7cIyRDgQmyzNHMLmCBWMEu4SO
+IBVx1ilFFWkgkJGPqvDpyMyUyu+bdqGxEPygiZqNt3R89O14kEuxGkiYGeYnV9i
2kLy174Oi0HzBFGBAu8TNZFaPsE7BXWNvtS0YqLLjTy6d0wutE1hYLAR6RHSBnVS
tH2pwmtRLkEv/2fOlvK6WvLTVJzgFuzP0R996+rhjVXOSkGCU0L8532VUN2iS/8H
Cenjce/a+VSzIHZSj62FFURJrfuPowjkxALFQf/W9yk7W0oVyynL0WPg75HoYJ5N
OOvAdZQHYmivDYtkE6J32MNH76GdsIMlZhnBmvqpAHaN1cCpQ+cpeJ7/d/4kecf7
7Up9av53Gxv1zfa/pRzKqcN0+yplA9pn9JbYV6RVBGGdNveuV1KmAx2/zgnmHA3I
2qgykYuErga8/b0sTYxpxwU5ZbnFI4F/X0z5wkxRLsXU1EiUcNkZWOwfCIwbU3qR
ZTRHsudUtb2ZHHoUPhXRNkXhYbDQOvlDO5+oyQwwJyq49Ig3cgeYMbGnS6w1C2nm
leMiH8EIrENReMghGGgKcqC5549Z+Ygp93waVZSrezCEXWvL68LZqeiJs8uDn5DZ
60pilZHh6jpcj3ZWcXfdH4i5tXOt1R9YcCgVw1IyYFbBA9ehwqQqAYF7NFIOKPPO
bszpzWXyEj8O103XkeoSHkLioSA7mvOM1DOKVKsYvUfVphGfc5Pah85FQPsn1AzJ
PfnJzl+MvtK3Q+slW+9ye/OpPgk7mRXpHvOHGDlrCC0+6ZEP2xPpKmrSpotTE/dz
sorzyfiLypgqELQ0l1MYpkDYdsH9PaV9rTZW+oz4Pc73N1eDgc1hf8CyocsQymPi
9ezTNsP2xYqTrnBHFueG7jJEicjJUupm4V+sC413026ssw0cEGbYD+GO9PcSzeaR
JuqljG+8CKOlZWK0oULW0Ye0BX+TcApnKvnr+x3S/0/pyz3Jvzmt9yGajLiU7rZu
YeYmo6qgO50NF1NT7vLSC+jLBc1nGiSG7ngSLqgSjGACh+IKP9yyo5LdXEj635Dp
Jf4I0+xrqow0eoELgC8/tLE9kgGh1ZNCBKG9zo4IvfeJJnnnmt7J3n0J3ouaFxKp
Dfpl4P7zqn8/JPBfH4NIc85orYuebn4EzjoQJkNRevF1gpl98C2XpAwUzKBJfxUt
BzFOIVwjopdNYvX0RdNaO38RN/eL0O4TGpElkwbZaPx09W4PIMSql627YARDAxwk
ZEapXJwp5l8baknIOhKi8eeRGepFDvttUsFByxsVN3jM3PseSQ37d5psVM88ekPD
BQQCd4OXWoBmA0yePHEgYLL74QwI7fn/vSr91RD8wpcAyUdnfrlyPIRmBEM9SkyQ
yv1gwCdM7o5DQXchm6+mmV0QnrNqpTot0Lj8UG9hFV9oh2pnBbz4x/FegKGzxkS5
PjQLdcTMlQXjY/b00CQPY/x1sjBLuTvNAwUmtAAKLIYtKn9KrISjE4NJMlibzW0u
GivG89T5mqoZ6wDas2KmCd+o+D6aIzaMqEKBue1Pl1QrcAOvdeyp0EOunc4B1Jn/
0Um3SIfu95R7RPEMtO3vqbhCdsgNRUY4duoVIheWHOlFgMSGP0EaMDfAMyz7VfSq
RzqhuieP1xaf1JAq6rnMCtfMZqwkAVJvaJ/hwktA7LzN1M7SiQszlYwz1MCAEwwa
NhEfiSYO1czr+YmsrYkDZKkY6ma1wetgWytWixBCiXzK+Ynr0jRomCOJuX5PPe5b
7gcNelIk8E2pW7lW+4h1kCtEtH9BGKmE470Vn0j0OBTwNroeuuNNUH5X8mcHyauM
sUgVo0EwnoCSBhJQq5URgOksTaVG8E0/avkzRVkaRIbBBoKE/Su/wRqadNaUXaSl
ZsDhppJ6CfGd8IUUjsjLZxddlvsn0uv86a05CGHeFqHrAEPWkmT3Niz3JW8NzhVY
IBWbJH4MHaiC4MC/5gWCTCaEXAE7SYhreFceCXGB0iW2fXtOxLMGq8iky/5jgyB5
7UdFi7ql7BAJG29vPKjIjQ==
`protect END_PROTECTED
