`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rjdvki61O3rMkUDq90Sq/p1+TDK4DQ3T6c0w46kAMufHla8V7dvL1DDCwmRJ4jKf
fMDbpI+DzbKEX9LQc/nUVUtVclrA3MxHE0HGlZ9lmvXoinFi192HpBxPlID+Hzus
o2Y3GwpvAWz/0PX0i6Z9jNmlW8Vy+r4Agl7Obrzrh9eNBH3IXYedoWh7mPJJX7pN
YGrqsUmGOJxTx1zs3kZawtcTssKf5OpTPaqeWHlXMqI8/R3rZmnEitGtbxvNsdLm
7ZrHqSWzBqPuXgka/wy4xeiw2mT5dZihGC77XlYE/dO2byKh7YN/mrmkqFykV1RO
mgym11oY7BguC7gy/x6rMcuPyr811Xad0wjJ+AMFdoOjknhtQDxZphjyJW1BH6nd
wmxHOWR2vjlLs1x8u3tGWO0vFtB3apa+Qv/2LGHl2cPL77OpGbZiF5FGMq5Oohe7
K1AA4+Bqyv+MfcbjtGvX/0yV9pGdBGPJKgmHuWAs2MB2BBINK7ab2XoW5Ail8HMa
GCs6UXMYQxAzgx+lUCuv7d31x+4DjnK+V2RhQVH/ya1AO/v13d0+k5sQ+bjvUHk9
GAWGw3cYAA2b3+QQLVIIVYh1F8VYcdwPVbgsegdHZNOuJ9151Dy0vBOrZ6WHcjKR
1SabC+M3QAkmdPFSlqPUMVK5PvLtDtaScjvt/gR5G3DhyeNCaU4d/gFYbZtM5OAs
vWFG1WINe+3q6MrWORxEeu/VQafQWR0K2eH/A5qclg2KYSsHB1zXdiNQmRF2+eR8
JArJHEAiCt/cZDOUd2TxbR2AeirUHRqAykaPjn+fEdEU/TVincKMLtQjX8W1SB0R
qOXwAnr21CP7YOp2CXwatnGhkySIEHIIxBQSZbctk7ogr3+OJaoH1fc+zxDhd6qw
fMtiTcaSj0R7uC2DrebKCuIKG7dmugFWfVFaEVhUKwIOgYvukR6dIhHHa24sjCCU
jVVR2cyKUOfC/nClRo63PiBzfzXSLG5RZN1U0y7Tf7m9Okf+KvfP3cMEVM77+6In
gKI3A3AOu6Nki1lfHbNSObHqfRpHVvXMY1j1U/l7/GC14LEqOLlXOwPt4/nS+geO
79C46v7NRv84K/nqF+xXwPi/XzxE20zqcL9jFrASGabSDWZCdmG2nuYEl8m9Vjzh
EGle43eBYi22v5GdOwR1l9VjPTAtAwKH2t9xreOSwbNbSh/272u8jPopym8HgBh4
4lVel+22yQD+2AIi0GkOvmLEIexBfdxtkZjOTSK69844wnJTtfZwRq28766iaTYp
kAGTeVkHTkuTU8CPuggga4TTi3guZVzGCFfCbyG33xwPpHqSIVC85lEYnCq52/MI
EX7IX5Q07Vop47eOfX7jVSLoCrVsOrCy8xbaCY6+lVMy2VJpGiTJ6XhgRN/WD6Qs
/EBDnN7uhgL47byUQDviVjF3ZHcPowXDmrdR2/sG8NSypHY1X9xaTLDqqjGiGk8r
IpMdACPQghDackd/XPDBLYcSGdREt9CE+7/dNaRde4s0o3yz1+Xnk732zXm9BleT
YEbmjE7p3fxrTWtd7XHIAOavWZm6+i2arIt+EkFvMcGpMnXEJUANMK1Z8yKMdIFp
/kk6eHZ9EykHh4QKeA/zrxKEZRtJxyEsaWEbHxLYIw7Mq0PJ17gIPyBuz1QizETa
GHHHwqFZ/6LtoQKaqHhbRzlD8PL/MA9P/oncHws0+pWJnOvRnYH050T1h6MhPfZL
z4kOaMKSqffjb2ZerEieVktiWD6QGcoJr9+EPjzXuDM/nrEy3ywND0PcciJExAhT
n/mu49ATpleRvpJauhk2MYI/K0uZZyZrb9Ux9CcQN3RBOD3nIhUxG58P2keppi3Y
M0gjoH1wKOgqbg5hB9box9Vq6+M0QkrMKA8PrwyHBUebRvypZDx9WxxrHw39G6ng
8TZO+HIj4Fk42KeOfW3QmTf84BjskqPGhUipmOWXEB56XB9UNGszPiR7/moxQjlb
U5jYCYIBV35D/WMnqZv5WlLSg6uKfOqeX2ElYU2FD3kYBMcgGsZXGwC2JVGJd7Pn
4mhlHpW7ns1xoiSBhaF3CsbFYDnBL7y9b+nnGawaebXCCBuYTVSXETNuQNEHW8Os
yhZm+cV1LTl9BnR384tdHzwDWn0PBtpi9ilU++S3EKM=
`protect END_PROTECTED
