`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Wj/+Sw13qZThf/NO1v0VWzVtbxdlsDq83O87aL7b9sdzBPm1l94CgC9emH7tUGr
Yw8xzPK4D0SafKbmD8OMPhDimmn/xSeE89LS+OoPFFTSxij6r16CqT1JB2HHatA6
4rPkMjqKSztL9zE9kLv7luSY0Xvt/aAypbNQQFyemUX5KIYDqi2QY4YYOyvRQbMR
us0S1/SpHFB35WS+5Zyi/vsTSN3TO7O//VMzA5RQhZWN03hCxVCXX5jg0++pUuJG
7sXc+c1BYh5EDnwmVhMDlTbBXXYYgegAG93CQRitTWPDRSdCTGMKadkeiWv1UjQ7
VqgbSRF7xIsOg2N8SCEXMsiF8ui9MOSuCql+DGWUytP3kl/thIaEfKOMgDZJNhXk
x06iI3LfNSq8pBEV2AcvzGCtyLKvamaQJdEw2pN+i+2Ox/1HAVpazRieno4myONr
yZcAZcjBZNneOCOxvV+8JQiDyBa1sN5vwgNpULDmuEozcDJUTF4WUCl7zpzTdr9e
u6ZaxMvXolL5x5GXKldN/FykUiPoptkXraUU+VAbIM1mnt4F/uDWSNirkdr8vbhd
bVxgypZFP6HCnyFx3GHLe2hLbM52pU0uqoog0gm0SmQcUfZqb9RMc2fRDTI43xt5
rYaXURRD5wAyaCa3t+3T2Bj/YftYqWjeCgedqmFFrwK8tBh/g3GhFuNmMU2MT80q
octsqqwlvED+/K4XU7so6c/7ZZW5mzGFTkSCtbTsYffNREcNUGjumobd9FfYbKAG
R0AVBjBbHR5DjBCRmzjFZ5JnvOzyIVcUTxrH6KkHOi5u4/GNc1fVHLiU2r2gVlL5
Lc7EQ76hs8D2GIFD3NuEitpblTYouL5mUfYiztTR0JJxYHHkypohwY73eGe/9prf
og5hg1ui/lByT4iHMD/9XS8F4TkUw9yDzIYXcKq36zy9M+QskZ6W+vS9Svd+IqbG
2FhMJ5CszbXfWqB0SbUQoLvZsmIN32VRZBbRu/29ujJ0lBIhNW3CHnzgVRMEwpP4
A5WgcBv9a5FhOSbt3/8KbkzneE4czspU14YCaG3JG14Cld90ycWm5HNLnaf9msqO
r3zQPuvqdGWS6pyDwu03gaM9drk1mncIpRy+aw6uMTOzdFwfyjoNQV6HlpiMpbmN
cJHkJGaWlyNOiXgmu3e+jk+QawaV+Y5c5/FWsOL0UNEN+kJVeTIu+duAZqCg+BHI
v9DHHlsaD4N+SZhHyQF4BkYv4IavHeAS6/QxofkTHjSGXsBf5gEbHpK2NR92bItT
BmxDL/c9gY/smBmkBlANVyaAPYXs1m7ZXEFWHUIf+fR66QtXciuNqd3O61KT9796
PWoZGM6DGfXYsuCdERQBrYrjiEA0q10CBUWce8gJh04tOk0hAaC6MZn0rCCeAijE
MY2bCVHsmML/tPsgpSETKWNEBffMnOZYUODJfKcHUs6VH8+WmatYgp6TQCGh8TIF
JsTgwi2YSLmyyClj322IXMHNxAfV7qy9zTOBKPJkGjNgcVyUl7fwyjLV6u663Zyh
fp6qX9J1eS1yr97Da7Hvk8kjKSm7YAEGhDRPNX4RihN1nxBIzfEBIg4G8sVNvN1Y
VVGUJ38zaJvnSU1OiqefZPLaFFe1aA7/bbvycleNfHH914vcUkbgSMHYCptmFaVD
7/Caumn0TbhBFT5VNbhkzQbwJp3qlD/+3KLIIckAlZtFyoPHFMjTAf0A7/iRXIVU
DwVqqSsBbrQcrqS0aTKd4wyDC1CAC38nQvH4ddsWDKsYSrzlUtlfzZKSF96kgpgR
vM3Rqytx+Ahiznf/FdciRRT/xuC6LJUvAmH7RR0Tfe+PDc706aryR/Xss9N6ZddL
pi86zQubkcz2y8H1RD7FQa1yH6YK1fTfhQiPsX4xORgUzA9P5xDhQMP1OihyVafz
eeQZbx22dK/5knq73V/STn28irE+2PP7aENNbRTHdgXGp/Mfb9dJvgFirbR9SOYq
eDzIyZDWeq0+4j/TvcIqIL52pdtHzK/xu0TH4t252XvOvQPZc6lFARgh3j7JAm59
sg8lPofI1MqMMPFrAFdVQotcNBh+tEozK6nDzOzwSmj3sbW0Sr7vNgHL2pOdSltx
fYvYXYKQafrOqFSyOzpvuF8mcestPoqaR12R4msfd6TKGcA+IqYfqNteE0bb+okT
w4a/+Sjh8eb30syMhLley4LJEMXgrN3DjDhei5AIiRHGGG8wK43rVcrRSKPqnjhQ
fnq6WOGv5qOEBdiCFrAXHqtdEn8zfHjRc4BtyabDEQq1bbAYYmnXhtH4MGadeiqI
91nzK2bLLif9ySoYFauP99s6ly8eYHZF5eGQA/nnJiFJIRZ1MYU3IPXXMPLgUdp7
5l+8AxCY1pz4+qDdA+bmYw0ZNzgl5+WkOChKavn9qRM8b5Da0eKAIOFlq4QkyGgd
vLh8/wOm8ozpUeWjlHwQALui7IMYV1Krvfa0UE/NGxfOckoBJr0yw9Q7MqMg9VAo
SR6X4Ga8ewqv8jrhwSzZCaNuPNhnPUgNYts5yyn1wOsmiGTq1bVrloevvHl5F+H4
LFU79dWQj4GhVJrLzaYodNg1GD61dHxraKq+G01O2JeiVLyftKblF7VuT4IYKOts
8a/OzZ/VsA96rAL/Molm0ntFg4ZfH9tLwYqb8NDWHsIgIV4QfrJShLQK3Tw5yVIu
RgchEellCHkUXTxDFJQJMChVMFHZ7SVXmwkyAFDltrhusgeL3PnXMyHjwo4Z2Ipl
`protect END_PROTECTED
