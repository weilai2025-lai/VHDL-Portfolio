`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNKVR6qOVOWGRJ1qie+894iAxLOiNNn6j6t/fCbln1vYY2+UfzfBhXZYsvJ2uwIo
GJ53ejVao80enWrkM98Cmb2Di26xiopAuQezu9FZQVtQ+3y3VN6kG/TCrmBEQD8z
2GTKduqotn4KvVM0SUoWNWgoGS0h0KTwC1jj0agKy/MC+MhfIxpxVUivXuuZJpib
s8OrR2+OfAyy0zg3MxcKLh2Gb+CE92SKt6RjDeiQK6mG9ylscOjsFHluCEWbjfgR
/QQ0g8t93dA/aRAkiIiijnpeHu9bBZBKfjnyqnsIik8g/H9orCxbSUyDvvLU4QsT
gquRxONK130vwUGdvotIF//1wvyB15kIKYjSt5VUXToJdC1ihrkamw1gaXX54Oyq
IFVMOoTQbGxGUvsxt+r7qs0EuMvp3FpdmLjhAWvVzfnAhBSMpT8+E4pNNrUnMgYZ
WTaudSYplZ7MLPCRdZxojPpZXa+UgJwHZY9ODJqg+tpVNxXBC7uUjqAuKnshIbJ3
iUhoW/c82w8wxTMdRXbP/0xSghONW227dmTtvXSuSsFlMmYvPuGECvPcuZm1N7YE
9sA0zRKjzr1Ja2NkbPzp0VChiJl0/wShfytaaTSJwgpoq4ieE5t4hGQYbOWPgeLD
apjdxvLgSeHeMhCHXHSUagZWckYsHvrFbBJa88GpWiTH8XrvsnsWRtGXqpKJrQif
4Puao34kYYH46LoLyIM381OW1cnUa7hrivSLMiBCUYoeW/89bSLMbnTSFlb9SDMM
vSV/9UZ9ZaxzNYswTGffQluMGlXOQN9gIA87nOKG8nlrQNax8KUnhHZB7X29APvg
X0BRwCDP7TDyeqLP4btqbexsUVjkgZS7+nqJPpBCP9ESEwaPHWXT8XBFMoI1OPDk
vYq+AX5PSQ112RZY1xQOVQwRBlp1F/TkYq6EnZaemdOKolBaf2saAq0qEG9Jfcmc
WnNyVDbCsuZeNlsh33fozdDtfsYQAacaGyzQWlQ5txaA6JFui3xsRjUL30AWqAj6
myovYeCCUBfgsTXKO9k0OFuZDSWMA9Sl+D14m1Jm39YkXOnZ8c1fMbgTZ01XeTDE
nLkFgY+9/2dceyj1P9vAvjoWF8q1AuznWNkSNE9nurrqAse6BT4YpVm7GmDZbJM7
QilNC9NlXcE4GDnxukMxi3GXCpiu7fEt+hL56apVgWo8i0SpHRUnq5at1v0NSSA+
HVbHr4M1YbpQgRit2a8jq2P1o+CIxyh9upwNgrCsG3HwQ7nv+ynQTuNGO5WcbO3i
ynTsgOv8+QH8E7sVEdNTcwragNOZ9nBRc2FKz/f+X4PKe5lpYwV/gs1oYyIlwxXI
/Mee/O/GlGYHs6p3dklKNRT3Wju6+WGsw/kSt3Jc7GooEQsJsBR+q5AeQgKg2Roe
Mt4IQE0Ef4kFBJIsps7Wu72LxAG5wT23u7p83Fh2TovQpJv0MCplvwseDi+Bva11
MGqrdr3rHeUH0cJ/jFHrL1jqYilUv7sWqGf2fq4sesIbtuDXxg1yWrJSEIF5n9NF
sTkL3uK3BddHctVETCIJ9vM3DUj3uDwa36h+EWU9iBdvzSfQtn3NiuVR/Ms3tyLa
lw977YVJuErkyCOZOpqx5k0Hg281m3ObRoKkZ5gTKz7i5ne2OiqUC3vxAQGOh6S6
F4XDoBhZI0afWm/QyRuDQ7gqcmHh3x7jtHqjaVIYI/BAXM27UYWUn3WadW1lwpFV
3aNYsI6kKTtcVQOvlZLHGDczz7+PhAn9EBNscYDTf/sUG1SD295yHEgPwIacv5l4
zp7R095LZ/eMB6Bi9QSt1rqngTNuldwpkMV7KgGC1bqo4MQ2zO11cGsai5hyYMR1
I1B4zT8ZXnfzZME0FF6cRKxToU9JrortUjoIh7/VGmu+wxXsiPMOSiKbhJzIZD6W
sSW+Mvic3uWo0oItb5vB7F4lPFu8UsYIMdCu+AnIvUff/HRM3S/yBkTl+AnRLPNl
2FiWOKsFsm15mXI4LLKHCHpinoKxeMGV4rJYIYObtoSdh9t2Nq8kI8uWH2NM2vti
lvX1bCeP+gpOiyuyJir7wgHcpx29+nvEy7VHwFwa4SxVSsg+OKBv+IKmklAYWSnc
AMr9l40AmvgX6GUh+MfRRM455RhAIkIzO+0gkiaIYAB0WGgnsLKeKt1aItYp65U8
LCs/uCDX5xT7nChSo4eCQXLmcRkzPNZAXjQzgsuqEwcac78cg5wp+V5ThrCiWfPx
11ICjiY9kABbJm2QOzn/R8fa93NDkoJ2mfPKUJ3oB6CyZgPgv87wOGTOtfSjuPHD
P9iLS2Z4bIudCV8lvxEs2epVy2rpZR3VpsFGNQvVBKkiaHNG0JyytnAgXWGfqbLu
l0SXwQf5metMnta7yLHwbiUdmj89eVIYwIlu6+aXUDDcg3W9S28XqwYTJ6/hbV3r
HeQGL9x0m0QPZOwegf2VrzfXyLvISRSq6uzYBv/vex8vpjsMit4E0z91jOjkNk2s
dXv+Gxq9OK97U5AU1JSzYG9eXthxAiQAMUOZSg3O+s5h8dwHFpII3hjhSkMgs69l
wztVEv9s7RIhcBhvtyc9QYvVT0F9z6jWhI8hZz54UdK2z3Hc3EowPisuu7+YBwEd
Hnu6x8/cIQ6IjeSKtNxoj4vaZO1fRK0m9A4LfkSe6RMgCWcft5oFxxy7Yjjwy+IP
alI33+xm7KxGhn1fSUyJjlB9UVAOT6Jr30rBRaVdLWowrkkgYEcmJ1nBYOJSYSVm
zyVTqCc9lyiEEpClQzClZnI3InEetNF2ISl1EjDJzYX45hVbWrFudMORajHeScyN
5FYd3VgnQrcC00Jlj/tPx/9QKBAz8Dgs4QaGtfiPkQq2LwaIVk2WddKW0+3QpQxC
xEA1CYEkBWtVKd/mVSbBc9nAebihS3oWBODUDTGI8mCHcrEMHVm3DovsyFOPtpcc
zcpIbm5KvXFLSvxbyiNuVAspoCDLE+y3vY1t3xftpHmoyytyVRDdjV0gmhjRargq
qcLFE3v/X6Sy+z3KYYCpN26dqv/kVknrK0sDGtwKASizIDXjcRhA+R171vW8qtXd
IKUWK+UEnd91m1pkERKl196/rtj+T3KRMWcsKNP2LngOVD7xCgIqhpfzQ1S+DOl/
3vRUfBU3bOf+Ee8/rOoUGTKg+uImjWE0aqbHD6QNKOmHvv/W3dP1NW8MPDktVHaB
s5lmDBUVnDHX4NOp4vmwi9XDG8pJhcpWA5JOfEV7dBnHOOh78mXSzsXZi6iXkuA6
0mDyIYwQioaoe8J3BEYbQfNrRSD2wuA/Pfnx6vZ9PfvBdscukLutM5PYtK8ZHHGM
N2x2NBBTCPKgeGN87teSfEO5rjtVfoIBiWzAyeX2QpZ1O7AdveO4P/Mg+iMqbLKx
G5t0g681GLNiVFQN8nGXlEBVGl7ljolGIcoOcHyjAZN5nOf+EUhR3Y/OnLZvXQIE
QAIprk8xhmqiMR/sFdLRaUOXCPChDltOx66mMUe6yKt0XSW5720W5iMSPCOLL12s
6KWNdINagYSCE096KYKhk7ssf6LCQ0p7ESd3UD5vcuIOLs1hbG8ytHp8Nwdpgjl7
9Q4HmFNeLpDhLQXxsgIGcYQbi3IWMq8UK/xpjyCW+M8NWjOlPX9bCDMq6nbryCyZ
eV6Xylr2E+jQ76Zt/8Vu4Gk5bn6v83k+fVe8B9r9/Odl+fNTXk8YgwBXiPSMc9oU
0WJP4Odx2tC61hRmJhwIph8O3TTJK0Ss6x5V1aFO6JsgO3wYCkf9RcX0V+G3+BRS
zhoc0zsykh42nIReInBJOMNtjsLAhWEcP97dhf7Hd+z2XkprkLW1gStO9+rGLfan
1efVDqqu8bRfEhDWmp5a+ZwBx2xY1WUCQcwZOw7J1ZNfYi7YQAjgVFK2ulDTa63l
9MrLqaN5U3docxmw7WzdcJk3kUNE1zhWKAEvrW87QzDAkC6hX7+lwO8aB9I++Dw2
S5te/mc39I/vH9aVXVFRQw/SDET0FnXbg0hdh8PjGkQvQi2LV6WyZ60dHJKqlQcJ
7nnDI7Q+3BHiF6OnXaPuJWKBWTPkj4L9VmFp1TcHKkKDKy6P+yBRBATWTLneycmD
LnWDkrEX8o17Zbdk26OWMeRiI/ga1PROpSx2crc1mPpcF59h+LjPBWJVX2V8QFsd
HPPZctHmbX2L8my7lVq/iK6phiTELZGyDrOLXcosyiw/7jR3bN+gbZVvAcNSsZJO
bB42sFegPGWsXpj7kU/taWccZ1007vSKeCTs8SFWBsaq/EMAUw3hr4LK7hlwlImn
8n107Ofk7sLyAX1CYxWbD4LlRbMHE1BgdNMzf34fhycaALqrn+5OY2Z3brx9Y9gT
8GOmacwr1AfChnlMgMYkvUEZWR7KB3HgOuQZAmvHhOq1UTr3Fno4rOKpy7GIPOfL
A7TrLdKpq+q1QV6N6NEVGTHHzVgCw+TY1dJZF8FUw3QQ35odNBxZg0E+q9Sqdmww
O5+UnfNk8zIrTaDH0ZF3UvSzQ4YYBasTg/YfoLdJziQuPqvJTbru7xlavfbsTxVQ
iAy3ehMdzZv+qxC5ipBXdzkgpd4XfOB0cLH03qt237v4YPby95v9uNAIAW0i15i3
Xqy4GefX/j1+06wvWPxyeZ0yBJxa0k0LjLjGnUrrOUgumv29Ut4sJ90axgBg2P6O
cJcqUU8S74dGd8V6b0LWtGFE/q3zFAxF2pdnH7w7vjiMAm5KjrNaEEG7A9f+hoUm
gXilMdmWD7amKgD4MLhFHePKRXx3sIyAloauDoJzLvatL6jkYvAG0FoauZ29W1+S
r0478LS99TU6JYIQvhAYedchTRfihuQpI596pNU421QulCZ4sdzZLbzy49UosK8d
RQun3svcidyR5LW/XNJmEP8XvGpgsHFg128deycA6hbYytres1dXtNbwiyNXOOP9
EYGYu/r0Pu6hINPYQZZAeEXkqiO89rWMY5aSjwIX06sYdXWn5YCnRscLCxbkZtlr
5FmmVemgPuq1kzejRTzLeGkqJ8kp12SLb7MkCXQecmT2oKZHFQT6RwWqpkFxQN4D
1oOIg6KVQmkcp7in2dYN/KflJs71Xw3IAxPNDeM/+qIdU3SfmieAt8MSLhz6/Uks
Eeuhwsx1ObIMZU6RgpYk2DWs54uDbwljDjN8Mn5ZwZ5icTAHyVmpUWOGaw0S+EcU
byaioqDJoy/2WoKF3s8NP9gg6J06XuZIVmiOUE/Q0Q1E6/MdJ0+r3E2r/BJrO9G2
HLp/nG7nGLSDLJHafGLcAJQIhoPeDcu14ELYd/lEoiA80Za1H1cbM+SePW8tCJ8d
tCVj3MtWTH4dzWfd2VdQxwqj1JTA2Jan1ZI4O/Euy0eWuX8Ue53AMSbKp8cz4D1n
jFZFASwvjiYXBYAqr4ZzrRiUaR7yrdHg4c/K5NV0Kq/HyFUgUA9YkDMmsN0qetrV
a9n0JqRMGTGiE/UxjHBTMidARzVg6mXfStxM+jWjClb9JC+pwRizw88qiS7USYYm
NVgoQTVgp7+0z76oKONaeDicPZPk+vd4zDwLWQIL/GXY5Rpxl1mMxGKjkD1Ohz1W
XZSrE+xjBU74Az+G8XvH24RbdIUA3LTttswllnFQcLWCOy3vjIW77cCDrS0S+cne
el3mxLRk6RtDbVc0u812RVPsWLw4Ap21w5FDsHI5rDQQwja/f/wNbPbjMT691hOf
zaQdgmqFj4drBFIceZ/FLDTwEvld8OEzQrMiYE1jjM5yfvdf0e/M5nL23eQEK8Fk
aQ7W5Hb7t6v8O0AJFESZlC7IXP8s6pEOmh6WBVgnhQqCu8TW2InDqY3eLztyHiky
cELKqRnoYjnBwh/fdH4gkVfzch3O/rATsdJyuUtzVX9T52xtBI8TfW1DB0ALPa5/
U0/jfoAUljuxxyc76arLJ9wsPo8KmZwcxy7W1ScbYKnCCdPTxd3yJAQFKm5oEzkO
cW4ZGuJvS0b8L7bb9z0IK6GTC4mDK/jT954HeVX3sw8t2NI/Q4LWPwMsqTMRwEEx
gcK42weTmr/0mD4lfZPiJyyZavNx3VHbKE7oxwyMIoQIllOrFzDyNeM8XtTQ1I59
+pkJ6Zo+UjjXSFyv8IlwrqVc+K8Bmo2QAitTFXwyw9ZREXhPkUTZ6XRWsVnfDAaD
9WfWOCu4xJOGa737hs2a7qwC61sDTSLy9e+zJp7Y7ECFrU4s9GLsPKEKjWj2C5uG
5X+lrQfb8szWIrJ9aFOrJtPM3KN0w9oIPZx0NmwhGcJDGMGwKDQaAkRQdQOsh04A
B8rQEp+xNQxMs+3msDdJN+PLGUVD5zDymb8yUNNk/Ezxl49aCmbUwPkWCGAfPwc+
Q+ZC2lOxUsIng9OZ+BGRrxFVLU3g+3BG71zlRp+tBxN0BSP3J9mfyBbLj+scIHkn
1ThJgF4INrafyPMrWanJfdAPlkc+IoGjmiqxRaa6qnCa7xbAvI2ij1TFt/VDuWn9
u78inrF5qt2UBf/9/i2/W/6MqbzcVmd3phOcl3Fqpvx2GPcxFhER4KZUSSbAtBHN
nRMUjhc53OpCRDpFcaWSwNE0hWkiUyc5TCpb/F41xLOLBq/0Tr8S8Z6he3YwtUVn
ySFj/LudtkrMWWkUQK60F4n/YTyWYliI5hkvkJnkcrr0w4Oy5qCMAYFYeR455dud
Zp6yNySTihNvFDab/YLdKbsdrakT2EXHQtaVEv0GGckIx1lmdkMKYGZpnAawCB7K
MeUSIkRVGSuZ5U/P+i1zo1DHNFLKBOOuQECiFnBtt1wv9zk/pQ2mRVbMDs9E3waI
GiQrjbdc+ebwBV5hR4eKtPbTQuUviZlgxGXcVYQlXWfMS9weOFyEvL8i5biZEPHX
dqsTBCM+EIHPF6ntr3msotpoS10BzM0GgQsoQKN5N790btVsRciMRJ1bErUqAts/
khpdPl8OEHmg0vOae0md7m+bn8o5YVeC8p5AXCKj+WLTj/LnbV5XDUpvXRtc8bOb
2VbVldYd5sP5EUTMlWayuqYR9Nz/ywoJbpdJ5zC9ABXRDYkwBYAgo9bGTljuavgm
VH19kvGpMgMXGilObXiuMp4kbyMk2pOHI8we1kpk4Ez2oOXdiLeTo6GryAbW8lkV
OqNR5PLW+hyzSbS+zFXm4oIrwwz/T3Wr4PN4Sgb5VPL58U3idW6W//lbzPlGEMeo
WhCQlEVcIwUBw0IY5cLwNBtceC0ZyyOxK3IvfP7a7BPu5BsEopYeCNt43D7iAR7u
9im/tE93u5nx0ya7ZhqaL8XBGW8v4kFOBYcXLJQZeXYCOhBaEd/n8xgd3v+sxgCk
z+S+mR2LY1jgxrsoLBkMAi5lsg1aOrfeXyAw++cuPqWHoNAZpju0AsQvBcEb0Mov
+zZKyS6nCouXNBha36yhU+xRQadA2z3A/k7wUDJfn7Vc/1dfJMQC29kXFCypRmtJ
meDgTHuRZOPqg+jaOEqkKFnLUx37Eq8ewAtiR9EJN04SIydkt5A4PHRY/vQ6MY2Q
1icpTKRsMBedZv0R9fJ8OnudhD3Zr8vqWTSGNARuSnFZz3VMx0u9Kbjp+12O6rLv
x73dTV5N9q91/3FHPJfc1b9AoAhfpO47V/QLvWgvICAY1UAdN5SdUFjFLlbuK2nN
FAMuPFgfj5w3B5QN87fU+7lUeW+B18BxR7sUqJ7uN7heMhFQXYVX7SOnSRI/aVGa
naxExFTaabUU9Jck3zgdahE0z8hrPGN5oy5tgm6KNytv0IRa2SSoYWJ+fiS4T0Cv
TIZ+A+xQdf6PQ7aL7qlzf0npGUBl1BaQXfGsVw8kRV9Uj/QCNnbtXm4SNY0GGA/z
a3l6c2Q3ywAcLmTM9ytjR8dqxz+aNgvvCY/o5BfGwiCRYqSdc/1VED4CPObm6lAP
JEcrap0+SGVzdLYCMT8iVOcXG65QF7YWurfw1usfTZsKEdv2QffOOdiFaYNEhLZm
1yUbHR2y57BJS+TrHA6sDqmN1dHeDminwP/6N5ZetTmrZO9pxJ+YEP+BBzHZDY7N
D2YzLD8/MeiNyrpC9LHQh9DpfVgvHbuAysVjPyuEurauOlZ9nnrbxCHWq2p6moBa
qLUPh0fWcZs+PBLzgxpp1BuN9LGvzuiW7SW1M8M4sVxGiRto1S1kPXEPjMcjzjTG
+H+p+WvkvWY+E842wN+XDfnMfR2QOw3ULqd0n03/E3RKLjkwXdUN0bCkeDHp6lnn
uc1st8pkuHVdoyQx2XxIDWB48Mr9Tfnr9ZLc7T+WXiMzVwuuFqZVpL9MjpyRFJ3Z
ZQ8GqrjpDiggofpfJfIdte/DY/rwAzjNycN1FBmwRNt1sFfuIunxwBcJMjslgVSk
OuWneGEr2GrLZUXIc4YAtk2r0RUqoBGKYZ9Obv1gWRp1120MLUHrhSDNxhSFOUtM
FgXKzo7rJWBZpzSXCrzvggFtCFZFNzAzNcp//Q+a/9u7JGyyp0HZgCF63qxLobAv
60CCm7JaU9K1jEVxHmOPLq6FMKRZ1rCrzLrpJiTjfdf3Bk8Sw4sbeEQOIDn4/D8+
dImaCwcJ1QSUaMTvOM4fXeHZ+s9rSljsc4hlsawbl8HoMXwtHdNzMCUmUSbnVkRK
7+6TR7lg5QjeysM3+OPGUgadQbSfalRNwMfvYa00Lia0n9x9jC9iVUcsZT5Lnj5w
6WuC2kU3XTjPSZfDQnLbdSVyLN3ePwk421vtWEvDMy4hKiOJalUoPamrbBmQ0hIY
k8J3Bu14rfVxrP+ExtaX1pWfZNALSVBDrLAZhbrEiF4Pt/htL+Ud9a7YRPT+mNEH
RZOQvVVsURwE5AUnpWOHSYCgBxj0qV9kPB60pTjOQmHkFxqsHJLXFGVO7L1XWOE4
O41D/uXjWnyclxLT49WGtQ0sQur/lMHVEO4iEDiBkIv444GNjcDvSpmrmXL0HiAK
oQ2Zj8jzYocdvvUyYG5V5DeWC8PZLXDTy1sQI4MiUu1sFwANqKa44ovBkVwIYWP7
GSxYYpQ5+erk8vEhLAvuTBHOLFFsg9oF6REDMmPRj2rSRhMyZT+fzoSypdggTgfr
QDYhib1gF2DqOxoFAoSFORvJz2JFlJ4LYsQiwfyCmIg0/QQ1JMK6nlJOH4bzHSLe
6KrOdV/Td45yZgmU9DY/P9eednfcKIx90yH+C/l8JR1ZeqF8w2L9kW+wZuG7oPIp
ueVchpS3lrkeAZZnhLqvvdL8a+C7iJmCfITRATM0748RO1kC0e8ykRMVdTWRImFl
sjRhhcloL3kN8CEbc1swAH653BjtQVUYLrmMYIir6cf7E0DE1jnEmR7e3FbAMDnO
W4UxrxHsby2Ye0gsBUBNJkp0J3q+znlkcB9Hv3S1Rnj88qXi4CrGmcxHlyMJn6Br
K0u9ePaMm8ycXRoEDwjLrQHzQXxSFcQiP6AqPT9oIjB8TGNSwQMeYf/gxlMBC7k8
j5pLgrwVnhMaXHrr/qVE/XkrVALK2lUSxM/dh7YkeRNJHNFTe0GLaqM4qJA0uzk2
B9y3BYbubd4MQs//TwGGBvStUz7aA6VWW86TQ1En3HYHLEgL5Q4Gv/qN2Fc5kf+y
05AIsq+URNztKhR+W2Mazue2zReo61c2+KfxH740MLrA/FAPb/4r8xL4zA5JepV9
MqNppMXH2QVFRnr0MVpzMM9k6Y13daOBDJwUi7cgByP8u5M31uqIqicIx7DUFRuj
XhM+spU7B6i7+iZ/YM81JZJs+LIP8RwAAtYsFrv7J9ie5Bw935r0V2+E246X8Cxe
nsCxWjOLOtDXeHKOK0olt25DBs62g48RGKmq1f31526VDnmVZDWwlNoQeNXRe+Eg
IcR/r+K63U/1XfpqyxqMLiU0oJn/JOfd4cVVvCI0bCu9JzgaYyJGI9JZ7gLUTr8k
wbrpp1h6FQ5T7VMwElJ4wQVbDYIW/F1VUaMvGzumYV9Q82eJ7k4/7BOO1CL/1l7A
vI3xES/vSY2f1Bkm6me+OuzLzkbK4ZK1L7sYrfcBi8FWkBr1vqibqyBMUcfUpmQq
tTHTvRqQO35DtsZ8b+j+pmxZCxIoXEfNWqtm7gbvm7VIwTWAhskPkMbhK0btmZkn
iTX1zTnVUhhnXdbY4Tg3cO+uSdmS8cpXdOYwsseglVTU923QkIu/NHdf/ngoDeGF
zA+VLaezvwEezmAZpu97YwOYXJFBFvsQDkTQJAFlVucxMfCOqU8d+pK5HFcvMdbx
Q4ueV+O6+XkEKD3PHJ6LiCJKADLoDL7g+I942O/xEubjemxjfvGX5qQRoDpEUTMf
bBP+/VDVuiS30pa9oNBgwa9SHvzwoUiIESS7dOwlZDcZLPZe0LGsji3CMR2EzmYL
1s1bV0HxbEG5Z3A2cB77IEHDqikVQbeu0ywOItfnPaD7LRCW7wJp1nHxUjxKQxz9
H64RAdR5CSGFprT8gXZn+AHk3Rt/BoB2Dv1IUE1WKrOjd/+7pqwz2v6Lo18NjjU1
5VE3y8CY+GlPc0NxX8nvw7j2ol4+BS9HoYKKMU2TICHBeZsWxvR5LPmqwDYR4iqT
PidL1a+ocIcLOGbKEFscp3MFBRouOp52Cj7Y/Kdlqz/QjbHCLOGCrxpEyvUDYThn
oBZOvHWl0uN+w2WKpygAW5TU5ObBWkutLCuepSC12zJtkU0o3k2ODc04EF6dNfW+
t+s0aNoBVgiqjL4iGjvppsnrQjK5XlsZ76K77h8ojBz/UZycVFPvoxRls2B1Ecef
B3xG4ocTZBP+8daOGeKfPST/+3SzQisvcDoXSE6tSr3APuPAH2Quf5iiT5/1WWpe
FWJKhy5mTMxCwr99stmFjISnS41rH4EmGUJpx+wcDDHvGe3uQ3zN3nFVawmuWEqA
aCyO8hcytMgub8qeghSYJLiJgYkry76CKNqE1BT+X5IncXv1g0C6dFETehPXA5H2
Gtz96NkF3NrB3j2Wpa+cySO1Z+n9a+ltgtbJrdMa84JPiQ9zfTS+WUpIeEpvaFND
69KGNGiP+H4mZXiV1SQBRTV3XIaytacp5BZAZ7uEcZnUEZVeS6b9vYMw4mEm7QnG
B/wH6mYGsdIPN6bY6HJByEe7a0fZj1/G0o1AkTAcbpYWcWFJD08/z5PTcRA+xfA6
iFFL73TghcpaAbwkHrVAdYnImC2kOvpVI3lyUEHse9rJUx24h7jzxYz/Yw3nOxXh
KddICLdKGPMmiPUv02qIO+i//ENvGbA2+ryFYV3SOcVuLbm5UMwhQXCyqALk0BjK
hUg0LxUBjCGCE589EuDlIHfBXROQED5MFhAdFab2/Y5HprmZpbyyLEHRVmzxfWd6
IgV4Ob7AQ2LhfPqOZYFiD1mdgTl6m6GbL4URBy5p4OWU0A8JZKno6bD6Vu8XzZz8
JL33Dp7R/ojtWsuoswfVYHS2JPtBpJCKmF/4mgQVzKsmU+oDfiNOf5cvL2mP9R0l
ktzazmhy012KzLhB3KiHK2g2pJVhSUJtL/iN8Y97wKX36nHOgNO1unBG4iKocn1a
HUVBNlvivLZWtz63vYALmCRsX0VGkG9WvtqvxpZfOEm4v3RUorjY1ORebGO66YP7
H2BF2/OyUfuhgt3Xhd2K0/Vm9zt2GkNqT8VXc1Sd+1LcWtxRxGhxQIfVu1RS8OQm
kNmodbo2jaH3G4/KX4Uiws5XzF7MXL9QEBzqzpkZOKHLdeeFUMyrShqpx/ERhDHp
6ORFzZfLEtTGAsI1TrwHlmRQa9HwPPalj84BUF1CTfL6LT/GJ/0TNk8TPqS5I9rY
olVHMy8ScJsy0GrxUz5YBuFbLuZLkzhMSjRWNK9kYkbKpxofjzw560PtIYbJIYVj
8dkX5CvVkrw3yODcIZbiiRr8uY+9xVbTlyXNY7VNMWkv7huVU/gO0LgTfofe6snV
vKGr9H1pV7oTglt128huVIiVXuMjUJYRdO9hhgrsx0kOYsys4FdQOHfxgzIK8XhH
VPbGUJIFiTXAeyZBOOqu6vqWQ/h288IeavKbNWIftAzGaZnX4HL649EN+7/Pqm5W
d816PyC75//m0oM74L8onMllkD/svYGkiNBZphnjUSDmi72wJk4wLNBGG5ic5z6O
1jKm+kKoy9rfX4XllcnYdrBr5VSR2G05WW/f1RMkUgbmUZGMv4dntA79yTmqBL6E
z9Q3oDDb60aUgzP9BM4bsiBzKkTIgJQR3zjXAdrM6WBpEAz8t692J1J23JQFyt0A
duiJ/ZuMNPtGjxybdOI1avoCeBgcpd1hKZcMYWNKX4cBNZlVeLdyyRNICrF5GeB0
IVwE0Q9/04PheGjUI0ddPIR8KWUnLa3DRnwesPubx8pDnDiN3fVDViEmtlZalT10
da50TKgTVjtJDmbvGbdg0ANm0tXtHl219SsB6e95kqQVA/GcJzlHYnFQLY5JVmkc
bGuiYX+X2ZVgBMh6Spcj0FwecGjUSNMM13TimfjOz/IYDZS/O97Cp8Y/hLD7R/Hx
cHZIfMPFnMsWJ6OeTJQtY7jwwfzynfuV4D1enSzC3T56P9YE/tmBAD+OrHxhA9ut
PAhCHpf2n4gfSNgy8f9w5F4H87HwsB9H59K3njm7dLI9OMEVBTZjhW/VVfkCvvul
g+ICkk73GNie5lrmX+go0z5kCVeq0gwWVshTT/v9MqJhVoqewN+l0La8KpT5EYOB
YPFAmCR7vkJEgO8EaN793ATOjbHzQvBQIlKUofpLbL3QHuits9Hxkmh/9BdnP9u3
vNVZHIT9ubIica3h3/KOFUX6jUL69zW48cHO/vZI936BO3DifU9H9U6n2S1vUp/6
Rf3ETIkribT8BFbMyh/49evVqx3CtMK5OfcwPyEhIG9fo15GOWnn4RB7Y1aZw8WN
xgsjlUNZsRHZplJM++6WZ0aQ7B4gTFALpFbFbSGekCHlkmv141h5R7QdkMrS3Fk+
tSWtoG8fJjzx/c7LzbPj8810yaENfKgeKoeKfIlxVuWHxUPQ33YZI1KqiMq0zUWr
ecjEYblPqx5vusIoWE5Ht7yib2duAzo0dxxqaQgE4YgNm3nVOck1OBEdbtERfKFp
V1zUJpvDlyzq0e93SE+3c+Zz/qIcxVWhV6W1bGIUG82+IX7cOq9nKLqAuhF5fLat
GmI9HFmYqIdj0ETlnEfmJQbgIVa5tpxk3Xky5cAj3pXe2IJkRT78boU+pxTQ5CG0
kRKcMjlhVX4cRWConiLtpC//AwNqdBGVXUjvtVyjp6B5797YZYsYLP77qtiOyS1g
uoKhgJSlEMl5DoUOun21kfkUE4kMGjt+SH9ZI6Fk4co5YxSXOjWbrnn4n1BgsFL9
/fmpGk0BXGz6XUMurZbppuS08S+1QFXKVTiJ9Qm92N1Ts9YfEzYiaYb+rS6kNHlF
oF1Zb9mHAqmclzJgQi4GkMXYomjLsbc2SyhBXlzUiVnoU6leI9DPt+ssUYl1vzba
J61849vHVVxRbdl6YHk+YUEGKx/w3l5fWNG8sEAaY2VlT0VsOjP9411Du4QVSG06
TEwaQgZj+30Lt6kRcS5YCnLxPZzAaYwaWQEixXR/yuDtw6Pmh6R+mt839SxmIYED
67Hu8p2Cev1/3YhPUg2cgYbiiVlW6uHBRjiO98dx/mup69wbYxgBHvIAJjHXxGU+
5n8OUtShoSxkv4N2E+JgtN4mHgDq5Qo2L7x8iIIuyxWNCwhogYRjZ1bfJrg7oc/m
Ifcdwl0lIYCMqzkgo35c69SPVGj+8oesiYMnq5RJfcLTHkiRNv0J9ew9SOZJYl+I
PcWeQl6v7CBFCGrY7BGdxdLEBWaSCvdM4oCut1KMW47KSsvJOXd6wS15qZhP6Eg9
g35X4tTlqqbUAb28XT2CuEeg+DUVXpG4pHnkdrUEVYImZk7joNJyOYjZC47uaWPR
ybn/6l72oeHVnEJG9+/1t19NOkTbUQzTlREVWm3tYcZAIuGb5jsOCCEVd94uCElS
gAZlDonYL1f7kv/gAUuIIaRI5TS0qRGFvvpe1DXYwhWMDkS1BIXz0cBjm7RwBqzW
ICquJeu1ip2ThviK7XPVr62M8K5NawhQRsDxAvKaxBGi0JpxpAdFENMWSSKA4d+z
DlgAyrZuVDfNabD1detNs+mGDj2We8kVywiE561+g2P0HZoKpv2WAwnIuyxZwURq
BrR3I39aBYPusbJ6k9vPuV3/i0OD9xasnCGZvhVj6JsviFERoIilzQ4/lIiRNINd
MvrTX57u7srQupKO3dNOPBpvmCT2KwHzHFO7hz6EPXnr4XMRZbGUN0M7ssfmGUTM
wRmylTH/QUsZkSiPFbBMAnGFoh34Zg4SxehcyVdTkXoBMy7x506/ny6px2lqgkab
T7GK1UZ7Wp1eS+EuLxkIyedW1Fug1sC+V8IwqWIjZcUnB7UWktjIDWeQNJqHZu9O
ApD3uhW/wLEE7E02ID0PY18qLNkl4uvP6zIIjv772YSp4TlXMJWe0bL4Ps9tLyPd
jb+LeeVym7AmWPkV/wb40gy8CMX+18slOHCXxMqu0EJknzJ61NMc8He0Bdaf+xjj
3a39T30EYKaN0/lR42inxZNF8t4DP0TNX1pzy8jhCQHftne1nTVK3jEpqE9d/fuP
D2ux4ik9Nf6nybE4pfNOyrR4W7q6zi80jZlYEn1q7PFsl8oWpotdlpmVZfBGAG6z
H8hDlj6071RiuLjMWH/5872ie6FcT/N0EA/sXEXFB5HCEYl5VitUn6ap6sJHCeGT
oRae65bz6gaSZKSLwJmEk+ei8TzEGIJvH/DYHXAuPybfqHck5R7/wo1My4TVjB5K
MnA/sIOdpiZzr+t2xcl5Thqu15iNKdIunZ5R69NE96HSj+EKVdNMNF04y3i8tIc7
QAHsTzUEwDh+PlCNy/tzv/70U+RavTyEfnna/LftAOjZ8zSH464rrlmBxzDE+J5A
JL0K+WcXXRzWBSvO55M86OMk392H+NxJiMLefZUiQahiAuHD8GXHLENsmXs3NjrW
3IJKran4kd9lZ92aOdGGIj1LdrFakg75vdWyopU8BLWDGBC666pMBh9h9quTFzFT
JAQza5gbzc2DzxJ0p1WYZxgbyskuuSpL1v4qCRW56d2j87v7O5M5wiXJyivel/XC
tMhob4/NI1tylmEqEKGXxWY97d+7AiHo3xSc8I7aBYjUK5ZTjvukz+ukb6zVV19V
vb/YmNXSgA0+F5wj6fIb2UNiNMDK0kGFpHirz5ypHZKwPNN2pmVWNsi78Ci1bt40
s1fhJXZxmndgVhX11QiT8+G7Uk00DbeQ1z/WnQttgFg0RJpqY+4pc6gYVEZZWQrO
jgKKx2z2HsgbUE0bZahujiCIGu7XkhrLMPLLqsFp3Gyjfk4l9++2/s/L8jpglC4A
pQzVKbufUmhVkbH8da/wViBKVzwvGiASqQHSvLYlFgM/+CLjX/XB5qzzypwtN1yW
ILD2xLMXt7YyLNpgMTw4Ye+yHUBuMppmfRAfqoss3fsrDWmfQVfFRC0jLKyiATkN
9PQUVNmFey7nPwXFItcu9ndhnQtBU3lEuB/b2UhFHYPXvo6q8CEDIV80CcIIVs+C
jw8lOdzz80fi5dVcnwdXi4dsSCkUfE3jIAzbSSa8cWr0mThvMHj2c72uzWKtz+gg
3i1K2ZDNzdd0i0WjiytkS8exGYSVq8wvQTm5amXa2GtWXeLIm4GjNaYpiNcT//LG
HjCZv3vcl6/99YRua+U+hK+Xze/Y+ou51MMmW1PwvjSvFckRPmnQhZmj2F7bvJAr
Ci4zzYB+bcMhq8X1mn30yh6PEYfaJDVkpPE+mdU5Hpad0emwJ8jrmAEglESJCMgf
vUlC84i1mxfjr+E7Buon90PcUcYPpvRTW7REdwzI/1PaFBX12w/f7dNRGC4UOtWN
WQVueAQxN+EhvsG8jcZbwZWwlryAjcPH3agOyG3wsQHeGsVshzMa6kK84uu2Wvcp
xgc+WZI0FVQPbZQcJNTWzEOxJWAouBscJGXENbJr/OM129juHGRftx0nrlBWdjRY
Zc2ADGBiJWVUOuhXBZjFZMRbAefqadrDU/WBaXwRxHGd3tnwU8hCg5wOljHOmp9R
qbc/2rLoVI0kaONFo/JNIuFUYHNqucWorB7uRH7z30VMH3Yxa5xthP0xwXOHZorc
MtQwwyQBjF5mEx8Fb9Yw1DeFMqXU2dCuMx43DXtX2b3TjOuYQiQDwZOlZzgTIqZA
kWCzVWjYw0WAUmdNdIMn3Buw1bPusgAVVF/yrcYp+T0DNvTtHbbEL4okaJg8w2PK
8wAfgJosSTzUeQLdJwkDfftaON+eCs4/+SQhVeTTMAiQz5EG5ad9mpyWqZ0zNJXO
dGuZzcbokeG9TEhlHeoh7Baoo8O+PdoEjRKkd6lizc75OtCtT2fmjtFGDzGgv90t
cRTmlJlA812LiVXe8pf2qY5C6p8zSlTyM7hYcFyYNdqLiuNfpqfEHtxfSirde2bJ
2LFxYMOez9WNkS+jqSZY3Tuulb8LJHAEq+vGeWNW39zjoOdc/TllCYMxN9Wds+mF
/CCPuCDEJfqjhGF0UOgd4ZfbEjrndsY86/7eLE2erSJ2aHsmS9pkWrOBI/cDnzy2
Uje4HYMDhc5nJXa6aBx6K5lFq4CicXmB6zcQZGya3J3pKYQ3iXjIFC+1zlxOhEXT
AV5vKtKAPu2gUgcnw9tALueDJJGQX+DHapRAejpE33v9HK/c76Mbwx8Mn5/oLbPZ
HAoNpCS4wRxni2lIa3AS6BOqV+nCGMTqrKkBVTpXtZWH/mCZ0gc6sRtyknAB06yY
8TZN3h6KfVynkObtF5S5FpeAwhkvPpXU16tnpb//tL5fCEw4arS0rAe4qzCpZM97
x0M0rJmy5QmB/8UgyjD4aI5V9Eom4sajWW94AP5RKwbwuFMB8+5Nu/U1A1svVXg5
U7RMu/n0kxAdBPjmPLsO+bnJGmuO8DUgVa+z5E5xCskAgTeGTrkWAHihz/O5JhcY
6zX1ttm4DYz0g5xPFYtcu2hNBgsGkKwpW4vfzTPYs28QjAftPxW+C3uSXv2tBYvD
EJvEDABl4FpFYEocuyYlYTqQSHafJ46TQBGXfy0o9iKoFOdTH2B/T53AaoD9Yb3r
VA8f9+sVoaldImNi8md6o67GOUmSypYPxY8cXU1o6SDh7c5i7zj3GzhyZXgwzUag
6cSNXD+22QKCHIexK5qxyAHQlE732BlLWHHQarBiSNTF/kZANcEoD+XwD7fmCI9f
iQECoTC+TeS3lR0jUQ9JYdfiP+dulRL3wVGjaIRjcJO10BYlTicawPHU3YoinnEb
haqGW2C7RSEjRYfIip1HP0hy3r/AO42LwJyQSK5Q/flpgEC1cnKet6aAGXJF/Q8s
pnU2bLr1BS2UZGwZLcv3jkyXVCn18Tf+fWqL/tUgrCqjTYv95eb/OBuU1vQhoQFW
uOunuf40ZMbd9KuPb+5zQ8ygQFEMnoi0dlm7UIY1/l93jq/dQmSBKcac03Wk1Z+t
lWyv+mmWCRqTfmk7Aey3+s7wgeITcCanfVCpk6Gofl0irJsVG0DCNBZ03xaWMyVx
fsW3e1ig/h0EVkzHm7t5HftLR6VnWEY+Uiv9T5dsp6ahCcQWxOxr+/rmONFVzSOk
jRJyDIPqMBK7Eg2AbKTixtqqZX3gwSbr2jnllcg9wfqaMl+R8Sf5Xhui4yVkLRXD
528jTiNIJNrQUeSfO69QEyOB11PsfN11WLh6aV7a1R6zvfnWITd8oI6fbtaKfsZU
S56p95DnKyvrFxNe4MZgZFXhZ92LfXpvj6EqKvwAqfLL6AOEzwcWEnWue4ib3bte
Tgl9gqf5ziRaLfMpexs8joTuxMhw5sjJwevLm6YZd/By7tddl/ltX4u8Dqgpy25m
H8jS0Ow9MLxXgUKaQVchjy3L+hOLSaMMJomXJBVckv2xJ8jXPfMxwSUzvdJruls3
da9hNvdQs2oHOvYK1PhP3xltbVvZqgCWLrltFZ9CdUeSRx5S0OPd/Ujlsbdw//Tf
WWytjvscJBgOYa1fOv0E9iT5+C+yHE7nzbkrSq8ejbvAS5b57j1Vy1slV69f80st
El1MdTbo7MhOB8tJ9Rflk74Px9JnBKOZyjyrCuT7h/O/ZqSPDYR6HRtUNYVEDP61
tk+3wNaS4+ixbb7nSdPUHzo7hhwXBcjsnFDrCUicFJ7QJGNDGqxb9AuoK0Oqn+H+
L8n+MN3BKSUJjpz5FBIR4zW5GB0QPUbLy5ccZII8QX2SouRCuRUD9VT71VHqTBFc
1VE36lnZw326sjnymztTaKHy/4h+cOBnya+B+UEQkyPjUOGhAguCmO1kOEOvCpI2
HZVGyqpxtOMENEXJlyTixbbVnvvFu7onimFvlbmytCrqyW+StHDBHpA7UbBgHxJ9
dpRw7evTHPaFwPR5VVby2480gsOs9g4fyX4PuRF3cyyUWtRrxfGBcKJdiLmgKMn2
j7pWE8SiOhLDBwH8jRev88eLrauZfDSZUnPFditLKOhFznKC8CBDOighqxAHSdxZ
15048AK4Az3YxQm5gVan/8qvV9lyn3OlBjOmoQQqZqaF86ttGnVrnQ/GuLJIdjxm
5WdGBHw6h1iXExlcCyVmQvwon6CSdy6SyV9kc8tEzLvtEYMjSBBmnABwmQE29Th4
Mru1k3XsJRkk47UUbNcLRsAdXScMHOlF5DwPWDl0QpRfPGHs1cdv/31t6pyi3q1W
Up9uDQcfQPHELx5L5rlwax7IXjI2Ap4Nvf+XjZtVwuTXRmxxpAUEk/21F1I9SkPg
Lzr9HInFlFqQ7m06g23N7JyjvpTlapsH3FriuIJZPDd6GqF4qqYEhoxP4kTd/M63
iZEhl5iz3PZfxlFVGX79oCuQZ+Jvuha+HN1q4QoLmyj9j56PCcNQrrGwRZuRi3Sd
1g+gfXVWs8V+GKP5sJc74+ki6SRKN/2p2AxSvLkeLQBKGk5TbOdoUiCZZx+ZPMwV
JtmNWTL0ARfm0xJDflz8/JbfXo5VHlPQGqwNghiig0GoHRq9pIMkheWRxKQU5YZW
yKc86N7vEzxFnNuPNttfDKJWemU6/FRta/Mh74Bx0XLc1eHw3cetdA/p9V410z4A
/2DYAFQdA+Ue/fCqBOlC3G5zy0ELbmdeOhegVxRJyBNOoRzEiA37ALNiuO7Ybcl7
QHGS+LXtzW25R5T2egCBBAAqUSDjZrkNnQaQNjVxuECDJmEOq7AwZNK5T+mYN6dJ
Fqi/RdlxYcS+fuKKKnpnnaWdDKrWHJEdLzGiXH08KX4LVgLVj9jkI2RFkIczYIkg
8+Sq2JQCoDXV/FZYWLT/TPv3nYGI72iuo7aRzMt0SCCRI7Lbug0OoXY9DzhCQmpV
keMGcgu9ShY3PmhhrNJkudTzFUCnUjINxkGTu2GyaZVKAKOm0zpOPuw84cnLLi0a
gRHTT2tiI3foQHGj1yah3LYJlIdh8pULt7nw9yGrUVBEgwc1NG8wGWMxPHGVbnWS
WjSm9t+fS8tJ0KFgYu+XyiJ4yH0P1Q3Dp7czxgR6ZFfQtSJQ4a+bW72rpfiswSrP
fWGbBmdMHL24WCEFo8qUJfqNetLmBkNIhAwvnQepf5s80UOTG6l8a+asYoYIdww5
AUn5LEV+VyhkFaqqTDp6a+SIB+PqOrShqzacKT04Ux9QkhfwRtOApBsOxShzl8lI
J2UaS//MUjv6qnuC7g6QyuBlFy9sBmLPfGwKuU073PrKvTpA69IsEsTRIPZ/LNx/
K/9XeoyYzuZlXRRqRkg9K3iMIDmFJ65FkjogUJ1KKxoccccD586/UZcEpTYFF6k6
Wuo+9ejjvCl7ggtz6m4dxB5IiU7QdZxPh/SizE23l9a/azq7uDJWVq5JVOEzcvd3
xWPT8sIEFjr7daazFJekTAcupIDJn4lMhr/mn8RgNxyGPWE6Fw1NhnbZa3d7REym
OsiTj3VakIcSSzAd+GU9ASBlkTE7G/esShNMWyCbEuVE0N+PI+VkxuapcZVqMwGU
TbGY0S3LqxDlY1tQkP8VXLVseDv1dhthz8VIi1v7OIwv4vx80BEJGyJfVs7RgNb5
TTmFt5N3fnkaD629N5N3zx2QztCKL3DSnrj7MgB8JyYT3/QzfdI1G4Nm61rW0Xnc
gGrulRmLaRHg8Hz5fpXK6cMZuGwAqFrSRQgwyBgxA+HGurP5hcHo3s5+KXTFMNzY
fno1S6OO4Z9z8PI6N1PQMHPvTiKSFOPv3o+QTI9X+YMa5h+nufEH00AHx9oAaOeG
NhzhWGZzQ8Eav3G4ysOzf3q3jx3QwApuE0oADcDRsaRo0ByaMYkk+DgCI7G2ArJ4
S/s0HiuAdzPfOt5DM1/C4DiD7AoBzUMhG/3/sT6E6VQr2F4ldrvjHg4Pqk02BYQi
fYwV//SyHULtNj5/FGpKM28tjCzX5GKRMs4sir7YSyJJhZhXJp6JK4F/GoQHoaTL
guUOxSRa9JepIxCL+ml3WagN56Mv0UVOrDXobnodgZK/MvD0zqtawl6ncSrbAosI
EuaSMfeCxNzJghFLAnsmygrfPpuKhzfaBdQHCftlO394SZ5/0OQA8hAZnYNKHXiy
FtSSI0KRKrlL2o/P1NpSic1eVsi/wXJ3hRIPL95lG59AJ7dmSjR9jUd2DSjueXuj
z3th/fnwEHm51mL0lJdaz1kAO6ibDXq/u6rtrBc/YGQw9wXDiD2PQ6CEHWJPFnED
PGxKZh7ZeVZGcrr/85+wDZgvZXC7nPBxZNxH5WkS9sZenJb2e+ivXJuRJoyYals7
uvI6GlYURgTHmWeENb6eDU6hkdm8zf1gwdfCDwpccXBhbCzmZvUkLZTFH2BM+Y8Y
FVUSiFaul8bxmFBqezsvEHnY9wK/JSoY+Ztv8//iCkigch1C1QEQYk5OpIeGwqE8
iC5Yc+706ULkPhf6cm/7Ar95Vva4qp/wWq14uO8qkNZN1H+SWbySxJDpuqY5+Ba2
gfcl3jkSfcx/2dTnc8DCw9Fgv2gmkqmHgrvIY27r+h43/ARxRx7AdXr0UB/6acKh
YuACCyWDP4Y1mmeQf1gEZfQiXbzcWoBVMKcdGnrt3UlSz2br+uJInJYl55M69087
Zfj6cEDh1JXrZKXazwLAGbG6dRzBPqfLNAAWEZb39yVbzC2Kzlp2nqg642PprdYW
CjaerqcNFOnvGzP9Nwc1F404tPqorusNSEYeW2ZNd8eWo8O8pVt1CokJgR1Cx6dj
wagY/W5BnxPJIPHUueDKETep++jDE+acSoqGyMrChsA=
`protect END_PROTECTED
