`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2U/zEGssC5sjjyS/gXnhz2A3CcbDqLZ0l/GeBlvP2oqQI/vqtbQGjjhAQCihlHIt
eBTJXeFJ36n3i+DpaR6FPM3zak6P93H0W/pCuVZ9Gi1l7uVgKpYFD/pqs1XyqyY8
XE32bOU2d7OgsU3Dnsykc2CIWo8lEyXrJGeQjXIYuYq/B2YbekDBsxV99bwwDbE1
ZvCm79yAiHqeOiK4GWV0ggHtm0C44m+ET5T+LYJY5QANbV4xbJR7Pa+qsSNVJ1TT
8jYJjbXiN064Jk2TpyM7rnJmE900eKPXjimvgPGq4F0M7RNnweMKWi2jY+fidNbC
JWpCDsi2HkZdwo4g22iq9h+AcmMNJhhkRYcKdOxQjN350s34CclyDSQ5clzw/Gh3
TJsyTIj6WmTq4kAxlVfa0pvt97sHszxIhWwCldLdzsCYgPDvQN215r6nxHF8NfF5
UIhSzF+ijby1cJ0K4k7IWg06h0iWiG1P3jVJl5q8BSdZgA6nL6vAC2d3nSywKlks
PCszz9EsV6GhbXpnxq/IrrzlXuiPd6+hr5owJLD3xokhl23Fdem5ez0+UYRXfORM
kX0R46opn9JL86rt4M7QEGULOSiCxVIG43oZM6RQshWLwQ1kC5iPS3I7ymJHVg0A
Pzjx6pyhpv7LOmy6RCWl7YN6LimWuT1S+aKOr65P21DPri0CbsGW0tsqgTXxLOl/
R015Au9QoS4Sc4Y0cdUA2cndKUw9qCBNfnROIQygJl0LgntdP1eoZqNu/twshQX0
ytqDUIEiMl4MDFvyw15NDSzBSthITAQAXAIcLUTK/q3wLnMCRdBhoWModEkZOUIS
+RKNjIbaFejRzwbZljH9DCorScYDnLF1z3ajtfNTl4jURrE2KEo/J+95E6moACFN
xR/6tM4ctTdGNxIhL4rKk5fWBeDbpmqlhpq62s6CuJstkAhQZwjf59NiiTV5FUOv
8OmSrQnGP8N0SL/FhqrsTfGDB10nEuPZXugC+F4y03Mux3cOWMy3xZaMN4/pYOHB
VEpEXUD09o9CDPwNPHC80au5AO4z5zF4eoqKFsiGMfpmiKbxiHwTCuEoeD7YGamH
cDCB6bBiC+tqP/vaPmK90e5ky+pat8DPHXXeSP8N9mBw5aHTDxWhRjArTfaPy2uv
15127alUz7aaXhFVYXl00t6p79mmFmMygj+SlXkzhv+KRg7DrmZ6AmGztA37rNbN
CAFWkf1ER48seiSd50Fc+H+BjiN1qIhxrUbIhyTuiCbWiXqhg39foflwQs5Jmcn4
ev77ESpFxihPA4kMD6JLCE2lE44r5f6CbveNnJl0OvUBD5NZwPRqPqMuPYdE7vLB
iK3NA7rHEm4nsdO4uFBD16I/W1vOvxN6azb2FTbcisJHG7K19lnVMd4P520SHRkg
YI1y/T9RrJBYcBM64/J+lvMehiMmZeXt0JfZrgJTNni1W6juSppm5awzfGBNo244
UaNI3AzDhb10uMM0QQtlQZHME+uHAxMZnFqQwyXSx3/J+Dl6bJv384Zzd42Q38D0
GSRb9yC38IFqag1uXAYL7jNJ+MDHcwG/veu4NuL4rJGFOaIoqhO7sGmy+IZ5JHYz
v2+Po8cWg5PV0r2CMatExMITXQKJKzGJtVV+EI8w342GDpQWkCQroUGtP8k7icC2
QSugPO7X/sEl3Y3PqnAqsUms3+qO4m9NpALc1Ik1uESWQpWac/PzRYorsVaVfiwR
JozDxFSp3KKQboM0HNaPDYgaXEbBGD7JHhcYipH9MFLHiQewhiCZxLmoscrVDn5X
0f5J25PEIWn8Wev+huETZM2dkwBOgbVaW1Hci8eZpDYCXYYo2HXL2NkXX6IT+jsn
1tQq2frRHmz9fbK4uuOdsJmzT8uGa7vk9TlqWOw2JQzDZD2dwl6zWs4es3zLNhBM
7r5mcL65eBfxrirJpqE1LA==
`protect END_PROTECTED
