`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5frhf03DGpGaUL3oXb1f3lB4kNIslXhLSgQNcNWj9iOjblOqm8fI10KhzMfKaKpM
viMP7rnYoEC6pb+B12tEfyiAqNFIimWcFgAgXAivnOBYqzYzZ0J2LG6SrgQ7T1Ti
kH8VplXcrkWq97pI4W83+YzMIE1nWZLldPVjlm8309rc9tOr3zSaJxhedqj2xZ3l
kV1AA3iUZyZ0aifCEU7iPLK64ZDQNbDw7X+sXr6DEyhRS4AH5uVikijTopG4Zcnc
s5HmckXcgypJu426IniVGY7ouBwQo4w++RHFI9ycIFA2HNdZP2rP4YvOlP26timt
I+SwIeMgM39DtwyjQ9NokuQa5XoShzlGaKQcLJM0frcRk2z/1Oz2lppRcAxVSLI6
2JOY+tuVY1Ggk8kx6nZV1Aj3waMc0XBOdCabeE6AbQtTl6s7Urf4UOIcdF+5dECo
MXFSXgqzSyV7o+7F2nFHqktfq/bFnHs/N0VJ1U/DRdKCnQwEM+e01L+v7UBjYiPY
vF+cgfCH0Hx04Rzg8jWwZIfgjVB2+zEuGWEU5jaz4H/HlWWsTXIdm/z8/qXgH1Ob
iup3IZJmbv3Gqr3Xh5PrxBY1kjhqZIxMhqo2C+i+ovGwyWDqFjze96fG0XuoWmpG
6bL3NGjFH+NzyqciD0BFukXiH/EVIIeZ21qh7VH/qt6cBzxiSWZdQiAKfo0ELSDQ
qrvWf4DUbG+qsyXFy2mS5YJXNmeHhcDrN1zCYgtBxI0JOK41qJOu9urFasrqaprx
RLEirFsocMa0cEr64dmsZOLl81EKurKPcxj8fdrOpJxMObcLpKxAcXr5Lp9Arzzs
jSHZIUpZigYyu7xRH7Tpn57/mvyaNuJA6EuGYp+FAzefzza5RvTP5rMNSnQ0PUHd
No08rQ5QPVdqgWXLIhFvwFoGFx0jdsjNXGLrMgNyqjqsK7r4n4FnBfUB1t+0wR5E
kFz4diwGh5+9v/2TFAaFMWzAsdJJBISBYK62vdphUzdLREj+VJbBYd587IpYdh6V
trz1CoG24VoA3hphBPH3dG2uZj5ohkzq9vB4kJBRY5+MfUF5i/ceAZ0bNxaIQdqg
lVU2HeSrIHM0Tn+APi5IJ5w6ZCpJbXcwP0KDlreEvn0IYDyphz/S1VowYf+EDNv0
SEdVEXbC66VA1Z9siIaAg0r4Z+X/52FAqe9dNJ++sDOZZkSfea6AcVwQivpMoXVp
sEZ7w1PLtadqivptNtuybqXfuwK46yU7r6eOMBBu48h4EUrUMmRrriMmXI2ZncSl
uVXIVGwu/DOy7zf96fBREtZB8PCrmJb8zYW5NqL9PprixkTaAzyK1P4qwridqWZB
zDxe8XQ1QFgDaTI4eAySGw6h+dI21btc4g1pU0Y2vKGAh+dULwYlV7B51RrPW05a
7Di49pP6Mue3T6eVMohKve1xQxWQjqkNu90XQRu+XcULwUdOhXz8PAW40ED3PWTO
cJqVqrUkxmc2HHt/26N0UVoB7PM4PBucPLN525Q381q9H+heIugbMUeyfwDXhLwS
bq0cFI8/dkAtf8hxfHd7KWeye/pV6N2yIlVIdeLAS7GY9q4DNCf9MzdfXVrP2kls
9PF/3OD7x1//YkfmiHFsUFdpuB4AzPY+o77RYOM9CoQX5dUnh2PzQ1s05ujlF2ww
x1RRNgmksNJkK2jKl8uRJeiLj5b/DGKNY2NnwtOQX08W27nSOLOXzMi+T4vvBZHi
KqhJ0f2O2m7gxw25v1I7AtGuegVR1Anqu4Rj804hdjoj82Ah1lOWz0pBTdsIeWP6
fbxrn4xlNcWHsyHKv4Evt+jDDp1XPHa3hSCU1iVNV5mDFmMo5oWlBcWUrFYwPfNE
MgvfaNy298dLVlX/w/RKOCszvNemUtQH7XVZy+QQZI76kCz1FLDUx+R3XQL7nZyi
M5eb4xB5We/uKqUu3j5BxXm8IB4GAgh1TwYsjTRUZFZCS5+ugVXjBS3Nhevv4goQ
d2BuZKbkTnuFat07G7Isxk1JHLqv6mu+alKCuiHIUivYHUo7oXb+sF1+LlSj4Pn+
DvacsofdhjuPQKzc36XI/ToNlnJUnKkFfdwxkpNElbli9FxQXU6IQ/WD9W3u7zBs
ClEDGtlTOGf7bLDPIEuPZM62zCyp2GR6LuOMYcX/7x/j9dXQZR68LUtN6bucXkHq
bUup2Dj9ivuiZgkD8Mfei+RRgHMUlBSWswyeANGaRZqjF5pxG9W35QaNm+PdlMpU
2KSsUMd98x+FNVZLZavIKO60Sia+4lOkwK9fBY6OOg9ivH51HGvbke73oNOqqYKW
xfj71ZhHVG31iiawSEToDCPaVNkrq0A7PckmiGu5W/x3JnJ/yRa1ewNvQ1bvSZzF
jatsOD80n0V8JxLQ4YcM/mZHk8oFJy3vBTguFedvEUlPp2yw1ACo9af+9cgBgz7y
o3I4NnzcPFvnbIxL2cwFChB0Vel6R4Z1DOFUH9V4RqLE/NOVbYqgryZfjNYiZsVg
FYvl+M4iXVLHBZgNYh/xDONDj2vx7x6UDrcGES6DuXU4pWvB3nA7s6nhUvtyZRpD
je6x7RrKaIVs0PlVbrYkfAC12TN4KTV4Xzx5S9RKrIHsDa5Wr+jyzhzOX+S0q8yi
Z+/76lILyXqAqQNKBclYdamc7AEs33YhHbt0gvATtpj2NVylSeo2J6LQufVtlLue
SeVZXNCvG8vHu9JCdpK93V/CS910ILcSycOBhy7hAXTmMdCqvHHqqObQjzf0Hj0z
qrUvKThcVq18wBAgqbX/7omCxsitxYp0CFHVvowxIrTDBrxtFG4iUoGeFtMD/aAJ
bcypgqFfQaTXv6rkYRQOO3e7QvQ/bVLgWPpwjER175ZUxajtoZmF9EIkct5z0AOu
ZLD6Un0aOauOo7r+M0N6GjNoI4bCjVjokvxPydKTU7bJ9DSAcMCwo+yBGbewog35
7svqAFoxGUpS3d64d+kV4PJ2UV+tCkppMFG0hCFZBfv+XOgdQ7VTwuECyv/zp1Qd
NL9ac0RmQ772u804rXM1rl5WJ9Trg/bggjS2WauStVfFpC343TExb/B86+/G7xBL
wQN8JtYDXCZR++o9Imd9lv+aSClTA5fFAZXsTnwd76mw4ni3WQhJiNyObfqfH8/b
0nFOS4KyKn1vHiAsf5+yx3Pk3fvd8ww5SMIlZQdr3P2ZgZfccNcKSwkz5i1HWVut
YzpmrWxMBIx6lmzFbde+H5MLywliDy+7fMkzO/Z3NU04Q6dogErv9ANpYu8o40Lw
rirEcyuC/4sAAssr39Ef+VAS7QzwxtPwmUqkxaJ/+JakoJq5xxAu9ZprZuXFuI+7
YOzmEUVz80SOCq7CKUOez4kipBroYxHqz27LNdlri1I8JIwole228KJ7gqB6iZM7
KjZyyvzVEZ0Lu2LNb46h69yJ/NDzjmKXq0KvkU0LlnPrqpobwoXyq4HWCZUj4TPt
zc+zWT9/si5Zq5tJ7FRCmJ4wLebv5w2pnL5s7epi3foOe2I1WD5nBjRfvSbD/+XR
8xXU65j67zjGlHRNdp4bUfWHC1ktoXjtVG994Tm8ZSChharK7U7okJ5TeDXxvL+t
YijDXoo3gcurr/gGO0MlLuH2PAXn6TjzCeUorccelZ9pXDobO89P50kgpZHmeKY5
4ttMDdQykZx4kw2Iro7NzeqOh8lAVmyj6w6QJg2tSu8LDCVrigxsXZ5HPtfZZVjr
Ed9LZJ6+OOCNn0xC/vOpDwN0J4reAgvp2mcCaD2eRLzhrevzp4Gf2JcZhlIY11+X
6XGw4tfgOaz93E6P1FaQY1wGFdLtH52G/yz6HMK9sv05UsUHSCjb0WUC8vigjnAq
zigaqgKOeGO++5N3NwkO2xe+9mXY0ccFXvXEhMlqHMNDuD1stfT+dYP3ERiJvcZ7
RG3Te2U7xwliZicZEnaU7tEDogkLvlEXxbInrxS1BuH/4nvH5UH1lgCu/JIZ7tBk
HhDgFk9q+xT9hWj4UhqvWnDCrGzl/ga0kZD2T+//5iXVcdMDfc95WImlN/XCew0v
ULhBHwxdAHVh8lXHJ6uLyd7WLkBOo73icGLS69NuAnzXZ9r+btuCBq1yAfMJDfas
3kbg78gXNTBHjISOjQz9dZlY+MhufH3nKKmnW3Qt+1u6xKSfhJsAAQEp4UEHWLRw
zCPPKuFHabLgf/gnwp320jg0f5Y29UzY3GKs5rvZxAgrH9sdegPJb+GArfEO0A6Q
vTLoIlXCeMq6c7SZkC29oBCf3tkSyEvnaFxf7v/pG3aS88Mr4J1K9bubKL5BirHs
gnTGBRvuf1sk3mZtfuNsUCoQ6Kg+MMODzhUQ7SzgeGCVv1N/Cm+S5v+JtxseWV1H
To6WvJweZVNoythnNJul+RwryJVHwD5K4fDd+NrkG3RsmMEJ9lKEZonsQeWTG8WZ
mjiM5MTE9Gl27PeDg6yflJIo4M6Scq3IJwCi7BJKF56bGFVTNYpyQUYjS89+9f4a
QG7s2/hH46hBzV0cHMIl/XuiYw5g5QxeNIp8rK3OviTJKHz3F8Yf5k7VCoKX/WFH
6OtdpMS/2Wja78/KegaNPowc2vp6n1z/8UIRkvLDN5cydJu6sEi+9m/fyPEGZ0tp
ibdd0Salo5F0mPH/+qPBUvCZtCMyBWGxsFf33mnHU+FeH/KAAUMOEm4WTVV4Kbqj
Ww0dKbiTg84rFpVvCCy9bzaS2qrzRbsDcmyc4MoKPArQYMnIG507O/ocAASLNtod
xbacmxakSkECjXGYMyzYmIteUOrxg3ynasdmY03csVWk3ZdpdGeypzwVRUyJVIcF
Hl429UvOjO+yN9Mv1xkBN+uniIs1yb/R07hKfuhS48SOVvd5JeoE1DGUAv9JwihI
KncVvXfFd87DWuBccoohNpJmQKsXgwsbMLl+Vuul478F2UH/1TwN1bS/IN0CbgMu
riIHeDT4CbTvgWBHqnIal6vnAMblZGexBP7H3Wb8ei/CTGYmLiMq50zg3RFOaL/B
++e5yDffJu+5GbpC/J67L2e9ZFFB+IcYKZIM3aTh/c7l1myZfPkVhfskmmpyTFwY
uUoV3kaUeXFg9jwIx2gYsfhv0f/jWfR03V1QGAkAf7s18ZZXcqBIKrK/0oqim7G1
vzawHjY/+WSy5KaUzGO4hiHvvwKCwaadS/uwGxmkPqIB0EDK0taFD5bOCIG5Rj6n
hmbBpVK4qDbQ9YmTmg4/klZNQ2hKkyZXRCpWIYgHq3LJkaZFZgxPY1XXpGTqIE42
qQTX1wr73u1AYGQlDPHs7I7ak0x99CR4IsAbEAInk+s/pfGB01WpPiiWXQVtpOuU
IcFijezK/PcvxJ9RIxn8ht/ma+ubIPs8JvLQEb/AtzyFLL2OA7mvJ6c7KfnZJgXh
BJJvr3aHVM9lePI8lKyhlvYewxOYdwXSKZSf6UqXdxcVsD8JlfwECiG8/57wvek8
kTzCmUcUnE7eV7QoS/oTXagOUll7EbRomuQ9ULvKO59ggzmLcmSeBnx7QlAkmsnT
7ewdav2NprZ97J9YIWcqFh7jvf2WEL4SFFQryxuPEteCyb6/HXixmuzcMfTnAhn+
E3Xg9m+Ogw/FuXYEhgvU37TYjBDAtCLQX0jW7UsCKtagntFPAiTZ4Eq4DvyQ+k6K
vJsHwicYae5Hmg7dLnkI6XbOkz1Ac74c9hQHwn0N0jLbOp8vjbpl6VqsRRyroowU
9CTq5qhdFfByGhJ4Haeted1GJ+gw1SfIoBJ88u6fNHCjwlYUDQEcYAqvcjjdhVUd
0hWNtIST1eg3oQe7/0NnfSEaAHJH2XpDAk7AAjBcBDy73Iu/f0ijaGbRyPulABxP
9dDwuKC81zxtnghRvFIJTcacv2vXaoUWWZQs301WUE+oyiCi8fXmsIIVogJDc6oH
CpGA4UpaVYmChOyvX9CctMWtvJ7fQrcTgPsrILvMUl8hqYksUPHn35a62Fvwc673
kht5lOoSBsYhGc0xiLb397S34wUOzs1wLYGbp/RayPNCYJWMkB3BJfmHlZ/dU4pB
mrR3UtW+Rps4qu66X7sl6ppkba/UY8bgr/7GY0PbQRbeqmqTXRHQFQH8MuS7XpOU
ilH0MfRWc/Gu6PfGEhfzDKgI1JJiQkb6sUcae2rJeo8G8pZEdg3xlf+GEVq1yZmb
boiwPXbaEDqcGen8rGPNkZtNL6CCeRbLECmv5iNvXTqdo0VKyBimukexoBnajY0Z
bJSGvXZCM8dIxL/eCZ0RmmAB/lRoWYJ4qP/XhqsjfAWFHYaNq8WpfEsSPHm4xDRl
xVuCxxsnzi3Flpshum+KS2UXOh4kBetiyyhy7DIcLFRUZs8cNWuuanOzHT2bBDdK
MpTxLV25ZZpNWf6XWYKJQh7Th3dWqbHfIc/lcGSvRlvKUPScuPqWy7hLIAsNocS6
wyYYN1Tl9ClbFJnlA+l1XAhnNhpkf9qa+Qu8+UXAiJWSucXDdCmzbXJaEbx1A2sj
RpGloVB9rcWL5KRk5yUT11HwASOYEDHpIDRGcfagHISEwI+7CbzZ5x7NdCWakeTl
6IVQyT9HxlwVf0RwECIL2v+OE7xma4LbsEjPXL905DJdCYfgFlYBLVRPHz8I43PW
w8mpEWD/Vtg5TT81B/2SIJ0l8+qU23RbZZSOsoo+rxCTgqaR9VILSq8yQbaIZ1Sp
Xa9CjHNEjME38aO0HVIdsC1yniPJerykesmv4P81UG7H2key55tkb5zdFQ2b1trA
lePnHBavlV8zPbXG3UziQpEQ9VSQPUimBoUMd94OXyNKQFmFpkVgrmv3N27RukKx
ROZ0EXs+u6AUYPzS6OMO9U1fLTaXK4m68tcAjNK1U96C26G9lzDGvz3zbV3m1P1k
L/aoWXtM/apc9O4/SCoQfKUoLDG4XOUDdQQE2YyeBdjZY4UQyB5F/xWF3KDKfxzB
lBVb8apYhdWmLBytgbjtuQ1KYcvfOlMQqwlp6ZOw/9KynXksefngCu700Ak35nR6
8iNH+GbGM7q5PXeFUTy5DKwkT8N5AhzKRWOiESzwXg3Q2gvyTlbnROPGyt0ZNUtO
BL5vgKnSEjXLuWiDTvkbvdAXsY45HJhdkPpGAAsjf6VZ2ZfNDAJ5CJtIwaSa5imN
t/vg66HNL2v0BBsqHm+P/WAoDKrFdRY90ZTgOnEEpOCaex7YzaLjUvK7iivFdMwl
WzomIYcLrvc2DBZjz4DPlwTPxkocXD3AXl0EiMmYhl6RkvcQirXAFB39TsesiRDw
Y3vTfZvyhhOQrlO/30zlAuVR6j0xRoxBdAYsbRuQONIBvtqmg3BDGv4ao+dCsRA1
fwFOic8ayomqFmomRH9AHhlLzjtodYhHHq60ZKrbxhKwhGlsuj510XuMd7RFTmfy
xX61II1BHMEHeowBzChgDOrTKDElvcizF0vrZ6+TMEdOZJnr6//d0fMvsYh3Rsr8
2ZTD9RzfSpOsmYBAPWco+ZBCqHxA5n9QydF058xmPpgjvASzn6H0lH4mzD5ocufN
BN2wdbQL5nsw+wZTdZKD1MYOu6fp3bMtyfc1GjNwJMzdWvbdV5JBLxot7cTc2mF8
YY5K7PaU76LyKlFoKQ+eW/8Bx/hFTVdwUoiLXQ/xfiNBVMLGgdfpzUgAZ6dF9mgY
LwP+vQfjGZx96GkPDTSXYpF2IuBGK6ciOrZBthGWvKpsYU0ZRqmZ9g1pCtP3zJjm
brLOYO70Y6foaX+RgRB0ctZsmav6GwbHa4GEWnNuRRLL+LYJ3dJMRCsm3s2e0NMj
Mg9HzNNnp/ovtzth9h+X+YYT2sPK67BkEes52GPVjX0ix4k2748Je8Zo4gKWZHA5
IurbU5xvuGhsNw/K8KCqmtduJNZZx9cADh0CO7OngX63L3qOrfqNek68PfBYW2+7
T0GPDFVQbkogubrVQ92env4nW1xsfBatAEOrK//2u9tzjbozPZJQ/tEuZNgmpl6M
7JIL/uSOYDLCUNOIfJSNuUllTBPHRg+orCOodpxb4OMk+KjSG8VQZua7ekDRp9KT
Mp6Fq9GsMj6YhM2t7ojn/aaQmhiiFRkRoLd3Wp2kBFyGUe+v3GloxJ/sHoZYi3BW
T4R5U1VirIDU2gjQt0toEyGuQP5w3CQOYBp39SwZ18EegRdLD430GC96aQU34ubt
SdcsBtLyWUpioOQuCzelb8ArPVsX8fNINrp1szzx1Y/UveJt1aWTVLErDN2Esxs4
pwTV2bjki5dLXB+C+g5uS1z2P5kO7V0UuSxQRdbNqoPz3LTDBqbpl/XfrdXkKvzd
Yd9OYl39suEmMPgaByr8+IgIu7922yh9fLbj14ECikLHGZVXb1V+QvY3USbmepsL
W3wYoDNrTioZXeEKgwD1cpf4aC7pP3/WhZ0fhyo7Z+QtBgRkTQofo0q/DcPuD9mb
t+TCs5schK11AjRvurlxV7/h5UuyS6DL81K0gaEMzZMBaHH5E//5zXDolrue0+A5
nQN45hm8/WzfC5tukxDZgEqqiPTNuFNpko7YNUC4hJOpwi0xNmxe9n1Hpe5nUxzR
vTnATABSKfjFHsbNXRkdPi9ZGahuzhGF2FqOHd7sni2dx5L+I0eKfvIAzWR65acb
QWIFi8YHV8c5i4T6PqlEpueqP+y7Ei3DtA1JHzUiZos9AHB1bYASF/fyimO4xLjT
HtFcStyw7EvoGRcHZZGAZmgxORJe3rHtbHNXOes0WhPSw0O4xRcLEjmMqEaIJZ1f
2RCfbFEx/XMdETJig9flb4mpRqH7U2anOgZyF5jAUurSUy6V5cGp5ZZ2MN3niJuH
VQ24c/EDt2yYRPcm0L1QRV7v1SeS2E7RBvgYHrF3MvnVjhGlL0iVOeS/9XwJJvKK
ehbGmxzWQfGKdDslpX4G5OqZgXxsRkXiDwK1AL/F4KqvNCo30+CcB7Loq7hpuzmN
4jRBKhC+5YLSv6K2/6oEs4xac46gC75soXaVNlCV3v3f7CVVBdb+oT+Ad/12j4Ku
OwtGjQa5sD/319SQP2ArRHF75ZWeH0IuZ09oaoh0N4sbOGac5qW9cVenI2fpWvyq
zzWR1l53io1aHnKMN3H33JSJEDKSmzPBunoOjcJjZipnGr81JHzb0mA1p68nIn8z
j8FibBtMHW7jqkGzCmrSKPC5eKzWMbcVHudAzUQbd2aF+oaFwmpm+j6JurwX+Q+F
I9EvzVYa0/aYRgY8BwUKyGzZxLd7DMhj3YXzzZWP9e++vKvm3kLmJinK3RIT7iRz
1BH0C4caK+PWGdCQSxEZD/nO2+XTgS8gBZMh8PG7eTNxkUrM1eRkTs3gJQkdguLI
7/Vgc4RgIUPFFO0xfyu2i/U7KSr6DXe49FheQ4wkP1E1YUHZfXOWij5NPQ9l6vbB
T79DX/LSJ0e+BUhPHXU1+93GyxEk4yiDO+HWmJg2VKTFw29hCRyNbfzeMNL8aXU1
d2QSJVfy1t8SU/Ehrf4U5CpyxlSuunwkU39GyMbTt9Dw/eNr5t+H/QgHpUoS/P5D
Rvyahpzaex4jQDZ3dbZegddKT5HB2q5EaA32j6So85lP3pB08pUcpS2jLuTcIG5Z
NMQGxC/xaiqaY7T2DK+5XjEFCR2p3WIaqQgfXXVJXqZMaM8k4htsQp0Bk3FtC85V
BeLj9HmyRaUQ8pSYP8JuARZ41JBKPb9OpCcZLUcrm8BI3NvVCix00VZzW54IuTry
3PRRtvE62Wxp9Yd6U6ZFPComK7IDCHQWgeVGMZXiYuA7NS3irneXaFoKgmSSeXfg
PRRtJQd3wwPeEFNISxOg7SOwA/Ft5j+GhXLjwbZc6pB+uUdFTD7Pfmiexvm02meb
fbhEwwm+er2r7aRldyB6EYEeu/pgddC1JStRXINcYNrF9uvfP7zInJz+T8sYDVVI
FOr553eQM39fQwSib+DXned+SRFu9Rsl7AztDb9A+4GsrGjO1KUpsw8hxRkOr17y
RK6OOu8d7C8vkgIC2mnTolk0PmIsxMAvfX+hqtVsTa3MT4NNPoRF4/kogGGDIS57
4ncNuJM1slV4ZtaboG3e3JuCsDPsJ5LPxDqqpEjx8dkYiuv6hWihynzqQ6kZ/5uw
Sk0HriNO1cwUcl/UsMUWe91V9CCmGyTTTtbPjVh4uyIgC/MzTQxgCHteubRLVqiy
zLVSQWMzWbnsfK6FaekAW92KwJmreaHyTct1UG1DfsEIcHBqaJlkkvMUIC6BctQ4
xqP4mwWR/EqUj8epuxtOPmIdCTlIbqH5bWgdHjzmbi9tmTnqOK+CT31wj0QaiZnz
dXN9dpt4ubEA4Vj8C+1hxYf6Loq33DmDsXCuiQWUC9nG25MHiGToXGpL44uzws7s
5mkhligEMm2+31Reyu8wuI9xXPzxBvL9QOMpBAV9ExFiWrRMz8V99ulNA6i6epfW
evExxv/Sf8wzhJW+nb/QICuK67MvqhJ1qbmYM9JMWvOW162a/qbKDb1peqUJZ2nC
wAweFkHJurm22gCDqBOf5l4UWEDOzZIl0/omihBmCs7xPLeZQRuNCVYMBlWImhWK
czu6KJi+F33BqUiAF2aj5FLO2mO78FP5DMr+NKWZDzsbFEwF6Z1sx7jepxmtIEWo
riUwvGKrj19ck+Da8TaIX9Nc4mFPdbl+vqpiYrBHwKhW3+QxwBz1uTdhvDjf0Yw0
zLJ+awahPUC8WCdE0r9j5HgnLuRBWPglUyCIiwqydAOqqQjRPJCpy/GzXw10NIIz
AUh89R7CEFSwCgLURnFI549PRsoQ2U5l1smGNkvfnuWR0OOj9zGqk04rX9pJJYol
1bEJdyoh+C4uiumXHaodvh5+PtpsNpWNOtBlSoBSratRxIruhGp8VmG5qz+B0QGg
qMQNkCPnGnn6lbrm3gmCTLmkQ5rxC0x7kcq8MwNp0jqIWxkaENnJZuglO+r9FIyw
hjoR/tuBQh1HdXk3FWHOCpyl9gdqZxqSm+VRNW6VwagMqgNJy8F5DzJ+g9mn+vpH
1cwUOtUl/JqgLKe0nazkJNJKEma3ldQ5ZUG/jAfbNOAB/NxEwmV7j/62lciSkIhj
XL3qNkeEXJbfgsa5oprcdA0MNDJjS4J+mIxidfVNWP6rZa82VtjdBjeBlzzGW2ku
oj+HfJi/nz0TJyk8kQcP2sIcX/D9UxETUsFZWKJS9bOw0+QROnpLY4qELdEWtE8R
myZGmZ52HRDEufeb5zHfZXj8AdvuJDnybKlR4BaQ12LGuEWeBndK4oWOTUjPnzqN
+fgrmN7ciFAuU2B6h54GGdWosg9LV9k5TS6fdjz77e+XBUnZvrt4rzNwe6ejKi1s
oUcef6OkHW+7R8gm4OWcDGvAdQoSqzl/hHjC5Z8SDuRGTOnaYJepTzrn3FpLWLBZ
qBjwyf6W81LSxggMb9cxxwYV1ka9/+EJXvW/Fe3XN8OlfR76UwI/oEkmNr5G8mN2
9h6ArA7SmBm9hbPHciBjVQg7m+mRgVrdLN9/BHq812JyuRTyWnPXizb7G+f26kXr
P/Y2bEcK0FeKaeQeNTbzKPI8FCkOG7yPIV8EelBokrp59JQBoBBNxlkhN7ci02Lp
GMR/BIgDUgYZYyPwY24Lvqisgl31RB5n+nKrsnI8yWalI9beYvb3Ew0vTVYJN6Px
C1T24UsE8ecNoIWU1JQeVf0BpFoPBS5Ky6q73FVfojN//Z4qafjQXPNx+8qKgY/C
k5QZWz3clivZm1NkXrKtBIWBUdNjiAMMveL2veX3nR/cBt9RCeHjd5by9mvjv3BY
hurNyZ33fxr94T3BwN/WsXL3hY7TlGjRzl2X931UPSzoIzBljY56dgdX79J9RRK0
B0ac+W2W/NN1aCTduR27Wo3yUdYu4mItDsmrHIj1Vlm/DlNoGPPe6EbUmkgBgrnd
NwGXUumM/MCR/QyfUr9hGnFP4Tx1dVjoUN8wG46bTLUbcVF82sXEiJAOCLPGWKEm
ro0Yi+roL/Gn92X9PCWpCjpN/Jv1RWhX2dTuJ1a5VG70sAeWXeEDnon03Av9EAeP
pxBShIJFTEF4ReqOHutO621FhhnE7+py5u7uilX7vxkBVcaB9V4W9PV6CrrpT1go
hrSGCT9yoQEJTxCdjQ16ckruStB8UNvQ0YrOKhYkNuzJq+NQ4Sm4Ztva4gmhziCc
xw+GP5g8TNXyluiQBPxYVN1TSEbtQeX6f+LUdxAn2TDTRuoe4jAZmnSWnhvYlXuG
OvjJfe0zQxjL/u6ViawXDgFpUH+0NWpSpFkIebtJGbWh5guUiqQOQR1eL91jw3VW
1LEXNngStb/aiISSlDR5qAjivkb5dnag5DdRGQFgnlT/HDue26FL8pmSSZwhnOEJ
CTEfgpOYXhBABKtBhz+BIRbVDaAu93TwvCeLqEnlxlo8f10iR+2txP+uI+E+cJM8
QSBInrUZT6bZwKaV2DXHVyGAXHN5prIShXUgm4+aR1BDZ59IZqw2RszcWc5c9z+n
STvGnAxvYUQCx/QyQETZVk+Z9UXuK97kloxUbkDc0aDozU5BiXbPBg6FsvDybPvl
PDQPNoIQkCLT027HAPziKBIUo35WIgFfHT9uH/MHjUS6hI7frfsYFIz3RNm/b0Oa
i3It1Z0JHyDnQHo3/CJstnRRVwbOVZOGh+inzGBGB9bbimV8jO26rqVRGJWr3C/l
1UxI7BTUB12JFuGK9/J6tpXx4bwYqpiAYolD5QWRlc8R7j3D5aa2h7FuAglPlfT1
sb92BEdSKpcIypqQBy0+eo5cMvaYyChmnKTxWN2BvwqNpVVJKzExrLiVpSMsAmdQ
3l0S7EdSn80FOLUhPcVfI/q888MBQQeEmg33dRMRT5Q07HQuT+kgBPae8Bn2Mlyk
zjEnumwk4jWC1xeiBgZfpVkehe7PiyXEBwisPEsbPDDmUtCCzUz6lXZEfOW5c0GP
jd7O5Z4IEphcv9+LWLGafFVYkOJ9MnBUqwnP4Gn8XxMl4eRZ15UkQcRYiQuWgQW0
o4R1XdwWmGl1RNM/itEgUX/PLMXgOqtAuQ8Ss9E46TPUx4IkxbOZPkoHhvN5i7F7
qEBOLDvGgEstbdWjvTPeJUh3aIVumJmpLrMh5WVMRlGH7R5SjLC5dq5LQCMnIibI
FgJVDY1wuxf6eYMavv8zT0nJaQ6z+0wJAfRi4kTYsYlGYOsjsd+LAyIcaZblr/S/
z1cL2EGtw/RYsseaKMxUJPB7tw2LllCf2vO9aWMxRTgfNmChxRa0o7A3FDLfnXvW
+B5gh+yeYDFmQygYQiSQH9cqdogSU8W055tPViOLFIx42v7OvfMjnU4k28jnXBQY
dd7h2aJDyEt/4zFlZyQqJ0KUYBIwiJ3iUMByDfY7jIX9gLhhlEpvXFZyOWvGuiBZ
4+HeFJn8RY//lp4La9RgjWETnJ709TcZV9Rl3cA739//cyXgplFdFUXbMAgMChF6
EQsrl8bYe15h0DaQKN+PwvGbippZ5iGAm72TVUt5Ruf6rkRUO5qaWqgXee3QIyBV
vmsS9Pn/8X994w4aGPH3AK4U2Xzap67fhs7w3ACuaxMNKLUoi7oqkA3L72/Lj+oD
s6V+qLTLRTCvUQTbXUEZaTlQr6RsWyIiAXQf6zZ2G280p1D7kE0qiH/6Wq9cSE5K
AaJ6Lb6I0IjvXvo7mJCwn9AeJwMFqiRj7GsNKA92VKqQknnbI9sw9ShKHdTSmyag
FvtvBLIXf/w/GHYDK7xy5jgT5B2CcbIaqiCRLsXsvSVltStk5LalXqy9CPCn3yTe
yYO/0mcBuTvvJEIMDftYBFQGS+S71so7ligiPJCc6gRlNOXxnOw9U47/Ij2BDNl3
hbA1ZFiaWdbEaJc6as5L2a870e7revVjn3kvdzAL3Ti9Na8BaJgCfjdDxsfzeYE0
E18Sj7Dh1D4oF3kNFInrhXJZW1glCTaY7HyC/a4JlUPpPL8DUnV3b41m/7zs52Fe
NvS0DIOryGEEEUIL95N9mzZt5YWR3iEDkNqB6+ws+PPpYNjbc5UBy+daiP7KQN/y
1/2GvhXNperEgQPZ81tuDu4l/UKVRIDJoka5jZ/bxB4/issXSERUDLfsCDzcmdOl
qImlOPxhfEBxiAL+idqRP2jcB0gV9T3pKUs2NUQbjfT96Ij0tIePT78WRe/Ph3Fw
XAklKJ4hZ+grC2NeueWW1o5FzUqBNkocaBYquWoplKYC3rGoi3WdX12ZC8U5Srhg
DgBfD4gsr2rsnpOLoL4ZV/CQybwjV55N9cvOHeMx7znuMPQk0a3o60OZ1MkFdfI7
ISdLuixbsw9T0+v824ktqeCw9Gj6nxWeV3ydo5FZEIm9FMYt4f1aTjpD5pdjbg9Q
mTpHoUyo6U5PPKCiFWwA/TbrnuhYsiP7j407niDOyRIOF370IkU8na1GI1xqTmw4
E4+nOBZC03oxxRp7JVyyiCU3sQmdj+uhSbCcQOEV/r3KIVaHwMxYqUU4gClSUzEt
Y4uoSphXHQHSgIUEOtimOhvEDTeqH33ZPVa/BnnMO1KDztU/i99P3yLYs3IL+9fY
0ddp/acCMrxJAxyGPPLuTkpfMe2P7RbosfDtGzWV8ebZYsJGKMMTj1H6Xldm9iB1
lM8YQISSFS3XQs/UN2jFLm6KG2nhkFDhNXhj85PKlbjbcH+K1q0Qmk7F/Zb++eR6
cd0+pUeWM2iK32RNu9wrSShRJqrT2XWKTY+YXf+eIc76c4C1GylWhl5KedJe0tHk
J/kKKosG6KnAQYpCGqQZi6TeYUOxgFsWTD06bQ2Iu1j3tZjpASdeBjgaEzXJIEdW
TC62tr5hrKYhx5mdHffPJRxkKL67q2blVAKSxTKOAKAKAR4rHqwpfl/tIr82FynT
ZT97+FI2xZIzjg9li+to2lUJm0xnvo/76kZvq2NyEpg64lqBQhWG4wuW2N0SQbph
YO8oyLTXDLf+5eYDnW0J3+ezSisx9dEoOXmtOEHKwzU6w1emR1B1N/VZmvSLoDAH
cCmNDpWyF3uCG/aMau9EwBEkONrMd2y+YYrPmml0RwOY12HcfptRzVswajsHNVJ9
VhyRi6IgNWXjON77m+ND4/TDx9juluO9kBBAby57sNLIA6E6j2Ec7Q9fU25MzT0p
jvlNdSVo/KDtY4bRsaObP8J1NuCEFUKu8Ydg/2NY4qhg+suvcMHiBjPAbDFMhjuk
DG/XgH86Yk7YJKFpYAjEAI7xzRH/ggW9FHH3zBOJ9EiKhgdrlR42bRaUD+pdNcsI
L3PRx7MvogOun7hgzAz44vgI53utB38w5XC0MTJITgFaaXtzwKmAA6RXap2TVfur
ynqcoZMwPjUk/oeWaQGnY8GoJUO797y10c+eHjRhH1pjBxz68zA0Ce8QV7fBWzep
s1Elrt07tAQ6hk2yb5L5e4trwr6aayxCYqSebyZX2LUGm9BM6SaoJ7EzrgkVDTFB
w7XDI3zDQ1Z+uF+phXRXO86tLOodt5WLQTeXnC64yYnRLXVNx+XCBE1TpIQC8ObJ
3UJkJoQoZaa+PxQDorVc7lTDdpaPN5hr+B/2C6d6NbQ6a1/eCG9oopUXbLd7h1SP
cTm4c59P0im+CgVwTiqo/tKlqODt13R4V2dFGLRpvQzbUA5g5C3yN0/n2L0kBWf2
DFXCSpxH7/wH22Ay8SjrgN2KSJtIiLzAqjKiJF/W+039hyrmMG2dnwhFpG9w8x3J
eTOsYbkSVPT0X1qZxwBvRizhO2wgz1f6dXqa8dvU8jV5lkdGYuzC532RYNBmnECq
WWe0iN6A36BdGLF6InHc0KDCfvQ5TT6dfNzvSNzAJxvsT2jx3KqmA9r10H9Z5ApL
e+6M5HGuOH23zNncW1j273NtFbQODMuSFX3E6UojLfDP0nhN4dKHXf6Djs2wNqd7
CTaveqE62A/mLRocG6+C3wS6ZEvFV8UI2X5gBLBOA94ll1Fl+s6hObkMHqGWCDRj
pcxZNUDVXn0hpd8SGuK7/YL4VOrPD9dJit0hPpPuWRwR60bYQmaTm0Dq5rKa6BAJ
7cj5eh1pQWKUx7KIDX1qwOZ+aOn/xn9RIeSJhsM8ZU8+YlLrEFnKITybZ+UM0VGr
G7Edag9Bx7NTqgnnUxz0XsF+IAei9YAtSsUTL2Bkl5Qt+L2gU57ZBHtKpPDQkg/Q
/X9rblQDorkAf0w7IxzpJC1XQbgPtwfcMauw+TD1D0/itbeGNXpyaHvaROcNbcLc
Nrktfuk7jKgUph6QSOIpTv45sCdWoX/PRepB85+sB7CV4QaHoPPwJ43kF3NI69kT
WyQci67h+gXcZc5m9FRX0qndKrC4cH+xLzoIGhJQ/wV3Un/AdxlCJDlQlDGD8zH9
f9A2P37TgJ3oKbXG7baYiSSqYkEkyXR4vXfmydpmFiXbeCFhxO1Gkfhs0J5MxUru
ldHU3woZQJdwEBZ3lv2F3DfXzVORFH+vcd+uDyDY/WiC7DJ8w3/XdFWSDwLE+01V
CPiwnozmqVQEqBsSFOlVWv6A4tirX8+jThDQmmERlWbIKoxca6xiI4BM6UtmI7a1
STu5Rkm8mybN9vVyUp3sR6rRe2EszWWLbtGLeySI0l/WqNgsnG5nzLhk69iEEn+b
zZLOXWuhF1VGHMgOESItJCmPSZnO1tw8bizsjl04HViwGiHcZa/+VBgjP7jWn2ak
C+3/MRslmJl/9QRryQU0Y39wGWdA3fIERMUp78w1GXI2fzZWYTeom/4fAvnjoKta
Z7rffKn2WZqjnZVPmkehzY5edf3Esnmz2+JAMHEuDcWXsgKjlJhln+e5MOl/gqCP
xzomLwocAKcgZUrUn4n3Q3XUjbF8x07Tr4HbROWt7gw01befILbLdnHQZKaFPcEZ
O1vWwF53mFvGcivJ30LiDuI+sWF+TJG4FOTRcWHLps+Ego6qkoHTAYiIgiymOaND
fC3UFHlstwFywPtAUxgB7y7b6t066cIjl/+J7bUpafXRFcccBHEYEKBGpbqV1kEN
3JYTcEyEesTLNhRD09Ygy34jBlaJ/BYQcGAFwoWVeVQ2+GqUf3bYDR20JYuk4dSD
QPhqMdfnOWysMe4BEZ7XWn2NEutwODk695AQcheRPBB6c83vxAUU1kMqoMI8sR96
0lndWEiM7/pKKF1uu0/0lVsnqMYEWB027IrqZ9hq6UxPCX3G66pRmg2CRJbE4JmF
uYIXGYB0yKMMSYO1CuZvnX6wewqN7+/kg7XBhyo59ETZYlrdY8RcmQ55jUS8vg6A
kSpZgEONzaa0HA+bRoRikxSora1PPESw8HhcIhzA03XIgq/RWO0tCWHwV5LOdJ5q
SPi7GzZrgubIIvganuunGjyEeOMjPu+tywPngb2rHDwumpenBye5SZzse7NP581i
h+oESGRkzWNLW9jPQanTZd+xwQ8jaK5Ps6BOqlCwvVXgL/YsX3mTtxKDta5/uMQZ
CNxQZnWZgYaBAmqtIZT79X7C+u8uIF0dJRMUu0CfR3POkTSvarxd1OZcKLVvTRMd
nT5mOpzytYJVFwGs7GOtZ64m4X4gN9qWX65o+89KZhG2hPZnWZIepsz6UHWpDuDO
5y+Tt6f6EXilfiibc0I6P5LLCksaxg9MroNzyy5+C91HuzvioLSBawFMetEAvQrf
ufRHUDTloPLZNg5M6QsrHRpUOfPJuNRToe7mkADTEYA79vUPkZLB+vNmiJdmZwju
8Lk/xKTIbDrEGeVUe7KCF+BBElXAogUjTxGJLRy84Hb9z95pjHC7UpVBMuuXfrOa
iZtM/kB0ttX3xicxQOL8s1Yhxx/Ukaft6hrrqTgwcilnZobEyAWB/qCfP4BrIaRp
B/uSmjVLLS9fxcXDSmNa/p6+1ZzNKGmZKj5giPpw60taWWZ6KPDSKm+QAN7DyUpd
xDCUPVt3LlqtdD4AdDjDInDxYDlBUmGQ07L7wZbu2RDJHF9tOYM2ukdJUzlBWSvg
w0IOv1kAGqBrsLhyRkYvtiR0b8BRx0UWqji5+6w3ZdpK2PIG0G6UkIbqT8YDjWJD
pyrrgbumkhSCgRbUmjXWHedkMfF5KdcMNX0lKY3tdNu6X65bDjXula9F2RYwOEP7
2RD8wCpvs/xAGpNkl2Gg/RYDyRT39738ePVg7eWxm/JqJhLZkqrR+yid+VBNyWxx
4g2eiKqW7A5WKEYgmfha8BsXuWvDUEV0ZC7uFgrgUwbR/518sP1DR9rwQeZpMPuq
u6gZ+68P0Ow9k2P/QKxKKbWqC4oUAHm2BhlNX+8zN0vZVVI3lUllWP+RA0tCIzfC
bxQunL9AEmq4RzrDygIMz4lKUzvp5ioZquAf+tiE34pfARPQ8aVJl8FoBzBcUi3R
fVMW8kgiGUZeqOgZvrkmzFXaZpcmdbyArn7sYg8wzsganRnADxyMtc9kBSohYibS
m69Q0cWtydzW92fZFHkf3jqr7M43AFZGla8uswX5KZNMxDIPBRdrgjFBuTV33Loq
HOXBy74F8Dxu7Na1Pbhh4D+hy/L2g0d5woDNOLyui3vpKAZMXrH9o/pZEz3yiNIB
/9Hly41C4/vJYptCqj5ze79+SNc5oFweHIADbYZO42Ac5qCCKp71dBZS0YFCetN5
YlIw/7QA8O6XxHrJg17M+XkQYNZAcZCdpMqtvWJyQOMDPIwdCc9u4JejOHNU5/WH
x28FdG7UOOh9thvB3KBcko1fMj7RxemUxjVYdJukaEKPtMMaFiyinG+I3xdHPm0B
d+5BBdck/b7bBp0ZwlP1F2Wlx7DP9AEdcmhAu6+bd1kiKIR+vegf0Daz0eg1wWM9
MR733bgzufp99wTF2vSnYw4haxYyTFY2jUzFazduPFIyKslMQIJpnpYGVvak4rws
gbDY3jD6LtKdbElY4NlWlCLD8Th3hdQUXLWnNwLDbUpKeFX2dp/okwHthyJJ7gE8
yWZEeV9KVe0KAERK6cQ7qRg2UnRlJC37fLJ21PbBNuXXH/GzcRP7uElYgvMXRVYv
ALSV8JBhbPZik70d0qkge18vKNgLs5H+MLS7wRdEjA+GzQzZ6WKv73AyISu2ypKW
dBtvSLrQt/Jz8yA992QzDSJmMeGIU6Sz+m82kY+InFjKKGRp16BtBsHdL+kPzkSd
avfkE7NaeLG4ajL3keocWUKaubrY2054sskzLKrN6vsWjtVnOJte66RB/oxmCAz3
TyaWFspSTjsVE3Ol73BI0pJcAGTUnFEF0Yo04vshvJwWc5yKdhihvr9iU2NIdrev
s4AygHxHb6QuW2MVsmu5DHC0Wtm0z9IUtmqAgLYDhz5lDqqOvi9NwMSfuoUMAvP0
2nK93D2TAopVpEIKlhaEeRTMBu6D1y2YNLwoVivAyXOJA5ZT38cm+r7pzeMKumrq
JruA1FJ4biqCee0EatLQalhfECyo9fruz0jbMdF1ny7vM/pB2s0WBVYFtjm2qeQA
+nuvKdCD+h0hkrebGIsomCTvcrBit13D7q8iKWCs5C0zLsmbvSTJklhK0/h0hvfi
WNMLiEQXh63jowOy2ibdY42dGTv/6BkUYjxCaOt69drhrqfWHfvfcPS+e/6+aOM/
tp+tOFwRMb1p1fZwQDaWaBauR7Ytqe+9YPVLhxzczR7RjkjvfZ5fzDB8chUg49Qm
pSPNIXLyAc1z3EXpdT79pRi3F3gWwc3qonWIljiv8WUBaFpQuXAkXF7mW9PwZkcq
iYmX9xR+KczWuceCkvDB8WpJE2o81n6N8+oyLrZZyNeBpSpT00RnvLg2Ld7BNyAk
bLIsUsCRuYbTEEztM6mVIiAfhrujElIZpOZFkPc5pvKaAD8pBgiRj2RrfBLVNGt+
3HWwf4/ng2Z3TjPVYOqKgG8GjdAtvPWREls0RUrPT0xSKF/NV8uK7q0cq94JKa/B
SqB36YduPs/H3LtjqnbMN+G5Z47oaf+mcxgGlT7AmlMVPjqpOSi8eaBb2ExdDJQH
BzgqXJW12CuqHEpZb64fBU6J9gplWMoeR86utq3FukVxDrRZxBL5MyL8qmh67XWO
9ONWaB7+MeKqrbN8WsRpEfqLAU0hV0RthPsRW2tykj8rQXsN1cmwZclJCRSC38Wl
bwur3HPIy6LWUtojfPyjcENpsRuMFFKKzUU7T9L+vmSyulv01rZU2lNGizaAEuBM
F1uRM+fbyNmfh4JqondWormPra0k4GPAZGIaqScIbc0ZqaYqaTXcVllsdhBnVn2K
kEJ3gGrhSYw090lM67pFdrkzGGdYQo86tP2I8PK+KDOw0FTaj5ENfjsJnCnO3+bq
kKq+8T1d40eompsKDyWSh9LB8jcT7uzSEw/iDi/pmkFiqI+wP45OzSatTRpurz8N
sbR+z/SLwdh70bE1QWJJeWq/+QegbD8Vc3aA8tJG2y6qYsgpE1h4L/36bkG27rZH
4v4nremS/FAsbV5TzFN0oayP+E74BgAx2e7q7yoEooqUw1PNbkh280YKlt8Yuzh5
oMdaqeytfEDtpmPqjX1WKSe6ctUB7iNMs3akyj3NISAfdD+KjwVmLM9KBIP8fhS3
se7iZuCxI8fomn5qh9IljX/z+rZVleQ3FbtOWINZ66j49sr/eHnBqcuY7+R0Y11S
lkv2Xv/TKx6R2mC4rwe+S1Oxo6EcnjYD9QQhL/guT0ig8nyscpce6Rdgniofz3aI
9rJ830Y2doNSPGzbPkBgrQQv0tNABsIY5NPXPkP6A8gH11ySNKaCRa4v9f+g6PGj
L1Etb0P4WtzrzMzbkMDt3PMykS8dm/6r9tOFgHT3Fya+Iohc4crStOMjr7x9Fqtn
Tl9zyZo5kArV7Il73uNxScwIW9cPzMxl3dkGIPEZlmKa1OKDzT8kyQGAhyqZySb2
TeyWDrkD+9buKOrQDivSCPq5g/wseLGuinFgpYJpX7GdMStvVstD9fdLFqCHHL2c
jOjjfgSqZ4wyvh4CzZl6CEs2Os//iWuPC3i6bIkpik9gbbDW08U++y99sDfggWl4
f6u0JgiZAD0GhuV2qUgi+gx1mpyixEHFw7dlnXBISzijBxuV5qJ8M5i+0A/KBJiy
kxMzp4RYzlb+ac7+iAUzbdXJmQx9PNLeaAy7g64BbTrU4NNQGRZtjHw+TKrueRVd
OB6kPU7jSsCbhi6DSkVNU4qbxqrLN8Dld2gybZvM/Gzmk5RvRithgdnIsLKkDO6P
Hq1hHjNW68oMSm7uEYI/LV0QKs2yTLVHAitgSeJvmjYml6qe9gD8DCYwn0m+UqcC
Cyz0cgb47T667jfBahjEhYtWDER5ooaGN7FOn006kvRpy6xwZzOQ3VdVSsHFuguN
wlt9/DOHbySDRl8eB2avu9HwyBhkHqurJVZlZ02E2oHcARQWkgXpEhz3f5ROZtPA
3RwJ7igLjDS/fewctL4cq+BLpJRF5yuKhkiWqE8Hn9S8+4KoyR/oC4n5YtmTEDPY
T8oIy7rxDBb+BMTwFNXU3p+O7ZjCdoyGiLxyRBtZweOhUkfxhcf/5Pz5V4DdN9BO
dL2TdrLPSRnmSGqX4jnMZw2GAgoWqMxQgzD/BD7+szJms3lQxnaBSfClK++HsWZN
rLsxabBkW2ngFWE0/fbnggDo/h/R6+j35hawBPvf50q3Gl2YmMg7Ynf2/a0P1tZs
zIk+wXVcADMrNkqyCpbYLd/P4SNWhit0Y/MRe0Adtbta7jwb0w467f4COKwxlgUx
TJVtrpV4gs/3Ecj5uIEzMgnu4ipfFYlQc9R4wGpGKJEx3HQrr2Dc9Hq/sUuSy/1Q
MIhMFyH2Qv5ZrqXR7qT3dkj4c1rBd8TXF6gm18WrTXeHid9hi123X2jRv3z0UlrV
oTVAYmP+UP5ryzzAdFQMFCL1YByoBViLy7jDaPbhniyQillPiaCvXwkeTWqg3Ezl
dVWe075Kz/miSyw87aZnbs7UyXkcLFTifzqAc/mSTClyYkFFCr23y/3WtI77b2Rp
GG2blQnvR22GH572zt/Jp2ZE7koA6rG/sgF3dja91wOTp8rO1jVln617fHJDLsxj
sWSSmMjGVtFatj9KR+xh8PbO2zwuBD+8JNncCwSbq5qFSOoKD5Kesqm5zIbimz6c
p/rj4PDqcgxAdEjrSZYWdLKs9lVr9c90vUPck+OfGZp2o/eBctBO2o1R8WAPg8Zc
KKub2mjdsvobyPWOZ6ncUlByD6DvJnavnFAYumNa7REDbLjphxg/udk3TQs4a5oG
edj2VZXzsQxtezjTqVNCpi62BuMRCbZKwePAYde6G/Cc60daxAAH9sfxLun5kJtG
9LdP/jGjetyNsh8sUTOdoLOP8Rkwz3YQPzzgpdchqKNwxzTtDIArk0xMPfeiR3cT
r+o8xwR21kIBnZWjcFzLVnozj+4GJ/l1ewy8Of7NVVbz0kz3P+Ns413w8MZxvaiB
rd6eH+gB8K4vR0n0HlCQClGOEtBsJ4f+nihil06qqratpP/vTei8XBbOn9AOeP1a
smJxoB5E/IQrMBucOZNLpdYO9P3Ydabrm72qxJI3bphWP+dW/jybsCyt1uQI3c3y
2hNwXKFE3Hnt8Se8c+iNUysfdVXKSoMvPttU2IcHoW49YcZzhN9Z+xb8SH69P7oH
AkYRoDYB0S6GQiADVV1uXfDm2e0kLjEagn9Vo1jHAhh+Tt7B7wEMdu8KRMruY252
fxtmiJVCgabl55Tcdqdepj/poeaiyLus0D6h28Z5TH0YYFgh10m8RZkof3r0M3y+
UXp+K8p2qmLF1sxoQIcXk2hPspbQC/CRPQKdeT6qApWLoJc3ro67kNmTJkJ83o+f
vLkKgzICj/xEY//EW9sQWaZKS41/2bxBuhrBTkb24MKDZ/wsT4+BqyMHzoYroKmr
UNb6jggxbHN1MjDl5XhTGU5m3fNqMd/1C7wFEsiq/ceON8ZzqFQvK6vHvDE4/s1y
wBgC9H3TiNkwkGEIT2G2aGIWoBtJSd5CU3jVfUMccXMkrKZ5gqESxdmyCju7IIF3
f/oJpRudLV4wOu6F37IveggQ2bVSdX8i6Nx8iKqC4u5v/pCzP2F6aKrrNNyYeJH2
hab4ica63SJZ+M0Ueo/f3oAidJMKSgqip0EJgN1ergyrkBlV+g+4lrGlUyGI8VJW
UFgBI1PSFNajtLWR+Pc2NPdhHZh+wtHw9ZwrNLzYmNU3Edebq3tuivIuPiwcZhjK
IhusbPkzw0XpOtO+M0DCj7wk//NyhoExGMqFt6twMH/is2OtTgT5gFEcwbLvxoWy
NuWGO0KK8sjIKyqJ/SHMDo6ZhVYCfg7h2Lw4uy0l6JZu8a9lD0keRnwCmGhIEkgX
rkyMZaYBCzGLvCad2JjMnuiDSrf3M0kGCS39wx1U94K/+3Ifl48xZEBrwA3HMswp
Yye3XmU8pf8mQo6tdB+S3cu+6AS1lBrDAAW1M2/ykiTdeIAVjwRYTk+u5aDbp8lv
PHIq8/zMFTKUcwYmwWJcEVrEJHKE+2oC+XntGusBRbgdgmlmWb6oYT9Op+KBDWTO
5qv8di99KrKogcu5vTRy9PkEMHskCZMOEJLgO5MjOH3XvaosdV1UuHD6N1jhfpmp
+dxhreliqe+YiwMWVF2qKQHnUm8bqhzOzldeTt5v7muAA5jS0UG+x4CDJKpKqDV3
xI6Fv/A+140l6OUjolOiznVhZ9rnnxiu1OUVy/kK33DD6JqBWuGvu5748tsXAunr
h2fhVp6Rmc6LE8N2X1o5xSth/NmkwGLzKhoicSs+IzzqCRDQWSME3hQr7KN9Mr7+
/ZBF9+d0VEGvjso7CXM1aLlhadzGZIaqAA0BF408UgubUklcsqU0xQ7h+ApBkNOK
L14MkZqb9KbjgWD1SCVztJMmcGJxthRmw7dp1iXJMPqzYqDkxi1Ea+L2LN/UC3tj
9YzUcvpQKnOzUTsQzijCa7ypY25MwTM7iXG2kzKvh0SxdbEbI9qMSJh4famrO1MK
gv3Cm6VUatIYBuT/8ik/2883zCJZYJNEproxOjX9+lTwILo0W3wYfRWwlJmB96Oj
ZeZlpF1Osp8KQJ548/DXXTi3eSFHtwiFRJXQXRlwyDUoE0Hr3n/p9v9miv2VF2xK
e+058VNPMo2/rWPsEeDvA0yYJjO8Ys02TnNnJx/EBmD8mlyx0IyoJrJdHQ9A2FZW
coJwIs+oarY2Vom/I5f8532IUEbFwMGfm1oYVbiy7+VvXP4/3yridQa9ZI0Hi+UP
CnLsRCgVWlf7I5wJojSRMOIdlBDkCQEr+MI7c7rWXDKlmqpRxVm0ob6n99c3dKPk
DahJHZ8qCa9t+Z5lGRjMp8XjWAnwIUU4kI/BN7gKm+H0lt7prEYwFWhYdzzSekln
8aizAZbxyHecOygaytlUAmJoaWsynN89E+Nv6Gi8WeDTbPaZKfkY7oI8fH4OSFcO
On9sC6EhShNZRamiJVKhlO/iBKuXmgbtvmijW6ftZ4iiVwhYT7tFzTgRKR6FQHfs
4+iNkCfJu8FNILe4dFNKupu2pp/gUY4nVKVOa6UMBAMrW0L2OoR8hs6mJpE5FetS
h0L5PFHSWgaio4XWuWNCKe/6sIPd17n5rOeLPDlYWVzHlpXVwrsAbasUHrdx81Eu
bx/u1np6q919lhAvPUWgTG26YGHh+itR+UFXyfLz4iv1SEOqflu99cDNF/ZRUftu
UAkpK9FCKf9ckE9/mubD37bh50gwpUYrvTEyfUQsBBra+MAlBGyNPx9mn443UrBx
PLK6a+5I2MTSI/Ifw3l7XfWh+7YGTvJNSsjoKFDMS6+4fFn4+BNv/ELS0Q59g8Rm
0n1yN1NV5wEiO2RGJCKNypathbGEV3tbUCMweZVjavK0/ed3B6uuxMCVe0PA9xiF
6Y46/cTJN89F5FuJtc2CUGhHvhSPvtaIHmxBwkcvMhlxyfBtNKB6pZccdm3cbvLj
kJ3clSTqjuDbxm9KLj3Uqk6K2gvJjZ04safVhnEMMYdI4mBpkTIzKDLoXq0ONdjF
R3ZFO6EccwNYjUNzVrfGwLFSOim+2Np7XLDn1rIrK2DmWGF/zmjyYviLvSSJSgqr
hsgyN47uCyDwDowLO4BjFJlY3ag9OiUJsZqOVm2kO2n8Sq/0oS6fVCoyUxzwSD6w
qZdM0PSvgidsyobM1/akhNaRm5IKqZIQFp2Lz+sH2DeWM192PNyJdTMWW+4ciJqE
9pBPmJQmBlXkmJfrY7Y+vpYt3I8gLOUsLX6OfxbYbh10Qrdxei5PqGYdEv/DnPiE
XDBsoeWB8lBVZNrxs7Bj3U0GUxK0hLLrSkobxC0zz9TUmzGhjPXY3BLEL+9JMvLx
eb5dk7vo+hrFIhzuw3vsUrjkD/QUMsPc4t4AAUWcQQxfZ/hoDEe06dbjXlnINKxL
1yqQ4sVQDQkPV1pquJtAYMnFWLIWjUuSWVN6xq1R8+8zZwGuQ3mDexbACIC/5lQs
xhR4mbsFikUli4QbKK2bxtZiUMwtsRJGQhP0SWr3VBRTNN3O6vT2VyAiPSSX1IAp
xSmhFEHDet14jsIDZtSCD+/s8I1l5S/StbsTeqjn8wGLYTzvfvejhbw56kYBDPp8
Dm4DYR/MWzFQaC4loVFr5Y/+xk/JIuBFMBK/7A+wogKf6M3ZQkn65kLCIStAlw81
JQSDNZlUDVYMPxKPVo7xi63sS2HeLCf9UvrCsSjMJlcInyERZdlJBdypTBvt1dqx
vUq9f5utBH+1iVfNJ2/XbINmeTGyOG/C1oOtxPKvK/1AgrIG6tJdAnXVdJlNqXPL
lpxpj/NZUtEHCGz2Z9ynEVqZuA02AzIGxMfGwTQD4OgKNM6MW9E6e5qjvHGIoeWb
gh18iMjM9uIHhmVoG1KPH6q2cGBybO/VcGhhFJeJlMsJIHl3+G1++dw8qNoTQxD3
wcZPVIha8xhFAbmB9j2P1LCCmNf3bPnHTWhDoiDNBG/GUrf7holcE/mpZt9Xgwm/
nBjijn5LjtVewzjgZc9lNUAZaIQ6+a4WEM99sPmhpGx3U4HtbweY7TC9DlK5UGS7
Qqhg5PkChtVKnjySWZrvn79FYYpLCsMdJpWKkEqXi2wCeAsjzmkFXbwWXFFVTz4s
U93OJtzg6MvWAYNipFRTkWMjR8NzPPM8ObttckdjmYY3oyLzu7YYh5Mn3k8rHhkb
+ozGumu1dznIt56MKV/g04xV6PALCa8EJ2NikcAFjoK9Q5N+qBaVxOqLCz8RBdmN
Wp061cRMtIvbPu8XpNvUyMtgGjYQ22/tGNpVPxjujOabKCWs58XrL8iKSISk0OOt
xBE/HU7QSzWISY6Ol7+lZ4FLBQLfZFVWysFjk05VTXaX/2y9VaNNXfi1tPc0X1vN
yGbN/Q0cnmUBktcvKYhSJ+uNL8sqSXcjpz/lvPk8wEZaFHKJT32dpH8mxr64ejLD
MgdvRIE40LkxLKU3yMMnOD0/0OTrQ5EYDeCVFL2hQixeXCvaRoJzHOYjlwsgxQ0f
uWPZNtiWH6dwSv846qYQ/0qEKJInhA4VCCr81EUrmz5YXUU0XS0e/UnwtfvYeU9I
3EWBqhd1f8RAN/qCFRzM7M9sVq1WfFNowJxUDgiJyC1E3h9FrD2IWemP6vINvv3A
OMLvaPZBnvtx+8MjzaFT1+SscTXwFijV5o7eTXW5tfF2dxQCpBjDpqQHewARDh9Z
susIyDdTjIoJ9/M8Hdp6iuRjbdYU3z+UVmflr5hWdLiBsMkcJWnrLNDMWNyIfvbv
ORuxToJjI2H0pm2tq6DK92yYXmszD7jkBMpP9VH/nFqoDoWPcWy3w4sMG3RoT/2k
vU/kP0zFs/fCiJfWXXIxI0m6nSPKWlx+LcDty+ha309zAzBnTaUXmzgZMdvwninP
gU8QHXQyjgjlXSeOCvG3txBAra1z4tnzEhNe98efXVME8+z2XqMeKZJXQfS0luut
bJYIR3lRz7Vbf6DucEexkbIH1XHuCHD1HV3NCF3MwS5Pz4jskxqG8fDiuB8EXdT9
CY2Oy1oUaqPgRW4vajMrzHrqm4qaSEbAIisPEI9Pghk/vMpgejlyOUjjkb7zVM8n
xYtYHAx+RrEVDyiokeCLdOqRH4XNXIi3ZbeDuZ/6Y9i94HgDjqHjGmFvtYCxY3Gu
kzyR8bHVRd8qt8BTdAUhbcegsa+6TUMsSTdCPIavBkJnv764zwQ6By9O+wAvf1Nz
xgbElMp0EGSnfE0ezwEsL2MGPOuc+IXsYWwljtIrUfsxp/BbNOCXBh+pds+q+Dqc
xNUmnAWpLKyF2lsFI0oJoCWOnFKTEMUvIlfUmIgIktPvOkbhnosSxsa551kZZGK0
Peb21yN8qfAXV/pABdkf3EdLoosukalX8qrDHHMlwzHx4di1OOxu2beiChOYrrj3
MJhvRY9+91s6mCKiRYp3XXhIUXkQ3LrQ6nJn4yq9tLLiFYvIBPr3pSILix1/6LWg
5iQg7A5AzJvTQuEBr7H1uXpzB0B8mvI4BzAtU8O7yEz00W7u9vW3VlJrQenUnFgt
e3xzDyzlMS5sal+kmQ4AEZ21/kFweq1mFn/g5ZJq2NLcqlsf2DezjHF64S9P4brg
5RgfHI8J33NxDQZ2zWLZDHrffdMXfof1cSfFnEWQeCC21Q8faco0+eL8A528OvcJ
+jp8J9CSRZnbfliSgoNdgT3ZevGlXOpfkZYFAR9DFFCfeYZy6CmJut2JQ39q6SrU
uamVx4c2oYOXaJ+SXcUi4vlAEuyUs19CAKbg39SbK85AlX2NIUGvo4ue6BEfUJLq
qIOLYl6HVadnrcglsICmX6L/sR+CAJw/nFYFCxyWXo3zm7Dw/ARPZB3aiuYw/e5X
DwpPmhULX3DNadlk9WxzGklWDmze+O1/i2Nr2bUazf8tK8P2QlSd2bFXxdJE4DSH
RqpsIgPpk1RDiuz91EM8nNg0tmV+wzLTx+1vc0n4ovD6SddgQWwgMQBCS7aM8wxq
RJKO25V315PYymGsHC1gP6hvALbqeG8wwHjZNTbaXRyFsAezlTjVSIRqsZk4eL9U
YUW5U0ZMaL6iUZjJW7ES72LdPtRnG1QTMCuWoJwhLGlfhz0xufKTRJPjM+9NAqgF
DmJkCQkwLjHXl7UGNhaQXbXIKNLX5RsP1a7N3thoghdXJgauiRunVeyW9tZIgWn9
jCG1sMe3ClQqCrFBHmU1O2NtvyiPacce/VqVK6I86PSuvozWdCFrj9bAKlMx5w0M
hGPC4vYFOiq6jAbRJjf+WvQWvzocN2JsWFOrjLtBq3L2GsQMZ7xV8YwpzjuLHClN
tXFtRnfiIOzsZO4uw08FUSczFTBDp9kcuTK1G24D2Anhhbv1jxbW1ei52uVA/Mnu
3H40V6DdcGsxaywCr5sccXgKyAvTmkK2yd95aDZt/jxDXDtpkKyguwirKYqQfERh
4FEqXjULloXVTtUIOXYxN8goPFlwnOhCsKsXnRJFGRDEbwroK+NSp/tHyogg53Cm
vYYY6ELC6GgOLwvvzrLUEPtCHoT/7EfUEe7Rfc0NhluCPE4zwaI2mvAhnzw64D+Z
v2wctAb3eReHd4JCXHbkOkCxTFNkvhKirew6JFQYIUzWPtF/pT5HeMGQQ6z3Ig16
jwbLPEtzfzwtjb69tqok5h8f5D3lyvO844IXJ4VShOYNjSeN+QEyZiXDrfQIT7JJ
wenzjUACr4IYBMPM56P5xSw7mgVALey9GHFecIAd0i3gmkhBwz7karVOx7GRXHAH
5FRMbhNEAg9myaFeqfyfkYdsq6QjVwVn0VDFTWM+dRV9ABpmAyGBTj6C2bonACue
zYxKhM9xjsOMkyyUatpdntZJrKB8t7TIHibLn0iuJCH37HwnpU29EW0riztF4+xh
41LZQvUAI+w28jGeCKJ/ac68hfecbgdnO4x/Y1E7wwVwBhaFEgiPOKTNR/Z9eppc
V/Fz0jS+a5fSC2/CuLdNpa5AnSg2XA+YLmN7oolEeJUUkQM4rTZD5WsWfL4w5oST
nWP189qXWcT8NnoOD92vA/nnxHzutCWU078BIkDiAl0t6Ddh4+TPreISrQiIsENg
tfsgdjHsSH6wXVME79rewtEonAf1usDmDMJ5HVX2/fApgrgO/P2Fx/NP2R4UHt+D
y6TydEtZr02ExGDY9UjWVYJwdINFGBJV7mSpq6jLqo+xT/cweYaMzE0oX+oWsaXL
QS/94KBZt13OfyS5nxQOF/hny5dlt78vHZmg8jrPRBwnVGlkrjXaD275kHIk2UXQ
ZwiuwTj5ob614VoD6Ncf+ISYZnkyhh5JyV7FOGOIOXyuab26T9jG4kT3nBsQVq+q
rZJYckl2T+VsZ17a+c5vEGL5PFfhoBLx1cr7QsHjCPB81B8HIy2saiTW+hGwSsHX
U9Oti12nJBSOqL7xFUb6fe4ziIIiJQIlyUkyV1TZU6oEfWEiHB4RbuEBoS0iPB8v
L64hfQpZQXiAiGOvP6zGTzm+FY8+gpdwUqXYgzW35f4kYNiENL+jmqAaNywzdtMx
JAOj5aQby2RRU7kfVHsEfrcxCsGpS0bRgZe2pwV8iFbCMG+jY8yYns6uBodXOCdd
L1wUAAEid9TkxnuPp6bcAkKpKog8zb6Oc4ZcnW2Mhz7Lx3AKY090Oq0c1K7/Wf1N
PxswLo+LksqQ6pfpCUDl56nmLctOgYtICMnnhhFe8bRatrBmfB7B5Q1C4itYdsHT
PdSJ5+VCSsFsY6WLSwmRDhwluz1qB8eN152X8TSayIPWWxSv84HSv/lS60N5jOVD
b3bMoBM7uqXqsK5K1jwlzyYEOe2R/A4F38Th3oPqOFlpVNfYLnH2n7OjQLDmwFwR
+WTVAIiEgXameq4FLPiIuC17oP8bvu40ZMC+KNIJBmBGjefbTeak/DMLHBMSIMJl
QM84xfdwjb9Socvz/Wdlzh+T5g8Qb/8igJ3RgN8vCSUPC4Uz63G2HrAOBFwvUz1v
TA7oTVzbyUnWVOxDTYm9ShWmWHJmEvKUGQQTfjrUnCAHweIERQi7S4KF3xYMs83S
Ynn42kaT2Z98iW01y/gTDagZfAuVACu7MMmItLMP3PAhKZiAQLPh7VwfKlktacxY
Rk2jInflfm7pCPYcon14sNwK7aAdE7iD7km4avu1EYeaeY9WTtmRz55PJoZNUehc
4A2jKwl+tJAiyBle2QgiQCh1Wl9iCYy6OFfIGfuScaVEYMXxOe/jZnQYAMLSbtBo
Ri3Z04EuLJqkHOcFIWro+C4Gyr6DssJd90mVuenG1o4eiSMs0CrF+zxnnmMvQLaF
/O8Ib6CTNDFKxsXNVOOAXzk+H8jt28l7LOXM+w/n229OoHpQEGbXD7JTelQTH0vI
B8w2f2vtk9LT9L0etqsf9CPLfq3l5Z8MAleIQWlOYjeCkSmeCR7v8IEwkqYil0QO
1rnbV+MJZHT1LubJkK+Q0IlP1JnmELfZV3Cu2YzpcdGHxbbI0zZobwfB6oEI8ruZ
Ns6yP880IamwDm0NAMkiB84nyEcIjbyaX4xju5bIEvpL5i8BEX5TQZkK0RJZmWCI
cGK8skTauiioV2KvLmHDQ5BSnTOB1AxYdh7RmtILhyFCOyebkO+VeFduLDqad7Ui
TO7158gPuWIGGQ54fiixHxDppno2v5EfYqg7A8Cotn/i5ZjDKuKlanteYaEfRqqB
2a/bOE5bxj0whMTMcaTNa9+dbFSMHz3KXWDXaCHtEuv0ac3Nrlonq2Ouf3oC7nNn
1B+AQFq6ZmIb8j3SvtwLYJEA25wMj8pTW96WZWMOEaqKVP4Jy5KBBkuEQPPupB5S
MvYMGuTbl0tldLFx/eLRCKBZEma1riE9D9Ph8+aJX+eP22kwzyjx6zcDI6dN2E7I
48dSW7tg6Ryz/4On1th8ZIK5iIH9mSEMaZD7HEZbIkdgxctmIfI9Tv/RyONdTECl
dSZusJL6a1YYab6gK9JFu6SDqkoVmBSv6B9zlnNtdfwzN/cxk4C4VdAHlBRxm/gR
eGNt/NvUieNXvaG8/Ol+Oi5EmRcodLZhLYnQ4HdFsqjXIN2WBkKhZnKn9uVB79zC
NYQbxzTiIOFcJGylD3BhEbNA4KJRiYgcQDIyupi/+wQ2+fa22mhr6BOU/bPeiTFO
w85nGuJvL2S8SreN7M1AE0RMYMqFd4PBZn+KW+0oWXHv9s6IU3cLjOQibtReNtV+
8d90McZt5XZVmqR5zrVIm/CYMnKm7AMBbxazVcSlQ/L2mDIRK62WyQSf5vxaA8Fo
0zMN+1rST9KG9H0u7Eaw221vRKq2zkW/sDsTWI5hA/y3nDKIlMfGoMLkrHWC7ks4
jtYzJJnPBCHRYxhnJGAb27v1Hdsjvpfaxg5J3/taeMJyjPMQ4M7ByFpbCDgpkXtH
MQCk7FRwOZziRPJpZro8DxDSQ0fHvAr0snna6beqMrDgvV5jCNpT4A46+AULKj4H
7YHRxvZmnJO9z9J4CbyEPVmqMBKzA2NhwR8VnocQg52I1imQl+4UcCVZpZV1ftkl
8LftDljtP+Y770GsIRdPNUdszx9Wc6LvMBlCEZtekXrfd0SDJlmbxdC+ycf4/Yt4
Ogf2YLgTx2/v1ZRMEQhS854MV2IFB4HpH43Vpax5PqcwCR8oND4POJknGPmcnPzG
ykGAhlQCRARs8BK+yDEfMrKfNpbNJJKW1kLJx75EfivVMwpbBYxuosPL6zvDEFbO
ecy2Z8Q7liN+DOLDojpt6HDtuz1FirF3hqIvdPoyKi8qu7q1YBTalXoBxoe62D/2
llxbgAiFmeonu4aTFVGAJXtvCk2F3pW/DTrarDXJv15xNAZKzW1vIAwaPyOqtG6V
9Dn2N4EQOI39LPqmacHnoKpVsKJElBzgGNy2BJDAXdTRlImleyVZLD1t6kZSJFgb
pPLwtpDdW+0UoVqSUr+nIK3bshJEEgGi/QKHU90zuIIPNoWs7rodJTbOZ+MSBHTF
eR2DZKTqz7wmKN+EeALXyn4kpBujzJM0KlvwYGGqw2MDMXUSkzYEH2reacjnfQEB
vwral1cpjHloBs6DvluOPBjI0SU2fHdlupQYJ2O2Du/DpfD2oJzCkAfS98Do+Nbg
4UkaGqsUuGrg2h1R52BCPAa5o8C99Qliv9lU2iYVjU7qEmrPs1NC5C7G4k8ITNxc
n1UAlNupiksD1urFnizlKKcDWVM+LoXGgzJz3iHBhG8rns8414tkUZtSFkMibS/O
hPMnFmjSuXoTyEglQdYWoRvzBcvvyZgmf/+M0+Wbi0lmvrkiNlbtviy2mzfP0HP2
l1cLduCqYlETSUqwUHXt92+zLcl/UOhCXpX5Of2z6sxOiZa/DuUycKqzk5hoGY3f
mOSH76Hp/DpzyZO+gH7hPALgj6Hm/T5a0NUAqwPgO9l53LYTKIdVlMYELpi8xa3f
kbCovTK68UUQfX9TIAlCB30U0lGoDDMlERjleDpBab7AiQ0p+IajkqeusvwNlok3
g9u0W57/Ekek3Zgq7LhRZyG67xN8kr2830p0hZlzocg4RgLwDfltGDLTKCmlQcfF
rdbBza4QFUk8bbo+V453cOsSOhBfBkofQeSyOen3rQP6TCUilxElde+DPrh7kw04
jSUKHe7vigQwwIZZGS1HkdXcgUMM/ZaP7JhpIErgpkPNOdhuvcJPX83xTVknYjAK
qWP7EO7zCR6IPvh82xyzyEu0GosZ00XSjcX0f4D5MqoBcjBfa+tgIdW2h6jEipQP
Zq5g8UhO0izMpSTfjwGGUQiqCMt2yydAIy3BKcKWxwVGSL82kwza8JjkESKOJv0H
jpKtEtMrEDKBjFSrZeVH6/c/phTqwHrlpEX9gTySIBkXacHU359mV4d4YfDBZ3MW
MB5JbQ5I0lbSu6ebjrPX9zKHHBDjAIPtZMF5ubmBgt1VXSWdBnKqc/tLqqnbyBu2
ivVApKjReaKKhNEiJ8lSo5yh8Ja514fBswUz1BSm/YDmD7SFrsKCnF+qYZeRMecB
3hENYv3ZNIhv2Wr2+bAhAcJTDjepgdRMBs9TMkGTXn9nFjYTa1heM2aDiLTmD6x4
AKqf3sb4S3vBWSpeDAyUNYa2gXUsbghBWhzCQnTtjtkkqWo45T/w4POZn2vZ2p/v
+YLvRaAayVNvcM267oFKB/swBL26VJph5FMnq3SOH/hv/7qLUW2imhwgDqQ25x+5
+89Stev8aj/LdSsRJHhtIO1TFkJt8D/tBmkztULgkBBKoDehEMBI6Mp2E2jg/wCq
Ctnq/5X8xvu4Tjgl0e2naiktw6oIz59pvLFxtSPmx7pdLVdN90XXEIcP+aWktH3I
qdqsi/ksuDhRYuw/FrT6jpmBBl6t8zQ+N+t6rrXSst55s9BBoDzaYPC/Xz2Oa9ey
xZZUmP03cEqaNJzYe2wbpxdNBlpC5wvYXCkeWTYhCpoCIneRG89DXkrnpbEp90zr
38927USzlWEx7b7zjdr83D31jkOoV4QufoGbEls2rwyRbM6vXp8yW+uxOlBRKYpW
VOCFIH6tx+oFfGji1UNNOMmFQDCvi+P5U30OsNeX3H8LuAfJh7SpqlcMjVZwvqr2
nSoBNES5JWdVJQtBSbVh0v6n+27SVmXutL6dNip7P1FnjCCqGVLCYGVLLS6f8Slz
wvgSKx9Ry8AOOKZrEwluRZOcYgNTP2w6uSTXdHqrsrGQHgPTIgwmSqOMZaGB/VG4
By80LIzyO1vZovjZILXbOszmoLhHzUVIGD0fW4xX965AC2T7chvMXyUIs2zmVpvc
0UN+Zq5Y78sYlqA5+xJMKrx1maJwnZB5bS6MacXlI54U6z052Adl0xQe7e3XDGc2
42jrHen9L8k0HEMN1stNnKH7IaGU9dEIP3tcJ8HYQrN4ZFnsk2l2AWqklw+IK5wH
vpQWcYfmWqBfn+EPFx0ft5rM8afuukgxrphsyPq4PUkq0lZXTksgvA/KeTT+7ZaX
q7aqKEddmTDhcxtOYUZkyy7KuFsOvWDrmErWD8XK5E2QjWJMmn0eR2bSTcbGcG2N
5JHWxPm3wWm+AZcno1jERK0B4+GthhGAmRFNEEy+mof2MxLEwg5FSuYGh76C9Kk2
7NpCdVddShAZQvJLY41pycIdu+ClhQw95wBOZHljJdnPrrCsJ8V6ACs9MF89qd+D
oqsr/abmQRUwRO9Ek5TgzTLD8vKTywVQE0jtv0830NzJqHZq62zoonHeJnnQGQl2
Qes97ndybgDY+aZXYaSWvJRw8RQFbOcI4LxNZHfbZkpV7w1IeHRzk9upguMLZC9G
Cw70iK0QHCqsA/BUkLUALfnp/sSgqLHMdut+i7pKF4/h4WcqiH88tQzlGtW+Mu1X
o824fI1JuWdUxCL+A5R+h0RpGby4JWqDPXvkg9SdORzxq4E+FOq//0BPw/Y9hGCu
m3A0Ey7Gdygk5gwx1EJrH0gem96NpxEjLWpaek8Qn+XGkxQws+ztyw2eD2syN4p1
jBtTsnvt8Ec4yY6G3uRGYbYFmkpdRWj2ma/VnnGUuKm2xuX6w77Sly2NiG2EdEEG
mlERN9iLpGLpGZPUGJsSUqHLxusfDWZZwxicUCoGnwEEk7Lol5OgMn1+eSkyBSaC
zpuJxx35LonsRGKVbS/F0E/OTXf0ZSFHjCZ0PDWkvHJA5ZeHKMfU5odduDoxn+yG
Qv97Gl1ueP0BpGr8cIe9czAj0C+uOkIelR5NnRIMVqqHlQyd/1coVJ868/QPSKNf
xbTC3k8utD+oBO6paDAvTral69bmFkQnQQTocdbdzFSCAVj7b2dsGaLGA/8uIjsO
6WKtLfn1p3DJwUfbwUFSf3wGn+we5XS3XgUcKU1QpD7X40Qj0x9fsYW9qMdVXuQA
9amJwb+45YL2UAr4gAZixJT17bUiGQ+t5VNKLQQGYy46Yy++G6QA9JkmDUd+NcNY
X4EiuUxH3/C5bS4yBJ42BeO6056bVmDBAgq8jHboRDkxNDbTU1ySuKVVhNcluMxg
JEQDFbYA4P6uidh2zBy3UtJufz0s6vclEEVrIWDHyNLY/zTWyph2UDT78FzSJL2m
mNoIXnMsYuMR9B4xuTm1kXTGeJ31YZf7n7LlE/JpjBEsVvZwkxVnUCVX6bo4FNZ3
P1NNHcK9hdYHOCQcE0V1nwUKQr6bzSY1QUc1X9eflBcrg7jVF0f8TRe2FsIW5C/g
6hjIser6TXWe7ITEWS01hmXg9VRW0OgQ/CA22OpGhAKgY3EGjZSaOJ0KwprKxzIw
X7ZGYSJpBl+A9s6t0aFnV8W3zxEvw21bPJNAXbdsrgFtgZWQtSPMIm8vg8V9/jiB
pdlHgeIhyEMGGBnZYB/2rTYTZUjwICESuxIIOXuU3LRC1h+OVwbtgNVg8mpbFtPb
4fK3FudxqZ9qFUWc8D81WclQM3+7dDum5/At7MiR6Ws5NNPWAQ8POb7T+ISsm+Q2
x0J1m5WJjjb90BSquHPu+yU63BHo7b7kXRk+fk7xG+DattP0T4u9jY3eJ+yhYzIz
rRD7hmX8rTaFffvBbpHtdZ0TpNRQxmMYO0PiTAnUi9DXEYy3271uiPSYXC13i1sj
7Q9jagOjmAr8oLt6mrfzYfl5dnSNMYhUMP7e/09wLAge4hncmH98RxMkkhLyuSsw
gf07ShjBJFSyBJ+OCYGvMTAv/V4PvjSpw0dZLB4IVyX8rJN69zyVkRPPqPk8wcSR
AZvNX5X0Z88EE1i8hC1l7utVJF3wkWxb0hsZAtAuzOJHqbDiosWUl3+UAxsCD8mr
GlQm6vpMn60eVVOT+ey0YF0hnjOWS074UwNw7eeX5qivrL36/15ZEhUwxxD1jxLP
voJBtevtmmkX3RT2huj1Kl/3fyDrm5WEapzyjjA8xcKXGBI8c00q2x58EXwKHaK9
9LEmD1Z3HJKGJRgY11Wt0OyMxDwbr/0S74nozKInJZesmt1xp8oi02qFlLqVDzkL
05ye/7feUYCl7vJ6kt3jo+8l1l9BNmpQxsVS0S6Kl3FeC8yUUrha+03n6wslKCgK
A7sMDKErH8g+3g8+aiBcHO7PV5/iT1ciPGW5ipktOmG6RcRKxlgksW1OvjSZwkML
aTgLwUGARir3VQQ4GAep6kfSNDAaXnBV3la7/3WgW4L1rbcLJq+/TXyidsbqWNwl
6byEVojbzftUC9udrPuw6hCwcvwXdu8ndMnZG2Y4pRr56CDSqyW2mr1JF2ZQhz+g
9FDVdFpLiF7qZyOcSHbI9y27DAFaIEJmwIr8BiLw4F1NxhN9Ju4roD42/GZUJajN
qSSbxHaHmU8xMWb+BxwFtxYGLqT5QUu8twmwh6sTQi43oegYCkYVhl//7PvLy/G+
BMZy9LaxyktFdt4/fu+UbWtSEYZ2jKS2TJ175Y/e609YfF5D/n77dR93yhGbJFY4
uAKym/Ulng1UTdtK8JfbWR4nA1NBJv4zU/NVZxhY+zLRqduFHTTnPkdwP/IRCKgN
9oJzdiurXwQ56V4b6Y42AHmVKR7vQPdFbOam/Gr0JWEsCJzZgR2VN/WLzmzi9/Tu
JbILBdiwlHs1KWFcd6oIKzgNlpXObs9vnQE4ml9IkME03fVPJXsz16VKQZDbGz8D
EmfvAt2uYOnKgDhe82kzhHwRN/0w6dWrUKH/S8PajNQ04mKXrEHmvKqQKrF5ZCyp
E7ThNEZZ5Y0d8zX/WFwQjhKAo4FRjLq4pXt6PmPUW6ZVvxtdiYFYPcvEbfZNXOj1
24HabjoRCh7qmi3zh0IlrmDinUHw5cuMabiWAmefvqD3AnXSXvbCLJN1K2bFOsM5
CIf5jjMRBJbPQRhIhFGyhoO/fdHvm/QyKn7Duelz/LK+zTG9MCPK16by2yxD+G7p
fkaoOXKUKqr77nXWv26xsGEUMXMQZQt7vb9vKjLHlkEGVIwwIL8E7N1ECdrJjxMa
SLMQc5ICm3opSkZORaqwriS0j63SeFZlW3Me/4ZeXYvIbqpVOe7UR+gK7dguYNYF
+qT16s6ygH5xWqy67BY7QdA0Eqkv5GAULaxD21db0ucYmWZE6LaTtRK5MXMpdFzZ
OUcMVhGZNw2nap8hF5NmAr2oyUsaCUXa1F2C+/j7cB186T3J/eCdG5pa1yZSrCkT
6IvawdWHiZaOz4WCfxnhXnUomne60OPXymS6Wu1OpvTL2D35mKOGSaryHnbruZjh
WT7fxtwBgmOWxVvug4P0pHBLOzMi4k9QhLRzEQWd8r/4s+1IA1xFfHbduK8TDrEQ
joT4e/XNikNruF63GJzGiqZbKxiAlN/NoQCNMJT7KNVINAM7wDJin7tc4yDixFgY
I6kQsk8/vybbVmOoI7SZ18l0R2i0XGfaGZyr2T26GTwpuWQwzrledDJ9QxSm0chk
4sBFWip5CpFXVtLFfAw4o+BgBcj9C3nGIxJosf9gzhNqVOUey1XaNOTBwIudg25W
cxrUF1kZ7bqxu4OxmP8XbB8eGiki3B6Zqxzaya6YPg8djN7YXnsaCGLAVe0Az54r
fQ6rjnNFohs/N6tC6xUYPRP2KmXhqMRrpcpUVhcqUWbLHbf9uxNvtwcMGAcOfuNA
wnzgxz3YfZ2K7JWOgZszX2s8eDEwHz0Qr8k2xe9BwMqwOPKYjYzllGMBul9ojxKb
Dui3kua4gHDVwEsUhom4BALoamPWuxS6ITu1yTsGJnBlPUsE7qaNuu/PwAnlI+Ux
E9lI5cSIsXASWskM7jyEJHkJc1igmiAcsY7gD9PoxobVsmTtuA+plMpJ4YrapzuZ
6GgmnEuBZ9lxUJgHmooi/0YbKYUbAOlx12+ByKdD2Xc3wG4pYTUd30hn2fG7Sih8
Nva+rYs2J++akYAePzDla4XYyFk68z8bg/DOwvzJL5XWanbCARvuilRjInzKD6xG
md0XMZ9T7J3UnbkdpmC0Hv9WvP8VBab0zvRYvrIoxoaZNePFQmGUdrw3PiWfhPNs
KWpbGiBE66kaIAaJbh7lUSi/NU0ykZBAgmf7kwUSetcLQqM90+5g4DN8ffx9YhRw
WTZBkSOV6cSkdpwFFJf7SDmT6X4W+92JQUJzsEGchLSQfEtkUQFAGhDewVEw1uN4
A0g+Ih847mZgCDTFXKEMISMowYBiRZYBjdDanCkZ4gRSqJGBzT1brXasJhF4ueqm
KvxUt5+FKxZFwIHJ1BLqmnFyD1q4qb7ucsq8dvT/jh5gJDJHDTrjMkO7r5fBVzQg
gVir7CP9TgKusW4JbO0NiDgmeTqUKXctE0A5Id14ufpqow6M8iRWbQN7KO7UlikU
DoYoqAVRhxUv3G5FYhsuvpMtKZ/JNhwpxCN0fwYnGt1NZYn0k4+5HDLmuOKFYDAE
j5m2viDybTM8Ns4Ve9kX50PVRJlxYtv8wNyD0vtfIajrzjiqtGxmolxJbCbWuKQm
gH9dZMG48K0Sr/Oa8W+3Ofw0/3NsoRkXOd2C62mybaplRu8ZDvjT4IP8RcPE1sBl
ha1pupOWXJzoBuaowVMjyFVTW9ksuA3SXCa4DXz9J0MSS5EDsDodiVxgY3lbcaun
XtVdHOLQ2FQY3AopGy23BpXtTtdSbzSdvH5Hgb2SLKJb8/IB5XPWajAyla2cRyCW
bO7WY/q/NvdICFKcbJvd5OBWtOD7FAiNMjtFZN8I9r7l9GtEeXOZfZ35MMByw5oC
2HwQloKlJUfKEiHpqbZbYHfWsZq7XMacowX64sEbChRaI/koPlZY0msZ5iF8/Xyp
TRSjeOKz3qvgZmtmNLJlc9MR3kqoAiciaanYcZvzK47cSQNvvVLlV17q+s6gWfAB
gi3cwGBIHbEWntVnBOxbOwoDC0VOSwbtCxHizz0Oy/nDOaZMuuGUUhRVlsk5GUWi
sIRgsCTLr5XqqxSx0qPld1v7ft/hi2f3pjLG5V6Mq+nabOY3gJRJuIBZIq3GhX00
tyJqjT220Mb95Gz2hXIXGup7gacPbKzA8cpLDFsuMj5lG7IOqUIHpbVR4dlIQYnk
zvsR1KRpZzBYbfh5FfgN+9a2ZRMZDY4rhSnxZq3it7+DhTxwHhjkJ+L6rRO1qdwk
hzzZ01t4XEMZfWhELVQkpON+YPsCaUM3Zjye3Y4pMIy2i6XDHgfMJRG5bN9fqo2J
GK0b9/puGGwy3nLvnyuWPJZC0rPStsnqOoNkL4I412TWHhKBSJMOMVpOJ4u5dn0W
H/JdtVv1bnhOrPirEtykf1UmXJKn2SU07AKjlCUbWLQ7yJU/sKfOGDLgFIURG6/M
hQqjzurkI4ClYD+FWDCBArdxLPNEhq94Bk+y23WuAhVFq4tdLVuUmSKnLWljyAUW
rK2sbttZDKvW2gzXkY3sBcAJFi/aYZjPDG/9cdNlk7zynjfkwMPyFEV28d8HYFj6
YzHL2XbNoAKPUHlD3oX78EgA5PfPONZnfCJ2zDs7P2MaCaWVsectc4UAuNNX1M8W
La/uT3ECaeC4bwg4myoyh8kCclSe/YGEBny4bguMI2fTy+hV3gM/0TmbaWUVvNhB
1Koq8OSibebsydJ0FpFZO+Y7ek+sd4LjeFQU0bXD6OyL1RZzPNdxuk/TQ8fsf2J2
dDTQIBn9L/8p4W7A66OCqiqSubybAVELolGZQC5F5Z79NW/vAOu04Eve5eIP5Fiu
kthW2MRB0ZgkUnM9up/5GXYKvbzhiU6IDDudvw6DjZYhOQOIIzDjcOFijNS+Pmni
cNXB3OLu/t7quuDc2sSkhHB/hPGB4aPWGUy2oW2Sj/4KLPRuPoC678Yh4+0goLvc
0tXqDnRgMAOmLHg63fR6p8JLP9m6PzKpAHNXruxyQ9YtR6Ig7s0JFUiPhD9iCb/4
ni3ehKXyNusQRGZxDjuPls8eDSMNgLGxjyE6awM9AN4RMVNs4pWZOpjzzs5ql3zP
Sxr1WxlvW7No+UrFnh0TMy0mens0x84uLyaH2NPC8X/MuYOMk6s1bP2EuA0hRynn
ZfVH2TH26LQUiTHa0ipzf4fzo9qe4Q9eRp3n50IHq1PUUVyIrwTJ2DqUr9LnG1fI
ecDIhaxuvOxTymRKuee738oZXFJFbVRDBGgz+pjN4UNVmIaMeCI589ZlewSHwvgZ
YMqhAqj787Ybh6+D7vhs6wmA74RNWQJznR3Qc4RkWeZPeRghiXI9jak/y1U3Uh+g
3hG484SB/3xPcToHuUh+3L3CKueY8Gwo7mIJqGmTQZA4bsFcHC9no/4ONz9T5qvz
XAhaz9ziqQESypTLk0IkTvXpXlUtJx5Pw6IjOgbBzPkaWnt80Hs+757IzChFTJvt
y4NVKH3l0MNJprbXG38chxChzn6Ie5x+yyjiNJENfvsFFvIjcXeqnkIFxlAC0CUJ
fBLV5nwGMkQzI3NqjcXa80P9LqOjd8h+JhRvZOLMF+M8xJmA84JhWMVF5rXTjBAW
qO9cs16K0dC7T/9xYUQzyNnp0KPp2VlBvo1lpZgQZk+GC3I74Ye2SgMQhPz2GCBq
hZh0wwGNw2OljGLjNqFCn5TwB13st3dbigxxyTRg23Ukmj4lW7Lzppvb32oJICil
vURdfA+d8O/ddynvNZ51f7XzCzEhbaUZE3uVDPNzekkhihiHyexBzdgoMOUzhbrd
7uz09XkL2G5ajG1dWN0pS5Id6MKJHWVVORdr9KbeCwa0IhTkrtbgAYhO3JEQ9h5U
R/XNsQ80yPmxli+F65jVWOpPwWPbKsta0iX3B98FJ2lpJmozV5zz7aB7aFedcbkL
p6MgH4Vl72jcNbrLGEMWUjE8687xmUd0ZYTwLkNB3jWxv4ugRDBSAoIh70jKzoiq
sEDdc9NLNbajUcgk3CC0+PT0tNPhqyeMBHyV0jH1BM2gP51NgnWJHUsgNiXZpVQH
IhfEBXYuPhO62Q5cS4b9c9itWcyJqwALuPKbLENV3pqfs8YIc8PKbI/MrXxpyN2e
cd3Y+tSzSPtDpAtmo3+/BvD/lVVQLmeJZF8AaP41lhmo5z2a6AD5FI92NnUPaHcB
iySlaq9Gu3Uh/WiXs+NfR1qB42Q/W7uNRN4GV2XUvBP7OZ2FbQk1vrzI5z68vc7M
YhDhmu+eYdRmXah0aOWwAofe5/3IBEfriI2gZRiMbdvXFhxB3kgpCwr/h8jlNjeK
VlJ8m/FpPXTrOEoYjJEjLYUyjYGDs0VTR4rcpplnsUUTm9hw3Fa4UbS0v6XSrtoU
Z5bFd4BARXxa91nvqvQWTk8NQa25oj+wkf6fouZxqKnXhljkpDo9dthi2tRWeoLw
5YpDrPnhFZcZc2Wn1aHIcinubpZQtR3aSYXPsuEik8RftghGWCXXQ8Vbf93d08pY
XqPkBxkaK+DJI2aaZroJWuvSAoccUjKlXHoCmjumJHjmTsCuBrQnde5It9S34ASW
SiinYv/QliqJ8JhiuxO/XwKhuTTx6AvGj43BeEWQGk37Awk3rMUi+U9kaH3DHrxo
F+6Mw2aXZHCVToSzs0f2TpRfvGu/uhrko+MSkcO/X9lp/OdibhstMTzagTJUUF3s
gNdfmnQVp/mKhNnB+Kd9DYn1UOkL5mIi3G31kJTeusyGgTfuETiBEsVcoOVT/Scb
oAPme0C5ZYYCAR7HkvcA49KFNtyEBWJK6d7jNTuK0kFI628uG/uPBafsavpSep9y
yBCr965qVK3RGuurk/bIprQXGHdfFoC9sRtkLFrIh+55VNhEBlfvBUgjXT0dRY72
TBujdpPKaPSqUwZAsnVTMD7PfAjGGRsZlErWcUX1KBGsJMm3TonUxMsht37VS9vW
Hi8cqA6bpUIj5Q3P3CvPn/dZVRLrfJAg/h9Gvhv9amLXcP8slCkA5c3eDZ55yO1g
iriI3G+8KiI700iDFgq7ZL0dc9dAXALq154BfOA7qrV6EUu74nprDDbuenfe9oM4
BuCVDTOtr+T9VGdgBvPAGPA1VdJLhklfT7BnUoxgAWsXBUMxDVk51zGhLBT8BFpZ
15ecqWZZk7DlnUEB2CEwn6C0V/v5Z/aedkd21jL6l0WrY2k14AvvomaMOh13vDE8
9qa5LQ1/r6jKT7++vnUfkqy8y/x/idId4rORf+YBkVidIYW+qeSiAVnbPN+/s4+x
a68Lfp55Rc66fyt0XV+2OBF1jOIYTwhW0dffzAY+1gVH0SdNOpGBbmZq+1phdb26
GR/IjXdpk0qpt918V3YPteoBZMs3MemU4beBlSS5hTReddyvEQpRBPjWopa/9Hx4
Qg+UQJa6uQbHF+VUV8GuCJeshRpxr4/yKO2cio04Inb9Aoa+nGt3TbLSlAZPcbDd
slGz3j1WFLoYvGx/0wbsfHj/z4xQL6aG4ZtOxY4co+EQdPe9KMY3kiG6/UJWw8Fg
lGnhrNtYgFYrCFXMfT/gMXnQ4voUy2dVa79cJgIFGqSUWuiAEboU2/NuHX8/gSyG
vIzTW5VmVYstqdyy4Pv5unYQrtZT6oxPqsYyl0i2HnunkGG8FhpSHxWR0oXHTjHx
IoT6TUPJtUDgTtiHlNx1nuO9GSpLdnrWLNP8NktN+Na78mxrrZ+YUkuRkQlOPE89
BeAQdRMlexTsb4qqMyNSHg16iqb57exUCKFzMQ6zIKYvb/GdgcUsWvT6tf26oS5p
WxDxiKDTVIrr7//cGf+JqYeM5JaMFpx9GMTWdOdU9oSEsbGsKtn+hLSyUWz0nfX9
ksYnGi26VB4QBboo5655LHtp6KNK0HWvyVi5wa/vatD2Z1WUbUrNpH6BCwLSerSF
jQd+sBT6MiuZvMcuklLb4PcYK91liV5C8B60Iwp51UFnyTlb9NkI0P6gUjUnB3/G
AJ+LMTt9Vs7pz5EVDti/BQsMh3Uc4bdnNyC5KZrY/mP+nuZ/KLXMMrUojIqjcBl7
x7V92OY9YQeKoepqJoT54fAmYZsZk5ArezFMVM4Bmfyed5azXT3ys4GFKFn9/Dy8
ecFFlJ29eY0+clZQpt1cQN1UQBoewJdxhrL/mhLVQktmSey9YN0gGsgtJXedB+o3
KA3wMfmoYgUevw1j7YaNJ36L6yAQigZYtwsjGILS0zgfvn1fHe/6LYqJs6/S3787
4zspZgfiWPXRhtSLun0g8T0mKqwHq/gkEb04Y0JEf5ZyB3zcewMK4c01ZpFnqXsW
Xrfr5t3sv0JNLofnTx8nDR/xufvXAsHYTYRZgbm+smg49ObvlGO3B87gh1o3UXw2
f/fAHWSEKtvVnAJ0YjIG0kb8F2b5yJWppqCMfuViwgtkYGvMU+2/QFE2KH5XKrYy
00HvXXNvLHSJw79Ol0r0WZwtD4JUZZwdTiNsJVcq+0+NEIr97EsuVj3xCSt4Q/f3
cDdeurRn2eSZsneh7Zej3EVJG+iWqKxVVfTaZ2dVd/xF4Ahcd5O8KTz0HnB9fkAk
khGVCjIUvs/EtLw1C44MtNoQpUmgmXyW40axqhsWWx+G1Fn5B59AtiKerG40m4oq
NUy40OySoVqGLFOhlxzx+B79DsqaMGa69M97zZkWXtTk5uVZ5KsVLeeYvoEInby0
XQ723Whs2BQL8hfwKDBOxODix0/7j5bLcvaz3RcgyNqYPW5l5tBeUw0LUQ15wEqC
ln933/pN2SgxTQOGJRw5lxfnLrt5BDoeY/ErAkCbSwOTcZ7/NIoXReZBxHPUPqSj
/a7HzX8hAuclfqDtWp8ATV8gj9WSWANaAJIibD7YWl0ex35mU6OEWR5Jnz2zJfC/
03FMUKbcLQDfE8462aYsUM0BC65BdqR3eNEwN1aek9yQX5+SMGTE3nYH38/TBehm
nEkHDZmZwD0dXl5E9BfrujMdjvJLiL1ZuXBlYM0nQRa9IP5HFa2KQ0VfOnyMWOiw
naAgROBzGExCdYQPyGk9NBFi97LoXVb8GFyA/6hMs3Nbmlc4GEMJ+IFDJKY1bovz
E7RjKhEcgG2XfZ9DT6CQ3Z/nIGvPrA+tvR2Z9rBLsXW+r8PwNzJkRPKwVD5y4VA7
OkbFgzWPSauKPhCr+lhkQCnM9ZkalR6JFgBshWF5aHz1+kQiXGkFGUM0smhXwgtw
RoM2dKCYXx+0Fpq7NzaScFivL95EsZsruQ+48BTx4MIvv4KuY1KW4ZmJ2VNH/NXq
xXjU0g31jUOB9U7BcdoKqZnNVZuIBF+4dOYHiXSXKhM9artLEso4JgIjsDlLecuk
Xe8YySieW+WR+eeyWYX97c/GTGVZPI8eJV8EPcZECzQd9UOgFNYraYnFLrSWBzFD
o1sxI5Dq/VOc1LyUA7r75SpGfWp6Y2IVyjp4rrVGIDjSzRue4ndllhRGZ2ZKWnOP
FtqbxESNEDPxDc3pbTX6i3Hs0I1VozmpvqHtJurDpmPkL8caB/Llt/gSJZlb1hZH
pT3mug6cAfVYkNwshlZzaP0r4KrIBoKwkFMS9NgO862JLcWOOatLmBwWcaj1JVEO
L1/cP3To7h26oGYwgsaG/m++0Rjp3l33EsqnPsEwNCvA1891+ZP5wx0uhZB07I8J
ySJDTj0sowqQsyoZ6eAZl2gB/v7wUsfFGvVAYMvYNiU+Izp8P8WmAzZW334jiFca
Lfwqchu6fnBh7kVKnPkvIjmlCbQKlEREztq02KRRxcJ0R85nmzAeKf0OzM0j0iXn
8ApvO+lTqPplBrEorrewGP95WqcQJ71F32aZGgHSbTrB8mYntiKSu1yLjkA9v7xZ
+pwVVgnNd12rx9I1s9SWMgjFqaYb+BtxuFuOQwnNwMlT5+E0sfeWAv11nAhoYP15
n/8tjMPG3SCN/EBDDq+5kkhcRfexPlmY7GHvgkQkxqnC0sgeJluc+AJ5kC8sUqQT
LVwn1hEAw6n0zhaUsfnUtg9xsikYAXxTmxDrE9KdiyFBbwFSbAnBYwcd6GhrNcX5
86jEIe4CrOqXVb2mUEDpSTzyJn6S0/X3fYlsI9Kc/r5BdsZZ6NpNiG+SiOC8L0qg
eDyw5EnJ+oTttJ6sF1WOqvelw/33CSTcRj3TIOhxV5N4INchd6e3a2iT++LL9wO+
UixNlzASyW4zdFU9v9zSRCb6+ksnJKkv3Q7/4Plwxn+WPDgg/4ftiENVniknmTID
brlwdn9C6pCeYswVuew49yDmhG8bj0icBcWdO9xWgsODMy25AeKR8cEsHD1OjQkI
FdyjdSyBhGAt9KqJui8rupReNU/PYdMZ+DdBWtI8nBB7o4Z3sIAXWbT/WpDB0oO/
kTkqmqFI02BIBTjNqigJbkoMcQCxeQgK8MEXo66gnezIRqs+aLmeVG/hCz6j+uRy
NaF58DyM0nWODruvKqGI7dVStH95waQbauSndE7ksIjEzR0FXtn5343yhWq/pl3r
dhHo0LRbNzYZdGlCWhNQORSYIApN33ZC3/BbExF6FRx9VPLvMfh0ATGZDYEq6oTR
LAEBPOzM/B730vTawWqaP8ISxumZ705CxbbZNX7L5jX0+PLDEgL+RRidmS8vCAu1
rZCebFnYyUwrpjId41C7g+WHFVe4OA3WddRv0hE4MvIk+GLd2rNkfWH7QURNk7cA
ME6guvsiPROerLzDOHAqh8ONIw7bQ1S9Py4yUt0HJ7Je+FIDNlcDU+/hkSZsHMik
kGPm3FDLuXQXLG89PCTxWHNoykcwFtH9yjq8gl6zmaGkw30APEHEpK8pyp6igcMU
00TgR74zqPjydd+Ws8pG+1FZqB5558ngpKWkLdaB8f5yw1ufkolxPeT7RRZE+zNp
8BpJipvpY1GCaP9QS7o1DgxlVE6osBYt9P/41akzWiicgpcYNBGMKRagYFnsTcOS
C4JvyKL9Wwe2VBS3BXMfW42youUb4y1GgNu0zQypWrJqz/2d2OqsnIPoPyPRA7To
A4venoDjP4I5IK+qALp+EiVbO3wirk+LbXaTVlX93KJWFh9qX1hayyNg5J4Axwa+
l4KdY7V1JjAEsux8m27gZDr3/i89LpXQbS1JdCYQSTY8Hnn2ndsa85Gmt/OJvsg0
+/3fzs/r4CIReTmVuh3p+PckwBLg7GyRVdcdyykqCsaPYuh5lczRKSLntcAaDRkq
j3G2UzaLAKMGlXc950yZCb4Mctt72s6C8K6FzfNOQHYXyqEIvxMXMGeLqr1B3lYS
BhF/kVgTAqF+emD1+rWX3bGOhlaOmL6EdMQB8g4CBZuyRtJ/z+dSk6LNY4lL8NsH
rNRcJmn8eidgEcW/ACHcR+HhNmPuf0nm1SZ+zY9l7cMvh43cyGNUzOxiPeVXRTgc
q9SZbQYYAHkKx3WWhhdZjZ9RXr7xF+0aJSjFLWMKP5xqadUjeKsgxSKDpcWm380M
ykxPFhHvhQO33XEQ75LQm1JiYGhVC0MJmydcydyvgWTlXB5OEBzV88X2+4vixirB
GbkvNJkWx5OyBhXy2oQCKPJjToBEhcoUZEc09QaiZ+uhw6Jx88XwiZzmBZTAciUW
YaWSYIlpUrUWx6GFmwgAhMND9TnOcOyL9E/EBRNSi3J3nMG0I+GbD123qHZ8WOGt
0LsE0C3weejkwe9fQn4iwmPu+fmnBeKi0l4UhsBJX7+9Bx4dxH3AaoQYIlh3Glrf
Dabn3S5mzzT5lRM65c59uv/EIM8Ik6IRR1MLmx7HU3HOFciXsOBz6tD/HZZipO6t
sl637z9a+xGhaK4doSEnb8bSZDm39c55qqes+sqCvlOkWWHKgcZyEckD56SvlgRJ
yCOf+z/ybXH6vpHyq1NSVzbda65qlrn6MsOTAUVwJTibBFcieQgVHs9kYq60E5Ye
ohThsOT8lUT7Cmb28p6Bp8xqhRyqyzYjuFinUbWsLmX3xDZw19gk4p7bApzaa8uA
Izbd/H7xTGlLthy9TbijK1wNbhHjQso0Fhc0aunk5IgPj44Zv1FPOlLEHjMOjzT9
M7RN/uS/WuLHjsOJeF2P+Qn9nKWijZl6lfFRpHRTJct4Q+ps6RCaneMyVmGsgw8y
2itX8rIryLJJ8EpcimDqWlsPT0X3QFFmtqx88jnDGn6Um/QWf1vBmJmNhRmd2E2i
fObNMfrgOwLS69d9mdkc1zSPZfBVp+CBOyv1LYZlI1tRPfcCW4k9TY89Z4eqMHk5
MlIExFEDsoORdA72szyAkGrMEu/htQ9x3hOG8Ec3PZfAUC1jXEil9zz/Rb05C7Xz
WNqr1uAOvnll2L0+HeishLO4Hb1PmJlHu6XYh5i+lv/OTf47CSj39euMO/KNcfUm
zkfb+l2hV/lpEhdUxKnfejs0oBcfDTMuwulPxDX/x/jMLDttE5McHpeAZctb+Al1
hz4Y6GqYtbSMHKeN3CDsOKvkhiMfSFZ2UmNQjwmP4lXrTdstUZK3OX2jbxfAYzhI
3F/Yqs3XefYsIhsBdNVTsPDWYlPa2xmR3Ae/SDRwuic1kK4IJOOM/WhV/BCYd+px
MXjdZtkbJNd6BP+q+C/n+vBGFIR9ufixg685AIwxd/mvhwwUIInjk1yRBRe6+QWM
rMa7c8I/oJgqUGVOdogGuKVojxQMNmf3t18EG/D9yqIA5nrFcqtU9yf/wrqgcWy7
ilZ8/BSIG0uS+yyKibfh5L4mCsWpWOgi36FFPSP27tvjaTBA9g+36wNmeKsbjl9x
g0+Q3fhLeNlEuVnkrvxSrXdOYc0kUuQBjOoQ+Ll+9/i3qkagw6EwcPDaanzNv1O5
BgOmAIKGjbj42ArnZbMtZazD/Zq4+8iJifRgcrgDy0EBSY9/eUz0htkiHQHHbX1N
cfE7hjmO0Xne6ZOOBNAKUX8Ka+ANNpgS0G8heduekLbfI09AeK/oSCsRJLIWSLrH
K8AItIjs3mnjAO5G5y5ZdVmekyqdq1XR9DBEADwksTocgMqtYc4HaaSCS4uQUscs
AhhfHKCzRIkjkq+QSjHCidQBmLyhd8ljt12tAzsoFtzI9ce9YV+c2JB/yIXEOswk
sxrxb5hPHbZmebyCqIObiC3dYZg6daa3HoqvNHGteA0+lio8msLcvdjnRwe8jAHq
MTLQHi3Gj6GbhLd7KXuVjlsa84btF/8j9+GTTDeQznW1ZRBUXWNpMiAzQRb5GSIY
hHplbllWtoxLvszLT0J2G7AAj5Q/8SyV70x8zeN2zTiQGEAzgnKSYeAox4gZ0YEa
uW9Ipccv2QlEdmxN/LhH/tJRcuOZBI8NQozn7UnwzTysHWOxSABIg3y9v+JSqP37
+wUEbDPhFddT3hmEZCk1EnsDRfytG/7IHtfMDbe05AsKIMxy+sgqAS19pXjeBvhY
JV6qqyhC5woDOIvE7RkAHTH2Nyh73ecyvRIqMuSoe/iHUoAwsp1+76oklV6yCIqn
+dos5oiZVFdpnoe8WtpyELYNgE2L1pC+IDvivVt3p2omY784hwZaL3e7/IxUdMK4
pYMMYp17JduMOPrOx7sRML+uuFg7xS7YnXM7OteQZFAphPpYrwJpinTQiCcaiqp+
PjzvFW40lX2i39Pg8iCtnIr+Haq8VvYne16lL6CX5sU3QdstBb5gfATtXfrfqMzx
+SXTm53XGUFjLAcxh6/RZCxSsvLKpcLbq9Gi16zICHqRNWGHxP/5w2CXZyIkqVJ9
HeuCnrQ9u3Do2aC/1zSgddTSMXvhldtK9PxlDXp7Wcf85FDro8VrVeNeDh+T7LdF
cn2i8s6uUv9TqrmfKRKeOt4uhK0ni747NFSURgmbWWJyy9ozRzsAYDl5157YQkDa
DD3K92gvi+Z770TFwicHG55CLlkOyK6Tdhl/5RpSmS5f0M/RUjwcq8aj/0xYKjDP
YYq/eu7zUPa92kg7uCkeiPSNQdxktkiFNmCNRZYV9E+1y45fTt0iiTxPRV2I29Cd
1JGklHd1VaX4RUqXe2MZBKKbE2nm6OPL7e2Y3lYUeq66tleik8PQWq8sCb/XtkBn
PXPzfATLC6J0f+HNyQEo2RJYJH6e4ONME3exOJe4e2qZCiC9FC2isGh+GOcs9e9i
iu8ulqTdA6xDwu19j0yyhWYCQ3FkWZP5vgqvriHO6OE8pRbRGR1MvnFyLfW7T9sQ
cCxXEB1dS5MdncjFbAUZO9y5DD4Qm6c04FK1pM5Z5ExFLfoiEhNS73gd1BcddRfS
zBFIkdjIj7/NBZbjPLVvgHsF5K6aA8AnYtSs8U/1J0OEIUBhW3lxQaFBQ5ysI2eO
0uJMRvU8gjswNa+H74kr+LFrn17WWgnmwXbBNwx5p/TiBwey7ibcFYRHRRrZx0Qi
pZl11hwXS+VwWFhQCkkq32CcrybdFI9tIr4j+kzmdH4H592OQHOrwV59SSIp5h2v
PRGpKN7rDo5gihqK1F3ILB3KKCUhlFAzRs+4arW4l0i/R4n1ep/Wvjwxwp5CGFS1
jbC4fk8nY9aQGb2JSnygSM20FOs+X2w3AMftbkx3SjuC2hiM4/IyOEo8Tnerqv8K
YmQ4Ex6KVubZiXNhWRc9vO+TLZqE6hGuea743STToLhwGeKjBVQmxeOWkqlonoFK
qIAtCmpsuH7fK0W447381St1PKaoB5s6Q1JAyOKPqtXnZWJ8LVmFdIJ/YHQ6ohn7
6XXcOS6dIPiEC53ovXcTX4AWrE5CDzcKZOJouZbe9SzIb/lHCJz5c5fmmy15Uojg
LD5Ml1bZHfx3qqfFRsQhLZzIWUMVowfxuCAzjnvSoFyBfc6sSYWaBSWyXKbTGiwN
JAcsIvRFABR/uylpzegYclkUiKVBZcDA/QZX6AdyEu6P1nTJKH2jn++25SvqVo/S
p8rcMXCratnMMoP/UAqMOYo4LAmBjYgoRNZ0zDkufkTa+YS8VrDEKOnXVBgYF/5N
zUtm5L7Klgj0dioXTcq/wJqFlGdLsjQF3M0J60jWUxUgUcxEavrYcs8REKKVMiiT
ngDXEU52FYlRVaIN2sMI3498CLBS8JM5G5ybmcICNl/6tOT6zRB1x7xrW2Dd0d69
7jZIgsUYhw3soLgV8f0l9MRVW9ff4TzIDLEj5muGFGAo35m3t894e4CbACkHwg0u
2wTxvaq5E1of1Qjul5gWJCY1Jzn6WFK1H7B+mqM8LksMvtzIA2wZoi7XewQ++nKf
9dZVzhBSzMKCZ/zPQB/mnpQEL4flJsOB+RP0g+2mq2+fZbpr4uo3oNqb90U+SD9j
v/Kt3LkBmGqkTcns7GSpwELR5+v02HIAN4Eg7l0t/xXwwQ2zTTZ9sEwlY/nKOJdz
kbsZhj7fbWBp9lI5+JOOwwf2nRlNWUI78GjjU1YW+UTMMizkjLCnhFnL0mOvP32+
EpVKMw+as/4atIcrSZkAm+VzDT+6rlwFQIFXjWsPiyilGkWBireEZB0pwhHs2rzM
Kx21+0G1U4P7KsIswEWT2BRWbHE5ikhfYZSHxHMNQYxZzt5wxkLFU3kwrDlCvQJY
l0XtxvWnYOS1C40KpW6iN87UrPKs426nSd/6WaGd18Hqs4iiI7uwTP1JZCxu8LAQ
ivrrQPpzLxwAyZU3SfJk4V6a2vgELJVcO+bpqTIeGrt0YWTWGoJT8nMwUZpJP+mT
UrqWskoB8He1Vp58+m1PB/JSh+Zvzhh6TTW0th1nWINFaOGnC79mjUjk+VZTafgK
x8TxmlS67QDnDBZNAKlgOQg8QT4gJPsaTzbpBwLpW9Y2XPJjxLrMlK9FkPQYI/Qq
XOCWgIDmo4txgowwyS23lEOwdmOOdAZiYQLIiNvLO5WKt28FAujynKIoiiyoT3XL
`protect END_PROTECTED
