`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uthLz7aIQtKmKQrmxvlyDnnyp7na3W/fY7hyh0bgJCF9RnmWgvOP2Cf/jB4dWT3A
y31Oqf9IbrhtCSmMv9oaVnn8FKL+2qFH4ysqG+Ued28e4r0fIPzEBzx3Wsir0NpZ
JVlXVDm1rZxCedDSJ9BlsN1EeyEYR5TuviEGrJLg7SqdCMpa8RtMT+rFM7bRIAIL
J93QNW/HmMvwvvu13LkvLyVb8mnTQsnFzeUFnO9EFPsPXjjzUFuaEYmc7GLk6BCr
La43p8gR6E+2gmqX9GreaiPW/IccizH/Z+h3akoTWjJR9P4oJsaBjtRuZ83heCuo
9U/IZ3y3kamQyIyUTpLo+yyUfoAGY0REVq0IJQ30V32nph92NM2jWK+oRo91pdjB
/m3ZzYaaP7ldxSSiRRQuSUqOLNOwz5C4Jvo7U8G93i5pFsYWoiYiJEqGQe7Eh3g1
vPM4v/4tn9CLFSwNMoNJfaDiUN5h2mUcC4CGTpa67oTljonW/rvK6hlEuwNCINb4
JKuBOA3S0Ko78OqSksqu8vepSX726O+Lv0kfn3om+ggy/TVTm1GGKmwWKWGY/srI
GDq5IPqrfV3u4yTBx65JT6piyl7V5v8Pb/Iy5ilJJ2cZIqnmLAoKy6xHDZju0OF7
LSQKLALBHCAdcegEN88heabL79HhQbC9encZTH2KkNg1kWwF9O15Wq+PAvUR0wwv
KOPH+LBjMoz06r77k6OTYSFH0HPYS7hEOXegBBu+GX7f3nIxT89wLl0tlBoBwkqW
s1vQxyGLr7th9hcyLAHCriK3t8wB+XTW2CDfPSADsNjj0xCyEtX/tdS/BRYlSQey
PFimqJitJ9AgU/LrDGzs/hcPAnpaQ9jk+00gMsqA2JMQ+WnlSNCIXmEyQmwLEq+6
7bNod37CV/VCwRy0VCRlf421ZFVxBhAf3IVEeWTRZswmBgP3DkE3dITODEW+QeD+
wYec/KpozIh+60uojfhDvqYtHkeSWFiKPYoCwz+KMYkRleJR2KCYMFkbNgX7FFrC
bB4zGjNGGM/QhliycqGigoDpNj+ARjDsD+GuLY10Ttc6/mwNhn57uyfVn62I/SEe
gyL0nyL0HHr75CbXwU8/xVQFpyg0vuAG4lNWSvhVT475TY71DrL8YvsG3JW5rpTt
lco6uKttuZQkwunHX84KoY7q7G7K/i9kjeddCAEkYKq0P7w1IcGygicxpQkCog+q
NqTbe1vT1PD9PGnpVcXwLrTamyQ8xj5XGZ4pZJsx5c4m7rLhWQ4fCod/PQYnn67b
WY9oYJSVJw93plONNpIft3Zj+jys9ydx6RaWrecFUuWksAxvaPWoJV48iZSPqYh1
3GQ8Wk11DUaeSgie1f3I/e1j4NU5rBUgx9Hg+zofKQtKhakMMsY/8quQPDpqpQIj
3VeNoNv89QfOH7NAUftl73ip1J9kncPKdVhhf/B5HmdCJfDtntkojB1QUUukPSOp
/sz0TiMg9Xs7BDKwL5Q9H+x+SsrO0bzS2Z5q25oiMX7gNKA0DuPlaJDKr3xFSXkh
280eg4kohyCOMz2hU1TH0Dqah0ns5ufedtHWZ4ur1f5M49md6yXGobOdYplsYy0y
J8RVRWqtfNk3kERc7aiIygMUXHx49TzXOhmk8PbpGXLS5ni0LUa8Yh0duquNoy2g
ZbUyL7tdZqygosWaP5nSmzpQYhvC3EUOGHhUTfwkINLcP+w8L4He+IFSmds4IwaV
yxdKRPqyYu00/LmN1xSZq6+HTLFc2Z3+8luN/I0KGpWsywox6I3jNi6E09zTcDcx
pfHB5eZGKA1SP1cTWjeaki7rotUEjSiZp9PFqfx4bR1mFWm6NmXxkF3c5QnNK6Gi
JOvzGZ1ACIkIDoxebv/AnygdNrDLkfd5nj7zVKJ/NE6k9AaejBnQ2IRsVhZa3qXX
lEYrjaBFB21M/IYI7w9k1+pKfOLaIoYWYl/oFrBMkOAzVApg4avqCQAoXMMgV+Qf
x106byREFh3Lw7DTh+2FRY5f6VS9clMCPBWuWb60mgldxA5UqqPaLK2LpWfF3kol
SCrEhphv73cnjm3PNYOc5BqTv0dcrIeSqbmXDeQUCXK4Foxl/0H7FnEACDLNt+wx
2k9u2J+JJXfG+8hMzjxmbn5FP20vSLHp8iyTJEFe3/s1ZpcNITSX4e6IuQT3iNpR
igN5sfm99FgZ02UX246Ph/ZwQrm0liMLT1t7SZYDclFZ/J0pQuZU/TNGpPh5xBQI
eLukUVb+RvvBe7nM5cTSzy5Jv9lywnZiz0gcISAY8IRTqFx/OMbIYgJGMg8TD+vi
QShqRxWXCbyfq/HSbTFJJ0adZpS4litJYtEDkaB7F+kATsCeut7su1wMvC7XtbZ/
22CVXaPi91FOqp2My3taK2N/n4vlPzaC0BWczSwHA64cxMx5fGVM3ASIgkNsJ1pR
BRcf4oaSGxAawEWSIUbLpq+xF8T61GIj5Rf9SUWebwJEmMEoAsk02xsWKvlz6DhH
bzMuyfSRUh9pdKkfp0ivsiYqzQp7HNPQTvnF7jj5YS14iCJPS6+VbFX6G/G0MqO7
0f6ROxZ5Zfk1qGehZFoEdsLsPszL7RBSQxb398+e+gokljvWMLcVNThB1UdaA16f
iGQ1tEpFcQWN5CuptSe96Geb/JjJgVYSJR88ATqnYMLC01S4rnRCRnzrlK8FQczL
LW5Lcg2XTsLP3ipU4dAU6UaqV1gU/MY3RYp83QGnbTAXoNDDsLQbCBhdHcHUupOr
7Imviwy/DMqQWnVyMHkPfyFePCJmeKtDS5LEL3iZK9ARgiiRz1wC5aDXo2mGHnIW
wNcGc1bC2kVSDR5oRi5xKDpIM4WVpaOsfJl0LviX+Mcaq4CLC8dLSXsozPsgNN3l
bUO79+FRHpzlyqSHrzp1ckIxayIC+KAK2Zx4hDnwXQEtmx7KqFIEBm3F1G+MDJcJ
1+BJkODH/VqG7cL+dW4Fp5V7IxWpupSVFYUL89EAvC5rWbeBPHfbv5t52kKQFuGy
z9PrdruNqy9q2OsbuoHEX6f+LocD3dIsXzeuSI2u2oaqt165zAItyB1FAiCl+imD
ozr95tiRNDD2nmbetUMp+58Q+5Z1z7FQdaYkrX2WVKONDbB9XoEhG/IHqGhXPtsn
stBOuXuJXcsuJaEWyHi5d0c+xcd1AA3bua1rSes+PLzqy9z0vMTeKO1LaqONOKci
oC/1h3CrZNkEbGp0wihGaywB1kdMZtytsDvba+tTv6mpSKA47U5ZB1vg+SDvfpPZ
p2yQ/pzln/L2VfzjR7GytyqRC+ShA9202ila7hKn9umaO8neUX78K0nDPp4e2CeL
F458eAAk2nACDhCQs6PtA6ml5cvBSDADpBY72ZkpDu6KRhj/vFu9c64RCA9ru/Rg
Lu4LAamTFrcb6VRsugJZ+QSUR2wXZxGddkv9RRsbG4GD8DQGLxDPCaoZ55IMQix/
wR/rHu/CdfcvF+b9kjH4eMEKMyIlutBpyWhotE+axOL/pYRI7cT/JVnhBCAHZzp3
iIeVSaXt5cbh4pSlyWhhoGnfEQ18MLjCAk4v63UDOZgpUVyjajRPei6Bcvq7qFy0
LksO3SIc+KMCL9tiEJ1oRqTKeBxtvN0u7P/847R9cqypa1SCAP9ytQJwd/eG2ECA
WoWLnlLOuBj50Tn9LEauIhA5hJaVpXrliFXPSG8EpzlruhVHZDIvkZjGhKc/BFNp
HfwYD0sDNbIBOFDQQrYFNYEhJQhnOdIAuDo0D2wKsE5HWtcEiAsjoK+kfAB9xQAZ
Cn4jDJFJlG8L/z57zHktT7hrYPF/X8A849ZrjoLFYUWoCdhzur/sumDlHFTKzIU1
nSOPBNT8Kq8XUgwJ8ZRgHlBdt8/IxpOezUH1eg5qfzJs6mTgXnKoGcKSWtw4IRHr
1hemFGQ7kfiBrnJoI5Pt33KeZqM3siYStM1sRSD3azLIo0cmL/rIKhPx0c1uXqAT
NhJ825w02kbH9Xhk2EmJPXnfZIskTJoRzU4CfVFA/3bOVv02m0B0IBCcvaawsyBv
Ysw6LsARWddQR21A46FcepOsYVDDB3oP9463jpimzOFi7GyOQ+XY8ZiRcHEKN/3c
xb4b454ZuEW3xWLw/QP7k0fxLeo4td8ITE2MBbL8lttpt195xVFlI8ek1MolNRZz
J6yXa9eyshpfiG1j5q5mEYyv3BiqDTn3AfiMSWb62iOhofUiqYfNJxi0LFnI+V+B
CrmSCC5sh9SGXis0mAd/mChtpXQd0qibfm22V56f5kxu/VFf81hClkIIFEYtZEY4
UHDxxWtBBpINhyacGJwtebCSyTieDPRbCz/rgdlu1Ur+RM4Opdru84WHfjSgPGC0
5yS7fCH3qiLC+NTm8ag8iODGWm+R4eSyLnhXUYx6MyNN0v42qzsPn7RgO/KDKqbc
W2cL27dvL5AYM2vkymlOPXFbKZh4UsZc2cqAMCv8tHWS1xL4X0BZucVImBnMgU6y
tUpO27D1Q3jqmT6IWfS7HYOuvURIQ7pFkS4ZxKyt8OXGB8MOIBnqL7PpQqzu8rkj
2vw0JSxrGyl9h16TlIWTZ27vq1NukuXYKWg7mMO66Sfpir6G2ygFsWbT5VN6a5KW
FXA9vPOaYPKbd9ba0ty3hAYYYiZHXAlBViNX+7RfWwKl4mkZMnERkB3r+NfUW07e
91vrUtqM7sfbEBvuIKBMVmFRvNwr/Xd66rjqvxD0OysqxW1hytK822KqjHLuTlh8
VVzp1nipQ8t0WTLi1R4Hw8OGzduicDaiGAidQuf6AdLl8zqQlhuIBXVcpLaN/kNk
NB4jx+Pm6ZvAdebZ/3n0PbdTt8xp3GeJfI2e+VqbfUvHPAzgZyImN/jFVCRkywLG
Qb3eiFy4UpPMaK/MvGWBOf0S1nXcNwJo5h7BIEtwKBDHKfi5b3sHxL7Vda59zqHo
S9HrHN2F6w+7yNw8qjgHZ2lUN5Hqarz34xoDZNcYpOD0d8y+xptas0fhww9eKV5y
P3g05jMba7sh7aez+s/MYPNSFDnNgsva1/i38dom4aW3ApO7yQuOePNJ73Tah+LE
Un1RqXUd1A84q+pWq4oLvvfB4VzyfT2aQiCQlHwz/Kw1kNur0B/VwCxBlx/3kvbK
L/guL5PvjFFowClgSXTYvQPCrts0kxtfw1HcreM5hi1l/aS2f7gpJa0DV2LSz/nm
w74F+gC2GUJT7MxGhOiLZgNRALEUHr/O5007sW+co2vR8KeHdxY7a9u7vOprMcom
/bhp1aD+pDTfnrFUbJN3Wm+Jb9DqpXfBSaREr4lfObe5577M7399yKvfKZyrVDrZ
mVrmx+IQ6hZaOAQCRE7T3fMgAL145MUu+sGSKT1aL/3srMV7RlI2EVkRnk7T0rAQ
i9TTDm4vNoI35L31jS8rUarGuW1NMm0UHAJ8VmgGqqfQVb21fmwH0pH85WRb/xzC
VP4mprY5EX1yj32RKp6Ft/teOLQScSAZVIkIyQ0zW2B0WFUniMDNhndeiODgHYoP
KVNj6g3E0pKQoarV2R51p3a729e5ukTNUDbxp+QKY7YbB8iCsevZjg14kCsRltwi
R7coawJPpjW16Dnwuznp73ZYv08dcalIjV7PBt5JqVbnvHsqFCteCW+SqbzsVybX
ZdPLH/nyMt1miAKtZunLkB4JOYZSP+NZeClVUpwWrLF8j94hFVGZb1hn7NTXD4ny
mMHIIfjuI5WwfyeRGb2AEDccZozJefBtzrSgpwreL/V8Uezakfs2qTlA7oaJQkVu
6s9hWmNXrInZE7n1+yu3q4SnNW61US87i4AtK6ZIPFBXBoxFNhdnZK5ulxazOLAf
vyFb4w43woJQN+QD8oo0ns7+MmKeFlA/lCmTgSIKw/AOGfj6z7vTKLGr1oyODcPS
8Nasnzu1U2TNgztIyWscJDzkdyae5ZYNkeuhtgBhx2UCeyFlF8QlNp8ybHVhwHbE
49sXfSVqyXF10Y9BsMa73iXOV56U3farkAnZ6vXm2HJ7IWegOaiPOZlMBQG4i75K
XHgVIh8PfptiWC15VHWDP1qbQtPTLC2lON0OSUYMUsCcubi6B6MdXI0tzKZtI9GK
TSAEk08y5j3ACCmh+47ewBktU+hcMkGzxERgWXJn2ArAXOYA9jXiYtGDzMvTXcM2
EpKzvaYerWCU9S5f9B5J6Jdy78lmtbcarh9gIlasxGbENDpvyXfK8Iiz0TVHXzwO
8+ASuLGlMAQ0OnWK2WuewJp6rl5rWjHQuo8V8jrbpHWPR6OzNHJKOHyDRNMLaTEG
36MAP7YT5AGx7mMZ0KrlWuuv0a7+DDFd+3ndFGjM8y8Od6YRwY2rkwR9EZixS1F1
va9bLEoxI26D+4qRhQx8rRjV+HU4W8zONtZt+mRlQRt2fX7gQQBmZ+k2yzSixadr
f9aMV44HUZ/urXIvwdcwgbVGWMDcY7yPB+p9SHxQ/qwzvSrexg4Ei3n+yvCd4v64
Z0rIUZAR3GMSnnjHeIWiKZDjyjxa5UDGdMSjRBp+gEUKrEK7/emdAqdNXHCKmUS9
KoSh64bNorxVNsOfProhNjVT5qk1YdU/eHyGzl9HeGXo6LUBrEXld4QifANJsnV/
0eQUAvQ2uzFvUr5IdSYMsz3SLv1lCi7QW6/BMSAYogY6HUBrF6TvGxC6AfH58R0w
Vb4ZZj+eoMC9Cp3iKsvJLRZxBZodB6yqSpdggY9/RG/LWhHipSK2A9LZGXZfTaCO
/X4cdBBLTHVtUw58oXAhsJ1+GDJONd5/UDaOHiomUcuxd2hD0vXZlmSgv99EGn1k
zHWWzV96Sl/7lsDgWBjaokqggQt1AuIU/Y3pAPAtGexbmV2c9DgPZKm4ht+AA9TG
ptQgGxtYQZINE1Dh5MQXNrjpbQwspUXpQOTR/CmyOVZmRtH5JcPEkd7foAFR4QPe
CFf6cDeJFqFO3i+IX5TREqv7RMwlffSwqRjWofrzkiLKuo5qpVpSPmH0z+Ss9cRK
3XFV5QWfbEoObAQWUemHiSn4BwddUqJlV+IsFaOOOm3cse863v6Tgupox+M+GnM7
9lEYV/oqWDMZcEKmQtdOF26A9pz7zgEwyDhS8olpC37jcAqAA+I3lPyTb0Z2nceS
Lgv7/rHsJGmd5OJA7hRr6YamzjQ+C+VDYY8Vl1JB4ZV7ZDnJr+v+esiAPBEH037v
CciKQzSR0r+gh2grAlxYL4b4KdSfOi0xho3VBEMZC6+/ZVmZcu3/pW+nkjoJZiLt
tAcModIj7R8JuDkficnBn+pbIE9V3jALku5QH0d8HhcRyOl8L371NNDNkM6R+hZ6
4R3/aIol59w8neajOAfLLSkkXYB1acyD5MoTYGrvIdCrqai3G7MEDZbYWNJgzDy5
tkiWupE9E8/2p25uTzA2sfKr0VX8EDVBv+MeBCU+6G2kaJaqqMsqm0yiMcNiVe0M
4SFcrB8NNwBneZzuINqFxp+uwv1eg8zpjjEziIyNNcCJ8vpEj3cPQ4xYQbY14Doh
TaUDcXnVzq6XXWQSA0OV+Ik7ApjAzmW0lWeobyGL8pfAYmAfUi8MT9rfgp8XHD9A
s42v0m0GKPKa80J5CTgKJRu8cK/ujrNpxPunqjhkuyy/AWHYTXiWkp8tcY8VFTvW
QZZK1PsP573WYI4iQWEdhdmKloojc5vwgDkTR8CHj384BQ9NN6wqQrSpSJc4bfzi
7FNd6CjLZoWmdvL8TV5N1scd8qQ0yd8xKoGLVj/KWtcfvbc5b4nvaXt9wjaURAsW
QqGrUYlm4Ojv+MghEgpGmTO/e6MBYiFAlphs7qig4+fBd8ej5WaDL3qcerTly1AL
VRo/HUdsHcoUz8nrlk7KxVOvpESjPOopkgWWnQB6XxL7oR4CYbhqVz0lPbAfOJiZ
BPFyJjhpOQtjq+5Mz/UXfcK74/3PUpNJzcHvwTEbnC5nO4/whnYyrytoWOGXOmo1
NK+IfTwTlB9j2K/c+gd/lMivMCgZ27Ga5dFJFspxBiTiTvM21Vs8H9eazb5qnDmy
o8ZEsrtCvownoeJCNVKQfMihkZlJyrMIM57vMLivrbYglnevij40SbeQhaA9i5ew
L2mgh+SnzG9JflSATKVoQfmrV+fR+S+lU3nyOcmwD8y8n+417j/C7dtrkBYZq68G
Y+NLCSljz+fI+TPbz/ZqQ1c6GQxsem5e3bGd23yMIwKiNXWM9uf/oOtdNGk2dUnh
OMmr5YvZ2sqN85pD+wEcL/HBQtXqLTJj4+pf186qePgezPNBgMdLMJkVOU4tzVkT
04FrPO2zCK54bIrG2q8MokIMx6gn6IMiq1kp97dlmFwXFyzYMMQe6i2muqKD8/gJ
pbbpkyVpnAvZAeUeOIMOmtHiVyUVPSdZBtYQjokTyWIJehS7btV4O6060MZTzt3R
JG+lWB8kzlf3Ao812upuJm3mfqqzXq0wEpj3kn+uQFPFqwhdJBQ3jayj6H9ENXv4
ckcys8ty1dVO/2RzZv6ykVv0NA+isf5v6/nyZReG5snVoOEC5aker+zounaKdnzq
USgFRG6k4OoNsbgfm2mMSd96RUOVi7C3Tw3fhvOMPkk8bDMkBDEmp/+4uDrRBo0D
YKAHON7XWs0dxkayd1Dwo52/ViopehSivqme2U0Mc9NGytog+yaDv0TXYQ8rcRZC
gEERsqUXvsOVKBm2a6S3zMvJtr71J4hccjqJlzlagxFeShUCBcowogmxS0qeAtZq
XNcovJtCgNxjBdYsp5Z8+M/jZcognj9i91OmEmPIbF2oQTDaXYK+GK4cZPG5rMDB
0RNz62Xmd9XtA2lt5IDLLUkBYwxFQpBPXN7l1gz1b9D4Vp9ucAqtF+CHG1bB+ihM
8bYsHmJjb1P6g5wVLKwfdQjsi6BuMoIOcGSKtgLPjI6k7MZyFuusoOx2bJmuOGjS
Eeghqj3Z5FYYjJT3+ITkV1MojFSYstXdZJpSs6BVuRFRCB0Al56NKyyEBmReEXr8
pm3lTQ2mk0FSWSyuSyANhwOQhy5QYKFkq70FbhoK7tUTPmUqRGXmYbnMIWyvooAb
Xqc5iyzdLOOs6NLgNdb2h8Htnt0pKtFlzVYOp7hWVVD41HF4I4PEbTxhJ2blF6R5
x+JaxJGMCAWEfhv15pQjlj5/501mAxUtKd1n6ujAlNmCR7D0GgJqoH+/ex9iPgGp
/aZWeq5Z0AJzambp7lKbW7Ubp8oWS/RtXNvCiw0S2ISuzRueVQ6SUQDfwKOJk2Bz
QD2QwsXn9/X1rVSzgZZSJvSbLkUon2lAJtDaAeUZXOyvuG+1WyZOJVAsRcg0vXjt
fiOPU5RbeNau1Od8p+MvSXyxQl69jWb29PUDj6qeLp0syX3lrDw2W+S7GoEsz/ov
cDPHsgrI7ie30uiHsbcXbUQiAVGtb6BTQgV4KjJWjnAjJo4F4z07e61VjXTfX7Ea
SGcfGq7lar2HGq0M3VMrxYolPdbUlXxmjAL9atf3FClIX+jy2NXxsx+BtSXNyfSR
uV3UdrsFXA/2FYSL7r5MYNiWSaEAm5GUuDssD8TKlIhPWHgD6arWSQfywx8V8eGf
1BtbhZ09LtBPJcKx0fumid/a9ZkuHWCL04xnJjqnjmFOy95TE2P1p/ZM50WTSh8W
T0KBAYPHuI/JbpRip8CUV/6joTK4vdIhv1LQNPQCWZkWbd3vCLIsHbNaeAnxEpEA
kuClIvqV5gkI/ZIkAHIs5aKNO8dTJ/pVbiCJvr/g9UryrW38eEeyvO8qedRR94VV
7c/es57wt2bs5ZYMg9PArxBdmyZ2i6VeY+uNIsk4SP9Wxeq+q99mTsVM5vzPQyvr
ZEQMwVk9+tpswOmb6WopSWyegbfGvtNJhXbkxuKSZ5fMX2o2juIAA0KSjoTrJIXj
ZbSiZbKbjTKqJakNFos92pXm6nKUm9H2D0fRpPMmgQFFzu9o8Rorusd+wfFkvQOW
XRx2J425GVHItzUsaBVHXhhkRJRBUTjm9FicceN9V7vlSKOPsGWMS0cFo8HyNKa0
Y0vbq/ory9F0KwMXWBsQXY51UJAuTbrIBp4PD4N2bMpP3pEe2Y4YsbheW/+IrA/m
rFoYbGnpW2YhopuFiq/iMcrR2alenjULgdnH5KTIQGba1eRrSs8rtXXRyX7pVv56
NraInVtWB6UIWbqiyel19o6Zw9edapUOMCzIjQdeXGU2p5F1zgCPqmQh1x4JiyF9
ZV4V4wSOcp3WFy1+gn0y2KdQNe1f6sVeHZD3163fokPF0iZ2H1QtJhwlipSd0tm2
kIGuQZsBzBOCuOaPrVE8hFkThvCjYmbekrae3vnsfNfwCY/nXnRyuWpjYcyvhfL6
u1wDTFf5HPHO2zkHT1P9PJg9r3STOfFgKlCK/IjzxVpSHDd/dzr0QzgZWdaeywFe
SvXJTNiw9T8hw2OwbzAKqjWrCcEbf0ad8FmzLqnTTFUsLnsBnxldCwOHMJe+Yvj5
Qh5G+1FRN4GNmnrqbsVJUfeiJisareX94WckS4wvisqZHeNyx9nGvOQr4KcCplhG
fzmGBUgMiqXjZHDtbZqVCVzT5lt5h655EhilP3E60n3/+8Hhv0QaZrIo+t/jGu6H
itZwUSgZBKpm5JUG5eKDIsww0Ja/Om+UqpVwxDnsM5KPBA48fHrugRrVQoE5v/OA
IMjkuEIS3HCswqYxFF8BL0xACJJcvKZ2cqulINkczx6mZJJvuU3Csaydit27Xsf5
Fdntnig8oo1HxNstpz3KxdL5kmC595JnDLs4BAxLd07UWp5ADupDl+SZuC5bveXh
xIVVpN64lrRLJd3MWRKvgk9/xT1KocQUP9dwW2F26+fxI1fh3cuqAN2ZoDw/a+Vp
GKt8A2ZVKdTrq0rRK/PnyIifYtHffwGt/Kcglbxhc/Zr/UsJR9sSuD0+xkTrSJYA
r88U/+/1tuI9gahJ2V7//YHNXmtPiqUlQnGaNCz5OCdYPj1u9dNay0rtN5ByAEx9
UbZt1xdrnnTGHyQ7RZdW7Ka/SlPt9PgxZokOf29wkS0CCI3qeAvhDAYq2cNw+l3r
GH3V2iEWeBv2kNMyWlzZJ4NobDA29Sen+0NQw71Pk/tKhXAg7XMnNkdEi9ldHVId
xHAn9thGuHF2Lv+TjiQtZCy01D+cbRIRKGgLBc2MYsEO9TJz2lYw5PaxCVIKFvVJ
TIG+LCnNruhXtMZrbjMBKoEormTMVGNvwR9tRbtOqJo+MDMBdIL9xZmvF4cGFrwH
sKjJHyl1A8Qha3WpgkqUSkdFbo88AcY1P4XpKf5FSjUBYsF59Pk0B0TWkLtTo9xr
w5P2kKwaQ55S5+c/FkACBP4dOJYmpm1xJnolNdMvi3dlKB7fp4LKgpAnNvnMmnLl
W+Ey8HB+8nBf4XlyC5SplKbWk5MyLWrtcRBgH7LIBppw4BfTcoOgD1IBjHQATnYu
EJF9xgVM0KVcc9cgktOkXVBb6CQGTKbocUINETmXPiZxtbhIlsTWXxRFeLiP4LpX
tWaTrELr6cQKBhQCv6GpIVsDjTiqNox/8gbi/3qGfh6EBljpXNX6R6O8GN7/uyfK
OJ+8Z1+0xw5xsRLFwv1kpEuH6S4R9Xp8hHhc9PikvPDxlZ95tBENbfg6WU/IsHR+
Au4xaTgeWI63WDHd4pYAhmOrMJKy8ON7abdZ6He45CJonD/Vi1rQXtx3Y96hHORE
M5IQ1wRoPTLgXVVudAreg18vbYsnjgpKIEFYMBJdme/D5RWh3NSzVX1olKi7BWQD
o1+N02RyqBLU1s5yFQOeENvursurt1A79vHvdhQTvb2CKoXt+Bw2K4/N3CJ/2W0s
+DxKbjI90UZAHT/Ac1ZRkHCxjV5qfoUN89AgfvrrLQT07HoLokDPHgQA6jLYBuis
6LUmn1JoGN98LyumHYnJPooPbITM9a4H5sexw5IjesK5Gcri0ppib5p41WlqV1JB
6haL6A/h6KA1kKUs983g8iRRA8NUdTdHZcMfzuQdz2uUe5sBH/8UHez7iGf2f9KM
gQ4e1H+CnUTQP35id24qllDmUkdcWmqXjPoboBzBh1L4XVv3ionXv3ZzKjvvlsYw
BSHZ1PcrOSZCna0bHdlgAqmjDpTazQgFRP8MbHDn8m56d+bq+KVqvqcUJdro/mgg
yYMVGUON0RkW73oUdPo+bp3TBHD0AQEVo+2q3mNrD9MOJa75xXS5uZ2vOfEr8qEP
von1shy91MsiM49VtDIinZyHOA/KNZTnNrnVu1NHAcy72jXjdj3M9aVeEsrHpLgo
RLuq+SOobr3Rqsu7iY942N2xZA9DVwvk3fwk2OBJUDDZfHnaf7NQIVudW4PkEPSG
Tfdofq+Nk5sKXtcZmFpXlJNmRwJMKNrJDTb6G5I+hOlfvXKHTWpNf5nRU/h+922s
DQHSWeS7fKLB2fEtZ+pZ5nFxOo5uPyZQy0vSLFDxT3NjMkDyYGyMyyiCyqFeeMPd
xkxnWrB4KOvDoSxKHzMIXpk3F0mqypf5Gd0JDHD7EPByXFq8SKpxSbICNKDaavqS
dfin6NA1gbSJg4p8tVRZjP2LNRs/2Klq+kxbWAt10YmWeWU47kf3fvGdbqLjR6ih
uKivVeT2oRri8EXa0SVSCAMgLdrjASWV1XJGJXB5CD9Qa3Vc0Vfi2XiydXQeIHjP
Pqa1vNvYtRo1I6Fkc/CV9eoSQEN8uAWe3n/N4OgdzxVI69FOqIVZsfvMtu7z8+He
m621AA4p+lcPLH55a8AKJZjjQ62B3/NIZAOleqXuZM0m7/dxJMkwiYkqBmSoBVBl
HVA5ygbkTixlkIjpG1wnaAmH3HmF7V+U0BBjAhaszsdzASytqVk7688N89cMV0yj
7Ol/DodZQB2dHgQTjPeNf9IplPPNSp3dOtOYB2Wwisd98KzwcX26yz6ys1Ppss3l
dKw5zbEgftpFFYlBMJytMfL4XFl6KE3e4iTMwbLSCd+IFRpE8Kz0bIMrepNzZYr7
94tPYhspqv9C1o3+BOtFxAhvQpS9pRDs+7cuXdmXiunLI+mSbc2zatEyFWe2UcyC
H5TPzkbqIrpX4AxYKbNoDUavECo8IstkX/NGgw/gQITURaFxkpyEfxjAv1DH24in
KpQpYxNiUFjAdhGPMF9rwxs3lQyvDU0W+E+MLiQmk5xYQ7BlhPfi0oBzhYmWePK3
JqjisBc5CZtt8poznGfhdhQ9XhrFPeZ6tw45ES6RCGcXeL5MWqUe8FpR4pfm/fPw
QL1AazHXCY3HabyGCppLRqOzUnotKVG6cBrq5vjdPgQRXK2xjGTdjjJM3Cp9gL5R
Czvgy/Y754xqvag8vzZCMRfjO2QoBKyDOj2VBJyS379zcFwtedT3J9TS5rE4rBSS
zCnVKttX8ATDkxDx0bP6WxAC8kxIy+7F39Ncneu2uR9bs/3jujHeACg7gpFbky3y
nrLk6tGEY4ofoVXUlIelrl1S5P/bueieAY1hGYcqxl2//uXwR+RqceRYIMqG0LU/
BtjqfOQSmZtbtPsdymbGgcuimuVMcmtsxEGcrebIHssSPAcPss4bCnA4US/DilWT
/McpkMJEsjv28M5jWD71z60VfvCvNz1H5UqWOmweb6ExrxvC4gnPV2/941NA5Fe/
NDWJ5PjeFgkMARCvRfcBgs2B//5t9dP3kFrajVcBr7niWeSTrkgQvYe10Sxh/Mft
dWn/oWQV2Otd+kTyU0FGVbciadMMB+NTPHI0CClrZX0Ox89BMwOeYgDAzSb8Lp6z
c/V5+pBYsi8FXwH8OCpppz4NHo3tQIy5R12uQuDsuG5+W2Mbt2TemSWPwR7aX6NP
a8Y8xb1eep7saoqZQ0hLmm/upyDXOvrhvPyLm1lPdh/dL/QQHU1MIZo0SHW1ZZnV
aWKgU0Dpj/ID7yew8Of3BUwSgpiWBa2XEsKJHCP9Kb0P+ukLSn5h5zl3/bXxHyek
m3L3ue/8I+9G9mJRKKPYhWX7qyi2TU3GfmBTBnCDwiTeRzjyFC+sidvaraucpjxN
5GP0jgakcutm5h6PUfbPmquxcVVDbeaCbEUsZPbRs7VBiQNrtVvoqRKy/ERD52+q
kilkDPIGZxgjknUBhxXUkSUA8t5A5HfNp54JnzIA5dDLHaizgeewKGNqmYD7bG9p
CktHLU0WAPdn2Sw40p9eiZiQTiivtoduLm6QYRBvdbPiXDy9G4abDyI+0dOkvwUx
BAZbLEBzaheCh745f7BZ2KiYkNvuiq8xdntGxtXBstg2qkKQc554b16Vr+Dd6vDY
s9vnawF8JCoejmpaMPuF5uMC8/XvjNazqmi6nyWHIHug99rbWW8yPoGwE0H4bqb6
BNKFTjfURTT3n1IE3CAUPPfBq7N5vaz2scfyCjpm+MvyhoczAYvdP/lTO1I39y/W
GXSyFbYuF4ZuLvOxdxODOB2DxBVXN66BrRn1/oQqGYaMB4Tce8NvOMuPrBgY+hCI
O5jzC1kQIEMnNjjZ4iQYY5l6+iG2VA/CmcO5SQuVaKG8gUDqYlucW9+qRZgEX3+2
jxPt4C+WVOLucYVw7JI04iNIJvppwcq1bzs0LsaS5UfNAgKZEUTvjEWh95xQ/cv0
4kHZn6heOt4A2pX2VU+GWmT6sfWK5qNf28ddFNWcNeoj8vK2Ek/v7Ylp2OdNvn+R
2PK+I2eUPRNjdr3EMcAXbeKWo01z561i2gDuCNAuFbS1zq6Pq7x3VpDmLffycE2S
pMuQBzPASNV7zfji0p+qDfWsQs6JbbFCZ1jciPq0hD0ENLMRmWq88hJByF17tMER
DlwEjBprA0w2FSKQtbWRRZvCmn+ZzYY9GrSdLmjncbcq2QmO7l1UY8Z285P+VNJr
/d4URXvS1zeVeMQ92quetRZlTfLT+6V7zHtBQTnMxl1IUsjoS2PiImKMjKIyAagR
CboPmZZKdgo7ssAt+FXLUriUUdsnogSm/hJo21KeMeD73OYwd2Y/3UXks8Q1CM16
7WwjRW2r0ydTU0DBnesomO9tUZSWsrs9AKKKeEACuW+JqalHdBfYXkCT0823ovKc
`protect END_PROTECTED
