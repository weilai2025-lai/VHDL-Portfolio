`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rr0cwjalvX5z8gNd+ddHMLT/EjhffxFKOrshDh/07jfDbjZFSwAwXCVIToNucePq
rJYrSiXjH/tR8FCWugDkop5QPpNUdT54lkMYBrgVuGNyj/JNbdOv7UvrkGCkikmh
T4fEsy2CRBSCniPfTkzFsTPoFlY7FJFnjjR/rX5HXnHLq0wpWzRo/08GDnL0ghij
pKXQMEjYOwT99BwQR3NxzxzOeMk/d6DUNEmb4pcHeJ1Bocn78IIkxGC0CnCAV2rN
0cK3qRY+FZDbKuIDQa5fUkIcgMKiBxzHlhux7WC9GVruuGr1UjydbdU1L1hpaURR
0A4xEJ7dawBiWwoPz5QfuAt+BMWR/JEsRDyAKHRmaGA9Ge/yFA33Sp/AaQ1Rp49r
bkQi1Zr66pRRB1E5jCRJCMplrVjJxLOXE6sh8cKLlTBntN9D4JsdBRFIMaEzRNsG
5UES+ufRyXvRDAyYNgGMvvfnxMOxyp4kS5P9FoJR5VhG/Xs175x44oQVxzM2FayT
19GEa+yWEj5Zr7UGp/d9HKA2FWfre84MfVIFpXFQXatF7aTuMoahWm7LDs5jcWk4
twgKTXaC1BNBZmKdqXN7dQMwy39GKQibYKkPPyidgabcCRqEn9WyimZoHxt24DjQ
loMpoHWJ2fn51D+b6AhPofpJ7MGZL9Hnrw/z+ODKa0j/UmamT260zO2cNOIdI/GK
47AP32t2rUdE4/hRBcjw0jTDjF1STThuonZvo56D7QRPzROB6nupX9BUgdArzOJ/
Bf6dzACkPsyjRLRFSdt8e2dY9eQA3HNGSp7pfr/AkXUQ4IOMCTWDAgdmHbFcR+Pw
88bkEUyGW3IQcE1da8A2tLV7FPnwwqcRjv4e04prq/OSYImIwtejbWx7xJUGuhsH
GGNP5BztsnLAMiy9OHEBnZ1IWkoqjVAd7hiEm5jbL7OmIHJR8fD3lE5JZIiUKzXA
EhnBBvUDzwCIzn2wDMyAaCZkrbLFbYRfUDCi0k5dPiJa1GTIJhOAPnSlRo66g2ja
985d0f3JR31wIHeZVRc6i2aHEqsX1o52TCa/a8NbanzfEt0gyVf61Yt28908uiMd
bL9d7onV6JS737OGsUoVfEH7AeEHyAZstJCp7Y6ndsN3mNrHPGH+9C0x4Tv6kaNx
keIht9Ge0F3g/ehwPkjSGBnnL2f+b7YDVmaAvC0i8JWeXKn4uDBNoofGQThqAaxU
jwe1RvTeO651vC1MeA5XTwfMe4glgkjyjq5oKP8nP22vksp+Cav3/J50C9RKgpgW
N/qqYeCXf3ZauoyfbvXCSQxVTMxsGQI/RrQINFCC+ilClLqnBG23TyTZ9efF3b0t
igMbPk8z+wLwc2RCdxnMrgwz2RYIyvErIunAaBsVCqa55ZDNknQDK7PBH1rU9uT0
hc0ueSfURinuDmi8pmYcgUwmx++PKrQxZSfkuAbm2173rcHTJYHgfb4Dxxnn2hTR
kslyvj57MwvQVLfprKNP2CgpeCOD/fPH4bavdj/Qhy7CwHWemVcmQuwN2r2nm3LD
Mm5EJMB5iLF8guZbF8GmC3PFfKB5G8lCDRsWvIrj6L05DENq4e8kiEwhmF3S6cav
g1D4KJqJeHCiIZqWSGrzBXX9Q+ZsXayyHUtdACQztD33DWnrjpRMKI9ZFfKaKMVT
wGr65ysc5USW0ZRuQHIZlPnN174TMDKfiwVNuGQs/afjbLOhkWZilEzzU+cXy3eB
YkuDIQKCTDzSgTEToomQpdyHCtAeaAhxkcJ8Fmgiduu0reWRySiVkBuTW9Ocs5Q9
HgZ2y/J4aE7yHG/n/Kka/CSZ1XbsIatwiwtuNbazC/01ytJa5nF0YDDwvxr0acHO
1CoCLlih+97ueveUzs9Ykn4kODx9a0Ww7+nVzJ59+LUV87FBwDKFiD0GdKZtw9at
DNret6pcBXDZ/uMdKStOm0rD63ye0kiH3gF4BHykG2g63RrV3KoMV0wt1ihlG5+J
9UkIfjfIVLbaht2D9tj2f6tmv+jJb5GGOacDmzxmU4u8ULSZSjM8sRHnyfWpZRVa
rm8ag5dsIo3blt/PVc7fuv1pPvpP5eCy8rIVDPuSE4xVarr5FyxhpEy/OFxEEkPF
CHsmfdsXkOG2/QFhoHd114rtqBuoFoXGE8VUS1qbcQznI9ZLVbR4StVpD/c2GXax
6kLZSSAQz/JOmPawEANICczOf16+MoSpZBWG+TYIwI2QaTC2tgm+rx9n7ZdmARJR
mEoSjw7sV0YM7iC3+X1TaWVzWZ/9jfsZ3LoPr3W+G6TcE7fTTHRhsROt+xjF2ZKK
wCjDnmTKcwFDz1FYzxky2eVddLivyblvSrzR0o/5ihRPw6ELLY4Tq/C7R5tGr3cC
CnO41Hsg4W8Ks+0+1ZsJgk1Mu+uyrPBSo7zDdjF3ERvniu9WBXz4QjoWQi5BS3vu
03IecWNSbNaVHFitdzy8IxwbZNcG+/5dMZwi/pOtfJgVMMS3Il037FuZXM16M9VY
d5/iSPa1K/x9a2BcFov9891WijEYDcCPHlV1Ljfy6D4bRTK0tTPJHybq4lS/OypM
vAgB+NrGs1NJharwj5R41ljc72s9VGnMSFOYOGh0LeC4K32y1CQ5xM52f/uIsgbq
5bNZcw1HPQIak6/BVZawupnZFewhQVOBgCHdM6bs3BrP/0fxLWILhTUZuf0DvXxa
CVOHCPXEbUtkw4bgURGpDVwomDpsjhw3Rq4yIaAfq+YV4aNXNB5XGfnWAsvdtm81
TuH8xZWybl8B3cRKZZ7F9Gc+jYOdBeSEITPF91XxXkWP1MhO7tJZFhVu4SlG3YjQ
zZRBfqNKpNamWwNk5NCHjBygMW2W6+bRM3uGLNpy4f+JB5ayKv0MnGU2512EeaNs
XVNFCjwnhgY4mkuIA6Si8UfXsXfNd1mRlNUIrs1J8G6d1e7XSQRcgHnzsKRdhdzN
pG3f5FgpkTln95Rw5lkqI4/tiKXtspCRwfMHHDDmI+kLI3/qPoF18lhbEOzG8zIx
1J0ISXg6inVKX1kBCD9sW/Vo4eBdJm3xVoS+OoNvHzoJ1F8wsNTtaNzTPZx6Xkss
IaV7KJmsdxTI8SrkwM1HR8TghJczYt4rtTGpkbjhycNPiXBO1A0QBBNzlfeD0NPm
SuHXjbARMc3j6vFoI2rGwErh7oSr1WQDGNWZu/cS+vEBEqvaoCFPRGOsg/euamAj
Q3+XbusjbYK8g8jKkRHFk5BEnJLOlxcRwFiS/zPGQ8iLGeUzYZxH9wPvwD82jd6j
TPlCqWyxHqsE7aBpztj4N5BzzkhbL53V/omnneSn9h7772ZZ/12+JRTkQSQbaIhz
oah8MI9xEtLnq1s+AHC7dB4qahDRskKAWYaH7Q6lSRsxc3RGK90nIwhz+MZupOWo
JKSlrH2qmidddTs3kjXT4lHRCWScRGK6CrLhW07pNOOfafmibHrfJ8iss9mbZVGx
Mk+Ow0mg0/Je/8PXa3ptO5m1QxDnb0zddle3z0WMG5VOAvQiNARJ43dqOTlgT/Lv
J6q8ObLcRh1XypuHeaU2UZg/R3wPWwmizTU6F3RZgywZb7fZQ5h6jB2ORATqnclP
tob1XJcU1FjUu/eK2mDsdrdO1nWZ4c/LGgfqAs3IFnHnQx798aUN7rZ34OYy1vnf
tjBeo+0pkmvkQWa83zoTbtACdTTXiZ3qzntaDkNDgo6HT0YIM0oTEU/IHa6OkFym
bMyObToA/W/eVn4Pq3Mo46ZsV+KjMsl+l+Uha+KeORh84DK0gJq1hpUmbID/2Z0i
fyiLmguBc4T7b34uPn7Vsg5WfqssR6CWT70wak0P0gTwCvzaoV5Cuu1+BSsIkr6N
6TsU/HCzeifYTQjOQRCYYYP+mgtROW/kNlkJzHwVndJIkNpfjsBlx7pvXdqWeyks
LLbGwFuoO2fihl0ldkgkuj2k3ihiprAnXEThUxGjK/V5ducSUUbcWYxcqV4qeIqF
FVZG+1AmanmP1UhJxiLM9hJ9JlgHI0xznsOiZ8N8+iQY6Li77Fnfb9T0qBLO7REV
tD94xi8Hc6zjn38Qa+pCJ/dEAkA9zN/tg4ry1wTSR5C5fawT7URA3rmdYtJYOyCb
SkyM2rS5Eq1VgxFR8h4ExWue3vgvZ5aMJlwIWIAnEPVxG2QhlpVPebxC0vHvWzuB
vyAzRRLAjN2T915VoGKTXxQf/LO33VljCo0++52CYTSzmrvmZQOsqDRPrBUgZ1lq
wUyiZUM0bFEU9u4jssgry5o2Pwb1wQeK6rUQR4EXYtp+tdNOiIeao2o6uWYm0RyG
ef19PmBqDhE1NoVOW8IkQiBD6XwOC2geo7auiE48MVJEIYOpHhf+5lSuL+ZhMgxq
0jz4qsc81YKfmrTMdPtN9DTaf8ZHlVP7T1+AWu4rThJOb4f3mGZY7c4m/TOLOS5/
tD1t/M70gt0jYze2rKISsXamyC2B+cm5UeG4lC9kHGrDuXHFUf6KYZ25bWzRzMmp
0HFNdXSuIx/eE6mAHZQcIzHA/ZLSJ+wQA5zYqVrnNADPjOUUTj/uaN6400zRrRHF
I195Llg/pkyuDfJE2y0lUny+UrfwE0RH2R6TCBM8EzO+m/3Tm56ktfOgky7Iyr5r
PFCAWcJjJx3s59SYoicHGYlMwgQmGy8ajmN0Ew1/vE4DyrsGagZjx60Knig0dI92
RudjWzDDx02ChVwhmDc4aqg8xIo7DqPE4DsWd1L7ykzmxNZlPXwOPYsrxRsluVYa
d6b5BbfHLx80yI0ldmjFyo0HR7MS83PaQBUSPpuEXaJZX4NJ/YchWH2wUWSJRMmF
i3Wbg9/9LcuL2WeltSII3p//Q4ec2wemNdK5vOKPPw31LQCl5UzM+RcXWRnEzGfX
cm9kFwpo/VTncONS/m/hCHblwBTXC2NdPTXhkZ6wTODivhhtQxUy7aT4SJG4bXXI
VFVZEbHAcWyzmby2nDJ+jvt7XmBB7kPRFEqANTxW9kvzP+SrJge3fDdJsx86Sw2T
6JLbz69nCfG5RLbvlJ6i8VitIMj+o7TC6v2f8z2v9ZVWLV0d8sRLGLccDc6Dl+6k
UApzJxlOe72UiHW6eNOGwzMjCws6HvxHZuYL2i1okd4Zcpg5Toj0o8/GgegBgNfE
I5/xifm+YnVJaOaXbHUs5frl0YwMrumTK7Bwq9CwFGdvquHir4akg1MzBgq4AVhD
gXzhVM8bkab/+o4vKCMA4La05blBGJkKExdzKYTU1HD8bHR9Aj2Tyvr4HcxMEGNn
jXzomc1OV6VTvt7EgBCrx+Gnz2gpYbDCoQ2rA7kvBIGidL6atAxmSszLuKA/gbwz
ZEL0S2NptQTtnGR2IMpzIaCoS44/jAdhtSNiNil1mdU3iCbnGN0JCHNT3I1aLtiB
MVZdPouVWK3K8wiZI1DtbDm9stWp4Xq3I/DizbSF0X32BCOR/GeIqGelyE3JxZAl
mkmMnlA6Q53M6+89uv6lAgPl5lI0o57HkzBVJpTn6k3CGB85YLikfIpQZNcU2ywN
LGrqqR9YejgRXu4xi/oTVVsNkWdtTbH6c/XITHPN/vjgxnBGDxCacC3/ne8KomZL
h4Cw7q/RVI2KGpBk4cOX8/h7leHR638d6Bi9HpWMJwjMnx+tJooykbDFKejYCrhv
uW4nS+iXi1PU08YBGh0nEG7Ysl7X0s3+9YCNaQpQFIkZFh/lcxW44AQ8esd5sXGe
SwPKUKBiYveduvcmXFmQ8WzyWBXak7oSZKnWXwIX2EHtqvq5js0/g3vDbwCtNVyg
rdkVaTB8NFw3Aok3oeTcZ/8PfTRkGyQg4nUcP8UlYiVV5OUf3xmwrvw/0pIyOzOz
Pxaz/mVFL1NPJnu3lYfmXlM97zLRjg5CUwjqgTZmQ0/qzMP5kfb0b2rl1IzyTkGD
teBNaDrVNOZBiO1tvHTX1D12PjRlVI1zERYA2Cp4WA9gw2rc1UwJl+djBPoxgigt
muB054ssEAimPHVxem6KmqYVj+U9gGXxB0oqWElfmRuQVAzyVUBhbChgPtTZUU5G
hNBL+sZFarlgrkyc7sgj1gw9stn7aZkNYqNHRAgnAPllgUgA3S6/Bmg59/iS3NFx
rioxKlMvF/0U+1LY+YYf8MR4hph/RthVJSYfrciKjX7nf8Fr3ym8lR6BseyIePxJ
DkszSXMFTrkMhBSCRDo2A1XZzcDM0LUPPT3v/0rmMnVwM/j9PdgrPwvgxB6+m5Qe
9K0Vq2xZR+ZMaNQ2b3o4GTpkCu3sfNvJP7ngknxr06cc+2H0zIB8S8RmYVsFitH+
vwyDLqUDchuP1tOXg/10/hnWk8Gia9Zw3Tou549/G9fa1c88siW+sV9wVVr70xGr
ByzQnXmIM/bue+Dx+/3MDy94bvF74o3rdH1fGwvAp8a++Z8JgebzlfFvWFuXqbWv
2up/Jrm3XDq0uoo5ydJ6EY6GIZA1+QbcpsSqea3y4IOQ76oBIixNl5R/xSd1IfpH
+ir7AFgG3175q4EBUbnaK5rVALkypQLezoI/zaNwzgUMgMSEixTTkUT20+i0U+3p
WuHcsEuniCUZnVFwiBrJR8VRV7zZXBnhqLMwGwU7JvhAYXGFVhTqfeIrXNVZcdNs
OFFzgwo6IW9frtlsd19rAz/xfW1Zg+VpDFduJbTjKfh6M4XLJ77BE5DQpuOmCPq6
kKGYtvrmMdCNEa1QsqK7P0Q5OTPYHQE/cd13ZijBqpmmYav9kiqzWVIG7kUWWnIE
f3KsyKwO5LTRGOfNNVwYAnzndlB3lzrPhGrdb+1yRSUgm3Lb0gDn14bTaB9sB6ue
qUgJjudHUrP62eYco7iH6XHMVT7cp8FMGxms/3dznhzM9GpE4u4QW+BQzrKPcyGX
appG0qXYkK1s5ICnUP/MBJpNMx+ajkPfK7iwJYBsXN1uKA7h6qjhkiMSeDIFUGFb
Sf9NMIQhzX2pITavnsbxk2Bq0y4E3ubZMXAjyTKbXSxBJNjwrtcRuIf2Shy6873o
dffPqCQb4IKI4aX1MBtCbhBhgkDBecgRgUvuVRk1fRDqBhs+dNi7caBjFsEvINWw
bhhlJ90eQJjjV86UAAdOHid6yfuAUm7tHT6WWSZkwq9ySUh64HQD8Tg7ZK508f/W
XOuG76XAOxT++KZdqCc3NwP5uW3ouTmsn8bNRwXBkCUIXVw/oUbSkw7wHppVsB/A
NcBhbhkp8qZButt8dC5/Ap0sqfABs41xaQLlpQ6vkBQWQBilFv2xUS3EYFIGMJ+a
Kn5AWpYQNJU9rmYnFoegqavftgAdZA0MYawsY4YIro1/eMllqG6gLl+1hEsgfrvD
3nbLdyc4mUCUEAKrwl++CBefdoZ23iwPlt+p/E3/NckzDRi8nOrbqkLJ9y/7w49O
Kjln2egyh8eExUaax3EEzijai0liyZw+7XdwmnNfztR6yASJ8jWvl1w+smumEZHf
KAEhAuMhbGHS8UZ7ApGBIpaOkESixGKWFIUj7jSQR5b39nrcaq0RiexMy2Z5jQUy
43+PB2kXxoN+gysGtPbqyvNlxQaqBuoRrWyZP1Z70SjP1tg8iZUCxsPABK0Bhkdr
IRcehMNcfDvQFZMjBveoSjItcCnshmWLrRGp19DTpmA6mtldzuLzJ0n4BEJLRIRK
fEU3zRI9RfNzMS7/sGQrYoXiou2xbbxrduvtgyDZq5Fusu+JLcKMxgqQ0uW+ox6t
hDEA8yVUiWJDpgr1pEY6hGJ1zrFHpHPv8jtx0F9SD1/A4M0aoVB83ZOytI92wI+o
qQSsRA08dwok+QT5BZ/SznOz/IUXIC+0YxwaR7IwQVCW3JK1Ww9xMtybYIUdCb3n
e6PjPZ254gg0R0L3tAGVr36HPiJvi+5JekHvQyGCnocMfeZZ0M3Iow6f1sRdnnfo
KJ83eKnivzQCG8bGtw9zt9CgDufK3JUp7D3gJbYFG/+NT9mDXfqJ3TqcGVmBOGk4
LPHb0xftaJ/XqAjEW5mwH+7jfGABAR9rm8uQkhVrZG8tX+Wbp+Bzx8M983jPc5xy
ES6MmArkcy+gpfjZSW76XHC1GBvZWFH0k3Hr2aHa1dmTpQAaEAlFnvJ63a1qhLaz
Chc96YKbkhUNOthLkugGubGNRTM5V0m2IhCN8THYtDAzEXdObzyL4oi6xj+SX38N
Y4DQrTUwQ8D0c8Tj+Ho1w/1o/HiTe+jzMLLzM20qexOkNwGOYlTNSvWAnIqy1S15
L0aq+3t7zZYKFDtW0uyJlAgU17X+Hp6Zky/9xhq/SZUZbBg7xVFs7D01sRVReUn4
XAcksf7dHUO+OLw40N4bqy56bZrjb9fod/xabNcybN6c5xyDiLRQxoSc/ddxTXyR
7TnnYtCKmL6UzC5Zrp8yZ8U7F2z3+UmeaX2XI7Et8rLNEp1uNT/HRmDANMxjrQb4
Drit1+8Qy9qIurRHaccRfl4Lgwkkv0wcMHdpQ4wr17HvwFLRRlI0nHLUKpyDbkEw
uYFgsw+lU9gmBgstdDsznvy7D63KhyHwHe1LIYYpx+L6KBPH3KFWptN1gM6v6K+u
g7meQ0eCDgw0PY1xS9HJmHwneGAPzTkfnkaUwrlzpIAhNm8XFb4KHC8XfAB/y+XR
TKeFCgX/wOffQVvekc3vQxaRKPmH1ODa6FYo0695inCDEQHq37DrrDOs61TL1uu0
n+zCitAH5EtqT/biElHJta62zk/CCttzjQy8ilFFgG/+rMMVuPqnXiwkgBRNRofS
h/7587rBMU86KbWx63OdV1046wbHq9Hkn+/mwV1rleRskt4rFNVG4y7okC+7ZUqY
kiNnrwXJIJLxOFQqUBEW+yuBrwv1HvgxR4ssXx+UkUGgcMKaYppdxUM/E3DzWdjw
kIUnkwRoDcVmgnavW6BgkY6Jo+NlWCvz025DkJI8gTIIA/C/0FbXubEuOX7e5siq
O4MBjUy3YsECwdLXXtjNzy2YjiYWxfWsd9BAAUuH8pqopEOUGt9w2/1bWbbamS5d
6/nDz8BTnUfuoIkUIunTSTPHbfGFGZ+SD1SkViR93/yBuvwjmu7ea5s8cseE3hIv
d450DkXMX6ph26CIwL1o61ZyitbgZdWJYJQB/yI0O55aY88WC6EcU2z6GhzjpOUE
gPhGx+9E97GxgVnw6Q7NCaqvlB42/sytFdJklB7rNjZiDJvL68O9UPF6doODYbvX
ZNR/1GhQLWBupl49XZmWbDcTNDmlkvbbqWlj0BRpKy1l5kGNNaBN4coSKRjLMhmu
ibkHWl1DIXF3XUIghemp3gAjSfw44kzSeg95cHtO1mtnNMQH6iRiY9aMQ9qmb58F
UBJ6Ol2CGqp1ipFZttI5ZD7UseuEow1jXpnBjsAE3n9v26Ln5Zp6nHea2JBL5EWq
Pon2FEBSx3LdqbXTo1u25NehXqRjIva+LSbPLt7HLxzS3AsV6wpLnt8RztphJDCh
dyS6mN8COoznii7rYLbAoXnJzXygBP5PKchLncbcvjxi4/nfz0Ann1albp6S2fk9
tsxMpl6U1yyWaeIrWktLj3oqiCv+l1+PZRw2TUm9GmTXp5YryrAjZsmJ4KPUayR1
/pbEQkbiQDdq59PjJ2RmJOorZb0bK31fLnYVRAOBoM1tfLZuAXfjZffgzxoL0wfp
LLz0lb9qLv8E1SQbw6N6GrMQYZbCGrUvtnqvqv732irnge8kQM4W3DWOxaFJXvQe
BANiaZy0qKgTfX6qspXyflkOMTLbLmsrp1pq0b11Jws8elCjOS5YlULTg6y45Sx8
GQrajgwTjXEQ5OIHURLgbwkLD85Zzk9O05JLx+U3PxRNy0hTc/pIpFeWuFnYSbEA
NzR9AyVomRiRu7YmFq1Ae6qsBqi3kfYx0lG9yHsxDJR0pgph4xp2LkI350VJ1/97
sE/XhW/6B8MNxbqCfmqgP/lwi9kDcUhhIxiJzGuHMCGvctkTSV58msCYGkBkx0fO
vQYyx1eRWBQv09hjwro9QHcrPZZHrX9jInAv8h2ZzTdb9ZzhY+S0lGlbc7U9eqcL
LNcFZLLCFb2XZmKHBGuE2HpABGjgD+O2u/kZBGWAmVPz0vC4Ke0jRQK1z9TICz7I
3mU2B61QD7fCLTohYNFB7qTPT49kBdwURNey4I1OIrx9Ch2AdrARNkhJTe4PY221
9AIIbN2YunH9amt2qgoChm6LocbOhc1Wty2VnlXPhPGy3OsdRJB9elz7vj0ygp3a
yUo214N4ypal1tqZrbDKJGYqnVVwlLopPq5Im8MkXLbUc17CMCSZl2poDlqnFXLA
Rp/Wbz6HHtIFOWDgSvzSvRIWk5rPdDeFyNXe8PKKffpKF9GnZ258kkQcp+7c5CNd
fPMuOr+s66sR3jrOuj0X3HToru8dBe7aFEfid4RsJM2/nkkyE5bWWVz3Hlje26Lt
TUocVgtLtDpGIGqfbJcCybPIpFWQpoIGAIC7qtc2BIS4+GBDVP3c4P3q/BPf2Qfl
puwtaFWuHGN2uorF91iDQ7LbBY/dk5x+mXiHJafIc1onQvQPrysPOvb9jkcbmAhZ
bV5tYHh+gUkcYSIUOE/rDtEYpBsl6QFrHdYoTK+bXM0JFtcW6LS2MJlcBXbiuom+
9frWEG0qvHanzGh9YV/x5vKHsYIRPmNOAFxYtGuDb7//igQfO/SbGrsCq4KVGgFI
Yt2eQ71EH5uj9m76oZF4ByrH8E/abhah7xfjicXCYS/yuUinJV6/AY4qeiaOykhg
QurxMfijlQD35vdSCC9zbF+QToWpc/ZfSpAVyJod3LKoGV5kOFX0dQapqaxAw1MK
FWINSL7apcVUQ1NwAo1yxtcgbK5mVMkzxAhU1noam32EA17ntu4ciyudFcOeYjI8
4Eqn+KV9ZQPMCLKNNRdSdYd8FAFCddLH6UVIDzPaDA2mNUdfvvhizRX0pawUG8Iw
gPlgmkePaTG9+jsKPDyYnCdR1EbB64WLh1gS5e61s3XF78EFUmyIJWT5Ek7Yxi4Y
9lNyKB8/vZ7Luj4PFD9fpAcO2OQJ0NOvYGr9fBMDGW57lx12vPTZ3Y99/e8SfkQ1
psF+BoQrYbD/gedFsOVaw44XM8dzpWJSHZq68W9ByZk28hJmG9cM49ODr1c1vpZx
7TaLwEMyOR1jm+iC6aosAbZO/0rmMrxYFbJ1DdVLJ0JBhoiK51jMuWRAzNj3W+Gr
9OToCBS9WAXAxT9Cv2qXcxEmbiBYqxbNOHYpWDF66rpg5rGHQBWRp2XMakdSG6nf
A3hFaA2deb8OhB/f8IiEKODXktaa1pJe6mpcyUreJ31RMRZSvwm7V8R94tGUYspB
a0ehGPRHlEc+tiTHbnsM8gpdzOqTNQfGjg9WcePebXEg8/ZySSfH4gl5fmlfkTEv
0o89KAQ5B0qSwDfyUrHjaEd0i1j/EeU53bnARvLnAlDH3NFwAh493uF/UyRIZp42
wcnt+aSQL9YYQPf6cUo6zZFn7upKFyJSJnx1w5HikTreg+lPpWRxTtkCrLPSVbiL
kKILSHle+SizuuR43aCiiN2blaGe9EZNMVA0rcqhoTOko0KftPuBcIMS6Ntfzm90
oZiGM7tuxJiL7TWb7zPQEFnjyMDkJ5X5af0VqEeG4k+Y8AyMuj8B401ttx2zfBQF
F6wFDJKgyxR0ACBosoB8k/sf4PfJ2f6tlXR/wLEHIxSeNwDs8kjQs9yHMauRZRbB
xgfJUZiIx16l+/QWUoh4GEJfQ06NB9Gb44qG5gB/aYUtsddn5FmO1dWMF+slB37A
ewOqliL1SbSe3IXfgk9sfgvXTEZ1KGyGNj9J07E/oDvO6WHA1L6NeV43n9s33UPQ
F9ujkFIjjv2sDUlG5GtvA/2IL29dEkHCkMpmIKs8wtPmJbY1t3ZenGCskmBlP6Du
rNrrNnQuxg3Ha0ylOgtCLpeemKApDFrnRJFX1ydo+XJwtGDbK+v6XCbsHNQGqfJh
dCBeBHKV/i6LxJuqzlInNC12TcZkcHnzwK7sKTR9M0xMpY8WvzeCSHnaBwjoSTed
aP0I6VpHY1v4d5gMEAwu0SrU1QF2PEDx+VycN/cS7k+NDgczfaAAq3Z7Nhdik8Lo
fm8iZXYaWRXGOoTf51Yp7wGP7C0agatqlWREUjB/m+OXymyvUWqRLlmiQ71Ndsoq
+BL75r+n3/eTu7sKwl2ap+FQZKNRJyJdXBZsc4vG3saCVWsM0wkJNPksA+F+WNuZ
3htJp80Mso8MoZNgYx/gR7AlMPF4g7fOIve7EnxTfjKpSzvDawtcfB1jfccZtWbA
tFGplU7c21GPEoJj3z1zzMMHOTaoD3/ZnyaavYEaln3FoMhzduSJb8Z/r6Y90iWe
XEEOEGjDx+ZMJQkhJOXXiQlHgXw4g4P3TFUctzgtJT02zwJ/FGLLFg5C2QjcIO/M
3NXDkDy+lwEDuCvvY91XrMKGB3thV59dkIkT1aS2lvzQCcYpZgSomH/ODM/pc+aW
mCe2EyPVxgIrhOlyRp5fKFPE4FV0uP3ISAa7qpAnW7XoiwCDGJZ5nl2+DJ4REArz
lDB9Zx7vVDJTGBB8s+M4wpou0DCUHXBq5YEe23FAIFkPmqSzjg7Q5sI7WCAbi80B
jTFIbtVUs1gtSUmpOJMi2QY7+cn3FXJfzG1WIPWsuI9A9QqWBMm0NXicFczjVfrF
4eP6CA6zfqpaX/Yz8Il21UzGF9Av23izFzny7UUxTg4vqDKi+eulC+CcEW/fsqLa
UMG6dz7HW+AjDIXfD9uPqqbbtY1P3vwUzLyxqQ2mozk8oJ2dsgM4GC4odzFkQONx
QIhCuIJYr0MlL5kT03HpJO7GAk2Fg4s5A3dUToQkyRw3fQTE9v0zTfwqkcrx3Hhl
zCLIsbEFo95v40xbBcZGVfkfkQwsF3sud2kw0uKcFvV91wbYtX8tjGf5j2GtUvLB
PUSeDynZIcQffwZ2VoHFhH3CbAfoQiDxbjAsbuheSrb8vL0e8w6LICQfdLC+ECpn
d4b81MExHknKys4KGqE3UzN8tbhUpev79ReaRWtihZAvM/pQBRKmpTIBTwn0klUA
oYgTeG2L/Rj8sSlP9kZMzTBDQ11CeLhTasJpEooRT9Tx7Wz3nRQS7rzlt1lF27/W
T1bTA5n7fG196fbbwyMr+8ts2quxaE6TiBwjTao39cezvx9M01etos16wJ9ee0hU
mOksXvhCYw2mJIMwINqbxWpy6w8ySwtLPaxPMZezZ/suthvsQafJ1ttr/PlZlrnn
LsjJlkN4UCWnBEor7w5ySVxfGAB8xH/c0Fegq64k71uzbqgYTtr/ZGm+LLT4xo+w
KdaElaD33puRhKuGv1K4KLEe51MSfKsZ4SCHKWhMGSYQAtn/G/IJ0auNGsuWimKa
kV3ciLwf2BM9AOf/vnAYCgIYAzH3mk1y9l38h9mvnNDx+zrgL3YaR2uHmLPs/8gq
cAEVUAq1lFfALCUgiivug0D4bHNjko/APY+1Jh7iAQfnIjgAAxGexf/lEgy7wSap
uX2hb0xg4P5q8wzOdasGDqLysyTn3x0e32XpfSyJkJqWdo94YKvn/yBWr2FhIQjV
T5k/8rPtg6U7aH2phkBJLvbrIbf18sJETsDw4RmhvPlv9q9v6EqKWkN7RqMIgjj4
oYJXcQOd7wnXOGFkQYQ2xQEUcRD4KJH8pLFnB0hqfTIpG38sS4c39hwrVksUMoY1
bgxTmYR04EPZjBYFOJSco47ZCBePr5di3XPtQWWJNKkDQ4+Bg0xSvDk7o0g2yn6t
0NqOtz8mwkCQCzEjACDgtDu6szVzCoqIXzkQZS6iNCJ2wWPWeZQ2hwCS9MUEgHvY
x3XF7KsTrj/tOwM2UYt/x81xlynoNdOpIoYljrcC2mPJBf34LwjuQkkhGwnDZ4bi
oEPnSqUCR5wzj7OiMTkaIf8OY6qKMeF3dZ1t3moTPTatV+eu2uJyBGl9oVH6WE1N
lMlb6go42Lk37lIaGSeWYmuwINFKjUehCQ2pR/53bkNjcVR6bfOiMU578YXp6+cm
N2UoUZlLB2A+e/ePdsdKXKcqDq5iUPT+eyDjWtoln2aAIW5nLMti2FWvH4W+L/p8
JDDWaaCMUu6CnsVXDbozzL/tZ8vqrZDdJlFc18zToSPN82nPohybRJqT0+VmDjC7
cpAJxvnHVmDRRsIA8Cf80dT4zkan5LRsRJKRP5NaGsDZZTKSL686O+9OAvFDhU/U
2rhUVh3pHAJLw4bMTVrOVySMTVut5bCU2xo0kMDHjlfTrSUMbnqrqh6bLhdOd4+Q
QLT2AwTZphUc24x3IXmhNL1nCVEocfekgaGPaZdDRDlYMniPHwqZvJd8OHeHnNKE
nuVgiTc3nFfDM/Ag+vCDjMkq5l6iJok8k50H6+O75PfgA57YgPm6iEtJ5pdc7qaT
SWOATpM8YVWAs6lUROdd2nSxd3VLtUlt03brBKMRqO8K5LYgpiQf/g4IlzEqWXzC
ISUjZZkWITQvh7PBmKAV+02fotJc5R6TcIY7cwEksDMzy44Y80H/0Uo19E6zvmXL
F8hkEt9De0IQ0kEeEjTRn8xOnfoVy2/lDNc8LwdLX0ex98miUwxCfA1jJOi+raxV
o7RwJOXwmT/rFJbx9GFGyzV8BDHFfdxbnUh5Ew/TeKuaUj3BIRPIQHd5o3rjcxT+
RzxMwJOaiZRawShLGyhB8dNL9lcMINojhJzfsjVWwPo4d5kEAqx8hZPEc51XNz5v
NDQGTO/TT4xM5fCBVj686LG8Ed3V+bVGEPhku8Q3vgPEqnIoC2S0rqM2NU07UsOX
F2FZK+rIvheVgn+qBCPaMR86yOuEufTQutQAnqGkL7VxLfy75HYiIUIQrukw3qL+
KjZP1lVGF8tmrfI4fQQZ0mQx+AMXrlryID1X2sUD2RzsiZJjm4FpBLEpIyIOk1Zl
L4VBgIYCysM8grXJ5bC/T+IbOUd+iI1AdMhha/xgbyb6zryQ0pczAsd0wrm3ZC50
vzJUtPq0vYZ2IXL4ffpfrwi2m1JUlU1LFp+FLNPMQIlO+tpCFFduIqjhplgBnTKG
wfPhhGtt7yFw3WDm5pPe+cSoJRN90gIImOtvZYhfIaqOzM68lNclUFUaMej2U900
8BrRJiDTpehsQ/fRXYRGFxQi+pboKaYX+s7Y3KuQ9O4msUMi9JQm0Zew3OIvqyZL
BFiZcvBZDWYWIh8rQUyS7OMEG44cKT/wKL0VIPL1EoCdYJQdB5Q+9msh9qFYFW8f
e8a+HgWficfci+bGeDav0gBE9kZjz68h4It/yevD4m0Jk+Z5n7LCKFxrAbCXIrWq
DefciSflW3KlazhQXUbgTaj4lviJqZlWBFiq4Gbx/bocUQpfLJjjN86PPlDlTCcS
mWKZ4GBj7G6Ggi30E0OtrbvmA/aU3NfQ/X7lgl4Duq33ciuSaPEFybeKu7J4AJ9y
renkQJhATHlVQSg0UDZ0vF8lcaHyxviQ7SRcB24uLOnfpNI9soM6eE66LRejB/sF
PUQxMMN5CuL7gyGNDDe2e4SggidjyHco1mG4qCkY055av9n+BCXgjz0aMjhuNBT8
x9+0pCbO9gbHJ+B9KmkhHw5NiK/MnWYLOhhkamxQRRotz2p1wbn1t/l5O13554Ts
7kx2sUFkYf76hth3rFafugMJ+/NF0YDAL8NYtcM1Zjo2Lluy+pgYnPR3pnGrtkfG
vuF/OaNwep+RF5KVrxI5HIGFbFfJeJegTSdY/iIjcZWrQ2t6m5vRfOHVShXMIkVl
VYubF3bQNRESJxinzI8zxPvg6POvBApkpHZNAaZhF2aElBP3mKiff/4xyGv4hrww
PYgXH5Ftz0/aRJ6kH1DDjOnhGp0WQAGOQTeFbjNHX/qqN0gyw3sXFMC/X9Dwh2os
qr9C2/K/UySyo8QHa0f3OnBSuTXxrE6gzdwPSzS73t7t4SOcDlfpWpuRS7AZ0bp4
vt849VThJJfWWaso2hskb8XlrPdiWRE4UIQjXr+673UVPmwNxkR23mhaFK63hIIY
5oIl7m8/co0QJB3RwXZsx0IuK83MJZSdpXCSoo50wLyUkuLF+WpxNIAB/qEKF72n
oG3ZTIhjp9HSHr50J+BlWlQ6e0b6+F5wkm1WbBJY/lIM3E4OmdN8rIiMahIAn2lS
zYqw07gGS5zCufYTQHlKw8FQWBbQaXCWr0KGYJFzbjoydeVAoCG9uWHhT/h8sfvy
Gh70GxMH+yg6XqnqFP8xylXK+CSGf6/7qyT2HjieqFTN5OuozB3IbLqN/Uv8OTyi
4bGUwN4BrIbVBapsWxUW111uouwjccl2FakA8VEqQxJxFpPujrB5E/onQtfyg+mz
ad9E6nkBJtKiYmipUJflY+/OSNxhs6IqQaaE3GmUiZnoe0OR2PN6Q7bmXPKfcmLO
b68xXqFBops2MQ2kgGKuklIvr1iWF2XIcPHG7v41vZdT+gm7hTIO2yJJMYMBOtQx
MJ5Ca7QTJU66nIU+hsPJ9Wye3yKRcyoMF9Ae/INYzS/NALYr16k5/7kgnNrPke3b
fXQxozjlPF8AjvEOeKPnuEg+y4ZBwp2zyLVz6ARO4gobClj9qRplODCj2ZIGKePZ
ctfYnTjEF4ZipmsJQ8hJYdjg9koUqt0KECO298ZtBzl0yMFZJWlXqaBkdhVeQx6p
C+dCgoasGwKHY9OwLCqfmZhqxg9VoLGNqad9TNdny8Osqr3yKnqGCR2+puDRPV77
SVdwq5gV+qtlljxSdMo/FD1LR2jugIQOszvM5UHxAjrtR514yyJ6Lks4589/ve4N
wnh2rv9LnXHlyR3BikFmW4pDrGCDV91U7N7yF5nlMculmipMX5dA+QNSBH1GdZ+s
x2itjC/cr5kEREL0ooDGXze9z1oQ1zsM+ZqT3UGICy65qRCF4ZS5JbYj8vnixCdP
Yq9YGOtkXLU0qBUulMCwfYvNT67cnqkbdDYwRHaUSJhpR+MkOfNpRIQZ5pZqYTDQ
FnHf/Gd8YyK0A487LZ+7DjJxfunRd3uLc6xSOq1llgvssEa4pbZW/7Ufx4HmdPdr
8dqCk8e57nCs7zZuDdq90CuqfODNrf8MLgytdZSxkreizzWkQJ/2N4TL1oqwIiK2
B8PKFyICq+4x/2cPp85tEbgjdDS884r2JxxfInffDQYxPK6lzz+fuABdbBWll8cx
z6j04URGFoVqEuqmpVBVMmnIVSiwHLydWB82lmR+Z9vXCtmUJORi4G5aPUX34zv/
puBued37aXeA2liG5a1A+yCwlSaeoWIcXhG7nua9kdKPYDAs4942kBM/K0pMnqAT
epz84UW6QgKiaepEbTqzTFp5iT1k66WX6vATJ/81cs8KwLZklrCmOrf3hJaJcplb
m2H/evpu5iabqWmMJ0zcFxvbCtt+oj2w1D4LAdVCWeGj6bolBd0pyBCnVBIIjtvw
JMggQkh95cLkZcipvr3OwrUgyxvT1wABaghCSYDQTjfHo3EopnBtcR94H7ivA6XF
Nn7eGMycuOUwxgCbBtkX4vp1JK27kNmdGDAs+L1g8ptqFareoXU+phyG0FM+NkOB
rCbYGDErvaWEWDQPCZNoAOu/IKRR1A+DOUYh1H/7CakxKpOJwd6C0xaJWFUd7zSv
ogfA/8S0c7IAVJ8yqwGwZ3h6jxJ1ohFupqFdxeHiioejwcKd4RTBjysbmDE2ioze
VDgO3ucY42kJVLAapwRDY60MOFY4q9XrGihRIHguj5H8dokFti/efFJcMfniua9g
Pn6zX2V/zK+trIUxGDXSpCqvGoL+3RqDU6+IEvP7Gw8Ixwub8Rvh/J05vr9r2IFP
6d3FMKb0cxX11MplqINIZ2S77xGRhBd5HpGSfIp6H7TCi5LmgjnibZZDiSyb3JCL
KdUDAmQSDLGulHCviVvQd+a/rulm1bElUPbNUg8JLzhYva+H+wm7mehGH8iWEpIU
vxmRt+MgLB+XQEAwEDvkYr1H/fuicGe+cAg2qf0fTGZzw7h8ZY+z5WjJNKwoTULh
18oUluQ5IzziF0fT6L1o/SY3I0KpISd+xLQO1SAl2/vkH6vuA2FwZxg/9VflLHFt
1lJ1muoJJbY/iFpgNMlIGn2HF9Zu44NMvTU1M0cL9d+0G8YzuvctpazTxpOlnjeZ
mUCylNz5bFO5jndntDRgDdx4aWzP5OcnPHDcPYuimRupED1v8jtFxhzRjrmZMh3q
yPpeWVP95+hAD/YEOhIeilwnXh6Rw9zlCQhuVtzkB4qkhWc+FLOlCJXodm790xgK
y+8kIN4WpxSJidtzdE85jm95c7qoZC4bjejNRekG7fHvYagQjveCfClPSWhLRxD6
lqP2C6/z2yJ3UM7qWvv97297+tWSgy2dUPSMCEsXOHUBq6gOfhfUjmEYDM+2Wdfn
B+nnoNAT3o+cLLGNsFPhPPbckydmaXO4sb77WOQmlv6boTaK5G7w/cEFwPboObVm
YwID/sRj9Qm/v/iTnLEXa55klqiSRhEVBENfmwTVVC+DBNmKE9jt74CxyEb52lUf
ipndUieMoqSmN7xI9dM+mDNGiqQDcOBdvtH5nWOTEKB8X6dOlY/gzIRKYb8M4Fjn
yRmxcDEnsiwqFE6lZEyCpkpEDJPbEnaTlks1N65DA/mh3D/2DfS/IxiEsIjGPjVg
8gLrUDxdTGcsZcAdQc3tjjtig9nyMs3QLJQeomzBkNaK7HPMTsoM1+0zPi5uTwMu
dJf8UW4tf6t6I8PFW+hqqx9A0GO/RN5r1aCTzIUeMRrdx82mdnXLeMFtfxL2K9CG
bG3RZ2+i0WwLpvpbrVpdZqdXFz6X02DF8VWbSeVYIAXoYoMEwuUT0Jxsppq1vFAm
8cXSozFbgJi0clW+A/agI0VYmUtQ/nQ7CC+4wzqNGSG246U5wu7oH1AnDSfx68E/
yxt1DYr6TvXKQLdzTtVeWCHOfWKFyCECVY1sD2Z/crDrakXD93RC1L5Xf4XJ8rRD
DIVa7uGflouxRYzlNfkoxTmNrlfphGy4rid+EG6r79N4vRH3+AOCOdfFPB5IZ20W
hUdAKXYZRrm8tZYfkzarzz0Pr3aPcTcolVPYKsLiQ3K8L9Up2N2wj5Q+CHB7xcxo
Xvh1OwZTcUNIREDFCq3xn74xrU4tskiIG1j/fQOUi6qb9/Hr6HRUf7bsoumPJTiG
GgD8TITSB9dPSvFBcj2+f5TNb7OjS/8KChzdz0O2jslxHOyJnfyeAegUJ/IpPq3b
mAZEIdaxrvYr8SE1JdT9jBDaiA9yRsBTGEft2rF8zaZhNzkHWECyBxEeNkJr2Adn
1DRNr+OlRSTpr0Vxe5IVkltJn39mdRBO5IlqPoXUVqs0OGEawoJgZ50482xS9FIC
ooVOuy5im7zTb1NyQxxXam+g7PBDN307zbz16Njw+JpxNmOvOLUthOaLJpVvDSNP
CrlZrgMMroxOBn384iVELjwtz3MRX3QuOjbkZ2mq90H1CYG9WnCTYJkQaqhtOxjJ
PNMDDgr5dvbL6rwehfQP2rWwO5ONs8z4VypvoJWDIaPq033jlkC1I4JeRT9tQRba
0Z17pdxCXjtXyOXz/d3mYsCtF0Bf+zWffzgfFSK07n3sZQ8Z1wr92qk3fvEJ1KZS
UkN59LtG2KUGH3QciT06/Hs0L09pUf6EGM5ZFRCXIBdDrLeBBpsrVuNorNirqWCI
oArqiQR9T+dtjekwEN+5/UI9Ug1Nh0ez3rrFTqyOxeyQwAAUbdnB6QHJipc708fC
WYiBQt+MGB/tgQOOntl95C4PIyUpsHC/5i9d/rsQBYP1GQnkTIn+0/A85h/5KCl6
B+m6TIwySv5cOBSyq6LQYZN7tonGW+UZ/aKZRbWJY1yG1JsiGQr5cT57oCwj3lcf
MwnxEDOCztSUPsCwt7rl/+WAm5n5mFhPV9pkB2ufCYqGl/IevNAyo4zE3IFWvdFt
CxKdBo3B2P3pw2+fEC9rI5wNbZYBaVdaQ1Yzn03jF9zyK12DEmyfgcdSdDWFqrxt
1/ny2fu30+g/LVQ4qC7pytMhctPbqe40agzDqMYQDRpJcZWIaiK+Zewrx1wZzmH+
+K429bd6li/y89U0SSlXiPlc5yMnoHy4A6mDDZtnhv2MqIHgRdg4nDVv+YXR183m
CUALsIviIHasmAYldoB9XinXwujl6V67CGUtMKw9fyOgqY8qprP059XcMGpilIOB
6N3bW1yzLX/6iPMVlb2ksXOJo1nGLkwIq+ffleNI7rNsJxVVykFoAYyryNOskfmL
w85hRyuKEzFO6Xga6lBH1BwE9YTPuCqK+HNDcRxSNXeDP6h3UP/BTtocpt8djc7c
iAqjrDo9AWmfaoGGFzMK1zINqj6a8IfbXWjU5TAso0j5ioUmhsXkKrzupa8fjtc1
yLnb8tTbFMdq2jESkutsoGPMbewmrlotq8KTHHLDQEBYzP18HSO1kYNfOkrqQJ8o
Zkg18Ggd2GLIKjVuLZUtaYWb2/JmUBPmlkK9ul938O1+dZes59nXlnjoa+DPNok/
gvCMz7bZcXV5lGJgGwOOu4I9Gw9rvQDxkxGnPebhRjbmVmV3RTGL+qez8xHjLSR2
Z+dHh/qAtj57UugpGxTFA7FtcEgBLq4Dl72lUHA6IPCoAEP0PW8OaasGzdt5qq0x
B00twgjaU8itBV0iaOhz+gHLdo+kfV/7LZNKPgFXFnNN90ZOtAOy5oceCaJhgzvH
1yBDcsV8zIwmZK/bAo/uACtaMfnnKZ7WDXTGqCEkzUL2TJh1lVxzb6ex9bZkOSgk
IRgVElam7mJrCuBLYiFoQB11/hriEA+eIYt0v0KIPiUQX3cT/JmyImIHLfX9rA2V
8AwW0PX6pTPQsLm7VQ4P8bsKnFiXCjhvoRXbau2hqNMPlg4qbYis++aiEfGADK1b
6MKBxFajmDL84JKVIKMLi5RoHMN0tbSV2bU5dhKFeIcGd09PyIj2sMcFBEaE0jFI
C5+n/YRLByY9o/lVCnBT6iPYz4V2shdjYNoI4w4R3b6j8uUCnme2D8Bj7jjuHMlF
z1nWFXwC/XT+QHjQO81/dMm6A2BhfL2HuqhGHqVtXrxUns5QWS3Ub/dJVt1g3CW4
mWPZWnM0f7bTXE3sVd+PYjpjKT4MqSYbLR32YTz2VP1J+sJt4+WhAWis35WdCblc
5o2P3Uph7HRTvksfok0Qno2Mg2GYfV4kLiy4x+iKmd6OyC3qm0ryp5uZbo+qZFoy
CmQszse1f9Z8Gr39IHACI1gXGyKmAxplfnawiDUOWRByq3Xx2tnhMcE432Fc3A8O
jlvFD3JBF78ePgYKvqHaEmerBQhNdP4h/7Ix7cEarIYZ851XhHlVN9eKhwvPXXsL
nQWKdNVSQHo6TAY8M7dSFb/K6c5WaZClxxYTaEKZB4sqRhlY/9cRdZN/hjpRo7UR
nIzM98rVaJPujYTQPqWtp+JaHXtpeL4zCKNii+gIAr5mVOIZoSqnXFD12hxcaeNL
8AhaxIbntZqSEXNnNu371EiN3l9NCGBmvsSpYmZLXcAlfosXHgCFeVZHlV9t0NsM
ClTeFvnam8Viol2uh8NgaUgn52mAm4kPN3r7a4VG8nCjhCpK+6hD2Y65h37xBRNJ
YZNiR6HpEubutdXL5H0ziXnv9Z3FcSICLUv0kdy7zB1W/M+ttPWYhEw8ROwqogDN
9qNB1r5iw9aaRrb8mASGb7x2Y160m8QrcnRL1uudShVK9ZjEWRapo1iWOWluoNRa
7cMl6VdSBf+jFUG+Ndyjb4Kzll4blzs3cbMlKc7mIlzAIIQwn3oYmbTyVneQsbEP
qInxxOOfX1Oi51NIKbQDyHtjsZZQjcPm6fK6aC/Sa+ShFWDh+NZNYYjC1Jb3kL+w
TM0uB/Vq88tHDBhpOsu5WzpoAApRIJIVYVXPOpMFa67rW38Ip13EeIOJpET3UC6z
7D6+utjf6daJGBVzoyxTfHlWZyuUgd5g0hyFfeAttF8g26dKnPbZPoKC63k3bxB7
2f5U8epFrZmA6CFrnX5dBH9HkAbdlQJ2b5B/zVVz3JhbTIXVK1Qajcfm2vOQpd+E
b9iWyayaf2apO6Je14/QkJNzpxs77vRnTtyZJicgaFgV42isNcgtxj9eIySBPRwh
e+IsUxM53oCFv0EyVgFYvfYE4JN+qzLfsFVJhr1znNhbhuTVKJizEMiY4yjd5ySZ
BpjMCO9FyLiMiiHvaSiVcfE9ox+HYyKiAbG8+qLDRIVaq4BmKMojtt2krerMY8mo
tXISJKXRity8xkqgL/Kkc/W/TjIdrZ8IDDpmAJm6toxkjHxvKFvNDQ3Hvi7poUfX
cqUW6vuwyDgNYSV6oUp/oBdTnFzBbifqa2lNAaakH2BE9Tr+AIAUcrXJ2SYhgJkt
P1oG46Hls6NChU5MmUA31AA/RPFhmqpUn3vsi4IR7RuHWhcThE5/q/sB4grvpfC1
UxZXmnG8NbWnuiUlS53Kj7LcHMLQYqLTiRztjgrPSsblYgbd/DIb5qjqDAaXgjvB
lOWZWoLR7RVaaA1kdiEGKkSUMtMx2Vfo7R5QnjdKtF7STATxcp2WEMkH/wss2h+X
Xlp21dRnEZe+tb2LlsXyJm+1ZL4dD0vf3qqtUWsDdSOBy8/UEBrrpR7gGWnf3Mx1
SmUeYXpElzi1O6wsjZ4HYcy4j/WSy/gtIuO2NDTZq8WK4GPOa7RjKTIXwyAescZS
lU6/gOmsfd9l7KXIf68xXOWCLXLBBSp1DPcIoXRA9PTbZhDDZ2mA3dRlBuVV6GQq
CsXG1cqvQyPtOu02GycLV2lSaqUJj9P5RtCtgiqAtHHn6GpOOzO9vrE2hEPaF6n+
Spb+QwiVdu9NswzK4DxxD5VwpPcKWyYFzaKMzXplfhZPDccsPV6LtwrL1WV/AYga
uamW2FEtkmmxlSPyUH4BtmR6sKSeKJZetBc8t26PPv+m7ZmUoW+mzwl8Nu8Fm0XI
+981SfoRG8p2J3wFH8aNHQv0xhtkfMmceBobQsMIh1bKB28UxfFssrWtOFVPQJ4h
GrazElt3g63mjwKYzfHkSZjcf1BBo5Mn+Fc0Nq4cLWe5tFFeFSJCu8AfkwE8Ak1x
nXxjdN90Z0LynAha2hgbpfjyIXo2Tf8CLzmoIgI+AvMGNbO5c9yq0TKXY9WKrVOT
P0ILKjLKDFMdnVtjTYXn05QVC5d4iMUWe9/DCLQDz58VgVGNVyMzDdVCgUn3yO+7
TS7771qCRRm6Qa1wcFVCRACeZ2i8MiKSUaBYMaWknAxlxez+CrXGnWkSbG787m8u
mA1VUuroT26UDMBz1bQVJSQyqlmSBJfUHKDtTUbpOxmlmXdJEP54QE1NbQeI+Esc
nskHIQrT1biXO4FDJr0K1Z8ZlOXGJKgMUNrIveKsWkkcCM0CE5wmJKlQgVVU1ExH
JM2mcthl12lCwj6N6pK5osNfuP5vQpOnh8isoHMRMW3IH4msQeIJ3eh31dZbDiQ3
YqxphnSQH+J0ZsIuJZSNsdWvGvV6tbNgZfjB+d2QZYqlBb+0RjigG5rtKHE5M0Y6
abMD92INjHJt5aa+SeThzdK815+pGy4dCH7e3CUfV8SgCbyFd97Un/gL7uSTY8GJ
//lR8zCONLOWFQLHKB3aZAeihVT/yd65R/77PXFexQuoznVzvY7FlWbMybp8dK24
7R8PrU97cie6phwqmtrTRghlsHabdY6qXN4fCctWkBE7NyXU6oib8x2q0Sa1RTaW
5mr0tKJdDLoKVfsO9k9V/kYMMkgCB2FjnkGGlv4EF1nGNRb26qPSVDS1hsHb/Cd9
lisKbElbCXiPNkEzxz6mUmR11397ouuNoxagtheiaHwCLcptGm35v+1DENJW6HCs
QFLBIhrsqZF2eZAxHrjrSxfQXTjbRx7c78YGvHoyfYrYSAdV68Ko1JI/pD86tiAH
gxIInQuuDvTO5qZXep2jwJxzHBbi8/VDqkgELjtWt9YiEgD7bCzjukCiIFn8xMgq
tcg/XGcXssOeCG5AITo//f9OxhvwmrHr2A51S4eSqUom2LLia5pQKohnpHvC6wsg
/IZxJNL1mqJNdv6SBpfywZ44OgVYd08iDSuT/cmL3fBIdRYNmOXiZNQXQ9I+jtXw
W0Z6hGBWpurKpFMg8o5kdRJeWop39B1M+V1z+Ma4IbM=
`protect END_PROTECTED
