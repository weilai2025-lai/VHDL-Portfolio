`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tewRc6Tggcj9BYGUvJYKHIz9UeFTyRX58joNKlALKitsSa74LdWPbgX2JLFk24IK
9MSyBhRsLGQDaCiP5K6ajgzX6z6MwyDphqQfYv589MhHblDPkCJkNwCWVvsj/10M
J/JA+Mrhkbq/ow4s5sv65oRTuir986UEC1X5CWV81EHHdlRo6yaWA0bYVza33TcZ
5S8seEpUL7JQF3zeOAJNDeZP59Atq5tRwziwC0vlRMH/bv6oTJctJy+OXv4uPN1s
GUBX3kPAhhI+hGkmjMJ4U6G0XxKIIhGFVMbar+Z16WARRSobxX5khqTPsMnimZ+i
GBfOHa675tIAt8A3Ai5CT7lRFli00ylXZhuRKHYMgrCQY/mS+KDT3qDuMRXeZBD2
DuSzWDWScqb1aHGe7O1FhXwSyRVR0xJOAnjpA3Ip02TrtBTFIbQHzi/z8I8DrnV4
Imv2+fVKinvfcemrjMkqSrOK0UfYItbnKDdQvXWL7N4I4PcGPiZn5YnUKP32Xe/Y
SqojJWmGQ1N2bAr4j7z+txdGetq8iRVXzu1+EUPrw2h/pG4p5V2XUQpwA9LhxWzm
NizPKDhFsPUh98Pu2Gj1tXgjvK7f3sbrrK2ocgThFbE06WhZZXRujSxiF6xw1BMx
bNcc8K0uHE/PLLKb3IInwagpsHG/QmzQxhaK23IujVa/p1jQQyBRruhz7PM68/Ab
7Jj08TBWVe4IrfnZmab65GloF0QsKM0Z3PtQPUAXmgO6qBRzqN6CGmoAFG9KS2+U
Zk94BcWqCSo4s8S31aUwPbj7+OV/Sj5mlRbtGpZWGVA3/AahIu7bshsWSjNsXBPi
PDJuhmSJHFZoqeCM4lW2tBjxAu6WKo7OoWBmWFUNZxZaFinJG5gWJNXhApdTzEwc
3GnavC9pr+/GAIZOHyoY8DDLULSegq87lwB4G2zx4rSf4TM2uUyZUzCVloEuSKDK
gdRSErWHPfWHl0deIRdltltpwDR2Mu/pKA5x/gBamGysZuEEv1u0mAerv6ZhNAE/
71gYqZ27KU4e0RVR6aVC6zCAjy/TscUcXSALMG18DL0MEp25N+OW1r9/OlpLRCge
FAyPzNZbkNtCDEO6rv4FSBxeVEiOWxnesC4cCtcOYhB33PthuEdE5+/zvtR8kHlO
KOgliIqz6ED3hvVasg/FjmckUtKFbHyGWwA4xWnXfLDWTJGC6L8zI82WTwxMkaVV
v7YItr/Ao3Alwj7wdUJVbCMhiRkFlf8T9e2d50gzvn560rEYgu+12qFXZdqul/QX
5D2r1pUuU8IlU9Tqv0hGWGt/sHcXzpuq7lKBgK9A4Hfl73OAyuSUF9NCFrls5f+L
8M7dnQS237y2Rbb4ACZBEJakFOKvJSuSmVi8dYSHULe6og3Gtrh5n4b9cxXy87VB
1dgmfR4fM1SZcHcMUUNMicdGDR4tyxzyuKs/salyRWENDObYDpu4l/cR9ABs6ukx
lXtek0L/EoOfjPHgb2iKgLcWBsk+KakZ6Ufu9vqD3Fy46W7HwqkyK47n2vgDDM5J
9O3Lkuat6ZImhPYjh6zNIQXvdnqPg3hYBkn5iU6ol9xsOnZMGwiKIw+XzzDnkLoC
innfPL5q75+Ue+P7LHupIRgwbpbQQoPG2tdkJFeGJV7+2swC+TOn2AskrTY5rBQM
InhdU1IHYQ5CeuUzGZ+K0owsvQHO83lsUHAeh0Q/2tFA3kelz4sjlPMInmGSjuBn
nC1ApXDrsTTrCyTF80c8lHoUPkXvjHXUbOwmEdXyEqW8qFXruGUYZUqe0AD2l3Hi
f3k1HU0nTTsnWjdnTn8q12FJExOwi7YpPC++rD9Q8kdGaxWgF0LIza5Sbvlc0H+t
hi+tYYN8TQH++msN7IShAYMUAsX3e/Q8DuN7vkUvDAPTXiPAAF84JoqPd6W0YhgH
cM/h8lYU6MLD3GMOQbBVlpAT6Ux8XpV9/JwQ1uCRGOTWSEWw77ZQWo8l3hf1HR1x
46aS26I3nM8LFB1lHA4qEkwMWSSh6Dq/XYMnOE2OKMb5mz+YCRxWiCiAVtYiCW4X
fmTC/WA4yUkdvIC1ioujH7Q98SK27T6lTrp+mP1vyqx5ezT7GlbAOdwXtv5/Pf0i
xE96NqW3arTHSZFF8TsYg3kxilhji18jHFUbtx+SYOSkdeh/sE+miHJHvMNnC+CX
0vBKP2jtjbXLg1bm1EOpari21VoSSQy4LDMKrtr+oWu2MP+stOAXQQUm0/CDq7dt
EGDPsz0OqO7uxPNY6P712lYOj5cIh7OAugeSxWEsEk5t4U7O3Vq2V2Lj02UlHa/k
bHuU3rctQNPwMbZ1eWd1AsxNkMqDYfBhi07tKMG3P7MWAWhlNVRprjb1bzgtCJWB
Jbiu2aenA5sWm+jBpNsf0SmnNlmbq1VeUUjexB042EeHyh7c31g1bzhG8M6FR/s8
tQhbk+rqPiXh/z9Agjcaa2zy3a6mgi2wTKLi23bvJDbVv8JG3ITTNe7UCFzAQmID
bwGUIcghQ1VxIT5sPH/IpQgXD7rtWIGR1DS5nWDZqmBlERt77ZXtqdmpC9xOc97e
Mc3JasyLZ0U8OBqpd4eC8aQEnZeda6wwSrwu6DWvpEZ9jrIHAquIaKvMdyIs3vcC
Z1cXFWOjrbV4iFACKUozYjE00vVcjY2Fsr+edZWdiXiey3o5ycoBTHiHCmTbd0px
XEtHcczAEPU9erLTfRwWGx96jPH1huEoEAe1QZposZ8cNYr3VviiQhRAlSy0aEDO
+kEDg3I1tN1IX5jmOI3y425V1Mn6O79wG90v95xYLb5vaTco2O2Na9JSJVZC7UqQ
XOr8yd0Ms5MtAngK6eu0D4w/7T1+5vtBFf5ybv9dHNTt3KdKstyVyndQrpT3MZwj
Vo8ZMgAbLYf6SKLiH5d2Jr+PokAkdfGUXVYNLVBuC3Bb9oxpr4uElbFik/xVQz94
zMLkKPEUtK4frZzUCuSFWzR4fYuAxcSrOgKBk7nhfVcjnodTUGKiEKz/vbfodjC5
WxzO6NOifuSMmK4raKGxvtDoZrdWy6wmPDf+EilZOUB7X3hG7dhG57T1O4Em7Oz/
LfbAVnb2B/LNWPQKJHaTunHG0wWHScOJQP9uSkpjmDqbTR1qsbouKGBer+76dxCc
GxUYumoVqVmeIo61MGbUIW2UCt7xfhmJZxKxEUFf+0M1wfD22RZQdFNr4jKeM+b4
ZXveomOBy3NIMnEyDZFI9O2BYVkwfgI6BCq2UeJx/lFa5tdSm0j7bUWWwhHrgHrv
Uo3st2D73Y/alZOyLzxSpa4ELkjc83P+vIWCGSnEz2TLeLnky8l7ut82hQ8Jib1g
OLO9uTlwnefI1tfzk0l5QwKASyxAttPxp3zl7qWIHCzwAmuHA4V6G4zR8Dtgs8mv
RzPbgqCnQdfdZYpXnsfEh+9rQTYrO6oXHRU7GaYADp2zUEmrRazARHR/8gJDqtx0
cgx66JPU6ybvxcN6bjWI1lATdIjCUvOCi1JnIbipcnskUnlGkXgaVzG2jwQdQpin
e7esKuGdAHkWC5DX6kV/sc5fPJ/UWu0fMVbZNxXvH3OiDmoxowL0+nNlAGOjWtH6
29Zol1YLySHk31ZozkSQ7Y8wLM1Mo+cUshFagyYmYgFbPL/vqjiQ0LXl3ceWVAQK
jxaji+FbCaXBJinSvLquvM40iOmSew5SwpOahlFCUGthR7r2ZQQEcXCaEZvk3tr6
ohSqXonzn9ksL6Ijss+SzeEEEj23Vgo2ssHO7R0mEkaiUkEK39juQHOC6IDW7ufr
uZtYMbmBldaW05CLLoDoI/c0XjBXSk5KhbFrsRvBljTWL1WVFW8fCkAnyWCPbMbn
QF3843Ypu2/A8NFRvi+cPxsU5oCmMnvLAXeBExJtdpcNCZWtIT70eEZAI0aA0WG/
t51cIJdNeGWcEdU0IAw3II1/9n9XofNk5NJZ2FaTkvtl0k0LtTJeMIUX99fnfqYo
zQP7goMqUtUHLY0KKtTgZZ0936iHHZc6ICoRxsydXjhfXTJEvx1XIZY2cvfEuukO
0KEi9txrFUqV9gJPf0xnHJPsI6vambTUXQHr2OUjWdYpyqaNuzr0g//Fo4uqqy7S
EuqHX4kBQZOSqwKxxKWlIRqsnXxymbOVsQgVrc8jNgPeGbKLUBJg5VMoJ1uVPsLx
/WbSq/OhpLybUSDKjVrimYtqlr27lz18sjE6ZKHHJIOIFyQaB5Etxmu/ZNtv4P+n
eH2zzpberUVgO7gVSoYLOumnufdYZB3ipiHPZsZc22RZg4BZXgO1/RPiblNdslI/
4yelegRghSTZmy8WdqCLIqQLNGjVfoedrv7BjJeyxmuaLH26Ngvd2QDwBfOrEhfy
mmCGFzcTqkMU8TN2I1ChTpqrf+ZJJt4ZceWgS6GSH4tl0aYerUO35gLQkfRCLmyY
jouFOiKOO0b/4asZgZj5FSau/3V4SslnZhKD5iA0/IA7I9mHu+mtGjVXPSp4Sjkh
F7T6SBXTFVsdNGVukcol81oe6Jp7D4Pcgu26A5zAaq23alcgf6j5d4tLbV6W7bLe
H/n37MsbtMFoWYTmGLF1kvvLAzdmBl7G2IwY0R9S8E8mNn5CdmmWiyR6YV5aIUog
dUZpNy/aHBiTzBuYwCJVUrrRRg0LigdgO0MniXFBq6nM/r4eHbNRjEhcgCFnIMsg
dMueMaBbK7k1BgnBzXrd7PwAyzg6K3kS8dRCFlO3r0mOvUNP7Cjs602v+I1tztdP
bAFy2Mw5iHtsq/QWJz2h/a3CcM8ZIwYF3mQC5rUAhEcFj/ql+5ocdHMphl5uA/7e
7VbGqDMleSNw4/cFrpYaYj1t+zIqWp/ACBRFiHud3KcNEfRz1g/V2PtLB893MToR
Np/tvNNgZIcNQOHYIj801UK0rKcnbj/3DTIvi1yG6rnlGg2DEMTo0RxwEH3f+TsZ
YEqilq1FLRFQh5ZML8XvNdcoxQd65zBBY3h1BzEH9q3GKcA4Zdoen3bBg9Xe6SSZ
ZWTi/fkRuDFN5k1puaeQV+15QFjNo9UYzC5GpHcZpzaTXxu5hnIe+ZoXdoDnC++b
WEpWfiBnTDqc/Z1TC0jCNgo05VXv1NUKm0H8lIhsqmhc6Y/NUroOylDuAANGCm9D
VTjp+g7NmS1gm1Kcs6ehjOzF3/4sZUt57u0VGuIi0pKd/FFjv7vIu6KZazDbB6cA
s5XKLiwmgEn6tZSbzJj9hP25jG5QEuYYHLdroGns4nwKcIWu4f9PC7AHm0OPZxy0
xxvXo2rlxoEcq9FzRMEKiDyHfDuqhVXqRPAvl3cWRN2QinrWxUTrqEqhhfCdbmlw
x5HmgI7uosW+7gUBXulbyg4wdQKfOD9MbCduytZzXEaDzXgWojMolj8BqJeZS/fB
EaNBib+8utf6fZ4FFoW2ECAlsIHM/8QK3z3i/YqNsQ5j58JHcXEnqWOJEzWsu+f2
x0gsa6w2ydaVb8R+Lw/gzpCNMydJr6vS8VPpUtK2cjL7PuMDNc9JjrJ98itbQKBc
tu9j8gb6cWIXidmYbuS18ZqFLK3a27Rtm6reOqas07nZLG1h1piQFZFaCSe+UupS
41RGof6ne2kcOyS8+a0D38fAMOS6WbfAcrK0rWE/g8xEC+ktnA5JKxWajrG31tMx
oZV4NV4hZeBoJ1WOVmQffFep34/sI+q7wfX0PaAtAHk9TDesICqhDaAutKebEahK
uR+jF0DkdiDcZCU3b1YEYwRU02mFKLCPw8PfKUE5OqmW4fJHHNZeZo9DcQJ9iWrR
dQkrYuCxDi1+4qPetfGuPLrQ3q1J8GN4BUwNfXJPeqfDtABzIdatCutjtO5Qnac7
LPCEkWxqFgHYU4J6kRern3BSUoi/VEe7iW47/V7k7xbMfxTYOnrzqt3dZyjyt/aj
IgEz6jNbZDJDRI7RTBiLLcMHG4jU7CsK7atjLdHEUzh87RSNg9dPFoXtpU4OyNKA
lreHt6OljW3tNo/0Tl0VbpBHGxu6fCU7hq2LnZudSLkZe1h7pAaJmCLA3JXvPn1E
wX7mPrDoYcgNBNb5zEC371voBdh9cT4touag1GuzU8fh5g9ywGpqCN/ae9nevdOa
mq3YA7cRj5RLUuVtGol+oyQKOWzvJsQVydxJ/oFjE/9lx+/tpecdZZ+cnLwjj7fA
+nP7aujFn7SpSegSleZNUKj3rzi2lheKrMSmszJm5mWvzuURzS29uPuRmve8bhEV
w89/71zOKwIge1nMNZT7zlCaANnWOQR26Lns3XxSEnofd2kqfajkbZAZDtkoHFu1
D9EFvYTEYNFkaVrjlsQcf5z0u8xrSIUlrwhgeAUcHQpYpFbxUPLsG4rLfU2pmHSW
e25M2cp+XPISpohI2eFWsw9TZza971QTmbDqtEMEaTqsVWvI+cVNakyJQlK/InVV
2ZvXWq1+4Cy9fS0XxeWSciITnD4n1O2PF9uONKcge1q7xT4lexzvTdBxuzVL3EVp
R7iv9mwVqyqudMBOTCVfZSiIj72lWKZvF7UdaaoXBVR/qf7ggSRWCSbPMWxACC6z
k3tP0Vt3mEnheAv7nO/ebzXkl0tKNeHb58/ijiuugUCzyTNZoe/F6JD6TeJvC+A6
WaVBOPdGXS8qBFoPqfBJwswPxq0BObZjGO9885q1WjysTahVOO/Odt3Am9viS3ZE
C2CHDdAL/X65ZKnCio+OlIGiX9f/DUf/+49wJt/05EnPt/f9yPVTjT9L0i0aAVy4
fVu2uj5rX1ZNJv1OylUQruarcgJWCsC8mHAY4C9nIqb3XXHzg1YWNEScC6AMejlO
9ONkw5WWs8CDy26pP2OJ350ffew8RUMJNQSnDkNk+BhoZ8t28dgm6v9FmBYCeB24
GwO7eAUrBWlVkIYZWydPfPo7LBm0QPzUEXeXm408aPqfoporpPGpz55C0FkC7tW2
Mf9P1AZmekaxWmU6eiClahb2U0h00PO9ZCEk+Kr/v6xGH/mn3Esq5EA/BsxnEUDW
rMkXHEQCjhM896ovV8i2LghbY4GaNGcWDdCrUToVtNjDnyzami35TQ7CfkgZrPc/
4JKaq2+Sel6CMwK3jUIgXEtO929cgUElOf5Z2MDJbr9rOeMg9xS6heT4GW34XNxX
ZgV0G5d5WRmj9vDSP6N91jb4DiKJmQssFBDYYSFAEdrdPb6aigxVprLAJrwGK/IX
s0xywFczxZsgHU/H/sVN6oi8rj2X0CtLSTtNCXmaHQGzbLjGZNoj+d23eRu9jG52
Aze0zx1kW8dIwMDCKas5UZ/HM1LMa0c+u9Ar+MuMil+kEVqVVUI84BKRedFF6o9Y
ybQpGg4geKowB+7qIYpb0w==
`protect END_PROTECTED
