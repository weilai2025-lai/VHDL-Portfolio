`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZRQuwC5t3+KnJjevh+kthCoV9vX+h4Zm8LuOzBoF0XMOFUxfhvCwDeBdtKSSVKP
pNloQ2NEymqalyHxFIPOdS+EzPhSfgtT6I3HXYXLnYNeI39J44A0rET7YW+nanao
4ISZrLLgVep54tXYauF49ScCYUh8DOQr0b//LflN4IFG++U5UBh4qwL5/QH1H7EA
B7eTvnVURzpq1/d/9dbFDJNGOHNOfynMZaa6VV/KaOHD2jJYE2+AZpBguM22llek
ZvJakXRoaCDQgnh+AUk6U9wexX/+dVxkestvfFQz4UihV2zRjZWnkKk0GoAR7j0l
u+AYVxA1jzDI2vAjNeuVxYmVkKamfEdIcV+YYv+LAIDNUQgju3bPzrLPDBOcCq8r
wRvTpW1bUdHQ3UyH4MqlM4ktNvv5VUVFsrFEwHhgRlqP/L9p23m5wnGDWa7ESjSV
upyNt/ejw6llOtAf+2Xu90eRkDhcOFPQL4L5h2CFuFz6iTyCwIBrR25fmDkezLI4
D9hqYs4e9ZPg0IgpJsXDnonGIApD6BR8T9smSwCpgyXk1r6GM2Zq0pkGs/glDJRQ
prvWW44jtsu5E1/6agYI6/u3xtocclQYjGU9oW9Xjn3F3Yhy7yPAqutc6MOL2I+A
so7jWPa9FFxPYtncH6mUvNCqgd8Xfdtnyh0ClXEi2/59CzwC860tslpGRFgK96N0
yFhd4jVb37c7yRDtP+GJtsBBwX1ZqLnOC1elbsMCuAzwQh25Ed/r/DPm+LTPrK8c
YnEpZOFnRiv12tRVPuqcLGUHyxqEosgtyG1q3FjOfNWCDahXYi9HTjvzNf+JjbW5
ma5viys0jhqiUKwcE5FBp+RJomZmqHH4fwN8b9fme7zP/19sz/TDYL8OIQ9FrrLg
rObG9Lmg8oT+Q34R6CwCYcynFNS3XirD33cSbh6M3GSf86EauJbhl1OqK/a0/ap1
LFVRka5QyMIQ5jzSkNFOdNFvZCgYJnpO6cFOZZcD7HkHI/ZICSzstkn+U3bOAph5
ZuDGfMk2G1GD9LJE0dcvgpuel+sEBLjy5cx8FK/vTj/QWxbpqel+FkoxDuL0gkSK
nddHK41xcv7H/q03dJSAnpeyMhTxL60UIAPGPYC3RXki6hoiV+KGpu2Hfoq85R8V
38mjZoXKcQLmneXHxoGyGG/x+doSDKvmGeCiv1AlK6XThopf4MFHQFPotmljZOAF
sRuQutXpgbyZtCni4b8L/oLIx7LkQQjB45sYsKzSUS+9UCxhFlflG4pxSWZpEvr+
eVU3tAdF94mrxHvC6YsOAXx6rTXCAtZ/B1zmAHy888cO+U+aYlcxMLuYqA7MbLgp
j4IUZGhrc7QOlnUlf4D3OQpi7xmdwAMHtpFgEI7WYaDfzWdCB7kC1YV+KY/lHctl
uio7eK2CYQJM8GJOc7sGQFpGvFx3M9oWZtIhTJmTtiu5Rb+O12pMd0nXZCk3xoIJ
`protect END_PROTECTED
