`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WvG+SWQvMQ7/ADGGQ+m0917rqFexXGJVz7LvHLheOdVUDXoIDmOZ3pYTMNyA+dUX
qh6U/m9h00bKt6DfHtGyO2L4pMPyaHcKfAO5fzAee9TJxHiadw23h1EtQnvT8Oar
MgDCjh1eSDJ7c43P3GCEs4f5lNcFSssdf50SXMSh3SxF58RiFf9/ClIaA5qaxzxU
sFwrfCQQiP6g8pXERr+e6YhKhCHINggpdDPpzvq90jM/r8zzYQDGiY3HW4t/cHCL
PYNVNhuWpdT/ZJ/ORZH2Bgx8m14roB7QmZtothdLV6bgamU2TsAXiIWz818wgt8b
Md5Nrj503+mkm/aL3MlUFj+LKKWJAIUsp1dDxDWpkGW2tfOhX/q/iiiJtmSZBCfb
DQlv2uDQ9Fd3uUS0k3LV4VGKXKiP4XSsAY15zQqfDCDZv3iU8dxMtP/TNK7hXv9Y
sDoaZfcus4cIGOY78sraIXLgpQ/qI0Z8SFMcNuUSQUzhLRxPLgMOOJf5UjeBJZFZ
Qjmv1OKPhEDg/SXWcy6Sx/T3vvmay8hqKVOHxdpvOOCrk/B3DO6qHMybVK1sMzUo
owASWP0Hb87RGGLqtyfMc5+ULplwto8MXovtIDvCGz/b6+//YgB+W31V9mJP0uRl
29k2IGTR9Qgfq6TRGApRHafj9LNJeaKjcs9shQz8mo88O2FvY//WjylozPKrCyc1
/LpNORy/gPsQLdFMbOhWaIkODmY+k87pbXs9HSGyGiq3lzEREF7YS+b+qVFbSdu/
27S5JchtSz3iWoYxHQwnMMWaMX49hZmAVEAKjRGMisr29wJ2nafqPe1KfXayzcfX
cSiy2bPrDAvJQSI5fhsL6FsqQG/nftEKeprr1MQRanJ3PwkHcHRRpJ9lU9UOkkBR
yTgR9KcKRkjpOumYxeHjLVsMH1I5ThcI6SB8g0e7LeVA9dEva8U7870JmYc2QVGO
cU1a5lPkYvX2+r99cdiroVxaMZbFdC1GFQxfGI09JRnsr966ubkfT3Nuzs8LIEjW
ENSlSB9zKuYThCkGsVdoHx1L1dEHnp1w9Y+b30LHkhU8Ov41SrCgyPu6WK2QjyJ2
sgq3OWsmv9Hj54R8jG9P/LiAl0qPTVaWIP3c8lgbQRtofJtzVebtIqsuQbaUAmD2
yVWGiYwQCo9mZ9Af8KPN2ehh2Ml46ohHILejFPf7leDlgGBiG9434J5KeT9MygRS
UTibfRQw50zHFKdKFFDGelVtd3qOT7Wt8haKvFK/PCRFmoxF8T4Rym4+eGQJGcT8
DIaKFcXfnuAYfTyG8J7FWmTEO43xxDj1lwsvHAiFBuH2Nl+2SW76x1hcCGYbVUW9
yT9V8+OK9LJfC0y6ibp11K+WRgrGLc0TVoV6gfGZR3B4OwNWclngyxtHdEIbhv9r
SnlVa8046hN9hZiGDybl8fL7JtzlpnhSNzAbWyu5YEFUZkOQNAxyyjRZU9vRH/FP
7lTFa/fqLv51Y8YYU1YFuu5+fCkcgzDdWjDkMl73l3+V2WgxWJVtTaX1dIRzxzXq
kzrIW/IONWm2YIpzKQ+wyfTUUxGYBswxuyCHy3ebdAG5JD5xFD0GcK8Q5ZnBDbEP
tmrSfVVFc+G+j6Gop4TzoPvkR7zzwpGvUCLWd3nJY3yCWcj1suJ/cWqX04viDLGC
Qtz8JBzVu7OleFw79vNvR+pngNi//JNgDfDjMQCms7etJtRcvOpGnQkjCWvL9zBd
Ut2yU10UFbGbe8FdB69tc3dz3i7Z3ksxwCB/HW5plCzR99YDe1AGNEdtNEruuBRm
bH7rRldArR9tSgY45LT4fm6RZR3NIJg9ZQ1DnpmERSkKJVKNqmBDRq4aQ68lvgxC
GkH+J/9GRzjfrZpY3wdVssda9rQYCHgApeHvVeRfcrcHfyZwRv2X0teq8RwyE804
YM9fofBT7Hm+Iu6u9ZCoVRCH+87a4/nH6i4MnF//ZCRSbBRAPlM1ZxvpjPq5H18n
cpPhSvGRu5nRZtxvgPD9MRtrFHsbGDfRxRvRB0UqUg3X5dkRrHgHKkr6agmghL2p
CIaPn6kPInANLdV5W4kK7S/r+z/7cg0/2lE1hfRjYFWPJwvozscbSD9YSBprojGo
cWGbquQifK3fQWEhlIVoQLq+ZaalXXHmIHDtJlGPD67nqeIkN8opynJnuNm9VzaX
Gp6z2ON+hO6vENiDk82PXFnAwEB2CkAtT36BZLg8B/FUGgbP9N1+umuQGcgy2BUG
IgK9eI8WEDhy94bzk17Ru84n7qIubMsUphC6FBUZffWNI/XY3HIGtvTOy2crb128
kTZE5IITkNZ0EmhgQo5cOhzcgzmn9lb68ZB19j9OgFb3hiNoAR/lRq6FFs3zxf8F
70oY6kDKvoAQF1pjJ4t8lXk5ai+9+DznPxxwHs5HaB/CJqrd8G5xtgZKmHugSVfU
5/tWzk8+vrAvQ513VD6oklSiYBaUJtUVSsr5uImR+7KaghRUNwDTOX26qtA/Ib8T
pGfHtviWEIqQ8FWMtCMWad6VLwKwuSlcOZOViNXXOrUwqOIE+Tg29bGKMes/cSLA
uWocnGGT0W+9q/HHR0eO+vST9L/0ViZlqe+LxAk0RONV84Q3NONrtyBBH3QtCvBr
ZXpL2iDZudshf7vUEuPkO96g7YEgexdl+OwuG00VyPM4fj6pdi8DNlakD9uqL1VA
EYYK3toC8FtwSGSsWxslhefMuS6fSon77EvOEy9vH+j4wRBXzxj6ulEm/qxWIHJb
YhRB0xO/3L3JDTU5dVwncZ6kHMZDXwreqmQapZG+kScbVCgxKgQPNmuduGJjlexn
Fix+9qF+cRhuDfCur3NdGCGqp8ZDzoct7/Y67iIXSdxq4omlNC3zg/BcYIY1J+wL
yh5pQpJ3nERcFMRqHE1kqyPN5Bp7rUGdly2CHKuJCnYYocav4hB+Go/PLgG+YNRn
EdiPpUwWy9Co0FaAbC8nQ0JRlOnfKL8A9Y1XfIbh2M1Pexml/oPMvEoDSBrEMSqE
qRc59rV4owLcT86zNKhVqL0yo3kDm2m6nEtumHhvLnarczQYm0PVfWjfoFkBtBCq
30QPfQRMZYfvuSLsNZvXr7B9Ov3lc2gSJJyE2EWGZxNAHOlNYqSvBv2Cp/5HGwXX
b8HuNJTJYYb4TtwaMvfGHMnC/hnAxxaFVJ8eXp8PxUI9TSHZEpSO1DuOU90O6XUv
HkOh9fJ2mKeDSrx7fNBGlLfBnZvxqfMyFsbmH2Kq2lJXz0v5JWm1LQ96yP6GgOuG
99wn/t/2VudURhwVOSyv51uRRCWHxcIL48gh2mySVrQDWPeZ07hMU3JOBB+/LCnW
3gQJ+q+Of5ouaLzj4UAl+Fsyj+TGuG6MsYxIzb2WleTUNiX7qSZ29R4yBbZBKv9g
v3YPEm89DadOfsNH5vYPHvC8SSar5jJL0WfIzwS0uQG3XPRcHBYO16gJ8D3jzzjE
yu6TS8ieJoeTLc/8Z1+2ODyEBjwSpEW45BVAikRYqXS0wg+u/ukwaapbzNY4ROiP
iz6zqo/ot1dCtEbci5nsZ9L3BQjVbwKNnlHToJZwqFcRA9n05vMMSChk/2f66mHm
JIzA1AkmcwJ3/Qe+wRWJE7Jwj2Y8J3KcfkzvCCAyzkxNpfc5tYUF3ficm7Teq0jN
Ta17h0i+aPyodhY8loO4oYb76WxQuIvdQTkJXWUcaqz8p+16T9PKg/58p+W5ALLz
sqCYkrAUaYICqB45cKJKGiY1KRDCvdBsp7Z83xOali8/jJpLRWpHd6v6VhHmOUyQ
XnZ7/XxS7TYxjxvLbAEw9VZLqT858+lIgYyrVRdMHX1kKdanr2ajrO4T59t5tQj+
4UJxHOlxC0QXOz1aKCbXX5a1AIEpKhQN0G0FWeiS6SPy6bJJ6OJev7vIyZJgPVpd
BLlQtXFo91W4elFYoohdlCt6uVrek11sg90zjhgY0Mw6pgiiJ6yUCfpRxJ55qOS8
etHe14JdnX8JblLVshDELGpDAuGkcR2h/M8UdedJWzNnPrKuZf21mFtyGl3IzjeK
6JUQZgqd4a7bkmz0ESMwYe72+vHmhzTd6A3sJv2gBUEghFAbSdleQGoVhh1yZq3A
xnKoO8VNoFhyAi2Fwfdmnjm5dT5OyqMMRaRbiqpxqzXN7gMBeRes2R99xND+3ZD8
u2r/Ks2tGZJ2rM8ec/279QgRL9+nmMnhsBOjFRO+RlUCDabVAU9DKNdwVH7RdCAL
VRYeTOR/u0GamlN4RUYEs0WevzJO4oaS3RvgOA5WM+KF/YLercCfafnQ+gek3Gpq
Z0EoQ6dVK3tANIfB8shGZ0xjioPeQKA0H1NXhZkpr1X3YI6tXZF88EN0d6nDVDN+
C1FplBocD0Z8dNkT/yd7mc1lgobo9/iEz+UDqE42yYhpLWMKKgipDQB7dVSOPjxF
r4WPNN//dw83vEl4bnjV9Ck2z2SNcTInPnC0OlRp3qqXehm3UQBByNvcjuKrS023
9LPDrxhEAIQKbOx79UwiWaH+tYu4vdOEo6b/E/c21aCmMSDENwmVzF/cYcUUTH2H
121pOyytiVAOdPw0MlaTTmwLhtntw8NdAyY9uOdO39Dt9ndCjMz0YyTmvayS+vBy
+RP1KDjoyx1BRWiwMlizM0GXZ8WHZIxX8dOZEemAeOolvCvpM+RD8R5ZpQsf13r8
4ESD0gjF0ROvgueTTPOmalwWQUdrxu7Ad5DOZINgMujIetOTnQI4+3H2XqtC3jdH
gEHKICVwR9kIxjrLxVNTn7Zr6h8KQ1D+zuJqG1L9eQ43fkemYHImuaJvrj9yweRs
XO8Lwna/DsJZE6IyCSa9JgoozITbKRY34zijwSJGING11LxejYICHg9azZhm6jDW
6va/HdcX/0ghvfLk6gXwRmJGp/hC5+MNYoL68bZuWk1Z8ubmy5NH9iNHbfxzkLQ1
0hJoQ3sMF8gce7XL1hVr5isZOVWSjrxujlSj5u05N5PgldeBPGsd3w/FiyaDNUe+
4XKzDmlWpHPVH2HtSyzifs37kcEX5K0zC9MYH9C6RGarRkmdKzhYSogGmFoPrGpj
DEmj0fvtFtWYr3IxqHdDyT9nKjHVSU/yM9GILsFGY4mlzlSIhm6iAnwQcGtu8EBs
bDTCS3VDEJZgmF+mHlXXX+UrZZ9iWhA4Rc7Ar0qGOaXr2C9ucbyexygUqx5XYJUT
R++2YL0qRHCFjdo2u2EfDn2YHfubaNfYZ/XT/mBHFl7INyRRilymYJgJ2Cvq9FNt
V6LYMJ5yYeTgqcEedJVCWN4RNwF+GaFWRIPMl8YZ0iNHjtDQjI5C6/oMc+0IDofP
9k21iUm28r1vgwcbsdk89fQqN+nSyTiz96vaGk6MhBaVh5fdSAAGiv6pVwiBn2tS
iUVOD9coQMsP00114Bz7ZXPqDXMrHtXWXbwjWPgtmaB4XA/vkuqDtx7ZSSPS5Dxf
O8N90eQBOYT147mL7Y7ai4ZkHDip7A03gKIgg66nLZ+NF2G954vzlcew5XFm4G0k
hnzhs+bEYQrWlKns7DPyFYQ9UpQJZ53mosgJO7fKknx5EwHl3olclOB8gZw31pgh
/og9uW+Zz7YdNohQsF4OwbCISjR+EjbxBhYY28q61xw5RN31F8ZhdwEDwdqSbjLg
6uixhDW7bS4GWrPgbFdcEAwn7EVjpR9tMFOfK/hC73k9qw9k72zQuKzRBxTM5JRw
2utHLoDy5AOTl139DRT3W2D4zwn3+N2leuk4/7BWT5XYu0MBLCzYRCTsChI+eBdR
HqY3VdeqUo7LXP0RKb7kzZsFtKE89gD4MMfA44NED8j1A9zTuKLE3ljHg+pOf055
Ece6OMG18OmdHdQ+fIvYMPYtPcrht156hGax1zY3+INqz5fishEaO+8fAQF4sFOS
y6nYQVD0i/uWUqdgAggtMKHdfkXTxnUe+NlcdfR6VgXkN/PZdt23AiLLv1n+NVDy
B4e+/GQQU2MVUuZl92/PZ1yJBBHMHmY7NWund2cXoU1TS73laGdkeVdQ7PaAzBC/
bJx8YuxTbMhikOJkV/Alk7ySKwTaL9SO0mXubPclWxrjky5RcMw9eQuQ/hQyxuuH
f2KSkx8eSLs7ncG9x9xj6HHumS7FlzldnIwSI8jbCxy3O/F9SukBn94IGvgWXvm8
Gcg7yzaot1Fv+R/5cYHPnWncngit5ShrdS46ynP6Ya/E6jChEWeTpkpcBWmHUMQd
pzbmSSxVZO2tth3G95ZdXkL07RBchQXviV3fCNDzVvI6AMERfivrtubJVTlbs0bW
3roP/NTaK4RSfRfbOIjl9DI07qIXklyq1dCDamYSmv+RVx0Zsj40OlDn/+es6QtO
smwA/5uTxacuPig1AeISzuDK9Lt1BDsfRdbYy0Y+NmZWYLG9BekvOnxfTf1moLlC
/VDGo0yxjZjhXbv/R/EDOtplSYHnYiWFxZAcc77X3GS4WNnWMxwbttDEJFwVAhpB
vCIkX/E4UYZ3uYcEw6ChIgngWBOudWi1bSYdNYXkkWVx7PZ++4qpikpLMf7TFQGn
XdcGfBRekcxASSh+ahgXGMj2oKj/yBDSA7ZUGBnMO8Yl5dTm4Kne9fUyF+eORlAo
W5TWP/btjY3Q7xnbbtgCqTSwccuQ3NdEGglMaCKJ3v/ngoAggLvA3DEcONJ8psAx
9xR8FQhuZwO3a5G2MVhnWFUXNLMmjt47nYDcgwoLhdkilR9ehcqgfySP7w1FKf2b
LHqanZq/UC0tNLwFEcEnlSO/kTyoSImRwvjxxWrNqARpXw2NeaJaPsK5AxbcB/3K
yV/7Jw/AkHVd6rnTu83Mn5C92yjhvm96RESUM6T2SPXkpRNMwplE7WwLCjBxKtu2
QiYHijpfxeV6dZhl9rHBRc2zd9IPIp/30tCSFXxeqQHKmQhoCpy82bCqQY4Jx6Mk
XnCtr2Zl88hya1IPOT2l1UQmE9cTk0Vpi2DPRzEua5aAKQ2PvUJ/ZktKrkqKMS+r
tPp7GsrxrDeYE0k8Sc6bRDmyJmBX0MGjQhmDozJKX/td+9CSY5Dny2aH4bYs2IOE
/kAioKQn5WP324ExMFq/FGjr4u2xzCR2BbYgdOr5RT72IVOFSscH3Mv+4RMXi3oW
I8lkBPRR9UroGrqqBfOmmQON3m945vvd82gMCid/xw9uy4r9VLVAXyt9ViqNFma+
GPjrI/LgIxe2myrgiZ/rErhjgZAkGcnHY3aVrYGKEnaZ9mR6DgOUXK/jS10tR7sw
WvheGsvvQD9WAl0A013io6IxzG7gIW01cp2M7vvak1AcA01glZKg5Tm4CI5joe0B
onHnP/4PBJZiUy1UcD4gtRDi2D/gm0M6sCkPfY59kOqFDejmN2VjoO9GfnjYvL1v
k/ACl6AylKo4+uUR2cZGdN5Jesff+uG18AW8zOihoAOVtm7POAo40fAHLiAGnCOa
rLLz86cYuQCcB0flhGJ9b1MFDqR85QUwmZVUJLYZ5jZ4n9iUtKM/ogalWdky+sci
/WTxozz+AdvkmLFkoyR6X9TLgSc0GSYXNpfFjK5RR1xUFRO+4coDzCqGTK3tG7op
DcU9O+InZGc6BVNPlrqX6XodyPeHgKu8anUqx7R8bh7NPW91TUxUg1bgNmNi3gQC
6gDf0cYUwg0oK9jNZR7la7DNRH4NjNelWuQYvKLL4utAqZW3MaKvSup27Z6rjMFO
TmWYb01ZrDr6wM8DBiF4LUDma/QI/K6hAMeD7eAXMb9v6PsRK3J2Arrxktb0KuoP
6M5L9tvnCufEHMeKge+0tHevPLOUz1IvfX5tt7AmvGoGKrkSNTauzN2BNQ++uUQZ
oXF82yc2Mk6cnqBdbtswSbEi959f+L+Co/Ef+VctC/QMDGjna4WbIoCqli70jdn9
NA3adoOjywnnIW/GvuuQQZKFaBaGOVB5WAYdYikfelnFThkbLpOH5YCid8Tb6zcK
oy7f7tm9ztBPpEsP3sK/ur3uev7DJvseTf/fHyTupsOeQbJon0qRjvt5zZCFKyuX
/QIsWX5ubiDeIekXlFcVPFLEP3qvmnUur6AnV2OHkdz6R3EQB4Tsj3tLSKkaWqhU
X1CLm3c8dhEO6GJ10nwwbC2uKzcypF6dZAC8tcF+mBXcdeMTFnjZ37qyoXNq6nJj
oEe25Zv3Zvvm/fSkL7FWH6CuvoeVAfaWzH7OdpVoo8lt05gP5HDO48/048oBJEXP
My6BNGSA3hSDQF+hbNhIaCnxz1+Cm+DWyeAzEEYfBpdNl+at9XxWfFt6HkUl66Ay
Dhpfwfa7Xt7C1IwpXrg9VwTwTu+ZBW8Eop2p9CdiCUwZ+pDNP/cJT81MsYVrH16S
zRBrKq4zzstthiOSXtZdBTmXiZWqnB8mBTaXXK5V0Iiy5gg6Yjmwpg+J4NkkzDIN
MttAb9x8+pqv/ztBComg/ucqc4zWssPFtX5o/cCzlO75rJtPKQqMDIJwOugSLf41
oTK0iRQ+CQQoFxhW7d2gp/PAyLK2mBtIe485yLys28zRHtIV7cz1kmy2A64UcFex
jGouTrLpGLjbcU5jS/3S/1CSGYEmcyyANP8GbcryZRhdiaDs5eRRtpf/NN4hCiKd
T0bzKwerVpUcIBCbfy6PMhMEnw4ydDQemM5ZXMOXElqWR+wyz6DIupx0+hTNi5tf
uh5iphoQfApbPDt+NsUA6YR4bLUGWcfJjTD9ZyqPw1vNvBKRWPCUyGecMO5aIchW
5kl9UFWtvJizmAPWA91NmLOfC1dnPiRPMkS/95uQtHE5XY2cZQCTqVRgVY1eHb9b
p2X9n6oeNbUFSmpxQTxq/NKiu0ZChgj4JvdFN12qxQg96/ngPNDRSuJIxYJ9w8lU
gP38n8ef7b0oQycP4awl5Yg+R60rJtjr6yvRxkH9vo6jmQ76Oiff/QX6mSKXjQQA
gahWEHv9mSMNANAsugMCXlTmXgGhzzyLneB8ER+NoMkjFqUNU46o5WQe6RV7FSS6
vFeJNCnWfOu+rRlmB117D5fdg2zfAvTswomXwKFpBRPEwg3HxCiT08EVuwUiPHJF
OZfO81pV9UIYnjytYj2a7lmU7twTNWsfkSBdt3Ev7kMrBcdH0Dk5VoQEIqULNmUd
pYdS03hVIRyd+GjvRSUNkE+UOp5rPq6WeFaxqy9Th4f9pNN3UgdLzUKfk7irNubE
y3GSmdJSRiZoqQxKSbroIfXR9skGH41qhPs7JEdCCm5a3NV8WEoB9KNqAt+Cu+Wl
QxY7BVG4tFTzHPNBpV2W9rEF37pUkxkTlnkbrerSCHxNO9IIS4nI6+CY6heYJ0nJ
nJWsQ8glp4KgwDsBPU0qo9OFvaXFmCo2rpLYcOv7EO/Rkk8Z45/LKfzIcLJZZNFL
8NVGMx/ET5fBtESxszmCzOSXVnkCrDq6PbUC0Bm+EDJWhqhJS2ROTNKcSiPoUeSM
a4/QloJ/w1g7OXaiaioEtLGa3oQzY4Dl/XMFJj+1/W7rYovKI4/MSizicgxOI0pr
oSd7bGyD/9EksNSbuKvLAUhC5BR2YewAxF8zH7JLav8i1YZTev10ANYaXESxszw3
+iSeivcqdbeo8AoEnWZBrtku18uX0gmcXqmUGoqWXn0+eHAufpVGScq3qEbi+RV8
mha+VcD8mJeV/BAMS1Ev6iLvAekYRnSrHaMt/+Brv+uNeTXjq2QgvtxNSIbei1no
RKhrowpzf9aF5HKE+TM0t2jiAmn6u5l47FyfuAUCcFOgEDgZ3yug6TR5yohbvm37
d9FwQknK+u8kaM0eB7SuwSWABUEmZC+6oXk77p/n1GLfzefebBPySNI+Q2a1Pwo3
hqc6P+qG58rnCZxJ/cRhyloe/84kxQ5inzobCz5QYmz6y2EYkQJsXOy4sUoQbmd+
aAb5S+HVq0dFSWr7EMjN+eXph/XJAxrTaug/VB44E8oS8rxL6HWOb84ny1acofyl
YUbXlmgOyfz6gIUDwyLYpVEx/IvauAbPq0EMa27kQaIldXptvR72TNvmHy+hv4+/
hshYiM1Ihdf9VIPozVekdUSY32PE0Ts3OqoOBbk1SePhBTQpYby+xI2oHPb3wUib
liAkBVcYA6aPXNwZkSUPsVe/qQ4iMX3UgFpcUvfk1C9kTVVN7ZIwMooUy/uPYxR+
Mz3MSlU1n/HNaG2SgFrT+NP+3ojioAzL8PFtqt8mSBFNNeOexRvybGSqc5UbqVhc
ARrTXjA0YDa6CvLutG10lc6sxS5r5F0bGnQ4+B/NFHfJkVYCqEoUPx3F9gmz0K1P
l1LIsdyRKKY6pM/jLR+AvofFc1Z+9tu0zTun/XlxRhKC3Z6YVbuBl8sWF4clLgZo
Up9I7ezwXdbdACA885lyh2VYotpKPI9lC7lQC6EHNsgSVIUo3tMe86v3hh2lTb9f
2eHfIbbvgsw1vqjG8fUisnudrtPrKd/CyheA0JSbg8yMSersEVaoHAXyDit1TidQ
dPxoTPAMzBJSqYfSEeYTRS5u2AUk3pXV4h/BpiZIjHITa3s/m6v/afBeChS4PtZP
V4EtscJZQDqnnZKuu2fqvrfSRxyVOPPRKEgorHUl84KTb3MhiQ3y62vcuOTrkVBA
XEPMmrN1Gp9WV7pvD8h5/3YK5Iw2MTytZTDLQln0Tzu0i3vRpbez/MtCn7Q0999a
16a7uxk4vjcZDkXwb/9nKvg0wn+Ou5Z3Yl+/0msT4kfqO7+vUYXgNiroTe2vqBzy
mGl0MI4fXpvTyZH9o8Zcf3Lp4bkWOdnc2vnsRLvpk2d1S9ztsH26z2HaKAwsvOh2
IRxiupu39HNGAh+tp2pb0GUaK4SrXdTV/cSu3swOki2Oh2ZMWXrUHZ0S26m3PVDn
NAu21qMYd+35y131QXrkP4pNIlroFQq8R6rYSDzmeXKnXzKlVSt5cwdDRuciRbuc
gxjpZCmIIUwYhkXOlUVTnhCPWk52ufyR5sgnAbBQYk73OvR97imtRaYJOMI5hFdB
H11DCQmWpMKf4Up/296D/xf0wh506mOjN5OuRuGfi1qY3LCyUKre00nhum95EacM
lv3CDh6Kb4oSjEVZADIQxUsrrn7+HMhubKyiMGXNbxeqJWbutF/MQU6u9iAcVRBd
Rvz4ohigrKJlQ6FWhPQ35q/03HJgZdRYPzaEShcBreKA36sIHKyfXwbGaLjwOh8W
3bxCsADBy9EyjmZixumf8Z0ik32pdUx39pZWrgyWxFAmRr3JAKdAaEX/s0WbzWM8
gcTS0YumRTAVONz4c6jxGtzQcM6GAH4QUWOyhqy65AIuSvciPBm9uBt/1eM5GFJ/
UnxsEAoiENArZVhhPOypFm1WcN9mFQLrGfwMDzRsZpM/rmz3DMdyYkfrgYE+C2zw
f/6e/ChiQ8iWiuecVsDyvRlbOhdPi2l+jjKugR+fIauYU2TzRt245WEN1iVSZQhb
eHoezUZqMGSl5iVqTInvitcMQw3m934qpbFF1fcDz+mnAWe/rn88uyrUbUHex4ld
qib+w/NRGRzE3slAvY8uxXYia+NgSkI5BfV5xlCepUaPLteXipHH29xqTam3vCOk
ajqKVhMrMdsLQt7C2ZWv2kiXtoGVoXldJ8xIZdkBpssUCZBm0l2x1LoqUAk3SM/p
PrH7Mw9Pj8/RBse5XZ7qfZ6lO6lkxATlQv5jGRutN8W0tPASXOR6eoPBQS9tWJlE
PuRxtdGbZ+ycjs5qfXGgfA3uMkUOVyigI4PVTMZUgel91rmOu+8dEc/JvCVwQxwn
rONCv2FhGRIwES89EbN/qPx12LMSKAXPUx4M84zIYKHR803yW/COYQ+ZKeFzBPln
5GhwT4vOBi7LFEdMD8qwGE1jqzi8T/npSeeyxdL5EacU9dEwPMRrs6+HNL3Zse7G
seUTKcKfpEk8Wl0zXXmQY8yWnuCJ5usLjdPKapQr6w5NrkIXPlQPuezHgicP4w8e
l4N6891WtG1jr4v73R+y/dKNHkrdcC3BubKG6HXTCJwwgiDFnE+xkaFXzQDD76FU
OotFhu1WJ0GN1EEiMubT2etIyBmMJ7MGQdnjVmYqzs1SwLo0bGQPfVNvAeaFlet8
8P8jMcHpSJ/xW0jV4Fs4xuu0G8SylljD7RpLv+FPcTo7yg+ECPSLBNm3/Q7ePUfi
nlUQovB0vI6Cap0h9EQw0Q2IvHJTov0SzpAdqnjOsSDy62RMV+BE5+j0eGHxYr0S
0EudCy6TyOYGPa8ohkpFZlUsY/AOkEUhNIYmknr62WXSUh+p9gbgfes101Oilj/R
UQBv2U4BCYjWi3KMGdQ0QjMfVR7Eu/vFZCt/pab0T3mp6jPIpd0LDWBBYh8gxDvb
Qy1/4lJ3HFLsNBncd+pVJszJYoo/PzcufCgnNiOcSc/wjhyeE0OzEPouzvBnt60O
vTDpTRqIEAe9KO9N0KnV3/UWFt2bL4Kf6OCz5Vc2C0Yyf8DyYuHWf2acwbgtDcpE
x8tAYTLFV4rMXRsWv7goAhFKhaQtWg11doYa77KuJKmt/1uJYT1VyCRz5vFDI0R8
dEB8JTIq28uKNWhsSMSvdiHcaKAAdvvvJGd2iNaAlZspJ2uXxb0Sz3XY43XRLwM+
Qvl6dAVg/b8HkTLx6aNd/wBMrzhfhE+eRkGwS5mCo01jvxwV69AXVvh1O0KuS5ON
Wtz772iuZAmuKjqhWeYzoFaOStFImeNujQ+IUj2sGzMQIhTZdb0VZpWrVEMWzV9S
ikGceGnW/YfseVyGodF+vj4ttUjUGavsL/mcRJPgWwoPnZesU0xhPNdWHFbIZq6W
9sXm/cU9vpCjbJ99nensQubXNhxdAYEw57FsMBjDLSCZzyU9ss1cLtF1ilACqQm3
n/LSvBgKNEM7wU20cxPLEBj+pMkYCSJD7o7aH/H1vmxZIkfNx+gGeOBiBHmPcaYn
5I/8KLvrV+iuTj2IKw0KoL29KJoZyopRSErn9vVm6MlZyVrL0sx/NMsaEtbJsHX3
7o79DhT9X3iJj5s17ZTeQJYt+/YiftziQPp5SLa0fqa2qNU5wQp2yLZoFEzqwg7h
AEJosQz/oxT/BRM6mDQlt7rAOupKttz6XSbhX21l6XLNTxm5IbEmgOkeFrckd9Z5
w6LP6qZNu1brtYOqATtwDL/FFDxauAOmAv0Qyzc7AEtNpaa8JJhiiwJ1RipbHkPB
e70QR5CvYe6wpQr2FvYb4p+CvH+4zwbjSf+/1EgsODe1HWVpTQ0JD608qYmGbirT
aSCWKbJrpgxEPg2/GNRs5T1RvlLTVoV90kH9jczMfMqXNk1HoGb+hrV4YF21tqFw
B9tW+2heHMgSZSCiN1a4UUQDR4m27yjaky3dqF94yw1fHCR4lhHo3a3iXPcAAZJ3
2l4mlmowncKlUu2oO/tc0EVHOku5b3TRVbfWwiZD/sZ9rR7iogFrgyv87TSuRra/
XKePfsuv38hCoRjl/4PQE7bWRzaRoWFBIcB5v2jJOAWvi7XX3JjV8L9AlTZIc8QY
n3V+iQfvhz/PE0FJ4Im22nLn2eWiZt5mIrHEvJg2kekGxdl+xy3fOIFEGEqE2l7Q
xutrg3Ev0FqAn9r9nXLnmKXeS2NDab6igV4MZ+jznn2jIajygBdqxu3opt2R+y5H
U4DvKAyhYqiQAYJCFYLXJdzSmoxwf05mWn+LfF+Cnv3qoUGgrvqhwcLS1RfBxHwd
+rIBVJvZc1bp+C8JarFO2gbo/G997sGzEojepdtdmM4f0OYf76DaZQcBsdPhGKkm
LbM2MSDlFKlOoT+ALFTlwT2kn7wKZ9kuGsINt9FEyHncKLLXOi+i5MnXczz0pLYv
ThGCYwkAHLuh+wPXfMKrLuo6tXO99yOwLayJ7SaQ86VaFJkqBoFeNbI/aJd7OXt4
waLhcvh8qB4mKzOtRtiDBszCwVcWEvUE/49QN5qxpXAOGeNeRECe/W7j65U6jLCq
NLMWaYNFwicHdCWDNUlGVVIw/0GU28f8NvsK8LlxjhiejzTfqdzCtvWC7twao6DS
a5eAB56f7/rCiNlwJxbgQhF9YV+GybYaPZY4Ygsl/gKdkj/DXjAAOpJfx7hxnZhA
7S0S1xBJM9ixuhC673P9yoZtpEAqpzxjx5LWsDyL5mpUz16Hv5Qo2Eq43ICN08pj
fErbV41YACgsyRqb/K9zaVd68QXUzeEpRxdtZqOlKhUxs6It6VrozC1GoD/9aL3t
slT4iWpp/9wd3IS9WQ7ZGvmaRuMWNldqKZ53K+3tXTVKpl2hk6CUnxehYYGKdI47
fCxOLmF3VqRv60RsBbtl/8trMk2qz9r8CV6di+kgMboH2zoYd9iC9nxTpDtdxDcC
VyoPzLuVkqG3lu+hpdo2p8qQjj0qz4qO4wr1zIQ/GEbTbvMNULfV97t34QF2+QfD
5iPoJgqUwMBs5Ixgu51tckRMtk2ykqVImFAvbDJXYiMQ2TsksbPbeerWfES1VUOY
tr2bdoZU7KNeiscywjKSbYNNRFyBVQtnm4ciuf0BTEGS+d8RWtZxfeg0tGQw7clV
yC1cuVmNcTIC1iCwYH3mqlbIfK3vAUqqYg1w9I+PSOqkle6/mfb2qGaeWLOsqSNZ
8ouGFec9E0H9Cs1nPK/+Bc8J7bsdaiuu1OEKuSdQ5Vyx3abje2fBY9kiX+TmBtLR
+vBDQf0wilYJBvqeRxlB0XXSZ7f7rBGkXQ3MAfTrcDyKpAquyKvodiwCFxtWWMOD
umtC0J2Xe/ik34RTtP2c2tyV1ebXUyFfvb1uHMhyNCqHhE2L1FrzRr79BZ+7tX6C
ROnHvoyjvIP8iQPMrt4ArbTHwlkipo+jG4Ge8OBqjjlkOb+mjzZnYWa7ah7+QRKP
IV/jIq0ntbNFvUMvruqKd/abWGDBTvM4TGI9QxnCcEUrmO/OgqJqaMOJka/bv6kb
kReMn6ED6ivEnwKssfyjKwcNe7QC9sgwBD6dEfRrx2FFh8kKqBHB0Yic2xPgqw6m
TrkZLLHsSfiSittFnD23Plix8+4IvUFhDi6bli0XZ8v9rCeyGCX4Pyl4yRJBXPQl
pKD8IREaAcrmlvH4psRludx0YCv2yuv4OOumPlFCQOPnrmqqv/295iIyhqaRe1Za
jY+1kxGeBenWE8gNrMb/kY5xyTr//6jGuJpyc6VzpufiS35WNnPBwCSQAo8MciyO
q19GzPo2asGBJ8It4t9jBj4xkG0Tcv3dq/ddJN4okMJqBc4rtZGaMdTqKtZ8YT+V
CF8dAogOZHTbvRUp+5ZQri81tl5bi5uvPlgip9owK/iECTr8G1sRB9VRPElrP4DU
4/jSFpXPvbRXQoA0iwXqSFkBOsi5+HWBWcJTulnmMQkZPSZZ96dTS6VJAEbnv7bJ
ODsk6Iec6M3BY1vZoOI4vCWj3FuaaBoepQZ1PBp3xKMxL2GQlseUNiX9vOaDg/YF
KQ+UWWHhkfMyYRWipiADd+yYQFYxS0ReoJShxBCeFzL8ZcdI31aJ5VFt3mdxKzDU
8IRtWvhAePvEeiPbZ34jywLHM4wf7cRI+d/B3IcUREqDEzZ7nrbMh/ML+1yc4U+H
1vwQHEvYbHgx6BPgioT7kCrzc+UqXklNeNrLa1ntVhYT3TPfimw+/s1qOv5HpeTY
0nM9VqeZfb/bXAr4rtVarb5Bv59qJLdSkDbeYMMLYFvIEXAwXY61YOmqUX1BiAxG
rxbnq3rreSyWsavfo2vw6b71/UFecrWx3/X9gBE3b9dzYxtU23xkKp6hLifCKx+x
cQ0Dj6tlkfPAbdV+OapyJuqlcrQydW/gvpY/F6KQ1ExoVQjwuRXur75sJ8j59R13
IZM2B8sEx0aZ/vvxiGyOh5H1bvafGyc5v07iG81jieou49qdDVKh+FGSIYvb3Tf7
pU8wC0mkD5LJAj/n1iT2H/hUdxMX8KAiX9kJ85yA1jsEaCEmD8l0lQs5Ig37/GcN
pHWu8Ev7ytT9vD+NhtRUAlhjwJJc1DToQdacRYEoZG493QKeJmRPqRGzvtQaV9mj
/cWy2rqLJnfQVtg6Ir9m0AW5MyI/JCUKvBEitT3v/g1k0IEjINM3wnnLHFaN2rxJ
NahVx0S5k5kFSz8OpFTcOiR52mYrpNsLAF0+NxEeU8yFANBxrQ/I7wMaDlO/1qZT
8yiJDIXjxlE2scChJBSOuUFZ5eiK0cDzMIJnsffxGRA5WE13BP8GYIsaGfGQHezQ
pjijeSTf0qEijLvYIuj2npnMtAIfkcrtv0i1Iz+rBIVpRC+ckgh5O7V5ifbSie6s
zec1b+6X3XaRFpTk7eWXUSrvzFMwVnJ+1ypHbOu2EMR12iKFp1sMPL+Z51pNyULC
p1NUKujjQdhq82DGGjwPemL0t8ezMYY7TAwJ6vVye4juHtfnLigENUhUwnngoU9N
baA3NBMzItpoRrzl2RglEnM5HI7GgyYCC/hpy7DxZ/cWJMueSBgT0dXpCh7Zyy1k
tZ0qHsw1JzvlrDdshMgec/o/ITgQCar6yNIoLxjSw7f58bvZOkENgu6VOqgPni/6
voYbZ7ncH0t6zWoWenufF2iAV6T+zzC56qubzQngrrTLfZNzRIPVLjr1xvwMMj1u
Z+8sJpoKMTDcl7vtPZDkzuwkBhj1FYooae8btODEPKyc576z4z67aPOpr4SIW8Ir
Yn3UPqYwl/Te3g18uKYigZCe/ktC22AqpxiUY7JBOtMVlREjI+WPOUzO9rQtsrH5
XfZY2pIqRqYi9sDIdEDaRM5cqYeYDJiQgW+B1ViJqauhC15NvSoeA+iN1CZuorTL
GoMsEyeRSltNfVkEaQoDDQJoBujP8tA1GgSrLMXKjjpRc54uoHw6qtb+oaqTBxqy
41hotYUKkobQjf4HMlLyD2Z7DiGG23ifWGk0s5062h2HM503GuZTrmuuaqqWvGQe
etB3/yJS1qDytlc2vtIDjVYYycEc5SPgJkzykCVm5KL+fxoOm1lYVuMBlbQFX5Al
kQpmSFRwWcjysYn2U4aqBUSPDfJEciAEraaoYF6/k88CEp/I7NjBcItra7yvSDeG
RQ/sKkvAs0ZAFwO2u3PDZcRJcZvriSUaUiQq8hkjBBC1AdEefl6bmaKjoxsIjQUk
1ySB4xeTHDVspK3N557e/A1cPDx0RrVeF4crxoSWrf3tigTW2rid1LWcHAQarAOr
Bro17r4hTUFYeo72qe/j8X1mSSvdfspCTG1JHNz+oVIiYwFUJnaxs+EQvvJsSy2q
vsF5mQpIM+QoX5izkun+VnPqnKFPSoLqb4+PDJc6JOt0KsNZ5VyAMKMB2HSXINqa
eFr602TZn59YM6pO0M8wDtDOPQN6tLffp8OaHNpS1LyaX7wETm3YWyw6TXCNQPpi
q/eDEQNnF9n7BTqyCIhTka50oLXoi9Q+t+KC16VlTo5SFTnLrjdRPAnmh1Hxk2sU
AwnKF0znl+R6cAPLXNwXA/yvDt6WnBWpDP5VSH5fLgx7w8319BjSjn7O/qx/3Hz6
36pRefhwMc9UlQ5/3c2K2/qgDXwqHnfOfzuka7Ho/kH0GDhM4UE2XvLLsQVsliY5
AYRH6sD9YoYU2jTXfTf5Gi3fTP+wgxybmkb/i4/S+03L4mYyRiW0+W+Q1GsK3ng5
H92x+FNsy1OqxmdRqqbozYoyk6T1/DjsGCTdr8zdndV1lkkd8UKtUXuNaMBfXb7m
wkKgob0+cY9ikCNkHWjz9pp74I0WiJ+BagnAS2dip8Gp/r7h75JKdV07Sp9XvJaF
hwHz0gGl7uHQ1H1041nbNIIPAcrds992fBzXIEjdvfo7AUfSlfZoL5elfaFG8qWp
QRobHE7s9NZ3i9JLnTpG0hYvEJc06V2nhPEaPkxpG5hGE+R6T0/v7vLaDPdYY8nP
g42fwwGpnqmq5+4GusuJOla7RAwPf9ozLX7v+V5Gk0sHhp663NMRErp191ai7822
hHfOP0+ftET12MtxZaVw9svZBUNX/xbe1/EeE3plIfvo9WEB9VBMlCkI3hgqlqa+
/ZS6SfD2A96h+MDeYHH39cgrHy1m5/oSBM2ZYqBO4C4oDyGgIZyihT8GouVzddOs
JgOoIZanSrFCVrCUOZv0VQ2zq/E9qgYWdyUMHwxViVthO1vAtIlnK3MIN6HYdFOq
jDU6g3rdDlarNdEg8DIGD5RnQWWqy9c5C2CzeVP2uwy2tu/Mm2vMqmwCo825+7h/
0xQ37qukNnDXHcNXVVjBJzTgiTvsehN6XOIkstgbEUnNvzOc/IWNONFWmIUo3dUw
2UkMVhQ4N7dlqPlrm96q2ocy2a/N0Zmy5815FguxpwDYIEhCz6k3+UbCl6CohIrD
IRYJkN0HgNAAQB9kYlbVDw20i9WZtNneusTO11W2FsSGAx95lB4Imha+pTrr+nV9
l7rV8yIlX6//HhAvFBslRudxpCieZO09MhOzwGoMMw6i16Y3Qc1A+WHFkziq5pUX
9AH1gz2Vpmne9A5QSDx134KHPaNGxaT5Nw0stQTNU0W52/tuuWq6t+q6B/+svzB6
qT3Ph47NwAt5j7av2S6AOQDCAMGkuF7eHSb2qay/kC9VzM5gNYYby3eEBP0qnnXp
sA0M32BhF2JOmNOAAl1HEC6J+vAWkQ7845rgd+EECvLEEj1gvvAqWLmyOgyPLsZW
0wzburKRo7y5wO62hKtm8cyesRwmBDtrSGdZU+6JBm80BXZlkFQ3PIkci0D8/01Y
3SJHfZt60jPJ8eTq/hWPREbwULNKTBWyPwN5eufnwRe6tUf1qLMLK3XHJvk6W0hb
j19IoXqYs4h+QStQysKkp9uKlZMIl5TY54R4zNOSrmHTvZNyNelROyAV3xJcLyb9
JlJgZPv7n8W90cOgt3BEFK+MQgqVpz+IEXfJQuUl4ogBxBHtY/pykt7cZY+uApny
SsA2mVsevzyWl8ilmB05a8S6SxHzhRhjRhPNXO5UPeFy2wClKMCmWM3kyvy8NmKu
IJVgwZAGWkq8eZQwhuwaI0g+ZK+04HA12maEtC2yXOVox5uwbKe2CLsgsgssTYgV
DGE6Uu/dDAqeoFNekLHR65SEaV+soX67PLQiVFur3RpU32W4GFWadpA2O37YPeJA
c/iJ5l2ols3yzW3Rs2G7Gj5eh2avoA2RKubTHwpvJzFbfraqEzXsoYIav3t9kAKo
/KiDE2X6r65FDWvDX4Qdu5j97DTMq7JBj7k0kVxfb7O7maO6XVK6vPv24BtpoChb
yCSeuyZBYWCjtbeA6uHQa27eeyLoeXAn1Vd1efP6ffNMgEaYkp3uZ5DYcBsq9NjO
ObP3QnELXKt4c3fSLv/h8Ns4+znENJFH4DZu9p0QLFNfKkP1gS6eiQxr/ZAWLctz
vYf7g3FBZ04ZyjSlF+NJgh2kjEh75oD3sAfUqL+ACH+KhHh3tssgvoBNrq35qR65
fypeQMVUz/exjEmNYQLBWgGXgArdEt2sr2nV23joia9OtRyMXuOmVeNmX8X22jXV
KUBwKUgJAw1oXaFQ78UyDJFBu9U7S4WH+ZFHHM+Ob+sAz7rA5mTs4YiLFWbxk9XR
2JURb9V9D76K/yCWWpjWy3E9Ss94aqfsDM2zSA79tdDIO0AeOocpCMbNb9L6ZECl
KPlP1umXXw7zuNt6CWkk+Ar00Uj5UdDYUobM8pG8zO68uabwZo8S6LcwePolZ59u
LeWkvcja0PAFWqnxQgu2ymWwFsz5lZQxLpkPzhYko9kChAqM0RrpgQW0N/rm4IWs
pbXhvzGVv1loz8jE2/RwHj/2PDk5FyF0S5Y9BVdJgloHl1UoTjJpPlI9NY5t+RaR
w1G/tCPUuk2np0wxENpKnOJPNpPEHj/9+OIs860R0+CUgUYbR1hAVods2wxTY6Ic
dsJKL6Ft/9d7JqSWpnLJYAdq1dqQVcQBZ7vatycQ5wMUxaq9QbNw0NJc8N4XOZnj
3u7XmtdZYGcXvSB5Cw/AHcYob79o03J3x4sJINjnG6or6p1o0ZIuG5/B+rexWsey
8/2rhS1JW9GZbec/crrOALLyBpAho0ZU4Kq903r6W9JjkY0yzhOSGDigbKlJ45hO
Yi2UQXXHJMPv9+i0O0o+MS0yan+KCR1+KBcb0tUgRR8tsvKwTepOw7zQ5jH9yG6D
ibrLFcH+0suCcBPFwA0NpEUEDsBK4q9WsPetkRkbSkYvFjKvpxdyyuTLx3TWs1AG
0UYI8l4CdkTK45q8ChMGgD1sT4bwtmYfMcXwEsP3DSBL5ZDJpgWgBizx6dkpsEjn
dHCiMx+rbJTc37yHyLQduPC/5+haaUMNszzunc2zx1LySi+toFCAXPHeonu54Q9Y
NaN5PoD4RcmyJcPmKSnYZlerpCmh2E11Pp3q2679MnKfZU0OWQ0XOlfGEJFG45Mp
2HY8P+fgup98dslyEKcZfjqqcpovkVXuLi7PYBUhvGG6veykd4TqCeHHOM/law6C
X8+txSAE+90akVDPkGZKLn2ntjtGs+6M/sjZGuJkMOFXJFwh50zH1wYf2/uNI9DB
xO0rwOiuJjjqUI34so5WShkji3WJrAClXUTo+0zVLOMgrTuK1Xn1ShW5iaMiFKNp
fm6g/fj2XaloL2RRMSscDoriS3o0703E3R+WTEXOj/h7R40uLSPsgVRwhFL/3cBc
IsJbxij5EKTnYpJYDsnr0esPDbVubc4u5uulIL/9qzNoIOaEva6Msy+P6fWcp0bR
ZegGiyw4GVnHhA24/PeQCUu6OJqjAbr8dXzAv8iKluzVjtvFrcn2l1hrKot5VcXL
06HLdbYcbuqvhtD7C7tSRgtGAZUrnldosjDKcFyOyWxeBp5P2RKslKhZOUzbXfJA
/0jkln7iica7ndd2Lk94uwCcIFAHlyYUyX5NcjfXQznWcp+gbbIxM5VMuH4+hbpa
gSjQRon4CBb/lmDXz6DvGrgcpBS1WvuFoZWXl8ggAp/RVRpGcP3pgyLtWaqi3Kb9
yJQB2Dwi5OyKB/gNbbXUkqAJYe95oXGmaxPOMWAAgDo/DvCDXc6DTJ2TCSWk7NoR
rQbsqLpzs55IeOs08f96Y7Lh+w0sEbB/TPWQ9FqE20Hr0OKg54SwrJ+Qqg348iG6
VNDh6WhqjnWk68aW7FE+6OeY8MnX97cR1CQJH5r2oihK4C2PB59xaOFdm7WevQFm
9JByaSd+PuVvsVAOo40XJSDhuzecMi/u4JTjtCH7cDqlsNZNdJnxDidBu95mhkHj
yjPEWLaOOI97REHLNXK6D2ztBsJstL+G3xVoAaUg9/AoHDAEXODVquwnnPZD5rNX
QEbVDkz4OwijicQq10cqLlPzu34bCjmPZlO2oigq9wrnEngMImdOyaMrEmdbJ+ht
2obQJa/P92ubSqsNXveE5ne/Qlh5oXugjgGK+HbA74ZjeI7gCDjfFECzSSmfQTkK
05+nQUkOr2xNqLt9p5DsucZKA22PkQ0aayXzHsE2qlDeLt0JdqWXNXT++0hxU5+y
FnddxBbZkUYDPfs+u1vbMB0GO/s9Aaybo96kR7rb5xL7JkbPivoFfAGruuI8+JTH
J7QEVRpEdYDKURSmtEdD3eT8O57+6uwv5Ol+RpOkmVSw7fWiOmtjOpUwI7hhK0oe
RVyRVAOfbPOu3bvJFtItuTOdkgF0+IBGmNoz9K5fNXGpU7+WQcbF/Q10+PpN69ne
xOQ/iTyzr4abCRNFm5BPt7sTddqEl9JT9ggB0FjzZS6YI+VLFtIu++qmT3lAvO8E
o9WP4I9nWZimQTbLsjsne8vAvcJKhVOM4/buW+6YvanZp/q6VJGx2gTazpypkyqb
HAG0SLyKdLDLtaa2jgBINHm7lWl8FSmLL952Q9d/ToWTeIIvoPP/0BDcN/Gvhhen
TcF1kW15OtGdBL9gn0GaEhAWlQUE2Uc+Ia260JPi33pRLU3b1e+QzBiBwLBzktw5
ivLL+G25MJyX1BrL50B1I7wrhKRHla/gtw+kxQdwz5QpoKZbf7d69p8DvHaY2mTd
GWXv1ea96cCedlTS9e3rgnRpSqe3Ej8wDBxOVRQg/v6NfAZ3YJuty2BLHoAJvpmP
gUMyWAYQ3sMt4r9ArvhOoyv5DN2vnZk2wa5973dSMlG6F83y1AodeeqyKh0vdlJ+
0UCLJHkINz3nMrD6D1bT77YgponGudUSsOn4IBl8EzMrCDzgMQbm6H8sy+0TV2Dv
lk2ate9cje2Dj9H5soJUSplVHlGIetKQSQOnQI/FxH9EabY2J49PVwFPeCClyDTS
t/EOZ1+4GTd0QYW7dcsS09TRr6BcJtNruHy/HUDirGIfRoIy7TMCZnL5GvddiJyy
6cyliv7x1fdLzuCr5MsF4zZKh9kOYLSgy05irKzColz14MlS9tngf01JWAn5sgho
MdqY7bqWt/qaJm9ZiWYCjdeJs5xut/5/dPc4vzfLXDtE0U7pXpvqTjmORK+2HLjr
w1XkLZqiQyCeeMOrxDppa5zlZ4qH23TJDbfYOomb1i08pbRLkJ/2N/aFVW/vGbLc
yk0c8KSR9hSXS0uDX+XT1d2QPEdECZLyuE5oum+raCTguFsshppu/dJ+d+N0snoA
FVxvM2damFBvfl2FWnVdXm1FWvqcIBmBEYfIyvPLgIjk2aXQdEaq1CpmfpSTLkIn
AeWalWq+a9hDdrcMmKKq/LFcldg35lSbmGB1H+quK3o/jTnsOjkwwcOi0TgD5JW8
9Q0C6l6/lwXX5UbnOgLciuS+ihz4ynqHKwpKT4CSWGSFsdnfYz6DzLJSkrhnWYtL
zZWkQBXyAmdkX6f3yXZGzhCgQUtY9RSvsBIAA61pN4OgT8s9ozBE5WpirwwI+wRn
TCNXVOsqXsXdHkKeYyCpAv8boHB/DLw2ISCdkv1cgfGEYNi+6na8VlHEQLsg42RH
gMrAE1RoX9KKj4vA7YKhuZU1hZ84Q6/zPK3xGCxv9eSYARkGps4PGlfHq6YR4zZv
vvG8IpdVPvTI5tBEu/9nuxrmOQHf0H+6Pq9g2faqSOIqS9tzL7nATHo17w4bS087
Xj4DLdWeqeiAJ3oE0DqDf4ttaAYiDW1nN6ACWew4pZPfxIJd31REKFPrQ3MDpnKI
sq8SmGeSvprbzhlZiaI9AUSeYpeFb3S7kL2NWLld3Ajp1KIDa51hD4hcx4uD9vJ1
7B2A00pveQO76fRkyH07hVo/nOW93jxcRTerFpQKbtSvIo3PwNH83Haecey4oWB0
LSanWGB7nR6X5cOCy++UnfRLlvuO97VbRHwjz4bwJGvDEZy9AGu5rHt1m6YNQW/O
DQDn5TJccprU8TSYgC5Jsxs+vdv2yX+xFExzDe9NtpddREQIfZcjBqoPgWaP/Qfp
LkgSRmDOTnc+bRhp7gUKmdhFYnm/U+WZx4grFKACsjMOuRtLHKLjE+9xYnAfsI/q
vUcn8+8LKMi6dDgSoqL8IXelOYsS+8famoL3cHaOa8S5bvIyGysG9W/7QEiHHeqc
s0Ajouq4gXYVolWES0ibWGfRDVO92Q23Xyz0gwBGaWtur2bHKb+wQjjZ+QwN2jID
La7KdxDJQgbWpJPpVoToG7XaecwrbKqAWaO6RDsWd3JdfNXFtVWjV8CI6sT5xWua
5febPvmRpj/keuSenbstRje3iRTV8V76OxoxFqqOugUZjo9S/kbsytBvkVaCmom9
Gr0uS4/GxNVKts2XS58EcAy5teh6TVB/6xPOopZiLzyuNpMxwdqCO5C8D9AUIUp/
QSSyBJrkUAwyou9Y52h+N5tPfk7Vu60r6Y8pLsL6UliCqmEZWfRoVACqSaya9zM8
8bIotnM1cp/aTGqEldILSUyC9BwXYqgGYJLsI9zh2ZUbz4BERNfWaz6IFp29Cvzr
EBGltRKQxbYONGcqx5rYP199Zjrc3blYE/Vf4vUeInTMXa8OhxJbIfaiUEm9/1JX
muLU+yRYNwvYQnHXPNEuNlWmepJrHQvnozmiA2y08qf8jrFkXmVfVdKTALnA/kn9
eakjPGgaq3R5Jl53+aYQRUF3/0Nweq0l0l0XlRHTFEWVvCgo4aMEEFNB2Eu03p+i
3V8Yozyt25xGzk+97Xp0q1p60Zwksn02OOmfuWUnFeErbD9yUBoHoKyyeLGixEYw
FR3VXqfYc2yvYxkrOpL4vlZkr75tYTw32Np7icw13qrmYf7T+kd7NnLKCGF17rWE
2K6hpAZk6JIrbJgG6fQQoxW/GTy/hmUEMmizrDYNz9Xm2tqH5+neV4uWZdowFyDv
G/9+GM33yBsYpXaDPQrDXwYadchJoEOSr/+360pbGGm4GX0oq5jWlxJjXbXZ4GrQ
LDnvdsdF95nngIiH0MUaBNu1wm/iBT4OoyKKcaE4BDXGyCISui/dHgjQaBSdK7qJ
yUCb+vUcYHyWifGnTrdI0Mz+OJcsHPWoWg9lVXi5ORo44ERnGagho0q8W+Zz6SQ2
zTMl9WRa0kHDnIHSJ4duehaHl4gEkklq4vjbrx4kjLq3X4ZxxgXGEpFUvHWKWUyp
Mj0YuRhi9lLtzYf7VB2IiFpcWYYx3A1DvPhpyGVThm8YNTnSPzu+XRULtjphfscU
Z3DJjY3VKglwrybTHEpc133MGbq2EIfVIlBryaG4EL9NpgSDu3/7nKr6T4PwusYl
9B+sfqsl84wHa4NmGyGPhgut4eWEbSRb46jndYc9R1qdB6j8nwtA5vpInqwulu6G
YZvb85OSkX7ezXwR13eFKUMaJOlshdbM1m6t0Nr0v/9SKPI71Kvr2EwtKt5udGAM
AgSU4BNlgY8WdDYqLWZlLwez1MRKcl0n69AxLiJde/xu6HvkSWycTZi8U1ZahKVw
iT3UGiZ6+I/YC528GTYdDGb/dJP/Fa5kpzCpuysjn7C81BWbbEyq5Y6fPdJ59mkc
v5JLJoyrpvtkw78Azi/eSm0tEwWnwVpDNnvXusMe7y9VSQWmWmFT6VQ9uImOm1NU
KfRGxK2Q7sBMJUtwukVok4L0aN+otxWkMaPMQFZxE3v7Qap33/CBcmolHLS7DZ4s
ciJIBkh1AdpXOJOXZwRBrwzxhbKMJm1V30hfWEGFawUWaX37HaZ+TVQc6eS4+vyo
9ajFDv1bEe5tg66rlrxtT6LM/tTO4PYCTr/nV9botwsL33kpz4E7B311BFcZvx99
X1yKBxYzt1f3F+5/DEmhSoBN1ZgBtJqCCRFt+GKY+JJkxvZwNmO6YRPbzPYLfLJJ
rbVowKFiTpcVDGHZnBrMdLF7v0bESpqqTkbsSE7bl+vqtuMxygUlmoLoESCEBaBP
WjNCkwBn6nfRhaRarT6actJI+KEawA69fIg0hd189gBK7UGGvAAXyNjF5eO0rC0y
qexLIyLoc23PqrwhPDjqLK4Xw8iEtCGwiOitSkYdsN5zxe+RK4oKI5J6NhAVMnwE
5Fqrrwn0F+oFSeDgCiSNOUDfcUScuUHDgR3HMMKA53iVTZM/gT3BpmM2bVqeAE8y
kwW2yWmBGd8tNDtxd5hX0oBiLRExHd2ZcSFdQqRIc5sQgDVrrE84/3Pcrh+T1igN
sIL3lvw+9KWiDKl9PdtZeqB08OaK+a0mwNvCcjBTSaApVU6oe4l4UlB8bw02/yjx
A6CvYSnZc3tn1lrVtTTZFFKYLA3RjotkUuNlznd75dvlyYhfCiSY3cBhQC+YpZ/j
PFO913Jbne3QgSzoEq/UezoVe8Z1/pxMZsx18wdOhlu02OHsyRPjtTFV2x5vSFiC
/znGfHmdGmGsKKH4aAbPcx1cRuhX/YTTGj2ZaGH009X4znBu3gtxXexJPYNlnFUP
suG9VPn1WSzjRFvv8S9z0b18USeWp3xmsRk8EaDeQvlzba6313gnb9nts6w2iuAk
zhYALkRMjhURn190CUqUVtlbIBz6B6w6F9klqXaqCbm4TvlfjKR5tC0rE4wWMttn
g3FR+kHJ26ooz6q00lV/K4t6Ct9VStwUMyjDHGCP6d6sJovP0IN6JhIrp5Y/vm7M
22YLKpeVrgwa6jU+wWKPDaI4wKM2SeafeiaINUkBvSj01XPP8Nnm8XmIN+1H3b/A
idnVtZrqz0qIJ9J0hyFcEyb/8ej0p9nLjuvtz1tx+LL8PCPOBG1UAKZc5HQ8DfHl
7be1JLQVAJW/eG9kO97AWhF4J/pH1Pebc5MIHhQNa9LiwEPTYzvT/uHw6Mqz2ZFg
i8d9+/LDiRBKr/wQfx426CHhyZ/qcK2r8ZiETv5sy9O3uqnseVvXSt6UFQAqga4Y
TMFmmqPNKhTVU7AXpXi2fKNzSXB7Adk1bjz1acoGcIQdlGlUzlC8nYPAWs8rpBtE
hCAuCfuXZ5KD6sbPCyJkgWkrQ+rGRqcjSG2Pi1j3+AI9RrgpAEonSXbM+1YOFRaH
TDnyxGus/jMIPLxDsy/5+Hk6aFPuSAnM+GDuBIjRKxATJhWCd6DGEBcBissL2ALC
E4a2yd+pLUFQZfQTZujV4UVubHyg6Gi0QUhyP7x9NvROoivMZxwFg37xlC+vX2jK
nlx0eRNwpxm1LjYjCpk2OGJNWAqvlEFUICluhjrPv8ZsBeTK84WzhMSLZpcsbeKV
RsWV5QqDQ3RuEsKW+QIeJf8UV8UrIgeW3psTE53quLUQP12cFXFOMBaCSsygizLD
rzKpJCiUCVuPL9H6raFBMXrQXrXoDgn5anGJpEXBjKXsdgg8TSXQ1R8DwbrBL3pV
jynC2CVL0hZ9qL6Csrnj6pQPdN3M/jHwxAH/NUubbCWwKIP+hVY+vKIvt5o4Ku4U
Udy6i92Y+rprbZqoPo23SeRa7FibTGaaBhOrZitbzEdtTXYFeq+9r9V+NvWBYitH
91nzgiVVb4s1ZEnRH/VkNBrkkndX2tZD9Ar4ILfPPIsuVulwb9YXldlte/CcCoiw
njol1YWWT1zeCBslFfGmE6c4KEgH+G0PbSp4rEG5Vihf7zaHBCJWww2i/DzdlEuX
/vUx755Ra45SBr8G8g7ri/27v37mCC3j7txpoGUsXtPb2DNPBjtNij/Tr2rglDtg
eb7zPXj78qyl/TckGYoU99J6iI207yMP3mzDD2MFNVWQk35wt1oUhA5Wa3nTmCBM
H5ZpX+z/pVYDdYa+rG5eXeavMNTsZ5NaQOvE7Fcd4+mQglg4isCbeZ2htL5pEvHr
FEeTHGXUXaf3lyoN860XLspTIa6jWS32Le98+hpjLyjb+Pok6RADVkp5J8rlgJYZ
v2kOrQaCP6fCd0S6LWGL31+y/v8LbPg0tUiKk6lz//ZOda8R6WBrIdv+tei4/Piv
ASwiy2VG4/9h4iCxxRF/DR0rmRJMxb+AJKi/k3BmXNeHiCcqahdEYroNkroeH9Di
3DH4vKd2c0Qnv9bRzQZi3vOAZkpa5I2TkU0W8uhozTWCdsIoc2HtixtKRmJ9J6o3
LVR7012qRJrtcmjkfWk40s0kG957xQQQwqa93OVoeair9xASBWmyovmOH4E0rXfm
5k3AKOZeArTUE7zbaZ1qUNVxr8W94ZOQlZcigs2cdHJ0Vel+kpdP7dI9WBtE1eQk
HVNBhqa3OIspEJivSxM5AHN5VBd3E3TdMdfQgQ7rMBHE60Cbb5vAJa+78sW4skLo
BKZqgufXeLRJIGojhQc+ai7hr3k0TadnJ2cvo3WWTRC9YHTt+F9ZL8OLTEqPhWyF
hhFe+yX7EJVb0XwmwAnAigtZNM/7I2cFJNfIyEB2t6p4T2343zL8xJU0nmzqV1i4
vo99heiCNnbR3JXaAOnUWHJdMhCF6qUUrQJiR5Xqp4c6kQxHE5KVllpuVCaQHgZS
NeIpdmzJcNPeluI+NfSiuw6VJuDKDvY96qiA01ARyXuUIaIkxWlFTqfMemXWUMhj
l41ydB6z4AE0el0CnxwUWUzRbS9E8iersByfNdMAil+9SzEa2owuOCbSI9YjU7z0
K2uYwUQ0TqoXugjg2jFyk6b/l4W/A6aoAjywVDoo0AsQjgtlNTDaJzESGEsskjRU
tza/h0Ma524aCGyJVxCvEhH45Hu6lr8G5+ZzGCjo8nss/CLbAbz0+VYB9UfS/hwi
4MJRJgK0Uch7mZyPp9hSJDHjERtYrQ5RbbNNQIgyISAsfHx5MIBwI5kj2/Jiekle
nkTSjwtSzmYkMzVTcESNiE3tBL8U/c0Em9gXTiH7VILt9H2+qmB0cgFgq9BoGiip
SXSjdxdYA7D8PtBGouxWOSBW3kvp3iRxIQU9CpeJ97cjtKvLuOyrG1YkqtUAi54R
imi2c6LrgK1folkCOYwHSyy9Z1qEPS+oCUNZAwOm3om+l1tLHlf/d31lrlcXg9lN
jnB5poAUrh9yywCzU5Pu6Lws8HIyieEkjZFHASUv662+PQ6w12HEN+lpSbN/QP+D
NbgzSVujkGvLgEUl+gc9kolsgni8YOOALwxPuhjmsDDt+ZyOykhtXbPngwlWIELg
awPGM3VdIbmqn5Mq6dkZFJYmh9hEehaITd6gQw+DEE2SsGoQ4R0KN/ULjsN3Rncq
xG+7k7gfpzjPM5y8PgYIHj2hfocnDlSa8yg4YeUoxbzNirY0SnA6ygKC4lloAluJ
LwGzGfLmdpGTI45wu5L8/WyUfif4UkbW332WKbLcwvXXCwCcmcnr2SwpnqHGOqpm
BWXvZrxh/rlnEzGgrmCb7GqpOmhwHl3oEMJGJrO+vJWR9kVcDpzkmPtRwDP2PvMC
yIY4i4mVw5OtuI3fV2AIU/tRko3FmBw1dKeorxvQGGJRMpNND0UwVjIX5YMeF/vT
n3rbtwY6claaJGdHqcamUuzex6mYbdCci/kaSmboact3QOpI5DO1wlAjwNOqKi40
fVJTxKOdnO6wTzjvIBcaNYI6UmAthjVMPtmdVnpQpK2xW9lIo1pd7aC+UWMaMdQt
kL/B9B/SRBaTMO3eGLjhTUDI7eKN3F0PYHOHjq2f70eKdTiD0AUOjgidxprN04vR
ceR5U89gE3vMvyjHotDEBI/HH6AXKxEgBJliYnGKyQlHpX0BcTcogGEyELS2Ltxw
OCVP3W5acW04itjavb8bQ1L3DriEm3fYanT8qPdvr71jGErlcgUtAhbJt/s8ETyR
q9zuL8moXJP5VlXlP8YJYQxZM5G6kOpHKuGU92X/cdrvlKjRMBvgXye9OcGJxN3U
2IvPJn/JgONSzzaxWfVLLeq7VGvV1JK6ymX+JG/qn09E3CsDMZpIU+Yl361XD3gi
yH7jTHHIzVdEhtlQCFn78eOHxU0RObHGgjByOiVgByb9E7TNJfZb1zkivH+d5QhS
lh1C88E0S4pz2tCty2r6jOXd6nvyXcjFlJV2ab98qnqVTMmikhzdYZZ+wvmEv8UO
9QMUMkWSbkqB1UiDzHz0jFeBVdUUWFDAEVC0snlegquA0/0DFAcHHHijcg0B/VrB
rtjZ2Lmmm9zSsrZTOOIsKksYYCKvV/xbRlNxaihu9o7shtkZ8PGClY7+ieK+Kc5D
nXU44txNxPc3H00HuOlPeUWJJwbf6tX6WSThUgpmwL1jXuR5JKd5nA8tlBXN6krT
fSSGA8swLW8ceP4fFptbJ98u9VA/fTH7FtiOwf9/6fKWPRVVTGAJHdXBCotfnRai
1keMjIBdPD2hZoDutJQaeI7Szpr4NKvw9tF+03z7Ij3ia8pZ4wL33Zn0q/wu5hV2
KMrLU3xVPdJUtxKM2ceCjgwBEWHwQBxoQQ40DAVKeNRysomCOSVTqFztvWRCfCuI
/+zwNJhIno77ggVh+17Vh11PeYiFsvCnTIhM4FxYvk8/dOGAqYAcFghglTsO8vWp
MI00vpNOfYGPlyk3zPlYxYZ3myBLuYP3aQPOFMFnH4mqck511roq8F6qV3Guu6qU
SIsJGmlGrrqwfPcZUBhHzPd70nhjZbTHb+LcX7U9oDl68P1j3uD2iUspHIcBlOxY
HPPFFxT04aGj9gXZhk0bWpTodDm/lycOwaKnPGgJte/wX8GQfqN8OQfeGnurydnT
t4FQ9yIM0PG5hqCT+5jnph2nGPFQyDdNT32oGaG1oFDfeA3U7f2XlMuCL2ao+NVS
/cz0DZnbgOwIM8oAZvIxSQ8Tt96rMJF+FRPkfNW5u/U92JPDuATot/Wd0oqUaGqj
kauT5ac0ITXvUDlHV5xGkgv4yKQcJd/aovb249O5W6/PBwPv5ln/1DhY/aNCkxUM
5Kc4fiCTn/gJeBm6B+1f2Xc2HIKnqRCTaoL85N4P8BJqB2dARpaEAQ5kpfR8zKbI
YcfsdUexx+Pcy8z4OnODBWKfR3y+ivKkgLNghdsYbLLZJ0yPiOmKVLAHIK5YnXSH
bNbz5nfgDuOCJ63wdc1rNiVqJNOh7/QE0SmmPibXcdpwToMn4+i76Kn7pN4rY6aO
oxvba4HD2y9s/IrCEpW7H8xgvJN5wAUH+izFVWoj8JTVLj9J8bfmUTe93d8bpqUZ
Udg2HsopavFzK2TEDs2k9XaNH4RDAyLA/8ikbzYT3lckA/26twMTgX19K15q6Rwy
L9Rf4jX+QbFi+Yrl8SV57RC+bHXrlKHmjsRgu5P677+xCahbXGvq3aQoJiAufo9M
8D72wSYwOdr19asy7YHECbFur1I56yFeh6rgdXPyZDC3O5gVAm4JzAKsEGSsMYA+
g7OFtixxym4C5UaB8cL3ZEAf3djAfvJHuyj5eDc1EFH+pWB3d9xIjzQdf6PlML0Y
5LftzZer/hKaiNmCXi3n5KaBVkMOEOmIEM1KKe79Jee+HEQ+/nd4+qpKzULQOFca
ymNqgkDDrNQR+t0+0N7j6kvM3XiKdInYDNyYQvDPjV2MitbTdO7x6HNBPYNUo5FD
0K0svvQCi6MikWgAlZDSzk+JWSdr/7FIR+LS+bsobm8PdYQ0mMrqYr3OlPD4szq/
l6he5U4Oy6lQKes2AK65vnXmwPo2l3yQUkydBYofm4EfHGNIEo3uCEKpag0N1epI
zpm2E1GElUHKNw7cvEs5SO/v5a3lB2IfJA80WOh9MiAkd9rd117zp08OulLsc16x
EFp5FIKd499ghK6uIkYVFy6qOJ0u6oEGTiVLRRAkhwhyOuGsF6JfBNG1FkinBmPp
f0juGrKu8G5/OTzzg/4ea3z9XijLQ1lttBdeIVvw/zGTVROFCzwgqKBo0Zb4uv3P
oZoFNnc+MEVo/0CDQu3jYoMfeNGcI1mQvLuhE+mlrKUtwIXC2LCllAzaq/s7C+AL
kUBoHiu2LT0XPFatI57PbAqMhBzxzpvCeOlKF+VIKSQUR7K2JwfmTiHPZIWF5eDb
xTxdWBhgfbIrd0HeuFZthV3Jst7qCvSiZihDJuRo1M+3pVCa8o/wCOrJhIt/gtoX
+v6Y1/IEGiluckHK/mqGYnHfI1UbNYRikRjtKL8Bq9BlLE5OIl/Rt5+6URriQRAJ
/Mb3Dh53vHf6hWf6+Gxke21Gh2j/zr1722eYbxMewsOFNqBQzLvygt5zS+IOHb3R
chDfagupz1rhaxlPzPY4T4Pj8TxEyUByoyD0q026v+32itIFdeW7nUgWCJJLODIb
L1RZ71TF2502iZ1Xqi7OPOIHZzxvvUnNal12D5LV/wjrNa+c/tD5F7UPddgknHu/
abalNJbNJ6d9itBllzwYi6DBu0fhaoNEZBD8XIVh2f9j2m1ZDCzN0gVBjBr7feqB
CyqaRFdgmE5HkgH7pKEnjiG22R6NF/qWo5dZgmQK5nqjEgEBFEQHbGUu52Uc87TB
zTjBGJv9eK9lXkQsMJr1pveJAJ8R3Sly1/zCVh92mnL41iR1d5GgKpUgvWLr4rRI
pqjGnnCaJcCz7u/hdByNJklfW9Wc/kAYxyulhk2do/15XSk9I4E40eziBqQgLdlV
FQo8FPEMll0UDwokTcXs7UCYW5YVyCuLYSw+IYjR4xEP3OSew/oLIBsyCFuUZCx/
y57WPaq2Ia0kAm9jQWfMuzuj7yU0jsxMPknaMQZpBsasnrr/QMISv0sxdHm2mrJI
+jcHV+z5xD0f6ProrkYA5oNe43sZw3C6uYWeNL0ui0RWcYCUk6EkiR4nevxKx8gA
y6Sfsr8r/Rate+q9YDfl6/i4yWBISHVrccqHfHyBtltfZHZhuHHqNxU7H6R52TMl
PPdxlPGztfbvJZDgPF3qVZK6o2RXUTRgJNCb+U6BNHB09ubNSugY+SBENKm15gFI
0lQLMyQBdyWx86Jqh9CMnsG9HHlInyruOQ0kLH9pOrgJPcEAL9ROzEvo5FTH9zAx
JCHGm5WXH3jB5piqvh7W5dl77KdLkx+DgpYH118bH21nvZHT9dOS4NVTshBSm2V8
62kTSeWNRPWlNGqgbnLP6zdcp1I4q+E8hyDn/T8TMkyPU6ozHtD2jrOsFA4QZgNZ
llJK32nBsUhNkvLJDGOjal4aeoW3cqVpdeCopDawIOnMMox/R3deIOMwNou1Sb9/
jRAxQ6/XPyrqhcJyXTkPgoMJKM6d4z+c5ChPs2paNk6Jl8JknNJLakUUkQMquck/
+p6XvgfkY7o1mYjP/UZz+xzG8CHaipneKa2YO27/+wM3d76t250ZwHw9WT4Yvx6+
5YChTEvIreIHc48zJzvU4N+CbNP2iOmJ/pIvZ/nPi9gNaregIdR5woKj/Xb4/j2d
vEZWp/wSfWqsMboirXxE09g5gl+3gusUMQFfrpvhn/C+4mgF12PD+21YT3XPaDaj
f0sAV9niODMXecEI8F85kxkd+U8N28zilKA/w70tzuCJ5qjlyF77bp8vqxEgHatj
8WsRhCGYs3uVHJp6vPdXWl9XwzubEBuT/mSjQfm1D16n5DI7ioFg2HhzgdAbrS/c
8U6ECbQwHWSqboSUUIv8oyBccPTs4bEL+S8DHZsGubQ4RpW+Ky0twrWkfY56CyLZ
z4RK743jpC1KchaPS4KW/TCNEFXX3YwSt9YF5knEdb6+BYCm3tTwBxGVThig3SZy
7gyEFvlAqHPX5bgk2CQeG3M2cu3MgW/aerJcUUX5F99KAKhsKqGgW4Aj1LIdRqHZ
jYS5bFslNBDzDbSzezQQd52KMPSFhcUDDnq2Z6wB86rZbA9e/ViH8PUWI3AyhedX
vcaFbYftWVEhQG5XXU/rVdhpYlW4DtesqhgFSHrygM7IHIHAlJGwixLFd4EvC283
Rb+U4ap8avbyc5tyYnlEfeP1yG1jnanNwdZ+f0v0YOIU7LRsEpTucnzsM+aSlsHy
nYXlK6Fmm6/Cb9nsSbHxgo22jCsNLcoLl93B/eEzx794SWIgvB72jN60cU56A8vB
0oiy+3wkLD4eHgGYFALKfYCN1nyKGycgF06zuspgdRalqP2Ypp+yWf5/KJfCVs/7
psypZfFDKuRHW4E67GQcvlnziYDfARc3+NdyoUSZkFsz9ymUhmB6uUqGcR0F9Omd
KdTx7OzKOVu+bLwTH6ou7iRwOyldN71vFJdRlllJIJEe1z+p3pvUFWFEoafH4uc1
Y81jcGE14OBUNocqWFE8/5wHXIWq6iS53Yd3byTbkYafVqOjDu6PLTVsPuZw0Soy
90fzPImrsMOF877chSODx6f8MW6gDp3jKbQScxJDcJLUy/u3al9L8PXc8ewgDI2O
lDrJfMfbq5ma4BQOGus5tSxrEFg/lUFJeWX4E09p1tqJRENT2P3u5xeoQQfbc9sD
sYXFQWVj6v8QsGl26aKppJS/3Blg+aeW0Um4jF8mojeDUCGG262KKXN1VUlbLWoN
1jUiAeqxO5nfufnRJY2vMCm/1KtyUXwQGGfmQL6+Ka+gtpy5uG+huyqXVjQxFstr
0+AI++Eq/Lre//sodJkrfM+snXfAsFDZh8v2juhHBjLhW93w5p8dayPmFbp95QDK
AzVkC3DlyEa5uL4zj3PbeH35FY7BCG1ctmWW/1NDO2zaX5yuL09e+0XYM0ms2zuS
vRQgLUFSDdpCL3Ukv8DOn/tpO+A9Y/5G8M1vGFAekx4oAOOgw0GCwFKbgxI34Otu
MzQSOcrmb80Fhi+FIvYlIUgCia/FUbypy++bZ8i4AWhg08qU1c9aqY2hONpPLbp7
7cRCyPiPx9KYXrnBoN4NyNo0kv0S1mu3N3E7ypP6VeCKE1DQxGdubuv25fUgHPGx
z9cchjd/kFw/tbFKM1it/fLArgca3vaNtcdrYXhQkBNZOEmcX/YJyMKUCnKx1HlX
Jf49l0vpIWhbewiZgauPqdDJRWE6O4Q/dcGwHy/VIPD4efOktdQiV87ksYJjxrXf
V3B0CE/3VHd7IqzKdHB/TyQrSYLuXi6hjUPOicvcHvB76m+EUItjLpoJ5L4zndRb
3Z+6fIeKKQRbWWFNw/i1nEfdhC3CI9ILMXIAyKHAz0QmLqOnHlGm4d/k3MATtYqe
64IjN37AiljvdjVMXhnfeo1+Jtfsz0ShcMyowjAyRDN/g4ZWw3xn6PEcAHbI8eIn
6QHYNmV6OFVHkbdVjZKrByVqNGd0bI8gjQSZfTwraZd36HSYX3Ykmmc5ruBzmXZh
j+j1YD9M0pgp233n6DPB1yqjWXoBww3+dLayptI3Zj3yBJdSZlgHZSfq1O+qf+wM
B5bZ/yxHy1XYvRO3cCZx8rfvUffgmM1hWZp9ZIDp4aojWyU0HXVOupqDc9uJ68Ez
bsVHSMddRpOltIdsTCKn+zRVgljjqDAmnVuyqmvh1ytqV8epP5S/KvMzVmFyLlNe
MlMObwsDR5xXqIgXSSehKEUcIyedpkdesCdIWYX9WHdBleoZqE2HuvY5pYrrb3Pb
Uj6w1c77Rj1dawMPHl2Hh7noRmjidrratDY8b/LaF4qtaNIVcSmgBsQZt3765d7F
YoKeh3ACW2NAGiqq/yDLUUiCROuzblVCkxo40j34X6N0DGHrUmFM9qC67dECC45d
jClBWzOBCkxj33sQACq7f0LZijm8sLu5oxZT3L2bN578VHYwcIAphhQtalDHKYZq
lRkyVACev4+zMi9T/tQLRgv4uyOWXygXvwHJFPQDTseiFRUkKPkJNtYtxyO4qBv+
aC/4tSS5+5ZGcflnRFsD4PWsyyQ1jAGAEvf7vRhAOV7ULjNyBLWqmiibOiw0niCG
LBXZUO835ODOyzqHIRxD+Lok7s2FYyCL9211BperYLrhxnCs9cJQZxK+c0zJhqEC
zNTBdT3cOa/uwdnHvwQhiwgQ7il09zMssoHHGENqtrurzgdGCdBQhBI2r5iR3No7
b/z/sgkcrCNoLKB63dSYGrV0vxvKVpjEZ2QdQiKtV3EZ/6OaV3z/y+VjwfGZtVgW
fJHhbwU7XFk5bukh4Vv13TOexpeYdE96cOu9fssYi16060pgVLcRw3zN8zjyyuy7
QCLKIZEVaIhRIbi5rshWnqry2uP9aagF6fWCFvP9V8A8dhqVqNueRgVRhfVBqCOJ
UU0mvPpvWDz2ib1iRrpYorhgLxbMrm+Bvts/CiVUZSKFyrouEOEtfcx6aY3Mp1ZX
1At2kcG9Pn4ub+Ft8RtXdrJrKjzlAi8oCmf5v+v+FCNTJjvOVSCeCQOPRsVhJOiW
Lm/j8AjMgP1zbGwGh3NQ9vR/hjRWVuYLL8YzgapFRU242nebVcFzfW2OryOi7GJ6
2ZtRLD8e4g7GiyFVeyTNNRHNL5Evc2wQIlFLjN+j/wj1BENLpWKLdotjAK71MoJ1
eXjW5H5Tne7aIVgsPUy9gOt25UN46Xu8NlcTTJQGWqXNctTRN4v1sy8VmrWndwSz
5erjqFBGiwCxs2qD9uytxquUVpTWu/Yqz9zHQXKelTKmzDDxvf3/baNcsEZMUeF3
sVYYrLZ7YyX034F4obEYBYlfWcNBia/5XZgg9wNzS+6QDBz3Qhe40bWejTz+eSaV
t6BNqH21WRz4BpqfBN+TrALq2RFSsinHIiNoxtJzgx/xcRTHEXM7wPqCkU2bCUyj
uroPqhDUacclCvoiBA7zhELUOeoD2mID9GlcxNkMRAWhJoD0KLK2mHONNgXkCLi4
Cxd6QH1QRLV/bnFGDr5BLmr4/CHQDbinwRH6iA9deNqBBvYLgfcPy95n8SR8y98X
XWZgfZiUjceJCeUQ3sFkJbY5SpTv5VeP8WmwtHQx7IzVnHbNXdnq6LNZBZfdv9iz
lUKaO5QsU181N7Syqd3XIeIxsOhRzKy95435Eais9SZaZmUb2Xe87Dp88BXbme67
gR0jIVYsWfeHPlBe0v5U7WsT+f31/IfxOCkCJGiX+uAfob7YurbBmjmf4QiG/Li1
m4PNyjmfnQCRzmrUNtsUUdqD1jd40ot/27I+beM3Ldb3pGTYsQ6ew34XzePQdt5H
0EHFfIu7pKhSR5Ql8wCaP0mguZtbQzAhH+Y9t6AvINcwKtohnvnzaucceBQTieXj
oNuoYFL7iJ+KCPIqgN9w2zsy6kMlCewiX6k+viZBbi/zv3skaEXxmKn9fdaXFmQ1
yZ5uDolkUc/L1MZngglCxlb2JN6Xy11oqZkgpIX755N3TJ0ENatrq5Y5FE0h90Gu
g4wEZ+a5NyFgDGVkCXUzIUmnYrt0aY9Dr6LGhDryDb/izf4OQtJvNCj+bZlR0fc/
8hrcIo+udvmKpZzrvroX94vAymI3608BJqASRfR0PSD1A2Lcp/tLCC97nI3cmHIH
PFYKNV+7jTMzt0x/zzMzdbbygeNzMtd+Ay4NxF48BIf9Fa50tCvXDcPiXdop9N+/
r03MUjdCbIIcOXCm0enbw6j6bP5UxFSAIgPxa3H/ijjLJ49qLn9zCBqaH0oSZnwc
FP1ys9BrBmsxpFAhTrWdB5tM/8BezSOPtKGmXudviggYuhGIt1ngoBKsCjSL9yBJ
fvh98B1Vpe+kYfon4sDyenzc/HokZK85LWu2bkPFw6kZkC/thK+a3bC6CgX5WU5e
mIhkwaP4nHHY1A50N3OW6Mo+rq9X40eul7LMVp0KiO2wezc617+hL9SoRRJigXV1
F5UhtlONvMIXLDfIUNkPOdYk+5R2AbB/wKNeJYY2ZDknCPGsCx7xMc3pjvUeAxYX
colVXgllrHkCay0u2jE/GpaplOWXocoYEa0acdx6rBxRW/5kfLsvPz1RaBPAP3Ko
BZpvuZ11Fxyn/Yp9y7cVKH1SD6c1JzJr6JdMVfQgEX1S0nZdHlqSDlw47qqJR50f
2qIusx2exJyFQguYd7N+Ys4bfN4RDBk+Woj8wFICsAomaI270h6gkropRrhNOuOl
ptBo2MQSdgzGbGX04+BJfXjwRXJHrU4Nzd4hc0sLJd1Zw8r0sU3fgS13pVZ8i2qL
RrEY/6Mcerxv/LxW/x7Raxj0ZyVZEFDEEfdueb/BU+dJcxfK7U6bayuLvRQNYPPq
TKnfZGLFghaDoSGKWf1ZVkkTKZBSUzO7R1IoGbHwgAfsxnoeKyyPqfOvgGuo/UZJ
EwW/YMhHOdujSbw5UQQvaxKAa8fzUFWssgiv6mXBmsAalvLbzMSdiiCmliVA4wPo
vdeRZoU1VQxHCV2v3MPbNE0c5NAT2ahq5IlJjcbUYUp2T5au1dkkuV43/wJLXngb
gXA+xHOUW4jRfY698GLQ23v4uhL/ra7EpFkKgvhABOq13fp8IgMsKLlLFfowQHfP
FDRrgQqr5kBrXjO/BIx7ioV15BIZIBgj6dC90Qas/0SalYE0QXA0z9a7o6MzMPDj
AbuH+/84CojrQYBj4EFCxrTFHgAU1Pj/2EeluNjpTA8lCk27dSwjQNzb88B5mqrX
yV5vn6f+Enpxz90SJ1wT+j1TeCeKYvcg/RuNkm40228H6SEbJE9T3cMYNErETlEY
zcCiMJs+mmBo43CdHjR9qBFd1CG6jqfrV+eymN7SDbj3k1ZdT65YjB/7eOsJ/dFN
Xp/zKso8Hc2mXjDsG3iPWOuJZcPIlfL1HbNyX7JM6GhpQADKBcQybE3j4uxz+azw
GjJkMsFWsym6zljMemyY0/xhxkj/0bCSdQ9PClGroWYjU1U1rKpNYLpT1yFaBqFR
0d1v0D0lAtiW58AVSazfz8tLaRuODrWiD5hEPhl+PvGR4vPpSgWbbF5I8Jz3Y+vw
ieXr9ISL/8yNlkmjY9NPBuz4i6PuSILVFQL+0azmJU9OHtbabmzx2E6tmYjSE8xp
S10cjuXx3RVJY1WXh3x6w+6ElQur/JyNX6hSg4UrHDGiaLxYlRQGAuAxyehH+JFt
01ti+ChUj0P5RwRD6A3N9zws7DKouuVBpMaUKbzeY29wZ2K4Lz2QYo++4zSyvnSV
KtfyMiWGMvarCu0PssxQu50pUEqmnn9Y2e2rGEgRfMqM6c9baPxHRzUoyRc6J8B5
I+12uLzhUBl/ogllNPjdXQKsRi/GThMm3AdZQKGFtdHQnPRx7uBNrNbfHrGdfDFB
cb1mfaWdoOqTR4UZh++p3zftQqDtDAffUN5SPfIA5gPmf2Jv+lVhUJMADF7/XkPZ
jWWArKHecFS6baAXNduwj0pq0FGGebkQfFFRuCXgIp5OCXwkBZ0NH12auQkrCGpp
O9apEWS7X5/DcysxUgHrkmd22OFb2QvkNdWveQPZjGX3SSWUTZ6j1UeCr7MKg2rl
liYHVBW6WQ192pa6ggz0JzCiMYGvAD0cwzBpm/LjuRur/oXWaaTac4r9S7xDmNyH
xuduSWtQkY0OP9ffOoP/f/4uV/HG5f37nj3voaZ7Lnm3zx7uyTIN+INnn5lgHsqn
QHTkIe52u4Cat5XgdwlewGgpSlr0zWU8UQw/SMWBj35gxCrFwjp2IgbXG45gLYvj
/8OfrIuZykFASowQw1XU9la0MVwGzZKKTuIrrOmVsy7xNuE8rwwlCRb9z/IuBduK
nCwEJsmhyDPPXz/Dm3R21+ZO8ERyKxD5y/1nGTf2Ae5G9jL1GJA5khdMEe9vNo1x
1wFelhUChmtP9p+eSUBhWyCcw4A6QtNimJnZz8pnCDfK+FJaXU0lsRatugaugnIS
nou3lq+nmyZGRDBNFSWUcl2/Van9lihDbmzWyWnD6p4wMPIx8mcQnltLWBRkjqYs
AyVkMEa4Xns1VM+M9mTKXe1UU7kdnAGMAEJQirjRlkmzJ/9+nHUnrlj490MJnhIa
HeQokgOih/+gjrlUf2ywnOD79e0oGORCLRwMNG5Y/dXmYQNHP3DYlzpN/AACca2O
MX31RJkeMxaFmwIH/hn55T2PMACkAcJ6s1fFdVQeQXgrNj6QDJaHAXAtuHrrhLHh
5sp2gdjmjy+bNqoOvXkQyl79jpKJV5dZTLwNWn2aqlOAMEeA8ZjitapKteNt/5ua
UejGZIvfzis0T3Y+34ouHRkWzl3V/52QwueTvQc7plCEWyVVOMoJpP8bVz+CC3iQ
XpjEDXtIXLrpMjeTWJCx8l+SbdtZPfhsj+H6vC/wwGRlJtBIUkI500zDLyy570Ph
5jq28F3vvwRshj1MpNqR9h/1/ev22gqVOvzOdTaZG9MJ8L0HoAgsiYAa73Ql9+Fo
rb4TFxosm71Smq32KaDsnMFxXna+q7eRZK79AOI2di3Acorz7TlWOaKaBUs1SPgr
4SUubaSaZnYGTjtzcRhFomh5Qwy8XlAHnToVQTcpMLBzopwF9QjOmjfAhLhZUxas
htV8uA1c5BWZi4Ee+jD79e/H9rdWMR30X6fqSyMym2d7Oc5OD7sm+Om//NNMhCcA
Xf1qmQqbPIfX/tR3+zOiPAdozLzOpq/+auAju9r0wCHuvvFRh7Y7S2H0bbTUi78n
gPoTy8wlMNBfUPdqiaBfkm/K0THPg901XoATsjLeygyCIdF8WtaAw5G8dGoyUWYg
CUsPOXHFdqu2+4VS4pdjOsO57W9ElPhh+u4Z72MvCiWUyaqMzu3Ze9Rt+PkfiGuN
HQcLbjZNJ1RFfAlLmgDqPUpMvCxHyTQU1FnashmKyD0la9zdpKZutpJt9uwNpDVB
Ve/aDAEp+TFPMADKCzjdx3YZ9O+gYhztaIYtTI9YQslYBBVkMyJ+MKEogvwNgc9w
26Q/PGtEsg3OXoTmLFQYRXhchHbygjeKOgfreB2lEi6rdtm/ErW7XLDpEnvUDvc6
qcFXMlg0glmWuxdIy/3ytKKSdCJnMcmflmP/LDwr5qmaKbV2UyNpEjdGY89dWA1o
4M8cGQjc49DbB4RnaU0kSV+3PXRh4WYi8Wim9c8Xb+Ucb0Si87Yz9KnzHVFO+XoQ
InwCVH3YgpyMN3pePkIZS095IFk3SbVQXnRQgR1i67YBMqh4TlDzbv0X1Of9PT95
T44DppxBDpdGhAxsBEhr8O28h++ehvbMpxb+dZ2/rpBSQffPUMUf2CESQzxPHYiA
rD3+PWApmNw+6nSzQwNYSzK/FZYV72bmYh7NNqbJ8jf/NHvdD9AxD9jVdaEln9c+
685wYK8CbSkZVU4J+hF44C5Z5jJ3acD/feAmrKXLOw8qNEVpLKnXExTLrtyuLMMp
hdyatr5NZgIA+ZswS4l8B5Xbh4hR0Ixqjouqm5EL82JzFAT21QpjX7b1E/gjcQoy
BysD1nZ4JIhTxIQLYCYtB+GbCeOpLnoo/qD5AYvCt4PmAUeH49ozMwKDYwBwXAd1
aRIMcVvLNeHW7oPFOubgUjCJV8amoqohNoOepNrf0tpGSAKDlOZxynmekEhg8+89
wf36OxVCDnxdLopG9721A9YimFMSau0IUbxsAHUGsdFo1xB9dl3zhMWPMwF0ks2J
pDK6iu0rml2WA+oCdMh+YV/bPWUzTtQeIin/P8zJJbgPuETfmPZhnhTiC41YMZtP
fMIQ3Sn4lot1ojUZaKMaj0mXLrhkSsTmdDxp33Ym7PT493ODLzTEWQ1YEf7Jv7Mu
ZXxst2X6SpaBLInYkS2pMq0BhF83doSZjtZRIexqmXucjBVtwl35fA23Asn4h4rt
Q+FnYDrMMFQyzdDsNwtEskAn3wspSemXDIOpVZAS8XAxahvf6edljEJ1FBn+jPiF
HiPAD8DHUoBsASVCBAJ2DEWQbOINYC5uK0SqnqPsgwAaHqU9/74imWF6nrT+Azvx
s296cWfEN6qvfyP8XUt39fzoGvPsz03Z22XD0gjJxoIi/aJN1KcTyLvreeRjlgnH
YkdBtgMVVNMafxbXMS64xDaO/NCppN0Y97ilh3P025vF9Jx/cARSSTHUzoviZt/d
dQ/reo1b+uPSuTIKexwEv9oP0e4xuDYK/uolGeBNjv2oms1Q2Vm0PMj/AjNwMQSv
G5stVM50/YXa9909W6BgbBk5ZYnh/PRZawOd9v9UcE6GiUbd38qIBnsYKfGC/n+6
A9NHW8Hx7uzg9c11S1CdFkm/B6DjzTLl2yzbelbHw8pIBLm71YlQlYDoJ7CZ9Vkd
FDoLNUnnCyo1unpdUOKepA4Qv7NLRc1A09RegTHrJHTMXz9vQKXolcrVxBcMQYlI
+I8bCyYB0OXAHrPuQXw8SR2JEemPj3fFY+5uVwxFeI+w5b4KR/POa4cn5/unFhkV
rVKrPse8Tx9jDsjBT3LGt9DxlYVsbiOtVRvOAZ9khshvgo5j5CZ3yRD/w9i3fvkR
l5fzfXb7f/vcNaw74lI/kRPJ+MX62BghaLePzDJiQI3KPDWfUASk8OZcl4dbsYmN
NDT2Neeasda3utbMrs7SiyI0kBS/N7GQDupAufCMM7Z9fSyZMJm2N/AEQz1K0aZ1
0exiKJK5YNd6o5d8Y9BIoDD4/4d/hfc8kwgpSevz96mf8O5u+/IXCLpUVliL7sOS
rM2UgUySNctsmtSgbN3CwfGCquOz1T30X+MelbJz7ehsQqqrQJQhI1sZKm70AGFS
yF1nN5GJsbEVmVoIZWlGIUxebVNEXRbZBcbNgEXMlK9WuXll02BXCDfimVmVGUGD
5KObNM5x+vJersJ3QHMpedLOz41jdttcoOJYUvRddapMDwFcOR75B96fnLCskMcy
vnCwjybe0qCaQDFkAyzuZHITGcFjF4HunQFZqaLG67kxqoekqYy8AXd6Tsn+CSb7
uLJ7Qt7VCJnY1/txaBcA9Y65kDE6Lq2wLV9bz+LqB2mAvppXSr1VcOQYwOwnKZ+I
juO+sRbNpgIGrTDdGrCYQJU3lczKnzdJ1QiXBF9qKU9H/c4QlWMr18soSar5fSpB
fMTUuNF5/jKl3qBU/gUYH8Evhe1n3tl3h6d9oy5LGTLsiX4aqgva4050d3AXpE9T
O5EF+d+AA4FX2krpGc+jT1oLlkMI8SiLj2d0mm9JFuDHuY4CZLdtZyoVFy2kH6w0
mOhc9f38IJ/F0ZDt0xdaBy7OBut21/fjolHoJA1r2ILs1dYgR9s4B5F7oefKJUNh
GfkvxlbVyk7sr6H+WVqn2dbDtF3GF2lrKMtcg/5MGB17YrRPZReCtGhGTGdeLNf4
olG6NunjBeNFZhgEITFWqBa0zRbTh0uj/HB0l9qcdn710lghytxV8Vu6effN29eG
DTirmFCRKelEFKoDHy3piu//y2IzL31NF37XY05vqgLiA7yji7eOFo2t12kYirUs
ZhPx/tFfK8g8aHHhZI6NM+7+hxnC+bTuqGR6Fi/ErCHFdV83iSrJx61wgQfsmUgr
DMCjVElIJ8VNqhX7zms4pSYUAwxjStBSZNWf7pcbKSFevWaO31bRClNDYESHvcyk
ndTKgEsUWhx3WXQBpxzvw9WxHhszQ7tELPgKqIjP2zBBvM8zHE4wXENOmsxyYdL2
LXhr+Cog+uKjXdEhwH9ID5pvIYKRwVBBhORfCLZvZjg1T2PD9dxcFMKeMJEjSYs+
NVC4JovD6kt7A4ClfD7ieNfrQ6LNMBLLUKWIjM+itVLh7cpt4p08vZmAwafdqYl5
Ta66VbMmJ5TpY7hMizheymfgryaOMbflQC/PZ+8EVKXrBDLgH7IeZbHDemDqP1sK
3FacExJwoP5EuPhIi1PrgkDHelcagaN+1HhfcAIGz2uoPBnn0X9v9qKtXK7gEL0u
4EPdDrvdjAHZr8jkl5eGXOazGoTRImPs5TBd5fH/x3oKYJ6UFf846IFGo/r7Zt8h
AcEpvNR+JEn2rgVhy6ouNS4ronEE5uUiVrxmKc2WTdPuaN2V7JJsz6OmLTXfuxFX
+56W6tjnbfrCcrJGdML3xxjGvPchiG/fZJ48PXgAN91SI7iVY4FD88kgcwvGXg9B
LUClj2XXL1L3LMo4AIkK8hnUgV6KV8IVLeQeKJYmQDWcF04CExSDnPf7UaZAug9b
WNJdj8oBfEoCqewqqzknSwOBJuIJiLXXYYW7FCOiMJ6kuPgnhwvbYWY0WBkDoJkT
Kzja06UFi9wBam2bb0789IWeZgby/biqMbqtm5mksLK8WdqgZnNKMBYeB9JKaW5u
NveHbPOW7Hbkr/+uinZ8Fpt4HnjkYqPF9exN4Ja7UK+vLeq2SsCfqecJ0jFOSyv2
Xa2hIUD3DFD6PpC6Rkg5Wq4GKqCaGPTRH34noNziqMy1zTNLCmUd0u8kQCwgtKkP
fGnj787Xrb5IdIHqc5o+TuuSQd9ZSAkSQq/Z/t56XoMmGcVji7/i0ffIl6di7QhQ
CEr/OhVdyUZI2u2kDSxGWREDGaRPkR++7IgAXo9Vr6/jHAemD6Fb9G3uaoRdcjbW
cZaB0vr4e8AvcR0IMMpYiup+mrO28pSHhJHuvBtMvRbItMTTrCUZoEMt0xxR6Xje
LAASsjlTpXVJUF9+1yL/z6MoMSGsx9LwP+gqLSl2eioMMvap72dj9a9ujg+iiQJ+
a0YtX39K76exu15YjHKV3ZldG58mU7So/GEwahrI2FJRg5xhFsqDZtEp+D9rxg66
AoX8O5azlbhzL7Bn4HovHQEABMOWJ6fLbmJlyIhVfvhXyXj7OYv8hW4joOksBObr
YzgssOBMXw8tl4hv5jETA6cACJVetfWPHf1Z1WnuWwSY/sqGZXAQ0iaSgS3zzzwB
1NrJmNaQz5QPtXK1ZlmVuHIE3L1egH+/SWk71NiVpPVJSOO18kxNxZJwMPvl6FCm
uja5ppxaTcLRMRiH4dJvfIz4i75epol2QCRTi0F+qDUD5zf+iymc/MEA5alzE5QI
EGPjQsIOS91ZRASQNUUPkTM4vx77/5dXbJ5jIFFLd+yn/QymLODZmKBCOOxJj2+c
M8pbQmJkn6Tq6P7Wsels9yXm7zD0UgOs3mduMa2pm224BsnhUeXBc6Oh19uw3W1j
VaqsA28mpsbJmwxJOSjUPrW8Ky0arczgGFA/01g1g/4YGs5fgfhr1c6FjXWTcIfM
Z5aUwQvwz1NTm9F6p7MvS+3pQFt2EB5i741kVfSs83UTuqFleW4qrSc3ZBExaJ8N
BeTXq8pwBCb3wDUmQUHe/jr2eiYJVCPPUa5E1G9MV34YqRh/d7kE+LixvqHiWMqa
bVvrseI6WaQ6GI+HSTXN+Vf6zvFFSwMFdIxNl2utpvGjMBIkU1Hi9135duck148B
TfexfyRlH8eF92TSJkQLdW4kOOS4zC5KAsWM6CJ92XJC7C5ChE2sRyrKlz1bGkww
dz0J3qw1gVxzDEwhGyIsLyeSqBH8YOfEji709WvYNz49BrExyAWMrywkcseQE1o0
tHcR0+XtlB5NhKWitqHUy02IRI9dROVdGuqU2Gzy0sqVQu/r0uTDUC2273sdQw3b
v8KXpJKE0o3n1HmJV/FlQGplZj7hr6JGTVyAGxr78GIuod6s4F6pDuP1Zf1kzd4k
RSF+ZvM+qdH7K06aHEHQsKJCF3n2jQ8nN0SxHdNYlSvPcipYA5k3nM/WnT+b1Yxf
IPH9YhnfCNU1jf7aMgtBk+DINkLIDiwtXoDIporZBwXUaQ16SXWYtDF6ch7CJg+t
m6eA0WTUbTvA7+pE42PD5ParPLNgkyJgYmDM4UWuQsYwJJcZC/F5W1btPibExO7a
9Jy3WD8h8OSKkBkJRRDKBmeLuZamxokAsRyi1A1FXUw82pU1xciiTcHqdnlyQxoy
zsqrAEKsXjAf788GSDoY2L1s4H6LoSKf16HyrA2yw/Pbdw8d5u/12cFXDauqGMeP
ztkpOqKU04V3f0vAFlk9RiaXsiRpdyroaLEB232WEjm0/5PiqR7ysRoaDHP8jaSP
svtEesFnuU9WC6d6O+u+yj2TaWU3tIFYT/9a45W5CAbiSwFTXrM3tz6g/ZIfcaid
UQIm7HC0Ktgi1sfTy8ha8tbGRdhHg077hlGQSahPA4Dm+VNB02qgIemiPqDCLa7c
9tiAyNH5vBUWdCZK+qLLud3s112kYWQPPtWEyUO9J6q/YOZV8ZAbni2PA/Z/oZri
VSu4v4SjXwN+lTWZkan3ngiFkFSb0oselD9BZOwAA6mg2HN7wkSvdvQ4o6sSYG/R
vGcIhZsbGQoAo/eLZzgNw0gFHsXhcIQdichXm+75gsruQ9eF79CnCSk0E450BFmE
gxKrHMcCXp7uQ0ur0S6uBPZIQbhlWWZyHaij7zZ0tOhI3+c8rbQ1XE52J4iY88ag
g2UJQVLfXcNhpZxN6dwglyc/2NjDFBKmPf2cCK50TAzVZ3yC5QJ9t5rD25jlYA86
CHifr/ocWnC0vltCMbEIDv3zqy/k2htUUyDj3k14/wrqbox1OGbbtSR4ylNfc+Rv
N0gXa2un9BNEmH7j8jMBLfegLUOMGYmBILUWqRLj3mWN1+ZQnMBuKDM8ZdtYojbn
KEHGFDU3TW5t0A2oBQ4rNGD/LYjtoVh8Y6hnB+QwCB+TbKfBWlQMIQglrLrtvh7K
yPpydE5CxEAMhwW5tzDyc+pBFtk+9QQtvZw2mSJj29Af66n8r/DBl6drDq9OoHoA
DrLmPSEceGNLck/j0o3VXwC7qMzv6kpIE+hNuaVec8rPJG8WAg+2/PrEU7CLT8mq
7iI6N6HsO6RXWooFBcEZ6G24rnsfoUoKatFBrxFwXAXNvjN3QB+NHy4+LN2fPMsv
5sD2Dph3tT6txSfiLtpjnd+M1m0dtQF4YALmhgVmEvdzLkT4qvdWDuMhYkqFrKMz
lKJ02W+HvKU3CPIFG4Ds7vEJTaNkZvdzSr4pZh5HrmeUZSZyJW8/2GJ9c3J2WlCg
fVOOGV8kxZnOcSmwVzfhnm4hAs1+RIMsufuOqW+Ly+hPvJSUZ5dgjV9nQKAkr8cD
AZiI+02qF1XJLo7xFNu62AoJ/wNNXr5dwu0KPCc2STwYdRAL1rcZkNjTUPy9LbHa
IhHs7B712iU8/I1ITldukk52JyVIEoz3YIjPeCtw4t+eaekEIuZVRuvUNOX0Nf1A
6KPrAggmaF4nCWbB/BaXtUu/C3HF4M8tWwCpUUgxpofRNE8vkPM4zIsmO2wzUoc9
YzgxjoDHo974EGNDk31M/7FDNWtKJqMKCDQkt2EzzBpa4OFiAaCZBTAhS/XEMZPH
NQGKZeIvM/3PrEmukhjFntuOdMgLR6tKmco/4n4LIw7reMLMIvFG0UTjNId2i8fl
rYO4YEeMLZARiKk+4SCD3EGEEzIkST34azxwbhRgR4LYP9MDPxRKaZQ2rU139RPE
bg6sQFSzfKqadgK2imAZqHAF//LZQbWeqb3u/crXuKmgzpjeXb9OaAD/+65plaGt
gHq996gCw5QCSDhpJvLx2nE3P3MrVzgpReIvTBSDZXgMkPGi/FKG/Mrrt5NvVurb
+EmmnnbYPERPzBQwlVFMduGq5ywt/MSebthTYEZha/sa+qXNTowGwPDfxJmLOqvE
GS7lLAcOpWT5K9dQui9JINz8A6sJuZSTqSIA9quokcv29WcZTf0UPXAnnqcGnqND
JHY78ozD69Irm+/dbXAzso8bSeBGRxSI3Y6K/iuBtHeAANNCQoIlqfC8zTGYWFp6
44fEXPY+R3qefAe2C/fdCKkorTKj2GEnFLKdx13m83NSX1z0pTKrbB5p5TLhY8yV
WdQjN+Llw/On9YV9kM3kh3vFcaifCls/p8GTj7bZZ8Erq49wjqYDVU0NOKhbrBq8
SL2loC+NuS6XK4pqElqp4ug54IIbuKWMCSrGe1s/DGiPCsfRvvtHDTl8U4LcoO/v
9lR6V25SVRqN7pMjW7U357RrGqyOYwzFS3tRPdb8SkCKyGxU9N1vvW3BpFXNy/41
XYJdBvjEoQFA9LTOW1NXkJ0rowxMQPsFaoI0WSSbzPJAiGa5nptX0BLzODO84x58
tKQlXCdQPNfOY18T3b9SowD4iL323+DZHad62OT3JKJYl4ihw1/wm4KgnuCh/XGi
jwWbNDVWYlPuXSvI+JTbujD1ZU8pRCUEZotDb+3miI+cunbfODBIfZujg/nWWgsj
4bTw24kIipR0LmcC16LcuCO8LVnkf5RSO9xQ9ZOvgQL7zPl40riA7uqgyq7on8y9
tapvzc3E0KDkINy8TYs6zDmiA8A+GzSY0+IFdRO/s0qal4TlQA+cfpe2TNfrDLv2
62ySdxrfjSk45N5uz2a5TsAmaz7Zu1WDPG7Nd9dUhOaZn0994uN1ISWH4877G5yx
f0slOrteUVSSiTekSAlzRNmLdDfnp1RQUmnwu4DUrg9zjD5jMvD7k/b8/43Gx1vH
8VqDPAiPAcaS7tY9W+8swhuwtEkYogb5xtREQuhdXsLII0xfcO+ug49TXgqVjSzE
O9iYkRjn7zsSDRj/hZ6ScvML7EB/ltRDVymY0x9dXXMuxBuCx1eHNbqLWYObld90
+mI2keclZ3mavDxqQ19Co9rIQOLsNTxyVjfO1+wwicFcbChZMhbtUHDtRD0hYNzY
fB3qsq4sj3+oljbawb5UGBbQBz8E/LTq1T9bsExJaKhxNKENFkPk008Q9Kr6n4HE
0bUUDfJvvpcIoSzb461Wg99+Unsh8nYTCfFqFrIe6H2DKMwcYrnuubG8yKDUdex1
XkMvbeugUv8EmlQZk/xUaWVG3xUen5CaufnQcNOn5E5cDQdpF85ewcMGIA8bp2So
WXERDtbrtLp78eloNh/Q2/HYAsCWh3IRIaUMd+dHu5Bc0+ublQDxivIdub8PJfIG
vfHm0jyro50ty5ZCaoOcNoajNokkThMboABHKgKMuxtZYtIjSxMgjiwGHyDSGUZK
qF3/IgdxFhKms+Jkf69ACKk6x5CMoJCCZ0QiEfZLqwIpa7kwKfyk/wrOGpUE7IRb
geRPGNnYJEYJULytO663nEtQBfunHvAsUCBQdZ8gnd+zdMijjUqFFuXnwKcOG8Ph
HfzHP5ys8QBTKmQpzvmooWxzoOANMHd+YF3nL+HVeJeE6TUSUhSpr+R9u8wq/7yK
1Tw3qjI5QE8MUs65fC4+/GAXOKOzk5/Yi0oosmCdHb/vyP/Q8gxFiwCDZTEbN/MY
7fTO8Cw7EW5KHHPC7oCC5J5WkdE/ZbY/bNmptyUGSqhAmwINyHng3k8E3KiSBdD0
tj3GTd4TpIvGO/5ahw1u8Yz8ed1hflvhqDW+XFsicCFb8F8NMKgIZE1iVH1XWULY
Q3glBF2g5Ndjb8ltseCiVwJxR5ri014vU9QcxZtU7Iuzn7aXI5l6evfqckZvoy/e
kmOIepfDC2gyP4es1sUuFapPBES7/3Ui3LbViMWhVemY5SWYAjLNSdbTkBaTUD4k
jMCoyjhUHCDSo7Q5m9IPJ1jbWmyMxyyiunYzzDTM1gwpdV+kZZneDMMZKWegiC7z
hgbCJVtbHeasYIi3lBPmgGoaBQwUhGgZga7SSx+dBhaQio8+rXoJze5oC8ifjozZ
hFfKlU3xbmFUQlCr3AIHKG5HPnztdCZ20PakQ3T/eIAFIf6KObINnRGmBFAW5KLA
LTgq/g/jU6MTtBVBVtPcdFeYRLYTMoxaRd2yzhU9zfSRpQVJfivX+bgP83BiFTB5
BWID5imZht56UWoF738SSb8gOmqZk1J35m1KQaoRsmn+HTa6OlUAAkA1sYIynOHW
z4b9/QovwrtdlTJ8Ot1lYR68Grh/Vjfd2KCDMcFce35NR718O8LvfQ2GAnQMncc1
8/m/TqXJnHOmd7fsan+RUG+ba4JdfyVcmDDU5ftTSAymO6CFer+rZYFBGLedb6ke
jQqxHGKdWWWuSEbRjGsgFvcVL81IYMVzT5nzisGBn4IXztzIBJUVC5+zwex2OSxu
S1SSCiY/BkcggOXwESHBqhYamvTu7ZudzDyVGLCYSJHqqm/xvFGjDRrm8ooVfA4w
V3vYuPWZ9it/b5p1scAQZOcSpTfDOh48OQHTY06ehAEUASVQa3nSlP8YgLfVby52
VIRU8b4NkXy+7JZHiTJGs/SGk+sDxmCts2VPJkpcVm1PMtNJghHNP1zoXI7kkzVA
pnMwpRzMVYtNhGdSiL5y4dOks4ahXtHj1IZV21OEfDN7Q8lAGF2M2A//U2MYkO7E
pHEzriLn2sHOx+s/p9CYtUTwU4LlPxwluFfDwsdRqVKGzu3lhznAiaWHI985+m3V
03G3xOwlDbcbUUsM0ODi5DXE8/jF7QF9r7GE9w10SqxFdxf2opIcQjRi2gdYXEtE
CpJSn19Ql8Bt5cNfIlsbMIumicaAoTtbNB3ykd+EXXWnlxWtApWch430ECyVqfCz
PH9qIiRQfF4WqXcxVxigZ4YEDVvq8hOcejdfc3OuTB3vgZ/6WlmqJSH+NIy6FKuV
hBXeaOFQUUXnh0mQXe1lQME0Yk6IQ3i+LhcBMtZ8Q/cqZzo7ctBtQIKoENn+kz4H
/xp2Dyf21wgVlcCd/w0iI0U+1jFI396YxSISXwbSbeQvTFA06B+i/QEny0JcsPAH
l7UaHbAehOsRbtsm1n3Wa4zzZpZ0s6qTFtDQZd4cJUoB0Oggoxg/BmzdkzG6ErqT
ijKgnN3t87cmPlLZTVynnDtZ8oaILgGi2TUM9OfmwKkZh7L+nDlP4Rsv0vhydW6p
zaaXRNNbAfirnW2gcQcq0RS+nhmtZrMb3TEjMZCy6x7R3+I0S4VrPEj1ooQfo/D3
5EDcFFJbcw8a/U/zNWgWxCtYM8NBX33oo0zNqB8OXNa3M9U1HcWRte5dyPSjtuhq
Dcp59l//RpcZw/mdO3oR2J9Jwcu/XeBPqWA9slST7RbR7UkM+jy5ZiFtKTKBVK4a
/jjYvc1jAOp2nxuy/99CWP7UpQqmy03h5tl3HhcPid6FZCmmsOdbawor/PqhdzDM
WyhBVDD1WNNaFw5pqSph/DjNK76iIZ9YM4LkzNfcml+83ZrAq2yPWj7RfUoLZSj8
rNzO8ru7OT1Vnpo+PqsBnH8M14jzcKhy3wLt5DfeI6RYFCCITHdttVclwsooCvDy
tp9jj99sB/yZWW0kNB2Bkki5ureGWmzytY+cfWofXw+Vyh59tzwJQI/6vjLWKlC2
ZHXAYNHYC4uNovbamVtUKGTYllpL5YE9pfg9YSU9r2s46MX5cBiG5kPPkssWKUb4
pvEW47DBVP1/7RUn0/1x/scS7qrJ4Fllkl6oJNTSPRzr/U2w5EZvcse9Y+N5gThx
k5JJvzDrEk2by7MWDqg6PZQ512P555dxB0RWS11HSDv3aZwPM0vm+Q5nMMVFEWWR
JCItm/fratbLs+ZhvkmLD7a9zc5THzisBVJ74OKWGbCBGlh17XNrvQAU1P1Cs3V1
BvQUeZX1FyIhBOP9GJ57pVV8TMsdNE91onli4q9spshORZtANfMZdTqsCFMrMy2d
n/map2xpbTJ5+Y9T5FuIJ1VuMg9GONKuvkSlDVApYVph+6vTy6QkzK+QbxjR82wH
YVRfK1/i/fUEyRv+dIkvuRLWICDmTy2pQ1BnuZ3C+iRYLouJ250afGDOmLh53FVS
gNk41b1HlfuWBbyLHYdv0Ubg2qZUxuNN/5s/L1wPii4iRnwZ7eaLhd86TBikvgUe
68paYyN1Q7SE+9EtyeoZNbrpp0e4s70PqOjc6OFew2YEdaJYrEAKaqYTfc3yaz2/
L+6VxbaIPPkANZ3D25RgyBjyu9os14CV+o5hBbk4uf/ShQlVCxKOWKJXZSeBJE+m
lhWiSLjr19d2sLrndp4/2VoPC93JhxRnD3PMQ8YLN/JN8f3AeVjY/NUlCRzcjJX+
05M5BKmPZdEczszlS72Cxqs1hA3vOqLTA47eD1GCPompRZ+5M8sv1rokyurjAEfq
dwl9tNDFytT51oCs49dqaHgFFpG8RS8wRQGBP57Une48lJmIrlf5rg4bbeTwImcF
2mC3wyEeED2O4s5hFblAyH5esnIUa1YP07C+kcy9Nua7bVD0erQHoE8oZB7ItM4+
Z898Hv5BIWtpJJzpZxiFu0yLFXqjPdptJjpZF9zBUUrKLzf4u1H4zhSigLq+uv8h
ItEx7nKrAw9V5P1ktmxV+wetzkT6OVE4JFcWhE8FqqPBp1lA5uY0HJKHgF/mzUw9
gS5Kw4Q20Y2qIy+iL8va6SWzOjfjdf4+Cq1emNuTGZOryvkUyGE4pVTK3HFtubpA
Zvujqzz9FhganTziIVHi3G55NQ9wf+oeH7LGp7FlZxRlro5hxVPugrpNUxz60qOG
UotZ+xck7phITqwP+fWcfIgMumQcwJqbCXG+0FwgLNy+NxWME5xBpPH7fsXRVmNK
Vx7n+qjeVpZN8I6INNo+OOi+pPZ3fvlEdIE1AT2B5HP25CB0V2iEYd90JcBSltrE
xmHULd6EHoi/KbYZS/waGHZQlmgE+GRm4/3ejVJEXE9EP8+rL3WsenytBsU5yFxf
a1e0Lw7mCjhk7prPEdB44cKRKgwBWh1igcIosRqlFMuF4G2FPV3tGUM1kXddDwnk
455edQQoTwiabqCBGHpGD4VnMT5M2b2hIr2197rslIFe6ptxb4JsPsX3mmj2oZk6
Eo0RCFgZQvxARAJ3tx7P1wgayzQQ3url7TrbBa4l8Ga6NmCRphe2a8Ac/pUeJDaj
qbKMSdRdKM7viWd6NSJCTUwfcyK5kk2BBefSf9ujmKEmvpqmXrP3z+H9DNLJr+mJ
YMPAvaoUzp9of2AvXVi5jw3keAxxzSAtH+yHxzXOn+ZNWYf7sM9tUHp0x94sW0MG
YmZmrk8Ise4zm3K3h/l8EEmEEvfs7gy4Sc+IlAy45I04G8Fe4C8CdR5xAnZXnO1j
8VWlNNbgUU0WJ19behePxGZWPg5eP6sp4PR3wxx09ML4RMPwErpyP9d+x2W2xRKa
6XpiBNgaGDEdxzWvTjTTzkOIM6KbireerQ1+04IbJnG6vI7zMw3k3SjHh+iWihAB
7030gmpz5WLru5WZY+/gRaofQMkVQYfKI6PJ2WVgtxs7rpBGnAu2Ljrobc9pduQ2
SDtLkvIYI4wG6uWGcQWCbyPqGeBfYIhZV7sHAlCktjaKHViPHyKkCMvw5RBfIp2L
Srhi4Vx/aWM2MaTjtNH9N4NpgqYuILXC0iwmK4GNXQg8L+F9bEsficSDavkJ7f4G
FrwT1xT57quGa9e7vDwQ/miI2zoaWfLn7mlX3EcftPN09+z/j1h2IEoQHb9Zr7+C
f6r8AESvDzCnjC4yXAfDlFCuIo9viQM+m9X/XfGGMBpj2j7eBFAmyB9gLxTb8S7O
myMx7yC/x143OJaZrG/eGWKQmTS+xjTMNp54v+mXzvRk9vRq6uI/dhzvP+NNSAZL
6B4nKW6QMg6m/CONQJ2gn44wmpgC9Q7gJwURpq7GPGnx6ltrhNeUmhDcXNSpqkAi
SJ4YV37eEB8pBvN/00dknKqk/S5pn32dZVSIi2ZOAA87La3FSRf7rRoTgotxmMS7
dmNHCidFp8N7B1EGPIvatQ0AsoOCEEgqi1wWRn87lHahCP+yweiq4IrdCUzvSaeV
5sVou/1ONC9eGcoJ8upunk+oVQHaA+I/piMJEsZKFZmudplWw/KQKwAHQ6pYD/Sh
+gryZASHj7HVH6lW/qVz1mPlgn5xd+2qNox3Nvi9ut7u+nx9ZFLpYS9a7ZaO/JIM
6uydnLNYthnqlFtexslVVZN5u/wH3pwr83eoqLk4STbRITfF2X/VtPqJ+Vca08f+
fLkyZLqzd6C0PWJA9fyEMw8oiUW/dbnhroGDVrIn1pQm+sibg2offRHuzUFPBqpD
U8oxA4BvoZd1J+O69zsEbT2k8RwJB6DWCHcSkJ6gvwOr4aF/GIpiBoBy2icuFteC
XltvBVarV2aeYGQlbnogcQ/M2TFBbFMIo/Cb2r4gEVEpDrONGbNKsrMiXH2vfGNN
pnorpS36vkbFlSDCihhG9J8ZjiZrLbyBMMTL44Z7JGmLYkBotTClqd0rkBlGfc0O
dECagg+LKygRinSE7tKzgzWj+dtqjoEKr1SrCjOLjfKYTYO8OUeMVp3eQehXUzeT
ysPIah6ci0MY2MUDPsyZt6e393VtO122VupbHvSn11PNqQc8c49mFfD4hCJBiVag
/hnbsDpTYq185p7NFlS/NejIsIyWhMWHLdlJQeoNwQ/4xOg5M2kXjAhieGJWNepZ
e98iBtF6fzbrrouxMffNuwRX9bIE/Bh37sYHUBOaYIbHAHQXx3QCiM81YhNf+Zcf
VAqnDMaxK4iIQozZyTfNni44lF/4q9/KcHvPANZNuJVRbk67hI1vJ8uhcJpayk8L
MZzBeiR2DtEJm4coYIltXINeuAklua5FQ7XmBTYtJsJsAEYpUEGswsiJETO8i5EF
0jcymwR08XwmfASrXvmOWPpzFwtqSoAPVWfW2mTunsxXiY3UtEPqQHNrakN7sCag
W+37I5VhjsyEtuptFHIQXcwGaRDInpIorB6OnRD8dIG7U30TiLaQ6cvSJ/dB7gNk
VM9jMKFEG8zCZnCd5gYrDx1SGtrrzAusCc0wlLgVG/3oBeMP5XBeyyeZOgc9oc+d
DKcwCw5H36+V20JqwOYijDJ1W2vzI7d105Xl7VAKd8zipXpC7iidRf1hwxqdP14k
sLTMAJ1H2RVrbK3OaWy0HlX0c3DnDN1xIpCGzgWkuP9u2GBSxf++FyqxTqAeeM8q
bgNgd6C1IVreoU5uY8ymwcJebPFP3t927jsl/FjRE/FhmTiswJOZTyb9DILY2WsD
PnYSG5hmxaaKvdiev3s8jEBbkgqa5jODitYlfrDk93uJmqWlbJ3FwXPhNO9UdhEQ
CTpxFW1wiIuPSx6w3mL3xTfQFcI8/xD7yFH+z8hjaWbQD/ThSK5MGmGR1ceOuaGC
7f4hAzLqJqxDgcBUiJxn6pcFmfkGVRtkBgnr3RusdAg/EWmNAO1nei5Dku754yZs
UGmi94oiYbMcZiFHy4sUA9v8TLfsQxmi0wHsWp050/VUj+6RDBHucWp8uDFqAziJ
VONynNTLdZFsR1NkUm9DClso8vpQmOqU/PsvIXMgBNV1mbT8h1Rl9novzgAR7ela
P2x4Y9oQdLGXD0tTpOasoHpEwdxpvpoYCB11c1Hb8TeV32zjYze41zDuJJnaxnob
CTDxQVfX83dQZspby/a34vZPiH85GueaMoe1syAjmRya7JVyHU/wIOncQqOx36Yk
PhtElnMxUzBcdT8iTqFZmivC9ND218EPuEbqfLAbOnFtORfqXE3cPYZSnD7ieVAb
mf5pJpQrHquPcc0Krg8FkKdDBnpyqg5jR6Lcx8HhFDsFb0FFoAYy8CYaRGWCj3tF
V7hgxZR9sr/YB41ek6MjgE8fo6uAgDq2XRazNUvvZYY0sR25RdjJIF7GaCxzWRFZ
IbOy5PT4RNwZMFrwRQZEEsL3WoD8l3PM4f9+XbaoHXPVi01CSnvuY6M/DZup1y1i
Nmmz7f3LKdah/gNWNLDtbnZ/j4dmetb+gdme5H04KS1Fis0jINY05NcwXo5kF6Od
XUTn0G1YdLS7y3pSYnturNwoEEpZBaUFMCKc1FmhZo23Od+SnjBShDDSXxMItjCk
KgE2ew8uX3tS/HbFd6akZdRi1lobpKaIbjtH/KWjYBfRWCbBP28XJAjDSqWJWOtD
B7umwHebBD/YahYIzA9U3zS+xOfaxeu0/o87Xob+ST3vbBbEZzRcy8aFzJwPbMwA
lzODyKNG7im9E1I0/3g4Wk4xPHPT40hWQSHW9pWR+7HEGq/1m0dubudUE/P6P3DE
FvDzI9qQWaNG+PUYtp9egjWusPm6RbuwjeNt3XvSZ7JDQqOytoqpAA7cSPotHWGa
lHzE/1u58OJJCvfMSmPjpxck9GQO1uZW/7rS2jYzOIMYa5gDoGy8UeszGFYYYQYv
B+QcLZX0j1p5/DBMzn4hIbbE6EDLTX53YYQRb+u7l8IR7rpyADhbnw0unY0t2PVH
LIz3ENYo/08bLUho5bW0WeXLQ60U6WCYk9xzTTwJdAZqNqtDnHhWBKpS7BRuODX9
yAGLRPH3Umq3HA18rZR2mf4mWNwsxcntqbubxSHgKW5tPddGH4Av2FUGIRFNRchU
83gys3bVrAShLQI9KSIJ0vRPVQJ+ZHHKfEDUjoDVCbg8GGaRMEiOCo5jHTNNHG1n
wPjx9xj/3fLBVlI0BTGGT2NfWIvuAg3uAA4rSA2fV+5o92/uaROC10MbsdKCBn9o
yytwOcj2VmJxnIzXwRwifGxBklALFrv5wibpNxXte1rP8Do4kmcQHxF5cmCYUFRe
B2MJtnUPPkVao96a0MbgKU+ENvtBT2TU0VtwbUzVUzsygth07VPDKi0BalPv7Axr
orWslGt8EboXhVJCWWDlat3gT3u0wtAuA5duwcj0AxmQ+nrqnP8xeBvzbi1a8Lg5
qFl89CJoMwh/zayeQ4BvTccHMRHiMN97ayKkA4MPRnnmeKJeR0qJrOFQhuBg9huM
UPqLSirWFrn9jn9LDByCOF/4w4K8Ag/1Gqe0dRkXMvK/V3dbcTaO+Y/vtfzR2K0p
hFIh4Oa74Nrm4TX1kvSIHWLTfuSj/A+UBsF/F2VpX30t4MPYBhNYLbLUm8OULRBr
azD+s3B1kSsvniRrrpWnl0hvy97bTpdZBQQPHRB05bqTEfQlrBVaFyT5oWrb98ui
m/VJuhopFQ9qmMOG4ZYnzCrmhvxqCUZedfI/E/5DhvWH0pqZJ3PGMlxThBzCD4Xp
0KTbXlcITmaHJaXrHQJLQ4FcjI/JzNuPS4eKZf6iwOFE6tX4XGHvbF75iaT7H72G
CCRPPTTPLi7a7q9/HXHVn+90r1DGgg69t4lMP2DaTaBp+649NYjPsdpmHwcg2VgR
loS7Z2qqunfQ6s2/ubYPp8WHavXIJaTzKs3RmRmqwhGDgm6S4D5pzvye3aqXYzc9
d9kDQsvvFhpYme/Ipin5zkoVQA5kQhWI7mepleplOsLn8oMRNV8FO5e/qkrR3i02
CF+w3cFJqAF/2phGu64GerTuEJc+BwKY3bRroEjHQdUXsiGceUxHSJ3Z9myXyry+
YeM3Hn75qmvKbNcj5pI4Fa1DZHf81N4qYmeoHvYyuFXWMtCdDA9XP/bzRA4CcBrH
7/UgUGrhnTHOMXD8Rm/XIpVsZmuyHxYGHagLpWzzDhN+Q2VFZizHPJ1EfNRNb/Iq
8wmsTRWEgS/A1dY5q17Fyo1fIrC8KqvMWkz5Ny7CyYDU0VOw4sAYxxV8dMO2CVl3
5t6iIs8VhzjuO2SRXYJJQ2SkEd1dG5j5ha64hqoJm6TX5kJhvExzM9xtN+v1HEBK
zPfqVZ0ozow447j50xsXg+DyKgD9ooJ0+M990iJdj+v2e2A+/NQQWu1e11xaraNY
oCSUJfrsZBPbn75h5QNG5ZpH5yuFi+8DrLjIrLhj0+uYTPTCVDz5UpmJxER0hEyF
Ggb3Xz7gxEgLgMlfAnRsJ0sE9MvVjXsFYJbz2XQugT6Mbd0z1/aKmK7sGkSeX59c
OFvmyuUz3F3FsfzNi+GweNN3rgFOfkE2Cl1r/prZcN/g6K8JOeRcsUzWUC2h0ddI
LknZKB68xifl9O57ihTXWRdvYNvMOYtpSwjo6C0P9IguTQcIn2+z6KEkDTuiB71T
dT1itdJTvti1pVAWohq6htPyrdGeu52WTFzOmJjnYLUiSUUOuw51BkjWPUGh7bdU
WAXaQY2fuQalqbuykGz4lGpt/WfrRdUjRJx31BSXvEN+97uQKeWHoQngrURDsI33
+bu1qLhf5UysM/nhXKWSPuBbosBnnK1S8b91LqnKPTSALkGqNXsOQAZb9yjJHe/4
IG/J0fdgz8kOWlU2IX/E9reR5T3B0o3guKJqmWMsbnz86fuKlHBRzRp8TRqk4y8M
oT+Po6g0RiyNIQ4GDhC11fhm9gkK+3TWpPuj1jGiPau2EEpi8XM3tteS5P5ckpna
KoSH8BI0oeSwrqUNNPItSDDL41pMPQC+DqPkSDr2uBgGlolPDwtyFiQCw74Ti9z2
FLmlBn1ta0bFLrB5d/AmNdkvx/c8+sX4RrpvRCHb7i8xog+JEVKXlHaWlnEWHIy8
EfNFrL3NNRWEXX6AmpKdqXLo6rtbmzmemUK2+c4Rnli3bbigsWB+ubWp9sqgH+Ta
Hb3RKHbZtt0KoM2395oEjQxDnMQfr+F5OXSzkayy1MN85FTjv3Qtq4EweoOtNIjn
53+FFZKndffkQhbG7O3IS3pvrrKzJnOWRNDsmu94h5hmtUnZUZHRrmHgUQvJkIWJ
1ZotPTogUAmt0pWsWgoL9f3/AM2TKhju6vSf1Su4Awx6NTUMj2wKXkSSIwfnhf8k
sSGng7TlIFSudTOajWWK5fOeDkKPhqM+zpjMgPHbwQ7zwaxrbs3GkFNvziEEmcsi
4sjuEHLxcIy54oZq09I2UXYUpasFWRJexkGeJJPq2uiYs3QMdjXhJANFlsPM/JwA
JynsMMIL26OoA18f1wrbAfOHM/hOvVbd7RYrvlrT7AXKVt6l2fD9ByLD7n5e5Hb7
Bqe4hfpwaxCE3EU4K0nCA2EV/DVRDWK/jPnpU+nakY3WErRSLI68hosrtpZxgNKH
frFEN+xz4MPf1O40DnvliOL5gvyXpz4fQnRTqczaCNR1Skmn/euvRPxjDBlYho93
8ze2TjD45kcXG/+bJUJIIeSkj02JfKXr0wjvtjP978vA8HJWo0ET4Ty3ZZYWe4Av
+JZFw1/h99qRFTFpr02TO4z9IDre1n05y8KL6LLj4YbVOnPEfnyZjJ5sfNX5x/ye
GZOEMy4EnvvwmP63yqG7bEAZqvYTKxSuiAfLftiebS5ZtRkK83cpLQ3IlFNClkP/
ZbwslXwnSsLrK509DelLDDgfVBNYYJccbklzh0/JgiCQUTqIUBeIVRkLADBrniHd
t9N8FwSZKM3QM1ZELgqDnDqf0+MTrJaubkdxlviT98DbffRXSnFs5FbUMGdfjQYE
ncewCwr9sSGApPdMqCfw81zrhu5AA1cWubGlkIkeGi1hYexMiz+MI7v2EDO5FYeh
R2/o9qfMslZSRPXjoau4nMyKSI1mX8RWffMQ0/tMZZYijU6GTXE5FZNo4ZiXjKjD
O3nGqVoQr+sHLd478q3Bk94WpaSGOrgjc41dPk513QJGY7XTmM57hGVyT1os6B9M
qLdnH/y9PlvolinojOyDfV0WdyDKa1UZidaLJbiPbGetIr7j9/SCx8vwseEfhADy
Z6Vd+mF6J1VM2FcPSMLv0OQ3g4hoUlLKAW31H7fec7Fk5e+oC0o3sf3koMgEpLQS
+xaML60nWCXFA1n154XOoq7RbT8jwjPl4sJbWHIX2ycg1jGY4gwfMDQLV1fifpPP
X4PgGf7X5uwMLPz4gk+NxcGkEoaF5FwiQ7y9NTI8Kt/h1PZK2kNU6eV5woQuR3hA
f12ZTXLgZ0HIFMxEVITLfzFp+UfKG79GZgF7CJADTN63KCaeKc/3LRoju1EO92Ds
A8I0RoNmYfjiBDpIDcWOERtX7KMTzF/GidqZqoXktii8zU4izLA1YLFRqbnF2JaZ
5pdVwN9tAi2Onjq9xDLKGiFfJ0FtKhy3l4nk6tLbt1FJ/rfeMa9nl6Vn4amsnwCK
bJBS/pcH4RzihLCxhMAnUTqjH75c2a+AgZAh1dfsTeSDuM3Y1+tjG45N53P56KMz
ptN1l6T/76RqG+Cl7dBm1KT28U6F3DQojl2GsHUVfFCYGLfGcQx57+HB+v2ShGvF
Owk0E82N2u5PgJ31xoDM7K5N6a2yDh/6eLaEPt38G0a+D0U2QJhMbS4+1i3jwC9Y
4sMWTTkV60Pik1g88NVjfyC7465MCz72cbj8uzF3KRL37uyRolLZAws9VNdPVOQH
ZEb24Ph2UqbQBFJN9CM+SiNi2l6MKP5+ngFTnYSKQlxtz7ZcSY+wAcWBCiFeHEtK
ep0ZG1bhu3ZVVYkwV8kg9E29ZWivY0uHFcycmca4h4VHtir0LPHsOSIZDXQE60Tv
+onGBdnBKARPIs1jqcSAu0YN06oGxqDVWdM4MLHMsxXa74noiVDd7lax/ofVxeuP
1tHAzowpHE2kw/XBTdU8/WllRtOablCCLttaavxprLANptBYtm+8GWOR11S/4iUz
xPwt71cIV18ah9+yHTFuoQJV2wOj0CLJtwU5WVxVh4g9hASIO9BxVWqXHXxyBNZj
yYwBY5DSQbxhwatXoJHfsipuoA3aMmPCyOF3m133V9EJKlG0DkgJ2CRTKhFL/xIW
+oVKyEwWEel7i5ACW1Qxvw+oj/wI4NNGLXRw9RTa5D8yiY2AnMXxdRj/7Lzjm/Yn
dhol+sMyy46RjktvGJp0gK6h7CBNGMu2bqZQv4Mf1m8Wi8jyrOMVR2MWTDW8PwBR
tmTSgc0IBJgWHw6UplG7TWIqVykIUDC/9xOXQoVSVy/mjWM3vKkkUdgDb5R1eLKG
5Qcoz+Yz6HT25g3uqGu20jHWBlnNG1nO5oNnSx2WzKFSq8nmvH0PuhaPZBU/dRKT
J1K02qcy9xMA+x7iPjYxQqKOhRYlbx5h6R5lIelrj+uIOyPVmhKJLyJ5yWxCjmF+
mnpvHpX9fOP5L09LxO74QEQskpohPEIzORP4o4pXAWLL+UU1ckhHhUySdfkOsPta
tfVvrxkc9abh+gXYlSNogIV+autyf9XUjJwFJEjGxZscXZR+ALi00uRFNiD758Gt
vUpZNbr17r3FzW4QdMDz+Jm1xtUVLWPSPGLd2kEZwhCyy5Edigz3Spk28NYFsTSC
O04nk0t7SpL937DpLidZfJSc+YUio8Qnxi79XdY0W5vHuIwUEDoEqf35Xz7EdfTo
bj7agHLtuMSJZxp6NCcEK0hX8vWVQg9zZiCdRKdL9o2NeAoVqimVfxeu1uywPBo0
JyzlbDHZ5aeK3FS56WHC8Kz9gW0LIKb3SvQRXMsVzT3GSC7DNe5t91AAywAzMEkP
uh1UrzKucfhsvgd2mwhnL3oT6B+69l8pDeSSKZkxFItLIXQu4AJLEweinEaP1ZGC
IFm2bWk/nnBYcpMTsCBmpoarHAfPwkAecRJ1DvZRir6XDPsv0/kDmXFwNtLKLrcx
oo1waTpn8fko3gd6Ebgj8Gx8tvsOtDVC0NEWJHZPXGg6IBGKTvLD/VjgawGNrnkN
vaXKzHVuZrtipHCE6EgK46ko/rkYqVp8Sbmr1FzD+gCi6KaCr7L13BbLes7LcyuS
o6uLoFLS8iq/JZ2/DIcUo8zZZ7f/k3EFuKYl3H5bJwsg1KlueKLytVlXJHXlle9F
9bdKyC8LkyAax6xtDDpaa+p2NAjdQ+N08pVGKjSzChQWpDHa++SkDHSuIg/w/LQs
ERixAXXpVQf8iqEsUJQHyDNE8Tsio0+3bP5+BoolsIvLIeZ4UiCcNqtFhdxSLkES
bFSHHXCSnTtBDjJ4QrNu1X1rinQnRZ4kADiandWpYnOm3CqWUzRLqj+lx+WEhcxB
OifddPkgHWe+9D6u65DRz/c96WntaUNIsaJq6h5S5Alx9ob8BT5piCSR1HpNSql6
iy1pMZDIF/jbnk77plMkz5Vsc8RJXRgmaZsjOp4XYxeUos9jYrLn6e1TvthRI/Yb
C+11uoH3fXa1xjN4ULDYs1f2o6OjLjAyqqHBK/k/QAe3+t72ET2m4HtkktwJXHFD
xBvl7Xqt1p6U19vuzbkCjGCcm1mVkOMxwBlB2i+5ty6e1bqjPyxDeGjKOSpahHuq
oJmGNpfJqCWor8gQXK7BX1qY9Zoe7n87O5SMebpSQcsoHwZcuaxfUCc1ik36avIm
jq9V1HqiX8RKkc+XrHD3Ju8Wt5YbtFhmmRKuBOnaWmRFB3HcwlGHos3igrBHRiDj
4yxvUCCBqnkUImj6zhJQ2tjelb2exw2JUsnxvph1iMK6DXlOITaa0jDVA6JSFgXe
4tFZ6SLE5Cum/9bPqdlnP+oufX5byuWxuhSXUf7xtnZXFD7AFZaY2DYp1EJGkIIC
fBm3Hc20xNWXS81sjFiA6Mng80LagvBct1O8frLWQe4oRNkalJ1uxfoleNg9E9eV
YbBJtIo9C8cXzdTchYW9hTViungrrs9AV+Oj07boK561AgLbMysdZH7HYiKq54Bm
FoTTdb2abSZ0smO3ONFttYCU7h17s4jHgbJp2d7v6oEEv39y0ScNGnwQoAG2DNVQ
llkIobRMRt8pn57Q4NL7AwD4Kg562afFcUUF8kpBydTp4B+VDKseBLMDyH9frS6j
+1vVg2iRXbFgzT9FgziNF9NnIANOwJJPFTxsgkVpwBQc6gU/a+4PMIWhELJEOXF4
mBWKNY2BWFA3FK0Ez811gFaHLYQMsNIbxoxHEdt2e0pZg5ifC3n0Xt9IU1tGgq3o
nLShiHbKcVJwQ9qyQgXbcMy3wkU7rWpghnO6w1nDGZ0eK30UE3s5GC0/1YVH01A3
jeYN4X9pImspj1hGOzYpzKZzkzDNPjhNM0UHNlmgyh95CdtXa6qsckuaP56wERiA
sOMylOEh8cvbvNpshhmfhk22mWCyOLBSqcc/admoHx3T4loCRILe6YliJFvXPFjS
WUKF5PXkZIY3SQcnx/onkB2pRGD5WHsdI98W/GAF8Fil1J8qzMXe4y24tusnGiu9
lhV+ad7BnWxzg8qB+j6zQ/ooYfLrLbgVvpExIBef0fmoFFj1tYnWmgZVKrDRY+RC
LvhVnGI8Pkks2zymw3u3OqxIuLhxnT+nATTQOmlxVmDg1f70L3Rmwg6MLbXMIu+c
/SBsSDmKTAiSZ/fW9PqfSuH9pNysxxpkL7KBOwoTnJSR4tLOdtcBsA2Td2y6GxfA
AzVDyRSuU/V+HPUo7EP/bWEZ4/GsK3nvrR82dFn6AMr2GscgFTAEm32CSzv459Hz
igGmDZkWs0G0iXMsDd5NHY1521GGTAvkvC+Mn0mCLCAJ44PeJZ7zhKQ2r8jlCtAw
VEcJW3YB2S5huNRJBGPSd9S0lna9wYKirgwvC/6hEjJaPMney32WAD2s+OaR3VPj
DD/3oDeQw56avfPhgaxhAgTSIHXHk+m/8jriU8ymzVDaQYproYrRu7tB7F4tl714
2+cVXCtvFhguJUP6OrKp0oTJ2fnu2tsW2ZvR4rY2dU4jvf+8BfU60lfnnOUZnKFv
PHDdJx1R4Uv46QcS+qtk2pVOUG4gtOh8AvFivRrtgjDw1VhVhc2Ct33hN6yijmYX
jRj76tH/1c/dopkTMfnoGb4V7yC3l6lLaIm5QELWHiHpcW2quZs+anDcNtV+knqM
CCxoHAU62UwvhS6N518c5DWi7s7Vp9dzu+EqZ51QXgJPZrO/zECmeFUCRMgNJH7W
Phus1OW+03o9TgTQIwsaveE4q7vL+mn05dfsvI3ooB+zsf2Y51SA8RVFlyNa1nrk
aW8qVkvhCEXAUR6UEtEWPHWDzi5u4jxHpKo93IWBEWx3+5gJTPP9ozce5KddP4ng
1z3S41G8nUaLDI3QBRUTrk5E/Mq/aflmszU/k6WRLCHXlf9q5Nhtx6JQICOVQImh
1z+Ow/L1rwWNqrWEJW4i0q3Qx3TcHyfXkTMTpoUQOPEG3pLQ3Smmlt4q/YIMW57r
6/ixU3g0xvUFxOEhTWRZKhqcJOowqbnP5AEMnGh2yCWcHjFE4EOEPiCCUor6wWcQ
oRJEF4wlAutSJnUQsAFf47ejv8qhTV3GaV4ojE30IkUnEHL8zcECifMtKp17dlE2
FFxA5hsX/BmfkFk2vKjYiU4hTtv+mKck3xO+yHohVNiTU2HdAaCDiyGsTWvuWC+l
XIKhA7wiibBlg/KbwFm7fpDuJVowSWIRSDlVWTnN4dXlkRtBUv6wfRDI/TK1c/tV
uHS4pSx8KyICJqjsn4QoLAe7QQ9smdXFz2FGa73s6f7fIal55PySMcDBgIj3+TEZ
3zjmedT4E/DjNK6Qs2HEZfg1J4xO7qFl0WvxY9WZEVaGjjFa2F3xNUVlOhq3lM63
6f+xGIclR248gncNLyO+x3/OtaDKf41liw23JQlC6RCiZiP4KDdTpwqsACHStI7b
6tKwfiCSUeP8hysg+G+Akqgu/ASBvBRtu3u+M8vsSpUZHNl5ln2uHhgi5CT+l/qn
kMIbWA49RhhOJtVxu9xic6vltTiYGyCQJkHg80PD6RAqLhI7qUMWqiQ0k8RNhdsL
A2ZKHGtU+tkwta/0LF7JzIISdlgIGSt4rGnuB8QzdmKTT6+KhT75C3Q8bCe9S1YL
uAaDgxvL9bjUkXic22UJexqgeRdF+XIjGx8n/7SaVhbHZPlwtTRC3s3uSsqB7vdP
IhlGKEhtDsgFZF3RmLIapXZCexr8b9MUYw7z/sxY+LNXmMcEoVNFkq/lOO5nuzUz
8e0/IIik+GylE/yE7GmaWsHmgeeJbCjSNEC1UZMsBacbb5nrsdADnSCr3NMvB59d
nlf7R4/OO1oUZl6h93qKjU2WY+8mfiY5VPt6jmTvaHaw/HpLp7WaFRkaZGvPfPxJ
2daFpweZM+5Ab8zMkbSTWvC+whgomnxT3X9gmv5CYKD2FAOiyNxPg1gKWmHLtdhG
wPg2QyhNbIheUI5hpdo7WnUfY0P66hShhP5efIyLWiIuE7n+V7pjXTuVqcAjcLPN
sfiGPpk1lE1Y8UYGqkyJrSRX8Yvz0Y/jRXceFl3Tj271jtwhb07gqDgDYnoj6mL+
NZT8J9EtyRR4f2NMw1c17KdV9R8nqmEWjg5Z44GGjeix9wPsv2hV1/6hIqhN3gGU
CWWJkIk8kovznlunDKl1WO01y4ndAg0rH/aaMcjLDAPEiRvLwFE///8CihELlhtr
ugpyjZePDYL/1hYmkfyDcW8/1ldGpg3KPWYWt3NsUqjLi5MvlPG6DBp4NIk+s9hO
FH6bzCR3Ye6241HwSxx3tP7dHIk4bt79RHTYpQv/P9KZpwLQwAfMvQH+kNKKkFWo
GRyODqlbx6P1WAmVLXoU5hdJKVGME4ylTUehmm7eBTAdHfxse0Ct8E5hlDQDxQ8R
HtCVmzXN+X9ubCmFJq7xpt90kbRVIcOS0ARfv2QgyI9DmDXUqXDwOW5W1APG1w0h
1MwCcT1wLosycppyBNK0mruNSkpUgGxNEFyiBfYFAoqYcwRKjbE36MRUUIJJvXih
PkbklzgnsiJEY5pIyB8EErS3F4FefFgw0WZQ7/jMiEswi//hMcpEJ8YlueaTBMSH
Sr4A7EMw1Cl5QHtMup38WfRb1npUzcxw5Soj7yalhL6eiJelACBRaIedBLplMvBw
xSvhRDPL7V2eD4NmtdohYoT9r4vnuSg+WfFgrvuJ3RR3gJge9hG55U7oJestT2/t
oLDsrVrTiXHgkNVQiVNn4X0u2nk56jZvZuTVHIywC47cyy47hFSc7qHRuWPQ4rNT
f5mcrkgDRLtVo48HUo54FlHZmhFiGjXABSHTBxaNEQk+lo3IlM6rAQRnlUigmcOh
JMFS7t+o2NntO55q7s3Wg2U0xVYytNMLJA96d9q9WCPuVX5WYGt4GUX3tVSzHwVv
fqVUnEoNOtZAKfA2MX1k8AlJdKPfNJi7uQ/oC7D6mZlmVoH03fec7VS/jHxQ3u3t
sA/KjhcxF0szZ4FJZVBshHrm8JKpXC+3ZO7MafcFOsVHT9lhAIbtXc7728uwt5JZ
e40r1j+j2uQXodaJpmuERPXZ5DLaHBq7rqN2UsnkO2fxnQ4FJX2VVjJ3trzH5iG9
5GLsCKjcVutpD70bGxzbhh3QZbuuRjdVkrC91gi3pHqEJsujEdZZzI/hbtximsFE
6UmJZeTIBLsrwANRTVCXXz5+DspSu5NBK2wAqpT50+9naKlMqgQwIb8UmEmSQIW6
+ZKlldgODUXC1LkbHXECPSs7ndeyW9hDiDkuLUmjVd/Xkp38dxP3ElmlXaCgYFR9
5Dl+Vlp8vlhrq3bHnO+LgwXhd6IFDUfx4ohN88r6EbZM4FYSZnOy516HiIjogWWN
z44PrbQR4GmYiCHOAqS/j4Y7U0yMB0cIp+hraaF4zcnf/Dewgji+WxR/jbNXP6U9
90ahe8bnmJ6wIJ7zZN2fAfTJtJpEa27go0ymBjO6LeCIiDAWzNiHwEDZD4H2UHQy
gsNFqCu886psMKpMCb50yH7dWnDdxvmlnN1goOyOMeul2wi521MCl/zYueMAH6hh
3maP4ny5x+eONg8rkKJnPFpPg97T4KmpG+gLkHCZR0NqD1qLp4TrdMt1DCbzXUNw
yHI9+URcF4vk5jYcI5EUW/fnohJpTkRaB06/+SOaZTEV3iMbuPptJN7fDx51/XeI
gJHf9jVHk1E7QWPtKLPqyVXPtvogZHUV53M1+ntjYCI1l2lMLQ73K8pVqJ3JzDZP
zZbGphoY2+ti3wQ41OrC2pKWGW6ikm2qFANjTxfuIS7ZDDN55GhDkc5OHnoNfKyN
sAL0GkZ5uAo6bhAOCbrkGUmuzl6fkWW7mkJBBZbhrqZc3O0K7iyB7eDFio23ur63
J4m6MwUqM5s6YXXCFjnlDedPFsnXsORKncjRN5I6gr/uMSxZjmMRvtqiygpumxNl
3ihHS+oOPzJs9+Wi0Sonc6iNJxP5yRiG718uu6gjC7vp5MBwk+w5Fqnx8g8fyXso
bYNN5oXLBGSm7WeHYQ3XVR+3MJpT4Dyc6Jmh00eC+c1SGhXuM8K8hndap9aIwoGH
lBU/IX+W2EuDfMhhbi8k2njWlFuu8cifNJtRZmKwwqs+b5KUXmVnhJGyTbCjeEJF
6e0nsDzWpNKZhNKK3SGHwkwLC8ODpVoJAsQ0eQVAS5X/44V3rbQkp8s37CKOm0Ze
zRpAV7RsxKdHXU6kE/WpaNa0xzBxxHJ1fIGTVkWgT+cyf9djShuTQcwbD3TGAyDa
Z5EZkMHXOqkRvXPBBkMQ+OWi8auGvzIn8zAVM2svcmWYlrVIKN3ugXSdQUAwqSx4
5FjfJcMWS9rXzj7X4KXh2vBkW67q46uevRWJZ6+Z/gBqk5rYxyArcAd7o4pwig5c
PIA3SKi7qtkUGbwbeB4zCJF6yClbqE6nUruU3vC5tzHotBAbkm24Br2At2bQq8Kx
pPbVSbsZ5xGCzYUsc0x3o0EC4cMCxCDfcl9TkYG9NQiGrMCQLdz1fKKtn+33x18m
qWaVML/HUPUYMo8nJNt2H0TJJUFGjWwyf/iC3THv62+CkyEc+Totsdn7mGA1R4On
DomyRrIh1SL92NrI5UIcmtwWdJ5J4PREv1Tm9om8wKjbxtM6bl98p22T6SNcggr+
4jCVOK6Wi1wQo0MVAyK7rZUQn1Osv4OmQxutpGexdpvdM5Dn40F2awh26JPST6lS
W24RGMKGVgN3EIH/B9GwT9jgnftvktiNH802NKpOIjtyV0JLMP84fZsGv29g5Uct
KsRMzIHqdX3xeZVoAfMvD4bY9do9ovKz1AR/i/qFCCmaLm6xEoOfu0oMafDgron1
S0722r3g7hX6litq4vs9yc4QIOf+E4qohVv/Qs/kJgBHGJ2bEnzAmEtfIYd1hswO
0ifpxmE6npONI6BblmEKAa04mbRToVc7nhr34WKH713t2mnon4CJyRupxkdWa+df
C8k2Qr34q0Q6wFkPE4zv9A8KmJeQl01pxjQsXgC9U7XYeNgc5nCBVegICfpGAtA5
Ze8B1a8qh4WqPy6RSXu1CW9nvCXIllo2jyMmZtdQXDWxyi05C/2INk4+vvL6S4tS
uwp0OLQZOBO6svVrWxp7JBDTHVSU9We/VAEnl5c4BpUJaIpvgdlNA+DvMPAzydwe
kUP/epMUNFL0CYaTf05PBFEZJjKyjSwCJ4OvUuOjS9KIVyBkBl7TpEkVSEG8Mrp7
NGA546gQpSZL2OgUzmrCl3kHzyuK9156iOdKbp38J9ecxTsihTU/9IxwYOiJpnBw
VcpdAN5g59Xb7bfqs8Q2mqrUhGjs3kwThPyzhErLcrKk2Z1uYXLcWv+SXc53KJaO
eNMrxFkS8f/QhJWDNzOgKCsnUHb+gYodheF77jjsXwfMuQDPE3ZeB2MAnbxDSEUv
7/0vG2/X8h1pHKMpPOjXTMC9aR8sVn+dsBnmFWA/hmxf0ZVAHH/QwWg8/+JDHPso
TgZ7CRusEgGlqOq4hlJwZDxdY719A7T04DeKhKuOak3J78bAt1TJqP9/ZKWf1/64
/3yJCfQXIjgdgjQN8+YxOPx+tvhKNMHZuVP+t3cfPMzCgs0hicdPIDgMb8eXesH5
AJDbn+P1zdWJORKOSjiPfcCoMDaDWZbLqrFowzBTfDaG7jnylrD/mQGY4bIZ33fW
KVzZt0bsvioeheF9NSd/JVuo86FNpAJ7lxnC3F9VSJmiLdfOSyz3bsossqTgb7YY
fx4G2f026qjNhYcZ1cQ/pRK0Ixpzm95U57ezgLNqGKh046oJX1TVF19csEc+N+aK
cden7Q8bXrq7Cll27RxAmNwuP1g5Du7MQncnn2QlwMiNT8peJ9rcsV2tSw1wAv1G
m4b+x2XU5ScfBxpFPCSpEXddGJOucgyUQxT8u57Z9W5MmZhgEul2QMPftxm8+IZw
sa+jMMxkw5xia5e4Y5PGDoZEcn7uARhyxHYhrycxW7zc/rztcivMZAv5sCym+LU5
PdSTDMZSwBcO/mDu9KRSHjoy2MuJBDS8Ec3CA43OT0JJqcNAiep3O++s6++Mb0UQ
MKF/qqvJ1u4HhaWP74zkhFpSMqdEy1JuG+c+Z2B6pDJ+W3VEDqe8ywD7dMVhjVaZ
PbXyugW7nmSOC2Rbar+aMhUv7F6HGhCMAVPWGU8N9HANv/dOvuC65MxS71BvT1Pg
mqhW9+hE56J0R/L2EJCp7HAaT4jt+dR9o6MeGlnBRPex9MAWV1nA5TZmf37PIUpv
MdyaMQl3ay1Kk7CEcHvpTQAKEKGDU8/U1IbWjXRj2Z+PDtkKkShRZApYXRrv5lSC
I4cwjlUNiJEW29afmRyJDhMkln6hlquOns2DmCe0CSJudqiGcCXO2k8KtxVWP/Tx
Rn+0Hf/d01ZGuNv1T0pF25eQd9yK0oSOluj9UurAUJQ1Z5D/X0nxNUAy4+TQs09g
lvD8yhZ01L2G4/DuDWBzG25deVEsiILWTBXl//KZgEzC7XpAlEdWa8PphKTGDKZE
yDrElbXKPjaqfMfRiSkWqqQUXB35SQc7AyuXOtc2aHwNKPMtUgO58UKhe/YVNDjH
L1QuDJD8FbVDrt8nozFjG20HWkv3GVn6oE+VHUGh7RmfZ50tuPffTfTWyznvGV3p
OKFjsF2fORC5ZTj3PjgfbKKzlE8K1MaYUiRyF/WW6ML4h6eirwJ4jYxjn6uXG3ju
Y3UQ7sLN9Q5Oabqvcqn1Ft8OksqQkGxv7NeoymFQu5pj2s3VTi8Lc8BwR6RhfdjI
j+yGym2apYDmSfw1YrzvZZFMJD5kO6c3N35ESb/XrWXtfof8cn88TQVGxxE902JL
UPjr1LL/Oh74IrCMj6j0Bbg0Ic0XNDMwEPB2ZtOZGKvIJKsTwMBbn/69WrCjeO13
pdkwftN/G/fRg7Agt1wPVbE+kEUYaS7zak/dWCUrP9bUpDKhC1jyLnpxMdmOArSr
OYcY+k0GHM+gtgZGiFqn/VTdnFvk4r4UKRnqt8NT+8cSgTb9Hv51JdLQD7d/YgHV
MF9g8ykTPO1fm8AThy4QcOVqGwBBsnmRk1DvOlqLk9fHYOLyPmCruO9gp+54E8rt
q2WyXOF4kQOJStIa+coptjs4Z8kDE8NeCfy1ZnwDCyR/JDJabyCA1Ni8FzdVsC/r
cTXni1x1U+a07qBMQkofpEsHBxyDbf1izU5+fz40Gf3zNTXEb10LW+CUO/p1g8kO
vlo+o+Y3PH6tGjEHPAtf9mrpeL1SEEM5wH7LZ4YqhiO4ZZlaDdIvBkNUZss62mh2
Zr2Ez9pybLEy04QChfjOKg+yIrcOzx0ZFsMr/b/7d7P21zdowBSJAvuaeBjCUWXF
pJySATt4Uyj63XMD44RLBPje878D2rNDfglLvfP67qK136QhwvBBPz/8hNvGsmuJ
xgOyJsjQt9l+tlTaN/nB9ZNbhVqj67RhvwBKEQkYAhX91rvekZDIsykgyZjtGdXM
to2hCQYS6WjS3z6K+w69SksrWzvYUYgUlKq7qj9P1WzxC68TOz4gPU46ZPuPzIsI
wzjBmrHX03VQv+oXjbQ16DihpoFsQCtNooLO5hCOLpgGhHqUyleIwHQ8sgXc9LBB
qjRQ3fKfdJHZbwBdUf6F39pLIjSiCdDA6cHG3AQv85zpCkoLyacfsn6qSfxVHgBK
Z4RvJDSFMsXJbl46zVE7X4frt3rcboSqgFRffqB2Xx57esxzILwXYPfdyaGiWOdy
qBAFz/ET1saObAXKDT+6XHW0d5U33D5Q0giPZdhBhPcKKoBmQE2rHiPopB1W+mRC
SMBvRY4HaJMFIga/BM9stNxnpzMD1UX6EcAPjGP3AG6O5v20ZXpKD+g9d3TSsFtq
CI3aVvgZnYbSjJvLIhSeAxKn9sih3nnbvVvb/DENPZvyS+BsUvnwfwM9JNJpnvNP
QOer6Iv5/bMaZlmYVZ2WLA0h7UTu7TANoeqK1G9TBcQNPdc3PGdcLRwgP6NRZSdc
UltUc4Qk5o4fHL1xtxuccVPbUcb3hCYIzm7nXyBuvBiNM+46WAzByKaLs0Y4TiT+
VCY7qHmO32GhAQIkxONo7dKTugntu9zrRBNT8I19OjnAOxdfC9nnZSi947RHDypG
3fc6MEGukLycs0aCRxeV+pjOTZusArxvpPc1RaAPKrIP0l78r/4uipf15sM3+bU+
5YuoGLO1rG2jYi8vIfw5PP9FlXBrHdy0spznb9Xp6Mml1AVnKcaCYkhbkCoteUyo
xVEqGpYOr+MOvuuO6uiKPCIdvtEjpJ2myA7u8Z0IMW37daiODd4YhL4jKfcEFAGe
A24rpyc7LjkoRIsoHf7hKJIaWjp0OHKeGyv7h8RWL6gtDhRbxnTfhojvLGWBnM+0
cHSISkpsXJ9U1ZjVYYtHYaHpYqZa7cG66EroSNLMmooz9fers9gtv29cxkNKAtYy
cq/dgkuM8yMJ4C1bjyIPv3L5I7zM9//54ZFm6Dp2CgyLBzHn0CiWQm43itFshUS/
VHK3UixPVT/LpQFUz0bKCYZjORENS5C6OsyBD72jkFF4cDc41SKP8U4Zt3rCmq/L
544oMQYzC9G4irE11lmrxFVP3OF85Wek9Gf6h/HZHvjAS0jsVi1Dlxqfqt7a5/dr
1BV4Ao0W68Pfa7iaoYEdxeHvTRKZk7pmNzeTrnhF0Yj0GQ/LYPTqNSGuHksJUiGA
JYc01/NO90LrYKMsIu+Er0hNQcv01TEAp0Q9JMJfyc4BxBdj03D6/zZ2hwT/A89n
WA6c12EAYvDRgkPABGjpWUZIbfWiNg57JS24SpKweU0nvmLfDan25t8fVHeTu3ql
kE+AB3IHpckGRujJ+NDhwXeXMRHkzZNfTkOmB6CkdbS4L4FQyh0O+Om4Jy5NPfHS
MfA6Wi21z+hDbsPOjibeQC9OYWh6pYf+gHavCD+GK3vZpiesNpjF/DD3K0mP91W+
jbRYaQL5WtYfCFxsCzaLM93kXoe0wN8007JoGndcOkFAnmx1XvOVEGYZCaGuekt5
RLDZwFCntjpuq/oNYxDJGhZuX2vBlQPiGDkFRcamUhUWvyEOISaY6wVv4C7ueXC9
zg7bovJLvQc2W6wki7d6VRYTsUUtcx9gXao/ptF7bcVV1kXA1A/tdNDS8brSUWMM
hTJZnTyVSRp2mbMxSTUarFbBHQ7Ba0B1DKT8ViMvW5di+VdjfhH9nzCJOtHb9TQd
DvGZrZKj+/IMLICbTWXKsJzbZXhAEMi7T1xe6TIo46+Q7IvpRij7smttRWxGpo6x
MQ9seRw96mPBDaAAVNG9ZorrQRWLKApjhf1UBVoEqi8i/NTbP1/ytjwAry91giUj
fcpKXZ0yiD0wMarJ3FlLs+wS1Q6DbeQBel6ymA1MVoMZgbhazF/+WPCMHI1nDe98
vrlO3w0S6hCi1SbYC05ldgMeFtJaoFqsg1lNwBBdlJ/IxFMfWVGtQMX3wU+4xN1N
BMKgitbCWjIHOhPKHZcVMfe7kgAPW2kp+FEK62OJJuros/7Fae2A+tLYBi29L4xC
LZgnWipr0LMFrr4RCogTNHicTKJnNHOedVO3ytivJwjD+2zS9Y/beAmFDoc1zWjQ
o63RHW5OWE9UFlPrajRwpC7R7759yRlGP5aFV/HiteXvqvywuuv/X8PvVwOo0Xyj
qhJWUFSnlsqcTPrUD7Cd+l4IbzBrq+XKUTwLnPQhCYSczNfs9Ey1pOrROERV5U6A
vPGa2k+2jT5ZQVjhHyQN6rhCyCYLzHtUWJsCBDgXpL2prwYYzGjvsaStIVTIRR3R
YirT2MWZOiVjWFNnZEVRyEqT+2yuOFH26l1Ssg4qL5mn8fWD/NXVYE7iIhVslWR4
X/xscdrCyRkUfFg1mD6k7LkJZgfqIZFR1Yc+uiYRbUSqfSqO2KV6zEnWhKsdz+Fx
gA/gKXtbMgi+lM0VQbrOVsYc8xW5KXHdtGNMmVriIBEitYtwZhiHkuSkz+ax6tuc
7O3Dss3m9ICgGBWoSlUy73DkdE6jr/RhEG+JZwYobpJGe5gQQ3lqK5/bFI35XFnD
Ud4uMJMVgIsxdueUXIetipGwQGTwR2e3DNh1rXMr1qiXd9VL0mjhZDIFaHGkm+vx
+bdVH2wTbfpaz7lIPY+C6JEZwnTlfJpn4Tu/obvDX1dX9gnoHePkz85O2DCRrGSw
Vo6kJc2vvs+x01g71dxyZqwoLvsl47fQg5RVniIxNLhkooFpOiy7NYwKg6e6Qfma
F8RqS8cNmpkx1dVbepgBtLC3wKTlBUupN8IKgw3V9hlKAmDJIVUGi+7W+gmX3BmC
jVnVbs7O2TWXBeg6hFF/E6EbXoEMt1SdqNYWiVOob4+RLHfi4eK2BgICd0BwY5Ke
Sjx8PmW8KiDzztCa6pSOrqP1ZytlhElYHI7LNXNTJ41em2ZuOzhgzXg+k+TRmOoq
/TpPiTAWKHFKf0eL9Wdf2hsiTjR4j/ZJHFsvQHdWscBmYF4rEdruhKzTJlsPSA4a
ltiNWh1TTY1cLVPvp89wuc2lt7Pn9ig5bfQgybNHTLU1+KfkM0yFavXblUUNtYl/
YsHrAwqconB1dEQxhIH0MtXqVnOeD1AreNBp3FSLCCdPVBiKD2Q9NrGvnS3h9vL9
Ro/HQlyZYxoXdLxkWAjSC3AIz5+Y6/tcM3NjVGQugTB/vxRc4KVT+Ar68GsSmBwP
pdaekTaZkOMoivYD9haO+yEwlTrXUc824IMd2UecylLvu33LFtsctAoEFYr/pxzm
ZUzaQDws3ofeDujZIhBD7RtglQH/jejSk3EXXpbpTIdsd3DsoTABvD6CBZ5/ytbU
oBnrBi8Xptx3nO5H3U5UR1E09nPBh49e2FUEKseJ/SLi6pA45XjCSY6q8oVnqo2T
0ojX5XmX3H4JRLN9DHeWsZrAbRvPf2qnz+S8bpAvtNwu6ypY72tjjI432pGE/9k7
KgvxCKlNMHPZXs1JnqB5VIFcQIW0iZVQe9l4QjSr+bS3psoYUbJym3sOxyVoBDVk
s3KyT78n/rv7jOXwiG7bNQj2mflpS/OBNDMKIq0Y29F1wTLpSp8PEnV0UHW7akD5
iUEP5YP7OIMA5kyhoap0/77llASt0LCQIvwpBUOxA31V7JDCLNKSMQINCrCyzksp
Pc8scpZNZcswH+e6kbGAWqCmoIdsognGAe7Zbuhva+cfgiYMQivxVgEM4ZJtGCs0
HOA1tzSNEDscqGfiZO2tXDvisU/vlfotWBRRPYZF243ZxOEFlPUpiBPPRy7H+WGh
bTNHSIjpS7lHt392FmsE3IhokQ0XdN4AqC90knZHNPs7AQkY3AX2ci73iB1736zd
JuazX6mNEoXNIIr4TRv5rWRSHYl2Ul7ZV04Z6X+9Sa2VPu0Krk+EvjeuDKQcbTn8
OeGYxQs9Ewb//TPwwsP/sTobsvDCgMj0xz9RNl+wZ3e/FAwtak0fCKJqc5Xr/mm8
U7cyhNZc+stgN2tzPmdVubRV6Wx7mfZ51nCuoKqerKVmIveafYrXlDtovhr7jHeW
+SyDv++6ndHpDyywgexq6GsFqrvS6AsUOVeRUREKz5vYzubV31VHsEptb2lDIXAk
2IUPiMkd1kTohdtWcjKNX+08u0QVgHUA6s5wASZfpdOdYbEGD8kOnRgkCbipSWBp
0qpMORXCcxySIzBae5oiKDz5N6DcXBiX8Y4T1RB5wG+5SPHz+wtVgQeC2mNtzqa5
XGre2q9ncl/g6KLvrH+FgDwFZWty7/95YxeAL5fEw038PhCiyFkO0CRFqn5RlDe8
0WjMtlZ7+ui+mbslVY83AUANjGEMj5VvpIHZevhcmbhBQn2Z7Y9dcGt+VlT70qEs
zDT0AIB008OsAOznk0XqDN1eBhoYaz6sDNyrc9pDDCLI5f6MgXC6+OmWdtO/RmsV
pjwe5R+HeuluJ2gXWW77wrPOywJyenjVyHFXEW1aNhYu23FOJorWoDiwCD72mbu/
mGrBr9Pjv6If6uoS4Kn7d+TpefkGSUNJstpblJ8AutcSuMaup7iQyUaRoMYQGqvD
F9SGbQI94Qmp94IEPgWUDEcdXWnL28lYi8xngMiNWFcUFF+GN+XQMAbff/F/7dLi
2jl8PF3eXSyEQxJwLaPYZiPTT8afWO+7qg9SM+zm+MnzpjSEBGvTLnOJ/Oa7/Mfr
Pma8K3WTVaAT+I1MkBOn2xf8zypaqane2ML+1gtIeDCbAYZnOtWi++MmTG9SvHLs
HrCJFM/UmtL0kf600wA9fPGINCB9qo+4RaiuLnYyjDr5WuIaJisc5wACOpx+1rVZ
gVE++aqteyZHL9Lq+5Zc8qzp6qHmmzZLQ89mht2qzFOGXPtn56BgMQlVNymVAiUq
uKFzfu9UK2p2T/mNIVvrfV1Wkd2mDSKXSJukBUCU6tkZ77lENdFFjLef+tFXPa0f
HDXS6UWtZEmV4mkJ38Y8HfcCJR7QOv+98BAWBdXwia6R6yB38gfSDGcQzIpaXVPG
pRj0VCguI8gNQ8EsqoEsHhvFoOgVTHtebbsBTalx56/MmFhdzx4W26pkJL8WjgQL
CP9/tFm5XzOqAb1JEZ69LVOpC+K4QjkP10kgZcUYlUAwu/qGLgdgv7Li0/UBjY57
yEjJs+ByuwBSgJplABii7rIMCARKZdouzKM/uGsYpd5ypxgsuvmcrcptqWDhB3lb
0d5siPiU1kFz3114EPWsTtHW+JJjwZurjID0ZUQI1WxfxOnzMWg9tv7bRuKTKnIp
j2UPwyUhkbSUe8ktS9Wby3Y4czVtZdBAl/6WtHnmzZilNEXCVj6lRnjMlyotW4eR
Fp/zeY7dURVgXGO+x4w1yUXgqkZhC+JM70zVUJyaoml1569hWVyWz9ZNcIFt/Bo7
32nBB6t9JfQYEBUgY9tsyE8eyG7AKteqxWM9MgciGpJSh5s6smO8gUiZ8aC8avG/
EtcXrUW9DOpsG7t66BN5d7rjKQhIVGb/DYv5+BW+mcqqsKw9FjHVvJDFxGSYFnlk
Ex/gDagqRbHQdd85I2Ux0wh+72Zf824x+A/fPZ/J+daHRP+BNxXbC+dHgpJ5R+SB
8evhmEKn7GEnRMLyDnVCzplQ7aez3WallTk4MUjM6Nbao1L0mOQdkJvK31UkXCIq
/uR0XLpiLYdXR+NZ4tib7S9zB/lac6ZkwYI+1O1oC4e3Uo27hEG+K+fB2EqMHowH
CWir0cLfQvsDgFmysAnI78TWJE2lbf2A1ZGNCIpdr805lns3z8mjCapbeCsH621h
gi/t91PLl5QvKjhD+H41aSN0Cf4JRY2ZuV+yLmny/up0/bU9+/0ZY2bn/p31sVW+
Vxj1cyuAn/ZeCDZzQ5bv6qr3CSpdJkcm+lK+4yqd0t7I/NMV8cmUX2dH8LucK45V
7m3OD8mx9+voSSH3VxP4wjFJNa5n19Bd3M3zihbZmTHkUOXDJaLx1UwRWjd6vLxk
SY6fpvGzm6s7xWWqrd4SbzZDgjC+KPaadKP3PjMM7JI0hXBVxsXb6VRWVIN/bIud
xVXdcru0yUP+iUqPXdJUmkvve8HwZdmcjOmG1PcMe7hNbRX+4l9ICDYteumNpCcm
KthGfKFu/SkTXxsJGdwv6CNjCDktnWTLWfEkYenHkoUj0XoWGBwEFbIB6egC/tmb
9hm70dP8rC1i5V898DneiYachMASj6Yfzq/1R6ffRtnNvv9YIjKclFqeBhtOh4P8
yT1f++xHR8vZyJi8FHAxu7p/vq5lC+YgqGcFNRBNWPZVntp+rjeopOtLj8trhF7Q
HpsAqKn0kWDMy/7ebE5obHIlc3W01gMcLER4iTrLT9TC0/rVpxSScMimkmmmMGNE
qe7V4wBX+T9bHEAZ2WM5oP67K+i5x83ZcLmI50sK007NTNNOnTrqoD3eEdkqIBex
XDVz4VJRihciTsTiR1LIT7NKxydJvfxrRdWwo09wkPqdJzbWkHm68lssxKDxpbQR
BpFLv/mT9o6l6jbobm6j009GUKv89hLu8AnCAAoyaYXjezZkk+kQ76pDOBjo2tRm
/oX0PUyCQ/layPddb4tKyA3kwBKmkpFFDaUmA6/caRvBfeOaS4O+zp0jtQzNgEYT
i6YY5DewwMJHfjevn9uC/VxALX2DvpUmWL4IY9XgMxTEWOg3XmB3pLAuuWtI8vak
f4SxYaGzt4qeYPXxO/ZnDtejZg51e3nqLOHvlj404Zge9UsuTVM8FIkU3I/j10cs
uCMTU7GtGrasjyU4xN5cspPNYTBkyE3cNE1sXhTyVy+l+/dN02yL9i+zwB2gk8lq
PJACkgRY7cR7n5mkqmBQEM+mWJySwt7DzrNB54t6DB3qawPN8mWP5GxzjViTIhuN
ut/fIEosD+QTgjX1+weK9OoJNtE9qVDTf1hjGzV5wCW6CDPsp3Z5wgEHSy7musk7
rm+jlE0yrJgahUklKvtCarpjcbRxNJ106/M437sh2mEWXl+n66IkqOa7bB5JgAO2
K2q++Qybs9dFTsGsyPxN+E8hthVhWxKAp7pF/G4yXPPdT9ZkZKbvH9eZM8dxlmz4
yZml78R4Eb2WbN1/+0Y6XLIZVCUcmoWHPy3s2zPPNh3PX0+y9Cx3tIJ3cscekX8D
zmP5wEdfDb/2JEj7HuUhZqv92sOf3YDZ76BYeCqisV6r14Rpuyb9cQFUqn77GTUB
0LIDyaNKcJQgeOp8qLYK97cAZ1/T/4EJ8E30J2SzbTmQLMad5Rf/54nf9zQgDcqN
BRE/C2cb73acViM0wgT1rNyRDWJAJFza0A+4vKCh067Cmbsuzchhdf/1Qg/XBrxr
TlNaBlAq5VdWe7/hRKjhPYZ6gvk2nbhm+zRsC1cHy5A52Ib0hnInRz9v3e/mcvlq
U72SrujmLLptEl4dmL3sWmdHDur2N5Ei61v/0AcSuuY04Pj7Vd/tP7zZXRKcjXiL
N+o9CrczzoxtrzD6q+CxTywQvcnhDnxK968ZrEI7hZS89D6XY2I1kN7q6JvTkeeL
LxUqrByaEQ8VH5O06WTbbzR68Dwho+PK7sMeATaZi+wn3Ln7KdMH2THVlLt1uEh2
qIMKbX+KmzwyOoVxWjqwt1b/jNkXCs5z8SOMDqJzHiPYD+NR4W+OsPOw2XYEaOYj
3HJNMXAsPjPv9dbwN4OqzhY26cti0EhvUL7oSocfhzQowHPd218eAzcMLzq3djh3
kA3Pw1+O1tJ8+bJKOhHY5Mpvhy6NGH1b5AN9pjeeOlSBQHl1RYlZCfAsjEEwq1Pd
+typ/n4KUUUSOxNlyWQsqILqVWUYm1L6aobpnY4rjWsd0w3OyuCAsIa31CVd6E5s
xXV1/6Suy7WlBw+OIaUHeUCHHpnGGmAhNMlISNZpnndgaAazuruwVul4u7UUxMdX
8BPPlsZqA1b1oChbDHfw6RTIEHRQA2LffQM+f61M5zHqj4YDx7j/ZJE5+Avbw27M
q06W7xLYKR2nycm8SZVJLJWqnDHvazj9yl+Zf+6/nqv5aGexPr/yMpqLyNUOVtXD
I9u86lTOXpyS4y78iDYnjQeU5zBX5Jhrja1GdIHNc3ZGRgCeVb+lLBHgeoMLPQvk
0ZnzaPNAchlTO8EJ1hBOYpcEjOd2EtBLPMp23c45Cxk5F03ZnQmRnJ5Nh9hZ1/iK
5xsJEH3G8MLrca02i6s7+GW5ogJSttbi7Rz+bAnt6ex6vT53biT+SH2RaUkYHHHK
Z2s/ydRL/gygl4hFXv1oXPBAcUM4K5wQbHd+2TM6lMSqmkXWRLO8h1VipL771K2U
/MH9j1roq9+VOy1vfSrjtY9hZ9GtqzcBRwFk6Yi11aBfmUx07exKTqSiUY3FKetp
9txqMnaC6iDYR2t9JII45XZ0/VvjKocWomKOcR+y8xozuA3mONaNxDSQDQStlfVk
JDA1wN1aMrh7gdrRM8KD9tFjTB0KIsoRKdXS6N8QTWyJeV541Kz2T0/Bd7nS2gkZ
tXa+4ltLE/xDuN2pWJi4GOPJGoFY2mDQab4K3VJFtLckT51nA0BVBp76aJjn9wYB
UXC8sa6LTqWDv5qpp17OBgSSHE35/IRiEKNwpz5jq1PWUTHyIj8qz4Bptw9CxAra
Cd0g2PSKZrkhby+J+vKqSaiDdIQbzcUPbSvQkltPKNi9v2nI6u25xRGkYMbDsZo8
+WhvGe/IQt+zPH+a7vMvayzSaJaKPN7+Le5aoTYIQb6etn7HvEERGh/ZhQvqpFtc
l24bPRnPGfmCFuKVaeS4pjwFJEMRRq1uueQxza86Hm/acNBSOQBIAqIBgAhUXkQG
OkheWZYq48nKqaTttsjWaNc8wH63TLaAj7N44qM66fc2pcwuZhH5kBTnXAPqlRQB
g23sYjVXbybflbgqpSGcbPuJL26hGkLm2L2WSrVNpRXDJiFTYfXKtvaVrUKtp5Nz
MXqCeZ7CXs1ox8az/rO8nl4kaIhNnNEBs7fKWKcRxeERrNVhgGZFyrrx0bkJ4mvw
lMwV+JOx/sK5jBBegsSbU+gQ97stXNL8ndovqScSsg3SjrIvYVjWhsonYsXl4Rr6
K/pb2tVHy++qzsez9RXR62EImfA3LLpDnacS3ecD8hHFgKyoZew5XENtg4xdga3O
S3kf+1FOpc8KushzaoD0/65Z0fasxkGop/eOG+7iEe/UlXWLu9uWX3Uf2fKQV0Qy
xIxqi6sEgG5OuKckqZZU1UK22c8Pv7Dv7irRUqSj7B0f772BdJtJBBMf8b5OFfdh
WtRasJsKQ3LcURWDqX0FU/Ruaas2M7kZE6CJrbcdkNdlza0c+LcyxMmMX9G6qtj/
d3w42w/epDyQfQJYqKpe2ijEAvz0EiYDz1PcsHjRur3TDOYC+zTx+9NFtiHsN+Yp
2E5UpR9jrRVaX6rK+aPDeSGqNYXGcj+GGNvpCQs7LZVU4hA9AIu7ttEfDJYqo9cm
z3TbsIPOueUu2IZ4KwLjvG72606QjEnaq8FrNdonjh+NuERhXLBNz9MsAAxgP7Z6
IUbE8BH7xO1uT2QtzBiyJ+PRHUvisxkyRPTfMFyjUmJRad1J7qZMSAxeQBZBXTL8
qDPj4u97soQNjwpdZzQRbSr8xxpwjsFzxqk1Tu+G2rLLGw560xjcxDmtmfg0DHjP
SYlpWAt/WPza0IGzG4s9wV4dM7T3Xj8WnP+q0qmT1CdmmRTD+Q9CSAS33QSmYPT/
sWNC1IVgYeRsx72aaSZECmHNClJAGRk9R0+1/Nmpy0G9MwqAF8Ec9jwhZB24Bumg
XMCnmvn+pKKX3YzG5M04Cca9VbKvqEXJ7JEoNc/a/8DB9y0xaQiegimYrakk/Mqu
N3pvhU/73Aeutl9uDgkVChS6T7HVd60iq+IWgt561WmKH/m155EgdJvPb8aTnT/e
z0vWcWCHWPbvOB86++m9CgP3Biz77gKPOMZ2BA69u9C7uwPZVsiTtf5jt/SzahNm
lM81UEVPN+Zhz++jhDsZPKpIZwYRabqDfgwZQvkiv/5Rrua+FzFSIjl9D1+UgZz6
AngK7o12Mn+ZtRWMsKShIMpVYyscfiQl7uJdnJikTqsZo8nof+MuOqmK4obWDobE
LS/bbDK3mDk3THa/gFNzLPfXGrz5MYcfXzYoyEDNBuioXEg0zyFN5eDEN7d0/th+
233F2xiBt5N8RfCtNenmViXi+ZDVWKbytI5DtlAksftXbMN2ogtr4JpRrGjCiNIm
O97eJF0pegj/TQg1uMgwxHDZkfYRLYr7q5esPHsKQHcSuwk3q0PlEjFcckHZRvub
63mdF0EfmSG7D3oVfiodArDEG8i976crIdiwNdJXd3T5mIr8NYU46Ed7Z3ekcXLR
IVFrNsws5qq3ut3UGUpxpCxiazr7tg4lt+zj/Ricd8x7Oor1XyM0U3f1X2HHdR8b
kjmqgwJ+sNZ++8c4FGh5z9KjORKwVPIxCJtJFMldE1EdcB/vJ07RF9qETGMFHWQw
0MobO2pmM0JB/eFdJj8SBFe8XnR0C9MfsIzyRkJrOD4R+OiqNgbGaEKqqFUMoG4t
rXxTfyPdl9a7iKZpQaRekScIy/vzAL6PYdA1O3ddKXIwBmLEjCgZnRhNEGj3O7Ex
nihTeWK7Mvlz5RDjoT4q5BrM1P1FE7Sw3CUIE62jiIg1WCBDaN2eTbO8wAas6RJS
9+mawWxblF1Nf8yvJgZGHsT/CeymnvQYxMTqWCJ47lXg+epF6gfDlwBBD7xBu36J
o39F32fvBsp2QuDUwsDFcC2YZGaxaG38Sv/B/6zgFK3Tm5QVBiucMP/4GKe9/vRn
j/xjl+xM3wn66vLMvd/vMxuJM2VuF/z3a+1GC2B8RVnykPlMXjKFMA2SlPxx/jdm
sbQoTqjNH38Jn49jE4zMFT1finqXe/RT4Ri4zt5rowF3FL9BfoeV0gkrvMW/EXKr
Q4cMunQqGGCjAboNQ5qqmMn3AVp1hBA2bUMWQiwP+AOW/RF0NfB1V1E9VBEbwfO1
n6iOh3hV1PMnefVt002EsqQU2pH8MZZX8Qx++T25r5/45jyRZGwUjMJMdpLOzvqh
djOCvIhUFbYhP5z439F9s362DbFhLbXdL+Ec3tkbXYGezMP6XNGQewGTwwMcYVvZ
Chr0BasG7uKBz0pTsGZIvSalBLNOZ+im5jIoCLTCOxmQs0IoPm3EXBwbv2B+musM
43SDR2kj8qiLNX6i8sW8x/WA0e5oZWmeEgZMQi+jCiIpMJEWiBrT4fxkTSOIS0tR
yayfjOpmBq1ZiE3Il7dfMSnm8YvPVjYYUvv+NaTDJNunKCLQzElbgchsHSDFEPuH
7oWA6PMRBBSwdk+yo2Vjqko6AX0qEJw3TvaHBJxJooAauC6xG/I+ua4CWuy2XBe3
amI2Y15Y9LavlB98unm76Cu+rxDfj53J23+uILegXrgvUTg9TiJcGF821B/2tLdg
Hcs5YTlVTfEzDT2QPUZBlb9GTfp6AK+E7vH8MnIn8hgZoYmhbstW8+d/ce9BiYOi
aSIdbADKjOEQMErk6o5IeuA7rNWvLu9YYVjpTxYirHUg0YdTyiiENMFYOf6mMgg4
76aemMGI5rKLlcqdkQNBzGvnctSw1JPgVp48rHHiwTcYBnWLOS0/F/xg6PQC2M4M
zinrFh5YNljnECclhSSXq1tGHrZitYTaGdvHbCSyATyMwPOofl5W8EDUKvC6vsNs
JGseB9Kx7lMWw7nIccehXWSy5sguYnFjanG3KovbHmIG14k1F+u3YUmOhHtpUKMU
GQFsyDcxF9192+DfqbQt5P+OiyBH7Z6aVF82QZdiyee3MNsBy/3RpBCOMn+kQlLJ
JmtppBKPyb1H5FdLh2pkpE8Gs1NXmJzZMyAaxuD1ngW+iF5euiDEVMKiXsJNkvPG
f2SZO1BV4CcZXn+JYc6ogR1OjQvSBP45xptEzWM5Leta+8VuTUVC75xXBitlRBiJ
IfKn74eUk5c5YKe99PIIA6NS7ls4bgwxYjepI4fiCDDeIjOrLbkd0guCNbu0gFkG
qqBaDv+NrY1tzxIundrBxd4J62VKgu6VW14+lRptGpr6XqfNhkRPpAoh2uPaPpjx
zsERWES6B5xbXUDK7RKGk7v5zvANr99MkLLpZND8/7vgSjhMVmTg0l0Q0GOPLWkL
YlWArdLslcBrEf5OBebp3Yo8t/50WMX6tmE3lFRiipxHChiLywovu6ZcjPy9RPge
Q1GM2phV5dFFO/z3B25HydOw6S/rfz9NHRt4GHQvVWHZ20aKX0W8BrwmUvs4tVcf
fiu3lpEGnwypQ5afZ+6GqIaarXogrzeK2RuwCP1PWe1DU4ydS4/+vxFjq2hskv6z
+FCMtEGnLGQWQ0OlHTk7nwI5cyeFNlVBeYIeHQKV2qRq/osMMwvCQe3m+BeP5+5T
oFhrNMvhn53iWQYR+LFhUyAzDpMonS+e+lyTcOe07PoSdrQfkRAQ9UDY0jBBjnjW
6/xa5EzM+Egl+p0WfEHcMWCMP1zje8ky4iBrXTR1aVvzPjkjGHzAaM4SpRbGkYck
xEo34wfHz61N/2abX8K20I08v/1BN7RuvC2Nfhs0jSzvWUgZtgzWVduMFjLMUVZ3
qwZr88ekORLg2fDrPOWlgX841zVE1mYHOJ8HL5SQZqj7BeaFZAOz5R1IokHukkOp
ohJkFJygUDS6Xd/mQEFO2o5bfzeXfjn+zvQn4qD5HgwoMh9Air3a23JYDvMe36g8
22ZWXDP93WxjfeZUwue2SpfHJOBtNwH/PgmPSiAfnd7bLAe786KCYGBFGu9nlMI3
QLjW0QO/47/5czwj/568zxsOKV7ftKstTEhFNHviUIXMwMbyK3DjpyXT3QbDubpT
dLj5b4ld1TN+wZgct/HceYordz3ScTR30ekUGzoy07pCJM8OqVOK+S1tXpH1+r9v
dMf6fPixIUj13kfeP12hHTmY8fRtChadLMkhIVcLKEmOZNh6fApRHv7kn/vLzKpZ
cyR3JawrX4Kjgwnl+PpMJnXGMhKDmcXAjMN6xPo6Ar6sgMN3MN7b5oy8FhNzfzeh
5DvpLmp6+9Xc0Qlit5ETNZxmCYCL4tdgxs9D/8f03MgbVNhyTnCE5o26qZoQvbzW
ekb5e/joWvuebJA7pgYzY74owbvfatN2HPHWyHBPAXSwqTTSlONti+Q/NxohSCKW
BOljJ+nBBEFQ4ntXMW/eM6XQwErXkDSgoIVSzvdAMKzOPKB+IBjE3prkm2Y4srg3
tcSV5+r+J5t4b5B083V0whobjXCR720eue7G8/arm6MbfY9r31+tptPkcPp+ZDmu
hi9wCfsxG3GoQe8TYpBH51lMvmAU5MaDrWMMZRz0WBhM00+mkkR1YY3infg/ZIvi
uV1/Dz9nW6TgSW6rRCg3edAPcRzZE0stwuvLZw9tlzdGiiJXIOw6WbsN0+8Rv1Zo
vpF9eS5z+EJwLj8hNttpYc5Zb8A+ySMrlBNx+VcJEuGfZzGzXJap1HCSOpSAcAmX
6xXUtsqVdAl8xxZj4Kl3iS1jx9lfxythcBTky4FSOLQIIHsalz7o1YgDIgTPcBEo
7DcKZthmL11RU65Jo+6VytPNEVptL2V0+b/Ku2P7PUJ72dC6v6UyrriOkWKqZ5gt
XaoWeFYxECtBL3CEpjbivZ5/wcbpSHI7C5mVkRFiEV0SjlWnwGqk06wzBAYjILKd
ZfWEmkQXa4QjtY93Y3PDQpHzMX7IbN/Q5Zf6WXruKRnLWr9pQf8gP/Lj1HtTc5rE
ZD//ZN7FkMr2fEXntOtu/y+lXD39XVeivKXsbrJaxlQKsbjavZjXr7pBiQ4oGDHd
kXRIMNJpRYlS1I3CqArEl+HuERLLZM0hD9k9GonTAMM1n9oeJEo2jcW+BH9P45pk
alBo6eFuZRNB94VBb2d0v9ghP6CNUbHVZg3UbVCkxR3Qw7GM59Lxm6bOwWaSe5pw
sNvcFJWNXagl4Zbad27wqwWfOg0jucpCTFFsDnNu5lCc7F+BNt4zYK/ApL0yJU1E
bUIDwMGa3YpyaAzjRy5iRYTR0oyIGxs5J+YhEu12dy8NxTKegylnpsILoBwkMylW
1ZHaxe9CE2688XvfskTjpzFx9FZUyLjfm2Z7kxK5uwZ7nwO3HHidxsUnPqXeI/GO
uPBzy53w6GqzB8wzjEkhgaW2FE35E1wYMi3x7sD5LxlrrHyRhQxBjbbXhOWH/tfI
8MwUXMdzl+OkK3uULgaz5ZiNJdVIB7N82xPRl0I2rylkP+PQir+odYHQd0ZjVLlq
+3xt+woNT9/iL2SExYxpIZ1JBkJsUJgBY6DfQPxR3LnU2dxwhr3JlC77R+rHHbHs
laJm+0fC57B0M+STze73p1QCHNTtevRrVkR8DAYna9cWhnQbJ+qR+ASCFJDjzeG2
u1h6iJkGWbi0Y2xUZM2IxdoF6kf0AZ8PSHZz9jm8RzBmRK8USbdugyOSUDZEBO+V
CXkbpL1Dq4ofXy7vkq72GglmYG0abcX3IpcS8vVdJZVztSfqIOe3tJvZE3+uD0G2
qxTtGn0VlyQS9ZCA3W1cQelXDquuuN7XGlcv3i0dVr1rdBUd6c7FUOgD00pR0Fkb
MWccLd66N6GijzQUPFfMBydUDlVNaQe74g/N2/ZDNY6eZoKTo2/kJDlkkSpL4gaE
tr09dadZI4uDMCDGBHRSh3w9zhqSUNCeTgs+4HC+rQsnHl37pzb+jqgyQtVNDCEL
aUnANI1FJfO1NyzAFWv6BZw32P5TrAlnZ7nyMYAddIt/m7Kd0R/a58s/ufR0k6QV
wmIMIYwShHXkzkGtHv+wMh4WiUnFdO1FYqyZQ2V65A47or0muGBjqwyvwMrBIZAf
os0ArdUcU13fqZdAMDxRMRP64IYQWphymo9GUwTXrWI66ldfp/q/3amcTOK0B1IN
qC0X3Oytw9xia0RB2r+cmlJCc+DwbxT8vx41tj3FjAxS6JY7+Ur4AvQ8d+K5fCmY
muVoOM1t+n92xiFEy5atTtANEHqxlEW7xHpQ6D38eOf+8OU1rTyFHA9drUOSc6Q9
WG994qh0lERGrO05S7kXn+xTUEARDKN6jjpADd7/wW087KPJanSYQCK/pOgqCiZI
FwTQr0B+VQBNbsr/Ch3GMVEE9XBSgRZXZC643BgREPLxkBUeQ85XvD7tIzoNqNOg
P6M/PSEUyiPjqs4lzWd9MsCWok0uz4ZrRgqLwxleRsTPV7wSGMzhknRCIoC8+D6H
5JwxInXu9NWYnTn9eqygz/d6JhJPm/BNWA4cKznHcOy+zC4mkzaCljqlZUrJ1vCC
+8p0geT4Qkbr9QkxsVG4Nm9SjVVB4fiUyAc+Sxlhr+4Rzinv8ZMoLKSa4zZ5G+BH
SjDwv4uMMGiDR1iCjgzBQEw9R6B4DydIskkRJtoPQNrFtRvFAC7ewXTpDbAn7YSE
Fk7jrD3m9c/xOIfSG9Tb0tCIoAYD5FSAfK/QuFT8tUd/eTErYuwLdxOQsXIU7rXY
MUCADGM/PJ1cja/x/fWxEpSDd+KMzKZs6SUcuSGKeGVoZUZ/koYuz0POrmXNGNFg
E5jevpgKVgNnLZSvDNnXQ2ZZEJWfsHrAS50snfZSHcjGvCAfwVQyxBlh8no3DzHZ
lIY/F6s5qaTcemSs3eRvCxxrd7cQIzF/61uuJ617ZpvHsiK5upkma9TUraSrQo4o
jMz45Tw61BnF4cVNop70FmrBjT9IPGLmvPSpUf52wtSbGtr9SJK6HMobI4o0SjBP
FsnWrwL2P7CY4T7pQn/UVt3tPWae3OUcOEydIBUJgeC/R4KMeureU2+jL0cugjXB
5DyAZ4hjipw2r1MScn/eFUv2biZI83AQ9XUAnFvCGZKhIGz+3NDYxAPA3WFChv1Q
7aYaqYdQY/Hmo9xaNPEBIslk78Jxx90CgU9N6HIqx6ZtWxaFfjBUwQcecomcwN1b
GaZs73z2YaCrXVPaPgqx3TFkfqDqBKC4WcAQxP0oVuxHgYnDPwC3BLWm6l+/AYC3
OxHTiEpeOth2OYxTSvqzqxss498/w50+0s4rPrajypV+7mWxzSd+CRtaFjYJ+eyb
mqeV0HwdY+8q6HM2gu26hoFRoJae/yIoxt4ah3RTWcYt7JT1jDSjzWxTc9vMY5Po
274+78qe89u71p4NEQGCifRL0q2V4dOOQNZsmZ0wxl6efaFA+J3DnhFhTeIGyi6n
qgfhC7m09wR20bSTeM86HPr3YtWwAVRfFPUEQAGpO8ACUwvSv6HZRtLjzo2APL6v
qQF4d+HHpiww4/SDWc8qM8WDeeLH397pn6Wyt5G1dHHDcsyX9Xp6BL/52BrUAQ8F
yItGKHlOCX2P1yWmDipQi+f4NJDzB6nsziFEOcRNZ5oDlr9P5KbKE63DweJ+eiMG
X8hDhnAzb4D6Uk7Q4DgC5rKjbEhseq6WGk7kEZTF1oVcapUExOsNpzhimIDSWgap
83M65mo6e7SlVJZkSH+CyyjXf834scITPk+PZyXLcK48uuW7b9Wxpwh1RvR3TK+2
066p7pIPibot4g/ml7BUetbSURkXiO5AVEQNN4Oc5zlBbaIc2fywOEFry0cIYn2g
QlxWBDRqgKgdf5KNbe3/CttxgYg3bqQ3JrjBaqtwgFjpJrl8dXXPgJR9NuqgQpvh
pP9PK8eL018MQuOHTiDueUfST9oVxvAt6jgPyOc/4WkThwWpLdPpywQQEBsRMlrK
22KWKorkwD+aM4Bex6RdEtjBE5uSSACvgKqjd1aOGfumzGCEf3MMCphtH+WEbqCJ
xqO5UgWg1qMMGxl1zcXofv/MTddrKPbJ1BV2p4JMXe2Jj7vF/8WZ2xIJSZteSrXd
pU7BRMJR0U6uzrpaOQi1jlSbBN4Kmd4wz0TTKHCIE4ECL4i+ei+jOgWEGhHrgllA
hCLJwnNEUhoMsigwAcwoXBBAts+FrMJPTVl6fibDanI0gk/494phko1p4hwoUAzl
Inqgs1lBcxq5Tyw+/7AHneC5wfdXuLJMrPla4SpU/nhf8XNc3vmO9079EN4SaASn
oCyrxHeFChedD3OYTxzKynErvgjZpvuj7n2i3NdPVMCoz1ttyCRjEcPF7EsFDpok
qqKVnt3vVYTeXmiPpV0Mtf3XpI4ZPTOurzzLcnmKifilwJdNGKvHmWJA4jQpk3vk
qJ2Afs0+ePZieRX0G1gSm5JT8ZHLb6LSSe/tRCiEQZdGBZBAucB1cl4hbYOTIusz
bQ7zKlQ/ed8MQrkpfs3nov17EkL5Jy9I6JeSlBef7tnHNsPGcMtaG5q+ATnx19gC
fmuFELD3NWRFybfET6TC6TrC0CDpoaVNU4ui8nv9d3zMXQJtQ4W1noKmRAheDaBy
37EXlIl7LxzmMRsk6L7ku6NQ4hSjnBQapU994Wp7tC0ZilS1gZ26NvyhgZ4NvHVr
Pa5d7APdjZntsmsPu7UlZGh+fNt4RdVXSRB3h7D11EZXOiUOY08XXkCBbZeS/pj9
Nid7x5e0uThVvU/TaochXZ5DzBTEBVrjn7xIQ4uHa7aH8dQMdsezeClNFwY5K4O/
fwovrLWb6pn9phbjngF5/6ZSJJHj97RAc+X4A8s1DdgXiGvdrv3L5jnhhvAc7FOw
crTqZH4oaYj482cqteGQVyFnD2lt+q+euRpE00OgOdrirK3erVzu/YlXEZpGQKCh
pB5jgL5Zc+AGr1dMlQ6is606Eb46VewE/Quh9txbOWapmK4ZHsWQivRwqKwr/MEn
2Z2i4Wy9Mk+nCI0ncYb1NwG1jo+sdlvKuRQWQrwj/mSikrg0vEn58DbuNRlbcfzK
W+/zgj1s4m9abMWgUt/4j+C3jU3VisZ9d7msUPf1jXCA/u7cyoJV19cmjbEtRBpO
62i1Gk4fMbDzxQPkIHtn8mxZ1bsbwLrCHe2iZ6FWkvonYOb5THzCEZN6eTQSAUGA
XvboTO7z2msE2/WNYojI+wKsXP2Eq9tgsxvxGeEI0kTbUu+hAY5HjzEM2zd04LhL
bBZTp+7StiCQsdTQ60P/QAwSKXbRNlnSW72lEfWPQJ/fFIeYPieH7YPVGG3KIzCL
n8t0Lv0zdU3dlQHi3DzHZyFZ9HU/cAn1cVDdjeWjok8WxIc09aQuLINm7ftOeny6
5xd1S9W0WG2nL8+8X9Ys9fT9j2Bv7/FITcO0CIQJ4NyW272YpOvJZWLk1MeyNAAt
zlV3x91mVn2DNqwA/49HsLGBnWarl+eaHWojWtOewFd7nQvYecA4NCwlFPji41Qq
7CMAjBlgRpMYPno3wevJzQUJFhA2Es3JsreId3NjsoB46V1NPZkRFB5hxM5ZOtXd
nh9Gj7+8j69Yy9rrTBDFM0hVqsrp/NvdwEnHGupjqVpWW2WKUYfoay1y53Mf+8RF
FxuEX2/0m0igRJ2WAxgXQTVLfPTI2gUXhLhmHhhY/fg/BPNJGwRQ33WSlFTXA2b8
hHYDkHRU6431/WbPsoSWqisKqwkv+8/7nIwH5T4WQ84vwllVpcE6HNJ2d2OfTc8L
P6uEblHDS8KpuRbQJ3RI5RPUS3qXVRNXOGII1juAmQpOcx2Zs2W0qQlDGFkID9+d
XY6MTxXgXExSRuuOal8vmk7RTBQMsgBei75jZAYgk09i+06OTvXkmbZXmb+UTdEr
N4SoSBZi7PQy8onbIFKVHB4WJkEQYt0QDXSB9G34wNFnsUAwpr/jxC3cp81Zl0WG
fYRSKfKI1CAEOv1T0+R0HKaZs20BjBkNNG3yck0lqK8XEr2zUxN1TzjQvY4ZE4Yi
zReZwCSM3xJc0XYsj9he4LI16jdz4PA1xV6oygw8w/VkR9pIroKJyAf745RVJAqT
QyF0/Mpe3/+9X+4oPYCACRqK9fkHe22aKMinB7T8jpGtgjLmNFZFQjwtQiOwBld6
0m4jp6wS9ff7Gu725HseB0RUkBXVIsH9PNiUEegXnnvX4+mIaNpn+6kCqUkuHEhV
GCc37llsE0q7Qm9e4sj610mVPmesHNxY9In7LJde/ptLCQ7Xw2Yt+TkW9ocC83RI
ZoYkFcwoZa3ADp5yWV1NsZPRNkjSCGBRCNV1XKU2BhbIEBJ+ucg+syvGvZfVlV6S
GuZNrdncK4PqI6JSzCf2nCGfezyfZkZ3FPX/jdIIoXZV7NO+tPazRSC14nd/ASy8
SpQRAp13VZPGwMkCKWmwzJR44q8IgP3wY3AUwrM+F3ole1i5wrGpA+G+7e2SuIMi
5l8MLI8a9nc9bWtMtOHYNjFva4WnPaPeASli0b+N0i3bJN1njiUbPEE0g4LqfUY5
LLuE6ZZnTcV+OkYzQw8Jugs9iEkXD1mZxHcwscpBcAjJo2QqPdMWvvNBZ+iBNKU0
Vj51gfEOAITsVoDBderrmox2eXk8+9zp6j3Vr2Z/Dmv5hxKGylnFa85sEGSKrH8n
t4BwJ+nbnjf3lm0PgFfS/jjZwI2qQ/jzmHERBYOJbaP2MXU0X83WEtCrJKe76vrO
yYcCiN0YWGCP0b5er/6D2S+SAQ6ZyQ+Y1nE5J40aijnnjWKr5aUnj76a5bvgrpev
YQd/+WjKSZCCGlqlQCEepUgMiFPczoVbFmxtr7pWZIf/Ea0+qM5wmkglIjIhW2bJ
bZ5Vq3fG6xH8LsbofCTILAd7LcrTkeim8rLZt/QAOn4captF0nkjLvEjaQ3OATZj
S9RIFCkRs9i+8wsUm8aWcANK0RJv0r3rM3ztC2Pbd77B6HZL8rOuibkkgDhrUnn3
VvKP2Ca9V2Y3bHHA52zdriJ8HTnK7qRU5MBJ3wHff5+DHKohP7Cb4J5fV9AFGlJz
oBCfpRg8zHXVSGTvatDSONeUlZq4VkqZ8IQdquI6LLWSNxShlL7wmWXG9VXy44Od
+W2JVALXcgQB874QSYdaTg1JKlLX1BSTCtTB+hkjVa5COui6pZop7Fl0mdEFM1WU
ic7Q6xQZRYurADY+TovfLtZ34e4BFN3n1fSZwaFqY4AOCkNbTHFHfEUCFlJ3SEHi
MEL0jQv0iLnMLaS1L/zCwJ/abfs9PChzEjXa2zmXB6JKaGNwVt1B5BOs2ahBeD/F
6XINr6CjtRbMRAxOrgRJ876SBQH1HEtJiiGSEIzEijVvnvpuHwvHAoaPYLKMgfAB
d5lWWHRLNVlTWCY/f1ZlmVW+uBK6LniQLRqPHYPc292+Q5cBxKmxoMG8XaYE2+Zz
0MSY0j2zTHDp++ZP8lRl2AnQjR3lKkstgTm2O+WkpomC/CT9Zyrgm3IlereFFmJy
iInXBTRbQX7ovZmajScaDECQk8/DK9tnfocLMmsaiOvtbggUJiyfhASgNlgcmfbV
CfZW49+FAf85xlf0qdOClsjE3zE4PvJ2AhE1WYCKW7hTqdzk9TSGaZTzWH0M6dbJ
YEpVK+DWusHK9iXYERZOwu5VIu33ksRdMOGta7PRvUHYNRd2yWQSsxFe2hgy5oUu
wG6WCLFiDfPbp1hpLv9LdruaJZkNAGGxv38kJlbV1BKSwW0m7tTcB1H/2UX3LmCp
Y7W3sY5DrPk3fRKstbVMe+blI1FVsqRji5Kbxumk/eFpNorpcNR3t06EXd5zVGyx
N0hJVStOPfrIP/9hiIAcOyXwlWwFkV141/OH+LfClVeN9PvHZN5OXKDKD4ytfq6W
bbtz0pFnVhEEasot6wSuY9Xhm1GDJxIXioA1+0nY1aNO+sKeHik93BhA2N7VJwQq
jTiaIwqxGKspgIRliwOocqVrO3Lm/JFbHipfra6ZMUoCSB8jfz/ySExkORrZrEf5
nAcNEnPK6AAL8lVCm0zGPh/llW+Z47DqFVd0k7Z5wrrsD9KFZUsJPlqtDyNzH1B6
wvbVo4ouPOxCsGMq1lqjfGEZbLDLzpmYPAdhWpyMkHtqaGADgIh71+9mo4H3I/lh
m1QcIhxqPSHLV1HSOXrazxG1ih1VrKN6/vfDt1DllFxtIwarm9n80zdReHZPj02l
jJnNvK6OXk7q+kMSyozO5ATZHzzm03FofZUDMCwDn2U6YVhBLqeYmzSgAslfagqM
X2vnrIdbu8K3K4ZEUMhS3+RKlZCir45Jf9YHPoLRmJn5tSx4QLWx3q13mlqN4NDB
IHcka9dkO38xE/qCUClo3Op6jwwmS3OpHM+RyDdV21UOZj7+lbn9enUCcV/3y2fv
u7J1vs2BFYN+LHxbyXA9RhZhJWAN+NN2CFI3DH8ao6ns0ICik+v5QTIYNqquiCg9
6XDQd7hiql7GsTz/mgfADi6zph8zvF1XF4NkhA8n06QUIWedFBp76TUStx3YNdyu
lv4nPY/FrwJCjAXYj7T4zI/ZwcwRLZKwA/R+dgAB8PXIG6pZWfRHdNfZ6ihuN11s
VDGcvGvjHOzP3DOxGMHeCpcXTgPjaYsan4M1M8m73oA8pNl8CRwD0JcpxF9jetjc
g5bG7eXYFQbVmY7sbfK9LnwYBjmZrkRnCOlpE0tFd47w2K4+UQR+JdPz7GYh+bCM
dFkz5MjwJoJa88exgGgNgNav8daPIXl9y2T2m09uUbYUVgHMH0yg6OC6tzeDJYTg
bNwxV9K7+7BjffSJxfTRLy+7/yf4PRs7epdN2Wn/rElxKl9AU852BhA3v1RA1ZqW
j5A1j4T6xprZCKKV+allkm2/rePM+FACvAP44r0GYdIFy8HApA3IfptRrkVoXiQj
ICcedOI/mn2/Hlh+vfupquCg8CwI6dWdCUurIMOyoYwww4q5YjH/Q7w6eUGSgbQF
U3IYHsvddOoBqe3zJVRnSN6KJKOcqXl7BD9pRRbUsEP14L6RDkhYj+2yLN0Vk7ng
LtGhh0PodYRificRgYVYXCC7APpbZVplDX7Bo1nG52SxjQo2Nj9aUtLpJ7Jr2Jzb
nkQ+p1bruwYEz+v/WQI+rrcvwUp1ZIGNYP1iWunnfZiL/4UE71A0JjxxC1vrX9GN
GQ8Ac2i4lAM8/Q/CIbdf7fwDbWPOYJ5oVvUdOOjpvu0Hu2I+i2ArKr+RDg5PWyTa
cwFkWeiw7C3bHSETBVRx89J6Z3Q2tbmBMn6HUJZXRrCg7pg/ylRnEwzSfxigCyuM
kxpeqM9zhqm/ZXxrsamfN0oWfoYyK5y/IrhobGq7Hh0uoQCaeoReFdKUPbzaOT1w
wd3f9xs/LnGxHscaqNp4dgXQpKll0luHg6f2sBFpsrim5/qAhKRCdUQZ02vAv0z7
CHQ5j2aUexSSZhiFEC/RXbcBgTjdEiz/Z9Om4Dm6XJfmQaJPqi5Uz6U7X8+Mbr0A
HbG4X9EZjuRTi+57ruvGYKZTxYfWr24QYgZ31ecHh8YA72NaxjPKmvqqZmkqcms3
ZlMB5Q4XtgtlF5dZEDAxuq8lQWulzq7mCKKumYb95i4D9/19IHNjo/2lw2TXWDnk
9gBdmwp0Avy1q6yPRe3bPgyQ2KD7zQqXmjcjts7uVq0xN/H7CwquGgJcaDM2Tegf
b3+6aT4rvg23mhZCKbKs5j+q5/GO4UJ46+TKZNmN8Wnv6V/HgoEKtiCjWFoHuaK6
VRXO7C8peOi9wtfAj4LqWT+VbqTqfZy951b5GgSYz5Ra+gVQwqnakWkLvnOpjOPh
wSm9f8xksS2fqphP/wh9rOzZah+2DS8JQUA6QT1fOoIRN2nJVlXjnni+qDrEVYiz
0aDoR4Vaor94YRzwr+4MKJHc7Gx6gjJ5LzBOaBoXiXcAI8E4sPmmnPfUTIRzrx0l
5qBJgHbxPYxQaZ8nsFvjXkOErmu9Y8sBmoheuSbUvqXmxkLnL/RF0fp3+jgsU/pQ
ob4iNUb+aWwJgdpbLrCXYcA8Gp2sUvTqgE7hcpeOt5lJn8KMz1EVB6TFBq02xN0+
okYqFz3nZWu0wdkKUapYPTu8JTJhiuKGpyOiPTUaiQOGP9Wk/91QENgIx5v5BjUh
o5dPgGGRKCiBa/PyA55tIILNPyCU+JZ22hznz4rja+M654ByKtL9ZP7Au8HvIUpG
754l41AnedsrVUVAcy33lToYvFFAQE9odEt7reizgn5bhZOkALcdVogeKAwhDEgL
wU97oPZVHXsi16b/eviiJ6ZnXMhk17Y4FWYtmNNdom2DUEBlcOq8kbumrGyme1uD
pM4kEP+HNkuQDAcMFmJkb9XgvTDViFHMvPXUopEjJoKnCOVNnuJt45kO11yDjjkz
M4CkKA0K80p65Dv9F3ewRb/6zjRHcL5TuX0YJ4uhalX5mW4au8FQj6udqauILwh/
8dSFbYkmkK0d3iF7NbXTW/2FCddvcFWuX/DKZ18dJyILji5Ih2B3Y+5AfB0WrDoM
iMntMCCzlE9c6qxF42VRASsuPaiTIf7BSI9oG3EmXWmSsI+YHQm25JxrlSSJ9mmg
U16retPL9l/YJjT2LEGoSqarVxYgGC76tjPeMnC2l1f0UjfVnIk7e9aBr+HGOfVB
4T9W3gKhv0stPbueLrLGLMyIloHYvA2h3pYQofaBjsrIVIfVc5lTfTiMqAv5mlLm
qbeqFWvp1ZpIsA1LBL81cWiUqbZZRrT9BlDbIrbKbrkI+rad5d0+vw9SZSU4V6xk
p5kWUg9ItimYErwt28syThKVISBJbdiS/2nz9oPoB6UYIrUVBuGnM3qoYwz8Oq+h
LFE6OTiC5Fp3wgziYRjiz4N22ppUhltrgTjYxae0zKGDF2PSe/yj4z3e8YWw1ODQ
MTbMxvz0KraFFDZkqJersXoyTj07ToM0WmuDEbFzMyX8zo79tmHEZFBAFMyqAouj
qXlJWL3rDbhFW+ABg73SdaenoWrS3fERAK5y4Vw5YnLINQxi2o+to0NFLFCqU2Yg
snIMvM3Vi60/TrFyn4+zO25gTMoScBZE3f3P/+ItF6FAt4HzV1AxlzfLubgIlsUH
5GCoyLblxvKiRByo1JULZrXtVOPxyr76eNTUypn19oTfAWQcdmyAcsN5zABe7Ox7
SdvzE+XNvUljsKgOZpus71C9v+i3+9+MoMoBmaESK7BS+G6KOXW5aD317ICHyO/C
4aOrYlI/En3ec07VcUhKrYycGklvknmV1/p3zcV41qafyMEiBqoYglnelWbAZknW
KaOE1KW5gQi5KDLUvNpS3h+q/C5aMDBpxc31ATniHTSfxPyJteJ2VkhTDjKO+IHR
zAy+yOCb3Le4hL85Dd4EmsZObyl67E1kX6z5quUD7TNPXMtKNXyDpXZ7YHiemPIm
yIuvtUCJj7Cmvhl1SdnI5PWVPojMRIj7mzA7ifggdP2+BDqbGmvoKbOUvAD1J1h7
dZ5BaOJcPjuiWmHcGyE2578RiKSuhiwTqWdr6uB1UrDg0ZP/kgImgiI4uix4mRIA
vp7EPPBgxEc1VAPMboCQG1LRmq3AvK6O4cmdAQ1ptgOlM2JyHLpzzvE+ufMb1i2o
i/Mc41A7xtqUZaoMqOcVDo7Ye33bbgnHD8hX/k0N7TU553gFZtYRM8ATht/9K91N
D1J86lFHpOePLdlPjlczv3/uPZqLy7qJ8SOvcRenzG5iLg87fuHI9dNndmYH+ab4
gKpa+pmSRBX7Zy5S80XeyYcv1rIs/+PadNHJqP3QGX0/bbxPM7/tc7seEYvHMPYU
e7ClJeD5yvsyXBJrse3aGUaJZhrWgwSBs5sR69dfbt5VTKiKJlo2QU9AQZksde3Q
LSGRLecmeXnApoc8PesHWEvKqaa/iMx2+cTplqSw9MP6HdD4x+tRaW4FyBKnk4kG
TxqaIpOzlAed0/pix5UaVZTm4znmb0x32t+0dHfUX1Bq/STghA5R56cckzlL/8As
3gkp9XIs9RN2OMZ2zGZ/c7GNIKbZqJr3ETBG/qOWoCE5fLg4ziQ5WeHCLf0rd8bb
Rr9EUwSUU0BIHfSjaj0XczWqb9ajmY27hTIH7AyGouHeuTVvsvbAycuD9mGEmaTr
pjEGbG3DIpPfgpnDlWiXGPPWiza7ayAVz+/pd/5iUwJ0hT55orJdA6ep2uQfg4am
rTgR+6Z8HoBpmT5/C7Mmw4EkxJcFJ0VGi+JrIEPOGgdbLh7GHIcApeL7kC6d/7IP
CuxZ58Av5NhheR4k2qVnaQXJtALZdMdKOY7ukFaIW4iSPYrZLYIHbhxhCx3axsMb
E2hyBzFRI5a75caulDAWgs55zVoaXW0aRnjDjyjTJZTTyUrggC0rCHaliYuNdQjv
X0t3qMZ58j/Mv+8kmz1SP3v0YUhFMOBJSMoSk4GkmWkO52Ne8QdmLHLNdw0jQCaD
IgHj04dN7+OSUWKwLEragGuoPUuQU2qjtZRStSrh1pnUwYQwUC7tmx87XskwiLkC
sEAAKFYkaAQwo3PFgIHOTWnch3d+BH6Pp1rKKMSc6XJXyAOoJz6FdfAAOdudn42g
1TUaacTj5gkRtJeqc7sPIcDnaTa05pA2tazItvV55IwH1ifYrj2eTDH84vB09d7u
eOyS8gp6eDH1NwWNmRDiUWhKVqb/bqnudRpnVYA4rdPxvbXgbG7w/g4Z/oFjFxu/
RtlO5H/UfHEDSHXdqc3fGJnchZuUplJCEXzbUaD8Ij0s1B68Ly7fkwd4T6CByYPz
X/PwHTP6vZYovGkmDvYCYretTFD4P0pw7bRHEltXlNzP/yHKXRJwGs7y6b6rSwjh
sc+lMsyDZIppALuEwpifdGsXsvq9p8SEMmzwrqszic6RB4jrUoH0evTOj+h89kLP
0y+5MJHINFb5QuflTbXRyFpm441geM6zrVzlXUn+m2S40NVXbvj41Ks6Cl/I9vQU
aGDzfxHF3BFqrpRHaWhZhkqbcgemtc63DNoCCqbSPPaQYwxcBkSaU03dYX5kIW7Z
WabtWIAXswaoxi0icYvnw2WLr7vLb8g6KTbCfUUbNICsc7sInddqDmvqDYMXMWwn
ndTHWqsm61a1493qBsXO4S/SmjCbAnYw+waAY9/NQni+5zZkok2rq6uMuNKzNNId
0qzhijM6OxepXDzMZ/MEx4QuT3Un6D7lr+Ru5WX86CNdVqiY2fGCKq7x0ZHbqpV9
E2hwketJjyJkGvS64vdB9kCC8XuIA0y8rfN/k5zt1PxJEsx21iZ/UBQhblqRUp+A
BNdKBAO3VWaSEYgDM8vylIdKcjC+kCoclxHx3+C0DbLJKJcC0MM/nS3C1FCqnAvf
VIIoZDuyOwsDotTTikqIbLOiahMhmQteEK9jpMDoQclkOS8X3kmPf0QJj9XogO09
kLBufYKi0eJI/X3IqkeG5RK6Hx5O2fSBNDzh6n4jQ81kublaruCTUGcxcVxBj4Om
GU6kTHTd/70rZQQYeYmTDdcbmr5LIFHmmYst6ijOPuJSO4CjJ3uZbfHqWiCwLI03
oSzEEJ7yDEdBwZbP//yUsI54xkfKbKEQQs71nuTwEBxcDAgHuyO/6Ku7tP2h1TkZ
NsZ2/Csv+P3GaC3I3qHLyDjP5xit5lwvN6kbX6chCZy6o1s7riuhHdbTeLKHho8J
YK8YaegMzqhQ4ZucPimiWXBpeBS5hcI4k58TKZXlMSQ287MHx45Z3uYF6GM1rZLq
HZIvKiujp+bg9v00+NS2Jq8+PD7cNBL6Dw0cD9pvh6DixoN2/020E/KX3dDmpmh3
tYXrLxujPweuvld4u2TvtvNcJeBupcyZPF++VJ74PCpyMmIw+mStCiIfSTIlyeQl
UgNlXBrnczErvWIZDhoOda79CVAanDAkSQNYGA6EnHznUU+IhoxgwiShlRXFY9/9
saJq1om+6+io90Fi4mo8PLQUaEDMLHB1pjwPJljaMBcRbmChr41ypAhBVxunx8Fs
rVKFm9xWU7LGozP9/2vu+/VdWaAsiQgEUE3QpPdhxJdZR9qNNeFrDYGxQxSJTDN2
vfgm6JP1N/z0n/Fk9X4JhtAwdc8r6zOur9UM7ZSRBpVVBnDVOZFaPUg/aRYOZ4rW
yTiebMcuIFZMS45coy0vw/9MAyAUGKOqs/1C+7rEeidIloeyK+h/Llz7g+lJ5dDO
fDHKyDFTEk7F27uQCR9KIghBlTBT6+ToPddFPntZcB8rd1Jr7Lpo/VZRc730RECD
XCTGYiZl0f15REtDh4MP1i9jNepDeOHyeeTE7kVXzUEUQYwMUalTeXmjde1x04lH
5Pz95wKnZV2eKEwrXU7scWTcG+Lsf6crv+KSUKwVcinHaZV0Ka/N1hlcJHP0P3hJ
EJf0WSB1049YJncsPFAdoQ+GXj4VmJqOVUhj1ixVA9HMQbXEcx8bT6xaXf0rtYYL
zHcqjD7/WURyWxeHfM9AcKdloU4ogAX0pOfexvB9hwTXDg9WG59CkVVP8i+2yidr
4oxg3R076ZM4sVAHXjSk+Sm27rMOweVNUyvlDsXZDO4SyK9p4RoB171PzUTiPmjt
X8SODPcVuWaTaMNMjsC2KS41iuvfwm71RWzyr0/IhbvcD71usPrg7oGq220fZMdN
7Q7gP2j+8DWYPHzQaWaQL4/og1igMBg/fu0pPw1d8kiSJtRNl1/G+F6LWwJV7Wo9
MjAWL5QHaiE5lBb+Lsa04YdzlBmflNZLRCibBI9+YbH1MUOAEttd5KCcJZ5izPhV
fNj3d64mjgJRg0g05fPlHf/9jAQNxZoMVfCtM8RDdJA+pi/5VQSyYg+jKtybBdlU
MPgdd359+RrINmMw/Yu/mFjV9KH4XGuwHgmFY/EC36Ipa5TSw2ITP+W+aSbsIba0
r0BxbKuwfltQeitUXAxXaZJ7pAhG2WIB6X/VxQ8TgvDO5tg52Qi8iHW0/og7FbJ/
rrRlZBzsj/MSezqmzmdf+JmkZJWnQw1wsvY0TJnDsF0sJRXN98+PKu/HCNxsVn3a
TPLRj8dnYTI3Nv/Ay9yQRA7Mz1bsOLbK3dSBmsTwk4OOYIH1eGRGDzw1a7IBLfDU
Vvfe+8am0gU7YLOYcHexVmQjMknI6xrXOokX4XXB27qAcY5r5hEcWkh1eGJjxP8C
3jgrQswj7H0zZbpnrVXJ//zNL4xwPC83P0hbg5cNLkcKTFj/pCaHOFkbBG6U9qs3
3jo6/zKKQPOn6jV4mj5vtl/X2qdn91H8rwgNtQlXPm9Om2/UHEKIjWByU6jn3tqb
xO5evTlGfBbiZAxclxCtGMNyd5Fv/tMpcsVGDYirVCuLJeyM5Wascf9sMulZclGt
RV7QxQR0lpTpvJKOOQUWRxKf0sp8foit/ysRUE73dQXP7YvXIBvaab4F9qVcV7qk
TEmWSWGAt0VymgL/fpIAo8h9hjOYCtvcYo4PtmxHlcZdUF/XQlTziq/5JOzD1mKD
MIKuFMGmwoo6Co4wobqy4lannBHyXQwtviCIWqxXTeW3TfDDi5AwIk6Dats6lW9k
IAwlo1owrLcOXvD5YcG860Nn3Ttp0Eekw7eC7yIp9oact5IGxsGzFbTR7utpyG0W
uiamsVCFzip/lQFl8otgD3Z3zEpSQpk/dPLAy1qc61edzD5w+Wj3GpCyVzEBpm/n
22X6V/YcjVdgFae02JXfC3QGQb9OOueEMZpC0t2YJeYiKsUjRIv8bd6SC020pKYL
x8IH4ju8wCCGqyufTHjHrTdjPp8p0YIVUkk9wz4QbCyPSZlE1qooO0mob5/tOS3Z
1QTl64lKVYA8HyAt+QKIOzmJqqOjee80/ICpIZJ+h06hHW1hLdR+jDx1wj5YTNnM
Y76VCqPe24gyx6/iTcKm+uICrKC9bW55+m6lCrOo1gN9lB+VhLVteWQH290E4kju
6fBK1UtlJJ7xJ/5/6ZX44nkwE+VIpbE6416mghcnQgSSfEv3PChaPaO9fh43b7XD
5VWLHChxEuAXMtsD8tm9/Db/tyLSk2zze43T+tRltq4ect9bRa2GcUABVsKlJhzO
bzkHAhMAWMviKdeyV6lSs2YckS8KGHt5VxarFTLEevD/TmvS6xjep70rKAYEj2/F
gFCS3ncFjXc/GvDsU4ZoB/OGw4H8WcPiFW6IcljQHVRJTae27FzWnXLRLLqygGiH
RbPB5XEqJCpsYdVavgXX1LArKhNnwOL0KIT3dfBQCi1nwOrpZ9WF09Cx0j3qbA7J
smkljuSfbpsm63byUnPYSVSUIbjT/fUuwA1DotIC0auPeDdZZ6GUHyfoSgQGz8KT
jVxkRvtNL55plXGNOukxaVl8ehplLw3jYiNan4Oo5tqIYZkiw97en2cP3WJhihws
6rkV4Tf2DAXIIvbvk20QD290jOQ8fgKS6cGgFLU+0ECdUd9gzydaAEnxUw12Bivz
FVwEJr94oV7XGWyM1T5XWO8D7R+KloauuJJfsO+GV8XR3xcpvmojDdFcJuqIZ2JW
KNP8BSjQUedLGQ7uzm+1S01GtW4ZuoWnMVhIs3oGjMAwoJr07Dmg623KrjuCS3eA
RgOWxabL7M2Tgrw55XMmgJdY4ge3jFrSZe2KPCxfyTEvKJiQH8EjmgKl1p7zx9Hq
hpTBoJ7vKdH+KHWAis/NBj81zYys6yS+PQbhQtzIG6dLdif9t27iDWn/uD+hsnZw
KV/+o44uxUG2uuOKXNXIPb7VdXUAwzYuIIU+o04HIBU0VX4nZRyVqW/1dRy4dl5a
h+IzrWAjA8ea4IMJpaBSeAJhVK/Z29BfrR2/C3+YVM81J3Vz8FOHGQ7CHB4boFAc
2eBZvImfMeFmhFnCTeHmuG7sKzPKV/zW/WDdh303CskyMc472lK+XZ6eoQhue9Jv
E/47QsctoI+0QRsIyL74Gc1DvChCdU86rilQIzAOUwhoSvt7dzjuQQut1BLtpoDz
kAR6OyqAwf5vJVhZPj9isr+WRBfk3eqt8glgZrZiJMORtssOujO3L41H5wUnZv1a
vyz+h6ey1V6HMquYsapR3ESYXpDzhGzsnW1ftK0yHktRUAKOqy3G24Qi6RCtP7jZ
RRYmiJGIEWWFejB3WY3qGsi4ssiYMiCrf4JXBSFUZHQE9TrNQccAlp2BtEifDHHY
bW0vvsY8gQpO4hjdBhvBaWGPN/G3A61btgi1SrW4b75Fb/9aHvJr2sQj6d86lfnr
AK6A425YfNkGrjddmeabpgcblSaMsBzSqvZBPL8+aLlHNbm+avm3+AC12sqAG1xr
Kbe6DdYDCo3+vBropS+KlvDqGSlrVDr26MPJOyXeHpl7NhhRc3vww6xS/7HDPVOF
OGcntOYzS4yl/L9JhcZD3582iYZoG0Rd0UiBTeSe0U/uHpRDZI0pnBOaYqqPvUgS
fRkISLDolkGbbov47xLQ462zqfdF7ifPelWil/fTLwAE2/WbRmiRd9YnrFlpao0D
NHwUr8ZlDZivZ2KLXiBj6+tIzX0T/tMoNJ0CaKm95NRuGa3IvvJFf3aA70gYel8o
ZsUA0rXPxg0ytZyj2ny5UYc3iKWUsafguJ+Qv4viNTCfIWCWh76WG4gphlS9KIU4
3UIOZq86BzTO6D6Olu6kfQuOFt791RYCGjoah5nWDAvPFftv1GVKYvUnnbwjxcc3
Xz3kIKleuq1SZ9kQN38j0jweG+VnqABloLboOoxhnjraOD3ce+KQsEmuSwLgAX85
Gb6MHDb5GegQVRMvfNq/wwj4mOlVkoHlfOctD5BEnhyJBn8NLeX9RV6EocmZYp3o
qOuHYE7GHmbwokv5hu72TSaiEG8Jy+eau1VyDl/R6+018UDZVrl5ZWNHSHH8/Ki7
tzsu30rs63USMZDJfqA35Wq4FWblhM2GEqL3ja/M3dzR1yfaqwH9+wJ1Z43w1RXh
HmdYFPYydADIdPkNnS2G3/Wv26vmOPkEaTzI+LfpV9G8R4cxt8vvkJOd6iEIGJRT
SuFczgfyZ9mHFCeWGv6UF/U57QbUwCpKC549FMX/E4qYQq7IKOrGhkDRKSMhhT2g
ENdSUW/OkhFa8mEGTdlcXYw3wxJXAqeLC4fQaitvtiatOLw2xhyapUfbM1r9LHyE
T7KVCsib8+jbwBJFjc5d8PUhx6TbRMcTsf2h9zGyBWUQs5wN3973Ncs+RLs3SU2x
/1xZJMomrnzx8bEXrJJBnM3xUD7K81v1SagrL+cNf3iGOvumRaZhTBAzmIj+ydLO
4zPoloX1pn6UlxKRPWo67W9HwO5e0vygSZP1vvD90q947UIONXRkH6hi0P6Z0yU/
4rMnsmPOlAcriOcQsv+3kkb5DXLYvB/CgRbjO3HpbwSzaHPD3q3O9WgQQym75CQd
/sXmOk+Dzv1wS+wltb4Wo0tMpo/6sdRuJWYG1KRPjKoOzbtuaAjPvCuwuqRdA99u
odioxH3FbrMgvDfvZORBAp8j6uqWpKiY+RcSSsde9iki3bt44w+MVpzthpOkPFH9
AoLp8DA70S/lXRwlB8wrSRDhIIIvWLzIOuQOPgU06zSYo+K3AiKPC41/o+azIpDo
ulqgrGxMQOql6MOXadMoAHUp2pXkHiJN7cT0/nEmdGIThkybRbiPT8i1wjvHIWoW
+axq3sMxqDONtrc6etFWhKcves18tT7UPxlEhFyXf9hrMItoJGIFJrdjncIBOF83
zKbzBuWkZyf0IPxCfZa/NNZSi/3gxXLjPiIMz57issrcV+5DmaSijKsT8E0NylSI
ROoLVoZDNARvUmadLI6tPrdsqqVdbK8Ht5BowcWHMNvsM336RdW+vHPqOCO2JOWs
/p6Aw3kUXOtZG3O0VgBWLJrZQdQxCXCW4+xWrJqDsbGtRNb7IptF1bJ+bvx4G0Kf
qgEeYCyGHn2OEQfnmrd6kY4pI6lPsbM9TcmftVFmIsc/UH68pChsXzoE/pciTMHn
za9Xxints8O5Bh9Fu51oPND/TwO3WtKRfcUFDLFDBIZunrdd3ESedZEaeDRvDjTk
PYOqDJCQjj/Q/zHnuxWj63k2drS3PVH3rmXe3CG1s81tk5oQVVwnRWqcwm148/CA
wiSSdU5uSxyUq89Y35KYXEsMEXCkkaCioR0pbeNODWiKHKICt/YushVA6m0Da62W
FYEcY7rD4knN3PE6Pjq6Y2NTAtNw+9jsqvUHFkf7+lC6mesn6WD6DEW4xh/fABhe
wnLTcFPi5xgU9wcXcUJKIAmuST4Y1TpvLJWq9v5/DnFPTyGwKjoRrtCK6sicKBkr
d9rWsKjOx5HNjDQiuWE/KYUTxHTILnCBI7CPPUersrXigmHrbGtrRYKon/WW1aXb
Zy3Q3rr1Ka8yPNoYx8U1j8+hRYitYLEIylBMk2+tzsXJFeuMMZqZtb8dEib3mzAw
Q+B0uIpH2CqKR/04CPpH80zo/KBiNHxI7cTjlJ5Ic9NJWbVwPKOT/XBirXTQsLsB
lQNvSif/VYGZeQIxKrUYsgv1ENBhpoOCTTrx2JHXlLwy6rO9/KFN2SawWtSQVZJX
fKHbxeLOkbU7kmNlTTACKbamnpv6gqFTn7cznQCigjty27WJGjBkbSIQJ0Q7DBz/
HmaKRiNFbkEkeFEh8H7uOMGrY0+oKPuAlpGUZNsKTrIb101MXfrjRY6uizu3wxTz
3gYB5FUbzp79pSyah8AvWfS2dznt9LVmqT6rolk1tQcsn82cO2TqAYc36zQ7eTUn
gDImXjtuRbe1OfLyMsN8Z5kwv6/9ixt3OpIHsZaHTRchGgPufkF/Avpb7o/SpERt
CuOxegjQoOhzCVi0xsdFCKtls9ToCBGJNexHuXHLoruNLkY/hhHfuxW5YaKc3nDm
Hk+wD1OjHMrGkLbkNp79diHy9xQWMN5QSRW3csi3LYHBBRfETS80hfxXhEtPgnck
cTYav2qVi4R1CFnAHibbl8GNXS3RmhazwjXKfLv+rwh1HGDhKGK5VK6W9VqagiPn
uIjwaEyANuM0G4WlwkLMMRZ2Fnna6lOUsiS8/Gm/ARBpKKW7KiVJ6o3roWnhhiYZ
MdumsxD45dXAhIf5fKTP+cjCzZwWJZ4+KwH5/3Nae3BlblbrfrRFOPSKj2AF1/5g
Lulqh7xW5g8ovV7o3WSToRFB6EpR6LMd2BeTB0wSxZ/lZYMed8TZ4jl0D1WBIQ4s
U5yV56Cr4aa4di9aWpfxCaUUN6fxIJAKb/oPZ19ZRZS679nv+Jt/gtr/TsjLBHYr
3tcufg88guh/w9mGTtPe4o0kUVTGhuLgi/0bzVARzfKm0FCQ+E7iwvk2sP3nHUFj
8ZPdvs8A96yCzvXkyw0kSkYsLxgtu/73IG3BfIs3+Hmw0rP3nM86CAzm9Z8tNdR0
GjQm7f3iIBkuIPLTejDbCuWsGM1l3IjLwu9JgSoMaHsPKwJZ37oUMqKtLfrLVqZI
/hy7LZNgXGnPgN+y2vBmRE2DJt7CXBO8swVBh5UkzEcpQP5XqsjHNItJUeUMLMOj
bt9hoF5xg4332lkiReMk9XPnfSxEhbm4iiIrTwluQIjRpBEgifkNiuxMvvmcLm2T
Y+Q41/17KB5G+TIbYjNg+8iFYBceA8s0fzZ1sKZyStCxqI6xIsRAGmRMfDb+kE24
WL3WHvu0oEiBoXdF1ol8//j3/OnLeHgfrI3OysdXAqaRtrPUJygx+ZtfyGiDjtat
uMh3eSzfA+7N6RG+u+KqX2hgV+wnYQ1m44qfyVx4mGDXXNTIm2D+2+NtSW47RT8C
27HiE02ElwwFZXq5pEAgfkeV+sEc8lRhBExTUzZVys9eMkBNnuxwyrB+UVxPBrRb
7GZa5BUG5t90SFzF0igpTOMSyxutcUaRBwkSHlKheuS/BsFxzdYuBrZBnd5yc2Ce
ZTpPuWiBWZ8gEQO6mQgskwG6SS4J20jUAAXP7Q7dtL55S00ml0qnGV4bew5Lx+ec
A5B24JNYLCJRIYm+zPKjtb+S4s2Rhbdqp6MSdXff8okKb1NSzX7VBx1k4809EQdp
EnHf9r9Le5MAyw8s7pgpcmpLNh7phlTOz9f1Qw+aGRLnVQGByROBtE12HCK0GMSd
3s/+2cgrifEAlA1KC3EPm5hbnti8qjCevONQxpVnL0Tz+eFzLIgfSq1pSJfXd7Z7
jve/wy3NTk3p7p2ahFjEaRiZdgQy4X8lQMr2brbM167181gUnPT2ejA6ZeETa9JA
D3r74VCb+8pjkISOD5NdmRCuQwXFpA0sBHf2zM760eCcEmooh2202VdkrTQPJMga
YULOPUVEmOh0PBTuc3x/nmIiYuhVqvDJqPzpR3fTCk4XELhWKC3bFa6kv5AIuYju
Rhu4l9brPiVr0Jmlh/d38ZiwRWFK4mERSrrD6kFuO/SSOqJoNdYI0niuebEmwRnF
ftL+nDPrHO7vaOeEXAZBUMmFW5MPW7HLjRy60wTBp+tImlGDvSizAPQsZH7AivDI
MnTIEQEdBlWJYbDbfWpzancygKfOLaT6zQnDCjgj7TDEptUvvu1XDfbeESVOGnVX
X64OTV0Ub4A3S7Pbf8lkfJB4AulGDRqrjaGorCGtF6SRKZsSHqQz2Bo5DY9QJ0L3
g11bBc2D0Xo47iqtDt7R6DhI2+xCjRRBSqxwku8Uf9JyNHgpZnVhlZKmhbVgVU09
4Xisf4znT4ERCuHIZTEghCX/NcMp/MG+CuHgZyjL80HU6kgZ9doLTOxoHq86mkiZ
qSWjHoABaixpglODdu24Uf0Yj5ExzzFGnK7LmKnaqvgP6E538U2R8D/4QyvEDtXJ
V8f2VvYq9xdKIOU/HTPBIpGWjtU36yS+N9xoH/KJHLeiaYzj5OxtD4y9VlwDrCz7
VACx3LoYzTSvrkFdsxitUSP/zHgi+Z7Q/e5MEB4pmXxP0NhBv1tym56ITBwYo8sl
x8M7eN0X1g2AManF+aoNvhKGzdl8LWRg2NTTCYmD1a6kww8whn3IBpNRhbIKOxYt
HxhP6+TVKil35pNtoGqHzHIskxn2mfQqQkJGmm90mzorngjIRmKRo8J5hKqlcQML
IhZpvGMYG3/TYJ/1Qc2399G0GU4ehRUQAeSXfKviN2d4/ZkWhfVmjcxmkxHTE5+E
66YuNmqRLW3ZX35B/RN9aZ/9tgsD3JTV+yJ5Sajiel8IVFCa4Jr8zdQU7L/ES+ci
AW8j9itf0p2K5V19YLpwmQQQgxT7MyKgqeyHysUTQ3IU80W7bYDFou1ABcXe2H3e
OfjEf8OmBnJnPHWqvufzz8qvY8y3PvGaVi7M5SPL2A46LybG3V6LjcDJ2Wh8Umbu
eKBwJymj1ski7CUv2LWh6s+Hp8fwJxvAvFk5Ya/arcS0kMvBImIYliLatnlwWc1v
9nxvj2jM3bYXUvGcg8tNmf8Zox0XKUCM8PeJoXvQOSzRQSI6SReOO4hiv1k6kbZ+
4R+74HmnG78c5qxQJXo/kv16jpfo9jSCA1JMfC2QspuPeZGdif17YCMVDia/monU
B9opRsSK5EEZuK0aGsQ3hmf9v9z0PxcNP91JpdSv4+dwIt+X8KWG0BgQAeNlVT3h
Qkh7ZBvz04n6jHM23uMr3PKKZynArHkc657XW41v/yjQSCEXNzPFSTFnitD1AUNK
uARbJyJgHVBg4qi0NLm29evostE5BlYST5ybl4Tl5RAZo5IMX3/Fs0MzaHkmgJCU
bm8Ia9eAtvzx3TFLI5+djrtKix13A4KqVGLUV20akYly7y8SKVwMfCrFXLBnv4Fy
Y2vxXdN6l3OyzVlVp6RmtD3vsRUK67QriI6gc3wqs2CZtK325Utz2a+2KJQJpOut
LzYroXR5bNTOsiHgwtDMfBACgZoM0dtUtjjZWebW8OnFu+uDvanb5NXA9qem3dMU
CklSaSDtUVh+pQgghHv0WBAP3T8lQ2JuzGG/+s/GzTUjgCIv1cK32eizdM8S/mAC
WlXEDlypxFQZf9Gg2fO77qRA4gPHAL7Ww3GHdRBkT0RS1rqZbhmNJhhyhPTOps9k
tlKM3nvRwa4uGj3DHQTbDzlGmnfwLkfxgItezewug8DzBmmq4dKIzL5QncE9P2kL
TXxQFnm+MJr58wRNlS0Q4FDu2Mv3zV+QG6hvnHFcSayTsOxjbiIBtepAS67Nbi0/
XE6HpkLyU1ighwRYCZovFSXavdFzg4zZ1OMLmwM2IkrZCIIE5zVJFPI8t3puaDqJ
mLhQA3yxhDJTWnkZe34pK4ov9bdIe8O7rQ2H9vC+1KZD25jg3CaCOzfs9d8/SaFt
UTkroZHZqNItZOgkrEgNG284vYeEeXxOV/ePrwxs4elUiZJE7AMEXiE+YZizorxq
AanMkwjbk28lNknSFXDr6kLMmAfsZKyWBEJX1vAnu/aV8jSH56bqr5RXaucAPTYt
tx7xRKZ+TQBwR7q2Zlp4x6g2/MJWoqSkLqxuLbR/1M5JwmXxCYsk3TsqxCgHYCrC
oxl5vjfkubHASlE9M+08gzRD4We+ln88fldCwxyVoeRhoLvfNiYl9ct+DM4/7S2+
czVkMMOwh3CJTQdmGLBD1C0BvyO7MQ+wqBH4Y40PUmxKzQdVidJaK4KAuDMTr487
5XXueX4+OHpHEY0pXyCiz5P9Wm6dSwaWyKFpntG7UsJs/0rbVm6b4fb04+ihQfYp
pCKJtH0xbFQJJOx9ETXAFneHCpQ9JsjIMrSA8mfxLlC9RZm4tIPDVb3w6uz5yrNe
tQPfVKdMCAIlDrJLDjYtredELyni7iWiPXIeNgiv8qzBdGEjpFZUDXUiudeKorH0
7dKRm3fwhsnASrqjKgRWcv7SmQVXPYsKD1IbdqvxoPIM/K1OmhshvCC7/oDQY2Wu
v+Mdrfn9108mKR9t3dbKj+92RgUNuPEql+/aPTxUbJscTdgDTpI3Uv+YG+xWb3eB
Rfgvhsr2HZVwlr7yh6uRgt2scgLjY5eQc8TqdIU0Dbj9AvpdvE+fp+q6Cd4eTmDi
9EE+YV1ExUnG5U4Vd7YJXpZrGUWDxDtA8pb34SSVeOeOv1qe9s2oeyQNWHaucFt6
MECnPX+RhJt+yGGfeGyj6Tmflz7sPjA0yPzZwCBv4D4uQNj3A4oqs9a7FGYHGKD/
jrNLzkA1bbah+TYJS+eI1cJpKPoc+bk642crC68bg04+OO5iTzWSjyBfKZV4cSZH
Rmr2RFSHN+vlnflVJsXetUOqjg8vPhBvael3yrzDNN5JZ7f5mzm8+CqEmJnLg01z
NXTGm6D0GszNbP8nWTTXWKXKoPugqYc06j9GRw9iU/6Vi1n+LcKbpaxg+hBBEhYx
IUFwD3xqe90O4lbWhAnJzd4ie5i5Y5sSMwLWE8YKbvDPT9xBro/TQgyMLBsC4j5J
ZE/BxSi5BalEs07AQSPVJrXTlYM4dmwOPi5NYcpvIKXpVuLPgvqiIYKr5mISiLsO
H588+matJkUNzOherNIbzaWScYOvfBaTNsmU2Q902nV7XFCEstyDsXiyYAOQUwC2
JmOUqeF87idAp9UJXA08x31QJNEzjNvB2cSVx5myeFN0h5WRyIm5V2o0HParh4hj
MBaozQF/XJsd34TSvf6afVxPOaxDKzdWJqVBWX5EEKbCCVRJVZ55/4E54BTxsy7X
S8jCgESbEAwYnT9xpguaML6NKYG3u1eQUZmb8NQjlzZjS7z9cTqo8uFFIwLk+/MS
vwX+T0enzOHshWGafDzPo1rr9aL+8FIlU7ptATyXnwFqcC2UcHvczb+pMsg+0HIX
j34klyWmhIlTY6CWvn6uN3bRslm67WQugCHHrlyxGHXWI81032nOnWQL1UO7Sn1B
q6YgDHHPtuGIPjxK4hSw1+Dso8p92sJ3HKG5onLqlG1g0Ce4i+/YZbDlYGOg6Fy3
KjHWK+80pRFQMi0Y6tRj4AzS/0KQ0V0b5aTPmOe0hJWDXqwAJxo5X5Su4fFqUtfy
SSe4RGI9ixlRTlDGY+PqakNS3krjBoFwNken1RIMm32SNYo4IXJau9GelM1/TXx6
gYmPhzUMofIl833WFQ+gZddM7et5phfWe7Q/pkwtXWQCGZAa6AdGkI8w/ZXN7sGA
DDMETTTDW7c1la2hErySZUCM320Aev8V2OpX3H39LzzN5C1DbibuFYTkChyAhDtH
4aWU1YgII0Yqkx1ARdPVAG4H+385qZLzUlTnJ5bZF3DJ6UrHE3AeY9e9/JnUF1XV
lniM5ssgkbhhQAzdfOpXFR7blBJVUHbZLxP4mGpStA7ykrTe9XwnaLbOP0snlue/
4wZFgJhRku+G28ZrkSd+IIzi7YMuLqmYGBDkq4Ynwe2E80GmPKoJ6NUTRPEVMHAp
uo5AizeAdEELFikKH+PCifGZUpLs35gjBKe5fCXQKCFp4/yPewSVC0VreTxkAerh
nohfBDMkCUgJsnFPD/9iIkA4+sYG2sRHGX16mrCFgtDSU9xo+c59OM39VF/5INXX
qKE5KwMG8o4ODoS9SRTVZ+0gKpLAzzI4um2XBXSYa5OU8LHSPFR5jUogu8WGlKeg
FttX0mLfVfvb6/O+gsF4E5VNOMR72joU5AZoZTjDd6sTJYy+ZXiXsD6Jsn2Mk57S
UcWuNNZPWnnXtpDh401ny92NI2PxxwtPHifLMRdfBtxkm/tiAsFS9kOwn2chwioX
YN4LOXwjZQdOSYq+Y3fBm5oxPCMjxBxoauwumZJ+VY+VBc4CeX2Em6WB9KG7h9OZ
gjwioXkU/cYuaQCx93R9Id2BttcqAvbQHhr9WqSpUf/5abuJ7ELZFVUzAfBkOX3g
NatZO8zKxqK3H2uJUi8+TvjdMf0v+o/IvXvBUhuR7qOxykrhWZNbYgSKKkV7+ewa
cVqz6Fh/2BRzivZxhOOvQg981DuyEt6Wm56JAT3n4B/rmTA5WtMERRszpUQ1jsSx
qXGMk5dK7XSAsJFtDgPYZUNMnTng1IydhlNXsQCh9N0INLy3N3s/NcIgjIEqnQP2
oMEM1YwioRkO0zDpLWbAmmt/Ki/voaidyxqQkf0GlAhgFwONnzXtCes2AcmY8YsC
twe81+KkiIip+0z7yRv7nYp5jhfwxXuuJObBBJzI55Hq9bahRovvNfdRvOwDMIX4
OQ1i2+Qf1aiNSXkK7mD7G89Im3ivLbLy3dyxZfKNyixwNsSufac7+UmHMvdUy/lh
x+Yc4wmS+oPJ9FClhnkHzs7Guw3E6rVZ40qssAS0qQPPpbCu00oC5perkDk3iVBE
Bp+vLFKcyW/8qNasx+0JtBx7qOFqZngHqnMJ50OV08GXsrLeTbmmYLnULMg7UBQt
cc/oE2OWMV1hkGPL3B1Dl7vuW4XvXe9MIKptFnrxZWS8WZsRwvmKCZEqYp6czH/0
3FuiEY8vBuQ/6uc339Tajp01urgMFBVRyMdSz/W2cY/6Yw/PB3IT2CxhxmcJPQQH
SQs1/kwZu4jY7f+69NJQCBa8xigSInyru0380Rseb43LNzW1A/Y//KDNCzoNDd1g
djXYGTPQcyIeZqPuOcJpCZkhaB9Qcd+i1gDJiY9sAt3PI9IvMMwXtGRqpM0O7iE0
5nBQ5dpSkAd/Wu05q5abq4n6RKy4i5ujEYXtxx6+M9tMb19V/TE2NJ+5vU3XGUc5
BOWYr6WYNDxZK76zoEPfWf6pn2iLZUGzQ0wHQKY2SC4218rTF3CxXQgYZZB2LCZ6
Mua4zAjYNxIM5SH6kl4owXX5GwKKSDOaqz5vNmgsY77JvUG/FLu/0/R2m6y34oFp
/30EgMaZQuefEejUM0bVLAxDnqRh+yTGTPwUz2Lw1Qr3I53+2gMSVE6Ec/yxOxHA
VtWB/OJPP/LnFRkr6l0/mTKApTNqN29NryFQM5LdQJ42g/DdcZFMzSjXLzqhR8hI
yGek2+ilKueTpNPcq0inKXOAhq/xBuc79pxBa9tx4zs6TnbGXSwif6+8OzVJ5L6v
TtmhRfAJVetWW0xKiQItGAqFEA7I+QTG+HBjwCmgnu3l60bL0hqpsHnxsdBqyqHT
thOYj2f3Y9g98EI7OyrUXFA2nMDIRTBD6//PQE/YjdBcMBG7ZiMowPUS64Vilvbu
oodvnbFnbpds6zHtzy2YHjImQs7tWdf4VHv3H9aAXcDry1EVm85jTy1/PRnNz84W
FCGLeGLuv8HdSlQaWx7FwM06GX/f6qIqRFyULikXJYKB+2AOGPlXyGFgKauhtuur
CjgaBEYhUCyT8JBjQcBQoeop66BNBktOb2GiwtqsH18zV1WnEBNb4BwS5iYpYJcR
0mdqgTWado0YnbftlOIrRm2hsrZVg60xcuUungX4ki5csO8nIDnitItEX/9V1Hi6
YONpYZADwoxCEY94YqSUQTA6iMq1mlO+zJVrc1wq+Lku+i5PlDRL+i1wdvFqi61Q
PljGzzBZskMB7Vy8pyfHE8b+Kfo/DD6mxmhPJrD6NVZI0ZmOl4IY1RbDRaCMDOBA
uhZkPKKMmEKNrhIyNG//EJSUuwM8B5kxeiwZYUYNsxQyUeYRWTq9xRxLUhiK4UOJ
Dmchehypi8h1uqxify+s9TKa1WKbCLMBtf0rN2s/eso4MwuHXbWBX2VRlESv10SH
wWjU/+dU0cA/7/ZoU925wEIpX16x3xUEUAeTdabra5O4Z7swkZ7pbSfFQdq4vIW/
KOV6wqCePv7dYX2uHYjWtBpAhPzAHJKq+si7vU8FlD4gpDLHnsV2hbwMIHOSutOW
ReRhO3YUg7vlBe9C8eVapnUHCqmv3gNqTPkRP8/faXqFrJ6tMcDPWNx09S0w8mih
6hUMgqCMtFIfRFIi82CpidIVwXrsnyIsb2HfEYy13FAE4Ou44/lvK1tcsag+cc0d
+z3iA6WtFkL1yqWck39xL8tPmkNHmnMcaEghWfAjMp2XEZnFafosa4Ll6xqSkAzj
ZHFDiTMIlnG5Gzx1YdYulaMKWgHhBymBumUVzUvoRIp5ZCeAKMntUi3S+VqGlM/s
mhfTOrJdaPGHo4DQZssdaSZaMVvsBl07O/I4JaTHeTtH3IcM1m8J9XaPqWB44igj
sc9NXOurDbq45NAnNevG1tYNI1486rKHS+CS7RCIH6fbotP1yh06Qq7IgE9BNIQ2
FV/sB/wXdPyuj8aojpEr/b8AJZr03qpqZntLwgIoeSdMhpjIrT2Vyly7iWL4765C
UfsyYmrwC5/a+dLD7EXYlJTM36nAKMpXCOxHWT/rnb1wfs9RKpDdiYfjMZ/QaJTB
EUUgZdX7VYiTxXdAPRAVv0Q+0bpstJsN4LiltqTkxdR3T7GjB4+qLz/c8KJUz3pR
nC/V4tqGm3Xxutzv+pvTF/FLFDrbYJIXUkU0UJ699STcYlKYnjHibrNGFpB4uS7H
DXT6yiUwFcctN+9s8al7PheS7zdUUhGO8JtLZiqpcY2eLR9ACgFsZKnXIKTClEfQ
y14S8Xp0MKSPLC+ydmlR3xhdRm70shDnDHFz7A5CxqzZ8ogbCW2kCd5/bHSaXfI3
19c3EwhcXb1fn8h4wXypxh0p1QfimSADe7TVxhO5Kv2SHR99LXHBIKM8GiPqH/EL
UuH4sZHUyJDnSEA0EY4LIK9JI52exdkl5gmM1CJzloo2YJhwvIaF+cXVSFaLHSse
G79Gyv2ZgEInTx3Jt6mPlhrzGVyT1oqtleiBCgxkclu3/PqiYycLt/fzQX/mYg96
JJYnst7aiKjEsgpd639xEQDC+xUhlRaNonkx0ANcX/c2f3S8oipmD7w8pTatL99X
FpEGAgGXE+6WU8fr7cY+4cdIZPKeYoNEDcPg6hWD9sP33nFKzT4PaYkgHav0SB3G
25NIsUznjgyiJzjvBOVRR59tR88VkNHqOa2P9xrS+XPNW19ahG23lsqL4KIef20x
ghCpqIpRrshaNe2Gb+5rWHBGU9JMzyfijDLrjWgOPIwsYaDkt1uifB5Lt7ad7ff5
KSso7HWsdxXkyCfuVekqctSds9yzzg2knMsGMFSN0B0HG1OTLMxTPCOKMXfAYduB
xNOVhCltVA6H+uy3vVEzuWhJUv4Qn2Ng21qYgoA44J8VTRohnsn8Il5s/VRZpoZe
ZvZ+QG/KFLDSVFg16QsWOsjFs+Dh9dhp6OZnkFmMlow3XBXkb7/mSfTXZ904g7UX
eK+4zWpzPH1R3QwyLIUma6atUXfYycQrc28ISnrQpoJxcWCbkUon7EyK33MjtKkU
xvWjGDTTBjfiPyK4u79gzRvKvrzRLyHsGeyN+Yk6LqQvIYYDtajRNkdiEjAgD/u6
Xn3UJKqH1NK+GVa2gTa2ewbbPLDTGfvopFLi2L+C5SF+LszhlfP0LBdmagQok/iR
M18p0Vhw0yRkYB+nefmBDqlePs4VbBTRdAi9rYmCtTOhCxUhDlBVHETcM7GLWG9n
cSUjnfFGcjJDx/IjLTLP0oDuWYbPf7Qi28JlSpZzkxjR0F1xggi8O9dHMwhAQjyl
uRgmZWPO74zuuidJSd9vRVH28MxEi+L08/RrCeQ+7jLcCQ4oMcReI1/oe1H6/XPc
CZfX50VqOtIl09SKz+D6qDxCZw+bYxYZEgyqLDc5XuIOy86tFOkc8WRPMd5pbTul
o5M8aQCnAyrOpNMStvVM+jbH84jTvsSdAAfVqs1Fcp0YrhckK+nDTuzlFsw2kV64
zQU0QRqMKZA5nHFT46IO3+So4dsU+hU6CmLpWVf6g2zyPAKqJU+hCi7pZvHpQSsg
lRpvRyxcuHxWXLwp4b6wogCLoxcdAwzd5EGGXi9Sx3iqnday7hvRcqPz+5ZcyfiK
AtDU9xGIIC64jVTLSYMa3eYo7w5IzKOLXjdsngLDo9gRs7wFYcK2kOho+VR9vaOb
bs0w2VTSiIEqQulOMD6d7hZGeXAOBWri7N2nJNfpHKxX3bGXXc78QYX3INaZBAiK
X8agmZMGHBlp//XJNLz331QREL9zfz1y3AsLZ2A636nJ48AwJhRSe/54jjw9h6p1
Ir+WAezFMMFR2gakv8Pwt5HSewF0WVdEaOFzT5Ud+5EiC5kFEDjFJT2KmiA80lwO
tkk3p/Jdbcl9MhHEgLLl4SSZbHPsctd/sg3yw2zsg6SRKxiXrhVJGX0n0QMIzb4N
rfCVsxywnDKy1h1uK2Zs8Pw5VfXbK3+nsVKZJeW3t0VznXo3pwXwu6WaxA3tlxw/
4SBUyK8KBmP8ydhEHk5xhXfgGtrpJ7JN0XXCbgISpsp5ETD3ET2ZM9/lKk7f32CX
EMH4eNqONRFHJZY8ii7+7rngjmkk2EUt4zWENobqoxhTH/3yiRvIWQVwSaab2huW
LjtIpm2mVAv6AHt9K01SSH/yga3pZPm0b07Ojmoj58n0TlEsSRjapB56xZFS6zA9
WmPttntLh2fHzZ8+LP80I7/T7y6q4QY676qQhJDHreb1+SSW1oNlCN3Cb5PT3DF7
S4g13fgyim2tWxj85pJlX7sMxD/DqL76NLkxkeQU+MLwu9+dCd6cvFsB9C2osYLB
MvjL1LKNl3XDD1sAIVjvS4kUTeS8+kO9dwABc/5hA+9/K3oWztV5zpoRDGUoLzmq
8bpe1X/0QdIIjbUUmCpKWo4WLD5d/rdgZbOAZpPvNTeC7/uefoPRnwdzwEst3baS
GyJa0VimqkgPgxxms/EcWUzOE1h4He/bUof5gwfYm5HIdWi5Jh5Ecu5dM6bJTcQA
g5H422DnicW4VOHxJJsPzSoUmdIPr0klwVi3QA6hrdGK5o0BvRWoWObM5e6c+MdL
sjqe/26do+U7BfDtQnTpdOUpaFgOBd+Zr2ZGYykzveVrDMc4YxG9X95Tpulw7VoP
ZYSg/nDjKstK8o86YqY3kZgUA6yWzuua/Jwi2WsZHrx0Y++5bEOKDCwnWBaOhQWm
6B9Y/oVs5yvp1NlgQD+0xUuoRhWmlla+4gy2ZbQo28SmOtX2odr2CnySV1mX0xsa
bStirMVh+2ZLAV9/+RRGcVIHRDebInIOPxKGvYKlw+eHH9pMpXDqqJu7rrqmjKC1
rTWeOkVb2+WuAxFwyLSGyEN5V6G2t8AwW3mcmug8Km0GFVrSaN26v4Uhg/FcEKKd
KFvp8XE7wUVBvew+6HCBjPc7M/mnxJJneUSoRUg8s2K4TQXn1OYlynOP+gYKKcC/
WocrAsKwJy8aCwjwFji/bTSqd2QwwRZ0JEYhmLk3uFthjF8vuc34glpd487aXv6B
xEZOY6WlSWOKfwpkngpU8oXRvyeoMYivWkuhIYsmyw8k35DnXmAev2xbXIqeiW87
FvRG4yWnYSyV/TWVwWEm0Cs1HZitKwDNpW01wkjlM8o19CGsjWIGOaeRBsm2oH3N
TlOwqEDNeIge1ZFmXDEHhJXv9S6Tx7gqFls6hFatS6+cgJqeZKvKacCVPGQk44wM
jHTGgr3pCIOC82TzVBnxoTemOHfATourSxs1dFEE3JDe3FFDlm4M4fhStyDCiDCx
APzpgQil2iWfIeZsOuuL3AIo4/+FL5xpN4s0RunQDyXUwBngyin1+8+tkYOJuY4C
TmCS4jI7656uv2A/+yA7Spd0OYe+nFqjNYgIROmyIrVo4Qwcvcm5D0IfyN36WRZy
aYMN0WBd2xwUnleAUIrmxqw/YwumjvPBhpJLXdpkQSb0bxu/tzADkp52VEMjYghL
JqhJ2H29aqcKCAxfpC+6zseXQqtoXHuOtfGU31Px89Wq5NJ+CbGU+J3DCDTIPRoH
EiIMlD1+vRLhbEHgzFJxzOUy1BNp4V73klcfsVpU8fvctAPw5fV6uDsb3hrsK1Ue
TXzobJ+D7B78U4KcjQVZmTixvRNyFYRF2wxPFYKo4ue/AZenPI+uFHINx3F+S8qA
fLC6k+qHOE6fYLFnYudw5LrEzj+wh35VSNPTT7rYOq81q9dftk3JDMXyBoUJNbG7
3W9HJwe1Naxec3oGSgAmbzyPCa+KzI3AyA0TjJUZe7kyjLwZEq/jogMgl7y3LABA
yX228tvofLK7V1OxyTDadA/4l/hAPPmITrKkORaXJMTiXLoDs3uzdmEFZiyj7gfp
WWtqEqsxXywlZ78X2HjkwPbYybAtrvZLoQT8g7NRaV7wIPb3zKaMVmxdZyozgHvr
vEpS3qJ9yjq7h/P4/ornmgMM9joI3LeQUQAiOPgF71In1Jsf+FAtDT+3QgYppYnl
QvDmc4ZitZhA8yiGV3Fup0xJjUC8GRIfHo04HzqImX5vFYQ26S1RKkLqIV8jLwFl
uQJvdVHd68dZbf6hBzQlHERbW8us46MhQH0bJAsj1XwsQleZfLbw0bsASGgCwl+Q
YRoRPW8MG4eB9FrSPoyeeURhNLKQaDTDTcIbe4ghICbA/S/Wbb7Niu0EyotuVEOJ
jtnXTkHtTlrWO7RGqQ0P7/E1hcFg62cWmt5uzXMoVjfTG6r2QdPXH6ntZbJlQlDY
/08gCnvz394OrWlsevRm3877/p6nRNouBf9X93Hz0i4WWqCDToqtRzK+JXQGIhzw
XqYKA64Cb4kTchDqQRBW+1Qb38VCqzjxCoCQ9OPVDj/xytRaaZNWhwN48lzJSPbw
dJkdVYiPc4qqIqd3D3ClkkSqhOHtlOvefs0ZZKLt9QBGA9aIXzOLMgbROnGU2dr9
hxrKZebC/cBkwi672zp4e4gkTahjCfsVazz81WkTR9uQFn0fAGLnFkmxQZwaP54c
KzSNnYxIfCfyE3nVVL7hwcziVT6YFG8/Eo+HHcGc13etiatX6hLzL6phZ09k/5EG
u//pCPD0MklckUyxs5DNtc0V7/ODWpUV8GvPz541CeWFvREKt4QsHrKcWkSzUyfd
GmIPQj0SFBm2+4U1okEIFw9gx/9KPHfoXeTQHk1eIShsqVZPU7oQTiSOj7V/xvFm
1nrBKFaVBIgxQoE0j1s1IPf3prPsxKxC17jJoAWvfNohl2gy97ZeDHikF58O2Ia/
BUEBLhmarVp46dYBEnbcty7eUwN5vWLHMTktkIUBCwKEcD6c11EUzDLeG/RY2x0B
c42NQYe3KVJDS4976teq5JX1XIajakiOZJ3BKKkZZjev1z1nSLzfv3RzXYN7xtcZ
F8oSsBMBQ3kZNCxEQTORF6zCYV2dEyByMgkzQDcQs1mIHoevwCDc45BIoHhddX+S
C19N2srrRjfpNL5udE+VOSzEKjQdjmcf+2CR1lIrRFGVRj7vNpGHzYyIgjoJyFjh
QBDmwLgB6oA/z5GYOQgC2o6SD9P/HB2QBhtgQXuXuseB5Up0THASGyh3B+QT4vt8
dakzC51kkhXVCP/XIC0Lm67yd8mmEZRIABSZgiWQq90RP283JSC7Yd0soZefTx+u
gaYygPVHwD1MUtsRdSOyBbWClEG7hNr7Q1zNINGQOXX663EFRPbYiMynoyJJg/z/
Gd6cK19rtPvwE/Ee/eVii06MiESv4Op69y4UoCrYnbp7Fs+dufF5n/ls1m5sbHIe
76vJdbM6H/x62bTC8+qn7drvCtxZ6vWzHtREyitvf0Wo1fQUfO0MrvoANKv+g9wK
aqoMV/dunUK3vSeVnPu9/8k/klVBZnC3AZGR1FurcG60y2Q2xRqiQEKgyrxXZcXC
E0JpvSGcOt8hN24Cja3Jh5iqmbsnWNX4c4HEGzqtHLE9EQlqX7iBdWSJIz8DN21X
bK+hg0Ypj0o1wJ3rNv2cbecgdNcsJl0H4RN1TBg5AdNorP9atYqDcYqS++ERgPcj
aRgKQwixcEeuJS9+fJmYPfSC7M1/LCv/AuBsgtyPyt9HjJvoTyXrjlcEoLrPA4hq
OkW5NBsoigPuuz4Im7kpsJ0QxtkHybCN32vWOwen/ujy0yP05OibEMU50f9HN1Io
8A9gE9zN4OmVJDWhiB2xoO7mHNF7Nvqe5AXGHzCAF7w0IUzPJ5VUHePfEzSsteBV
OMmIFIm/CTUmldpTs6s9rTxz4cGgHaXRALssCHACn+JMVP63IiApSCTsfTKipbe7
qENIT2Erkxf8B5RIdlD/plFiXXHNbsWmEVgF4LlQMUwpN9L4hd0AdgDqgaAd3jdF
wtY7Ct+ssQqZRYdWRL54hgVqjoHA9jPLJv4/T8SPqtYYYBTLx7Y5NurOhJYJIY0z
fK0KLbMZH6KAj125XtCbrlKiBQuPmZrRjv0MLSKebQiGdWcpKICUxzLpbCvMTMYM
2afiFgS1+Mgqr6B5zncej94bhV7ego/ie+gCfziuc7OIX7uTckrpuk0AyPTgM8bi
pb+Pp3gBIxhzDev9f9W2SYoa4UuI0iSL5ZHwoFW8g+1sowK+CAXyOtrlLPK2BDVR
JPJp+vkr6kOGA3/bFkxJaUxjVXqeCdR57SP4P5N2oyyknGVkbj6Mqc63kN4beej/
x2R50noL7I6SJf5GHTJBTzdbG0r8JbpQUwxI6JH+kA1wLPu/ULfMyIMemgBKozHF
I7umBYEM/ZL/Fe+VskWCTwXGdVq7Xe9Wd2aCMclNebkoiPeAVtyrjOl2sJsH2MtJ
Tvfkova1B01oT+HRBxN3wmzY8n1JYCDNirk9kfoQKOG/pcKYTaOJtE4Q4ldnpXtS
NSLoToH4gAI5cKaBkSEljzdrmIBaEhzkvCVXNEUzJlSDTOKIhJPTRj3rnING/E8q
mFGG4p3RVCVtTcAHOEISLwZTycN/WFI+ic4sflrCiIEDCk0fAiNPlli5B0AYRdlO
Yq8J09bTLpg6sCe1vuzBXzz0nwJ+Y3+Ml5RYU/9U/+6iY2JO89t0mMHPd99Gy8lu
eePoYp1M7Ll2ayDZqSJi3ootru9InRPTacUa0AN4aafy4zjJDjxM+vKf9ZmqZCl9
hsrn7IbAlZBqA7ZBwuroPhzjEgwHw5NRBjfhh8hyfrV9CbkKXW0gkrAgdLx6rJCV
ZlIi8fxoY8npDqXr5YjnDEVl2T3KbFsiNEGGqnI7DHd9s3wilmOrITXQlRC3uMyL
peJSN24tR+eFjDQyXYavdkaQVmpOzyYEZkai9D1w1q51QDVHz608hukXecw9nUAs
4/7wqwN6Mcm1QriSAzERdimYnrunVEcFzTzVqqCvWiMlksOj1XFSjwtY8OG2WoiR
VgxPJLhTes7qmVmVtCJzv5PxyvtGpCM0KfuJZHEviGs7E3YD7Ox1HJETdoMyrTau
vkSqj/S39Ok4sEjgLt7aPMZ10kZWebpkstH6D+TnBLSoK5LZQl3JG15dOyQhjMzN
4M6Xd+wKGZFZkt0lOjCeYJrtNkzinrwloKL8XAuqCc4DC42ZfFh0AKt9ubLKr1h5
dfKFXcQ0Ai/jqTC/PFTWXjK1qB+4YwCf7PunO5amtUL8CZuvZU+KegU7ah5Y1JNp
g4ZpQS01OF9qqEDg+j2G2o0Rjv9XkCdnukjp4BQROqXRW8olVTpax7qLQQtk2JPd
B8aZcFE6qviaxb5Y1vEWQBS7Flr3t4+/Ai+yEKd+BoRkSrVMEr+OU94aSfrKooco
79bUXoIEmwNgaf2GY9yinLOWXg7NYqA+r1SoQj/+z38lKXWniz7FFF+G4uNTtYd/
KNStMEKmNxaayOlQ2xb3UpCde2HKo/ZN7BtlkBHmhtxygt+xD1EUFXUxNfO1lVbF
giSUg55JeAxcVIptx6551Xs2jFBOOJ40QrYh/BC3RKfC3EGi8i6+Sv34y/HHTlld
cxa+5ikafUojad2Rc7DewzLRQwqVyr1v5Qqwvj0gal7VuB+TUNXmruFyJpZBDQgq
ccjVhfhzy4u8Bnw0q2s/Q3Y9ztnehXTDb5LJg4brzErntmEf3FPSgncMr3rPnUYX
h2o0jmD5Zsz25WK4zzkecG6WUbPgUU3JnhsHjD1WT40Y1cgdkpl168F06BtwoPMc
5zn2Swyvjf6Qk6aaZCGrk2MkPw8z2Q07lYLBOJ25jrIHeHvvJv35I+hYw4UaGXuV
1s+ONdp2P7CRc37mnIQU71zEds/od/xfp7ck84MtC+46MO/RbNuDfIYQgbqLf6b1
y5txy80F8agpXdzNEWplAMHx5ipwg5LwAy/bM0GWBNvH1YqhRKOOyUORNWAFOkE0
EmjkXpDhmqmQ3vQb7n/JcRn/pI/Hqfi2t/1C0E2CuXp19wgvtryYdC71Kj4zuo73
4URsWKzVfiYvcBIOdWMRSjBgesQPNF5w4aivGo6SDgLWqV73N1WpnO9fv5QSEa4e
NXONZO5k2LAMcPfij/HsxEWoDGDKWzuAi/gvzIwA4XTnOLD0PjARbfZBZwLP+F/+
Jn6PY6uxa7G+pRsZ1Br9OGttl6Gq5VdA6Ker5rK4i1T7QNFky1A3RYXgxkT3NbV2
YAoQq2yBggjUfJsC6CLF3fHJ0JsyOAkBSWXijDMCHLEDfXSY4HgtUgMMY6Iaxrwy
FLlvHtjTKh/z+l8GWjsrdSUauUMj1OrE6BJKdVfgCK0NhwzwLFgrhRi3cwcKUt8Q
MZRCJSy6lfMeTHejIhyM1d5KR9qonaTpAUOtkHPaSHOC7MDxJZ4ngX01lozltWM8
n04Zc5Bc3wnpiMdZ5nuaeEYlkpIOa40UWk+ZvGFvnAG+a6ZWzAYBe1uw4AhRDZ6+
bvaw/2hS2oD3PiQMCpQ5/wjNwm0Cfo09elLHqLRuVInV8s3DMF91kYDxlTjUVnMo
Q0AoGyWE5RDZd1my8XCu8twxHaBDIBbmTTJHmjOyLt15LTGyvtPCMu1sZWi/AwyP
KpnnogcvkXEFZv1SpmHrvrbPiwIojd91j5VTLHs+3LYy7KpB2To+J/ZwMuu98Y/t
41+w+lHhZhCim3wm4DSKxT/Z5oI45RjPCJzW924gcmIGDTKZ+0ekKUyjqIVlLrIG
yPHl8enwghXAXkVOd88R+/iXlnixkGT3+COgQ/x1QeluHOW238TvYR/N89Knew2i
WAyIanXR9oPb+mzyBaHoUt801PfjkBsfnaG92S3mqrIXwq87xx2NWvi0RDUHLzZX
pTe2iz3R1spLSQfawg442oUwbnMeEcsYQ9pD3vcyRZsiyNBr8CbUJUHcmc2IxZEq
T9P3tSwu2Ydbo/Hgggkw/4nNV5KnnV3gtv+9CSU+9BppKf3AV6I/YJ95XGyleswu
BBByhLk/oQjjePBaaqBo6Io54psglmDzXpAGydGFkEflEG5nsy4SEGljlMp29v0E
2HduXOaPCH5RdpC1Y9LllNUOlEVpjlHBRZZO6N5CuPb0xbXCTJnPrO30gMqRgQH3
embMLGQRgl7Lesgo2uKMRSL1UkeZAj5VZ05QwoN4W2TFWexC5AEEvUREOc4GRibv
vrV0OdIhtAMfGveSvSW4+Cgwh4YQcfY4HhCVD/TSNmQ51odj3WlzvYnSjGKSFVkF
DaRelSI34Uqopka38eseHaF1D71diPSirBXQK9VuGahWRtfRbq9L0PoLRnVizuaX
jVHBmroP/FLrMtVgWVLPTIgYs50IbYPrjIM3Iqhc7Y5M3NraRLI+ZS14VRbsYkoR
NkLc9tDGnlhtpvxtjtIw0TeSCoH94JttahgMkqMINV6TKQW3BP9vOJWNz0AqRGMB
w1T56Bc+cGxVjeEV9oigtlwupCUS8WU8uNSANF6Ntawe68otlI58JeSqbduo7Jcg
bleFr5nSOn6N7xw93NmPscMc979EpNaJ3MnOYwFGV+KmpmHv3+m9L/znMWcjokja
PdWBWsD95ab3BRpURpZx8f/5+RH4o/p2Y5ALNQy2IwTpV6PEWyFQk7j89mR5wvTK
TYhUhdi8KWU2R1f1yqQLGKnEeSRbcXuTHz+26hWfOwwuyfGeXINf8PM03qnQiUco
rcGrVh9uDDpGIPutd89kPzk66KGAyhJ9JnlowXcV/R845ar3YHApi9kU2EJVxTuQ
5dmW2SJie0D/ODmq2/pF0MBW3VxMT6uDi4xI12mQCey9lHamSGBrmMXW8TvbNK8c
nl6i9rDSK6RKtn9qNxqGplS56eZUPVNZFUncN60pnjqJMZWzwHxrx0SYRs0vEhp/
pjyoYt9MtEkh32hLLtAc1idhJCkFlM3ipFeA1PpDQzfcvBuJZCx1L+Z0wQFQeI6j
Z8sCYS+3gWF3yvpeDXLNZFA0yaBpVVyCLoGiUflMqQBXnYm76PUo1eFZqF6f6d3N
5rXhcT7hwRV9FIZ5JJLyF/0ydNxINg532qEC1GwM0Je1Ju53srisKDh6EcAOMSqs
yEU5PxK3EapcWUiCftjP79X62OqzRLuEdSVJOu+GIX504MZsMNq8j2sWwl7ALVyr
nmjrguTVZDELsf/nU5Hi2IxEDaR83+ci4xN4rFFc8R5TM1jqekxGM0BHKliGwyQE
XnFTd9vINqgB75+pJ+dKStRpGoMEWmcUML4A+wl9nKfvcxaUEieteXJE/yhX9eal
Y3wlfZUisi1BrPmTa0T26mvINJwtqvpF9mvPuGM3R6sMCLCjHQEF7U5aa08ATifv
H0eTLwG40rPbXKu2SaShx1/7Z/2l4OUJXoDu4PGGxH7q5l3vutnyjoSGzyPKy7VO
XsjfYG1EvurVz/ec2qGm08N1m9ekMIVb2Fk693DmDFO2EGitf4dICilnJoHPkaXY
jPkV613fAAQWEJ+efbuDa+eLy8T9wFKI5cYBCrSqq48dVRu3Lz1f5wfszSlrG+sm
vzdfUkR2gNRX+IuvjBS0hZk58kkX087r5gCcgZfWPFipDTwPnKJwptuqLlCfAonZ
lYr2Abb7k3NGh/1m4dFAiGAQqVN6hm4IIwH+tA+xjPDDycRnRek4C6zcYgS/GEnP
W7Z3LVInmuJWV7qoe4l3Jp1+urAqSBP5Tk3u4kPt03wt0ortVbK9xiegoMVmut8M
cJZ73US/P9+3kDWuFbi+CFx+EzMjQQoz9y9U8Ip/DKayhZlfNza8h9cqLKKvpOtk
RVh8YZ63o6Qx5BjAexgA0ZFYlIgTL4ro1XTd6FQib7kgmU7ttDOhM92Q69+SDc53
M56ExGuaZn2qY/f6aLBRYXHU80HdmeWWrki4TqDju28SqImJBJo9jFSsveWXsFbD
bjS+57aXg6LT68Ey+OD4+iswJ5fOMoBFwDQvh323NViDaV1bQnbAr6MHCqrHv3CG
m64j2Rz/Stq8Eyin2o7+nesBKT9C4NGimvS+zeQvYai3CjQl0G1mgK8XsmHkTJM9
0ITZ1ReXt1mJ72oX/kVix4mzh6iDI2wWmFQPCH6CCXsDR0FMP6wp1hUoAdl5MOoE
BhBeksrwLxc4ssoUe8Oc6DapT7pZkLjGVjdDurCcmdgIZXNPy+s/6S0uZ9YUuUh/
qtXIrVSWmvqX3cs6oVQDMd0e0Q+FldyahPqE8hO58F9Ogl+t3UN58D3wILaRJHve
E7YMPnFdOdHHePGwtZ0d5lRQRgdrWjMAVF6MviysnjWuPr9fM03TanDnsLFOgpka
+CM+LLpOWEOkNAhF1gZ82CjJ2RBRRZG8xAptnxZY1l8/haVshgcjyDy6i24SSUXQ
U/KlHqa1Pba0GlKlv/nM7RmaF+9OUoCD8fQQdFKq9gKppZl3Lx0YeTor70Pd/qHF
NtXESOQADbxSWTvZxTJY+xY/EPdsLNCr9GY5xdTIptokjH/auy2Pa7C3iM3L8jJL
9lWIw4gYcxKYJIqZS/nPifOKAiao1gNgxvU1tv4s9CdD1VCOgeMV8TbBGi0XjbbX
6M25EMP4V6A2OGGT8P1sDv1osp0Vi68QQtBtco2UeXxQn99t0l0Gc7tBCgaKYa1F
TDZsBQgABR/Ogn6U57ydalKNqDlyUwpcDtw78JLLnmdheJfyrU3nDFXCY9+fU/mS
+hSREyrlzmjGA9o3UrClpOoz4mFJ9EhgDbMw8pDZPH3nowfWzTSVt1Y9wNwsLe54
6ZDX1ZhNxm6aG+/L8jr1bE88UP9DcwauyGhivOhGOsBae/FpEM5yUVdRdjinpKoJ
sE5BDUlq05E/azCvEJrD7R2/WiVknDc2+z2xJTNBeQTIZBUNXLI/qw0h4O+d4613
xpFjJqM8FnuqN70ov3BKymkEVpKOfgbyeXopcdpqolDjS6cC+Vz0bvII304WlSY7
8rPWE7i7/pvYwCyD7CZwvKNOI8pt8urTUm2lbub00VnNG8bv0cQ/Obn308VNIn4B
mio/rGlq0rXo7l4jajaagPP/QC+Yn6fP6r3JTAjdlH2DBVBoPjSMyMvlrI+zwrAq
lCx/x4vxXdTYP8POHdTjb3ksKLl5njnYF3QeeVTyxmkNFNtqClSz8l6cDHrJGAUT
6MDkQynihQLdBCS3fxEu0MGzaAeKpcRtWsIQYh4ruCvJeHRQJDLG82Dj0VEzEhQk
U7wjDjMKoX/8cHyXbZnzGiiiVXrBdKlHNc1XImcSujkqn9nwTc2iJlLLZ4vzrdaw
OSZbX164Dxaw233nBs5hDpaiKiJ2JTLcTjI3mW80QE7PSdLFEtRa8JO0shrI02oE
VghvpDK8Xnd8DoWJmQdmHQzZWQJEJt/qfU66MDjJS9daqbtv/dM4/bofqBI+qgtd
TdG80tvdHdMTdDI/00Gd9wxiOxd8mz98DK1ZuUXuOslyKuisVeKQj1QIBlxmUeQO
yZRod64CAkf28flzlEJJVGC31X4xf1+Jfr/+AIIul2pDYaIjZr2scTnjEdwvUOtX
WqM5VgcH/ssUoauuM5eP0Pu5NV0qXlAuesISox2ezOLtOdGKn2BVAgNBSsg4+Lbh
e5P2LD+J2whNEAzccjrzgZIH4kVRMM1it/HEnBxXwDrwNyZWT4UI205l9FhElfri
Bt7QRyqlR3DlDppcRXMC0vAgxXenQ/rFC0BYV6ziSSOlL5ZKDs8c2vTTdvIbkzLq
6PkYIp9o8GJ3OWaMjgNirxZCq3K5KLY0GBXFJG9g5iCweGrFbQrwa561LdoYvxhd
Jj12LaTjTmRAhZpjaAGj4EHhEqzf3IYWmXvFTrCqy11KF3OLWmVxYZBggm0Yozd1
o3Aka9B53nT+bQZVuK60cNXykkEF6mKR9zCzhoKTr8Pw0gtZzD6yauwyh/B98GFr
B0y1XUAVlwFZhxITqt28hjGKhN839Rcl49X42F6sYQnWVao0gfBDnUUeHlPZnDbe
e2zhMaRjZw6cgJAZnUK/Z67I89ahyQgLREic8eiVnw9rpmFdAeX9qywupCoaMlf1
ap2HT1h63e9b10t3CeRr1AoqCNLfqVc6HagX4hwWsl0uuYYZXVjy6ZqXG2XlLK6p
X/qw8ny5FYvBHsBRYRa1wFHCZH9V5SZPuCXRyEbN7mL/LKn3KXaBmj0/iCmg1RQP
ccK4XS0byX0jZfVTxpNqSMU/5ZETj8ONW88GZ1H7R0xc3Bo4JjKszB/IOSmR0BIT
JZZYK6Uz+2+vX3DgrJEVjKiAMCcR+D7cZpDIjR3Sw4Vnhs63HEJ+f/YT72T5tz5/
UMWASy9/+vd7IhBYT4re7D5loKkp1xkwPaHDikdD5sAJU1H2M8CFyGDluk/+RmGC
XJJOaeYIxPWAK6ZmX/0AZCnss55hRQGr9AfjGo+uNTEZaGTxauybfx2Dh7coM3Tg
AkAr32v9ukrm3tZhwOdpHa++8A/0nrDr15uto3SGHDKicUjmvHIcmieULCSmYxRw
LDsXouEfzMMq6Oy9hscMjSw4KDtC+QVVAL9PNI9btwQiXyn5jgnt4rO2FBe82Sor
561m6LfHGGjhoJOwtMtXceqotlcMy42uh5n03fS6GTJXCpYUxx8g4vA0wY5mdXWY
NMqhpz3ZDwvpkCPgG2LfebfOD1J5lb/iA8po5UTLrO+/JWtdvF1L3HV2FGMEIHDs
IjfRiaEggcNBeGUrIdSVwc0bfRKwL7yKVWTlo89w3gZZtVBJ3iR+aivFj35HU7aT
3DlRQm7ypfoDyaOaDt832c7uzCtHDEbWfP/GsOxgkXa2XOfBxMuxGCHCeh46K3KY
gb5qXrKkv3dT8RagQyVpM7GP0q2scfnSF9CYGCb5QOH+Z1NqbSy7BzplvN82Fzoi
UYDDwac6w33tGQbNCx1CSRmKKesdV17gsqjtJFGbRe6XjCSkhzKpWWU/x/RBApPc
Ltj4kAQp6yIXtCEjdPTVZs7oObYEx1uxbzXyTJXQPaejw2TMmxgO68Alk1Q+n56l
LcTyVt6Sw3AuX646fbA4lOs0+bu4zEcoEzdBeFsi9pyaAfkgRe3JjKJecp3orm0+
E5K3noSFGmDwYWVx/6bO9DKfDIj6k0wMl9D/nIELZWQ6cTWuZ8+a43XrcI/2n62O
KrfQdtLCEES6W9+gWvR1emxsvadMc4ugoApjS7WCCmw3z3mwq0FclzjCHNFSOnPo
GEU4BGbLImRh/affCX+V9VT+PDykbCWwHMozwT5DzrL/UduKGfVPMM1fMI/hSj2s
u8SVlyU7tvE/G5KuYidc2X0DzfMe+5Uh4pKWxs8SiQAdZqopHtBFO1DW/hglEQXN
Sb3Cha/Z5xhvdgXNWyIkJivZf1kVyr5z35gl6U9sosygqkZpY9BB91y47r2wv0Ls
PPsiuKkFXyIKY/xEG3o09VgmRkNq8cPg6qM8a39hhoXyndVapWAq+cjqoLcpWUYX
8GonQuNL5q34ryARDq9EGp4veP8koTiszgF/W/Pfsac7iVjaCMbix+ADM5PjbLVA
3M1F3jK6yhe8uAGiNUKgJ8Spn+a20K42le6vMf48magD+4S3zz5EEnpP11SihYqy
r8j5oLXON9+YlRJuOjpUO79VOznAGPZBXFD9ePll7ZwD46qV02Ul8q9ndXANfJs3
TL2uJ4jBfGQNoeYFqGo/L1yOymEjHjZG5Tudc6q369RLEwJMhDUvzEBaj/emfFdg
CRgbuC5XeSHzvjHo6wxF544MChf3r4STE//AuPdIQti11q5FupREPSyfPOTpDFKa
uViSVFgmIY5kdMZKJM9B8OQo1zEEfn08qfTXKNEfJ4P5I3J6ukPJ0fsxauHiz622
6Ia4pFgFA2G621WUWEua6aKwp6NrtNfKoshA1cUDSIeemZG2YCH9RxepP03XJZQw
kxx66fvzgzOWPeR/oaABW2D97niBItYpeWEPoXRVdPYNUUoYe+4XuCnKmxzsEroz
up/4ZTCiHaHgtyUKniovWwsK+MqfPJo77xp+1ciBG3SM4F2QyUc17fSfnBYjU/zZ
kLL5EEE7T+gNPUbyhooVVQIygZZJzUFkpvnrlkfxo0akg2DL7aImSK4+Y5E42aOB
xaeOwOXmSbjWwhmzL0tiv3Vcih9KLSk2+V8Jgz5bY1yTqLMxaupNFF6v8pKG9Cbs
Wv0xAoFx1cTF+GMY/0zJORsskYzzELKtasu0gdW7JufPmu+bsU6qyXu8rbq+RvRJ
DDldm2LMqkbk4xsHOXNjiYcQADL+lwWeO6zgeW2Qc0xtZmKQkz0ZkBp0fdxIUllA
Rsi4AUNk02gsQQgjfyD7twLb4ozFjHU2ruzcGHdzkv2D40Psnhe9klpNrXROvRTW
VuXcmHErYwSMR2Fmw3MK8i7begIRFGzi5w7F6gu+QPiFMN2wQU0FOX8dc8kGHRXO
IZNv4xHlk1+jy2kLa93esJopoV9rge8UCIygCcgsDDiKRlDIb826/pR8EKLEGSA5
D1eTRr+e0HUF3r4j1EbOB4RwTzaOJ8Aqh1TCiEr9TNqs0RD9ahBp3C4eKkfIkWFB
H+OLnFbg4j6mejYY6spW33CxRAp5D7G/q+6ix6+Z7a97AhetQcpkduCxJ06/Z6hZ
OpYbWgZk63FmOp1ahb8KbLW9mlipTq0w68vO6r2PzDB5EhwAPL7ALlKkBhgFTb1r
/qdhz2MPQiibWvpIeIQ9haxNYCbwDgtnpbC9pO3RMCulbfYPkihV6JYFDEuqkKoA
X/RQQFr2EvrPc1nAy4VjarrE6Ome9MdJDQad1YS+e5pMq1QFsD0XATa2bfPa9uGE
0QJQLQILeOkwJXbCpPuwNMR+Rj8zZI+577N63O9b/1TfkXTZPCikkBwmy2KVojir
5k6rPA86vIC3BKRkyTXJAyy9wjqQFofh2CX/V5wkrKRvM/WLnOJWxV5QcAEhjQBS
tUXuDvEWtrhs4sJoRrfuyV9OVQmp+UHpKAnhRnjs5zQR3FdE3kSrNaT/BW858k8f
zERGrQN+uqMYVJhFU+wfP0Ho3gvEZzfGvL+PC7GPo8As9O430BKyWB98b0/0juWX
QArfjN3GMMvFYM0YllIgtianIjV28YwzwukWFgG2iMtQteNE5YLuFxn4NZ1BZKMk
eQf5eFVd3UFx1Irn5GLNr9lVxMaY3c6rZgrTuxnpPeWjc/7CLUYouGpl93dmMBC+
nQyOHPbuOVMirsi9hCfSrcvmNPTgzNz4mrg2Lx3GxFpGfnu4EdjU+l7xIi9HSXoF
KtgPiFKU/SXj5Cj/QDyIbkjchu2WLtGBs34/2jjbvnLNXawzcbizZ1jKkCaCzQPf
Ma87ADmWdk8l5eERZ0IphYu78blOnxFRwUXJL9vuH2PGJm+IlE+4Yo+M9OXFRfvg
rePaJTFcwZJNilub7MQ4VNn4fX1imctHQ1PHnrBeEZjkZMh4XAmu4ge85mSRu3EE
jR1MISTwPK3IsGWkrWpWMTnAa72ngtYT9X0M69JLfYgbxb/IYdaHJfcqoOTsbcWZ
J4BLT9Xnp9HQZ4I/2VVV0okJqi2ITol0TbV6BQCPPrQkzagCDjuGbZ+pTvtppIDa
UehLZwEWRe4AVnzn6OXIxTV97Fx2jn1FZKJlWR6Y76Yy6WcHOXMMWTxD9bLhThbb
VRXtrGamlIUTWhTB/ozt0k6MZpzIKDZ02dT7RGCVGFL/b/bDDDqEAZ/B3rQoJyS6
UE8g8eb9onZ2xr2Rpxs46txXyij1ZSHvF/Nv9yFZ0OZdmMPiMdY/qPtSieQgdaRZ
Xrn9Et//24iA/jkKMWU9lveWopirC0YacNkezjg6m4JBc3zsf6B8FrVea2YhucHR
oA9CG0fDdY8It6rRvRH/ub35Vc/ZYT7FU2MPMgwM1nqW9HvSfLyJsU83dbTb6kw2
FaU9DrjgsI3mgzMIIMS1P+grGT4xIYRTfMqd9JO1J/O4NTBfbz6piL8e3h/Uac2X
Fm+adjWwqH39fQFpAEJEEj3yGmfvecieG3reQvFb9OUlHywV27YwV+DatAAwX82t
I2u9Rlhj7ag1T5KdnVBRE+4UHymYUA/5ZIS/q9mTd30EN3A6W5Xv1zgW/kVUn+98
Xe75t5OErbR0MTab9floeXiUo4eXO7ENd+cmDQF3NeaAlRQDlEWFApBz2QLOUjSF
+5wwMnRkZcSMa5BzvFhubyQFETTTyBGGosXeRv4xnvFY72l+Zxs0kFAXcWu2v6eg
EoZ3iJVEfVsD5Lt9ZJIRihUCvCVFyHPUfo+p96/TmKSvXO1IY4tIAKhUMROTzNE3
ab7KTtzS7i76juPI/ny+I4xu/cZ/aRJxMoOf6FMzdgXnDfdhtgab1m1xHJ07HVOp
U7FpZntkj/Vda8GF+eGivmxcEU9mPaBK1VJlsEztAS1dpu7W8LX1Iq/uYU8+NvO/
8D0g0IBZPg0PPLXE/UqlEZTjlCeOumzNj+Qiy+HqxhJe3kMu0K2n4mblmAYFrn/C
l5ZEq1uyRHmXhORczH9toQFtkfbG8i34YVK8LVofjMp233Cet4qyIpddQMzlJpel
pN9yZWQaU+ia7rBDkhKRIOyr3azbxMFFQ7zDUMYDI5rLdBNnHrdUYbDki+d0RbkF
7KQY2zHMlB9WN3CDMtKZmaJwWpxCdF1TLvrS9XXZkKQXy/sb59GRw07f3j1PKzAH
sKW19gKbAQmzdm67dklg8Hy/GWjqZyWisdlMT7efSI1l78ZlzPylOLCSq15dz5pm
9GpJ3MOgqKcACxSnYiYC80Amsz6VGPK23XeAe7mQD00hPmKfDobvWYm7M7mXl/gZ
RckcqklydB2QEaY1OWoTIaNqA+m9VS1dNp2mz90b1HmVer9t5DESpIg/cRftzXvK
ouriU48jSHvzpGiRv+JS9kPQvd413apapZoGrNVmtGUUbCr72JrbRykn2U3UV5jm
3J9PZhE96S9GRpAwyFNXydEd5hl5iDWhI1rZV683LjFqCLZctLs+SfCzshoR9sa7
OLiF6VxHwwHJkbR0dozbF3QGXXPlc/QopI28NvTpcQLfCrMpXVEp8SYhlxBA8UnJ
XqRupAOlDlt9L5qis7hEwI1sbD4JV8+oPhVzc1zjsdUXmHDwUBydiosVTxUTqVgH
IjPEUlR91W+LOICrIOjDh6NYWCEPM4d4DFjUVakvlL9UBz/umTfYWY/U85VEv9KT
sndYFD0AqdhZWRHWmu6xFhG+9bfs37Wzy/g4xV+EvqPBC6tO6GI4dK+PLud1Wv5T
IQfHKfPlGzpGwgSt3rQCjpAzf3vaNJ4EzoTUoVcfney7vSfANLCArP7YikB2exRU
JNWRFsju1eTBwzgFDHoXI/r2riTt+gxrdVAQX+HLOD0zIg0+zzM5o8D2Y+gTDNdv
XWpmZGF7dqWQHuLqv6NR2WreXgN52pRuhLvYglwDowR9S35yludjI8P3oRR6/8v5
rzH1bBFv5hLHmgXcLuEj0aVAz9aBdL1MrG3KTRZswiJH/OcLs49hEm5gSi0wqoog
BrReA8z1cl3qrfaifOs5iJcUscEgcWfatpecJZf5Yl3YcwDG9R0/mJNSMTaSTRBp
VFvit/nM2N2Z62cH6JeIHmFIlimjYGtEAgsMJnO3/FamjxwPT2mL8EXYrOsAXNmA
oD8umGEKTdBnmJIGk4rx1pJVwet9zT2+p0xZ0jdJ3G+0jWxv9UN88MAfbOBF+5NX
N6Vs5JbGIiOOpXZJf0RHnNnbtwjA7prsb9DXunOU7L8daHTnZtmxv1iw8irwhBLX
WzdyT1A6cBf2XdVFoaGuTU2/T3AHFymuAqQwmc0UGQ+dw5h0NKgvgrdRjZDF2E8/
ewCnC4LZ/mZ+xe4udZFrv+EFpV2K6sNzBTddWflUFiP8atOsgdxZNk6FKSIA8zg3
8lBgIuJPelzTXhYWxUB/QRSOBgAIun4kulw36W3mfmrLLQM3tJaL2RdHFg+WomEA
nbbDoP85sL5McdtxmyK+Oxambbs3ftiYAbLsw069oEtuoMSt1+2tmtHXdanfZJ2f
EUi8IT3tCd7PeDKBVKMt6/WWTdRGoe4Wrk3D7Fc61B2MayycrIumf1A0Rj1HMehl
/msi2VLFVUxEm2Xy/IFA4G5Z3a/dc4BM1qslmgM3M3NvTWBWe7RceBHGeWdan6Nz
3Y8cGQu408EaiTiP7L3mAEOxQmwmiJMhuSXU/zcumU7iYmU7HFIek8/0vKr7Qzt5
vDOuKZuqTxAjp/lTrnnLV0x/rT8MpzzrGFriTFaSl6uT0nwJIR1oCPlkG/5byX1y
0yeMyUwv5sSFbQOu9r+I9Ab0n7WnyE8JBvJE33RB+UO2lI9kuR4QdpmUDpCj73UT
bL7sCRmWh06MzfctEqEIYmL/W91l9LIHa7TCPt43FbNa+Rcl6kAC95fY9Lln2AIt
YpuuM04fepBk51ogDGx8Yf5KNT7CvVk2as7Y/xPIcYn4/oCw+VzuYJ1DxsZU9oa6
FKEz9RNYW23yljXDDmqCFSLlRGc45OlgoiUZrYW41+lLwJJBbjZQwuBJAK8TsZgI
wyMFXyJquvqf3PbT9IYLzdhOXpFRGz7IspIlWQxRSNTr1dmJ+wLhRb0OVQMsnGbH
xxSAvJusMjG9SKpgl0ewYOB/lh3/ycR3PCaSBOfNQWZkUlprMpASQDauPIN93/c7
PYU5pX98iw5bq1BBLi0bNA2Bi8OkcC3eZs3YSWaEm7vvcFEWRBZvWc5lD17sbIDd
7q1z8kQ26EIBQYDwGJI+LjzbWyDJiV00Lg00sBg/vS648sV401USGbzKsAXPnQU6
93B06Zot+RzrLtKYSifJJzgDi9K0gy/fY8eVzlpjjqaT8gxuV3X72l73YsVWwa6x
ZDhNLVRfN9sK19a/XIxG1bwWuUP8GcL5QIq6LTyR2bbvH+EGicvMLWAeAnBaqp2Y
RrDJ5/psAOsrqSuGUxsRtcqGHHUIDSXAucbbyE1N9ce2dGHQOW6pRhQ9tQYbUJ4D
l86jEUbx63VPW5yS7muPPghkLcAqSy2O4ObBTi2lUGrUG0rrUd3xwmsHsWsnBXr7
QyF+xyW13377cFUQwZU6KC6dLthzHhfljXiOkZuAgc4aAuPHBIs8t3OJslyDow7t
J4HaTPhOxIQUG37Q2UW1nYm2NodQAiBxT9eQ/NGtKpXtp0Wnwl1Rbaq6rpgk1Mk+
o3q/xg2PtxZLvtNCFwPXmdjo1wTaT2FT1FWmTpM2fMW/y6xyuBoECURYilJAAdOj
twAjUYdyEquS4LUFpxExRXqPTMAq5Cr88IQTt2Fn6oGzgnu0TJLqAXPJYwnWtSQ/
ExYofssCSA6x70IEJr65DWeWe3eoAlx992Rp74OJsZ1ufMddiJN99C8WUG/Mhx0s
yscDNwOxZKcKSpsPb8ulSD0nvccJ1QY7R/7GMM/QRu8hDqmXfZ2NusD8f2c5dLym
fnATDdqEMju0LJR4L8Gm60Vx7ypEUISpwahQXk95gJibY2hIf1RJHbEBwXUGGItt
BOUjRJkgXwLRJqcRtj+TnbQNUkb8K9sC44VDUiQVyGlZ23ZguJicJrhi+vKnKJvu
XP08WDPu0ngROlaIFjOrZKFPFzT85HRAfzyG+3sW04CGGG7b2PQ39EESHRqagFXb
dfEGbPGTKQUKnQ72bonV2e8Qltq2XHzDEPPcAWbbCpG3lyiZMk0UuV7Jd29Hv4TZ
lEZcKkP5Lu3kUJHJl/ffNbdnIuLT+Uscj0sN+Sra9Vq88gSydAH+qRFddDLyoCDk
fQV+7q+Z0W6Bl2AlPc3levIJng0NwCUH9Is4lqllwautfnm4pR4/YBqZBre6JBl3
e/RP3Uw6ZgAzEiZjDdR6x0nCuaKsgroqaBsKMTBYc+UTAcTH6QWj5z0vnqnXU2G3
HZri1d8LohKXOiCN/6PMIMVA/nXWXxlzpHH/12rJ24ybuwvAGBovM/6LvGlf2zQj
eSchZA3lwAh5IBFRdw4My6630Z6VfPCdn/pQRjbiIGxFgl1ePqscWHrfpFrVYztn
1mat8SVbbejLUko7mlcYC+kdSOusVqRcEz29soiFBv2wSiRDVPi2rrDSC6UrE+Lg
f/Aviqrxi04x82BqhIbDOka6vbD4Dt00f7u9uT5OaKnHzxkwxS9Yw9Fym3phLnO9
gfgEfbD0XZmbvIteecaFGzlep0lUQ5JcE9g7f0PXwXQtndAS88gnIG1/1YH4+RBE
ynVP4Hyn/ZrXgJ9qol1sT0+vGyTthQ7W/1rpbRKaC7VlPJ/uiqhKKLEPQ8/5+afB
HA9zb27dLuRbcpK/Uu2ADdI80zDA4XR935cRSsU15y0ENfDkywyuEdmK6XtQ15rm
5XnTWrklv9HPwPx9UJjvgeDZ1EOD+qEsEjUBewAJ7X2txtVmOYJf6dpmoR1EZJQg
1wuPNG4IetVRtAb19frIwkgHCoNpCKAE0WA0tfNvKBwSeTrsb10AdZJDQ/2LfL1q
rq3gW+2qZIn7jFI/+/UaQM/O8uHR3ccNkUMZGOFIm6BrUdxUT+hSOTlK7v9twLzP
vN/RFYJTm3KlBmcsmq1mslksItWSph95BZQMNcX2jJxBdvx/hRaWKkMv0Q2RJenf
KDxUD7lXz47eNWqoA26ufKHT4DsyU+hi0GUGeN031xmMAJFGBzpsJS4lIPiHZBbl
ubzYSDK5N9Bwbrk3Fi08IeJ1YDs4sQZmEUzQpdjpLyEuY5pymMT/DCCDSUIvpQ6b
SQybTR4KOK/0z7qKkqYtDdyS++kPvPtoXfklvOeY06umvgQI9407LFJ3VJ/q29/r
ksIvlE/5hwr8C0pmpNfECujWERxl9aPeawLkwiJa2F68zvr8TTwkUZrv+6rSoyz/
nzomEKuWCja+lygc6yrsQlTgTN9deH2dHAZOBZqb8Bku3QReutekby/kDdtGfQcf
QThv/Zqxy6XTlolkJvchYZVbd/CqcNMTqvmWOB5SBBgxmN8s5qr9zGcyEbU5JVQ8
FFz29aELuWJ8DxMRm9DYpmVqsazQkiZpQeb77SqigUKNt9LD09uUYHvDCHp0RTk2
Vbfjx8VY97ZqREGnjhmbiFVmH+AW+ho8XgMPpahMoJN6uQgQLtdbkWKgCbhiCj1t
7gMJnU8dEXx8uZJpfGNM/2dhieKK20BJK90aASWCaaOLlIQ2ds8JL96J4psumXPd
NpXCuQ3VVbEMfJhHrTFWdMKZb4SK2BIZIQdfCVaGj9d9AjGD268Apzt06cTGTdiP
E0fA0n6yJeCJSa8KaM5X/YF2brYRbdc6HMt8M9YDsTPbLyplFIaMKEKSRZ4fv+D2
TzpzXr1q8Z3wiGWfYot7Q6h1yTuobOxeUro6QSl8c7K2uAfLCHfPFQGss2TAGB/9
6zTGe4vaQRIzabr8Sy7X+LpyxP/vmmFnT3p7kf2hnuBj1LBm+GZmUgYrjUGEO6u7
OVNKg9Xc7LFz9DJEZ+WUFhUh9cILk1eYA48rKX9CAInv+O2qDqvBlsAculEJJc2g
Gl6GbrG5wSVAp95HoUqmvMOvDfvYn8HhKdOK4ukpTkUZuwW6hEKFKsZDi8nz2G+g
A+WtbvwXp5rmnMfp3KW4OUouGrIfVF3mxY4SkOC9Y3us14oic7fhJCMOZF6mNHt2
wyYU5912E17KtvMFWCpytGfVWsrM7l3zMZj7+0ZFCH2Krc/3+OhZGrm2D4taNt2L
9n5+OtRDaae2emQpHaaH56JjUMiro8YqAM4Fm1IUo4mwSAQMMDqSei8ibZ2YD7/v
vY8ocyHdEJvv+zB7R1hd2QRG/PByeVNE70qGVSzreDaAduRJ3xKGQAmdHWVUiy+E
Kk3cZuKapTSk0J6/9ve+muIh7h5udbjSUXrRGU6OqhcUszhkWT8RKcpfX0BJHFL8
Ot/mdSkNazzebmOzVRcKntaWSNuo4ngYwOA5kd7QM/5V5DBDXnQpFvyw7wOKOBES
fPR7+i67Y8yAWQKZcMwqF/fEu7oSgKDnlklpMZaBGdgIKIzuk/RXqt4Bl5KmRtuF
9wXmGna7MyRpG8G2r8BZBfnySS31Ff9UjqGaStZ0Yh2OfZ1lt3kQI0SPxqjDdtiR
YDp1MIgbyV2Eefse48cJvrMJ6tULNPsjboXuI9leM4M5hxWUc5jdEVBkuPYz+TkV
U8EnKtqXg7Q26Wq+63QG9bzNwhApYdNyrW3nItNq0iBl0Qwk8e1y/OpWG6JXqiMh
ktxYH/cqBimwcucVpdCXWEMEj4GVh+FVIHBtzhG24u+RlNGdJtljKyakfJRvJgf7
6oElFIb/OTarRbWUtGgd1LKlhf7RCQl6qO3Z39m9VVXGAem9AhR9Py+su0qHlkW5
IszrEp9Gme0o2WqxuIZXGPzSOrvipTyx4uo7wGUjUQ/yQsj2iB2+chPFUjtPf2uy
6xnIpZanW6kwKWenbIGlJddPqLSIThZBpzD+1MdE5VGUFaWMDwtVeUhOydyFBQj6
MQLH4oafmNRX3Yai8+/BvCRxK13/f8rUXxXNOtJczLZ/sanTLhZ5AqphB4vDjL15
iDgniuZkGUSzpaEHvGcKVQPmqktV6tPkNA8CZccjDcUzssG3cwsMCAfnWyveh5dO
NeMxqt0yP4mhdDko+RJ7TGgiuA79mRRICcJtuBpUIEPBHPHtsqU6CmHvo0ylnVBJ
oaS+1r8gfsODbghpS15457yk90r0tDkkD79h03hSDgY0YjraBxhiVqyEa7bU8lFR
qn+cMUHeuP8RHN78Q++LDqbHHIQvRl6HXtr0HwhrIMajN0dqcbfkqUtvWS+FT0E+
uhYqs2T1E2vH7oiXyxgwMwRC8VzoGrP/YIfJqOgkbxTOT1obUtIBZV5vpoe1f/JV
//1EMDckKKQjp3KbzSqlL2PmCUJRCntqlvWL3GXAdii6qBXBb/CcgU4Jos+v5zwZ
e/7wXjAOPEn5wJGF2ZU12OErjRnK8vW1NBiATvvw9H3cv34l5k1+Ix4ntPQyjzxa
L4UUj5OyN1uIwGgWe5wZWRLkV5KOKQuNelxJTZUlvr05g7lHzLvqxJ4YPhtIs9Ca
kOSf/WggY9r16ME3xC+CWaMQB85SVtbQcFLzJ16OpcHhKgeUjlAkpF6E1kRhPOCp
9kaEfll3TGycMks74KMljzGbLjRWBMefIp/WcAaYurH5nROE5VJlumjU2nSP0vbd
7vB/wkhKx/5eejfsGoFq3tRpQJAbV9lZMW0hiemtMhZ+XXLthuDs00FvAO8o1ip8
K/0M/rByGwDEi9U9wWp4uTXcDMLOx7PTLqs265k6GpLytLk6942gAtr91kvkAf4p
dWj9kBSmEuGrt2NtNC6Slo9is9n7kV/dyeIGTPfYaoEDJ4tz9UbJs8luhzQ9k9tL
mN431sJjEHJirLb2xrWVI7FFHyFpdIKPiX6sfSRQN2jITKFY4PiyMnq8cn8leByz
VrZ8Ws87f64xNz2aQgSALk43w5WPhEKOjW82f6Ma8PQFM4shXWeP2P5nnUKfII22
0FTpxXcfLsc9Ozlq0Ek+p4lRURyEYFn/1sDqGrJFwvrteVdX80i0SOhnPj4m1VWX
ezwRzg/rKwd5QYkEioxLiUREaJfvISxtsZFNyOFgvNxVN2PSs5DaHCd8oBX/l1rc
ieuyDVBnpohKsmcn4DydPl83S5OWg+IGb0H4HhHKyzzIjHp+3oG2yoDHV3RhBFKQ
6oVm0APmqFgPUbzPbAjlXNvAlJGiJjSTPaus/EH+d1fAkeaazkYuequzN4FnErcB
/uYx9RR+5+Ty449HP8zjlSYJTX1JIo271SdSH/HZeNImmAm7TGZ/GCGla8GHKFja
Hon+YAa1SYoa6/+8lKyyyB5vYA2AeH3GrD3khv3X9kb2OmqdRTs2LyuIOBYuqqcd
REFMU3gNKLi/5u4wk4QmZqY4gM74MLUwtABB6L2TslHdo6QFMDovkjg+VBTWlG1S
U8KsLCpZV+cAZOIA4rOPkdzwsGLA1WqjHBLnP3vfeNbekZbLRII9wxCyozxnj7D2
lHcZc8wEnYPvbdg5WUBuTUA9LbyslpfhTY7O1qqYzNWp9XIQJihiRS3Uo3ScZdTj
DYkU2dz0oBv8k7rQNqzCKGcWwV5Oe1Uc55af1n8IshqOw7M+zZH6+n+kgZLlCgeu
2X/jZCnrg5m0hPgm2o5I1yzf8/eXBe8tn3MlKqDGCVZv0rOPNEur8hS3CTylMcvH
BmnF751S2gMeCmJ8rW8idnXOYOrsjLRrhbZJEPvlSUHSUv1gTCG94cTvlJ/bxtTh
ZzJviwPp8D/ngLJmzdkTq+T015wWIDGpwmjxjS/Im7Kspjw6C6+yPKjj7aahHWpJ
+8dQt+cMFkDZ4DoYuLj+DVu1eYcpKMJFYvqxCQWBM50V8fnQwOaeN/5ieVcZN5Xl
e71aXceEOCzsFcUuXlag/10+TQC9pYODnpjJs3u5K8CuJZ0sdnsLPwe2cRjNuUFx
rIlvNlMb7XXYeQvvkn6J0WPcuOXre1QU6mIjAzEERaO1jqdgGJ2bMx4/1EA1aDrq
YJMA925jncPT+/ijbleWQRpFnrhmDuzDHUcjn2I5e5MMmVVxVhAOxWynRn4lRPu7
Kn10znDOR4MSUEdJe+O44nynD9sshZNLGiJXhXp6T6K+jhz8aY3f6d/1m+0QbcZ1
MWoD+3l0Ao9gKRc7/9SEzqrOjGR753Ofgz+Wh0Dc6QcUpPtSnvKofoegT0tHWEmt
+9JDSySb1B2aYfu3Vy5kFs0VALDgJmEQiKBXd6BAbengkeFws0mjeZbQK3UTQ/Et
Fis7rBGks2CxZiOsCXsNwiiNtirSiJZAO0ghzMkMbkK2CtrP0sSbJeEF/jLAkhVX
D0YeT4JHmaHH+1DIN1Noin7AU6CpmBP6FUvy/Gfey2bbN8rl/3g5GiUXQFPgF9lR
EXlijn+PPs/o7XtesDieObfHItR38hqLHHIuHd1bBzgwBTMjGtZYbMckN3l+LCDT
bQTxkRN6Za4OexgI8+TfAZpARGDPYtOjFEvt+OKJGJIwbfx8ntSSRENIC71K1ar1
mbs5B0wLhSzzk2NfaaK1u5FCR3vRf1JhRmTmrHaGrwmgYnz4T7w+pY+kpFoDAZc8
5cYQEfPuEt/sijEqyoxh1muXho9CeaaVyl8qoZBAQVZtSnGwQMLKqkfTpa6On98C
Hk2xc52k7ct9CAyZFs8wKxYanjNPu7ROq0qd4wjZqKv3NRCFyhDW7yEEIRJ65dZe
R1BAxZgjseJIh+a+1dkyasOLjJswFFAKPbR5V1QF3n0qfFWUu2p+NO8lszw5PcD0
Gp+dFyHnWuIANJZQKeN1+Y4cHNw/av4r5La4fxXY21MbGahkoYSo3hvO4NnYGWy0
uyH+Orp+18HQnNhY+8xm/Og1gJEnpzPIymvnkOsa06baI3LfEl7ZmPuqXaKiR2r7
HM45MR4XGdm8VzVO5INSOWFazUSivEh8eVLc/vLqcSyGIcidUe2h/pqyehQaFxGq
uXR9+GWjZler9nxRs3svDmNTI6pnXos/UkuV0XNwqFq+Q+xd7x7oyDv44TSsgjmP
Vk5weo1XvMbdBfyyuV5nx8SGyD709tDIIdaFcOlxU7BNYUc9N1t9n++ZVijmpjgG
Ptj4QnCUI5iw71B0iP5UnD9m9ztMLFwdKQ6e8OlipdMxJW8pLbl3blKH4ZZCDBFM
k9P0r3r2hkSTwmidhACHgCfrkvBCHWr/6sAmyYV8BceykE9MTrsdjJaxid9qCmQB
+/bUPbcSCwavnJr3Cp37flEoFLdJm5li8iz4ro/UEXONQ20jhcjSjkdSnR8//4pC
DCRxR/PpUaoKIUi2OXBY1R4ZdDIKLfwfvZK8bHpy9U5UFAhnY7MrTJiKRw+duLpG
Acg81EVvPbeuMCldVrM0IGzRtv4gP5z/LtmmRePc3QVBgBEKwZmifOhMHk7XSirk
0wr2pdt4Ud92qIz65XCUFpzCl8k0vVbUuFGpn92jFVpRXdZTuzg56ZhFjjX6jdtO
MQZ7HtyftiAWp8ljcnTKcRplip2uYS7Z9Zqdq7HYrrjnrNOcja1Jmg83FGkdDEJH
o08jsBra51vb+uVx1JcLzuUfld+lSxcpxomozO5ePFaYoJ7qTQHrgMfHGYKWIVNz
nLek1/EickYzYz4KSfU3B7ClDYZugKkZoXhXXCkpCHNrIGGV5Ns8rMCm8qcbnEAm
EOkM3K+HC5c5kTgymOweqPZVbzoj0FzI5CWRWBxG4MZ+YKj4LFk14UYQ2HjSXpUF
pwRWV7+ncFrmQ39XU+P43xhH1InQt5ZVwmePSHaFEeEeHR3gFIV+oVwO5/ISdoPs
rQ/5S4ku33swIYgw5f0ACmlD63GyiKtOJ2IdnxfjFlqeXG7N6Ig6u5a4VC3c1ijJ
SXIxXoJQQJEvny6PLEnxKq8Y/Nos8c5NCQPo0UXMzs4KFQD0/yx03Lzt1otZtL0l
8bjougcI2jnfxthzOkt00HTIPN/wzQ+AGJoqUa7CqbVRRVE8w6C5rXLQhgX64auC
2FnNKn4N7U7AwxoAa1WCUVkuKrlQnh60J8bSo/Vx+Cr1J5M9iIJx8d8iMPNTO3Ro
9Usn/b3GpxXU1CzLkmYVJmZ094Dg9vM8Gb/y91kiqjO9ERzTR5NzOmzakfgvK5W+
Swezpt53nau6NiQXQO9BfkOjyhsnBbScsl7GfaEsetCwdemd6Ir1vzlvdOug09fx
zBFMpAz9QUXJDIQdVEaGyYSmsPvq4nkZC30HKHIiwEPChTshgfpnac89mIWp9KRV
6svHq83bIAfa/1wLh2Aad7xRM1C4q3IiKu6GwHp/UwftAsx6MalIDMQzksOKmqTf
aVvRmsCI22lX1ZcfsB6ZgVDKEwqIxCUtsibeLE/F0+ZlUCGsKx4ZYhAlMAxNRCRs
N6vTJ3ZZ7GCUE8+LtJ+JuW1t3HHa30k3Uzsz+wQ6GA71UbjQVAzQck5wNEwXggX7
M/v+rJDcPd91SqnsukFK06RKqtWtHYLThCnOPKe6AHZQDIfmAM5RVF72l5OGdkjy
Rsx/Q6nORpZC2zYiufaDguttYmyd+kLaeQ6fjaArj4/BlomVA0LJJB8f2R6+Eth4
DG1sHWgOE4KB5ha8pZxJlVidE12O7/bHydn0h3q18A6AmU8Ax9EhG2U8zGg2kvw7
aTquD3pN8wxNuCwxfKlsmZ/bylnjCbfEui6IcBR0zAzpSWEMDz+f5dQskzL6aUzr
5/437gzVijWL3LBLPk2MzISEF7YPfgwoWOxH6bw8XqHQe6w3KvheEJ95sOmyEBaZ
pBrDAGPzfpMWRydiM8cSMgZ45chU2bw+Fy9xH17o+YpjXelD6AdHgRAfEAsPwskg
P/q7c1HDeqCZhgeWdnvVCGdfSALjFC1hooAlnwXC7mIEGYlmdKELkvYwdXI9iZ4A
TllXK6gDUvFHojfhLpBUi5NeurhRFzZ1njYR3yBBQIheJYxYk4ahSGv82Uwjuz7f
cJ7fGbQbh1AW48V+1lViyuNobLJKOd6SdTS2HBDgZDS/uLIhye5ylaazgIGLTeex
k8MiODgsbDNdEUqRNlggNWi/ziVvpce+0TAhbTq4d99QhMMqVwp0OXVpgbaaVzdf
d+DCbCTOuE+xLri/GSbGVg342YUk78e+3mfn3ZcZdO50iC1qgSazwj9Z56N9gAnf
6oHw23SWaqKQPdgJckTd5cJeZjS8NCEZsae2I+ykvDqyww3ogsd20GH/iX6eUFwY
dIxintvB8d4FSvK/+vH10yvNc+oU9oA+o4ZA0BFNNEI6mnM4ppj2REtluTusDrS5
jiF8XCa7Z0NUDYDkG9YvM7Igr7U3W0OqbJfanDrA97WuXDcZCauITjag1V1LBeq0
JvEJtmebhFiR+j6VQ5K9b7tDoBIezXqUaxq+DFbgV+GZuHgjzkDHO+Wc1g9VFBSX
u3JvfFTR/wqCHenDKc3mNmrV2w/wPYB9fKV0cd+OucgWUQ0EzOc61+B49+a8/C9d
PxWmAmHxvlkxCM8WGjLeZAxI3Z1aucrZzD+9N5r4B+HjQPbZg/y0tMYqQFMWMxKi
UdJSuMQH9ru2WO7ewI0WD1sFLbGROvioJQ+5TrPCAoHV3pwpqtmGllj9IwFGZzB4
nJv/dxF/I97xkU7vzFehBsRS42eLgItmlLEicEMLlHDEIVBK9NlapID21SFWFz13
vWDcucJg0sNr7ngfXHR3Ub+D48u0vWGmA8hMBttbHQwIS2eYb1fTBLfFcxVVrYIu
C5noJ0rVXGGBKQLBqcwZZdk8RG5kXu4lapU94lfDRQ6V1EyBO0b1NkKTdfUZye0e
LJrHLuRuCu0zsg9oEioUYfo9OKrPiin6woSiK5kTkFtEy7bXfIt+A8R2pIVPE33g
SQbh9gn3CXDxwiUEEg8ItWEBVkrhe0XsTTq35DXMT3M5fDPtydMcm9GraaHqsok7
tvrSVwTx0T7cAOv/X/LpBojk8EZSQTiZsPwYGArKthlOVTfOO9fe5Q09ZH83ZoHp
mW1Wjb/XNiLTdG1LGHk5A3EveWMKnNZ7WJpJQbCmU1uv0OIva1GTxAafq+nGnBTh
t8dysaPgqF/z86YKxjkuldFOQV7nMz2875ddpu0O5T9xm/qg2LMgLISNvO0RJ2Ec
54i3wzNbLxxzUjzge4aaSwElVcWkOXc+QPirhIIXniJQwkQsc4xbUYbRlW/eu0Bj
vnndPcaIdzNRxodgDNMJTOMF2t2HuQcinG0i1ZJKhnFfOwc3aeJvlt359dkjk1Iu
qzNWmjgpzdlSzbtZ+0+DiHHh4WqpBuuhEwNMENPr+tVCFgFq39bwX0P62Io0/YAP
X4lVjdumTbMoSEzlgdTLRUnTF+3idb2u9+D075+xSO8oUtl+0rt23uNq3/JKTGUg
d+Or0AE5HpCbsVrmcMuuIp9wMd5EGusc60nJbG3HKB6mPNain0P0ZHuerilNNaBb
fCN5I8oR8QZH3/MffwI0bLG/B1V1DWZR4PtLALIJbC0iUobDgehJvNBvHsYzDfW7
dGfaW4yfVmj7Dr5WTRXWPWOKKxR6uEAdg9QR5NuBci6sVyaI8vMEELsY9yYNbk/c
J2qdp618ogCBp8KSjth4outbg5oVftnlEsA8x65vHCYncmCuQmKYiAzEu3dmCeXi
gx4Vx/FYjUCnxZT6mQsOUS6zRwvgi+sXj/BWEHzchGMxge7rN/1E2Aa21akrIIhq
7K+TJZ64n1smsGiWBOJDiJWoo/CigxCQuGC9LBCTeaaAVcEMFQvTOkQ6urVXVkdf
ELxNuNOVc7oig8vcOhTFqTiewd8LOchQdd5XiSCP+cm+KcgNt0eMhLh+ATbPIo9a
Vj0CAax8tgoIlNtAL5W6LC2Qp92wyzzSzALrCBzemqB13lhOrKpetsWDWwRH1SpD
KSmb7hepnJhB+inNpzN8nWXT/gYCfCuviKZ6EYPykbwiaUN0x0N/lw/1y8qfLrfR
6xknMSEPd9DB13+/kfcLHP6yGU7qh/dTHUvBtdInlvgBDp9ahXfYtR2IZbGcMQrV
s8bCHoR3MDGKUGMd/V7uhI7SallhZPSLuXbuSudkDRdqQjRkvOoA/lbKWTCHoe+9
XcJSpXyMOqJ1TlP+yf8V/ML6ssX8476fpkFzPx25sYeRzaPAcAYMJ/HPBtRrj9fM
0EYFJgVJwKh+xGIKvyWmxuokuluLDUyp7eW44bAqJuM1zQPz9ObAuKfNgsLSFnUt
N5s/vJg28xr20STmjktV2u5l3JKTHVyqrYGjqVdhBxW4K8q+ezvIPe1mwFusjYlR
z8VNpJZVVWkpkpWexuHCsd4uPXqedVis0aigXXH4zADj+F14EjmySgU5toZzZhw4
1R9jNgfN1wngnQuu8lQebmZe1fSDcH/JeLt44CvnvMVfRHTkpI3kRAdOxtEVCMBB
LLBW6+LT6yP7C7PSIy2gOEbjQUbG5UGTXotka+zuuB1/Z00OogtI2i8JqVZJ4N4N
NCvYvhWyPU3uggVF09opz5saDaMMwAGtQ0O/3e1XhYQDF/P3cXHcW9jzWRkEjFRg
huPOMGQIMTUB4w1ynSw90ttpkkZ5JXMxcP2FGTd1X1Yp+Or8VgL0JUl3C7t3ZSa7
cDOn1m/z3WzGdUAKlOMC6ir3GtwkAwKdfNUH/0y/iSz6JEFXL0YMqFRuufPfD1bb
NU3Ea+IblaHiv6M4gGu7v9EVeak91wT3qzEjus0z6Ixz5RfMpNtJEyTpp6kFsfkd
gEan3LItQaIMjy/kids0us2xdr5mao172S+6ZYM5oC6iJzRX2F409xJJfijoqmw8
aB3rOJdn+0l2Obazyzd4O6Daq61DCppVGwwfwWLOEgCRXGV7QpHvGVrCkQm7jtH2
IkpOFcKne+Kt5l9W8sqV9S41JDEfYZqKlIfyeeov6aXS2Z1Zk/dOj9LrA7rPxs4h
2YrYBFtI1/iXQgkPYq+Tz89eNaLBFBNlcq3EGnkgagG/jPyBC0tUo5jBKoXZ4v0i
o+XuuTfzT8IAmD3Foux6IYLbm5/AX8IohecVNARo+G+bXdWQuHOhoypxWz/wE1nz
nSdUJvqTzGfl0T1uoOlJNpi1d2XqCmjpsCCVMkhzweaVibz0G2ssfrQmsujVrL6z
kDD0lSwx7sNyFFjVrcTjjUv9QOjI2+2mkuG2733wZMOBNPCG/hw2j81dO3NxjRMt
FDukHdB1T/Z+E6fvoZ9hWYA9BuKp13dujzjlHNtOaKhy7qqIBDpx7PisSyzMjm79
SruYLhGgCTVrfd+/wdPP6jHqWBBv8IaU4BeQ2fYoX6Hkb8WDoWRyid0gYsL/Vd4X
ARDb/OzyJgGFwVI7g5sZQR+6gAqVPZYFI3HTIaoW1SZArYYdI9sC7zfXQFZjPx6C
lUhlgog94d3o5M32nybbkA5tN8kCU1tLhiYw0IwoSi/6i3P0SAOXyTjVBjlBI2Al
GDR6ymD83+jpTzpTInrFkMjCNBsfjaNc8/+rFP8Njv6+k7Ng2zlZWqnrUj1brqeO
1YsQZjDpIxFqV5pnr/sxQQZXKXpVe4VOiNbHxpH3TBu5sgveiXhodl4cJ2Zsrv8d
NT/YfIilFB5wQrkJkN1YjULjpeyQugO1tIije0oPshxTn09jhxuV0/b++sxnj2ZP
n6mqi84mZQ59YaWz3Boenw7M58UDtjOunzoZkoFMD/UCIfzLbAOUskF15xBUENjj
4WYcryhneugmlkyQYULq0hHSjq0g2QHyuTqVe7Bf8lTFtQB960vVV8Vmt7n+UFo2
RiuFhS4mGTKd45J42+7EtIEmy+3i+ynqwENIcEec4uaHPyIa1ZsltC3K2WBz346g
wPl+Cegz5xE2u1l4/JVkhY7Yq+yIW+qmMsib6WFkLeb1sU3B7us8mOGQoy5KMH5X
LfIslc+V7hGYeVBy96jH6iPX9zoZ4T7sd/IfXchVG1OEKPkwmaAZP96WSJD5RotW
ULaUxgCjvt5t0pbzX/LjezVSNQJUEJE+NVLFDfKLSTE918Dvj3EoXtshVjeYJn5J
pzmjQjW8TYoDQs/+fe/Cd9FUxNlliDIopGwiFqPgdUPkz+4OxZLET/d03+xwA4U3
qDM4t9yoT9UcJMxPd8us9iqtKC1jO499gBFZAaIy2wwtelJ/MYDmdh1OEDAWgN9e
QEjtWs4RHrQa20pNs2wBH+n27J9YIOxoxzv/kyxM1l0uhtKOVeWgNSews1pDiE2c
08SJbOa/pXPZdnMy0FAJVzA0KvKW2xwyhUkoAZY3uhn2Yhy/FX1Xu+4l2aacXGlR
BkhH3IrHMDLeaWrq5i1JYI1pN67roaYjQXqQ5+Nd+BXf9Rr+Z4jfdsVanCOvZN+I
mMJVzaRO/1oOwUAcnwwrwV1kjCyl7otUmVfOaT3FgGcSH3+iO5Ig6kRAcLHZ+y8x
b/TdUCN9Yt2ytcUN1GqlI8uhNpmMs5sqFNp6VktF4Q33SAHIlo6Z9DSXBJwvtxNo
jte8I/toDprn6n57c0Pr/wsvRh/Z1gNhRz/YlWB43kE6zZM+j941k6qc/4C75MIn
4+2vtg/EfXzx/Yn2QshceK8L0PI6gfX/tYUuxX2H6bOuaOg4kGaBHSM1F0gv2WxI
ffpmMYpz/FsSbMo+cjHw9zHP9Z1NZ9vHXyS0CkoS7gLz6RvwbXQoOxlIZeIl2fSP
wmZkJ21KlAAxVW+mqgBGcWZMPaMzvjMwR5hcckSWKd9CZ/qqb2eP3SBG+GhmZOw4
hrExmCPzprJY36jzNtkn9qKODAcQv6CGL44Z6g4Cb5Quyho/J9nNpLIb5rnx+Qex
htp0SvGXQ4CckBMSG/J+Mk6teKL5ju1yCRdLVmpGLvmQkiXfqP0xP1h9Wxs4CyOk
LOk5xMQO2iMaWkv69a/k4v6UbLiR1p8s8E0Z8Wy8e69jVC8H1p2MSUXWC1/zzy/C
1fCfeEXAfWJmhFqfuIDkKifT//1j56mmapPgunDHGdlPT3p0uM1yUFZJk1RvsaKP
XCz6yfIA83TBwDniujMc9/6fhykBy9MMD4Jw9f+uYr4FfEVrX9khr4fqVp0+Qw/R
aunpm1YTlVGZpLNcoGgQKDwLaKK/VfBPSAy0jLVvmsfXE/p/rsVPhhbIPl4SQoqF
2bPIaaf3nvkPQ2Jg5toNYAbqNERAZplUMLa5vhOSia3LR0zilhWlDXT5Q37117Um
huJrsRzLzfRb1K1HoI9RT5JhJsE34IyQuCdKF4oOUW3i3C+KEQ6zE1asp7FAfWhd
y/dW2qln74mheK8dgZW62VF0kjhcxV5s+jxhkPZjoPR5vjSqz17X/A/Z5NVp+lUv
5hHh5TYwPcl37fOjNLWNd8+v9JM3QPOwoCvD1sMY3OixQLByGLI5LyMW1ZeNQapd
sSOZGtNvV+hRiqaO3HIehjYw7IcySCvqiFAUwftT/hkXy+jN20sc7gvPGbKXkmKV
tBqG+6dxxlIjtXsL9IaisccIKz1seSS+hPfM3eLlF4MchlBCgPNJp20xJE31UJMC
QrZ2A9zCVFynwLCJiVB8t/G6lPgrMInWF52denu66BebqtGPPtfi7s4CCAulX+cW
rWgR2Zoc93fvZc1u0NI5qr30lM+bDcTn98X5CsyzVhAhkD88SJNxodGNKtimOLOS
u43JEOWxu5lq9jY8YCmxyS/wbie+9Za/wulOPqpKRJpkIKprCViLrNWZKD1r4Qf2
xIVPU11/1LU5Ei2d8adL4WlsrkoySQZ2fW+CukMY3714twbbEM2GLiVy0wN/Sz6l
w8ZACB1ufb5oCzahSMIjcDbx+FEhttUwkQuwmF/pST8u8e6k5SaIWKEd7fa7CqPf
6pX5W2qnAEeUAZEAJLJQNwXpkuGwM4duWTscV2k3EI11bwUNIm9qAKLNu7UsDzGQ
+F/5ruFU7vEsuykDUIaQAwMecV4NWcWeYErCzEvBpIjxoJMvU8AA6vnbuxswpHbt
7TNf1j/uKNhxWYWqhtKRzfaMgw/0VMvnDmxy7srRb8btIGM0Y59Z1+BGRmcNbpWk
bXM7ND56ephuWGJ5/njXN7/L5EfCyOLA7d8HuDaaIwNVSWfcyu8uivAdeGQGrjUj
Yw/pXhPL3IoO7Fo0yBfJLiSeYlXI3gAW3PRQMGM8pbsDxf5vHXZ7XQRXTyOCuZzt
iy5kO1o14cHYTixtb9Lm+5zKIs+h32tSEnx95On4lTVOlJAgORlG1VjTgOp/Yaum
wizI6u7+tzFD7eEskfE08mejN/SmSedFPKRkUvFEzOFKI2CZthgTY3NC7w6u88aJ
qC3qBbaMxCElMTVOh0lULk5VsUOzdj33DMvqHZI5lARKrWjypoEXuUZpjzFODcPt
UCVfL+I0YGcYa1+DV/vlw118jNJwdP3Zdgm+R58bYFWytRRfIde6XS21BqNXWLFn
d7AYAvXPjAcjLqC4BUAaLxQN2d9+TxYiPyQxdn8VrUkWcoXnHvOsVzjReYTcIt/P
/+paalrwGyq0T/UksadlXG4wDxwQgnLWaCqk1xv3VAD7OZ7wYXNub0Vl5NDk0nSI
RDZMhZaFfHIPDv9LnjILt2ZXVV5/g0IW5cJ9XcYgBw3vvJGXb+GIl0QLXEWgvmtp
CEc8BNVbOuyr5YFFmuvA2af/8a7V9w1EkOi0MKxKFJDJ9B2TK200Gx3R+enhR1/S
BzjjZzLCyrsHQuDGmycIzwncfVLSj7ZAY58NtYsbHu/hRmmPB/1PAKX7m13Q9ehe
a6E73lEe70gkEinQpUOho/RuGWouuJgYFBzpKz5B2CHaVjAXN8snB8h+Eidxz+iW
6VVEADfBXYxEyBHmwFnaAYiW2sCuXrVio0OaOv+eNcXTxfRoitpN3KI0aig4YgN5
EB6j+6ZzFU26yoiFrVrYyLqVyXKjuBOd/C28CKwXcafkAU5NSLsrko6HeMF69RPe
w3SXEX5XgOa/AV8gnlUM+fblPZQvDaO7EVAF6J8cPrBrle8cUNzuK+yDfRrLH8BW
LxlnKGHFpZcIMV678o+GM5TIqO8b4lWizL90PHU0Gj66oRr1rLjCzB6+cUtXepBh
BYjEEH4/tzfSkYNdCR+UFhK68QAerscOysKBe5NeNdTNXYmWJrEs+vBKZJ1MqPCe
f4sISTmAvHVsuzyaA4Zq0PJYyPY5qcGOaIYhXX6Ti4a0FHhj4+zkYoRj0L/L7cEa
sutTUxrEMBvUAcz9SXk0VkR1bNaZAfB17KV2sj4IGnNkt3hgo+GrTHbm/u3b2ncj
40+gSg3l16yE6RtGnhAqSbTSczGvtEav4QB9eHeS4WJdhLrEjORHfhY340+Eyjqb
RCmnMSC3sRabF1uuU5fszAtPff1kNFjW9IZizJOrVKb+vQqZOCZ2aCi6ftbmX1c+
ayDGTqh/mJ7uyXCYc1AmMpYzrq3Q4K5nztIqOQm7ltBt1rsQ1lpg4XDBiWiV46bP
83jzwfMA3cFvh24lTTjgt/yY0ev8PQYiiW/j+ozpsqqEnw7AfAoG9/8K4quE9KRG
JV64Mu5uytwdEBNmx71J4riYUqgslT4KxHxxvtL7gkw2dMrSoA4GqLNYbDV9riK4
YfN/HKvbPxEaJhxTcLxv0+4k7K2i5tR6RPCSHzKiDoWJwEClFFRbVhIDDSGxODvC
SKg4Tdlz4N0qUK2xKPXV7uT5HkWC4LIcmGM07w040N/14WEJxOM+xxkpEsMbEFur
Ztp/Zg/n/SMIeAaFTFOcn6cjhsSBawHcYyZiTDFWm1+wwr3LldGvPnD6GxJ4PkRo
51rsjoT2n7t6BttGW4ABisov7l9acJgK7x+ZjIQk1rVXnJ/gQGT+a0VaMIt3D2sZ
gUpmDH4R2qq+9ae6PEq2Uy5pdxwoL01CcR/+v5aP9bz+fvp05Ca6qtFfjEdGmAV9
0FfhXX4oXTOzoIWNyTBKxN/1rry0q8m0GHjiFXSEWd5+mBinMstoVtzUOA/ItMfv
uLQT0MsjaTKE1Zm+FNXllDPHnkjs1/C2irMKtzLEYiv31qswNjpgZIM6bHo/brFD
JmV7MzKM7CKABwNtb/dW8Cbyo1e3X2XJGaTNicHVzB5kPMGdN8QOrynCmqHIt6fy
LYk2U4bqEHVzUXL3ei/39AKNMdXkCZRu9F94f5bj4X2umdEffaBzg1k3s2BLPdxa
GngaX7/G8ly7z8OSPOiUlQXEU0xQNsFRsfw+CNqxO29qfAqUzwwoRsSq8EuySxW0
4vGjxLquGp51FAwc8HJgE0GUuxusKe8/IxLpnCE8AnShwu81De5OeVGjseRwrVkE
Pb7yvyxAEKwhIfQuWTQWBEuR2zsZV60w2EzVaRq0zzIx5yTUBDPq8jKT2NTRAnNb
oRRqhZaXBKBx6+wBwro9TZGl7XPnfskSx5Xmbzjh7a8SOHrSJYUgwgY+oD71ddhC
WKoZ+nMLqre4jU1NRBSx4Ab8LlKnqU3IMtF7u9G7uhkuM4hV1yDDbT5q7INi0PKg
hKhUU8n5DrdMmzx0Sax6vuoNVzqcyPoa8g4d5UqRuGFvHqnmcPNlH1pZAlZE7Y2x
5wTNzpNCVwtjtbDjKargZkRtzmPCphBsGLiheKM8nzr8QIWvxX1UjYyYf5kL0p2D
S+iL8uwqAXSSkHh1HiWmKrovS8tw4i45c0xZTBMe3DuyUDebq3z8EBZfyM16XLK5
kq2U7tBMDhQkXBVfi/UNAmT0FZ+McBHvxdWhDhxmrXKogaXfpWsQn0fCchlKRSzr
CRyvgXb+3jG3w4KKVy7bpffvcsRzYy6AOoaoqEATi/IGN0v9S0Dzx7QwK4OqRVVT
HFIJRo5z+a8DgBTEHgb5BlGymfyqWJL7aSmJ5axlukzg5Nh9pYH6tw7CZ1sNCYlk
1hsejPoiBdcxubNIouxczHolSVd2QHaQUqEIOVt5+nNnj8Fl6rZOslvlHGlHkEOo
fj4X6U52P8Cw8cha/ZCDHsREyH171IWkPkZFLfSfdaIZfZrOnVRG22wCHxyaEflN
SVHATNS7/Zb7kMFsFuf69HNV+E6ubRjKng0yTkYbwG+poQAk5vBflsKcKl05zeJb
AKjBJn7bmMYCY+8iEJiAexGG2D69KJny4OQFBBwScCSzT+Y5TPs5uRVJX9dxN1Ab
25t4P8AcX3nMEpeYP6HIIihWoHjuI2vNtaNGE2G1BRSsZV7j/+bC/FSwe2++8Jah
Glqb0qVw3CXmHqIucSoD6VtaykMQGH6olH4XDYiWnBDWaEOwJ3ZrFn4IqL2T/eXZ
cU5t6KTGMjwhUC5K3+oGKpakVa/3jKIRdO7pH0hchoKX/x6AvvDQE5damoaR/uq/
dIuynHZGpIacjYJ/QEQHYXLHu4O3rUdN9nu+lnoq9/nc/dp1wn1kZf4C5GQGrfAU
wgByrS78w20xZCQBEMwX/Vg+NTbGZL7mkbBo8CVjXGZP+fcVLzPOzdT2Zw2/xOfd
xdKThcFCMMwxL5zq029hKqdRwvVV0lyn9RcUwrAAOUhY0q/SmP/KjcuubfUGAWFC
6jr7eOsWHEwlI+HJj8maYz8m1b75mNBT+oo+ECXau7RzVgMjX/RlGYoQLvSGZ9IG
Qz9k3UERRe5/Ef2AHX7yqQ5h14vUPDMP6b1HoBDBc4pJls133TUhW/0TCnOMA6j/
LsX1nCW9WHOdVXmbEFbWQhGi1GJdUa9hEgrkl4f+yZb1h+lKi4o//cQlPT5sjrbq
xRfQvajau/fEo157MzGyqlqddlH8l/Qsc+PUCVVWaSMqBqxWCH9xlkwx6/O5a+TB
je8IFm7G3kuMX+w3mlarb+C9BRORTOJ4fLPBvtDC5F2WeEo/IaPLz6FQ6UWawjaQ
qxN1skaJ52MBwgY5sYF1bhk3o4NoUxdcHVWC7eoPe0ITSiPhEQGKryix1w3Yc12A
8wSaoFpoLv0HYAfjgh+iHVgICWbm2b2FQmEvHWU0XJmMpSkMwcD/6Z+xcNPsjUaJ
elqRfxkksabQy7dG99fJ2G9B5Gj6qa5TDPLCqE09pbKMHPcUzZNQNibh/x91iz/r
+lMFJx1xH3r1a/PyzRv9jNikjUaeuE5YE+Au034aqumcAz/T++1NsOkl08wKqbQG
Mr9qTlg2VhejBD9y2vRFMPggQyYbMKx3GcL9z102gC/R0uOibiwtU9uqscB7DJqq
h6Mu/Y6Ein9/eS/ld9PVCpiuw3z98U7bSpxPxSoZrbrDC2VasAR8IRyEuAqdvXJ1
9YkMWIDpcuQ3c9Xeu1fX36t9m3VD6T2XoDBQlVigQG4SaNoiKXBTXw+TyAcr9wdY
i3vc8+BknbbRMCo82CA0P2+7EIPwHGtMH0/jKkOsRKHivFiL/Ak2l9unfro2Y6oX
+mFXxvEPeAaC+ITLBshWPuNroqA3fme/KJpbRqRMJf0W2QYHofpJUVLb5ghItPJD
HN3CikSKEZzJjKDpJQhJ83w3cYWNGGrEpoNDkdxINvwUPlw3svoRw0i2iIN7ZGGH
JCK6ObaDC6qkoRtS5/MM3AHuNyAKQ3kRFriWi84kPFWwabv3UM7V7UM6R9oryQTa
dp/rGIBKQSSqUHHoYTt02NjXSbP/60FhjRaABvZwgHbL2Ok8nKd667QT2EV0SGVm
rOD/hpjFegMmgVEG8lOnWY4s/b7admibbKOtP4VZVb53+Jd2xfVPJ3rd9TRlEgl+
sEt7NXYtubev0mu3jCkxR1m+MGqe2Y244w38vsHxkuUOAK/5VlF0LaYyTwcnSQ2z
WZBphQVOJ91qDp/CYEHeDdgigMuvrsUX5d+1eQZGjEFHrh7h3PoTBmmT1pjkT/6A
DYc4jvvzonA2oJ8jA/d2GnI07jAb93ScQAF80lcP6Pc8OYsAAvEnWiI5wclUUWHs
I313ewXZNCC4oNJxiV9F9ilP8mA++PyllFTkeH4YFQeN9DDSgrziAtpZgl8dzxz9
MzPS0DMsrDVP/rTi7P1agf6DuOSYqFTc0CRpD4Y4iii8DoO9utSNtUKE8ghuQYlV
2X1Gd6ojooaiSu46HYY4Q49+AatfoybJSS2qnMv+WDSO3mUr/efHNRqgtbSmQJmI
eOH/CffF8lkkAL2I5zzCbsWt0KEB/RC0GVCKj9RrBhFREoiX/LA+wyr4D516vRH/
WGdNY1zHMIi3i0KwvFr7UBR5qaVC00A3aJraUbpdPWstr8fHw5i/KARJwXlX6xgX
k3EO1d9bqqc7GlhiX5DB0o1ZiLETTRDkNAqK7uhzn22PYb5bozDO343S7srdlIgT
xFwsxfatYLzDqpl+S3s5qWgJNEuvPqF8pYBZU9MhH4E+b9xcglkbhBMoxrGuthDr
BGIMhLwXSlVqZOSjt4c1PwyJ6oK+TQ1W/FJi5gwvYn7ja30UZzC7R+Yz4D8sT6Bd
NRwg3gAx9libcs3yTEEST5/SGxkZ9OJRXvroegz+kaT0ET11epnngQDkNlC3o7Ab
P75YXkqB8lcvtTZLb6j4WEnuE9zaQYi98Ie8Q0seO4o200S1Uy7/N2FaSUqMOW3A
Rwairo+YDay0LT+HcU3qoEW3bLNQ09BTE2rqMGcgA37/rwFR+nQV94VxgGERLmgT
XhMDj3xEYc0VRqW+YB706GO7oYXBtHnV8UFyy1vPCXbw1uZUhcOlwYlPgTpgTxcV
macjLaIhMbZ4PbAV9azhPF56PoNZ6EUMvU+BLubbQL75bEGBzVs4FAgKYneBmSZX
xriVjX3PNg1W+Dm9Yna3bx2qLUNhIKRqA4uxojZuyFu+gssqY2+41+PLr5Oedgya
rFcRh60U+gVdfemMLUqKOx0iuVRMpPfCTE6GkOgQ4+X98Mpialvm4+sWXl9dmcZa
jOU5AUlSWwxCT34Wlt1+FqEvPqQ7m0Pna2gxw6KsPdiNMn5OPwBq95SaN1D690x4
GMBF/GE0qn/DXLCt9byr03+o7S2/L8XiH7C0/Ye1v4YO1DnuBBZ/24SId4QmGhW4
Nxz/uI7lMBG6TU8SEIJMAkEuo+GYiyfC0sSk8P2pXB5ZoriuqQ/XR9SXa/+fupE5
imfPKKQC50AhnSu7MT90E9T9tOrYJvm0QbZv3hN9A/ErCcBMG6TBaXKZ1BrRclfm
we3Z2rs6aRBaRw47CL3Mmq6EjC+4pW3PG0pF7EL+gTuCK+rk6fFikmjteMABdlV6
d2ko9aTNwWXF7VC6WCK0HrM1kzskHBbO9nx1OJNzQbugYBCu15DaObVOhdL7iwBw
F1RWRLAVOpOUo8B1CXcddeNzmtz5ueTKsRvsXRCoGNaR5gfMsosEski9sTNoToY4
ZyTK2KsUDz/Hfh+bNx6vIhnwvfbO7I+EvgSIvsv83J05UTikPVWVeZrJ80/Ac8BN
YV1zhKfygwlH+/XXNz+iJvq3Nr2oKTQXRmd08wCXcETLDAsvUFyyfxW3bN49jdue
Tf+Q/ToVH7BsIDGsA4HWT+S/wqkGMkDIQw5nJqivpzmz/8OWT08IRWxTpvWV6I2h
DhUTMnAG8ecD4UcGf80dtKR8abvjtbNaS3T2mBbUngOh18gTitTkJ+Ru1BELBGC7
NlPpLkEWReFSnHcuQayy8ZaApsOY+eSJm2uAxnbTStG6TAacqogoT/suC9X5N6TB
yDJOwEA8Fc41zxtm2kiG0oqf1OPMnqQBsAiFBOG0QAQ2JAogeDGijNuCAys9H+nN
iEoZkcRzGP74ceDnzPbLYS30vixAMwqwKJUbfYojxvRpdVOo8S+xwwYGw06VD+lV
HWXY/ft9sroTPwDG/4cYKlFLOIoZO+bSrpQEpRvY5+s/7JnWcYazhdxnQgMiMEKH
72Nfezucf2yOlI2NRXQmNpWraivRtujMgMATnm2cME1aGhG9CTHl+JCyhEQIq8GN
ja9p6G9orGtf+ca75SQvnAx1rpPjtpu7/kwzFBN6rQeLqVfuTh/EfviBM3a+13Ki
0AVjDoNYwavkJHIkv3s6hdGsyhXqcDbVg3ZF4NMPvsVCl4qkf/pGl79o3Y3mMlWy
R66egkFVB26e+TJnusQ978y8GHGWMr37e3V6atBaBediLMc+OxeFZv8fiLsb+apV
Ga2sBQTE+E9W+TGyQkfkMhphEov/a3VaQwco3CAo/SixhFfAyV6UZ8pE1x3qa0S+
iFDTta7wdqkJWeyDfnaB6KEiVugMerHKYX6qAYfXLSoChKx+sZzNg7+83KjdFTGE
kDSwp7mI+U16yE6nj0IdMBUysSvgBiu3YsCUhvAs2a50+DqyxnUJRO6m+ZrGADmb
DCbIEqJV+gfP8v6XPVioHIroiHm/1yihXnDYUBOvM7UjFuFBBdhqJ2aOpOmVvCot
6JJJKbOzg2SCYLa2NP/FmiUkM0/NIxj+iIYKTCO5Mo9k3PHee1QNupAErS1g/xxg
Zro9fGDJsvXVYywZOZBq3ybdLRpj37R5ijysq0YTR08zB7vfcg3OCIlDWXQxuqIM
ynrI7CGpCVd96Rn/r4MMFIh6+6Elu9TR9rNWiLak0+L9CduZNzqjKC6UunIP5pXS
QAd7wqN48jotA6FSMZLGl9kT5oulOtmdmkLApn/isFxDncPLZuCcYb/nr5/SgRov
ooRX3ocMPGGsAKXIgUIOJ6xKEmpu3Ltlx12X9U09pLTb+KTjAtjJJ7ZKqnEh6VoS
o9zIHPa4YOMxKILQzfM1NGo78YZs8YU2NEN5iY9YpGuhqPsJsAFY+y8KrCrgSu23
kQSpru9yeFQf/xuZJZOOqqKLVfYGmTLW1pBeGuZno9QOI1tq1dWl3mmJpKV1UnDX
V01kwWjM3vyJxdkCpIX9hHun2q4cb9p1FiivPsD05G6KArOmkcm7U7CTD/M5cbHR
kiH7OldugVAcaN9Dgknl75C6oVKTPNMrywSdTQ4Qo3xsvAkrpxxcoLxeOKZft5nQ
w6qoHVAEs34gb6x6uHgzxu1jmqVlnRzcryE7ugUf+TEkKQQLSTXlOcHtylPsSrmf
x4yrekaqvH0otHdGIXKfnjJyJoQ6rGbYqvSD/fO/Ox2qd2C3tsV/8E+EN93u/aW6
7kXBDLdmrJfuhum015CGv3wzxVGBGAHeI85/O75/YfUEc71vb0Dt122Pu/jxnk/j
Uc1r116vWVn2aqLCxq3NbLSh6yMTgZYs5lUOwlvEu0+g8Ia2x/Atj7kxCQfKpiFi
wr2idBrjPRFSvTJDK5wgDM38kgOqILraE/j73tCTT5GIESnAc7SFuC16GODqQLcl
dllDWpwfpFX9H+iv4LNktYeigGxiS2B1SFav5O6zClbBZLqnl82QqX/BpuW9D/J9
lsm4SReSSrVGdbdIeTmT8TzDHGibYNq2XMV8jK1o7jf7FTu4XXlc26eGfCKANuVH
zNhIBQx5sF5+rmozCEN0fz/hyeUep17NP5f6IFYaBJK3pZ65ZRnjZvY93Uepz2Yp
i97mDoYi1RIcd3pN7cBd8xxEt/LnsBZV7fPU3T2MQ3E+kCsrYh5ca/l9rISWgyoT
5C65CQ629Feg5glGJcdXsxJ5g7+OHOWEkIXAJUzFMLVrBPNsqxr+iPl0m2NW7o8a
nPPu+qZnv18LDPAWOmMKwCvpXk6sxQpTH9lccAmM0WQOJJtoRN+K4V4llceOXVeQ
XkegkLaIMs8pnoOVfyXNwG4fe1rw2fokNMQf8U8H1ZL8Mh98jNbaZ2kcvAoDN5gh
FhP3u3zbz6eVEOT4pFrq5KZb1CtEu5kNUZHU7oGpojn/krkJgmskgX9tMY9S1I30
c1QuPB2YomwvIykrtTX54CwigXXzzLeLVKzTq1uFH8dbdz/FozD9sl82rKeSLoUQ
NMsFkrFf52WFvxmn4n911U9vHcjpM8Y96CuKRExEhYk++pDTrFwcWfdephYG74zU
6QUmciLh4YwkZynnBp2baBOwadH9l7ZxP1IcUB8KfBEbReSfAV9blVothyb/2z1I
Gdtsz/h5OU30vNzCi+N8qI//T0aCWFbQEGaOFHRlNhWYkguHjT0UtA0IKOZ0BUZG
5Myg9P1LF3JlquiuYnK6lIMbGfYywcJf2XHOQQrvqzuGXmqKFlMYzrJw542sUCh5
FwHHNAuXTNNq7sj23UOjhRBv+ArBag08eltQ3katRkwgUK9rDGeztecBKBH8Jkfs
T+nRfs+H9+7oVKyQJikPCFqAvLZqe+75OTIvsEc+LmJYckfZZtJnqACj3KuHIbYx
Yv2XpcxE06eHu0DiWmTOWxL4QX063B+ZhhlHrduAX0otj+OJQAxHO3nXxsUe0onM
NiqHAp7faPhhBL6zlvkyKHg7UyP0AeSUYuYAqGQQYE894Oem9imUfn81xRXsMqby
c6ChtjI3waONsXH/UQgX9U7ARS0DOjAAigu5SKZNulUeSGgffYireovJg6FWH/mN
hCFbCCtKwh7R383KfYokTI3UytpFp1FHlCJ2ByB7oOI2PxnfDCI14ux6bnmXjzbb
0ZKsYstnRkzo9n0NOpjkbUg7XQutUcLnGngypwD5Gvklcg15otdb/FoN9sy2SQGa
iJ4csgWmEov2JBKDXkAp2E5gD37tfEaPgK6Lx1D2Qwgz7u/ePO+IHPnm/mNhqA6i
/Si9ZIbGmEshe1VD8Up4TdWr8zS3yt+5x02MT+s+tQgWLd5GsZOBgjU0i/RtO6+O
8KQ4d/YlAFskO63+26QKAX+QhY3u/DSEIrPBBc784+1uYIr/Iy9WWAdV2vnYOpuC
4Q+kf1Ies3iMoyNQGPh6JafyHzcNd+sqIcHYzP6DRrfLyB7vEi3IHTOcjG42wLRP
gKpwu5udeKMbUXtWM1QgyOCGKmGgTQqUlTzBDm8b7yokvUzPYs+Wih2L/TuXWzhc
FsCCnX2Hx5/n91qOoJ2rGtA+2hemxFj7IMW7q/WFyQJfqjpuWNzG8ah0VXQtnh/R
oLhsmKEDyHhmGTv+2meRBkmS6WnlQRNM5pyKc0/j2tdfP/8QimCLHBW9H0lhrx/+
VXrINqdoAy+iK81UsB2D8EJfto7LRIGUJ2ShCp/u9ZrfiDvspl1SN6dg7clhlWvr
50puRWwRUBRAjak+B32RTWpFPSuA47+ljRGsFQaoTloAbeSUGlcEDjma17Uf/PM0
+EH2zekQH3FOSpBJvQtUwqxz8J39MZrfq2We7d0/Sc46x/9wf2/k5sdcDfqQEEqt
yeRq3Cfqr5qiY8EF5Sc6oshewQHjXl/6W6tAxY0Xu/Qkm5UPC27SAJ1xkxLeCEzT
RNDAzUubdIU1HkhTem6WH6xu+EYHKu/fH9yVomZM3zslO5C1izWUxk5gZY2mLFLc
MjQm5rjWElaT8elVvGRFUhwmwB9PRKqIC6K4JNL5lj9Mz3T3Ed6VpxLAABLFvHO5
CfFvo2+xbt5CHwoNo/SOn4eTG+YC0tEKJwxrHCNYxywHx2+SJi5dcE6bPe4P2gn4
74dAHrebul82qemcVPBnP5hetDc/nqrX4EZqP2SXUaSl917WI70xGkcrLZJCpMmZ
yypUlGyFI5XfMCmZM1nqVulztuHXWUX7gena+9TfMvojFEEprwWe6234v2tFpQ3I
ifIB9BFTuw6Kde3coe1eyPlqxvZar10Vq9bL3o2rrJVidLt2y8rexjpcRnCckmkP
ZJabF3+WMqtPk5jkqqjw9lVzMNskctxnXh6ip4vxkVl3w3WuSxH3Z7gPcr8yfYkT
9DacCzT4fTCnA/ecEe4l6I3Z6HfGsxHxgs4ZJ9eZqpwV1X9w7X+6hjeh9yHw9EmN
1G8+oV1joBBcItA1Ysf0ZNBIrx2X7NGYeN2qmBqwhbbwQyaKZU1uTUB5tPQasHjP
lT+CbyKI85HhAyZSof/UV8aWw57Ut1YXvviEHR7Am2ic7T2My1JWf62vTaNNtZhT
gFHORMXi4oZvQfgRg13LG3OvKe0fOS2P2HN9HKSFk6JhN37K2f5Bulzgh04cpM2o
0R02/TWRvQ+TyA/uC1E3fYLI+FsHOHTQ4XfCtimKsVl8pYYVLx8HvFkHO5dAfSpn
OBqFHQe51JmUs3t6gfkAiqh+F+fQ6BQYVzUZN206iMcfYXwTY+ADE6TUD9VVbkTQ
phKd+epJ4GB7e9GvguqijP2iT4EyNvjxgQ2HhQInH1JJMH3bMKW9/1bKhnpAPlkT
WJNTx1PMTRki7laet/jkccRG0eyMrbh2+ShX4/pg9b03ziYhH1lszCCRL49K3ATP
v7fgi1cOCLrTFwV2zc0VuwPeDl0gzIc21D5f6/cpyT+nTfXPoGj0njr28c8xfxui
sdeftTOyBdui/bfgF3koLau1juWfzR4GMLr6+xN+m1SmJ/96QRP6SJls49/x7R6r
3/8kw6wePMdgLDR5CifX209Jy/mBnv44PQB5V/aaPGdHaGN3X5Br9zUpCTDgLNHF
AFGfQn6nvNh37HA2QmkVFta3RjGUCtp7m7S6EtV4VHyQMvUoHN4L1E/k8ee39WBl
zif2lAvSj8IIIgyqj++hNe92Owe7bJ6mUROxA0p0nj3mPPNbd4tmhrUln86afQY0
Fv2SIdL2rCdSnTL9LgifYE3iYqg97m9BK3lXwJcqdc9aZPFS92MK057SCsLBS4Rh
/MOA7ZJEwZDee7H0KH8gTQ1+TW1IO/o8MvqUx+h+r9lBYTFwoP1Sl07y6HKx6urr
AK5hRVwKOd+SnpcHq9/Ffy2VHIdtJclXdEHvijP3V5z2L20k3p8teQyM1meWWAT0
nVXSOY2HXLBmCFyq0D/B0pDjtrdgAouSOvVZiLihafW7Ua8SLjo0a/96I3fW79VF
KQ5aiIZLVN8D7UkuJABfTA9DVBj2vHcxdpzCEohFRwo8m2E1JuW9wSq9VJfKT0bu
xeSroULfkUaDzyCtRvgBzclMN8+C+Bvfsy43CrcX54+xssdQ0PxmbRShSG3jAxDv
X0QRb6Q92XuncplPEvOLZK3HGJLouHmeuYgzrCitMpOHDAiNO1/mFkq8KL1z0f91
dG/1BWfIegEd7lydXPipugWu36Hb4WAWygYhAHH2ukdao4ARZXlcCbpsrKdAF9ex
DJuASLkhR6HJ8PyD+66TZvh/GflY9cOjdIhkme9zXqOAHGMGYCxZGX0tgUHHZTca
bwKYx4D9sJ+dT2kxI4o4WWZWseqMS1LfRRELkGq8PNm1QvGADCSoedl/PZ6ZaIQ+
xUnkdxU/+W69UcLfciTYBl/RvXWuUBpxe4YOTND3UWDRmx6J9qwNwCYOJhfnVp5R
N39OaOLrG8luq8uycrmmxqk7Nbpdv1Wl9JqtNZ5iEgwOxzGgaG3x6XCmQRykZZft
vHkOFjpeafrq04qodj1UrMIm5gzSzgM5LiOEDWc9tJFhnpVCuWMnNXsf3OK3NsAj
sZgzOl2M8v9LBKSctl0ktNcRsa4RoboLMBhQeadl0/vHfabeMeO6077aCps9lQz8
5XPbydG/81ura2BOmyCsnWYjynApXtI153cV1x5AxyHsa7XGU/WrxcHaovACTajc
OYb6RvFYJs/4QqhcK3GDF6cAZ/iRQnb/NsrI9KzAuCfDmW3VG2MSQgoNAt4m12t/
89TTxJvLr0bbcLERHQN37r4505haAWsa9ui09l45chmgax1yhKtqyAxOwZPErAq7
2lUKRJ1rHgtNhp2F8lzkR+O7C68GRirG9jZ0HaUXRf/2+NJpy5RFVUxx7hqDy+H7
IQki2UhPM3U9ScWRTm+3KdlCGAcuBFLBLrZ+xPRNFUyAbvq4JEU/kJc5/MNUE4yk
+BDxbJrYajmExeXfgfTTO+2LrG5/3pi24JfZHiL66Fkg6/RxUFfJx0KqST91l8kN
xWpcl0Ez8GOTLdLlEDU63O0kASMhSZRGTYxAiSN2q3VQ5E5s64mo92RTCKoImTWI
fBOsDSrvKNITGn0fDxCDOzf4UDTDjsAYQIwR1ccKM474uJSWI1B673NCa3/7muOr
Mzfdb3l1nqwo79gdgWUQJhfM0Q1DHOW6KL6kwCoQ5zYrc7Ekm69VApaT29gzOkTC
o/ec6IYWiz4xqp8GOYLDN9OcwZATa/7h2kLD0+RlC+iBzA1g1SN4cr0lIR16jwdt
okCatsrRMaDLbwtDJKANJV3QJO5SCfQLssGrzyI1A0ryzqeOMOU5qGXRD/ti1o/f
EksxaXtjcPk9MQz2Excn2NB/6qJ84/SQnFT20BGW7zXbMtY0hOXKIcUp4lwqXspd
5mVJVBGaa3GG0Bq2oBiszRyb59dFH4gU/Nikhdu9gSKvB42auzNWhr6UxBKrXx/U
8fIX7teHs/P7ctULKrIljwYYb1zkZPhek4or3X86J3mr6hM4UwFBGX8uw7+NP6pk
KX5Kmd4+nFZ7NHd3m3f42Dm4rE4qXtjOSf14uDj7NUVwrbmSU6PQezd6KyIGY5cl
OHMxglRW0Kfi3lXrxDIwdZ1d6i9G6yWs45kKDCJp3/6fjRqquvjcALlVy6g1xo+c
CnrnWFlxnWPLbMfWONrSZXwOf1e9A0TBpbwTW1mYpn2suQ7mDPLthBy9OYwuA0gQ
WjUqxTLWGlFKdIExX40VXEcVRgvq7tB6Pnt1Hk0rJa1y8yDoRp02ve6W/uur8y3B
H2E61X/bleTn8GTwxcJ+sOvvXLrkQdFsR1oj9quO4lBHgm/h4/DMK6lUXhU42wkO
VRHeJu5ZNW49BAXeAoq1NHDxWPF9mVzUfJ08aJbJ0FdhKuBoZpjEUprOqKZvAyXt
PwrpRh/E4HYrqWSbzioivCiVxk/PtHqHvKqlvneG8OREAxI06mrLPT9eK6uLNcbP
5bKeEf10sUVQcN1c/hftmhaoqzkpgndlikr1P9Ie6nAwpud3/WvUg+JaT2ecTecN
9qByQt7SibTwA47y01lJW2NbLMbJAKPya2R5ZFwtTT+NXLTzFKydJZ9Pb+HOV5S+
oZFl9S3CmgmRZHQGMr1cL3jJU7b/7IdCEnhc41UcWlaYoI8aF/vX8tVIuyO+J7Dg
rCOLyIAHG0hAWK0PkYdQltDcO9lmuyecx7X/hM4JKo4hb5aCj+F5NTAtZhSHQaRC
geFRurG212+7f3oetLpalJo/1FAgU8bZHf6ZLWILs1Zgctg60vqAIlYb/kW+gyYu
8UNVRnKDB2+TfGmzPZBaihDo5/gvzAxmYoUXc5VNBrJcbJUS+Bq2lnUugBPrUZrd
ozX+gChtDkKRg5j5fFAkcx6j47vqh4XVJc6JdwtmB/0WJsCfObaTX+5xsY2SAJkR
/Ni7Xum9reuV5WF+LnaVxtEWlS5iE18qI2wsqzIqWcY77stZbUM8AaUhH594lJI9
Dhi4gdniJGGiG/qpo4jzxxVZj68WxIBpOe40Fh9k6aPtby1br8cOxcDhdJiWGfi6
+nOyprdGS7fg/bV3g4+XhJpBkZgsrxpqiT52qiqsnBOpWgVbrG0znF6biJ4Shnxb
DAeW+lECmPd5sAoNlBZYk0JyPXDe4+Q9s6ASFbI4mazZM4eaSmuc0BRHZXhghGPm
OnqmjFvx0CH2nUDPvsKziHxu0BlJZyLZKdkOasx4cbD3RfDQZ0o3KYpdIEamJwpM
sEarvVUKECLkXkvfO6MYon8c7TPstsQh4n6B5+333aI3jEq9X+yIwBvhPuDcxwAN
lefwu9LEanm43EJvNXY8tWfNSyOWIH3K3PQ22ftQIhg+bNqc9FSWwxdRC+OonyCR
yCmCmC3JZysLlBw/YqJNAon+X2pZWkD4aERD9nuhusoGEBugaui7avgfkunTv96a
hnohuWJZY5jkNz/evpoCzj1W3SynPs2PLpSxg//qkuTIikVzk2AcqyurGcc8vSNu
qUtLflMautYz23KQ4e73mZgRmVJHavMopJdVWNB4TjksVyq7kkfk/Bd97zW5ow5F
gtWyuRrzCfqh05bHIfYox/aOUsgfoUEF9A619EQ8Xk71O+xb5GzL2RqILC1Nx4q7
I5LvLr6tk6YEZV7oXPSaYD5aU55jcoRfNmLGDkmG6E5Ume/Gscs1wUOI/iYTnz23
KuhNrHp8g0hrXufAXTltxRuYCKvyK/I9ClyAEsVCaIRl9JcpMax6YC/0z4ekYCsz
yQ+Mvztvv+4i/58+1R9kXaPk3PjjMi8owoB7xmEANb8E9+g9gpNI/20/2ujiisv1
4dePQyeMXNNaJAx7yVO+gLql6/6I6ritB+/EggZ6ItS8T5XWCB4XrtUZ+Sb7+r70
W3ZLSXvh4ZC2h2qx7kda/uvS6jq5zCirgX1Z7VksAFyoJTYg95B6+YfhUe956Zz3
cXvpPYX23nSqMIUF2+faelSDZ2F+jdOzYGWOa+oEwqijELsBNJMlr8vkVracJK9T
94Y8xMbAxQPlQX3R1w+YQE26bXWvgTG0ODRJbssCnZMIUGd7K8uACn5JRPXsxPlb
U2gg9noa76DQBeK6S0P0MEqe0IVYoKq4BWQYUeSiJoN7lVhYhTbMbKcARZq0Z2l6
8dFuztwn47/leY3S5HA9UVcF4vVXslhZZPM6ZnjUUqDUwHjh7ce32oDa5wAxPc1X
MwDG+NjpErJRa+s8bFz7mJH9fCSW6gJjj5hBHdoVci7ASuQjuI99hJdA1iXpsmoC
XHUqxYuawnCJwKMCEQz/JBFv6BgmttMVWgHcEwgf64Vpk3RjbtEh1IA70BqUp28P
k/JaSLn+YrOqjKCVaEEogrI/xFUo93HVMgpVLNJa00dOtvYWmgzKJKwOI6sCUPs6
31i1aGkLcSDkmi/iWNiUa70CF19lKt8bjVDcp4gbNME52eCmyBLF4JNc2LVlH3xT
ozG4zJ+V3O7e4rcLDCUg46MbU3NHjdUw6i92SqDnXacZTI4Y9y3leEf1z6VZczKQ
FLzkoNANjp7QpXVRKok1K4gbDrYkbgW+madBEyh8oZgJmDr3XmIo1qtybCKchUCg
qZuvz73Cb1c332Q6ahrIAIH3kfAlZdKFb45wuzYd1CH4NM9IqInJbJ44fHY2qRwc
Uz8JngdCcFoK5fnAOROOTI6i9EGhrxhDBzH5xVOH/LSh2/Q9qSAk6UNMN1e7Sp3x
/r2ER+aHdvftCxB9/J3MrIOIiuofc/V4dQRs0S4mrj0kg1oH01hmZsLOGh2gI7xS
ABgM0+wOB3CO3ro/x8yaK/HKzP0D8C788ZUY65RWUlZfJ5JL4uuV9NppTJsmwxlb
MJzqwd47ukdvk4v1j6JVIqnNULF1RTScAGZDvh/swxX0qFaSUP0j+8J09+BbT5p4
H7sgYqMUdTQGXps3QmrkpZBWsRxIZPEiom/ldfGWPG8GfL8NmXz96IZ1e7mFi3jq
o+xgIbx2LAeAu/nkUWFFeKlELXbTnQM22AVSo/uTFTQGVuJHQqgX43q06E3dEb0B
8G/5Tt/vvACvDxMNwt4xxLYF3vPxWuzTpbkBPYtShzV9h4amNcMAAu82zWuDCxky
jMKD/wQ2zw5DLquorS5xJpXt1D9J08UILVIHxur0LK90tML7TiREfW3iXF+XSblG
2JCe0NkPZFjvr+BCYIsYETMUnpz1ZA6Dv5NPVi06lIi/6R+5OYshI/JZ8YkHxdNC
9aqbtKDJ6OjwhHD9tDlhWIUIqza05HbgatxbhZw5hB3QRKoAoz3deWnGgYtc4gEM
td69aamg17EY/ip80ceXmwkCEXoRvtPcSt4ae34Xu0da7q3yHtRx0K1EVdnIrKVB
Td5JVSphko/N1mKLmn4g/2q+63NmT9cdI/78Y8uN40Ogwr+TcBmh2RNCrtmODp05
/xtotzDQbuyrJVsXiOSqFuYmQ1fD8sLaK/XkPkOKDobUcl2XB5F1xTht2KMnXeoG
dhtjds3Ihml2lq3zLzuk6rSxASoGa3uMl9a7idlhnMPffN6SITA5FW5Bq9jWeh5f
ye+zlJJ9lyXWENOwMHBiK6Dtqiz3A0awxqP80mW+sQdTlu8hqgXmRl5PNPP9hiI8
9CHHPnPObWhAh16084l0wkya5QlqAe+amnOTWS7qDA0StxZPmu3icap59Xyfatv/
rNJEnGW/8d9lP62xTxvvsZEIoN/dAi7xMDmPnR73Ed7Bt0RixU+D2tyDA9a5vaFY
CnMtDwUSAQxU4PpCI2avOUFbmLuLXsmtvLxjuueMYw7oE4F/KILHCBBhmgHkfWpl
hDAdXu9TBo+ks4r1qetDY++fOcG/m3Y/oOkjghAbhEJhju/kXra/USUn5ea2uvo0
5qSs0uiA1In7GsMX0ABKsCX/XLxO0zD/sNYumAZH29Eocte1XwZM99YHPo4NEHyB
ZmOlwsT3IAHfpzQex1KGjts0oOos2fVWx3zc7Gt7lKjvMrZBy2SluwdI7V3KFg9E
l6rL+adjNc/xSQPbfLDUGPRVhs0IJBJVhXPg2NE+bYxJVUXFZuJfn308BCZAN+lS
1xJ/xPfv9r6VgLpqY6gNKqc8BFT2BlRVgUQ49bdCJnTN4YPSUwxgIRncCp1MsOJA
apUAujA0l7kT2DyQnOhutBqSR8w9diLBUZOKGfqyvhuznScaRi2jje88SIh87LTt
YvtDp2FduMMquqhooBOPYw0Trj4I0lU3/+bZGOrZ38FsSbs/U7BI6omVG9rLIl3q
o9BXSFbvTCdrw1seiaQEJylimHkFMYixTaMc6WfCIrStYfGf7TXzbo/m+7UrTwY1
ygk0iY53wDdzS8hGOCNLHOW2r1nrCSLvnPn6PQtlQ+bIkA/qx14UgTXu0+n6//vU
S8Zfc2el85vT5NZlb06+A4BQUhPkd7D1udrqu03i4/+duGUjjHHISov6txaYFJcY
ZQwhhDIDdpn0UlKKAnrYVAGl4PUk0kkxxCLSzhabg7J4pDCxbPseCWSsnc9uZTGo
Rnwwy2PWL8Zcry4CdgH31duD2T/O2fTEUdwj6gh0K3WU21TeMfFDBk7Jxbuja6EK
2AZfge0VF9WvKLCTWyuxJbZgWM7LV8NjOu3GSzEyTqSxl29o1IwMhRHJB6HAgkMo
g+dYRLSp6rHbGc8L+LkBbpeZszNGQ04lfjIMIxk5gMTr8kh0x7/31/9Eb9h6A/q6
Y5qY/BA/EmGMnW64VBOHxe/FlEj2LSpSQdNu0SLkPQdAcPauHO6AJ+atGcqUhwEK
0X1SkXQWA5k7j1xFW/r22/RCwrlY3X7zl8AfUEJuDPxGIH3tC3mebjJYEWxH6MdY
X+ABGbF9xg4st+QGfvnr2B9uDadYpAXrH2Nd1SDoAxvyArGAK9T/KHAyNJN9wWS7
JGYbtVvIz4mnts+VMwB66718GtfugyuLKGS2tnSkSLCPAbQvHa3VnUXFIQ/AtqAY
/qo/BS3YdKiddR2FHfqrnRosJBbdV+N5FXen60BgukLobIp8WaSMQwwnwSAN4Pnf
Vg6EtHDyjz2vQDr8KweI9gQQajKOH1q1uP+Dfv5pQL9+S0ieBUJeG+CLrPMHZ9MB
vYs6duxcHas5bDPp6x97fw7mriyfe7jAoeB8HXQFsWPraNVGhwGPJJHmhL6Sjo9A
woNnSU0NVTxOyl45iMJRMLkMWDgnOQ7k0mfEFvcXut/pAHinzen8ySoEh6ZlynkB
teK7aqSrDTgLchDv6aBNRaJuxvsZYyboexkGdvWx0M1RvZ473Ylrrh/Nt2OgM8kh
8RC6F5TprGVyCd+2EsFVVqVxm/dtC1OZa7yIQSjNZTHSHwUBKTo0UK4xL/dfFX1+
ly7zGbnhjRhQYDBRZPGsEHgPbd+jhp9+HsE9kfr6/09E1ipQEb2Alfd1E+firBZ5
4frRRl1j8TXZMLuwSdllyUca6q1ZwQgWbkYCcTq5YgP1zsbmKJakQxlOdAvBDYCB
Xk2AheKmHLw6UpvaazXFCiNt0KdCzHslYfmIJYkFCnx99D/Pq0fwovISE/mt1LwG
g5yXMkIHpJDUOd1HE45aCmf/u6f4zMkyI6z+VeFjUj4+i+M6cZryGXVxhnhKp2Wa
HW+6DdnFxzxovh0NOhGUZ9VlEX0WF7X4t3pI8S+tPB7OHw+FS152Zsgwhtcd+6Zq
1Ax4ZO73e5EUo3JyRgb46oT9FMDxzPuaLazymagBXXYmMHJ/GI9O6NNi7aeDjlmQ
IDTaU9jkDPLQ0ORE4L2QubV1V4xoKPO4CtAyiLToNQf1jmwm7jUO1r+WEPTfs2UW
WI7VeWTJ4SIJTXRD1XX1esXOTTf5c6g8wO/mXgEYQOfgM6+hVuUqJLUrEOQELmvi
OZgIEUS44TOoqW9SCBba7g0cFliPm/4XQCj6I4Fkr+3+ilSglP9pcz0zrh7AHz1S
QaEuwMmitl5tilYKEAjxgDor7LJIRYIIxUk9omc5hvdDncJhZSq+41TfHgURG8fj
zsyzcAAP9coQqQICBEAqm6Vlua/HIibJEa34PExF+Rpo1qaWgvFiduA5BZ4eCcpd
MhoKBuj4mB0ac0sooPLzfettP/TG0nR1uINB+dFCYzVKv6FoKYKcsQ0zF71y5vkD
2Z7dD2Ru+cAU+ZGWagwdmgpo7ImidV1F2sr5GM2bwgGgTZdMecTDEzm8afi+DoNw
yAtlu/UhB5ESMzcIVo+DK0TQBiiCwoeaxBkSeXQcaEyuBIcF3OO2gv/vxIBVOylH
sKeIqM8lCoxGC/4WSGZjlAOKae1p86PCK7q8MJt+VNjXfwu0lOa1dYZY1EsGF34f
lDx8f4jyZcP8aSGsf3v4+j0B2IeEXF/ndkibtkJips2FOXA/OuhZjNXOZWDm7+UO
TigzUV8v87GUGaUu6hZC/FzVDyr4bBxGqDkSom8INpFMAoxxd6fC5t4ckDr8pvXl
sVI7NDJVElInYbAwledu25PNCw3mcmCiueQCfziq/ZNdpJTfzOcSxdr2c+aKFzBg
o2hDvwFqkLGw2DZ7tQjoQrv4eJKIM5edGz4qLrtA2kDgiCtISNj2KnnubjgVmUvr
6YNlzABSMKIrqbyIonv1bqyfExUUwMx/Ct4N02HwcDMYTDZFCYEbi9dmkGalQa4D
Umrc251dPyWYTBNPoOU8POtpUfHhRsTyrmovV4gPWcDPWcuPZSlU4qRlRbLWIJ/E
ZO0VUIYAxQjodKxpNWwwydcjOkik6D0scwY53pkZ0ICmThhjTG18o0p01U517sMX
++9MxoODr85istsAhbRcf87uXfAH85njSbWGgdgI6peVsZH4XpKUHhq69aRwv2lq
J71QWUFSsyd15HB6SmiUmmaZPNzzz7iV1N5a0syqGLmwNzkAxnSYLMGEPb92JnHP
wRAE7me4bcFdrbMLOtw/YLAXzyRycXSfEp6Vd8xe0u+8yNEjIUJCxQIyaCHxgtpy
lcheYwYZ1v9Wuxz7q59RK3HMA4mA1cUugrK1ndBeVtQrwTaW8rFbjaeANIL8RsUB
AYua3gx5nk6Y33pXXMXj7MiJeqJfXMmGN7sBaZN7rONbqkYc7AcgivPE/zi+cq9Z
4Wj9W9bYJPOb4XouekZ2r+cmb1w+W1lko/zUzOyPOisAJ5YK8Xc6Mh8MV/f2EgGP
CFmP66CIYNm3VFtdE/wE2hvyQe93S37GljESBKf67zUB4cpH5blINmKM5pZPxCWW
dPUhM+8+YREagvUD/saMZ5VplX0HXMe6zpe5zU7fCMbTZjyqsfR+Uv1exW2J8R5e
lJY7qkGHo61pa/gH1/ThNxJFNKmD1fI5Ggwp5zPZYEWxd8VjLZg4oxzi3O/JcGlu
CLCdtgW7fFjRshdxylce8KogBqqhDMr2iEvqXK9xIcO/ltaVlkV3n5F7bP/OR6W6
WOzXmFbE0fNjU1wSaT2lyNLC9VuRySjtexZQXtiJeF13fP+CdPRmb17O5H4ZmXf+
MDP4/+9OM+XN9+dQbDrJ5SAqvBquvAB0uYjlz2PHze/rxSt+c+j0mHsKvbm8o1bF
vYET3EH34Tjz0HdXJ/F8lopp1GAcGqFgQ2jINLAZKlYWmoelkB13Qq+4MkkYGZCq
8/zy3pTwm+Rnx3WSchyAQbb9VWNyleX40NaB0bVtPhgCDSgigFVugMeYBrkFyQLp
fA7PXWQzqBmqXrEJ6kdd4VXrSJBltdl2kvdkkpjJVf9rTVdQ1m/NSzpkg04qogLM
J+WTBNaBCdFQ0RTGn/m8js3gfD6mt8GKZR1ISwX+9o9cVp5WC64u6yPuoIsAe8mC
sgrhcii7AqEOxqaw8ZMctjPWLX9a7btaR2aJoJEMY88yzcjOd6SsuKrHKqxCVSpY
hGwD87s1P6L9AGVCX+y6stRiZZ0lbrII+0FvkoaV3nnl0Xm/+8+1gqiAG8f/s1XA
FgegGsE0YXfMVvofS3sffHvQBbfhFNmEDmqb2UwHM+QmlbmMz4Vz2+esXXsRwuXs
65ZMEMnho3gJl3+O2kIpU5RWMMQ5Y0A/7z9gG/M0RBqZWvsbC/MgMpxAY+MG9Pm/
H9DqvfVEpoKZiTvp2MBOtKlLLVL/y/uM+ed5U8tvsmkTV2t2WsXWHU84x+TyntJt
RqILqX31SWvjBLQn4VUCx0QM1x+ujVwJ4EVSeSRcobrGJfRi53Cz5HQvDht5sEhH
+DquUm3VQCebNmCAHsWOAynP8ZJaW0Ki8xVrpQymmjqPYNiHsSqKrwWtkTOsLuGS
aZiOFwtdoz5sYAZG0fFX+dKRVQqKVih5espLdFRklOS9Fxjzs1e3ir4w+ESNzWqf
mO21LcBBdGSvknwO0lELoiM26MCFINKbpnDduuMiMw85gMvGxmZaTOs8aFoJGSQd
+LqWtTDy6kTHuTVlR2U174Ll5M5yP82QQWmV0SKWUSjCMDtPooVhcrpEW7zRsEb1
hcXG3Cuav3T8tdjhRp39s/Kzm6iBQmle5RJbdq6O83momOZtmJEYUzCFOOeVlTsD
FyxIFsti19EALRTwfB+I7RS0SFG3hkMgEL0mBq01+H1t1brCYVDe9QHSd9WFzgZ9
cB1AstMujLJ0fxz1RtR+fumMrkhM3N4tS2NchaOcngAg/CuLWmCqh0iK/uJmsjYK
l51x2R8Oe5bYBr6YqDMoHoaFfIcLW4Zjs9j/0ij/vByfkU7i6XAnThur+yXBx8Jw
+FY5X2s8i1jP5nn6SES8pY0Gj4SSCtiDPtbbHmv6AM3S0KQVZdBhl4k6L82JnABV
UdF2QhXeSw4WrWI6z2c1ZVx0JPHsUY2zy5oXUEl1ZfiAQYHsDb3QtIiFwXY7/Bgo
U+o6rgoO1Bsrb1EytU1+bxOan0GwM+BSs22ClTYuwWMsRnteNT1ipS9f+oQzos3w
XIo7Yt7f1/bTBOM4IWGmOPKodELSQodkthfpn/sjkOgfjJuXuwQHHHeYzfsQgf5N
HI5f99nskvqVtuOoogmbK7SRI8nS85d14bgYsmlHjg8otR3aulOFdmP5HyCPK98b
TDiP0VTqGoCbD8nrzjiSGWgcGvQGzYcqVCXww1PD12AD9rsrfi5CuMNwD9+oqoRd
uCEiaYZVx47vH6jsn44S22Z7SmZWetwdnEAIEE7IrdteExO2LR/Zjn/iRxNm9tuw
ve1Lrb0yKorkox77o1PrkrwOD98qPZfe83dIwoMK87zQxhVRRANdMBzi+u4/OKYB
69dx/NccAcaFlh0L4dxsz0moPDFRGdlt0f02OZYOoJ5aH1zLxShKOSvNOU90qnR4
EBfcwxOa8Lbucx0uGogMdqkfP6Gsq4wduslG46guKe8m5HeUjhOATWg+R47+b+ln
UDD2SUfShbaI1vP/2Si34EVPiQeZNzVLqnOv/emqtp9sOtKa5JJpwfhvuqIuWaf+
VAeQHZUG4mCJlF8mGoOppXhSSd6AffAEd0h7XLczzJzzcJ7lgeaE5334z4jYfP7Y
9GAvOIPYF8YNXff6PmWHuOxAS4/tUOg8tv5oNgFzS0CUAiVyAGYmwLWZAlc1EiUt
M0CvT697bs1EBwK9wsfbRrDFCIY4AI55jlbkEGeHanbMi88SvMNlbss3WpkwoWpf
PZVkBt4DPyvlZ1F8V0pTOhnFhBSooe2rgN2bgwcaJcXmJPcgloBVb7ZKkg5yD8Pm
1ob65RCOyzJFGoZNfExcoZ9CDp2H8r4BrpXVtwWu8Fy23M9DZTgHZboA5x5J4AMd
uzNCkG26MgxNbdqNaWwwBX05JuRm+iXZBODMGit93Y4iJEl11WAcVSje8Cn17oQp
GZxXJRPevDtmVPe+tUv5rTuj7GV64OZp3lo/LOVSAr5/5qH8dSrncGst0xlj5swP
ahAwwa87Y8ozpq9QadIOG+ZRXUiJU6s+/B8zMAvMk2dzpXCYSt3ewSO1i+ETnWle
yjXGy4P3roQ/djceMeWPL0Kxz6I0QTXLeKTw5HJ/OIv0xl/mmNlp9a7xaJDlxtqh
/xtgOxPzTR9LMQXKoqQDoX3tlw2S1BojKFhyGLiDcdapI1PwVvheroHSa7OW6bZq
pWCcsFYQicN6r+Xd0kV/kfvQmP3CRE/tJNh9nBuvBj7JerbW36QZK52rdqayOVKn
wj3NVhwJNjKKoIE+DnVWJp1uS2+3bgFwechBl0CqF9TWTPk5LdDOAWhq3t91I4Li
bcYscjDj+pDI2RJ7u7gdoKU4EdXWp+/pS1mAl980OsWg0TaHl/WdwakJ5o6MHggY
42Bfllek7N6XyxxSlkoXz/+si/86jdhb6Jxqq9ZCNmIuRDtHo6xhIdKiFK/kxqSP
cb+nS3VVy5FnlelN6AkKzfj6yaET4AjjQYVD9BFbobHBG/kIy3/dZWkoYWJQe/le
JssQ1r4B61q6NC8vss9XVkZmVPmD1QCx8EDzzawWSyii9wVomp4Dy6ia459CD4oR
7tlUzdwy18Z5tkKBzKK4fUKmpKDohx5JB0oci7R76T2drXfUc6vQPq3BadcIK61s
jH/HB5JOCQ5Q+S7x6BOOc1n0qBeFKph4bYhfXb82dQmvIRKVbyB3vG/j3FLZFHNp
etQz459w3sWCecalcQL1Hq6uL+hzQQc+cn9llUkhagSff7p6A2D4LWmxwUpoHxnY
Bo5P+VN3yLE020FdljEBGS+IKZ2wn6xiM8h8ARhnEQ7MHlZC+KhdhEIxKlqv5YQa
f1R1Ve/0ucZBuxVsWYGploiU2WmJ3bt9hIHFGgB6IwSrkMpVJh9K/B4NDgP+lAHC
WpfluaMSTvZKyIXUSD0h9COUDkwshEC6J+Tcq4ZZxvHTetGzvLOhCu4lHMCtyLX7
kwPJ1DgbktXdT9SbSt/da+25alIYmmtkGfRHsbCuWQy2g+EiXN3RFf78tMreDx1G
pdCv3pw0JeFk0xEoQtTpKzCT3oEk1s37tYgifDwa7fXqtvcleXAxk4OS0zkFzT2r
DveXrhiXJWBTDMpzU7ntVzlKdOKltffZv/rvv8mK9dRQj769bFqElzHIu0TLeFw3
9byIAcnid+JkvSQqIN8+kGKfhydBmMRqQp1Q29Fc1Ou2N96ODjUYpJHk3P+Pb4QZ
oWN4sYMn1JBPwQWK9JZ6SqI0VpMuHn88cSbcvtuMu4rsyVHxRzInmjqt9KqtXQdr
yb6qWmKedBkpjbaJRc9UFxmlG7quBf4Zw7KXSU+YNlApPt/lLbIiLnBmyy9s1XpH
2TbBhvJS2XZQe1F1lrqWIpZvtJMx+yk/ViW94vo2EAbVt/BnBb52AjHQ8Ctl9uN6
M8NkZy1tmSt2mbi4ltx5cztk/g7sDDFRarQeAsgDM4U/sbOtPW2pT71SCxjfWhSG
sEt7whPBfqXrJKNRVFR5kaGXzVTrBOg9te3lmsLUxncTOwNvsyRwKQcY8tX3QHvo
ikzrh2Vo81toUr2xmZlI52pPEXi2xGDpG8dSpgYBqb1aDJg+/gKA/Lj0XiB5REXj
hLvKeSS+j/TDCKhUkdvmCuINswGQ8avi8IvfIFNPip+GLLIdk2l+bKjLZDE566I3
fh8fXAPnIqHA78thpUQqH1KPliH5Em0giiwQfqCO3fgTNVb0hQ93fThDcZ0p8rj6
osaoDogNvBfCneZDRjk35yhOS0iPE8YYYQDCzLce5zwQsZ+oeq0Yk2RgA3bHpAoR
I556zpTHg81RuRKIYbckqJUse7oODauJeRV9eLhOJbmsbVM849C4w956S6WZ+PTH
DoYWn1Y5Zzw6CxrzdmgjVpsDSLRQweyW5tl9fNQIkdEbvWXAaoGhso5WhHJJDXBy
+2xf+SAUjC0hWqop4zX7YHDp/NfQCBrXOoaofjaZP2079AKUnU8PjrnoNxnuSzeZ
AmZHGa+PVBLY5skc9+89p5PQYPputy3gV0XPwnabyZ8uksS4vWhUgE5cnXNAg/oE
lIjIFikjB/37rfV0tqvuCRfF4luQPcpcL+//z9FBS8AHuM+YHABuweHbyz+Sjxs7
gaPfG18G9ylniinvgqYhLoCC0iM0Q770vnL9FVfKrE0dhMu9kNdxysIBkS6PHean
7Psin6BkrkT707xN1yi6coZsCajAA27EIEZsNjzIJvVIbvC4+aiUuA4iygwNR2vs
CRAqtAxcNm3bhUaSjYfSPR1F1UrjkZToc5Fc1ggiZBg+JWvdP2odG6IImyGT0zXW
qCmWE7d8i7MyCKpZJGG4qa9XSoNnW/KcER5c2jslGqLsijaiBPVZahcc68QA16x1
y9ny1JqsJnD5E6qH6NQ5YwMUHjpW3OraLcdpnH/VrlsLQsB+7/+mVMPFsKlluM9S
a0hrIqdyX8dGx6VY4+c4nwxhOj7pbork4ITyZY+FafM7URv40LuO0OtetxOa4byl
sSn3lrSqPAJp9f4vMbadcnVprkRLA/egABrhjxo876OrK21HO0h1tMnbdSnMYu+t
3vvEXiofUW9RMkOgoG9+XeXbglh88kyhRjlr0RCmkuYudt+6QcL1Zk88x2Pr3dC4
Vfjqk/FQ2GDEOsVzNs1fNPbX01TeCPT3wMvtAB9fW2QPBdRj5PnUUbPfgP29JaBf
wWe3LEw/sdoM3u4h0vejoGvK/v2gVLw1ezC+AI0I8WqmuC8JCKG6qqzM4IOp19rE
t1NIs43KAq8065CdkCzcomhHJfysuCTwmYxURKvwMiEYZ1bCq81wXcr609wHO4Mt
T9lGzm5PmKOpLnVlLEOkMUfAdhVypU4pluoNnlwSzz4t4aSETICC+q5qOTuPXQuR
1hLZCJJ8R1fEeQDegO0+hQHCdL0WsNYEHPyFS//E7PA3Njg8gSjP2oGdOs578AQG
IwbCqyElQLAaPtXdMNw63++TCVpuwslNdmOn4IoIimCZAUwh7ejIN5CDtPmCZIB1
jNxS1Z+MBnYPBS2BvyQIZnZQkrEvz7/qHkwDjm53nMQ0hUjiMbV/nxwpm1hOEuvd
vF/DdLycmNDENVjfOE8/jpwP/dKDQ47HhFqDRzHOmJpS3vn1n7zQ3uUMCttftHgF
UdI6LZ3lYFbn/1rH2P7wLaZtCvK9OHiEvCRMB/VrVuHRRQqnoFwjslHx7mjUhGwH
cK6Rdp2/5DNCTupbpmS09z/FDn2x/UtlwIbhOghB5/8fLpAWKcm6f16Q6aVYRvey
uNvVF9woc3WsV3sa4l66RofrnecPw33bCFFrL7H7xZWRIV5SyDr4Aw2ZieFgZ+vG
dfP4dFbvY0YuBlhu6yBmEHwAs4Vj/DBjloQFzaaWCyly8JC8ZCWU3DE0Tf7Htmiq
LhnzEE9XN+5W9lqEKiKvSQtqKKxo55n4bb+uAvRHSUVw/ql1abwz9euRuqBDVSBn
QO7AzyosHEo5yL0bnpWOXrlgRjepBkE/8JIj7Z290L1Zt5KM6vFJhIJuUh5e5Lje
HCqJMjGPA/PQ8HQlDTRU5MHXqc7xoS4XZn1RyKfbKb8gIyPiGujCaIakQ7paxXoi
ZvfpCHInvT3WzivT0JVTkkS/wdCx10ASQijYB+DhF7HC1v45MWKntjQ5WpGUL3dJ
gYgXCO2SF1nVIP8Kq0MjFJPXK+x0bvK0NLt2cOA9Kh4FpzLFz3bjeqhIp6eiCKSH
nuwSUI4eCjdsbCNz9gUtvhRTyEi4XVMULcX9uU5W0OUeR3RejvS5WTcuekFf5Uer
EX4ryeLvRIC2H6x+EBXS+0MQuNvEz2kHVSuoazxoKs20BrIMkdwsEO+ga87r1E8F
wIGo2/jNz4u5C3eAqbsRo6Cv5yHy4hOorJgcQcSSzu2OT5bjyrU2+KvqFWk82NFG
5cNDIR1Cmqjk90z8w0ihhw7725fLVmVaRrVKP1Seie2xtdmIftfHJvVBDFr8QbCW
OuW6Qp1yVEW2zcmlA/zu05YDQIRFWZOZwEovH6yKEBbP8BF08Bt2fuWIpC+/8nS8
eouwnhXCNVlGOd643P7w5YQmHG3/PwBIaFo/ysHBQW2cXfnmrGPhMd2TsIzjAp6c
tkp3uQDi79XzjsbUx2Y8c6RUdxWeOsUppVN7x6LoCy9H/4OCTO0zaguOI0ej+mSD
2M3TI4P4M9HLEChvEfEhqB9KNup2ePHRn+UPrO7HG5x8BM+NjE3FsyBttIZiulxZ
T1+TZd+hroPjCr+IdcT9Y/SgnWXS0U2dEqOfI8slyoC4GhzhG6wZ5mxN2BQNa7bd
USNq2H3/mGqlr79BDbcyfSyWDIh9KSKIFj7S1jT1tGl5+z+bhVSRe5PFIQpGoGw6
2PHUabzvsh8RR2SswnR8BslyK2HWqSOzANn8bvGXUgXbfNDx0wdcHU4QntEYBMIy
fUMY9gBUC8MBP+JAFE6mr3AMyrhYr9P9qUu9yyKrP8sW11E70b79z4YXNS4c9Uhv
BadFbhrcfB+/h8B9RsZRUEiiWbp66Suy4hyeP2OyKPlsybarlRzXsmDB8ytW8IQL
+ak/XYsWrg+1B2t79EW1nDgUMRb3eT6ALULHOjx0zuOO0sSWPmlqu+QD9LmyBAn4
qBk0Mk6zCzrzBh6z0piNOJY91IXrhJy2oP6ALZp5OLiJbPtO6rKrO+d47d12Jfax
ZOf3oLl5iowKoJmSAD+BtEiGsqDFyJs1EPK0+c5+3T7LA8zsV3yyUCCMeXpFCNUf
s49nE6b0VVMN1EQ/TCXsc0PB/H0xw+NfjgHD/E3wMwhWpA+cuVVVkVK/jK3LUp6X
NDgShs4iDbbdqe55l+lvB7h4aaBAmW6jKU+fK3EHo5j8Vj6AN9Km++4gnPZPWoYS
1hIr7SdxHQ0DIvEJyzFqMb+FbUIOkbca6Bj4yX6uIRILD/PpkXYcYcymtFhGJ0ag
plkn90JBuuja6F3g+g5YOPJHNGukWl8eLJu0YPKj8gLOOVj96IOkOKZukPWtcMQK
ZRs7gl4AKxG2glnO7yr3k0iP9eTEaGgG9iy4RQbAlcKoZApcsyp0Jy3mI61XFZ9n
YvpEG1DuggTl6oKHLb0FkAXjzA+3mgWV+eFoEEHcAE+3o/qO6a9UYtR2FlZagQX3
aWa5LKkCdVe+kmPZAFBP3AXCEI2H5eL4w6jJSs3zSpjVB7qEyKP0RvUB/jqu75eB
MWuKFe+L+NjOhR59SFUrZAoT7TVfeWz1fAGnhIVodVnftxz/hXUKGiwUFQCvStad
s1p2h/dR1OdahWdVB20pOmUkx2cxRCe9OuCaDzIu1DqY3e1BiX5uYZFC61rYYW6W
tv5WdrBLi1Igw6syjSC99MxOIeDO7kiQtihO6quAGC+7lGDcUgTggsK1Qf9XqTDg
rD/bCJqNDIjCYSxJxgwidWaAIOa+4hyY7Vzs2TIFaqt/5wbtb+ZoCBPNRppVEJht
jEovNFNJ6wXjfogU50LTq1Tx9/G5+va+PhryApm6y2tR2Ib4T+V680dR9JMxhFjT
AocIqCn9lhY7t/xJs5zZHYtWnL9yOFlnXdvRiMYNOdiZKfVD/CWw4YWBzafKZAts
sM5WR9DVYf9ViH0SnIMxLr4jcNjvZEM1Q69Tl/+gZ/GmiG3rdzLEvCOq7vV4Z8Pt
pNzM4mURHXqjP/UV9RUh6eF00TTILMLRpN9MVtaC/5MMwSAN8ZzS3oQxzvn7QgQx
a2GJA533ozZRreGmgNL7lwktWZGGb8xXv3ag29PLvBRkQj0SbEk6Ga3rDOlfNs8c
2GbsCo3ebEUXuB863TS3VoMol+qhH3kgeLSjPNXnhATXT+XQ+0sgZhg3gpeMLS8I
F6JuLu53Q7YNdTnlXHh6X+YJVnz44QmlMpr0aaLTDYUzsAMEFu1AJ+ORVfuGDz7q
Uln/7Px/EQC1oaqX9wh8afFTrN+XvqCZ5EFAJM7CJiusSwZNERShawxiQtZ7Czdt
NYtMDGJyq50oqZOMiGVSX91jJXOa/ek1aFIa6vHwuDKZ54R+ey8rzBtaX9qxfbxt
LukIrw0aSFHS2q4930UuKtKPHEQA1IpU2C7vO+V4Sk+X0+YklHdYoPUHVsfoj+E8
tFb6wB/k8VqyZNvXW4tj16G5feBsmYqu6E+V8AXJYnWx8MytkbqYAGA4cgYZFlKW
3TgeBEPik+9c7+LiuYuUb3K9uH1aiQzMIrlJuEoKkFrtLVIjK4Dy8m+NqqAPzqz2
ueUgM6q16hQNfXtHsDPHFiS1AiAu9UEWPu8sZkneVIGX/I+katiP5wFJHMI45hDK
9hYymI+RxvxhyzeFyquwr7FzBRSBy/swsHl+5Tk/k1NJkk1gCxZvzabFSjKVlR+O
UCrV1HRO9CDgQW2VVrC8SHoiXYHSr+OClgot2qbZ8IV2Rpi+KHKA5uhkntg0wGzY
3Hk65mEx4MRTXulJcDELSuO/IuJXePDyzB0gbeO5vMyHqPvQId2W5uNnV3PjWVXY
jV0LUDWfSytitFS32o3d29/oze62+q1eLnKDcjE7kWYdG3RMsuJdwMEBb4y6hYTN
Mcp+2sbnUwAhsyJ01lbfjN2rDmIiLZgbMozTgDHjzClBFe+OW7wgNLLLSmXVMm12
SYmkc+tNSXAtThxK3JuMLWp7CtJTdECgGXgiQa84tjhG284EEypVK7QVLJfR2i34
Xm5qqsTIvoYJxlzfE8no9RGM4o2ZzPG1a12W1FUKlS6FkkjyeIDQ0Vsj0X1f82Xw
PBWg8uGOVcSGAhTn9ZQySJyS2+zQaqks9YHcIcmLKHopUG8ylA66alIcwbRQ8YGj
BPwtq5va6fRICiwMAhU3FKodOR99I0wzaM+I7rtDjNSWRt8syfhTK7S91Cbgrng9
gkIwLQizDvuYUjZD6cdkUC9im9XQ1X7Dop9jePTGgOB4p+4UhnJlLNn19q+Qfh0d
m/a4kvDhWt8D5yoiGApT3HlGK0+CJerZofTl2KsUFOjtydTcqA1heKc6OUb9Z5C1
LMkjHmLH9c63OepvdpFZWTZhTh6vHwm6ZZqg2B71RnWzycg3BxLpciuWoIuuEK6G
EFpHRRkc+xFKOOg2pEpwLyw+WFsviuxiFkaDZQnkE0uyxXi7w6ksyPzrBsOeDhMp
v2HOWtO7UGbmWgTnUgQ5hsGVKcqE3W6cKsCNjZQhdkeqlngYEfan4dUwNVHiRf4I
J4cPTJ7q1p0vbtKXdWqwzmQuqCC/bcj8YZ4xuUgI0rfzI8dj6lJdjZh62N0V0Vao
ScfahaCSVf0ZmNhYA9RSUCftODoBZcVypEH8pWmN4JIivkug0fRRrO8Gj4SRhaRy
FmiQC+uOP/ngDeq/pzD0jxSr4JMzefwrFjw2ufrfQusBJLxiXq1h6gjlRrl9WaD0
n7HUGUg+iehRU6er0ah/NzVZGfZ4hBG75QTkI07skCAkoVYa2eOVNmomgOJIZAGe
CO89UUl3Mp0UFb2zTpv/QiKNGMHif7CuHecCrmZ6sGmWUn7RToVVbO2GWdtzmiIb
hWlrbyIglaEAVZ1R/rVXC2LJ18GwigpfAQQK2bSXnvDY3GUHaOZcv0Jw6GEaQQfd
zhSPXXjmCVS6FmiBUS3ftJwjG51zrXiFbeNjFmMXuO8jA3pLU/e5GFi0qVHcwYzl
f4f4Z92dIun0VBzjXA6+0hozSezcmXPfiLN8JqC61iJLuytRnuWG6UZ+dWDd6Zao
oDC5p4ktpNJQCx7HnCwWeWF3R4L7b5D6nOV03NCZn0v1C46l5o35wIYNY27mvEdO
/8inD/APepHzXk5nSIsoFT3fVxrY/VUfniLTaGYbrBoRMHpsc9DuPa11Gv6rGf+k
73ptXb0jpM4az7r6tp2ZyIXUy1xWZixQEbnfYLkBL3Nke0rN2LPa04CxEyo2QWod
x/3rEom0m9S3niHsuyQAMVjhxepWWv0gpDU1jM8b8L76H8L8wPNZzRDQl5fFy4jd
EW+4xaTM26MYg5RzzrUOFB7sc+BhhW23JuJm8p1IQGRjGdseTWIXsAjwKLbq4SIH
WFBtN/429GnYnaz7NjrY8zj/nvKxMZOtsxtSOURmRimaouKR9bhxG+crVrLVGoR7
drue5I9kLetcISb15SnHY14gSFbM4vFTJ2xieHoeWqli3fVr3mErZPQx9zgwD2tU
4VxIjDUJvjuh4O1SPUy5wgh413sPkgfKcLnjGHbVPOuGxZjT78Psb/AnIsHpZ6c8
93Sg0VKkh2Jh3hqfzJmYzc1Lq8Zh/WOV6wplaYe9qZS4IuqUV4aj0LF/GIMc4OBh
e4SAF3Ea6bg6JLDEjNgQSlSCZqyRMU1R7pZCsUTGE57f+GkvM1HyR2at7kzoRty2
1BM78x2XhhobjxEYJG+P2+ziRA9j4083MSkUzy4pCgg2Sfrl18OuDcDvxo83pALI
kpvGGWHwVKzyVuTdBUt7wEIMV8t+CQymAXvCV32g8nm5r5wCq3qYFLX0d0GGlDKI
kSoiLpbj/3Qcx+Y0aR0SaLExeIUiiwk39yocXlF4OZLDiFqDpRn2BYCvKp+n9QFc
CSMNX1ED4pdi9R/r+gbOLDpmlvZupRDwgxgIJ9kmAUN/XZylke1aqfxOd3YmKaGt
Y5GNiFcnvI0p+5ZqncW0bwuoP/2A7kjFFk9ca0CplGdBI1WO+6+yshahEUb4fjEm
cHTewdt7k2naL43Xf4WhWi2Dp4M18Vr+4HY37hXqN4OGyJSLyKv4Ob2NXFJsjCbR
fYhXWDN96H+Vf2tP071IKT6Q9YrCaBgguQgdTNOXSbHBaQYzjrwP+I3QF7usZ+az
0r5Pf8VD1CtJn3NoH9XtP9gbf2kUW3DdnRrtuqWoi30jtTgGFJW8tt8us1NbJMRl
rzE3TZwiF58YPivm8AfjiLhHBD4i8Q+owNrXOg57QkPU8fk+gzcQpjcWQf9E422K
IJIfZ7rIIW55vv8b3nWS+R1kwLEi/U/rdrSNKqndnmrX/yz68kQshCmSW4vr7Pgo
tIKXhW39gD5S9jT9JuFza3ltOsypQIEHSsZN/1TkIBgVftn8qw+qLZVU9MpBsEYK
oSh7Uowf9+dmpICOhNMeVp7oyTYQoAmnUg+sBeP4HD6fijdsBMKHljSV+bYvylvA
OKRB9YZpkimHYUUcjHs3vVQflpMdRLlXcYfP7Mf3JEByWCEKAYttWr/sckW3BMHX
/ovgGSuUFMdpCI/gJDmVW8x04mR4i9IS2E+Bvf4MgETaBQKiG0vaRRHlo7u23ejB
8BX6rCF73t8xG7d9hCLDSN6WOOWQGKyO/GLK7G9DSGMti2J2fOPDMTGyxXY0lUfX
B7ma/ZnSvg8bZErrHMnFBmaS/NjBuhBf0lxuliK7VGTnz7PvOriGR8vVUSysNpcz
tP1lC9uyKnm9CX8byv2o5/9eoyJnwqmaVxgRGUSYyuTTeaA5Io5ZJIlxRsf0vA4x
Dl4ZWzsf2sRNpS+xBJpDY5wiVMg2Uo6cE6kljPHAijJ6DOxHDLlRkWJIa1sFNSaM
DsqIZgmku5Jg6AmicLod2ByKATWWvEQI3Jer7BNdpAbSShWEcIFt+JBUxjU/PM0N
czXMLBBWvWTCnkftHVEwEXuQtSs/VmhiZSbJuB5p+VpxRVNFE2oi9jLCSWOOZ4mG
pSrRP/mqdiHcVT3Y9sbMC3luAzGxSmiaMLrcaHNmb/zj6Jgj9UHXJ4lHcKS8tFVM
Rij3IIiOBScAfc0noVo2IpAhp0Q02ock5eq/NbDstsieShG0kWj1Er/vWyaUKbfw
o7AAH/ZGve68ftbcOiicmxITVdYTS9aj26AnsGqgThZP0f7djvpkQP0nrqEQAIY7
lPjLpFgdBGKxGtrbajdIxWajTfoXQO1zJzSHnH28FXYOQP7hawkOvHKoAlCc9gBe
wS1LcerybCxij/RFl40eZ3xUhCDVS1ZIIxw5U1PweuVsvolntI/5/tDh44hus2CX
R+2p5TOlcqLlhALYgUmhwDNuSetkF+jMGLCOczmeGpZ6cfV3gFvscdcMk8ZzGDp6
Bp1AL6ct9jmo75c9UiW0meNb2njCm8hoJ4Zj695UlpPz+0utTRoV6sHsnXLVQrNo
aSgnoVVzSAYLbAlJtzf+NkQVeb5uh7wUmK4eo7vcBTcTTkdi2CkpGMcjspdxpPs4
YLJy3A9skcRYtBHC+xN8HZUFX8e/T8HjaqD/Ck6mkFnrn8Yygjlyouq9zX+hcv0c
1/OCyVOZw0xkiY2V9D6ZroGFXYtTWPUf9cRh/Jd8YLzTLwNqkL83YZklxtGEQmKF
smAq9NdVgUefmTLmjN+H8CfKLDkD6eQKkacGaTjLVYF0iq2EdBdCXtDYJmUiXv3v
sEcOLwaCztkoB2hY+Nxo+fAb661osw81FXGsRdJu+WI4Xh8ILRFlxy3kAuwRH2JO
1uqpmu+epxWA6D+efUglW/Twex7asK26udq6TOEF5s+v5+Lf6WrI+PlLhuIfGPMc
O0HWvca+winuTDbM5ef+2AqYA4TOsyK5TIpdPFsah2kNiTI4WLMWEtJQA94LnHy1
xzb/EVht0S1GiQ5y8r3IKzdfPo4nT2kYDcOe+Blusirmj1BG8y8ZJQHgROG2CmHC
QmFcDssDLBnmi92lx+efsXYHawJ3wB+/TE7cQz3EmpThT1xJMO237vPtTxsuLUTR
n/g4NQ5CFsW+UMV+GcQu+D7sYCpSmTlTtqfUmMfv4iMFxdfsNpygFtOeVzrvISjg
Bsei+DhVJFXUlSKNis1qFIwWtFOB60LCD+kwHJl368+6keiwy44RuQ7xFethh9+Q
mMR3/3vv8ue9uIdsr3+sElz+T7DfHuwkyR8Zk0Yny73Nws4P2HXndGb6iWcjuJDR
tp7L7WwOL2lbe1C/KRRcZRcGRuFMxdkVuB9nRmOr9C/McLlOwmLmlB461x42/qmL
I8DvMTGIxVhowqqxmhpagamj4V6TaazGMJT0EtOv37Gmor1LfD9eEGcQmY6mskQg
BVE/xSxmV9Gj60bREBIgTIPL2QOR3jM0IbNl+ugy0kyPJMNRNGqL/DurOzmNnegO
WxqrME4RE9mrfCRV9I4vQ13LFvbkzPs7c5Z7LkPE13QhOufBkzYMhAwcqIOgnZPb
XV6n0obh/RliRLprOO3EltVtTwg/c9haiGdHwy7InhQKsQJV3IpUSfuEjUcr26so
PTOAk2O4S+CBSoaPZLOKAVZFnoIDAw57q8zH/ydhdrp9Nhw8Q2eaWk4LkebPNUyP
vZqFDNhbXEibm8oQBHLjlnzPI3URp/iBv2nmDtLmtys2Xvvdf7w8RS3bg6yPBRdf
F+1mgcyZvajbKtTVlsrUbM+dbQi+Qi/u0rGk/Guyj018HVf6n7odbO9Yx4Mfo977
QdfYKCv3DoCM354kys/DC3MsbJhTXGeXO2YoQpBMkoXaWvDN9OJTFZHpQFcCJGS0
tvENnm8Ry2+z7F1t9ZmlKVImIDW2WGkS++dL3PB1OJe8XzuA/ZwceIbMYej4VvYO
+VpOyA/Qik/WHzbvPr+0johgl6m+GPeN5O5RF4ThZcY5KXPsP5vItGKANWwIHY20
5LDD/Qkpzu10+TlldUGS5YAGeWmYzOp10lm6oHjQA4j+wPkf5+TF5BO9je9c6GaJ
4Isg9CiRWHDzX/d4YqJNS50UJPCpdrTRAqYvM5Poe5vVMuDuvHz1DWAhUJGLw1i7
KT63nOo5WEfwQSNXxwjgX25QQ6jIZqx4A+HPQEvQOraEkGwXAKJwDMfC1WdHqtKh
/OXAyMJkvgLAYPn5X6LJV0ALjU6Laevfiz72kqG31R77iqO7Me16IRWNc2mQ64m2
aJYMMfZMReKv/R7LSBOGQddMLWuLOqh0aaaJK8f1CDDPj9YSsrG5+W8n6kQ5+CLh
H7M4vb+hepJ3OqMWsORCnbGf0WDDHStXiO8WGIKxOtcCZz159x6AGgpLdjMaEBxR
/SmuMZ1koVvM4sVdMaDDzcr7h/906Y+c1QzzFEdumyACbTvYvkCj5IqKgkQn747R
4YYmmqVmUs5jWmrzf4EPToKqzRoLUyjNijtoitRnhCsMEsAlFe8okuiNPhtE6Ixs
NelVjfokn7GMfuL/HNKQFaoPMYt+bQjujcwZgJNg3nuwoNaG2D4rD3Ngq/uQc47W
tiRaTV/9MBy1Jg768rOzalQYqk3Wc8aGzdWZQQfirMPyinU8zmR6S1oj3ZvwmVff
kwAKzuKJ8AY4XLP/B4soY3bMRYfYQD5OIAGf7sDBDdt559OquQc1jL8MORNVG1QP
IZW/0/Wzp9ib+Oqx3u5mmx48zU7gHlvXENGw0IERoSb9itlyuYL2mqyi1vbDtyt5
nqDNf3UQMDjIcawTgyOZGw93jXVnPEntfVnur/RRD5mMvCkg7qpj9+PHonIjlaxx
TABn2HC1dPvzj3t0Q32HeXHE6IlLtGTFX87jTCIaJSOZDWbGR62MljlRtWzr1uik
LB/pdhGJWlBh+8wpEsUvoxGOi18at3lTlC6s6ImFT04j/mGWFSDdXUJIBCuG7TzC
XGqaXyV1DdiSH3X0egSYv1v8bIZgfLkhWmRf8TqP3zDY88sMX0OXHnpzwXU1Dt35
KdaLKFDMdof3iGZaQnrPFcEYKzd0ngRwihx0ggoFqFlxK8L5yU5FUN2cY6fjV58f
Vd+7rXWyAxlljmMYIdrRHWzjfGhrIWyPCBt5Dc9MxQ8bBDrYlddq59Cng/E4vcEk
te90rJ5+d8s9sgSkJ8KGRytHcH965vKfF38vcVBQ0sy6KTr45l/kaniwBKMAa5RC
A4PsmCSAoMmizjcINK+hW7UVsRdt1u1ld0k7PBtsdRag3koIoCgGRjjuyiRnMoft
QSzXtXPdkfM3vFFti6ueqwJSUvIS/GoD/X3KRLzWCit3Y+OxtQuVTqQ4SgDGP1Xs
V7F/pVitVkJEKquzIM762pXk5S4ogsC2QRaMXXv5FLy5aYNYidnYxl+vaoNpggK6
Ja+HaEPu3Jl1rp/xXCtgscz0FxUK1sIbZl4MR5z8SU+8gz70SKtqtXA6Xi6VdN23
W62y/yQNURieUGnAWCf6eVsru8KhdMW709kzbU+YOf8QyN+hRmA9hRCh+WwF/Jf4
+O4DLWxSwcs8manl2dqjc4aPO6L1uoL+WUxBPfBk71xS+YIo33+EN3S2nkwrt2+N
vjJZojNvltdmTbvACh7DK7UONGrz3vfIkwgxxf+/fIRZ2qDo65c7PXfhddcAwQky
9lrOegX9+x5b447g47kVNXQqpbc9ZjhtSFZNZWgyPza0k25JIp9bteGpU/9TvdFj
4rTmTXeIyUxlDvrsGm5I1H9yKVBYwhlsNxHDTMIhvJk52NKp5teoFwpvFazIHy5K
hAfxoMF42ZWtdsFnvO3AsIEE0viu4dsFIOLvcRQsNlvy/jmEvsXE57cZmctBDuuW
OWS2oYkoQEDH982CElNfs7y7Vc/p6vQBeE1tmCiHaZKUUR4SsOcZSEL6AevBCUJ6
vz8SQAhCrUYzkArfCv9O4agnxhiLi1eiR1GiiqNKgKJeTDt8WIHkaclyXZSYieUq
Yl5ZP4Z0JsazIGNu+f9JkM9WxP1MW2qk5vaFgY5WbyQcKAl114f+PVEcDh3/gZlh
qMJU+rvD4imBaDeLd6fM2fv1iaww04JBtR0s82eMJ1LFBrV2vImPoE06vcTbnbtE
sg2TDLTy2HB0+B1Fs0fMufCK+LUAEEq1o9yFWh/04fEGMF/hXnwk95uSCyZSknoZ
cOvSxLmzKscKNnd3h/GsIaXFv0l6R1r/wkVNsh4wWZHMQeQZJ1I1Pp3R1nAZaarZ
BY31FtdGYgohM2HuujOWYr5J79TVKhKZ78J25t6+luwKtxxnfsrRf8zJbJzUwc8Y
n8ke9kcTDEToDhvnWDkM347ygyZa5l+qHXS6EmA88Q1s1ZJ4287Gee5i9ZXOvC4g
FifYGY3SVZrTnnLdUMcGPxTyuQOwcoSkMzVom5MbAfnCX3/Bk/O+1bTcuE0ZmDc7
BO7iTvgS0fcPhufYRgOGZ/GuyVsdFWgbrQfXpwNmlOZg99jbOuSkY86V1zdDSsLI
CWnD3DNDKqQb/eIbJgUeE2zfWMyEyGWDhNP5U5ah/YvidAVXsy0+qtynK2B8CeHJ
biA6cRJdrg99Ie7rPSVNZHuNw7WayS0mZ3jrAvHd4vHwDY9+v2ORmUwUGMJLtIr1
qZ4UwaamepYI+v165Z6spOpKWwsfNX7YOXURQ7L4gM//l+zYIKFyclrRh6l1zdf5
XF79vw6aF66iDgZv9OiwzBtW+6hd5M0DP+ptWVRcrdWnm48cUCfxD/czOBjNtB85
5pVtDvta+wHZQJBRghx6AzRZFWdYyFKk2udvx9XmMqDSeqqOi0X0IjQSasc5hrMe
yqohbF0t7u3zDQ/MpGBAOlkl7T4E3/z+z4NqI43ff8lPf2glJw+5GpWzka/4NMsj
ExooKOJMbvxXQ3ZuOG8B5qScniewrJvjS0v+2hY6/fv27KKrY2lPIIa7vc4b/m38
jPuVlJiSC3vC81z7s9A17NylsxVc6VHX2JB8tKvhLolJzG7X5wdYb39OeJqaDnAJ
aEJrJHBOH4UT/AtOq4JGgPbnNjFdyAOpxNeGU3jGGSJx7BwS6OLRI73t3u99xK13
iPWht+Jf+T1uddYIx4QH7l41scUYkMG1AI6xJA8rfXLePYTEWErq27e1bOEMg9bX
bbOPNphePFKjRNoYeVSJioWbVWRi/oRQY2N9Nu1lLRECDjlh9tXTlgN+7P+ez9fP
NxMS+siZm+vDsgslTW3aZ4PFzSHIHG0AJ9M1G8o/B+sEyoVcb62ZSpSwiBJ4LRjM
EFiS+yI499oVfex+VkPVogxckjGYA/eEt90ymnwtgd5u8E+P+Hsn4oqvvwX2jJk9
8eGQTl6h+1R3VgzNmk0zxEfTUnerFEUO4pksEP2NfyATi6H0mExWIb72JDXLxaL4
R7OTfPQQa2mmvIJs96h2o47WKhYrgpDffHg7X2M4eBTrIaUGaPgM/6k4tqzTiJ/Q
CX3MNpcGMGc7NfSmMLZ7lNxm5S6XX80WZzmTxUwbdMXZF/kmbC+XbNo5nbwcpCxL
/lbaV1DSjCkI3BpbyLVHK1miE6hQ0RXGFKwf+SMRYw5SBr+xyixiBfrB+wVx8DdX
emslm7oiK0nqeMRy+6ueKrW9t1Ycp/Tvm2jHFIZGaKftS+JTen3F39PILYvX2duZ
qK+ltZcoIQ3PKlzDaCasqONFndkAMDWi7++q3KSqXOz3lZyZeyKSmEjtYkZsljDE
0/5zYSXV20q0RgOwiAkfZ4aLJ25U/R0Y8f0Ci4dDt2Qgv1F/qWJ5wgBiQVRmVbQx
sar4G24OhYvl2YLhahQc9EeBo/kfSzZF0wCSntkoKOAqHce58p4JYTK/ugFdHQRx
DwlW8vu975DVOlQGAydlIsaim05XGhq7DbEeelOxjWyKwcIcJojCtEt6+Ca8f+Yo
asj/tbPWgIQKhzRChTOXgixfOcMHB3/5iDqb8mXAFySOaNlQPJnOlc5ckU99rngA
ZlyW7bA9ARBl/f69G3xSOBlVwFX9OK69Pw9/mHaVaHCaDuIvGi7rseGAAmqLvThp
MdsOIidtUcZ43RI8ndNFUULJb/dL580ZNO4h4EqNquzliqJ0prdMrlaauH4P3y2e
JYdEGjcNGq6OFjzVDPVWtdz+wdo6HINrUVef481nAcrErqvEonAbZFfldzekkAQV
ZPyNi4HDi0emk9fuEUyjBnfHGjj5AAh9YS7FiQCEJwhcxSNqMftn3aw+JL/6t5Ww
sjs26VgQ3vvov7lLnEjYGRv5A+yrZPf2Tmf99JqMPr68nHy+WxFFu9DFEvSVFyM5
MoAFJLWxiotyce4mFRer1VHN3rpZHRp6fBc78bjnabwIByg1M7h0YFBEZYZRgo/q
RctbCP1iFGpy+X8rmdtnToY/xyjpve0TQRZeIfNVI2pBHdMzAGKtI+cGf19V9D96
/Cf7z3g5TtHjgmwqAIlqfJRU3kdyvN9B3OxHzsDT86XbEKSN0wxBKpdEhpgJUQls
puLbW65AYeWjQ050rB3OGqSDD5XeeldAvXtuNAQUWcRVjBSNAC6vveY4iVVtusSo
/V0o+BFGdMPy5KT9kUJYIst6NDuwhZGjUHbpucu2Q7/7JuyNJaEwPWepK+2oIYTd
UR9BW19obn+VKGJ1lrmchc0qtYAPHKCQAAFug8vtY500+hM0N7fn1hcXZxofD2p/
uhHhlTO/gnVqa4FK7riaiNlsBHo6TzlP0ceLg/0/Tjom8stTJJ190vZg2qrGMIvk
MPEar3wU4+OI5SWgFKVDitXiZrm/zszxZoe37aHNmM0pBjWkwtBRNIFdA0zogpjE
zk895S8xW+W+mz0WUABs8C+B9/OZUTATY9bWxzTg5DP7SDfSkKlRMemYAQgff/KN
yFqiB3CIbXYB7+UZX/2aKRFhR1p8hZ33BZpcfjWGgiXv1ag9O+MgnMciZAAG/zWm
LNtSUVWNxI5inApaahGUdmOmNuwSP4VEcd9zCHNGIoUzdJUD7siRee051yCiT8MS
mwPrTXdKCQ0M01JySDXdNrEYrCS4VwHkPDvMb52X4xELx6V9goZaEdeWKQx9Clev
laaRvaV8FZm8Nh+1sW33ajmbERxmXWhpAcPJKiUaX8TiTnQp8RR7FhfvLgVSpz7m
sukJsyvCzmXwezhFxo1QfpNLJwsV1NEEoNqtU21LGOT7n4JRBPO9SjyDmf8kOAck
Y8vo2VH3t4M6vtp2AJ48XB7Bl00FEPpsLh3THgAHBI1qP3egpmr66O3+Q/qoV7HR
FCr74USMZEvDMSLunD7gX/1NRDe8J0C+220x8UtWn4XvW1K+e3/bh+eWov6K1cV+
8O/kRhpjRFD106jUxE4ZojrhSdM/0B25NTKrtDn9lxlb6oUqv99AYUNzLLyKNbO4
yGL9CjIbYk7Y3rYtg390V8Axldi7H/419Pjd4tYsa9YJDOxhV1ndo/t3SvRDPgk+
xiwNkXRcE3HfvoG4qoDwqSmRB/YQlnZu1JMKcOP0+0TaXCC8nB9GvYTXMTbfxQ3Q
EVp3sp6XdYBXJQKoira+6NRohGFhbGlxw/ZCtMCa5SD358PQxtxqkgbU5g/DqXSg
9b7Ue2rI3oy+GSburbrOnzMyh0rnrLpfRlcfQ45QHS297WcUdXLniLCrVSfBpS2J
6tGuqxWoylDmfGWINZ85sh/IY3Y4djR6GKj8Ie7Ew5NhNCY4CGOW+yZnox7Ehvpo
NiX7FQKG3OLSQEPHgncU9UaLE+FFXpk8dqdxDL2qsgTcD1ILJtQ0ATO0oAHX6lGJ
5OPFGJ/GKvUa4gcN7fMzWXB9QjLfJj8lAhYBEzComH5UIiXK0L5Qqtte34V+NpBD
Y/H9aKVD/DOS9qi/5EiHmhjSgqi9EJJMGIM+UIhGWE+nsZ7cWP03MTWaJWi1RE71
SND5LA946wxCB+pnMGgScDESzqi/EN5XwbMB2TJwKgVcDUTW8jNCszvNOasWPwxt
ykJjKtmvKV7nGbfCG8DsJuVmMKSDoxiZLrBHP2x/IVTRB07h1fJKxFy933mZeiQx
GTd7uTCU4Xc6f/DMtuN/sR/SGwC92zBwUwGFMfvKjlZwNNbnB10UDiEw/wEtgWyy
l020vAfqxwfZBUPOxHqMDmp2m9IB/S8elKniv+IxwZU6hj7X164wCH03+Ct6jFeY
humRaRvf1k/IP5ethwwcMC2IcbiiWIbMXP2LGFxAXGzGEY6O6macuOKp1GMF1xJF
a6fBiCUvcvRWmcN/O6Y6PouZMDEAYvggrQalx5+zO88qOvY3l6D7BGTS3u1ZH7yW
KGpNUmrdb2jsj9u0P1orhHZzDHwfFvLWj2WTKqi1tKFQt3cy0BnWQn4Yj4xi+NJ+
huu/8xwakzZhhxUGkWplX1qe0rlj6sLBllEMf+Qh5MAYlFoRkO8YlzodIzjF67zL
UMbKWh7/xqo91TchhLPD9aGumb3dDkAuRrQw8aochfIRZvCL6Fn/sl3c0yJGU4PM
+ImKyriU55UFxdZR2I8iG0/Ub87yQ3Dsrv79zZ9KrFj/15hld7DgEeYIjW07HenM
9ygkFgvERnuMDrb0JtVo4eyLbMvsz3tjHfB5nuM74Bwcn4VZHbj53i+Em9fqxBzE
nZkZNl6cWkY3o0/+mLCsG5oOch07XPFChd6mSRpNc6NJ3u8uiRh7nlQd+7PhCc0O
mVrkNc03UxvlvcZGE7Z5lS4aMkZx13+Ev9bhj6RD6LFeIu/17p6qdSVQHuYGRb7+
aN9LZx9ixqgfxwcZw3hnin0qULr9cDFUhJvGR+Y+B2ZWEFH5a1O8+HKJ0c4ez0Rm
HdpRdO9dJVjtUGCuGCXCfs3eMiCnxd4mWsRQh51QJ5lop2Q29CSrtaPRLpVcIJCv
HMf+VlzvMu9KG+I97Hrd+ILOa2Rwh70IQlUTLLEmP6UoeV3YIp2DtF9cCCdyN6DB
076S63b1PvGry+NfazM6x/aAPphhcxN6B0sWHZY+XqwJzNitIheUdW6xA5swKySv
Otih4yCutT1ZkhlTfXb/hxJcey8H5OCkZQkwksNjUat1V6c1dQvaRzdBDkRDs590
XspUl/IhNsMK8FhK/CIIJM3bryIzE8dmlJJG4JYv5X+g7l+gABP6144X3tB2mX9T
NP0KdhNvm1oY0vQaC/NASv3FhHZLgPntyl0Qszo5/yRFzgXZdwRtklm1Y7Bb2M9k
orGmDMSYyHEQtPzdUsVU66qSosYggZ+XxQohfbLnaz2lXywbW8LSqXYzWNdGDcLm
Ms+bHwe6gccg/ClpZEpW7n4gyRTb0VTY9ejetk5fr0aTzYdJC0lnuPdDzwPoeZjB
+6tmQNIS8kV4eoUe34pv6iwM6BlUdGgzvwyThQxS1KZX7qRE/XIJEs7Pu7F3at1Y
Jg1JfeixKe9+MAYcHZ9rTzF2eYR+k4bah3J8TWMlGcmIu09ffUKaqd/OLub0ODU1
yFzmgRqStkONwnoajFK+agOg2iDZH5Wu5is9BIquLvF5Sz72KBF9GTYPMzKn9tnD
xBC/GzeGxMGIaML3dM0Q/zgT46wyTuI+IVG186JHXrlUjPEgVuYHZmDScAH+csCL
K9t3h/UUhW95gHZyglRPVsS9W6sJ1k8WTgYYWz2v5TpL+jlP55zSA8HCugOt2qPJ
x2D7LQSNf/Nhe8JS4g5wgtLC1rkB8c+2n0QO+ysFDoY/61t/TuQIFH7US25BdKiA
9BjI/8BnWasgCMriMM+7/hJvJQZDlLhkH2J24v4lwUse2+BsyJC0PJuJ4dVIVVJZ
oHzTtk9PK2Dsb8hMCS2IOvGqgi+ORVMnmifuQ/X9knGXiLcfgBEkYq0d+24nUXdx
vLSdNaMELW2e5/JJEyS+vLkLvjZNbntzW/nfK9vpI8kP/vbQpoisQJnkpkoFUZLI
PawwggI4KhpJjXzmqUS0RHw7DRnC/byPIaSuyqZq2xI0qJ0U0p7XlOoM80mOwpkX
mRaOhoNi6W4w8tox1iw1gOydlOitZ7Bdg6mB4zBVTR0=
`protect END_PROTECTED
