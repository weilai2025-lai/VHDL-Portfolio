`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHmjX4XFJXXkgXWoVuI1FfU9+wcNP1dUO5E9bRPvjwWV8ZscJeQJxF2hUHNXkV91
U8r66RhUg23en/5YCER8Q4CniMxHCJXirspaJ3ON7Z6MXh0Tq1kt74JVoUwNHMED
oknZQZSqpQPbOhLwO5n6SIUmvFtYMHGsIzm5knPM7hBkx7J92YykclWz1NK1K2gA
o/9dhAiQAPPb7VPg3uzuXzHPS45pYOZOmTGj9fn2ZMP1Ob3DCCK1KvmXMlREn0ZP
d0gKPdma+RkJfO95DAXbv9SoHskgFIkVOHqK+z/98eIizHSJn9YCfDUeBdz5i4hY
g9e3ZwJ4ekK4jClEoXBuvgZd88dAgd+gaoNeGCc5eISGpr2qdxmztB4theFKjTqN
G75ldfin7QDyhZenBz6nHge32+X9hl13ylm/0XrKdcVU/C7GMJNB3GYIP196ol/S
nxYNuB/mBgsh9NhlHNlSVOq7P8zz3rXCH+WfpTWyGI8/nMD7uNNdrs0+HW8a5rsU
BRhft/9tOEZCd1ORxMYM24hszR0lD+Sm35mN2xEUxqje8dwmkYvsQZsN1/1b4VDj
pICsjrJEYDnJArEml8L+h+3PKKnbXXu88p20N21b3ceRPb+JSM8D0OSy8Bu9BnFw
riwBuZ+xvHSmOeRDpWZo/+VnQTRzQs6pON3aRLBb1KkSwFfZXd2i68E86gDfUhUi
JNRGbngaMK8JW27WKB0hUXfM6Ga0i01TXSUxQqrRwbxIYfvuEpI/302zBgEIT4M2
tfRq92GAtb2ks5SCtnKh0XjIJeb0ljb1mbAVfrTtE/TXctmnw8tbLP0rXFshXdQL
ZB04Nid1e8195TPMo5WlyGWRMCeF7WqIw1xog6TS0P7zRDHjmNHMPRLIJ8UXAqqo
`protect END_PROTECTED
