`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPtQG8gHKLQAN7CT753JoPbVNaxilnJrSc5Fgu4OrS6R4rKPMM4sTya0B8oT/sT2
AAC6SyPdaIUQyz++coyPf9BWwgVTBpa2Ay1zMY6drnZ/tBYpNCnYZsVUYEqP3XV9
gWko0e7ZVrbD3YMqJYBG32SsT6VeQjuKipXG/t7W2qEKhsp0JE1RNYYJXRRmQi2J
c81SSMprzjQJIk1j94rTfyzqJpiF1a7GuKnSB6NV1NGD+Iqspb9UsLGSKt1ChSxj
NHTmL30BiOj09Y+wTp0IVTiQ9/cyEsAzWe17GLmiiJ2av5NRN9k8kTIYvyaBa5W7
wR3rK38moF/P1ijyvVaRC8x+WrySGICS8s9grqNwBzCwbikNeZiDM1pRtlxam5er
C32xbt/EUKIlW13vWBy7WXzaHJWGeYJ/G5dSWNR9L3nUzQ3/3KWlTJbFtIPlCl7+
+whnEKC3A7Kf1zi3oDaqwpv56PjbtextaTGd/Cv8G9pXBJz8qo9sjeA0i3nA5/Ng
tg9lEBZsF9OiBgf700WMLQZ2+wKCWEQ+HnelpZrm6KcnpaexVBvPzMfiqdFOYh0m
5juY8z7S8VFFbuXiDcWRPrhTH71sPeTUV+O2idxHYVTPB+NhU0xAlPabauFbjC29
r6WBcvvSoFc0R1ILVA9KBZDOQlNCeJUcWhnEKr4CZppR2JQupSblYMvh4KiNYOYx
AjmYr6lY8iv3XAW1ectp4KXN5l6wQmP0qa7HIadzbm1HWR89bVs0qiBLHQo0B6G9
8MSgmjekYHFJixKDH+9UcYY/SbtTqhtQ6GPYpqK0VlXqUszP5VPyyRoLRm8WnJUv
gaPAJ0ROFp15Nma3/0CjX4Aa03cwolV0GtXDBhfd0FXLRtdXwhemvtrcI8iAZYd9
SECGqJDI2jZFs9Mm8keB4FaF2bwgdYttZtpG651lua4p3dO7xpinRWOrnYphPPaO
OsO+d48fG2tBx01F/oaWUm0rdEYHo4FomT8yiKXiv5nZs8X9odB2s39n8bo4QxzG
mkN9mdoPMfpq7k4gZrEjOsFijOe2ghHrGwwAXaGWSwLvKZ/EvRo3e2+dDk56zcij
eElrSHrybhaA3b16BAv+sEnTyItusAhBOcvEfUA8OkMDRe+Ye44bRBes9U6YB4cG
ANV1BEU0GTU32wMm+tZIPkhSIG0dlPXMW3Dv8jzVFx8Wg+fzxjy6WPoDxcz/pg1l
/er1GokgCCs9Xap9D6Wd/DU9SBx1Gtfb9u314J6IC48oORK6aImI2o3sJvFGX19a
MZif8TnF6vBO1+UMBIxIRP4WHIj81mZJ+cTYonf6YM2BC8nawYSGvGhBKjlYOI5h
HPgV3gRQvvt9gPV0zqlNoVSyTgSl88WFvBfDDYBl/flNe+UtgyZj926fjftEw6yO
5vu63UK6A2/WxnLkf2mUPItUUQR3eWFplmSXw7QAVuSEs1A7LT5OwV4oRagVdhA3
XkS7tcKZTbRxUb3L1pI15iwwM0h2deTFHFODla1CBS0FcXSRbVEqLp2O/EDfn12O
RIGqyeIekx+yZWgrXb+h0PyaxSDVHCxNWUdnlLrb+CBKWjuZb/PtVHEazFXazQW3
mq2/tY0hrfdchYM7h4EMEJ1w8NhnUkCgEk6SV0Rgay/oKOZ1BLto3vdugwNePoMx
HDpeN6KSEJLhN5xuUqIXbwDVM6Nryy0DfGbWVZN8XEyNyfR+LWw5wSfEbX0RE5TQ
GT4gmJzvkfsFYsdiTXk9I1qJrwxjpO7SvW/anngTgL4Wgbmfwf6BSf6vCVlRbF3y
3/Bf0CGReOKSi+IKyOFK42zlT26URPKBrGeQQ43hrValqkMvQb6t3dVbJE/MlYJr
tQ0wtTgGReNEYno/wl7NguiCf9birLqEgjlXt1x4KEtRndGmd9OOf841ID/CJnc8
WIRe9wbZoyQvabfpuFGOxUaMz3dLOP+pkTeT79vTG8yGijP2eNTSL+J/ILZF1gC2
ejnsgOzrTp2sIVLwYLjJVIiUdfn6uhBT7hE1s0g4a9HtkCpZoep4Pn7VrsHcNtWU
0iQxJpGuRaW161zlPZ6Op9wAZwnEn9mnrjVfRkIiTpTQzoSF265viOIWV/vLWK76
5+seSEfDgNSEXtJ9+JmAR4VM4VtPeOcxbnIlaYsG5SZ+cf2OZSL4RcYw4SIwFxXe
gYLVmQ1aTX1psa1rjJl8GkWEQEC4OhuofuXCfg3Zd4/HO3iVpk3xDYORAw9PHz0/
1HZWxEQLVxyb8tH7EAfWrw==
`protect END_PROTECTED
