`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYgI3rppml2mFtHrxkmmwBwO5Av1mD9IGTvyfT3xjJRtk0M55F+U8U0scli+rlaZ
VkgzdHQ7UePsmhL/HUHK/63Ww9YFKa2LgOOFPcrUhsRcKf7XXg5BZqo3/bf0qE1/
jrjBD0DUbJyg/nVVEh85xQo7hec+tmQUGOZDTcGJo5d/8nYo8H0DCQLgzp8O+tkT
JCVmFiaeABi8/4Fn6Vd1V0yIlH2IAvK1WnOHhN4shURMW8vhXK5XzT7Lld5ppC9b
AeJ6pl1/It1gv6Jt8stm2F76MZ28qUg+ISGseStc0BGVCOWFpRzItplWADBT6VdI
YuEHAXN4FrFyG/6I5y9d2VDgrrvo1+Q5B4zd9I5s3UPq52cJP2Bg3LTScAkQ4ti6
YOpQnm59ROnvUaJsMGtgA5L+YO+e/6bjlBr7JDJXytHPgbtof1FG0TyG2BPBu7wK
9XVecLrkFzGLUQdMX6ncYCXGd5dOlHH7EfaDCmyKBUk+3xf2WMpYR6/QoPtp3y8R
NmWQJoFKdmSwOPjXgaaxf5gPhop80O7ufPUEKPgbY+T4/F3qcfyx4UJmmEjgkeWG
Fbsz7dC0BT53DsC4T7yuP2VjOuX6HPWy6kjWuKma2gkmfKwZ2kzUGlObRNG8kxnv
ZHM1KMVJkqdye3mDN+RtfvOIJ6AJFuFgf+f3OMjggPfyfljMZQESvSjldwysaOqP
RpD3a76XvVhKe3Y/SLXAA19o5BIXo73SEBqG2Tuz7uexi07mdD8jbOvBx8gEL9oF
PlIe8ZfhVmQYf5I2dwGugfWDFXdYR45QGGnGtalVke76YhYeCVzsvVMLSxHnQU8E
YbYYfepZUiAh5+N5fRCKGuEsMT9HL/T4QO8Q4LSA7z2soZK3IpSiitzkMZa38KuV
DjRGq7WdffE0ym2JMf4D3cF6IUKizF9I8PBxxsIK/BNtWugTzVbGusZeNWlMwls6
ItAbY3FYnEGqrMm0R0rfL2BNfncyj+DE8cEfzZ6zNFYFcETmRTdALLx4BVEdVASP
UkfIBQ0SsqZ6RNHAJNaQR5sXP2W+q0R1GvudRXvx12sSRDlp9McVIXSp31hfz2b7
0nOVOur5ruMgIWJrqnaJ2jyW6rPtNQe/7n8gh2pFsEO0zshRw5OeDZNNBvV4fA2y
FU+3rwPBT9/tee0BYYN2mXxTkiX3OPoXCMVwqRGcxY3Y1vDOCRhN0olxjRem3k0/
gQsdE+MWTIjunFOreqwWSOBE54HtrIlYZXuAE31O9dOq6NmrP04GvucBGyHTNVAg
A5VriYAUqWEMTTpxQB27A02nrSRhpHi1KGgCwPRRUm5dBrV7lTmuXBXpdVtS1P9N
pgMXClf8mYdCmaBUimmI5NuqjjbQvbL4qbLk0y9ALDE7k3yR/BZu+5kqA5En4nqm
tn3D//j1HpS6EvktpPVZBKcwRUhBGSX8iDPAWZykvNvEfv+zvQl8rfy2qx7asfnN
UWdxyTGluTYYZ/iy0BVD6EKWqselfUceuQZ5m/dXAGJavGmlzMLivV/ykl3UYOWI
cmc3yphpFwLq41L05TeiKic+EbEy+rp3/Gf2rtNSJoGHSm1/z7YaacPHNVXX/dyr
6g/oPuJ+G8vjp8e8dSkLu9L58JtIcmbaBL9z5ps+4MWUZqlp37Sk3X4RciR3E+Ge
FikXyuLBnwn0yhKLR78TD8NuFq0fqnVHx44+UTDcoSOiJINuIyrVhI+pQ67y/9HF
9iEymw1ZytIj2hMaJX5QWelxy6E98Mqa9xAf/RG9hAu5yjOrJcfKBaj3w+HMRRyI
69o4BV8zyPEGiohXjI+NdzGIRw9zCN7tkpDnQMa2cRCZB0iecE2ajQLpQ1m/vCkx
dW5JdY8pQeGqFWPP3HfI2dOii4YqU5f3B3G1xxtx3rOGgabHCXq2UTHMuzJvQtHM
RO13zXd+cQxppXoGoMBh2R42eLfuma07Wt0Kw7jpdpaQ05KarE8TseGLIlnXj+QI
SJChqX05J0BuMc0CFqyOF680PFJ6fBEcdzSvQRV9eJO24DloCL8XA/afuEFb28HW
oOma1piy7LOzlWWJVHd6QRe4qvDIYwP+wMrNq0w6I9ogXQU1I6QAZ4cNVD+rVPiE
1scT2XdgfGRBRc3jVOSTK7n6nMIKZ+Z4yBRJG6uoav/46+uac4Qh/tZ3PxKvx+93
lXTopA9w3ZlgPh3ZVewGAWEaP3lYQPhTuclRAWfcZ5Vf15BqNd+NyYONCJ0XhulS
R5Y9jNp0eZQ4Gjq0Jcw+a7gSlb3Q32ifnbhLNexP1/Vrk+fE/csdYQcjF9+TMIVR
UsPeTFF0teSAXqUw2XO1WcjM/n5AMO1VmzHmsoapOxP6+wqoK7OuX/KR72+9zW36
d7nE1EjxEpTbqM0ghAVm2MdpLanYMQvGihD4VznAmT5L3q2XeG2NmttV5uexAeSR
Sp8OTFsIqh8CAwmfmpnwKXsVT5ccAxVbmYBzcByfSVIotVf+rxw/5hyPCZODGlEO
HNqLGyu4W6mjQYA4EWy/pgbR/RaA6a1yS57fOfgxmknoTigiOBIc3QvR6723lepT
vPCVerbH7kBQNI/NlKEXjx5sCHEUpmGtH4qek0HcP0EdVcgw6gOILucAeH5O2eWH
YA2f6oyjx6kjp2wCmDCtWsxcJBS1ibWz9u3RmtzBV/cJML4GyMoEx0YlrICWGdm/
xH/AbQzvxBmct1iPkHU/o29c+D0L7PNwYZ9WNKidOuTPhadUd65D3pHL1Snda54M
nw6Bw0DteIRZc/VzMIUCCRQibas/0KobYb6i2MiNx8akrYemTml6Fq8t7GtjGI2Y
zdJOfF9wJSD/tkC2NBhO5b8BGaDP5A6xfQ9SD5ZApuLwYAIgi2oPqpOQvtx5BWwc
DCaNWY2IcihbICqrBCpMF7z+XM8NRyUCIAPSU/2pAqa6HDKSIB1aoHwbCBI4fDJ1
5mMhbdXjYpVuFiwHer8klDwQ5+jYiuN7ZUzj69P3hiTm7p7VLziV/gIZBL1tf4jy
TvYXa3xY6cI7fY/v1KLt6FGTl1h9XSAEb1qD3ORHQ1ZbbmmOJp9lXyBcsLbS4jDT
jko2AfRTj1QDC7DRtR13f22ZeyvRg6tWxs9stQzcP+ROa5iqQW6En9H2a5Hdpngw
o6YdniP31uedACPhIqrxaMue6npK0+oE5Mzc9KgupeXlHIyfEuThXPyFlJtri4BV
QVHHqYlm56qHey+4Ot+xR9rZauTBvIMuhdwZ7W1Y9bSYK42oIj7W9e8AlMmwwvKB
/2fTrYRyt+11K8bRTZ7XdxleI/3GR/QSgSdyYMkke3L48NltPAis2JWrgpoDckRB
l97X4cXZOYJxJ2J7Wt4a5w1zc5hT5QDnQOeNJmg5yAD9Ait3L8sybVQKqZJwwqWA
OqAw0CxjseVJBZYXMCGmMI2xCqATXPLTaguh4vF1YsTTM+OGvhUs+dmsd1GkeCdJ
/Mpa7YaYxWRQnZrMoleNl/i7HRTbh1dzMAEthSC5L/M7M1QAEnJIFOn9wc2/hiFQ
1TeV34Fl/JksHt0+JeIvnxm+UTO1kKY7vlTsk+Gy8l/FaMfkhn7aVw9tM0V4sVul
u2tMVKeuqGQp2pW2BFZV/uED2AJaNFxKhv3IIQY5YLkCYig6CwNg3+o+1SfIa50/
gks4tqAF1kIS3lnwVfXNRS0f9S9PqJNwtb7BA5FBq+CI7qXuS/5C4KpM+sVL6MPZ
Wm1QGFXQvjlj/6dOgayM6CdP67HtPIWJ0mxFLsExWHObIoEPwqoVSEvvNDrlnd6r
dlj2Q3JFwMxkCtqtxlsVUf20rWwDW8+pt7AtHekExxAgr7oP3s4S9NKWpQuRWNGF
axinVeeZgdtfQCwfRgoEUkLzHyvFyIrsIgxobPfLmgZSrEkemW0jUULqYI+Hb0vb
tE6F0syUjXbxDB8m0ZjCZVo6IOV7DydMYPFCqMzjQmRvaI946E7MNkPw6uETt/6/
sPyxacZOkKg4E2IXl17xVAYwdyKt/qIosemKyvkV1GbMeTgnBkaWNNbr6iCqLI11
9By+uzBQSyQ3M9Gkx+7FRafSAjW4zSxEfyKWyAndTV2uu0kKmhzSouagKR8KcYMj
u7aC3pBWWiZ+nqZO7znKkfoQIbaQD4k1W1bFwi921rajzW2yunnX2NwSSEysa568
WtHX6B5sZ1UcVQ5QO7FVedY69+j3CJ4EUfGwA0OiPzF67rV1FtYQ+cG8L904MWh5
+H7h4oqBXNnNB2tDTTtijO1XWEWvmv/Y7U9bQ+ag/+CW3wFaTWf3AMnKCv5yIeni
MZhkR0OGfWdw2QdwCNGumO2baJU4cWOghyPAP494P277jxtC1v3bhNItPJi/B/6I
ER3Qc2M5jL5nCYwOilFVpd+ruPpA3r/d30PvcElz9vZ7L5y5HQjGPOBMJo1xdcnm
EWC27PXVHUVwfFr72JDOafVefcpYoqoohBd0WG39ApNlWGyZ+htXErPydCvm2gy6
97Z6+L/AEfEjwvbO+vWl+UbRQ6437THQEwoEzLUlzbkeT+N+kEM6dITmHzgZsq40
SJz2iOPoNGAbgC/GznSqJ7xrXE+habzfL5dtxusOEcRysTyB/9ThDDyz9ESDxtEN
3tiWsvJBglU1LbV7qgEvtUMBh2tlBU5NDQegMgja1J1Ds0YXSk6bRl4N1jPSSWxI
S5lCNChx2+9NDCGGpogc3GobFeuXHzp/+7MDPf1DNtHLCwDzIsXGPlC5bWKSNKls
srvBzD7oii8EH+azW2O0HDz1P/gGVjRw9G4OI44U0lmgchTidVX+T1e4dWWC065o
gTKlAyKuVx8PTrQq+HFwrbaraZSUUak5nb6ksre+6vCHcwk4EbynMbd+O/8IjrRT
C2cyq6TZmZ2gdENlva0JKZAkOol5QEAm5InCLDscJsjjldX4A9XTZHUgx9hWe+Bg
jaBKOmw4+iGN+s/gXsDXfXA/9sV75PYd77lNU6FZQfdyfCdkIezcUbzuuAki7zGp
SjNzggWjPFeLpBjBz9EE17iQ5Dnj5t7RV9cjHJD2YFJqyC8A+eBidouHGEvRhDYR
hT7bRDEgOs3uppSwxCqCSvdiN7CNdmf4xprV4xtsJ4okYwatQDUXsIompC+unV6H
PUGjcFTWJ1qZeJgiczsaCknwFVDrAYDxYMSLo8U+nnklLjLx2WLzHrgOv7wh/MBZ
5XISKRIcS9SkN/NBHYFnULdd1gVyMmReyE+G7Gxf2iBIJF8Gm75L3A1iJ6VVebSW
TfCpTp7qqR2uSN+07A4/c1F0H6RrR30FDkYbmSbazxPevzXB2EkR1wXAsDy+8R9W
SBbEvZA2KV1gmYf8PWLGho+m9yNVy97OP6kMcn0jDfugHv3XFIPav2vw2wXtCUQW
SJVuXxsi9cv1x+1AdIcd1MV8bmkJTHxFxVfjja9jmd/rHegrxG5xntnhKk72cEqq
F7Juta00uKeN6lIu1NFGBjN5Q8sEGUwEE52Oua5iR+YBDWWVjUIUx2RpbQ9DYsuH
cQooEaOL/W3GzSddUWGj5pbj/jYOb0WAUIdG+e2Hb0RQrgzqNaQCwHGTcmChXKNu
Ekq0WEHwlcZnviB1EmixTGz4FZs0csqdyDsyw4JU6eviL8iuV38NxhhqiX08YwUw
X7fTny7/el1YtrsaKzxBivYhXNlrp6WrlE2i7lfriKkpJhBin7ygASojK5oAqb5v
QcWNKb89YIdq0YG7hkE6BO8gN7fyz+w/qQ2/BlVfypOpEizRNcNjuKBEgLBGwQ/i
6UZGWmC2HZkWxkfGCQDKpwrS/70TCK8/T8obmYTDAJlJ3MrJenDiXi9bS8b4BCra
hHkOToNyS8v0pvP+Mie68oDeUnq4TMEeEmgbXnTZuSApsHWK20NnnUaHDTA6EgQg
/mXzTWKBTP9dL4AArfc9zP+Nyrd7p69PoBfIm0hYA0K4S2i+WvP7JK0PwUmyt6B8
ia7Ay9lblGJurnBxXkZVmWg0c7S/95sCUyr6lYfwWpSrdc42flv1IU9/TiOFERB7
ajpEBBGG8JyGy5nabUevLFm90hv60b/B4TPfaqU91Hi8Cb3wVIX/1OLi/eMp4EI9
akpXDc5a3bWUnHD4fcIG4elO7QgynNs9cMQUSN0j52JWFxbMsRvv8Ec7f3c7AhU+
1CnQMCWE07njpmThuMSiqGHQlMR6VwDbxy8KEpai/kfppjTlgD5SZuE2tkKywEaX
PB8h+oSM3jpV1HCi4iArcL5lxOt4Qt4ZHAsclEW6wPHxAdw0Gbe7bQAFPpqgdavp
BzBBlWstB4/U8UFK9u9anmnX9T3bgJRBheFVF3REW9RO/zK6hJvpzW1Ng5F8TFmv
Qz3RtKozMObmhbJDU+Gu6//qNyJYIhKoPTQm6ZY7SXBJC/xRItg4MxYsEs7Pl6iM
AdYtxidagmsTUqZ7gQes7HQG58Yi78bGBncz5LeTOGqWThXPt9sqbB1P1CoEVU8W
wSwZO9aVQWZPh9q6r+ILYDlpzjMltSnGJ5O8oCu9Z9LA58KXYuEpxNrQEJO1+GrU
54WI/Mz2OO4kGI/NcNbYbrq/clbANW9YzfYGPvcE/ihmY7WqKAx8rECN4K+AxIk/
vGL89GOTpG1SEoy5xAzDapT4PtwiO0zwvsAxrl7G+GBr/W074aLcudqq+OyStjMW
FMNtVOqdbWfyXWQFJL9+16ev7+U6XVaGbfJzGNyoqnXpZEdgSKe1HPNBQMPeEDRh
sUTB16fIoEESzCvf4ytkPPRpGhrqrlPwtRnqu3nSaPBr1Guw27DwJbgPLIoz+Vc2
8Um3GS2ktgClrTRVaSlIXMxA8tt3HO/nz7y6yjiLtSxuMoTQt51RjHGEVHgu1XcR
arxiTki0Q0TB/kuM7Cblcaq7kW1XWreq2CWY0Eh8cPnASokc5cGEfE/KxbghrwUw
3sdxYR7Gr6SUGdSh14S5E5Oez+AIWacZKrR9E7C7GwY7Ka/UWxP96iy/uvJztd8A
rL06Yc9k6Y0LZGiY7wEToBjdF9YpNK7p+ztOC8GnOB2J/+HzAr4vDzDl3MCgZVAc
DNp69xYdcszPa/kEmo0o1jpa3TVnkvPGLn9N5YE6jjFoNQVou7bIY6HiZXmUovsq
nSL8GIdEJWSz/ICYdh+dBP6uBwNH6izOo6bB6DDOiDTMQKnolP6eXIA131BpF0L2
eSJ/ARtHGXTaAV8EeuuqAA/gVi6GovVBpyIID8KuF/NtDtP0gP8tfqjeVFvF+xJ5
BOqX/7EZ+N9lXTEC8ySG1pRnuxy2qrglPSf2kkN0AbLQFi9sNuXqCMJQEnmTR8eb
U8q9MzYvf12DjEnGIN1p+YOR6qnLN41f9moU5Bstj9ARyXCRbPXsO6bn/BDcEQxP
b1rwg+lafrTffsJ5xOOt5BaYz+Ob+zT3dd5wBv12HS5Qln5wdhL434JjeyZbvIzK
JniEpXLCyNkE7TvFkvOgn3v/obx1vRXhe+TU2nU4/zK2AbScnvCSSceNY/u0+tPh
sVmfjkE2YQZanajT224FUDnpKoME7tZXNfzmH3G4X2TQeKYIXHshVNVXLB9bm29e
Jc/AVcfERseP8LmXDw4qagxxO6ihTW8u7zYqPtAajrW5UkQ6RVNeLUxJmt3AQW8i
qiEw4/ipiq25fsFYKuA3Dh2Me57Xq5yAij6i1BgclZnXjTYIFlqU35+4Rsxwtegz
qiH08qc1JzfO6+9VFc7Vq8dFraM3dQVDIyIxeKr9AOi1ZkOGn4iipzFmDMajTHTB
C/w7LX5NGGh2w4Iq8B9kNZdQOMebEs84aKFWImW0tPb6sRe95ivYgNXcam+iyp0j
47wRHt8fa7AcdHJrlBEdugcWdJbw10QXONXJGI1VOlsqoOg/tK12V+7hfYhQmxNT
KgkvCV1itojg8zglKH1qu5Xh2Ltp7SJk8h/HpQDsu4dtntXQcKNcSd25RgbIxJaP
PvTCBvUGe25fF1GjB5uLKtf/WIPToMkbGsVerLImsT6KqhobdBWO7QJYoQ6tU/pd
kw37WREEgqYUg11pLEWEeT0geCN1IivaWxrWdLUvZN0uoMaGybD3XHY8I877S28c
CmY8OuKyBW9L1oKCx59okFA2XewM2hW3G+A9u+59yqpfhj3NQwAGaN1ZWEjYBDXq
IYG5Jun+DL7AP44M+37LrO7HpcltEROsvdACiNKYiFBmbGCYzTo4+rTIEQPIwfOP
n3SmcDDy+9IBYy0vAK3/Wr1QXJSlTHZD+bzBiYbrfZMEhuBYKZaRTaykZYfZUS7n
VLCtUOWSdzKqL8JkK2pkC5IyZurabAehDF+qRqXBVm+NKM9GYdInh9vtZzsebdEl
FNn5N2EXWY8Lcd4gSwfa44IlZLb9uGDhB9bAKgZvBLEV89oiOkcAi7jSI3uVpzbS
uzjCaCjqJTWLJ45ODZNVUTSutagDPtw2uaN0ff0+7A0q25l+qMXIQVxYMeCqWskR
niFcjL6Kb/W37SSlc/wrqKMbQ9CyzoQvfNIPmn1cuM1VtUfu0o62XR2ipIjyLRQL
ivq3SdxLYU/aA9l+RVRiUGlcq7piCTY6nLPjxx3Icxt8Fz7PtIruaerIiwsn9LQT
cHN/nYQpTgk51ZPwT4N3VBmJ4cjv9yhfozRTEGQiMSISDRymesKO2diDgrkcsYXK
b/ohd9P0LdBTAmK2ams43njA5vXnftweqVMbbxN78odDf3Bw6WNWn/U3rNtRvucv
ykMEd2Kv7mFCfJlwt9Lbt2PEeYrDQzASzwANNJbp7t97NR8+UV096IMJzjdcc3nX
EjFXOXjf+NyowCkiEdUzwj0N32+kMHud7xJ3BZciCtjUGpspy9WfEuMS25XNmtJw
/ZcUkQ6VDxBPufUxo6PTuP5JzCzxBEgKUxXUrwws8zsN9/3CtWWaQGuyKPJ+cWUU
izmV2Zcjix/sKm20EN24nNVePHwvir+8gstYrbpt+mibkdcDE2i9uyWGsnqJHZR+
8BMNuz21Zy/aWUDBDOkYLg9VtWrDQn0sJJgqdqM0FwD8R5m2GJ7kJFafy7/Cu1ts
LpKe8ev1NwPFLgbTjKZAC3P93vl94wQlHdn+78K/W0tU0cLlmHREav3BWSfd8gCM
cT8Fp6BrAchOqa9GmWhaazw3bbY975AaKCwRE/mHheOwMTxWxFfzso4mn+dUDuOQ
LJXjwQF8//PwKbKahtgs4C/xmQjPnYJhbS2UCePIuu1/BEsICG1kCv29tgGoKcqp
+pEMqxf3ZL+PqSti756mRAkdcPq67EeNVsSda+ja7Q4ksU7T7zw67enmyb9pm/zd
fIiPVvojusVhUZmP46QM8vHF2VmqBdNKzsRaXpG1pUUwgC+SxZIXhrpgxp8E7jeZ
+TWVC81dDjy8TVBC+zqIRgaxzd1N0L7YUCBE7WmzElgHlIlP690IcKMmjCDLKOLM
MLQzCjfn+hPyrCEI5q5vJEU4mvQA/1nTBaaCkzyaYJjKnvRe/8jb+rSVXk40K2oV
sm/DWmm4cvh4FPn1O+PBGXYlwJ6a//b0mPA3iSDgJs7ptoUZewCidYNNrt88xL65
rWAaKeOtvwrVaspNUdJge2ACGgZJPAo3KiX6HspZKq0CtoUshjjIMtOmsTr71gPs
x7cbOQ+jx+0QFZU+3a7s/FCpxj4JQylNMumRGe7pPlHFgY95ckyhg2IlB7/omgXe
7VeSyOhof0MxT8LdmglMnjPfPmOrGzM0mN5Wpp+1aok1bBBEI3OKpMyUoCZrTHzy
PWwtG5krphmLiMfYdhtj33enyFe4iDaRte1L8MBnISLPD/zwsCWN47QoEoMExAxO
E3l4qPDQtIJgbVNCXztDGOyW+N1T1ePfNIHW7hy5ZGMpFjQqVKgql4CkgP15z2kd
i+1WZ1fM1WhLxQajVgHX3QELIn/rh2j6wEOCWc68jW/Q6ME7CcTuunLb0TuMCHgE
epg4MNxcvl3hs73FftSCTF2KG0F43Qg0WZInT8IJGnXZkMBI6QjSeE4aTLOOT2aT
nFRaysh0+vx7eYumoWq/rHVAT+VK8lm2ApP93V0o3A3LAfgl62yruKLNE84vud+n
BuDciVq5r2ujIaRpIf/1Z5vWKIxhczABIQXkrEAv0gQxKOHnLJ2tFSpFezqX53VE
ek4PlfF2gDui1lyv0FTIwGznMje2ZurIqKWtRQ/ibvXqAl3GbHS674ylJV8WZGXl
VkqbbMaqRUJrYJssCunnvHodOGDhYsIynnjaPLWPSNO/0JGnokBtwHPjstPjHGm9
Bi5yxBHv8tCXFSILtDcHCBCCtxbr79zrmzITrPv6zPi0p40MY7RHsh2bTgLsyD40
ABOfkO2zbsa6jIC+eTGJlFG8iN0/4seJnmbdezvIvBW45itZQVpN9FStRAzrb0xa
TV4bXEEuEHm0bQ1UmGGcyXJpzzCjhWzqgHOfCYk73+jdtnuhRA+ypMiUwOn4IAqL
PWRdEJCXu9cN9dHkMfCx9YNuDUVs9A/1U0rJbqPaW3QrPI2JiPys0CskLNK4BjLZ
fdyeG3olHRmlBuU5saZIKedYy4kj2ZK6hS2dvPVjofIqXPF8YuqXcG9YU/y0CZZz
BCefxMN6m50sNa2tGP/lG0QPvupFUM1t0py8JbDuqK/c/cpF/Puy9669QxT3+4b6
IidKmfR6v6WxgAdAXeM1s986IUHrqgUNMPF08UremryjEwA22tKvxY0HfXK4DfT7
SqPITCPFb8CGxEJTBbIDDK9Sh1/Oz3hoa6kGPQnY1Cudax22HXhAfeHWS0Ch2R4f
gKLFzzUwK5NoiXNQZ0wycGAA6nqzObaVqkNfrwBcjCGcJu7421sO9FUu9K3vP+sj
kbsPFLH0bvkoZiArEctw93hKMbGJRYqdGIVLJnDogFXTHeTWNVFGf/7zG8Apg4+9
XJwaPrS1J5U5tLKSQ+zj+v5/T19SjaD3WT1bEuA8ib6UD5SkBCRaUrhj4LmAfoxx
pZPW9VlWeA9mCTOcpbDmDBzCY8M66L3d9377o3uCR7Yk2Jd0H5m6lGvbMPDKO3Rl
pxuR5Zkbvx1Xztd1/SfoSQN5sRkOCmXi7P+YzJkw90UD+b7vTEH33eRfyWadgUNa
l/6lKqfDijRdElLZyhypXn0V+MLc603PBuBwTnua3nEYGBnEP4gpUax/ytXQ83Ad
KyZ8if0CUvUX8diRWPBR40z4llYn2gfldIR3QLQVnEgYVumh2t+dmesXvbwE+k56
Ml8WgieREoiTvSo6RuXO2Z1hFD7dhBwGGastPgwhxO0OpZMuzLxvdqy10l9/1zhg
56kcdT1IwnofHW/+OscZso32XFRDT15VLapNtylI4rOyW++45idsgllRrNb+P1p1
WpYUH3hwbwEu1Y2HLv4nruJ57tci310TPZw8+DgXFlxi0G8PwEy+uR2SWh1gzQo9
00NA00FkL2fVD/yShAmnoydIzd10kHon9UUpueH/ON5QrNXfqMLdAW5cE2JHmIb8
580m7HqjZPB9+mxMYbC4rx+HjJCkbMxMsVz8stYZ2OkpzNb4cY28x5hUSa60SHct
01lTcauJTLv+meiY1W1/fGAl//stw2xlmEgo32yFH5Yptj9mFb73p8QtPCuMSnlz
6vAePNevMvIz7ylBxnNvhDg0m9CrigAho+8soDL7r7uQlTa9PhEENLm7gHHl2LU9
MYP46QYZa4qdCLTyX1bL0rce2N+ncDMy6a9DVm/JpuZ8SiHxXm3WbPz5QWeckznO
0r0MPFNnOc/N2GcWTvcGmvQz2DMm8c1Z34spArOTSU3Nf1Sybpjg/gUzo20AQvgd
ntLiEkVK41d8Q9JZNu/Y9F7Roq/RXKc6BY1QuNaXOtseVrUJbQ1nBMPOsrmLRTAK
YzTOgXEOrWXOwt041bwGrdwL/3vpLbFwGJ2iA+moKFzDKhTo53D48c2URSDB4a8R
al7vltS9nIcMiwet8Svq7GXspBsh6i3KRd+mkouycIyxh6eEiduC/iKv01luV8QX
1XW5cccICPuw+xGJAvbMaJKZnzVDeuUBVDxKCgh13T7ShM22vq4NRKIsUYxsKojZ
oKGUx6QMOviKUFC3yQn0TfljrX59zwjJG6n0QkAsjhAghpPm83EsJtD71MlF+nJG
SemcWv7hr95NgW6XFEdCfpRxo9vbJuClTDB6S6uipe1BSvP6+C+VQ0Itw99q4VDc
tUG14pUFS8mP+flUbaat4v68kPAbD6CYag4zKvYi5Uaz0QXXyahoj6fXc2m5ydYI
KcMewGc2PCe4EY8NxvKQa+9CwClk9LwZRXBG44VxzgKLd5AU3Xq1IoytlTij/ENZ
o+2M2f1P2jgvU4UwtfBdKG5eSIg76NAq2Ooi4UTCptwh5dKIHNtCdsVlSzngZS6/
LxCrNrhSkkkuFlt6ZGyvuybgbN1tVl0SZo4FmVBeXpQ3aFBIDgnpXlIW8tdaZ0sF
gjYH8+loNmg6W3uF0xSsT73JPF/TXUOqOV9FiyHKO4Ea/hRJubQ+SFqfQPoU+1lh
bq47aMD9C1XzJyMiTDLDJWM5U8uoScVAUwbHqK7CgmpKu3D8V82EkvNShb7ICZix
c+KDrmOnxuNFLb6SsWNrJunFemhhY6rRE+WHYmMY7YJQaDqp2c0NnoX9KuD0l+Ow
cgYEguxPcu17aItxTG0ehpsGEaxFLPHv2Q5n8xSx4m8CprSlQ+aV6L9tTAUiHw4O
zK6tb6yd+Jh3eymTqQCrfTWqMQcenY/Wl0bAzqW5ytYzoknk1G247emWEZTwIrir
op00b86+gxSo0NejeH5Rhh3Nyqy9+duIag9HJ+4/oB7cCbkwtfA5p9EE/clzGrGi
ocee/j4CBb36VGZqSnaTIPXDBNyXfCNRiL2tGlztclSCNi1OUNwEgJSUGTisThEh
2VmEPUnx4B/Kn67t2bga1OuoOU3fy/qB4FIacdSTN1zWS5FPhqCeDaypzyMhfSrc
T8gwPZpgrHoLgYkw1uOmxGOJ61hKLrmtyABvE3Bb3yWBXCKegM8I5xx1ZaULC840
9YpVsoRRKIaG14Vh4S6Itff6aNQeJK1aXNLERWveQ+6TvgWDSWDqWhiko6FW9G2T
YouK+BCzcNcLxnOz/HDzw+ifvgxRJ1xJgJuFeSyDaKirzPCteLQrLRUv/T6fR3BA
HYhwTqcBxIi5LvQAmM1pbmAE9WQrVcnIKnXmJ7h7gzljYLPCrG+r32bFTE2S+fCI
6cwjrzcb1gbcD6Bt9j8+MENvOn60iEkK3CW4HxVWWSQhdV6tgEF04bByAtPGuGO+
FLfjwawHccicP4Oa+CIl5QI3WbSxIlC1IxPmRgd2DI7pDd2O/uBg1itgRYcPa7wN
OQ0A4JRh4iCTZJSqpt3TXVANkbNocWlchnQKVe6ggD7vyO10t5JPgYiUy0NqhdMt
cALNLUpQAcHighYZxjeODY7wz4AY09UJ7x+gAEqq2eIN28582ExEYnliCcD/FUOf
0K+UWNzNJTUA8yhl4o6OkoEKVIn+na07+wmybFQTRUWqszrJKKdsx+MFkqo6bjJE
Ebo9IMTaE2T0dU64NL4iy6De3C2agUU02fn0bGgnP7hbZNAabgvIjD/4FWMhMmkn
IssWxJhYsZOjm3bA5rqjqGKnL1i4tU2orXPdM4e/mODSpoj2tsoIbSx/iNDPSLKL
CW+rVVzGotD5CYJIYug4sZpVd5MnnOo31W07DJ8CpcSiiB1f1I711g7XeGuHNSFR
1QXo3bvugUvi1dfXDzWWgD6AfiQKpqVWx7EysEcMQYRvyI8j90F4mi0YQ1VXg1hx
ew728dZDQsYuxMdWGc1vWBPJsE00Fjo2oI5Lt1cItlN84K5n5Xz9nMGec1Nmi3G3
XioJySLf7rkrUWVJOGUdjWU/oVue9wuU+ZAcvyJRSQ2Pgcnd7L9L1Z+8jwwx7/jC
fSbdh7EVj6ffUPM1V0w9IOu+YRVYAp9ggd3At7W1e2Yo5CzEACx0TeySOLeG+345
UPLOvTzLwOyt/SFbyXRNJCFUAhb6rWMC1AewBgjWq9hsk5arR0ayS0quprBQ4yO0
JWV+BYe8bkAswF9rPQ1s89n+nEsUWDchfKv8z6FpseDNbq2up0GMbfBFtwAYCXyE
MPzIDrrmCmOa1gbEBOjCSKCDbciGXlKx3yprx4My+F1+K0kvdNIZyO+Iesl/RUE3
7fgrhjGxQUhrbScsRs3nvzZrt2XvvXbZnWF36u+8M8wMwYX9WcHMKLTps6itArMe
YuWHZ5DoTjaOSmcocupKufks9ljZJJaWv9QYpWMCLNpubPrPwjC9uKa071/lzJmp
rGnp3nT7urFLtbZFXUF0gCtTQB/07TczK05qSq0L4B5GNLMSKzzR1SyUFMqCkPKP
Dz0NX15m29qDch102CuxrwOqnCqoN8dD1DG9rAOLhchcotBtXFP9jMJe5ZE+LJw8
MFb7UBKl+Eg/Dp87jjrpBaq8rWZ2TgVhnBd4P7lBuh/tgIzg3P0acu3Dm1OkgR5p
BJXZmB8nTRsWO71xsVJTnU+TBWamsX2CsIXqUfl17eWuUP/9sjdvHEyXyrq5DA8e
4222IQGXV5ZhrDMj4MRQQSJUpIZXQkkgTak76Jbp8lssvz41GgnmSxARVRHC+2vI
ypcRStPdM3wvtkE9cagp+wPWzkwXA0GGFVrR2Fc7vjnvi+YT/+kBvpRxk9c9vk1k
novFAxR4FMIT8Vtj+1uf8lJBAjnj19U2AO5etSU6qriDBJmystGURyAapOg/Eium
K1mtdj0dTw0noSjYsqQv3tQi3JZAjcuqzm91CZUcyCb2/Rnq2QqaZZfrOjuC4HHM
vK0VVRw1+xDi92JVbgMdCEPjgBKsNVgF9dGO4wy8HpBt40UrLc6gjj700Ey+jMLk
boXoQ8fyKXjA2g3FozQHvAF9x+Ex8lCWH20oLCF3xKcWQJrIJnigEDSqwnCRgz1X
Z5hBJYECdSOp7W+o4lIq/4nHb1JsdAFUUBYdFc9cKxGdPiNYMUX2/CrZW1wFo2gw
SEQyv3BkZFP9QgNk3jKYUD7jpt80HQvqwTyM8QpKwPbPPjlR9dmuiLKzBUsouod2
VvgiDUwWtAIXjq6CjL2HVn2O7ZQ6YVY2gE8ncI12vTWNyRf4/pZ9jwpguFLXdlxU
B4qS5exj2zk4QgFe/6zhK32oniXwgSoys7RsICK1MoweDHpOsHu6iY6UnzLeU5RH
Ed6i5n8/iI/xioE2q/x9ENb8ehkJBp9N5wZUnnkYrOBrgHWw1Cgx+30O1tKwBTDV
Ri+EC7p1gnyAdzbEwZAF5JrD/eSgyVAjJOewsYRSdbFVt6T0Fqdhjaghg/cdzWDR
zYyId4Aog5up17kTxjzbrZ6hLPeY2TMezCpGjaTLOZBSH9kPMGp0K9dqztTAlGk3
xxrSQecogqhy8irx3VaHM9m+aHZN3DBYyh7/GUHnqBJAiQAG9PEuNEIv7bxIPW3j
Y0nHzrKCOMcDGFJdRPmfOJyBaz2jrmpskNcbkihEg0yHpJ1b1cSxjamU8hMfsg1O
7S96apF6dh5Xz8Xc1ULYQTQbvRdDczib+LBuNhs0OUNv9XmvT9KeErVgKTNA+I/6
TMjeVw3qOVng1qnrcBgP7klUNY+/K6PDFiHzExmyTGdbdP3GbVOKcGGl4wRnmsCy
YBHfdogCIJ++Iw6Vi6zfNYYO47zdL5UhRrHJauUzA0mlgUcbMWge5c/75Ony3dB4
0PiX3f/nFHMVn9yw/3feZBZ9nfbpB/2CB10ndain+rkiDieffWJTozT6dX0NT1rw
Vk9G/Bf+ovGLZSKNI8Yg9R9x3h3jo+aZJ+zapKmsoGKrZKdWzbEZ0IYJgqACjSyv
91DTbtInsBYrCpg3Q1Jv7PJHzFkd4vkL4Anbd3YZHy9k53OWwcAEmT9dv50h3bfc
YRhnP5Ub3vNDYRqWxKHpLiEx6bnwu5YWnJCk7M6x6n4fcni9GVrmvqxumPDXUC/e
6c39DzyrbCvNBFupUntsEBkTCwY04D48HtmAuPNH6S1hYz1ufrSy+R49ssNEx8Ds
0FY1+36r7uDQgyA1HORIh2ItN3P/92OnsTqGr0fR/JnJmosO6bBXyMROYTpEMDNZ
k+3XiGp+2kbHombuQkAdF5TmDdL+TB78gK3HPgPx5zF7Kr81uocQQ805oeNNd58g
hzLTCBmk1kJ2N7ArC9jKnhobaIWgcuwwo0XunOuqY04Rt3OWeoX5NhAwBF9HA39m
HBnpKNMxnUWvQP0HC2VVH+3URWhvCAJIJwKbqeLQz99IC+fH6+OwqF0HIO29r1mT
M3g3fWJIuELjt06K7JbhlZDxTH6qrax1KNCzSvo3o81s/27EpUV0z9qCsP4ZvX4E
0kFb0VOSQINgPB/HPuSo9HbRpkIUCugJAYaQC8a/CxVGe+Fhz4ougX8VjRRaiY+U
mLypACth85h0O2mvpBTQbyQ21ePKBNnj+gXYxfTFvy2tDwo9uUx/kU6OgVCCNow1
YSmUazsx1TO7CLEW7gVCfTsrBepEE2G8t+7KAi/q2rINTF1AFirBoqN65qkmltt2
j6UdaCDTb2mOM4e6F2P+hVieIwU3/H8FQ60SGSBkiJYI6yAGdE67Yn0igQaCBm8K
doa40DfNqy8UazcGYqT6brkBZycHXymx97BS5AHCPi0CJtv4HqmgvLtVX+HaMQm3
HOtP3ICpb8GzB66IY6KvBMpfHVoepGpp/RekQXKRJ6Os9ZHVBQcT8xGd2urMnh/9
BRNyERvN8mPOjWk6BVSEixuydF+WC/HyzKizd8/cnxGTxdAn8rGHrIHetJWT7yhR
GPyVL4fEsEH7AZJEVESyMO0fVhoKMNswbWBg4TIKGMh7J8GLvJ8sPZLx5ImQvrd+
eRU3hygBj3dfAGBe26AhzCct1BY5GsV+cBtiXbCOILz5EJuBJP2APJt5biVmRoAl
4ZHYecQ6jrOkSA4aFx8S9Qq6Upof0ADMjYuulq2H5BT+ycYyidtNKecHBATSJ7j5
R3l5BkJA5/6tX7IwzYICI8MSxf6y8n+swjl1zxOVSnVLjV+27FyzFkg+zr7UxmuQ
gWk5/fxvkApOS6MzwAKZWzWqWy45vG5QYQNnxQu+C7qwxEiY9wH91MVpmdpU+Pdz
QVTCvSOpn6TJLxSIhOdAz0BgxzBgVzKWGkXGQVcjjzrNNKSWU/AYPe71dgHLyO0C
XX1IDxeoPI13LTg9A27E9GAP6O+Z9sIWXx8oI3/M+1JmJAhTsZuXCrBDi7h/TCVT
rUsuDMFCBcXI3ENKZhzQLtwU+1lPydfBnAuLh0wsjONX8Ymq3B5xlF1yogakRAnm
ULtVaWc5DOLnyeg1bdF6KNBFb5cP4zH8U1CYsX6hTVo4MS5l2lCVYMgxFvxAkY4I
S6qEvfMrS5jeGZDLmBJMO8Qb0FYNIBksvBEAxdRzlgbiQWKqPK+Zq+KGtNBkEei3
vacgQL87W2T7YZG3UmAUY1djLQp3LBkZgXmS3WZ7vzj7klh3AnmWx9bmBIIOHaYy
RKxoHNiZYwuRQQbwk1e4uxc7cEHXd6v7wD+o60MS7nHvJMVzWIuv7qgEL+xFpXOD
0j7WcJr6pLSrC/0ejXZ644lMQTInnrQTnylsXN4z9T3zdb3LbY8WCZE0CiBMokRh
3epKj0Krq4ANUuQuYUpOmG7y+n/iCKaU2uunbp+nCJ3582oUPHvF5vf2X4xTEB2t
fsR2zPKksSPo6DMmAVVEe3Lb1kLP1xBZPI+VXuDN/Kz0X7aTTYEcL9zVY/pzjXFq
l4vM0qQpmiQfjPhgpnCYEs0M+PePu9w3zmBY4G0kznpi02GUHJg47NuJinN14loj
I4tIKC3w6D3jqfyBf42uJJSU1/8Hd9zUGiZ07DWD/ELl+K9T0XU8KTcHPfXp5sfF
KzOaP1hBgSnJkKxarUhiMSoleKXDTpsd8yfJCEM/MfOgck7/nhoIK/sqAwYmVf2p
QMTRa4RNq2GhN7va/rEsBSxIDpK7kyC2QgrywG+I69+PwM1Z1A1WpnxoF78ezqvP
h2XjU88+vLyN/7E250m4NZtr8p2zRjtYAXVz9ZCIYhItpaXKjsvqlpm6elA1SjzA
m7tMgqEyMluswzjyTorVzpN6E4aB3FXQCn8OYMjl+/QsHgHy1hXOUyVbAveIitJm
IFptCzqddr4Op6ksTybjQypgn3FZxszQBkyQWZA3T8VDIt78U9LyGrTlrPsKjoR2
7OJVTs6qZHU8/2HFrqmA8gXskHULbvDhv3y9LVsu71bapIdNXJbOJGPcAEurlRVe
zrJzHu2BDvu0HouCFsvp6gD7Wk9zXrkGgpJNT7jda1spk2kgMI8Udea30l5/8i2R
v6boUiX+LBJYikDLn2HDdN3qnqxCvOeC7jdMdXgsNZLBys1V60LzvWspFr7kfsp9
u6kPoM9NPvXw3jBC71S8bOoXmTD5OfyRjTKbEFq7TneLAMHY20PkM7aeB4jAXKTS
B6Gi+3I+eY2L9WtkZNY/lbJvvvEHW0ohn12zNRyq8CPcK8KCtGPcFYOKX7kl/C/D
qxct5g12pibjHlV4b+ZJl0avuNeLJ+ycmX7+sXyVuPcnLcpsR9jpvIbahlUqXSkQ
6qBTMeJEFih1FqkAC/zNgcEcIwvsZBvM7f7R5msT8r1cVOeQQr+nVvz5IUnjQQgQ
UuErvuWMp4HP9JkegDNGjZ+Fn1TpdwpVywImp1OfVG1MF+cFmUVVNIUJ3aqZhfEc
ttRdCGOlvuN+7qKhSbWMwfhMAYnhxhsnNyQt1CLHELuN0muAKNfU0fLJTUvxZMis
/+ougtIw5jLq7O0OyvyUI9IwJhsESBWYu6y1NxHJXWXv/vbUqLJ3E2a/jEzGmM/W
JXnqr1UFiWAoe2PrmTm1+mkxeUwHqYduLYeNKcoTP059bhcX57J2V7VqlNJFXvVq
1S8nGbPMkQiA/ITwucZ5bW760xLuPUim5o3Cdq1+CdsvTNuTnHCMdSe6c0+KHXUd
dZDR/9wlCl5jvMpvPA+/Xt/+KyRemjQq4UO4qwU7IVpAA5Q/RHBSnvjBeuQa1P7f
ERaGSuGnfEFm4XqXAwLdXqj0Ub5qyFJww++d4eM5Y1rk/XsOtBRjDw6DDSe30tTO
t4P0yTfGYWAR74meznNWjt3oFHOCQgSbFqBHF3sqQM63yB9F9motPSZ6zqokQqwq
x6FT7vBtECGn+/NaU1C/n0Kmnu3l2SjOe5NdBmoxAJRMcaLmBTXy8ODq2slh2PIt
680zjm7q5FSgHQ//d82c6C6v/vWXwkAFA4KiDjsUOnXMjOKgHkHxl5H7VChBdl1R
FQ7bDZuQqV5pZMQpaNqfvbXa8gdZa9V27K02P6r2Pjj8ri3NQHdr+EHdTTJdpVgt
FhPEseLbRgwz1idLT1QKQ899aMCXkXZp+kBjQEBhJQU7hZ6Nxd7XDSIYTkprGS61
IVnDyPi8oQLrYgkNwKK1lbGYEOnuwepYyf6uA+TQrD4MMFD0QqXdbrgGeS5GbP6K
EuNOVtyMC3hi7YGV8daWzljXDYGmNERlJlVTQ1SCjdYPeWM3bm9WVV06BBycRCR+
EKOTZKHALEJK6NoDhdAHPfOPqQMPXU9E4jkBcRD751a5HlL+KZvpH2zOxHNJMX7/
OgCsydgOUhPllMEzUThFVYN7nhzMm0FLY2qTZCLd+0is0kWfYa6Mqv77jvWwx+K0
bj7NNJVo5izJfsn8jPDobJ9csNSSoG2MND7ub0bslDQivVavCnN8eoTDojmRgNZA
t16PZISxDXOYKbER1anJi75yrK0EErsq+iaRih1IjVYjFUQqX5MO3aRAan5V6d5S
VivHPbhJbYbvaoigygkkgzte8UWMbSueFdb5GA3ztORhLDnBUs6obAEVP4RWRXfw
RVbJknJR/H6RuPsf20HRbwZemy4jVyhcwiHPMTdJ5hoW8NqcSN3VqdMCh284jIGi
QYW5ffbmpfVqiiR22rzxDxcAQEmWZV8NIryHZCaqlNJgDzO2/xIjVNiUNbUr4LZX
D0/koGr5OaeaLuP0q4CEs2Qxcsyf0TzTL5wHT5IgeiXEbi7FPI/M1c4S1qX9et2p
gjWhcZkOpnrWV/v29rEdBR0nrD+s3xM9tC15vMBj/LNsFGi3X79RJRkWfSduQY/H
7kscgbmwJ6RhlS7y0wWI6MkKZTWLbKNiyktsHb15Ih66tQLzW0mlqkGcWZ82bgtF
HF2g7RBqE7VzGJlaB+ASUUGjU9fFAtFHQjNmim/BVrT6ryfi1vtGh7lQbTZ/mZTo
/10BDMZTz6vmUsP3IkGwOMs2P7+ZIcnGjWERXqAmsN6eTVCINbq0d+p+7TQ38nqk
Vx/du4nSslME1m3dyJL4L8RpENBFjqQFVmjQ5OnBgtqhqM3VXsbJVqMhj7pj7QK2
kq92QNqLBFPOpeP6w4OqtZNIRfEO8dte0EO/ogssYuHqotdSzLVy6iSLHXBXqRHA
9OOP0DHfdwAoEjkw+Q8isXvioe7/oXibC7vFtwtK6QR+N2yXZENF6T7FF1L8+ilD
Qjb1im1/ehnOw0UomALrlk5SCrXyDKUrURpMYq7xgwdv+hpCYq58/STESEoWj1iX
qx9rK36uLK+SDyncFBALBMJU+pnvgCCh3PtwFLZfmWCmPexkAo7Z7Q5qugOG6qtV
yP8KyZ95MwF7+Qoh0nUu8JYbEHzmUfwSQksk9ovwBUUFvDrq/Z1Eyd2e8cy0Vwv4
83ZMuczQeynvxGapoCvNYQAJekiOtQHYRgcoucym8//QviCYpL2/uecOsmR+KHya
io9+eXF3SlKj4Lg3gfzhFj+PlF4PXLjEjmH8Ihgh93hQV3baGGi0VS8eGhzUdHQf
AxIimEZhZTllmxBpu3wYXOJFlskfA1Mwvc+QNASZv8tGZbtTPMv2bssBRqGd4L6h
SG9LGrTjtJD9XTf5je9EdYlPWS33/PQq7qedJZ281Lh+Uq40ZquHViMzgvp4F6H1
A31R90tAd66eDp4Ifr1hK1d54x3SXnW1PsazeyPQcJDd1o3x5AEqVbGIB2ypPusJ
GHNwR/mPesxV1zbmHDKv47Q2w4rQS3v2FUTf0+aqo7o5nHjuRvabQ0euDen4BU57
Qi24+HvWvhikAulaNfuz5Y+TwPdLA2xhYmLiqobsn8qeVFZXGJo2jHE+Me1IyJeS
Mt8RA7p2P2uyWTSPuiNO7nvlgYRF3fREjXIZbUDTzDhFUbXtIfwU9XX1ZKc7Jnjc
BvACTjhpUgvo8UaWcpRUzYCO+lXNcnSRveZiQgpV4+Y2rV80cY/8cUXUVAc2obZS
3i3ltOGdMGctVkVNLyIsOfgmudD4Q4gaafdlRSAJ/Og=
`protect END_PROTECTED
