`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SfNWlEpq981yGyoFDskWa20N4+jvdTPPRpRdaBqV6iAt+iQcdFAK8kFK+eBgVdYX
320MsByF0tgSlL4RAemhnJe1V7d3Ht2I2PafocwEl1a63CdSiQd6uUjvdNi4yppL
RudIAxMrhrP2igI3IqbEJedYHSLYKWe3Vyw/jTe3VxaPF0+ym1x8Jtlm/bM4zTc1
+4eA4IOET1lN4k3I3Xwq+Xdu8w5rNquX1cCJHCn1LpxP0vYmqGqR5W2TqNb+I4eo
J6bxLhvyBu496s/a4NEV49364B+bNyst/gvBI868EbEXTs8T1NAlgNPWHVDTxpWe
KFdhAvW61RjafTkOu6ZCU2FZvxr6lmLhc0MPsKGq1Pa/a2o5A3w1A23Rr9dujprq
pKhJ5hYiwhmZTiuCqX2e4MucHcwbHJIUbUECwwBrJ+khS3ULR+8WDJjKfV4Obtc9
Lx7jQ5nbwJN9ue95ow3qlhSnUTmQVob/TmSMtwM6eItAXZ00JNbMf+ykEGTQC6xP
xeU+0X5bpA0uxa3P2EYD99g1RrIwd3C88dpC4FPtGVTvrsUjE270KyKMzTwr5F/A
pzKbOX+DXPuKiBvYklDND7PX+tAWh1t6VCK4S3BkmaCK0L/EQIf4hApkps/4yBfx
/JAq4uh4t9Jt+S1S8pYcRWvBVjoAR9HUySWTJVbFCR2eK+zDf6ukbyFOgJXR/+9m
wWvOaZMNndAaW/h9CHVaqAlwTdccfyCzHfxGWct6GZE5V4k8KFNNP2F4WIKKvCiA
ce3ktDn+tmnb4zRNed+lKdc1UQ1AHeh9rHNxwcfkVrtPoyDFq7WAgb5Lct+x/ZZP
Wa5c3nTFzxYziC4u8oIA9RqxzYVZwkiTDGIsGrfXp2UU8JqKfh3Jb9gvBdJCG1vX
JZbI65r9XBfqLN9KzwHzsQITBD20lFzwz6tQy2kv1LotXHxv3XSFw6uGmwXAh4Id
EeZPa1gApEEYPt/EXY9eobopsoK1O/qcTkjYIG6AK0NKQBmJsKNZd9k2YY+Dq8YL
GcCD2pbjYFWgWXWhK5LH6asqCt/jdPmsMvjOlhLS7XKPe31NTh/MGzYerFtSUIHm
Ij56vlG2jVPKB3s8zWtAl2Rel6jXoeDDpm8N9wGSy2p9ZnOePIDr1oZ4Tp75urSS
xdzYlJxoXwAY0Mog/m/zPn3tiDEfofDm3rHonsPr8mUJNooAtHb/vd8I1g6/wi+M
CEHGDA9JvrTBIrEH9HkmSaWL3kgmNV7CPXTwLEkFWGF77myThoc2hx+1jEOYDcSl
M1/bpxcEOKiNGmsfj2nfSF6bjHIT/xmAt0x0+NJksYrklezge9p3Z50Zj56Syw3x
PAdQtKmEflLvys0fEJ0tui0JWbUd+OxsTA6uhbEbD8WpjeBSMSSXKDA7ZYxbLxqy
mayU6Wn5H6RE4BvCyEGje5hh3f9XUiXkGfYplkmc8AxMxGrm25Wl7/7iqJMxkvnB
8lfs1efJ9RB8Jz4ncc59S0oBbi9sk7SdJGO5CrF3wXLGfBmRZj/U/0LWnhGcX733
iGHLe2TGDHwhLrCe3t5uZ4pfm0QFvmhd9EM/tyHQ/HPXR+2e+BazQGsp3IWjeNe2
gxDDUxzfn/HCOIjQcjVOIiAtRyjZD5gzm9+7KR7+9d3/SqBGzQEdkBKwP2cefZV9
2qBx7ePmh5Hzm5XSPghd1VOiRr1NSrsV9N7Y8daYxFbuu0plYsZbuaWJy2p5H9Xx
KVLSPWEQtPbeJKFnCN6T2YfJJFMsjMmWSt+NoX47ntAuN4lc7MG9lcJXGW8Yu7EJ
w+gpcdq1T7dcWdmuQYT9MOBSA34HNp9iVm9SqxNIn/zI3Y7LmHfpwF/CpA6dcnTO
9+060fxnazJbu8SDRu4oTvqDLCpLX2iumy5ONt5KfO4Rce9Ikrimxo0mXA04p0fN
eFe6ZYC6yM/OG5hAa4m3Rg==
`protect END_PROTECTED
