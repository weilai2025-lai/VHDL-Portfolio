`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzWu1ZQLrmCDC19fBUAnp8RY3Q143iSPsk0Wsks+d1WIqdf3YkaYW+/MfZ5v9mUn
RwBpgi2bsG8GkkUyRfGsw6FwsYb8dD0jHYn3SK+XQjJJ7WrIQJRL5b260M+czgXj
vcfbifrZQ7RtFVrfyDLQFxpLdVPjAYdels6JcEla+5noD5GEXCDL9AfBqgjPBPIh
aIQopRPLNqxPSC0DO2n3ztArzl/1Yx3t6zQRvZW/05BGzdpBU9PO+bwX8+uHnT1j
0OP4dA40xo+y5SMTgEQWIBhMOOI8wXNQ0GoWzrAnQ0LzV2/V7IEmLixOBvnGYERt
4Fe2oqXBBeLymk+AyvRz/Ac5TCdrjNfAgcI/PcHvsjdcGYV3jrS9WK006kkrSeUu
ny5MXqU2VPfx4adCUzi0Ask0q2g++Ck4W17BVLv7lZtzsphDNZiXdGlqoEydAEoy
MMCMlwMBf2mtOskYw44+hR2raCA3Uq8lvy9YdfAvrQnTFOdTmrBVZZqhrpmZcuGW
axOomyTeYWj7/Ki3dcOKGz2MUA5Nfry6WlHNmNXoE2/TbukgkvRDqM7oLMucy7/F
TFHlkWWRb5yL7mkZ+DQ0OwEEkkhOyeUPFJEyr3tHFT6FfIl1lUQWtWvEfjdM/0d+
lX4jy3jGPpAgVa418ZaO55G/P3OtSih/NC9bVUogVbizNflV+CUtk3Y9+FuTQrNw
2OFKUuedrtX4blSBPgZTvvy/uTdIq/ZXGkktMfsbuWJQDvJJ1QSEO3NjiZrldBmY
0CY/r1wli4zAvM8f/DWfi6cOoENdsWLigsvr2ZQqCR8OA0FZn7Rixr2CLyYNk/QR
6MhI+wVOQLS0SBt6gYmkj3YcPHbgTEtFoz1RW2lDWgzsW1QcgwHzwQpg64y9gp2/
2okOEk/OD6oh+BI3Pc0+RePSS8cTJkE3EE8YbYeftVnNt8u8Z6kvVRkNaw83lOSy
SXirmF9hgI7O/qp1DgR8mmChS7U/ac0UK2sQVdg6q9Wj/7te5uBJWCbo2pCLMlPI
Il0WnRRvoLoqPBbHikfnJg==
`protect END_PROTECTED
