`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eTsRRsFslYfgnKV/qDcfvjSF6IUab8g1qGaTs+lZSIkS/OulxFEx6c3W5totCof6
GjjBTMakvPx99oDlBjlgPi80NK/bxa3FROoBx1BipFIW791vkxYrDz0zynqZ+KWX
NkWxTMFCNj1tRkUt044TecKnXH+Mig7BU+/lkeZRsKZUygIugkncUQHPoaFKOMCF
Pwpyb75yFAhTN6c7vhh9zfjV/yUD94wFG2J1ea3PnElESRHlT7B0ZCUrmfyqTDge
wT5tLFpr3pkUou7MCHPc6ltLRIxfWQjr2IL0PdM5Go/Mffy5jC0b1oN69RYvgw9/
cDf5fHOdOQ1BzC4yrH0Sv7m//sd09a2TRCVa+iB5+wrjqxgKtwS4VKRy533JKlbe
J7ny+0NXvE5XExSoozWe3khDmKFkUN9u0r1XcQbhyF8bTwSgMJ21+aE0TXtOrTW7
R0eg5sryAZzICkN8cEi6CySLgVEmHqoftl4eH9+AtHHqpp868Q35UK8RDgo9tyfv
BZq4TQ/EtcTL6OJwt5blA7qRM57ZI/M3KF8FOwRklgR50m3DSyovYg803PU4ToLl
qXxG6t/uaGVq++4C71Prq4AaqqcPNLLiu409Oi/J/5pVeRFY+uVzGjoHTfdTqUIt
zA8YAsjwdz6B7+S6Vu3EuKqljY8iPJoYE/WV1sqKNe5BkQwyiNSLx+CE/q+TB9tJ
OFFQIylzZQ/j1zgUfK1K9DoS8he2dPnSHTHy+uqTwsPiV0U7oNeFHx9vo4aysjqv
RgNsYMZpfwkoHidAqlATtJE4fR6289fmihJ92u0IR/v5bcug0Zp7FQGB6L/EAcs0
GqxiCd3moob+cJ57dlOHQrBooPk+XnFrOIynaL1q7mG90ZsqLRk6REXp60Uej/SP
q34ONTxzkdLvPt890JzmFMNzvhzCg1F48uXVTMXFHv4fYnt5sllBkyyhKcH57Th5
Th1yYAd9XLpZ1Ak59lfaJKn8ootxsNRM3YsoDxbh+dpDfIqCfBmtYo48p4KZEIec
HGcjHwmt45dcWxcF0CKfKOUMyBxZTUKXIWI4nhRl+vrtjzoEn6g0HftsmtymHUDB
wsQiLqMyxlcfbCOhhNEOOPScbqixXi4F+Vb1EVXCE5gyYXdEiWbAZ/5ULH510AY2
3Cd5hUgEpzc3KEjidi+5ZbHc752K+aBM0wD13RbbkEi2YsEPksqUiyYIJZ4ddIWz
ondbQekVg96LnJynMzyNAwHY79iAHsVJrQ0hiN71uGhHeA08RkAG5whNxqZv26MD
xuAs8q4+AH5rEbjBcOdbkuCM2t/LSE6p7g7t2qBzPzU=
`protect END_PROTECTED
