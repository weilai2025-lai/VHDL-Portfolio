`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26lCecr0WYDXzEmNHep/Xt6wUWOIRgyU6JErXExA5aogcq8Gk1Se+DOcU3xvd0ds
HDmhynqb3klD7jlL0R8Gb2tYLaeEE3eChPs41C9zLnhNYOlxmrB9+DgSZvGxLYkM
vJsc5+CnwMT+DyfRJt5ZaB3ElDY8HMS+oWT0YC/cAC6DP/wj7g4XrKAB50AtVFV2
2Vr1GnNy+g/jl2XnQnpWILMWAzCVmbcHm4v10HTok59VW18gfUqkRl9Wsbv8CNHn
q+25dybUulTjrkZkdLFHeKJKsxBHq1Ak40m1jYvIUgynvOWrkw7//q0NDaTga6Nj
HrRQCLIy7lHT0FMUCY7xD8Lt7qHVu8Hri0ZIC477NrnuVBpB9V9aZExJ+5hZ+W8m
XyPvfCi+zSu4hj61/sni44nFSGtN4cNtXd016DyW1O6YheN+Z8yGfN8jnAJkmQiu
/oNHf6VZt9saGQ9wOHX0aQlwjfse8lhncMFudxiPuxY/m2pYSflZMxAEmOAjfS3S
6jiMcEJPk1Yw1Orhp4PbOB8ZAnOucYJWZZDHkKdbt7ogcuLLiIaXQ0goU5WMz6Qs
`protect END_PROTECTED
