`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNPXJfcplUbImdAPH7ycNlqeD6b0W4pqQGOaN7+rKDbysOK/Qtxu/6TyaYBYPALY
DTLe8Ueg8S6xOx9bnERW521r7PsGG/EdiOOrQSaB3NnocUaoym3j8abr0yds9OJy
q+9ywmHZwP6Tx7k2RrRuDiV4P6jO2ZuJxBjcpAbRq1HZF3CNdfFKM+7m54epx35o
/dYRGvayycIZxpUV646y1C/fnnXUbt2b6cWjXHmqjaQDBqYU8kiIkLWRJwHWRsWO
WmBvb+SPE538xEDqMtOrfsMm0mJeQjJftuKptprf8jXDZnTOvxW3jB1nm2X+WJg8
7jeGjViii7VmKbSLizeO4M0Sfd9frP+qquGxSRMVwG6isdmn/XFn18x/hbqLrMNx
dw0PI1fr7WPyDI/xnyBGybDD++pRJN35JG5m5rjI1Xms4sY+Do/PzC7ZVwI8rn1q
1jDCK71dOU1H8T7Z72LBq2N3ZOovHc5EVV+cJcFYVpyJkJK+t3NFpDgENYZ5y8YN
KLyK4NipE+e1PZikrawoFpcclxkxxTIjU0QWCxzPjYyeU9hQg0/BNDX+R/f6i2QD
nYs6F5WlK0sIUmpv15IYhxfkeeEBNkfqFXp4xL6N6a2B79pXNC1KX7mXVpYwYeF5
Y5A/vcPEHX0uNkrENsE8B1o/KCYJU7r9drspM+QMH06yleu6VFE32w8fdYQEB8iB
ker8JXasHcgJWI6E1LCocpK6wuSJHy95YML9gCRe80NG/Vm0CBT3vE4kNb8OdXUA
ayOrZob304ubZLkehNHcWXom+2vGBB8ytxzCq1WxPxFP/Wz/uBPufdzRWDuk8+C4
nOthOuK+pG8V7gM7PTqWNuEA3zARqb1OtWeldsnTUS947ymw8FtPr1lgmxv4lSfU
BE0U0XrHRpY/QYWMBlGAty3D3ws9TLb6tL4CtTtKG2RSr/jbDLEIJGVhFlXJwcGA
bxUHVYnGLp8d95uZGGkD5j1E3VsjwTS/JpcflrVUfmyELJTO/KMMtAEpYr1bhe/G
YGwZiYrr+IrLphFLMp2qp1fMnHxibG3LbZpftMuzBpq4MrMOX26xFWhBOzuEHCQM
dcnfh6hX2akmww+eEyKNVGksTcRnsLFjvSENfeNII6ar2SNf8ixgE6gGfiMAiHaH
Feq1FNuqTwXvIl1vZs/T99exFLFtmY5vcKpTHpZBR64RjYXt1yCQablvcETDbd19
Jg958hu67ybyXEzcJiF3xweOwuQp1a3Sad7/Q5WLs1nQoX/9RAwZa+44M4j3wppz
zlU1QkUsEkwpQMonj7/lItYvZUw4SibD1B5kylz1jMv/LdoWySZkaeGh9sTRbZMV
Yl5rdEOAntHYZPgrlsvPKwpBZShZKOJM3s97Aj/Wj9hyguQ5PmE96xQhttfXnbsF
dCD35xaxdFQZ6tQna44pNHR69msDSmPq6RB/q8+IGMHeIX5a+DmFZOjomDZPgq2J
fkKVnpXN01oMdfHQ528tfHMnaobChDMQKxIXyi+6inQ8qoAfrN5ktdOoikob663+
V7tMsupYOCq9cNQldQDW71OWnbLO9gpUgRU/H/uo7hsu1HepHcLrTMGiLARvBolG
cpEfgAxqJCWvF74pTcVAMT7P/8DsfjZElooENX1CjSqCuGiL4YFfKD42obO3Kebj
SkccuvHejPTuS854h3lvDj63+3vlzxX9nUIGyCwiJqyq44yH94ghoYFs/kT+tdRf
`protect END_PROTECTED
