`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxBebQpOpVQR0s6IYGJnKWF1boynwtpUJjEbmQzeZtx0NI5wyTT703xsIeFhckPw
5/f26Gmuf3scrAvqEUzUJaIZ5DR8w+eW6Nagg+T08tuWJhIiH2iWI/1Cm4/pPyJ7
To4Qb5UDpLtrlbUVU4ivSOszhxHjuLOphFno70xl1F6r3x4m9HWCARwMCkNFeFzB
l06QiFJf3GbdLEeR66GpJ5/+9PHGMqTJ2Yhq5pdICHGM65O3v/nMGqGPoE4WBPwU
OzocBbXhTjRKht31M/ZHMdTm/MwPT6XidVzKUEt2TL16Owc5CagxFw1OTYs+Pxu+
hTTjIO48LUHb5PyMfom+CDbtsTTQVxkj/sNH9hIjHH1YsdNAywB2e5CtUecFHGo7
OdUdc2yzahFzG3OsWNjaOotG0VF+bWG5VKP5KCx18Xxnl22e2OWCEm+QtX1MIcWQ
dMHEV6XMymUgw1iMXwUUYO/J0qr0amSgFejRfEUSOVK3HGkimNNWOcgZBstvvvHb
IkcBGWJSrd+KMdG4SF6OtOJ79UK0eNqSSMNrAJZ6xQuQMFJ62blQnfpInKK6XMrS
fu7trJrRByNbJLAsbt0LlP42hMxMjbwdn8Lg4G6ve3HWH745mlpVUv5iOUQLYkpx
iV9cVMUiZ2BWZDKeLRC1ZLQH6fq7CgbTgRrfptFYKIlbkdt0Geu6p6hYt9JOn7NG
Uk39GjvQvMqKkJbVjc7MIGCg0fysC4T0+MsDSd7dHZcwbz6yHWHl5tm1WjSIDdTo
jx7+6lLvbl038wPZsMRcFkTR1yacGUXkzvHZvzEyUjyNADl8hUAjgTVnWntcRkoj
fXH85vA2nXAZcNkYg0uuQ20jYmJ00Dt/drZFjm989gILAJskO5atsFFVpJDSp9P2
BtdC4PXNWuhcIrFV43GarQWBwGak4KGB6UL9V2SWIDjfnFG9vX0g9f4mKSxGZ+6u
77d5Ey3JVmRie4ymADDmPPsUhME0xtcHHUvRQIRkzqHNoMMqanzU5pqi8cjEqzb1
fpvcfGUMhb4nPHrqkbMyqEPMX8JhChmprJp4bMDCLIi4bXmypdk+pUCzKgQOS3nM
QaJtKhgvxxumVplKENkRSSBobqniDOnuqgLLaVKt4scNS6A/Lu7Z5ODuEgp3bkZp
5/N1AbwyU/N+DJb+4/bcmK6A46HOfG3usl4Q2ybzjZ4vyOCgzZJ7D7XHKBXgMQM6
Ouj7MNT8QmGxXJOIpiCn/2RkYfza14zEaRoe06zAfwG+HwqIrRi3srqmDzpXX+jt
czsA3ePBSQDEz2Gx7hBmuAf7uSEG/8/1kVs7XKuKDZiCCu2j0Nbv+1OdxBshq2r7
sa9Y+ux5lJSk9W9MWymge/TWRIZ9E1EJmDCOvjfda9VIzGppbcN37d5w8Ekr7nHn
MgEceTz4MENYJp6WSl4Gl8Hq30IitOarYhXM30neKqvhCo0vVUKMoUJX++ZnkFho
qfH9Yy4IvYLDqFluCITlEFextHirRuWC6VGDlwIbXsMW+MD2sIs4z1r7bdojnxpd
VXa2Ysppe8eq31uNnHWwcorMtjgMzrHVTaTaq25hs2czXyCMmbFNIFqTMc127aJu
8LQOJ31nNkssh3fn9N83Yu5xty+4ik+XhmAkjNYzLdi/if2v8LuDez/vUGa6divK
zb4cHC8GRfbvb7r4RB36XrdvQa/Zzw6DR1JYD4CIiIuR2hUx3PSFNJGnqVQTqS9g
FSEnu5smbIBTpaIIPCGgnyEnN/6QVX5N/9Qyg+D4K6JvXpp1EfnG9XwYs79JSRgQ
wI2YxIAZc5iAHnRGIAWcbl+tc0a9lD5rmosRMa3Bh5I9X9XQA1y6Z8pdOxKj4YkN
UVDvxB5fZQDyrrVQr4lXiuuNjcA6y/IZraxQaXYUOJRpkJoDIIfEpLWEutiXcs7H
dfpyjW4u6n2O+ipNmj4I5/SyQUJ338YEzV19lqNWM/AkY/E1u2aV3YVO+l+5Oywd
1v6uqy2JLx8Ns6nr86mm6mVm/lYM1JX9Rc/9hyLyQ3Z0E9kDkqVlCh67T+5//QHY
zbZ6JoofmWvieqOfFIOulH+uVynYXGn7v90mDV2aLxKDsd3+TyYEYaunTLuEMwyn
ycGfQrFlfj7kiIe0oER1cKfx2uctTOYwaFszPnG6Bqwy/1PVw0tQpaF5h0KhesRx
qn6A31XtsHe9UPq9YmPm0+YOdipmj0nyoMn0DWDoKpkRDn+uQb4NMjhkfrVs+FiJ
jsyui32DF85pv6myAYJetQkooOQ/eWG4jgolZlzwI3VevWMpv6RoaAULr8oGHDaN
4sJOSzM3arw7TjQmFAq1+yFy264fX6TLVOY73qbe7RTDeWPjZT23ytdB/D7laORW
6j6Sae0J8Smg6+Jhqz0GiL423w4CFZBIggzOMdVKKSak8vm8jnehci61EizjkbaS
shKDK3KiX0rFHQynUXbMUeSuOZuJqZqJgho4UilY9d4irIHLSLU43dRf3F9a9QEz
sDjpxTXkDLsFPANjktC9xRGhRYOC6yW66u0ZulbHvNxqtDAAD2TQ8ml5QW0rtCeI
22ctHSf+3QdhlYl02TnnyfASgOXdOlL3vax91esxUtgGzKPAOZm/UGR8ezYi8FGP
n9Sbh3mHgjpdXgeeNK2svivu0qVAa9o1LFgOFcuTqN4gHD8bIVcIu4jC5lBjSjqW
yXbjPiyrsNhjknJY4qXXAUruUV6nW2e7N2rJFATDmw0KyDY1KRu9l1f88FVpqgR9
m9reE7ITdDYYuU/Mn3PaUXTkfo46769qVO+olTWsyco3mi8bSEyPjpxUVq7/yByY
8tD/ww+B5Ot+g8/KpxGm8RpR9aGy54DYv+SnNcqVCmdInJjCEQH/dC+rSKdzAcR4
bzNQl5bRtYIml01a53OcFkz0i6hz2L8BAkgELUTE2Z4z/E155FB1xG3MntbNpLIN
/aDCCi65N6oOx7rcR+ucOfZ40fLiYxYX3IVw+Ex9wd0L/4cAlnD57K/Shdwk9Xic
eW7TfxwB2kLPrcSmUihmW1odnyHlKEcL9AdvYPKNaLFF0j4J/oaDS1f3HvMhwb6w
3e1OYj5dDfWrNcN0TzixzxeAPpDGBN5Io7aBQSgsfjy82jPinIaySEfcCjGBuwNl
cteIklxUAmd5X9fKGh51ZJ55A2IspHYC9ue6W5NmPC+jqa9xYhd7CNs9uAa/KD/M
M9Ii49atnXTeOoD1hIzBYBG9udOOfNRVj6U2VI2dM7TeoQDI/5tGhW61ftAiazJw
qAHBHn+9JvOIetGxgPR9Idf4UVlCmCFLfC8wlcAkFulyw7ef8IfwsFKlbjuPFiOk
i+6lTghroOsBTBuK/mXlrY9akBgsbjm25EMYbS8JMBuyzbId1TheXlppEk5lkmXF
zjS0WmvCO0JE19ofN8r8OYfwWpoxRQwHzHZYJ/JnVEbYjhT7tzyY3Ohl7PXch9PP
JGMs9Zja+yee4tIJqCZN2Cbj54Ai4L3rikW8dShihRIB8ZMC9UIaiQICCoHpJWtn
VQJGrxu0rLyhyPSGDI5U4qm+X1EdR7Q19lR+8FYa9KhsqKrWhlk/PuWS1BDEnMX/
8KAfXYMscyuJb9vGio210yKP58QPj1cpPDek5Q4AqgHkSf94AUSvFpJ8V9eUSXPk
LNhyvMWdsy60v63C1EzF3N9T5aksTQy0U9mZreVViKrx3ytCRHoxbIzF9zeTn+P1
KstJkFIr+AOywxA55l0s1KFMTPOE9LrB01w73M8jVEBFsCRV7j1Z1LtlUPvPJFon
6z4SUPMyZvaC9Vxf5okxhfN4VyJwN4jkCQgm9Uoeklban0941Jyo//6Y2qWBKeUt
F8fHgjvrjhLt94EIyWiblBLqfm8uj3CDKyJ3UHcG/xBwVLH1DqLqCvRNyE756W68
oZhTuQGDkKTKZSU5CvMBu5j3cJH2QkX5Sp1ofKvpPkdRhbVBoQOyqIcPMR4mfcMR
NGMJ1fRV1gByyuqslgrp/dkMgyG2DBMrB2yz2PEdoWCutCFcSgxrXE37XGq1LOSA
5fg/0cBVfZJZO1K5WaLfyTDKMc+KIx9OwAxlYKN6zTdtzJnfCWE0DhA7FvnnZDnb
`protect END_PROTECTED
