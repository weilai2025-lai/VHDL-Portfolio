`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z4Mj9k2CI1TxNvkEPojsv3axFKJaZGGSjz8hvDEurvae+pSh0jqfKq5Z9cLeg9Gk
mkKE7DU4GGN++PuBemqg619eXmSy5FLCnRMuQ2dIQ0PL62u5FJmvfql43BeOiRY/
ocwUE+1MHG6LAKzK/D4qMYvXsFZ1vpk75ug8irqlugEeptuHaIk38k7Z2br9WDdw
HmoOVtkpmjmlEttg8fo1MT9xjzYe37qydig7CSDIiSn23Me3ZxV7N9oj4Vz1nCqk
aMViruXEYv+3hFB9XGF8u910AvQNROtIRbiVtMsLHnuv3w+g9fMYVl2M1KPWfh7e
Hka5rGLCbSeEz4tAcugp9jRD3ntlStGHjAPB8/QloI50N0x0q0Pd3jssLImORuQj
s2UsSh3R9yp6KEeOrAJ8XfCuivae8nzK0BnWRS4MXQu+psPV2zhm/L0T24Hq8/KB
E8F/fqu+rGtxt/HdUIVVJ8mK/wxcyHtzl+Je9vHr1ZGBnMdEvgSA4rs1whIotafy
uJJZmryrGyLjGp/Gugd5ORBO7V9osq6ODk/+jxfrA2SlbKKdWznTx56XL4dlZVb1
OiPRDaE6piIW4dLe0j3mHYhtIyC1mbYquNgGXbzQ3VlK8+yN2Ehg7RHqGuOnneOI
D7jv518AnqH0kWNJWu4xIHXB7nkW/PT+vDpgzyEFezcznRsbRK3tend4+lvpSl4p
zS/7g3Q1WK0TdjUIcRTgQ1fHRtVtOC+Jg7lG5zikmdbxGqm7JNm2aN9HjGlClN4G
OVRWXXQ0ihUft3045YAK4aarrZ1+mALOXuwQk0TpAPiQ15Ukl9EqCOEBLq7gX7j8
`protect END_PROTECTED
