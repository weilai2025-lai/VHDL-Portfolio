`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fz8tihbeGfRV0CXjoS5B2gKVXWI1fRCvMy3pH7z56Q6HHL/wxopXswCiYPrYkvJD
eAMfurJykt4KeBJBE1ZeFa8g3x/Rdtf+TYWEv9oGsrUgkmTo6uCNowd6LMsm/oD5
JHr8q7KTHebdzo6p1iDq/zy8YhY1yIGNGnTSpJurDXydOjNWjxVDyaUver9J9o5U
c8xAqIawF79XLkd9BVsaB53VjO2SoiN6z3/zeC/FUX1Mfj/587haQeq7TRQq1S7M
g/w803PwlAlFwzysCPIqcLf4mjqJIThlNM2pd5o+XXMmTpGmhq6+24H/RXUMGXay
2jRFgZcMPb9PDmmdwO3Vlbj7lMyPQEc6QM0OXsypNcu0E5M9fsPiCbO/BuRaNwrV
z5lQ0hMPSeaZjskJxQIRwdU1OMpNSveuo++HL3UIp4aSL8Fnx3/rEU4KhYmi86+V
zjsCnzfCUdjUIMctCh43ctmIc2TlN/BjxLh6U0ki32mv7zPOFSZDprV+qyMJvXln
NkdlB7HSsRcvK+9X48t8KDpyHV+iTWZMHcF/3hGh/uP2LejPGge8Og5ugUN3SBan
rdiz+dhtnZgvd1FvvWaQZHeknRF7TAPtKzJNhGKk+wF6WKDf7EaDf8sB/ap1bi7y
lPhrwt4Y/TvY9yiztKDM6O0pKmSiZTGn/5raCSUM7q9UzM9HsuBgm08dhCpaHEvi
HDTy0OaXoZHHGmfuZQhQ9kU7i4+lvjUNPzgB8qVGuA+zwiwm/lIi2GCcoYPZv0pC
GCA2/rcQJY4y6aVrtMab4o79WNo2SDbhM/eKgZvSfrsfChsEij1meR3hOInJTkvw
pFKpp6NeKc/268ydE29spVguDiHGyvY5z09E79NzTHsKXnZIV7C5D6QMCGj+PtkY
mHKdZpYQ1rXrZXk3gvRN1w5RxtQVxBNTgqc/R3Ju9SCbsYbyD549Zpr658wVuonS
`protect END_PROTECTED
