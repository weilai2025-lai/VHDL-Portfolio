`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWdijubT+XPkIGxqqpa4LexO8bgLVyrdspSHtVZoIBvVygxvxE4+lbfpvWKDfzyP
KjDpCT70j4qIYsGSkU/2dKI91uvcfpCjeppJp9z9ctD/UBsOSQ10bAcslc50LG8h
s03u+AJImri+vq0yjeev7kI6qhYZtgWazoJ6FizW9/jniBrE1WK1+IuHUrhCV3sm
T02I4/4FG+MRJOfUA/ILHa1FE7CH8SZ64a41gvXsVEqUer4WnKKCfX9xuSA99wp4
sxCOyu/mqh+k++lbWCwT42pWuyQ/IveOR1f1cvXLqpweD39aZbcBmnlNnjWE+E/7
FqvSXMvVC1fMig8Ela8z9+GPecxHZJIZQSq34u0cgRZEzQI7+JLHZW67MNYU5Ma8
44euIgYJowQbjPRaLOY3xLDnjnAhWxGzuP9sC1V6YT8T/7q49jMVehZrIQhKoG5F
nLSZFYuTdfdVh2DZYO2B4Fq/P8eY6hvxqZtsGDMAQ5y+XpLZYUiLOsoUHCraiQCX
NKMXl47eEujaEaSyj+Fkf7DxMC7qa8HMrl63aK1v3X/86b6vzChOELLbITkP+1P0
MBHUIfiJcbBxvTVmyWTrHxe3HM9C2MJeqnlwCSDxdUWC9H4s4EwOLOpAWcupgLwh
XgwT4XW5fYvtcSGrEd6l6++srHBEu3A476Jcvrb+fXxFpmPPuB7jgiTtvOtv1GMR
C1G36l0P84qKJK90pQSxQH6SDepaXrv9u6i174QmwhJgieLbD6YW4Sce+b+1uv/P
uxtPmFJUzwelIQ70NNeAw3XHMsPQ7Af68tMXGx50qlnzzXwFXElqAu19/HQttUbm
F9pHobl0qpIVHSTdg018Yd+jXDHG5x5xkZDp1q3ROrfXn+Kdzg6zxgFD/sC+jzGq
1czFak1rq9nBe+6X6G3iCpqMGJnyQr8IU92GC8d5SwrBPzNgXmWLOPWb9n/tOx74
ZkC+brtR09+AHsQGRdajKTCiUOMnyN+hOwxvgtfSFopy92/TkLmpcsrhN/0JQRO5
wZWv+q9D0aK6vl0utsJTC+r7rKuSoKi6BVsuu7Ze9rNcLwbOgEFBG/dVwXCA5HNp
ygqWVSjo26JGrwQwrz8VpGqWMRhymZfVNt0lejYwhHcGFsXL2MiTzr9+ynxd7MKN
NeSK5cSWdxTgt7NOOiMjx8wkF7QYvH32zjkOCuPmowO8R7b/g+dWfEo/jmHVL4Qb
KnXZP8t5zkwiXKEsC95MaRsTjbQmVmEyNTS+tQmz60ll1R0z51woccociTCM2UvA
zC0T+8YNAufuSFKQkAltunOa4Zxl2NWOwIvmEfgiz/cDBGwwOguPCpzl2qS0s1Z2
s8Omam3S/wLOwqAsFp0QEYRqc3f2Gejvj6tSQAZmmHQzjhMGIL1bfrgKSekn+sKl
D33FhE34HjUhyxzMMDPwE7QfOtkBYbygZ/0qMPzMv4oyV8513J/ZV7o7wBTay+KW
ZObHWl581cVIwiQSZmbAc68PxlqVEsWBV5MeaDAg9swnNmqDTZm7OYf8d0e6AuQw
Yzt5OTMYRbSg4Pz9GXhKer51h82aouHLvq/o/lQu/Q7Ft+Khed22jspgpqxHvotk
cjvMkjE4xvjoHt3KzI34Cx9or3kZYedGZemjZ7zOHveTfcKGnvwVobsA4VrIx0qu
w5kZS/SeS4SxbOb/J8YwVFuG2t1uB5X39JyOHxlen0elclcE7b5lfGc3ipxNEoXi
`protect END_PROTECTED
