`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOKiIEEeysU6y4jvLVat1q7LtWCbvZZb6fETaU3XjNHlH0NX8OiWu90+00wXsVdW
RMgHtHgioEJeASjfcBlgcMci/pzYw16dGi8KdRe6thwwnMHSNfqm4hGaEpw4ayto
fgKqKcDiViKo5Y+0Sr0/0fpYh3aaJ63Ikwy5n8VfJPVNacUu4FprguCB3FtxYz6+
7yoKukirCj0lLBmKWYHDRNkKR80jLb3BsWf8gXmQ6NfgrxgozD+dlfJ6769nwU6+
1X/cRZ0yOemvpgjrGqHh8tVNLGSob60Pw4O40heP7GV2KzwWktukuiS83t7a0rjn
k9fuXwVPuWBdgQTL5ScKgo8EylN6gP3Kz7Ijps7n140YY/PihovIYmFUm03Am+eN
pv5ZJwi4mXfvpsPR2LOHdL89uerbjGWKyFohpZjZGwEr1Vst2V4pzXhgZ8XybKTt
cYq0s76NVaApHSNSizAISxEDg3FkQ6McaI0OAh55ZS3l0ZtoGUt6Jj/Q2nqjPW0+
AL3WOifS4kTnyEfb3rtVcQ==
`protect END_PROTECTED
