`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOG6UWZ0OAQpFoR3+nEK/Q3tEWtB6oLil1LNUlgfoKdqSKnaxzUBgzhlxPUDFULU
qH8UA98R1kw3ydJJooLrelxE3swG3SavRx/tc1NAV2FFDm0JDNlrR2S98r0DENjW
2K6e7+lpAXjaS4+tMWaT8iRIk5Cnmw/UaTNY2vKmvt2H3ljDiHvR463woGgQe9oK
+B1HKr6Sdk8TB79Y6xUOoP12phVVDzJ3kgWDsyDNmP1uXPqfX7/byz0N0c7NVVJe
K9xT79VM8hLbgm0JNYZfmBSsYhhISeYgXr+obyS2H+5VrH8rDDsgkK/oXE52o3qv
btKcM5kFnw8/OZAmaeIgJbZnQCrT9dcEKPGp4SJE+FMv80GdjPivK+wK6f/XjAkX
thE+mlXrRhwWefIj3HC+BvhCvVAnkslu9csnqL/2cC3sl6c/5BrK/k3XhZtli+FR
1d9aZ13iPRyNMtS98PvlX7Zy9tMd/by0JAJCbG47gR1anC/Zb5mcSicfNZVIBB1a
/z13liwFc1pvE/1NeQxu1SmTlEUcUW19al0UjTH5FIBpxDs/AoI1eGWTfNhqW5NU
pZidr0NB+SucGYu8q8agcBheQg9Dc0TUxXGdpkN7eNnXmn+TlGl0WOmu/qaD0O1z
BpXoulQfFV61r5YnVYbTi/ZF4KRvGFdveXfdUy7QqBctQ1NGnJJBhhVc+/mMGygX
qW9dozmE2Fz1i2uqhTnNscwdDRs5FB8yGBI8s/a+YEIH2CxPD8DNmYqh+TxdPzsp
Ys9hsoAmm0zNUaE5xF1k7PCjcHOC+wZfPoEAA+tiBlutv6P+qvj8p2yqp7h9UFBN
obLX/qeUQJZDeJt9kAJfjw==
`protect END_PROTECTED
