`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8nGLyhp1PrVSNp347jNYA1PnbGrrifiYWrnGXEza4+SHVxqsf3Pb3+xfERC5d81Z
aW6hTgncgQtczt38JuYX/KUauSFnyIqlebfpiounok79yJ8ZJElX1eEC7htgkR4c
HDXeMlLtBNhjTY5HKk6ElTUCRodTAP2UTB5E8wbOskYE2WTlOlpqH/gtHwI1oyNk
1IonBb1XIpdnm+gMq+/VlBIbat8sFiClonJKgyf/mw9fexkDX/6gbHEQaxBy0Gqw
sGCiodsw90QmBGZq6XjSrI14pHI8cjXv1qoOYG69DqIhV/JJpvNabcf/iilhfccU
rVhS7ISV5TgPQG2SXJzLCFZglXoxnlDMn5UE5vUKIzWrqzd3ZI24/arMiiZgWzV1
61zOZW8l7lnqQdeT0WflLYoSs2qJEvEM9POR1HU6NZ1g5+e9Nztohfa1XTqN9KAH
aXcIGJ5WiZp+9U1RQjAVrUGsxdAzX28Mi9QI/MUvyhPcV2bQnBUvwKBqEabqMwix
euYynkyK4CF7DGeREmLSKFtbYJzcm+N82UccYkVbuXfapmbASj680NLkgGWoLCaO
xdbk3D12JZ39XRfxC5Yym/UKuUOM8MXhP0JumLQ7gev8DXZZoPYa28vFRExgi3am
lKQPwkeTHeWEDsFWaKkB4wUkJjVPVpzMXc4mZ/MNwm5PH3OBcOy3Cx4EZgzzKCdz
01lGYtYoFvq4vz22Kp/0VKRsEyJABb1jIRqAEHvfw0Vgw6FDzrkWpZINJM/Vh0t2
+VXkObeZk+/FeBwRtTJaQgYmrci7+5qjkm2s3DSWwHFao5bNCpy39qItPHGrcoFw
DzyyKwrPme4liHXjku+jBUe7fDvshFXXaJagbwDzdO+u3gPPgV3ACsPBwrIQLh3H
mjFtKaYTBijZY7nSq1b7mTZIjCLplvkDvJYHMyy5WmlRqVIE/5Z2mlIA2+8iFrUv
Gh5arZYsmI/xhZGpZ/z4Zz2SRGyy4RdQnFAyCZgdI3oNpU4kxFkZ8J9inpislK2m
C5Uu65Ynl2Q7B0kwP3APB8CcFcoUviND9XJRvR/AMUf7M2b5F0WPG1m4D9Bswm1A
nTSPf6akjuN4cpn0A+BmytfnxJxT+7UdDtBwhkx9+mU1qozTwMGFSX0oSG4kL3WU
aUt2CUmZU91nCCq0WBE89kxPsn+pI+0pKsQjtiCXTZCt5Zz78o9fSoNRyOXJbbpB
nQlKgCAu4oIvVEJJ3Ro7u8dhptur+T4YUVvGBj1elUHEfQEVwW0RldWZfz0Usfn+
YJhyOkKMycWUElbOaxqkarmOhJohEsZIbXH5+hFPX2eSWgHQiULhV8quItWZ3ZMX
z3pcOWDG2eegc8MM3W42hztZjtmxbnLckLm2sHoTomZZUnK6NJ0BW7gzIeTtzWsj
vDbfY47RTLzv1euVMdmPRhCelb1TSaLUH+hCEkq25xdIooSyMOudFS9Bg1P+rWSn
kfmUl+WMauN4JBGJI1q6RippMM9X2rm5wPoAlHzOYETu+SLdHWk8Y7Bn+QPX9Xsv
uAdC3BDdJOjNPsdF484VN3FznDgI1Vuw9nBGL72sXQtK6yX/k8tVOiyFoWRt9so7
ZAcPfx12gecCeI8zHxY2N7GhsSqkKAm0iAU3aknpt2rsstawTQrBn041KPM9XkOi
vloiEhQGUakqHP1r4q1A5QSH4rIAFKTIoh4rxJODHpm3oK8i7/TO30mug+LiBNBQ
79MmFhbeBvoDoyF8JSO8hoa2yyV1DgMk8lnMXP159mbTK9a29KnNLn4oSny3hhj0
Ks6uS+/ZjmqSmUObpXL5b5KPXVUg6pJTckjopKLor2oq/Dj21aiDsDnQ4I44Jb8o
g+56D395h6E0iLibq2rMD55Q630mTFfmddohUCXVlcDhujT2VGgp3nrwLN7NnPe7
gKnmFAQZd0N4qf/4g7JMoHRrjKj6fxc9oLeNdLTxfM4sUn3I3tnIHq9lI2ckXR2l
XWtoTG04yQxybx6JkjetbhWoiNBYqsgr6ZlaUIZCK/nthdm4wuU7C6lzelny6zFh
MoXsi1+MADA2A6SYYEfpfG8Nt7nEbB5tBxuoDTewBhQoAeZB69LTRkaTBEWn64iX
9rGN9gLUYHbrfP8Y+p+/unSwysfUEcAzlU5G20ZrbN3KuyoE44e2unGc70t87t5V
igAiv4Of+sw/mkjwCX81CJCtfro9NBGANevCXehJybhJleI7gkNK19c4F/P3LcnS
gmMn0vQqHGvHJLlyxBXYZ5afBeCNWejnwGhtJeLkRQlJk7sYuf9anko+KWKSsMXD
kcr5o0oXgDS+FPTC0szxJVO6pQ9Fnim2XM1YIrXrszuKs2bP4zqcowG5GgbHhPYK
lNkDgyF0X6qrBnok0DdqrcPg3TGqsmftklpSUM4QyZLfB8N8wHCku8BaKuiBHG08
hjxVmslnrJ7vOaVZBC/tp4SZSuS5yfaSF99WqshxiX60MI0fSmNiiPeJH6NQV1zn
jkUDUuId+OYN7LMGOXzyDGDRXqxZl+5qGmSqIeaLWXMrsfJm377tBp0RXqW2Xe2l
zz4ulxjNbOmCL2QCv2LWjKUEx8f+SxV46OaWCe8wuRLj0FC0YW7OiMqxODS5+DTr
lJcf6yrWzaChWEhJfzHvD87/Na4DiuNd2cE7/3AnfMfYTgx/nDVCXyK959gHL9TM
vr23D86/phzxLApRwhl4mg4OyTO3cdJbYWZfYlMFOZYafw2VpIXnOiCMezxH+u1v
EUxjk3zGo4kP8cv1bA+5iN4r2QY9PYMdZ2QElnS2Mt+grroAla6YIo2FfizGHCnv
n5vvm56mZz0FgJLPXeVpWC5NVmGelG/l93znXfKf2UhxRxXl+2TYfnMQJ74p0xCi
6V5mZeuk6hyv0SoXiNlPTXLyEQ1Ow7YsuxkRyzsCx4jKqgsC1q9Pet8tb+rENry3
MJrUs/+PhmjwD16AsC27WmIwT0WAtrdNRcL4n+Rpp13sxUdt+H3G3SOR35NReSQK
NtSGeGChgFer3J/fjMT2ODg1JUKL3/KGFgwsA3N85fs15AHL8OQ9qLb8XWqD1m2Y
Oa5+lrwajPSEU1+atqghn/oPqRjuMA869cqsIiOIb25RBEVAs/1bWE0LN3BOSUaM
gXhaVM3KhOHZ5GS5QhnTEDsO3zubvctGFRvtXAabhP1TudOteCDMItAtq9W7IBqS
pSbJzIFYZyyT4DBRJG2IW4ifFzp0Uyi93GawLNLGJF8gVbNqXBIip5q+9bPtAqD2
3ehUpgt0MLsv4RU5lB4Wv9247PZrz3F4I4ocueIfXZFX8WMpX31mdH5mpVw+lq70
tvkZDFxEp9zF/ANo5iH1oMX/bCUExQIAhHTBhCXdGHcuzrdMBujgOiC9bJKlcZ1S
ntsVQiY70az9FIo47S8Gj8BBu3K5ZAkdwmZyhISYdHGQlRK88y9lLoqy4W/8XcM0
ZGR5+KXmsmvg70HWXugE9Gir0eeckZjHqmWzFSvIxj4+IB7I2fzaxsB7GHYwNUuB
SNNxb8Hbnii7mDpF5yVYmxv3e6oz2GOP9uYa7ZRdwntoYxcib/43kcGlS0dVwih/
5S2+YkZS4ww5hasdtYw/Udc6Vt06aahhyBubO8itDi0=
`protect END_PROTECTED
