`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpDnLqQeyP7iHVlUpIjQ6YEi+AMIH8kYNLihnAnpzb/5+47RkXw2GKDXx06X+Uod
NXxG/35qVb1qIbCi5PUSOMctpJaNsA3rKnswcJvbtTAOS8p+gxJVqyHpx0RrbLAX
dLdyAsyDZzU4N3pqGBTGH67o/X3j1qH1Dxo+0yOBi3wo2j1e5K0RgsqWE0PWxWeF
xO3ulhOJ2CsH/gj4r0liJqvBmZAIA0jKyKTSFRCOHQkm47JKrRwqqc4EIFODyIRx
YphS/SDGTfKB01a2xawfb65N9nzx/pq52MUkA+n5beZQvENH5+YWszRHR3z8VvwA
Uv7JrOuoVbElwI2fYFHj0WloNsE7Fj2j9N0N/smLYw+cnI4XpJC7jGoAP2QURqim
cdz7NWuo1W3zRBrAc2dlGStP3PLxXD2fvkMC1VXVv3n11nzdMyo4IzG6Uz9cEUHs
S6qrbNnRBFEZoXnPBbLNm1oQviJaHHqUk0eF5E5I0oGF52kbM1ZXaL2Ob7P0OidV
827ZT7bV2hprpFpucdo3GQMFiHeSrg9cdxmxICYOV4Z1ILi2is19skbwQniJruXg
VIvlfGn1Tr7XAbeAZDUdnVe9mbexyGPszL96AI1eA78jjDPUrUs+Pv9+12lGV6vu
5q1kXf04nkzoSwxLJ+31Iu+QOka18f8t74luDv9nChIkyOhJPydrb6fYMePdLeHS
K4j9hAvm4vUnk3vc8K5rUmSy9ILsydEz/jCt6jf//3DmnTfEazw3ZZnHBCty+4XQ
hVxQ2AF/WtK7E30Glti658cIaPPOXYNvHlFwKlps6LcoQSBhKKRFRQJ++wnuPXNr
cXJseD1iHfzkQxqCK+fMncmTZc0tWz0t5VtPB5zzR2Ykwy35kGQ6mCT7Hei8pAcu
0xHnFE0F4udtQWVgprpmwCg0cVGVcX2cxmFU/YEC9fajU8dUypn3EQ3sXKDWZIGT
olAwTaVpd5w9p3MC8bsx/04MJ/wM7H3DxC9s/C/vUHCHZBqboz47bowGrvmiBc3g
wfhxNF/docrf7zPTdVyLDDEJjCmYZFmWovkCRJ5xxWCQHxHjBvgWDkUQA381XgM8
t/Be3uORRADNQcqsFKOwi3Xrsb/mSAJ0Luj0zbnLB273VPoGfrQdGk/HNPy8GeJL
fMp29Lnhtd/qVyiN7H6cpfwzh5U7mVpcP4Vmoru2cX/oQ6KgvCT7WuWSVrNBjGdb
+NILENdbM6x4Y9nEgFAJVOttjX29bAbNmYZ9W3Mq7uXqvG9ZR+W1Om1RRSgu5wpc
2VyQAffeDGAunqDhLOMxNwB2+w1nRygBWfiK+Xzk6aguS9MP6G6d3VM0yeW6bwAh
KzXjWJr5IEKxFI3chsT/nDljjduIsiG6hPKR76kDDo4xOZY1y3waqPodLMGrAyov
gXVcr5hqdQ3jgdc+6YNg6icJea4qrWthIUYo00qZPco=
`protect END_PROTECTED
