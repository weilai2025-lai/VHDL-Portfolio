`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7dAGOPvwEG14PlF20QN6G3UVzU5zUUTBGuFmkOIU0ajvSWE3GwgBbP+UXwj8Nq+V
heYMUtZCWiwD44bw2JslS3op3XT8082H778D38eQKh3eIyEPBLH8XTuTQQrxr22b
0P9ZRHE0ZGiA16KN1Dv1KgwIV4GWTJVOz/J08bjwgG1gbTqjDravFinfj9EkV3tY
S3gDmwOoihRaUKKOSdG+KQn9qeqJKYmPMkdzmd5WhzvMr8Xv4BcmPIHpAenPfK5V
wrSJbGU97SkfByz9iX5dn3a8l08FxDk4rJK6eoPnfXlSWkf509YHa5c4v1q06ANW
YnM5IA9pOIOE3t9ruO+728MJJYy3EHawtAtqcZu7m85/7L1Awe9i+JxWopiEk0tK
Z1G8CIrxxhJVbYidPqDJ5EpgbgBHrjffg8LksYnBdemYNkAeSG1G/oXz2dLVGY0t
XWLKeOu/1bPfgkJYsNuzDNrqdl3xyFU2YL/MFs6KMGjuZ3y82ocxMMQKbqStesIm
59E92XqNs+vTGp2IHIEPtVnnEo5pqtl+Q9xa2yqqrAFPjYd/n9rEm10/p4kdBq6n
kQIx5IJipxXhJIG4S0zZo5pDjfCzmXjsee49JlsWSiNQH+IStqjYE1Yrd0Dg0xGj
Wo8jcgWZXsG6MTByPwAXuUn5wgQeutBUEt4NG7B40CD1STCE9AOfBLJatBO6JeQY
xOjPsHojbniNt8Bce1c94eRSFZ/yytzqV1e5UHqb8IcjHh+IjwQGNWMBXfZVYU0N
lmf31Am+0TIesDKMqKp02v58DqmPk/pPasxs5hs+EiZqgNtxiHLrVPAScfjUtfuL
nVxxPImewYJZMPRaRYvM5bydESW68ooQ83y21NbTP0vvEbzqODqittfwO3joKjUS
TDfdQsGpDIP0m0+nS+0vSfHoMztO4WOWO9QWT4wRG7q1EZS7FHzXZfXmhKb0kK9q
zcoX4UP2L0jB9Lus+U0wyQB7U6sQMLixXsn9lPh1h0JzLw2fCGDSsCOIppQQjsro
+7cS5kl8xMuZC2ZwFx/zTuNEQN39PcayFU1IIUsc2lSJ55nxQHSePM+rT+PY5FNh
`protect END_PROTECTED
