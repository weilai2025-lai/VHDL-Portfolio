`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYHyh0pOpkI3/GaOO0qb1/FfJm+WGKe1jOUV2H4fyqEp5G7YPVj20bLjY3H4vw6s
DSqTv6qVyna3IWHOK9LVbwxXGg9M5OZQPACjML8udmb290zTAAdP0X41tscmsjxa
F4NGKjtDbIsDhcRKdXpBmMr9kQhLkhvbRwtO1NzMwQ4EQ3NDUFYz+5FtntKmnR8c
fZxDA7WE3zRTLCgvV5phR7Tdpzl3WZ5YBQ69tE/RwS8AFk2zwejZ9zpTRcljxgPM
cRCbZZpWpp7KtRqCmz5j8+7BcSaDDDtqa9rGk7RIy/xgqdx58rF1aHuzyKF5wXlE
TOKc/rdLQrcre1uzFZ4+Gn+bEqmq3QmOkOomqrIRNGGtTtrHjec7MbpFIh/AvOwR
ECf2V2xqIfRcEaMWjRA1IxAym2J33oTMX4jIRD6JOQf4YGAVkAu1UxngNyUq32yF
uTMjWV6wLKDNP1kmhW6vPvX1Peb+kosjs3V7Be0l8TZZ+kUYoc8oSKGbUqjONwB5
HBduasW5XVzU6EhiE3IchR+kBqor4X8p+Sts8bef4cPge1eSOuDHaT68htAAt4wQ
XAkPKztIcMBXeEfwLKSXkIozRv7oQYq2lK8tAz+Dls+BrgKexciNHdd6Zv82dvAr
CNo+9ilOnkQm5j7Ttk8zL+c01T6qLFrrCZCxVYDRrVUxj7Yq1kwiBx+/H6pIf1n8
MPJt0B/XuJaXXuP9+a6MbSGuUZU5jZ5juknJu/aCD0qdx3mgnXftDwBJaA5MJnif
yheVxVk3BTVkuTSQoQdLqM+0B2GWgBJih8u1axWvuYRrGkT/w0m5btj0CspAo00g
kLkncG6ddO3FYkTyNL3zVzkF0lRGQpiJv6fmaLGLSIgvkQoJz9UNmEzhfVoABPqj
9DGW+GWS89GKBFa3WEM7dxcrg7yx18BRPc3iD4OgCp8wOudLJFKLnXHcmdqavDvi
qu6HKfvbbIJLRtMH5DIfBfqSAesUfvgWEwBnLu/Kcd72sru/YgEviZIdSPkKp7FI
TjxstfY9R6MoaYV0XRPveD7oRHn92YFFvhhQYZSHetFL3D6IBWsq9mtGAyfuaSVP
+UqMl2k006sz9CXVlyt3sQJ2zWRsxwmED1AqdtcEwFRPAbFcPJuZwtn8fF+MR9/a
XiMBKqDlmRE+/utzRUKvwx5JkehMr6AIxQGglzEbGJ8KCBfO+9Q6RO1MmOb9kljB
tqsGOrr3RsiwsgsNzmJ+ThTisXWJd1sDVGpVXbM0RPAhK0XdD73ZXQQwZQWU0yL7
d2groJgMGZkNNOogUeyf3LSpQoIaBePg21WJkbG2acp7FiYbv6tH9ngWM7n1dooc
R658lP2DdUDPMUF+nUZCDtDoCh/wIpn9kB11BviWqP+UZ5FEsxI1Pxu851N/uWfP
xyuOmBbrQ99uwLQij5aX1Tw6mtMGdk0S5M7b2q7skjTANLkovhPEl7vpJu9bgqnm
5dbNIcODlnzOjzvP9KuMsyuvmsfztYsB30+qG8IYNho=
`protect END_PROTECTED
