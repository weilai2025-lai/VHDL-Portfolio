`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9J1Meygb2kyNfCAVKxucii3OzLlqGaTNi1YehmEhOPvpdHbNNFuvE+nsdGA1N8I
LI5tO9z8cn52XMAHdJVdJT8LhxJABeX48SiDpjVi0zHsE3yGYQ9Mm5QvExarszI7
Dswp7jve7JoWHdDaQWb9IQdBFFeWS3j2sm0vb9qZa99lHz68hFBIGIYiQDqqeuIw
me31mWArzmNtefcRS9RthexERRXa3F1aUG/LFVsrMWxXt6abAjfjfUfBIni8Zg/6
J//glIuJjap2wQwanElLBdYb0eUR3/rtCNLIN1I6eDjv8Gl5Mpgmg1lVjuWrkEd3
9mg7u/F5oEoKa3ysxAzZENXvn45oc6JcbZZ9eZdN+xdcKnkDaky/jHEWs+n5HYKT
plUb16O8sJLFksJoLjKPSRCZZE0Hwxd1I+Sq19qlSkG8zbmK508usQD+mDKn/+me
1fdjr7r81dXfbPFGUfhZ/JasZomtKTwFVIcWoUEb96Kyclw5C4lve8SRDLOZE9uG
TBEeqHvqttVivOBNPNyT72Vm4ZW5BK7IztCqpYuViJSUjmuAAXJYHb6H+Osq1m44
fHnKbeFpCjgrmUGXuhoiQXgbqHMZBAZLVclK4z3qmWpj3N2yUHxUg3S+pIz8WOGP
ROmU12l57ayrcscqFlvRjK18aegCKu7mDW5t/D8zcgHQQUJAYWIvE3yQiKadbkFg
QIedS8iMgWGrMjUL56i4Lmhk3XWalQZgYdABpM2EeUr301iOMY0mJh37zpPm0kbR
TRaYcS0+LMya5qNBjNWDYlH8F/RqKv5Al6wy/dF1c5dC0Y47Z3Solpn/Ing4RFIi
+1eL6xxsQC5cJnQYwaDXwShiQPjs+rbG4+HUYx9A9G7XNT+GYWzKDhrHiPlm/EgS
rUVNZYNe90qI/dukd/LsPJ3/Hy2XxDWamW+WtEvXrynfWFHeorbOT5VapxVUAbcR
T5AHu8zKLZomUsJr3UQ/+YHc85czAY8TwhLB77yO3EnKU8MBnmroNfrUUINMmQK0
exVm/4cTQlYX61Lqq2EQZCa/x0ceuy6WgQyL5wKA/uj8rhLQnBAHB3hDeMz9Dfk/
KcAYiOmUC0/md9g4gNUbAJsodJllbayZCrLu0z5f3k1AkVOEyRfkwkcNQNW5MXHW
RYiN0THaYsO5tISnWtMMNcUaJNPG2/Mtx7PdGW5pnqng3A/DczTXE8uj8lo9Bj7G
AhLGpgEHA1CPaWlmrPuSQ9nMyLjvIbrtGxdQtLRSefWDwQaAi07SizNfFWAzrCWf
w/t9wdpwwzEMscpHfg57NCUiSY2QcF3gVV/dXJnPhTXJqJWoKwA4VGSTyTK/SbiG
MSyC6LAw8z3rJKIYkW66NKkMwfXH84ZOqhl1IMGC1UpGDt7PlqXqii475ZLfbNoT
ughxkQrbv01koZdLi46wBJcTOq6g9LkYppygKFm+3pUvz4m++AoMvksh7mCbzU5o
+ya9jFK1U9Bi8EnxE39+X6++SyiAZGEgGAwaxKcmPrELcaDQHGCEH6jvSP+q/8nW
NuRLGMZxsZJHtiDj65NWgyxIy2CQATG9bz4acVA8JiNfD4w1J33UbQjxyX5g+e/7
c2fnmT10wW+GqsqOhpYsmdTi0hN1rhjV5PZ7jyitcKDKij+aRxgLVsELA1fNAg6T
eeC8t+f+XpLCCKsHINZqrnV+wDIIayuOmgzN6dxVWBnH9+Li/+/7BoUKpjMmLvWw
jmGUD/IdEt/cZP7CtgSOyL4LMYykU9FttltuYkTSXpZy8t8W9cOsOtaynAXzKBqd
xemQLkiD7Tg7McUHrmlypOKhwZdpzjlAEYS7FTjGkG7f1PLEEMo/2cex4iwXdcpy
WGt5hQpbh1eTWXsi3lDcdw==
`protect END_PROTECTED
