`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zgPfXazZ/aWEiUCkWYxJ7lnCrRyf+yc3d8T7JrCDWSefuH1HGUKsVIh2uBTE/p8E
h4h/rhBDqwpkN9axIsT3aHoLKf8BMLTzIbL3VPVXc3/pOtWsoBGiuYNivsQ7mY29
NuS58KCJ6QUHnoHVQKTxxueOnS+6ImkesPAY9ZmX7LUK/VBPCySouwxpmoVjnGnG
I9x//o6DTo1eeTu44uno9qbCJlU+C4SGVZjvFDCGkot0FnAZ4Xj3HdlKWazm5ZpI
LHinBdkMNSwPJ7Ld9ta8dsdXAB2q3/gFhIJb7l53gESV2zz18H2uyfho+ltLJv+z
nrdi6yDtojDXm9tf4pvvFoUMn08xr/DzV+wJUN/AF6P7nNCyPDhNka9jXHgFjcaR
AtUXS6TzYWGe9qW0OaxraA+adKNgYdAjsGuVQ9Be7fEfRHXD8OKN11s+spL6RlCi
nzare2B95FAvAJ3WbKDPGGdWEZHKlpJfZKpREbdArlhMd2e+AOY4RHWL6Xtn41RL
eaJaihIz51gNW3v0V1+cnXqA2jB2WueTASBdn+u3G7PAMnbfstnghtV1rFhTPtXB
t/V7FN2XqZt/o1irtft/EKAcl9HvUeUpPtI3D89VdVVIPbIZ6W5ypTnLXZomNjFn
QGj3iyastD5vQmPjfr36ZmYcD4jXeD3wTjDVxwMSHJxE3kLM7D5L7YNlsJ4gTwdJ
torc06OHxEsyH0f4jkER+3fpJqN9VELD+jr68P/uvB3F6MsLk5XRvallYxHQlp8W
Ohctdb+KXztjtfcl1QQy1iKJElXl45NAfLRdaErtJ+Vm29F3Spx/hzrWfCsqHr38
lO/WhB4uz6v8HrAi3wD6Z+Dbe4lss0wp3V6BmeNdnX4VaubT7rgv/dqLyKPrSqiA
lP4qJylhB7/RD3f/kKaxTWDCqO+6V0o7/RIUD2rJBBFJfcm86Z0fndoNiOOIjDg0
7SHIjl2bJDT04LM95n8WL0dEBg8kWwVaNboegT2UwfOJlOoKme0JHryhFfUu9TjY
JP+oXrotpPyvvDn5OK9wrlSnjUDPrIHfZialcg0CpKoJgHUXdHKuJ7yKVrJmE+qy
QaG03z9N/BCrtDyF/Q8JxG7qJvhIOVIiRW2eUp2JjE4kbU2KpjkswRxyG/6ddwuD
1CZQCmDO9q/kJiPRxfu8ntp+lUSRnHVgFpJMEIuusmdhaTQO+DMW3NniAm9LgjoE
5IWNFVOPgcnIZGvxrN9+f5lwcWgmjLlLM1GS9HLJ/m8oPy1EBCpO076lTQp1/AuG
Zkg+VcUl70haKyZUOYRs+IBuBMxRE5YS0fZknRs242PViVV1HVESq6acYVsZsTBI
edcQgqY1EapmxOkw9glsUdc/F1OpHQcQBjYlnrOFn+AdPF91QNd/QxW6slSKEssi
8LjnQ8TcR5X1LZf5GpKIushggAYz1nMp9ZbhDBp1E15c9GEoNh50H0+0px4lHgPe
1avpJ8UgX6ZSHNrshNSK937Ds6Rxgwq/rj98CWCrUJUemr+i5VhQu05mkv83GUXt
z2hHLRedNF2XtEcgREMjdrqcv70xFEdyKOqsEDTNEhH51n9PF0YTh41Usc07l95F
3J2LewbenQ1alL32CSQbWzV5MJS3BNZYGSS8914uNmVcI21+NnXooEubeyIn2tJ3
Pvr5pZo6oaiuGCNF02h5Z83kFaZYtsUlxEwzU6xmY6ULXMcxrORjJkPeh/n/4EgU
iBuPkAStCz7axl4kf2mmNTnsBszZ7CPfyJPKcCN4nJsltoMOxwRrh9CzwfquoApS
b0L1QI8V03xHiXRhTtr+SdAkgwBHV5O9466Y4DPjHeEgVpD5BUCcIqEPhhHv0ysd
oQSgHwoMXc+Y/I/aMJPBZK7YHs3qax2Xg7I+MYzZbNkGbK+GhCH98m/2UIkol+Ng
8LcsSRCcF1Ubw01qA01PEn0WnX26r/TSFc81/Vf+d33j5nbcBEb9PeizBhurFOAu
GhkPO0A9g9zQMwkOLMAdqkHeMU2QcjVAOWkYRg0f5gtk2P92S8f824jMFPlgsbuh
NEHMJIjoC4CbhXQ4v+Oe7R4y2X6atam/rGi/7YK4uR23t40ER0bR9AKyEq3R48W0
+w6FCBV5O4Z4xWqD5b9pICJKOECBvIGiwyIAtdyTyqpmCxDqOgj05MVHLZ86WN2F
gAXGDLrzc7gkBntExEucMS73+qpkrnFTsAMXQeydx5/Texmqu2UDLRbzhQf/bCum
krvTZrUQVxmQaIrifs4Dom2Z+S9j5FV6fTEo9Zg1YEY7eoS7NUdQVI4pGtnDd1yd
HieWedcz3mP7sqM4kNFlOMdjr2bbK3KO+jd3O1+YxEq0f0fXMXb9a97TugFuFSNk
/YhZSHigTCk5q/oYHc7+WFlzmLLycopLYdMx7wgIaVVNAHIUvb8rU1WUH8KU5pOY
kjka6mTiFh3y6ZQ2ABIOpc2ByoWmSQ8Lt4LRF+eSVyG3nWB1JsS5bQ5Ym/pSPIL5
68zaUWcNL71AtODjpAVuohsVZsfOliU6m02PVYX9QK+n4HXiliZf1abg6Oz7A1O0
6Alxx6/xcFDQuq67lyw97zYlO3zn+Tp0vJAbvknJ6IcgWWQ10fVQGiGmP8vbxd1X
KElVmrrKzgAJBTlUYt+mnRzIU7oydQ11a/LhtgeJgTEQ/6DQ4gUv7ayvjxt8sCLY
6sNq6l9YtYkoviVXr5372gZkT4fECY4LnvS9eYVzWn/F47kOd2xMy3f0FFO4dcJD
NVX3Nam/jzhEIRAxclbxqiRTGwrZxF+SbTX3npjSJrzQ+ZMrdpLvFdYHoThwI9aF
oSVkf5GYlOTgB28wLkEQvxMXJEzKy9KaktVtTb5QVbkoZNmwmwRm60bPBjo6gUNZ
LOUc66f5IglIuK1OwVX0lT1DrsDg4f+0lsEzHf+2lmLCEyGJqCC9fQs4jHdpCfdB
lfAJIuRQm4LCBbkCEbWxcErqjoLWg681P8ff/SDvS2oa1aK9cuxeN95JJcmlE35n
P5+soxb0TcXCJhVv7bywGPZBdXfM1RNdmLa+vF56pqa2I2wwv4dVbt5gJGbGVuXU
RrZ+62MswG8Wi0cSw+XZg9GNOEYmZdSsQ+F0itp7PJfpqErV4JB5J1ivFKFVHuIn
FkbiE/cO42MbysqirnpcYkhM/56LAg+Wv/roIw/3Zzj6WxKSR2dmpuDgjS3tcu/Q
ctGArFaQeDB1tFSCjFOLavcReD1jJeWBvbO3iEB4GhNunD4gdnLia4S028rZp+uR
i5oSeovtd6vRaOKfwznputvCIwgN+NgU2CsuUeDMWktzd8y/KR0EA8KxBpt6BthK
85X82YGYB5htN9NkSK5PBqgd8L9pIAodKVostAg/6J+lw6ymnWFwsAuG3DyKGkkE
VsqNBZaVFEjMzM8MXQZhvARY97c49D7JHpZg/93wB+Pem99Zq9RovAUBFDfVj66Q
TKdawSiMoPuxuGnZ3wi7bcn/7PIu/+PO7QEe+HTwIjTJZ3lRShMufjlUnHJEiWJb
yRHRowjPTIL7+n2O5Lgm+q9JpHtFbY52VYHdIpy0ybXndVXASmLirfVuKPLWsDDa
bdhzcVVox+q9lX0ESZPVdnPRrsRwLCU34ST4mHKMCf+DwpazCyQUngZT2jIdSAbh
rZiNG/drY/NjqHx7gSZ+p4JdD6FWPGLThsTGZeEAPgCOjOY1R26H6eKpncIGqp3X
mIxQWbYT90uRPAsu45hs8Vr6lw2W+MVvNO+/n5x0EYzeDvvWvsqR9idb7fQ11cWL
Gtp7USHKD+CmsKNOTncoffqPcH6avcOg4mCyyyMlhEb0bXvU1QPxvsesqmJmpKPx
h6fEFG1XsJM2YRlE8FveXRya6F7RFjSb4TwSc3g5BtTEL4QmPHDxUf8s8BTDFOea
zU9IPsq5FxPiaRLV+X38jsS6vDRGHlBf6+0Ifddl4EBY0f+PhdPtaBF1YEj2iZ6Z
VU3PcW7QId8PtG5LT4+cd82Q+pnmHlQ3N6zxlmLibW4TpG9VtIoH/6j5OEO3crk9
uEX/z3xA10e/3uvrZLrlDfjl89SoyTMnpsOfobwu8ck5Z+i/A8OfZLn3qozhmGsZ
s3kNMQhCXqWL0CnJJOwxGigkpmir+TpAU/Cimnxs5jCXdz9J0gJYOQ7xXcowm/lf
4YvgDTAcPv0Xx7c52HsKht6yFvqT/eRz5P+NUV1yqma2e/9cqWvfKGYIAMgD+E7i
isd3puD94bnoyyyJAyANEihJPYYgcopmeupHZHzQBrIQaYjbezWPbtteSHL+uOEX
/lZHJk3ZafBsUGK5ythyNA0BPpH2EkuAJ4Y+ZFAnHXmfvVQf/SdvU/g5+bhEic2j
5Ruj/WJPlvaAVZlfqsMdP5TZMVRVbHoxHNWX+7uN8yWsAFO9UIucKYZKz31UvuPl
qzY/j1rhPkcgKR+9if/z8NcWW3gsd7UYkywsK2h8Cwg=
`protect END_PROTECTED
