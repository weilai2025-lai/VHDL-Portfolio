`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/Lsl0t6msI9nO3vv1a9P0FtbeWYascfpQiNqZIZ1Wp4CagOfDoBXuV7W/qqERnt
badCgbnVMN3+W8eFOOq/4psoKlbm1DtfzYVwmWbGkdnyJtTDg6pLz2FkA7+ys23o
Vf3Ul+n5ljeASAd8N2jVV6JCeS4yoOtVikE9G4lUph7QPTBBDq3JwqRLvPdpvWBl
NUUNXHuv+OMG6tibQkAh1OGASWMcrRU9qeH8MO3nHMCp5kqUp7bIlXSX2b5pP0It
GMmxEhSAMfF9d+1JZfc8L6JP6KW3IAepvFKpMsLKpF0td8X4FVpciBhiaSErteXQ
AZi3CqJCLW0ug4mtK4RORC7V5k79il+fSKjXZAyKQKmkQHB8uSVAWRwWQU4aORlY
UOTiY2LoAa1JzIKFABm6fYjMpXaLlkADiqATt7sqm7Tz2ZJ1UWiDXDLNaCesOdTW
XMGin3wcAZWcwkx+4Ykn6af9DRbT+wPBgF4vepBfsVbrdzIblgHneaUNyZRtn+4Y
Y1UOIJ4sas3e3tyPcngEnYwSL90HTnHarj/LqXJTP27RPVS7BwNb+EftD/bL2kaQ
wrknN2KMpqthG0noboDMtZrgS8UeEGFCL5NycPlxQ8cnglwnIk7GOUxXWqapgmSk
5gPyM/J7t3szrpK7kCKx2M8Ob82mJajTGHD0eYiiXUq7zqBc1qgluozKSHvsInHk
`protect END_PROTECTED
