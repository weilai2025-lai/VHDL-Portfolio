`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUu85tWpKtHhDivuX/3S8zzqJaYBAAg1KhOwgNTMH3TdV7QDMifvu3ZGar89wucN
PC3wwT9L4WDTdcO2MG7kZMB2Ka9rHSuLRMcSXvMRuPiWEefxl6u0kAL+gDrWs/65
/Tgg+/dAXBg2KjBtjze+kaqtSbEpBXygJLnlOTk141ffoH5NyHCDNngtVYvwsETB
p6/wLjFfGg4wAKGoOXusWCZgpMXN+m36PojbS7Fji9CX9g6ZvJ8fpYucZlBk7BuR
Q2GqAZfK/TRD4ZYtNGd650VocfW8xGs+gVXc+iJWK+tQWposnfapf4lU4KpSQdmA
+MrMhy0ue2cbZSMtik+Hti4549pPIZJWqIAdNhL3NoLbyyeEH0sY4KMFK3/orT2l
78G8FIwMoOonQkk/aMUDGPFEih3SFOGmMNwg8IWDh3oGlacxjzN+mLPt1dnNfGrI
rglz4TVB9KKdfxIlvhWAyLQA8zmXWNeq+os+3grDttQXC/ChyJCDlGdPblb+4fUA
mSqre86L2tGFempeKALUwnEnrTCXP118YK2OIrbDHdkKeb4RG+DH0u6hIXkEQHAt
7YjRWO1h5KXmPP9290eeXFd+IX3y73wVMzcauyo0se96Np3oTaCoiOecejqlIZkn
hHIGYiQ7CEQxvSlRBWLQTv+K/Kn1j3uT9qwWzLPiQnBOrXcgYhzffaOvAVkKMUQy
x19d7JOMg1fu1Mz4d5D6IQMamh/bMYPCIB4PjxslJtl5M6w54lN0fD7Z30gsZ29c
jlGQ8SSUWx44C3gaDD0JcBKPAWdWAntrU3qnhhLRddoUYkrjRpLRJHMKPtoZJNWM
WpVDSsv2gKqMsW2+mv8J26E4/uerrdngFUsfiAPDJODBhrd1B0djHfU/KrLZftKT
3OCKKxXZS7RQlv4Wt4U9UCJqVrJ4cqVdJTUgv6zecYDb+WubBjODhiQDnRu0Adxl
x535Ah1WQ2CUBGfAyBnMk2E0b9a7KhO3qSIGgydt2lF2no2yXV9Ya0ZsV0uRMSXv
JOzJ77CNr6MtUd9GCKNmvbttMxfvAI1llbrnfWgUCTTN2uvQwAajfEQ5/zkVPAEp
qaTw6xNprGa9l0HLHxNyPkxlqBl/J0971d9D9eTKoDm83WFGyJzA4XlUjkVFsdJA
qee5rSM2LkBO/O4GbVoYHfcbMIAOnhONhpsGavoyRvHg0462vB4S2p8YrCBKehCi
NEJpcvMRvfLpTSHiQ8dGZSzzaW4zzC0BmylLOJBBaFEVvnALQc41zkMraE7wEdlK
0JMSQ/DKwlj8OkgOdR6Ob6fRtXyduAO/fqywNiNWi5wTiPUK9kIgyKF7YTfT9DQu
7Xm+2PswqoOuoNUZhllWO2HaRYjMXDQZLsZ7jKfwFz1o6u/NX/8Fp2IKe5H7HxXy
VTum3zznT+mt+tbDMIX8iFFctalu8dPQsa0LWofniqQHDqcwHJ8lI7K0XjcFEHOe
It3Jy0q4pAlS3+RtfjQRwsjbi9ftDg4GmfxygtSrrTE0d1K37Kvbe1UFf8hTYM/1
25mpmvJEGgJ18TfFWhK0lzYSL9BpZZP9YkmCb9IuWZrTavJuNsHe4FZeSxbCB1sS
WhEKeyqTwfJ6KD4De5Th81fAToe126gZQbqzPY8dWr6n595se6bRWL2sQbMOWjeR
fbTTuE2rttWqQkVT3OPt36NVpp42TgdUvq5EnVLgrsIfA7LP8opUiiDIVpP5OntO
ZyJUpsfORJ1Qm+RjIxSYgvG/qIa4d/VwBZk3cV1K+Yhf80tTLcEohiO6LQcgFbSm
yt88raLfSU4rHkBv+o7fYpWvtjVIRpwEosfYSBoKZSF8nPn/iOTIhKJFUhxHujWE
erv/zokrR8Ez64UG0rQdLw==
`protect END_PROTECTED
