`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pnrzZydEXA1NTz8wD0wE/2dcoj9ozB2R0O0WRLyoZDElDjhCwh4QMrpeI3qkpp6s
TkM9IesoOApOyDzkIr7TFi2AfQQNHzEIDICp5UVfTfjIe84Hu4g9EDIQ9cZFGu9K
rXGAJDafhrF0aax/vKNnsz8A5GnC1dDb1LCGsjL43oI1FPfoBwymj2cXBn6yMS0p
8JDG+Tk6vzAKxtuDjJnlxY0huonZCa5jYiz8FdDfeT92VVc3T7mvz5lcCBAjDmv0
PNWHbO6qHSialywBhAtjzfmE/2k4oVR/sCwgv/bfwLzt5GqZTaMq+4k3Os1Dq9tb
os8sx8AgRSpOowNhZL7ijWitw2FLJ47mzFAa97T//PRQWNc7B+vDld0YZdUrvsEU
xqH/lkOs/i3VTq918FCBHVmDXw14O/osi77MZ039DwtD8EBcGBZhOeJPKeWGY2Bt
FSWB/QQNohoN9uqb2Irk40udY9KfBxxu3Cbza7O5kpLj+43M7tU7Wf0EUVgo1Oc/
0rZrB3EJLd8OsNY1OoOz6IX6+MAen9vfxhe/7M3egeFVnMxwoSB2cLWsond6WIBg
ym95ROgaEjK7sEZcubYArCd8hRUpPVGEnCDUH5LAB1ld+dLk2vs+qGeaPmWHi/mF
Bevi5t4EBw/TCWUXv59cnwUFofHo71Rlbu3p5CNIThj185Mfl8oST7nkgXB1h1zv
J1EM5Xfn96jbZdrB4EAP+3+vmrgIsxP9GLPa2TI4NdmpbdE2VM0spEe7awAk1GVy
olgPunfIc606HZ3lCdhxfMruLVc0bKE7GryJc3c3QbAeQEMcPvhUpQpYN8u8/m0Q
UFVi1RB3Tty+NW1WKgKRelFd4gGq6kuCi8Fzvabqlyv8+QjiZbwNE0G7V6SYByXz
2g2A5lPNRuD8R27FdQzrPwQirAvSxA0uee7b4uUloOORv3ArDe56c02RuQjtMjJT
E17aMq6rhMkMqqTb/t7M7cXXzCWlZUZWsmoyITiz75mzDwMt95E8T3cEBa9q/WqF
jnkccD6GtX4NA9QQcbm/C9KPGjYplLg1P4qlgzH8REKPWom+02SKOed7wh4eFdt1
SRDeTIFgQf/bl17LvNOqgtmonJkyKUWoQJTl9iCwKHb4jgQek3UGjK3tDYOGo49z
+g5WC0vcPaQuSHNnHjDh4/AJIiFUAqQHgDEMccDTSdRN0AOfOtgeb0QtgkkPXDbA
l9KtO121MUSTCaHtUo9WXAsDVyz5cHFlqt1661/QwmFR8pTvMTxA3Pa5YUpicRjE
eBV4gffx09uaJhTsoEmHUEzebiegnqQHxbNtPyQ2UaefTeSEyIYlmeM/NNxDvdfn
SjllbJSa3p9XWm2i6LqUQcH47hxmuedMGiV10x0zoxHe4foYStdA8KC/7/zKCX1B
xeP6FNjiYaRVLJnxLPjfS/Vc7GWh3iogduy3CYacLpgc1wL/EooIuOEVB4XWxW9J
QWATx9CSv6Tz8WIvJYwp444SW71t0VmKpiTAX01hN5jXQGARr0RtZN+8t/Ibz++F
v3oi7q15PyHj7EHqZoveZApcFsWiJHK8/Z+2zaTTZNqPlZVs/BsSfKh5/K3LhpWX
b8Todshq1ZTOu0ElyO2rpRABIRPABBf+Z6BWEfRzoym3mqFqjs5iWMljruFjs6KS
RMA0EYiZjW8nqWgmNS6FMvoigwjWtUgENxgnoiEK1akHFSC7EyENRNQmv5U64Np3
fTAKLG1UNOLdKu5e9eV/Qq3+VvRnXjk2v4AcNqucxgeXalF1zJZFd3YPtJZlzDUa
156KDA+mhgNi5Z+rdSVELJYEd+Q4dfI7hpLWtmHYq3QexdlglTjFhDiZ2fLmruiS
hGnqsg+Ft5QX0JAedudVBPRBjj7fpbpZFSVvPwelQ5+fRhD91DsE88kCnPUukQdD
Taoar9pKw8s9rErMAbOfH5ucgxldoxe9UQpO3dRSpL4RZ9+yc0pmWXpAAKhbDWMV
f4w+IznnaeD/0yYp/amm28Bj4KU/SSKC+HJBCNMqfMGw2kr86IdpynSGU961IXYE
l7wDXd/aT6lPFPyXA1nxU2MttyFmJm+FEyxdbqSuBlFEEUncOlPpX+ROd4PqVuG2
NCLeJjUBopS4x1Eh0JU2SoVfQXg+1IuZF3wK5Wlrvh1HmqLW0UXUGNG3gDeLh8jr
QDTOi1OPe3H54DL49p3nXBiWd2bSeKKsngEvNc6vaFecXfA4WFPnBbWOEOiBGsIS
7PGjsQWqnVg7nUjKg/I8IrdeS2+v28FbUeqPLs+dwaS4Eaug/uBAfN2BYQLT+VXu
imA5bHSWjKU5LCatC0oMVpdeQBBgGXdZIWBYBhr3ExHIsTDeROyaiiJqHhsHJTx8
mT1H7s3iQjwE80s+YcRDGV71bd/Az8C0sG6anDtxaBctWOAj0cUCNMe/B0IzHeuy
VrXReOLMrt1k6EisABFFjGhIUlnZr6GJIvwe7qazWLvmbFW35QgpK7PffsbVwxrd
dRaJEZXFz72yDyAESUxH5EZ1etGBa7yyisX0XVM2g6PipxNIOVZDDQCfwijIdSCi
YCn4lezDDBeqzqtgtZZUJdrZ/f/0eIvNnnL9u4248RpwQ0j40SKLI+RmednVG5Uo
SaxWRJ42FkDU9RQRkagljhi50UcoExwWd3JYvhdixSjx1MzH2zzPBD7kXVwIvi1Z
N/Ag1itl8e1tyhEEw17ZhoGOCSorW0Oz4ujYa+iXQyOT4UMNXOOucO8g/fb215kK
tNqcCr+1MVh37zcEsD1QkLeE/BvmG2e92zppRrw8jqrLiHUiWzs8YHD4bITBE1Qu
WPyGU7BdeWwnhpylx0N+UApOZQ4hqZJ3J04dyXElNpV7j8gDMx2N9wcy4hm68HC6
BRD61jaXxtjj/l0AYRtPRNENlpHnvJMiBdn/J1HNfd26ReAlV4zRemI/IJPNzD4w
yTZbsBauFb/ZMAja4T1iOK5cRQcWPfIIusn0ZQqokKOTDFcUshkRYd8R5iZ3+kI8
XHBfKDnOttqi1bjPi3AkoNt2CNx4G6zFEuyOVexlRhiwPHPVOWFoXFuHYD3CefkH
nr9f85/tSApI8PEYBDUcbm78IxPONXcBUd1t7+LrwP+y0anPzC4z9+Vzig1gdH1G
45oCinV7M7vPQyzwg8gxLrYbojZRm2xNC83kv/epziW40qORL0G7AGZIYyXN09UR
GpcB6pSbp7ym7yi309KwYQB6BIi7/I0YNP4zwJMkXirGV14C6qiHnDIM4dKWZu+s
Dacrd6SyAT674eCBH1xv3NXp/huqcOhX5oU2KqaOAbhumE/RxZz8jKtJ/3GI3JOV
rHKZRlqVCy40OzKiM2hszgYC9UCPSHWAtnBQMMOVSc/dURIv/bWXIiKXzv/OjNCA
1G05JZ+M9P2JvR8VnWLLlbjUGSFpGPFjH0maOFTRAw5wexMQAokXNKpFlIjF50JJ
iiQc8ayr0B4fXGSaAGRqZ7ezeHh+DFFe7KrpFRrxnxZZryKtysV1E4yQEhCj1rc1
/ayXVuCM3ZmCSQ7wfo1pwhUy4heyY54DHJ/ao8QTIqe+ZumOCJZETrYff6aZVSD0
7vRqoC8dETQqsai5cUjwEeuXO3gUm4KQPnSB5iGuy97lTrzQYAAMfWMBKd5G+AXj
XM1aFMLvLjQcm0bPVPffDsMAqCbFPQe++tO/trHPSCcS+WqX0M1mkFBn/5bOHWp5
aFZmlx0h2Nah7wJLT+JMEiE/LTexp5uZYo+F1lIYNbYlJaujhSrZknYi4x7RpZ/0
HIy/quLcft18T058KTyiWMy+80xUV62gvofZTaieiSqU2+V4C8RfhXvc4PUf1pf8
yXlYq0C2lw775M32fzRv696xYThkIusTGfqKkmXkBZK+EeX+wRs+DfW/K9IQtNTr
TLO/iPdxM7Ltlx+/hTD7G/XPhzWlHeyXWvgHEa1HlAQ50NzQNLOxp3K4ULgR6Rkx
kcqbWzW/JeBtI2sBJFpNXa7HTSBvbl2Anx37mih9/zu6/KqmufRFuZAHLA3xOoNy
BLhsdzK1y3HGpuEDpBvdb8YrmwQlDDFatsXq/vedaRJGfMRxgyag/ycyEHMEse0g
8JgJ7Em9mbSiQuKzTtXm/3OBzL0iOLnAqj+1E3ig0h/Z5HvdlluOr3pS4FCxS8JS
/j9+3Y/1dFOUHtc3bXdoAQ+uMNMhgzXfG1u6dRdhZnAYC2GmJVnU3D3pdpErcpVU
4Hl5ZgzBIH1dzU9u8Ne1kPfrz/Kmc2MuCg6CmKaFKygHIxhF2bgoGp6Bvvtmqzvu
2E3j/ZM96moB07adzOjUtjRQ8hDWhEMZZ9bDm4JAjmZLcPE5mO+3wAjAV9wywKWy
TRrxWZcQVSSxskqXgl4rMEwQT/hItxUON6QkORba7oHQLrROC1GwmXcv1+Zk+evu
SKn+ReTmgyjosI/fIUm9fJEpdiWV3kUunYI0C8SbezcgFF8QbMgdnE2LjThX7UrD
68YV60h8YsfVqxX2lngYPUK0UVAtXVCOoPFU7OSqaeJjW62Q1tfTbzFF6tOP/f/e
frZ8OxuVlALmlWBhF1zhO2gJgettSmx2Z5duMkfDLdLBOl25ETcqrXOoGZD81Kv6
WfDSbvEWTh8KP2jDWB196sf9a9t0BsarqvAM1PTSqyTIPHNYcPmyre0htjrpg+Bj
LEUrPHKkvrzzSlGRUAOxevMR+z+dvbni7PUoJKkdkf9QsaE6hHOPHsO41gNQgtdZ
qeXC1EAhM1myB89RLyR8hC11ndE4vEOCU8tn1LLEIt4nod8UdOYp9Z1A/2LYlMBg
i+Yga1QkfAsJjk4sG5Rf/7DdXW7H9Tie1kbm9D2mqIZmi8UTkmYlKfdUTRDnh3ms
/iaWlpiTZdqmGnZTh0dJwa3hI6WXMU7LSzT+6bfWJZazvYCgFQ8TUlpJegvm+WwF
CtwC0BG7tB1g4q223gmJMaKFBoUfBYI7DFoAqFoRsyFbMuxMFDD4SW3YopMlF6f9
C77MWQKroLm1kjrVbTLkg6naZWvG6WMvFzqZj6y5jx3SN4501jyuWIFn/QDqxL78
q18biDwxZxxCjXc2p4YD89Ou4Sb3G+GuJ+4MAwjFAI7Krdn4d4uBhGmlPYaAljJd
noaXBrcqdlr4p8fFiPdNXG2j6cWCoEpiFYO9msnjN5kCcDCyKMCiNckrjv7sB8lj
oCYrjyTC7uqV+BuMvV/z9Gvd0M0iJ4vYBVYYVqzBZGJtCqYymT1mW3aK4HFWOy1y
F1+eL0oFo12+FE0OKU0p+trOsPdZXefNtcM6vLIiNHPJ+B9WlTMCcTwzOCkqY1hJ
vp+j7NOJOlx2vlPIkrpixySaOg4EiDXnuFY/mniwFfPT616W7Qpjidh/HpByz8NS
PAVhfwNqfTNfh8KmpsVi21hzM3R6sjwa4MEYtKkwD5ZDlu2yXjFndSEim7JbKsml
F5749hPumGwiKevYG5YUDgXJWjN0JtzdP6B6C1z48gPQZGUpvbC/9lJlI4K4OQ+R
vEimbgQTGs+BWtijZItcp7SmtbNY+Sc0oHt7gUdSm32awxlcofDNI23QYdW+phYr
6ij6cYl6wdfsJ+zx7XBx05Mlj/UHO8YLBE7DTKqT+igWKiM5u3AykiYXu9NyYTCv
9NQ6UtyhkwF6l7MRnBTk1YyhoWAaPFuGC1L5NYYizsrPQaGVP63eKFldQH9I4/78
lS5WhiUu6k+o/8NMtO2zqs/YcSlX9mUDahg8GySU++TTW3vyJLEMteqg/ovXHFYT
cCjNWpGcVMzXrH0hxr2Vp6nB5DyWl2XceKvSNL/I8YuGieEspQqrA3+uMSILzgxP
alb+yPwfFre8RhzC2HDxLnC3O3z/KU1PJ7lPIStpnAiNOn1O7Af/dr1IrOAZp3wv
338E6Goe4Kwyg4rWHAaPlrQabbGMQY6pN072k0uPLQZYV4idAIAt6kqSnRoAGODi
3yJRihPunAosalVnPMX/Q4TGc8UmxhdApBjkGbeM9m2glTWsrUVEHL1u/0DIJs6V
ZGqO8+oSiEkXfi2SnCp+mWG3ZA9vr3T/ZcS4W/RuCHN77F1l2YgCEpi/+w+AqMY4
F0y/ELEJkceBvz516cRfidnGA/FyeOJk4LdcB1DRbQNsSkHqo7po2TrK5oBzxAd3
D1lu8BRjNWRPYOVvuTZ7KUlQd/cgfnzaVZvG+0zMglDJz/Arp5QgrSQD2O5sGIt8
EzVd5Wsz24Hp1ixOStIRhFC9tgVy1PEcvavHFluokqmo/Y9RNxrTorqdYfsJPs4s
IXlhMUZYaLiuRMzCM72fPH7V+XUWoNM3oY1mQ6lmSmyZBmnurJufzYVxnF0eQM26
dUzkV9elX/DNka1StZGtXs4GfXYlLvIuo4/j5qi08Hk+BBj30Jbp+krE/8y9UsPX
cqzSo1U4hOGudtfqr9pNnBnK59FN5/+VtpNSqDA9s2LAr34wG0Q6ze9TX4PN+bSz
+LqAEXm8olFEsvw6MXgJ6+9FY/flHqaPI052Snd31fkl9tYBrlsHHUtBtoU2MMgp
aned02Xfd+fxdAwuQI+iHUmkDEordk485oM+IAfuU4kOGEamamdLobgwIyHpHlJc
uJ3wUE2CTRsXVzqQcyzUhKpK5WPI5bl1IRRsaDq0JaJMI5FED69hdynW1PI/7ZU3
CeRzS6+Gt2n5GqtUcrqbHXhKMhFzlNl0K7ocrOpIXB7zNPZ8Vkp5f0dFYTs/Peqw
72Fwv4h5E+qLYegDMaYgyHoq4MDnu4/zBvrkj387VjPu66SMAGsr9/OxYSDY9Cwo
NoiYf6e1DSUPwq7SWQhQ+quz8qeVMH+Z/f/V2DCjpAnzunX/jIJmB3wohFjKx7Zn
`protect END_PROTECTED
