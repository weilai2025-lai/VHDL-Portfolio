`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ruRu4JKKYIU0cl3ajnVSVJ9qVsjoVK7kcY5ptCwrrCs5anpKii8AWbwQEmLB6Mf
W1iuA9FaZhHi9B7FqWmcCuxEDaGT9OWnIx3VGw2lrIFjefe8tuSJTvikWYfK19N9
gbDjD2qZISY+BJkjw7f2i4i8tbIByLeI9Q7gVzq/QttFRAJ0+YhMV9iixvLLrSt1
moBgeyxc1uT0cEI3MogXSfGxUAnHZNNLmIJBTP55Iq4U8o6Jkv+YCwDaB6fwkoFD
an7qkmQhP+Jw6+D7ogNHGTaVv4Ax1J8QZCnHwFFPJEvAhvwSzoTgly7ax2KEYQs2
JlafW3roXWY/dBE8XoTaG6CVsVQuBO+26SmV3LkQHeKjhH2BWYsyj3v5oUV71UFZ
17iGCJlGXZMgGBkdPi/rg11/3f/PslPOMJxBT4dMu2GlN38fIiLfeUzIuLkDjWD/
dwWg6Yb8ColrI5+bxKY59hNkTktgfRPYNmscNOXLj7ZMf/30jDUvX/Fr17Oviya+
nJrx2XpzU5Yflv6ELV9S+xHOkTMZvOdCLaBi8bMIkSyeXFoIabvAgevwtu4Y1Utl
4GcRs1EmPhyb/YXx2Vxve15CSQYsbzD6j6jhgjXGmjWh6Rq2by0I9d8Gt+GIYZly
BdDYrRmysWkoi/41CTJz7PYTLC8zw8f/LpmD9soLm8b93+it/8uSnBcK/tKjS5LL
bWJhZ4+nUsdoied4dMI/pjWU+gESqchKnS1s6Hg9SkAUXPCpkzc7zHjOEahNMS8o
x5n1mAGc4MJcWyheXuvMWCy64rh2BKCYFDFNnXnNc0+t4wQ2nNoKSibWg9Mlvp9m
Drl3EAEKWlBh5W4z6u2FDNdfq5FG7ZP3yvsNSLb/E41vCnP1bdpWYhfvbB62Wksc
SBkM+k/7SKO3h1tLC0u3HgKwdcO47muIEVi6ddojimjzBGa70WLJsOyxbb60/1qx
Eg5oVea53rS108hDShs447niiBH4aAPx0j0NCNoMtG/cSxkmkEbngp2GQogCAfEz
bmviCmRJfUnZJ2FUf32yR76TI+FBvFMHLlDnmSgdVWETAb+asLism40PrvQmUPc+
wAnSBcpV8ozkqvM/WYH5UYamCYFqqku4wXFJgKEfhDttFAV1g14Hjh4D44zWtsGM
97zuu2Cr535FE0ZNpBS8c1uUbFPFqgD4JZP6zHPfHAR5YbESHuzYYXqRIT17Q5PD
Mo4OwWFKY7/P7jSRH1K/VqYXNlQMbFEYM/Fq9BrEAZiQ838pfNwYCPGTuolibuy2
KnvRwN2wnQHFapHIAdaEg2QoD25Cop47YH8V6vSN1T6LouWvB9W5ZIWA20lxjV+W
uCQxZ97pOyqCD7SYVZNdJ+yeCMQXNQDH7CXvVpHAHxWJRSrNs0nzceooRLkbMm55
MrVYChhJshAA+jIzzzsBV0lfbwx9EulnjBOy2ED6qVVclugO/yKPYbPMKo5X79tF
Fym/Q4Jwz2JGnZC+9bXy+PmKwIF9YbaJoL8iawrJm0mVMljZZ1EKevFWlEexYkWZ
nDpber8XEvehWI6GpKW6sSUSbYr9MFKv6AmT9cLysDnGsj+o/08bmDXawkTdwmn5
S2CvuVNiigRx9ZRNqXZeKbpYfmcGiS63tvOrz+esHqUoEkL1rFroacWJHeWgCXa4
IvXUbnhHfUcFyI39L9VQrMnYvi9rR8cN9kW8o9K2XBiGCVPaGAdLB/CAzWY18Vqt
5RIJEYZhDzUoveLisGfGnfy7B5IuktQFf0O9hB/BWe/pjQjhdrTXU7rLQuCtwxKy
xKT1OOTDqpbUn2HSPuZG/MH5d5MgjjX0A5nEQxSiexBZrEQGzQ/uUIZ36tl4m/eI
bsw63m6FFu3tWTrzm1jTzBiFQodXloBf+BUX3MJ0Go2dldY2cWFqw+CTLcncg+Ja
2daivwoKCpWglzB9Lp8yR+MoLsML+q8Xm/bcJsY1HvafC49nr88igjlsIUxba46X
DqozRqTL84dZ0NulJuSaLPuoEk3me+EMRoSAVmF2akTmB7apFOjK/vsQQW7stFyX
GVx5KZbJRxcf1/8SiclkwOxnR8PeWlGT7FFLYwW67q2tTDX/bf0E+hDG61mzx7O5
s1G2nBc46JFngZYr0wIqGIN+3+1a8V2dG2dMIkbrtI1UdQ4sTtl6Rp1+uXJCXslz
CpOPT6Yyrrmbt96vSqOZ2MkNs5rLi4JHM41UEG4Q2IQCWDghW4q/QNsy3SIicQeo
527btdfyXOhMHWo0mq9aeBR+RuLEjsrqpmQqrPI9hKhklzRpRFhlnnWhsjX0ESeI
JT4HNx5nQJrW+HAO+PreHc7Qttv3af5LVLN8thDyKF8K7kLBnZHbFZPFLwYDK/KA
cHJs3o5qRZvXdljts5TwaPEitXLia2XNkx2OAwmQGknDZi16A1+YBR3O4S7unI+G
g+5NloOTiw4nriUAc1ZsHA/xIEABnpjFGtPnAhAqP1WER7Il+uj+lrqn1PCeDHPy
cdxsR+BRi3t1clszmP7mV6ZF29uzEuTkjOU8Nwl/GSAXk4TKFlvKxp2gI4s4qEcA
gjzraG9Ku5Q9RKtlnHmSekPRDfjPmjgvBdpbBgmwWmg8bTT2Q7qOihETknmWZArv
de9JGw1z9oZRMY/seBZr/VCtt+mMRevbLITT1amGgz1veTIlZbUrHl4J5YejYmlR
usOGLqcQQqvoAG+QDPhLBOBLlN6NgQZ7DXlx/bEmXJRF7oo1+uJ0wZVJGrXvQWpY
a5l0pSyMD4MaKKN1rmB4dnOhiMFZhA5RKz9YECsJX20XdBJ0HBs/OglejHajWFrR
tAg7Yp5WmdKcffq/96MNE2vp/HuvqzzINDuImCZAEhCmyxI/zlt5D7zAXufgAq27
DxEZVZ/ILAW2yUdKozbKA3L05hRUSIm6Qs6RKtugbfinoUiCOqynmmd/uLAzyJcI
PZfB9Sypll90j8fXAkprKKEjX6DZ8GxJgZ1Nscl8W+AxpUSs1vWNmjv/HNcf/6M5
CRRapZ7eRS1HB99iVpxUBbDvNnb6pWFDgTnK6UUPpj3kUIq4QPH2N4i0fD1VlL0S
2jxsh4WGG+j0o9AYbrzKQIPkVytL+mAjNuc3On7GL2vuaQ/VVAcIyY+H33fWx5zw
U7RX2qCX8+VDcT/0mxK8spOelrg4udgwrFXPGMzIAz+0OREH21qvrCibjIAjP4Zh
+ZOazCBoEMPNCjtYWP10aZaqyMYN8lwLb2LV+yPXadDMnqIXeIAalFgI3kygPAjo
7sxNsYwznGv1q1OjjR5X5t+VGdPfqrUTuUmn+q7jfw3VhBBakgBYtslpLsmUpo1S
/UV7chF7PCpowzEP3ffmcEHS+ZmsYeuTxCR/yjeMuQ0SorIdTUegmbNfrMAdT8Zg
ahZLMcenHDKrb7HWg3oNfWzFwYO1IGrgkOuUg3uuF/zq4BIkHDzT9PRzCQXdCMJ1
Uxo5dkzfprW2qmjMyHjKRh8n/jkByz8WsygHbO7rrGOAXwEcsieSThmTQJSvFCwd
rZ41qhMbM+R5tyChuYKRtkMgg5B3kk4uIx+zvdy1sAp3fEUvuucsCpGGT1NpIlbQ
GEl6n0qBhyEtis+YxT2/+fJQlls4nSBi0Zf2AGoFmklfRGZSZgUF+aWRGO/sO4zB
rLEdBOhIU4OD47w4ayqmZWOiOQ93dvnJbJrCS3CcRImMScPTSipztFw4qpqnQ+Ne
BxmFKTMMGMN+KmQiDgLNrMqrdxJLDfrrrN8Hy7oFz1q7pA15fXsrOVaeZW4hgUmV
fcQP/V426hM19MxsbeBKcd07Eb5GByREksz0/YGUCRC3LfzuzUcjucJl3Z5uyLAx
9sLhT/iixl5NLwkclH6VBQIx1ubXwGARUdxAkYBmOXWAT1rTdzJPJ2HqfSeVjvSo
Wlz5ws0YXv8mZkIdFrmScNkZGVmPc6So/eni1E9TtnxIBwz0Q7vt31NMNVuJ/ev+
8vRs+7JGWNQRSewTh6qF+bzQYAGq5fuYays5bAtwuIE+jKnC0D8J0nV5hmLsqm7U
IKF/WmHr75fZSNmsAqouTGufu10xAf/pZ/+u1rIj7ne6xuwxsZNPKMJLZ05+uI5m
WzuRBgbGF3FUSGcLJoHLCEqSkfIoG4nadYJ8FrJb0v+CJltsX5k1q2d9ovDVcVSJ
o4enmMYPi7dgAuiB1+RBEP17q+7pSbJJlU8zQcQnlUqOWheg9Q6YrAYl2atnfvYR
YCWohKrDQH3vQj16IdBe+IV85duNNZ9jR/zYZAQMqYbfmfuOBQiujof7SzRx5AjO
T0FzyIl1qJOZe99uatSdnp8i3k1cSd0wnAdlMj7T4JLXhvxslMn9Pwdx85P6+q/5
IrGhq0Bq7dSjTNIxBejGdcFdoebFBe+LUUZlHQ3WjsfVuX0K3Aw4Y+qPvH9wI3ad
ObXDqtp1DvRU/62ELW6pIB+zb8191Vfc2wvLd/PYMqwTbIdCA05ZyuqmSb/gdvXc
NyXzC9eQRoBJEYcPmBTCw9LseXSN5b7GZboLMTwvBjE0qu47jYQBolhHiEQ2mnhA
29dV7y0zPwfssYRa5LmdMuyNcuorvoE+PVnksri7/DKrIJvCZhP8JdAXPAemr6KX
HC/GAfWzkTc7TRdWJOhBh94JNWoiLRQ7ZXQD5cTIALdQBNl5636KmcBXjPBM9HWQ
vLMZylZCXv4lqHJ37dn+Vl/oY72My3OYFMGmiNZdQ5odzz2wTs5jKlAo69XCPk/H
IKXGsRO+BIVmxmg8ciIrga2CjLkKfqFFStl+wmZ0B7MQ5UpjEdJfAUHUTXwHeQF6
e8x7g8O2qhQfELNupoIHo6krSvNQ38yCu5sBTtepe640FoQdAFvLlKr5L2ybP4yv
yADOaDxe/c5kolAUFkELY3vBWco4hrnO21uMlFeH+UeMV0eMKuzZsN5vZbhjDxGY
Z9Qai5fXg4En8pXzzETL7jx+RUczUwRlF6YsmsOJcQhgagI7FVnC5soW2A9gBDJ4
415wK0GdRV6GSJnEylmgPtGaQruFvSzndZNQfQMwx+27x48Wiy8B7dhUvSP3fjBP
rA21qNCquvuItyKePNk+LbQicE7P002jrjwa/gPHUYk0XF9m7I1r7Z4cM/qKLWFy
5uJr/DsKKZ2bO+xsmufIeIdpTj+7+rQVRGAI+CMNH3qTQp6nPQHj+kstle8NpcVp
+goHMopuQLQygVJTLffwcMqxNhIiO0hNjwI66NXqZ3OSjwgf6j6+NKtu1/ZBNmwS
U7xHLOfCDBTfakwR7LEE3xKMONRWCIY8Hj3fsfzdBgVtChWpoVk/yqActfTZhOLA
m7tuK1vVEEXmeQLrdHsyIEdy/2Hz5WLLLXfA8G/e0sJRZ31Wke42cE7K5K4EjLT1
jXTi3rwTQJKj5bHGik6Da2WCf7lQOl+bwCfG97az5DKnFLyW5vMW0nF+9WPZYFZy
xe+aXCP2vbkxH3rGDstB8VHUOzLUcawiykBr7zAmJgHNJjTGNpLWmZ8rBv3Rm1Cc
X2Z4a3SSzn2p+1Y6JfcmzAjaOfKQsZDi4Pve4wKJBSf2ddyhA76c5iu/HmnHUhAA
zdm59m1skt6YfIRhj3wZvYzZ5ZidhgDkp39/2yBs0N3L96iyLW8EgoQXG639EJ6g
WUIYz88rVhFZMoOe9WX+K9f6ItEZynVTsnUdkaIc99CEZif1oYe7catvFyAGqbfK
n5CS8qTGWrOXReLYX1uF7ufmt4vHBTTAPGKDWWFR1WP6iA6X7IY79IEC4vzokdtY
M9eaGMV3dHZfHTLGX0REUDX42vBS2YT+kY8Fe8ddHbFilo0GobnfosxyfIJnEqub
Cwfm3jQNLQ1ihQ65E/v2wLwlQhYr4bDIg+nV4FF35Q9ral4xrbIl8Nt4ikoSO6Xr
oqG1nv0V0WJxFstBct1VpJo2HgLqu/vCT/GL84nqfnRJdOSoUD83XFsUlv6Ax278
Z/v5I3xlV3d+GP9e9i6CKJ+jZilGLRRih+GWzpPMGiZHZLwm+z2VQxjGWR46IRyN
BqeJlycHR1eMiajFw3Ss/kJETcEOFgKRndeoN3VdhZYU+sjDDwejhwwppsjny1fo
0Ylnbkavdq9DILkxUT6w6jRr7wiNz0LWUkf6ZGoTLCAYLvSFjiue6hW0HFuDu+WQ
QiVP5POoTKiFCKnxB2pzPY3OKSL4G85pu+2idTt7xphvU5sVxoZ7uLtEKWGHbN7I
/m7jiyZjdD3wu04LHn2OehigF7JZncM/KWVTu4+hOYs07dRbGOhyfUAiMVhyHK/6
A0ix/ukZqQyJSLgirQOcK5tCFQ0FjjH1AY+Z/Ry4QMiP1GqiRABWP9dSV/ewoyiD
785VPEqZYx7diF+tXh7HavolUwQwJKezqqVzjldIkdXxqz6M0LQeT/f6g/jDSkft
3zbbsmFO49+G46Dt1TVjFO2tDFtiVJy69iXKewPk9gHf/B0fZj24rwQtU8xRpI9p
x2mjnjt+EegaESOs3os3EldE/qqhmeKJJLPXUW3rKLF5pdS3lwPQbpeEPXUMHQxF
zcUPp9BHZ06oxOuTvbEV7Chhjqm8rsiabfnLJ28x5Te6DCGpY08excm0DxpQqIP+
xvQSSDkh7F3BdQX5DepHEc+k0CXsd5e5hAqHp+2axOasOmaTIoSg2lslVrxaM0AJ
XIp1vLqcGNlhAJ18cyLHVVbT36bRJpQXATwdvhGNfmbiZKvGmI1wZKALrrciwblz
CBR9WS0gn4DLMFhQWNpS2wgcdJFEBVDTNJpUybVlWjbvK/AW1JTh39NobQC4xa42
XclK2v/BT0FGfePudj36ItJzI2NvUMUoyuNuqFgMBTcf5FYPQL4GT8/Edl4sMiA+
qXJyRiCQMbrN1UTGIeQSK1anrNHMPbVwhhQ3CbORbfK07LvSwb89LtWL1BWkmlKD
WN9BGlUXquIZHVwh9HdubHDvfUvcRJFsob47HUO+QL2PFVQz6l2z/m0ZP3D9nj8X
NeFlcgKfD2KcSFeMMcWPGBpK8c1kvnUC2bdUUGvfWy6DE7vDpSDa/vtjSBHLG7NN
k+NuYqIoKwBSjVxwes8J+OaJZRKrB4qBr8EgGccjryeUakgr+4K18S+LCa9OqWn2
IQ55mYHmfwV4+nl92LzOUfwzJqnyIJhuSDQ93gyXQL8aeTIdy1oTeSVdJWC7fRD2
VKRoCZx+aEIfIF2ArhYv0txLbtHtVOscwtanVlbLOahbZ4VzxTX15d44xtKSBqgH
7YYkHXPbBpWy8FaZwobpWxbmvOV0RPhNRmGg7jdJvunxOuZIZM7Kuacuuua/rYp6
vvJsQ3fPwa2A+Ku6RBt7rDr+HRbte4jnGipKDZ1I6f0oiT/ZR/6oandTE+Veonpq
WboAPD4TWEjPSYyEdamKIYff5yH2/sCKTcgjk7+Xy0cQynV87juwwRksLY0A5D2s
8mnsQx2zdyJrmw4jz0ERfoF3YCvuSxV4SSPR0exWWlC7KS2BimRVNVFLb5NZLuz7
uKFGI39GIoR+lp+GIrmPgJzVBCV7cqC7q1h5pomj9WTFGrY7u+ersuOgvrFpXcx5
R9/nfdXDdlsg48CERHW+1f6cFZCW4kU5+KUQgHfRGTcrQJr2iLWui3Z5W6XjJkqG
4+93N549ReIRZ1JFn/79cgUKNSZz1Sq+bGVgAATykO6ab+5WKNuRnBmm8OKfsRGT
UnNfQWT5geGQsPHw6QBrJ9F1gJTRd0GznjDBqzdiJkSS0m6PS362M7WgyKvDivGf
AoL7Rrg2NF0vAxutIHSs1H1ytw3rqf65udkHYEa49Dt2+xd2jpNExY2b/psVSLL1
tr68kvCj0o91BVFZe3VVh9ut/CPG6KpWdUCkHwX/NQeEjyZFVaIWjPkw8eujRlog
Y5x9rBEQkllRvseFyqBKDioAjOcMdtRLuxQ7lanR1kIzCEhLaMr+3tpO/j8IC+Ev
yQdiB04+syjN+V/62VDWnAHA7oE+c9AGdBchVAeUaN6lBWxnvPBDVzQjoqhxjyHO
obDJ/GtuklZgfunjN3SckS0eLpm2XFja7Ppo87DR5a8H5d803heuVhk+SqKGAlla
8yZZ+Ni0NTY7jAphRjaWWH1At/QbWlZezAxj7yoX9zB3WWzniV+QA9PiqCk/ovmw
zKMYM7+fVSwqxRDpTnS2As8sV74qw5ehY/WS4wbxRqi7GHtay8Q3xup1l4YKpx2b
NkiufHWcCilAGXNCAEVCGNODt0GQJWNyPnJHq5FH+jdfysaE/mmF7qd9FqgB0XWQ
bl7Zk7iI9IufNZjuO6U0NYQGCYkmGGYW8PGCrdN5l0hC1dvuGcGfrtIfEL7+5b8N
lOVexcSSqxtGyJZ+DrGQ82xni+yozcdL5bNd4SKIhi/YrS2Hz3ZH2a7sm8zTH7Sk
txFNuhgmTk/uDKBCpsbqgFf8ox/Ukdh3eRVkS7amFHSSY+eweiGZocV35GS8nq16
iV/VOpRAmRWW/0Z9vBmS/17bVTP5vESyWlQKepb7acUNKDxEFx0GWkgU2xoQQGd3
t2Fvi815rAw/rmO4WaL3alsKKYkFZBRpcEJSRUBD4dw9FQG8EH3bSA8TL4fiscev
aoZfL51HvBe6GdRPBQqYxCWMofJZw2C0hEGsb8zf4umpQgHEfh21Nc11X/VhBRs0
/LHvpymamgC4ylMT60yR1Zum3jPgh2jNbF8w9ZFGFpggRHSXK8j5cnAAb4H0fY10
RlgOpfYHFrSeOl8aKxC5HPqKwb2fO769A9i9LrM/PfOb75VOyfr63Cfk1JpFhWEH
ptVe8xt+lTm3Hj8noJJa/plfLk+9aeT1k6KlyxpT7noGUjWUzH6Uu2qaN10avkXN
EE0JwCpn6jr0HidEKxQ9FEDCRnuCc65F/yJog8G6rvAGKvAkMdgl4gGLxMNxs+ml
m3Y9B2qGFbwYGb/lDyaFdZ3JFMg2gxYHUXI+Nrt1B9V0/bVlZ/2bSBn+dvCCws9K
bdoakc4B8hBcCgjzXcBX7qnI5ciN14c6qA/NCjK3cEB9ZRstPnxnzfoKmObhNsfl
KQiH8zX3YpGTXAbaokiIWkPR52G/Zkgi+ms6+FuE4NYkA6YAZla7Rl2W7PyLrgfR
ueugoVlR+oNjoXgDPbQgDCa/pvkK7Y5S47cxZeqpgEUuAkVhCCaXjVIex4QNZ9Nu
CAUgLqvUVLsokv7zp0Y7vL6rNvXIyUB+6OGAtsxDfU/biopsrAh8x3Eufp8NXYEb
FmIRh6XkECNfW44T1IaPN14kpyacsrJLJxwjzhXC3HeTUb1DbW1kiBnKiTZAgaGN
aSL8dZoLDyioxDr8qcQ18uIF1O9K9xl1KCINQJ8w3ip+ndrn8pAz24+AaDgzTUJz
mbWii5OLm4Um/XOU2Avmc/9WwMIZ14TkaKHTT5oguS5GYN4/At/BQHg4+VU2gXQE
bTXStx1p9BQXq2fp/hjSLxF8K0c69A1uLjgYQ1nyJoxZ6OG/STk6VEC50WCFmGwv
qS12L0Rpw/jbRYjWMGjxON8AKM9U73xNnSlV3I4yVSLJrDaTEEASlg/w97oel+5e
ZElDwsnsDjKWDIlWrQGy0ikqHrg0VB4fS3Td+GbL1egPwH13GHDFTXC3p079KDp3
SKb7gIYH3gJ/gSkH/zqUZco8dzqvrtSpkIO+J76Z12osp3XTmFWnmnjnV4XO/gLJ
zL/C1+yQVRzQ+Jp8LerAcsTSoGzAXZRgODuwwSSdQtEqwH0bSA//CHWOYCXXSIIF
utzaJ+FjLuf4bWdW/7j/PzfjrmQbgwOfWb3PJrwUQxeGr979cWIv+z6IRW1aCwaa
1BUZJ0YIiECln+Wz16+n/fB9kdPQ+Zp7yYwPx9VgxxMrvj5LUhfMZ6IDCjcGhqLT
xeH3NB+gCxkvFXr+d5kVdKk1wCOfkGVec1vqTjGqva92WhTHAJvUhbR6OiLocdpW
YgPBpaZvND9XgY17UyzrapMErt8yHRmRjVPZSJgUiYycbEABT203Jx3TXyYoj/18
z+WQsu4bP5zs7M1cSzlafnuTteHLLKKnFcu4L2bqi8guw4mBbZd+IQEl4MRAYYUb
Qlz8oBkQcaRRpUOQ6KkSYO8BZC6Fgfu3manEdOUYwDFQK1VuUXWJm/3dN3Arf4C/
b2AopF2Jvw4IpoKf+kpJpo3f1SPZfzs37ArqPjJxs/XzDr5xDbxicYNPIEqwK8yS
N5tDaM65cV9+zEc1v4a7NzSwwJ2SytXR3nB+7eFEowvU4fwL2U6a6mJlueOaP90m
CCzwmOm7TH70FvcVk+qHaYzACVnzV4zd+3jJwnaYAO+sk8QE05EjLGOGMp3emYne
nJb9Qs24YuetZruPCt8cD5ayT0qBNdVuxQaFW1xhKChlIgwWFeH4hi4AcGY2GQPN
tbfzHGDSM01/Nh4UrBvpXBFwcPSSEGIuLEyXPJ/gSWLInJLGR9dR1AeP1+uXpVBF
VGS8xjfZ+5l8c+vVgZspc0lTMRK8eq+AtxggIl+NKCrAmyXjjKhheTLKKy3aCVqd
Y9rxw3aabI9D6ghX96/zpW5GaEyaakopeI2noQ1/EMC9WJz+WXCUu6bMPUhuyOjt
40Y7MAHghgEaykNuvubUZt2w3rgPu7Sy2bO3N6Mr7aLmwLNco23xhsStq6YhJ04v
2QglAzKeigFNhzQz+8DkZHDIL86nE4udPURmV9GJSOkGbFAuwUyICESVYdWB9wGJ
E0yhPvPenlwCg2LfadAHtMzAbXzKslQbTKHkRU+hsAaj0KxheNEqaKEdjGCsQIrc
weuklHgHOw4cOIvLLoBShACBvERgE3eEnsgnJHxR3FTwlyAUtmiA5VzgwH1kLcyQ
9JYyR5f/+qrMn4O72wKINLt3oCisTV7UBDakvB+ADgmc5dI3AIeJd3TxfcuxeYWP
X5fflnYX18HDg+eP9xOOcks6VdCIq25Z0I4A5B1g09K1blkB+6v2KM60xfWBLrNb
ujLeUFqF8ELZJgtjM+Se0/9F2zTOVq6OA0ehzMr9yBvZSfMih9PS9MBPE6wOX5jL
GE2+aI8pXxizK5ohLVdJx9JMkBz33XsIb9IGv8araspsO7WSfGBhXhSGKu7Tnejf
xD8qBLx/e+3YJ1Nz2eKk0eoq4PX8tStWLMBwyzt3V5r3iX9AWuEnyEvmKSKDj/NV
4nxkmVW77KD8dJ3inHPiQHhC4ah7V9/lTm6/AefUtKPjHeg0WjX/mExmjzQxx5Yh
5IbpRpBZdp6RC6zHMpp0YzccC7uOygeVa9noy848yBs/Sgughzz7rBRAWN/gVvuW
QFAlss2HIBUk38qee1+ferc+NdvzpOH4zny8sy2oHv4ihlep5tkNFtNGDxPz+9/e
p4uJfTVd7vV3JDao82blYZxeS9fdQDOPcuQdXy5QhiahYzJ5wRB0kYDC6GvJxHAc
CcGXL2vSiMTAssLCzHfe0yw8a4iShJ2TFyoE7HZVUmvZybZGktDgZ6SS2dn+hivE
qloYEAJSEAIJZ13d32H/W8SZBDt2z+2pSyjy2taxCvJxYkAoITj+7+js3LbUg+nh
gl1RehnQF4wON1BW9ZFjAKl0UF4ha4M2Bg+iVqtbeQ20lnMkAXpMn2aBTfY+2Xzf
zAkOshne6l/aj9Tu+h2q2fUx1AfZ0RGQ7JR7ebX8QiOzkKvxBQRD7Xq6gnkULCWP
QL61by1UpBvKF/hQSk/VnaVBr45zuAcBkpfMVVCRclbhj9VvrE6+DBlLEER3vqNn
GlpTLqfc9ffxX9Vnh9MdnYCO8/bXI72ckfhv3mxvyz/CEf1UpcB17H3euAlYwEsU
vXkUqRPBvWCacuEGR75LN8vdSaz7eVM2W1K2ZShuLWLEkEradcwuhk9L19zCXfHa
Z9dL1GaSu28P/yCpZZWcIkNIOAc7T07jxCxPREtqYIjSku5hdge54ECRU0adny/z
1e9MASuHdYuOnH3xej70W7MsgcW+T0sJHbxntQMkpx1lDw+aH+VeZktANQvL80nA
yI1IPV8+258evNvB5oqVY+Pv/j7pmUGM5tV1JAmwyBreo3OwkaKAxFu9tEveIMHd
jAI+O3kjSPJD36b/+U1SGvbW1f1c9/7Qy1aco3rtoUg5/7KuVnBA6Fy2gtoqAAt5
ivg3UtWifLYivjwQkpECN8YXYZd2Y1LxmQs2Lwreq0n3Fs5LVdEeN3pKFB1E/StP
wDfCU35U5JZD8BTrN6+lNipG2j//pyXkXPv2Eivy5wlUYW6o1bl36yTybyPKIg5Y
4ql9u2dXSFsODIro8VZ5JATJY6OAuUIeWrPQ9zNANpELGOievHVMbk3OiLE37U64
Lg5okFajE506QkHX1mBEMl2k6qA57ODUgEtcHCtFI3+lFRmX9MBXXeS4d0b2lHHL
1RCbPtd7KPtkFYLRbIw5u89KDotdyOBR4oTdi1FJsiRkunXVfPCMhgMvKBnrytYi
5uJzgcYkNSJu0Z3KVN0ej5Yf1EnJ1dYQuRlWjon4EXkRVUtOmwz39hVeG+eSy5Sa
qVKDtpYmuiagThIokvrVZBgniY5VEhX7rrYKC/jmvzwJ7QCPS2Tx3/ThbRzrt1sg
mku2sqzG6q9JyL4+LbrerZ/nqMmUd4uu/Y5zL21WhLfweLERvUrI+7q/+Cn1R8R5
YjX8XXt+enkAA3dMNSJfhbqqudRnKUBCezaZ8R1EgNrbLMiNsMiLZnN+qWtjdxjr
fP53Ff15m5a2Fs0oxlBb1kqapJc46FJaAyR7wHY5OMwUnY1NTzZz8GB4N4+zkQLw
eWomHNUFXTfengdnPo7aOme+r3/aq3Qm1OLWdze08mXVhEf5i38sGXtEht5sAHck
Aq5lQmf19+/gIhCW+1iGmQeCpmCIARtG/inyVPABB7LsXyYhwD2VPqiFg/yTlByS
epqznyQXIyS4TbD7ynd2UVAvCj2VYH49+EZQ01eKIP66dbN+yCDt19mIjGikMCl/
h//wmQuRL+RsRUIJnqBgZF/Dv0CU+XnxeKVavnWrEtH2HcjHhlFKx8LKRP+7AYIE
uh3GAQWCSwAr5vRrdGmxsyrbGrPnpayCI/JA95OsF1GEebT3EiEuLqYv7fS2ZMzo
hgZxT6GSAFMzkfF8LwBpiDXC2TPqsOXAknZWJ6Kby/fpwQERVuZ5fcXRuobzXWJY
/2JCWau8wECoF0A926uvvU6E7fhZJg1xaDYV10+98zHM+3pwHjsuQIlBClOk5QUR
6rkEHMX9HhRLUpqRgolI8NO6Y4CgPJmVPRN2fYC7G23QmZ1h/O7IlNBcz4TqygxW
k4RaSENu8TLPPCOMv/wKVJ0qol5LTiRG9SjZwnzPtSxSR9dDwujdjwNHfKKoM5Q6
eSbZZOtDhPwVYU6jNR+v0OURQcK2t0YOoIEyC0Cb9EuV1k/dxug7uRWgnRGMLWVH
kx4reDNeK97zMGrALa2Lq3uem7ZiBLmjaRVKahR6cCT/vqGQmYNbsLY5KyOuDRlo
4HVWr5dhw+zAGYROOi1AVu5pnR+8jaFghlLroAcItWNYbeUj/o9WhNby623IpnDV
ttEA9KcJ2hbmjb1Jy4eLgRUX+ZHdWHPPf2YZLAY0/2h4rNhoojbay8GJ4EbtMaJU
EglPzTHx7wdjq2Gb8V0CJdz5d7e5onTeIcr1atSwL5q/aZkYs+ybG7pCtV0PSQ8k
NR6rRfQw3CtGBGndGR7WwynkoATIYOGBXpPANRQmYMd3kQcANIzZzuwuPAZZHVQv
d3xe0ZagOWYWSdSHutQbIfWl84vk31BsoJHoHeNugff7BSh6uhSsHJez7en0bP27
/IGPF19JARUcK2yXKg6yIXMcpjM/tT8zB9GMIrNNt9p+g2mUv0gkryDS3A4BOU+N
CUHY0Zsq5E072ugFRz41mQZXl0zm4pgRzYgF8TrdAFiSY1SLKYNU6Z7sYSgbXK+1
RDXaEyr6tfYouJ4d13wTSC6ewaVHWiAfw3oxlJqMiUspPrW4EXpDfGxd4yh27+iZ
o7EQNwkR3YDTAsDdSmRvn0dbIN1KZkev94xhPA3fhm4F7auUCsYdMwHtNpxdOO0Y
ej3JpgXgGZCcNmw2hO4a5fT8znxY3hZw3Ctk4lYn/NWwcK5GXK2nZJHv84/lFOYo
aVGEMMJ49ZLSe26dM+PWbD0djHs+yFSSLzAeISfpehlj+c2Vh2dk95x6WsoWG7dm
OXUhfHHcHk7EGQbd+huiLqfDwoaGFMo7j/8Y3m3hvrtXElvtVMOdT8PwA/DGoMPd
op2oXZ+mrIX+75DGLI/gVX7fmqsPTQDC3UjrF4d+R+CVWbwAznCf2eUedbi+vBVj
HoE2XYkWB5sxQDHXR7WcTB+3uFWX+1ZWxsobhwBP1X8koZBH4skrt0Pa+77ywsHD
uTySHRdM0oHDdF3Cedg835Vz1mIa0JNITu2wdHvZUjauXF7UbngpyHdGRYGOR3TH
UsYP5gQ8uZtFUnQugKfJkgFHY5Ep8jxR6WgVQfFeSRpaAHrxhGtTnL6Z2D2aGlyr
SxkcrzPPzauhIykoCW6TL2P9CPoYC0REcnA2hcVNion4p/0nrvPGZCOuxPmmFD5+
djBD4jwGg/P2BGLqyPgfBa227/GPuktweUgZtlbbahZ+VoMqB95KBmnucHibCmSE
5axwj9Agib4mybmMWKoLxNcCAiZ82l/f+j1BgeHpFcBqRG9NVEfyJ2MASObBb8fQ
+qMLHTtYxeVaX8LPBjxiUSgDX3rlR2aFGbIx9gFOW6VK1tN+DovpdK24HFDd9vMI
euD5yTtt/pGGo9UqW/SVohDWH+uzVlK3DtnXpSUd0ioZ497V6i1nVrP2rLcKnRLg
yN9UFyh0i4CdsFoHl1zIX2PGN4wOr2Frwte1F3W82rTYy3VbInbxwu3H1mHhyKpC
3WFWaOEeN+3uUzw/Wu5x7IBj0qRcf0aD0fr5CxinRBaPmwwM5/9PPKcEkgIbNP3P
M9pHagU2Kz6JBN30VraroLN3EZYQmN8mackt89/GcLzwz8uf6I70Q26NsWYoheyi
+jbqI239+4XlHYsHQWEiU69tqK2dgLnQAYQQv2exdZOJKNF5sgKAC0ItorQTTwnC
j+3lVfKD0JhSi8aUwXbLbV4qJmQbGdF1ZlxMHpfB45VcQnprlTCTDSStVc2L4hCc
43/nSeez7oAxAK/FN1sa3d5rpqruXVozZw1T2PxD4PoUQdvD4EWPB5/k88+EqPBd
6vNrakc8Uk8sZKbnApBJYLo1t3Z/njlXxarhbH9abG8XA8wbgdlgvqWbFEtjMBX/
ZNBqesqAvyewsZjmjVLOOX9JzZ+73KIKu6iM8avvNnucBnQOQJl7EihhoHHNmv3M
gnA4JGW1wkLe7xIX8P7lac7npatErXl4AxB7/C5BYBQbqOm2uajpmSRaULsWlZ1G
/7ea7+Zj4YgU7ZW0qirV7znMa7T2fABnVAXIq+PZXUQsFwK0Z993K6YyTwNvPpkR
LD7otB+IZFqywILRDyRIFNzDTqRzUbl8B5OIZhDEx3uGy4wdxEYF41oEny4t95fn
nFf0EUf1z7d8iQ/YDkvGpIE/apRL5/0NoPDSGLijbiWzPtgVwE0bIuVHnpcOJDus
3ug3ToyD8nMLsTncbwNnLIonRRSJ5F0qiqg5NAXt4N2zUbrPt8/tKBUXpZPkDido
rtwkCDhuP84Z9wgMQz/zkqEaiIw358iQE+gXgQhTCIkwVGAF7rqyZhM4H9Ido/2Q
EvHdMUQvl/eone85n1xHQGlRnEUUpgV8KCRF4ug6beDhAupZ1q0JdiCy64SeGJYi
ZFTECGsNnThlARwyolR0ol/08Kx62N4UNNbfD9UMKiux5dEBs8+cn90Hf4pzkWip
sKAzT1qOGANt9y3avwAEg6u6C1XL/bl925z+XumO/BVSiawLHRmeNWOksc4NxRpa
J+1ubhIsRFh4SEJy3ERdk3tqgnzkXEDmFhjyniykcO5jAyQLnEYaKwnOA0vZv+N7
OwHUj7iBzqJ/0ZrQLSoc34f/njEU8EOgEXq5oQDgYWg6A1kL3MFLtabLRj0UoU72
8o2+QJXdYe36dMpxCKOqqKa7HEvICbbma418roSDCYfNf1dv7Fxz+y+XYl4Grcq/
0QHOo/1/QERNWpWsGDGrV2OZ9/KdUYEt4skifxSCdaFI367dcFRJHyG3ZbqlETDF
ycTljGAAFscO56xmvVlFb9Zp9HanTK3bkOb5LtYda42r0VgSZfrLttx5ZTz2PGXW
O/hirq+qCuSmYk9aTF9R0q4j9KLWVuMhyT1XiIxyXn/NGsZLqoWoqfEFTFPMAEIa
sP8+tmYrTVO7gK7V4cxQQTzXdazkrRFOuqWj6Hbx4sLjB23gCvSIvpGYPr2qGIv/
xLA50KOUN3/RFl/n8soPeiVzI3XnNipe+1r38bjppvKsVlyV1pOcpkVL82cE1uVK
ncXwucKvd9LU5qMKnxUA+aA1U3Q3bDdaYm5L5Y/xfbQxt8/dQ03gShUns2ZZtrID
vHBlvfxcNACqIYHdxQFzXKK9S+iD1MD11HbOZpyjWUtkB06LV7p3LemjspFAPIYS
WtHMYomP5yj11LYigl6wdud77Ck8izDMj7OuXhmTOQMdYd3I4DbT/lomXkpt9FoL
5hTsV1/FOmuvdHQ7ODoGUzPpfmWM3i6kuXKyybqd67fbAkWdzveMKqxli5pRGY7u
jvoyY2k499jwCpGD9w1+yvbpd/EQb5c+FSxZn385yHj7Txq8+FDQ1IB+GuC2F78b
yUdQ6fJ9gHcK1xakqIZvloHHMYi5P72KZCli6i8u79PkDfX7318w/pRVctGTT3Ij
/xRgEJ9H/jJ5vgAr4Vrge8yqEwX3FyRvu2DTslSp543VxEOIFChOls/0VbkhYQ/q
8F8of6m691dm4FYfX1bKTS910s23JV5cOMA/pDi6KmaQ6FiXaAjM2oJZVj/BSwnY
98+UxVeCek59r1Dggc/ERd/R4Js+ZAqj0tEQP/jJcwJsNZLdonpbEqHN2BQWnnaH
9lXENjkFARKjGMX69j0mVeIbF7vVuKoLuhqeqc0jgMqADvF1GEw0DS1pnrBbWfJH
VYNB34xgxMPE3sEOY5eaAr4xjy9++1PfzC3E2FVh62ZNlDfWhGDFiYpI2aNJU4Wg
rnxQK6M2D0tJcdYo57fxTt1ranB9QUUQoGlNA0EJwqzHDuD/kRCnj0D+Z79qfflx
VhXQnvPzedykrnEaEWAz3+P81ZSa/gTc0pJgaMiMXa9i+py8wUfO63Nfktpgjqp/
/Rg1QPo187SNahA4F4qQ7qKPTMo+I4ONNH8Xca0hE29kzGOwgQJfWWMDfKoncIxg
DQv5iAa/kkLvbDX3kJojZsTq2DOOrTccJed1MeYiOE0JMBQ/YOH28uMhpDyqWQXG
ehR+jdrECxGquA3j9pteK0fyYIgBHVQn68pbz4rMXDhuxxkXj6TrZ6E2XjT58yrD
VMSAGI+LtxQVcmQwkZ6J3wTU+gbUAAqrsNCq0zumjoJQ3ubfwwyVfzMSNlzkDfhg
vrBhxpl4Wtoa8KQknKO4lA0+ywyj7PyGscxOpScaH87Xp072jPZjRD1M9I6MV/7V
Rfidi74wA8hLiZuA5hwWl190Nmy9sGwSXWdO5GmDYrFK9DSxtws+ZN8FDeUPEtxF
g53NLEw152hody/s+yszyXXa22tgE08xAhlAVCxl0ePeGIe2iTnjqAKv0LghFRdj
OGzulC6jSpNCnsLWzyxKjskKk/tAZJXXhpQabELsdBIF24s+MQWrvW5TJbiaaITa
i71KB8CWQSzq9hxbswD7Cv9NUiC75rMl0CvLyz33/ZcM6JWqLw2J+Pl8qCvNZoTH
VSMz9ZOs0/yc7gZPg9C0NeGPJGzMTdl/E1GmCuXGs1UPhJqk+d8tEbWRZoEWIsCk
DeiJfy+lYJBLBtyBM0YAM1TUAxrNTitOBMs81PsqXPS6DB9nZ0iOUMa+gjTiSMz6
xhgSUqQbsL5NWTnOG6PuJ6bImc9g7qqbsmWpzklfow3Ley4/K3gBuCAHoQEUYSWt
VqC5xKwEqXQyk7Wd+ELTYGCxrYLEnG2DrgilRlFpwwWWxNSuRg4Rfgn1TRJbvdli
6IDnHS2FlX073fmntKcOK4uwmLy0NyrbFb2pdIiFVE7WuSvr0lAKXZUL++QQ3a8e
G0ZOpiqV4cuJKGlbKOzYcZ2QdKaJzvrqnuTLwTOwu8cTOU/w0yl4y78y6KbQNWaB
jR5oShQ2VT9/fa9Qa8qERyWSU72bgEuGq0OuIiUXKCUqhO3W/a4Z2SdNCWwFFbF2
q4twj7VqHEcs+KYrM865f3W8hnVqSkSnJ3hQXRdEkNKSFvgwoAQu4UCrB+zcXBcv
Fkcz0iqQpI5Arb/jAyRNI196UAiFCIHn48I9ItU1qXD9qKx0fDo7cf9O1XtoATBy
ZHK8tWX26EjYK9OHpxD/pJRp3CHpg8KbbvvMkVOfSRwz+9XimQwpKiX28yekCJxQ
8eTsBKgJ80AmUhecHB5jrT5IMM6SiILJYcIx2y42MuDb/0WUnHDYrPwou3EAdYZ+
0VmYUz4gx3qxDwmeAvcMtgPIiMF2Dnf9YqmeLC9BlkQYLiieGMONY72HQgEShXIC
jg5Ja1wXwKxKnpG1/AaV1CIKJM80ByFkiplKWWEDVFGLk78T3mdzG5LSWBi40J1L
y2fVkHO7WZW5b04lXbwcjF0JdPpXDXK0Bc9SRaCCgYXqZWouHEW1mOJmIFsaGxBw
Ni8KGh84gvfliFhcJ0kpHvK0kl9oWtEwzQavcotLzi8RVFlaYNy88T6LGOlMlQT8
Ojp++CSwQt4RNDLA3YPWBHnsTNn+OHk4vcjhUBIbqCMCzhApxRDDdJueHKNLDvc8
G2lxAJcBh6GKG7td9P/r+fRiaiWa58q/M1MZkM4zC8eQ5eoV836CED1pzBS7pG6g
HYQ8v7MhTaXJv+5IO81WQC7OXorz0sX806CyDPW1RWgr5Q/NX1fr4T3CXSNxT/AH
hXhvQtqddDpNu8wgTXKACd2xVzMOeLbqPJiWp69akxQ5A1MGiWSF5g71p8h/5q+K
1E50H/tggI3LI1wiNjEHnBnGH5FpmOSDUhKgNzRZ9vwmtimqINsSBNi0kcbJXC2T
X1k8TY6CobKPXi9Uz/Gx16eqpgtyPUXb+g5W3Eh2mdiTu7xi/z1S2TbYFEWbyrfH
bYzOctxTUAvVMK6NTePIiTGyru1QVoOE5shZb8HFHPjmoYLwqAgsiB8m4vpsZ4QF
t/aYq1Xpj/1gaqCXQR6cBUlaB4z7QD96NXYhV4pUuFm1qvjhrUrfs4CpStXvuVi1
26dD1H5Yue6EsQhKydjLR43kp98ZNfyldrmOdEcsw7ytsRSwxiMMApr/oR0kEKLJ
YaWopk1vptSPZYBCH/aGJxVqWxU5eNt8kj0XnkoL7mmW1JUKBx5xBGT4Fw3hWGfd
9BrUrxs2jAelbHGcJhBd74lR58D5YkGE1QVrDA/bOfKtaOzTpuZc3NZWJiJUemNt
oQYQ7i59nSMfv15mJtVeP8D7MNIDESIUQtSL58Oh71YXzdVoBpnoXPFVxlM5+b9X
aoXjdJQmcmZdSxoxr+5nAk8t7BzisTyT7puRq66BV08X6z43dAuia8kxXI54sNsM
Qnve9eVbAD9DnrntDvUTPWxiR56XXnjAAMJAUg+hRd49sQbTeOCUmS/mF5HRhYN6
F4jVA9NDlJ+SaNilIHoqeoyuWiu+YBP9bZpZcJ06ohGBIxn5EsFGAcq4UtpNq161
kkRZvT9lNSBlRRUl1WgYNXdAqRz5byGOcjiHPLxCkIXdXWQBsLLOJzsPdNS8jc7c
dj4w4AEPz0MjNu0XWTkr1LZjF0SWHSIzIR0xMC+jgJpSy46V0ZOg6UFiYzCifVp0
FVkMyfU2PqEM15jt15zVGviBM0C36qEDzsYBL0j4UPLPYLxBdeQKqJfxTdqrFOPv
LNIj6VRzjAmC5RgRhKgbIOWirk5/GlkTlijZEtBPEinE0JmovWxUNyipC22DNXiV
f109PABmUNbO2zsIFNkb+HNI2rRtrJrIsruXKVEIbqhadACMxC66ssvQVSEJPD4V
HIlCShTm5dJP1LBxHANY768hZVwGmshoHpyooWuFtWPKJUgrz73xeA7mSp36HAko
Hi04JBRIBpjFRTgIl5UFkiHdUGmSw3qcp9ypsoMfuCTPy+wVArPOtqC81uqUA+ZK
HA8cIZAy5dcSGCu0uLZjVlUelBRunkNryFx2HXhTSAum7AouWYPrMTnbwlfkO8d+
ScuO87KJnb4nR8x0YYaw4vOloeyEVFdwLKviRo0rQw9FtP3ade6BjFXecTOfYO1V
PhnJdS9907a0FYCLFi4N2NRiT8NNge0sUAIodkxwmb8VnFTEtdHBRobkgBIpQaLS
uLUdB8zvtpmqOgQBiIT8okiEMbBs99uzN43lYs7UXgrdJwDZjs/+nu4WgibVtjdx
LyLtF6wm8+FIh7IiStkAz2ZQRmFpXdLyZudjH9S8fgtXgn45ErgeyOiMnMlikYYu
pJsJQQNBZbAubnJ/sQlyOIq6Vszgdh6RPZ5Nkdsi5VJZjSyqwTF7UOzpEpJcABpi
aZfTn4LgARrT03crx1LjyoZ5szcsbKHMDSbOrCh+efZsaOMSSxR+xPdR2ujB0kv4
Zm5vkVvHhEpv9QyULgyqGz4Ha1hzuRr/f5LBK2fivNnnC4xAdpzgdiHDqyNON85u
ulE/7SgtnFMV9cjzf1SpYn8KFeFgYuE0H+aaK09bqLSMq7NnYHoWi5XKKqPjJbMl
KJ1yOAthlzk01tfqlHtFqAwzW14wSrybpOvuL39bopSXXcbwYfS3j5gm4yqYonsk
aOqTh6Fz7ZsQbLW4STW0fNRl732UzTW+07wiC9tP/OE1dCrXLnyrEh5dvsuVozDb
40zKWif2byBAmpWsHzFNOmyeYIxLIfpGTFv05YYPX51TwS7hsBdeKcKBqgvz1s0t
0BN5d4cJvU70g7K7VH8ugpTIzS1bM8OMvL1YdSablGghZoF7bni6W2JUCpBDpECR
O4uEn7MZM+aMXACW2Py9k+XFIaWZ5UqkJ7Xj7z1z1CnwXAjC10FGrGDtWVua92le
xszNKiL/FJbZG2+uDuwX0nwLVP+5NKoX3AJC+GuZ2yEcIGQ7r50wJ8htMunUki0J
NRIijp31NM5v1rsMKfrZkDYjamhQgVw1SmV/+4gEefSdbt+cn/wLv1zCUBf4bTYa
fUsBi++7kFwSAPGNSD1OQ+XguP0KqzYmyj98UQYxfjhbKArlPD5EijTSew+NzLpt
mDk+bUvDyFsCdgpZG4DfJM3bU1lLQ3qzDwg1VQ4gq0+EmGXwfDexJptSfqcaQhfe
VQAutG3J5J2EeUQAhoqRFenakaWIzFhbyLR5sn4HvABFGn4NkpGkAJcEBhH6FAcy
PgwegGmvyfGg/AH5XOj/TE8OPatJRS8vrDug0c86HTtm9LSpRkI4PBsUHAfDnD4H
Zfha83FYN5sC7235tRT/rhYz816lUOE7jI/OBcTZUZPZ9tCnu2v7C7zz0nIlbNxe
fVLepnjNLLqsDwhi6Q0PpOIgJMJVnQl54UDW6m2aatYgUD+ctu8wD6aNslYqJbHE
r+7UQkYCgEh+tm544p7TpYbWdtef497nMOS8Wi/TE3UOCHHKToYSUybO8yE2k98B
s/h5yH2A3148nrHPt1W2RbuLR3zvS58NgsW5o2K0pYSqgSxmljaAlF0cOtOAltDY
EWc1onWMPmRGTJIGvBfp0EH+9nnhRnKSPxA0Y4qmn7mtSD3PYgp6DQkTIZ/alHLF
TvWEPUTh3aSeBBi4G8e6EEsmCubC7viR7Td7/rQeSdbrHYLDEVWdvdHUsTXtsFMm
JmRNK1lzOZDkPskjQwPuu3r5alwwKCqcQnslBbV23MOQafJiNniZuM7PZIPnI5DY
ThisNK+V/UVc1tKU/8p/ggFqlSJ9kodW7D0d8jfi264oFVD0zdHIkZDTzZD0Wm1p
svqKv1C9RED1LjAyHzJoRmNwqXvanifDQRyp3ndIeEKZrjdnkC6vARH6MemaCTHp
KeZfTC6gVmB70gmCwoqAdYT0vxbs1QFUbeg55ZDcp42UkYwph5bOghmHqSwiSiGa
0Y0nPcH9iDXeDC0ywt4qXvUArpCGkYh2TXtExPaFYtxbjC1jSDf7m6EFvj0c7DCC
/BHXuyCQ3qHvYG0nmTvqgB1I6L2FF9kkIzRX5u5tGUfxBwbV0fLDGJGoCVQwqirk
zh+4gRiabSOKtDc4FjidrQJWdsGWgKb3QHMWXc/VvsMFbcy7/7dcBwBPs6hPbkvq
evEOKPio4ZxCf1iuEaADdEKRZVowWiXjPIQ4mGk4TqykSsqA129UDAcbiVZQ4mea
UzPozRZhCQI+bV8nEhRydigHfleBXAyULq198acxBW64bTxkTRpsNM8aTo3hPXoV
QMEPy4FSUrlrhy6Jcvi3vO4Nc/3GXfTGEzGASqZHSQbNzG9mwUd2iDKCL3eIlgqF
R6BkdOnc2Oe5tx2Sus3QzdbDiG74tRhpYULHha++/M+yHQFZA/WA0pUGnGQGo6xn
ChrJhGyEmXnUVeSoU6Z2NIBlPGGJ0Lj18TqZJ+GhKp02+oJcpF4Zfioa3oZ37RZT
lG0R6J+Okv7sMokM2K3p3yTiutY2zrTya0defiBF8MpDUF8FtKhd+qimzLW2JXXT
5yCRQl3C5092tGnxwgoKpidtfVTiG/GugdDVsS0/Sw+PLdm2lzTNaQFhWSfUuOtF
UmXkZgf8vEVSBWI5cp7AOHNlzUmdLBUf9nENSE6Ce60KMpHv1WRAQbAyyZoFubQg
OZ1mwGdOKEEpwyrdRDk/Os4qBCntlmwP3UFiuHRlqGRGQdFhU4rL0pmoYri9jk9z
nnyjQCvxdV2n9dnDWK01pHaI24yZE0pv8ih0CdlyRS4Q7abBTFZI03aSrkzQhCBb
LZT1jD4J9fvn9S2HGsBdVvHXAHI6olaq8K77emFGGZ2jQuQ2T4TkunOfPKi9V02O
b07h/Kxb8t1WpW6LXYM7/oxJmnORuzjj9UA61u0iaRzqeJrfnZxxsyCJprB+OpCi
DfXk6Bl5g01DMtTcnANaXj7NrulEHY27xgbOWTeo6utDHpqKnk/KzTxn2q/Vjtoo
373ipi5UNNT5ywY3+Ux6+rtat2AuAc5xhfiDQ/UyhH42gXAxd70PctAn8TV8eASU
CSrKNS4eOg6DKGKITHs+77+QCR5yxWGlfL5ddjm9+/WPKDMtucX6I6D5vR2TVGxv
3IeMd3k1SRwuJAteqR6H+gFdIoC2Lq5wEiRGcvY4ETx3eFVgNie9hFK0wGuF7STQ
C2Uj+7CF/W+viX5J8FwzFEECpWPJiEjwtM+RO8Uh5yPnpheqWrsl92bmbl8KKzUf
tmU193A8LQZ7d/s1+uOhXC94osWFbvq2wLe+I0Qor+e9uTAjQcjnZWy7HLej6Ufz
F1Q+Ia0ic8tG0TEDRIt0jmFLPc7WWDmw+yvIz3L+KFNs9jLgCkLyIwNc3Mb0JudL
CUD86Skuwj0PeMgj7+pXNr2nn9dWuBP81skgRfQStnOwSFYQ3glVOjeisFB8Z+mz
kn8DvoOux+J0z6z45ldBJyIm2wSWNITHFzfe9dlwcg+QFzXS8g9F/vEFfVis+p7/
1Ds+oFL0wf1Zyx6rryd8+Nh6f5U0aF0SSFEV8iSc07dHg5Rfqs+CxZvAOT42RkrP
4aWOLttiffXepM9kCylGUzRcZOWbyD1WfpoviAyrLI+8bpVEsWKpZkNIAGUdiX6D
OgiS7hTccRWjIzwZAmXhxJCKUebl/KA0LuY2YId3k3/HC2vJOQRAeEjb0P5iLuuZ
fMer00+eVT4OeXa2gDwfUGcEf8dt4QXoOF9Fp+cJo7Dm/YcDuPUVHEPmYA71QMNV
pIsw1dFETeLUHYouOkqNWe7WlDoxx9QpxNJeHuoomiL2peekkEEKGyxgPgorMM/a
g4tTf3Qx7iXmsc/GjzXnV5UZaVi4vQoPdwfHw7rkkM9sa9ukQcGU1M4yWiKeqKk1
antHVWYxX0+nra6QP/vLNoy4y34GaQ/Ojr/Q1YG31UaBIZC+oFg96rlsIFq3nzMy
dyPwprMwywPiuyS6uOOigixowkYQuGmMgokvNuA7+hyNb+Qeud3JrP73B/XidpGc
Pvl8mVQkdm+unro/RbbP3rHt7+FQleOA8HcL4SEknLrSGxKZqTs3Z8ZUhui7mJOC
IjCwm32YwXlJIx8fIGUntvTdaZFCHRA5CSYg8IyVMH9Qu3+TUER5bRmN6bVO3YwQ
DA06IxSC3PHExoea38r1tV0xuN81O6bYH+F0mHAhS1LDyiXmznmGwT3JNEB+C3X0
mQb7Ea7WbFsH/AbNYNcGEEvi2gWSAcHqMgfmG0YLMOg/2Feh/Ary44T15iaG5gu2
lyv/9EHfMLO3CspXX73l6fjxmVYynzT31JAM/xLVp5nwoKZJ2XrJaHpEewXjiCl6
fUtUzqaCEFC1KKV8K2I3Qh6J16jdXBYTBQaqpNzc4q4V8cGZoX3MvLhlN779uqRr
lxWJos27OskoAaWow3gEABi3gwacz1aGHKn/+Fzz1uwDZl+GSL7FrbDgPAnWL6J2
Ju06Kp68EHn7hw+WqisDXnRkwLyJfDCR+0nRE3P7gCLwsV10Zw7V98AGY8Q+exki
qH+rgUg1xAaJEqlD1U9hMQSTNJEjka96OZ4nl5NIRWVRIA7HP833ReTO+NVvw15O
k8AFTczfwDQgPbVTEstPlJdl9eMuU+IOK2VvtntqNpu9CKHshdQnyBJKeWdnEZTA
Ko2Q7E4wmZHUuDEaaH+hxGW3jvhRY2wz7U8HznuRwXfmIxio4xrOZJuFlkeNhPGY
7xvBpOAYyrH1oG0pbVvRWkpmhlS9WqLzvJ0llZyU8i6LYrfpkZVZGYiUhvOOPx1k
+0vI0p67P5BDUUgZxwJVWbSuCEOJhdicJ4+KjEZxCM4kg0Lwwq5DS0IWrBBomtx4
rqej3uJQlLUU2gMglfaGwAsRST9vZfSVE8WfezZSbcgj7xPyT7O86LrtcmXpxfcq
c0ohkQHRrHP90Z1MhsQhwMoZS5LeaMrl1PPdhCoXfttQNZuNSW3EgBcD940BiIoG
Ti8IZARyiAJrEISIXLaU0OEzBdyEQzAm+3HwI3e+DmqBBQMAy2cS5s+lf1ykWFb5
c4UVeT+xkbj/dbuuquK/FgJAA/21xIatrgD6o+5vWW84+X0iJK0dMyyn8RjI2hGN
AvvQtKx9nJ7+ojDslSNcgHDqav6w53nCMfPRozgee8p91QlF6iFiECT2zoTJ/5Wo
GKHcdXoWcUJLctRxP1+Yv6hDJVqHRPqXStaN5wVDrknkZVlaVJKxLQUtaF1ZB3Zq
BPX0mGAW1CAr/SQAQoVc9VYlOCFNMJegwgIw+JEGciwEjeGux/4uvQuUYT6Uc/A1
0sbo0EXR3weHYjVmGwcaqvC00/c9QVxjCiHEiDInh2PUFkQJ/O5E2lRXaXclrf/G
2P9irLLMujImHdVHQggcmUWTIjglBAjaAcMLfsuTyJ4wWJDN9CuuB1ikdXoRzyQg
QBR1+Z+acwg1RWEuC0+F5o+IEVWPG5kHexuqbZ+44J4vCe9qKFdgA8IZZV0JfTQY
fzdSJEjG0rrCrImnW+aSnu9PFb0JFPR2p9G9LfrFjoX8ai6fdSQLZ5+rc+R9kTRQ
4NlQsikOpjxoPvUpXHUk+i6FBY42uLp/NLqEeuZ2kvvqnUGYXktMb7xQCtuvFfrf
3QaRTSd7ppi20+QJzeH8v1RiFHpvkpmHtHYnCJi5sk6Y9NguQs1+45cVPTdThkIb
EsXCTa6CFM71KW2c7oKOqzb56lXOX7oqosYMOIN250hBMpzXTki26c2iaA1FRNt2
avM0m1GARCz04zQIuCqIyT5XAKIH7F9EGGIAt4mKpWAjbDeKHuW5rN7izIvVjlX+
Dc5AHBiF6qD09VG4zq2KXeCImiEOpoQW13xCiRRA4tCWdV174Z9c+xEqJFNVRk+N
hoPckLUmdqGeJwbU8CycQFnthY8nKkY8GiSFHW7+NWg/5iglguWmVbJYG4Wn5AEb
FRLEfTnlCcYM+8cirBibQ36UK+H73KcDXRKC+WoCdR73+5/CqK8T1YA8yAuE8QSc
eHzrKRul8bIRsj0pxfJuD518x6nrNfgx4KlN3waljmfGDFV1/JvFGYHzRyl6SSDT
JNRipwoFCWRWJscctv/LuOtoBriCeF/yk+fx7vX1ldn9GRju9mlxj/13vr5TI/59
0RjRoLM81VdsxAlzAlIUplct+RwYMlO7H78YpZF1t7QDGRAVhKyVspMvmxJxVarD
Y302z6scU/X/S5CumCtRbBLZfdhKYloMqHNXiZMaOCvNlYcmQxBRGNfGBlYsAcro
WA22KAQL+2PTZvZtqqcAekh/H84t9EHq6w1o2b0UWysq/lXkojn3o6J7umrwxGFF
iTm6CyF1iUc8ZBZU21O5NnWeWiZHVhCi04AH0BiRPg1wfsNnqNHu4CkTP5x4eXpN
L/s71LLmT84k39VzbF8tCUva9DhpmKeiqF9DihLbsGjpWZpRSI/DFWbGpXHDCgsm
F6bEI9kjppdbc5dSQjxfx9cgVdN0h5sPnRyQPPtJvRa9xy9rXd+f4kHsIm6zh6X7
W/xOqhzrxXf05gChWF4dpBiWxZVk2hFoqKgJN+iCps+FSXms/KmpUhkm/B6PfjjV
dXIPtibmXS1RiBdrOKyDKA334mGtJtQ8fcBaLPHuyK1yXHAgHW32vmo/Uatx9/v2
67Yqg/8jJn+SZ91BkKuDoQkUWAO1KXTdcjc7h0dyybB/crgcVWE2eOGZkNdC7kx+
CmFGQElaKmPNg03nfYzvcH/0/X4WVqhALvkSV8jpyck9ERcvNIOatgvirqy9Eacv
lPADHaljYEroQJhr/cd3I4p3gtl7EC/UOX4cuu8aFRNvaoHbCWdA1Z9Hogb2X3aw
cronLWZNpK/r3R8wqEKRUC9JrjX5CQH1Y6qxt1rbbfII1hwoYR7NPq+CHnXRN3PM
M9nAI8VCiph4Ef9dMNsjNCPIzoMaIlFRcfx7H6qhPVd1IY9A8sDZFDOfZ+GHN4GB
O9gjt4B/g0N+GOO/wfc6QvIY2SFZeqwBoOTABLBdw/TA5NSk96G9XYorgotdHimx
7hg/+CWAHsdYrUKDQCs+TnT4vUXljC5f5QzhbydOiyD9XKhY9FMJOL87KW2ozv39
H6gIZP7OaK+agsLFRRYwkbOnkV4Cq778emLlnhHszCKiBohGcrJ2qjsoa97Z7PPC
AknHKeP0EBw4M6rHlbUHQ35s+DDQ/TSA0Oy7eA9xE0Q3B91aidOipD5aRFwCiSgs
nuoQeSxKL817FGNZSvLiZOj7MfrXipGi0UOc86aG9ESBd6U9+R4VALfkKFkpOBlB
0tIFK77PC9Np6MsvO0xlurk/Dl7yNVC5Ih7ZAs30weN5sQZZJ3cStrfYdceWeNbm
nNrZ2OcR2h5SWDTAVOMLf+jMWi1VnKVjM60/q3EuG9EisIOT2yw96rRABT/068cK
fICQNSzL1N9a4SBtCg4T/OnjhZD0uUGUR+YA2CTxmwVciMlscaaoyWaUJm8TbpfY
kE6LUL1dfKlV+5LEWxlHZOxGMEeDdXUj5/fj3IIR/9tpqmqIH8TrWkdxv6gRydqc
hiSSALrcoCKUubY94g3QNbA6tJkcLCSpBgk6fAwv/CmTPG/InHkkuxLyuRRTH44H
SqIlQL5rtpyyKeaYMUjpyOWS2IPEB98OWJfIQyOZhU8+dtMFzTdE7bpsyXtECv3s
RNYgJ5ZhqJ1vw0HhLnbk6Ef/7HSnPXadhYDWes9KzOgXbK3swl1vlq93VDcGaaT5
Mzf4KAUX52pN0dmZVehzOFP3CIPqRIbbHiSVTgdKMCJ3rRLSne7wc0DJh2JfQi0d
dI7eO0tteBBPgt1zwYuEhCrBxVOIAjts4O5gL8qCSYcRyWWp+Tb5moD2QrGVLGVM
h0atGJ+6hXcjx1fFQtR2ZlPh8OlYLf9qk5fXN9t9V2R2B06nhOlc5qctNPZQK2xM
qVFuo5lmKnEtkxg2XXfHm9x9SpSaZ+GHNsh88DzMdvpD5xeShZGpsmGruuonv2Y5
EeHOSUiGTJpaP6FZmT026fwzO5Oqn9W4O6QVLQDmI15543j0iqu9lurEK9uhCEff
Q4AjpxGStRB3Ep1GFnCS3mTuNmL8oaAv8ceBcLT4iiO75JLeUK/yvmQ5tCF+u++l
id0mjSF4O5/4OYtOVMa2IJ5/IVcZptoo8kHAyailaeKZ64r4Xh1qfXvgluRD1clZ
vDir4ox+uQVpFu2xZWjAWaBLcK7sNbHaSs0B3mWKzOAczW8Ns/czA+AGk+CBMZtq
aZF7e8QiagIoFpjMSuUe4VlYJRszIYQ0Ou9ugI7QP6jonQcm52cMVsNRhZ/mM2GN
cU8gM61VOO2DY3wrBLBEQdZiyc7dnTEL3W+NZpA9YKe47j71mHeSGP53828UdXUQ
daKkXxOg5ZHI1slFSMDHW18CTglnWMyO9kRk/rETJTop4HWJUpRzCAQPQwsTEPLu
k/aZ+G+7go2PFC3fqmdu8YJXobFyl/pO0LtjOFJ/ua9HvN6rWdcBvCheaiMLjqd/
xOU5rN8FkVTa6IU4iopG3A8JC4zIwhADYWaAEgMsT88wQ3XGHOEFTtguqdRMHe/4
os7l186YfmPteTt02rOM9Zaso2uF4clUzKr1sq6RPiQj3clH+gF2ybchjUOKCuq/
lNliKedaTMunDE9HiRK95dpDpI8q8JxkVhDOsb4Gr2EQ+56U2qxguT+0rH1gUBDo
N9RHXmKaD+PdFHvFxmdz0rRb+5ScqjgKXIn0fBa33ySVkn0KkAu6eEk/WWJvqWb6
j5Au6oQuEZCdnT1504NItjc4C18lodMPAYQi9B/20u66nQnr68sQrjvE6bmHfe0k
QcI6xEItBUg90u4cCm7MvU/Qeo/RBDI1rEPAJYV4MnZI7Tq1gCTHiLXWBtYq6tvn
VqZ6vOUEqF6vVg1xN/lrsWKUGCR0wEAjyJYiSLFkDugMbiveJaDBFdHfEUA3DE52
CK20WFIDahCWOnGDpnPnOqBI4VO/Zc/ck52393hk2Bbkehp3qcgx0UuDQyPFA4u5
rBAYhspuSfAnBVHoqFQyw80qB1Id6Jx1k9rFcwR0AjX8mXIl6xECuoru/PSxilFz
2Optn2S3DdaIHKdXzrvgqA+Kn8qB1YAVP/4mGHgiII2UJ5b5dJY7BK72z5J7rFD4
D6E+3eDImpUqhcxK8p2qzzLQNwT3OGXB/QhkasWZL+4uFqNi49Fbyb7C04SQrXYV
chboBSNYeCbwaODaWaHVNYG14wo1h8o+J+gv9PO1HpG4PxMGvIwjR7t3AuCjzpN+
HlcYqwT9czAIFSfAz4eAP3Ksx4vjJfKVvHCeHPYNrRBdsGpk07Vpx30Kvuo7RORH
V1ScPWTa5guSB5Fn5SUvSRMQntd7SJVwl8eH+fbAbiIaXfP48yFKJLow4zQ2xB/e
YyvXZM2N1tDy+uLVmC3nIGy8MK6rqgz+uGRiiEXMjlvz08Pg3SR+VWf17KdRrVZH
xD7tPWis7J4RAMEPi3DbqUhGT71e0qM2sxO+8IEpzoafVS4SVNoY9k2v1/wZ1EXy
BhSYCkiAb0DMx3+R7u/7mKkK0aLNIrFHy7RnW9/gJfgi47827I4EZD22kQE+e1DO
J1OFglMf/BsH7ice8buQki0fn3P0CiA9FAWpPI0OyImOCrLWOgc+q5pdVmhGv1lO
CbwzwOLxydCdieHOOAHAfs1d4gHDXr8AEInvpZc0PmpC/2eqw0qPFAYnO3bzGIk9
PEmphPl1FDV11BvVPxP9mi/YcdgefFtLS+a1iXntEBApBQUuLW8WwnJLBjo8Y5zB
7IB7DDsJ9StmlUbdmT27HD9ZuNqlB7B/CGpyXlc6vKdAUV/uiRUIImVYx1FY4m3W
YDpgDo29eolYp0D0oFH2F5urgUb706Meqf2b66skJ4oYpMlPcQLo6fSBoVzHVvd1
nTpv1MOQtYLmJFIz/Qj26vNuxHNRuEdzkcgNlXgA1nDeqR5A44aqq8Jdo1w7QmIp
MZ5pD/X0ACmGphfbqHpCTKroJer4M3Fo2DKn3x9UjbQrZpbidM/sO5MLopYL80jU
0AAQhx544smFB5hLQRoW9NH6nuepX10HO7wyT5TxMgUDh53UD6n2vR7emT0AUtMa
QOTTUQ45fr5sVLEiCd7hBhB1wPuzZIwTPIqDL4TMMz5hhkoKviBQNRaiUw9vRo7p
ZdZxzR3qF8E5D3dLar/pgsrQ7q/kTK6ZJkim/n6+ufOTBk6esDOiIIwi+JMquEVJ
N++0pcEam+RPpmPZZw5GRhDE6g59btTv3QizrJRETfOUTLjDaA9K0f3XiMlNurEh
5DM5IPcTXV58wYmDtO6BU7fDsH13CPdzzRZBS5wdHDff26qj8NnTV5LRtIigyA93
fooy1EcagH/h+dUZ8S1289MrUPqvMpqUJWaY0g05LZQqKRgOYHFO2gRoczLok4zv
57m9Y9tGwi2BeJb+46oWklnLTcrQneZzHfgoieiCriZjEyldNvPddUGnPd0V4Ytr
ADJhrFVm8ZK69eIGWjTMR+Luo+7t0yuTWvk85vCbM2KSHd5s+K9wDyehXo1ZaQvU
En2lykO1mo2/BlwGmTY3OoIxClc8yI4ykl8sAb5tVV4Wt9z7j+b3VTma592Wt6ae
ZNjtLT07daCc/BMqSd7rCd4CMDSTiEu9kmSONIJcictcdLVqjZKi8NFWxHLI8xgL
hhVhP4Uf8FGRTRa1gLDfl4/ud8x35of0byp61PfphtvEDH502iCi7K1u+C7Av+zm
qhejIPpOx5ysggvrO41IFv+9gvAYnrNyXqxhZIpNPUx5K1Sbi9L+RNv0qSfnEVme
gN4/XUf8SW2xsWlw5Gca/BocKFidSzIbVMgyD7J45Kk7iNtCPKto6nAeiLLJFRG2
Usfr8VM97JHrPhFIyzEsUpFRyrGL0mTQRB6sXSrTumWw+OmO7vJhUvov5tNUyCMI
QGgoOJMl+RNFnxc2k1/sIAxiTFug3dY8cI3MBTBxV01PfG+U4scQWKj0cMAY0N6Z
5nH2eMZ3js4pSR/ZQOfjIjQJerh6CnAziPt2VHsraJ80SYkFlpKvk7HcC1/FBeAY
TDAWSe5VA+CPl12Uub28V5wyJ6DKOdSGxutGzcn1dzpTBtdtpilIwdDeXliPM40T
BQTMbwZsJnQIjSZsA2opbZSaMesNfeZUGwAHPzrmY9twylAo2EU0glw76qEwqoF6
GFYCmgPBUF4vJ+zz5t7OToyPSkh2jDbLoXlo/PW0aAG/dXtiI0JzK4Kfg8sy/F/1
4JSmVIsrFNSpgF+aqWfKpkBPVKbyxEY+jRWr7x1YW0WatToEwuH8xYR/kV/5qkWe
b7D0uQQRr16JkhoA0HB1gOC8exjYC0YgAdAE9NPcD3ytgIeOfpQygi4iJQg3+qJL
150gtwuJ3dmSMWwreot9L6d0i1bfowI8DAYsdybOszVJ5+N7Y4LrXWHaDVZRB3H5
k0oLi9XLB/Cpi5onRxS36YbQif/wegUZQ7WQa1gEbTGUJ+h2pPXufEXOaLgjrn77
1m5NX2F182IT4y9S2TojbRLWIQdY249WbSowWCQA8//zgHFySTXbGG2dKHw+zaoZ
SEhl+jIiprePDka6MIr8OSfVp9lMOfj2SO3iNoDUj56F5Fhrn3/P7/N6fkef+yqS
XDVOqe/d/YhQ+2ZPfQ5oFNBtGICcJq7FpcLePtf3mCTJI9gICuHTU/RBmyHYfAPD
AJJSPjM7mhW5CGlj11F/HXDjKVHdvjZazAgWYwlNgI3kWMpO2Y0YG6uT/eR+Ly54
R03JgxWa0pZxsdov4fXdyKNVOdDt4R6nWuwlVwQHZcRBL63r8dnljYFH3VArizrD
fVEcVru83yE+A0qU27ODsTNIS9LQX4APvd9C7j6JUUPQvYLC6YMtFberM5Twz35V
nQTv6u5oyTAJt48WP1ymyWY64YqFulFb6gRZevMFzhZD+uOK3HoskxdWRibkr27Y
qwP9YUlmHRvsTcXypeBRzMwYaUqf/NemDnfxWa6Ct1lDPfQx4mK+oKs5YzHt5cZS
4jmziI7FCXAkTiWYbO4VKfLmWbhKaBbYw0/rZqZ4DiXryCyv2MwkEP/Q8e7Ofl30
kSZSlrrXxLrPOZzBijBvvzfAGQFAwKUd+2U5ZehR/TcZ7BHMut3u7yrrJaImqFxl
Q89Ug79SW+EAaHqxsYo1owYwN0FX5ZbIG078jx/88zsub0Lfn0uUMKAcMI9uQFXI
FTbc+j26GKD2wG6BXHqI/W4t9sn6i/eKCCt2bG1ivMcK3/8lS3wZo4AyMKKdPazD
+KnC69Q/1YOo68Tv19YkT17PzCfN24eUhS8vyHy2o44l/mm5jOkrxMt6kr7/cWHW
QnIMx+SAXUiqk9cd5BY2Va8/r/FqmOFZpt2HRHl7M+UpP2N4Y9FEjBz9grqc9kFL
Tai9abSDSB1XrAJp3A+McBy5mHgzVNfurZK+frGvmASX/0fycUCK6EqXN6+FF/d1
nQ6l+3O09Au8jgAkP+jji7PI1jzk37xt6NnQ7NahtyRQtegsQA9MFLsQOSm9cB68
boMizY8HiSM3gXLyQM1RvCap5LvF5cPyYJCFwl1x59M72Ak7AkFRPgJVkHRRe3MQ
3UJ4jLraVUwsv00qN4Z+lrva2VvabnB8CWbBURDVlLcJdEmNJRF1K4mUO0nk5tsA
E44te4pq6s4FaE0Dq+027JETxj3M6T5Bnao3YwZi1ZUju7fiv3KptruGQ58Edefl
NErK2S/JvxxXMt4vQ5cW49D5us+cMZ3Y8aTEtkLdmb2cpiTMlIaRp7x9re/gbS2w
tshQa7d+epGMU8mS+oFqr9P8T4khWtbZkdweZhwN5HkjackvRDXjJ7lIeBNAJbzX
KSP+XPsO5rB30G1I0Q3QsDOiZXH54AC3Qy/j2GqZ/FEelL93VTTfj1ReRUffvEgv
HNuc/TrLjtPsZ6uMmkhIr3R2fLHXAEwbokkoQz3/5g9/5PLwuAK45VLsRGojCK1v
hVbCc6I6mrHa9VZYX3HRJ0Qct17ZVeJCWDNxjTW1pc337GE/gGB8Zz/b6MfwVV55
M6zDUAzQYywrhnCzYKYObBVe9rt9zk6xrfRnFAhzTaJ4AJq8GrZyN+we48MXIGP9
GXo4LbsPiUf7Lhp1VoGYLG+GgnIlzFd//rEWw8SzF/Yxr2WJ9kzLHtKxABLCo0xn
yjjDXJxJap1AaSCuADxIh60b5kPIhiceVc+Y+pTuqIIOnE82mRd4c7aKfI/ols3M
/8eLO93CmHeeHg9tpIBMdxzVNsEsJdg7GbbcbhsfvO9B2+Sluaf9VRxqNhUPWl37
ErOMrt7w8V1zYXq1kgHDyKbHA3v48pS0SXiypiD83x/BN9VZs8Kx2G67ANpb4zQ/
Cj5wJs4caYdnbGkBYcHyHsA2J+N5IpO737Wh52KolEszmelvFDldkPdTG/QcfJ4P
IhvQYmmmF+Jt9KHD5oEPAeNlM+BQT1+RBDHQEDreNtoFyV6nIMQcJu9MKfFz6jQz
GFhY5caQEbywFs9roiR0DQVHxcQRp8sgxSM+fXGtsUqLu3G0q8PhhIVS5+9p6O6y
CWA231qT5JIcWfTja1jimcQ1iHs5/IiZN0sdaBgg7rVRq0b2gihQEGpN71E5JJlZ
2H2kDJ4bPMkLhbGNwAyNLrg1XAveq4fjQZ4KRj/8AUL5EhgoZK9CyPtuSqIbTKvK
vQK9B7d3Q4TiyeDadeegILAzitsjJdVMXJfJn0mJOLB3QXix56/cUS91s6YSwKGg
x/gklgZ6J5PTuNmif0teogMHBxuTbMCl3eDiwFoLZCCotcZOlMyoQpj+mCXVh1RF
+F3CtlLm2YRC4RVjP+fnM7QYNO2j4Jz+dXEUqMgTRka4MEAN4cmYlvij8cNAtJuS
TFG+PAHOd9Iwr6rKvgrUsNahDq2WV6Zax+ZpGOcJFp8eN30BZnyMpNGy57x4RBW1
2PpS8QlTSWXlegoHP6fGQfF8M3rWtLnWz9VRhfenEGpYJvRr8CDdpG8pcfgBP8E6
RiuRQI0OkcyRQtl7FyJFilvLcChJtBJRsJVBmD3GYdpD5LmKCEnMx8KhSxcY5eHC
f9qH6pbSza/b69D3SOKpvBP6p+ug97dUGzC5ix26NnGNJnbwaQoVoy1TxVJCZ+zW
rQMPqe0deqsZJACVJTtevkVrPGbPcmt2ZjXsDh1/avuRT5HHdm/WmboL95B01PdX
g1nZoQjMTYhPCfcGUNmJpwQNmnuDzV3jl0ReYahcxrtA+ld/x2I2tSDdp4Z5jssL
rxaeL+ZX6+8N+UmzUjnAk+0VhSbdAWJfdxlmfDVPehtzoBqxn5NiyhiSxViwcjck
QwLbmFnne+ApXxBW3qsb2m61e40rZeJp0S/ak3zyhfJG0TfsThbMPJkS2ddJOpBr
0XEdX8JO6F1M3dvRAyrCyp4fspLIgeC3GwaZPHNYafcuhWgWZ7PxtJkYLP0rjiz6
jxGKvFVXpLBgTwyUBpX1IQAA7IpkDT3m4UTtp/YeN0pgv5+iY+P2U26GvB3sbfp3
VWZHV1FEDrLYNZRABvTGRb9Ag8faCsMGWWoniBvSoqVZOpKuzIpzWrQx7F/2c1yj
rTe9wM4f5qxmx6U/NS+uXZuxlBJzL65SKlCa8qmgsvcOSVtfVNCF+rWw74EfglMa
UpnUd2AiPPeySFeFQ0+bt1uc3M8pMOlZzVntdltfOS1A88ZTq5vy4YaBF1FFLZBV
nomDfZeiRjUT5gxv2UPzuSHBL+zXn71egU8DPbRwVRZU6e7lWdNgZMO00G8fSv+d
1tRx0oCAXN1h7K0A3XlcwyPFzHvOdAQ2Y1nbJW/9PdoAJI2XdOyPpMvt0EeiXxp/
yAh2KMNybCUui0W0368fFr9+FEHj3LMrSVkvsqbZkULcqoXuIUI4xmfTOeqQ4sPB
n/dep6HCiaU6KFaPvSGbUQirf6pqtsWGzyTpFQiDImsPzWR1rXLzr2RFZwbMPxF6
BVlmRZXVpGdAuMBpze6y06yehBc5cNsUp5lz7g9MV4S+vLFkDGlty2laukx75vj1
nWK36QppMTOJ2nRWhgHWKuL8gqzE4zoTTc7bbLSMw6A7EE6N23RUej0GI6H6sFwZ
f0/xWdIOpr+h9EOPOajCz4xZDlf6ADKUuBO7S65T77NqYgtEQ/L72hRFSZMBI7S2
sARSXyzuz+HrSK3xplqzPO9r/iQKnYZiBQsZPrpahjtghT1FRgh0zdKoDdtinBKH
KaEl7vTBCz380EsJbfMd439NwXlV1fJBJq1Pu+j5QrWvCAcZMhN5dN8nV+oB1SHs
KOxl/+SISowNIgMss75zL77fmk++2nqtYfaCEvHvvPekRuVCOKPCzRLe28FXoDB8
AAExaREGCfm8TRefe3HQK8LQpF8v2m14MvYIuy8oFj7imkcXKa2r9hlRaqN1XOjl
survHgKm6D4xMu0QJpDY9O5YNNeXCZsk+6Y6iIrSRgm5BfTF/jaNR5hjV6EtNKOQ
Ubt1vNz+DaRdtQBLLaxLQbwYYHboeEZemO8jaqgsfcYGLcrnVAe3EPha1tzQsp7Z
3YpnXutLvONeSOM3Tl54l3P9wvX0BOCkKrVlWU7SGQhpRY2lMg93mAog7Soesjfa
QvPfn5rcOd3Z/h2td3Km5qFDQryqtYrtIK13+Pjz46Mks48fehb19L3oeiDp0GnU
/5rKpOAyUZMjhTGO+Z8rKTh1vJo72eKokAtb39YLirx+trV3ePMRiWHdlyOBC55G
sQaniYga4oSl5cKsJPPaaVAeCVnw3vXdMnfW4/Vs0HIVajO1s/xWA3gXIvpYtrXf
OhfoaNjE8nOJWeDjB2DB9XnKc6MHzFneU44Gqk048PN2uKQo8eCjui2tx1eTkwNM
oqLR9K0ki0RGsMxVj0iv0HOp5P28I9Yn3buZmVNPVgLvY3fEVqbTSbnKIlXzPBqf
1wU3B6nmXkEgzQBX7IuoZNCokdTxCTdToHWYNzjmGfQwGv87TQ8OnP52Ivm7sORY
kxBmUe+5baywpjOXbFVzdmipnudUcTI32hOsc1u2WHsAi3RsMzUcOQiURXu9+naG
hoDsw2zGInZXPkxJa7fbJHZUICuLWLAkVymR4DGFufksqIIFKZJF7lVBQPB4JvaM
Mp5si2bPUtPgFR71K8up1s6i4ZEvrV05DXl+v4adcZJ4v6QfH3UCdHm1PYVyj2LY
8H9w5VcW+ih5M5uTK9/YOhyLY3NtOtwuL/aH7YfN+WLmi97BTtWKrgs6YSc+0m/M
VzRsTt951QRSUu/IspeIDwTQUwhNttQhlplPrAi6IrRvBAnvMFHtMmyPihbJtPi/
j0T06QOcWALLQu+NS/otpJ7z5BSo/dnln6Ssb6T+wXE/trSeVZ8nLJFwTX7kNEnY
eY9tkCxtMj2+ostfRENLmI2S7MgzlQGiRSsD8drxKda8cScrSAa68efgQljYAWjp
71KamgeKi1jjhbZ+VTpzF02HpnHce0GrF3Oc6NYnWrHutPZ4SZRo26yhJSpeQr0L
5TCixojFj+vR72PwYzgCbU4z8Tn3vH0JxOAGOMeMRXILYx0a9W/8a1eHn0ciNCeV
+Y96cCewzenVBpsQbxlCSP6MiBm08vFDEB6ZSL4t62PVuUdQ3EJ2WakoCyXUM7Ej
T3HD0UTtXT4F8aMUMo7TI553crnTGsdiL+S5/4h3l/kn45Bh/vny75n8c+KF511i
ZstktDJaHcM9lF8mN0T24PbiNoe45z84koUMvZvuAg2LTf1sqTEs+mCePeLWbQ+0
WPA1O7YnC0xyPE5UI0GSx42rFC1Shs9ddNjLJDgtNZWrORtWmsUU6hODPbOcX0uG
gmWTvLMe3PNIuTUQ3Au9ITt3pMR7ZswOKTd3DJtKgv6qtrjGLiMw98np+1Q+IcCg
TzMQ579DputhL3El0QAuDQTQtVyjANlqtNqUQ8kIuT/amD3G1LXHZjhjknAF9jaz
pwT5J7K8oY1PX0P7vHORcyYhOTYK5fjSrCQyiqciSoj3CGvtwtpHVoMKyy44WB7Q
MwqZwYoThaOPzpxfpGPE53JHMARbP0rFrpMhYJ5je9dYK2Zk17a/u+1e2KXQubhx
9mePCqn/aERmw/GJE81hhnlGVvwFXoysty3MUZEbdGGQIpcfZf+OCKkGjvPfUcE8
QNoshal7Ll1YytxAN3ycQAi8iM+MegAmEt3mh59HWRGyCAs2A67ljUjr7GB2QK3R
gZqnzt7xgHOE8NJxgkMdJ/tut/sCQsR4KKRfGBpFbsAnS7vhVn89KbfaCuEN6AHl
+JeCqWEarcC90ExQ3AFcHe7E5qqT6Ekdtnje72bo6vD7JrtFuCm/dFczq2SU94Dz
blDNsmi9Ou/dL1eKxGJukB0ba7STAEDXZrpxCz/OMe/9Qtj8LhogZn2IPDF9PGza
Ay4lgTg53UMX4iHFiItjVd/vnU3pc+tcD4NDIas5TAmvlSn0qhQMp2pP/JuAssFL
hJ2OBg1wm+Bng0/rC8G81D6w7r55ZuL/dSdOUBlTSpLeFG1WuMxMj3KuWVn96iOu
IsPoFjzGzsUf+dReZPFYSS4Th/SF2D4lB2xu+dRFNhlZNMD/OcrVcqL0RHwg52NH
orQXFaJhjjSotnsR4V9nNxl7UHpyrrL+OKWwp25GsEfMeLAYdFJEtZYc6pJsawx/
TFBAtwWR/j193xGyU4Gp5GtxK7EtDLeCZYTXqY0jU6DAUDIW02sZk6dZTMgKwaSd
FTvkDnj7Iq+fKQtg12d4Am6i/IjvGzzqj58DxEw9uk3BFq3m/CiCwCEIXeAyQlhW
+UzNRHM7qyXZ3nyaII3TupbGXUeJG1h3RUCag04P2jhG6SZF1CYXp4oJs3ANjwd9
5pJrJcyAsc5xmJyYMKG1vOmURn3O8Fa1bOg+fwMRym3DKQqLyrGq7XL3fk2G6PpG
40/UXI+hJGG7O1z2piluBQ+qDseHO1kCokubQN7k0jGv4vDp+hV+jjfP8My2CGjs
tpH8IgHJIe3SY0imHTOqc1Wzsy6yr6A9Mn844sBptoTcmB0t7G8pNjiyszQdWKdS
XYG9g9H7Kb83GZixXJeAIfl9UmLXtlvTvM2zP2ojXTfPs7n6CgcWzfbc3nD1z0Mk
Bf26CR7qFLvoXv2h3xy51fn67x9RWY4FCyySiMiinpMyZVseadM+yGkQdKk8McNz
CwudKKd5AkePK1NuO8apT2FZavjbCrgCzoGpkVL7mLk8P1C948G3zW1Cv0cJx2kd
Iokv+HOYTBQoe8kJXVOz1L5f2JjRpMgIEP8AW5nDCfqVGlXbMJQyUf/MBpcpg3OE
qvWlEQHN3kgZLlckqD4BOGBS+8TEegAiJily8NaF4kAd20dqATGhxUVjV+vbWjZe
AN3g/L4OZRgp2EY88u4/doyk8q5w03IvfdNZWzI8ZqW/OE0G9cmVnIm2hWTh1BRL
oc5F9sxji8oSUNyETio0hJh8qUeQQEHXLT8rn6HhMYuEL2B1dhxUOfyfZLRb7QwD
O+hhCLOU5QAIPxoJP53shcan3Ua6GvV3rixew//YiRZ4WqASLbWzA/P+9jxPPqcq
uAQw0p0LX4X9AdlLWhAWmlzd2lcHrSEviyTJwAx1RGvJaeLpob8ZcekeNT74YyxL
Hp7FiQEp54Uq5yQUpPpBinADBjPURPjGCUMYbqOQEGfuSoCCeUGA8WkHU0zLjFOl
n6ALno9f948YgckSQbVqGM6HkYkD2gViq/DjP5A0jaEcjFh/O1AvE3rLSl3RlevP
xsn9iFgvmxYnGHgEJQtinULktGrabiS8B0NyTFlLHy0CvGDLSJeBA/nsmNzgOFir
MKrPmNYDFe+AaoxFt875T1ZrzoR3gtVJkAao50Oy6vkszn1IyiuMcViRdLW/KXl4
T791DMS9MRWQMqtt7xEG0sDIw6UGKg7aqX+N5oUImhc+GR8utfJsPDY0OWOrZWxO
nKb8sAdXXEs6ibWQO7071c1xlF0I+eF5sfyo6ldrTpc1GuuMSSrnUjnw/P1uTEGO
uQXGGtsRZlST1aCADt4vjIAapdz2LgLBVhhG/abwGvccUwmRRxhV240wjJxdOWIo
SbG56peujs1oFMGRqjsm/NgV5EfB1V2lQth2V1WxkV9bDk5iiBoT5ukK+J0jBM7P
Oxddw9Rj7dKxVKL7IoqjRPrFVVN9wU5g7m3r5vAuefOoY00kPdiLwIMXlx+4i+Ho
ZJ5QtsFA1tYs1XgiSUaBhmMrsEwFXrxJ5HLHt4VuCnaESjEu6toGRzFdM4I13UDi
9iWRNLwRUE2lPDCHGQfVxfUYhUUc4Lhb7lkl6W3EZpOazy2TZmgISvDcFyAbjy6V
ikC7pXPwoO92K0Zjw2gzfKFrKWSVjWzWRq2BidktUP88wkmNVVy0N6eK6dCBmecj
dyxw8K+dCHPQL/PWGWLCY/tGUxMcKmHqeIhaWxeiWDe4Ik9WAGGmRGvklkaAigKJ
ZTfBddKRKPeLp6t6vV9Kkln4vbXIfGIJo9ByHjnBGxjczN41IsesRK3iLaMkLgNE
ZI4ButGKiayEGdm0FneseqJamt5NwbtVJs2iSwhqA3c7MTLn/FdERJvrvGZ/HtAg
8WwlCxgrr6S7dEjhifLelbOj9g1MZes0Iu+zhU+DBycl8tAHLH9sYos9OIoFyHl1
UD8KC41GwWv38Y01b8d/c2cxQv5aiLjhanTiFaInQAIOaQngmEvkQtoJmmOF8oSX
ibDnNEWPfs67K8h7zAv8IdP5nBU98uGMdikArh/JPf67MOwIdCe04yJ/kuj4TXoI
lpCnwSWrPeoWlaooT5v7WgHtdqwhJGXOO8eTkFTWK8y+c49VPGueA7ytxevnhkiM
tmQRtwqTUU8xvNd2KTBUXcO4nvd6zCt7NJ+CzPWCJUhbJdSpaPp4fwCQgfA0EeM9
7Q5oUCy4zRQME50ljaO7X04HCEB0cKyxtspx6LS1eoZIlg/ys/YgRemqZylO9yHW
WbRKL7B57aSqCnIZmNlSyL0w0OJujoEsM80i8moXg5TQdIbLC0FhF51GanjIbeVj
SIJEMivc0WdBnRaQlor8/SXmiQm0ij3/FJAdWvGSfgtFUASEqqBRNbmETaLGN77Q
oHJuLMqt8cF/VbBWIbGsYHtc43ygxUGEpfsYPS3L11dcjaXIB+cltJD6WtbvRAxC
vYZSki86n0MfFhgVTuj0KjPBnysmhSEewCn5i3dH7tqUfMCy9AAQ8KB5wX4IuVUW
4x0T7b63PITGPYzOau0HOzFV4MRne3+xdZ7fm9KRBFyB05+H9Vd9KUBL1Q0geoTC
PXL1K7zoCAFDyatUCBemOIGfQ30duVz833wF/jHSeX6fRsXmnrMaXZlGW0QNlDSS
2O6338MMvaOtEAFR4/682w1shS5JuW6nJdiZMvjs2y985YV2iD2phymYRVvxVxvF
VUp8zMV31G5p7PWUc1ZSmTsNIfZ9FUbhw7oikx4sUoOKvGw1Mv5tK/EgDYk01/bJ
TgibQNVASirQCQgl7jn2J1MK36y6wBkKuzWF3rfTIcyUvLfZipoUKaHSROMZiaEd
NpoRqbri5iIC7VemdMqDBT7DctC4SAS7q2mKoMuTPiky9WAXAshHO25gPZNSyGhe
o37A4yVRzvbGJp8osYREmelwN7jV7WljGfpuHBCUbW3JHggmS8iRL15GpIGWXDtu
qfXoFxxMA2VkwGnC1t8xvkqh6pbG2tQ52DyFAs9LNQNwYFP4N+5hf5ZRdU9OO1qM
ART3HHb38Vm9pl0xP0b86WF5qrKy/0RgFrHFJpeX6Ycac8qcZTiXNnB25nUovxJq
Qv982WqsY9VrlJ+AVp36nkb4ceMMG/obGdzMEeiMy8DemZfD7mzhiaBHTnwugene
KSg6u0oq5K7Ekd40iI0fcBa9iO1/LKrPz8lhyPvdXZjkZecSPf6jElEdWfLkVjx3
/yjcaQUbQ61sFWUBMlEWKwDRLV9+bWruILKJvRQFj+AwuBHq2HjpanLke8JZopUP
4e+vwgbiadx1qGoKfqnIqroJlTJHCyuH0mUhSIgSqXNRW3A/+YPF9q+iP+g/O4xT
soYW3ckdhvWME5BxWdNhkHRYRNYFq3izn4r066MATdCVg9IyGJMQQxVSR1ZEEXqz
5luc5q+zAnJiXYOcMoL8Pa9+dXSzwqF8W0tvBekUCFYLVZxsy2rfxDIsS87g/645
hz7y4E5dTufsSbkCS3j52V3js8ROx+hOIxtiHCeQXKgAMU1srAkTc8KTFFNkLc7f
h7AdPGRs0NfS+e40KAQOFBSpiqZSl5/uYJJ53wa2eIXG60VT6uG2dfPl5IfOVREx
RklZGw//y4BmMOrD2+Y41mdQzCCGfdsdke+98cUMYtdem+1hquEpdiAKvyE+1u0q
NzPkEgR9x5dqe5Lk4oq6XbbPkXHDM8Cnr97AGjZFPSmzVnZrr8Pj3F4HyF+lf3l4
Umaq1XeKZT2hRQTcbyqQoNipJbyH15wGtfCc2rBvaAZ16GGSgAathObNpgMSVV5w
sa8R3lDZlSSerJdUoali6PiYNmmuR2IOiynsrG7tfa+fafRrO+q9qG0qgkh+FUC/
ZCp7MtrBYiTKgVsRN7CWXzW3AC7d/B5GtukoYjen4xHo4vptku830vxasNerZYCN
jJ2uEOLZR/ndpL+RGqbI8gWAaswPS1bAC9Rz1RKrlHQzHzHIm7HT1bUH/WEWgCeQ
6mR5jgxGvLWJl/BJ52GrcuavoyxEfSj6MtTK1+q54myH81GNckjpiVPlK29pvmF6
kvJ8viWl2QYof/HY5R6gcyfoG9BXLt4DKK8wL5djdYAsyPwKvIFsa/IkKoVerYdz
SWGZBxOnUgC2EEL49oEIdw+UtEEdGCpW+ZKIqlznuyfEhO4i2XosfSFJ7glmg3V3
warVRVyT7s4OZFnlSyDS1rKIICZhO8sfJes38DFAQO++n1EHWPjGQ2Em5Zd3/C4Y
F6wbghChLg5vtVHnxYvvnskJuHJkJdfN/SSCs+IXSbXyYD1Xnfci0MJeD+9Koxbo
NOftPnc1+6ExLH/uCjWiHTm0V/LngF2onv8rSddJffgsB04RxqkVrhXnl0gOY05B
meJLUN5dbHabLsv9F0jukfxt13Fjk648OW8faMWHNdpxBCuH4Eku1zjlN7Y5XKae
DLclHP9P0CslOiQlEmnP2K6VwUZRxjal+aCTXAFkKelmKiFee06syFotOIenlHx1
YyMB3T+e02GHgenSG3Pm+pIp15N0DFaPOqR9yb8R4lknGpscuauVCkze2N2AbVIq
eNfQG8dt6Qp6d3RG2HZLw1d9fct9rXPs3sl63fVp+ifvEwIKz8jb39QED0CWV25h
yGB2kooO+zI3NM8KETAcfVLfj96/awRXv26Kbr6eF7iOMFqASrWGdFsye/TQmGk1
KUNzd4K5LLkOeNbJt/FbH9MGVnQ9RoPj/AumWycKemEYQ2HR5DDJ/ti9ZTV/nBwz
J7tdla3KdDUVTYAKRBcMJwDQ+MHqcJwWGjSzftHEUPs6SFBUuM9QLCfFf5TpY4oD
eS6TNluvQ+6K6Q0U4brVpiO4JFhkoW+2CN7BlemYe/gPxgO5lsyXbyBkOacHbzK1
OVRuX7jkX0ciSyUQTpu1NVZOSTbRNd+o9QvwQcK7pQBuopRzF6agZ3t7Hc91nk/O
KpB6na4+csjbhOr0rcoDDJZW08G/cRDAA0/UQTnJQSpP4dA3GVyf7mPUdQbigiTp
7GPFoThIDfLrvyv4kvTT9QYPx/duUQUf2PWnG9gJsl8h0wgBKMg4sjhbuOqIZObF
/dT4I6Os/a0xXHdw4x0JkK4gilqjLUe6ls15X10iyhjTwu67OrX/dhrwzjKCkBq6
nUCgk0zztjCXisbb4jnCC5NMT7MIgTvnIPbiQTFWCFOhBi+qqwd2o2GVws/284Yi
bo19g0PdRGG8Y6MR9AXx6IPJRg7bJwng/TR4gTkeQz/RSZVtrM/acpBKTjBNPfJr
CHpWp1JNynXgsE9j8kjOeKpYPYjsFq+r9YemcD+HOchkzidydURnGVCNwbMFImE+
RAWMgMXGPP2pBt8ZM6bF57G4dK9iTV+9kMBss2YRWQYEJNbSajnsxOWVGm1sgdhO
TJt4oa5IvnBED4qUpXTOXcWUnHEbyP8MzRfXSLTWmzt0QztLielBQa+rC+D2HAjf
arWP74CCv3aQBy5Lvxecn2WauslpXesO5/GuOXKUv8AID5kYmkviEKwgGMQVckp8
dxgwr3fQDqXTLRttGKTaoXm026Cekb+FV5Fu1PRVj4xlPa6Rrc/oh8y7eSNrugr+
HP4gMt1XAJ5wf5u1GsL3UyUMti+h63guaG2XgRMd2qq8/x3DLCWuMbfCr8UtPB0E
4MyP9X+2NdqIPFX1PwRfLGQNCDNbQg9waa7cpNILZ5A0dafC/qJ1l4uPXQ3fRTi1
rbAQoAAuDdH1PQwCklzUY2PqCkaB2SbZIp70Gjv4JLva4mHopSrZZ0HejvPWspcM
KuwPYyV0YwzT4lg7RVl/8fUFHAkG8rLUqVDhRkw3rGH+BtE+zEeoiwCf3wqV4tJM
HOUv7V1gouJ0DmovSWyPZh27TyfmEfg+yOYvA4dE23F1hfgP3pSXlBi1GN6TSucJ
971Ph0e10W2CXI0bhr3Z0UdnTZ0l+QBDH3ePwumYxs2UHHHKOaa19odGcyiGlPVP
57k8Q//Kz4FqS+L3CkPSMtpm8KDy6gxngYYd+QEPv08ha8pTkwxYW8OCTaVpAKn7
z8l9hoQr/moYB0lI/NMcD0Js3z1cp7/Nw0cM3LEc1LErepFk9a2/RKifl/g43fLy
zN6hAqUa8c6+R6IpuFUapybs9Q1D9PJQU37V/Hv4U6dMiy/KcdgqFO9Om20M6bIe
f+/D4NWO8wgt4YiXViDY8faUj4NADRuagMUreavoLYDlTNrbyrgBZekr970k+zna
5WokTpRDcp11GPEx3W3oxl5MxrcF4inR3aKFoUhYpLWRlCHCFGplTJVh/OyjMWbk
l/axGHfihTfWLbKjtEte/K9FUKCcpIXlvBgi3vfiT5w1vnQkC14UTZUDCmj6QbCA
k+RmiSuifXXUEGGeu5+y3hxNuEtsMVhb4D4TeKm57mJS63qBn/HjVimw8196CKv0
mvTn5zztk51c3hl4+I9VdZmlfDnfp+eVfQi6pPaJZfts7So2/j11COz+8OdgrXBY
Q+Ae+5tZw/149VkbHStuz9C1KOnTFZlfyN4yDNKQUSImLi2lprzd+WInDn+rdFec
1yKgrsFwJqHRh/IxJmCrCxkz4mmrRkzqrjN0BJyPeTDljuNFHig1nUMYplS5/HAN
TBoYTo9PlqNZeEm+rjWjOPehc6Aswn2wjSEKJYzioPTWlCW4F2tzJuPTCITh+oj6
47OBSjcbNTohNd48KnUnlJeUM0DpKqbPhIrKqZ0e0c0g6kQHcePzh0vn3ZBeBJfa
91ZleXoBLqOMjGDImm9OsnLfj9gylyXNGwUbx99ttaPsvI29vmPpEaZz3kQRq+56
jPWhmWwuao9pbpTDLA5Tpjv0Y3VIDJzbscxqNoYKqCAYonV2U6Oeow2IGsBcerMB
jcPcOUH1ArnRtUK7z8Vi6QZyJRE4ry3MuY9VVNSLFZ69dJTcMSAeo5J+7S9RGzrD
+9OS72CIKyhiK8k4RGqewlPziF8KJUn836izBDc2VgDSjb86brwzt2nItu+KQb45
xA6FWdi88c0oVyPp1++BThYcCW/vOlmrs3qjOeuwIV2BZ5gET4H/k8BNRueU6YXS
LrusOo/QtgITWEcC+bF3jh8528aLoahsXaFBWTOw2h55jQGGlvCBuu4bK4nTEFLc
Eo2dsJ9kZyuDr4QPnXKBg2YHCy2ikRhi5klsOYZa2jc43T0z6Ra+bcDs5zx6mYFX
JUKJnHXFGtYBJtWvdHYPmL2taU+uGW2OKAIAHtNtkVFPdtKKLV4lXS2YYrYpDGig
His1wr3QXHSKGLsCNbm0YCdeeg4GcdsjabtzAsuWjXOXFkrNJTntKjwRFM5P27ww
YxjI//n05bXLsIxPKyIM28CA+kiYYrlDKMFh8xwjKkcbpCMYIWpebthqXZzb07GW
oxbd6qv59RPCwFEoi8f55nV0X8YgUYbP7vSoMURw6lXvTdniw6JXVXPNtIjr9/3p
rkAJZJPtScp3Po7DDM+4R139EQkWSlidDN8aDP5Sat5cuDevzkXV2YmsRDkiWxyL
ZDs8XPMXs3EhYHxffegfMmDf501es16k9hKI3TPWOH0DVoGRtz8KvenDz9bubE+x
4BbSCmaUExsMPymdaLuhhoJQoNKaJLblElcHgHR6osAFzvxQhpEpC0x19+CWtqOK
ttbo8AjlfnRfhYxNbnS/ry/n2zD/qvQf7kxb5KCBxCN8GTi78Fm0Vo21sH0bSR5j
DYRABTVIaS89iG81ah6GBnNwmmd6IYjLAfNtiGQxZ89PrMYOtKH+Lskxyqtb7scy
5xMGHNiGYsSy6yf1pSvlHyqN21fdC36Qaw5GY8gEthLp4wIVT6ttVdBxaPLhbyN+
FO4PAf+7A7wIM5HllDXBNU+FBLP9jRzI/0ha7BhGTVad+Kvvz8MzB7KMyMivBUsQ
5sMd3+/ki+JQfqQzVA73xvKy5K3M6BoTq2taC//q9b2PIsJqAOJhdI3xwiHOqlof
h/7jy3p8Jo4a9WERz4hliF9lRF6V47dNXt19hf5obgF823b5ivQLr2qlySHFT8+F
8FWcwkkjsbOZ07/vMEBUIo6JioBy9MrkEblA9lWsgDLws+41nhEoo4W7R91zreRP
+3FRzMcaxYuCTNT4aVIUF8cVreJFEVyvpC1Gsx6YslULITXAASBlPQT3t7wolOZX
Wjp2U6B1aL5/iEzowd5gu9QsChwKpIZQvSEvUls69zsaUbWQk2b4gt9s9Gpw+mGa
V6A/B7q1AVfWDB5Kfu4J4if1N26TEL5BAUG7O+HR+K3t4a97I6SsLYXdldAIg+cw
NeaemY5tDyEmDp1ve57iRy1JfT/rpz24wOYYpi30Wae+/zAPCMB74FmG95Kh58rw
d+aUeHa+B0Dicucg8ySiqKKSRPULI8bi/aS7KL6Hd+L98mWkjFgXvovesD6e3AOp
1Z/SdPXM14FXRfMEY+Yc5OR6kEqCcARr1nhVQB+X1tgfu7mCUHFdUc6E2SRvPJrT
eRSfx6DyuS2btmIpHO1mZP3uA3Tut1cmuwPFRGxb+GqdAVOYM9+lO4f76VAKFydN
ufoThZ17O2iAMvnceLYrV30VHzdPaHeVABaO7DKKxkjPTiHpiioKc1OayMTqbsyy
Df6Wt5GYhSv3iSv/FkzOXEiWs6Lwi5vA2w81q0LKJ17euVeuvBAvFdBy+vPhyz0I
zxH9osJllDXumRLCVVSeQ55ZjsiGJ6us/8L/Xbzmb9ObswSjN4Zk6e4hgEttc2+f
ohBzfbJTBSkeEXCDr2oLPfpf7paS02G1UjWCqg/zPhUrZgAS5p173FU2vbJFQLVn
fbMyH6E+auRQm9JiVRpWRPijDSnxzu6K1+Y8+3INX7nBS4tFC0ztti3ZA498ygMt
aeGUHYBhT540lwxXCQV9q6f3a2/DRBK1KpMGk92USDrmEYr7iFKISgas3/YKVgDL
25Ks7rx0pZbNaGo+gN2WhEFzN8tHVTy3PGGBoEHdq3aNZ0Xd8hZql6eJEO/r0izQ
m9EQ4o4PuvId6US+B8NgNx2re3ugLIsplmxYhzreQ900NLzBtKt77wxvMYD15Dzb
K+5a3EaDYCVCeYl1p7d8ds2UXf6tUVKN2StiTwM3k95bsDYdbzNBYYPHw5jvhGIc
0iElWqaXkDo2iKbDHECsx+AG3joN1BgYGcflO9/Qy8qIJfW6ERFETYf+kpb1sTc6
HjUMHItLnx9DM3oDqCELLk4rYrg44/WkzpFA0tsRveEUKgU+P22eYfGi9lVXBtSk
wm9lHAFAkFIUqyTHid4zn8+aB9cqo1K22aTF/YTQytEivDfBNDmNO/f3804y8agm
YiIEoWFN06SdLnXeb+BQMw9BX9vy3tnZ3sX2GUnzAENM40qG/4Qk1dlOw5Mb03WV
krC3CDKnRXpRaAEOsj/dinkeh5G3t7j5F3lXC2rjr818xauWViHxJAaVajbdZI+B
+4eYYEfGYReNRdh/4u6yzLU4iW4TLKaQN4q4gKJcXdw8wmR2C9NZdJ/jetzUUwUk
VOzRme4ck/W1tdxJAt3HciB27thjeldnh5Ru9Kz4qNTpclqF/hLZCehgxIulZt1Z
Ahsd8N6B6CKPKyrSAoVLvlqAHag2x4mgmS4m/J0cs0rMZEemUvqca9zPkcQWZY/A
YuFC83fUjXNLdKKG8kbPZIGOBYKUNG65Aw1UiQAWONe7t3dPDDjyhfDfWuv65gdT
0zsdVhP/SghfMvzCR3topU8Wt9t02r583SRP8unaOXUHOeqLuRjaVBDT454HduEZ
0we40oVC9Lww/fUAuVkyVjjDJydwmQ9S/zuhqxMsjXb5cVrxGkg9X3aZ7YVoY8sS
LgnASoQ0+hQsDK5/hOlmy883W8o2F3+8WBwJOKZlHbod8QKQBttBCNm0Y4+0yZvE
H3QJQwtiNYowaEzo8K9OGZ6y7ZNyBsl1srkwkJuuo0EbYL6ZsltnlpTuH9kbMuSJ
QoC4gCybzb/mCer5PaMu4Yl/YaOiL7YFzbuBwH3DKbn1eJrTR0HhPCL/T0i0Ne8l
7HiDS8HVKzS62Vcvt2BTdKMPUtwpvJZ37AMewj7Ak5zHHy7voELpG6kR1M5IoUfe
oUjtwOwU569qz7OHLnsMcAaSTofaD/1PzOnK5ZjOS9wK150J4qPYRdN7ACKXp8K5
oDqeK33uFzCNamxrO+WoQqpkDp9/qjgv/rP6K+fcZRhTf1zZAU4UAsaducdRLr+n
e30MQbIYFN0rsIdTkvIJN+YxFqvBA9QCUU/FXItLTIkeNg8r9qbVP9lqV9+QVd8Z
sOl4bHLw0CEWopMUM8ZjhwC831LzZBK0Q9QTL795NKY7wLOuAmAOgiczoLJKM3sh
TrSCWiOF6GjtmvDsw8BMmX9LqUWlwrob0LUjIHy3EynCSgM+7+k14HTPbthtQPuK
JB+6x4uOsyf2fUs1WeoxpGgDzOgmzAKj1qAtec+00xTmr71rkUN5rDoeY0Fd/h4T
E4NKll+NddYEzszdTAqN/NN86DPgobRIvVi4zxFmYzDoYvV/L5IRymMnJT6B25Ia
4az7jw/63ssPaWT/7t/tT5IM8D/oFGviBk40eUxLjNCJxDaQfCAA/LTtlu3wEBJ7
6OKENwqJumuTlqSWpgAmkoQp979Okk3vQv2OkQRifEnXMPB5JC7TVtzYGigATDIY
PA1KgsD3gIDBwCOBo2LDYmmiIBlUzMucdhI67x9frCofQTpcpXXBkWGeVfpe9qTK
2LsPLBAg+yQ6tS8o1B1/Mfi8+daKBFxg9G6WrlJkBJY9Zz9i/4obrSxQPj4U5WW2
aY+untQTVjj2iZtpVS/Eq9P5ec07FO/oU/sKce6L6/14LaCmxvDQOIXxbIuN7bH8
9A1dMe+R9jMmlWFbAQ3qxopU2+Gmj0KZ2vsC8a9Vb3jC6Sk6rWfb/7wjGJVzeA+J
EmACkEFqL3I/wbBCS6ACqu1/TiEV4MuyychgGVleGLnv6MgkpH3P/ivVlAA9OAFb
Q0bJqXZbWsUWP2YeH9WgCwZQ65atyIFZ/MbDF5Md0VOg4w+d8IOrQfd1jWCJHhLh
zzWbF1s65GrVjCFZCjAP5w0CZvAjwlPsRJnX7WVbYuoUY5wJZVVKvyWBU0iL8T7l
JkdsTcmjW6TeAcafVsOYlno8ryypT6uulTwe9XvyPb9rDBXtN3WlS0KzmlkAKWwr
tUkF13ilJsoBy/QDuLD66y2VIDHA84M2PzTkhDq6i61Stu33DGSlpwAUmOq0F+Wv
NTbHwspF8+n12qI8pT8795FasdiEo7s3tlILCZv7xM6br0BzJCVXc4QMGq5mtixn
ur3QCTurQnIPc5M12M0N4PtDai+EQHy+CfMbdM+0otBBJAbQHlSSPrVhPDU945UO
JVORzPrPq8moo46F4LW9goM63H8HaOIQKJAyrFJNBpN1/MpX9fa2Bre07Xi/89Iy
bFlOfGD7bQB9hDUytFqThpPlZRkb/sACXN8fkaL6mCkUrQ0bUUxmY+crfz+Y5jnM
8824LTcyaIhUYl2QuvZFB98r5TXFsGkUJ0dnO96CSS+bThNHhgp+u8yd4U1BDVBm
ZewYhzMlNV28g2cMET7ajXiym9TQ528gUa1CA72Gs9STZi31URNq7clxUi2vZoan
D83rDb31TbuW2097pwW9wQDSCeN2k0Psaw8Gz6BcXa8l975IE+5J7ULMVjaUBGea
sSc3d+7uKAzTGxqKJ3uEUQlkL58xc3+4Yh4iaC+vBoIpMbRMRjv1R55KuU6ISWzE
w0MjWau5s/3pLrFDZs9BPTn/+I+0ASrBY66809zwkUzzHDLT8ZfqTssRFm58Nrm2
rEbRdwxn68AWw6UuHjLAtboMOcZhTI+4B8Y+49YT+Qvw/cybDB3hKBQNVxQ6sb6r
JWiHirFGjXMpYPm8lTsMcObRuVDVHY6S3YUurE4/op5Uasm11niQ3QjQXe8QWC3r
zl8F6JUcBbHWH+oKi4K8zq4lnwFG2OqfZj/Lx2/EqBlKdH5DQc+ji6vlvBkzM5ZY
9BTdwirPC9egkK+rkBjkVyd20F2UOX1OO36ZcrYOkROBIm5s0i+4dh4vBpj+5+oS
+7k/YshSplM00lBETv4uzuIdoR6pVdCMfkv1ja5wiJmnVoe4xLUZ4DCKeR7OUamk
jbk6VsCuRVe1ZYO9vkU2m78DFi2phFkFQKG/Vv/QI9RgZQZEWxfVuVMMruVLHaL/
SnclqBER+KN9YKSqK1YdwfE6u7aN+ipAyvkxNf6XYuF6lq87PexATl66FU8bBlY+
K7XORgRmgO2XFziAeiuK18J/+v76hPrAX/eGY8d3QfSsKMAEElcjNwIrinNJmn40
f2Upg7k0HNn3Xxo+DgNjJXNkPc5ZT7LMkHW57GnDBwWBC5PeGzOqHuCYu4EPq5IR
KkjscOfZMdlnbfFPTjOfOmjskn+/q8+PIjhMxfUD4oEQ6CoeCG+Ue61h4YH2SRn4
B8L/WHdvzLfRjhBoDOsTQ8k9SJndqNs30HePwvO4ot9m9VIJOHUjxIeKyy80P/lD
kfmY9A/T1azukc254kf9VY2llRwBccdAfS85eSUAgSR4HyTbZwgi42IKsTBCHcz7
yneuKoFDHNPk4Ef2UynHnoZKmkkzGNcIxxAC1pFbjloLAvST5UzgiBvl537ZM8C4
yGnN2zjNnKZgxursSY1ByiaZ9CmFG/bDBT32hd+oksUXdRqQbR+y/jLROaBmuZbp
cZ2u82fMhLGaZM4nl/YdhT5rX49duGKop9HnWmYJDtoZ1wRymV1Z+hE0nrgJbbEK
/+9TDI7LaS01NF/MI7tH3WtEeOU4H8OKvxs9cOgqWv4A6DXZqRocvGCNkPaDgdIj
1hai2L/uCrw3xds8IelBVMgA6UA0KlGTpam5iZJcLFsvYm9xopj6a0UaQtCPyT+o
rqfyFuu+0wsqc+RhOevD+ZzWy400ObVY5QPyWvFQqhfIxmuLQclCXh/wP5b+MfcU
R1UIGrtgWtJNqj+HEdXJ1pJCNBenuRP/53WrM3+PF1RFmAMWY4XlF4/g3ykeoNoK
LcOnNprO6uQ9iPTTJiX6t0Iz008kz60i/+VNMTCBubzBhUEKxr2Q99ZljkoTBVsA
NoYeb2TjDL1TcxKsj8mw/YLZRf42J0Sm8StjYX4Wkkxm/e2nZ8QyX2OrY5R4OHmS
ALoVS63AjptmhALicEGZc+lXo/g553JczB4WmHG4ZZtjIVEPbp5H+qJ2A+9downh
i7C6DX3xQ2wKk2zF439CgHU9UtMOaQEqbQWMg7tn6A5E67/o3tDMVD3QR4natJXx
Y/rJZCT630p/cNDMcyd52Miz8aYwTE6f8Pd78GD8Yth6bxor6cMtvdA4JNNKqS+0
Li0DMUqMQTOcYO9fXef824vJt55z7NKB3fc89P1Xn6GUgaKKzVr+Q5FPUMITU2Lh
yD2w5WDHcbrbJarze/8GfX++lUoomW/imuA6s9noE9TqQF7R9nXP1R+qjBQrB1Tu
GCbSY5vVd7hVtGQNF3418Nk2KQ4V+zrio2VkF1mAV27gCtoGLe5qm2NhYXO3gOD2
jJS8V58giaU3ufB6pCcqRpN6+w/KeTVtEdPd9ITNSNj3wrfDUY8Ue68pinWt2/i4
5n406QdmzPqfGQocZnic8JVRah2Yn/ZbUXFyFbuIprDCGmQM3F0ELAS/BeA5ZiK+
4qa1stUzAFDwet9ze6mF1W/7LEYxLo5Aw3CTSnxGrOXYBl9AWkpyfAmtgFXx2eqo
gBSdzWeLFzXLPK3+armlvqK1+QQuR0oYR903476bcZVU2TNSlTDrrxL3G+V4Ve1e
8cC7sQqSzJjB0tMvhyGOgy+b9tyYkzWo1JKq2grujkMYMsreNZBJE9dOvMiNZsKV
qjQqRcWyp8ghbvkJhF9snx79zQ9vGGFW4widFJbRj3F1BrrRQSVpZ6PAolmqy5sy
EkpmsAQ3bXVHwCDPH9KlYpje0FZRm7Y94V1jm9vniR2WY27Ti+bc2Cj5S8z+nX/p
GkUCa7SdNd5SWhnHELpWWHOuGzbmEWnvKkINzBQmT5YaJvkkf1qpOmta8uZclIQ1
lImKOnM0f6NTRE2faNC0V/9aRPR3eybPwWjM88O75BaeMr5rLKnKo0YU/2RMUgXm
iw6OZNnWUn+fUvQGn1a1q61sfqS6P9i3pT/Aq17VVY3wCEfs0vn0hMSTX/ZVhFSg
XxiXxwkfdoair8iJ/lkb+fLcymDO/CSRqJEPXRIACNCeY63B6XN5p/KpD0MvJYhr
9YEM35/Nh6FCzV/5VBdwLMpkAgWOBybLLmxQHSinaG45Cao9uBmlcuK3yok2+RlB
IYzC/DB+YYiWgrP60jF5HNBmojTM0D/lihcO2hEol9oyEhxUpSbfSJ9qoQYnHreZ
SpRzkHmoUcl7Q+aaMgC/nHTvWfvzYNpuogtpOFImnXrH3mrPLsTWj9OZAxNOqyMJ
6GspThcoh6zAQ7ih4WgadeqaBTVMOuF6lKGRUcwODG9DyAxXgB//JbE9LVtK4B9z
L+qwb8fEPNP+ERFZmZuMSsYjAl+y1TI7TKJNhGnipuHn0MoYax50NjUt5gZruqFA
tjYG9qRP59krflEuYsH3LCub9+KdY+BBDxS1n69+Gg0wIZLgZ2+J6u+dNmcCmXfp
mCNBlsFA5Z5WTFw9pWVpO8PckzbnpFsqmt2jX3TqubYEHjAcGNjWGH/FarAvNpS0
UmqBrjvar3OTsTQ23W/4f0YPPT/jfVJVN+fAsL89TNXhXrwEQbKuWZH7uX0WnTJ3
aSo13RjJn6LAdLm1A1T5iw9FiMFvIt+BcbSugZ4B9MngUDahoUTp5NTy18JSPv42
RnCBu7mrCD/em+157SgUQA66mxZi+25VOUulx3QCcg1sMRHR2ISWNYcvogARAg4Y
8q3hQW8fuoofahDNRrN1SWyQze5Wtgv0BrRqEZBxzCAi9TEVRdzAjs3+M9i91dtU
wf+5qFblCt+zk//RTJrGMttofQGQzfi6CxMRxvoXQO9FFdE0hlt+rSfeH0XDj2zW
5RKj2zPxmYU6QqUJArfJE/zp9Dg/dWOkJKKgUI1A5Ytti89oOM7v63LHqGyU74N7
uRH5wlV+yzJtqc/P30TqedF0isedk6/DyH8JoDgUbGOqK2AsuwCVKc/niQDbGeOT
pkE3ZQtzR7ZDYojVuiWn7BQEBUN25e+YV09F1mVGGn9P6OgHNpIdlmgRfYaajNXe
znPO+rHxkqGgPKWStZg3XEuW0AZLBFjuEcnGwBdhqvr8+tZxwFsCht0dkhm3CyMC
Ho3DSMVTvl12vgo8iLgSG5WQaDWk8x+K2iGGW6NL7UOLML6AP2CrhSDLmiOaSML2
pj9MoOklBWU8xYPi3BOBrMuM26igu+zMGj3rTxKpDwV5tvhp2YLOh0TgkKe4TPN+
AL0LA8ZAVzTcXkQIqTsA+wWX/RQNitwXh8XONOUnWCCogAYQw2QtlRStfyadwHnI
HzC2Sn0gitA2s19avFDyG6zCpQVkTZUa1OSI1NPAWxtTMRbPOLfiBFN5/dQEArxV
/FVKITHd2ngGyIDaLVTcMvu8N2weukk9PMZFbm6XurxXtVTHWFA2x6Wto6GCmqci
NOiMYnJ2E8eD1VnOvFrTwebEUasBUQ3DfjyEhWxl4p74o/toiM99P/sQ86hCXy/i
pPh5SV11GI/MJFoXUPEY+FQaLVOf2gjGIOup3WeVNcwSWCTDAV42rp/TVjAFUh1X
/iWKS9O8zv/NmXBpjg4VmHg81JaO5tJSk4DvNkz5SA8x0pD5zbo5Ijac0G2Em+vJ
LQLf3jJLhcWzYG1sOHhCEstMWswpu4JBJPspDp3pHp1y3mpfrvODk9qYQz0xNyZk
rCOUvw1lP6bBS5WU/MIntLJ1payqZU7dZfLB0guv9PNY4VPCxfjs6HRSvK64D2bl
MvSpk8dYEoezetVfmbB+56Ck3W1oTrvhxGhYeHHVLzhmCxSlGGJcouBzEE5JvCfR
9chikJiBZXj+VIFvoRIGVOideDP0PckrUTCPmEyH3pBmLtNyUkGd0Fwp3PACJyRu
Xo3BkTAqT6vmHSRxXdowZ7qkFnfZs7EHNZtgqj+YZd15z2qyho/i00g0luQYr4XO
IfVyBg3zLI18pMvFOZL7gD+VA2CtM9a7EWnUg01KMqNGG4MogSXz2RQkg7kAQkqB
tgwKlzia5ZiKnuo4yfT3TYQPKXLt0Ai3NTZGXDNcvFohLG5GCRPjFdoE+czRlH6k
H3I+PjzKrT7nw4jHkH15I3k8nyLkH2Dk01Q0rFHgu4Avwn0o8ZpD4KIBRf86zJU6
W/+8uitjKVw/V6JNRFHie79j/JNJq752q1zkw3sxyZ8hTT+pcNxcLX3psSHt6f7c
oUbG7wd9YSiPQw4nUVsXL//dAtg5OpSJNk60SiDNGRlCc2nVOELA+focQEyMFszN
W0u3ibi6JmmHQNk5KU/g0H4F54hs+10fu3MoOnOyVZGfyrWsqEqObHi8mpBiQ49Z
WrelwR1AGnp282wD1aPOsbON+esivxybl8iH3TeXOsoxfFwbS9GYDVlwR+GybmTF
vMVEAsLxe021LIxO9VZK0BRKTEOcxrKc87bdemvxWNLUAu0JeaXq2MlEhj6346X/
icTkjQm/ZMFzJ01qP0l53my2hvnpsH2j+QuPWFZboqUxFGYvuFzcurFTsoxAFehV
YIIPG/LJ6+SuWrXM2cc7hPLGgqXN3OHooyswM2WXFek2aa0e+Iu/+4eIGZu3lfD9
nlWyt2oS+lTV5+60ZVydDQ1byblQqyAwSXtX0zHnUwePuM6legavXU613uJ9inmd
yp2R34JyyQTRRoDs7ohOqsTVehjg3+bRaHkVIVnClRVXvIUwhsoA/CVQWAOMH4eK
UakQjDd+d3BKyFg27UTDRvEfAacgQS3oRmFRyZPfUjeM+vlTr+7sFfFrP+1WGqq7
k/fkWGL7XdC+T2H0duvoDLQ1FF5Xf0reeGacGOqUwfHvWqzbcNv/HxgZhxZw4Qgs
t4d/xf17jajifUsu5F14+gLK/AFY3JWFgAnSlC5c/x6sSDkKzMqnwatY6yNVDab+
3GhM7oZrH3E/79iS9J+rxO+Q81pvebDZJWwyo/JkrIAxia3kqc09cK/oZ/HnuxM9
BiU6+rO94Bq4Tm2WTOwRBDlM84ehDMczsyNGO1y83ul3gwzSDnlcwQ2/26tYdMaO
pE9ClfVgRpHI3anA1bQwemY1oXd/TVuoKkwmwvb1d+VhYOzruxBWXmhQd8R4zfNN
jXYcWwnqSYRXNZ4AGdUQxzz+1yryKsn7dIiqI30eEAqy/SGBYDX5iZa13c2eRAdA
6VGEjrNBDQR6X8sJ9ovIfpjxzkZpLwUs4SwPypUgXhKAEEbua3LFJ/J4aCfdVEHN
8aJaP2AZJVGSLCUsCKAwLWTV/2s28vcM3dpn0ECAmeXY5f4/64/LfQt18lInr9Et
hGXzegU4bV0K3K8/4kIyYJkW3Z2cPFohMBh/49S4PxnINoKdpLk+88oEz5vXagPJ
wbe/AZn7epaJR7VGovYd0E8nE0ZmKJ1aZckccXG+VCkH0eNPtmKY+gpx33A55wW4
tmcBNKaCwnOczkg9oq7lvIuYnFnIgubEm+/VPFwYbHGEVj+kHfP9+V1zM7B0yTHd
79PejYnmx7Zesews0Swy9Dj8dTWMfgfxCvn+D/c247vrcLkEinAby2ym4ij1kT1p
5VZYzDteSAC/9wjDOZ/UEVyq47Anqi6Tchbehy3JA8U7GVgqeeq5N6l4tJ61CGjA
GGQgTqEh38fcvNfamDMkEl+I59lI4RTN9kq4n8AzrrE6ZNIHAaUILdogI4EpD24q
n0WZCmFg371O/c1lz1iI2Mm3DZNkef/Nu4O0WKIdIzMr70yCGuO0jXSBoN6SVUI5
G5wzzykUfeIFrL+PzpjHGMXlvtqSYGeqS4N1vy4n/OA4UyCdqsAW1YIvaEDBR/um
1WnhtQ5EVOxVwYGSSXqwlML2xGyHmRxbvt4HAZoVl/mE/X3x2gWkfKSt80ss0EWF
JNHpK2rw3h1gZHHwI8DqrXRPglnR4aQRMG8F9zNJLNqyaAGs8NWqOeJft2gU7uM7
NJ8Qet4jkN6HuvLPeocTQx5WwFPbtB0eDam1b9AoeduzvLgptL20B8rSNpp9QNn0
Id8eIkjmIyNbamtPWxW2+qshf8fIN89kOiP+CJTJIeesEM9zEUUbS0tOnN4uSrDV
gewTxO1UOo9loVGllcR6TeKt2o6U/23s52sEyAyonXG+bpq5+7wwHJBNLVFBusPv
OOt5eVaWQX0ZzzsXfo7rHfVB7hx6YJ9WQ8Oo2aCn5UVdjwNzDAOqRRKd3lg+fhvB
awthQfv2hqcKR5MnGHyZyY0tEeyYlM7B7gYPL6IjQ4/2J6CHXzf2VmSG/IaaECaN
XqCpKAhtfbPh1r5MO8o13Dd33vomQUxUIR+P/iIu1Z+/5qY6PQ7wNxYgnGvdOpQT
mqtuJTUOkTnRRHHAFqw48bXDZwy+tdErQ4eJkV/7DbXZcuflSjmT2C7v55AATvc2
NTs4Q1Jqy9MPBue7Nn+UnB6c8gGbw36Pe+Is/rglYP8gA9w18UcCCzO4Y5ZQy+/Z
4vs+3TCM7itBpETSVZzi6I5rm7nVM6dne/0u3u2VNa9NGEfyP52NgqAZHxtnwPqT
AOl0Du6msjm/YuUQOs3Etj1M5+L2bVxA3pBuezi7dtM6ud7pDTM9FDVlBo+csbuo
n/gITY9fx4hXUkYFriMg2+FLSCEZ+JbHDbTAfieHpHOx9AuG6N2q+iB2YrwQdaWP
J5OUWRzCEeISNri3ddosLbWmIUI0kwy9/3KEIsRhd0B+oUsd35aEyHlwo48tYans
d0flzzhz4Qgq3UsP22JX18fyQuPpkVNWm44jjEqj/7OQpvtfvhn7IbBfKHeH6HR9
9Xb1uz9OuKYPaPdJqsU9Insb5b424uEH8q21ocoHTWfRddXWyEuJ12uidsoN+HKw
meid58X1Iqk3k6kzDv7jLnd3WW/XzMXkLhsaAfUht2ggYP3JyMU/EwNetOGUfPPJ
ciIBBr8Llho5NCmRESa38sZHOXVygeY82WSlGm3OyFIdcJTetIaQJzAm5H6iYBij
lgT+0SKRg/E/pCea3iDbUs5bvY95e1qpbqsgy/UEpS4ZTKMYZT3DRziULpe70tvF
rBZBBNgN2uzi/whPMEyNiU8GOniGaFyClNzpWwyCSuIRsPbHk4rPWYn7pe9LE9nm
hQ3rKQLsaB8bl04b1gHSf9aP8eZVVp3ejAmU+hDckuogQtjW8iZAw5oio3Il6S8G
rPpcDvntcAJh2PokSXLhWDyR6Lo9iUUiaSSa5civh3I2LTl2CJglkDVn6t/7RxWz
Rw0xeuQ0FgbbLvGwsqgtQw6iHyQI5hDRHdlLgqgo7CF5U+SVqct+4Ykdyg2dXT6+
HeMQQl7mruz5iTdBy4BfPfPT4xyNvA46OKk0qpOxLa1XMuLWHcPYzxvlxxCvAWFl
lXx0W74n18DFvi5AXeRwhLVWdPasM++TtR400ccDW/a0GEfc40/tClg+/CXDvz0T
ELXPs65pi3BPx9Qno7KjTP4khi48IrU8QIy/snAvaQQ6Zi7Gz1N5o7Opis/b/OC2
XaKrA31EZAKm8c+ilGytM99AnIL92exJwoHkHYMRNIaiExuE9MPUG77KDVLIyMO/
HnrA2/4cA4NzZ8Q+5Et4QBGXhbzW0DZA9FHZ7JHBdnKrvOX7d8qN/fFq00e4cgQh
aK6DpGo895vkpPrY6vS5IeqNv1sFbeL006EBpi2d+wjm/iKJ8dANiqjvo1PUmNiV
CMy58I4FEKgN5YJMRMAxT7ZNabhFZojLBEq9AGtPMeqnq8DJHw5BEPyE6roTs7Pr
c+7IhSwITvvKdGHtx6eVX+G0xtcm1/qVpOkjDLhCZc4oTmcY393cUTqS4MwdhfLS
D0xvPv1i5jfnd7jrGlcAq3H3BXgULwTQBvCkf3QxycSADal6qIu4CVTAsHEZoM34
M872Eg7t9pJyNQf4dQ9s8pR4+88PrfupwVS9P06ndt8LopKhKGWSvag7stAytrTN
1H4PgBVZzMoNXEPIq5WY+XGmVAPvgKArpa1dCENZdyz7/RKvGKvf+V6etwXBTo8l
OR0jdMNpILyj6Ogkf89NpCNnxojP0Ev3Pd5lEszXM82Vp/4aAyaVQqHvj+NzWwMl
GCLGpicjcjoZEJCHalMoQ4s7ryOsfh5bXKauCibS1F6azjmAZf8YKF9OEBXn7gDP
55FuKo5Anx8gi2GuZ0s2JySAGKGt3C5m8r9RLsI7NqOFYoaENnVkwgeT6f3nepxM
/tEbu2gvJx6L6TDhWavjrADXsAoOfnz5yiaqX7BFnnCvoaZKv7rwP7JosZdmd5Jx
b0tHWJL0o9uq6f6EB5P/r6rqlO5Li27c3W/1muI46ZGAe2OeWi/XIsJlCos4RnBJ
hUhNUVQRwS6OZspULuSVFnqoVcUKuAE/lrBmT3iu4urI/kUsfN8ODUNmPhWEcDrV
syRi+RCiqUn6AYbsqgRpbgG7V7ylb5D+gBMQGZePzNJ1z+hkoUD8c2AH3XK8MF1M
hxO9XXAwaWEstOJBiI0Z+1MCI02/IzeVS2a11JLgNKKbc5DAZTKrjToT3qjNlnxV
Mrl50ZjEqUdT3otRuzJPkaBxvUQv2843K476aJouwLWCH1xCWU+UvWDd1IAfIWnK
+hcfHKEzw3eY2/0/cUVJPZbhRXJstrAbVcaPVTsc/e8RrnVER+6s98Xw7pLg+RIO
rpZzxfHi2K2WQxCheEysf8chtI3dShG4zHej6KlJIflXUivnhEgiNFIaFMD1+J7e
0V3uub4uSrNFivpNE4BugWzz99apDMdO0x35rOZJlYux1+E3RUO1wTiQMDKcAniw
yfb+DclxBL2flGX3g38noN0GBf4WSGZiJcCUWAnNhZgeWfC7KThuK08IE+HtvVHd
AhpBYhLshBBBN4bWnViRgue6F4EE7M5ADwz2C4VMgUvuEaDvfbhGTuR6BCczmtDY
oMFC1Cmnt27GINN9NpT5Z+OIEdvavDUEWdq3g91vGoCqgO5wLFBVC/isK26YOpCf
70fcNLBN0ZyXg/K3L1gSuCCAyr76ZFKwykMgH9Np8+vq+C9A+2UWriNXmQ/cim8T
Y7jHq/ivD2gJs8sXyh/8eFAtcFFEy6h0aFEMuiD5U1oyx/FXOw8yVUQ3twlr7t3R
2+lJ/2/uEOYfO5WE1YoXORtI0FmXIuQ1VhB2KtGq7U9q5oKAT6iGhhgCKMuC5X3s
zIK/vcTK7MgoG1n3qRy1TEgTRmmksLYl71LYjrWH9YoQqA3jzwG24spOL4XIn8q2
lhPOkmhJn8PsPSpRsfOOiGNXIlHRmO7eZ+IZ7elpY1pDKzS/wnHT4po+VjTDMHqA
eqOPBFeNc5fiphngVo20B2wHMBQr9aojgreszeqfBbKhYGzPMsS0WXHcnzorhB4p
SjOec2rRIrnT52pKcBX5W1WRnJWhVq+w5oqNQVoXmVQtwKhklVHyyUQA9xAIopXB
XyD6C9t4hiOcGYsIleqqYB71MSikKKfFMtOQU2fO5RI7mCQp0jwmqNeaSJ6K1DK4
PyTBJr8P4fFLRGOSc7H95dOZUCXmc+ynz8isuZe8TYSmpPLaNfM5l3e5aBjYSy75
Fj9ItXlTVDvrgHTKYlyUIZ5ru4qlHamdyYeIZ5CIaSVgThOTTW+VHcDDBzYF0SbS
MPCdsbsohiHiksM689L4SnNJ2qWIxoZ8mlXYt3CW5cE8L3MLA3C4QibU783CMEvL
i3f/na+smPnxmMfzaIDxGy+GRutL5vwtvmlZC+6MJWrNqzzZYFMZMThA8aXuip4+
X4d8bjHaJAO1UGuEUMbKzCov0EMmTux85Rx0Ji2pdRd9oqkufNjjZNAuAawrOx+0
ic6l3Yc0g67Ay4+Qu0yB2PoRHMLaQiO7MVwrbNTiBEYQj4S4BplkWIFzjVVQxXsN
i5VMAlCnCoEi1Yo/zxAZX3u0mah7IaaueALkb4ye6dOvUhg1rGDJu6iqD19ULCaR
JmuI8MBoKCEAk0IiIy0qo+gIC5TcazfaR/qGQv391CTITiaz066mYTk2dj8Wn1D9
u+/k51m4LkbHR4SzvvDwTIVx3kt8saxu4iMfKpap+U617lHik7jwYJz4JdwHR8eq
mH3+EPu5auPoaxrAjx380TxXePi3AlzEusHC5h5HCDMToaeLLNoSkEFYfd8pkuY9
M8KpBkH49+nniyKdEYKBHiCOf7GvfkgDN9Zua3XrjbGVYoj4AuvQA/ce6CXvDwnJ
USSByJ2ec3JT8uy/u9o0m9Grrqmvq87uRGgCP0BYcxMf7X0e1V8cJnKnUuDhdbPK
QvJoE0DOD2rh0eoZIuJw0ybTnU7fWo9a0M/lMiWC3lhAPebOB34JWKJOg9ZFDMwl
pO1Dx3StYGLVfK4hy89dY3wIju2VntcRVXRL4RCREFd8G2pK003F1WObTvB77TSn
irWc7ahUxjvqYSGejas0hJZU5CSanlpxRR71mQZI17jwiINC7KjG0MuzbWpMbbbL
is/EvVJU6PfPvqoan1iWyoVCHAphzCO4+P/QG2Vp3mGafQ7e5RrQ/mtEkDXsqliV
hXPRRk3/plI0SYsi853P3OS6mP+b2W9crBR5Ko0vrIsF6Dej4L1+X3O0oOo/bUiK
hJDdSOlerz7WFQUuvyar4PlvrXjF4oAh9VrbkIdH6frcXITh6/9TNT7mwzUpCrKX
EWg7YfRp0CF4k7oMU4rrb+Rh36kWzBgefTrJT5NZvu0XwDWg2UkNDXEh8KLCf3xF
deEIFWyHtpcYXzpVg6j80X+qxZSKOQ8mw2FbLymJkbXIXtlWPsL015yBYZonkt+b
B5HNXmuxU+jZxEl+2OUeXkAYKmRlzydh5L2OCbrDSK9JffFrIifYVC0/d6eyGGhr
hmdgRVNwrlNZ6PJr80OaqLRyJnQz3ysjGEAoq8f0k8OK536jFGdAUh9g/lcc2Qfd
lE48UM7r63mENTeVAXy+N4r4duh4KvsZ8DgVfCH2qgxHI27OkVjgBGXw8HkscunR
9RTS/UnYdpOpN6K0oh1MjI4lPofYjcCgC4J8w6qY/bid3UimhBnDmczbcc8MAf2E
h+1dpMPIhrBAD1cY1xHM5VeyEZ8d13Bs6yDNHrwubSHpm2JQzypsBPm0ClqttCd9
oQmxv5mY1RuqnBCuYx7KbgfuSpl0DeuVic7CVlT7a/Y8VsWA0K30vddA62Zg+9lD
Jf3hVyISr/2W00lNy7QJvM9fF9+dlTssM5T4Wx60kpIJwKpxU6KN1zrY4syKlfkh
7RpwSRzD3EoJKDhsK982WPB48v1fSR94jDBMPzlhLPdBFp4ZWcKCeGyh/WV8K4BF
iDeW4jSFyg/xa4H+TfuFNaxUrK028Cq+VYXE2xY7antjJefS3ODE29AvecMFeh4+
CldFBazqSMT9vjbmghn06upF2wSEiVcSdhVy22vett1Eo0Vpk9GK0WwwYvf30ii8
vXUSVtAwk6AodAaCZpGuCYpnMbFUeBcSnw7BfZVocgPq6J3ntwUEyj97nxkDGdgA
07/gkt8oQwFig0l/UdY3OTyKZ1t00OsgWlUWhP8YU4dua5ZIbtm2LOc2TGQmZZfX
FCFFYnX/smsqC/A/C6b0/u/WeATY7x1KOZd3GxEafhYje5s6qr38LmwJHLPhSBlD
V1kRHdKZqbVI7uYg4UldB7ZKDhHen/RKokLbfiW0Wtm3NciqoZg2cYMAnV7WLRnk
BcsU1oVKOi2Xsz92g97lWk40wSmXg0ncsJfaH88Yo5e0V2HGJ4yMlENwll3tsBES
5P7Cffig+PPzxqofAQRj94ACwuoLJOxcio8JUtxCUnVQXrejvuqnsCRZ8LWyB0t+
/xFm0ktgd5YI3WD5LUX3syiAf2YvEsdhsPDrJziYbaWY25QqsJAde8bMQChDf98x
bdoWLKC+5AjmACGcl/6wxB3qragyE+ckw8rqXrLIp2atzTx+XFU0QdcwRCaK3tgE
0NOVj6V1GmzJHRRV3voaHQbC3gWjXhKYOyZkehUEo2XaoZK5rpv18mBeOxgIKOOs
N9Rh2gu/R70N0om6F2ntAFFCwQb41vjF2SDpcQ4/bPjZOJSLzKQD/7fzdYwsowXJ
X9xjhXWpPEexOJuYQYwNAUTYJXYF0Z9rnrkCaOs8r3futB9BHxouFdGHeXmZfLt/
N9qLgVfNdqFo92rpuAhN2i3BC9WtStfURb/OzblWiPkb+NhT1X9VqviP3QmctgsS
gwg5C3ExkhQO9G9gUfI05LYK9AJZz6E+9tB8BB6/d9I8IyQtGfszD+9V9PppuVvk
84KAYW+2stnQ+aV1NcjF0LOFffzT4LGnasRQih8N8eY1pyS0/gAHT8L1THJE2Jjt
cQal6cAPTNTn86p9PZUjbMUQqcJyBA04SSfvDqMuxuR9ieqfnNiSA54nh36XKOL8
2hSIj5mRIis6SMg+5llj4yoCn9fGcD57QHORyVAGzDrryQd5KlEIfe3HFcZ3iN8l
1rHgdKiNVkoXOnkj/2YqkVOvOy4+paox481cHBKNQwjXr7Bigc53uMi6uG9A9Ffn
yGa/Q6b0ky2rgSDDwAIo8LuMuJwKrwlYA6epdKModQdqySLdoGt85yKVhOKwijEV
X81ISO1Xn12fLcKlfIkffpPrGqfsHkYBY3Pyux7ffrgSt4tyIA4G/Z8aYJiKsTwf
ic3znRUmQnjZmfucuZRH9doxLYfwXsq610/kF8tDIZ/XVF0XWmPH+WgGEFavM0BI
QclKsRBQ3KowaocJ/1Gacu/G74lxFS5luFbpBW2LyvFD0cQMAuxBZm9hCKaccW8X
eQiBHnJMIIEtwn/661upat9Sd+0oCsx2mKE/5ue7QkuK0arSDkmxXWVuxLFBVMj4
AbzIXwTmo/Dk3ZgRO2ZoDQkIaHO8FegkTy+R8dxZ4kdyKjB+o3pK+KKD/ZnFp6aD
ilg3OybkYqlbLH4t76ymNOe4XcBzGbv9OwB70RfFIDv+km99qxZHhKTTLWQfQM9S
fpnsqKf0VngNabjihNEIiGt2WWWrwOq8eKL9aSW5c2WrRHb7PXjLFnklp8GrnhL0
5+k5Ne81qifVMQx9j44g8f9th+w7VZbITghE/qC+thzD41HcAC6A2dp0Gb4y1lNP
GYg+Vs0x0/oKCbFSUyG1H6l7f5P5+8svWRTIahxWoEDJ1bta1m2XufJgWVOrrBKt
65smgksVK4gL8tAFK0MRWajW/8EgENPBvg0fIRsNbkK+Mi410M7rFEhqPkpT2fhZ
X4CVBRdcDZd7sXYD4SLziYH1z6goOk5EccTInjOKvgavbOb7Q5AM2c3UPSL2v+fj
Pb5sifdleY5xRKrCXvT6SnG9xEmQ07Yh29t/LPdh6ArEp9JIHbztbAzhp37d9eV+
V9pqV35Gr6PoaoVIXLCjsjYZ6Sus3sAnv9YOZy0BlOoiMHvsi4I/oUH9qDRt9THw
iCB9qsawM64rfL811ZvfjzbcKjNEx51VX4miYINI+alrVUfE7MHS4xUKm0HuGQAE
zJC5FqbCI55g3KCNfVIFvL9KlCn7a/BBaR7QGKIAE/N9DnZAwGGg6LGGRnTGcQjq
OxKu4KsPlgP6Yz7ppC9xRsiJGAWTvkmWwgYRpLKS+jmBVo7VRhfLlQR/uOmEIKq8
35syV6XSMYrc0mJZoUwnkKRZNzKqlun/xm1yYyiFrDDTHkWl28j1Ax2rFAP2mk5J
DEZ1U2Z2a2+dAaeyc7rTw4ijsBARHWjbnZTVoEqsTvFvKmjr8JAEqhIjVkdPnCVW
gqp6C5ccw6id8f4CGBHxXvQYNodWbQxw3+xSZOdnni677PSmFTfK4Tj+BWkyELg+
HbVM0x/HwbPX3TZiXje+ICZ4SXjzs0qkmZ9Rxk9duKFUPbJTsJGl9/ITozGYKMo5
UL+NblyV9s49z1lSgZUHlzH8Kb988xmz9jx+5MYn3BNKgRJRhfK7CuTVuwETKhhc
BiTQJAAmad5aV6D8uecOg7810ov4TT54GgSubbRBNv9eLCa21/dOQ0h+S7XhB+kB
4XZbngmB0tGD9oT413PYGV4PJ63ncnpbj8Z0v0YbetCJYw9845xByCGh16hbCBbP
vCNztsVzIiFCx3Ez7Fel2OXRUe/Ym0oe/yZJIFP8XiMdztHerseYV4d2r/MZQnEC
kQp1F8Uxf62uO7i1a6l0VQ0fGMcCnAazGfYe1Jb+mAobHrBAHvuGghkxXEYjsfka
af3hcLyDD+LPjSyoKjtJB4ymBVvFqCvGyFzfhZntWCBD6TxxPbJ5mYMKOZ/99UYW
v2QTYNkMZ1RB00MtxLfQYWy8ClwSKzYondCu7EXDMwU/HCXQziRY/AiFjpKhsFkN
ImrRTHetQnsK6cwi7ich+7OO88n7D5MhTDT30r/XMXhBF4pBTfONAjSPBSyCaF9Y
4yXPIIcrHr5Z9hO+CSXsIKPpEFWaV6YFsTuTTY/D8/OkiGMRzzdKHCQPGGpsBcY1
hMQPdNX58XjRmybVUEn8yN/0LafAXD8BrYfQN+LOFbCSBJS3LY9JtktkAtJ3POoL
qzDIBMGxg77PKqEkqiZ1xRtWC/TJo4Xj7soBmelQb7dDL/vkBC7QWvtkK13wXBCx
IsNdhOSXYUMItqJHnXPtzZbtbr+lszTWoIjuFgwa5IXjzgSxpkGNG54SseVSmlpK
Jjy9l5DaUxkO4OhRUV8jNSBfmSuXztZQYS5c+jNLkLrhNTFsAgvXeBD5lu5baZBe
T4Qy31ZPKd7aeA8kLYd9092SMjQna7pfhJHKIVjbPBqtmsBgT7nGHL5WYMGCcyJo
q90neOF5L/pBVzDwam9EZ98UJQ2C8Guak3VnUS1NqlkY5jJmnbIb1mfYZ7+X9x8Z
GI51mhvLlfx+l08a2LcIcyTB4JrgMcj5iainjAq4SKcGipZ1kDYcAazCZdXvJyrH
N084cu4zBTQzPR6hBLI2U1X0Q+sTs13X8Agp5e/JtfLY2EY1AABPN/EKCqtvW07L
gaEjjGGxbdG7EWef/WtQ6MdDvg7a3j1g0RWwFXZ9tAZi4K7HbXig/YTpgVbTi2cC
xxUafentpWGcOJE6hqMAX+jRuidH648rM4uhHB2ftRI6+hsmktyrQYvsfBDtYBK2
aEzDpCStdCXX1qCVAvThgKquv5FPOZQyRfwHXWCFRbPk1XUimiHIWLeU9Z4E6PP1
7IB+FMV3B4/nLyQZDoEltDchTMGfAkwkdrfWlmn27CveKBWFoW9uG70KuLb4CLIo
OHhMnAfCEkeoKlLmk7tKVLSlauiARL9qTz0fRMcA7TGJwCirsdMRhS6JmfnqCmVV
gFsLWmKpNgPV6yDDkqEd7ioD2vNN3eTsj8j9jewsGPWlNu94Nj4WyWxiKgW6fIVt
hrt4rFz+vAdFnWJ542gS8Dgsh4f+xa+YjRIWo6zZHkvcINGTVjLJNX3+n0xfKnpK
Wphh+a54UCHKY1hAniJR/v2Z3By1H54xn9Z+a4siahjCJo/15uJQhc17jc2FSO7i
cWK2mtwvRZ9zfgYcZWXDqxL7/WM7KCQSho5z/95RiFqJfbZ8niFyjVVH+XXRYHzS
Xet6AiXiG3Rcnseb2b6DvuEjnb4vyR9Gv3Nf8uyf09LUF22zi9a0V5rgCPExvCYe
2vw+djKQ55P1rw1V14U90+PAXzEUZ7NGzzU2CYwzDwr0Ij/2FkGbS0Apwu4ejh6+
dlART2ABVnO79jA+2pv09K/VeZCv4ORviKix2geiUC0vWCyNzFiFnFn0z933oKgU
/1SeHYii4QT9SNSj8NX67jMl4B3j33xtpNd3hj6ZYjF0wiOWUBbbwhiV4yusyfwz
o8ICwZOQz/UKzgO5bWsfFAT7Te3zhwC5S2bXb/oxR5M8dClOoxxEvt/KaTuZE4AJ
fhVeu32r8RR4+EaKZdASAjf06zkmfQuRVoqFyHWjCZzwsqAIcVcTG1I0ZS96bPIf
74TPexD7FMKgAc0sMP+lPmLLvu5MT32XE0vdM9MkEtfw9UoB7iozxLdDSgh1lqmj
Jmmz5ggNvd2ygW3ntdCBhX9P4Fg7mmLPAiCYfglT6tmRtzOcrYmIaTgp4QpgG/zm
9v3QeY3lXDucXFeBmBhKLhJG/nZTYLm9UalsktY71CNwwssCkQolsKAYcvUkPDIB
JL3QI1DoyW09Y7PFquP6ptjUvSt9KyfSlSl9Id1+Ys4E5DqXMYh+cdnWphkdJz04
E3ixlC3bKm++L6WhVk4p2DNifYrGZp666fygYQc9qMfAxsQSdpxU1sXiKfLBT2I9
tSe43iOzYBWAAWJh9MEN4FMDL26nvs++F03NWCCnmQ0jftX/TvSCaLf/U9pfkPfH
Os8M98xWnhmniXVSXmpCX2k1EqX+pQ+lRNqOz6yRbhW0UZrA6/fKVhuaXMTCQHgT
AmFUS6jUTRBOwytur2l5OmNzQrhT3GLFbotRj+rxmlfX3XGcplAbz5gVVqry6LQ9
zGWgODSYZzm1wfHKrbY54QMqgiFp/ujEbBNDbh0vnlZ35ogX4M+1RWUIV9Rf0AIT
66kB0rhbCcqv+9bjas1NyKO3CB9zoE0o1f1DNowu56oCNeYv1YrAF8OCb48sbG2U
m2ecXqZTRqof3MYlsp0hjzSpKVJBHz8gbzXcsjfUD5Kfin9beFmLXZNv/kkp9zfi
uO5XKOXehCRGZxIHYCGIJsa611KU69J48LeVc+xWDU+WWmX3hSfVvDzw/oFiz35p
gQmF1gOHrGDGzod0LDMhjNsmM0dr292ANyzOeoipuFyaZgrxG9JalvZZz6GKCTSu
ZROKp2jM83VgZgHSB6xrvUeUBn4ft9AX9cJTes0b69XYjcRNfBm8acs5IyPNqe1b
P9gE15kzYSIHJxtTCWn8dtgAim55JuILlS4+K3oUyhecXEnvjcCK/FmGknAWgvfz
t9/bCraNbZlFF831B9UDMv4Ph9IuCmD0t+T+O5/lnqwp4j1dpR9lT5AvkZCMQahW
fNbSMmBA/Pv+bJ0Nrp0uJhfppQpZQpM1zRCNtKEkGabInG2ohskXK1hvUORSCocg
rgxXNRF7Q75f2Vf7hX8xAyp/lhmtXZ4bM04tW0o0elO8r7WOJIiynULnfxxjFosq
cLWhR5XA25UHtbXaEjN5MHCs015xIVLemLDVshe7nw76apy7VY1G1EwXqXrQTGau
Cukw/2K3eeMMcwQfYkjH1KTB2DNafq8LPm2gP/EA0Twshse89T6U0F/QyjV03L+q
U6BZAdqsmUC5zYeFJxR2zGS5GhxpenkQvqCDSZXLal5BFJBRkFHP52duWpgdnrDn
jJLzmwFeLXa8k5JTugl8EALz6OD6tGV05i3wcnqvLcBJVWZvdIB2VfzNnyyhUlCJ
tTdOxqcep5POIske5WOB0ZlOQtDCEMX6fJWvsQSmuH7bPsz16Exwa0rFVxhcLs33
VcwnUlLQCqhn7qJKWTYCeXgkjVqq9tPamdrkBLqE9QA2VPWX1AjHxd308ciZwsiK
peNdFHWFvue5+0Z9YCwz0DoLAgD4BadAlF9OLjnAvG0FZviScp8FS7SZSaCtGyob
QIc1JvIyJwnZZpigb/4OtY7VvrFpZYuQPRpMX6bYBGxtRUGBX2LlapuBo09g0WSt
uhb9RP5DfK0/nMtkDoGjAUF0sGlgmbxA7vi40sSRAYb+oaHjO7GCveRpq6OlsLDP
clNVYRyZ4Bd1aGBTFb/wJcVOzeDrwbcYjhv7TkVW4XkPko8nFqhTJGM+c7V0Xd+c
vesNvW8rE++lAureQtS9FwB2YL43jI/9Ydvk0oP+zwZiqfUv+tRVsnm9apLALXKR
ihtlahhB0HK3JorPm9qbx5+YpnYNKd7P38LiZ0XluzSOEv6AXxHSed2vrVvKvfJN
GJ6qh1W0YnWIShONaauo6zbYn3Gony6Ivklw47+Qas9RdUOJSs+Qd8O9DXvM7yel
wDQFqfumVm5dLP7ChW3H4y6YZFybjVMA9tNFXei0EUwKswtNpS8y0TCS/jfmhrl2
ODKgmUBuyOIKl9OgIwcibm5OCcB6+L3KvW0cdIaDjDTywWtJzz71KtkVMrSBwxdm
83HQN/xA8JsHw0ZzvBJiT05A8qwhR6aKBe/zOqyjdgyF4WSo9qE0f4UgyF7rWZOw
5wxqID9Z8LByjiwmEOLsDttLW2vTw7+XyGkEB7Ax87XdOwheXfnEqg/6PjB6Hofu
RAjd/EJkm4DBooayrI0NWC8nWgJGt98L04EoEZLmcphl7iQ94mFi2+ntiV8VRKZ+
Q1ocGKsIXnkm7KKuikl5k0LEFKCZS1V9/3LgtWjpKdpHKkyX+xz9mBOKYt/9Ao88
mDSoIJRy8Qr6rIWI+AYmHAwcQW+1GG4gR5yQkBRJ1aiVYV4q/V5sGNJ7m2Ypls5o
x93OZoQz5R7OwUAxvWk77ssWkb5xTtZA2SB3OHCOiChm/N+2ZaxCU0JpFoKgUWUD
onDtNuWosBBODl8K9x5q0y4xzWBdoGgkW+wpSp3frgc3IaKv778lWch2yKEvbtsD
+CqeP1l8mjqDn3PP6EYqgrJZv4nrQTukAv2L9bX5HdUB0O6SKLlyW5bEkZCe6I+S
pyVMgnVkXYQQ82KWQ1luJrS+87jDGFfkQld0crHaXuufwWuJuleQajNU6MV6962r
d/vxjAQ8L68JSmMoksNrT2+KAaUtqLb1/Tiv8YnpMhqHwv0ViTWnw+ln5xHaWbAk
jiWkyx+GEQjcSpNf3vLFQ9zb8ZGz/7SNf25Izf/EsmgVYi9/+IElJf/uxxw7MPLZ
hPcjl8xJjwqr9eDRSb+GVxbIJ5Ny8ae8EEhpRxvMuPYtyBGWuQM3i8gH30eZPJc0
MKcBSjrB2fGY4rafyJxxTovAn7u8EjHhbfs7iysgdi5FjOz/DKNh8rTidzECB2AT
x7Xo5leBgvfrV1JV580pZi7bD0l08FxG92PWXVFFUvcvE5c1G8PNQ9HZ8HfupAB8
nREd3gHzCHwDbifMF0mHSTBf3Zy3IL2rZesEcvhqrUO3D7yEVYhkbpqWDRDpWtQy
IyRyuikZZeqpnb9InUmVJJjJ0b7zl6X8C8hpxtMg2zwwlpHLY2b5KQWRqdiwuBmI
Vn84OsZUFX4sJ+e074vS9DKjY+fZ5brEE0B5z6JocwnkKNNwN2j8TM6FcSD7rcF/
yczKP++IcsbushpvPmrdg8iazVNdtR3I3Ewrdmt7TMieOv6BND2hCJNc4aaE/jtz
la6cZIL0oom/ppZQBd1+rYc11+WcZysVPnxAgQ/L6QvuIDj9XyXEQw9DEPbbhrZd
p5/G7TX0zJO1G1jIuUo1i7N+HgrDymgkGxntZwjxeWzDTck7SDzQ9wwqYzMID3lH
l5nO2Wv9KS1GJEm2Q7EjIUw7KtRC/lHDV9BeTNbxOrPfPAw9NUT4tbboneqpgmCt
1xpwOotrs85Nj9smxDApONozzh8QKNbzmIJLdzkxDijMIPRZjrKFq3GMFijgyCzw
3GLYWT4vHoTez8IFoWUGLOqDjv3nUrcD2xx2vn6L1GQLSd3jRzrVZHBFjhfNZ+3C
SJhGaY40X5vXlwzexqD5fez9HAYfjtfvikY+DPEpiccxarICN0BMtQr98xQg6WPo
l+mYYooshTSJpMnRdreu7YLVgKbPcs3apKspt4JQbol9YnC7ObROO2d5l4uCu8jD
xK/ukaeBFVm6bIghEYtKo13gQ+2azfNCTKKIwlwXDCK2osOe0DIybEVn+pFDFBIt
+PrWAuqBdnWb2aDhpvDdFsFL8F82zU7xY8ZE1JklHGQHM5r/DFDfMkEBHraLttCN
0UvbV7kMF7lM2NEy40wJVRqEzqhBONuOozUWPt/n8pybAQY3GzCQL/jpVL8pdRFe
XqiCYEC7Dw6z4AsxfQ3kb7zOf5k+AhVz0Pv4WDkKMKx+aLi63/pHdnEPyvzUXt2g
FyjAPps8166DVsAtP5V15IMbB7lX3o2UZT1XAoHH5ltDsQDJ4XvriH77UQ23HAfc
WNOEvJFN+jeq0x6c1vOm88iFhEet4+jRha7dxr2uveb8lEgXiNoxDKVlNhHglr4f
ZYFCf36gE/zAFnJkjpmRTZi6K9NehOKX87sqZuXDInxGMSL9LVB1C0afLRpU6t0L
ibpFcec5SuX4bUQzrNvsy5HVM9F3FW8gE3j68hB98ngoZ3b5GrZbF04yVriMxdU0
EekZhz8RlkX05PrFFlNGOFC6Nk18XD3yN28daMOKLX2RxjgfJ0N9Bs1Jxtvv2Q8w
rtBP8gU4MM2/w7vFM5g+u07clcewIThuECfqipbg50j2AQNEJ6wFUcFEweAVvvfZ
HfAPbzsDlw4yCW/4cY5E7Zy7cxtTOfhXwXDycMsTLJNagrvIVL7POXfU1uqBSgit
nNiJ9rso28Qvj3LJwf9SSKaCmEgWZKz1NPtsK+hmkRHeo433wBZ33tvWF0SYeSWQ
Yy5WgnTGa3uoIMVZzWxn5/tgPyS5FNK+zjA1Ki+BYx75XIsObC0AaZ1TglH2ANj0
DZPcnxrpthOPpssMoVpY3/oFUWAW61x1ADSVDsob1y+vQ3JoS12kOPH5L3wQFv+L
gp4ycYajvlibtN370Q0J2b7nurh9e+GBjKl9qck24OEbtMqRjRPIQYoBUZ9CyKh9
w5Bu9jcYM8otSXnshNhLy1sD5XFsWHUAsMLdpFHsgFSug3HkCzfaXBVGhhB9UXV7
AcJmeBbe9/43ZIFUzKtl/8J9v7QTdtmszVActTqd+Z8ruS/bsC1Hvm0dpqp4hK4G
gCy43alrQBdJkqc14hAfYvPej4kxBvb7X2sv7j29fMA7yqspBHPOl11D6LQANj9B
MB8SvsFDlIW/8JTV5G1xw048Eh2Bw41iY4MBr9fGrmcEr1DOW9m5iIbchR7izGju
0YcLFdaw/lVOQ+4Pmnotg8NfUOIsgGBEXOIxdNKUPuQSQha3O3CCW5QTB4HcouxR
ZGzVVRYljJIOz6H6QmRRs68TQC9Sm8FgpFI2YASjJEYHNs6lfW/enIMq+bXMwEp+
JZNJYZDtuEf5150p7sWGTR/CZS9wZlKZo8b2QPyvwxPf8ocr16/gkpCzw+PiIQ4+
ObIsTglI41PWHzLWa/f92X5jZsC++f4e71vP6Wut83IbfSFLGMuWf3yCuLkyblIY
wBn77sCiMWw4x9Rng1tpL2G+wpzq1ZqKdD4CeywTG+HV7YN0uExl/mX0HWc94PMs
zZwpi3e96vOmGi2WOE//xwlA6rRz1HOIt1fih3qQRkofNyjFHvsP5NgxWmUG2V74
1do+778JIZ6F0fj62VHSu/kRbZ9eCko+t2wZOj+zAbccuX5p5ae11zWonqmH/R04
9PMIHpYD9GXccTkh147g9URptIjjlm7B4tqe+oDqHSHulrkyLR7KRxryHdHJx91h
r7Zp47giV46+PNSmAe4UcvaMVUEo4fJ5wYVjuf2KohfdMB4+sxQVTLIPVVwxnpIj
cGk36EjXvxcwASQhyMGehfTdK61pm6W027mVk4jj1X8h20dixRL8B8k0jwxt26qj
dclvt7bOPkpMLzGkXu6CKmxc7NMsvRsMojG+obKrW89+aoZdyBKKoWU7mANKanhS
TzV8T53u6VbSL2UcWDOuFar5tGQTg4jIpSfzTGxrDSpe/v3f7qR5IL74nG0ppuW9
seO/lf1jO5UxJKG24kMRusLV2/kjA+sI+4KTRkCTHGfU3/qbwhq+xvEGbXZRUmcr
6DgmFz9JZIZM2LqYACr5/DdtB9pa+CWcs1cO5nKZGjZzbXQx/m3mIdcPuwDkb0XM
1CGyjkKoKfhU8tPeBL19ODfDSg+h3by/ssZkblaPuFuGNzDTDgFRLfL1Dmbz0mvz
83+ZCvLTCppzhbUStx6bTzraGwlZX8t03DNvYYWDFxc55zFrOATzJBYabrp5ceV4
mHhlh/rDKsTbVwbyQ0H3Db/EaLxV3UJTtDCxQZzPIrBvxYxgo4YGkm3/PgQKaThg
nm7DhHQHLwZccfROa0oa1UiPDEay6Kzqvwat7EtZji+RyVdtUdzfrl7/Nc+8NonL
bN81h8DZqZMqqLXkye4B6FIV4i5kGqFrFOpUp5/fFxhEuSw9lTfyt+OtXuCBzBCj
dOkMP8pNPB3xX1V9+VE2uivfPizOt0WTZBtzowj/rxpwylRyrRDD/f9nj06lOoP3
nEBM36FNmMb5uUC4KESiVEw9WMqUhaXl3ERDcwgiiKxtZ4xphL7oF/z7JG2y1KYP
jqdzIdlf3yST/2/x0aI+fMVgKbclxOsvRBso3ejyssaYntfPawgwnb04EdkxuZv/
Pr4mfc4OAw6u84gGr45VZbUKQa+byATnj8aUuYKj5WBC2RIDuVPN15VKEKS/EtU/
dnYuDf6Tj80gI3SMC9XQKOE1d5DdqMeYSXDIlTbcBeKxwaGhXnOucdJR2wDAbHDJ
dZx+z+YH9lcq4/VOpUxgWHa/6g6L4Zav6qvIqiKB31C+sfx9mwR/DeCR9S/O50I+
28rZVwl4asrj8DJdpY592Xhe9uhqfIVk55/o8JrScXREY2WLDxQ/U42UENDuwMuG
EnB7F5nj6vXwoDptchaZgZX9FQlczh+Ip3RuBtytl5qDhSWwyFSxf3qKMI1lGr1E
CajenvquHynQZbzvfJPcXpEi3taE9nJ/XPvzooj8ljrE3x+SSlzyy5UtAb8Y1zCm
r6+2G4Dig1Qfs3J3MpTjGI5hKBOsXJtPOlbt4Wt2ftZXcFA4TaRaSNIgFn8vWn6+
3vuG33qKje/adCB3zs2bRhEUphc2B3CZXVKH3dO6/LcLonfYgUXUlq9+A7TIjduk
vMpvrDI0G1vOSwQr5X0Xjzjdx4dtzUdteOdu8TVH+dyOPOlxgL8tWTptzlCfgGtn
8XmprrWtfk7saCdLIPINzoxMgiMW9XeDohzR2hhlARAl2JKYetR5I4wp2+Iu9lyW
sGChKrsoAR6i1DoEtdsDKausOeBkhlPIunL35J2VwzmlcansQeNRCp4mpt7S/CYG
ICzEf6ldxv4qDu+1FMogRTrx+T41Dv0MYPHDZUaU2AeT0vVIMa+mK+JoiP+YEaZw
0cOprVR2ooZHAdxWKco9CW5cDd8chL+EUjlJdYPGlGj6D1KEGF/tVkyXf75wfHmU
FWJGBuBID5D/Ru29P2mfxY0qn7sqCn7hoDiy46uyT55hIT/OkbqJM+hAwMWnNO4K
pg8Z73gZcUApXVZwVSiqhWvxOyeFy/CY+o9FaLSfkYBwwF4LopuDSrqyb1R2f/Jm
+Yvmv7Y1mBdf3WeowSq54X+tC/Zx9WvplDoAQk2tQ6jsMFtokWgqrmQ+m/0jjVv0
oLMBOIG+zeOplRSAXunAx4ZC+B3kJM5IMdegRBu9IcX5P9qWFZZlrLdHpCQ6K14A
UGqnF7rneJAsgQ7YFHGAWyrbsqVVcqHqzXckR+cvPIPwWKnMHtWOzo5+XQQvcS1p
86tK5JcSg6+6J2Xdc7L+b2px0Y/V7FjAB98qYEDtsMein5jRba57DAUACZAFiDGy
mAHkg6OcTaZ4qWcXhKJfoXyG1ffsQyltIr0SFhC/FBTHKOo+eKV0iGhTvNRjr7wa
HtJ7aVRvrXRJCBFpgXb8gyhxfaXpqPqQvA1z3arqIWbpL5R5QO5vJj8wfLvrs8ve
OZGOqYeOqDSyj4GhYgCAIcstPQRgYbefgoXVM1KPgs5063+GrPApnXf3HfjpSL6o
cZxJO5USeYM6zCExEszf1x76KedmPiCp0mw2DnjRo8KUaz+osldnvJhpG9vV2zoF
FajUtVIzm/e+N2gMxjUB6Clo9TMCUArN3STUt32HwzeSsUSVMMUiHqxgkKyy2wwS
bBxitKYc8gNe6/LTCikh8beSTcDIFIuxHpPcpNOF/+MgFceKZMl/ORvMXEUEbk4E
MiGELfWSqZ781Qhg6IFnbJHC/aeYo+3HOpn/4QRO+QSSx47TrKt5EE+yYqxE1ZgZ
jmW4TQp9yLcdACwDc7UcgYm4oAjOHQjK5y8TMtx7cQnzYOK7tcYVR7ivYEPhVLcL
6N0piQglW6Y2HHRFW/j104OeV7tG9Ym2OgVHmp6+Y5ZrcI/bdyplabCLfBDT0O+F
6zdfuhMAcSJ+MeMvdRRJ50XPIieo8q2lmnTNCbO1emgU447a5NdL+722fYpFe8ZP
dYnN/+oF147e6xEuLoV8DRDnns/TvqnumH26S06jYWrYYA/6RYG91YCg/o9mvj/S
wYdIoUOYjfOLjgWQffPhDp5bwFnU+cr7vZoa/faxFbyn621UFuRqHjSeG2/mGPZd
rLItsCt8onZqD2SvWH8w0tOCvKdnDysjgmlxXBvoNhvUdmbacnzN67CLq95OJ+Jk
ytOrA/xP6lXb3zhp7Xek4g2hy8lPJYifl4nSr39o0FRySQcVQmsPu+CEUpd2gwDF
cvwb2O7FUURdoaEpgabFONkflzAa9MYC7OXF43tWivAZ6YxLQo09hin1MQtNZPSF
bgCXdXB9Tifv6FgcuhI+qR98IHgS7YNXk0WIXKQ3LKP8ZO5ytvfSW3axS4Z7OHn0
b27Ug8OoYkaFASvd+NBPDrvD5FY0r+WlsVBy6d62oZwZHX3S8f8CVQdt11orjPbC
Qf417DSbc/4Le4CM3t/40NISWlaKdIrWVd7xhHfFplai7m2DUlLxLEo1MYahOsw5
cE6iy6Dn1v5oC/He4oshevrtjQR6L1Hxg48WxNfruYhahdepH7/7rxTUQC9hXjwF
NmMcDNAYI5N3vQ5E4/7uGKK8QyxF39qJrrVYRVw34rbHSwKVYH3CAAl2SSALKf8q
peXTbDuuP8KonTL90OirPDHSgrF2fNfX2UvnUmRpd2vUTNdpDztXgqxV+P71moEm
zaKOp91smRaIh7R8G3Qqo5sKxc7qN5xRywMKJSs1fUTwEHDOsZVpWC8/Um6DFlz5
W/mt9debCN1xl/MfsM9eTy4kpr2e0RDy6BYZtHWx5jlXLnmAcFl5gU1/7X6eHKxk
RXWKTepz1btAvFcvO+R+5w7a5QC+437AIyrbok+lzJpr/ycgQOfgEFENkF3XiFE0
nx+4WGEuBVmnuA3RO3BmujukYrSzoGkAm9Y+ivGFMXDfOFhMPdTLH3ekzeQH9WNv
/X+YvC+M2yKbE7Va7dLZrU+FMbVYuofy4ADvzMvuvGETvs7DHvxX32w+QJzx16X2
CmdPRk3C8oIEwJ1SMf1gEg4+GiuLKAvkgx76U89Dko2yt36Ay6N217wTR5j5leif
R2U/IUQ5HA4O9Slm5XF99zqFx+NRaiMP4opZsSlzTDyCnjk6xctCEQ/RyV/qKwoM
e6yogbnQh38pRzpGPApmVncpxs2KZk1ro7jel8BpYmqqXDuDlr/mmLEr83EoHozX
WEUxUNKQi71unLJ88vdQUvlY69y0FQezLPXmxjgFTrb4zn51suKeFIah72OqGtys
wES4S0aiueFQvPi9YFWjhoVaObLWD5ZjnwcqBufv48JsUgIoQockKrsSOuJfB0L8
k+pBnSjq+9PlXas9Gv+d1isIeM4nmWLtuK38ngBgiNw1PWGKyv/fC3MPUeBI7eaf
5LCjJ+p8PN4AFn7nVs37bRm4vUfMUnUJ4PYEjNi6sjr/Z5n4KGzDGfacEHVCTmb9
mYWwQFwGaZ9sUOnoWYCGncIZ4EWBzL0bHd9EJ6aQv4hGk3YDYB0btzCwEfn1btUG
NTwIAk9c90sWYRZW+Ti5yPcHqp75ds8URZUza5eedvTji+5heLewEBwu/NhGFeyL
kfy1Et7RQOCOvl1w5p9+/BTXyJG5fJoj6RE3SS9msEHgU5wl8OmL2H6rxYHS4SNr
8Ot/P8+ncPzQO733NhQ2Ot7R14yXQjt7Z3rZ6zIqfQeZ4WI5i+CH8HZ2C/c8vhSw
b3OMqPHd6e1TCOnpGJ3d2DdAYI0cptcIku/coRHSojQa2040mVgE4G6RX3AI1GxM
qATInWeVCRrF8QtONebNkAFmRO6f3WpL3TwrrcIdQ3InsErS/YaNejy0uEUAVXIj
+LnCN6Qzwe+iThqMZUcAED0802UnHk+bj1GIiPxprQvUvODyMURsKb2UFe5OmBat
dfZ9sSfx00VmCnZucz2C6imH3YNX/axZVTZsDBTsctCOwrYCPrhTSQI3JdeDksZL
CIy7zxrb7MCo8ihM4JNbSiVDtooQLlD5KGobbuo+TiWihlBOvMDHpj/w7688y6Ro
T5h2ehQprFpQh6mcEzTLXNvafRQRTno7fNjKCYgKMK3yzKAUXoxHomsySEOzVUnP
+Fw11Oi2ElvXWdhYoHHg3t1XvvlF+ey2b4pwImMoGRfCl2m0SlzEXBhmbTku02s1
91xYlncCLq2OQPO3yV/WCXO0fTHDnVudlaRojwQdKKCAolRXXOlb+cHN2NzkwPw7
kA83+6dJgbWaioPsG8F381CR3kiKfhJWQmxXEMo6JNpow//DRg3rlvYWiOQx2R03
yJoy/BLDnEFB7+hVxM7kJanEgRy4l91NqxBakVanpVSK97zhW+cbDEcOMJkBe+bf
EAn9j50Wt1MrHWqFaKSR7pOHkbSX4kWtNNpZB4sW39DT+t+NvxNe6/94W8l34i+y
vB9t3EN8ZHU/ilpWFvtLRzApfIS8Vv1E750WgVyazd6t9O4QYEk1GD346r7bqHhT
7qOE4ZKF4W5FhhbnZ8fwGCM/NgZFq3n6Y6IJtzgucBqxq9g3ARPVsgfqHHgr8E7W
gakTjD3AVxT/ffqdgtERg91RcEg5I0hKepLiVqLwULG9RTiVa+/DQoMCDyItdO4z
zLBon2mqp1dbUb1nPxuyTgsnk3EHvVB9XlUM9pvaINSKqkzUCs6nheaRInkm/Bfc
6CkL5L0HcUM4TpVvfuNdJ1yfksxmVp2JOJrPj0ecaennJWEm1fupv78zt60zjMhG
ePOd7t9z25NE+1DbjkQyW+T0QFNJ+AnwdDA/7TaaSlCvH1IHGXLFpsBsrTlbNRQ+
QfNb3rF9Tgo0l73FpOdYG6fuEABJMd8ssa3e2Jnfkq1XYGV5zfZkUnznq1wxRtil
wfBSj55QJNzWp4qWOmj3+IkgfVlDtJj+NNDi5ts1JqejoI+IfXbixiTxWJblPhF8
nqa/CJb4bnzgDnuul6+JvaDjwFkL7cox85bDWAAnRklSBI5cTm+Prwhe87h9Ukhl
Dk8WwDVtTNvd/OjsmMyGjzK+bCB1tK8lgcU8Vk0bO50UeEEhcQVsSWvCk9Vm5Kjc
sePH528l6ilyx5Ps4Ng1axStQP4hZhPG37sDfSGPLqql3h29dO6aKZ+WHyfzT5UU
GIfyvgLBVAu3ew6AhW+OcLnM6inzomq7GiOjP1EWjV1I0ytVvhU87tfrNOiqvGHd
ZQ8EpxgUWIVlw1p1ESgMJ5rAuE6U2pF83i7YEPUs2VD9n4vyAxSsHJxs2NpC1ApH
dbzsIbNnvrP8N69A+jGGvV127qhwhuT2O5+v64N7JQZvLHcwTvpKhMgHo1aGozcC
hSjoulXZhEmuGsPQOxBEXBYO0qGHmEeEwssVS5VEonLHwMGfk4cXg0sMh73z/m6r
KypkwVhVIg1leEElTMIqPFJH3k1/AVDAz3iLSrsRkBHR72piy+YO6WUGuk2gCYp4
yTv1wL/9cicOuwvJk3D7xEVePBBUGN6ItBLBXxZA9lR01OoVCfq2rBLyhPRXzryt
2Fa4GFdAn6ALTodSQAhGmYibmhAfaog8QdIBDH4Bj6Xac1m7Ozg3q5ZX8sSFNqcR
1dOCFAjbxn0CS60mKywq3/pRCfP7He39Kjb/aSP/0hLT1Z5hX3oYQ/9USanmO+dQ
8nftUZqp8mY3mpK95wAk6NUcVO7zThrsfdM1aAPDkWrcQoeyynWX6vAEF9Zj1KfV
JBDGITHWNbIm7K5BRGceS2XaAFjCgNwbGCE+75mhI4RHMOYjpjzsOO4v1wNc/sUj
FA1xh0HqnKdT3HwFsDfpgVSZAhF8Mh77Cx8QH6PrjhE4a2jiJ9gOG/jrwnChRjVr
F832ZKn/xzfS8TLti7bf14odu7qibSp454WR2+BH36zoLp8EpRhHM1fluMLBHFQH
9CQGoFyWTtnVCnIKxE1I5bFnOmN2xEUpQKxDaTZjy27YoZv+2Q/bt9MIzk+5A53q
kHoXyAhWu4nj8vZIsUSL8IECM06qUefJl6yd+FpkTUfEJRn5kvZyUXDJFhswcKAR
KXpoEse5wJBgF/muz5OCO/Sm6CGnJg8ecc6957vO+dNcGrJDNppBkuYGJbkEI9cH
rqRJqQwVMTO9GEuQd4f15w8EpcLdxkCNE8oNXQhK/a6P4v52oZg1sIxnHFDQt5Wf
ZF01jYoXo1R4C7OqeCSxfvMmfpiTb762U9RHEHA6DbbJQhtTt3ZluKd0ec5a2j7b
DwQf+sK+ly1IQ8kUCbtUE174Ya7NdXGHeeNydR7kgqhHzC3LTG5G1YJpbOoNStDS
ABt2kAgjw7xJ4Pb51SO5eyrdsETu7q3PvD+qCdb8kHL6kchrZOPMzay3Zlx9Kts6
h55tevVl78U2mS8J75p3t5qUWhbWPH9fHYdt3hRxDwSVqGeCxo2TgLI7GMxlXX8+
fInrhc2TjBu+AMde5gHhgmC4sHSFGBAIQ8ALAC64incmbPe0n+tRf+2by3DD4U/Y
4WdhBA3acK1W3iWl8WcUQzVUWfvw41rmG4o81MsVLlzuFXOuUvoT1imuq8xWIEkm
ML+cfqau0Gs8qdWzPUcLRLUXN58Jr0ftRdXLEnZOUNOAEsp+qffuQCAUv128a0wt
cJl8txv4KrReqC9KholI9lNCvLEeCNff3VNYPnBg7wwgyujXXmUNr+g0GuGzm8FS
YTQwCx0XhUp+Gu6lMelSUqMIbpWHhmQlOB9y0ucZStFBfm50ORtzK9fIyt3FGrq2
7vy+BLSnPV3gYHm4U/pAIYzctkpkZ+6Swko/3pgbuxNSPRbG4fqIClexCfpQGBcG
RccvCQYEF6ionhZt5t8EiQ4cC0HNwBLqxqJgPzqG7WwaOQfJbuRLm5MkO5ppDYTk
Ygp6UCjkog7vMlB2V8pNUhCUkaLZWPCrEJ3xGR195GN93/7wKk9WuNyUMH4u0pIS
17VbUhSCu4enlQEkcLPFz8ZxQxvM5x4Pn/UHHYX3U9B63etzRYxCEJ0TVFtyhZOx
Eu6LCUdW6v6DJmbz6WYd+lwEfLlcFfWm3V0HuGNRoN6N5EXRBDojevdS3/Sxuk+k
CT7GeI71dPEg/gY6wig2rzfH6lC9QcY4BQY7ckoBswr48MymNUBMuV+AmofxDIQx
w6f6TugXvcMl6PFhN11xrRl+XqSGNrRju0QCyDDlpsm1jChvh3X5wAqSNuxJUfUt
XPDA3DcdkuxqW/bYIJ/Qc+qJ3n8R69JARkubg4Mn3vD5c0VuGo/ZeY0Ml+A3VNTa
Rh/pFob+kTIY1M3IbojDOvr9myWMPehZZvZHPRKlrG2RKX5v6XNE++COSqXlVWoR
oZzAV2061geMnx7YtIK/WTDo43krBTkJwXyd5oNkKt7WU9LMbSSJ9EaPUzwX/RoX
GymBsG6Z0huJps9gDqVs+p/3rA7crNg0ilOJZ19M3HigTRttNyk3OTQvTygrTSZI
LKcZBqPH0K0psT64R0fZ3+hlrqWW5b5W1SUUlQuZ3BWvza1v3kecS6vZnHIVntZB
VqVXpQVoy+oXb6K8TKAigCDwdOaXwTEhIh7PsTOlj5VIHsB+yvdZo19geG0p+YPY
/x36CLFeOgYz7vKis3yZxeS7Ezxaxwd2HekuD9Q8UiZiVbCmgI6mrQqg4/U3TZTF
lC644nPPl2wTWRqzYbsS7BKV5ZVBH+mFdmz5zNXpJCM4hJjYYD/LrQsOVC8cN/xX
3uuniKTvhqNS7OAV5gscFqil/gky7ZDdlqkSxIkO9lbbIiCTe34kpSgX07hLUe9D
Dzr9nC7QLBNlT/b9WAu/4J4zY/OY9I1iWg+shEhe7pfJon00JGo3CD+S0qXHl6A3
bg5+aqeiFv/ViQYVeXr1WvgWygxQkLqwDDKEhBn+WcZ/8Gp75w2MvTUhmv7KHDrB
+h5PBSBFw/5udO/K+BPYv/Z0bJIHc5GrTk3oQAnFacFr+RGIvjin0pFSf3c4RmRD
wA8HAkyFgJhmc3sEUw0lqXs/GzJndArbFoRWJhzdG26xtJFXXK2KpE9kzS2PkipR
nu6rIuM5tHkynalkEa5PEVIVdN541BdYcX3j29KHSMXMul7cckCaISlrI8Qcq56N
/gOKubIT0+93lNPZi68/O1kKnKexLcVBehWETkHXoCPgvVUNDy1VdT2G1xEYlLPu
BBxp+bq2mEtmmLxgjSAQDFIS1NQXfljtcz3Z90T+0rYyE5Cbb6JNMdMy8XJituap
CEC9eBYACSP0grXXDZb22hIMv+NiTg/Ve5io7BPINemMpQxhqOtBouhQgrZ+nPRD
Blt917xDYyxLWktDQghPXtJzwxfnxzwvAvBQ3hNxBzaXE+yEmNetftV04mG8DWaW
8zOVLkuJkTGAPOGVMZ+GuRSVZ1I3fQymufhKwfO9/BB9Y/BHbyETv0yuTJ7ZLk/Z
3uk3lXuGQDPbfxaIJr5y0DSpyZuc8O39jABT9O5sGsFVlWxdjfJqy35bnsValsao
2N00LuLKl1Ta25a1MwpM4QdQ73WW9js741P6J8jpeggfH/y9dsXOtAovBMKv1Z13
52MD3e0a0yVPYBvIpeDCvfB/fjVpgEbzrVgbOBZTxNqRwlrORecZ3YxrMfg53olQ
70XS7Jeq87lfMMdFM8ZGlcRnqZOL1jNS1SNFs48EkdP1EZgIRfNBFbGqtnDDXuJY
0xfKTRwvFVl8umt6clujnnGlLtNuiLvIbRvbiNcJ0ABCOqGrwqYwN2RqMt6v+mPq
sX1bw+EhdkyCiKlpFY3a4XIBAKqYqwUX1dxLpMXSB+raSB1oTMpqdHwsa6TnSaJx
zlQaA6XGNOsPCt5s5A2XfKSPeA3QWl5Lqrq1F9v8OEbeyG58KJZxWc8wufNitOMx
Pf7UAZe7RsmE2Lv+2MGm2hiUR+YhPRA0ybhbLzwBsneNgl/oVtLnWwBCawmcyfMZ
QXH4s6bnJxzZwPFgtbweChZpkHOBeGcP0Ti6dgeIaYMaMbXTYtgBOzj6ROYFjWzo
5oVpm9wtgYy5NlpjsvjrAfEsz6ruBfmRwBHN38cB8WHWd+Nb645mqosh9V5T4JiP
5VWglpVXqpbdfXFrWddfRoFX4emZ/ZJow3yIyV5+2rLr/w50OrjYghxDk3ud07ti
GnBpzaQkE04/TyoWRGnYLdGMlScCseFBZXsbr4bFJ6MdUVUVBODBZUFP1z5Son6N
PVqQHAi7XqNCXRBV8ud68lfsg5Vlfe6HQH1iVsNsmbJlRav3fl+XSyLWpYV/xVWO
AJGRDwt0iIEs7g9WCsBfov1Yg5bxW7bCYylqhpkNBZDtDbGJ+ak1DKNNqMNrltn9
ySdM6bPEDKPanfOvLqdRN0z4D0In3VhtTmlUDZ62+QyRtQM0z6S4fAQj6r7VEAzI
E2ZYPEiYR0F1D3S7DLI4eFGL1ObqAxj2JUqua9GNFV69+AgIrlf9X3oSCF1dQZbt
v8AURlQvkrsULkJMZhWYf9Pd1TzNo0g1eBX3kkeGnSKPvFbVVk1xE8TAyyvvc29i
wA2xKW/+vTVcPKbTe2VfMcXbhMW48pvaKEw6WDmJ5a7dxxe5LiHHevL8zGo8zvRn
1CzTuVK6VIiPazL/68UJMP0RyTNEKgu4MTeYxKIN/5/PT4nq7ZwLW2YoYl9MExDC
bZW4PeCdWYEFiRInrI+spYLOUmy/A09Onk5St/XK2jx2QYEIvjt0nbnHn4QQ/vZT
rK/LY5DaCtp3S7mPjFLpuEaBsrOb5SBhq8+5r+CbDNv8LUq9Vd+kY5fU7u4tPzaD
jQWPnreDpLv3hBKRraleRxB7ERYv4SIv7rd7egVnqdun47xhFlz93l8ZLdtLrliB
uhMbCcbiJNRJ8uPcF3YXww3lHzmDN6Cq96aWi4sdZepoceoD9bL7fCP/1TJw7ob+
CNDO+L1xtIv13AsZupdAN3zfEx85LRSYUTv10QZNTclD6BzWYQopQm4oKgVRwpIX
qW6YpQPpLBzaMOHekLOoQyhxarHGr5Rv8FpQOdYiz9OL13g5rvzJfmkOW9tYDPTo
cHFa8vyZLLPmJTThbD8vaowxPLt1/+8GEjKkSFPPrhhyDbPeN+J/eJ36uEafsdwi
E9LvY2/HP3fnhlYO4zG/3EP8PLIM4nldcUYBPQ2NSFi/vMhaMeQ13N70vVsHRAcz
wgP1fxhBLLMOvqVWj9o6LeqwTqsxOblwPlJXrilm0BUuwWCoQfuwrpzjH4F+9MNu
UOslbQjfh7K1xvZYoUKyWgV67vVGH/DCiHdukeiG0wURy3cOEp8eOjQvR/UGCqCw
thyfklRRuj6m99ewhwZUG606W2J6gQHs8YpIou5RmlKMgwVAMWSIW1ptGqvBOwGI
r91LUR7/Cai4luZ8WsM7ieQvqRtRYLKmhWxp0W1RvR3D9qbKBL9pR9I1mSTP4XNg
GW1tT3L3g9X6hoDQUeRhJGeec9AyJI+QzCVA2kxPs7n+FidEupOrTNgonXmefxGP
qXRioJ0cdVS+RSTUCABEtdWQgwKmI1ZGteMEpCW1JCKTmVIz57hmZQHjoFEsxHAV
yNHzho3XYPLQaxTcAznk3HLtEneBK7lh6acmqzaCk+U/MNyt5AN1OJWhXCE/eiyN
OHR5WJcxWP6NtPrgrgiPLrFxNq6Q6Aw3KnYNqLyHNeUXVVTaQNvkedO/qbE+jUTY
0SALfBx85/aiACSqvq2Pi8WY6QQgiKUDt7hBtD6Ig39KgeEvaBgD5ekFvUFtizHl
6uTelelNsEhNaHMR1w+bx2GLc0lUbRoqCJq2Pb87yOZkVl2Hd8W0Ng+7dalNyytY
e10N2mweGgIDbjKToWkrxLFVdHxg/3UhFJY4ydQeza9JD7ZXFzOIDymb6CKgSBfR
IaYXn/Tf/KvPiCR+7r48ecg2UgBCULODNbMMeEhaE9RrhzMowlBxrIOAq1NA7nmj
fFIcNSKiJsM+Pk0nV9IQy3UHNhet+pXXqopGWPqLSOGc3m1Gh3RuDPasSpmYR9Uf
LWn0rB7aOAthennlhPoSO9D7qHD76nJ9P8v0y07rnYZspcxwhLXFeBlPARlt/0MN
PYknR9yTfC1fTIssz2xhk0yDQ3kQwLBhbIcyABifkAP5bkmjCqskNVc0LUcIXTz1
cGVvWHKNAJV68pNqMas/eURobYlGQMH/BAtjkTKKrJeg+UG8by9uoVcXdxx5MGst
0dbUVnOiSqHWEd6mptu9AZagRMtssprZXef2dMTwpJ3QMCurUr+niqY9Qivdu88o
xujtz3YDogJWbpsZSuWHfJ1GIpKjE0Fod8mykH90g4PiXy0SHXJwDO0ZSiz6wBlD
acSuwysWXG6ZIUYDpdcwT4QryorfVn3IAorsjOmzU7+UM/gC9iz3AxRHF1HGAqJE
3/seHtuPUij3vGCn7Z1Q4otmd7lDgYS1fzCvO3e5Jv7LJ5ZCUUfAkK4+5r2gPVJZ
RVQgRFr3W1OnsZZpd7LVxss+kjLRwypsUV/yIoUIVO7FKwBD/xwGVeR92yHMge9l
o7b8xIOO5s+OWcwPdd6xJARHz2BTW4daagLzIBVFYp9T+DVca2ub8AMxoVi0NFnP
GsCR+I7EkRyP/+hkz2K7aBBkloIIp91wDAxwlKIH/T/R04RVSVJPkOpE2FURh4j3
vB0wWyIQWnlqeSwaFLVgk7g2WlrNpM4lV36WHFUllxjYI0jlxteNkUHIS3UJWVtF
mMCzgjjf0vcbnL7f9WCz0qp9aaAKd/JxUmahE10wJ9k2XvicrWpI05EOVMkfYItt
XXSYXrM4KDoc1Cg5IzSKfWd4Qxjb5HE+zHzcm4oBk2tKizNZTAyJ9w6rgHuZXWJq
TMgWSt4Tu8SP2dVVH0RWJ/xioxRmPCUUFMDcS/aT7/0GFgSxynh3sdeprlqapdcy
jlGTFLhWXCn4tsaTnGCfiXSQ/n2jBoax47QIo8jEvDoYjFJzytn30PUo0VPMqUFJ
rEI9BH8dDkH3ktnwUetf22gHXJnLPah7QONAlME6fJ7MIIVpHMWYLSvUZzUn5n2r
xhErOCBG3Q46DswdsvdNiGlwGHNExhL8iXkHezFNvkxd7yTrDYu1Wq2oSpsIootc
OJDm3sYCo3msE2lBfODPrZemH5+rLBd+KRPLgLDrHTtqTPXPjVea/gJZXb2N0oIE
2snpFrVB8kh5+ALCfBN1PXIzr0J+RtKnrhv/9vEhFQhjz7NhY5JJ8C8zf6PBmyO4
Y/yzGzXss8CwcttFeXzLZKbkdAegRTJWMQl7LRQq27V4U7sF4wWkBTKFf5ghvnht
CKUClm1Xwyj/j1M48rRuGIvfU4JzmbFa+GJglazP548YaVXpouzVqnI2WYyAkRJw
JZDX8l2qSY0hOXJ1N0791BbxNDI6BI2arc0duvod5Mq57bpzALuvzRBb8aGo5qIC
hao2cVc/mP1tG0Yqwhht19oit6tjffL9Tal1Rpq46HABquHnIajRW21Uv0t5ZGe+
ZE6Vpks+1s6cLj6NaRg7eHDJm4p6kIAyDo8MXQuCNb6xnEj5MO2cB7AU+xi+s7xO
NOumTffYscLCLAx7gNt1oSBAKoVt14H3dFM+bj/9Vf/3AR3q5DQImlQbiScuvG00
YCrK+fDoPTKq/Qf8rUHNcUkJD3pVYA1qLXz84kQyDJUNKge6vxhdpFGANUe7P5vF
Yj7cwhkKTmg7wQCSkVu/nsTSV0qyaKMGmy+FnvXUZwa395pCMU8vViXRd1ZxUrOV
huOlaowdroe9kfZOvpcujXr+kn3wq4egfudCaFL7jgksdCPT4KrJq9KLG6AvK4H1
mUpFXCtv5v6fpB1tQOHSppb9FDBohQ+ZWHkLObEttsEgjJUwG4ORsyV8KihmAhgR
5fHtMFTxE/w31xJWFXsb0JK7hAjpNmr2PXf83u22Sd1iYolUUTemaMuU9D992BwT
7rS5piGi0e+pgxiRv+/fefWzPAAVU1RI6zp4hcHjDNfLe+GNgRkhJtt5epjkvfnd
Khtger5obvAKrywlwBUElO61mEOAhggWLGLDzRLCQ4/NA0y+2t0qFy19Prq99Ckw
JbiYJkD0GCh57GsBF963QHUSYB14J0gPEEB2SH+clQClvPMEQyrkEKT/ewhBk00+
Yb+I9r+ASzu6V4h7dfVcJCfs93kG0U8/kxyrWBQ1jfgmc/aArP36prtOEQ5ia7N8
eSQ7UUuj1Rm43N9Ou7jZceplip8h1ec0TtmrymNdNlPMr49gbD26BSi0lV84Edhc
oC76nOypBcnQwiMJRqyr2vpSo5PhHwP/04UYZVouFRmJngaScPqUG16sqQuiJhHl
jB+uAaHjzp8UxhFbDzrWNEu/M/4/mbSGfroc/YTLVp1a2bkiMscb+aLb+ngcKoWp
ts+kxu4t4B0hiBpmRPjO3B7TRME7zvsCT3CT4r/5SkLoqauB1hipX5SZCc8Rf3fk
4LW32PFqSaUhgfEnCrSCkhiqPV9nwZC11r8Q6agHPJeD5qR2OrrDGHLNAtM/y41H
mKvpWGF5RQj3Z9Z6bYgHd1gGtJmz5criBq75zvYer+8QP/jUj1lFn9uPE70QGrXQ
GS79gsWCGqGQQibQvrVLtNmE8d8+sh9Pxl3Zmei0IEVKjiUpxlWHCSYD7AWOdPwg
4bjOU14RzDVoGVi214t60rQqX27jf+ISNWfC+FdeMLbsP9h9npkGYuIQuDCYcwgf
MKL9VlZit88JfURQrKhbXiIAK3alWf3n9fP7d+RYsVd3m6W//lXn5RxVyxyKVmZL
GuErYntHpohRgKxBMWWbbaNhNKbuJjzusJgdM60EWd0zIfumkoC0HS8eGLumJi6T
CvO92F7Bs9z2vqsyeIfHy/6CEvBZuyMbypR/vSkacBQTqDuYk4uPowrHHGx579pp
fmLiNtIHH5ovC3YLBPOTtP+pA4Nwv8lFBIRAxJQ+OaXNRWzunzsCNCnzPTKkUk5K
uiGO9OH7aLQF+3Qeow6FCiVtki+1mgCBa7OXZdQHXia/Ye3umiEiIlNhDeTaMmgi
PMwb7t6MQipojZimYDrnYxHZ6xh9MQqzahHcEWVHi4RqVFctbWsBwU02B/a4TrCU
ZtmuCtWKORBac3KEunlka4c6WlN3Vs1m/8J+ERG9clQupqAvzAhawEH9hr3TdtHN
biGHmx2BvPb9TViP113nBL4/gPwtVEYH2iHVbWIFq89X1BMuKnRPrWnGSz1PUzfq
i4FuytXGqvd/EW7+IvQAIFI7JX4NjOKCO1aGN6QF667BYPeq3f7ewHuSSmrthlla
Q8zuc8w1lSRlnTL73KMGTx+zenAPOTNiaPLZzjId6xtq8ojYL/+acKP2Oi2RRB+e
h7wksU0q04+MFFrCNvy/jMdP2dOfIXUUi8ihoWB5AeSc82M13RjrWp/7EElHf0/S
/VbbwNoJOuX0R0ZgZklMPd/YmEsClmcwUFCuFs4uRxDBDi5tQnHeTP6V2MKx4OvA
VRq6mS3Q0NHFYMe+KpoUesyxhrbAj5YeeHn4O6TvuXl4WEqfHknZsb75dhYQJJIJ
7OfYKNHnkEVAk0+v9wrO6wBH5S6I9YfwgxCy4ytTPXW/30ralefaBhxs9xZ+u4H2
idXTHkazHQLsmrvO/zzY6ZmpB3XyKG+6Mhplubdwx4jiNFbyhi9jXtyyRKNF6VtV
ljkJ0M0ReGw31s6tvGk0xd9KZJjtwvMXc5FgVdsRZLvErQmt10zwPC8746Jh2i0l
Gpu+63Zuhlt5yHKlOr/WyAiNbSTAaOJRpjxqY9sRGCK/dYz+fkOUwbIGUGUwot+G
9SB17sbJQPNrUWtsifEVevRxh/OqwIo+toAyqIMvhPYAwDdjpNceK4kZ/9YK4SFK
xfMm3H3JPDT75TZ4r+ahPTEmzM+IY0SsfbL5o8whpcDzTVRsKa+WddmJHvYVyJgO
r6diw6g1ieR/nqn9DOCrrV6IkVcxK2npggmZVTYVrzc7PFrTjSb2uH4QUvsM1bI9
R2XPMKD8fR6vNNicoFdDHwwo1/0wJKuglszbrEab+o3bqPHEWsVT18xxxvEkyJVn
QbhO6leNFTcqw3cKIlmkrGDKrj+HNYg1vjh8HP4kUS8dfikK9DraA9WlpFawOYrA
fpxMRFCt+nHQbyvI4Z49VEaARVhNODP4crY1wcVYWelKz57A5NoBmPS60GAk4HtC
C8ktfNV7HeXK99g3fBkbHYpcFryTzramux5QR1WgN/Cd+jJCAfDFgAh7cvasPq1U
Ntg2DzGbV6Z5zouFo9M71TvkpSWsi82G/w/GI4U8XM0t7lDz6WsQPBtTGMaFNwHQ
+5BoyY/6SEShNBy/SqFePziYuAiYFz+1hEdC/++PW+bT3YWNCRwNoldmdohaKwHd
XwJg89DeQk/4lnE2uJDpvw0ITiwJGWrn4OzDKd9NtPMUUm0mbHL+rT8lmy3M8Nk3
FXJNK7TuAIR94jGy5Oeef5bfdkx1xbkOvbK4fXzuFxujs1QuxRIKRwwwKifBtt58
k0n04pZqJltcSZ7zNbvzSm6Qf/sqZzyZNckA68kfKLVxRljT0KqlRMyBXkSMwEhh
AiTDFeFDpAkWC4tqy3ZFm2aUJ3pKqQm1z9GRMDjpQ0NQGdCuHiF6DrLg8h2CE3Qj
TbaF0SZSSRZ76f/sP+Cf45WFVGcWeJdnd72F8C+FEviCWn1sYMxkwaIm5mMlkexY
/S0H4T3vWuTg644McpAL012vkjmPcck0hZ8aQXIeXlr55eLRoqsBfzPaUzOV8XKE
QpG1ovfxDj9H4fiZ446oOGa7vfyFJ2ppIa/NPUhry48PHldYTGI9WI1+iPUxHLUb
lZIVCNA5/fFYO8GCayCI0KHuucuu24FRBXDQnqK3r507nNcsrsuAgtMsdRjqJhsz
MyZmwfYl9ooUmEQR5wiQiRGokHsV6JW5bwwCOvz/semYjm9O6psKDPLYQup8hcUx
FmmInFWfnGSdoqA98AE+A2TxXpvrxRqDJsv3CpXuVaX4BcK6kp/hyt9s5LiNAeHb
MRmpnhAV2sP6UhAH5lDtJShHo7dnMq+WHdv4vfH2pypSMWtSJJPmg98xeqTm1Q78
l2pgR+QQ33Ul4PeEDKe+EjIpM4XHYlkBOGhsIvZ9bXyCELjm7QLeHKsaM+muIeu6
Ws/Orw2v74Mu0qrTyh1s5+rLXwfiYDpLpU8unENmVoFjH6YjTWJ/fTprGcSbdR+Q
pTQUWanrb4iGQnz6ANekc1z8TXdkPcV8xYnYto6YH2gpSE0u0Dlay8Nz+A1OqmCk
q/kgtw203hxRtBc++QubQ2gUoCrE2NBic1oHwjjQ8x3LJAvb+Ro7IcNZbX0sg51C
/kIX+8aeZ5UMhe4u4xwkjGPqsAdIN/51DQSOT9uhzz5Va8IiZFrTDyOayzVt9+kU
uBODL+K13QhkM8UaYBii3EYFeEFW+KRwuZ1N7U963tNfFPcqt5LZ4lwiHzC9xWQA
wLIvxMPUmQvoSMatIyWUjE+vUp2VOqDh/sd6Ph3QUsBXDDRXBB0fidh+jxJTXEY5
F0ibJV/7h+nUuHbkgzvKMmwIZUDV3++CCjpixy/oj26bMtN5q6cCaSLczEztKoF/
RV1IIGi72EQO9qjGQtRk7ZNrPOTbyN4OfimO1RuAxe7FqUz6mOU2xPnc3qb7ruu7
7CN7Q18wpOdVT/24LrtUHjyg8Jf5I9F1Fk6NV6Mg3ybG5i59Vg827UUTYdCD7cDM
dyo723lqwsSf8md3fc0LKi+QMIA1mo/RD4gksQcltykfDCDRepjqZLoScI3zOv2F
PhP+hRYl14awmBzIB+Qj2O4T8LM/CTWNAJDHFKyOxPH699vIcssE2IpAVdWAQAlm
2cJ+Bd1geY4+muJffVqxtgxbBl+Ax/BnEGfdHdyztXCFKKn24LQ8NbYhu/a5G+1L
IRPrUbJgIWnSWpNiulNuR1eewCqLRCUGGVW2oiJ/VVIPDolTVWsaeS4qyc0DTId3
YuE3uHeJK0f1tes5V/6HYRqWUX2VdRXXjWZ+i4HEa98126bhCTyWJcZfFL9dyWAN
zLkyrPHnR5+/8eLeKnm5tcIncUrZyolFtBDITa8YQk9FgHcZJVGNOiJj+8Y42FnU
jDF/q3841JfeCHt0/kI7na57T6dSLOLYfo3LgzORrqtNCwPUeqe6DhtpqhY+pb5r
sHAK6cDRpfKq1Zn6WhRvZyuZx7mI5k3wgmNgzaKEamH+SECrMx1UMp6lUb1HqBaN
ZltZOR1UV6lbn884v5rGlyggfefuyIspCQk0a7hLa2Icdu7wQmZHC4TA1Ht6off+
BuAt8L92+9BV0LVBkb7Zg/okSkQTGxG9+ZVXs09B6vJX3hhsvTFAYPFjXldHtKxq
wo6CmuymBWNe13OWL/Ajpacs+Sb/joY52U7qMAuCaQK9kK50WWvsSoHTLOeje3rJ
jhEtuikjjyE6zwE3PjJCBxkN5pStnACMw2UN94d80za1usicVEvm6mAiQtwFb7dY
/zN9oHfXTHlabf8qpL92yNfLkGg303NZWvkk2blMwJ7z2yEtpSYuP/v+wrfGztVE
AnTWH16lp6SdpFaUeH0yETOoJtIhEJPDKukoT+08gM5alRixm6iBfR46tf3vWeC4
92svK4kiB+frof0zgkbdXqHk1sEX+MsmI0tWwkQ5PrUdjIq6BKJa3a+9AmzUWIRF
nWu+zMtsdLQvjHg307sOwbXU9luQ/U1eRJrudqG2IEn2Cr3TYASiE90pERQzR35V
P5UMBwIHjdI2PzCkTI5C/Rws7SH4iVaJj0Fog650zYZSPTnk5y3woIZASlW1eM63
9i3ixgcTJFKscFXPuaIx2v/Zse3RGRMRKGidxn0/GTWNJNSZU6oqaPC3dj3laD4Q
uKTId+6K/LGJeGm9a0l8uhcVO4RKJmQHldlvAHcIOEcepm6EWsbiL9xha5In6PNj
jAUK9B35aFa69TjXdl8AYX9FW7rw1YMMm/glGrSkxp1286np7x6A5sut+1YZdTu1
+vXYPtGF69L028+eDY7/2aeQpotFSx4fjfNhaa+pSEr/TWY78tFyBJOk1+tUofLf
Vv23h/AVSFT8SWUZ0vJcCj6OoWsnRHjZ0Y7lsTeBy213zvJlyHTi9BvhFOsoQuTJ
0mcF+B1ArNR8d7hOU3HVDz3JVJ53HNS+BuX5JCeI5QZJC2VwvpbRDqrlPAaiynv4
4gJtQCbQN9nDhNUVMCfFGTupgpN2+juN0BP8yMzSc7CyHo7RrcFlXyMNOg3RtHZC
uu7B6CtUotkooD0YCbcX8mXba8ettwDQKkjpZWIBPurbhSvoTx18KSzmAO8YzBW4
ArGSzMDREyUlTaxdZD2oE2QVjwL/Qbdr1he9CAIEeNP3/W/qxeOG+bim5f77bsK3
KTFrm4IqPhQXEQ6MfaD1Tcn5PU1uvH21LAFTpKKQOykRF+exI692ozLOQfsOdfTB
GgssnQm6F5JR2NR7xAadZ4Aa/3TyINUXvdUbFe6eJ3vg2tawXi0mHCEKgsuYW+Uu
OPY+I1N/ncGyUejjUSTdTT3MkvDyJBQXKAaqhywsQYOeABEtn9bP9LNSj7e75LFI
57WOO3TCRtR9xgel3rgCg/Yh54HQiCdbpue+yDO+z6pmOKJAdI678aVK7q1T9ivA
xiy9NHQQx2J4l3LdCpJTqLZET2sZ0EvJ3Gd0wJdTmdCJ29GWYk3bBxVmqNP6YqRH
uFED3/dQ/RTyZHl5N6AVlZhMMLhQAtMBOczlYAH/gPZcBqMD2ho5vxUC8y2Sux/d
Wdt3wla90sC9TSCJ2siDAJKqu6t2iKNtVFkCnzmwLj/WymOsY9CCE0icBptwWh9/
ZjTT1UV/vuYmqZPp0VyxacbbWygeernv35DHPMcZZpRlKZ4oO0OzAz+idjLXF7u6
SQyN3/4fMb23X4ba4zbXrV9YnEiAyyCB5W0+2C/64JAjjp84sqROhiVchsDhbJRe
Skad3phEWcvZ1NW09mOYcztfBjQAbuCZHDgRctTj643DcmQg6ixBIluujN1rrfyz
a3rzEXjqYjJnRGpZDQcU4UMkhbvDrSlfwjE0VUkQ4cdnsWAcdJkk+DCr5u9NMN82
UauIjMVdRdYn8BFTMbodPD0h2wIU6OZhqIxt6qiYeao/BWqSL0dDjT7kkiFu2gb4
YtxVsbW9yw37+VwqlqQxwGb0BKaLswS+ll1ks1myjADs4ksZ+JSRzITrhQ+v7H6C
MUgLFxJfsuw+YIpEotgzwKx2aOwSrOa2tPkc0118iFssld+HnTNMpV4Oq6rpuHiw
j1bw4qHffMHCiGT4zuqZ5BgVuvDIbRu34bCyQDkJZNSeT8v0fgFBrJCNjM6JaMEu
meu0GIqMZU1sDwJAg85HA8yS9holttTQKBNG93dmH8QEKGlfC2CJgmMvp54Gdf7G
aHIxM2CbuBgpsJHhZDkvJWIPavgAtQfqDRCW94GsSPGe0g58G8upCQpCfSdWO6OT
b79dKr3mWRN97xQzJ4xphuy2OJfUMcvtHgGE8V57LMiMA0cHOUbIM4TuSajByAZ6
6BFfEQDqbeADLfdzn1untE5yNUh2PhEa02wHA/mU23uT2ut5RbdSy0i5gCRbwrkV
PFKlZUiGO3MpjgBKCVEw87ll3KdoD17AxktWn4jlQLQ8rd3z0uwRZZv3S4eyUee8
NBd4r2CBLx138HIU9bgx9GQG9aeS3Ch0f1y6TEqK/V8zNZBZb5imcPEjJe7wjCPl
Y3Ov+FHhWoe7T4aTWISGgOkGOuJsUFzgHdYGZ07Hj0vpK4QHWwaRan7OlTTSpJii
FgAFUe1irmzngLS6pYhq1za65wD7Ak9NhjWyF6bi83MDz8rKjlY9qs0klfvNLANP
tI9exn9ENxIn3enj1mlqxZ5a+wAsPTG8jsnMbpwfeJ7t3zV+pViBzwJQi0G3/cSE
PQ47JfTIx89ol/qnvNNfgUkNQsh4bOiRpTkAjYt2o5SkzBSilR40QreGpS0O4DJA
TRg/Yg6f1/BSpBDzLi20lIeXVxpAv7nIy84E5wzmLZboqR8BQ6VLQw4qL9sb7qKx
2p2CYrWhhKN6FFOwzn/82nRQ3vlMkduqMqCZNfrohpbrxYIhHT1a8SG14pvSkLvC
RCi2nusrK22hdvC/8P5l61GhgDhPJnysl0p/p+ecNabAZA0jOQSNoHX+5dt20mH/
DH0CjZHSYSrtgrucsJzHp5GEsHm2m3WnIG65AfxV8LlCHO5O0lDYKC7FJCYbSPxX
x0TwKEp5G/htA2WUmCukv1k6/OQbfH93pdSmAJWrmqMIKe3yVlVCoWcXjwjfx0Je
3X3lplALMtZrKH+Q0LSBBLLfRuB7Fpia69IykDmgDmzdSF+OxIOh2cLNp+H98523
9rn37dDxwgepY+NUOoxZANcdbPZ7NlFH5ffSwe71UpYD1B3x5palVxyMp29p7B31
KpzsDjdsUhmZ8YyXsLA4eVEVl5BYfCpf0GmglTZuFLBCO2D2ipJAAzMTGaAiSbWD
yBAd9mRvLSHuLrLUI0IWjYIPJV9hOKKLXUAjJ8QVCjlSYb8AeCja7n2SelwwY+gn
LO7MW/khOvqGx8Tb/0VoHUIibFWkTxyxY9JSmfFIarArfpvlOlAc/D2uaCzbgSzj
On3rCR822A6ipRlQ1Gkq0HiA+/IsfeLnsNyQxhOvqdZ4SKxu2cfVbiVoytru4w9i
hO/fJHyB64Y6lEcW8L56ygSH9nSMx71ZZcjIiOMS4kkFU7KXNGv9CirM+MgmNtF5
hKw4F1Ugs8cS5bNRxTDbIZuegkbad6p2z6Vzs/oflL8KUF37FV0JxMVVmwycx7ll
sGW2/00kcjkmGjEwg09bQFZMQEMpn2N60tsqrdvzixYRt1cNSSGcqyr5ho7y2CDS
+65XH3bIFPLNqQlje1TViAqcNZ1mSyB6d7sdAOFelT1gw0l3zc2jsGTRTOpVH3SO
41nxXmUpyzI+E8N2KR8Oo3PDFeD7xDniV6hBbPtN/pvJktOsyqxC0LQnSNriWVly
EFx6yrgv+K/BmhjVVO1I6dpyeesRsh4B5EnFa6jUi1+4IJ7+xz5n00kL3tLx8SLi
KOXSr7iSUh/jDT7ZN7k9soePV5W0zCwI8RCQa3TinwzHH93qtiIt/IQl/hCJCLwC
Uc1ZadTqAY6GCx0LfzX3juyzcKrAC2nVOkPsfzawT8uNcMZBngffbRIZIcD39NK+
pSDeXaP8R8EuRi67IZUO23OQIGDWm57Ca2wJT2Xems72j5SnXqSAJyZN8RdfksyE
xZyFnC/OtzdwacJH31+4Acgim/g7d+ugIq6nILQTPvyorpOHksEeIlflbQsUjm74
ZqCpys5pNler0y3ClAN0BDoKecvYvp5CgBiSu4S69jFtTjHTB1AUsb8gcTuZMb62
f4ipjkcY7LEbsCvaShTAqM/R/nNanDeF1Te9x4PdgGxllRnY/y1ZYT1c9/R6fHjx
DIa6q2TYKlWtHaNFRgbwxdLeh532ZpkHjJzjqpdPjrtKfH/Zu54ok9keeTaG4hh1
PbPYSmCksMY/GoOeHOtYfA0SmPL9Olw11KjMlgCUDsg1xENunzSHBPV4Th/8Rk6n
D0JKaW5ZuWyD3fmGoFRv3FNkwCZfqv+al5izL9vX8GndAn5in3QK5DbJq9lwYD/P
XiMUHHcyMcrmTMq4U5LBiqbPUpTS1eKMaePxhaeVyU85Y4zxNLR00qFB0yioIos/
U+GDzKm/lVciZlnIFq9UC39FRjv+ukcPkYtScITA1Fm7s2vcB/h601ZINKqzahom
+JUZ8mvjitCTIXleSZlxF1+ue9ohSxN36gX7Dm5IHRrg/4hC+Ix19LMf3Y4Hpwxw
`protect END_PROTECTED
