`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRuaQ5PUl+N7HjpaxM7JrL4+B7WwVBnnIMSUsP04ErilqNuMuMwpB2HGbbGKabei
o3rAgWvKqTLV0uBx5raPqkqERDzzswX5mxN9f4J+66++f+JXatj/bKTe1lCUpRzi
IQX9R5fyYvcNDsb6djCIIwHqVKi5OL+eY2gSKxSBeVXsbGqdFYw0Ka1DSS52aK51
rlWef6RwdGMnzUcn6RlG6BH4GT+S170puoZAHU6uTvsgV0GpAk+PFVQrpYCOuBqA
rSwvBrPzayDGH0Dug1P5/uc/9b2KFPvTvYvw3/1PiYI1CCpETIPOtWRB9pQ5Es33
IY7uJ+bgry/FVq4abIckES8yT4kzeN3g8aBxuTFjmXb3rVmjsGdtz/rBQIG9x1Yc
PYjSk7U+yomdPlaHYh1GWr7iyrhprCN5sSx54YZSS+9urx5pgamamSqoHW277hzq
qBBBH2YhDM/DeKt38ObjUovjvLfHBruS/bjMm3hkJVBt4nlYFTA3RRjdbSIlvKi1
Saty7qRsBHDlsEfmwIiXDGxvfZe8cFDA4d9OvQ/DjhjLWZombioZRuJ6hjTMHTM6
XKPepBQ3Uyio0LIKCN3V+YldmbJd2+NBDcuIUUG/Ag+qt5pivdpa4ZnBlCpT0AxY
DNRB4UgeYTz8ydO4cqfoUT62aK65OHmuoDt9QmSV7WInGHel1vdBxj366Gurg3UP
LwfcIkY9B7+XwOmG+Tq7Z21d0m05m0WRzs99ayMUVFOmOSj3UFm51lRbQ9lOssrP
vYoKhbQejdhU4ah6yTDBQgBAkTnIvd3ueb1NsdebOvYyqk+s39j1Pbfwr6o7WYk7
xPpK9dfnYlqZQVxXlHPCFJfoL29nSxvTNM6Bc9Dvut4aBs+M64RrmoSjC1YsTvWP
JQIXSfPAa+VmRTVCL6yztqPHN4bgvyDWPJrWgdAuj3unu3UFScLD/YtKVogAA2Fe
vTWPySVXUUyZYhu+yL0G3Bpm/X7D9iHCWqWhn0dIEiN1RXg83VWQVflliqCnAS5P
7yb069ov9jWbAFL/qlH1E5q+hshU1x61u1vx0fbP/ZJ9kf7pT10Pt15X1+c80SER
K3pMbiXZXZGKnXaQut2xZwQvkVh+r7VlAZIv5FEEPhEg+hVko92HdJFSUBDV81nb
mQVgEA8bgcqfn6rMfyeNbbC3zbfO1FmdgnDUDJh8T4hwmsm0uBR3cWV3NF9izbef
4nPtDyY+hqNXHyHGqxt8Orlch6UOPOtGmbTf6IYXMWHxWux34Hf+iyr46+N0bp9U
JobbzLq3U0Wg91T0J9upS4twSJ9mIxghrVxNHRdGgZ9lSVX8riNRHb2AzLJ/szaw
cdct1VrCdZ/FuUgFlRlQZFWreScoQ//TOTjtHfDc5wOu2T15lMwcTkNt1gHiaMKH
8BiWDNYtK2f/nWz5mdTxsyrl0r3MzTrCmhcDaBLnB6pFXOLPvIo75CpV9WGKp+yw
VOSYwYoJL7xD5gkH9QL8UkwHeiB9hCECKJ+pcGIog5NKPSBDDZw+4hH4FSEE+ITU
K9MDU/qGGtO55MqyigvVJwdT2OdUqilctfwyrHVuDiiQ+EpeuFsNVyLcbvBWT7l1
ZfbpqLJBDYNJFLq37gtCdne5Djr2mEiQc/I5ACefGar7OxJGkJ0A5Up+X18wG2yj
2etKZYESo2y/LUWje1eLYECfcj089Tefr2JfOV8ttvUMdtgJx6kbFJeApCMQA/O3
zAwUA7oAooGLRGS4xqDlnBIoUV9aDU4Epo7kW7TSKYgwJKsRhpz9jnCm3XHK5JPo
IhcNRxzKUvg9GTUOXKW1OnmVMEMqMPrjmwXroQMvbl874mb/kuMYuo2bAjL8SMnt
8MxAOJjmHfrzBK6meViCAZYkyJKmLrrVl6p6nDjqb8zqWDygrZJsr1q6ob4Y2gsJ
4/ls2cBnYxQjIQ/esGsK+VQIxmHqKPK6S+kRKgd0We0/c5T64wikFaJ/sfp4yBrk
OQ9QPpWCD7r0RkiVTD1jt2dT6FRxZiNkgy2UYmcMvnCCi6uPOtgJtBXZ+PC0+kPW
0XNajvN4fwkPzef0HcD+X2oSnTBJ7pkp3Nh237+o0miMR9/V6Fe7WXI4fxlq8zkt
gL7XQ3EYx6YfzJdhSLQfxU+Xp1+9WgozeRswnBdVxx6of58sPHxytfE+CVniq5jA
XIJQ1TlMtra8/APs58+X//4HrcHcavhKu/7Y6HYbcP7v8ztUAw0x/1R+qkPRZ44j
RAnGtJNW6iN4PvVvD0StPO2yc4JrF20Y6dtzjqbyNzPMHIkuy3lEHQVR0KX+BKNg
N2L9U6GqdPCpAOHnRK43qAVk4C6CO48/NMVHrzH+ybes22ZWiNVniJdpAz+LIX1u
NyIS8HOIx2V/yOKKwU4QLykqzkDWQcilQ2olpMM26nQH0T3L158kqpBIBmiL8b/U
uFJLA/Xf+niIXL89P6o108xIZS0EdqW4orgf079kASM+DLTIVGCpCiV+Q32TVAuH
UNTj9oibciEBPmpX2AmIuWZH00w441g5FruL87I2W4ZcVWAggaWwJgPcGfzbRk/k
eA3CjYeIzEPMhH+iH8+Y81FL9At32p8SD0LeshTRJ+U7aH6b3VjFkX0BDFLMV3qn
hrSo1RUtCYUycP0gEFVIMFK9XXwHwAM8LPJysRxMhuuD4O3/P0y3eSmZVPR/pdhf
GDyv4MrfKkHthhMTAsv/0hWXOnH06X8wbjFq8k+er6rwi7p3j5HfUKVEVGcVAFcw
h7L5AWVv2JoZMDx3urt7apsRnYqpioEUK24SMT7XyA0+SvzB+ysyAuiG9ooBFyH3
dYPRz0oxI7rDAjenAsQ+DpsJGpjtozahWaCHJipJhPn6dYlXVu6rJlm/ekAY3Ysf
ysRb0jn9KEvDFJnDDFDfvu039y4uQK0OS+ee5uoRBNRIMzI1L828olLSfp+iU8yL
P38tHHSJa0P1l8eqjTQRfUDV5O+b9a2bPCP0drbBn534ERUoXUNWVrF1rF0foYMD
d0AV5Cpa6L1hIxHl0w9iY1TjwJAcMGWYaUPljdh6cGyvpMYYlZYxgDvko0n/95mg
7OrG1YLFrvdK1r/HHcibYfjAGqJFagZvx2xJTuDzX7r39Lawz/yVQzExn020qAa7
14rNGZ0CnYEiazx2fSZaljm+IiNcsek+vSiKESGBj9AvoJU75ZkweyP9sO+GfvY0
VW44aQP9g/iFGD719CvOGxlNznIcdCQ1nbNMq+AunENjCH4jlety+IR6qAHZFF0s
lpIyMwZh7N42NS5U5q/XVIYUv8vQlcffeWJ3+dpS7OR7pVppVFKkwDGXEHRsEWes
8JXzd+IxLtZmEMkCXrynNjxTm0B4sj1YBdbhp8VBrzoe2Npgjjgw9epN7vcOdPip
6JZNJvbI43KlFx4TMd09gaxJwvI1IZABCYRGlNrwUhFAKuWFaTqtUKqBb+PKIret
N9OVqGz7GTo+asxrTFmykFxOyIoFNjBGyjtV944aylp1n+lfaegiWEKvB1UkRnZA
c+K4e8lesR2d0D2LcZvmKdyqu+f6BpPqLGF3LQP5cwTaX5UhoOUGzDYP71+50hiC
7QfFrcOIJNcML1Cfhqzgq5qd54EiEGbylR+NzDMgk7sW0z1fxf94pPCxZcd/0Bcs
trTMDuE7FbhUVq4Rj//AjraZJgRMF3yzkuuYRIbYnE7loYceQYWGqAP3VXVwjxtx
WaDwxDqYou2ZuA0i9v1iFpSHjfMV8AOJfelno4AyL9ElVT2/2dIAgg87wfe0NvfM
1J5FAJ8TuU+MXXiUTN+eMe9X4BxfedcQ6ZwsG1xXCKBeu08YA5s+Yyk/6p5Zky6q
6SDgfinHAOp2K5bWt2M4eSohxL7t8bN0BKk6hU3m83tHZKLe5izJmuxm42Nxe5hW
niZ9DgJHBHt5M075xGfsR7eDq4ALgPltI9Q378ZxL0bF8gnkNTz3fzwmk926ikC2
tULk8QmA3CeaK2M8p9l5bf+UkBR+3v7xq/4Z2xkFyHJSa5/Ip1tSLn3g+bi5b25Z
bmu+0mzZMNAxwI23lhKkJz+KEvY43QEImGuMycNF9Avlx7L2ojD0ow/qUNgyqqdn
doAIZx9oCZQtwqTm7QQY+bncobFGq+mWNYC3T6GZ40if0IQEuhXiGE5TJSNfPlsP
m0aUL5J5TGpWYViAtYT5HXoIQtZ2I14ZrpgHv2Oq8gxiuQGYvwYwQRHtLDYN+E0U
wbMSwu4Lb7FmxExZPHZ88osZWv8PTV6zSV26B7txhFlkvoyZWL8iDD6zoteG8oe/
kKYQfj9rA/FzxGhej/7v086FxKRHIpcRyuqtxk71LF31dJ3+9xTrLEI+NRUfnuCs
OxKjnkAXZc6bJuLMnvrPmUHV/cPWrIxN6fH591Aw9cUWBTExJTIQMkHm+WqervJi
v3fVHAXMMKaElpD9EMYGXJvwdH55qZldQq9IqOsb6A1ZuHPI2+NTc6xcYUBpy1I6
u9xfPRr/OCxsx+UB4F1TXJWENDsH/TJZecCcGkvurLEDlA/RnsQb09VZ7PM6KrCi
1pP0HBBxyOSG58p6Nvlu4ldjZ09F/YWBWNc2Og+9uLTqfKhCFr8m8nqSJKrzko7E
6wZIa3rVYZyo8NLaGnUU5Q==
`protect END_PROTECTED
