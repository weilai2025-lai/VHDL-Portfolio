`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8zbDGkPGGVJRE1ZGnGkyx2Odyu4uOg0EzAWuZ5PIpTMNdq6uyVBPVHeoom72sg3
FDwAfCQBi+lTt8AJfqG0kWpfdN1CZ9S6vbwCsybIsh3VcddfBsAIFyIOKbjoulON
75xn4R63Afyy8Uh/Mhm4G/inVa8PCt8mjPGFZ7/aMuQqzknIygack9HSiVuy68jq
LCkVyeTjod5kQbRkW2IrrECnb3dpP/tef1epY/IihmWYqF9Jy/Vf3B4qFWhIdkMx
DJUl3RwTD2BAYNaOoK4LzuK/pFcx1eFgtRU6LniF8W6wyao2cZ5nLesRcglOfz4/
jk5/W9vcEt1ltV6TQC+zN7W3f3O+CeOlr4HX+NOSuMlW0u6JUwQz2CgcW7aHCjIr
vqB/stPIYBYI/MDgLgpBqEDo2V3ua2Gn8SQUmQTKxJ91IqL3bzLiK/2PVClQA+YG
9JgfIQBuyMqO2nFfavflBGh/pFQlHbuWiDMMizzLvz/wCOK6BG9qcQwsfmISUhko
OwE8f8jGDnoL7F4fv/JzRrFzO1csiedRrBDdLKJxozXsB8bEIUl4+8dSxd4BAKha
h/KwUG9qSRnbjqjzGe9lu0yjRyIl6dxq9FvMCNhe8hRp6LlfBkXTxSzEbC5O/gZK
H3fT9XRRDy3EQutSrz9RdukgZWabGEf8ivbpRoptfGJX0s0OITWzT1a2XNnZPFDZ
qUbPhMASH8GjmVn7swmKtig4whjWg6OyV3+/cQBbEaWYVttseqzALqKIi6QPrvNb
aZqC/a+ZADBMT7XbI3WrxxnaGLd9dzXrtwsyYw4g3G4Sw7ABegO3hnxZSC0xggqI
0pBsgQZ3XpA+BxF1r6mXIQSUlb0Vt13e8FNVmHU4e8n+vMfuZ+SAG2oxkA/GAIl0
arpE0mHPPh1mqSWxAidbHGsecnlH2TkculAGA+TLW1bM7Uxf9zCQcy4sezwpzyDD
wtWNps8sLzHQn4HqOih+aS9I2Q6TnX72ludeey6SlVnBtOzXnzkKdefFvspscAqs
avwiDt2PyqjYgGwiV681GVVU+lU1G1SA6JsXYIVftjiFOCeuh+arUdPulqcwEWYt
ynVhuUrSqz9vA+mJOaVSRdvKJOP2wbRHvQmRCrRm5YpifZhydE2wqGDpJ8Nvyibp
HgdHh0l81uFLtroMfswNgmCTcS1lwG9Q/H4tjAFsbOtPoLj46jaIKIP9+JAoF4z6
A48r1/6ZR1YyOcO0urGN5KNc78EcVi3Iteeeyhmk3Kaa7cr/eUF7CKM3nPyAInkY
SDFRgnC21uGCPxDm/jzIu+cjm4vYLGfhFaJYpROV8xC7i0peqtGFcp+qJWsC89SA
ya7lkIOMOkrCIg79HtLn++IwYeJcgLoZYxKlnsecMKKhcx7EPrYO6RJfPRm4YK1a
MAYomW8NT1JqX6AU/jRN7Vjp49/YrPSAT8BCHgh3sLI0WQh0sRrFXO8FvUoaAYOA
F3Z/33rIyQYq2rC13jpqAIzUn2EXGbyoArjNcXJrv8vX6NuG05RuOdcQ8XOVwpFu
GrJTEgt6wy3qNTW8KZYgSnG/79aFjbJi5KtZzqd4EQpLg3s4h9bz2dThHlqVyiTA
dhYLXy7fxR68puAyCtfHHecbj+DBYSCZdnyxRs5wCgHetPdtBhttQ3NxoKV3D4Ol
mDEkLK3ai0tGnd9PP8qgqitgrSUZJ/+MzHSiKDd5pQpxCxXh5ZeQ0u01wLixdymn
quOGm/losDBngg3mWYMVMcuxppqpVlaNwqYeWHkUMOW75LAlxaflIBzwCt0e7So2
auZxCSAMN4i4F0QmpGIcOfjJ4xC2g9LkIaSm6Kkuuu9vACuHjruL7/98f4pA9xxh
wxSwpWSMijz7hcibRh8tMILEsH40G4zJmGi91QiGfFCuVYtZDyWjzTP7dBhRv2Jc
0nVDI1+9aIkUoio1oOhN4civxqpswuD0AJV1xSQVsON28eNNbsIvjnu6M5+7qzRv
uYbMkCwdUGnGGzzdNoPOhN9AbVmb0PwkTsEVNrEdde69cQh1TziEZkMwbEYG0uFP
79gKfL2SHwMfHV+IC9qL75oCv3UCMeF+P+klLiHS85wxAW6LYkxzr2DzoznEE5N2
dP3WYgD/qtAxIkaO2RXOsszq3/4yQsdmg7Rpyt/L95v6K+wGQsEbzbdcvkBUSGv3
6hj5iFolHE5qAa9HRe0bdcH3Ej2wqyweQSYa8Jh43JFfjLBuewt3Vdj6nXoy1k3+
7tSMEM9VAj6TgLTB6Uh2WAV2aFj0i/anOypChSs49Tos8Srsvf26rWc6z189fXj5
NpChSXvrLupPH3fD/kcOtAaytGXL8IB8z/D43ZFlZ3QE2m7nbPsf3dvi4QoEt5yB
wBZENKX1+wuBLG8rF5BJh3Msauf1v3/yHhjm3jZho89ux8KlmzPrcjLRghQhsHIe
58XmpGce97OeuoLL1rK60gLdeisJ/eEihY1MGW+LkMLe1/yqXG34q7m0kzM9O+PG
vH/Mq+hR4wo1imMFEQMQl00b+2IHGJGowAcuoiYICJKdIQn/lL195VZFKrUgjTmV
CSFxPPFa+jfi4PRiF3M3fpRy6R4l0mY9v19Raaqwn06UMJ4yuSf7OO6I+t3AmcNE
ifiwZ0JxYCUKi7ZTQGMqNpCCkkydYHlf0xyR29BTfd3IlFuVNiw4l2/JQSuQSUai
LRjNMU52mM+Wi773vn55Q0smqVL8YM9ZDlY6sbjFtgrmkSCmD/EmBO/9Tx4BTYMs
bkBzB1LPMZ76hybj3YTKZenl/RVKRvSACdh6rXMLHTKH5KLKC10Na8mrdjWUp1yH
M+CaFwt+KoMFaYKn9pIftwWu3tSKyYXPCuIaV2FCab4aa4qGiwBm/sjxaGTZ4OPY
sMwsNCK8veW2T7EmBX8BRRv7KsJ8v8oA8m4Ss5Hh1EEnbmDogxk+Cl6HcJ7ptBzJ
8Rfg299+sGsvGdi+y1+IUp0FcklPZOpsFZ0u/fe6OBpV3nulZokhXIgZg5v19fjg
GG8Y73YUP8BJKqxsyCylAtKdOhEKkn9FNqUizpfh6mfk/BVSl0RydY4aAZhvBcyG
4nKba6Kk4seSoqnB2+AJIWy9amvpwz1oPBunQcHeBpUnCMmQkSQS8u/eFyD2rutX
fKTy8hchcU5mU5N0YQm9vP8EoQMfQXxd1TAtSvyK/aIhu3GNHks4ej5d0O27Ej4r
z9u9qoK09KIiWt6MdjxaUT6stKPqP9lE57eXJlFwUDv8/QG+wAFs072pCPUp3dJn
4wdBF8g3FonG8c7zAKbcYlIiSnearcbAZRCkMk+HiBbiAaxbrr5+w+bUmdWYU5z6
tbAjMyEGbObzHwNarvKxku5tp+82n8+GQawY+HNzfnw37ght6yKsEp4H7D0GRZIf
tXlBzMOlDvtfahn/S3zD9DE6KsuYA22/8YcgtFoPXKYMPnq4Amtmpr6R1k7Pt5SZ
yNb6wT8Jsp1K4MvM8jvLXNENtm6MWVhXSQ0rc46Z5NIuqfB+LDCfdU+UskuXrICk
g7O+PKXiEn7JIPHF47xEGY3F5eNlY9Vx1YL5QAtzcShgzh98ytpd3DELAXrf9PtU
xbkLvwCeaFFFAv+/vajmELO9RBXSuqlqFMh98VyjQo5H9Do+9LVBxDtNty7RKtAn
WKUqQhfiddd5DvhvdoPQtpGA8mE+FNBomxl6ar2u4g8TCs5hThL+PzXCnYlQnllQ
t1kotzxeBAnPVUSkSWbvpRzEadbBQ+wz8a4hUwEsPw4oMPqsQ/L1h3VNsKVPmIh3
SxWhOz4tFbKUOQmrWtmI6397fZMu9z8Z8uBFKblnvCtec1FZC7sPHMzCIH1JInOS
kB6pqrqcx+Zv55sdkAQPOmTZqmAzgEuib07W4wSV+cXRhAI88lPVUbXxjvqbh9yU
5DwPrCmQd8diH9OGzOQeTeQ9e+I9Yferpz4CN7mzpnJACDmkAMwFLb1AGXAO4kwa
Emz7719MQyFoaWgVuAnvtShhAnhEyND5DlJ7U8uryNSq9OOuWRNUD+rXdZz4gF4+
elY9v82b7c7SXym8IYyfnrVtw7qKGqc1iz+6ZdNUH2EbfWx7+GiHoO9Dsgwz14wZ
Ci70t8EhcqFGqa8YP2VaROClfHReIij0CVuqkakRTqwUetjCpQ0s19kBJziXTM08
KLwE1cp4dSiI/a9Tf6CRzLpwqqi4KveZv3IVSzCGHh+zyXhXKlFe/+vLB9Ikaq1z
HH69YCMDN/rY/JWNzQqReYR7I8wD5ho6viAFHanFju5ObUifAugrmDNjxtKIorzA
y0OykcIwuQOiH6DhuFU6rOJV4+2LcSsCrKdPlGnXEK25tIUk6AxiGXNF/dtNf/st
rhxnMl+Ue/QtJJ28yAC8poDrrc9wsxCdGDNG7eATOfuAMxGnf+3G9NWTnWHgFF4j
VL494GUcPTmlNVU0Mz0viYAplQfM9s3GHY9fcAn0UXY5+Uu7BpmuDFiBm5Y/in80
d1Vwvra7+3GCfQ1cSiRR2qtpCI97HVj1qUyj8MnMCv+4B1z8rdphhjzBPGZ4PYf1
tG/RovxuUdCvp2725scaM3oS2AbaaGkriOj4sDYHmMD0ZjyseF1mdMiutbFRaxgi
jK6Cigbi1iw1zeH301fIYzy0bfn1roYyKVZA3eWhD19D4um41ehMINaQB6hGfkdT
whYUhMlTxyaq8DlGRAKIpvUbx4aUD9KUG5WKI0l4uxJaKH0h7TVihAmhtVcOyj5b
THq1bLcptgg3Vc/AiykoelrUAxley1liBYoYuwZzaNJPzxEhzHC84h//ndknVbqo
N4mYNr6scPbt2CJH4XKg384X7f926/OIlw3B/ikCndF4GW8TILr/ORSENhwjJRg2
OO56qNQmuS1K9oWUrpZhWAbv12V/sFtPZyDQzom0Bm0AON6z2sr4gjMsi6ES+E94
4RQ1BDVDAKj890zylZqH/zRIqQ1NiYqIc8uYrk27BSHRJ/wKgR39aGKHRST+eORT
1N4nV7du2PWc1ue3rarwrjGe62CBtIDi/U9ot6mIQi415RF71phA2JW/zjb/BBoo
I57Xw02w86//jruxXpncc4SD7lwAT02wiMHn0m57DOeOcZY3yr1mzmlZGoBo4s+k
QMtkQ6ASd4X2SiY7B7lJGty/6QOohsuaIk7XoamxwVEIZgpwhvafxPoNVFXTz/gk
g8UuiqCmNTS07KUkyj8jieFsUHVuPuqPJfGkeS5f4qa+VaKEvUIIXmGBmnlvwsWG
YImMSM27JKO4aU2qXPfZ7TAlcmyB1yM2F5k7o6Aa9PLRA5zqAdPMrT+cURhYeXky
otJC1/DeQqhWbrrXwEM9M90eZhrZqn7vOGLzJ92XDaz0GSHyE4I2LcRvVk39bAJX
6qO0AaHE6jyqcHbfXt8TGiZacfFxAUa7fUcjkT10u13nMoLF5Qv1U9VNd5cO7JyX
9XOR+7xWUAh04f9x588N2s4IrisPGjfjvBQgPiOPxlabaxf52y966cqL3yQWTmEH
UdhTWRP2z7yUzqx3n7wpVE7yTdmS4p+koBOJZFnBEdMiezWIW3RAK7HaCe3OLt5+
Fy8I7SfFpnu0BIzgPP1RbZxsGib6aMGTaZKxmYYvZbfdyGTUgq3Lmup9NCSPaD7k
IDOl3TrBqZduaTHuxuJg63kxnHwsMA8uj7h8X0J6h8kH3j6eWIT67h3lRhmU/GA5
mEcvx5gW1/jA/FI7ntpkzQxxgrfp388wzAmDDjY1FPd/eTz92EEMfKAHQ9JyEZL2
ut9EJvfPhV9Lg+s1zMp17kDlPzTo7AGaCad2N5IP5BtL14jLrABxIdPk8p06zkWI
XycVTySAxxH5toQGWBwBpprnZF5RUO/Qo9t1L52AQBlNTSjnd3+mWZoY0MTiFpyl
h1id2zGeH5LMTPlzFZGB/MX9WzLtG/ZL8kdnmi0uQDccKC2iveBAFIZbdr6z4MSz
BgHgSffxXiahLrSmBb/yvntMwd7vIT+RCjyHH97qrxnd+4KJ14QyqAN2QF8K17c+
icxyrQu1ahZWgMJYpMrOgrdgbCq9RqRehlpJ0D3xQflg+BpS+KSRj69z4U+/SxCU
Mb7h3qqzVMhlpP/eHJFqdMeT1Unu+XM7OreVa4VJPUlB0CqigZne354iJq5wteL7
ab1W4trhkd1RSv9uuDSIwMGEYQ0SBHXGn95IhPH2ge1KFUwGHFGrYrK0gR+1MRMk
hvzZWQzoiU+iWLKZta5ENW20DciBIJ6wI422j77j+0WPOnbsVGC9PGIwLXko8L7+
2TBgo+KHJC9ZOuXn+BDnGVY3TkyJPcgXjmHpF6W9PCcuSlQZrKh4v+8yrLTB8PFn
YGZoVP033a+7kxu/Agkrc1ZVT35VOwkLb5Yp60F3ct/Tcw8Mp1BZ1GUuL/hdbNGg
ZXteyPeXxrRD2ls2zOKKil2GAEXljZ+yIztUxmvOEUF2EcrYsHb/3P7YNrpuPPDf
QxrhhNm1s+jzMAQmY1M8WcjgUq974hTBmXJuIQg0oqHjFUqOZynYD8Rrf7IA4y5K
n4DwSo8cfBewRBrnWVU6ndG7Gb/0Z9qvATqttVzL1OOndlF2QaS50fwTP8YCSBmi
u8tcxA8tYXq5sZp/C594IheZ2YgxnWj8duXsF/nhBBLlUjzBovubgtTfZoG6zm7Q
FGOftX3fgJPPJ2Znik6r74JlbMz5SEGm3/ir9ugwEaZLLmoJDnC0h0zAUwVmDPjf
OBhbPPpN0l58xD3Q2y1c0BQiUgIKF8MCL8Fk5K1Yp6T008Gix9BFljwcXP6RTUdw
ZS9PHzunuqQ8e8NH+ijF0jvx61017Qi9SK9MKJQP28vhTAf2Vm3hbfrt70R0qfIG
a2FzT5VZR3IQP0dTTrptFHlUqXMuEd2bpkxHKS31bikhSD+7pdNW072p5AXtnpdq
e7Dc2rPNs5JrCmhK20UCWB2+wTIZ4fG8VVVfmisUdsjbXLwwBJXFwDGZmQSwm91b
gJfHV+/VSRA4Hs5OSE0tTx9yznHCBLpVpAFFJdBB3vjsOR+fTJwZKBpVSQ7WsVAy
XSpjpwyjIp2FCTePdXETlV77Stwdu62PxocpDSl5Cv0/rJ+MeYpoyD28IlMZMGAR
avccLqHZqD9Ns1dDbhgEd7x/v5Q7bMEyuDCQxlSxSfxr/ItKG49H05YdCcIf85Iq
Dgjz5a5WZRshchSs26ba8vUYETos1zMmp2quNXEPMz4L++Xk13WNQ9qwQKDXmGY0
8oaydn+ZIUDHysDEIbQXHw+bEyAaqt/9g3rJoEyH6t/2fxyoRQADfghrmRE96TrR
YduoFyxwi97mlKExynXZCIYs3f7eMGbMg1OkljWUlu7bUPcdPbAevOlHNA5h+A0w
NAbgzQIb5n0T9kvWZ49EJNu8kIljGp8rmJwFlRWeBsFBoOb/7cB35r56D75KkJ9o
lcGU0vIyZ7yfZcHmALLh0rc8K2PABX2ZSJsrq07dOMAnXxZ9pbYUg2HBak9p5pfK
ERuFmMoGbs8coPe8UwEM98MN8Nt1B+FC6ihV6i2fQolse8eUVeAtd0GkzwwMT88S
jOWL+NJjGwjtCrKqm4VVMSAnsBQdao9UwDvtp93b3F1Q7Nqxv5MeXQjla4LUwwwx
/I+YatIAPTHy2xedygalJA4hgU4PX6fQr96brukOzhHpJ9pbamqN2EF9kAANqF5A
af/Ji+aNp+QDN/oG+nXgSwCIGg5zjGDuUmoJNqbh0OdoBRy3RsyPpjf0Bv1NUpi5
80lhGXl8pHerySGshHsTedjBsy9Gi6+BpbSCgl702IL6Yq75WTGMnRK8/kLMR8f5
lUD8FeOY8kJ+1MwE4GL8HyjQAwwcWnb2xnwA+QW6Tq3smCKscQYYfDSY8e8fO133
C34Yvn7R3c0/tnX6ZheNBVZKaZ3eUK7MGNC0wB0t1CaMMLoDLkeKAWcicNPVLO/u
IgAObsIgDrluX/jb7MSWATMq+rwt9fd9B1ykcRGBm4ayuCoxnV1vulNTRtDJn5X+
tYsLZTRYDrPg3TnfiCd0qdBf6KGFUF6JYZPI5ps/5axiUtQZWpGRIZBrwb1jHRme
5JDKdDEkb2WE0sGx+BXczXVTdqGva7fo8VhOF//3UopzxUEPXxPP6F1A9fgSQjT5
ySbG8QRYQx4syRYovZ4jJB/HFvHrOwvwZqTzWPX0cOwX8/LuyUgC7RietX6F9sO8
/V7dRtgcxm0muBfi1VG67VkwqLTm5whdpFkvo6doCuXFSXPx+ZX8us7W4MYSAfD2
H3EmDKZz+mSH42bRCjrNMzCtxAbvPMScdQWELO3kYn/HjUEq+laJLwoFNCTZzgeB
TXue0p1wU194LSxyCNLABVgoLVPbgMbyFwDXOh2uUWDvTMUXLPYyOktgs6JJVjV+
vYl22hHkUBX5KqIJWGgXRUfPb1w86LIN1dipdrYVHYXI51UO6gVMbkW02YU1jdGD
dbUN9gWtByNUF10XqIC9GQ4Fz0becLLhUJSNTV74RyxAZ2ybyDWb+COjgYvd6pmN
Z6+ha0DZYl154La+MBAG1/xC3SLp9LLJhlTzuCZYw1mGuHghHwKdVVnU5UxVtvQT
F2JG5HQMnmLyUmB+1GwOMB3Vc5+xgVD06NbG2Z9+YgTAPiJGGu3URkbU6JxfXofk
4UxCzVWyMlVL9C4ZVrITAsia8sJrFNMLSA+UkcxFP69ln0B3ALrUE7wnvKQj7Zmt
aGT3nBT4v6XIplQSCJ/6x03Caa/Rj1t6Emu6ubq91ybfxkyfWE2Js6wlulRH4tWs
ySy72OuTi7BPm/9lyvPed6ncT0kbAzmrgak4n6Qw3ikaze290wuM3U6RPhSvDyC3
1npcWhqPeX+xDJu1/Gonwk31tdRO2Cbm3OsTraHE3Lmpy7PQ+wETX6ulfMIzeMBu
B/x/LOohj11yjBnpWO728LzMlnH3B4n2zsnglyg+f0/7bNjWRR9UpGWul454Qm6m
H/hO1Eh8UShn/MzF8M22Jpp6FB0JrCLZhnc2NYi8Ub+aXMgiU8NjrQNgooRC2L11
9FjGPKNS8dorWJAlptc3sQ==
`protect END_PROTECTED
