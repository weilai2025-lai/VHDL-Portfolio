`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xhs31aW4oHPb2bxuWStv/gJgnVZLIYBJrYzu5pt2xiSkKPfuAnDDSs72REWgymZw
8fWifNYDFxWuDmEpq5UbR2o3SUl7vwTwRJZOjx4qyJDAdsdJ1WbpLqqNMT2/aRF5
MHAZNAunshS3wEApS4yYUv/vqcXsCOZTEsz5gyaruVSD7GyfTRxo5TJzmQxxd8N6
ZQ/bhZo6cbqAXKnWgqZGoduSdMtqa5mNQZBr7DHcUy1GNoeu46FOvNT1Lr3xhilj
PkTblF5rfFkStNNw+IdAUPtuQfg/J9A0Ql276nygicj78sg9kky0urULNf2fjYZg
iG+LnxpJsdgDx0daH7S4qwEG3ydolGqoX97RnKcQGt2M4OVGmbtE0kVeryRpt9Ty
qfaYCqaK37EWRrqwb1c8dAxZb3a7cH1HtZquJP9x7M5I/D1tXUavi4X0ylYIBmtS
lNrvTedi3SEW9FkBm3ehj/qDcEWSis4Z7YF7K6ZRs2wsSd8DUT7GuqHk5F7gjvE+
rwjFyJvZI5NYQlwuiUGGnO0fur0bFWEWwebhJqgcv1OUKP0Bv1CwM7q7jsQB3C4X
rGbl8ig0zGplVrxgu5DvT2XTRkFPucRvEN7ZB+CpYKhyZW+6q3ByTCCymgsx/AyQ
cMFNR4hL222REgWzkfiYOsnOO+QVSmRkTlZaBiqIaV2pWau2y1Bhsuse3CAPmnds
BUnwdTE2FpK7rYWXLTLNfh1RbCoAdm8ex6UTHjUPbVxwYxkdjTre6bsXDIOT90Lk
WhpJ/RbIgGmKV7sqUdCwVLz/tLBf9Kbciqc4e+JLJ35lJiKalERh8AQLJHvIARZ4
JgCIOtE+BcH0TK2hPXVzvlFCgi9Ewx8Jgi0gs9aZvzWdPFOaQfKQ52bDcr8Ktckb
z7LGOY8Np522lTAHzH5iqx3T0+Ly0U35yOReAjO9SfCtiP3llYgesUOcZqcbkXmO
hPKTpw54KFyUsi5iYB0Rfg+sIQPWlVcz//RtT5JPrgnxMuRa63N+imznI85Mai6J
iJ5/ZelXkDfNV7hqXK2Fhmq2UlruI8w5lpYlfT/koDq+J1kbqD6y6ZMbcXlCe8Fc
4tdDwRb7ZweMI9BsdK1q01ae9tjAjNnLmBbDXAD3R7q619bWRIsYzygTbnKQnr4G
jf4zptjXQ3HdQBEfEQ4ozs0A2p4bCdaeLyd8OF191k7/iM5pgk6C/zf/aD+quSl8
wIIvHYTh/7FH8uNVKtcLP8hIMBr2quH1LdBnnqhrhEsaqx43M2ztdxf5Aj1q0JkQ
d7juREAFl68/oaHlQBxSflv29EkpbU9A5vj7M9HLp+ochBA32Nwb/NsthsmupU+F
QqWxQoBC8leIbo8/obKjUzGXbudFqP6IZo9bZbrV3YDoNHb30pIvH9AfT8ZuzvJP
Kvg+2QlSW4J1B9l4/td1GebeeavdiW7y2oXqLzY3b/mQQxnTR9gJXlN7joXWlMDe
yrMv4Xl34TzFbdY5nSx9/ZgqeYlvNBBL+XYWOzGR/UyAG6wk1yN4mWLdPUOH2tNq
yCOgfRXLEeudscaZvTA6uEfjIb/fCGgeTTfGPaSyQFh+DxdYLccnC2MbpG3Qab/f
dhqa1bVSDWUFOYLzLvNe72QFitYp9w9ei4lVvR7j6vF1lMJIAKn0OjmDYg58NzXn
kP4B9vvMeTxdHhce56Mjf3C2WHAVwJba1bIotDYs21Hll1FAIu+CMF65XAnJV1yi
ma6UwfAsTCOnAqu8pGKfhtleiL/RycFLD8sSXelp5tjeGwVJBF6rptlEk4qj7fyi
5DWuLZxy6EDg/EiTOP9E7RAbwBv6kLceNUZLSPYxiFgHJE2HW/mdJYBgloDgnosS
/9n7tmgORGvzFW5AxFp7DrITlyzXkYOMc8xkXXzF2HiVReu6eWjbshzNEkNysIw8
WayTfk1HnTU3F9aFCYSgTkzhxLzIctHyrKb/u/CZBOF/NpnceEiNaY+qgs5+oQlR
uL5m8NilQMDwRDCDKSwprThXaZkRpirtpb92hGvHjc/BwxwcJUaxoT6wgfHJv+0Z
cZB8OQEvQyqIVoNS3MUTFU+McUcq3lDB71FBo4yFW7AgbcDl53J5KTPgLObPDpW+
rUVelU3ao602AB4THxIh7Otf3RE7FHBTlzLcSQfoLxGwW6ZW0Cor1C+TVKm+n0QQ
G22QlqoYwpjYUtr9qgK7tM+HXqqQfls6emMnB/s4rfW0PdGrJaueReWktbaFkh1f
6xzq3H1onJvVjFUNC18usqgHwCCB94GS50beSHQ5m7UqrB1q1336eJXTfeWXRRZp
TogH7+MBtSb9g1QPqKFn3H35u33UkMYOBUN4AfCBUtmJKeFzjX0rD6brn498IR8W
zY6xA+jhsKa3AAiviIG+Nk9DnELf6PLNOvSJttDX/QSt5P3o0LrSNG/uDw64qE+N
Jzxm1Nfh5Z5mMM7sRs2ZKuCYn9jKwpJ4ujpBi5p2ggvHD/M8ivsZThSJUZQAdYjA
OAWpsaNiiHG2+09BTaBBNppYuMY8jv4HVIVb4yPPYN7oFnLzkB/0pVp2DGBRZMHj
XksS4uREgsMVmsFe4KwoTSckGWBFlH5gecmw8zkBnZ7fem+LRdfFDMjX/b9rt1se
xPPV6iyoshw4PFZiJtig23++IqdJpOcASgQVnyfEs7WJy5CUcvd1tbuYc5Lou1zy
y1y/Y8JKOgURGa7HxbMgLwFjihNwg+qkbnsfHh1LESNopzxycRmRPLvvfkLjWVn8
iBqNcbZuPvvmlddz2mof1GYXAyTYOjyzhpENCFVr8IME3K1w1Liwt2L2KGmUtmfA
o441rBXvb6m2oHTfo30RodJLupSaF4QNTMja+11oBSAHJ9fk5W/XacR/Fpy5FiGM
tFD1Ohi9LeQz03p6LBOYII06WrwsUmpZRTyriMqlTz6+7HR5DcPmAOot5FcLkBm5
OZ184aeGC+O17JWM6qL61tdc2deIxtUnh63CBNXEghI=
`protect END_PROTECTED
