`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TegD6ntFTDkkCswf0eKbDFtcLCHX+H7yZQhdz+ig62bAAUjchPO/ZUjyYXtvJWdu
fF4VUnFJ+nMkmZIB/HaU1z+yaCnAiFXh+ypEyEQkcGSAqW1Zx5v7cmgKVqzVbsuJ
3jZ6fEi2u7mesBJNQPRraVQiHngoPz4NUkXLJLSpSwv27qpbMv9LcC9KcEVmqg+o
/aH0Z5B3uNIjgpW3lBxAjivzkfE77txpoOWlNR5GQsYt/cH5UFdy2gfdImgvcb+k
uRXrj9kOFF/16EHVQpAAsFPrn3V/BzH1R4RB8+ljkq/G0kFdK9K4RgeasGXiSwT5
uXBDO/Au0Kj5akXiXjy+ojXFr+Sy3l4mGkpXSvwx1UdXE9OsSNHEjaR0AWbhOS0S
4H2EuGhkTdUl3SIdGUqmncFG36A4i8OuYUpuzjU3es5x23lpKZU1B0KGLuLJ4Dc5
cWcXX0zxUZXy3AsPPuCMq1qDlr5s+vj1O48QGSotZMnw/JIxQe7q5eXcmlaAnTh8
EK6D4ogkS/kVnCL5uk3stvpnYZM8XGoXVH2/Z1ixLVcJgWd8YZcFyD9bpvI2obGr
FAvppVBLq4XTdl28jeBQM4JqFZXuKZ38bvCYa3RyD5hOSt60+EF2FfWUbE8Uv5rb
kZsTuJPPznWW0S0ELAe/+EEFz3ZVFT25IB4ByRywkKK/KG0m124WWtwmeVGGux12
acL3Yvom3ZFS14xD0TIJ0zNXVeVOr5YsoaGZxpY4hdrObafEFvBgDd+aoazciQRr
VFr6lzXCglbsjBtzgEDS2dJd/q24yqt/PxGXt2u3ylNbDiNvAIZcrrNwuIMUPM0o
lCiba4ns41pMb8f3p1FbK47iZktBtGuXZ8EFZKae2nhSpZMrjwaEnSJwDLDIthUK
a7HPbn2UF4TFPkxebAywknVCEC/V+Po8rIP0EETUZZfYOkAj7vIMOylm+kVa5PWW
PreasvNqrLXADaSy0IMyXIyccS+fdeaouf8dbkL7X4n82w64dhOlbLEgHUssjymO
sE35neAcLW7nOihyAPwMa7J1SlGo7XprGFLoaXlEnycnYz6p1IWGipNumSciz7kO
xwGguG3LNxZeC+OfWOwT04bdI/QHCJ+Ov+neHFrmhIKHWymTl6R1t7/rJ8zgHS7Z
hWAwrFsD83mSzq45CQfsW7R8MqxT8mO7hYHJefRNmmkDdISoADBjb+j8/UnT6DsL
7mo0pccDHs/cbbga+BwQSA==
`protect END_PROTECTED
