`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDYXO8NlOln7bua9l6OgInWeuN0obWrjrD7BjDtFAmJW/1wR4BQv2NOOFOO2Kjcv
I4GJxA1RGTXfgtTZ11RjuN/Uo+zrMbh+P3+OvlgOC6t0Ni/6Dn17leKu/gyswLde
vd1PnfZxoSLkZ+rg0pp+wqhz21sugS71LTgTWzJCKMPHNoqXFFFZrE9jQkpFYE7f
jNe3H6/F6JxkqUMgbv4a8Avitq8b8HQOPqUau1HIT5hgNCbn4maxhVi/SMGV27+U
LriVMWD0eozUwjc2ME5Mz8JPVuCZ8kxiKKVNjpIqZ15YfLPBIKb9d5DX9IoGcdLa
LiFi9b5lfuuIMF5M9upbnaW/6006nTiNYjriOGrj2+PI5zNfdihcSO9EGX0xYQsF
`protect END_PROTECTED
