`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3MVK85dhbrr83GunPzZnJOJ7jNphqBBVUGwGg5y+mru8wnlc7SLnw0Er1ZZmby+
E+ezTez5aBzmYPUaWVknKW6nMP8zejwl0k0QJF41Wzpe1MecMXwFqxmPQmLkOtQR
zi5I1LqcSLazfsWvTrmHdUqeZ0GKlq0thTw85sDgDQUwnwRBnAbA0Rx7SmfdEo7Y
BSMEjRWmg6KfoEJPXkAd3lqUyzGH4UNhkNUO+XItwhpxnZCRPJbmvLA2ktbFlrZ0
aeFC0eS61erMlVY5wDcZMTv8h9XrKJMjSMG2wRRCfIpJvCc6awmKRv4xQ8zb0mqO
HxjhLr1l6msq5eiWQF+Ly1WewAzbbmd0c+sMWE7ONsg8MvrVrsIfhtRflPyERSBA
oMh7vpJDvkHAiLXhWrfs1vHBHcdaudZYswI2v15yon7/ncwoGE7ZxsmbQU+TNvw8
x0OeV/sjSfy2PKd2miKHnq2Hy8y/woQTwS40Sa3th/SMUAvcuuz32qlmtoMVBOiz
wWRonL3a5pzsH4sIsWcMTxFaD3WmaE9yW8z8EqDvvNFooc7LBb1t+gVLCRvBQzCY
uBq29ilqN/PpLSJOgDbC6K6c+8qhcRwGHEITCWFRDfsrbBDjdhml+NsaEX/4V6VI
wEjO7f0Z73Ea7P6BmDRkJds6PE7Bf0wSx7S3Kf/Ho/OnEYyuv9tHebKFNEFAPXJL
dukD3vj6XNlqKiLvfBnJu6+cVoIudb7abZ1TfB2lbTvDbAAOP8GIa2M5BLgETcK2
`protect END_PROTECTED
