`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9291Sq8V4pPlmaFsH5IVMWn0w0pytYmDVHUZgmVQswR9T9KdvWmpuzfy/sbcorj
6rPtOQ3dq4nqaZCgNs0MdM/0RPZel18bca+i/eSmdTBRY24zHmWfkMkHARdONoOX
GhWACuGaO1I2BskIpjHcDEQUgHGRGtKn1pqLMsyovOjvnfKl+rn/xXBkHEXFZ27W
MZgflz8mUwLFX2RHjUe/he1rE7Qw+Y3bLJysKqLJ6VC19uj59a34ICTYXai0NnXy
u2wzcxEnIHFNtNNh65XHY0P4bPCFmNNksBancp2A2U9eaunhSEVNCq543YEpseRB
zItYzkGZa97HjjM20kAbuIw80jyZonYhSQU8KBywMi8hhKqu883gKsJs8fAnN8Hw
m9vjNFJlbsMVOGKWPAGkyMtWVTk3z0YxxKGMNPijvQ5sDijFiEqGMjTPfRo1Cphp
LntpwOMD6B/yz6J9tk4mE5Hk3dTf1IJvOYOSTRLO0C9yrjUksBbT16W7omencHTh
c5IADbEs9bcIbIiD2POcgbZoXhMTqDYh9RlBw9efw0Kovduz4yHRbapYbk5IzhKu
Uhk2+zaWZ2ZcP2chVT4n5J3rEh06OYrI4A9zrcm21WC1f7kFcmc7E4XM8Ase6KOW
2rJmiWdNdkC2Q4hAgw1OFRzJstpmjMXHRebR72pvCUBOZtTatdT5fryrDFsyxl+M
4slz56CLjuGKDR2eTsc2qMYm1KhwX4zQqKziM3RyPuZS+aVI/fyozzrPGeQ7cIo2
RgPrJaSUSepN4ZQbJC1muljORZWXHHnqegMIaQQsxGo58X5GQPkvlrdNEWppkER4
KmN8FuDD1aveD6AB00eNkPzGf86H37oE8mreZoZyVGybp1PsYTpYSZdpDouPqcaw
TZGYr5Ar3XM+Y0nHMFFeqj3zyv8nDyE+o6/m6m4cAM/4VtbJ6GXhzK9upz+pxCM+
ibZsfvCXyCztnnB8Q78Now0mTu3y9EgtaROJdRebWL3uciNLqDsN0e7R5wWPgboK
aDgvS6kYel9JwCnKU3jxxbqVToJVCt/w53j5H1P0iLGIg7y9aDR3oecbRxZY1vQj
fhmaPin8eOvp1JSgDsXPpaUQg6CrPldKOTdVJxGMFwH8q4fi3uvfaY6/ltAUcANR
pZfBx4lBqzEXAJDS5h5m3+DLJZh0P5nKp6CdPnM3WjA0CXpCcRrrFQG1WpChvf0k
qeeOFHEaRkP5Tv+1wP55DbrBh7kQ3wJ7H/3d9qVicch5/TsKen9kKWxjBupp7FbL
GDwYwkn7UCd1gnTf/IkBdbZDo+4ACeTf68e8/J2lGJtqm5VqYvukINkrGtoBsSFZ
3kUAOu2lvFXoZjW4eoGc+lkmQ+UrR8mlMcjgWobfAvyjTBwPiCIXsdZsTMqRf/yi
FRbqCDAq1Hoetoii2lZbNuDcPnemTjpCFgKOpumKJPAWk0mjwSI9ZxmPT/31Wzb6
px92HRjRol/nsxh2UlfRuE4k7NZ8GSbPcJIeoaRr9MtZ3GGTYRoOBg0wEmth9QvP
Fv6Jkk42ymehHgcuM4p7x9rmguJfU+yXGv9o+Dee+PTTKC6kJ9sRcxWuvlt94TNa
dizuwb/jg32a7m+lcXfJz37DpEJzMBdofP377zdkIOIe1K0S8Bweu4E7+y2NtPgf
AxadOw0BuLfr3mgqCDU9cwnwbvXsTrG8djwITO6H22Q/VttQNzevLajV9agJd7Q0
v/G4YFqjfUcxV6frXysEMHp5s+y0ekeCVGDdJBsQw0B7BAEg8+ar4BX/B9oQdgOw
yydWdJXEbg9oJIc90+/gfWhJC3hUBW1YCtE8TOIFf5/9/Bp8YhoLxtE2548D/XP0
x12TK5Ri2ocVnhprSFkmQYXFf7c+bqsbAObmvqETazU5QDIvHaERpT2rrlqUaoQv
/kqADkszCQsvYBe7FgoyO337PMffSOJYxk5RYmO+imGR1fDhhtn5hz+zwlX4ID36
uV+lgPKICph7EJ70eE5X6mGQq0WERHRS66EeQ2AJPST90FVzQDNGmljcEuz4pJaE
c+193PixVAVR4XD9wc7UeBTES9hnwnatL1XlQjvnu83tBNJE1UQM2YpP54cuhJQJ
rz7fxHWNRXinkV5/74xwE8dsy+Ol0/w6wV6bCjLdBoLs9PiYh+bcY3uFsl36+s54
1ol/iulktRaF+R612gGeeg6bbccQPfQzLNMq2lcwrx2nIw8N/Mg2S2/DTrYL94ap
X7t+Qt4K3yD9ws6ce2FNqSuiiW7lRgGBDNgtYKm3Sib3KATV0a3f1VMEcuTz+zcz
eQTYKW/NGb2oQVYIiR26z0bY7jIK8l1PTdIT1oyrMc0O86YUXKoVOH7MS0w6/+V4
Yt9eDOvGIhwkGTMIdtQYe+wbowKDm2qB/XQMzF7ovhj420JfFMPbWXv+Yd0COHW+
Kjg4V1uEVXCRZAasAmQsfTusHuiX0aPURsV6u9IVctVymRu+SHqd0jCuu+NONBCx
u2sc1iGT8MpStvK+nxldbqHTxe7da0ouatGbM/C+/QuwLWfqyoNM7ep1PQCa0Rm0
aEzVXKWAGLqOMMB53MgSO14mR0a0w5zqSFIrzIs58bGRrC9lcR1tW7toIpH9Kg5T
40NzOU2RZY6x3AmZAUobUUMgFPlNf5N7tsF5huziMcNFXY/fsl0u60pNEvd/JSt3
kii7pH7GUcHxJE1sHgQ12/Hz7uRr0upH7cRsc9y7i3oIC04fUPQteUkOi0qgXQqo
UDX1o7rOhwcmzGBNItu/ZKL5Px2zvZ8UcdnHkfJdP80amNmrTK+C9vn7hwtt9gNn
RzR+2OC1/Jl7WeLHIdGYt0/GEWW/a669LEm7v2nzWsYK+ZBEqq9lCiAGeTlEGV/J
nO63K2TMSngujHQOdPketMU6heoYI1UE/8wPmE9DsiDCaF9r+woicXmqpbhjSd5U
xA4+yylQDuSpLUmkofxLFTv5MeYUiHi6GmpOglYFhAOInsMBsrkrR8hlHsZbueye
9G+0M4B/BYoql2lN7bHWpP/DTbulT4p0/ldJdKMxHj/zoxDXG/UglrflOpEgcYDD
gySpC35gNx6V8pc051W2LwwHNUDbgqWY8dZ7tIccEgb0nETShSBfaAGNsVwgaCU+
oIXfDx4CfPm7XA12syVMirVOcTQ0a/BHWy5wXEbu2VtIVFH+DwsBkHkkiN9EOLqW
lvZOmcqRSK6dHqCKrNCt3ZABkrzyYHBiquw1325Gvxn94hDdIANWSy1Bf0kFsB2E
ijYOmlQiGhElgGcwHHgMsBgNsn6vvJHa61yiirMUsiQAE95yR1/SyJ41swjxU+Lu
nJg7VrVbOUU/GbGaHVRNGNe6GQwu249Vi5R5i6SkH1HYHhG1zX0NUAlRGGXQawSE
/daShSVGU2sPNawSBr/nTkmaQXA/ShC4NwZ7Z9cW8hRRWL+k6HJi0CvEt+KM0M4P
pwUCXG9cHEMo+1UColDwczVEhY2cZzf3y9L26pfoJtw=
`protect END_PROTECTED
