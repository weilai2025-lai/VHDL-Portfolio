`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWhLRybYpBUoI/d1UzXUKRLYMAkS5CQ4WlednPs2hLkedu6LwegFzZVckFlR35l/
52HVaaudw62PglKDUhsPn6uUpqMqdS8ZNiBtEr/Yz4Zr7I8myj8mklg6X/VmXh24
cnk/WTfeFn68z7RXmdDQgzto8KHeuQmv6nvBwE8pwnIYKTwN1kw33Hmc3rbMV7lg
qpGtIw+MRJUOfh2mAt4jef8Mjy8OZwIr5MpA8/zz3AgBweJXFqZrg+vD6UoD3mPC
KRrNFMwupVYJAmcDZ4BaWw85pSh7y0Kp54N4UYtZv6Xn5/iUKUlrleT8g5elYYQL
xYHoNx4ChXlb8nJq1muAGO4gahwtTGZf3istKha9Pxhz+GKkAoENKZ9Tjt+RkvHA
Uf9GgBiugdwL9gvI3TA8dMuwNtl6snClvkQ2yxcDR/HgTG2HSE+fXhFVp4jODakT
kyuL7MG+GFmLk9WhIK2vwPNSrkTwf1ogXFL7KigekdNyHiLF4PMBGPlDz9IsuL+O
iyN64KrSktsmNOqRbR0PqMasjM3ZrD8Gj+faNcZpzmL31dwKG4+RmSEPi7GqISHa
ZV1BH1CC9idoq1znUuMH4euwq6oecB5HrcpnkBPpZ7Q=
`protect END_PROTECTED
