`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09Dv1sXW2avTGAdgYZpowFxhrCDC6ve+eMZ42bcmVdO/F27pX/TYqMG78z+HQqB8
uRuf/rHbSmk92nT84JsVktcpIIflQuWrnX49md80UVKG2SnLVdOItEuAKPK94ExW
KQeQEgEc2COWtMYHgRgtSlGGXRGvkSGMJiqUV4BQnhpyoGZE9C/lSEpKVHuUB+6h
6PWAKWUvMyJODWH0dfbYqwj9kr1iGyeKQHXbj9UvEgCwE043Pj+fbbZ2XHPrieCQ
afXenZh0NsUpZN7nfzRiUdsMF84gixNOZAKO98uuGrsH0PsN46V+/N74ZGUie2WQ
n8NILqNrgHel2zhtPck/3f+HG36yyYxNyYbM42gxPaFKLPzqMIwuSkSLE0WkJ69+
ZKVCfmmHa1zdkdvuCH3skLh5olEmdSejQe+pe565/ueN6MsnyTK+wS2jHb8kdn00
98NnhTQ+ZHK46XuDD6Z6VyHMk6+jN0uWrfLRrNq/ahbpFCj7S/AOzxLbR559ekbE
BHCAPwuutzUJOQFMQzDO+mwV+LArsaQl7soxWqANqea9LnY6I/YI2k5HPa10GOSM
Y9XYkLhiBEc8QNqRR/atBrJ72prrR8LpL6/gvQAmYM1Fk7PAzSqfzlxT6HoRutQr
/VjU9ovel0b+nTqf23mFTCLdc/BovVKvebpGCGskDDXFxXI3dnqihf5tnYY+7VxD
GccXOObCNeeopuq38RuEFEFjSAcGWecyOoQ8aWaLTfLNtw6SZb9cnKxiKtph1SEy
6kd2nL0OFvfoyf2ncCMa9+XGhzASymMwNYbeGHTH0f6r2Kk1BOBq0z/GqUydpKUN
tB62sf5PMzDwRVZdVdIJb3tZ9rCAzUIfjsBipFAb0YyFVvltwBFeh7tQxj4Ir+qN
weo2RXdyX93fHSEsm1o09E6w9iTlNh7hj8K6TKISlQGe6JzDEq8is5XXTBaGe4lL
4ZpibAN5zNkPrS+RHj/qjg8aAC+tzg4amQ8Uglzg4D7cdCwnwoVrOwR5UhaA8EJD
jm2H3sHtSpdBtWwSguadFPkgE6w6SAFNxUQ8VAON5Fb66vDOl/al0pdIKivbdZUX
XBkO3B8VWyjORBVidUzaIenTcT3ilHRPqFTud6zDEoRvrJfYnYONltxj1bdLUqps
Z+qdN4S6MAR8B5AVDEGO9onq6Ef9JZ1AtXWmVa3H99jm8jpTFw4QvrDv0Gga05fA
Sxv4xYThfKlN8NNXlQSCZ7eHc1ENNY7W8bSgeS00cYO7AP7N9QPk1UvWOp1yAbAK
cbcepxKiFnpH9MFoojWLsOvAinyV1UVKX646jYum6IMoTJz7bKjlOWtOa35DD+Mh
nckiDGGDSnisOCmzoShvf96AipqLw8NnRKK0w8lxOkL8Vl+o0dfdJzpSyZCBnd70
KGYFABe/aLyoLBdVPxWxf1cD4ps7BmaRGKFm+ZIgc+TzwEf5Y+WYm5Gbf+B3YQhf
96Sx3bU3ohBJbW+YK7AssEXaFNqfZkzuVO2NqbxWc05m9sX/fl0yDtn00QNDuc2T
hA5GUZJ1CDGCSpy1DlCJdMUH1ywDWa+glQEn6Liyb7ifZ0h1E7wYQsOLWcX+XaF7
9oT9sRNdO0HijeH7ek1JKFGwJxr9zI4NqwA62rpahBB7a5UaFokyCCqDUYGYSUSK
coYgO42k7JIYA6y6KSki9idHs5wkyPxQw48uGZFgcv07bz6/4JL/fK0LWxY+WYxo
+DERfHz/5rX1ykMIYBDLcCHA9HdwDLUP++JXQEPxb7S6wqCsKuS0hHONCflWOVnn
XiMKBalWdNzXj33JxMObTl0VfFunXemDG5XQJl/TSd6bMO4GseE6CWKfAeaiBtTb
23G/FdxtD64+xZlxldlzSEFTrYy/pKwHHh/s7fqEaafti2HDcUxNsUczePmAbCZj
IEc2jvVnKe1znJuGerQS9tzsO/ceAwITpXwmK9tkm9I/1ln0A0p5rSNUUyTz+mDM
V5MD5aS4PH4deNcqSsMlFLpog8vFrl0Gd0w74L+vAOkU8D/lPW+L4c7o1pih3uRV
QD8YvWAbRcDo6K562EYboUae3+7T2HMFtHsL/KRcjkK3KCqmPnemVm03d8pvRMS2
o4aOxQQufrddgFmqsfBUVrlMrbOmr2aJekwnn3b2oHe4zKrQpBKOPP25a9NtJJBV
7Bc7pcBURmWli7iy2V49KPy7Th4VInXiFfLHzG4dAF6hqsB36KP+LcpRvHWKAgMW
g8Uapn57/6wEUEQ1dICW0PYyRn8XgeYcioLvpG8G2S29+rr4qBOzOmRt5s0c+ENa
CA/wB3xI7GO73k3uygDG2XqtoWpX1vHYUgOGmxI3uUTssFOKMG4/0/YHtE+tBqRP
qtWaZQV+sQVgVCXdHaY+lmGcx3JotENJbdb/78Afim5avcsbRBYmxAW7P/Zvy2c5
MNOOFtI2VTI2x/uuj35TnKsTE5yEdCY3iMWRGmgiTUzlu0mzx3xQKRv6XcIVOKTY
NH25z4EpPnnz/qyTPtrDMXAYT/J07kMRmCcN2uijndcD0h7GcnhjySyGxvlb5CRM
WLLpMiIB58RCk1mU04klnTMHpmV+DOL1R/msodrZuopvFJtxadhT58un2purEtyd
cuVPzJa/3GhM7pLT/M9bhDT+kN0ipeRBX0R9jmmilx5yPAWBMnh00JUzE0X1mM4q
Xl9lFM9v7+iD1LzurZQaruiJgOP5zUj5dZ0EB73GqV67r5A4sB5d5K/UtzO2TFRb
R0NQnIh/IAtjZ15F0hCkJ34bsWhTjsJo4AUufwmdRW9gnd0grAk8s22KZbfjfyGZ
OtJU9G3CHTj/enZBawj6BjrXlsSCene22yfNwlU7bpKrljkmnJSBZkLtAmqL0EOE
`protect END_PROTECTED
