`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uT96wHUjsaKGSe2l/nCx013G8DNV9F82ILFHos/ILJmG4fnwyh2OnvmgF/GmpPrJ
2PcazsLnHoVhh+V8BoSRfmnp+nj8Niq/8daW44Gs4vWbPUEvxX30Nho7P9BfZgSw
L2Q0mpP2l+/4s4vquIOHb323SWPsdstYbgW8pFupogyOdws0IzIJmlY5i1fTLPxx
3XOOv1Xwj2n02tRpXQkUKaDa9hay1yr9lnDiRsFtHV214Apv68pMNZ0/l7wGjKCl
HCr5gb6fSvRfH3WxCTC2Zn8cWA9jKgzc8qFbu5+bJ7Rl/VupfJvx+NDq+iU8mEqg
qF3wJIzUqXDAZruhFkjP8LpsjuI/MMVUW9KfrpzriDQVhUV/pHHm4nqgdkNgj+M2
NfLHuJUSWdA5vl2ed1PplsxmoRrRtF1lqLZlgsOGPPzUBdcA4I4AXSO8Ho3wAtsN
CjErx/q54oysJfiryC3UnWBL+3QJwqSeanYQDXMFkmUEHB18xK13lwGBDI9Mt1T1
VLw3r5qzKgDUnvIOlfc6qmvfV5DIjQ7cC6f/S97NGX3FmMeTgyC+S4iFedH3YIhJ
QXYPuSzSqLlVM+6n2STx/lPqik5n9G6C4yw03EPJdqb5Ye0fanC6goT8CQc4Yd0Y
wTIVVFsG1MrzPZgGV2cLxrFl7zG2G6EyoICdB/GjP8eAujdJ/RwxI8C08FveAANU
5Uwnw44978k+9+o8j0d2IB/sRfncefPTw6sCq4VLaThl4tlU9NyWAAOGOX/cYcVW
UkWfB0qlGiSLlhsRzyRdQi07FjEDWJ+KigKS5OAcd82zfvghlHl95p3G8Ccrr+i+
t01JzcC6QLp27JCADNqDAcfPR5yXYBWvxe6ittdDJ5VDCuuEvbMSc82ub8ElJ1QJ
fXT+xLzsvOlJ5zdN7ap2xnPOSmPio3o3pPTjhhuyeC/B1PINC4HseZopJ9wrbYxG
kmA1XBc6MDdpyZB1a7v9TEapgL0ncdjFcGV364EhsS79QwkWQzRA1PnYHZGsgJe9
9FJXK1MeDpjPw7pMQuhBUstTiUypZExReokMJiphm7oj+dT46GUjuRG1MqgDpkRv
I6A2cmhJPrq2OHF8MLtBB4R+HWstO0Cm2FOrVjPugmhXA59+87JwQRdL5FH9kzQp
5jIs2XAQascYMgAdeeCVWSZIKwzXF+A8gB2MspxCB5sLaqwjo0nImdgFN1Fmc1Av
Yza+8qRSrPE+clAaNNMMg+OHTtA+vRk0/kzYIDlstgrwqqVUOI1TXSQj/LDnMim6
iPbyfMh76fSaxqPZ3rhLYDWR+T5NZ99z0gq5N/2Do79DyimQvQdJmdG5IoWZwKtr
sdHj0ZIhKOYri2Uzkab+dg61Jcda5eWmoGgn/buUswNqHhwQzOvmTD96FQaJWjqg
yD8PP8R8+e1Johyb+XQZ3txWnplxhXssblF/8UKPOI38DFxAHEcwkf2tbapCwTF/
+FdEl0xnqgg66JLy1dQmVGLLgIzdf+1k6CFy6zw2TyGuWutcQ31e/ibsrrR4vLhp
tb9iuWH6XrGeNdX+gmc0FufT/f8P4i0x4wbs2EO51gg+Y5zMEbahGHOOf385vALz
R8HMwpuGKMiJ74n/EiFqvyaWSdtLNTD1GWMgkRfgmnQnfsR9fB9W7cs8fPLpBgli
SdaN4Wk31d0LUyiM3jOV2vvt/wTumblL0h0b5XWyu3/9WQmIrqIposIovvY4CAHF
5G9e5KqdPZXvtF8OCwR6hPyt2IjulRCSJ1yaY3JCFMwMIlH24S5IGxN+LKyAjwTt
V9GsDsGmriQZqHemF9pgO2DIFMgoLuEomlkVfzvsMReYmQHLR0l+6XVOY31+q3Pn
B5wKPje4n7C+SRfJAjwcylybwoYxb6HAnSq6bWPQNBcfIAmBobde12kTKfCJfz74
fwQfasRhnTDr6X/cPFNKiUQ6FPPSRoGfFCySRHrdWBrqKm+RBLVM+q3kaC0+NT8K
30WtlLvwYgVHYbjHhdCGk7wyqgr3UnkPK47+xE0jzsCzizY8U6imaJNgwJT6vDfx
H9FkOmsOhk66ocQYmCMvjC3VzDkXQmwLvf0KJlGQ2Mk8N8BRri3zCpENnknHbVbR
AbwkFH7FwXrhVACIemSPiVT6zOYJLf6QFl4CBC3sA1epIkG6VhkzadSIn7TRip4W
yMvuF9BCbCFvnQQid/DeB1Wr6qTdtrmn2miJ3luA5UZDNkwZSRgvV6r6WX2txKma
fL/G1UMv0b6/4W+QjSE8VetOU09/XBoW3HOLbmpH0lwf4GEH0JoLiK0fuDptKEWg
eTUSs3qsPybDUj+Qbg/JKKT362moDQ3rfcigm/viqN+kXMtEa2neNzKGaxqiwPZn
yriAXzXlrCM2r5mqjP1Xeq4H2pXmIgODsq04OWQUJpRd/uMRzAT2+ENdknPcDqCW
vp5BZWUQ+zTGceC9haIzglZCZDoFBR0e0VV5wGuS//fMXURSHMGeNeFAxJBzJmmp
bRj5N022WMjIrJ4G7rcXHl6XAlSgl/hZlPSEYlNq6Gb0movTIG85pHggqtvZXYFC
CUloHydyyphBzu/LBJiuao2fWKszHQ2rgAozs++yfGWJXpUbwHLqbjKeUZ3bcKLx
nUrpnvhiZOINoaQgrIz/xYtqRhVcQGw0hLPmaJVnDgQK4TA3r2MnZxIsenS8kaP8
vEJPVwI6+AhyvV+yEfN9g6GFug8eMliYI+MnzoWPxMmanatuevG1fSQrlCBTIz3m
Vlj2D+bgi7FBTwG3huN+evL7D0ojZgPjLIKyaEHwz/LgJWY88WufMrT2BKTFrzCa
h5TeOOxWcfC9+KDDV6krDuqMHh7ZzLtPwbrKEiZWM6TuFJ2IA8YIenZvXdXarkpD
sXnJZhwHn7spp6jfSaDMZ/KDCWz49I7WZjK4yafjPF1OP8Th7z9OeS9RjJU+jbqV
PY+yfSjdxrTicBg+Ihpkx37dhoILoEBgjb32+VfDAo5dFLr7La5XLVHMMcNhbVPV
wbKqKcDvifpSA+rQeqTg+a23wpT8wD5w9QpqDoDpOkEdvjFt5ET/Zng5wl4b3NC5
C8AC13h4n2vncAWrwrI1foEUHea+BN4vKfvBsPpA+CBBlRDwO9LtBcTHnwbgvw4k
vhOONQggUJkybBgtEaUnMv9Ki4FlmNg0/cIxKkcFrcBX2XlviJ40JWQ9FZvMT+7t
8flWeQOB5TaC8tO6/BGlA1z8EucqwGsrqo71Zk7N40ba17X7kS5l1rcwBNZ1xqgZ
m5D0YHejQsSLiBmyJHfFONz+GnBB6ecsrVtUaf+XqPhVW7yHEPEjOT408Lssh/NP
k/fg+67gwU8WiZeSLqpClWW9t5uNLGrIaq7aV/ihr1eord52Ll1Aq7pFicF86PZk
XOp1njyDyJyCraTpLBSVyyeYfeIbAzcBlslHbFNcMWe2229rwnDaVOaF0R5YRfRv
e0Tr/pVGNUeBfK+BooJmAmbU20AB5amHS8FvyPVkJIDoX1QHcDLfgxgGrHHYiv65
+OwqGAEw3ma+FQ8Fr6osKEpmBjZ49rOH04G5jI+gm7jgpxUZSvXSZneoAgfFWe3e
V/6id4r7Mm3hxoktAssqLME1js/uC/eBXvwE1TuEPb3rIzX7Gb7s94Va2KmM1+Ta
8/6xKainYwRO4J5Qu/K95HK7G/XY6ofb0w1k8ZpqVqptKTJLUMEG/NeW8gp+KcOB
yvQ/V8kSmDCbkn+gJiQ+MjekdHCLzmkPiMKEqEfrbEnstVnNiXzdCE0XFGt1+sMK
SV7H1wcmu2ChsBd4mBpitU3zjYYSw9oaQgq1R2jX0jxb+QNTGmsaF/z675BGoSIX
yOPbE7pGMF7o3UPp12pjM3ESaeo6kaEQgzjHKHB3P9zWOXH2iX+PgS/E72tHS4Xh
gFKfC+u8rKTiPvlVeXV5RBoDdaY+gqrKkLPVfStTh11YGyL+JPiV6idHB+3+PehT
Lv3Beb0v49PX/sIUnj5vBqXBv6Uo+TqpDfv7a72nyEYvBJEjk4qjD9e5TPueTkKW
x11/baACcLhXqIabI51nmpATfJxX1DJ0hqcr5QFq3T9yKouuFiEmrQo95Dxq6oiV
B93Vg5062wmk3t8pa7JsVXA3u/uN/mgONiQGPKJ4dUjRNCzP/nXe9jn5jH9OEVhA
hbK96PTlPUJF4TuD43d2cTV4U/Ys1XJ12CBEr5s3MsntDTzO7WgBHEhEDN1CNrGk
xoVVpFgmYhbJXeCzPuCITzozyn8/GTHzffPf8znRDhs0qUsnXTjWVt42bisrudTq
SjsppfglHYpHzts0lf47AeUQBS1j0GQbzlBlTRL+CvPz3mAFrCHo8TZnKh+EPi4T
8utpDHYvpjfLYX6eo1m5u7sC+2EZ/6F1h+5PM6wI65rWVSUALbBeN/jk6vaOA0OP
+OBZylBYsL8wvqzMagjF4oUFm/0lr2rqt2I6iItlQeYM2t43QMhK+hNk99q+URkb
5oFh82TO0nXUm2LTlIu4OOPA1xqGzHhpknWHBBqkjZ7vJpOp0TxOglbA7wc2I2Zt
1Bi9SCK0K2pRlVg67iJqipJ4na1sTC3ZtVzSboKHjFklvh4iBP+0g8TbId5K0ZoU
GnuUsqN9tq9UwphmZrhC6SHuPAy4bZNgQncyB8Id3lWp+Dx7gW6QT7BHkie5Mudk
RVGemLD/jCMj2v5RgUaKEwSVQKDk69sGnH1cxRdQPYVsYwarBumbWnv95mjgaWNQ
LjCzYOQh1qmzW97rTKBwB254xdSMP/dPM1eHa4oxfUjZnJkMdMqNTJVp4+eWjc9k
xgNV3hwvBrm84/NrFoAfU2RJ6cfRTQz8VtkowKog36hNH0/Cpvlzyo9wtS7MmJc1
OVQuMDpQMhziJGQeC16l8Noe7U+U0fP1H/vp5remTokfsoxr8mN5RnsY1WqAO703
2KSnftxerdtOXDyrLfDFkul44C0z/tbHsi1x0Pb2apKGZI/tG4bY4nOxCnk+u36k
Ryi4r6mIJv4ZC0G+kLYzGfRUtSQiP4W4SutjcWbov5g9Vo3Eb/5IBok3NK5L3YqI
c4vJWycvf09dOvJWpFYuRVcin7SFMY/JYjihxvS8liS6y8pvdcGG9fpv9JvlVPxl
skPHZDruyMfwbHCVfQVcTUw1uQHyDPTzC34qWf0H0OlgSuEkHaVuBUrfJ6jKDr6M
ouYC8vUfu31gAUtsfFZrODLLcQ1HkIuGALOzd+o8sdNGqK87AE7OP5QTn3UKDDA5
FxOV3s+2PAxrXx7JXrfZGzWnjgeOUyhT70Ho0ABvB0YVV0bkoTKb1Ypy/KY+jVQJ
itIDSG2dLZXpOkcqd3Y3SobgH7XVNNpBEXO6/YMQq4K6YyNPpTLr82RwhzF3+lka
/eOPi42Rvcqrsfrr8i4yJOKkM0AGDBY/rTrqn5wIYan9OQXIKX7yIuumykK7zQUp
RZlASky5mGAAyIf7yktzBJzfFAYOvjO9oQ6kbCyGU3vvtbb2Z+a8xrjY8pCZh1wP
YYFOPexdR8sDErubOOgmXtoUzvGrC6uClJI8qSMq7Bs3yV/4gsuz0THTMRM3OhW+
1LIPepdh+ymPJ8VuX2farapByYyGEMGeTP/JvpoyQP2/aSEU0kkUFLQkcpJ4YWTz
kkMMXDB3nD1obFu67NgG/QKro5un8DYP489CsSzVzzJ7JGAQGKB6u9KrPnA6IFqm
7ewHPD2pHsHu8s4DWK4c7F4xnnHB7ZE/m0+MCMkMUIzl+j6E58LXXBV6BWwmUjk6
YaRyNU+fFUd/CeHRvJjSrKNAmJif8ZrLW2uF3ZjPBdNqO7gCuShJ7ADrZIo+iO+V
Wciy0DuWY+BZN9QFY4BihoewpLxll5dLXWL7ZMNj/fIB2f0NOTORnL1Izx239lpH
lDB1rfB2eRZSFPS6joEuLed9Eg2AUry01rtWZTuIxjsXA+26C2npVj7hsfLp1dlI
z8ilUWQ5CRmFnrDvWT9kB5uSykSRoi3nFj+F5lHdpNejbGA8s/y52Aba6N2znLab
P9icYruehDNw/+ylzm1lXWPHq7EQahgTM8+O/s+OPcZS5R8Bg07UVonkrTewickj
pUB/3eLTf8+TnJFmQSCU/E54bWRUNA0BZlPc2SzesB7to6zgiR4RWw0/vMtwKsey
VgW78d072rEeI/mjb/KoksS2LJ18QsTKmnf+Zua7cuOFFymXM/LK1F4mQX4LO18c
n6n14kNSHWnOSv3DNqcZBgK4+eG7mkV7U/LwozcdpLE3Za2196FaYz+eRy1DmMsF
4f3vxjOxPcO+LvJ4I3WKFZvSG9E4dxd8+AceyKswgSAfWL5+kcxVPIXovL+oENii
PVQkbOW4IRyG4j00G4gWTWtlTNzwAr39gobIwuZGtnsB6rb2oIZmUlTOnMYqlQO9
IMQlrm2cH1LJumYUOpG6lsSAhVPNrdxHXHwi1uxHMaGA2RI0aSWdrsvgRSQuN4EN
U/exOvKyr48UylgookCCFYsmK/XVBJKnyHAdVil8LIkemjobG5rA+ebRmxLcIC0Z
OayikWCfWNocpUCohFUfd7q74rXtax9A9U2LePbZUObtmID9NIDTirN2uSMvkvEw
CqWVMryACs1pwy2XokQ69lRAuFqgBLoNYgVPl/Gs091P37NXLyseym4Yax7KZDEy
/haF7XJvBveoey9j9qq57Z0zcAoWmSsAxTPKrjI8g29EJIvDagt4Y/Ez8azjfoDD
SZbGwVnbcGcS5Z/FRk41Xagq6UeCRfx9ypHjqNiZzdn3ukknDTY+jn/X/T42RXyC
iv7hxaeW+ocaRnYKnwkb/TRTdzFpnmqSI3/BuGyeoRXBx+ZoNPJLctqKkBy056pE
5MbvkLiy2GFTSdoqZIm3aYIOf9xWJSnBlY/7zi+WNgp+JkGG62yDN2aVng/nLZxK
5N4M7RC1/R9scFnLoJciDV8RKsBDgEBPo3uWPYNU2LwGzZtw8Rjjv3KEFfnwhbdQ
qZTTx03JxfJDucrTklOLXRwgTcwmr6WE9YUXrZTxPD1MpnowYyVpYn8eu0Fy6aZp
+DBOzGp24vFQqe2x1raP/f7YVAAKco9k7eBT2ACAv9ohsLXHrQ3roaU2iBlkR4KQ
7K41SA2JlpBg7tVQABcVh2NcBwwEtotpfVVlIAAyyWmZceqgbURgmXYHEOTLpxWe
Ea/6e04UE8v1Hs1atbBzILfJym1SnNLRzE8L1XbQQ9i+efs8xZy9hnvpO/h6o/nH
cVCwBBkRhNx6JHHEgA/0eFovKyycKqVBvD9O3eAIxYiqFl83sIvmHDGMLPKLQzA/
r7kJ7ukXEFyUetieXKo36nPsJrcEt/YRskYPhBIzxxm1SVqw6cPMiCaReK/LBLpI
SXznI1zBnFnA4qthxBfJijE+5mXWbTrl9lZcWldJQVA6GjGsQBrewe4xFshotro7
zBgDiVNVekdAf2cHbgU5Nm7JcICQOrLLmpIH8fI58Y4Y5ykOCXIgH/umOnfs+q/S
6Ax18VnZx2dQ8Q3+X8wKOMg+w+USRz+bdtS0rv3tzQpdpZr7yS78HyN5hPGCWJ37
ERkxeVlIINLfSlxZ/5dTD9WsMjKsq4jud8bi9S5l3Aq6bYHDu4W/ri0L2MwahR9I
PYXgwvkHOdVrxjWdOmr+5dRmAeXe9gfpdDBTvooCwNStC1klflJh51Zqp1v6z3ce
0+DA1Hwnl5bfIEvKeBbO6oWvSclJD8oGadGsExrzhOl40S2V/OCzreWCw/BZ7DDI
JQaoKRHcw1FREY0l0h/lcZT5/MeipjbmBX81lbXi1L1RxUS/xIPKM43AVwbWX1Ea
77ojno5znL1rM0NBKgBXkwmRMcfNwNB/8M+RWSavD+EP1daWXTE10lQrXV1M4+RW
t1Q4AMj+Cd4wAiGEx88F98/JJbNOAT0nPDH+Ty4GDiomKswBlop3gVxdyvm25BOx
Rckp2WonaDb6bji4ynmESnXlR2RycFFmGEO7/J2LZjjW7cHhY78Icr8Z1DpvZzh8
58ZOLgOm1qJfNF8eLbnz8vTf3bQCiD+O2BsuRYznhbfq7L+m6G1dMKjN8BYr/Rp4
iEkukL0ugaNmClbNqMsX5LNWj2TGVdTzCGjW3kIWpcBO4ahWsIs7ENdJGbSB5A/c
Ku659GLKz9fuKLyunza0Yyd0W7gDMrpKrkbNJW+1W6V7xPwkNo/LeGn/IbrbkPw+
hzD1ujgQE9HMJP2/K6noghgnfKpUd1YqMTpUhMAt3lGANAhcP3Is7EfEuUzRtCap
rCKb5gIs9QmGznBaE1sFYo5PRwV+iWEc3LVvO2nJTvBFVCG+Hw65t2lySERziFPC
cgdAp41CmXAgI7VVyl/KqKQVqnUbSdpvwxsoN8eVgb2tGi26PCyDLZaqobrklBY7
9xN1C5CXwOotVch27drMH+fm6WZRIHch1QCnkH2Tsg6Pb+pCqQnrNWqftEai0IsC
ba3yV1x5RPRld0qWAWqgAI/gb+342a2JHGTQm4laRu3DkMHg8WG7/QStaiiS1nZV
ZO5bPgbGQmL04l82m+Aio8MURSR/A6PqGl5qlPOxKbWrS4y3q+R5BjmdYy+I/96Z
QjhY1nXbvOy2dutjqhQEZ8mOZ5gXSox/xEyr+wal6qzx11PiBR3MbMciqPM4YcPI
rsX3hg04Kp5qFeX/Iq7xgFILcBLmpyml5CAXgtlKHY62cfmHcx80FLw6UUXXgumL
vQB2ScEXeJ2Rg7F7YVCvrBjF/g1QcEviK1tGoNRXAoP3nAyZ5ZG9Uc4d9AAdb2zH
bzp/Tbsx3skqFuor/BSeDHf2cclVWqHv2cD9i/Rqwf8RApwPd3AQFQUnJD88qZd6
7iERz+PZsl+5McltZPpe5mMgHzvOfFUmkoL3KvB7SHTxT7Y53WauPSZLU3dRo4d9
BhiDKDIMzLKHbbno/iW58WgJb3kZxFiImcKpsBiNCSpy/8MqoMSVPrh6McsTXMrR
ZgOqpq7bAoYVdGuoFI1OScmS3WpYAXsql4HuuRFj2T4myhj2JBlQrAOh9n4K9qI9
A8xs4DAfFy3BgaBGX3ZXTVpljKtASW4m/sBRgT+y3e/Z2mBxtD5ynKPCCBC+lJpt
jlKyP6eyXLVOam1Fz1k0If/hC9KHWcI+jnwUSD7RX8gQpKa5qgSof7MncImAaL2t
gAwp+CCX19dpK4rBrsj+Jb8q+usSHGUL1DXA45zTUB10TpCdvS3G3Ae03doHe8x3
8gSglXJUJSbhGJPLENU9+vO0WBE0CNBmVlEGwqtCfQWlT9QQ4zFgZkyR6BZIHdT8
EJ37pjWLC+oil38p0VV+Mpik1lA1NZ+8/rm3Zod0rgcKEJljLrlYZGMamdPX0ZRN
iI69UBO14kiXp858q1DnaI69V0kI3Ju1Gz4ZaoAqmZuNIuFFmKO67aOQ/ov4xOdf
9vn1PnghVcFCCWpTNTRnGXaLwBtqhUfBlgx6c6UTcSLJTetFb3VzgHWI+nYK65h6
JTY8QL+j8W5cJjiMQx7EZzWxwbgo97XHDqkzVNDQt9tBcuQbC3VRHfYDcpEfnRvu
6OAk8tUBPRPpHmbmyvyWgTWkg2owyNeytSQNiAPK+3zTh7Hv00UOwOAV3iLs5VU2
FEDr0KvWxr4ZGWio896uR1RXSrJTkEcnCzJAJFv4HxYZnS1lTEKPLNJXfJb+2C/k
MaHmmzGym3/ayCu1aKoiOSxNz2l/HS0IPPtEW7pSur2bEDsh3RsG2ShRsf1R3ppw
sj7V72PVNbVczwPU0i+p4wYCjpkcpx9dZ/QqehrZRKNNlQMAy1OwT23dMM5d31TB
NSI2XkAZ0/WQHChSm+8qWPNtqkaKy0aCr8UoyuxlVD0DOY/rCEJdaCUEoaM2v2Kj
ONSeFesRb6b4eiHrnVe8T8bAleH/kGrx39uMT6gj3F4sfiISPTkKOPqH5qsvYAt6
gQ9iaSXVn8emXpkM6Sb4yVbv/4nfUJ7ylL9E6k5V7lmzJ9pztGpuXaO/anCCw1pp
k7CCHOljPMQbIA5atepxhWZ/fDIQRUIzj0sOTW89xihTkyPqFB4FDzT3Q3CTbmeJ
MVEXNa0EZz3seMbofCQoojjSxphGlj6mXAmd0fXNYxQK3C8KE/AW7czGHYQsxGEY
9W9sTd5UyIGeDfj7FuI+bxZiQC3ojHtRzHOqzaRDU0CD6SuIJRt+l5MLVZCYuZDp
pBRSnOoK4rJ0z51mFsLk8mI+p7oRobCnAW7yzaCn5275vm4IEQbw/Rc73SKrBk8G
LJIQJVKT6Is6pPAimuz/NgtKEISVVl6jviEY7rcQELIjG6yG7LJoZNn0DTBkQdJt
vARd4FbjKXHp/B6r2vHOoZugD+WNUxUlbKiWjjtO6TBYrgIz845PxEuoDDwt9dr1
oMRC1vclmhruQ1MTa5n3LN2xFB70mzhsJYcARiIqyXKm9Un6OqVXYngT8/2boFGY
M7hjL0jRrJamna5yNRmBtnquCxs1DFSo/e+S0SFK6M11hGA5Kc8Mgp/pGNjj5qvS
Hbe5Xgqv51OMXUALJNmroIVUZJAP0zgMTyBwF0txXWUZpRoSdCTVvxaAeAeB8AsG
9m/1QuAyybh5Erv/40kP7k7O2aM/kWX7TZWgsFGo5nnNIaBEsHH1xLsh3Rn8O+LH
Sevr7bjkN512NcKmoND/nn60AnFEgPZSrorV6K7DuuPMu6xKalb+I5QSbcxAWir6
A2n7hHQNTRtkRXoy/AUdu7hPGGxp3k1YvDij0/wHdrXcRHzcYBif1+ieQBwnsGZu
Azysi/U4N4uyy+mc8pvVw2V14QMv+iUd7bV2x4VTJ7xcPamwfTO61bntIk2qBeh+
xF5LfLYYr7G4cjlNI3AoNOeHyMSeCYFsoBf6m4+Y8ZONAjz5QSGanFNhkbuwH/Sy
9DqrfIAx6Lpw3MZ8RVdjtQRCvZGBW7T58xbtebtgr/AAigLBJFx6TJ/FRVKBQmkl
et+5hTJcIXugNR7M7gwLzW1Or2iHsK/+LTKGcvfm29bFN+IQ076MRSSWgKw7Brzr
YwJVrxzmDW4Yad2lxDr3hCqNgMb8yI2sv/5r5btJryE8akWCYmtsre+RGkKLtwmS
jdk4SRQ12i7YWMKf4G2gCDLzoQWRdEm9QVc7Z7Zhiu7htN/rvco6RVttzGWvAGy2
/zT2q+a3+jpTGGvL0+cPWAOWFLDyfvNEE56iTz9eYj/WMLxS/pkHtPSt5t8HPOE8
GGBqY0uu104nyhQ+2dMVlk2c80MQds099cbSWrvyek+FEksL1vMQADkl+kWwNyeM
M/vb6g5E91jtjc5KKFFcyvyvV8u3WRO9zAfA8CgFZ9OlHg/qjRvEh+tPfD8QSt9v
uh+tcq4Eo4I/qdaDkPdtPzWefIjZl1ykDPI7ajAj68aCp3GoggjwNy/tg5tzLpFj
+UcE8wPyg0DaHfRv5q4WSpwnjsWi6Xej7VzWEb8LEcDZFjJs2gmct6ZnhshSwYnU
nHZaEkLwPe6rE/w8DC0/KkEe9cVxuyzZqQNjpcHC0oGqkVzfm+fd/7Y6H/Po7mJd
HfEA2SsYRm0Gk4IvOxrCQTXK9aPtp+RoacYzoCtU/Lt9rQ5lS99ezF9DLX3d8/gn
KsEtGIxUsHlU3DnkLihg2AIN+9l+Tl0nXSDGXtuSUMsmUVd36vzhixuMjVxrdMUL
nnJjkI8isY8bFJ7/ySg/hRswXkPZGoLT5JflKZmr3i/SNyO61wH68lXtS4pxefNe
aQndmrAByCuKN0pVcrtzq/PHK8egcVFr4DzlzhclWgObliMGRNn2EOErINdZ8heH
q2RcHreH6bRoMFDOJHMIxh8fCj3w9VM9HPRkEARFk1IUqRhUokJfjGH6H2+QiN75
szFBGOP71gTjNtZAG5fmuNaoUmuCmRVCuc9tyqrSFQnDLJohwoYZ9n9DtbdFTtBW
xXGLY63CXX/SA7z+a0UfP8XPP8lVTHYOb2huyitMX0tqs11/h+0IFJ3Ov1RZrnHF
1JEEqhUfim5+pp0i9ut6YtMnNLp3w/yHCgOIY3MgmwsepcNeVR5fd/JuK+fQA4OV
sCpi1Jj/bfFGp4TH0jAHM69kVF/4tXWKa3igcTG+bW7+bwovUFHJDEXtOb28ce8e
UwsIAfHvUX+SH3Ez+3pomuP8NfnNHt6IqtfGMX+d1WAbDgyNK+64T2712IzIlZ+K
yv5G4y/naI1yUdwBoWDIApyIlc48RzvNvXfVwFBLPOi2K+FaakgthS5L3dlPwYjT
5EEqffqZy2b8sOLdGXiEjW5+TSemlbDsHkeqauKQKT2SS9Ggu2NYINkYKDr6oWE+
qUd7+OrZdRFYRisrh60WXdBT/7H1kPjNKbfGEvgna/4XWAmvmQ8/b4eLDh5ez/VR
8wi8+dvMafQHPTiPkNt+4wisjNTL0VLubRjGsWe4fDGvOILntihlJiMwq0zuMGll
2ZnRaBmvd4htdBcOu8dWu55CKHZxS3NRqSg7VSvMvQUaMD2LSNJrB7HkRfj4pw2b
ZLR1qmapgHy8jkDFTu7/WXoSzlUsLK3E550eHIJ+FGeVdvXwWxmgCtkH74Yyq4T/
C7w/sjUDkyLeNAWfnxAFkDyiPh4HO40zSiuUZu2oAf1nn8GQYDLG1STjZvL/vnhd
aDTcGiSYF+z6Xh0oXrNvHcSfLPGJH+d4g6Xg4s7POGQbJAiQ2mdspLxmJuxEhqnt
V1gN93wU1oAsJtSMrjFccBzuw2xfPA2RMcunlEhPlXOEJkMFHHkWoIBY5qdIbe9/
FspJPK4fvVHdM2l8BiHRRqqWqoITdu0klPKngcaTWrkIId9TzWD3sJgr8fN3KKKP
CTBksszsMvxoTfB/nArbSqEFEXHy6OfG9MvdRiHA93nAMMWc3r1KmJBA1CSywhae
sWySQw5yh6Y0i5oxp7eM5/DXMdDJEDVIqUIuLH6daHVcSF61scWRhxg7O3udHALJ
ExLABcdAYZlzUHTTW4gV302UWslmMscdzKKqk8s3er3+Qh4Chp1o7gIUwOo+R85M
iYlpZ524oxTJtQfr5An3a6BGXaSDv+UnX0osRyaD79aBrCcwf1MK2j038yfhWguy
ov8l3utE933vs/64jhlaWqtipsPFXzYdqPNSikDn0D/XsCC97qag9hgcQszdkLlK
cgQm34H9Krjbw/CZPipPH63WEL0ERU4Htu/L7F34ANn7r3zdu9qXbalArb+LevBl
LMS/BJyh57YteLFrOXZhjGGXMAXdfw4DmSFC17FEsbkKmzYE6fjDat/2nEcH/p9g
BiLN3y/XjZufRgmN46sHrV/tZAhhhJ1bKeW1uPiRj1YQotMpdVdyXkybeXDlYu5H
KryW1sNcVWDBi3WiuOHDdBU1yoX9K9R9XPHbphnYUzgpDlFkE/2Zc0sWBa9tEUDK
Sf6gU/a5EsD1O6+s6FDUxcC/n5se46cRPmjK9we7y/c8PNIsc3osWrMrdpNBAnoH
807ug/9YPEwlKft6MmHMYew8IF8zWpBXfQwaaKX4HCxTquZr2Qq8PDb2BtI5CrJn
5HEMmrmxM686qHztokjd3exLw5BbFhbwVuBx8P0o5PD4yY9lQbvrrfAwB3XD0ZYp
B/I3e5fHjlcSnT+5Qbf6ohexwutgjSQkXwb8trj2DxnTzdEeJiRxP+XIxK3Nlt2B
QcWnvWaa9L/9j5LJaEzOCGbiYZHeUrtwL2qI37gER71cUxXj0yAGxhEJNR7ZQkTr
rvbkksVNED/hxeJphOpWjnXA+z1KKvMnsEUNI48a35hPHrx6YXOraEltv7gVpkxE
3G0ZY9X/3BF77jzlp1uir4ShwkcYGLWvkInVWWtmbk/gLzjTuzMU8cwpmMe0XkhJ
EnUM79O/d0DP+jphP/MT11A0KgwBfwL5bMd/VuFpECrJ0ugF+ZiJtm/tLikdaG5H
hXBl2rvB5YF43C8aUgp7OOO6VPkw3FlwPlAC/fpZ9KXVbeMALUNdIER91yQycRaj
ckpOUcHHnmgsQ0AOqDWy8RQWf4n/M2OU5q6UWodiG/ubeLJZ6X2xb+BXXr+eXxUN
IqAcdUVreGyfls4BnG2+kF4MHAaXErfsJVfpDvb/RyPK4tweCdbAcqg+9TGKwLtR
thLpkenKRHeh8PAa7ErUxdi+mfXY8UfvYTUK9o599ooW/rEzixjqX0d4U4eSP/IC
DMjJcCYsFYFbwh30tSwlfVYxkTQAPdt13R4blq5F8wIARQuADS/tFHyYfFv+nPfg
5Q9JwKYUWjdZizkIaszhEUXOSM1ME7L0Q4JJ/HaIMfyhcMInajeQ1cVj7fdEkKtF
Niie7nfAtFpLMUkzX4rhWDYoNFxWxCnwEXatFoE0eJdH9OtYvSjIzfFhvG7i4DOz
hHH81gpJCIB6S+dMMs+BHjNUevD5aRcaWr48jEigh3wWlwk/h1rP0EZnwjhg/BA1
z/0A8Vi1hby8b4oTsT6MCVPnSrapOfXmq+RJx0HdFOwUqk/auMwHg3C0ugeta0+y
KrxYOOH70GwMovyh85U8fKtqs398E4KC/gs/G+CooYViSpAIQ6X2ysPLCzeidOD/
/+RN1rNtR/Pak32x5tOebcyMqRiNKW59jZwciypg9CHxy79uxy9bRfyaAoGFCuIX
B+cOVVzSaPiO8Tge7OskfVrokrNJnUPqCLi7tzmQ282Yhaj07gdY/vq2i2ULxg23
D4w07ScOIL7BZsnNYZnAmKb/+94BHUdias46JQ6yzzr7A3P9bp1gJb+R70hBhDfc
3AOqxQatI3Pyc+7xACstLx8rYLcX9Uv4TAivL3JdM2J7e8YYMSuB9hwd2WLUkUgd
RNu0zGZxz3OPs0FGBeijqaf/jJ6XYjixE29jHjZPl4HVlUn0JPbkKX7yL7RLWoZw
0YwaKsDKHO7meubyl+QFMAK+aNiHKsSTqMCRouLajoevwpy0YNI1bQatDBV59/NE
m+EUKnZP6PJN+fpnPlwTWkyMw72+aDAkep4Rp2VV8HOi6cE8BTm3aFJNwxbH9uer
YN+SI8oeaABQr7mFu+qfMGRKIfJCeCxc0SjH+T/4p+f/znTAREVcOYnb/1RDREpj
DPVaNI9/td7Ul7CYhRnQNqqTGibpHamx+Rwl5046/drHrS091gDe9jY+kwRhYC0U
pPm+xO92k4+UM5dVIMEs0xvA92PMZ70n99aEFZXbckG5jva2f6DR3uGKvPufdPCk
7N2Ete+d9dTj0sNvrGGf8d4TRTnpM2eG1yqObV+a1LGkHNjEWy0BpXqwonAhLa+M
yHZ3huQpECkuZo8NlSaG8uNhzJrm4bK/3/6h0Gvg4dZVlzPNHH/qzySuqC9zqOEb
QRoxLY/dJ9SE2PLtCe4gXuw4aVxvjOIAoV5TJplaAjj49KFSlTMq18YbY2TpExMZ
eoOLrshlM1FFun/jpTwxvmlWu2K0Ddqs3MuDOtYrTbTFEUF4DOY8GVD6iQA2J5y3
XQat+C9Ha2n0RMlfUn94nXD+jmiecpHuYlFtRT0KydNPrCjrMmTdZ+Y1IIsDVrsh
k3cHekVsly4ElfG3XBaL64UqW8UtIIcYVbM+auVuzBK029Z6lhaHlNhyX30ke+m/
Tifi7BV+KLAnOEHt6ocXtFa360RU2OPGWBNpM5EAg+WzCkhktJ3e13sSS86KTQbL
cV9TbClR71y2sgNCt+14HwN86IcRrgw7ngCq1Sz/cehXOwJjvTW/KAdfSkJoyo8z
6BTCuDmH0s6G1IJXX12rU9OHO4F1CHSdRlZrqne1kTKhPkfSY8Z67VihNZQQ7q09
1nPbIPD0VA0NNoABlDOdsmkjDTFGE2IBWlgFBaDl7Obcw2K+BrVDbKpJZ1Ac7w1z
IFIcF3M+O9OZ6848p6H6/ugAfemrOIVc0B7juYScJjuCqUcgiTT3JKKpkoYI/TS4
tmZxicxcltZkPR3bIvnXgSH6VlHD7StnGokg7LTypHVbyc+d03knRpdsVLGaK1qJ
eJxiHeERULhhRZuk8TWVYIgCKqHUsHoNkyc6JVJhzOgaOIUonU1+dfMwz5L7paMe
jZxuGbgLuSM2eE6jWBTWvbDygo+ajcxvO7hfeKAn4btHONnpwj04PVTBlXq82Rhv
C42GyJKIqtHoVnexFwMRYLtQQeO2MkM/lqNrS/LMveDNIdOpoUAw0khbixa2f4BZ
FVV3b+hveE+xLr8yC2jzAsN1JGq7SK7DMlASlL2qn94gBAt1lUTcJMx5wStfbWc3
Ys9u7ZaL6+qevpXIMoxX+UwduaALVlK0aU+HiG02VQwLaq5iCE3Af6RMbQZNAmAZ
H1KpSUICITATL+S5/3EpcoIKyROqTgNAAW+8GDafazNZ0fYzoz3aozXJMelFhShD
KL3Zesqa1lARbTABjwPiVFMD858KapUGNcdhhVUIkgI4fNk0RNQIxGRz/i2eqRwS
PquKjEhxhdH0ORvR4NnUrBTN5D4xaGRQbthwMNwLAIGfCVcJiidHV2+2qG5OggQf
LGhJ8CZv4CvrJnOLRL2kux2pSiKiPfQw6LOldIa0kdLob8vgIqfBgfHn9h5Nsfgu
WAgwpLQTiD3dcwBIZqbLm/oLBcJqSu8PhSw3Ql9rMSc1qF38G9PwpgmMBna4+WPT
3DyGpVd8dH9RDpFrg2zG8UEa9j+mfjR/AN028mV+y1ae8cG18NrjjpJ3mhVEcuEg
nucitd+Gl4H6ppU9rtE/9KBTsC2ORtesnb97GBzh8bUM69GG+Hi+pg+CnG/9EeMn
7MwE4CFq3xBpp8HxseCnTTepQnJlHHdzTvaPTfCc89xSBL9LNfJAGRTry1FCHa1e
2f8WFBDusgmznR9hzgslQSlP7le0NIQQQ0ex6aVwOOm6j+CUUri+QITXjjYuB8J7
LVm0ig1BOW8Sf9xM+EqxJwp46u96xH8IKb1qsf9lDeG4BRuaCVUynvSnrMF2TCOU
OCB/JNvxhE0+2HF6k8lbMvW+YHdQTCvhRFmRCy7N0ReodXEZb88hC/gk/QYBZ5f1
mnlAv+tPTZY4A1DdfpUhiD242HrRAvKOQF/2/g2oV4FTvpFQiwfxWp7q7VLyzrm9
IrFxDsuhg8IT4WtKQ4MyJawaDxJcOOSOp1Orkmr0kRDDDVcREYmyv1b3Y+LzErzF
yoXqh+1G6+M5dt749p5CUBen7AA5TgUABfmDcvRxcmyX72d9ySKvNK3/ahsQ9n1F
tzTOWWO8Aj1ZHUpEXVSP1W3MUFreA3Tmmlej0Sb27WPaZDEaZXSeF1/3p0ij7EhT
/iHw3VSX+ofxZ8k3T/J/s0aVIYlUpqINN2zAkN2FcnJ+08Sf6Wyxiw5PnACTmANu
StEKnj80T2zJAUMm+Yr3NlChdZA4/ZuqhoMggermDhYkQjP+DqFK8G5NAmavrdLs
RiA29EwFpNg1MPlTe5NOi9QtqEXgOVPd2eXXYz5DMlLMEwseYx1KGBAuin4Sp4UN
FD2F0QE18nXpa7Ty8dnzuiAvjU9wxaQSgGNIlDXKC1qp+Z2nQWH3ha2HXBGo7AAM
F0i+vCmJ/YVmr/9BCRAzqfmfD1jdsYf7ef/QCseGjIlrsRhSv2FPScB5gQGTkIlX
gwKwQBzOD/xt3gqGCvTEoCFgIAyOxgrAE1fECmM+tpQ68ywI+Bqu/n8VWCqRhTk4
cUSE9ajYmk8q4onajVYmCk6Zi/oKR1OkR40seZgv5z0jKBFIXLOZJ2LuJ3VQdo7E
D59wqmzGTLBLnZ3wN/TjOAly4vIiF8qYOIJcpPgEiVXneMYbKnoFfCUR2NlkB8MI
/RQHadE0tnYF1Cy0lzdLODKZ12wVdSdBhO7h+N0vL8UxW8xj1Aj9iWEcQR6yATgJ
5pDKa4K0lJx893EZCXfQZUDzWYPHAgs47wwEgYly6a+YKrtvChsLU14SViqATtHU
FuYbi88CvCIIH3ZT7lliUklF81T9Q7aWJYkRKnWguCHWGfBl1rruiHyyhHZyfWJf
crzEpxS574f9l3hiv8/N4NQERPagEjPyfkqgaVqEoDpEuW6dnQY+J8CIePV7Y9Gw
zlIw3s4Jci61kTdpH9muCFL5+57nOkJ5rXttyQBhE8jw0FleAJgvJ1JTopuAQifs
oeD5nH1ofaczYWPyGRPN3w2fpcRKTQKQtZzygRvAyVdQbG8OPd8XEhs9pCX+0mt5
sQu+B965NsA2RjFEAEOWyJ/qxJGogh8vDNnXStSTdKUw4eapzoSdTcCAGozboTiW
Ef6BqKPThjU1zzICfzVhta/2rYAm3JB6F8kTvStNYrS7bKnUwKKtzZk/0u3IMVZR
jzOWTPkw69RdaZO49A8WTsoEcixqS2FkJw1lC2GdnOlT0HXnCX4J37Fke5kqNCLs
cohqCc51JZCwZOt1/Ow6uXnewEhTH1yxqFyra7Ph9CGnrPa8Yl6NaRGQ7hQJ5S2D
a2cATnR3YTpaxiGvlySYq0Dje50wsGpeYJ8G09Xr0irNru0N++yGyQIh6+zKOpRE
Wzx2zHsqRLka0e+gJfwSUqY8Yz85llfuVJGa1YKX9aGIDUh6kXssayEBanEDiD8U
aPsHiMiX9L0CXkHJ7e47O4gbbcGnGBo9BG4Mx3/WXRU0Vat0iXBx+Xj1fywzCr79
Ti9DVgCiQwl38DTF7m3BfAbaS7c1HMjI6MU8dYnUChSKqyz8ShwepxwUwqhhuV33
ugv2SNmIuuIFGvePPhrVG0Uo8xMFAfGCyEQsmLGsjPSeXlMAzMGr6lcjnyxSOBkV
P9GBhg+OH5qW36gzc9CO/NuMPm80EK4sNncoOTZMsOXj05egsEMC/VJOwo2rKlTT
00BXo5eOvcUjKdFW0XNvFpCtbmHpoFVbl4Fy340QIY7YNVU8xhhPMivb1TdXkrNW
zzuAKcfys1SeRXfBqYRKzKgDLyieD3Y0MUi3/dL2X1Ys175UW89C9acOdzoMQeAq
ZE3zGCh5/6JNQUktoRzExgBNr2Q6YnGKfVPMZlB/iDch2w2s4yZKCg2nxe/kErEq
S/AckMvPam8Qx906H58yvslcRJGY5v6WFJnjf7XM/dSLx/fbgbXeID/cORyzRQeG
w1sRVO3Otw874Mju6Bg5fFnxgcoD1yjSjEL3DnAoQkorAGxRbxIpdOtAhlyPXJV3
gvHm1lqu8t42ME/aMiqHJCn8fsQ8R+DxCwpU3bnDo8G5STMLG2FzAq129gleLBcr
OP9Yq+HR1ey6mPg3HL7Sjj+YjtSjA4eY6tbOWPKbuHGwcyK8kG6Rm9RNYVHFewUA
P3dbUtpOlRCoYiM23zQjWLVCGs2pMUeb9XlJgRshMI147pkdjmMtV7jKxUfs5HJh
NFX4SnjHvt+RPK46ppCBSskQezLltRcF5As0eKfhQcQZO03WGiSL/sUnrehe0QZk
WXMhEfEGRayk9t/2pc0kL/928ZO4jJfPOVvBTVjzamAkIhoebavLuqF3pBPs2xfW
X2BhU7U0hDQOSiAcAyB4ryTty1S1TKTWlXNZBJRe0E2tt+YyGRoODxpF6HiZsQUh
UUlqN5u3sIuo/i+iK0v/w60MRDOgXVIcBBko1K0RoeB3Amz62BlAkS5NBs22RJE9
ZipHOijfgsT9QQoo84L8UT8JTiuNopNuSsYNs+MGok3Ipb3kBCx/t4g48AaP1Adr
e18t5MY1SpKRhplxlK7GycDkIV6JwI0e4VBT+1iYdOuISg2Rb8gEWcCZ1SSG79Aa
i7zXqlzhaG8y4vCMW00qlw2f8reEGCQN1Nt/gkqWAwks49XoCTq8NJn0cWgaVmed
B58NHAcG+leb+Muk8D7qEil5hTo2cx9NfJ6p4C7QMilS/1But5fgBZwpFz7rWor6
k/WHUcJMWM/dxtpor5PFmDvbWJu4ZmcWfjOdKxBnjfmSzfd5lyL1Soa4Pv2cr/N7
U1kogT+fzjvGwP7hWBW2qrwaH7jh3uMZrAvedJxVexmCZIpx07K0EIVDG8x25CT4
xU9AoRiQDhn5iuGm+CO4ylzOTBDBMglXmp4KJSgJUGomSB+x7EQCeCFx52bZLEx9
EDK5sujR2sawg8e9EJPYDrlnwsDseX6oCIbu8f7+HSyDgIWCnRY3+BN6yo9f8s2/
Kk63geQDOKIITYjeuCPQE5pCBj1hGLmQcf02MtiKfn8pvwy43OMmXdW/IHOnncbQ
8Vl64CBKlAKm1g4rJsmS6WJpCNCmYkQZEiPt6OrILQ/pfibm3ICFLoNo2QArZuDE
hR97q+qjcmJQ7cNfNi7RChSWQ7amXAXLxV+/5p/u2B4oO639wLZHJw5U6Xb4aWL6
BRTnEsWgvosHZJLRJGkBP6yQ3eg8ngqFwVYfKRrhZ9LlqKiwTy+DYCPE0/OeJ+1T
XAAi3JjgGXWIoDq5V8m2X5VxkFzlp0yyTx4Iqy8AU5HMygHy4Zw9ExurmRmhZfTF
dqUvqGK7K7jA5Tkf/9OsvI3vmQ/h8QpE/H+NnLVPWh41DSJdbYPRCtMoz43q9ebE
0SjVRFHweE56T9hmINQahhFUKS96kOYWak+qbjmtk7Z+w2JoA4xzZ8GIUTBqkDNU
8anH6lurMjNYTWvhcC8r5alA6pKmYG0tiyaMcayS5luOntWSEZFnSCk9lF4MHqQp
Tr9QAT1ygYSMMF0OhMHFs98DIQhdXBsDYIvkqEpudJbYnYlKLh+WjoMo9nCh9usK
qAOpNbg7MtWH4LB7EoBvVyOHhv82cLOZBXu5uE+4XHDZBYJ4QBOIuWaKVjCmQBaB
bsfJLs/Yry5j7kL5PiCdAgY6G4U4J5GK+wxR6AIio6ktpr44T3Io/0fsr31/X03b
nnsDlbHNFUgo/gD4QuEBZIOJEIw6vA04GFmwFXQwrWlbfiGFXaEXdkOVJgnNYLfF
LOJeYN4ZmDV4kfAvBqe8Fh+1O53Y7tDZlHniGKM8ZnA6ySx9NWdK6bDNriqLPyoN
WmYmlBV08MGJuyzMP7eEUBqt9yi/bpLI+5m1Vqk4atKYHqthfTkoynyoXdeELaB1
hf18q/Fnukqf6eeTlbYhfYjxlIc1f/aiHjIqEv+uHkZLQO5LlSTDGrVdVswYzZyx
gn2NEUAHUqP1AcQARJ1y7p2g2MtDLgmC6epJQQxTPQBmS9hReZtWifKjThzdGZmb
vsSDnzpnnoBd85gVLq95moalrXXSOvY0MgHOYiiXdTGLw6YM75v8qg55pMSMCuMY
Ea63ANd3Ojv7CqSxLjHLi2G3xX+U2h97ubJTknY6bUbSM4A3986fAUCKghgxCBE9
f+A0q41a/qAIEpKF/GAwerJIl7y8Opsjs/7xhkx/BS0bSo7bHIi5mPCguw+A93+w
3/EqRzc2M1KnGe4W/iib2nP/ScvD5Vb64g61tiSyN3Sgkb86klSLXBu0S/M3/ZIA
+otHhwX2ckp1SpLfQuqAfT24vNv2atMy5RvMaq8m+kwr0Hsm/Swg9VQwoljJJHFQ
438mlLDLSmC2U7buNieNvoX/nfH7zMXldEGmnT3ln+JZcp9P19rx0JsCuDnsbIIt
K6ofFKSyO3RgM+lUBcMkjW24yJfloKu6VEqls8zsv4oR+btOjFj+qS05ZAiIOPp7
ZxErJX5tTHcWS0KiDuI5FpCnr7PbIw+ke4PvIuo3b/2RkoGZ2s/i8OyRAHnH4b1l
Qx2Gsj2lg698tGMkMmswixn/psg1CwK8Rt+QWkDqM0J+64FDIplPbDLJZlwQACy9
jrT5yY5W4mv2Rrh5r9bSBdkT6Lz9I3HG+Rp8nYt0P7PiwQMJcXp9xzzbZWBzNUjr
x1Fhi8z2JintW3uJirtELrJCbpyJT/dXvcrVk8nVGCfd9mUEbDdPJQub6wZrYLyf
WYPGn1m5oLpHpHaqt6b73vtrNxTfz1h3zxhvwxBxMzUcz1iP2S0hwYvjbeFGmLtC
+IG8ajg8muCtiGnPV2D4eWxoTek4NlIognFCKAF3RuRh2GppW5cWwuPDWcwZgP4E
d3kFjtNq/OH56Ql6hhXPC7Yt7S09vlMikwDXBdb9o81YRyUHuRm9EgCJrap9epG5
UPckHGxoWHrJtwcr4wkFOJrOy9/HgODiTGO1yKS6P64RKm2VaSwy/ML3UNf5x+mw
caEG91Ht/mznDcpeSIltmWZ9ZXuHqE74J1x6VKeyxWX70j5zBdM4Mqg/D5rNdQnR
oa0/Ux+fx7F0mVmoqwfRC2wCeoGCMZ5QIS3DPjO3pchHqo2WCz9tTPBr0jztfObw
+lUhFAoRP9GSZpgfMGnr8t92oWddjDMA8DRRsrgPyRgpfxcEuZ4gdQbqPrBMGJOJ
XQv7LAG3BOoviPCcamOFpmNlnkiVz9WNoOdlWkeYvZtK2bsVgScrMEpdoGoQfC1S
prVinQglr3y6GQKVFlfgPhtAr/ifXBEZFTjTHOtno4hnisQ049LK7FoKQ00V20XT
L58ilp9pveplC1+c85abXp/AmIVIaFxiSeM8W5tucRJHtzFUZ4zcOwP2qL/ESAsn
nBSnWhbdxzdMSdGoXW5kuAJZcJUd1Zi9873oWxoMQBq9VAY9xLYzfq91bDNVLYBc
ulqjXoCNajquYqJ9A+MnSWvDREHQkMq3UXhufymn/1LnXZlVkznEv7ste2MLz0UA
Bz3S7oQi2N3HHuoxiPkQHn1PT5sIRfSQ5VFQeiTdjFwlkvCvVSX917ztnKiSyLAx
7w+H9RsMXZKQ6PhHHPbh/Dx4QpayiUVazvt4CmgRQMCKJxgF2Nfl0htB11Ca2XL3
93fKXG4I+17WfYHaaNfQbnIql0dBqGvZ5VCKpFXJCPrdx4Yjby7GKSbvgnZkzISo
MYWPMAfCg2N/AsQfStWdgbr1+rM72muaNwfF74l0hz6tT3SlHvnku95Kx+0qFGHM
cYY5QudWxMaRG/tc0cjiwD7k3HeOOcARI45DHzuJ+IjbocF8ZAv8xo285sRKrie4
mj17jND51Egnyi7UYDK1EXD3xTXMKLH1i6olyNkrY9MNlyOdqlPGXEsXG7bHWVgE
l4ooGgEUqE7xjH5S3UdksB3IRUami07fckj7c6nuV6H3zmRqaqBZ1knXOprNi6JU
Rg7wJsHmIipI7E9i0K6E+fgscr7I5yP0r8ZrcK9/cAhh8x0+eY411jwEje3g8b87
B5HY+/EuiBlYqoZNGE80myrttbXVUKBPAgyu8KJ5gH61HSwUkfrzAyGwSs9hau+d
hlLyWtgfgNJ//D2rVuuaYPidY93gehTBWTL7YoWPS7lBn848VqgSioHsNKVMKSxW
VpxlyjawYK2WdlA5DhS0dhJiSiOiynEdDi/ZtUgn+ToCdDYFQPRDewTBNmwFs97V
taY1nSYL9Kes4PEMBua+Qs+1TmfcfxOFyfkgLhDCI6cSs+9jYtI5u24Q9gwhHTlx
2HwTE4TXCPGt+fiLVLKiJlrjr5RESfmyuHFjXWoblX9JxqJaX6rgNimGKBNTeXtb
L1fmAdwusTHfjotDKAwKMTyIB80LhDWl8MxiUPE3iHRpTz0bij5l9V8f6cRI8aoK
9Z0ioOxLUDHcwatFW9ock89z/gxaJElt8p/Uj/1R+XivK6jxGncYEgN0yCx4E49f
9AGzOOh5YOX5zWxtfHJ3RU6W24tnJjWVs23dVDxVRb5gQkDEBowsWE0dnEQfuW5z
+1+VNNdq1/DXHlU6Ec3a3HfevNWG/XnUxQWXNAjUHhr/p+X7tljQUqq3s6NL13Iu
QUIxOrtaWWiSPZlhtLoi+c8B0tPjp7si1Ey6Yyz4MHeziIld31XEL6dQQtR9CZI7
/XCIrYOEspTkVIimbVCE9Y5gr/djr8781ahKAAoeBV4TG7yS7l+DcBHEO3/KoOuL
vwy9d2AE6aAr01mvfFcmDbhrQK7plEOT7jb2YLFlNd42ud3EFeevixeHwJi9Ebra
5VRXvKXl9CqPCh2POUAGEphzhHGOB0zVR1n2BmakkdKdjDt2eedjdBJxcODz1NMy
oOurvUcRjbyC4WqGxmFDWb5zQOVlQCTJqaxsMH7p4pJ8BQB4TCTO511omLCSw11L
eTn8ljI0LyHLJqSYzp/3FPim6b2/oz4ffeK7OGqCaaw5RQAyCi+zKrw+N4Tqb5fy
2MlQw8HWF6EuOVXqSmP8qURsRVsO3Y2LOqsV8el7jQcplNNPuT2MB2ryCJCDT8Tx
6fXUWsEnrzwJTAS3bUi5xn4v2Qhp9MaXtnfZecb5qKWFS0TcEPmyJ/FKJryT9FAK
gfxIfgyOzAHQM/I+pPmnccC8lB+R7UWVFHdC0H4RcNgjQ4+7UlSBDCB2lvmzhMy0
vYZR99OEIJYkZPYF8fbwx/8BGtMsiWk7PdQkb9zS2AK1+FVHGnLzdVJigXUb86NR
Tti3hkk6eWfMnHB6rgovPTgLZTgwOtzSiLdu9Rr0i3uxsx1RR+L1N3ljCVd4TGmy
XfGA8pA/GGMADI0ETjsCZqTdCV/62IVXgxdwQe8mBgJYpksoPc9j7vAtYiS4hrtP
NfTaDZx74Op0ZhMa+qb/ABQZ4eAWPqSglAF847CkZ05jEo/bpoRpmB2VWiD3C3Nw
LhADHaZvamk1hbAxEa7aOlq6EaA+vo9KBC8kca524fd1sfJndatM5pTna4UqY9G0
2ptFsBtVkoWHWrIcBYjHZH35J0jDAqzrQe+l7Xokex7P90w0xeskK/V7VGQSPSNx
yif1wQ+0ddW8vvW5FBit7O/hWgJvakwtZkLe+2SyCbBHTATIyoVxTePw1Y3ML2lU
5diS5mWgR2/UEM9f7CN5S29esx0xbx973tAPclKocqwp4AHWrH8/TQPofY1zeKPJ
hKXIEPGY+58Dl7zpr40FtybjiEBWOmDMjAMq/cylpEdtsAYvGvACp7NCZ80SVpoh
5yOiC2yuMTwCdFwlonmaEuNN+KBhqTdHjHLFdAs56S3h5Z1r95sn6K5z2S1w4K+G
s73EEh478L1L4Cyd8YpoNRtOkNr2/GxAZv9JIfXnsjJYr/o6JRyhbiUbvtv+TbTz
Y/ksZXvGgJmmZpMK+c5MO74KD81tCkYlsbQZDGHXo8EAFRJkqjLVJOiBYzqnBIUs
iuROZZRjijG/Aznx0tpVNatP26AMcB5gIYuFM0qBNcUS3WJ+JYuzRrcO/vt1mv6j
t6qheSRghTHx9w7sPCQVIlbOzXjgD9B7BWBI4ZBX9Xn1LnRU1L/1hR37BYrC3OsM
tpNb+sGdWMAYjhu6WbqIpmVmk6Zzdj0BewAT0HTjXyNBSFvnGsUU901AYqB5RZxI
Ua3Y5Ew8o9UDaFuu12OIh9I8Ij+BL02q7mfZGDi8tfkKdJSWNnsWXMkqQldZnhjD
HOQczPVBMpIEF8Pv4R7URb5LdReVP8Xbhr9iVOuubXLaGDHVENZrzqMVaFfqbdlf
f8mAHP7H6gzj6emPZjd9bNQ5/pIMtsQE8RPEiB1swSt7pEJgq/b1UnZ8R1e0kuMp
BtEWwoinOMxItU4qfEMfWAHNNFMaAj5vI5TQSIhvKNJ33VOrIBx47PGFs7XqduE1
BvOSUBKALxGkjk8+BsFhn9+i14ebCl8qkDJvkPv2F8zfrTC62Bnb8FmyCXoWXeRc
+xbR1D3c7QEHy/2QlQAErsmD/ijacFqi3URwG5PFT/VLircTLsok+wkJqOQ5SjBG
9neCTZkVH5XIZFP5kM6yI8zvv6LibLvAVHE9S2hqzkqyWQvTzP88WVntVFovR7dn
g6vqkLiE7TzLhFghbP0bjA3HOrY9POfmLIrp8Sr8iBTC7amGXYegVpz/z4LY14N2
Ejs1rwdayvcL4hykOY9dWqGGcg2UtuXxUC3I7mtBaQx143saPROw45gPhmRpfZ8P
ek1etnEedsw3YPOTy8p8Zb60yPBf6kHcXmbP3OMjp+c1F8tr3kY9aN36iWIjNNHl
fGzkS60dNPN8j8R5Q/H8o+yk9MQablHh4AiZkXLt1KAzzvydMNRvRgsSeXm7GJyd
haB0spTZeOFO0IzYAIO9e/k/XCHRPnORYzyUEGvxlKLnRnBlZC9AGmZ7KH8Ka7fj
KEl+GhgBTSTTzb1wRxXRefuNIvoTRsricbCMuEEGjsjFO3Ac1u6MVFX2nqD9Psqz
Q47z6f9bXW/kSdPJGA7pQAG93Y8qkbvIJLjt0RL4JceTkNPHLYi9Jm//EHi6mRTy
PFKWPZ3MvqEvyt9p0xhe+11TWUzC1fb5cUM2kUDmLEUDJsySNvuAgp2uCt5AsgVq
yLp7iF1RsbtEV6C+NKLlD0uSPgTKXVY2IfxLxNXfzXaWpjohpGYSR+VJS28AFiHY
rYUAG57NbnE9Hjc5cDisGprku4MX2NU9KpjLSt3c1M4XLSYTDCbmZ/jYGrn/0qmn
vagk9wSCnncocwe1qqXIKhO3nmWszhlzKvJGIaBme4e31lY/Evsmfyn4J1ikVNmv
8JePwYdHg7qEiYUXY842r6NBnt3g00zqPuH1s6Jw5OfCkTDb5qPdrdYlxb9q7+YL
G8yEWfHOxiva0vbHssV7k/U1FeQrL2a8rDkFOZubKyZpt+rMwR/YYpbR/bY8Y2zr
DOM0pr75BhKDgJSXvu1DQL8ljltanVrDL7Lm/t413TgKC831JsxFJL2bDX38Td+w
MqIGAbmP0CQXze0VEpwdmZGSkpIzJP12MUeC2H1PGErcwXWuyC/dGHZTAm+HVfH+
2j3RbMnYwBh9yak2CvIJOAb6+aGUz2By2a2TPNkzBPWcofcdTOIt3Sl73nbSMVi/
yrXbwBlg73yVX+R4+kCF+b1Cl0vpIUGJTlhXWh98rTBJSTBjTV8F5699oildyHzi
zyJ56EaAYInUcqDCkm2z7VMc5SAVs6jKNy/Ned3fPNYOufWNjYK7LGZY/Yoy8GZO
SQyUJBJ47ua+SMZkgBwzRMorXa04SK0vzh/v9vkKC3Tsz6LuhenkBsC0pm8ewHuW
EgckCNvcJ+TDcDCqHhTGkSPkljeXn6/11Jc1HUbxxo++ESvQyeYPTfMKptfSwDOs
AtRJ0UGLouUUUQeljjCGoS0PJzJodQUxNErB6GL6eGESk/p4E0O5llWnYDsRF69H
qzZgCHPSEQFZ9GnHvVJmSOph2/P73VmWkQ79Mg3ryR7A+zwUmnPFSg4khJMBte2t
yKMo09qoluuv+gMOUA7XsiU81hey6aYvdV1UFNOFbGtcBpHY5RocX+dqB2yWMdHq
Jy23O8gm4CS3Ic+Jd9OJnWGRGXrP4WmjwwN7P0KMn5K2oucZXeHiY6jOjVrOFXi7
9VP+/J0fqij6U3vICTUoGkXOh+f3zGhweP1B0+OV4VD9lGZbzkKPzPv3GzKsBQ+n
ZT5Nqiwu/gUq8wKD8+bVsn5iDhgaEvt4vc5wrPdS72RDlEaOZiq1vF+JvBxESlV0
BO3SuRzgTq3n0X01AIH5xPmDm1R4BcfzIK6/6qdKTubXhctjPY2hpnuTrpivdgrZ
NXq2xM7bL2bbhUUf63b8PgQbSo0vTjpO9oLErNJ5LKG+hydnM8djB+MiSB12P/om
+CLVWnjxXhAPB1nNsOjC5lmwoPwtV/yiR5CBjncjrEvYOVV+5x2lPNuagNw32Vzp
NiI1jJxY1CMaB4CIfYl/YwFXCfl1Nk4OZfc5r9P2EA4AhPr8WBNIQA1znidcYhrM
tOf13Yucm1Cz6TBX7CG164p+i9OfNOsi+BvD/1j5plDdWKbjtx+GpxyxwS/Afn8j
Qopz2TTfsMK1azRLgUt27MiXE9sBI0qy9VivxbaETBaF4zjT3aX+o1mh7rQdla3O
yx4sMCV0RhyQQp9a8KXp36JFIx0J1rV3ZZNOXkh36L9whvdLmYAiu7TIaJcUkxdo
hOZGZEeLKDyIKU8VvNh7WSuylILXU5UdxzDPS8+CRV9irP0JIoA8b5PiPbEn1q3A
LIzK/XHaJOepYSrSolkTRR9e1EcovQ9t5Klw25LgcA3L1XiVtqopjhAcKMgU/o8d
3Ctlv24BoUfpgM0evmw7ZAeeQ/Ln91to6dYycbx8jNqJgalyJiYrduxDbX3+DUnW
y+/ymtVkZ/gHSMKCEofj174t/+thWnKOF8NxB0PPIgz7fNeFuB7Ft8vAO8KXOZJL
fggMsAJj5zbh2pcGGZlPjkvUEjkeTNg3HIhUyvyRUtucUoVPa2Sy8Iq3/k1dlpW4
yOpmH/uE8Yx/Adi7gPEyctL6yn3eQs41jJosuu+bGIR4yxCcnot0vOcdGzCITioa
yYvUlyp4RZODHG+g7TB8i5YwqDjxszXV7f7JHzmqIJuWlMAH2kZ8mSM88iRNVlYY
ZAkf6eD6xF+a04oVCxc0FHl6VTwWxK8vvldFkUZIDiwK12LJifxYa3G/R/k8jgor
kYalQ8KDrt4y4IEFSnX9+H4CbdTGJitB0T7yNVmUqV5yvVD1KCHXXrxB27uC+7fc
twNUyXJ5FKrv5O0frX/b4RMRpMb7RomNbKJQiY5cunIJyPjtSgVV0GyiafUMTeth
hNvOGj2YLwDIIxOX/3LuD0Pb6t98d0iNTiyppqv6r/JkjFqXu07t8L0sRi4uZPN5
tnGI4atQTqIyjV8Qwk7xOcpm/YgwwzT0MRyfA0zN0u3K1NFUXAqoxlRQbc3ncW3K
LyOnrYv2atoOxiRcdOZuAtwWuVdSygCPZX6fmGb9wN6wNGCA0kHFWXaA09aK+rYJ
D/IBpEAfmcv0QvbV1NdE76pBLhckqS7LqrBR3HF0WEGAVSlQBhI88xy5SAg/Gaul
AwkqqAwkWYwQ4sQ6/g+AzLYD6xkpjdhcZ9IK3GEBAJ0fF8+949zSG9cRuEOYL6m5
ayBwrbJ1Ff+QKvLyysKY6lv051JZkRPI2XCBEJCitMXnZi3iGb9IJFRUdNNGlKWo
0aEAWHmiiQLsaw9PupH99xsIbOt7vUecP4iEEnHQaIxXI9bIbv/v2I3wo5AFiqTZ
NI55+ABVQFYm2aj3obXA1PcP2c8zQiipL9xyquIVMeOwu2ajQ7KA4rgMr6RCJ37W
LVvwae7pQGVLZbE3kbt76z6bP2fggZ37zWrd+8Jqwjl78DTx7ibRY7dcJaaxwQc9
mIzGuadErjndSB9peTdQicZNe+TqqJsL4EQqPNjFN9n1Z+/0UwRgjaIoqa4fs/dT
7HMHh96uBTgFkYRfewjaKTz4+LZkau+enC/hLuap1JssLViZaF4h/bvDObiCPRos
bbu0l/6sR3w/MYS9wqgoxpGQ5YbeHiFT5LfiiDll4TpfxKZNg4+dd9DdLDPXRoDJ
+4XOl09bmblmr6E8Yba9O/dcrSEqTVObYfyHA+2PJXABo0mYFRk5jp88CA0NkEsM
eR45oVv92LFKNJ/Zou6vgU8GAXVSgD0MQtmOh7jOdPhw/JFz9XkHJsjJmRhFRoCR
6LblghdEieazbXKgnHtj6iGrGFMSXQ2YGq3mXyEAPGrR/kIN0mKXDwS6nzrTGkak
wexvxLr06mvGdb1BkJZB2QRzpnhPfk2q1c/Rcda6quZ0wgEl9g6lfRZfF/RVTqAF
UcAc3mvxr2yShlQC+Dmorflni9lRXk0QJ8ST8fDtN3ZXw26iWVYHktSGhF2CUzOE
M3sM6qeEddlCGxEJNOBJyRQHaH7NeGRlUIojK9JWGZhn/0cSFlQ8P5+LKLc0gY35
f4Yi+RS1WPvzNwc+Dr2gkqdmNXks11ytJGeKEGI3nbUfAvtsogjdQJ7NPOoep5F4
WP6KnnCmRPmP+nTgXzpxhxiGcJ8TmPZjaze1byMpVJ9l/+Lqi4mhHvTgEGwaIFTJ
Lhw0iNiqEY7ajDuMykI/IX1T4+xf/pcbQYujivJY6o7R/odeY6IoELccHZt3iDcJ
wRerfi1dl37IqX1YED/sjj48vgAkI9RHiH2LuRvLfaiH3vqaUKnkNugFxwKBOKDM
TPSCri05pYQF1wq/qz62QT+Jh/XLntiJRyWJcrgtPfLm7eAov8c6LjN0rraFQK3y
BqpsVFrdZOrCU485R+maVARrBGbMHGqIk8vf6j9sVFM2kRWn5q3TW5fStYJH15jp
jBXpHFd6ixFcq4qtUrO4XzFS8fBl7VLE3tnMnaqMxkxmFh3brSufGWhpo+Tdrkkl
fgvwLfPCnqzR3Hxuh1tWNQ31VyhG+ojyKlV/9lFN29J974HFMJq9udzKYc0X3qan
Uvy7kqIlLiBAWJhAK7KIfYJ0Mr9UNC0t6mOmeYWx2vZhx6gbbaUumct/l5+AXzRB
FlOq7AdRPEKKUxGguKN1+J9yPwNoy2p1YpbrZ5NGD2ZHNPE7OMPucKcFNlq4FRcs
BKkV8BXrGfnm44WX4E77t7IIlMQu1Lt5EAl0qc0XNzzuW6kMIvGb7pSQoZUQ3kNb
VgCBo1j12xoJ41aEB3MEOPXlU83JYdyDwVP+eJrrhQgmAX+ZpgJq4ESo8VbhWkBf
M2YjH/emrDRRBjK5OyDqSHVrCQeOzx94iZuw1rHc7PjFKhPFTlgYJMvb/kmRokIj
CxoYJ4quiGN5yGVRSKXhhCIMxVJ8K5D1z7u6vuZ21CkBlDCQfw65sTRN0M6izlaw
ANxzkFDCvh2znowJEvgTan8174dpFu7uCxcxcl23H3RqdoW+8FzXfYC3UsylWo/H
HKoAtv1Q++uOWNZHWVWhyt+SiEW/MBLd24TvxGcY8OsnQ7iXkQT4dH0UN4dUhUbZ
d5ihSBe9Zjc28hqUzV3/XNWBF5A1k444oUOVCTrCs75wlVICna8no+wBd9XC1TeL
KCJ9uTKPAA5MOIjRf3XS8RMS88QnlWZYJdx5ZeNMKqofDqSLI56ColnV1RO3bweo
ECvIXC6KeDMbWSSinf4DFx/So1SIKQZsPSWbKWF8+b7KPi17xgoo2rM/DF8iqmku
Qn/lkjVJl5cLdM3RRr3Gpv3HTJVP6jPl5qNBp49MBYCmVGY8nhv9pClpy4TB3sd9
c3eK15espFhVulkAlZC1iEWK/cGQnBcOThQOVYqTX9eU5eYRXjzgfjkZZOW9t5po
iZAntTmEI7l/1tclqN+8LafZvIiV7dSVeTFM9KwNXI643XOyy9g5+Jis5rN1vZQ/
ocsFNu6Xlp61CksgP0/+0o3cpABV2m2FrEjQaHYL7oXP0FFbTP5NCbGZWEwwHWin
EBehuO519pz5M7H122mhBCXpDlTVDGCjEv8C47l0dGjstrV/fyq+TrCbKtqpB+Re
svAVusJwleB68ZiaYwiSIczK9I7i8oEVgp2nrNZGNcYnY8DCKg7hg4Zrj7IVORtr
Ai9Dr65Pyl0SzBU7TBc4cZccqvkv7SGSlTMjc6R3lJ7N20aNbjZvUm0CGe6qw/mL
GeS0iUIC5QqBL3dVFL8u3H+c+f22JFOo7Ip2r9OCU+pZIJXVQHamQTTbNaWF1OKo
EeJpZyNOlNOqHy6i4dx4Eb+ErE6LtmYvgESvsFSVKTh9Tt6jTxKPzARPYvDJbrkC
oY3HnOx81RwheNS3RgWFb6FC+y4YbRT168jkmMCNRoFnnuhWaZMppZtrV9wD61LZ
Wsa2hJkE99qcK8nujVwlE4ZtZZ62sgBNr/+XtbU/p9l/SqkxuPFZtiw1/4aDt6Lz
8gGUA1d5MwxP1A6DyFpKbIRXOC335eS+kG8e5k31fgBN9+D5H39cx2amFjSUcKU5
elnRy6Dnrp+8k8vRklen1ZLBvD/45XQkl7luIvzK86XLjwrj+Ktu2qAn7g6v7Sj5
PkAPkpMk5XWZIzgDCSGmk/VK2i/kqTHqeZzmJY1eNVds5tNQOwUfcOZ/6LY7kaAY
0BIFPOd/HZH6s1pdYwcNEPiifFxULL96rnXwZK7+C+hVDQRPfo2Jj4PDw/pDwPP2
pur1lFvWg3qspFrDdQWXnI31MPb6DmomR0E6FCPBLn2LfclwTRuZAMzW1xftQ1L/
vBoEis9ZFWOHBrqCJGb3w+7FzD9gQF+ZZE+qA6gUDOyHIo7f8OpORI0uh0h+7Zb/
JIu9d/7G8+kt/ArrCKO4T4LLzabPzFUcLzKvUswwkUZmx1mSzju2oGhV/i1QdXGP
x3Y7OlvI+gEX8/jZdyNAPcxp7U63jS0CwZC7BdtVeoNt2Kx46Uk+3SI47PLwfXMn
5un9Gn5NLpq/9e+bd32yyfeR/arHldXjR2mZkYVL1HHWO1Dr/+7asdM1tqgLVLkj
ExQu9XFi8dXYFmbklQGcb3/KH5oGyrhgjUso10+GpYtK/InnL8Xi7eJyPpiBTy57
hDCu/DobXk2eIpMqhJWmIjDHWFrS8BUIznTutaLNmJiw3xqBDmstgg3lN7Wh+PNf
qiHe8+OT3yPlseMKKUoF9MViAHtzsJA/y4tmoGleNFIPNSr7XIQ4XzKSCcP8+yI+
UV/J8qP08RIbFwShW9UDUcIjshOgAWHh43L5qgGIg88beP1WQODq3Q6Hyt2cO1aE
24+Q0mM1TOm7YcCbA0rxz+y/YcigOFdg3lcg2SqR63XJ0MNoWj/UtDL1JQjajkke
VWje40PNm2yrqKRaSgPfnnIsDcRxltC09h7vJa9pqeNGxTQXDIVeZHsCeyRDufoU
PIF3YzTm07y/ts2mWm85X/r7S20fzcf3CVZqgCE89INIH7V6lNHg+SY0XmdNqUPv
a/yhxUdIfbzZveTSwp8QMhYcKcEW3YWVdBPU5HqinZdknhG9unaX1Qcckbk0b7m9
c3Zk33EAMn7wa3GKYT7ddPlEwVqeAeP9WLqiAaFjxzN99eNN9Vzzrtr0wFnSa9UR
AvCSnHnmHq9iyRaelfKZ5tZfkUcs+Esr9hl8FWjA6oDpyyUOefA2+QQP4Qxqj2MJ
OJaiEB1nSN6avp9zuK60IAexU25Sb3/Zjfe6sVp5OV+MtQ7bMwhxl4DthG5eXPJF
SxD3ZwGLjiDCOA50ULPUVDfb7PsWU/qcBU31OBXcDWuDlaAbhXbB6V1BOOH0C5b7
PtB2tRwUfxzyc2RwsnsR0v/4gJKdLCpN1KIq3LC0ZdMg0YiKoqdAEEzUUguOF8mp
h3Jkbfl/z7o+QLDTcmN9tl7QIVxjRaAd28PHb6DkU2tMk0H1Qm/3mSl7Y28Dwfwm
N8qH8AQ1OmRyA57pDMtQOwUSUKHbIvHwPGrPATJUrgYI0btV2qKXMW78CNcSOOXn
qkFlu8LARRrRh5JcGi/W69wW5Upqn1BMLkB2tRG48tHg95b7TFetA86zTEH1XDx0
80lm9vAysrwt0Bs/0w88UchPOlhOCHEElDgbBqdONJwVeQC5AAlkjQ+G64M8OQFo
szYGSY4pCwvpXzDi7lm1R7gqw0lXINveJA3SgFL/PIPkTeogOTf9V9b8ic5qdP1C
P8NInmk8IS/01HvUM6ydGsHyOjnJXs1PYy6qw+FvWQ2j5LhwQxB7eiqA/aTY8Kw9
vJDNg7Kv8Xa8+PaARsQzXCpLcEtXcQji1jx2T/FeGdd8K95vHpT3LX4hntU1I8t4
X2NX7DbWrGW7hzotS1BSjZqOoMsfnBT6rWhr9MFn8V2ZQqGkv1nZiB+Ep0AFEcy6
BWrFvc/g2oQnoRhiJTgcOD9V09i07uG1+VGcy11cvXk6nefosxOm/FYxgblglY/L
qNRPsQ7Pg5nZorZmyvHDX7T++3gjp4bjqLLZGQfQEhGRhuMVAo78tyrxgl3NPCD/
8t3vJCNO6b9Dlmz0IUl17BanHASoblugIhyO4E8bZsNY3VvTQ4sCLuMiXghLUF24
zaJw/TUffBe+H9j3ndRTowoujuNHjzhxXihvmDSlK2CDrxEAS+ZLJes13G9bgf2n
1mgxXtJaifyLhPw3iVo1XTfM4qZbi33br3D6Vl8HD/ZCMxIPSm8kXbm5TJU+XUN/
aFQB7HPxHHyAxWKXL8kfkFDxGYFGAexic+bpKEzx1Xz7w8BpL1jBcqncBavB7BHo
WJkfTNB0Id60e0On7L9/GdtBr211MaXBCJIXiiB1wrLjgFbYwwCkj0tepnYeBJSt
exRbaFxvLE1q7urMw/QRlpbRakKGuElcoCAbsmJoIXstwMUbaCJ8Mzh+dP1BjXXX
vDefIoBu34gDC6zdblFMmGfwmc9BDvjhrnjUQgqZt31JIZjChEqZNlMdO2g1cjYT
BW0phAvG87w5TTpxpXQWOM/pRYWYI3XWubEIEs5jfUoG6NwwIDcAUa3C2wmLWz44
EV8WbarYGqHYNrUSOS2dwYagrC9H3wuBAYY/xDSxj8yzxZ6qicQxPm/+c5IG4Ohb
RuVVcq+sr+Y98rAguiadeklRP+IXvj3CS9SqAXZu27f6ACZ4rVJX5tXeqc52Yxc9
59pf/p7jRrkHh8z6N+m5orpuM0zbvCnOxdzRR6XZoZhtKZ9s7SJBTMBu3+pKEZwd
E4m8OuV/0c3yOpZyRsnQghyaXkz364qhl8k2zYtI0N+GwyMO5G+MIDAl3Re5Fb1j
fC/OXVp+SXRFhXS2hmE2dBw9M2R3qIyLWTkFy0CeSfxAy/0qoeOcJqNGGKXFSa3R
8RPzNtjPGrYKUNyL1x1SLKzY9hP+v9hcbxhNAozoro9NQDdwX8hMh56L1GkeWEQm
q2Bbn1YK56e6XyWKJQ9nHSXESKylVbMJoIhBeggWvUpYOL9fy1VV0rkoM/mED6gq
qJ1rg0A35Z8SPiNEZZHZzYLisvD9Oi8JjPWtGXo23dv4xuT5yvPw1SnBKI48s6Fq
kIojgKB/OCJT8bo0NOBlR6rP1VIBl88pf5L7A9a6b+KMk14R4Ky30mRb77+o2nH+
K67gDfCYo601uyuRXVXcWx4CGhCAVScEnKG7VtiOrGAqJkYCaJz52YI/zVRIk7ur
wtJtdL+5ztJ1bvpL/yGPY+H/157H8EDZw6D72sEvQS07iQQ6r4kW1J23e61pe7NU
kbFOksPR8biCLsGK8FDALswHgIKu5nzcO3u93IIOWuZxaGGIDbklZYUP4CrbrNa8
m1qibYxerC883BLVSYA7xRgnGhr8dtpbqXFWOrN5mQpxT2JzRoBM9n26qZb0G++K
A7H6oKvqNMUWSe8vX//EA04qGanVyBHxryXkP93THe65bN9qcZ2SfyL/yY6UAkZl
/aSNjRPVCXxL+quVsc1YvJWnt6ppjPiuqaAw52AjThtiGQ2rDyngPqNm9T7bACKj
LXnQOOL6nDlpePWkDSQHO7r/x4wfNnYXMdhsNcHBCbUJDlm+naLax7bEpFGA1ycv
frFWJmiwDfUwIuQ9IBtm08oWZumg7IC05vyo2bqvKGQn8sHbm602KHQUHicIBxF+
DOKoSfhGu3PyuiOiiPzk5SrNCTk0XHDtV2h6uKuWC8gmqwCDoadcM3CH2bsO7RCP
Ch6Bzb7EDv5OW95hBioC8V66Jnfkw2LKmsJSQkJPY/JJWz18ljvXncJltmmbF7bC
evaPXdfjmbwY9kG2Yopk4khwO2aFasNpRB++jt689v6KXLml2P2Ty6KLieWMBoHr
dNFwDBK107kM3gby9QnTHuXuV+Tk6EJ/wv0sWcIb27hxQ2kh3fp9n0j4zJo2cT9E
q5smaszqSFT4O6iqK8u2/D5xX+C50MuyiBftrNsBU33jPgwRYr+6ffx1qJipe4r1
ZZZO34Bb85UtdkLepb3U9H6QGxJEbjMIw5N2FRKDy8ldvyU8UETUIgYISTI9HXxn
Y7SWZueGaUazKVQ22kNhYaBkVfUn/LvnHDXhZ5YptRZIsTWbr/OL38PNmNs1b2Uq
tnSSbq5N+9QesOLaIdAuHDqGSOtMUJF8dbRjKzaJAyzJA1ln4KSgAw6fwtfENqcS
5TpNMLiFrbP8jSoK45JpcFela/Qduv3Oy98HBwnMQi1E/MkayVNVO87VgO5cdrkD
7x8WVg26cECGLGLBXBaa5DLZLz+j7MVqtC1drkWHoqQOR+qaEYC+Sb66SO1lL3+h
yzO6SfFkSERrcBTQvcwALkM4ZGZa2FEG9VKg5mtCGusBF50vRPRL2s4GOe2FRNL6
tiJCQdc4pMrriz2k9alGiRmy2Rf3Q5CPnokDGvBbvykf3IjKmE76qiZDaKFUj/J/
s+ShJ0Ya2WepP9MkjiOB+An6iyyU62+BNLOfwszkXvT4sL3ihBvPDzhJUT3Qrfi6
Q/Bwm1Wmo+xzzezfdFkmy8tl+jzViZGUldny/K/sbX4+VL1LphUhlz6Tie8ygzxu
Qe5paIZuIVTC/OurepBlQMNsNn4F1NqJoflNNZYRxOYnTX6AzeqdmMnpSlXQA28e
v4V3yCMMJlETuCLwVLkuyP9fValxXXkB8iE4VYi+KLYHsYQjkV/p6UrcYPwYyKK9
W8zU8uJbc2sWLjQLw0FgLbUNIULcjtWRV+PgvPcidxElw6OiuqkIRmxtXKrvLn40
4qffvJ1L/ZPn0kzbtlAP7RHb03RQMBzOnJo7YW84iizOyhSghwBX7+QuYFgwlKP6
f586ooznOjg2Qi7GmQHSS+3RFylPjBcSCip8jFtirIhZLhMpkqBXW9GEw+tl++gv
skJX9BcUGdCmjv05HH0shBcb+9w6ZclUgRybFo4lrsYfL9xKzhAiirN0G7ln8yQH
hx279XfEyh8pavYssyPPRJqM+w5vkZYwWbGvh6VG0ydMCmosAHsGXfj8FWabweOm
CvEKe6MTI1IxFiwFcy95LI/E2b4akYavR230Wuzwb3MmvaIt/jTiH3fTh3kygW4Y
H6oQWgx2iEt5Qrgq079b6LNQr4ycLcaJR6St28nJGRjtGyUMKS09pAuBkxyP/HXa
YiX0kECrK8MaK+w+plr90NIpViYvhon87IzxE+KDrSX0FXzcTn3NaaZutQOXjZhB
SzMnwvB/Hinlxi+8gu9zq8XF2LHFCMwbhJg7if0p7riz4VlUdBqCfE8In81U7Sas
vRk21b3x5XBTCcSWBPC7usyXpaTDoA4P36MTFYDM2JT+k7bpbiA/wlKncMGOfbvV
pjIQhIKkDaCmcgbomEaVo41oiXkalRSyHSzubLN3blpOJVU4kaNMLmOnLxH+7ANk
jTOcxY1e/FdS2UUcpT3yXVlA8/FSZWludGfJhcei7Zyau0r7fXz5kRteUtdqfcYd
rPP548QWGRERho05uEjVCUtM3ryrsKQmFtMOABzuKZNHXRFs8/GX83LXAjDAn7q0
YjR/32u0pr1HRS2HKbRaKuzD41AS4KBEzqn/SGHQTUhOvG6+3yzBs492a3hLSK8R
pVcQP8WJ3cFjqB0yWJiTOa9YRacDv7HXSv8zPY7StEsoVkKqi20kALSVINDUk0L1
Sc06L8JkLiBGS5BzJu6voawFcNGdGYSAQCiUEBq9MBRJYI99daxjUu75PTt3qADM
xQjWooQZg41yiL9NYBxXT4+oOvCmyZ5c+iEMmndpJdGMLX7uV1uW8AiVuRDkLm8n
bwBWUB+TtL1eShqL9clwPq267j0mr4HShssAcrBLC9h7qhFF/ENJcGgmZZcG3TVz
kLyKnebaeimUH0P/IDY4PAuaE/WZ6ngwjh1kAiTeDHpKQImxWirO6OXBcr2XvZPd
0KgLbglgcCb/XYnySoG5rjYWuWtTa0gukMtsHATBL0ACbk2W9LUO0X7MvoIQkRZ6
Pi3ZOSpEJCVEkVCqeo9OTG3KdB2awRCHkSpf1zYsOe8Cyn206Z3JMe1UxbsBh2ip
/wgd+NkezhkwKb2N3xO1v7PayF1hBzmYXPg0InUtM5PPXgRoxV5KwY7iCN4GOIBy
mimui2MFZVVrjknR3jNzAZQ6iLjBUgI7MhPXXmw4oi2hfwBelJWhZQ5CCclIlNYN
6FmqmBVYOtjQBhYL+1JzBRBNFO4yTJBayTUE/jXGhiFvOcms00EMfs1hEa8UI0lE
Y+k0auVVZ2goVhyvtZOcp0C8bVCoH/H7uDvx7hu8OtrDOqxcL7po1nPnP8DRVYSA
ALnooAfQ4cRKEU7yK08YA8mPcnRH2FsWUkcCctfLWWnnFAJ0WiWCZsKORAUWVUOG
JUwFofmO2Oi8yyWOBcW56Y6oZ0qTlYw4Wfqis4I609zK4IOPfXf2nEyIF/LJ3J8V
+hmblEPnbqlhXxUQbuk4YyfdAFCGxmUofn2Wx20bzYocUvQxHjYX+4XCE9IYteV3
Qmabiyer0Rb6KL36rxsp5MAxnMEOZsffZB1ASjc56n4orvOlNuE7bDwGCCxGBJUN
RPEo8OcM/Jt3uBq9ldj7b39cXIlEbM/XNYW96qrXDyfLJVzuETXmxGyasxPn8RK5
x05AuHYE/CCb09Uf/R1IWRp7ZvAxvjrzqZYHoXUCELklnUXOrhNIjZuWxDGAYwW4
5PsumncwRl/Ei1/oWaqs8E2/mdn61zA11TrknVkNVDZT0DSMk2IMqwdIc9TxGzyu
UF94GP3QPzLkBH9v/OrgQg6MDB6fd8ZOg5G9QnIjMgXIiGhW2miqKnGJxjL5QgqM
iC8B+DhQrYN7wa1P4tlKMKURC535HZjawksy3pOCtydpzajZP8sJl5K7bhvT3r+c
5xqaAWwBcvEHU+YtIznXch0sSYS+ToGCBcFQgifJy/eqHLHZb1Ddkkk3aNPIrsxo
8GPzkCBC6hszsO4yTngT5NMFS9g5VmTa8Sj8cPRKlfK62iO8OEwcsJVXDT8xEG75
0hEUlWvqqD7yteCfR+Ss0ztiDpwtg9X4WvqnN2baushNP+4qqcjLfkkkJFwiGbdy
SLBHmaKB9qwq57O1aOz114RYb6u8oInp3x4gJgW5bTdyEIxbNkoEur1IvkYbicVp
PuNXUizum8UKJGvMcvCffAG/rkLoQcsoI/eCggWKZ0BWUSp52fNpaHX709v0vg+F
W+PHM+7bjPkEjDeaVe5DcNo8k479KGQIuO0yzZxDZ86EZVV8kwuab5IduBgvW/rA
Rqdp2l0l/m7pBntjr1fJR23YwTZzQqgRs6JQnVki/fScVnIyIFAFlCW1G62VFxMQ
eAr1e7UY5USFfhyISZEopjsR6g9ipSmz3ekxIygdZ542RkVOSUG1yJWRqFsY4lmR
ZYZx3QP1EmkbMk/zW3JX9UzTlC2Dhdd95yw81RFJzkx6UXh01sWeXqazAlGj+zgl
mlbMLx5KmoIKcaxukGQz9laMkzSrNDz0tqRvydEAbn4YUKt1t9OoLVvt0MzyEWDp
yFxhC9lrVjeSTsj1aP6HY/ns+eeE3bHSW6JHEQWk2MK/IaigsdIqujuJKfixfjkN
RFBHyb7Y77SdNAk/yjIrKcJpP0d9ISsgX41yifTK2puYU8jyb8wH2JFvqDp7AQk1
cSO7eyMsUwnmh1ubPuPCL2b4TLDbbTwZkhbhcS1YYYWUY0U6V6OCTblBqYnxzb7P
f0IRnNJMI4Bne8to/Ay4Jkf8MMK+AitGA4bsEXG3+EMwXqq8VXrjnBjBlsx0sNQy
7SRoL2WFHJhnFQj/Vbu3zZR4rEaxjFTjj80ZqNhutCs6q5TL6bMlsXm5BrUFd7pF
/v7I5bUaSGitv5Of+kPTnDSv0LCNR99FFG8x7R2aHXE/ClCxqEXIei05ojyyZvOv
QpWPD2jqPGwmyhwkc8TeKWPFpnrMO1XA11IVbMkOZVQ2dU/NQoEary70LYx7U85N
OGC41Ys5hYOtaNuS8FePH7lVdlm72NszEBiGURJRHAWEWvFkJeudfakt747ViHfD
gimf5WBRIQR4UqJfofcrOxQwhiYyWicu+AwXuZQXcyOel14IdDzihnbX4QZFG0SF
3ROUim0HCeZj9U0t7n7jwMzognNu3RwVJGn3Zen5Uju+evHxM7P/qt9Rt9iqlOiq
iku+zawCdEfwUgToxgFkDFcs53haRK9iSNffY6IZONmzNsUAmTHneMv2AtsYw8CR
vDb8dLxqvS4t2iH87fcXOZTdrXQRsyiiJbmeAGgbcS1asVK0y63+LD+RWjTSULAb
GaOg7PE+DUKPN+3MeNJHiD71TjvwOBiGhcUwSY4I2s6uhkC1q9/EayTtL2ZCFVRr
TZaBuz2EbushKcfij1A2BpBEVBCrgKUfDyU1H+hiW7NGftynpLLtlBGq+3QbZ4HT
fPXyQkcQE3A31AsrmgTenpepahe9K9j+etPl/tRmRpVtVuzBOdpyj4aGXlkUt0Gf
gYbWJRXubs2KlNkqOfHumnj91sUCTBHifDMaeJQNSNuvrX9C2fUrbVuLCxkTJ1R2
mBB21zcWV1E1TNFqBItFWMsDoVJWOwsJ/CLKujt9+DngpPumG5arguYN3NGB7/Bg
Aiq1xeDwUF8G2z68Klhg6KRpVr+LEyxXoFkIhYUEYcjiRKNJfzJr+EfXEvodr0kb
RnHJ+RZQk8sVkPQybcVXd21xNanAcXY6XDGiKvK67kvBuY7JxMR8Q5sZJogAdW2t
wyMno195/eaG/anIR0vT7Iuu+nuYmzXn1iHfMqF/PCxmkBcZmF6cvjQktHRtXQk2
awG0DjN8Is6ba66rAi4LW/+sWP9nGn1N49nfF0sqigy1FstM4GY7DNOuRpOLhoa0
SpXiqztGghqOaaPsNGeCihUO7giZHeWT9nyTHlKWD3rH0K1ISghzoMBDDKsMMtrA
NOAh2E0gPvpBCxh1VDR0DIUfXgX73mDY6oKg7GmNeI/W9aMXm2hUfV2RVLnXPnbV
56Om4UcoGTakJrt7TCn5m1Yjo/NRiN26lXA2+gZe37HCWq9b9qFtlBDrGO1jzR8k
jgi7hxU9QVMFxse0gKD+VwZq0/TXJ39PJsyF+f12Jbkge8+lVVJPh0+nQBnmVPUv
OyD+7TLZe4lAy9t6DIeQ/CQrFOl4tW1aFvPUE0QXzG7/zr2zfulR9t3/azWLGaCI
9MrVHCBJp/IiFKJPfxpTqeM+OUsfN0KTzQY+LowSuBb1UsSyDUOZNXppVIOUR8tM
AjkKRiozPKslho5ExOG4v8IxasX5tHanv+kpwxb0S7rwY6gw9uLS8bw1eW0rx0GA
qR0b+7DlQx69My70jcT/g2HPg5zHCGtjOhhdt3+KvXPfFWRTsonsQf247MD/2Bz7
PojePJh2QNNdO/4nYsSKKvFSd+tRjbiGEhqSvyluqoJNBh6arI11S6rr4VUxnMFr
kDoBq9PKpHXvuxiaKfrcuoO4RZZxL7p9FR+ow0gGPMSCcN3pF+4jERh8OYPatgaf
dV3Ep682HJFyzS09jutvrCe+cj536WZWF4n5VFhxIVn62lwCnmBYGOKfTIoJZQBj
Eb1YqDZxvcKeUsp/Ck6Eu4nHyIOpQjOLuTvIM7vsb0c//KBoy8WMTOPGCcmb5U4K
8oQpe501v3tKOElfX6axr45qrh9fn0mo8AA+gxTt9ApVP0kooIlgx+c+qsJm6Hc8
gBNMMThaQ6ukRuClCSwdZ8mgsBHvp9dVZsYAiW+khf1q70o641lEkIJoC2f+WfCD
tWtGl6g3fMDvRww/f074fjd/P/YWC6lfm9zGLqyr8fWlfWkl8o4aDwnGsQ+r5RRq
aoONe+mutWvKgBWH+7VeSuKIzHTlaCeGZAgb1rAi807RLIK3yAam2Bz8OUjf/9zR
ZRTqkbjEUQgo7TpEGJXtX3Hqd1hJXnbM8sCTHgpgBdKvy5B0BLmBfFHI35oIeFxz
bi+ZbkvEZR5/CRGKFhGwZyhmQSK4oemXVI3j9I91BiKH/mX1ze1ioO2drkYPFDBZ
BwIdQIQtqErtStPXEy8SNcOxAesu4iuV0OoYLeZvQv/aPfLoSXgsr8mm8FRnpC/p
LBWQfjYhRBC8m2wnv+306DiTJZ5UPjPz1+q/IxDFYTrED8yv26Ho5BXbm3iZjyfc
pUhWyZpg8+KhABLgW7iR9VEDMJqfd2jtOvARvw9tFDT2uHwhhN+THOi6Orq7f1rp
6YrJ0PQsYqVOHWToTEG2WbJM05U7YnY7Pz+qb6F+2Ute72teeSErN1pbglePD9Ah
zPr3oJK57OAioTgHik/KYUUnrZzFJWDHu6s2aFiuXBOJfbzsaKgCHb2MYho7LuqJ
kd67y/RWoqArtX+RVCqiBLAgcB/izHldQonp1qWUhtRIORaidul2Bf/qm05WhTgG
WH7tsVy/b6Xkx2dC9MBdMw2m0BlXv8sq8Dwjg8ey5O/tIbZplYq1AXSDJUVfg2yo
ggi12oHp3pTQ99b0yN/e623sPDS/AOU2qFTfk6T5wznuT8z0WtYMRIt1Ro68Za43
/5A+HY/x/5WK0KryEQ8Fx72MKe16WF5NK7d3mIvmSWPH+IXqJ4QV9lj8fCeb7OJe
PHLM5oMIkAX5tYimkv4QezAiqTeZmDasaVNQyZMaPwoX9m82iqkpL2/oj6HeSC9B
ZcWZVEPQZd1Gbi8CgGfko4NdWRWSiMdrTJ5fN6VarpEm2TGkBnQJJXwNfKlUh6sL
PlYovqLZq9X1mGaGs2Q9xy1RcvASc53ZOPcHKbvdxcXOv5ILf0bp3bbyCbhqs6pt
F6VleKA4RLhfzhH01/xvY8Tko7ckUr/r2RC9ariWSNhbnHnclbrUF48DjsFxQNPx
dR0NGNYm/wVdFBkFpM17VhqF+35qQpFNBv3Ce66MBg1cG1Lgki780UvldpN216mL
mstFVJ8BtkELNs8Wt8u4EqeggK/AZgcplI2C5TFS01HH4il9tYOd342ffqbwO+Oj
zvkDGwqSKgnjW+6osMgwj38gO5oIT2Fx49MI4/kLF3skrWVXtIt5lVtdj4yZNrET
i/7hXnBsrCOtlfVNLEeK9nLYDwxHtNUgEZX/VV06KT4A262ZMj3vKVOyTschyyUy
W7/isyxqA+v4do1zez+kSJLr7nYGBbOKBLY1XqmHaiv78myNbNiMNkPDUydwrFE5
8O1QL6UwNkGWBs8m4Y48NrzshoerZyoUwQkR12eGZM86rc2C0StIQrXr28Ly6hhD
LzR+nTG3/4mYcTRTnz5CClsu0996BS1trahOKp/0LBfPzCfaXOYMEmK/8qZn83zF
nQBpXw8fenXLNR2OB/ZOQCsslH1AOCtKyjmCZqjjUGhkYYQ+estLKx6HwbnNVHfY
aoSFwoHjgmcU1SkDZjpqBuP0gB6Qi2j/0m1ChoLgD3cmcoPaZrrosvkDvPqGBOYE
4IDFDTjbid8LuhFSYG3Y3w/Xa6cKY/IeZmIEaCrpNVSzZwLa90zJaC/tJivPYPYz
/4rToEPW7GCrnnufYZMbDyyPHLN+Xl1WrIhMQquVujJ/X1kRxpVJ00JDtOjQGuug
LvcqdO0IGfL+hhAmlkD4U3441paaMt6//NFj7w28uUsQRh7r1q3gBUWz+zzh8+o6
LjXqdss5qoS/RRyrm58bMpBZuYyD105kXhuds4R2wDXOeqBmDrU2hsMJf48RHBie
gxHxWPK7gpvWmoU6RfupU+T+TZxPldzws0kTEDSjDCmmlqqmIjPLoTf0qwQIHY3p
fuomsYjGbBG8IGIS2+UsiOCpzhSi3p/EajDcp8tUFIllrf7KU+n6DH9ShjJi8v5R
3v64fmiVfv6UqDIar0fa9ne3hrw6JexH8E4XuRRFqoN4aKZIcR1w5ZjyD0lkOzCr
Dr1YWuAdd3Zz0A2D82TlRb3wuH9oEBTgyiuoib81RrW8vujCBxdo2jt88d2JIia0
jXZauAH4RWLEtFWuE8AwFiC3FTWYxWsGcxXIi8PnDibgc+SDtlB/fa25FY9IZJrQ
Lp9tX+lE9zFSz/UBxGm1QGSykxq7OnAO6ZbQQCEy981AYZP+vUSzlla/LJ+sBRs6
nnlp8sL3QXWRpxnXLTNt9dI36nnXyu8xMwEaIVPGxFwQTegBXWECzeYJ+J6eFj0l
yyvLihfliYm5LKnqCDyqedXYm0ZTBBE7HfS8e4yANn9wKbzU3kuexfnJ0IVoYn2M
XC2du6NVz528G+N1xD21Epop2sAtx9OhgsrsFR5VgcQS4PoMGTuxdZ3L1h+HgoGz
nMgIN2ZgJiXdPcP7+WcefRMu0v4dXMivZfKFHNTJCzocZNE/ZKgZxMYpps7SXR1y
udmZgIwlt+8tfGvdPUPD9LF8quQD37x5XeBDkI3zuzv6zZWP/Z+/gafX/hMGy7O5
jEgE0Kr/hSw94eDr7giOhwC1slH+1WCtysNKJgV0yWPTRCIsj+1+8mfCorElwh58
lru4wAj8wCtkZlKfUKsiZwAtku4YJHG0cMdJehDPruZb9sAOZQHzVJ+/oA441cq/
1orXZMm1M79groIxbE4FClw7NSz0e1+Zt3ILkYGhY5civ7fHSubiCP+Pd/l/Rr8p
Z8ca9MyG/CMtY7/V+3aPNtD2W2dy/LhaIGtXdCDJeW6nn3o/7ktcjidJt8HOKEFy
3bZnXCamHA07K3boYQ6bcsbzq4tuBuahrbaXZ3HiR5hv0XKAptHYlYNEc4MG4Zaz
wqYCvU+hydPJGm2wh1DmQDnZj3igka2wIMyLz9CO7xyuXYC2IdJcbPQvcKMC2hSi
Wl/QXPSyXr1hhE+8UTZ6KtXO8wcaz5xgEcbL2Qqylzh52y0lly6RofSAkaf+N1Eg
nVrOKlOcqiSecATUcpAuua0Qb4xx4T0jrGz/UDgBMu/sTYQgNrIP6Ll9RnBRfPUH
exCNzfyURMTOhvokOftJAS/FPsHPx3Rp+jKFo+2H8rIDDWoDEfd/OD5or9W+/Fqr
RvobOo8s9ReHCo8wBOku/iLCaL/+ZtBRUaX4rDqgTAWR8C1Aza44Fgbfrdp2XJpO
VSr99R4Mpu7nfI7jLjsep9kBu94XO/Ovo7QJYIPWx2U7FzfZp+ff+P+P7JeqGREc
VO3a87WYsyuEnJqmccTk6lMa4dDh18+pjxhFfVdBup5/TrWbT0ZfIPiETEcdBY71
W+mUY76ubhFx7WeRQVl0Pc6ph/Wtg4X2b13aJ7rqqFryq8hVHRQR+MJS++Rg+nQu
9yzSr2GGu61qX5fyNF9P3Lr0yJg4ZoSqRUcFGjx4It0/AmjZcrPDiIYdRoJ5sInF
At2sylY2BJArP9mMLpKWD3BlbwUmtzhKPhDnaKA59xpto4mucf2XkCeKLlrA9MVx
OBmTj/Dlv85NsEwSL//1ypG8PLYuJ+ETrqylAF4fjRrUMA/SKAmqNpNa9yM20wjY
y2MrFh/CsxXm5KHX2b++QfRazIPgeT3n3j2IY1+ABNkS+6WVK8WDLkUM7JYXgMdi
U6v7BeEwr+59Ey5rQFGgmBr/rRfWD5sEwq8Db7oJznlu4fDu7CL8iu4+2CfEVQ6d
eOTsN+BLCwwryMk2LXEAusUdUwG4eUHDHRyZAUPt+N/3Liiee/KaDziJJRDLI1qz
PZvAbYleR3k3tEEQ3W6LEpeXlrVZOo4t9mQ0M4+Y7zkeQ34cuGHXo+bE3g6vzK3D
8QNKAEr6seCXqZnfeyCHpC54jt/St/hQMxyuGxMOuAW5UaTHvzUr3ZgUJH8drWRz
SqaimROnPXEMdoXjFKrVVXmyLl/OdDu82aMHkT27U+eJVOfm3a5v2nVxch+YCBPE
5UUro0mXkWbRwaZ+QNzp98z/p1GG/RbUQ7uIVBOTeAVSWzG8JNoNbysnFy0vOSoP
+d20voyKCOxiTlboIV9dkQk8ZEuRjc5EFpy4nmxBDyGTENQJ+V26BPOm16eKq0cX
XjegWClzBQu7aqUHPIY0rM1OSA9mElzUzDckJynjbSyyuKmxrwtbQsUyASxL0jxU
I8qEr6KZYJJKIuvj30gJ68pGB4X/eRbfGVM1Dpfk7rdhUx0Jk1jf4f873/QEa5MB
ZntKZCbrNAUZ/7raJPnKhjH3GjQdIpCAaI4Zso1fp4OoT4+ByLVSC+diJuoMTnhA
4x+bHZc3z6vRXlyxdF/8B/bWC9f9bWVUbIbSCGv3OHnVFGo5RAIPaQDU8mxIymNx
CQriZlHkb+C/otoP031asvMvnGYNMgpkPjbPMTkQonFhjw/eHYlgqW/QldniZ8cZ
m+61R16khkmhU3rRF7GpqKUccVaw3EdQCPlRQ6EesmgsQarxSEigUsVmsVjmtGrI
iV/RYCt1s4YydVr9vxuemgn8xByn2DQytzG094S+3DArvkEBt9hQ6/lUufWeKW9h
GXcsrN+icZRc7E3oTmLSWAdQ5xHUjQHbeh4eUZR9arUv9P4L26ae3w/iX2lIXjiY
xuoTqeYOTkJ89AY3goqmLsSjMeEDwev5IGZsQDepnco2Nn2c0GT1UlEAxbrH50u8
2Janx9/6VF2jWxlumydUxBHnLiLsuNJYUKuzcpNouvxBmq+xftZ/2TrIQrW2VOpj
hPVaXzMCap/gPImBvnLBCGbOrjiTrgNX7mYNUyj2YaBDHrPpjB6onHkgrZSf35Zl
HusEPhjnIKlrSFnVGybcIhj4oGsA3MMLdrKRuJRYfTRfaff92aapC+AwPzknMvmx
ATH17y7BL/2WwZfb0m46qZBI/nv22F8fobghH35OMAE7yLbSO8cbgX24u8dyTmG1
+gg6Gjiqj4de0RMQAgCLD9zUeSM8LZfgJk565hY49WE9Ftdlk8caHDATy+TwDLEx
IDV1qWYPaR+NrKuE0zuyTinSk8KPuUuaXauntPFGM1veywfwGj0ae6lp8cL1PzuP
FEsLS1YUJLwtND3Ss3+8FUHEjVXBkRiXjbivzJZ2/Ai/S9+uTtg2HjG010aD8ihs
jCIrXJ65QgCcVesj/DTmsda7aqToYTxOq2eXWXu15BN/ck8QHEg0Qe1Zunngo68J
tWvs3VdlN1g+MH6CuXWWypfBAuGW3DbQHM+rYovbQCUS/kPQObJBMl9cPuNexLuC
gdXj0sgVVesl9ln9pzjXXapSa7UiHWBWtbCzGbDLj3sTn3b/SOcVQW2SxBNfrbpW
a/xbtEX12p4w+eGqSvdfI8xsIfsDuceC5RQJyKQTIKeTqLSsxnLknJY7LAsta5JN
mXyneWClo3LhxAKahtW0Dk4XkUWgJyBCVIV26iGDrPzQYUeB5bngPjma+xeExRHI
Y6Qh4XkRlMxRuOm2CanpnblRfAG+Hy9XQlZ+jNO91FSuZ5VW55Wvyrtw4O8h2orz
0mNlr3CW6Z5wv3cFJOzWmsTXbh+T8HwFxU3Mz3DLg/M2VPwh4LvmSy7l6XfsVEr/
+Sj8DVegUt2Juvo7hAMUn/Q2J547Gp91M7q4r5z0kxBMR7F9QCf8RtUfcAogvdOc
1pqPv0uUPm7H2oklfyc/ojrIOMSPQT+BojaTznq6JGZreqAuXlC1T9sypgjbHRvL
p/5x3UL0ZegapegDouE0RBuA6epLeU7n95KCuE3rSlGUZvaEG/GaI1KQp3vKERMh
ewzCn0OLLDfmfIijS5h7q861RKWMoSQmwIRaPNVX21TrM43iQjigbeYfkGdDeEHN
uxKIBJaTj9DdIi+JoZ4fdHD0AId67O4659KVc/9ZT6G8Ra0Dt31OQB5KOzeEJWFL
Hpe5aGIKHwurFubNGoGsFhHFLdR0YHqrtqcRoBlhWHqyVckU8W1ZVhx9U02GLl6E
2HTeWU1KAavKmJwzoVTn/gEyBXSBDv2o0BjvnCkNOGVSD3f6b3uugAEBH7B6qfyo
a/kq0YxNhURj0+zIQA5/PqavyNx+3lmLL01J1R3+snEVE9pjowzRqqdQ3cIWziYi
+1S1R2WyzUFCfauGtCRniC4e0ByjML8vGXgT8nE0HBm2pjTMNWB3/gDiV9ihn1en
Vr/B/T1LNNqLgDjx1kppu5fHFWwle2AUo5SiEPjt41r6JqnHKi79fboCP4ItHneL
97JTILPsLqiOkQoYrdtKFLJ4sFmw7oj16nYi7oh085A3alyyQojVUslKA4GS1Ujw
eqbxNXdZoMb1cPm63DhWRoYB8U3nYrPVIYxbzs+g6Sktw4lpgaL0tyeat7JcyKjH
9SjlaUXXuZ8wt2/X4yuw8JNBeZtS7smIduqmih/HdxuUcarDs6cyCrXh4DAxYoBf
efbQ0ZRijdnGDPufzzeLeXTZTyXQ9ceJga8LY39P4T+1cTWfvT0gDZ61vRoc0lJB
8gel3Pte2zmzs2vBrQawr+WgILVqisqXnQ0RLka250VCbSXcsceblNLZs9fg2uAq
nmMoSJUyBxRxIOfmqdL6hmakmaB5FHgyJsV7j3ULOiFZmptKe1AmoiCUpjIYy9J2
pvvmBFqLxkQQj7ufI0H2X7gdE3W8cda64eejxW7n5gZt5kZz4+gakmUcuv6bubj+
A9rpLPwx5apfvHGrYhU1J4ccZDd32xvrjCOCvbrVvfbixMXpIcTGst1J+w0eBUkA
eAcjEbD7E5jnsxsPY9JE2q5DzXI3rmItDlo6qaHZMChAoYfdAbgvYi1sg6RJNmpP
eWNpIaZkLexbXqWppeaLqcw2h6blhCzRHJaSVlSolonQwEHwvaKtk3keCuuWhR6R
c5Pth5jYrMyIeYXMneUqOkX75G1t5fSv8Hsu7Jxgvp1wu9QdbJGd6Vvpq323KNK2
TzmhUjyzBywbd2PVvInImppwajp5Rt1gMZg2DfJJt2cNlciZc4fnqLfVaV+mdC/m
tBCegglI8pYjk7yZb9J42i5KJwve+Fn40JKtoWbGbU34KZhp0ASW305y4GypGow+
ytqtUi6ngS6xqqUu1FIO/qROiQIJIMtTDsU1OQqsV8X8WRs+zcKJvHBSCJVXXjEa
ZSVUZMCNIYZNLWi3SELWv2k9WKDXCmwsomxZMn4H72YQ7rteh0zRUFIrOkV0EqlF
AsbrIGwQBaI2TM76vLUcOFZGaMZyOotGWzzVWb8UhGvjrlqNRDaR+dkwh2GZsSTw
rEEKfKe0ePtUDCZl+68KQLDgDJpIlA6XhCq905Kg9jYYQVGL4W0TEs2xa/68DA8L
KcgPsG977wQ2t4xhfqUC42+c4B7z74vtrVd+1MThuPm6+s8To8BQNV+fN6SoSxGB
Abrekzytx/mW64qM8AFYxrjDvkucy9B/fwf/VQankt0BNg7aElTJeIur5/N/9LgZ
stZk0j0+D86hPC3sdBfVtIjcYwhRzBKoeu6OKuqnzrIsnTG7ZakSGJAWm7MleS/J
On1QGnR7bTlPQWOIBE2Qv2PCLBq6e8F1Rq+ZxUbHKrGxvIx6caBWZ6dRHWVrSWy2
zdi7yTbNMU3PFza2wanVU+zozu9I1C0bc9qr7jN8nq2pBJ8icF8JknA77Vbt/vgn
PxMbS2stdDJE1hng/7K23ZixXRRe8h694RHnlKikd9pnQIFkwA1iXSd/UaWl1MOS
HG5NA0q1Nlby+20LjRiiaV4FPFp21D3UcUufvfW2zVfyyDbAjMG9Gk2D2zy8NM1h
RjzbuMwcoCXzUkL5iM53OdHhO8bnPRRhllgP3DuVKCzE2vTADV5TeULwndEvDVt+
4ff4STALYLIOhmIbIfIefRZxJ8UC6QkSMOe2u4GC7CPZS5z9TmerpHnBueWmT5A0
T1n77df3/0dXXFEfGj/+MKid65F9wqgnJS46Acab4ilBUTRXQ7mewrt/mdkv/+Ld
M2phUTapCrR3Vlwefr+G8BIk7TFRbvXcpR8+XMRKnYgXLmqazGx+BQW/eet/WKL8
3j4N5FdtLWqkY8igT1q8CRUslNxmtWNI7wfPgzd16IYYBjWbsyMA6RdbXiuksSSp
vjWnDwh9Jd2mCTtW9IzQpzHsLs1ZqUcCDDFZLk+fp49jkGXtyG5tr3vofAU0htDg
L9//ee8ulgarqdPJtbP1IP+I/kAwTCmu3/RIwK8QTtMBg7zbNHbp0h/5LMBu5FCJ
V+94veN5jBdOUS6vtfB/15LrQDj+p6rn7gluVY8iV6MtuQqsjadQkyXoUVXvoBjG
TskTBC3LkR/+BW3lAqYLfyWH2Dqv5apTMMWryjsthX72ScUzKTH8AFb/XFGfZt5u
8RZvXIKieNllmpwLgSbho7Z5Xvbc8xiKxoCTaHUcuJg85ZWOZ3talLr7I+P2Crx+
PeEMh5RwGBlM4IXe19KD1cM01mwPHaSd1VjhHEvXH4OYPwwjpe6Pv6T/cHZTHVH3
pko+xL4FCArGyrFhBnzNxjb1oNrY5AnSQhIHzgo/FnkxuXlzjdYQYA3uvhP35TCm
BkvywztjYy0o+SRW2AL6qK8SqMFcy9Atpdfv2ufZFu5xGjXa9uZlJQZw11FOeqRM
FDkzUxsVWyQH7iyMOylLcX80bYn7WcanYVxkKLR+wS96yaz2SdodJPPMtlSSVxiM
rawyvM3dHsJHAzMZ8S2DQtO8HAAFmKJoKA5qKldiiyEEf6E7ubtbSAfnO2r4IeTS
AZyoyhsJiIxGsPiunuxLbAHvY5iIDZDwe/du3ohu12SoXSR6ofcEqHp73ff5TwhS
uT4DA7yIcU+sl91OE1f5jx3E9Wijyy99QSrX/aU3zhBdoLxq4m+hwB59tGDlY7t4
aAr5i2lv+D0tltLxbfVczFmYWF3pbJLKYEoBsrlVywUXsnzPLaGlBlnHoLozGsCB
zNTv8QtLa+lRFT0jwx1JDTPD68mT+urM2+5wy7JEAlr2IVP91+gur5pSDaXu+xGa
QHZJzWGxeWJocd5eQuBzUktfWhX3LC+qzPJyTU8d9jL5TCU4a3aQTg/KT+PbX8YX
Xnszw82lMFQMke/C6IK5AW7YYZ1I1gGS2iKlJMfo+hZqwKTyRNkY3cz+alNNNtSF
AsVbSAH/jUBkqry5qOqrSeAZ/kO/5bwpjOrxCeW7YEQ63qkiLKH4CmXxnS1CQbng
8CkRzg6lTWq6Rg4/1wDuG0RdFiDl1zn+dyvb4QhBRBIJpnV1tLOjnH6piuR9fSP0
1pD9SkLQwhRtPynEc19cDy0Jm0KEPt5EgqYBUxv3tIr9C0obIn/g1Bw6h/iSDnmI
XpR/pI8mxqxGXBqTDXJpi/Gq1/InRMgj7x/qpwvEeIOjQmmtppE4rDkbDo41QZum
HSjbb81dKweZ2/OUxhqNm+ekp0S7OvwzETGY4TYcvjefZj/OyPNQwINFoz7ti7ym
W+vGMTJwZx+mtOPEiUl8X+s9vomSAIYz18enrteETvPIjMTa9LYNTHOdCNwgzwil
3rnHrBJEsYaMKdwEU3p+8IYoI9X4EYK3LnPGPP5oPlBN5SJxYBe1lTKqG68DTk4C
NlULszHOEHE0xlyHy3B+nHtJJ7P8qnlHiGz8BfDyVr/jg0bYxkC7gAq7ehOg34cM
ZHoAtMldoqwJnbp5LNC7Kbo/liN+BSBfIS0TmrHVMb4SM5VWw1u7ZRjUrDck1mxW
CO6MWDsNzka19keBSfevImS6CJIIYyXDYhw/ahlXGUmno46JG+r7EPpSL7vamDIs
ybIh+RCxtU1YUrygzuOhTSTb7D0WYwSon5sx239ixEWog/kK9XqIIA2U6LX17p6o
08bxH2i82HNYlbTPCoxCuim6mXHjITtpLx+xUKnFoOdhbMeZUobk4ODf9q/VjshI
KtOlfzvX+iQkq6L/QNNDD7Ozzx3CoGU9wpRTW4sUp6Wc/gWKrc6RcFxSN15+NKes
/9GgMSOgB1g4HFj1Tb7aX/Infe57ObdkNGZnpo0Jd1L0Q8q4u9fTSvTxf+JjDDyw
3N5Hxi1CkEm+oq1417rN6i7eriKtjgNTiQs1zHzsc5rN8Qv2Eil/3iK18wgf5gwF
+6fWjZz4xMFiR6qsgBkDP2IZQxTWUs0tEBVUBHc5iNm//SA20qJJf3PqXbLaX5Vs
+SkeUIe2cGQKas/AbOzzI6YhNRkOTfzuG3Awtkf5XZJCSa5v7yOacpER0sk7u1Fy
HBENsnHNeRugQYiW+esWbPHW8YyqDpC4THO+7Wn+1839Ui6XmZSAeof9VfKN0meL
1WcEW/7sv+GuVIcdI8dNHoj8u3wTprqgVvULoCU4Cb8YOAclHc7Twm/tMiIzqmi2
Q5rnmgsRGsLeT3E63b9m/PBwRQY/lXtWiCe/S5zbU7nmD4Q29MMK5Q8P8uvhwlC2
zL2fK55Tlbv6G4NHh6MqZ1yo/ff6s1Zpz1tWuTs7IUsqopfWgO545Z0OvH0Msr0/
R26d0N8QWaQnG0l4SaQZIvxmqRn2qLmTe5LQSJgGlcfmTcE+VquW7lb/vVsbLG2y
EUbz5UEMrnRM9P+jy7L/FCTyyxLDyTnX4AyBLToZd8O1dD0RjLtMupHKUeFPFyFj
gMED6AeApDEm3TuUFgfph6u/1R1fApL1qydnn2xa+d8/c40OlZvXbfUSbmIoQ+lD
ThDffVimgg4s254K5eE16pYpOq4LnSp1md7lqUYT82tti1UYpF8OAEuVn4EizGCt
zRXsmEILhJ2nF5Z5bopmg8bAhvtAlLm+4uVp/HIiJGeiXMjmlf2BZnv1DPiDp3yt
ErjVugDu3YmrOMx6ExAk3yslT/J0alI4+LeuBKiiEGXbIyH00ZUUNDef5/RkLLVm
HcLQ8xP23ahXViDka/6mZBga8EoMWG8l69XYs2x8phVtRuc6GanWFJzFhTSTJikn
8f4lxx0T3iQge+sQEIwBVlt8pqJncloJaNPLFJBeySY/2BGvMSClsoJLAN/93u6e
7ryBeqlQfIl9EkBOdcqhP6GqG1aGW85csbv4v+4hb0ZJ8Lb2Urov1AY/TIsSTxNw
jwi3nVHUV77vDnhDnb9EWeJ53BU0h/y9y7W7dSVWm0DeSfTh8zo2MyY25Qx0jUws
ta8RxXaGb7By4qIKC/dh+GhIpjirVlFHUkHfEI0Td1fXO6kRVEUjTn+eDghGH0MA
DPaBHkw9+scYCzan4aRrTUQNrzh1ufd4samnufsQgfcdvfEliKVm/4JFwMgWyfNH
fQq7DeUhpjng1wF3tGSdTXwUQg3oO+GzncqVrqi+qP6BXla6g2J7tqsf07STQ8jL
/PGxA98hR+LtqSlFHTPKT/J/Sgg3GStkJPYyl4zbdlQIEXvcEFnQlqf5o9keCdgn
Oo3+zX6xghHZdo+OzrS0dgz9V6wsnD3/Ni3HlLXKyiNvFZp+xRLz6LdOMkk1N/07
Q3nYo0MhpESfaS2vzwAutymy2q1/YQ+9Z5wJ3YkLSbRZSbACkl3rAVHCmGBwHDtx
sLAnhjGrpg89yvEqRBB07Kb1m+BG9Gz6GEWYYsxW+BMH/w9yACjp1WKdTDaiVr4H
AnKUmDHyMMVswlekn+RcF0PL9lbMgybLCaK3ibSSA6/6oy9/LP9f914xfq5lB4h1
0Y3+VlZPWsrh1Ibdl9msomIijDwQvbKWS3he5z54WGSk1zpJD4Ikw0vna/KgRw8U
oY6bblHx2etqXwUG8bj8mQOTV9gJJ5xWXe5dzvURK2sHqZKoporZIx/IRJdOQ8y/
136J3rRiqiFsjoVlXwZ6HEB/H46krj0WUgwnSFRbyxlYIWgWVAj7va/3nmyysU4N
ZcWjRIFkrS3iPemB47PjlQRnQJBlib9kWa5CPEZKftD+oxRsdSNMapAbSaKbBb0X
3+TMNxGxMvVNlD/DnZMe9M8qIY3iU+JSLRMV2AOAOeUecwFhN0j2kGBEkG1IsXv5
fCnJqiTbQknIhwUcR7DJDTv97W9jhp4obLjKizQ86qyKMsxvO9HPwVpny63HfO6w
WxUAkHTkdpxvvcv+jUTSoV8WtCSlemeDbwN0iZQyhoNhKjR3gIMBMjc1BPlelUR8
hJ9wjfplvZZlUvz3VYL6+Q/aXZ9kaA1wuSJ797xcoExbC88su4GXucj5a7teMPlI
iqm8JXiRt8DbGetWcvPkhj/xfaLZoqizTRBwhY3zQrySf2UPlwcE+nnbRDGUoXib
q6ai4x9Rpf9DxP9GNm5BBOHdKKnfOhfGkX6QJk7cA6bDMfee/vu2w5yE6fYNbXjz
rpHS6dYU2kxiCPAeErHlBJgz6CctoYUWsavV4MysPMZCnoIezA/xZRILfzjvC+aw
CgGsdPyvyMGZpN9g2lpVdPSJ51wkhW9f3x4VxdFmJP09brfKb1rSMX0c6sN7mTAN
9togq8DxlvBgPPF0tgR8XQKTumhuyBFQzOlXaW950/PCPvXrlkOQguJk+2g+AVVt
P42pNWgJbsDSipzCismPhimIESAeZ/ShX7YgNRdLyBm0xBsENapjdChN4jM34oGm
QngoVIsI96dGsU5sJ2uarmEDdJkkn7rhc4PIKW7aPcNf2ujKURG18wC7Srh/MnP3
4W1Bt56gel2dGCW131gPzSwxwIM+Td6RY3dIgIiPd+/DG4oaYwFHVWGHG/Uhi+kO
Iok6ev6KB/9LUlh6M57fNZE05Ano/V8jwP9Z/2J6eG9+tuoXyWaM3AqjLGcJ/1r1
3KfHEVFT5evie/zIvGgC3HVPtOQ52KXFo9C4qWNVMHXmTbBJUn8JvT28LO51bz0I
YP5fAdPCEtBTYQfEKS38hfSvgPxTA7+KnZ/uA5XH59iD+EDr7dUZZWXC1hZ25WqU
T7L+bWsDINNpDJvENIGzYyPvrCWDKJ3wo2XfArn3tKtBDR6qIHyH/zaWDWwI/rze
GuAmOiKvhRLitzIU4HDXxIiYuIG9lLw7mr57ghqm5Pq9CJw+U7C3K0LbwJlSfRYq
GFzmfDKRDvbgnBYkxNZFE0eZiV90VblN95V7DH/zIKtUELaVisnF254xdcMNsxg5
Hf6Hx3Q2oCIjUaod78OCLws/J/z6jHgbMfOA3nTAXaxZfd/z9ig5zZFQewAtO1zR
EZba66leP872bFpSgJwHLYOZb6AWXlBC0bSVX5x7H6C2S/lCAOXFe+N71EfVfzqW
pG+dJ9k0SRuWJ9QBetXOPBDpgwSzTdgnVt0EABBWtxocrWHPDBtMd3hSgZ7SP6lE
SOoZrYsis7JYfqj+jIxfa7JHThOmj13WkKDCsANvKOiG2vEYHkMI5tDME0iK/Otn
aTkmBSOPVt4TPeda+0S9E1JZMMZPcKGSJzrhyv+/8rtX+a8GHiSw0yJBjQLj/ouX
8bgKMWuqCc+jFALarpcDcb+ExVPktcLm/kLVEw+IgtVCB842958ft+CSeRvdM017
qQ4FLIfGZm2RV7gopV4PKKpqJuzq1lEsyDRlolqkmvxDD1sF8B4i9oB9s3Y0ou0z
mMTEYYGlqi+hNL1h9KSq33Iq9mFBYvISvT1vpGpG2nZ8P8FRInbEJCRDFf50qjyS
ZNTkb21tZfUZXhQhuiI0Iy8PJVpaipMo32lJrmhm7xzFJj1y6nhjT9dZ3luuWBaC
fesDMOHupGcwpOC4GZDEt1oWlJSO4ZkvM04ewPiJ912IbnvD+EAFvzfjIGBcUdOD
QDfAJy6kDJI3ozrk8Yp1XuqDOlEbHN8W7BmVJQegQdcnHMLnHEp6un+rjQmasDop
RwdvOZIfpjRFWQYJScpvu3BLonMob3BoDpV4uNS2VCPk4iYCQIc5ctUyhzRHpabQ
2a4hYTv3FfsclcpYABvVy/6P/844+wAeK9oPAEG5XEP7F6maZsi7vXSlJz6jNgfg
KhYcJr/1mkm7VeFKYQsG973cN0yL6Pw8je4btG+TGPa8q1hFrLhhdwvh4IimLV5a
osJaXYQ07GLV0XnD8P1NaCVFsNwXfBpJONsOrHXOcd77+3xruF5KgI+nNPKMdppp
3Mz2Q1z/VVwM4FM7DcN2ekEh5va2QduuHCJMOlFEnNBi5NQGE5Cc9g1DxH3lCfng
dWRdhhvA5v+Zn1fkuJZ2abpgeIEqppfhFwGrvataSCb+BK3ucRGtRv78y8bR0Wls
lH+TmPbRcTM6jv1ENsvw7vOoXWn7TnX+MugXebnI0khdsjFNp+Fll14pbuZZ6bRb
RPqzMdDIvNvCBJ3Fxs6kDRAPxKH9c7g2a1KHWvjIvaGkz7KVIDmuVcgrpvhArsOW
kIRJGFOBTM1n2bY33gVNVg4VQrWqC49AGLkKTj5+OxU4hdmDqplR5UnAfW3ZN6N7
gy4Cky5QVfp0XbaLO0OePC7kg8baIcPz7XRETMteitYHs6aokfOzTbIq8enf1eEb
hU9syrZ7J1pI8d30o5rbiPfAvyDxltrOTd5AA4fUPAYBsZXJHLerab6grxhKkf1/
xvGBrjOIGeW+4f+8JyPLkQPr6SuiapOOL5v76G/RoFJyw1S+iGwCx5dZcr+imx1+
wCK5X2c4aB0rmTEDiH1phIzY3VzSUIGmHcM/BPwT5hW9+j5oCnMudBOyPwDKFcFi
QQdfNdp2bRU9Gy3rfnx5LvBTf7IIr+DUDA+Ivw3PP/pKRY3NWWh+qR6AkO2uP/BJ
hKftRUhqNQqe0aD8PpSIao25pwSIxHeZowAvyby5dpbxyjh9OcGNIP7gxNmBMses
2jS8+jfQuI3NZ9Rx4FByw0LK8JgVxRkUoMrh9bohnax2exe+vacXhWvtEWBomnCl
NqCEgZ5X5PdMqQXntJh2Gta2wtX5eMvpDoWFluOg4wu5PE6P9LmKrvLpq5MFT5xc
8WPHslI46LlU5Q0x852gp+eIV3jhr2UIn4HoC+z2XQuKVnHdrkex6ObxApPRJVxg
zQBXABSqELuzk+iJqp/8SlzTHuG/Dqi0vY3uwqNAa56wDGjHIDAK/6gdX9KpX9bt
b97IJ677bT2vudA4rX1DXty3bQ8OhYw1ky9kvIwgcbEAPASzclunChzqna7+b4Pl
YpttO1ebb36EJex5S9OB/szOLvsTfd1m6ChtoO4XXnpiNcgtnnOulCyoD2oNGU+B
g5z5SKhDWimjDfIg/lLThbZt3FzqEncpozSCYvjw7CJHnGGiORfw7GayF3w98VUQ
0Y75G8zJmYLK9bXNjjA3habVHJu2lcGY+0jlMmG1CSNnMDqreVUxr9GsOVLmLXrq
Jdb45Wl+dj5F0WQ/CzzQZN7HgTWrQm/+vaIMpqpYatQsCtoU2jPVd+jhL4XmUpPk
HGL1IHt+nNHuDby3UaGxTOFK0eGCSo4FlvwJH3bx7ye7YJL37EWYLljA+QiIyWav
6tMEw5Qwsipox+J0ya6V6VJZfpjHbF7ip6sGDnCc3xyu0SKpzyCFqQyF8hM6Zo7n
J6b4RPP0HP8zwYv9XTVa9dNBZ+OX3DgaIeLjDcQtP0bwyS1mBs7fmCYVJji7gYhm
mPM0HA7r5wmknf4Vqqq9oaXidB5tjAvCUihCmtSTQEIxwsUvtj1aCrcUfCftZTPe
NW3juc/NwP2pl0VmkbOugozI+PicKmt5qaK1VpEQb9G47l3yMuFp5T/5xxV3uHwU
wuSwa6r/SpfcXRCfIWYdmxBGt2zlJp0ZwUz1LOIM/zLYmIBqwKF/VaJFYRnjz27e
dkrQt+MmQZEgWdT4bTTKnDqh8Z9CXBnwPoQrXTEOVxWl6wqM8oDVq/ZxbMnWIuGm
IwfIlvmoFW6H5y/WTC0iApyy8akPXQmzqiAHxbx7ctQNQXINsv46bcqS9oUUw2fq
Du7xcjC5M5Y+SVH2OJeoSLg1c6e+UyM3l+qffWY1S0vA8iDeMReysV4v1uVJMhOf
qhOYywXz9BNQciNpOAWYydBBILZQLrFXrKP/Yps7G577IjU6ZBOJa420SRtDJ4BV
fk17r3BD7x95/QnIhUMRDDZZvO2jF76oSJ9pDOGBgIgR55ESrd3EK6Ngn4EO9q2b
Vf/JO0jvZapBx+Qo3VyOishIZXM64bWTMw4ZW184jHb4Ed26JCYLG5PtvdUudNeM
MoV4AJhkJ4FfpOIck+BEgloeofU2n+VEfhjhlfIddU9VEjjq/jGqFfG4XUVqHjAO
7FSdLuLDrn1q4IzqYN6ycQ8Jcobgmu0j/ODJe6Q6v7CtRMX3B1s1R+yovYUUZGBW
dW29yb4P6JEyIboA5BKix6ORcKDXouJH83ErQ1NNLH1x5We3IvQghT1FppvH0uBT
HvbuZzqcCs18HpD7dsWZc2IGFexhxXWlEfOG3BOPnq3BSisM/G3adv+IGI1TvBGJ
h7+W04SLazvcw7Q/rGhNd1ZlUq9p0ERImzbLCzBItrPWLcqtWtgdQI3gfcc7Ruel
z/Kyc84YakcM+yIDr6koWNuj2TLS6bXni4iAhM79UWMRE7EQkw2EfWX8QXZde4rE
IRH5Umkhi4vSY4tC2ihuC0AbjNnQTP2EKifbsExYN7J8JX4irvHedZc/pzH9AXd2
da0JpjIgi2b+NIHhxvuEj6yuH1p1ZBZp2jldXU9j8GktBR6KaOvQyoeyDGm54bj0
d6Q5p955cyEHppY391G+UW04l0aZwgNrAKt+R2xPtkPSIrfL14lvm35xcgxhfisy
XWVXJVzWFQTKSvNy1XL6rEi0F1DrrGEsQArti6m4pmUur8UbniwTxwFyRdU1q8l3
Uwxfx5cMdozKJm+erRi2DeVmoUotvf8ufEPoRVtkNdt8xIFFimxeeqGU8DAfHOQk
wSqnBzQgOToEYFNcYjX18RIZ4tiKHshyaRo39AMyYfN4xCBrvygHoXyzdauWMUc1
tK022s9KNJkKyG5J7o/I8Pm74fkLIhSd4dyOvbtv/FDC/oPxiOtn0lyEk7cZ22vl
kKnhCWggbGSz/rtb/UxTqkiH/C2rwz/CAvJLzJcDKXwX9+Ap/+n0hKMm3R17qz+7
iap5Naf1AzgqJ4U+UQV9b+jRl+5+ZsJOVyyf8U7kL5qlim7l9Yy8lGKlCxLQWjzS
JeydOBrRc1LiJ1Ki6xGEV0wcwFqlS015f50e594gBm6qeRJdAlNU9HC0bqmZZl+P
7F83N+60kZGmTOyHvvgCnn33xzSbpjWPXU3W4w/PBq2n4AqUpEpbG7rXcPbf9Px8
5ydEe4Ezys8xoj3RNZYlIcyG0DpzzWePdfopEUZhQCp66hcyo/XsAVO968BhVstZ
9lzHKjx4rWhHLaFBWQ7Pf5VGwwMoUa80OFOgMkzesjqTdhBdC/ezuH+eaBsv5Aev
Trxw+VutnsF4sQp5QEhCwWsn0jSPN1rnpvkVdHwqO0CDxd7bzK5aEYylerRss4+w
HX1fYK86EH69koc11wJYqMwfKP+VeY9Gl80D42crLTMqXJmwZERBp+NWFq/FiZvt
cxeTIKF8GQVYz2TGuYAWGGrZHDiSw3hmGHPRq5xj7hIc6PwAxZ3d5f90Bgao09s5
A7tXKezCmbSAEjJb6RlqRUf95COnSqN/y4tAGIAsJXelnw6eJCMMJLm7hNbmyaHV
/7SPDMskgqRNeJRYx64fTZlDBN1yFBwdZZLUg4SfA3iz2c3tMFbi/KWGjyT5BZEi
XuCWpMoz/Pw+hMzqudIZl7ux5v99zLUSCLFQ3h2sacuiGHI1/Jksi4XBl1B2sMRJ
Qb0HVcXc1VPgsgt5NXCWcT2hlC2jk1znPXoO4aj//34eZ9uER01YsfBELNp39irp
3t3qEv3LPxjclugyXHjxVV6TL+4aydB5WGgW9LuawxFRqI9G03VDiHyCFr+HFlMt
2elUWES+YBLEjxnX0d6hh77mniCeIEz22tDrt0FXikVS3Al8NSOcjVWf7e2M1737
4EgHKV9B5fdxKS9fRSWx2DVeg0d6c8SfSLaSOqKmyqekf2DPm8uA1J7gAq4exhMp
/VH9YWdDIGqUbgQnHdGFLVtxIfmpwxHImCyNoakIDx+BOcNFybBlb7MZfnpX8OJL
LCjh83QlACos9RQqjR2yqI9WbFY9lQNtBvKXLWkxNEq3QNGxau41JNGxIgyjyeii
KHkLHrXoQlpkp6RW1JF5UJORCBTQ/1D+Ol7Wvk1dFmNzUVIKXrHr+qH/LBGsJQza
82h0U0EHtbgX7VltNMjfLPG0MISOH5nrKO1uKdKJIIdvXZESQe9h396LIOWUXEU4
FFqZyMhv30DNGomRhBPu7pHcSdSgaDF81YLHF6bBWXWktNxec0wu4ka3pSDl0hdH
VKRJn6kpuo5vLCpPH1fOh5Kf2QDoIXDDh6MbrlU9A6SKTF6yFyASjAe6gq0dWHJj
ZkezWZaStYbPiYWj29WQKwBSquG4oaJoDCJRbt8uvWoeKMr16mZhwszsoldL8dou
2uMp4lkhE9NpHDVb/RepFEOZyK5qGMKngiU+1lOi7b+lBYbZA1c88x4YuWH+AH7b
DVGVzdhqLZGmLsAK8Yoek2Yledj6nHf2PXXyM/hNngaCnp6B5jehaRh1AWbAVP8o
mRQw337JzrHcLgOvdPXmmLo4Gafp8sOtAOEVYYjaj2SGDik0eHkbk9xLu0whCT8i
ceYZYKWRqVP2TG4Mgbh8WONiPXvZ3Zf7dBscZHF+WtvEhz0beE3ZA26kZU8srR1U
VYoaN5k1Ee3F2G9YkXa57mPuGQiJN4Sju3l1nhmIHLM1ohpFn2Vk4GSBLQBZV3/w
+4OFuxStJ7iXC/IUpmxIpYSzYQKoAivMnlHj29P3sqAHA2qnX4S4R0no863QCbtI
nvDJj638A/0fFbWPS87GQyxefJTolU3L03EPcjw6fuLyXZpY3Plp7opukTZybmxI
nMhR/0VwkS8qxUZa1S4THZTcbd8ZLqCTKHUqIV6ZDDKo9uuReq8UuueyNX9hMxjI
I3uZSL106yoAcLZDKWRRMP5vZPuuchBDceT9bQyk7wh3dvyyuwqOH4Bqg94XaCn0
jf6EQinZ0O2S5DzAh4Lwf4RHSGTokVsqIETN2Hc22YOwtxptBXv7B9y97d3HpEPo
9b7xoNQCSU3o8JRRw7K516u2+U7lxeP/L7grgVE9OV/hO1msfSc7RZ0w3BKE/wpb
26+Dm3ZXc2v+ew9cV0CfCQF3DhKdzyxsiZYuAEdUzl78T8s255x9JopbtkDOzUoh
Vh3jSdciJV4lQ7/+v+YClIjB7GlvQvIkyL9+u6mrNhr0nnUOISv6cD7Pce9oMcsw
dz0J6nwNHX4KavTntXsqLHTI9hupJ6c/aCdtwYLn6UCEf8hyO77KgQs93TXMpvF/
O1BqcBOVfvCFXRds68JB7YHEpGUeXV0abK44sn1Oi7xfOpcYXxzFzu1xVc6BrdCF
5q8UD9G7NDX+PAuGkuCpSA8Ba6h5RnETcXzalD338Oggi+mVUb/6ArcBw4qa/F05
dDiYnW+EaG5P8vPTOntVOvezdZ2JK1ifZIgSSyw25M5edrVql+hCSq2MUT7ynmop
PjaxFCIHVo4ajOaMDX2sbcikLXojlJ2+R3f10zGtpB2geV8Hm2mFTyvQw3a2943b
5jhxtv2EHeuSNbheEHZy58eyqmn40kC+wFkUh0HZ93xyXZ3KvFxI2joZvkRATTl4
l0ViswPgwP06LYaXRNiCIkZA458ZeBHAUKMewvDY/4T59lSwTFQFjRJ9OW6wKgUa
MA/YunHWiBMNE7re4A7YPZ5HiCjID5T+GV7T94x7tHjjffkMiddmJtYGajs69ZW9
AXFo/MZ3xQz2Kal7LCiP3iyE535qopgtrAM5QvbidHNfg6P3Rdp98e2W9QhED6rG
LAw126KjWfcmKqjr6YowXBmD2h9AxLhdnqmH5NyvAeEv+0P/ayAuudF696h96K9w
mpK5OT+FQVupGB4qOAtYEkt6MEiNheaTe+PmRxGrBf7lIPIMD8Dia71zC2vH7lAQ
hMg+tbMY+OS/I9nDcB5zjyQCQiQAxqOBMWzmIQU3JDy1D6ogfmHeiISJMhoM7sA9
2BPPpivAB5FUYHds5WEjV/2yEciOBWJXf5aRtOih98oA++n+dPz6109c2NHIl5EI
bsCiNXW6OkKgtToJui4UmyT4kUYH1LAzPcD0ArjV6ZYGNsY5Xa8KNsgrbCbO87wc
aWmfI3tfPazGuSBRydqLMHju5MfV+VKKkkPaem59quyVnQe/BGRz7k51qIqg1F22
+cV36k8bnfeiL5HiZIBmLWuSMxA1TiMB/RUuEpjaBE36GbzTsFGAb5F7/IIQ8EOn
eJvSmrAAy/7OBajJ5JFpzuV/C3aPCIjnkGBQt0K/qCNw4c5K7dZh/cGIIB5uwZJq
2pIMO1HpP66b4U3x2KbCoQ+Yyf/5lZj8hmKXiqwTE9jADD2cTb+pIRR9tvHuLspN
RICbfIbHteuXuGlgMHEwjFdw8T7wa9OQWpjEUoeC0gDnQmlNdcegsOourcsagBVV
Awa624vRInPy6h1UhK+fZRgJgpe6JnCBe3Sznc4UxlWZUPoDfnmMzLwcbQxPcbFv
wRxA42mnQ3QACCiIg8EUd8DTw4B4dzkwgqIEWjQw/rl4EFtky2T+JhLXuFx6Gdl2
ruKANIafUhbQz8SHfQkyV0FZWSwM9dgyDm4BCE/aGPfFt6NvnwM2K4jaVly4jlTD
OLBNHPG0BkeApLMkbZHA474jiJAyrd+AFulW+JPbQSiFkyu65mqfR5AbEjBRxbu4
2sXCZiNaz64ZSI3aWSo4KrcETd1xqe2eHjK6iZ/Clb2gQJmJvigYukiCwxVg3c1/
MzMbVje0bITjKocujhoWc92R+tVNQiTsW42Ci1JjQ45WVGJFIxFF5+ZoxHPrj4d6
0VebTQ+8rejSPAh2xuIkyR3QZFmFyvGmh9ixl5h44uBCUMJQM4zOo1wf/miGTTG3
l5oETVnhSgWPGYycZe8E/A5+pTORefUHuBtO6Y2K3fXoFfGoc+9AH+PjFaItG1IM
Q9cFAF2xg+YMv/HZHYhcC6MWSx/g9Ny/G7C62je/mN8Uy4GHPH/eEt47bCBozXnV
55Ph60LglS47KwmBJlDpy8Y82u5lYFZhnQvkBqxjRrq5YCjZ+ynXa/QOXgbCAyjb
1bCrTB0j4w7dl37Ax3Npe5NjSZzmFsUkzKP7bnZDzNvel6kCju6Tz69UcOljeoAU
W7Mil7SWfz3TX0tsDuQsDDVTkmU8wJzjpPngA04AG1GFZ1kAaeqOrYXsWM7c4cLN
Tywtr/DfI4d448wrXGsUpiX2V1//zif6F/v/rGmRsu8MFwqRL8amr6GywkQ9bB6z
pe/4Xa+NHQ45gRSrDce2KB1RJtNo7zWFXP0SoU0i6KMRLWOIR+d/itwTpnWLwnR7
Lnto6VxGmWju+10aGZzy46N+rs+A3sBCFJcjqZKEzk7/JaSz5pQ39gstOclpXSv2
L0I1BEklqJRtsaih4HFI/5Q8DkEqda26ub5XoVTpq5AUG2qdKDItqUAnx8mcATBb
AfZGq5hbbWnilm+2Gzxz9CLfTL/FJDzdX4m3QBZLy7Ry+nEBNvLprylHW9k4tDS/
SDlhmeJHNVTooKXYk2r44loTvY1LC/ZY5pUMPgevznkoVj1juZQLviG7pCtImW9g
0hlQLX4poLCK+4jtb05M1r7OmoFs6RSruNs4+rJSDekw7FMzqnrORmmJwltCmmTE
k7ljtxUFo9mo1lDOf2JreIZKb/7SHW4tdtqyVWMVEglv48JAK9gp6NZ6O3fkhHec
GnR7FDFHpXwa+u2GYkjCHiSQJMjPYdlDRAXKTipzvtFaOi/5Ye9P+ap5NuqQZlyy
Y00j86fnu6d/ZR34WmDupXh2d1xQpqsqpUf2ORBZBwoOKNt7rgM4dfwW6c0xgoEK
BYBSm5uqxGcTcmR0TYXvkoutG99wPvHG/3qEUHwslvGW0Itv6HDu2mEMzylioI5K
aR3DoZDpHHjETv5jviVvUax8zOtGFAeIfY0LVlKkMsYEXFze4AV2tyBsHfTsj4Dl
XykcJD1Kf8cUs0JC/GAGc26AeiNaOl9fgqrv6gEaa+sV+QFTWLNd0A0G0nz8wGlH
kzlxIDhhWxouTHDeela1a9KzZ3oV8gw+SM4ZW+z2y4S7PFQ2FlpRuG/nikE0WW6z
TQzOUeW5Z54MkZdJHY7kINsHQP5WSynf4GomTybLRkS3O3bhQfSRXckuwBPzFtnB
+Thy4EtExvWbW4i/1piLiOQeK1VPwjo64qAznvkll8Jd9OJ2E/09BxhMN6RKFktd
Gp3KQrUABEAZMpB6L1kCPx5v9wYgdAxOY3RE1YTmIVmjzALu9gI8zeObPwf01ga0
Bm1spj9VlTMTPXVj7CmAbprHIpWcfNhcRybkeSsPuDmNjN2r9DlEkfz1tOUnZ4jA
yixSxTAO7FbaH8rEArKCFQ32cC0CEYCAqfVYJv/leuuZfht+TG1jZ2KTo8wb8mN2
idQcn0QXSBF129M9PNPYlHinuGbnxgpsVE6yCBcXHqDJlzrkQNHTHQu8gPlmsS9B
ZsGrmnjMBNo4OSKJVMOxnECOB5UGQHZsk/bZvnZuL2seODmMJcPZg14LiXLQkpBF
CwgAUFn9fL6TCuPeETdNmZXXXkxOxj1XrR3rJASKcJXQjLZz6i8r/bthxBFOiwZk
keyJ8yeCi9M2cwmIRLAFsmZE3bcP0Hq+Gbmsz+Q3VMMlMflInYDIwCT1Y3b6MJnU
/dYoIl+GpubTXCFmpKQNwLghp+9P69LLdeQ0UiUxPKXmUY+d6B65Iy9qMWOWDlKe
Inu/Ww/+XtcQbrVnaLmt+gzf9zYsR0x1jgnQbioJFBcy580kaop1asECJ06nlS/c
Vm7K95z1m/6m8wotY35GYQmkRKcQa14J9j8ee/Cj7zDMlNzPNYxrImyfdMaqJ1qn
jiun5dchx8oO0OZvhD0eHJhXYPn/XAUBnNfyUAGNpP+6kMGY17zcNvuA+UgxfRLA
5JgrcyaGc81+oqfoV2bGccN2SXdrdS5RSjxFAoMpaqPcyYJXkfpJfe78X5VhIkNO
FXpkfNdBBFZSj9f2Hr/mAgKyqjdJxrARoAdEPvtYp/465c+7KvEp6oHv4UsU5j1w
85xEAZNlBj/HWYHJqy2/jItvMGgCzWHaPvnMjFQ069uFQIVLq85K3ViOYma6rWzC
MNRP/NmbNu8LcDk4IBwV5JrlorotlDnNp/df/7s3A1EQq2a1rDWeOPvmDCB1PADy
CvH2kq3mVf+MJ158kwkaXnkgaXUeQ6WLINR+CqvaOPskCVJAJUk5GXszS+DwWzjB
WY6YjkG0XeT7fiuJKSrbOdzCz4joELBcr4KsuAGW6G1v0yU4azXVkNRvjpq2H6nC
R5nrDxuwHx3fenAdFbE6Tdz79L5KhZWwWqd1kJ5871jF0aCgbcJDoxDfvck9d6Qn
s2eqMbq22mgyH7p9eJR9rO9ryrPg9RWOzRH+SG4BhkN0L79Co6BXq+AYso3RP92o
WMspXj5kL9k5m9RTnVE7l0ZcOD6Q1/gV5RKE6pnSwkDXpp8snuQNlvifWZkRX/Ga
ekwqvUHh91lQ3Lhw1fGusVHj+bIvOYBwsUuEnpZUcxxeFoI4vShvPokWPWPFHbBJ
Hp91hzRbzE/rzPD7OT8mGJsf3VjTQPPBZli60mhUj9i3yHXSelgbNVZElaNt1eBP
DjA9fS54txX58UZiJYxNJWWIGMiXzD55CVIxKuB9m+4TbwY/ZiwszNrCtjK9qj6B
tH5DSpv0+sCf5GrnRaJefRCxRJyCmpWLwEkM+3SmY7m/F8i2/QwawIE0uFpAv8m2
XVLknCdiDx7ceJrJtPulYaJrezz9esS8AO1/Pn41CotfLJ2T4+cEcRrCp8BL7fWJ
cJKFsFOvAJ/rfYJjUXzemQjHxOoNiSBFpIKwrWfsKFjBiSlloANT4d2EEz6tbPMx
ah08N2WPBCd+gwcdMKFMzc4Jj/kIeNiFKLk9iMruSV3vDcOgEjzVxwiDwokNvhqP
v2IHXNHQ0nulaH9jRkT0f7N1SyOpURVSnm/6AMl+ggJIfk9bPiGQmsMNXt3uxhLS
UiIb6qYOI80TYI915qMwfwBR2aoqqHCOFgOL4/gHaOdwz7JMaa9I5K6MbY745tT8
oyJHRm7ke77ZpI9G4igy6bBmaZm4z0ClAXTawRozo7nHd829BSqn4pv2fQzCyQgk
fWHpTc+9HdRCML8E7lunAEEZDIFk2CvryzoJx6toWstjSnksYBJgi/OP5kGpNGj3
AE9lz7mOTf6A1DVxI/edwrhYgCEPOA5wMuSPStDFmg9HXZRzv1AMu/4Bgt5DXsFQ
ZcjBU1ldq3f7RgzSgBHRrAOnMMfnwqqIhzUEL760CHCmtm7QBGAdU3M5JOTdofNl
C4uxUtP6lGwUzqOCJJuuVHjNoRfu8IEDoWsS3Ft8+Gzh1E5EqvYMU1v46xOCddP1
Bl6ZT1wfSmblIUhmVmKNujLRG2j1/0uCEjO9+um3n9htr+oyQdHWTRjVuuFsxWtg
p2CjOk7kcxV3S+fLr9LRdyhVkx4ML8UTOzheKouuCzqcWq5AyeSrpIaw8YIX+gex
b8korsg/14gliXw+YXGnWfahtFXO7UvjrIsTfAylIyhGaLgJXTJ5h/B92mK+QEOr
e5MjXRxjQMklCu5oVJxt3ctXsSaQb1PbTpehRjX4QegdFrFGRMW6sEdj1EaHvoqs
zTHpFp9PN/XnSkQ5/8vHX35qkDfi3mHLXhv27tnUYqTz/20HZPWS+oHbAB+RxG8M
WNXom5Fv0bYTFzNQPY9abQY4eaM01SmOLTunyOuC2di6yY1fN+AVSWwbYNM0VJKQ
KhM42u03ORRQ/Cy2344NnUTNhU5vUISd4TBU1bF71rcrZmqxdeM8ulo3uNqW54vA
Ph6t6AoIcln6h7/vqBu7lAqszU/79bYag6WncPJH9jhNLH4piX+kAVMyI8LD0Bpa
ZAM/wwBgZ9D/HCGIO5maTSQlDhci58LSGazU5a6fAO81ufjSwvANQfBoBdEPyKae
0V6RZ25X2UVharIL5Jpejnh7myTNaWgrHhkPy1CaibGM+gVfnvsnU3YtixdENmfL
CjqcgxFeXOK86Az/u09h8RTk1pla7my6HNSSj3QD2ZsC6c3F5FKMXNumkryBlwZD
fI8tdtGMzYaFXi7A4OC0G1Bgxyh+wGmcfoq/Ybj4m01TpWs9uZmbFa5tbpHVJgge
UmN+J+tqtdm7OzAaq6zCvKnUwohTdPCt53vKZQCwECJDKNhT4ZVZ6XORy5uJJpLp
s5GP4gzp+Lxd12sW2ZyJWjoWgRQw5oxnaw2vY6AoRGoFG3m8VIddS3NWEsr/U3Z9
9P+7F0RppgPNIiXQ2B/wrQmgY3oSof68AncmdIYpMuvjizTZ3aFB8jWXkA6SVq2L
G+By7EckuNEW1KMFcflwHbDJ/9knk/JIuAn5xhSW5FRUaigyHH2zPg1BsMjcKtm6
w1hzL34YLSkAluyEig76IPSCZTHAu+AgiTZXuoMtbRnnId8gEOdpiEVcw7+IHeVR
8Hs635pF8MxZyRpzspL6xQ01ZE8lJAZu8Zpb5KDPsq17KCrT31udOVTH1kXTWLCU
3FxAJVn53L4OCC0NoHeAC9z5k5/vNxwo/cXUcRMD+eabLm4S/avTm5zuRSppR9rJ
EkTGblsHYvbtOICNvXX6RVIuKhsvg2ojaxi5QlUYlIq9E3S0jw1wdnVaN+2/Q+vn
56B09MZvC/L6JRogCvkG0FnPmR/dhOD4EVpRZnxJ9958MtGRcazzAYKcJp9JE4ym
ldrUSHVfg1u+g9/kpztBLSuuYm3f6rkEziTgO30vlbs14aWYBdJywHUS9N5D+sTD
9yZP3j8x7LjqzvuJrITDSfBUTwePVpzg2ItL9bcbGBxACmQtHmUzunO2hCvx2GLN
whZZYSoCorIMWnUcYIPiqOIUIQAcLU811o9pFN1W49auMynHL/osLqJGRMlkpYSp
ikZisbCGao3++ZrHadwSn/Q5M0UgLhsVfdYjrqO+ynhhL1HLEXYl0gJIRNYcXbtv
ATtVMUBD+xHsop2Oe6ZyHMSGsIfB+8LuEDzN9U5jnZxLamjDeDTLcQ0h7FqjP7QE
dradpminabwjrc47Rb3GoilpIgCyZDM7p8Ck5GPioco6H5R9M3gVr8MA4RuLQHAw
vr/vY/wfLbNqkGrM/qItPpZ27ANVrwMi6ezw1xYzHNXpnOx5m7LSIt+9HkXhHKDV
aci+oNoG8dZ/WoqmiKiGGXNz/uiO0RNa9Itx7Rm7+kuqB+dfao0esZRQ7cCRGwVR
JcUfhCWGX6puN0dDxqtZbzDGK/AnFezzb07rsArm3dJOP6qPVLpsh1M8Pxa8FWmJ
y0QM69SnXd60sMDxdsTVZaNa2Gfiow6eHZD/15OOQe1lGwtboAqSlO6IYm8xCqfP
W3hieX1jKv8j2juKXHeRtmXZiEfXg6XD0OwdUl+D7Rx/zDsjyq8ONKVVii8pgxq6
J0ZGH56HfWIgkFZAhphW0MAhsLzF5XVNzrT37oZ9Iiefihj5uZBTQmlxGLBlJMcq
X+WotuINrsPn28+btdaL959ROBYuLqbjlBZwnK37Dvlgyc+oQNyHIHslOpV9Fgq1
4a1HMmewrwD2pJDYCihaR3uMZPLKM13RkneE34XYHOhQmgt4nCjjrlTacXwie83S
I/zFyWSp6I//9pg2vs79IlBnIJ+gQwDdlNdApoKyPzqzA2ZNYaC2QB9lrSu2ejeP
ysPa5rKsAt+uYvHIJbb9g+fWs+lKnPmbfX5lyENt6cmIlbi3BzJjdsZhN+uBjUc+
F3AdUM4tcDQT0/7djC6vu8150w83/cu785nOlHWL8w+aeGkRBR5zKEojcMvAO5Jh
5ds956BrZIMN0XnUExlEVkf4vqOFm2LetMecLkHOUZccc5L6xlNNXzQpVafmlDyE
5vEOl91cwkJ4TYRyNvo9VRh1BkmkXgGT/moNlidxd7luOKa3wvjdSKCm1v5H/6rY
EXGPPGGnzGBlWgIE0oKrTYtfZLOx3Xw51IOI+NjHOqM4t2SbdaemjxiYgC+sqb3v
Bkqe1ITf0r4fVEVfhoP3exCvbqNbLtP/6JlDIp9qHJV7c51BZMCAFdM6FLyUnO1J
5GB6Yl8G7EBbRTS3gG+mljWqTFtdZg/5wDGhkeJbbEoblrINymXxNKsM/TO7yVps
gYyCRa44X+UVcnUGExS7AxAuiWzcaJBbTwD403Jl6/xck+PVMMwGpuKNUOe03pDx
7vp+YHQjyGRZ85U4JlkBkoIRsrWvsw0kMUZwhjUpF+Usx3Yq2WEOysCmKlO5J63+
9ir9hY+ROo+aRNXoB8l69fU6i7rqRPpRwM1pN+G+LDjjOzhuu3TXlyDu8MKpnmBG
39crPr/mna2d/WUDU9reiiwX7E2wZNC60VMDnQ4R9i7yn1tl+QwrNNx79ZSZhnFS
TugqLV0g1JXgJJu4Mn2lCP1wncf52tLYXJglZGKXDcK4GrNryJQs7d5aKqrWpsCk
GDxqrXaK2lc0Ha7F4e4MCXCj+yTMAJWQ0ejlfWs6aqxlVY+7sWQaDPUxmrc+wYQb
coKhRtF5+K2X7CBWGV9pnGNNeLR5t1LCsxvfZgeRtW4ovQ8yk63PzaUTvr/GQ91y
3mBXlL9My4xqF8NrZwv8o/iN3FdLNSllOO/WaZtJ4YbkQJuSnCf/WqIhXH0gJ5yn
uQ/9NoU4e1oNh5HRRvazxSt8a/f963RpkC7dIIvAukotZH2rsLnJ53hH7EChOYzX
aLJj9t64kPlYfRjdDKt5Efi5crBh3klPdO0Ril0BW2qk5sHkVL1Gwhod6yBUZClt
Y/t4fMOduyU3kbju/wakYe7kV5zpBlQ/P1oj8pV7V2hFxkMl0hfB+w5AD/cGppQI
tyawJl7SDAysJDnSmEIPTrJnF5AIDbi+sDJcN1wWOoy/Od06vmpF5zp0p5/KYysL
bbYbGsi7qx5m+I22/U3xni4vzmq5vSXVRbYXq94SGOcP2BMZMq3Gg6P13zrQLCIF
8QqJFIi57bzgePkigk7bAm+RrP5mh4syqFiXSDI7TNWMWiNsMIGlVUmnc3AH5MHX
r6xUoV5+7Ecqfet1h4J1mUBr06QPFlAjEdJXivGr1KV4+Zqrm2qbu4/NPcJ0HUFh
WdaICe7/wncptPSl5d1MRNuAkIhiPTMfUd3fZfqow7eFZfGCMXMCf2c3wCuQzSyV
fG+v0Ko0smMiIFnkZZOyzbLG+xHHBPOGYQaIJ56G+7BV80qoPMUMSG3PUW2jvgeu
UnJPY0PAufCw8vxZMFyl/gV7ebwppfuC5qrhycP2HM+rBY4b6D27twE8UqmSsw35
r5mLInBxtpca/Njq16OofpicCab4yWYM6M3ou3T+BmOOIl+G2vYuyURzn59+dh2u
eESyVOo6fw0KfS/dZ4fTagw1kEMPRZlFBKc6PP2DCAIvS+7aoT7gaNoN6n8heWdb
TISRc0ncU7Ndi3HdPMqflPHZNAiFs128iJMWbazwC8C2H+prtT6L+FzkJJ9qg+Ah
pwLUzrl50RA9HwBxF7qv3e4orBdI3+Vatm04GIwjV0OMEinHu/4+ix1VLqJhOUbT
/PUMiMBsLmfVRc44klOpbQo6eEFgNdg6WbXK5xEHGlHnSLEvrcVS6jwjZQ61BSxV
1jyaXUk+0wt4HXVz/UMwloslmdl+gXM5vFqifhUxIlet35ExTB96fyynWOSaCLVA
VryIU4VpNTvx+lcJB/r2U9YCWv5ZjqCZ22Klnm7igu6KXAP+8Gs4tlSgTiNEEySS
lgXi41+eqDxSyvNpvX/wk2i7c+rBtIkRoKUQxlkDdOcDXDb/uumzx0L6Ei4rsmDt
CRfYR45p+SYuasWQ4DqgakbGvXbgZ0NacNNWRB2hzbYAd9Mm32j+GUd+9lZxOQ+r
vyPQkgziO2qb3lJhKTcRD/OLoOH2bjm93pTx+aULgiv0YzPTxycIWjmuW+mKk1rX
b/0xYa+rAYF632+GtqbdOhDlyyz1OhVQ/Cp7GSkKS1VcHPRUOTctxnaKjBZvwZn4
HWlkfesC3Uz/IsK6SOw03bynf0T9VW5wyuMvBt3Za0I71621VoZGn/J8ebppp0mi
+G1LuHMGsJNvNN3RExMpvtT7EnUnmCdQaAsbSqxQJfsnnaNv8YyOzYUiWdUlSTqs
OuJgvy+Z83tcLZWQFr8jxC/h6ENBGm/0CZTs0bNqBi16DWi59ycTU7vcsNf6iMId
Fi1ohvX7zyIgZD81a8vGzY1l7MUlhZuY0W0qijx5hve+sP7pgp16y652HAyNAHk7
6fYyFv+9d70WilOuCqgZ/kj0ICr77U1yNGyZjk8p4maqP93xpx3N+1L0C8FtLfUS
D1ZmYamQdoyP+iU3Gme17V6qzkUM75xVupVh3ZdpoiAZ9QX97ZucNl2vvD66jqEP
6DTiYtBisIZTnk1ZNWJBpcsElRwTwEzx/CYVvr8DF6oUl+Xssm1HgNevBxTmqOzO
yIhho8NKsFQw6A8TkPpr8CfJ7T37w1RjHXyBUXFfy0VhXNu4rFeAOXb6yoLoyd71
uY2b4vhgvpzSnLGndjP0J91gEsu0tFi4dClH3+uQT6io2mdkUaW/miSlK6WB5H4J
02JCzxCmJHNnsNfvv+lT7CyqP0DAT5qJUZSdU1muRQRko4/raTBES+8m7hDuQBZ4
hVtnGfazLZqHuIODyJ/0kKHKaE4zc1cuRAE7Aq8+ALcSzJ4rjz4zf0+g6paMw1pb
b3IxDtLwqfU+bcBxIp44B/e01LPMtyqY4oXroYtA9q2kRLJC5bXg94aI7H6WCKMo
F+QyFOH8LczlOkwILJwexCsW9QUYzd0gJnPPDlPm6bo/RlH53GsTuxM00AfNAb3l
kjUG9atHsb9lnzhP1EArEODwFImhiDGhFOCdLtbCdEwapOebqeZX2+9fq/03IPDK
J5WHeHjLxG+rTW0eRWE/bvIrjArV7KBucXBKHuSkwadrNjydacgEOcIrqzrpDcAP
q+3HYP8CE06kh7pVU5SSYfMEzXojzyXDPp6zO7XJ5a8Qu57xjlJxmCuwo0UQ3OOa
WlJTeYxXZ0SBjpTWulpPjEUP5y1rwATRI8Tl3fryzLsDf0SCptKAWoRN44bh0G4s
7LjVPuZ3Ap30kCHshKdjpVC9lgmORveJU/XHJ+8qeiuGTknU41etIuPJQFtpF1S0
AkiEqobFXGywiZeb7Z+wRQozaWBcEHD6UQTAQhD72qtk0UChIT42C4lWTu7HAE15
9oi4pqw1nY+SGEy5qsva/82JB4B3eSt1/QYJc1mb2z6JiO3JzIOqjHgGFsdrFwzn
PgGmmi3kC0r7KCA3bhLMWvM+vb0Jzvew5Db07g7bmBSw3QYRZiy608heV4vxX8cI
vSbfz3VuuWzw80sazUk5HV1WZpwCqdVQ4TuHqbOEk7skRPF69blTECIIipiPV1sd
ljyWMVMEaT5viIgFyC3G1ZJvboceRfdQH6A5bsEiFOjM3o8U2OKYaGZjxrvkfuAM
v8VOAe9xcwAeo07/gz9Afz7v6yd6oOaamYm0hA92rnfT7LIxyNqJp70hze5AFWfG
E/c+8qSchkU398zw464skoqMsy1q3XfzXxyEIEKk5QwvpfBVxNV1zxg0yHbp7nif
ilfofffdATUyTbTwebMYryMQ1K3uZylrjTDLXQHWkWmuI2HerlrsDgLDT5lfixAC
IvfoCqNBdR819Dj0mms0yJ2OJpDdAgBa/syQswCTgQeHmprB2TgHhWhbH4p9s54P
tsxhVTNv8NtPk/ID8S6uDTWwWzr/wQEohn7OAV/rL4yaQsJ4aqq9U2RciA+VBsIm
/F4eUzJ7KGL3ze2/aUYQ8f9KzROZB/0qp9njy2BtYDlVhPUgjIf6iypC6wVVHS0K
SZkfvC6PSG4OmkWCkkewkrAT1lkPYaE6vn3kP8h/JC9dMI/PSk07ZgC2JeATjOMV
IJoiGS7naMShHKHcKf4QHiCjWKh2vs3PNFa/CkZPUJ6NJ/7DQLygndF+/9cQhvQh
gOKq50OGRsbePkG1mUQxvUqnOuydStVyjC8MEP+uQYPP3PQBB9jdF2YNPqBu7hy5
EOMsT71Ps6RHKHXCmqQ+eUysCxUYcx/BO0jFZgx3YLZt4MkbeC7UTcQ5tnyCV2wi
cikbvIWzwFYW9Cf7WLkftYKUCDstGazv8/MItA2WePLUftpGy/Viq+xyPOSwkybd
QLl29/2IBuqEzbwXZflnIjGkd4MNnMv0uXVRoqhav9hL9AVAXTJAU4umcvJLuZ5f
hXfJXMc3psdaQkSKyQaCClvzawxbRdSqaw+SwMVFjdmnt6Jwhso03QYdOwEqueuN
KSNjBF/Yqa+skybPDxEETPeSJxdDiwFFoCsfKq2BfyXg0cA/n7Xefnu09RtAJ4L1
tc/7WR8lqox0dC3efbE9imXTKo5rvncA21aRurUYedWRWEkE5jD3W9mr7YbQXJ45
3BDJKiSjL4jdIH6Nwp1PscYGDAP4mfUxqA1iO7Lp1WwHXJpqyMuAYU8bd6fp3R/V
qEbhVVc0B54GoF4muYsJvphLiOysRqzcwIgWpisDT01NRq6c31n4fcW5BaeMgRTR
t8p+QYFvUP2q3AFT/AMXEVELSh1AZdMIUiDngOIWsbbNIf5AszJx+mxogHmGlqoA
m/XNpAQT1PEW0soVFnSjDUdHX4C1uX1l4QHPu/tCCz0nMxvDzgoCu9AH3Jb2wWrn
0wSMHqjjssgW/tv58XD2WfjaQx8f5nme5+2IXj09kCWxPK8m9yfGrA53oaXOya+Q
fWJS6OuCxQD91EWBCoyBtug0TUJ8ERRyHCFzl0X6jFKMUFcgdYRaMwQ+doImSeR8
JVCkvsLIDbuGpfLCmB2hScQvAoNgqFkbhyJgaMT+Cgw/sBlEyk1rSmOrRb2xGuKn
Nc/sSBMpnfIZxvWbJlvypJCOSN+qCF1HEOP/njj/ohdy0s7/wKFuNcMZGMIMXawv
TCGkkeeC6MbyJGY475p2SVNWMl+WB7RtE9NSj70CVntPTS2wZUEI7AXkswvQRZS+
iloE3fFsrTwq31UA8Buou1zvRKf6SQrx36oAI96QS/S8ZM1aTq/DX2PrdedlwCEW
SrBn1lJcST2AAIJcKCFEFJh6HPAvo4v6dIkHFrziFT4Vk/Jz4A4WZTrt6mvW/c2x
TAlt621ZhgHcfmdH0P6BEgMdb6+gaqSnWA9ErMbLGQ4ax/uFPK8c1a24L8wl73k2
J4HBCsbk+1CnMwgCDVG3Za1PaGuPO6oOn8OnWkWTjP8nRkeo/TJ44/R3P6iIHFD1
jG65s9A257iaUtvMkC4THkvE7DGm/iJWANr5tb1B57bzmszph23tOms8jFLcNXMU
jVcsbnE8AjXJtre3qm48wDpQagvl0vt8nPxCcKekLPM=
`protect END_PROTECTED
