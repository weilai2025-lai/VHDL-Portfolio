`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9yA7UyCREoudY8lDKkLb6BJB1Yh2vJPPNvs3N6dz/7vKCmL3dKCYszW6TVRLs1A
skY0xQjw0UYoowyxdTm+Df4ENKK3ST4I5kfThmvDgOSSNutk/+TBj0wfsZDFrHEr
ltMG+Im8M6LTfSJRsuQWMFTw2bL5/nx/pI5hs8lJdXSOahdy6pwAGlJsr+LY/x2i
5ONYe1iVHQa/GOCM1o64wVraaph5ezoEWeEiDGNQvawiKsWzX8UUl+BiZOxkp0GY
NZBcQtezFGEnwwXB9aQQap4c8Gg5WpwXB2OpBF2QoDRQMp8DR2wVC9UQFfy+7ue5
xFZvYPWzwBBqN7fGeG0EVWobo8zPhg6SavoILJ8T9fT09V6ACh6EvOT1lKc+9i8D
MEP7ceuT7NCYFwrNtHoGshXDU6GzQxY28UNjQsYW9Yo8nbhvrchA7gl3br9dBJS3
fW4QRacQWHfg4PYuX+AA4I43Ile7anavqPMgn/XP/0Roa9aRXJ+BZ3fRl1cH0DdX
ahJz72hKUHdODH0+JKwJXVhjEsIACdkVrJJAD3M3f1I30EALSZpQniQT89umwTiF
PpksG71IuEtbLg5h4spQcVal3BR4/gnxolg1AsIyqp4NduhxGwODLCyjIi/Y0Vk7
AZgUOlY47LwUivIEb+CLKid+zerG7AAhkCXXTCD8xgvOLCbGDbRvawgbzeN/4mPt
UqUzB8CTsm/4vIUL0yUAeHOm+x2bL33PuIi0qiyGVEp16cHrdHv/4XVO655KmFR0
0y2E/IAJ0c1SAxICpbKOtONGlUt4frPHr8NkTlpSrM0DYz8K1aXR+TYYfkSQhHsd
Vztqsmoy4P3xGZ0Q3481gPgzAetZM7uEQ//TZ7rbiZ6Z1VLFT7cEnU6xkgriSrx4
EjZsyqsuuFMpM7d/pxAV2nLjGeFKUFTQdLvOK8VTcTMRTATzraA9YUXLeu5NA2NW
1zW2Qd5rBBRicAMxrdBONcBNgMgI0eAwJX40D8EpBzSiloeWJ4Z0dGTtvqTeNltx
9AZRcHioGNFGUVJAM631HAieHPj34CtbmchXw+cmJB/6So53UZtTNbg91UgqVj7Z
EEzhs5ZYSUoJqULZSefYr5JRJYPDvXH4xn2LWNG2739v1DuJCdD/fx58Gr85fnEH
GsQgdfxtCZKGdeHwGV+POaKsBJKa+mSdQrh56WP5IzcGQQIGE1f2b4Yxi42Md1X3
XPUg3eNc5LWvyU7uBfkuY6z+amcrVZpPlHiIJvJWbX5Oi/WxgRdKYFFC3zBgeKR2
+Gx51l7aPC03+rg6WC5zPLy7O+HS2LKCt8Whrjd/4m3MG43qvpIoCQX/9Fllhhvl
Am2XGSSTJycLTvdQyy+SrXTyKDwNdBTUPU31n95aXv9QXxW9B17xGYvLYy8tLvbD
g5oQK8cMoLMUXM8SyJZhzW4Tulj9L3lIv++ww2UHqz1SVnmXYJb+4Vc5Ubli/OG/
H0r395UOjKgPAWyx1yoEFp6DBko988lssEE+lRpN7hv8b3wJ2YAUcBXTA6dCQkH+
sWD8W+qWXOQWXCb015qTQ0U71FQKqVD1ZlQ8AFBeA8+fAHr7XNdplSsc/QjqgSfB
gZHWIRDBer0mPB3GkhoAx1MtGbxDfQSu3N2CO1cCD9cOh9KzyDGQz9NYzUasqJ5G
c7PlY7DHMTKJUVez1D+I24OjLIm4y1EZfvs0k2bgiG+vMCRDN0g9CLjfffZfEmcz
1DLQPL+5oHbZlXqiOiWAv6fyt76/rmozAvlrcGhzA9vZO4ZDJ+m5e+9YWXkroghh
kYU8TmTN5rox+wbM/sLM3Ab7ExHuR+o0XDE/hIAp+DtQiFrpQ5rZy9JA5tf5NeXj
8zJqcPzj05pEbrN7c8LW4G4MZNrvZ75rQSF5UM1ye23HY2U9OVdv2pWzPxNZ5rAv
l1qGZHD37WtjEQJGOQAiPWIPfuFIC/xcDDfX+j2XCqMcf7pDJRzCnL7m2gKguRvY
egj4hV9EWdDS+9gAq3DlCl5XxANtOas34dO0a5mVaXKTG6npE6hYvWJgsoW8TvUd
Yq3rCZYC+TFOYf1K/2dCIsQdW2kb2WhBNi0vgo63mYq2GH07MvQEiMJG8UK6q1L7
M6w1yRoMgz43hpLRN+sQBuOlGfDk+AJa/QQ3Wc0JWKewRZZWmKchl63GMTYcr3UN
nHF15sBGrQc7WcvvCfVKs/m7RREBtIgnpjhT5vDgLe44T7JLnyzPXFPHt/Mu4Cfw
P+9sknJLBju0MVUT0E1dnXDhV8ynkMSJPAnuavg5659UzkiERwWdOGWNZRtG2q8x
wxNDvRZ+yLpMcmUcVXNGbvGhICDEZixy6Ibe+kAM6CYaX+B0UfVyIW3EvgJRj7EU
`protect END_PROTECTED
