`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+BoSn85655VOK1AXXosdaJhFUjy+rcpSygXD1o0Q91J6RyOdgWsuvlj/sYh2k4A
hpj26SOKTP8eNNdJi4DdGoAt1TSs0nQX84Aj0cgGzSynC6jc2gnpOJtvN2TlPgxg
kj1LNik+oouhASNDKrGhVYF9TPSafMjC5g1fFwJlPIgDuueWqyLjA+gj9w2I4AFq
2cPCe4YMBfZHF+u0QFCcQ7eVfPcjYqx83W6ALfS2APEsilbDjfraUCXpNmkcMwRI
TdTwoe+xNuWya+J1AmAThv76aPwF11DxsutLRoRMl6ftkBU8V4M4Bvs1qSsbX5K4
A0nsZJff4sAT++gKgz9iWad8C3/DFhZClm5a+rS11+qb820iVRk+BNy9oD9VxTlH
plyFVrZeX8pvBrjSKfSdEtarHN577TkEHFpnNV/9ZiEXjq4X5Gv7wDjJVPicpWPu
HfJY3lXDxp2D1qfSMUgN1N1S8w0/85larujR7Tco0TdgTspAlZ5GUtILi2ez96IK
5GQ6lx6gYszZ+PbUOdhTn8C2cdJKQMXLeYMegTijiTb27KW895I29/7waH0DkZAB
n2rtZOGC5E/iuHWBOVEGqLWGAJ994bzbPp/vyNioXi46xuZ9PW9gvFq7Ig+JaJip
cTDi1UtVyAwZHDV6H8q6WecyfI9D5JVwPIWyNCtStPJ/u3OyHP6plGGewCNrTDzX
M+vi1F21VK2voLkYixJqHn/tXFYUxyOAaTYtGT1bZw4=
`protect END_PROTECTED
