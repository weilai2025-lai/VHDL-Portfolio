`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1WGZxy6AoAXbVcfgRg2eL+8/gdIF1LXE58uP5frciKw47pBG7AEzmNDo+WXrb2jl
UkMWAEbvHp06NrQ6sD/oWV+L7iZnCGFW7UItFFZitjLdMgyeIwq0fxlzSawCZ2II
ylf73BU28a6S657WP3Os3/myQrd1SjenteipQtz7jg9TkF/rNypta/wObhlspPfw
7j5Kxo5fCvJGXoVR/D4LGC6eXOnCaw71ZqUOd8knOuuAefOe3PgtMdDKuJM/eopU
7fcO2Shg+rpM3nN7V6zk4UOpEnw435UWd5A45FJjt7+myFPYIZLUy88czKcX5kVz
/tRZVoEotc+/62BQ8N4ZqNCl5tbZLAt6hqQEnbtAZ7Yif+nPqaWyvuPqtAgw2qci
o7Axr0re63imxJCQxhB2ox7/VyHvq6F/nvCxHb9mjKYI0xPw3YVrmFfIfqK+T5mJ
Y73zgQ3Hy6SG5xmh9d3NOY7OCLfDkaPRSmv0ENjXlQ30Jetyjxan/Aly3jR9QVbO
jptJi5GkUvTXwSFmWovQzP3hyeot33Lc/KXT27OF+sMRGY7SK+KDRJV3RA+6rviv
lRm8it99Wos+IG1Utyz4C8QDnKOODIxvnXM7PLYGRHqe06Vd7U9AgElv/dfFfvWV
U563qyjPHeZYik8aUmBf2f4rC5lwzCoUzXCY6s0YWn8cG5671W+3kndlt5xgArmk
4sUf/H4mEZJ6oe1U8/v3F0ThLKN71nHRUEXzAWXZzDWaKo0wUYN4N4V7Akpvbz5a
MJr4eNEnZLrB1W8SRMqkAM+EAV4Sy1x0cSTXriyWNEctNGDmOok2qZRosBU0YcdU
LZbl905N8MMweEIaBWUSxjUjxA0ky2dlgx0px2sWBj/r78EyLxoPwrbRDvfEjtiE
nnplsU4xqddMCWDjxNgT5i7s5qHbuySPnlkRM6Kls7KUD/yqK4CSwikWelVJF/Y7
bcLsZcLTaEaSbZgx6VZY22gEwlf7wVb7YQ2cljyPD9Mw3c7EXvCqzyzorVRZ5i1s
FNKpSNNZCvQLeKjgkLllXofiaF4dRx42CpPlo1mKAsCaNc9lbOaF3hYY58J7+fs1
KEs2EpD/T7RieyEvCZakPYk5+cjyu+ix0Mksg6H4b9xXsPgzdgbNSWhNetPsZUe2
YFlJQhKY3qzmFD5XOIIcFW+pthJVwDnOoGUb1Bt7kljsjRuY+BwdQ2R7oEts52s3
DbxlS0RmQT8FSESwKmXUKV10So6v4cCbzrxaLmHmJW8O9RijNmz5+2F6PoGX1+7d
3zuDU8EPZnkglrpBZHCsp+ZmdCSvI7i0VX1xk98AAi9TH/MphRIVwynzHkzWN3iW
aMfM1+1ECi1EaRoAYzVrWRLijWhZmnxSK0CVJgJRhJJXXdpyq9Aj5IiB+YBbBQEu
RlD0erBBRbngHhMTiiq8CuyhEQIRQMCevPCvXPjwq7WDBTZPLAPqCVkCFohip8m5
2R5x+nYLmw1cI4gq5l0P2urmGwaihfVDlP8dmLvT0sEeg1V6ZpD9eIf45gN/MhD0
0OlAZVi9xsvcf+yBGDAdSoxAzF4C7R+zqf3Uk0Z8r2Tgd+xNO/nWx3ZbxXjTetw6
uCyoVrCyTIpDN2vSz8gSijkLj1Mog/zjESAXPksnUf3lUFIqg8EwXhr90Uhj+9Xy
/ISizqfrJUALJiOBTuK18Ob246PqdFMIRVj7hVb+qivhjm2XYml3rgYPpyldMSsg
8wCQ2XjMSbXxS3+2g9nG0HCdke8NFIbqP4td5udESuzTRjK1l1IgGl0CXqjOcFOS
kvOkTc5xSjaK0ebPwegEFFVjzDKqecIrFPu9dk9R2ZJ6OHo5SRubLs9k/4ogC8KQ
FxXqbvDg++sVH6zNcEKoLRe4xG9X7qMWIo/lvlQn9oghDUQ5g75HW4WfKKsY5Gn0
cIRQB2TrkHho2+QDiX5tV9RsMf9QXolGnkuv9d5RPuqSGAXA1ofux8+tSRFrQsiK
mwZoQM+/waDRwz0/ny4PlgF3+6TD+A7qMxCUKisdkEhjISy38qIAkbP1SdQZ41Z3
+XnZ54ekvBn3Rx62rMhjk6Tx0hmvGwBNBZ/sVWXMPBDhOqv5ekL3NCe47llMKlQy
BAljY4uaY3Vp6WqDK7DPqiXt96XHGHJwTpq46PSgXOhm/VW0jBDUvdsEk/aTiHFL
VdUbWQJ3fy2cLThxhhzooBYptj6AImzipIkmgGxIr1cPlg2fVBgCuTIXpcsS9xVt
mVLgLHRWPvZffRwTQHCNKqKXNJu0rHu/qvwYM3OR2xn7T7pM6Xq9zsyRBmwrm36q
9U+CJgWCzWO8SnAriUujns/8e32p6Lb2c6jjriY7ymorlyxOGjnL7rBTA3qqDbbP
NQKMx++Dwh2/3iVYdEP1cCBapovCFrK6TS+d4rGnmeC9Mpx4q35lPnaGou7MMLKV
zpIJLcb1x0RirC4KCH4TAXKXv1UFVj9mANnM4Pjjo4LFfEXNKwwoK5guGZMsRlLs
GHqAzhQHKCp+dvHMkY6xY8/0d3dht24o/u2QwM8HLyxITJ+cHSyClmoQYCviL5BO
uhpiE+0oq/BwJRs3GwiNk2bQhidTQY+LVFDRJhNZzC2ZT7PHkqaESVakRBMC0gwh
LkGQXHNQAxYZWSLSfWlq1sKk1EEEwTNksBQYJYcfWoYKZ8/lhFRKCjj7dnnkHb0G
2jOj4NsqUqkQkM1pLhmwjILXch7vmeVQOg0ysntzwTl+94U2dpcmTE+Vv1PHUAqG
ApYQ/6J0Z+AoCj/x8chDIc7qzfd3pau0KGa214lH+XN1PwVAAvMqdUYQLM2YlVzp
ycbqtS6qMvQG7Dcq+ZUkJpoYwPypEVI8ER6JbhLWHu3TzMpDguec2hFJCzZdeHWr
mGjud6PdmGEaSY3CyAcyIZZNRQMvAzmmoV7T9I9984aQ6nQ9ikWGMAJWWpba5N23
b18q0HT33K8g7Nn73wyiaQ94K3NGwsHlDsEmM4M6FuaZmTfJL8WvMdgZ1u3VSENV
ya2yp/VNA9+VWaLXPOeqzT+8aSM9CPnNY8xD/zJgrcFHNkUIBSyFjWuLsd6xgMAP
+cuPwf8LlqJtLXMdn1R8ONBST0BhqRfWGojk5sVtLA2ccdvwW4P3XXYDY6H4KlVc
TZb+Qs7LULPL9k+4rxbUQx1dGaCbQ/WQyO+mYtwn+dpVZ8B4fK/d30p9cYWf8ZFb
FVjXBKnHXkyDRbmpwk9/BXNlm0Ff3SAKCL2yrkv4sxPqKzQ8kt6e5+8qRc0HpwVc
NGDN72cWE9pvExx5jR38bfkboRAG1PvU3lLtROJaOw3y/dqyahxPm1s1WYLl76Vz
/4xiLESO7dcFhh2jv5FoXLZYp2Q4uJ65m/YS0qE3r/OJr13SIWt4PsYLfF+EjpXq
4yWrYDSnLycMVT91yWZCzMQ3GeD6uja3vtQhrVBYK1aSnGLv/9QzvdIl0/mGTAH5
qfm6k1oqcPMnBanjvbj0vjVXu3txh3vBCMGIyvqguePM46s5QnE/t/VT5fxjRb2S
AYi8F8y/aOGXg+cEUFY/djQaM1CvAmMg55e5gIHBqmpILeQa9pvfoS8Pa0THQ7q4
7QRv9uic7JVyfc3lLD1QL0yQp4pOydD/KL7HuuvoC3FYkIFeMzKMmLWho4xEPwXO
8JXfwultZhPZ5QKsU81BMtv4Avp2S27wW4prJmbCTz+qW3Uy/+uHBfmW2wnYOW99
+1mPAs+ceeQ9VDZJNX2np9/h6bZTYK0PVvcIh+PLTiQxlO1XnuEgYhhiquOsZ12g
1/cRKFaze6VrKqBneqIW4aNq+FzlpAdVV2BuMDVK/EzEofbOqtlMzywIg+Q9nA8q
lUwteamsW9RIh93BtdagOrRwQVbOjGXSGPwG/nOojRKFs5YioWteG1ocpnlZkT2e
GkpxBWi1SfYgCntiDt8beYInnz0d9bhAN0sYA1I1OumxT5N2otYMDvly8iA91GEG
YFK4gtEZHFQ2NuQT7/K9G/8bNcEhXecEru1zQe3rJUQ=
`protect END_PROTECTED
