`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PijjVJVWgy2RAz2WGlMaQIazaxE4R0z0W3RU/aDxiUB7TuNbgtoV/FWwiXdpYPeY
YmYFqoPPyctb3Rpt8yfbtmVkd7So+LPWNqm1YSF0RGKySCVQE0Df9yKEJwZ7CVjf
rQPQKJ8qGsK2KdJcAaWDfRslybqS4vMgmT+9mdY+MQvVOAS6mLNaMiZjwJNWwOEX
1OvXwf4H9HgZOprgTCBw+AUFGF0zmnJvLmM6cbC0LK60ZlvU2YHuiCn7mR5YYdzf
ySPgkpDD8MN0rgERkcoohudtWwN6c9Sleje+K91Zrc53fBTsF6L/X+V7RlKgLF7O
t/+CKe0FSD/ProJ+l07XR04bfldk/m0OUc/WVzhLP++RqU12/67j92BSkr0xaoTQ
7rGUQuK7wbcgrNTVsEEw7ohFPN7m8cKKja7IhQ1mbRIKJef7qWoEtr/hkyh1kR/x
c006b7JzidGKarsclSLwm9wn3CzljaiUFwn7g0seezoIOM+xd33R5XMSArimR9RH
vIodSAKXUSXNcn6jb6c5oSJEicvUhbxQ2PuI5KZRSCmvkKMybKQIGQOeredgXEUr
9H7JIeQchs9YaMJcpE6CybRPAhk0uuvH5Zm8PCvAv1lKUMSlAZwCnPXeGrOqRglG
nwhaVO5FnbLxJ7VTWJeP8LPJOZ6TkO0L6fLpdkMzIGlXgfh44F4EibECHeiVUE0c
E+qMCygkGLl/JYhVsxw54X4qxe/hoqyFsBmJ8DKRIwyowWFgvIU4lg3x7bEtdZ26
cB3phu7RSQ8SBk8yjCPdrxLE39MF+8YOR8CbvfJC99gI/d4KeRTpyKKnRzEqgBEk
Un/xAFIjcZEBJ5+qtBS/Xw==
`protect END_PROTECTED
