`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0LCgqWfDw5K2nLpSWhPD5ZKR9mY8ypVrYNzCIdTlDvPRGosAWE/X46j8vnEmut5
2cmJR9LrwXM2I+MqEa46YiIR0qLZvKHOzrS5AnB5mmg2il/9e1Wo/Y5JXnTC8Gqs
kX0fySz5hCAp4gNrCnlwQ+0L1YrHabMgmaWduvsc08rjZ79SJoODHMQ69Kps6fcY
DtgvDYp+3CRr4ugbdOa4qMyX8CRXZNZL98rGz2ob87l6XNZmpjoeedpMsS/1B3Dq
U02qkKF8P56Ar63P0dxo51RIcS6fpzw0J/HMuMfbA16m8/932adiHpbnWGfrpDy1
xBVGhu5y0DQN4sUfJwVQ6kfZaaEJjLeb74vjziQpfnPFz5Aqq12jKk91uvb7x0aY
N6Nu4E4TFU57zKTga/klIw8B/eOrJmdQjx/zLRNZnGJKz4nljBtR75KfEPMy3CrE
bmwsuxzf+e1chgVzgkWiLUqyA8xAQrcWvtBv1oou9oHGVcprQqP7J+0SIg2QfVok
`protect END_PROTECTED
