`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nEvAVzXrOnTiXaVH+dMgKBqnfef08TUA90TXXFbrwy1PmQCV7IuMafsDSW2E4NC
ZjhKfhN6lgyykw/jjRqE9V0b65k0Gg8NX+bxY/FfUqHEl7ipJMmkhlxGWf/dkUgo
E5TZao7UtlVXk7IwJSOYH1FxjqFzs1zaKI+vemqXHNfgIWN+x6jNT3jFxJ9t1+cN
wuAf3kCobdUu+kAXjHV+Y/32l2LBx0tuoH/2nI16q3edVyaToYZQgMCwToRmQ8fX
djs6hotZTDlDiWmTNqWSAlQe6Lq3TQQucT8sO3JbOPvzLiYjP39DgEtSkHgefKVU
+4IpUobnEi3LtYUrle9Jf1Oyzc/plRsrILJ1VCMMhYR7r9ueoISsSl/+OE1m+MFE
D9c0tbeUBsleryIefq516gw5PGeopZVCgEduo016deH7eKRQ8J9f2r/1HSdAkiVq
E/ekeUPm4qDNIqT/X+OGKgdyAco7zRAOPEVz76QV4Zqf9mv9KRrz4uxoEgBmad5V
0/iZxgSG9BqP84FD2oMUKb0vB9lW0+uQQXgsvOxoDRcXBubrxczrs7aa2iVYwHdZ
D9HUuSVv6LiQyckxw1+goODR5N9m3hq/gTsq+d0qTbLQn+QijcoMB5pauvJ9Kxh9
zj/r++MIXBFpQGmqig0lX8ObvtcvcjrI9FEip3uBalmNq0Y9Up4TMcFcrh5J+vJS
4xUN3kK+utMbSpseOusoKIALmKYJbi6fC8s//q0HJ2wOEev2wrW43NxZQ+rWFCvl
9JYQ/Zlygu7DRvzj+Tt+YLOGC1qRZURcv3V+q4FeUGXK8QR/j4M+RLEIAPH4f56e
w28ZwO7iDfUpjqhYiDcM2UhgECCY+Yg61g0Iv+SRP9I8a4vml4+kXJhdNrBv67b7
IP2IHbAxpRN1xMSwEIn36poLEVpfBi2gtaDoeCGPajw=
`protect END_PROTECTED
