`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lnrdbQl8zGM5La32vywZiDE+o03SLW2JUBgqV2notBaWjP0Wc3GI/Ifo87xVCJ1c
h1PikPJ7QWtDIhO57Z7+8p4tiy34CrKrwAYjBL4waDPpaJMGIZzRQFhq8bFVujyd
/jDIIjaguEGleQUgJq05a2aO3XSbKmAG+x2Mv2LmVyMjPJvsNcQXadH5CuDBPWQl
Hz9Wa4+m59jPr2dFVXMzbLw5fA2q79VJtsczBvsitqlZBoq2DNEAvb6WhPw6BVKL
nfGRTJa/isRxjnpYnkG1wY+snWctGpnmLC9RnrQnxm6JFs5rbY3J/gb+dA3PF67x
hHWQcAtzX4QsFoX+bUITyXSBLyrTDMEjjjqrYWQUpDY6qXw7b0XEsH0Hs9jIAmVA
1oasSIdl4JHvSnNEz4hAg3GiOeAXbVsUY8ykW4GUHwnA8xXS24D4CXkFWNBIP3ty
eFx7uF5GPDCQK2vm4ZVGfYCQU7vY+Y7tGV9abGnnSJeAuKdyAL2cRIa5YMuWvNQa
nHVKeX/nGGxqZRiq2c5oaRt/PCR0ix15VGop85ALa1O56+Wc36RbwE8Ui8h5bNMt
Ro5FiHmD8hsOBZInrPFtWAAlWfKEWwxXjXIFEIrmdD7S3qhI0KxBxg0yGQGF4lJ6
niEsdOx3g4tP8q0a3GvLv55xtMj/pdfUSZ0I+sDgupHlQdr757VmosKayEZy7yHr
Vkh0dd43sU+EhEJS4g1KfGzu4sAqvffnUyfy5HExmMoHLGVucTLbH0Uh2m9O2ytc
acGoxmERFKJkEiaKL16LRg18VyDT9fgBROllnsZtCPMJuXAP9FBDcMRlNJtCNHjp
54Y5mkfQ8wX6wEufDawr1eYpLKMXW/ouuRDPq6dP4sQ4V77+8D7gPC4/OyN5Tz9s
Eolw5Xaz0GaNp4sn1QzwJBSv+t7/SOFFHuELj2fwKNA68bFsAh0F+MlouHrdAhqj
IPMPSSlzz0JPPDhYRRVhwH2LwS3m7nJqSiDDroesfGIUonLccHk9KhiTcUTueNq1
RA47MlDfGl6gVrDlKpoeOSDakMSLrIvdf6ii2cz91HEN/KOjR85X+99Gkh4CJZgB
C952W4634W/yFxAxms6mIOPDodM44+8U4mPb55h3Hun25k4qK1e09r0t4WGJkdyw
gziYRcCwWnaD1KAwBz5RlkOG/YROr1RZEpmVZBYrIr4pOjWHHRckfN6bG4eN8SOp
sBJ+fueoZwcfbOaSsGTHlLdnALm6DIYw6k9lOX4N7uODvwrLMESyVYvyFVTzl6ub
XqWbTLdGTYjqLVpvJZbNIu/YEagBVL0w4bg7AyK6UwIeuM/sTM5Llb7S9i3drIf0
K241vJcl/D/7Ezo9WSgWIcFlvhTDhtpmf6b5pGFW2wfyQ8OOKdbDT7hPKr7DOj1p
3FjAL1FZpNy7qIlZs1DqlYr0FTP+pNdfDkBbDTmfnrKJOJ1qtfewC5ULPUngPG6L
vJqW6GlRnt58hkiSleXfav5vY55YtHZEHwmLB5vgneilFLBkmQYqKmAUUzPwFgw9
btWRwPbuG4qRJBmUAU8ldx8qTysiXnuGbTi0jdIHC9Xd5CX3WiQf1LAz2ZXbdmgc
03q/iXNSWGY02jxHEuZbPgCaohDfDREd+1T9I9Oju3SKEF6pePwP2JV6yAYKjwbK
9fk6TXY4CSWUTuJM+kiV/14uMd8UCWlhz94UC+QJ4Uvdt7yYOgBRmWz6GEONmlfJ
KfjRXxjPvKK0ip1J8Hls4F1vbByl8aYE617ohvxnFXy0o+PKrRaa5tJsyBUBXsd+
7AQdqOS0VuI4ISz7UWiw4xEgKa8evj+2QVLoJtIEVblp1cxl7Vm42S7+p0WYkijE
2y+JmTvsGxhBVERbJZjH5aDxtMJI05z2We2fdL39nbPx/hOs6vbcdclHcwpSWZkZ
VEd93wZqlkcpGXbR7ZdcWwpwWoyUKxueKUwA1DYPR3nrpzHAm4ps/r3Ah/7NnEC8
+DBJTbYNLojtiNDiXRUG30DUfjAJ8XcUTT/vdguH5ROBjLjB19nmuw2Gu2f2h3po
iF90DaGxzmrVqxPs1tCMLMi6UHdBKsHOWzfeX7PsxXq9zOyRWhLGQxd3ng2ZE8I9
khxKZXzl8rWwd/bn/bDOMrw88piAoVS3Ak9yof2zBns+Y5kmLdW2MFnHaYB8ZR6M
vXcucPRBiDQ55jLWDaqqPUxa0qVEWpbX2b0G0r8pHmx3NuSCTjERnwf3CNQhURXO
k6HYLWWx20A3Ck6tSbTv/0xPDaDJhWRO8mEwJp/vTxthGjyK26cPowdup30U/Cky
fPE1HHFoyFQJfmEQkSHWUyOFYBWhhhdTNrlcWEHbVJ/X7ruo8ySDrhwdJq8imyN2
BcLxQMwHHbg3iIPnjp643/Pzn4fAZsg8j+T+m6THKgYDUCxLeKa89X49+VNRhW3x
D3dWdve+LaL2GGps5RWT4B5drNRisZPSsO+IYesKTvKAsv+vLfySyL9K9CeJoNCh
YMi9tqwEuXe5TVRCCcfgHLhGvcN2P2dUlb3Nd1WVJUtEfImAwwYIjujFUVYzxxo9
NTyvUgPRAFCy41cQ/StvHwlTEnuhsjxGaOK29ng2W/lvsBjgg6wpbI150g+cxgEq
SeUomwr+B6AcbTaT46LRxGWxRXCHe3GNxcWg65ZGJS/Ovgd8UC4oX5c1GtiyBzVl
RntMseiAhh+UGSXS34Lq3b8hPG60LHHyMRZ6VrYZhNfdqUttrrCVDeXYbz953+LU
5WZndKunb2TY8Ht2MnnngEOByW+oY+aSFJ5ULCF0oq99DEXi4SC35HcdNJek4RJN
5Dn60r9oIwbTqFAHd9XWEhydnxgAFH2O5Eb44KNfZEWdes/E13xBaMN1x1B1ltpl
b7svHY9M8ES3H1xlQwJrP8Vv8ezd7+sDtwE8OImRVPcGNzB2AbVmXZMpyNzjnDNz
F7Cj5e66AFrWdf72ZGRYr5tCbkukEf8buNWIJEQpPxk20nhdYgxKSGKy0IM9rhiK
/+6sAj1wlIQjMw0obOzMvo+trm7TViBOz3CefCXjelfyWCuHewrDTJsQNXb40qpb
jQZ7BZw/mfgrrX82UPoddup3NH5+eSXHJR+sZLl80SuNnik25EYN3w+n5swJAsYa
8kJhyq3raJBINxivKsXDIS6T9LvXcmpJqHx379tIo70nEaa8Xvo6yevboHbOdVwp
UDd6evkI7gqmcb/u7ALxsSmDD02b61r2GIa74bBH5fZqrQ9d3jJwGU5mN8mH7ECY
1peOPcKa+K2h22goaB6pgKQYrlXWz6F/gIEPhzz6VyHUPKWzyuoEtet67HBIzcZS
5tRgwrHnrzpZkYwIEHBaa3Grq9NHuB/hDhM7J7khjG/pv/5JTvsWa7wUF9vbef4X
iQlG1js4zT+hReNO0qXkHK1xpEjE8KCB20Mg/QCqgfz05mZecJZM+6sRmTghA5rE
CneSzGVI9nOAoYjxTddy5Z520SIMGmS0TRwanGVTKJ5MYUGEJN+oen8AV8fkQHtV
JW+bLYzQQoJFtRXUQLLRlDXU9vXBvSERjvBcCdIMFpP4we4rEerrv0ghmizANwHF
zmm3dze/8iU+1KEMoG3UREOMkXreyLERJV+IMlY5Y8gX54Pcjx+GuocaCIcNXaY1
oP9u5fqhlvu4r3wpuucSJI+/QMeLvC8V8hUYsOwEkkwSeH/Usn3MVKk0MXzgu4eR
23h6Vk2ogrdmES0a9aWfo/5T+oUksqQZCURoYBqaCrVJppdR+UdUfYJzWuAs1/jY
zjH+ViU/yRdRadqssLtTnB+wdEbfXTry+rfNbbniSJtcJLOdI0spZ+Hh3/PGr52I
6jLNGX0nfFD3xUrA2r+ANVQkVcpaJVXqTxj1LH1YMgbEkVKUdL1tcO2Fh4O9zCqm
TXoM2epXXpCgNJmvkQDLCb84jvSixkwiOV0F+qfIYAFRFv3hiyEi1Fo+y0r/WRcW
Qysw0NSKdgi65L/4JsdIJbwqv/yFpIbXd75gsJMPduuI3dJ5iSgj3nx6x+y1CfnV
R1j+OzfB/alVqV6k1lSBxeHK0NU5fo6XMmj94KSS795u87CCQI4w5WKDyQoQLe0s
WwRAhdim8hRi8pyW9J69W4WV4egHIJTqcY7rtZtL+mXD9yZ7GS+P9Db/k5g6VB0J
MRYy3PMO6dlgMQQ/sSzTt0w47NdWSut0N34n4YYTxVM5BgdNPifDELrGpBmP/+hV
dudQwcEcYHm/OORWL2nOSrObymqyOoiv+oGKwIQjJ+SK/+5RpvLzMAB+FgDUpBXR
jB7wyAicHlDtGSuYpOcDiJ5OXExeARzsyq3OSa06kU6z25h1nDG8S+wb92HZaSza
2mIR4esoDTV2wMMAW7v+z4wedEdg31kfHCL+g5MDE+FH6WPHMvIc3H/65hbW3VDA
grHztt14WDvwoWGZk1+xcbAnTX0RIrc7r2eC9lPKHX0HAw8Fyi7UpATeGVOJkQEl
IAl5U2tfjjLP29JxSS53Or1BOWF9FwACoborTNyNqs+7Xpk1ppf1QeO9ilPsCeeF
nQvJp3LqcnO3BGgwp0D6/SKFLHcnn+MtOX3oSh0MP3Q4ZyyYZWdllkzUMnVmV+Eq
`protect END_PROTECTED
