`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q2eyC9+ss8hqouk/zwiZgHCcOeJoOklz55N67YuTO42Y26m0xH/ifvu/6tDapfi2
NbHL4KHaYhQFdft0/brVJFFi3I586VCGq/HJWUXJY3FPeGgsaq0mjFhKck/zo/im
2v0r3bIVloVIPG0ZABT+ztLWGrJDt5jDcqzbClCm8LJc+pTbqU2604rdXhl33Lt6
`protect END_PROTECTED
