`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrK81ntM/mvxQ+8yG44z37/qV5Y9hozG23KR5LmXqjPhEgnAxF5W9nmOI0Wx2FKc
dgsN5sD+9OqW2ZihpiLM3n7caUhOJR7PIQRQ9+iRzUmsUTy/mLyNHpx+r1ZLoLr8
H0R/B33hpjpcx4lrY4QUlB9YwSxO6+OmZEhAR1pya4BbQ/UvrDD+hs9hIHXOUJS7
LvhwpL+FbzgEMKs55Rlzz2dNEz3LlzBZdHqEsgjm4NlNPVLtgdU/4IjxGQ3wi4BY
L+NyOBmCyco/SFKAvByRyLMiNG7OJE+7yz605zpNMOqvyAs1g3uYDv5N3wyqxbq3
24LqeaJhCStPBJ9yuo8rkJheI8RL4ohwzpvBlfWkO6vlGXXVhMvhV32fBtnGqUlH
do2I/y5ImwGXt+Ke+S4zF37mmSRo842Ev+jXkELtp6hWqdHOP58l+3e+zjjUbs1K
9ewJFcvmWh6/pfIshtBY2wTnmuOIu9lmwtgTIjbuPIF7uAT+c6W13YtAGklEyNmc
Yvd/RAGNOUOS1TSj9gOMttEoARquZvnG/I21WMcDWLeKuWfP/CurTaUAh8NN+zQu
U4IIBYc6Ov4KPCXnE3O0ZIBT3ewoGR3nBTM5gwI/KN1FRZrHzLcxybEpN5/FmO80
tEsH0ce8MSy5BqZNWYrKf6u9b5gP3qyim4lf7p6U4IHH6VqFBxqkkXdgY2R7bSG/
OMtnpwbX2TICUIaYzW1f/RAW1I+8n3NX0YalsZodduWp3Q7MtGRRz7z+jOqnKZlo
1SRVvyV7Cb92iVBlUetQp8zbSqHNo6znKmorMrAOJGHft23uieyZYjT+BjmnFDa+
qVL6iL6SaWVJEYNYPciEzOvcG8J7wxsSmWQ5PRQegTdC/pbJ19Jsou7aeusOFe5u
l/DWnuz7dGJ55O/GQWQjw92ssziNazFZ09gdPnGpqa3uJ0hb8J8IDuAYnHRNXjcC
nZZhxu0ImTTKojzGc3vY5hJ/cLi64bk3s8ZwRLg2rGKW/Jh9BaXYS+M8txoYg6BM
kX0jPbp3NCt/7GEMTIS0K7juwFffuNqdYtpAfA1j3zp7zxrqWEsLEMEQcc6GwYy0
9evvyuKMhlSuY75tlVxaasgq761CVITror6Bs0PmBtlmBN8IBeKVSOhdZBPF87nn
DYbJIkcxmxHuZGM8AtqFWgLCFoTwX+kP4x9kOq3CeC/iFzj17lCd1KX9XStHrWLd
PMiL5dK5zuOIZqNvVMG/lrsQOqFkEri1df5BdLT5QKZSWErLBMpG+eVtjoWLM9+s
UCqr7iqlPqiasUs0wiQPN0lHww1T/x/rC5S3SysOInzEpSj2q2R22/XuEZVYR1JN
1vWY/UW+vp+NvyuUCS5zdWHNWUMy0MpBvPabIBpESpqjFwCJT0fwyba2gEWlDAo2
hB10C2JPJISRC+rvjgchVlY95TCohHLwv2TqCteA3gCIN5TAkNveD0GiHW2UUHxP
eAJ9lFnGJmYE7n8qnPDttd1e5/UmxPEwW9T3FFcda3fZZnmjBt2y+4h8N9itgbzv
1qX1NSLSu3z6EeFEbGcR0a70ilXCUXNGrD+Um9x2FOhd0nJCOFgzbNxNXFpR2sAL
cPg1p9HdO6T979vWZDEABuafQM/6pglkC+6xJkWy4wlcsUdw/MWIgfrojMgYcbVU
bZc9UGcVXyh05eJqZny5O2S+aWx5vz5kWCFN5HwkxneRD35K5N7evDjyqfd8tWlz
dh63/KXywaPpfp0olSSaznxm0B6M0IeCzk0B067mA6LJqJ8YnYaLNPVzNclLXSXY
ElT7zAvGRqWa1ZRzWuiLCsMHdR98rW3w12hnrXGZ7S3rDXF/Y0PalrgzejM26vRg
A+SooOht8oKOAEURQXuH+mauwWvXQ0ewp1QZbx1QYl9Q36sxujyoJUKmPkaSACP7
UcRVeCFGA9XxNtf0uWSiK3jF1ZwD6D4z+prz3/p0nq0vYpZp/0520TQQfeIi+6gg
l25kWglu1ylj2Y9FNWk+Jq/tIAuXeUZUE6QwXXpmIo56FjkZNxI2W26iWcGn6UXA
W/PODSURCdhsGSkqWXnCYwiNKwyG6DauoTspnxG3MvIGrIrGZ7koBcDGUVke8pHR
0mMvISdcuHcm5RmWNCTzBP2MEeum3mdGceUHCBYUy6toXXqOSmU3mYeWWzRSupYU
f7FnN4V9RcezU2XHoUXZphosfwb0UY4+3FFbWSXO+FD53bjrEJg6NCw2pcpGOgMO
MXNpJoyYxJXsdB70kDFdMg5t4gEa4ZK8crMzG1Vr6T184Yg9IeqPmSb62Uoi7Gph
3AZk4w08OLf7xCgED03+9W+aE/8bDssnSHKl45iV612zLtVAu1CFA5kE+oMg4ZRM
rSyPhQYmjeV3+BxsC7Ba7yVrC427Y1isXt3BbYjbiNG7/7pz1mesiTJbvxeVUsUW
xGxamNEvdPjZ2jePaQygjAmmFFN3f2uTckedieR/NuU4QuGmhP9RUoFc4VSrgsdO
PN8NzUmhK46XQ3eb6HkIGehOR710og9243j7ALKLCG0NW4HU80sjQ1OAqmhxobSw
FiZVwrWgQmXWaHwYiG8El9Tkm0nE9KLoSUlUJKvQEA+N9ADatj1Rs47tfViaK2nE
lnf8MRkM2NX2cj8MqoXsko4HzRtD3MYjts/eq3BcxpkpRU0+pbE27ehl3TdSBHPw
wFMP/JvYk9R9D4y4uH1eTLISdPMbjHep1kRYQLCIIKsgjbVUzh46h5ywejFJUqEE
HRwbkEbo4XNp9AhUEyeGnRkXrCbR7mdSEdVgpguSbTHCQp8JFBzM1Mo/FdCnvAIi
Gqj/DvNEsPL+Q8MjLHXv3GheucBdM2CoB2D0oHe1W7cv+M9zlgu9fVgLEsSrcPM/
AWKMmfIKlJzA0EgX1vXy9Zwt3l9sAsu0UH27MDBEZr4US/Z7p+hdTIRGI9/yEbJ5
FiddpT7rWrvwVpo8J4DF4549HXVJEkJgp3CZrIMYSjVu/ZyAxH/8VyoaaD9AVQjC
ntSXprAroQ8ezbSpmVHGxmVA2jmAIehCi3qAPWq+O04mro+9Vjz63qsQOLV1aLRW
A9Xs/nysF6BznxvIhzbyDE65IJbBOF5LFJIwXNbdxnc6ETbPJDTo7OQhzFBpQ/5x
ddslNEuaDajDLJleQHwZ84O4XfzmzYSTG0Qgrvg6CZksbObg/TSSZ/udauB1GWCZ
OdCqnwXb0tF33ghGJ6Tr/tgNNoq4607H2TC3X4cEXUKrRP5IAGfnpTsCrV9ukRmr
uuWGeSSDMnVx+zSBiU78fWvTWLNHAAkTrBfRqVzCpXXCj+XCi+jQyJNZ2vHWAXaA
JPZbNSN/c5ibxx1cepfxDubm2bxr5EycTxbhDq6E1ZuUCLwXeePefvuiA/8l5Fk6
KVDVDYMnS7v8TfcI9/wvOzN+a9cyYdEZ+BkpMZnmwZt/7jieoyC2y7hnzu9lCqww
D3SBUhWBXGRoqxRJwlcnYFRFd45xeaySejpxg/6WJg/AgkYNuJJG0ONSywDyDDk4
KKPewBCy9Fu8CYpOGBZgOAJYkxGvgAzzDFu2XXr5S//g6WhwDvkkHpjj9mrNYjt6
JEQZwNYTzd7JMngJ6KbyS1ej/ncVLR5h/HtXsa5cbVx6y94qlwCr/TUtcmTDKqDt
D93nnWfa9GWv6o4XEqe4w8J2OzaSnx86CHD0ZM8FhAERTuZqnBm9FLDycHj3XcIk
/NGhAtJgqSKGpsFdc6DMEDqXsZ0X8OUI+Bw2d3zYKlE415jC3v1oK2IP7CC3pR9W
f+xzML7Nk8VjFlfrP2PVvgXpZatqECnzTn3TufqRkiHbyupktYey3i9gHZN+WalG
Xli0wtTWWY/AO9j7WYtw1Isnsl7V/TYs+0ndCaDtk9XoskAsXlptiOMLAfrt+nOg
+lTZlBbwGP0oF0Oh9g/Rqw4/LR48DTQ2P38672pyLu4rnAiMlEPKAW+YbKDh2yfa
wKbAnc6gqpohD2oXABC/qQ39r6dBd72aT8Nk6gDoHtb2RgPfu3ko5vVvCqWiu4hM
mSlnOL2nH1baTfRbu1gjWmkIoPxhSYz4ODYugBXQaUHxdXmEiWCbC51xb0gKBu24
mB5djDGKm3pMafzc2tCu8hJLHhHrDtEcb3h40tsHA3/Fz7e4kgRcy6Zq+e7o5j3s
WOIOzEk10f96ZmrLKeCP/Y+NNBLrxWA2g5GsfT/AQeXNY6ufLgoGdSPzy1nn0qMn
YbVU5fLA3O42A4mbqKFp+yeAM1MBKlolSRnZ5CtWHVoj2cOmvfAK6ODH+S3+E67E
0R66M+aUAUPNXJ3SKWLtDnin92XEsSZKlLO6yI+8tEwSlP722wtlDUrXOA1QJR99
r8VNA8Wv94zNBk9zeWO7tK218tf+09tSU3oB+tFxaqeM5EvtIdLRSl9+7WH0INLm
PGO4YPaOEI5dzVB3+Xmc95U5gv9WA4Gq/6eIAG5WXD/OVRLBS+OOH7lF27HkInDL
qytD31RCuPQsWdYcPnXIrGYuPwzXQvUorJm8dXSVoO79ydVRWStqvQSrqNQpcBfE
7YDU47iL6xkzu84Bvbx9x65CdmeIGCtVWQrTXgKEnobs4d/zS9XtEH/c/9548m3c
/74bnMJkfTmB2a1IX0JCxOgxlsUK+9hi2wVdXq80twIQwqdP4yMvPZSOqCYLB3t5
G4umU3gk5M9+YmdeKtKZfJH+ZaQbuZ5OKK1RUEzcg60cb/WZbUwoyZnIN3P1SfmH
9xIHlQbUZQ4HwfeHINO0OCt0CEHP8ct5KhjxoafmDAjIQTVt4a9E751cdZXY6NLc
mxVVoUF26ZCf18YQcjcS4TO83KRjBPKYICRIhOk/YRDCb108YK0E2xGnARqUpt5l
gQiQSQLEfSi068p3G6D+xdnCGt6by7XRx/y7xGTy3lJX96x/XpkjwinVxWGS+Ymk
84JFQ2VAc6Tc00hOHhYBHFB1jxYatfK9XfG7SHU9Vr8RDkBLS54IbUFkh+AWvMD6
eA7ezBhIoEipwsPHh26+AmQrENFzq6Vew5yH/OPxCdlwpzu4ZmYCp7+aK95bMoY1
aHdzNvoTi60URpzG1ayjJ0w9G3l8rzR1k45QMpKLkp0G5B9VlSwes62Adol67/fq
CKeA0UklJSVkkiD7BnzE/1oo3cn2iqBOzaoNc31zZv2Yx4OND0Eprs4eNxDIwiUp
sOqvgxju/1q58g1WA5QJoASTQLNKYPgWLsaGu2kAkiwNlvHAC0ZsqVuS1TG9pEAJ
OBW2GGlJpzvZarWpPGTEh21fFiY8eMPzWBYTZMizEimW9sU8AocFXFuHUtm/zjFD
i53ax7EnNwDYCAKImeAYuO9Wl2SEJWJ6Q8+i7GEa5Qy03Kp3KY5dQhZeHgUEtFNv
uLk16kjU+WybBDu5/t1Hg7kXzkoDWe7jSXpCeM7VSjo7gycnnd8KEoFlJR6QflMo
vwajsqM33wpqEzLrggefa9B8IoW6FN3rHbnQLQbp8TVpSbV3FYWvc1LBWEbthTFR
MBDUnzlN0PXquWFjKQWtYrr/Tcb6wmmDkpLjEDTgQ13j/02sirs2VxSTsIQoTtqG
mQ26gh4SNIkfBqlsap0VBAV63n2rVVLTpePPNjKkZq4BOLfSgoUi8qCw3mRJbvRd
MSiMTFS6m/006Zp5dF12o9TORW55zUMrPpQhfxj5+Y9XwnJcdvu08XJ049OD7kC+
ZAb0W0MH24GtoalxO2/U/oG/ETsDv/o/OLXgZa4Tb5CTDCYonsBQFoQaaIkIzgOB
JJr61YON8An0Kfxm2JBo6xusMXa2oBXag8N44tA1h+Uc5oCYBMkICk38SnLrql7Y
d8Hb0xkD957lEnqeqAAz9QBuGnFTYFSaMd2e0+ekeCfJEC+s7isCYn006IHZTcfB
lV82cfExQXN9KzS7UcKzkXmVnmTeypAkmNJB0xXcV54tPStPOmq9jxqsRlMjT9/4
e7Mdoyf/N2JuUxvNxKndzwTFsO4mjFcFQM0oh8Jl8IahiSxhCfaHvmXR878LhN87
ViyGbHXz8NB4yBSdXjT5BwE4E0yIcOioxOhr47NeELh5ss/s4C+/2mGFLxIgwhRi
igd7di3LrBluUgWZnzm91zqBJn/EQbjNVG9qVH4UNmIREDW14XoF8Fo4lEML9Dz1
Xaeqp0HnoAiLT0EBjpZ47PTeHMy0wOKrRp5c6DQHfhoRsD9kXHmYomkDJHrWRt2M
MbplmjiY6Ibh0UDLZAhs+hCo+w6XyewOwTGmw2Mr4zuYobSjnOJ8SzNr8mOURwzb
W0VCRHIPwlpAOcrPnc56Rr3wovRyUmSeg035rcYW7OfLGJesfPdPxb4JfAtoVXEl
fVtRaH8+sV7ReYBNFgciXiiLhPPcT5lMbC9y+WUGFbAj3X5eIlI+8/hoykfDxdI/
LxMr6PudShYFiWY21Dv6uqWgfQhOpArejRjMUVkTSgi41zeCLII3blq8awrc6fEY
aWvWLsR1/gF5BZgKfp6q4dOfB1ZkJ0I7aMfLfqOxkM6oPeiQP0mYs8REi3zIrfcs
s0KqZ0NgFbD32BLiULAMzDPwLJK67MTGa1GkGm/67Cp9m1Ky0JAnVQO4DC/AzxtH
DLrZBKzk7eo4ETltXzXDtwG3ke4MEri4PDpqWdf+A6WmIklNN25pwSX4NNzC0lm6
61vnshOBB8Wkb+SzQi1++tjAy/oAsqGt8i3pCkXq9syaxrkjZh5+xMU/xCNCJ4eR
gjMvWVXOTMPRa2UVVy4aEr+iQ5C0wfxHhWG7DG53gkQHQmmjVfA/msIuHf6RbeN8
61tBHi6laCHI++Obyrg7bHDJdW1jZlOIa+LAuhbxlXKich7b76tK3HC5OrCqEEW9
kkXqya2id69fd95chSW0tCy3d2VEBT6vkV0aHlvZxr7VCaQuqk5fzCO2aoFno0/S
rZUu3vyF4136yeTTEj5EVVGTnYJ55vkvNcqrRkTauQxiqPtCZRJc6vrutRbE/MwD
ld2b3UYckyJ8IJ/ZkbRSXC0986D3ea7x3HLJ4VmoyRdA14p0zUBiKlv1BNFYlaZ+
+hmwsDh5mNDDomzWyDQvxvqD9daHl3EGpq86wg2pTb8Y9JPZL/UIjM7HMdv7VWBd
l6F/6r8KGvgOE+vE4Cx1GrFFu8++NoFctXLWUbTiJRsxDovsH1vgZ/BWn1ZTWmC+
Yr/xpe1bp6u8sVVLGCDasm75U7mCaGeWo6en8qI/fbwqiDYqInfEt4mPjnry6G9l
2S+hqdqDZ8FtNUA9cbLPn3xwRZI60YlF95PUz32vjLNCDSlu76o7N9v7VWp2mSU4
M0WJORKdewgfV7YDCsdNh/EpKvZgUzsaiHujeunb1Y8yPMqg5YCsJaFhQ/hS/LKa
YfJ8SYH7E8JvDO0195scyeFQ7WSV0wdSRB79uMxi0dYU9CmgNj/49guRnJSvgyoJ
XD7vIYPHldro0QBf7/7fgTavl13x3UC+N/NYWrFbFgxVAvQGoNVolS1OXBDqUzi5
cieVf8Qfg72FHyW5v1wBZ+3YuaY2MtmLCEZz4+GBJ0XQKZgF56m0K9XzAoNz3C5M
roZRrtINUm9u/RnXK0S5+tCYGzeg2D0zNRirwZdOs5CAn/jVgtnGxHm0koRP2vCb
cajNI2Q8bE6zYnp/Ly0/1EWhAekNPRj3S18uBtzgfRVisTKRm427HhVH0ijkuGCq
8TMeh6QEPPI4enuU8GF8WM3lOuVu9ZKrOJsRMJgMyC+beT7QNPTHo92Q2MzV20Mv
ClPNNb/j1UQb9PAiGIvoeOsSqM/nQlHNN0JY4sO+fpOku4RRU7t8C/g3uQ3nK7uB
P/xh70JAWdkIlBFksaTv6XX/NWn7zGVs4qfTDlPp9aSHU5XIv4xXrVTZRmYQRlf+
Hfr13SE+FVmtp+z4qBZVPfKuaWKALNU+9QZEOszYE2R0em9MihHtOSd07mTQ1cgm
3hYTm7ObJhsV4M7OeGJDWqQ/ZFI3gU5Fv+VWVaZfvIf8K11oRIH3cWoAwnq4DoDn
/CEMiwgzMOVvHm+RmhQhwaCmTSdbrQ4b6c499OwCmPJdgmhwdifK0t7r17tEjK6k
pBv4N+PKSa7ED9z2TROYxvvkNBXHeoPYwzGNBC7Cv1U3bXEv900knjy4yLV9y46J
Qi3y2WR9PY4+NuVxYw9bG73fkILE2yNOGfJ381K0rbpfrZ9o6KkgCguqB87nTPg0
0Kgn+RUWy2JOiCynfVRcnq7P536gcGQCKIzgYU9wkws6VHJpRUKG/BpFe9GpYLQy
GBELIKtStgSN+NjeSbayLWY9sIrsPKKG3TtKVIbPXz+osW6hMfAWYP4h0pv5lyZJ
M8sUAmZc6YLXaE/F/R2T5MDH9KxCj9TOP+/LtgLmF3hP6y0crTc8HCRdlRkLanRj
HttURO0E0wGFy6y3YsPGJpAX2FHpJpd3LszYaUOmFji06zj/9oENova8Kfk9GZCo
QtoYZUlgMdpBWlRACk/byaanWhvIlecj1FdGB7+VYQPgCwZCETi273Rs+wzw/xrg
E7DfCZbUcdFKmwKyu0Ms51/ne071PU3Bq37jZXcSSL8UtYx0FnV7alu1C+Gc99mw
0KOL8FRfhQZxGIJ9Dy8AtEAOcwBxdYD63Te7rfhNAWgmsividltIeshfvpvNxsbJ
FLokdVsagehRyfQzodC9tDJABQ+FTnAB2FjHdFWeysD/zEFW48eDtOQnEvOtSOWe
VqGWsZJ+KG4aASp2246jTj9qwf4mqABL/BqZupjPSBO0ODnrqaefAN+f6Qb7vOnr
FI/AA0rrzpwUe92mEX9PHPUvEh95rHYVhZ2EAMOiimKHm7GOdIN0JHnkk+OTciO7
AiVJRnBZ94iyRCQZQcmB5iuK2xU+1qbDX1M3nDUtitxQnKkys9s1BkcXG7HTicd1
JshD1EYaTwiuiz61ZNukU1www1uBWQwRhRcBqX4slAGmV8q3+2+RX4MW8dDIowJX
SdoxEzF4lcDgcmK0gkk0IP/zSeOcKlKBrD+dV87szJiAYg7frI2RjaEYQhCm9aG7
/hmX1Gmqxfvn/Mrb6WlNNpLBViuMGIFa97B3HXSG69jvoFfpEI8ak1OMwgi649SI
EpEC9LmsEhnqwUzUHb5LQOCyVmOu/ykzMQwprmhASDGs67+IdLnaBKoVZIBYB4Xi
c2wBaeR2bA36OL78Wc7Fe20GFXZDOZl9j00BCo0dDincJIRoNCB8XRFiKHI9+vY/
aainBgmyN/sC5WKGXDTZ9TK3OgRvCRwkBOXCb5JS2tVdLJWA2x6QctY4Yal8QPBT
/P0T6jRsvV3+4L3vEizY/MESJT6M3diQeIAFGmEJ3GfxxKUmq1dh5jfiTN+rGOb8
zfMoCEeD+8TEE1g7HLdM8oqKNC0X90m8vB5say8k3aIU2cOfen/smiVpss9NvVGr
etbvGoQn8NFLI1qJojoW77e0SHBB0iKtRxd4eetDC8jvKQxlc0ORxZ4Dt467kcul
BHkwV2UlnbznWrY2FgUO6FFV+hfrcIjF2jiJma97JD95U78CUc/hPzZBSOJXl20I
47v0iNYGLB/K9ylH0D1QykjY4xmcqg9t9k4u1m04VYdlgjWjBeVgX4/IUC1fAwq8
7HnvceMZPqdeYyfYlSEANpZl/13llkCl0IMIxhU15qOqkMDZpbn5dVY/SFTmoakd
X1QXtrLwy3S0/O27scPO/rSxQ040B9iFJ7Z/Do5VWJdULal6Y7QYkwztllZfvppY
EeT8T7s5iw5FFvewVAKQBegdbM6uoCnvqB5OCgi5KPE8wI4emn4uCW4bIbb8qpFc
s7YDdmbFAY05igacYSzSnkXlzuSL/0qczZed/yieOReFRfuJbqQONYZ+5e2ysfUf
/kA56I6mUqafutkGqqQliKQNybeTF66P4EJgb90Qj0jXiqcAUh6UViYI4jlG47rK
3hhFDgbRVZ2iiwiV85czCZ3rA5SfNEoCg8uO5gpaTYYEYoTiTi9wtPdKPgbMKySr
fA0kt0SBdd4X0wBKKQErei6V689OlMASzkyPw7ODYkMNJowJuzrHYVecJlbgFcVf
UCAO5BtGNXCa0BIpwxGCvlUw8kDF47vJGkc+8N69x3mJD7hNxMVqS+cLsxW+jWFn
yTSx2Q65GT3YkSV2rrrstRX5nDYLajknE8EOUThiWzuw7D8kOeo0dJE7NegCRHCi
ZJcscsTrMv9zFWhgYM+x3IWpNr+aihNDySfteyiXHVxiS5CQ6+cXxrFt6A/4Oall
qyDPWwjJq4XSFhUBi9jaRdBj1nwjSXAeUr2nhZ9mlwVUjS3KaS0jrR7NzBmesKj/
HMR4tX/LNXqs27KjzndB/wmVjPoYXLlRGXtcMPexo683HtlsNAY2KniemLiWg5ML
YgD8rfZovujK/JrMzYAQaMI01odY5Q2HTzBms75Dfp9YxraKFETrBCpf/8MFhhR5
0BXxZFtRta6922GeglsdHXRTBZIeUweZMfDLclhek211gqkIskBEev8SrOIqvSYM
+Qp0CYv9sVq3+D1B+DqV40N27VnhbpKx/VUXmC3iWOtMSwNG2sL9F297ImSDtaP0
KPTygSpwpLj/7eDaKVTlydoLH9/tSU6muIycjxOwPLl1doQf/LqF3KcksmFHLqU4
MNlnPULa6FNyGE9Z5V/lq5Wq6SuxLZ3FT3GuwTA95LXYGOANRHcFU0TBzrSyyE9o
Ru3ZSyLY4FwpA+hH8hWGacyc04ihr6jXnbWEqiikuoZtY4fXNXvSHrJzoOrzKLcE
+K913Qcb2jTRGtum1NnVMiYKXGIVbIYceVuh+1B5GIN/XJcwRlVxpC7yIAXQIKfB
+xJ124aHpcpqzXyQlwq3006w3vD3yH1+7fnjrfFLc7dwggNrKyzC3+vqfpvBVxhm
0rtBkWSKVpr0CGBVysCNQB8Ov6QGgyFU54TpFozVUi905mTRTD7U8qk9oNntk77A
Pmzx65vIMR5ytoWP/KWiqMOyz42DTDLOAGCK6neV/sZRPsIGGHPcmupe7KtnvJDe
vNFh8dRzzg/qmzDqYvzqoNFZTgO4jxdRk0xBtilTSoFbjBbkuaRno6B2pdlV3PM7
MDTWSUSMkBflLFAYEiQRE307ZRHnJHTMssT4mqh4m44bblN6Cd+i1T5OhkLXtTf3
NP/YpYfDsX+wZ9AeVwLrNzptBJw+sPFy6W+NdBvmLz/euigq1peQVD/k/kLIz8Aw
O8zTTeuufah9MHvruJVwfqKaM2/U1Face28ru+FUCkGCBX/0EGKmt7lVLmSaSCbf
SmhCirn9NOgeRp8felupYjamJEKs6DALWjpxHxtES//8mqsOzXpnIXOyRscaU1C7
sa06UgJObjyAJ/6hFBQBR49mob1GgcjL3aXafSGtBjPk8mxVWs4xt7PxwtpE5xJc
iDjMo+O46txkQpmU45azI6UGnr7FI+SPgYP3SHP8kWgrK5AO1jRcZzxn5JPXwagy
OwVXDcxNpGXm2ed15z0YJqyjYt5hrTMm0km/5VuLiqGqZvR/VfBBWe9vmSY65aQ0
zNu2Q3+2tYmb6kC3+Aju7u1L0Ji/BWBV8Sc3dTSnNDcb/05OoG12ELrkGJ8XAXHL
Kc2rOnqlBudBJtNcj4P7/vdgxAQ3qI0zQuPH41YCv/uLwpLgGSGgiLzBZ71TKqRl
wssJiQXfaztJvJ/wM2YErGElF751zn2vnLb9zCx60FOXk8PzlSwsqSCW7BAQxFFK
eQUpqLGselNkx3QMouD5G6gI2CsXg/+29ZMrafBwSPUoN7EgMU39R7q8W/oRSoF8
rac+PUbjF7VDmuPMZqJud3Zo5JF98C5WuH95tUU/pR/AxMqtaDCx++ekbLiU9RQq
Pk8hLiCTHXgzHSAYMO5vdLP/SUDc2Qb4RZtDobO+1Jt5MicMMWVs+TgNB7TGzvyu
i+3grHRAv93NxzRqXUO7EGlFWeeTJGQcnyIzTNVABzoa0/ilY0Pde7ZX+XKbG0DF
RO88HLC+UlAx79YSLA7XYZXcghoCjHzAPN8MiSS/sVi/Y6KrOGV17cFILxhYsUpr
CK+T6NS5UszmXXenplIYS6mlFndeo2IUeRj2sYkfl81tevarWqb6ee6f4JjJhw1L
pnjfe70+qu+7MnJHhSREATnyPxLlv++nrv09PiRyy1z0/pRucuYx5lSdZeHtQJXT
EV5RRoNqQCwMhCxPxW9HbLOb/aKnr04IWeg1ys7a/bNMd/u2OjHP8lyLQ+iOszTn
kcR1vnBA5zxCnmwwigftqeXGO9wC5WbSNVidyxKMpAxEQ26l6n55SqsZ0Z4fOUXq
+92p/B2YsGtxSakV88KLVm2naM7waIrJ+o0zyt3KIxD8OxvKLrhBTMQJ+NvXuhp3
QYR7+zHkiu0k0Znr24nTOVhvUtYtAwUJcd4BH1isUECyj1OtjcsXvoU1gybDfakZ
pOKPFp+o7MCPl/zZUJUcWf5KPe1XWtIU6gYEnjpOLx/dQsW2V/h2KEPvveVP/pKY
STIiDlbmQMz9p/g9KWzlIA==
`protect END_PROTECTED
