`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DtCU6WgjbYJqNAYvhmCDy2V2sXn91aR/40Uenyc4qXvAx0+R4Tsb7Aksrt43D8Sn
wzIr3FU7tC7msNRr2E/ija2HQd6zZ1LEHxMmuC0+X9fI0If8PwKFzWjGoNDuFfNa
Sbx4xOIA0JVS6GGvKqSPPm5JZ7gSRjyyKNZOqobGCmMkyns9Gmc7PJ3ULd3J/2Ae
76uYmUOrqFk1oMkfIW2e6KIqY+5HC4Wnlv/FphfBILwsna2neIZKTnz1PcrM36Qz
JjxJRUrBnVT7BFiU7szgrNL77lwCWKTNN3Fz5mNbGiLCFt4mkAWo+WiEruxoGGO1
HfJA6qA8REpw2kzIW3+T043iBFFch/azmWyJVkzQkcl/ooslxujlbRJY6boIo3vU
QFP6oqbvFyRTeDUUbzZu2hA1jFECbtw+7y1IJRHbyDSQ4TCoW1JdjeGlBrY/ssF4
+Dl6HVrdkdnjS1GhTg8OibLTobjSt2sFPe5ipihCylDM0/gynUsTW6P9xCQH/VXx
`protect END_PROTECTED
