`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLzyHWnA9zt5jg1Rp+DD23D+HoktCZpq3/0sqIMPRG17n8p9kaz1NsBvtoQEkyW4
CfyIsNCJGTMzFsiKEnEY+fCiyteRL12gSRTCBxIOrhHQf5JKMxf+NzgdQtOr0VfN
uMn31XprdDnaszZUCNyN1QzCUre9JbTIhr0yelcjLkEnYLOleBrD1OaDx7OAq0rv
1kPz2hU7Aj/O3WA7JOcgMwPBEqlfjSiI5iNiE+2UbaTJ+y+njP+zBGd+PHrieCNs
S2pbIuyk6Vdx1RZ2I9NxCWXErfxgv4QxavQEwJ8Rz1WtN5vXe3djoc7z1mA15yCo
2LXEcZ62IQX6SyqxKbsE10ChQO0bP79dtr0Bs7FbyCMf+GEQ2wY8cVXL7mf9VWBT
vEjUvosYtIXzx5xB85Uvv9o9a5Hkah7zTFQwRy0ANXO8ZjCuwHNRwA/RmRekaghl
rHYheZpRZnio/29Os/l9Uo3QzhbMNpN5UCiZ7EWzE1kfhLEt0/xvKJN6Oc7tNvLP
5z5Vmo9/bKkxvGKICsiGscRhseu3tCPMrzbKZj0QdJ6M4tNUwFn2aLY2uiT4r1wK
PfgMxOI4nSNFYQh3ag3b05v5AVRrPE+s7z/qCTWcTgSWCK2RRbpn6X+Q4t+aKkcn
J7oysE4s7/C+Jr3fpg3MOT0rSz6p0FRCl/h8y0zBub6mJty9zxK8SynnWsw0Nrqt
PNUdiSOO1AKngcDsEnStrChz46i6uAZMWitBraU4paCDP4Oq13MS+Pz3Gsvmhsbj
YaG31zbfWe3LrluyIXNHtE72AXXVEVE+0YH401A5SIzKy61+ykIL3Ot8NNwvcAaW
g3ccq8gHx5omypXqZqNZ297BSoH4SAHdEi3fFVr9YxEBpcAnR/5shywhgxFEMpDf
4XpyT7M5CQcQ3WdB2gw/7kt+FaGsWlg6ihmgk+hXjVCC600k3BwTiPTZEjvq9kl8
vYqO9wtY+X9YRWqiOTDc1QuEt+BtUq5pCttQBnYUUEhkSjdbuJNg447Iu3PLxVxT
mNfZLLmnMC+1jd2cG5FMBjTvLt7Iw6fwAN52sqOUFi2C9fwE991ZKbeaiuAE91Zy
brj1mvb3ouo+7bH/KiExgqVszonBliJn6EmrnKwhqQYwmKsOoD3PJJpmgUO/4Ain
/z0LBb3+Tv1A4IEApbTmcIVdZgQOiuYpKHgxWyJCVt/XUvfaQnpC18u1CTOPU/cz
`protect END_PROTECTED
