`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zb4EAorbBCAE5oF2Q4vo498Rl8PFzgoEeqG60sPWkULEXSOOJRTMC4u9DFUJGmdH
bUHkxgOwjVMdbdWKUrrchbCSCZyTBRodnIfT+zs5TaeqxXgO7XH4w1KUMNrLsm3F
DO10Y/L9Fu+vR362D7eVbwpprI4uHNcwQAew9in5uzqBSpKBXoU+0+jt/Xc53HPy
VocQdgd/SP7sLfBujr1phk7DmiISQ2066GDMljYYiyiTdJ8UvyFsAnRNHOUXyaiO
Pz4jq2AD3poLGteHejofGLjFREFvep9pfhwzj7J90BSZs5UBGBCRuc3ryFBFd880
7cjPP1RuxcJqPF7xBdE92iWLMCrsW1DfzKXwVQ7qliHYBKecZdXO5/vc8x1mstYf
zF5FVkw1D6cDjtVuvQqpMRn47s4WZ/dqZ3hQG6m7A7SalxXW1TNU3t0lmJpaboDD
3JY8C9keeBmDOJDDfgBGm1qQQF6ogR3kbYI5+bbJ0zi6hhWlF/bHC1eIuW+/4uIj
96QGraAhpQRM2OgxoKFc+1JzcOEIrSrsyw1mbTr14RQ4UZgc1GK2it/kZm0wIrge
nuLsmbAg5G35xQ1OZov0qubZVCxF7AJ0HwHjqVswqBet9YJLMyed3YumRWVJHXwm
Yrjn79NXbYWMsMmls3IVH/7O1WDs9XPKOmXr0WLsegI0rYIx7slDnHjIvkcZ5GYo
iuzIrj7AW7pfhprUsmSSiAMqOmZEW8LhkD7iuR7v+TZG83SU1QysXs8nuceNSFmt
QY0ZF8dV+W3BXlHFZsftrA6bbohBvFCyqB41IHtMWw4Gp0aFrQT4ta9aqT+hbWiL
wf9/En31LNgcal7SVu+Ym8HqfKyUnOYQYMeqgt3fTeH5UjP/n3rrM4lJI+PgWFFr
Q8SXJxttmxAU8dja7Cpi8qnB1SziO9ZrUTQYQlQR31PvSviPjT7rxoHGqriQlxvs
IUITdxZQqCWYfiRic+837NDBnxah5jLQj91gE2ec4bEj6cfb9jrkkkJ2DjFiX51L
mxsHfcvVeTGjBrkQE5UZNwG30JA8zdqCC3MiSWqepSDUw3NxLJq/Dte3qj2qXcfR
U2Q9lySut0zlcFGJ5q5Yw/qpf1ivGTRNY4WVzMgpE4uvxiQTpCb4L+qSa9rROo0B
ZVZceFlUvi5XPwVCGc/XDb42WN6yri2Bx3HRioL+OOWeUQAhssnqXWLGkR0GBh2j
qiUdIWlScAN6BgGHWIyB9lVFQ+/CsqrFMFc0Y+fa5ie2fM5cmmIFIE8NQyFGJuHj
sP62ynBu5fUIWm7MDaWpb1GwV+tCXuaWP4GESaZFEkZkfw5IXKAvQEa5z5EWg8jk
7VeO/Xsuw0Ivqy+EREjKqT9jIIdfkgNyM/ZD0b0AYIxoNSSe6eBiwCoYYuEGpVEz
tuY4vVr7RtRI8JW5XYjiklE8ogLyNTODpL+Wscbi9Q8IqW1hrXkPgbZVs0qjqQ30
L9mlcAxp/PQ1atrhnmgQ21T9dumObje+iU/1HOF920+hCACuz7jgWXNgTc3TJ1zT
zp2P6hPIR9VV7ga2gVxUSgM12dd6jYFBi3QfKVjZaDhV3TX4sUbeFSC9N+T1+9/A
gv0k4Y/ZNGgBVK0g8/abBrlElIpQZaCHjRTUYe3xw6hQQGCJhfqBs0ezTBRo4NpN
8YINn3aniLdxe4S2zCSQ7wby7uwL3IrTe8BhRQpxy01GXTJJA6ay40JVVDXIFYPd
/McqnWcNMmuq0vAa3cT8v0KEOTJpeHUzd8dIQMNunfPRyA0hLKDhR09muFXVDlPM
yD2GqgG3Wz/FeBgPb1BdY2Al+M7SI/eSBM0ELc9+O4CffuFbxB3xhI4vA9X+ofqv
h2KNji0y3EkToojepvLddE09bWu67/7IqhI2IUuZUA3DYwnj/nehbUBTnVuOHE6B
zFV2ygTbilQJ13hax16KBTReUtkflVC0+xGmogN5YF5U6QINWb7a+fpwWaphealM
nXpnj8Zs5Hd2MAlpdG06I8bQjjFzmlu8AsOFl72oJvgQ0dZCLbg02xUVPamt27e3
KXRPHa2GSyV2MwomLWfOyVjsq9Ya0bqOnauKD5AES8bx7CXdN9CQVCTdeg1I2aKH
bkWvacZic9qG3bv/j+ObC+OGX+iBZ0vhgxNgAkGcpRrG0kbkXv6k84mjCHwabEJ7
9/KVUR/NCuFcADdZqccevuBCvwdCNTJAIiREiRtxFbewNh4+ZbduVKdSIfx9JQOB
7Gq7hygs9Hpb3IcWjHbPdulhm1LnOprGT3aN6BLfk28xpBvTwjp4Yfwhxt/DxQZs
zvjG7PXtS6p0Ci/5vSwk7KqfK4rPv0OICL8AgKnYqzNDv3BtGdYzctXtVzpSRowa
z8m7fDS2eW04IaeNMaS4HAtYAK2ckM+uRaGPn9+qr4puI9eEhTZtLUql+G4m1rI3
wiRrSH40tjbPPmC9eeSh60Ow3GLm5XZzgClyhqniwX4nGgKt3DlDFWXXfZryp+5I
RqS2L3fBeh+hI91Cp+c/pzwDVDZ8eM8gHOw7BjXJZkKlsVNnGxY1NzSv7YI0ZS+b
kYhXRqPWOX6lLTMHpzUTkVexUExkguGJ6kkJtnHOXWAYvxjPH7zzUtbncPD0tTGM
0f/HCroPWuw36wfudTV5PErbxx6xa5Puiu1i8YBl4OE=
`protect END_PROTECTED
