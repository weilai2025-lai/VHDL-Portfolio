`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjYzRxt1aKOqVf4APVw/WZB7UBl4YRqSJ2wKfLj3sH0OnBXr3C6YnIfLGTYBiv1u
MO0wtmJ5+/LheYV/ryKQip/Xed9EFpy4aSUgaaljLWEb0lIuUAxMpb/PkkW+Y1zd
iC7QQgG7Ts1un2Qads901vv1p6f5hABm5Xi5hmAgV+EdzXIq8a2hbQqZ+Lu+Mr2O
J/14VUGx58u4D+YWcfc0SzEgEQvVSVIlLa5KIa62BLNofBa+N6Q/jr7JNtaDSeOV
UdrCwK5kjXLLbcdXAcVeik3c0hSTf+9o0AyZKMu0jtqBXRRMzigD3idM1Tvxir7g
8cwWRfO6EIqgwXcnJwk1uwgs9TC8emG0DBxfz4Ek6f00sC7C/xK6ykVeYqgVUQ0t
scWhEQB9HbatNdfSo2ZMeU6KzQ4tKJd9SK2IKro/EGMNigC/MbkqJsXs/5CxGR5C
1YLfvYmzKUaZnzelxbfn5ftVYvOcL4QZuj7Y6mZVrdm0umdWkgbc7yjSyKOnlszC
2iRMLT2LpKcWhSu0i7JPIUdIXYTZo3K+8uW22C58qaMc2D+Gfe/wTVO3dvf6Jsiv
691iqSh/l7zZQz/Qolt9hbuOqjQtk6Ju6sM4bqQxENrYODeNpBcsWWq+V3GiyFhU
zNkFMmd+AI7mlcbWC4rxAcqXfZCUWlsJtQLyxax/6zSdslkMFiTi0dwBINVHNI2C
hPSN7X+P1Rms1915TPkYOndloFUpf7+ZBHXfi7p1l95ZFmVMurQjV53CKDV5fObi
Dy5b5sjL/qPq8zJJ2mJvALKczR8YeW3BbHpNS+nkjlPNPCxd5E4JV7CNEAFrgUfo
3IaPoNIkihHoipQ8K+092KkSQGXQ/NJ0rPHrcy51ZdxGZ4Sxp9HtxUnw0M8E4b3e
5HWhVXi2IDSLPDuQNz22Ow87+v/triQ1c6+MRvJY+7GOKdC/RuwNz4thQ65yL0Lj
1DKn6j214eMY+o1NnJAexDfDqbZWX0AxeaxYFOWITgmnabdw0hGFDGmkD1yoOZKn
hHfS8MbKqJ2npOslnOXPrGb/ft3kzcx3HbDYTjbJpFbanJfNGu4OUNgBI1fmnUAg
5oOrnmu33+5zj4Aiz1QE2wLR1nUwXo3ntedfbre2q/cfWIH9c3XHjumJO9EzDAe5
ChH7l95Cb4xw2hwOQCaF6SlXxz64Q67SG9mqN12XKBhVxZsaEFvnfNa5y3EHLVZq
79snxR5zUOZDSX4xGc/h1X7WeThjIN4VLcYivShihAdc0ZGFen8HT80P4InK0dP4
X6cjKhs5FUdlCWJWlMTu0rDh2pptC0bdDUJL3HrXCzm91PXrlBqZdaERSuMRxc+a
Eo5pL8JJ8AXJdKds9Aq+XsGMNzo2qvhC3P49t9VVsyW7vOx1otHRkLVduHzibJjc
lAMEoFUN6zmjb9h6RidJIJ7e8RasItlV6soUim5/3YEm+esbxuyXrvOLFt3k7o6t
nYBa1oUAUVXruB1lisE1EiCexHGeoGCEbEzM0pCauIYJcXVSm4QXzgcz6YVRmNIM
sI0jWCg3/YYymEVmgCfJaFHvKXsWZ6lnbPD9xMtlp7KH7ZEmzQ6sg2eF5ZijqKFx
ypE8/G15nJsC/WvweIUXPu5fpoZR/soiwQHV7jkHrLEqZSw0SU2GT4mWQXFOinAa
Mu3xSIJpXJ5WIdGSEyWaDPLAUtxHfoxn91FqgO90xNvyIoRb2UPv23YRuhYsFAvT
OLfNOHTZa72mSepex4yak5bG7Kr1O3qN92J8x8pMtAZ0qkbj3gZTrtSbQtqikZX6
RjQdREHHTdCpZ5K6/+fbPbqTKYK6xT5S8vYl+7+4T/66JK5xt/VSNhNtRq+BAiGW
kQMAvMpTZdq+q7VIICukfoSirJS3JnXuNPYv59ETJau654p4YJ2s359Ufg/nsG62
ZzQ8nG9V7lGnVvq2YykKtgbQtQE1P+YunXNYdSafKshBOv/sWm0X8Qv8J8bMz5SH
5VLxhMdIcvTm4EDbAXQxtOeSKGOVUsJKv3q3QuqCKPvab0ohdE/u/XZLcenZzMW9
ZoJdm6kOIPOu66vaOgYAuLMWdFI2BD1jnWWd6+5SX0Bhk3cN98F4cr3JF3hAXwwD
zR3tmyropuCkrNM8zDkOYJE0qRBGCAEREIbyWesaQQmnN4FJYSRJzsVs0BCk/skY
7mq10h7ssJBPd8qLPL6ELe2LlbgpdsEbrcUz9pCjYWXM8wz5z3oSnb4i4Vift9ZR
MExbzN3wdZ+TXM10q8+kOMZf/Q6cMlRvYdwNfyc2NW7ns47poeqMTLeY4xjy83D6
4EUpJuxdiabK2S4aaC4qgjjWDLNdJ8Doyboley64sbMMjUJImb35PO7vdbmeVGYo
j1WzB0pkmjJq7EnnKxxhIDexlYZb59U0IW7K1KKWwKWb+MBsq+Gfl3Q7XQaYnve/
F5FEsSUS3QQsjPTaRmsaxatzcBeRCMNwlg7Iu95rS7IOo3k6aPMrjUztFowNzhFi
JbhL76kejUCP6B4OAS+bek5fHhLTkzExDdrEYp/xxlIqHZuQwamI7jDZCeZ0wsb1
F6PGg38RzWwK6RKqTpnD8L/TFY2Yz/7Rd+/gbA4XtqljuOxQrb7dHM4dn2EzPWaH
N8eAq6nKKWt8FwsLVTMMFJ0j/0LwQzbj9kCRxs9kBsoqFWe17DBuKj3r9QyKjZT4
cvVcpk0BTMJIgA4fv7dtwh7jVrMRvyB8eXIPrgf5E4xodxmIHteU1jU5aynuAQuQ
VGtkIySu/U0CHwMlcCuQ8A==
`protect END_PROTECTED
