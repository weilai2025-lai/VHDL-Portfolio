`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xI/vCI1kvR5ltH1jAUxX/rg4TnrmY39ARXIDomRYfecA7xvQs7vks63vypXCOtH+
33bU9vAxV+lsAtSsY/cH9j6VCLewhjOExJYq4IIhH7AGC8VW3TtJHRXMISoz1/rz
+9vvwFn1ehF1xlDcqQsihOsgWegkRcB7RXpxTBcn8p4sbb0kGdBHmFvvSycuKekJ
`protect END_PROTECTED
