`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kSaywKM6WZt1ELfi8n7d8t8TAoXbc0iDO/uHUcGR2bZJAQ2foEsN1Rs3GBZVBGH
qw00a8UajmGavPe6754COYgZBFP7eyeXkQVbTfdYuGDPWMDNu74lGatl62zncYlh
t1kxreD78MGu7fnh5ckspKTNHEcm0jgQZKyyvlgeGVe24a+kH5sQ3uArdtZ0B2zN
+bZdC1NJgTsQ8yGWVxmNEa4jpTinqzwXiygzSpJtjxKNfxhRIEmP2g5LT0rC9v5B
V4MZng2I/j40TBtlzUw1sl9T/zYj3fUBaO/IVSkEBe+WL7Vi6TSx9w3G9wEKTNR7
mcxFgYpZXK+lFXYOpMd4T6+ixYm0cG1QH1nXNn25BecZYsMSsDPOecvI8rkXzjxN
`protect END_PROTECTED
