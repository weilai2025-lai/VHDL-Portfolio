`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvIGWqV3hKqljLxTDLlQOgzwbxAY8TJfr6XXkIRA+FKHjwhpT5tD/0zCVdlF79rh
GLK2FBmQAE+LD6Gror3mVsTFFaTsRoUYykIdveT9Mbp6+aPFFIFlPKr1s354C6eM
rVkkiVMneFR+QlQn4Zb/bKrk9S0bbwrggCxIE7c0aQDmKSoFS5NgCdFnEnt4F2me
lavKYm6WLNxEXBPgJt+KkvkmvkFkFgApMVxWAIDkr+DxA3T3+WSCUsEhrp4vLIqL
CBZnNxqtOVzCGaaJ/lM+9Nk2bAiMIu06pNQluL25vMxZw42bdtMVpzxXYseP42rG
M85JGPSCpvANP6Wt4IRmbkFQ4/xaUYEfWn2dSFfbWcSLk/kxC3LPXtyBBAj/QIFi
7504AgEOPTesnGIZRAWyjSn1znVaFXyqHBIEyXUA5Rv7Clql3mD2jAJhrBb7xUDa
3SfyVmeb07k4XxbU0cssYekqtlct7VnclhO5+/my1ce9gAqUPgvXXm1AhW37tAE3
OOP/V5wv8VRcO7KgcENeJb27k+XiLeuiurlQLpUfN6bYqTpO+lJPRIT//EcVHZL/
RDflMr8gWz0m+TP0fnh55QJxuZnpOfvEA/g5J8+nSkuriMD5UB9gkoEEvt8nH//z
+SQb1hCqrrsYF9IiY3EAJDQ83tZJrztGwQxmNbXUxLIxAM47zAt4UVnmk1VWmqdK
BcOIfLiHJA5n6pSd5v5Wry1ttAm26WsbxaUewQdLBe7CGVYH/lG2M6dtP+/3lGLQ
Sc1BvWH/oYVgmNNqDGZDtOi7/TooRnwtyJNMTIucybyKdNhIcVkoQsOMlOFQKiH2
viiQEfoCdW7vMkUQAN8lhCv5bBYAgKtDUqv9OE7mlMF1xhr+QWCgoTO9p3Zqqv3x
EAb8c55JKoOa429gmqr3fwOLk+bQPCNi6fzR3Ya4Sa87IBz8jgORaQ8KM988vxme
eKqNj1EhlFk1Puk1x547nOS3NG74eRMy0UN7awEZbvIc6Z22D0nb7jfVlC8RlJ0a
A8VXM8BgeFyvOcC6IZSVyOJumwd1Zq8qiFaU3QtHWbw85U+ZTWCtVWkFr/42TTYK
GJkVxvgqxhxzq+4VFnVPmBgz4SLP3p6gVU4OOTT172JG6zEVhzfsOrZBmtOqmJkB
y6YKOPittOIkMkmHYol9HRJSz/hruTMAssnXoMCYAJQ5kT+tZ6nq+Z/7ETSUigtB
UsDHdiuubGt1M4K8MpY6BgDt/oU31zAyrRVTUIgwOzpwYrYe+ivEKftTk+kdCw9E
iPXimfZXacRD/d388tqEkeYcxYHsTKYvFAS04wsrs/smB0/hkeKESzMHmytMX1di
iqnZiXpn2mOf7ze2kO6kf2wDMYevgpWGY8kwhkY1hWaWMpHCFi3fOZPsQGjhhCqd
8hldg93iWHcB5vKd5lQgbftjHqDc0VlD6ah+fHw7WDwjS1hQc1uJcHD5jEFvyxHH
631GAIXbEyD7KDHY7H8hq5/hpV+fMyQ5dfJkBJsfl5CcM8m2MTOXk5+Zyk3YfHTs
6e08HKC2LUfYa8X1VKRiMg==
`protect END_PROTECTED
