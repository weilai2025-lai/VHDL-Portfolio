`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uy38oFoSpOBA1tYol4kH0TJ0WGuwEaIoChO1GIM9JCO1N6fozvUAGEnAF07EXbBc
OuWb5WesWueciUu941ZiOR20ITmBX8L37rqgianOSMvixqFc1rZguM2NMNWjZN8x
LqgG+I8DVbetevsN0ueT0ks+7Oo1YFLLzjcpViE6s4OU0+40MdRE3eb0J6sJymdP
+w4PGi8J4Rf8Mh0eiZO6L5nYXtQrnMcKctPBGzr/so3FVMOdHAAQAVakrfoH+ht2
3tRxf7f8MICS5plXv7dT/vkaaMa1sZeMy31he+XaVDvf0RdVbwkIwaDlG8zDuDog
0PiTKJb5FgtbKC9fG0Y/QJWkULoSPZMp4YSfm5JQU8VsdlFxjcUN4M7DLHjVZKHz
8ib8uJvaKnKX3ieJkj1naXrkU5SiNjL220HiV72jea9sBoUnKOShPkEPlEaVW9Z+
M+bCeAbgzOfatUk1AJwpEQlMkAVp7QuxIxwsHzBw5OtYKV9ClLIcr3CsZcuHtjEh
C0YhjA7vytm3snSj9DHCAn6jhHHxyZNhHyHSrWWLYLPYbYhMQjc9yICnTb2T3s8E
Dh1uOHin7ZTwm6NiqzjKM03Xq1kskOCrU6Wsy18CuUJWFrj3AXZmo29uzrc9meiw
eYabt0q82bmzYgwVAD6Zfu/Nom9diEgR4mBi6NBPErwO+Fxm4qrmKxDvc2Wuu24I
`protect END_PROTECTED
