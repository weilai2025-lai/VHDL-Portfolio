`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8TQ2TpePEFpTJ/1jISq8X5DTQAREOWIXiAIv6yCFIglpk5/2n+Zv/M6MptFDhMa
8ew4tFQAe1Cxhc3A3YrZ+VZjOGP1oLQXoC1hBsgEf5D6k2LgxuYb+wMAN1BZh3uf
O5BRLUaS5ac8LU5r4yRlBdcS6P3x1GZQybTZQ3aIKj4WntYq1PJ/KOnWS1jSxpbW
GNY8jGkLcGw+qFuJyeXpj9olk4E2mKzET9KnXJw/resqaEXCNVD+Biwq2Xnb5xA2
F6wN7samLT3AlMch2aX6jhdAxZXKgN2BJQcHv/7kvfnV+clTEoHn68i8i/1epd7t
UtVgx3FzIQHpCGenq0Ie9FNAKPE5vpyKZ7FzrF1nflX+NAydajJj4HpjkuclgK+h
iueLjZFjlPBky/GjEWXvF3UbcuJI7G6F5StLMOZWL0NDcM2G8doio0hp56F8ZHKG
5oEvQuUhNHBCpXGUVGMpcaK8XgmpnFyUZu0EvDWtw//s+Cl3cYEjKrfIhXTsNo2R
VGe+mEgj1SKnujtIyVQn9YEDY3i6+kwsW92cPrKP/h3fPaTbYdjhqa04PqsqQO2i
Fv6AzMJFPDY3IQU3TvwgZ1qxhN/MTmHjJeN9GTwFWKJskPAHhHsYzkEaRxM77QfS
SRVI3x2iH82rTFIQyaOk/3bYe6OlICXvaw9VDPA9FOZpaaAVvsw4SE1OtIpZxrHS
osE+N7PqrK5qsu86C6C7n6lVcLlCFbZKU2c7CSQEX7taNbB4O+ldaHVCci3u8CdK
kCin8ddrSjiHeyxALt2sw9ZMmTrCcePek+HN0/VDIO6OJ4rsMaKAbzJ7kKAwbNRj
pFEmpsvpxQkPxZ9vSn1wPO2EfOKOANkZt2Im6uOf0hHa6orhsEcXY6IjmawwvfXJ
U0A8kPSvFZoxR+HsNwhH46CkHlqd3Qf8iVmnSb8Uf0e+WXll9KQMKFiyMs0FlgCR
Sz7rV+qV71Dr929eAUmloyDJVfxIJp0MQYTj0mrLVSxC6+nh55PIqepdBbbkhVjK
9nO6hP0/AHmhM697IojYumRPUyi9k+nLEFrZ2KSX1Ef2BggV66E0+Yqt1Xjl8tFd
K1oRb6QTl5OEAl46ohCaG6XE+yLEo/VtYM6czW2iqGXvw59wSUyOc+5tc9z3DEJc
aD7o81FHcQrWbDsyJTrbcMvsYvdjlAP4jcA1G1UbQrGkRcNZbokVikHU/vftLDJQ
1Nowkx1nTU8dDaE+TJJyLCwisduPePsuLIlMZqii1dMfgg47nmwEb4OZLMh45DGd
+vf/jX9CFNxaua3QOn8ZkQC4AFeKeAwn74gVSlqnH6G+1yCddGUp2Zyxu5CQz804
8vz/WFV7RNHQJs/v3T/C2NKOFL2SQetng+Nyhv8Rg4gkGhFvBZ9ieqnusbOBhP2Y
7bMER+3DPpgUygGIgDkdt271ju03nIzO94Aq9CgDhwoaJNWup6/520pxWMZNRUi9
HAOa6zvxC1oH4dh48XNlWd6aGUBxNaGaNgLII694SDNrOKpgHFlVOvQ8UnR3CzG/
+xZ9NhyvkEN120v8kWqyHPYSRnfWK6B/Vz5C7ym/Ffkj4C7fp2isNMbOEji+2ZGi
kiU7cI60KjnIzpTv/l4hQqByZyyyc9X1oJJva5pT+yq/gA72MwrpTUW5NeWEeHp8
oN+Gu9o3oYNYoyQMf9gDLVhdXzTMkskBBeKSJaBa2R7T0mbPMXQSKrj1xmSON+Tw
alws0hetMa34L/KLDrnkaFNXrhT52Wfy70czmYlS1AlWubil9OqRltoNwAKk1MRl
`protect END_PROTECTED
