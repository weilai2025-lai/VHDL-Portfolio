`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o78xdrMcrcq6Oe4iwfsigvYbmmQYw9ehgcdYs7jv0i6Dw+xxETklz0GM2aHeqn9S
XXE1DKY3ADJw/BHgEVHNkUZWtuEU9QX4nGz972aYQ6HSROi6iLKmPFEOGrWEkvif
6FQhPnEmqfbrOLFli1+XAy7eKybZLD3zx3vZHTiFS6Ds5BEICRLS2HCoT5HNDAPo
arg3ObjwYCc7rH8mB8uNAHFxZ8dcNy7oSJvYpx/8FZEB9vv2Iiv6PqYWtwD35B1i
Y55ikLmdBz4gwTekOH55T7d1AIKmOy6hruNS+FlP0B3R5tfv6AyeYh9NHWz5nV9m
s+IULrqkhSaPc2nbPccjAM+NSKxYlQFT0xJI91DgPZI7wZy/SujzyX17RZj5AFYw
PkWr0JhOIuw1RfRyVd4Syl0D4HnRjm2d/nSrq6Y8VzEn/0nj+Kra0HhLtjLQSG+B
Ol+fZ/h1QeEqjZ0l8pAeBQY5duppSapqljjb3vuGCD6Hhowrhc8bzzFFRXN8oOzd
VtESKieja1caXzbuRPYsBo1NX4kXOgGJElJ4bO7lg4hKcUtOzIoK5FFQrb6v0be8
y+GduaypmpnI8Y8ybGpCz1yFvyIsqymVmvv7T6z8SmeOtqz9NkBkZD0kIl0o6J/z
IAlpen5PS2Ikf9Waw6wruLLaKv9NYycgqM9gcNTu+PmBdJMOEfBTHGoKUOjBtEli
Lv7okjjOdhvefqSnSZ6npNnQYTNurNqtDsXR5q2kYMm9hpxkPXdAymCqoXC6DzEv
ySllLnKbmmcmejbXpZFSJNiXzktbfY1MwlfAAnECvMc+OP5GGlIBgrgYmOd83I73
`protect END_PROTECTED
