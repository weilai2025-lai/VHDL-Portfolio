`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXgMxYC7vACOM1tXu1ZkvMi17qNhjtKWk6SmeAmA8hrwVoXT+YwDMHeQ2AlT2mc+
m0YG4iIeUd/tnOam7jqkofALMSrDLqF48xVNgUTdlm/UHTBCzSS2E0merfMKX5fV
ey5bTWlgcUMgPZ0JDmqEzXOWQoknfR37p67rXM/eX0AMFEizMudSKqoFlrnEGTLt
5xry+0tI4rbeBiZp8kFxgbu6lo7Ss9JyHDMVzq/v+JrIVgXJiMS9e9A+Uq0oe8Ba
9cEP8SaINqtOJJpWipmRzTK8cdL9W6yK2gWhxdNP6y/jBB9sVEUP0/HDx0mdLYtI
Wg0hmO+tX5gKdLTijPhDpE0YNE/MrWugtNqgUgzf/6OgFQw/ebV5Z1E9qNHLt+WS
89uzzVsWXzzjzhHAjW06BY1esow3Q56WdOWI7AupMdcjqrOPHw3Wvaus7psZeo7w
nZfhfxtQ1sxM7KzGBIm5wMfWGGfUaFw9o8k/yUHrY+BsOu/rDNLbctaKBtL1tWJR
rBg9jWyad2a2ULWsfsjt7iqC0WdMOBqLGMBvsN8sFGLfY+BkRaV3m7X1xfAivRf3
US05DNiR9S8UTwzXBIPnXKrQibCb24XbpJ4BwiAsli4ZIfDmFqIamgjJfG5+DL0H
4kLEnzXFxVbVt7fy9kv1ETEFLeYTzUkG7ewh7Isg7H5UUNAV82psYtFvYwvTmT7o
tXK3J5Xx10fDFTWbQIEw+sZQHjxO5xlXyVGoeXQKjstR9wGuguF5yVwuplPHj78t
HDl9g1iVNlVi1uf6EeIZIpec9u9d+9zBSFZ2CGa1iE+xutptrScxzX83891lrpJS
sFwuvuuq3g0hLb005NSrVsOkvtaCAi1yrPwxzlCSVPo3TpzNPFjCT5C4qjQqMQXs
G19saNRRqbEiBapq1SXxJr+yTFinCeNZU1CTUuRVVKVKdA2ZGobapEzJyLNA8MXs
FDEYvmleos7P2hRRs3YwQVDzH+tdQI7SebpWkbQuGl/P1RAoMIY3vyN6zKUXuAPp
qEe++3FiIJw/lh0wF+fTT09lRmTqcHRvan6eGENa0mMyulDlY9fr7A2E1c/1rTkL
DcdPIOcsueOp/ddcUtqk4rvjQ+vplIEbkwRiUQAHMzJCpRbj/7itP+OzoiG22ANP
G7x+0N/xG+izhnYVe4AeXqYBXFVI4jqKUe8FIyAIkTkGMwSCNYceh57D4JbC60SZ
epMtjQoiOnV1cH/qQUNI+vhQF2z5DXgK4w+687nf8KlDO35w3pymk7gIuzNsZSoX
ruZIyUE3cPgKbkechtBseoEVYYt8iKMALNKzae8/Fvgs/MRWb2NVtiJJlSjc+6zV
ytdK/AbkCUVTzRswunCvyLTAzbnJgKpdUC0VFW5CajmyfpYWlHskj3OFygH0Nh0p
chF0SXyVEe46u6BGNxk7+FKAEcDYuDEHph+0YScr9OiGtUm2CM9difYkl4wzNAtR
cqGthLk0TqArDUHzajqAvV2f+ZKUzfz1rmW6pULbFf55425RGZQixk8zFtw6aUGS
FsGe9Cd2oChp+1Q77UZBwLG5keo8mlExhetxsWMDOiKnc13/91L6fgAC5+OXFqHw
xT5bLF6pOev8ZBYWwwIxVruwLvKvvMtcHkiEfBWvg0mOWujx4c8SLLPQPe8g0jAY
yDYloFg8gG8zOla3GHfT0wufhx3hxsBMfBGyw5hdGpWrY+3wzYfYkg/4UrV3rTWq
a8B4qlcNbiEtM8kk+PIeFiN2kyh4IJJOlzv+g0R0bsivPZZ3e3l/hfRd6AgkuLdx
z0Ktpn78kTdDvMJOj5Ma/SdRdJwBUaiQ7EI4OpIBX2zhBypTEC84BGmUhP16ANjl
/zKxu+Fjs8PogQ0q+l/KfVpP+l7GtlaaO5ar92gN5WI62m25T1S/athcVKeyXUN5
v4YzqXzb3ccNgHJTE1gs3M7c+GC46/mzxt4ZcNrlmJc=
`protect END_PROTECTED
