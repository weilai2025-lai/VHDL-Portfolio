`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uT6HDst9PtRuGNuxFUs3d6LMKyneu352ztNpVy0ZRm/UCpYRkBPFrQdbxjFfZ/Ub
T1I9H3c9HFwFbcVVhA1kuOQHo2jNEgPawqJ+wawLUdlFHtcXXgCwl0aite+wu1JF
wGptrrKupw2TC1JxvJgZbQNhysY9dkd6Fh8nbnNvtv6xJTAY5dOXmH3n6DEwvLal
ffVYRJpHvFfj0//rs4mZmsHXNHleFSTFbsEn068efZ56zpsILdLaTtg8suShLdYk
pGkxe/YfXFvxaAUfmXHRXIpQ+s+LTYwURFOtZ4HvyfZA3zna949f8qaH4TBXHgVa
08cRK9iLlvYUCif5bIdfShSeV/SsQwQF3AFrJXWtnuMK+kW1KW/frDqODqhRuKN2
pnnPmDRGx6FTOqABFyCeGc/kUyXzT9DzvjOLW5H8FwLSHfvp7gWNHSJb1l4HMs91
cizLjwnZo+f+8KvHu/SRynAc6jcvV62lYcXqtB+4humZLEBTRvMafSBrFs7PlCui
xvHapOgKG2Rg13auzpb+1zdCfLlc6hRzrO/frhpmdUZDMnn0P+tr5cOn9h6B99pz
EGHtzBT749FF+aklqWbFjA==
`protect END_PROTECTED
