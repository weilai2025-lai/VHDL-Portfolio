`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VH646N09u7r2OvwZP/dJ4evjfoTonMdMWHi+g78Q9Gw/u88qYDv4WYm7yEBtpjJ+
JftKtMa9QuEECP1XNRf0gDrCPCb0wQ118KT8okbLiGKG94dfcehBpwhfBTCVVL/n
5vnEiNlT64gaLFrkpEa8IaFmW5jEHwAFMAMiRE4/vpGfWR9G/Wpbad2Q7DtKzf/5
UQjpVoyoSUJikormlpNaS06TnxOEjoevmiHz37Vscyuz79Uo9mZZFQGAqn+GBnv2
YS3j+ER3KBYqGACSg8N9ZZVKZ3It2jXAB9fXfN2a3yjVtOWXkgtu66wNflodrOFH
VApjKpFvbNAq2owNajnDheYqntZNYjMdhxoFObpZKUXfRgq3vTJXzWacKSor+FsF
jWHhYwPkZpHLFTbsYpghwXxjUP4lWxnAFofEjzc0N5NmDgVLixhEu2hPY36NmfM+
qNV5/2HtUsOSJjRsbjhZ++r42Epc5QYGx4jvo7Ws0kr52sXdTFryFZI8PM7o3ZoI
29aliRKSbNmb5EBRA6YEK8XksrZHRZ8X3evtk9MKo8Zld2qB+MSDt1JjUWlvaQs/
2NCeHOAC3qa8P7mpIRzEvFvQPc3jUx9Q37+YgrtiqJAPua42bQwLbPUMkyUuuWUU
K/8Ctst5ggNinI8KQ0pSWe1PmnVZJUb0J1UFqsDo/gcMgxhfXTKYF2SgjdS4fLKW
qZtIyX0zqDzPfta5LFy6xBTfs7HzZ7iAQMzOhKK8iDK+oochM958ZMi92iTcY/19
r4HL7T0xd3WikGoaQzfX39PmX8hIuirJ2l1nRJJwhQ02Sgh8CrCvHALtWSwSYZni
fvNbPD15RPJPp4uteG+PmmfsRwEE6mcRpr7t34FD48rdCnLDmd81ikWgopaWkJfb
XTBruDS8QvdWkej49+Yc8YxByNjcj7lzvhc0d+5u+IX2mFRieawBy3bvcH1u0lw5
c3Jajqk2p87NaTNUhgcCpGrkjPy5zhBQXJKxDbJ+CMilrDIf1V0CyjkgYYLTfSl2
YuANbwCB1gA78yYjNMuDfY/Z0+2HeOvXX17v3Hb+fGFRpok0J4kqG81s0PIIxlfc
rt3SDuwI295/JgCR+lXywEb2fo6fdAh/+HfOoXvVRKGlBFuLOzWnwGe0/w2vVIw4
Se5IGA6KZxKK6YT6LFnJGX9tGG18awV5I9rxVHHT0wzj19F+W3p3W+/myqi1hNxD
WoZoFPMMaOnjWuvAbJrHCv6/Iae7nZgcRD/DvZMb0zMN+mt8H8WeyMJpB/Zywaye
SBLKBZwJ6uiEXyPXH+FcGR7gLuyon3hI0zD3reqt2k+vb5fR5gr+JENkKgk/3/bK
Zyllr8E7YO5ANCiqEstIO3iMru2gBMiLC7GjV2UaUAQfs2KE83gG/HwznpUEDejm
kXC22SU780rEJDnjUvZWHWWGib+kkqJPiWK9Rv1ObZyzTykGFqzzweLzrBELLWSL
KClj5W0TRM6VI7EaKC72CBrWt4AdGwTSPX/2D/Z0fXTT6hzEf9zr3UbGEmoQ1pMl
bzy8lDTXC3qcswQVxFVTaYuKt0wPwCwELew10j6D4QDUHCQNeumVgV6T21Cg2Tt0
EhBpnRQOGM+M1a91s4ZKXiWSXJcm49LqNJJFEpITz2+X6Yj0feBEUGQ/XZMIGtIQ
fh+7dJd7ywq7t1EgbcAR4tXcoc1OAaKwlHy4gUb18+cfykYWGVCE4j7v6FhtreA+
TD2NvqtmOUXLOjKlzvXZpkN/PPx5a5SlLuLlqUwyVYaL13Oik1A1F19U+yaT/OqD
kerQxIRPs6xKBwbH3FWwydgjI5Lli649TCn5IRSTzlh1Rg8lyEvNUxuwgAjt5d6S
DcY/jfiRZ7S9NDjjHmNZZ9kogj8TM8yMKms+xfcjpGJ156zv8/p87mm7Fs/Qy83R
uDYQxgKGmp3CGegRBJCIPspfLFebyZGtDEXlsVoUBCadiLdvz26jvYU6YzGXmkvw
aqL/jfw7BcVpXprhf2L3sdglVwkaHbA+32bJX83RMqhHbq+8/EFq+UrNtpTISCux
fgarApjNa3qScEegm2sm5BeGAEMxCUagPx1tsfQqbsaMR/54/DXruGVoYhLTMi6h
5kjpfa25W4PN9+Xz7Wl+9yhlIrRKTBz4NOYLvjapdRs6GY/SVXjksOqjEfpIWPKO
9c7OdW29n3gQdpMixLFhV1i1EZBP7xme7MDjkaHSWengeIfZxgpH83nPWL7M8Nu5
Y006m+G5mJ+GaTxkPOMyIjkMARG+iqXQYYf+lFucVufERJK5gFoEdTY2cbTRKZ+Q
e1opzhvVo+oVfX6z+8gFZflHMr57DLg1c40YemkkdBYz3HXqcrs0sLTNOifO/8w3
4Mawjmffbkrw2j/ITLkeA/7IolI+nOhMfzNsaGbfsVMo/Fr7TDEG1X3eXLRCEfIJ
Np8ohIUXhSNKpQ1vlXBhBcXy5P8Wubp8JJIygyi73qb0BLftgQwnUxXdqiwg4l0z
+gdsLNScmfvDvyamNxsYb69RmYQly1hZE5evkLVdSdqd4qFu6ZtPG5fectx7sFhE
ACed97ujMFfnz+tzag6Pc3hg8MkMHVWWgXEpeARrBt2mWRAPy+1EAIMUX7S1aZYC
OOnmsONU/doULWNm9RaieaTpEiNvecq5eSztMdL2WLTZs9Ah4HhqG8+pd9qC243f
m4vReqcah3+kgYaR4YxYK69+Y2FdqW72arAt/kuYCnO2txRAXxg2I3kSsy7lC4A0
2iR82w3DsI74eyqrUJLTo6dLIJHaOEag9UACoDryvjDG93P39Oqp/RZWDy7J5qWv
PJvRk4sn1k3qpcLgaDjhbOydVKfEl2xpwVuFPg7LhEHVdw+skxUPWHyxNnXM1G52
h22Vbk6xpqxny/d0qcoptqofxM+mlpbT5sFppXtsD6RtjNbeti63r5K/hZYtGQgY
0+a3Ce2RyRIWYPQvVdB/WK6INS9YQ77zYv97VIMBonrqn/vAn6Oc4ttVui9KoR1R
zl3d8Mw6I3V8YLh26NjqgFcdZ4lVEK5Gv3BMH+0GPcfbIoR+SW/F7gpc8zC/xakx
dU2N04eZivKbsVr5UaX9IeYq+7CqWb6+B+SYdT/wRifiDzeI4zhiBhNUDterlkiD
tkgwfnJuWNd8E4RtrjRq3SrIaSvMexVotWgJNSL7mYlDBj9/h+Fcj3+hflgZeJfT
b/ehzPiY9AD7hPjD+5/MAayLa3iHESBGex/gReJm4rG7rXLELyxIqBQT2Ak1Hfe6
irUmHUexagtDZrs5OS+8U7Lklsf7Wdv4P5aNWY8n+nVKflSu+WFAQDAyk3Yq2tqO
j4qQX8wCuQInIjRPXeYHhH1yDL+Cm3dg+YGez/LLkfXRFPrbfZdg+FBCz0aa6bcf
qxIfG7FENLcHmBfCZgO6oN5y3rgTPZEzVIqIuEQtVAF22T6zICQqm4XMP3Xu94wP
86BwBndbZLPWuSC+Af2Ujq9hsPyzlARDM7oYtss5q3mZbK41myFutMwD7tNZPLRm
kZ7UmEQgHEgEmM5e8sVjmnD7/X6Lnd8vM7AZ3XJ0yU/UUkfXNgAweLH3RfD3NREy
X7iz2vm2cDVeCnvSuUfP/iaqAvJ/spxXJRdGL6OEMEAChMx4HWEavBJk2BXpPzvB
9RVOZGili5JH4uTh1r4F0AJnWTmywzDTVQvItv6yeqMiLo7anHlC50Ww97DSHnup
B63PT7sJbtqrzTUWCMzaqWoeXfGncrzdCzztAPD8t3n0LS8oXBKRcoOCOTzsmr+c
ZwJAJlyzWEWEdSiw2ssCzW+nhHjQOxhSSNcHmXB9SjATlY25mL3x1sO3KIFA4yiZ
MoeqGKaqtceVOLRpvmaKhBUPY3Ea/bqTzQMVYxgHAKP5upyCXTz6EJqDpRPSY+6b
4cOnmrqhS+Yd4ocCRlzMcKNXSOnGhqFcYqK9h7TnQBpcpZdsvbNhJKUEMguVzlSb
Z0c0kRtrw/72t2i+5OY9ziKL71ie+1z5nnpgaz+ic5yqLFKg3V+eFeukqXRJFgx3
UdFc3bzG46mSaWN/popvTfRb7X6G6WdGrI3X1h48iO48eW9aXMawU6GEPWKy8Tyi
1fhPBUB9dyumAOFqxQ5ppWhLctCh+X2aLQeSy39alM0aVROuoNhBE4ef7k8dYI4O
DG5iwpHuM4tl7F+U8wqoX0Qw+bdMY8mKcSPlZBSbsBZevmTRwhQ85hTvNwrMjnS5
m8UJ/AeKyhOwCqDa6QVM4fzQxHpjQ21bV0IAtmlN6xeZXoty/fISv548ubGBxHDF
6S6TG054QIn6iTrFJ22hrzPs6+pIxzceFhbe6bNKwfY/evNB7i5B6jbbQxS8Y+M8
lHqK4jCmMlv2XYSlmGjnxpFhAvqX3aXllkwIugtGefjOdKmIqdgXPwxyBWNuhi/Q
MAGTpPt90q80FbBb2Xr1coRqHZPMOzsDnxNGUhRIZTLTYLHb6dWdYaLVXrhuYsAI
fhZtYYPRX9KcJdGaBqe49SuP7QQPKIsVWEkN0tvD9TclYkA9Jygcdppu6qstfbF0
Gc6hKH1aV6vgHu6YSnFK07KcQ5qh5aVh+T94JAulRjBcHK0W0fwy0vmB/GbNbKYc
iDDip8ybIiFCHpFeDsoUuTqdZ+JWfn54PgAmHU3F9hC+WwneITprNy1PFxmUAg0W
I6T0VK6vlM5dJg9G2KcFjZx99u4nJ0NGcuJhNmBSuaBOd0ejM77BBOH+WhntBYz4
Tf9cpok6Y5g91g/c3zoUYcPk5FmAEqti8DFqYAqh7ZdzpoO5Qwi4VubD9SjY4fxK
a7MJgAbaDB1BvzWDieKM+LJWW3I2w6vr2/zOkJMu2ALrBefB5Qu6FoX35sG3oE4d
aQ7Kc7NcK9UzTn2WKs2ndCzjEvXY/VGU7enMYDWlnlcj0BBp0UYA01za6Qho15Eo
8BnsVPBDZKtb6Q6Hn4IUA0PAV65nNlpwrLb6jbK5dsBnzlBlHuICFFUj4n9Hzq6r
yVi5M4Pwmx1/03M5v3lGSEVNiDw6rlf9h8gNJqUzDx9TIDZ1IJmAFJDOH9U6dWX+
qFDD4/2u8B2YQyRG/mDFNfhBlupC7Xwt99QWNRyjGadYukut/ekn+ywvwbG1nWdC
MMymeYexexL831gIkWDAxf+4b7saZj/CBrr74bUL6jI1NwsKMjCDd1NUS9YVl9mo
SwZfi6G83eE8jpS8Y61XUHF1NR4gnvx+jggDQ/b4DofDqhrnZv4cP7LjuxOmGVz7
zDUVReSyG9r9tvtQFwTwLfP2Gq+si4U7O12G8CisF8wFrHcsXL3xlhhm2noG8bSV
6PcyWmpIkCPQ2WYAMtNQ6jAldgOP/C3grNbO1u7KKbbv7uAru2miJ0bv2BDbslqO
YXdDnD6kkXFiffngO4kAeUl44bUGqGo+g1y4du5WOpcMzMNGgYNh3U0wnEQKWJHY
cCRopxas3bdJcJ1IxTm1rIQe3PGemLNRLuCZ9t4jdcAttR6B5QT795jXCeb6jqIb
xHK8paGW0u/z4y9kYJmIFw3Tm2YfwifE29VlbbmHiPLJKptvYCSCdRI0hCOKn29+
4xPgm2tgqODmBbKMfQYaouf0/LUQ9K9yY5peWhLYz6CIYb6jNt2/bStdRAa/E/jP
jVIN+gAFqQhTbwCcC45Eya1URewHJMEvN5HtR8xNFlEgDVS+BGg+Sn0aSRPYWsW8
gdZ3Le+GgH9d6cQXFYVUAVPhQHS9pqO3jEoFH4zanN4lIt8fVbWpz3s9AEUwzTP5
hy3uNwLWr+J+OxJ6A0QqOxH10A3LTcgb0Q9Zar0wEfUTXYbJlPKMQcXgOd64fzBb
b9HaDmG7mWUSBtv/To73/6R7T31Uok36T+VPTaF5q9TUxjMLoQs2ChY1zb8daeUL
AE8a2fBXdnnMzImpqZGRge7FY4pRLhnZGiRGU2aeTvioO1SDgw2CWFq02S68CoBO
hPM9d06ONlOZjQkdkvVfdClPz3fxbxrPBjDAofh/DN75TpBEjrOBmowJmS23PpT4
NesC5X3MAlH6vKy0HC5ym1UfoBaLO5Evh67sloZAkkMaJCFIT8kixLn1u2Sl0+Uq
E0hGDzYI7oCodKjWl+mDAsy1uwMyRz3CHKdV7gghjd7lA7HvC1wpn7VKX9hjbPVp
6ac2udPmNjPDcsl4nUBW5uRpenbKp27NfapMbLdpovJ3ucoVbeZRrgoByYxIK698
6w87lEGviaGcr+tQBFnLPRKaDDHKKhTIIOcSyuYnN48cCF3izy+1PaKzItU4I0bS
Ha1EIEGTYZU/x7KAMVQLjMyYdCrpRsrH40hxr+xHEmdb4e07HEDNF+XBrQrfNkcS
tXwrR3F6GHmXtByIigJQRPa2Ns46sdzC58vg65Y2nf7CyQZ3wk7hBX6U7fHkATEm
aaiZH+kmjaz6wAveg/sJLnaUqX8EkqUtA2B7pBRcmnusL2jhOnrt/eXe7e1MT+rt
DhIUiozG7tbAw6/IOXEDPgz6oty92cUmiDmmTXdFSR95CASH4C0obWClaIzqyThg
fSNHBYsTfGjCxB8bKbf25v/A4SXySBKe6EJ/Iz9hOBdU9ZbKrLB9JEXMgw+WNJMW
z4ZcdN3eu2WPAIBZ6p8PwRGjj3pAvgk5O+30VarQuw6OaMyPSc/LhsEEDs+MCXs6
Yt4fejPPFT2dpdVrp7bA+j5Zo7lnF0jiIo9WMtqo4Nb+NKUHZk/q/8KJReSZe7bR
37mtRK0h6x2VznBc5+rymbsKPP/PwyKt3PTW5r2eHGMF7MHeB+9hcrUwhc5XnodK
xCckFwi6ieBDkps572pEv8yk6wf+KHczKbUYtieMXoOFx2HcHJcIyp2WXHl+1AyL
cFsSVdlCXndM/wq7WmhCvOWO3Bqft2Gog1yFq3ywcJl+O2tvbXaesM5t2oPBJPMQ
+Z2sbzQTVxYdsvNz/yQpMqTS+QNH7ix6PWNZgLw1l5CGDDQ+TylNE84iD4A0fySe
SJWZ80hX9FqglWeDy46qoEflc41tHBV3GN++AM28ZcYGxtJmPET2grXq4b8tw+HA
4tcbxYPYydXFafe1IljzoPnofBlw1X7muKOV4qf1VeAjSiYZIDroGao55/mtVIF0
JZBSHm+WwzM8neRtBU2MtfxgvqI3hTPKWAJd7DizjJUxKqVhzhAbiqlTWhLRtkne
CXu/cTMG63ur1EPOXrrQJwz9u205v89DT5C5KA2S1OA7tI6/n7T5gSptMsrgu2M+
DUdP3XRQxCvetIxjeLq7StulorU+tr+rZ3MD2VgS1SiFSPMN+zuUoFzmgfirAzF7
Fv91upojA3z67cAld2g0gWJO+Eash6FrCYUCFNPoL573F3LYUuxkbtyF+LgOfwoO
l+/I7j1ySgzML835W/+mQ9SkpXzyUjFSNdWZJCspR/XVoJ1+UrNXemhYjX+RthNY
ZXj6h7BW+a6QV8Yy4meWGazf3PHifLWloTnMEv/TYDZX72QQWSrXq0aC+0MymTda
7yl0TAq/EoDfyCXoY+sUoMxPFsDJhnOX8M/sRdGqscFQjdOs4t1wE3mAyknEU1Fy
30TUKJiAaP6cisYQRLOS62+y7jb3hF75kRikYyR0lB6+a4zCy//VbxgzDSKWYOkL
jZyoRaetxtocCzaSdqFKFlNSkvFYRGIICAKBUf5ydXm00Zsy9F+PUfd9bu3X17vU
m2UdBqAT4SFDq7iiOW+6CgYQ0xlD2HlPClZgU/TaJgEx5wnE7/i/A9R0z96Y5dQf
aNiMon4I4n0W/lDGwZRgU2wY7UB1lIOu8c8EyndWQO/tR+QFvfhUZX7vNLOUzNwP
7gTTTiatek02R+Q9BwcJbNP8N3i89Z+iCF0w8xRPRNlux/tRF9+vxjW4YwHAV+n7
Gpk4LV3MkLYsF3j4dQ7aztBrjH1i1kqIzNvxRiwd7PAY6k10ZmQn825qQSlLdDcp
/qRTRoNEpLlV1qxAtNgYLIAub/ENprmtkdI9QS2eGJzQHiOQnNia2Btvhx/upS0R
7BZZErk3YJf4nZC5ImzoxNTgtJCK9WQTDP6lN/bVsPwnRO/MsYwpFVbo6I1ZDm62
7SkaqtdtxEd3IjKhh3tBFGZ1/lS38eXiJxtVgRgv/7npwC0Xo9qP+STosdgxG2Co
IlJrv5Ilqt+s9erskPzZ3GTHsp/TakYpEhl2M9Ar/NnluSzpEni5QZD0ilVz+nzU
iL8oorlGu6Zpeu7nZo4Pkb1jLVDWGQ18yQ3ow10ObodzkUEhT6zf3y0pe8UE3FWT
AZOYFIqZKGY57dEpZtJc9nslZHoYgGW3tlUjbqQUCErGO6Wp7mINQBxbpJAb40AN
1C8bS/bV+l9ReEEJKYk2vRIb3A4Kxj9W2GVrRuPidkkfsSYYTpcLQMWrQRk2/fyI
WaKpPs+6omF7WeRBAYkLcig7drc0B25XWOzc4xHxxfHMstLAhQLMSKzKhAurgac9
fexJ4BnMvU/Am5nJZY5vSgEesGxhHNcJWmlJsOeXVBKIUb12W1pbz2u1FROlb7KZ
qPIU477XVhOahu14Lh8iRC2FHvKq5wRy1cAv3qAK1W6v3HY8kRiqA07fkMJniSXE
VFfzivFdOGMpxxNYUfvRWY+0muJjITI0Ocpb51AQv3g030HcGCoToPNqlTVdAet2
Y+wPLAND09G+C6l/dlsVW1EZsgQOdd6TydywsuxN/GnSaWYv2c9/dEM2tti6OLVD
tVtQEs8aw2LmpxDSX4objdu7wMP0YRUXqH6cazSSal/81fQMwEWYoU7dr6W4um0K
BamwvpwMWU9l3DYYJvYXqrqFXPvesOJTzUA5YdkElJTN7Z5JEi7DhTx5f2RS0knf
bnnQ23HhIyCT2yH2RvVHjfnCfPCRUa+cLwN2cOkvlSpIX1oi3VMHR7tXlXEmMUiB
zn6XGba7HMfl7sy39YnKtUaMIdv9fs16gN+5LSaBsHrrvi4+FfP4fALtkjf40+Kh
w47vBg0VwPfRgTaB3tF44ZaeQDCm49UG/jUr+9NrvQdX7sKWq0PaYsTSs1/M4IXW
JqUyOhB02qu6zNL9y00tN7N2MQv/46WDIQEAlzH99MuTl/HPiE14lO9Ak96x4X1v
j1sgBnBnS+C9WayApllXUysJQ5FesUytAqb904Fsfvc3oNxlQaCDDccSvrUiuSyY
Frc9VQWw4PWYi5xgL4EolbVZYjHbF26dP+l1qMgWKj+CjYXwNWhMg+uZMEpUUgM+
wGIyd4Gm+5BglfYtKGQazjfUxbzgC1rABvketAR5v0LQZbA2xFk7wJ4kfw/Cj+B4
aBmBoFuZUNfILKLhP75LheiSibh1fCPsBLDZ5p1YHKL5ZOlVtDjGXckEk319uRSS
22MFhn7qR4DnBwAfaligsjdPUjwL1vji8sE7a0RPuTkoM7Cq/hWCUWv39/4c60mt
`protect END_PROTECTED
