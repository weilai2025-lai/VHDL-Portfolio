`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ij0bT7a5rjCOgQWKDkmzhp0c2VSsu61tz/xY9qvrOvHu9oiSXOCwDg4rMjT1rHMl
Gik+9M77MKMcjCv/yfHweAb75lMDykB5RGhlJRPHcxnxCTNO9YXvut5RxsN8tzqa
14K5KzUH/n+b5jlEIwLq7g/cpAaDUlspvXnzVB//5osaNPSdN/hYvia+Y/h7Eatx
n9IQexRdQX2AnOXcFA1EQRj1R+gm9FsYbmXGBQDXkEGKwqP7F0RNVcfd4uWZUSCO
jGYX1DWUN48k2VgXMuJQsrkRhG1gCr/dUnviQYLRIXLfkdD1BIBJ/z98Se9vX2QV
y6R5HNO1TNuqUQ9MV/gKIoeoK8Oe9+45Q+KjKlJ3TFki7Swq8xC9Wy4ItQEDJhHa
8OtKU647IKARevTrb35UVtgZAcN2VCnCtLehLB6UuBM/mmdGIJDsa966yivoe4Gj
JM/XHqc/D9yUU7Uddeh5GxLt8BWJ/fT0ZdlQxSYX1a+UvR9aSCGMatywSoixT0AM
HQGSDlk96pp29DL/rgEm83k3++47qzehr8RLbAIsVjqZwOUm8CH14zkRw2M0OJjB
Zwz249/0rG8jTPHpZl9m2ucz9X5Nu2iM6aErQRk33qCWvrIaFfam41wnhZZUzqQu
GE94MZId8LppfHYrMA7QRIgSEq6rcJeH6fx1q+xzYR4iDxcKMULS7jFMw67qCtF/
ky3hNgcKfu9M+huITXSP0QAY7wAIsknDKkzpGiJZd5KkPSXgVM4/f0DNTqophs8i
HCH8pq0EMZlcgAdvvc1ngPmUFwd+XNI6pMJtMDFt5rIudPbI7tZcSZv4B2ud6UkG
1HU7u/5anu2Nfp9UZyFLhggsA7wJq+tGE/DPchYSeVUpA0AgVhJDc/6vcn4JX9BW
6LCQOmGVutQ0kcy6KECCL+IXhWpI+/zC8oZxNdHonfRn3pyPOQzuZ4Im6aqiFC5C
yQZNv66JJ1wFxJBI2OxDP+zj6SzV6vk1hB6XMt47iWAn52fsBdNH1DkiqV05UkMV
b/Y5IgKGTmO/VOr/t+/aVhRfgn1KZHK5JCQErei8u5MVpOjPNQRmCCpLW1Rul6PB
2k6HW5v24DofWcqFM7FEWrMVIMbLsMqdNTilFjQIkYa7WuVHFROIqiKbh+g7IoW8
p+aR1gdzgzmrgrktPGn3NKhqGW5ryuijA29ZXkkDSHw0TBsgIS61HF+eSLoK4Yc6
5cYVTWHMqTolIkrz2j2xBhR5iBn5FgKWsRB4H/em8BUUVZZeGYOEuFG6GTd6FAbE
Re7nqPyP6HolDZyqG3+nLVcMAamsmF3fOqLWoxoX+lKVvbiDDsOSBdPHJb8NZZVT
JFUSuyao7THnSIOX/ezKBmMjiNmtW1uTVzUbf7XhsgxdhYNl3SEOlKCwOR7YdR5E
63QtwTrAqh4kMPWI+kmwpffhYjzrtMiu15nJ9gS337BArPHmZwtf/PlJaP6iPfjg
LXJYa4Tjr6HgAqkN2rCX2bzuNX6/diymvD/oVviUJ6k=
`protect END_PROTECTED
