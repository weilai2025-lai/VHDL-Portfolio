`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
00QUshye8I8lrduL+k0VSK6q2SfxsqMgoSosDVazzii7WgUxda+EZBm9CueSw1Vt
MCAhEguhz/IwlZw98h8t1zuywxIX6cHEWdkwwg+ptrQg5pHmprdS4zHSuw9gtwEg
iVdtRnYDQbQ24dvJNXhSJ/Gc2sBtP6r9VzRxmWrh7E0YsnJZblFb2KKKWmEeJm91
vqnHlkzTsR0vcSgfmQdBmM+qoZpnEqQfV2S14wRmbGqSthvz1Cdi0aCZ+601/mOS
RKQ0kyzzf3XbWFGuf+VW6WKxV+hzQWcK8kuKFtzkLANi4VO2MvVLx57ugzwu/SGo
zguunfh3jx4PpRkaKD4F+x7GI3Vsy4sD74WJcX8hD+Jm4zm87gWgYFBerAFHAJhC
y5r2hsZrdypJ97yZqPVQK+9d2Dbi3B0kzwIvwDxQFKpgHy2mopi61NlqgMKRpaSY
zPlTiW+3QVK5rbNtir0nDltLGsKDsi1XLHEWVFof42if7NP0+r3dviBzqf0TyZYy
hjuvFEkPi0jXIBqljGrfn4tZ8W9D1mHRLsH4R99tpZG2quztUw2VMicpWAS+k2+L
3dYYrwkdH9F5go85DYrENxkIafHAeNhF1ntgcs3TMstO8tDfqgfTClRXdiqtQ02Q
KeUu+5pC4jvosRXRnoRFzdyY7P6bSZSV+PJ+eE5E/WYcQdW4wc8bvAhrk/dVF0a0
Vs0Ci0QRdGvn9QQIv3xsN09mR+JmgQuIeQbATAgcCoGQJxmNdCAFCyLFnyGc4Mfp
eovAiy4yMXazUuj9a3a4GcodT4RbL8rN6Ti0+N/ZwaL1pIrba5dcsAyUKCc5xcN8
KT7vJvd7W8l0WDiLK84/R8QOo4AZ++rJYCRlsobhmRTSQPa85L7v1e18cEJ49d7m
qxpGzftOx7Y3WIqGbCHGkaRYdLQYB69kOvxoNjPHYneUz2IM5eiOq7GAH9qfdta1
2aMJ46pN9TBWKTwAMgrq7AcwJMchBW5lN9C35xhnJ1eSE40WPR8PM1GKz6h1Z0V1
/pLROCMrhxFeBE31VQ8S4FM+SIjQfEypfLo5dN+vbTuQsVvcmZyEra9CVGqiIMVS
vSV8cHaU5VkAhqJfTQRN8yWVXpc6fnMd6/xajgN4aJ2cxrubYbJ71zdG/bD8TFnw
kNEwK1zMZ+EHjH5YV/B2aokB0fRtpN/Coi49A72l1KbwgXpvHkvo7QwKgfqT4FxR
Lnm3EzCUGq2GJu/a7DKD0Au0kIeNNDJJDNIpbi9MmwO/IQ5vgP2Sf0ZxsMul2qrw
UkiNOEKDgQ+de2UtV2/8EInPd42sIvSMq8KCTU40sW/owG2/tzwBeTlit1UqbImG
znx27JOhemWgYax6csZUV66NNXfKryM9olDqmMatnw9qQbW9v6On867yKoXETG1Y
PcI1Im+pj2CLC8RcRR8278gQKjXHSMH5KLx95eOBzHkAKChGjpMevsJYJxLeLPWh
wfXxETJi8cPMuNFqmeirDOdUGR1s0wZ9JD3WxXMj+AHGl18EbAGKtoWDbhbpzXRF
AFfePWHva/EA3lSE29RPAWVRVpIgkGjZCI6QN2EgYFMM+PVq24F8epJeLTgt9sEC
noyrWYdlPZATjkJOLflO5kbxoEbwK0j94SAGfdP7alNhwBmGt4K6ml4D4WUuUBaD
hRvsmSOOL54gTzBx9US1NOXQ0e02KSn2sBoF7c+pM26MsU/bpPtn6eGtrmzF48ZU
73U3YphtQdcM0pQmkeoCBnQErAN3z8dWr3jaPK6Z5YKhF1feOO8gfLoIpSfGhERV
JIhl8dlohx9b+ixFRrbCEOOSJljezkkrneLZTYzjsyQ5T+hCIEIQ0XE1V1HvKp4j
dSejVdrSjj31nVZxONCaazlORzgaNTJQfeCuBeyAOT6km/SqKOE500uWdyXPVjc6
qi78C8gpqS+YhqjG+0JDIqQK5GHpf85c/X8aNCaQmnOv82zRVlL2sdbfJLZYthmB
Y72ZOrQjBq7S9deqi7hyAJ1chyBj5VKzmbt5gzMkaQNclQu0Is9f6/G+9PClPR/F
eNrDEWjYhp7p4AeObUUGnAA2xsugBBzu6JCAqPx2laBgnoNYsJCoAaWjBZTj1NG1
Ku+SvUibwbGeiSEmZnkjGKdE6EQ7GC+RyB6w/hsHlp5s0uJ0Y++vZphtHuRx5G5D
rViL+zsy2kS+1NLxlW9nkvelcNK25QkBeD6vSeWQI/lltTCOKDj7kqS5kzKAhVWb
9hDxGYy8EJt9/4UXKxsQ7K8B5g0xAFg1WEJ/YR8azkgB0hyzw1DP8AK+RKmKOsKT
1k7W4AR1I5mJRXxzjMi0AyxB5WpOjKo7Tci3rXmzlcNEY6rTcTTBgjyqoprxrKpd
2u9S7lFJ33sy4e3FpydaxlLMUFlsI1QIix0BVl2uy22OGh5YR1NQosw9OLLwvdGT
381NOWO7CM3iPbCwWG3mzCEdxMOyPHldr91GDdT0H4hcln5YNYCtmrrEU8eJ1pjv
5OX9KGVglC9Ww8WCX8hgEtXzos6KIYRpXkhCJTfEXd/sIivu4vBRAgu/o84HXx5y
WahpSKFo40hDX7zX1n2M0k10mG5ernkdDDOvAx9pi4us5sjECuYzyQclEpSGlMla
t7HpQYsiMeMR3U7Xs7ZapiLiRZPmUGzzQmGadphua/scGZmHs2G++xrzhcMYEnTY
ivHozxfycwhpbvFXBJmCocBYaDBYbAsEwI7VdnF5bWh9hgDOJ1FwwV5q1u6Jl4Ad
esJnktQ2JLZEgcQOwuZ/9bSw9e2sjlhbMc6wXM5JvJStXIzMDInKcJ3pJmIdjqYr
IrFk5FFtXd2uSgIyTZCAaAnnFFLaXy+PBcDNJTPa7Km+hW+uE/CQVvbVGC45pYrb
OV0a4P4RTgstLuKRoG0NtjFnH7aYiUx2Bq4pqHcTokapALgAYCehzdTRX2296BPE
/r9aZaLwgbQ04dzLBwSh4cU9B2p5aul085Ck4yhPmnPParg1ZflYqIAhOScYJ4QP
QQ5thPa//Npku4bzzu9xhc72O0WW6Ey9MOSvOj7QaTkoGCTDdBzDvb783bSlLIIS
qhwDyfuF8900YxO7aLC0aejOH3/e+XqcCRVEU1Q9zG4uAfwfLgBRCvlIhC2j/27v
5WIGMJGyD2pj5H8re9toiMb99ihl78b5V6qVNVsYvChPC8hg4A5M+0I3upAWspKp
cYWR17ff3E+z9gb5Fw4qDVkivBasFpXQZ4h8X/GoW2eZ6TzDDvMdQLMpKLpyHsJO
/2qaluoCEtBPLJ8JKE9noMZ7L9DsOic91EYmvpL+f8BGVwJM9xToylGztgPWhG0G
Cx9HGURAsHAmYfY3GFKE0X/WTlxuNpL0fJYDcnIkn3iLhcMJmr8Edv7KfRwYT/de
moOQ6+kKkESkmveW3FpA0DLLwkPww1jjGHnareyhA+cO8U0ijMeYpoAYaKrnnlaj
dEOc08PeDkY2k/gak0ofyE/J05GhgZgx1kkdTcgjoZU3/SO8f8woRHSiJLNOn5By
KVzhm0FkPJvKF06XjQX+QHhAw8XMseHvbZOeaAwYCzF6xTaOg/DS+8AImqqn/XnS
HX1R636KLlfFEganU/dQVq+kx5xM/rDkV5dWOXRMY1huwE1IK+Hkhln/mExgRKCA
ax/B03Lc4YnkzjMaHQH/fiubfPx4y2ktAMuK4+8xIku9ctctDjnlj3LMdiExKu/H
nWVF1oMsU1iJcqG7Pk8vaKv7WLoBaEvpqJXFXJ0uFYt4RnRK4cVx/9UySlb+4SW0
IOd6Q+HVNhqa94M7DoIs450OL6P1cQ432rU/gJLa7jCWon50Jye9fcf5Mygeu5k4
HHrHAGIHhonavrc6ciaLDMB52Ra6CaFB/g3tiLmSCJvZgsOdAIx12/R28h3FU0Of
1npW5cHv0nU9SeeghIpoErPSRaQnT67y+MeMTS/PLwkPzk2cgIqbrOOkXMXQm6Rb
Mm0vdQ2qQiGlRG0x/co+YvssFGJPFAjspifBh+BnUH0bmfTOC2tyRTUTFP0Ypane
+n0wHRvl6Bm1y3AQQqPyW+b0bldXr0BcWGw2q6TTqR7Ul/UXxvpTk1ji0f82vH9r
3Ef1Eepdd61fnINPOKNxfgZy2+5YngEf8akkd/4HtCGgiNtK5zur47oOeXwMw69h
lxHhRFeix1Tcrtkh9x6i5JdnuAX7J8xviFkty+MhB86deIPHOsZNLJo3np0ka6qr
qqpFGUDOHmWlF6wKrS3gtTeu+lb6TZWxzXmt6IcmS3qzfHMsIVbSlDzmQDQZVpIE
Lo4WQXr604U7mBFAN/9+142VytqexBNvgiWU9+JVKgmrvWowtgkPToGMJAWkJ176
IkFEjtyGVsJaIozpkwEIIpZw21WC2/N628LVOfAM18qFn4uZHm+GUM9i2+TTWWFI
p5pg22/ufxvjTp5eBld5zSWDOTymWMeVXKtLXPyTzKTcc4B3P3mdvg55Qxg5YRj+
mC5XNfSckEzNREZUVopYD6kk7WyJfnGMaqj9NH8N4rihGzZxu/W4dctPmxFtiKxU
oHNu/ANDBwVK219b7IHDruuPjAZRqBbGmIY0HZ3m+hZdQGuUitk4iayWbOO9jmey
Q9wDWHeuPu6brT/ilJTTcLRyywjrx2APlRC63mByJrHjUPdbEClnmLNLbn/5eVLs
Yj5sy9AuzIu4w/sXXJdn8QzbYyUDZq7lzhZSQj4mTpoNTIuAPsSk4NlHORwhOuD1
LVHBt7T9ISIXvSYr7f7fV+ZJSV2kDysOetE8pE4QKEGJDQuskOvLrIq4FKATDDrA
6JbOq3tTBM4oa76jgFyxCWN8knwvOJoL3t7VR8Irnkp7uAo4rgUZqnT6r5et3uys
ARm/y904gS1jjEAce5eu72JAeTVEg69VV+/f7pZPoRHBNWVyPQiOgSQok1aFyVQe
o2xcUuNzRXVNpwxSzBfdJfO/BhoPr1CctRouzvMtc40PHflvXjFaMAqhug9eeHH/
YHGCL8R1nOiFk5uKu3kAxiWngJzLcsQM0mC1njZL1UDp7aUAoQPGSHT6RJ8ECSvA
hkpchVbTdTSGfAKOtv6pL422Od7JV0T+RpO5GmXKUMdttSFwGX7Ylnr/ZsZK1I+A
Gsu1Nu3tXluGIit0Wq0epzXOVIzNISEcvroPq+KBXustXUNnOugEHkD4cG+nwn/y
EL9iIb0tBqRjyAPYNQ88gHpyDKP8ps7LykzeyRZ1dBzeSOSqNE02JdId/V+BYZ4v
0qbUzWHsOzuaj8V55hcIDEB7CJukRMaWcFxArRkGyid9LVkxkc6FcWqUs2MwU0Yb
ReuxokMSlNHj7YbkLODhKImjucKgo+mYbupwMXnzmp6EvEDZCiAiWLfG6yz4WECF
wJaH/+ClqWFIQErJKlLzJHlSRmHPg7uPlHPuqva4jfZK0jmwUJbvU6v0UReBrBZH
TzjambK0iY7Nq50dRTjfDqQtoTXyhyzw4gRUW41o7my8lcQLFXS/AI1dI92kK7Hl
aOUnG+666NrB1W+TieX1umomiXLqLnjzKN/0U6emo+DOgUAhR8gUKdgZkQjS6CjD
HAQe5fQWcHkAxku01zcr8GEiKP48t9EJUyRCI0x5IUGlo7MRyZTA38uQ1mKzTkOp
xx8+4Pxh4yQgqfCa10/CeURFUknl6FdtLwIa14WEtcv8/uc+vd8POMnKEx1j4llU
8U9UdcvFQKlJrdkVifM1utIz99h+n23XmIqO2jyVLtRGp2XeH+F0wXeC5fU1ACoa
4rvsdd8FRrsPxszQNSn/CgxjZRKPUeaEXHJopqDsTYf2aN4JhFx+Qjg8Dhxg+E4f
ioHXyN3ikrxeMvPBDL0Y6Mu1lKbfpaIbFgcnSR4LjoPHrI2ZRZ2B7R+pFXiVkx02
rgCGv2gspQPldYS6Xz5sRK/kU2+1KlaFi6ezahySBOILjpmV+RO/ytUkacRGQnlx
qSqTiU55X/6s2yd4MzZq3CR9vuAwfdOCszLKvg5ZLhTAOh0+pjbUDMuhFG8gGT/U
aQFvFdkGd/vSNS8nN+blEhnxxVo0vqSpRsVnZ5mZHJCnYa4n9hL0fhbwsGbfQzBW
pT0hlsmpthEDaF0hzm0Bw2cRq6Y5roqZzAKR0/e+l4SEwUd1ChYvQp0DzIaqXO0e
3WYmjmFVy6dzWnhO0egS1n1VHqUSMI4WDKSl7wVYM9YoHs0TiEBZzgGBeZieK8+U
pBP/aj1w231qMEcUt05OLarWiD+VeHi0E1hduZ8PuQsHL3JacgzRMxTva/4wZsrG
DMyxlIYLKCZ22XGIwrEkyruwYffxf6l7R/I00zOjKmUWNDfcbvNuowfwAcC+wL3z
lQKbZLsqVvGUk2+6jkbjgzcgsE/pNwvle/uNTYo4s510pqU+5vlACCGHFuJ03sZ8
VtglTf0sxhjhCczuvauz5XqI6R+amtpF3nnOSZFYyWqZvoHp4GarvbcAO86lXLdB
rY6ghNpqVLRraanaDaoYc1IOpwnlKQJh6diusqvhJK6j3ZWgZfS73xUJXgHoXZoW
y9LyDv6CMVw8C+IAUAV9xzWapNicj3/jALRleTF3YAyXxd2XSvGebNo3MotJrph4
CdwrAprn9X/PdrI4TxoI+KAtCyAKfGdcEE4tT5P7WxWdGp2M4ghTAbiUFzLmCIO9
Jo3EO868XlrGUsU/WHyiDmt10SFhCbeV5lUJEMr/SWqpyno/4SH7ZAy5h6KmlU4g
gmTmqq93Jz1Xva5vSwl0QZ03eAHqky9pdWBzK/izuIRL2jMHlTjsSbR1lhiA72o2
DKHPXo3pq8DWIDU7ERE2yk0UFqmHEfNEmnnwLMfH6pfV50lVPjBgW3EfpSscam72
JPxQKY0uQ46qRst9VYnUTQLHES1pJazL/3hv9VXCFyIvsUuIr1aEvGmEJDsh7ce8
5i1jB1AHSzGC7b2/r/aCAarw+pKZHDLG/FsMHJx3n5ByT5t9+qwJCfSD8h0h4TOT
toM2cDAJIt4rkNeEfq9eWQp8MbInbwOv6+uOQ2GIpB11lp+btFcGGHmLdgCKtBHU
2pWZ8iNKKH9Q7LIN4qX6U5pjWoRzNeVfKKDELlffwTMFFibmSO38++FXqoDnNg04
cPlGhqynWAFUt3eJANXyZnOgtd028p3+N+FRn97EWYQ/mPPNi3EY1SvoUwxdQqHW
dxrZ1PFc8pflf/Djmw5eVGYRsUbB4i2uufC9lHPZzYorGPAp7EPthFnH6AbPJL/F
QRbXnXPg7ESDYUrXu1RNW7JDwotAoJVOMdQ1jhrx6ErXTT8wGKbzJ0aCNuEto9yv
y23ZObJjNTLyRqYo/c8Xcyg9yg/dl7JCuGD1OtkWV3alTaNf+rP0gOXI92Gk/svZ
ibiBvct3PDftl0BfsldCDWo6lWXiVAjrpsyHWO1Wfg6/6yaV4hayGyS/yawL9Dbc
+Xq00UY6Y5q+nZX2jJP5d8xHPA4MVdfVF+zMgfjKgAvLx3RvIy4gX/43FiYJXsbd
7ijnlGOm8yalfz8xJwivK3zK7VdnlbCEvb25TR6pvOcy5VCd+25Acjva2hMMWYGI
0SoUUOYfvkjcfuqc8Nl89Ii8kOJEOtZrq9enNVCh9m4y8G7FprH+UyG7iavqSKMN
5h6mYeM+cQS2FN4KwHfXVwkVcRkqm8Lt5oZzj1p/D7J23NIae2G/jHWb/4jjSLU1
jMf+s7homFAVf4PzC62qDrqFWNkBXLAV0rs4adjXQz6HkE2gihdc3BYy401wRRnv
apjVs25zWPIvRag6yI4ITjlBjSCzI31+0lKV3wHtnR9mg6iwmmQ7bvRg3vSTLxBx
skDUBK/qE2Anm/xFXX5uABmcZPclt55BmzGQnQsmtJM0xUu8ff1fJ1C8AMGpVLf0
jLkurLRyaxvILzKj3Tb/9bWSQEXDY0i1TFDwiHE/40JY3mqdTr2PRakZjRMGWgfi
rLgKcHha9mKUhY+23VeLEdqw8mmg7po8Zv7ticb+GLN86lI0q/d1HqyDY7g4ztt0
kgLDZCrGaPsgdoOlzBt4mon6g+hPHLCWPAspCj/8WUJYBqL7S14TkKOsXd/vycD5
VNP0IpUUZSBquNylGhR4ksy2QCqYfHeDww6KAkuBYlZil+kUCECkM845KEYOkHHC
gjkTXJcZrokmTjdUFbyfMRb80HY9QuascyR8JmtjkmtH2xSzDV8PgGnWGTfqYDbK
xoHFDjHSYZ0c9Qn/hosX2n/emC7T/31eIz9K3Q1QJFv3Q8UkA33u8vxyUaGmR4xE
Jfc1fXalG/8fAJg+/S5zmibSwIAXBCI+8LWArc0XsdmMif7ibn9ybjrj4QasQZ02
NxRi9i+BWsmfIKF990lcpcuJH5E1q8eyBVbJ2nKWDpubNCCBfXrsUuIh+wH4v6n0
U9DIK4nu2hKvc/8O6t6Ror6Nwxj+oGvab3m2VLNf+fvRzYZXm4YvXS8m3fEGOcrF
2XbRBp9003KTz6fU7fn+MXWn2T8mVl6Rd2OlJfC/zJWt4tx5HLmPUtHylqOpe5AI
r4lfs5cMi36LjaxLpPQCD4QUea49a6Zr+P/DpHFgkIRWbi90PLyy1id9lQzQw6JT
zyNpF/afbT0dKI3QFFAn1m2Ag9kCK4PFuCL9dGE1/HYAkzTzC9hE8lKwM5BFcQqM
nr+zyEHrOgBCWktY4d6pZ28/r5qcuQJ+pyPGVLx4BeAMiYdO1gPWi8pYsZf+TwqU
k1Dv3TC5XTK8cRMWUlxLqvF1Ihbckm9zrtXPzFqImZt1BsL/Ln6LeBe7VYyoOQTf
WBorzlbTl2VVyNaOfi6TGvVInA8PpX15mLkPmEBQMCjZLLcfjw3xBLU1/Wsnlhgu
2Jkck/YXB6fZW2+sLBgP0rkqnT3yGuy0FKlD977GhmIrVqgkbGhYEY9Sq5JKqiEM
1881mSsinb2TxCb8t8pgHQGy2sfDgxOF1YhqWYTny19cz/NzmQtfOBbcIQuqJFbz
I4Nz1NHMztqcSgLbSAnJuHcbGVBB2O98SNh5j89dGucqJVXN5a7+OhGEIYKTrH41
S7V47QD2o/YfC6sJ2TlA2Wlu7a10wyGa4McgHlN3NXJkopDEj003B3/8ecCoaCGM
asKGyltMONF6AUj1GLqRXMgCjjgKVpvHyzhG0mFdfmdhcWYkga2zrsjK6C4i7/rt
ECW8ejtz9/NzZupxozM4zGmaG0TCg31NUf+K4M6NR23HrBev9jbGx98WT7uISck/
1zyAzkX8hRVqU6n//uNHt3rM3I1vyi50ST7OL7qkXRU1p+dhn3dQfHg0DIdhe6B3
O6LdfCxA1Oe9wE9mNjN9rBnvMqeVVvtBM+4sLfczRJGC2ymX4uWL5YlBU9YFu/lP
t1WBr3Do4acdSze4iWnwmSg4Xy8XZlWy926pd6XN3QTOpKH4D/WD1GhqBuUR1Yvc
beANJQ/bhu03YxqkiHWNV9X+CxmCnt/CUx92vG7Nq8vr8uQLwTaae/2tgFp38Be3
euDiYsAPjEDM6RjahAyDM4YEVbuCKb/Ee+qAgUZ02ctGevitCXiWRiZF9xTuoTLT
XpLXnvpI2w5rzfzkON8RYIJE1K5xUl8EVPKzhaLY0UihPSR7inlM84PcGUVOub/S
tKT/R3zDjs3p/frMHir971I4+RF/kL2zjva+kF20EAn/MD1kzfdV75wYt5c5CSGA
XCkAXFdi05vwwt7qF8lCncEvLi+cutTLIAvpoM0iBubLI1+0HE+ZsrD/MoQ8PByE
6+xKmlExLmXL2BHoL395Fk8ko+cRTwdMf6BVwcwbu6M/kBflH7AEAPJaX7QhTk7X
e9QRs07RSZkETaVH7z0f42s0nXtIFJT7qzlhMV0bFZ5Y+L0f5g0hvCmxxK+lEt6h
jDLLRUKtB6zh7e3IMkBpnWre2UhHC87GoDW4o/rHtmxvW6WcGOJmgO7uyWYq4jLi
o+5dGD3xMa3/rRw8FcrQMFi7/r6BfpSP4N1z2He52TM3YYV53uWBDfyjTAZS/Kb3
UC4UpPHnJ7t8xHDUVjIaVucFTsQe/htSR9wndiZvaSx0ZwkUf9XBGRA5AS90FTMc
OG+k3wbhfq81xY6CqekAr0MPlX5Z7QO/7jLF9YWVEzkSviVnszH1V9zjaF59Aol7
kFNv4JBo9+uGOyWWx8OIvQagqaEXPvWyVa/0+0hvhYC0D6bpb52EkebhZm2dr/nA
D6gyEseXCPbLI9GsH5mU3s0KaYkvxlX05P80nrmOawOxyjgjnJcNztQUMfwDngJj
lkSy26KL+fLdL05qT+Yw0XW49lXUsz9+kxk4nxCaNg3wakqIIgAtCcUbHqlQTY95
E843+IGbTqzwaf3Bla7nuWtDGoZ+vKagkSWrKgkdtQ/y+AYwtab2OXT9WGhdHP6W
XuEtGH8p+35+RR11t8yFu/EkfWw9NfkM+4AT+RxpJsTjbVWr6/Ab1R8zxrcUULps
4oQPXc1GtiRN3nBPbwft3Hx74VzZEx5+NEhaSqL0fmwNHhywV+PUDamXx1YKluVD
14MaJDqf1Y7jfBhZNy9jg/+fmR4a547zMoH79tQ6+svNB5FWeR6PkEMdZAwQXjHJ
Vzb4vTpau/7WQcTVMDcwDGSwvl8Gy4OMe/UWLYLH6+vHxfKn/53gILrT7rnJ6fMr
o0XcZxlw9WutpXQcYwOrxfKizFIj4A9U0kvBlizBjlLRolMbRhBXNL7xUoJ/Qs1l
s6huYMcPXqGSxdF3Vv6zDCdGeSIUZzzYz3udGmCjfnKBASEaQDKKxx0zwQ36ZhYJ
BfS6hLrLZuCnc/JbCpncAlQhUYBvjQydklulosmaqT6I9Re3oFw4PFpzN/qXa1fw
2ETsJ0AxUZoAb59ethcAMjSmFRQKlELlE++OVPJld5TueEWXAO7agVKMHZ97C8ik
Zyuz3KOmzNxc4DQZhLkMVQXZkJ2mZmpxUs3WffCjUkkZ85fTqLsQjdt3UOygLAt5
kE9Fb5PPxbprTftQPlxc30uLQVgbnx4oRaNNHyUdg8ALUYxns8a7aH4GxqQKJl41
vZEZHqvk2PgZoujKhxFgZJovPa21SzqerwQBHFQQeSe4seOgTl06ylQVLbsghl/s
HD6NP801zvm/Kj77NX/tTBj6C427XpgKCN2C29JxbOR2rCHeiq5Vc8zn5pQVP8MY
gvSBSXn2xkbYBckMxuCZLk/IocpTfcbP5deaJELjw4sBIUtZ/NXK1Mm+O49ZA3Ud
He9k/AHfpCp+Uxl7hAt15F5vUM3UxNchBlgk1THgLJmeVfsrlEIeqGPsRRaTxX5m
OCrWih8j91zOdbjt6T4E0wp7RxCarjLVHJn/M3dYzAwy0BCbGErmODk0hVkKDZr3
5lgYq/JPl55aIidFK2caQ/bw52M8WnP8BnzDu99RinMuSIKVFQ8EO0bMYPC0LbiT
xF8Im9pN5jTZm1K5+6Vnb3bkM0ZKet+3vzjs/RIadq9vnbYTL3hEoRiu/e3nQYfO
PMxudYfQY5RhyYddZ6L61qrn3RI43V80uF1QUSIsMvb8xwM2/homyTclcJElYone
/KgYkCBa67Y3R3cXmLNsHhlA53f3NVDP3Tsyn2hiTNFgrVQhzeaV/INbrpEcb/VP
AV5DND3QEhHYHy0rl9eaIdh+gkc66PDHu+n9cudaoX9tcu5RhrKITg8+25n5oYo3
UpW37zdwmIFDKaSkM2VZksulDTTElMWbQ/nQKaSIuD2HQtHkl1XY1JMYhiHjp+vz
2mX+338sa85llvo7PX6lJe4hBc6ul1cfCFnD1KaqI8FW2934qeTaDRcwQP4kdv2g
XU7UXN9WVtS9I77mN3kK9kT5GqMl/IplWo6VtHTNpcwk8rWD66R6LdqheSHhnV2J
r3VH2H+hxIogF4w3QwZK9JM8sdJ8z7h7EybWQ2iJy5uBA4CN3Aa9BZQa8RggKAPe
4DumD+N7X7lq3QEl7zTU28uDDY+Z7O3tZYDItCGT2JD/SgX8xa9VQZcNzd0pMZy3
DJJWrzLSUpEbcJhJM0mfXGpfClInDyN+XXHqm5iWuQgeyF7kpSpI+yLOJduidSNb
PKQ7JfokKYz6CWPz3+Q/1QVqZfVxzP9KCIuhldTJUwsmNuzWhZa9kHgRV9a3/9B7
eSp+a60MXWnT5mff4M+JAi9fz0ECS7TOOXtA9lNiYp76w6sbE4Xx2/Bo+dbaameL
lzVhRHoqgl1Do1yczqWwv9uGN2B8pF3BDr6eJ3Y+rq5Edyc2ehB1WRTMeZ5O7gA1
YCnD5HQK7iX+bmsuucvQszpmx9bcZ890HTaTTYqKqX8DSdvwRQoGY3i0zuLjAxOx
UuUtFckUlDpEMO7gHV3NE3dXTmt8iBcFW0Ym8Dk0r8RN0gGt9XxAWpAlEU8Y40m5
l/qoi05K2go6j2i3zc0D5xqWsESiuLfi6MYnyd5uViLySWtyfy9paYRr72o5qGQ5
CdQih7zyV0CKeMRlG/g1d28YjmEAkpWAnSf9CBeMzLLMD5oIfVZIcbeZ9enwGXsd
vJ7eSiH//qn5b0udnk20GrHfSap5Kt+KUrFD2RSUAYcymdQZ36H9yKP0t5lfwBX8
HTUfkaMnmoGvUe9dvqS02K5OC8o7GzQ/9TFRuZxVwo1aOSISR1+8XFn3tdfqmJ5+
OkpWJjf6XQZjrkm2sdiuo04KsLl0gInunEn0enAxA11h82TeRqeIY5IestTMikjD
OxS2Qq+y76wYKkXSzEsQAnreGdAHIuuDn2+VTzV8INTWT1Oxm6YFqgdbFpHXKrIU
oc4qkdVIRIgDoe1LsVHmZDrXMnuMVUnKskoI6gQPnvx11fvpeUlWg4c6W9r2ZL8u
aPzkc9Rcx0/7I5iUHjFvMx7mzSDeNmrh6Xg/Oa0V0+PPL9aBO1NJuidnOtaQkIIQ
Aknc+Qaql8k+K3pXCZv3FJtxVIxUdap6Bo4BrJO7f01vMyU/By1P1NhPVU7zrO4I
g8wjcdnrIs5CEyEA8h8g+/Kd78MRpAp4CbuFvJcDg8+RdhIBR6XFpo5q7TXrNXcQ
Dtec/j8RX9uNpHiu7CN+s0qT5WyhAe9Emez2hz9nGrZMLlRAXI5MYzanHyQqnH5t
YGJWzB0WMvKY5M7T316GmjDcAaw+jv50FffuqGJLv7tTlVhbX4aQJyOSS9eBYtQU
NifWvvq2uy/o4M79XDrOq1gTlFCDWivYzFRn3LO6ppWeL7HiOOoLB+gz3r7sIYw0
LT1IRyE8U/XHX6E/KcDHyspheAP44bouH2XYIhp4y9cYF5S5ZWvDeM6y1AXk0Xb9
HOTbUsnK7NUzqbpz8uDRS37zB3UkzocXSPsUUSVU73mb/ekMEKYyeBlXowmhXTo2
keH4G2D57gh+Xs7LZfiQPIJEuKJPqj7hGLweZEnbpTKMRh9qYknXlFb0nOs1NV9r
3W8C0sIGtu8zbwbbMr/iDVLSdkrPFkHZGizHFsksL0Efr8kDFkuAUC/17tmNQPW4
Fl9Z/h051QeIfQ9WWNan2a1FDSun2gs3JIVB9M3s8VpGwVVBtuk5bZ7fcEDA+S+7
g3pKE7y0ghTHbKpZT3x9JxBBXWxaeZjv5DiE7A+YEqRji5KjRr6JOSDeIo7TphDC
MnVDKTKvLZWGz8ND6JXWQni+WM7ei/44v6I/kbW98qcZJwP64db+xmDm0kcxx4gU
s3vxT2ZIMCKRPXNDzC9byBvOZ+mpxKsnBxduffHoEcAUA79LvQcLA5zyM8BmPMtZ
dpizU5+ordg4jDgEI8pWYSaOFkmPCjmaP0MU7MPGnmw+e0LTaXFbmlmvuCkF2gL2
Z4dRnS9EfGFNNlYIK641+msjRtNumnjnaRrLSnn5EgiQtywu/UOpnT9e/FW+BG7o
tus6MH0sAKDpWAebsvf/bll+mUebObJX4unb8pHipMLcInVBJ+yeq1Phe3MBKPh6
yq1/KKjSmE3LLqTth9XeSP1MuPF4vF6Md1XrQDOFXtLUumeISxBQizQRA3LF0UWm
3rKKYFep/YxEfWouIvitVsFtqrwabFgKJfBt2qXV+TFPVPYxiSZLaGE09kWOW54i
Bve/8A2xWt1lkyBh78N3WZmu0qkY2H0z6PCG+WE1GM9c9DSppvM34eULSNLxNSeR
0DUuAa5p6ojlJ6mLuQKCo5GpAXhWIoA4Gw/00E5IyQULG/4QmPP3/JXWbxugj70m
bFifrDmZOnQ9UOy4d9IrLxgCs12EKetHq6Tu7EZ263cF9gV71LIO6ezjHWjrt/Rd
2hNi/bk41TV5mfGfCQI02aTE2eG3E78b6PUUwmueajQW26aHjlueUA4uBIPMQu7m
vFW98RK+9s1LJ1bEfQqZl7cjyctjBV9xf+v5+szhlTipgkGpuMLSluMhf1A0pQwZ
9ZeG1DYodzqVoYTBdSaW7kjhi2Da++lM2LtaOnBNqBPjZ30+tqG8X20A88J0KMgR
H06TdFMY4f90neYb0/shUEJau8xR4RKMD5n4ZlkWx+Etz7KE0lSE6plQCv2YufDn
ZbNxN6rp5EvSgIN391GdId1JXemh/8xKfPm9OCwGru7Fu0ib/MxuHdyDCJ73fACB
Bw++FZv3FUl7twHlBvclwNqagzA07MU07/+xbaQk9hd2Bn1/YQgGUNlOJdZuMojq
JWJ9VbD1J1bPTk2oIM3ACksgbtV02/BVKHiGOVlDyErylijPXn1KtC/0L9IWFfWw
ghPDcv8kJwBrrReJS6D/hZm6sDp8f/0QkFKIuouaUgEDhBacyRGRjkmdvT3zis2n
2og6bYK+zh4Jipqonm2/nR1ftOj31gUiS4Y4ZKdHrSbOtRywD4OFx7zoyBC0U8BT
Bs8iHHSbDJ6RKxuLyosPVdL1CKW0KTzinyqU/FEIczBasVtADk0ANcn/PNbMYwba
C1vodXF4iaYkI2IOD/W3GR0Oa7MRg0OGWBHWIngHRPlwNfutdnk3fRe66M4No58p
v6P5z31XoboNNi1c/my/HR4EqvWUsPZzEsx4Rrlhg420qTmF4BkjLvLJ31IfwEWz
lu9ptu1kxtej+84XjhahyvQWVDb825b+EXN+aimcLaB3UWM8L0/PeBi6szzzCUuT
sNgdTIMr4UsRmbzzIhW35dRTYHCpKlakmys8NRqQfmBtuotLafLrufYC7I5MXBl5
TgUemuJGJsXOL0GaPnKn4sMbrfs2UTapmPmVMEQeMJND1ZQ+eL5eP6ZBxgLWPnVr
Gic/+zow/IQXo3Snmw91zkNndsxAW9g2fQs8KlO8WoOOWCP/IyT++CJFYwIktDpJ
+Nnv4t6FwdSiFTdKWZ0KP/BCoaOkTS6ptj8kFmc1VwWUQYONozWIWSuSUUgL4JIB
VJwe1Ktudq6vl8ZbuOBIjNIV+AFsSWU6HdkzckUsUQvlmHbX0WKIRDLLsSPMDFH8
YslK9vySfsTsMS4y/DKubRYzZCjpa68gfR0rIGW9jNmMINzPpust4xXini5Muamb
syc6fn+ziKgKYMU6Qp8t/JENa/9eyICm5HByIzm2tO5U/ZTnoIIWMkfkh9SeCO9b
SZeTcfVzH1shF+rhYJl9oiFFNQNsKZjc3AUryzsj0pj9E0nKVcq4ZVceH2n1mHIw
LBj3T1Kf204Kzvgs861IjzyXNSfnsfA87TnozeweVgIhBqCcZmJWKW/Ej/Giq7i5
1+1NsPLQ8nSnVOVaSWugILtv8eT3en/pbfGak+LccOs3oL2uLLKpzAw2Zp5S99Ne
pZyvkH2OtOe3mfi5N1t5q3A+sNtRP5sA3vNP7a79cyj8kQtQwbCEeDIeoZaZhRKv
d0yE085SW0pN9MzNC6i+1G66g0bW0Asw80ltKQz83P0hJb8V6qMjQ6X0oroVs9ZK
p/1Pyf81vujRLm9KYPlTeSCQb/wln/zynCacfq27BmOb+PlP6toT+uUppDrjr4AW
PDMc0W5aJ5DZSEhwJkyfFyBQ0RzPcOPJmbeUoaV9jcRTTRwf7JJjq64na8aiByMv
oWHqbsb4G5NskEU83m266ohsODvJ2k04I7PAFU1E9PK94sPisEHGq5137c656zsL
WoEs7v+qj6CRW4ZGfsoGeuGe3dJnzUNGhtki/bFqQdaxg4A4RUvziGssQ6YHql2n
usHnOPnVbiMG5AzHrWVj5V28xFjlkCT7XV7MU0deCDvVKyhVqVvT74NhCIsE6pbp
ECTgH661tlZi1qKtBpygLq69DPwf5RL01ltu2SOjIbxDGdvy3Durssq4yGYu4Kw4
xx4HT2Ql32FDCrrnmWZc0nEbByKXqoia33wgu70iV5V9zBzxdJfyDDBblKdktCFS
5zfqYziZ1T1KhqHhkunBi0lEH/7wr/OC+5l6GWa1qP7f/cR0phDrB7dyVLLIgnPJ
WX+Q0UegD/b4CAy44jb1ktBFxuTSi7dst3aKlGURnf9aJt40MmupcghgdT+R4lml
KxM2msCattDqVtsgw5n2IyJy82leFcOC6POrUgDVrC0x7BXY8rqLJOEx4ARhrGNw
qDA0Y7YHczboUSliBpmVadWK3DuVRURQMGXCHAV9v39QU3MvEc1eDVg+WU4M4oX2
npV3mzo7SdXiGfgEVayGv5b3NAnxmKhxXavjMB6wf7sTB0JzkRNlbi2JAFeMoM7w
F7dPmWv+Cvc1uQpjy6kzdH3Cv3UYISKKG97q46HC+NzgeLfXfBEyQcqdNiHFIYTG
kPCyiPizoWbcEROz25vX6v8Rv82X6ugC7oqkEvSQSQskHsxANMLiMO6f572k4/Yv
zMkEjMmnFNqbB3p9LCJ+1knopv9WpQ/w2zxlpzZHUh1ge3Czb+K7kH1Pic91Wlbs
TCXO2CBFDrdbdQG8c/ctusFtWcoVVZEY2BZEt7o9ArAHWLOq/BGFQTNm0YrgTJVZ
76v9vqWYMv2RKLP5ij77Nx/4it707UkeZYAWbYKSxSgTkYvKslXeXnHfKElSZvTP
GAY3Pd5H9oihaaCuaGL6b4U1/1WYuwVnzUnOOW2YahEPyeITG8hCgKREFKqv4+0w
IWuMzCPRSfwxh0SmYfIzDzT71ZAmM2i/6/FghmXD/I6MMQDKKB1leR4nCWfetDac
q+qSxjUu0W+gf4Oojax2hHRY1gBaTS7wvTZlRidT8LS/Nwh6KrkgiM6S2X0HTIBP
DBavcAMDIQVVqSmnHawZz+GWU2cSb6U1BDfJaaNniOEUgH0y0q6Zf9NHqCkrJRdN
4xr38Pb7KlSCmgOcFxeN17RcV0Lgv9TVeNZS5w8UAKAl/I312ZR7LOoLJ1/jnWoq
sVO05AtiB8Y9CJkVoOLAiCNnyLrmkYhWH5aNzB0e2ciOBEXPz38sZov7Hc+X3BE7
HGdtsMpo5/bDuWPsAax74VSeUsOqr5geyVnXEEr4D5bV6Jp4brTu5YnwVctO8YAQ
xbW11QOwt/D5bcXHXlICiu7xPv/SRmKZxxt0N07WTSTQ2J6BYtY+YpyNMwV91jn2
TaWAtm87TkpCAjSMLtfO9xYO2H15ZtXZNM0zHL4nAXZPBt8wPyRdQU5Cc2RJ7H/d
++s42XEESHffRkW5773f+gb0QJ5s5+yR2jI2U0dyJwLuGV19fYklaiW2gjnvfYY5
vEkPvUVUu8VWMPaIeFJPpE5XmNJe3Ug3vebISHQa1lQ9cksK/Y9x0AZ28w88NxDr
5/wH6VsriO3C2iR33X5UAN24AKt8O9oicM+Ih4UovLN3ftdA4NyYDE4BXa10PRWa
B2WmODTmJOJuU+9/SjA+cufppLKOZ/5h3oS315o3ME/7d6JM3diMlAo6nEyHdk1A
m7qmyoS6189wTWsyc1XW5c25InhGTNK1SWMCgTbmuEEaTJOaIkih6SGs2UFB1/eR
0X37Bx74hk64rY3mm/cXTbGHzDgVJJtAradg92rTD4vEWtywfSaPNTKAyXnyTvHZ
HUY/ULWyuBYHPm3zi1Y8s3J95XmsLCI7aO8Iotq+pZTYoxFdk0UpIty4eHNMm+Mj
CulusnlXuzRa18/g5cgIzc5K0Wym00CoVqUk6iiTdnUiEGZy+8Fdt6ONfmAGUK9K
fk8oWJURiHZbFn8l34S0dn3T20JLLJmdH3uf5auAbL3EArkqlxTel5cIhJR/Ks9G
hWtjvgAC5QHyeIqAU3DfOAHw3d7E/MHIN5sThWskFKtX2ycPpTfMWeyg32rF/6aE
jMaEiARzvR7AD923PwF4p/k8ESbD39H2JWUh639vTOT+py1sk87xmwMT9fGsjO2+
I6+boRj61Fa7PFXy2xNXQ5k5Us4MhJxShAeeGqwv9w6vKZcuv4TMk+jTlU9tNAcM
oNaHFC7o5n1SX8FwZMIZF9fKFySpY4xDwV/UPClCkYmBPF+I3hM2O81hARmss7be
JSnBpHULi7Qp3K3PUBvzD2QyWS490w0ndu01BMQ1AsVhqMJgsSb2s4Phmpg3RVD3
NwjLdOk10mTcBSNv8f/3Zy/4eFUXkQ4LR4hDEb/fUjiJM7zCF6jO/Fr6K89XBcjK
bvpsZmS2jfBrYWSJ/60rfG3wbK0V/EtKIMj2k5BsQ3R2XhJOYWSORDcRZaJgFRID
LmjPlYiUSW2obLL9DtKnp1B2JaXS63ysItGpx4Yvu5Dl8CmQI8znYdkdj8YD9Dys
R5tzYmzozsgj9RNIqwcuaIOMgcI8dnxVvZ2pc1p1kus8dubqDXmYlyaC+CmfXJht
kvQsC44pQ1N2KqwM/mIUKuxOHObjtAOgIVPSdXdWtP8JR9/5YMsnQBIsxnZDk3Xv
iRkDscnLr/1RF3WF9z+RK5ni4/oVOqokYeO0IMrKWsWSt5OmYFSpkca6EiznDWXG
2q9DdOtdx1oOFiTONeYCU7E35ktUBbHqClEdhfcJFw4PyfscdchAkZBmmBYx1i4N
/cDlFCCDht97TsRDwrk7De5A4e73rKrtIurq2AmpGRAMnZEnF/LhdGhW55TWwdbn
c3Pm/jLiq4JestSEXgTGY2KL1rq7vWq9RlcAYP9NDix6cRaXbRl1R1eWKpeCAV0M
+xw8bxMiy8hUp/bCzlCPlG6f0lFLxSRWeNHLiathSqT41JxndGasOw1woXvgPNju
Uo4qk3EU0PF6SpGpgeVwJCnF2Kp/2CC0SAkTXRl2F5pOf7XnSCaBCV3IzaTF/aza
jjUKY/OQdRH9YWzU/7sldtThASAsNzYlaOoEWDMhkK5Rg84jEwLoXMVnSxDJ52ob
kQKXmjui23I6UeCd4xUuPC8pgisA4lrghxD+XAYvZ5U69CRvKn5VpIlogn4+ysLV
zF4Wd4CNH0E6srMsRTQErb2L0Z0fLU0Ng+0WEzB+4TGs2fLJAvSZZjC5ky6LZs7h
L9j1+osYQM8437GhoOtPujq4IfWjGCm0YgSLaIsw2FVhkXyIgiOXWCbOCAAbKmVx
Zeo/FJYIko70xgZ/h2hXl0jX0FB/+U2aFJBfouM42CdoMP46jLd0VXGLBlSQLs+w
mzCOV8FcPXtFjUtGfr+xYCYWl1jlzu2FT8ZKvpMkO0HbPLUA5JVdGTLVRLpMFgaU
BhlBsf/qBByxBHTldciuDKXRKXzuyAlZkl84qM2hYaUd9b3Z+gBpq0CAl8lqgZlJ
j+lwZoj3pY83q5G0KlIuYO5NFIfcGnIHn01xvw2f75B5AMNAyLijjUUx49rNs8jV
vG2Hr02ugO14Qn9wyPg7yM7ItIgygW2bCWmtPQxiIhz3tKZdQwEWu92CrOM5Dx9j
QSoJxsjKIssGb+d69tQCPMypD3XLnJGH7sTSuIzraPWMYCDlBj78Cgt8A9vugqRw
+EZcinjIHe9xwYPnYZMf0VF2Qbzm319qmgrMAoZb1eDZ39CFvCwo/kB8GS7iacDc
kEsHQkS4SG5Bh68eR+HY19ao39ZOUaA9/SPO/cwdc96i7OPzh+NYXrb0GC+0j+Bp
7sPQeAzQjehlpK6zvuORlVmf8mw2szmLKtupMP3U6CW5vXxWxN3DzKfIMa27n4sL
UbBpyyGOEG8GkCNEOtNy2G1zI/k/aPjbQFyQ0UqDwpVPK2PSCV0Cbs6JX3GylCm0
ePHeBhT/MLEW/g7Jd0mFnT3oCt+W1gfBQMH+LyAyJssCbn92A+91iF/sfviIPbyf
gDQIOxPKMsJV5g0gqTrxlovYTu/i1wUS3HeUDIxsVP6Dar83GLFFwqy8ZCeVt2RI
yf2NVuVaIEWGyQ0QhTTmAI8r6OFCV+ZKjrWXb0IVBGLDeQdm9W3bY5lre/KlVnkP
SNNNPpLMwv1BdgNgS6c1xIWSBiRjUtrW0h4KF52PFG5UPIW2ZIfqs+uImzUQ2HbD
20348aVEi+hWAqmqW3AHaTcJ8+BBqvkeDMRswSgkLqbWclgU60dV/Pp/tAgJox/x
H+5KmOnWNSGCkQRndUEOv4jUcFUZXFaIHtMsNtMOc509GYvsEKbV6EBDv0N2m3R+
Xq3M3jUg0paRfM/mwH8FZCTB1F+7S8cvuEwN7GvvO9RTtbYe/5m8N5qEZMdSq+Rj
xPmzWQh39+PyTZCmhyxeamR2Jw9lLlD6k3lQJGzJOYwjtOvgNv49pacXy8qyck2Y
Hbs0Oei1K4xrmd9yJERVZkNgeuiaIVOh980T5KYbxkQxWkP9V9OzQT6rzNmuZ2iK
o6gr3ywhVqAuSINY6y5NIrW+ojmQSHCBCIT205PVIGNzC2CSed4KecyARo44Yssi
4V9pmmW6QQGSeHEhyt7Xpw2lXoNY3Wl/o+esXMii+CywmHywbqU8ZkUOAy8ZOyWp
58HE6iaXeFr7/WCc/yeG80k9+1ikdWCfRH8mUE/9obxGIKfJXWlskOspVZi0MNAy
AwUwMa3la/Pc5L1/2VtVus+0QkJmGGmCS2n+OKsBX8DGFSESUI29bFxZhJmldu5T
FWXG6e9KKomUiTb0QTpfpxNs/h68OFXnCxdSIvRL+2KySRWKOY1bbjNY2FzTYEgj
lIr544D1PLCmb4OTK0rykW0JDNbMVrd6DkQPzKiIDQVZmWBHG4IighFzSxurUwJb
1zrjkZX+mRrl93WLd4z5ks8lA0xtwMoMGlSZx/o9gmn5fdXkhESqw0LnLE8Wt70n
DuGxlY6QoeUsU1kVBBmgO6YqhlhOI6G0fWPcfRU+HgyJtbZfjaMwgZDQOU4xQfBL
rWGRmpgaOhC2Ec/GXqAWQd7uh6+RvmDgBOxZhGGZ/tyviqUYgJM4ZaUVNESyHNEN
i/P+I+YbArvoIDqITeuNGqEz5tMkeRAKIe+t9BwWT4ImRtxYXQyb4hxD2IqRxIb5
J6Ohs+6f0mqDoPjwXJ6y587L1zugm1GujbFrkn4QIRgiQ4r6XfMfDW38Rkbuovrc
9eRjYcImQBz2uVKfHISVqy9WOZohUWnthAXWRbaqFMNojev4ztYi+89EV+zgI8NX
mRk7xKJn64SX0ahXAKGH4A5vheLgdsd2ywx4gkbBI6o5AsQsRoNWnZZ2cRHm4QIB
fOw/n4wqdrL80VzQT1+W1pAvBZAwsQDNJlusrhH0SvEXWEF3/CAv10kqgQsFkyVW
DMfeXM4lDIbIagGF/QbWQqPdNn187FhxMZpDs05j/GGjlud9r2pedMfYI2HaR+x/
GGDKrkBjarOoah03rnekWW0/tBW+27gsjHfoPepVcFLCKE02Zns0QQMSfvjZ3kn1
vXZgqr+t8Mc7t6POdYvttxDXI2OIdUHbl9pCakJMV3jZpRaw+WPM6dqN4glp6ynw
TtVzkx+gvEYgoaDbIRVd2jihJP+2yU2QyUT6feBOSZ+UN7KD3lZREWALljc8t8Rw
WDya3nPJxfR8toC6oFIayKzyt+EY19zTn1MSwwKu1+U3XwyYOFk68uiKxUrFDFdK
Y/uoYv24B9U4UhU5HQxr5DHngDePHbttWWouzh8s+fTvfG0vZYb6lfKT2PeSaIeK
gE2sOHgl6jOvKgCEY4KB/eHdbl76Po0cTdRV+TUfGcG4o/Rs8b3XWbZfhUdpKmnx
0xDTReBNAdFiWW1Pt8NAMUg8hzwNR/QQFk0RHZDlLb7t2gqbJHr0MPALfaoGDdR8
40QvOd0YjqyQ4Jrvu2xXaed24G4YdwbA18GDAaIr4gmnwubtQwNaJkZIjrIxVx15
JpyxUJBzL4tSsYaGuqUzsbPdZEetjjcaEx/3wMs8cTsaiYXp9b12ax4ZDye5T+hl
Cg2P/Z0ED9E3twzkPdJJ8APH5JCsK3XMuVTyGFuXj3Rt6EmiM/VCllTg6aZh1Vls
qU7NHzm8MWvf3JJYc921E4OB1XEvse9GaSl/bLkYTN70Q7rnX/knKnfNP3Snuqgt
avTZHaqqKzRco6TRGSh3OMslYhu+oMq/Sji33y3eWbd0saNWFVtEID0j9Jc8iMgH
sjbM82fYV3fLArlChvPlLC/pI7m5jr2FHRV4D6GDCZrFS82iZQa+2Oq8W3i+sOzr
xboQ8bPfWdTmBzWRrXCD+7prUzpc92nJKdrV4tdPueG8Zt5hxX1nXthoTgT/Ql4i
LDGYjYW6dGsbOhw3K0k8b5a3coRBDoF8r9QCy0OT+9TRWofzFUEclfGtiRvv5jm+
lvvdN2/8xJQr1Vqp87mhpIMHJhR1mG/gWlMdHbqWsG8N2bBPQEkBGphHI9f/7IeA
MBwJS0HWabC265mxcVlY1FBYzEwa5y4a/ljZsffuIODCrH52+A16t9e0im2Wj0wj
jNVEYt1Bzxlj4tWMOyyd5+KUbILAQHE/CRSnijFs1kb7qzJaMp3XifIeQ/UdBM/K
tJQOIYWmhsxqBFrb8hRS6BppgUZgDirInvP4gq1onWlSTgDPOmbihn/n12J//9+L
jZ1dRyyKTm7nhtYxMx8C7PJpDW/gTjnr0jJf4MKYoAbRGEhoTfhCYKFU4jpUnXoj
HjvzCBfAAm0QojMRkpdZvQFA4mrELqcI5ON9eU5YflZF6qh0HBcXneA0Bv5OQNGG
h1bCvl9gaiDkMhcpmo+7NCsKvRQWNcCZGoUHych+EHOAYyP3carsnAS3pOpH5NaY
HKO5jMF17TjpNbwvN51+8g+vbnNXHmGQ9NaYLjlXWQKfdvvvuFg3nYAsF6f1Z3O4
M3Ca3R1/9CosKYbRxhyoQHYeEac4lbn1rNjINpGv+MJpvMVLWwTTYd++dSTg3T/S
cazuaEWDnDtrmYfJZCFB5NAa5yCbt9ns6MpK27ixdma2QpbU6hbMol5JWC6jzjXg
+e82FeR2njaIgciOdQPv+Ea0G8fKm3O3PIKzNpTFIDg763E0u998uvnZt4pOVGDI
hhX9FAIQUn3qxSLn3JAaiks4AukeWv20MAJy/IYriGrO86IfKzWIu/aofRJnma5q
yWK+jtMME/1FgRAVlASC4LgQg81FGbWODAbmL+IJZ/GrHBV/6CUL5abcZiyej+3x
cMAdNbfRKFHChBpeY1fEW3IOGZoXTKf89HVPXz54AgKg1nCTVRpoNfWMUmEYVHrB
CM6X5wBwi5IG6pmGZlnlwFaAxiDYkZN+54RC+cynI90BzDKVAPVmqyfcX5eI2j97
LZKfyvVCa9UhieCXQnhAvyfFXWUx5/FrkVHTG0Ho4Re+dE2OUJrtOj0X25kKN0IW
e7zlCD8GFMtff+w51GOEYAQhJPOo2GaqhWJBvM5i4x2iWnp3KDRquwLLT+Ve5pvF
/eydGk4/fyKomB0xBEfqeh14QlWK0rHU8WifM1MzWa22M1C5KwbMM97wcG09nuLP
7eeTAIouCRfARp9N/0zDrJbacuc80sjxjfxflbLscAtARjPgTXuPHTQ2VlhX92bi
kQVS2vrHKlGm6PXA37wUKxnzTm+guB2ZuBsbn/86awr3o1sQlXSpvbAhL4aaMO9R
CkZYGmoBjkVX/QB79ubKfxEknMIxgb4luKLI4n8Ik3rk2+a+Qpkhf0c6e2TxWEC5
A8qWtvs/xPV0sKw/r4OCoyygDGZgNTmbSyj1KOnR2LJdRBDH6jSBdNnrKJ2p6ZaE
B5YcQL+E2xYMKStHLLFb0VFdHb/8rNz7+RBT5H5/J3wNRbs/UvJbVs1JTxK12mfI
wTKiw6V8u4jQtSoKu/uRopVrJasz9x8pf6mAuRj7cu5N8mbHDw8UuR0uqWyECaYi
8I9BSpS/s/B2vsRTnOZU7KoVFUVYuxKe4n8dGtrt2VoUb0kltxue6BI1OWbiRgGv
UP6Th5vrT+Yq0hcAaHWMkS2JWrM38qN6FnL1ATfclgXN038tCnkH2ylAU+GsVJht
BzhRlbmcHWZN9Trkqk2aMXscokjuIOs6xKzmdhRSX17c2xPQUN4r3IPi9sJEz2hq
pKCN4dg1qLDy5Kb4ddikeuM9VNn17Dsu8UoHnsxueMXYM9dpPQXrA+Qj97BlN1IT
VBdipFnOZJlBYxsYUJ9qhEf96K3gAtOAI2mJAlbR98EBOKSFjc7gZq6tWF2t3QS7
J8Byv8fVF1JtkubTDnftuuSkrE4m2VQm1As/208YpIT48VRXYF2il1XUhiSCzVA2
RDWTF22FyWDYzWHwlWwKvg4ys0WLQfD19bkUuiXu+pz93YYCyrq4r3s9kaB7HOev
hNjyUCrkzrg6MZkOVquOodJGiFyCvLrsvysd48s64GnPIAtlTiEINQAws9jLjY4n
OfowqpGTeqMjqWvh5cBYlqGXALhgtK1tKLPmG1bWYIRUosVAn6Ao/U0M39edelA8
ZHx/I6oA+m6IXVE0H5/MVwzkGsmUuAUIANZC+aNk8wDPtOFlLeWyom0lLLvYmSRt
xrHFylOufVgEdRqDi0+v8kCFU4vCYAxmXJMq5WfbqIYRwS0ZTaK6Zc1bG4NIzUIf
rRsRQ61G1GbTOcje3pd60fYUjDsmNHXcvKcEhQQINWzjwrfUn3w7Vx+o40B1nFdb
GVaZXWYaRaeiEGmIG2xnvVFMil66rD6jK7C/jKOhBLKEyi6wotK2tE03zZIunnsE
1Qeb5Hbh2O/+AeErMX16U7JlFaCmB6tgthd+APE/xjqoc2WTPxd3+6d/gq/Spqm1
6uq0knjvFee5STzcnZFevUGtQCIStgCT9ZB/PAK04qEjaDF3GQU4zfzjN7x+MavA
/U+pHIHcp7vf4reqJEpM3ksjIotsshXUTEXPiGCv8WUDB9eIcKghYrK53S1LI50D
1B6aBNZ7DmmskUYvsxUcVPej43P1iDCpoPNFYrywBXNaWHF4E7zUwvA9IgamDTfd
0tC8QN1IwDZCEWZtmQccb1ENS2I6Gb2trwEar4QkSE1Jg/P6bJ9xaQgX6klbY8wi
gXj7BXBh0icMAFr2F+Pcj1BEhEBAhU2y61tLAPESfj7/addCok5SgMrU2vt00wIj
2BhRz140OCDC+A+aD6aJuEHDSup/ecSOrnNOkCLBBdpnXMQwywkzaRwnkawuXp9Q
Qk1ocu+Jb1ESLRjTY8SkG9/kG/4adm5r+MG+yOyvfLvCbXeLxbkz69Dz/l+AxjR6
gQG0cbHq7lDL7rkovizwqvgWWWJKrOkW+uYtTzryZAsF6nzsD/+/k2okIGtm8OCX
QTW1NyZKKcA5al39kSdMlFjNjxXq1HADBhKoejeBwA/nKmBF8EmVVubl89VnnTNF
AE1+Bjv9kRHT14otnei1URFoClcYEFcxpwFYBWr5JhhaXgIcmL47EQNqE6YV68TT
f2cWfuA5hKhzgTTUOmWOWMezwtmBeYd4foyPoMzX5sG2uRkKumREC8YEEf3/Ej4C
MgLimibVtzkBTo9ZnhqwkL3KS0G5QI71ksCZ48KnhTx1iUedM4Z/Lc3U8pNE+nAM
kCHAXHGkicgHeov3XC/Aa9V9tB+QaU/S4QKgX1xaBYtdsLcnHfQpfM3Ck1oZp57S
+Kdk29hsXawxAyMVmEtPAgnfcWYMyAsCXw9PwXCgpkYieY0wdAbjs825wN/Bq2Sq
Qy+R2LR292jf7B3qXzvYV8dBSGXjhCoGEfcffWzYhrv/m/zQJ19kMDic+hiG4tHi
k3SWokzwgZOP0ycgcvFh7At7C41krqDJX0oEymb7vvNoYY05skOBBTazLYKSuiVt
A5+GvQdH85kfojLusCkFm/9CIbOIVaD776POWnoJXy5GjFsEHswT4dkCLHqjph1t
fSMv1bXGv/Xa3pJvbWdTlwPCSRBW/aUunonMp8umWf00bntlcDlJ7HfSHEWDsJJr
eR3F+cTJ47DkzfRFlm62FsT3tjrudNRgmzx3LwePWSYSpBuR2btYnhLOZcoylwiv
H3DyygcT1ssRjDQlZput+d23sx+1I1bgT48oJvtJqOHeI7kw5OKAZT0ObCpHGO9+
46SruOg299Iwy635IsqxYaXj0PjXKlrnKA4jJNxJuUtK6/TlfAO8SF5eiFIi4NqW
FzO2vOnYe4TfB0TI+ZVsdBItubGbVcmC0fEtlXWyLvasZqMF/YNtT1EQDrvSExRL
3gMBOsHz3K8tWkKR0WVzv1mwCX16VFzS3YktWb755X/YldVsvzUxyM8k4OqHmJRi
cl5aLWe2Lz0TfVbSeKGW5CrmMBwe75y7x1nncdjROPD4WAItuucG0CjYuccg3aG8
7Bg+g1PpUql5yQqTSqhFWtiVx/GCny+uE1B2HNDmULLOm+g1Ffq3RdtG4e310BII
isX2xCtUeUD0h0ywjCVeI4f1UwsIcW5Rz/Mxkx2dtHyFQKSGFw/Qd3Mcg3pAME8Y
SpwIJoiCxr+FfVZGmZg9HQKg1/J2SB6BTNsHFXVRvSYVVBLqLgJBuoRloXFgE9tw
7AaVyYWEigtwhVq3zBV929iR0loo91k7awQv8hIMhUWlu9/MKy3Dqg1RYzYKoEKw
zq66rYiyC5ApWrqXGXUcXLNoZNiaHLwBflu6zjzSuhGHQQW/1fRBGCHbpVqCWzFV
YH3piCGcoM3XTPq7QoZEvUM/HxPq7z6Il405VjMO0xiPBYMWx6yKUj+Vf084zFXe
ilme2DVkS+bHKragOmzsCa6WpjJIOqV2DNjpoQNB7EXAwvtFAzwljnLveQT6yJWZ
vjgr7/1hId5fLs3yjr6p36ACP47tiKhP/haNNCSVhSGDFZcVZWQGq0DDb7LWrxab
Q98/VbU5mp8b7hmVrCpa3NoPRCI0yRpOwav7ljP+2dZa+npD0UbTKZYoANawaH56
7clzgmB1N0aV3p+Ul3VsxTYZmOdGyC6A+/g92pJKUYVplwEgwd/OELq/ZHc9GwJK
OdGRD5KUn7Wxju2ip2k8U05a5UDF2IrxkS5WEJTHmkFxLRBpF9UvREriuPAOf8yS
uPn1NP+YhtdacKyywAXngobttH7qKzwqNUjRBfUIZhBp1eVg5Iay3jffTnOv4x2q
yYvFiIRFEu413SCJMZBaHiZGsb1x1rr9MZtKIkIKlYE4lpRJfCq/lQNvmNjDPapI
gqGwWacmqo21nE+T75wFqGMFv9wt5durkSgZ6FZUkGf1XUOpUmena5198z62S399
OcA9FehPd9X12bUpq/K6xe9KMBtgIX+HjZGZwawJYViupLAEpWgm82WNBW6XV/W3
IDDkQ5plZPZSSB4jWvSt/QEvFirXzKqDrEkink0OB7Odb/f7yYtBy4qThRK3RcMQ
357zH5GtP0uUdxwINmELKykAe1RbS8iMHwtQk04wWXPfCGDm6NwR1lGu3CZ9ej6h
JAObZ2VlSaUGAqnycTx8CL1NAIFI4kJGK5EqbUZrFWQo+i70YknGbbXEqft9UZ/A
t8CXn/WSygf129RZyTYKLtstoWSlxhRYOL56vyv+TrCC2siEJmgVT3s3qHS+tbGI
C1PyG0DMFgN7corao0ggqhgmmf+gh941vHA2veOUYOGdOa6r5ier2ZNQzbIrZt8Z
YtqTpf1O/pvs0UeXRRips+AyOgC20BSEiEXxpC/TeLe6I+JBk1pqHyzdAdY7ZVvK
htn+WSZlADBaf/ARrKujqGxElg5trWNV9NYQNF7aIKaQ72Szupkde41+V5xcq0jW
tfcu8LtGYzNswtjV7Ui4hkvVZNt/vyZ8vRl88Ud0r01GIcYz7h+uRYDi0Gb8q1SC
ZKCufzaFwr6nhQTgZ9GEPEhGGG468s6AEPh/3rH5O/8WyvO68DXeA+BN1wigvkF2
9zC9nYKMoteSlMUU3gllmA3euCRmrLLEzUQFhkYvqAZkCjnledHEh515FVpdukRL
bFDr1PyQmawiymaA07jTbRp+TEEdorkcV+lXBzrshE5Y4pfCnOgXCub3uBBCLGOL
5V2wwv93EEwuiIkRKOx3Y9PDCGsmh/PoP1iOc/QFlydcosY1rAjP5TBqD1WHKmNG
M/oLI6A+k8Z3q+/8HSA7NNjS+t8WIgA8vEK8FUlJcdApy0lDU1e/DoKkhzA4Qpz2
UluttmVmBPNCv3XWGSGLqM5EuMiHoFfS3f0vgLirp44MBtPPE80Kq3VKgS2WCzIq
4XZyZmZ01lk6TmffFrJyrnQyZJJy9sFdaxvQHLZq9NusWc37Tgq/XUIoWSAweopq
XFglaTReWREDl8yyQqkTvF94djQD+kR/ANEkuT4T2sGD2UZNndOUxTsk+FJvVRn7
PTU9kapiWiIOncK92WUUPdXU70tvHYF96+fRDyiJb9gtsmZ9TLIpDR6qoq1yvBB0
5JZPMRdQiO/V/FaC5YC8CmLE4j24KWr5KNf9DnaUCPp59v2oTmVLM/PKVK1f8O7l
2/NaGtbEL8O+jcxD+h/p+T3EBJ8SkNkLeGbwBy/AYx2FNpv7pnInz01U7A4TWGN+
Ev6bGwLSFlu7zOK/JBWnpESq2CYeCNqrOAFZiOv0l/8a4atGUsIh7Nj9DcCF4yrK
ZpkYJVHIzVPpzgnZk6kFsPU3Tqku9DkJFLIc1OfxKOVjKeFx61LoTL8Rnm+MGAMG
Q24Yu8Xgph0WnhklKwPgwh16eD0gWpJmbXDoZgVuH1e6s2MZcx2iXO+pj0pytV/v
0HKXFIChQwJnRcObWpyWGp8HsMkUHCvr2KlcBF3zZmEshDeFIwbcr8u423P0Mm85
E4CSp47DV+HPsdt1WpsaDDWzP/xoD1kfeQauK04xwolWRLUykxiqayIrjqPp6Xie
G1AYpgXwTgrgkJ7jIh6NkMVgFQYbIj9KlQAK3N4YRANhYzFfg1EYanxYahf99xPC
9RSFkzKGF2qQIBMZZ08D952dShipJNOBwM4lnBg9GHvlafT6Ql/sLvV5s6aApIGV
Lejrc09Euuz49b9FOuF6oBKxql80F7DOuzlH0qHB2s+oqJrNF/5CQF7TQnlo8lMV
z0zKbhoY3gFuCWE7pDwu5D5ba/ZV0Ic/yM7VOElBWbu+C3I2UmtLpgj9ah+Ipvgp
dlu+fIJvhD9uoLwEypUeIWCPZf7HQ4oAyqpr5sYCV3U1Y+mZQg9QSRtgp2qbKdHp
Dwgd5h30GAbQAwxyXtupX+xTh9iCk41M6lS53WtpbcXWOAgqSsPdzvc3MIe3f8/G
VVSUpB0PbnYKxxM7zHLFrJYFBRCg2PEeAOUoZuymtbtJtHWBX/ho5OOxDb4HTt7I
xbe3h9gCNU5VXkxzBm4o/4G1D9SEIMpwgTF68d7FhQbgAtgVguMztRjnsEg0yIts
YCLCe7X6+IBrjbKHj7Rl4IVWJe/PsENcOrcYbSH5NgSKLM4fhDzEnOrq1Pf5bh04
LMSvpM5YeKte8SgJhBpnSO2IUU5b+ozsDLn0ugJcfRAdm1b4Pz33E9ZGxB2XiT+3
TMZsQA7p/WqmEtS3FpI70Rv7/r+95SmhRQK/DdXp3EyFTzG+9n2i+zclZn+259/f
aD0FClVx6m5IOreIAeZKmHmQmtQ1oeZegulL9YzqBVAozsnGrNJAyctbFTyEps/h
Uu5xeOrFf8+v9L4zXeCy/91NmIJaVVol22b6tOMg224ViVE/gZq36yPftrrj4Tad
OVB0Fj0yQtNJhTkIttNUZsMGdmGtaf/4PkKYad+rBbskUbF05u2vP34evNVlaFiO
4Zb4M2aVDKXllP/aujOlE+GcOJ8SVL8ZiKnvEg9/Zq+A/QBLgLiUsg0bWtdQEndx
NkNq4etTiFmRN/d7S1SPoFmzPpuHNn4kYrgQ0iDZdOcOLNVhqKbQOFqn1lvv+Xh0
aPgrGsRCZfwukE73CPFISAGoQDXhLLyRDDQlVnnDAIX5Svm2MxNm6Zx8ycMTIpIi
g/xB0xvkZghRtlp4nMKujWaJmebw+9sb2ppfhP7XcNiZgtpmYvb7YcgW6gQbpZQn
wOYnuYy+ZZiP0+OIqbvHiPQrN88yQnvrDm2BdhukMqFsxAH0lMr5UDwym33LQhXJ
pz5sIF5Q28vWptD4EXoZsAr+3Uf+5FJSYS0htljjedMeft0546RArC9rbNYycAh3
oW15zrxNE1tWE0eWvE9FPlwLCdMPfqL18GgnvAwdNlB1QjCrfvEmUJlgFIjZzk2c
IhTBKTqVymFJYWOkOCXcmm2xFqT81+oqqLd1GKb+nMxhkgX+1ExvWvX3BWPWweoU
M/txoey2RmAUMTuXgxSwB7rHdDdH30vs2af5E5WsIS6RbRM5il1R2NKAjAKaWR33
g7CAJM/zi8z+SMiIFw5blTLqjgyceXcBQ7dkM1xhLeKybCT5DoutHh1pumVdlAKH
ux/rrdaryB/9WemyzZjoJZZoA/ULj7P5VznZ54NHegLiJWdK85E1YNBCYm7S3sOz
phLK3r7XsA6jWTFcbjhapCikCoeZPmvgvhk2VoP+Kh/nWY08EYi2EVn70pNm4BZ1
KiHzKmuKCvya0bXefLsclmwTA5ZJQyrSh6KjcTcI5aoaKfuquXf4B5R78a+K5FdT
9Kyan4gzgLOvHLUE/x1dck1aEM3XrrHnPsAgaY9XsaVvkQnifFkMGJVimSmk7FG8
JkVBN0XcxvhQfUPmZErAPXa6Wg47PRsHpYe9EbsGIYwIooHDguZJbQSK0SQ0KcmK
QJTEyfIkexaYBWt1k57FshlV7l6n6i2bng3figF5XXBG0McHvid5iqe2ENawfFMK
Yl9qSDQlPpwxNRsm6EIqhrmkSaDgLCrLhYLB1VBX6XIOOX6Qz93RFfrVUEHPm0Rs
lkBSVFyYkFy1FLMOt7sIfQ9JElaFeo4BoSrE5iexnIAwm+SQEvIhI4hI+KA2ltz7
Oah5Km1q0vyBSJgvbkrVgCyTN9l3/ZeC+ZPIobrwnKKAR9Zo35YUNMKFOPBy55z5
yzVAXfYme/4VsKumLtmzhk6RlqiVH9OykVH8F+vWyeROpZn7YXeBp4qkYwry05m9
2PUiZrxt0gyKCy8nlV8DmsiIEq5/5WhecD9EpVtNmZ06xuUKIlnaYTc6l2CQ2uWs
2MicLyNRaVyOmMakXk45EIRz1czuXLCwemg1VHF4cGMY3f6P+1yC8fgtZB8Aat7o
nXg9vRSDKme6xvYJPii3BYtx5j9qR/QUz2BJPUFYhu8Q3EtxIX3aQXIsvs8a41uM
iqgTWKmDQxPPumgwmAS70B8CTtT4BtBmwk5FRJM1UgVwhqgkMI+W+XeFa9X4Ev9k
8NTxntkCx0pN9Gk9ZukAJ16Gj/DMvEim19hFS5ro71DYlAKfpy10ez3jDdtZ9+V5
3LIs/f61zAFrM1nLj3mzD844l9f9gncmEg4rTPED1OFSgU/xVGIZP6RHU6m4lDJx
xenut7+6HGvBKrFoERoJD1aUZqMQFl7xz6Q5iQKmsROa3R/G+vl8xrHtdCDRfJ4e
ZcTkR70LQ0ZSJ/WeCseqqDinNci+Dc6Hl7j8EYJlenqqd8dkujO8xPsymyhst2gf
WjIGwuWbpRH/62eqVXZTKoPJDfF3+eQobm4l8x8YaQcZTYEcH/4kJA3B6spfGif9
NEYS/pN5T+Ep0g0YJAd0R2mJScl7+rAOtLEJgT0mLQ134HjsHaLbi4AzzS5qIFkK
JeSvdpJ71Mb/UyYppEkrd9WtHz7krmZYjQ6fa6lNPpfBicHZdt6wGDGb5sb+2u/4
j6ve98iPp/acKL76CaPmCWwcwJNBODenNOQLDv122Wu6PeLYXOFBksm4E6cABvqe
0TCLo/R4F/MTdTFpfGy1eGyKPXfgDJygwWWTOhB3Mqq013MOz6Q9IOlPzBO8Ka0+
L5y6CQ9Ktk2xMJ9nmxF0mZPIgwYjipyq0fBZdPczunfyRPMcrPMOcALqYNTkA6/d
dR2O3BW88mzWOKm+zVcDLaJOQAuHQC1Jg1PITojPOAFXzvcCSyrnxdefF6KBWb0P
vEW74FRh3hPcqBOUP0lMrNupC4EqBQtxAE9mugB09NhlyFBmp6TtFaBZwCm8L6Mk
/402syWix64GacBgSpHH93EeqKpCa8lTUAX9BktHPWa5Ej68chowDQFsO8HyyYkx
8wAOqZp8cnX/Zn9Ml9hpaFSjjLfpXGY2GxgmjXXzwqijaFb1A6Fux3c6Uq4xXEsE
9Mj27RInX2LB+tJqP6NlMGzX9GLpYxVuk9ydBdarpu5IRtNWqm+04CM4MKEHKSdD
JWz+Cfhf89x7yHuKS1+QjUbS/Ug6WPAv9VcDCuzxlILqqA0PtjNKLP48T4TkcSCs
HPgmBrqnFukB/O3ymzduURSuwbjQejJcocCM9eaiDkU/0ljUjLfr7KrZqr0VlQvK
hIRCDnJU6bJkkq3pdRbHh5c3xlA/rKclq3WhEhy2e+8s4TRRTIrW/08d+JqcYGLr
JiVAJufxTQQikO6HH5GmufGP2Uff66U96E+FnIVm79gjTGXez1+awi1meK/hpUEZ
brirsi643B5rYMYgAyyBi6NL6koqPQCvf8rCmHi4vi7jfyezu4NX+lHCa/dM1yuq
tfGP/TZs8lPM+ZvrWOL6TZZ44v8R0UcCsGn6z7TokOpdfpRvroz3rGuUmJBSy217
aTJDrHuKLu3huxifLG27RGgYvcsSKFSKDRuvMbnGlF47eBij6VLxVcwUsBoULPYm
HNfswgHX2vMq5OYVM+oCiIlOgofvqkSd+EQmoPVPNHXCSxZ4Urk/n1vPfKG3dICF
Aho+PilTWgW8oYnDlhULdIiDgCNBT3edyO/Ezg4DtlxUSwTj8KiJrmll1G1yhlTS
flZb+qgo/RjCe/bxsnhVl1Dx9tsfHdAQyUyXqgz1wfC+aQxPsZkEVfOiHI/xv2CH
8+FvYQkOfQXcGXlXR9l4EpecllHF6EB+3bqhUoMLwhVDIpHA5MuproEf2XN1UDNo
+n5EMOif3KvgwkOAqFI+eB1HlTJMZlazgt9s4xEgjgLKtAM2Ckuv+1rnDbdIqumv
gqoxuoduzT/buimy2t+LKeUeSkNoj0e0FfFK93j5DKS/PqK4sdrBYclPaJhDgDcq
kQJO9gstkkHoJ/rb9WvuFlrWfTGaNPRY033iQkAZj9EiSpWsCZHF4Nx/AHgwXSWA
9ro7K55c3WeXaHsXyM+QUYMexTGrOy7anF8jFObRJR644oWe4D7g1qSgg6pqhDlg
IjwMyjgSDl4A9FC5TUn4PLM1t3IFZoa+NyRPwJh44qq0BvyBu5PrKrK3fWAfancd
Es5vmXoyCRSql0ZK7gX+hTuvv32e/jyZrqIXCV5Rp+oIkJowZrI1kcGo13qXwqdG
nQJVzPSaOosU0o4OeqofMccjQvSUvYSUvv5NTtod2BiwTQrzpcAlUs0mCQHPgF8J
62nvGqyJYn04ZYrL3E+OEfAh5kPM58hoxbCAdSCFtFauQ8hu1k+A4dr2W58ZQiOF
mxfJFpSOd2foJI6cOOcDDbWvc6ICH/gUUp1QcmluQT+r+OWaSjD0wQE3qgomzIiz
8bCZQ7SuPw+WXmytZzbl5EXh7637UmZOorQVPyaApuBIGkpqkERk+3dq3TYe2KUX
EB0irbDuich4Fxgiyhj9GrTrg0WgwbK+6TOmozLWkQsiS1WfOVLkwAu50pqpNN3L
DQTnbM/ubVAH1enpHEn2rjLEQF+QJlY4zWFnKDK8dMDAmT6cS8exijO5XkBXyCoq
oJ/P1VdxwG67ngQ8qWxA5XrgX+RR2DDFBKlP6vdJ4yqDhkZKdARRCHCcHY+0gQc+
ZMS3kAvmD7FDt9AB4rS77raHIwQVErODTpgkqE2CjIX/2TnHvpnKHKFBPUcGH7+B
Ue6nfdo8U99KETeKskcavX6noksecRdSG0MWMS/Y1ydNynz6lr/0iGWYJLJTZPzS
9eQLD9CGEsp6JIkoXhHe4RKR4RT33aEGhq/iNihjSK2PPF+Dg0uqvhf8cVL4WDi4
Zm5g+1qPwV7yMGLyEYy+TQVPRumQadIKfnemr91DnQnzyU9tM6jensyvx7zU8GYg
uq8ZMEr2YpS4Y0WJ+DL14I0RWuhgBujts3ugmoHkHpKu20z0U8z+C4hR+eepbc3V
tu+Qw1Uz+ZVcsGli8/Uj/FO97bGVA6nSMW8OKFOWIxLUNdKwrXDYxN1w48m+7X2Z
a+SXODz49ecktr3LmbY2Ty604ukgqKUez3mkkydsPEQTu42yCwEJ1vHa/qfMNgM7
fAH/kqza3F1Hsb7XEq/gqWDlo7Efnn6pktftHH9rtDIoZFoXQwJq4IhNHS5KrHAg
maYwaTqf7prI1I7jawcIkPTelMpilbZJbOmMe0VAQK2m3xjpk6NNAlJhwKKuvSKB
37ce8ywg+QI4/z8abxZ/md3g99TAOWmAXLOmlEhPmMMc8t3OFPjtje8J8QLdV19V
7J6/UI+ap/vRsRXHz7MZmvLvH26KWLmUaUfusBko9WffJVs6jw2kSWzELS0mqvek
RMXmVymkn+MjYJfCOYTJzUYH8hP33y39xRl0L1CpM/JnQnkv9W3q4QiXmI9NrMYN
uCvFQ1M/LheZOa8gZkgLnXsNGHOv0tMU7jbRlHZK8yhH7cQvlb8p4pGBlAYe8yXY
Bs8G5Z+4JCkcZWYpwT6ks1ZspCSF0c8/hWBrEbvmqhON8Bbpgnm27pw3lZxLbq2z
gLKZjmi4cBDMrxWppEKFRyUNRXNpOvzRcLZREemPx2cqnDwzE7Akjvu+ROoplItB
PxQ/jydNM2buyAq6+UlxkdxvFCc+eg2s5t8J9DtJ8WZ+/kPBFfmmu2cSSKY8nGPv
UPMaERTwEzCTnm8zxA5PJUZ5iCTVcp1WczNgD1qUDU5rj1RFeE+eT1ZOpXp6N5ZG
ZNUNNlal0nF+Nyg/0MGx7UZ5i0tFpb8YSAMClO91xofyyti88RGMLKqEmhOnyrU8
/PVppxRkQduHgT1Z+JAoLc00HrSlSR7lX4FmqM65oS51ADqJxgEQnd2C9LYdlIGK
e7Ra0fL4m/dUM4SUOB7SWJX9nH6J8CFhiWN+mY20pxvbnX9uWtWKJZsKCYdQlIQw
KCUpkV7TIBFSVuioqzJElkNQti2EVUzmDGdnl0vubLux5XLq2pzuR5rrCYC10u8Y
oZRTlI8bEHKTtwM8cZN2tEHpALad11Sy8JAXQlWmYXOmb6RVLOhUcmRXwtgfJf1V
PtSzy8iGGW+SMyF6GhelU/gHRSS4AMK+Uobi7GOqZY0D7ch32zP82on7ezKCdCdT
ruHObt+oAC+G3QuRml99wLWEs3uB3ywSPMoUhM9poA8bNTPN2fE5XAIEF0sG67TL
RgMY/+TcohQB8ai/Vorwpsf970i8d5psPI98yq63v866EV/NUjwQ7f8uicSrYOst
OiQMRJXe+xJaLK98ZK22YKL8Mjz0PXnDf/3KRciuaSAb1gc8oIxau+U+npVbFJHX
PEGbMRN+TH2w/bZ9uajaIo4qKKcMXaeEfexFOrqH3BzWxvtSDTTc5AySjH0o0rd8
23OHvcy4lLna+iCD88+cHa6i/ocjLwSNrgUIEdtF4POCOHOX6AWIbFxkokd4Ub/p
BLw1PqQtRd2m4EBNTW2DCQKczZ/eR+HbtzaLwfHmEiE4NG4xVTiq4lka1/LeifiE
p02OQKwVZexC1v7PGAJBTRkJQl1tLhJ9vYxVN+BVYAQpeXVEYBOUrXfKRo7soFNf
pVB6dISseYnp6WigCGvRPsZogSWupeTDdd53tnZbOSKkcOGxj330bXUlD7O2q2vt
WwZcsKdDah2Z6hd3PX/vMtx81yne22U0wKDv8KFj8UbR/rgm4FYLjxLMAElickH3
OeHEOd//pVrQjfbdqbougEmNYp+opOo3IAaiy//kkIiV5unOdvtAbqRalUDfPy9U
lzUBlgnSSkkTlySI5fu/AZmp62MqCTI26V28G+Mt/7fnHdlRKyTwPDTGyii3z3D5
1XY2PDyK6z8SsFBHIgZ5OEbq35xdGAkc4cSusiss8bn7Ux3mK4vRS5JSosESi5Ys
vPg6pluTQenOrMMGfnkwY2/Y7syLdyhfR0qAV4SngENtUzgugIis79iwF/mhdNkQ
gyDGbmaZbTe0fVAV7U+SgLWYtbXEbuFRpFBfsD8I9Zm6CkyDqZCfnL33FLnuAU7g
tYUD+RBlnqoHQQ9C9Edkv1WsGYdvPlBdTy4D4S6WG7/dQHt9mKjBaWREWxtKr3W7
P5y5Nzm2vEQrd9dsHbrDXpJL8TMsRZCcLzOUgpRfSwcQqsvSCJERUb/CnRGlkAdl
LOlv52M2usoVPj29jMgu7zQ+0L+M2blTfRYHeOZAHWA0AAVGuwAdyd+Bsxf7WGGF
6NAg0TtopSNLdSVlyXjuBwLMxdKNJQo96H4EWSKf3THAvYdv/8ZRaDgzupeyuCQN
+p8SQntDnRfsi1nWc/RfSZCG+4jb73lee7gvmdUn6ToD9tb9JunGuckkAVxDaN7x
WJwcn4f5iQ1nOL11We0wSHXDSjY5KL7CuWca/bp8XQ8TzjbDAiZ62YszjKGcxqxn
YF3ITcnCXsFqDqL44nrzQkoJV9qDsyDbnMZ2eMDHOCVsuOQZedY24hqfE/FnoB3r
Z7VdpK6P39Aa7PuM4hSKRnpiO5V6daTe55Qq65LZXPywxS+FLtdZ2RydPoLJ7jzN
2s29/4rdbdbiUwPxZqdPyAULWvAZ9eDsKiN5Okhk9ywRz1+sN0uUk7xbMi0yH/1T
D5fB/B09mOaApUqqN5UQhcO+nTB4Du4hyBldcVv6SHyQX5CawiPrSsaBn3JlPFBQ
6LKxKeKWOTjI29zSJK2Zy+XUfgdtUIWh5AdiJougUpmL8Qc6Zvs6fH5VQTnloMqW
nVdvWMXh1mgqvqOdviQ2IJ1gtjgwZLxuVaby6hcK2B2XCRpq6yYhMRhpL823i6b4
i3xk7SEOFnRuo8IIwwHqQS+YQyuARF6faEXx7uy4Nmtq/ccBitiSKMXdOyFVX8Cb
SGSMgFoFKNa7UJSfazKnYxLz5qyasO0s+hU7y9qoWdq9m/fDgi8fiTmA7ykmTU9r
4Hv47Wka/YC2ReEJu17PJdWiv5lJHqQGPPkKyZTMNuyOlZRkz/CPN+sunpBHDOE7
RjSRbIZgA3zpGwxKoYShOatb/D4IOXImst5Kb3JVmD7iYEFSrs4nMVJceG9q/unL
O8as0z1i3sH8kvUu9a1qF+N8gA5Y7/Y+fpmbIuIX5moOF7395Cf+0Y2NKrZh49hV
gELLp9BekPt6y43c4ZOwGbX4qdMrbbVd7VF0+pkYRi8MOopFQ1qo4w29315Ahfem
Sln2bBlpwok/0xpG+jIwVj1v3oNHjTBmiEX9tZgoCAjmZZNHCkHcwNnrqdVkd3WO
v0NA2fATDY673i+TaNrC0T7CZF6XJxrkMBJR1qxnZH7CcUcJfex07/UZRgX75MeY
XUkpkeac76DyFXIKL7AYzvLu3//Wxip7bge3I0oe62007K/7/KxZDhCXKMUd98WW
34j8XP7k1kREyISV/i0so/EMYsR2mBr5g35P05y3nd4oOQahcjIZbVXyGMutB4fZ
Y4G3nApm3Q481Rnnh9un3VCB8UMBqAP6Dq2exFEoatDMPJnMdQUPAgIQek2zubHc
CQYFVrYfa/3fYTHSqGMDyCiEJb3np7YDXbTdr50Wqz/2crqr0V0faOKwctY+1h6O
voimUsTgUSR84VSHi3n4HAv6m7Z1y2C8LynsnEsyC1oXJZCwF2lfzt7k+g/aW+zP
SDhbMfl309R9gjz82y/q7W9OO4m/lugddaIvPEcOoaMLVOxZGFfkZMpNdfs6prBu
QRs4uhqwVJUSdEABQnXIuF3NEOJXFUFMLWjM8QoF0OoeqA5oHJLZHpQCMVZzk+yX
dRb8x3RD2nwA0Dra+Df7xhXffGfonxDXySwOdK96LqmTvvMhZtuhRSBlY/HJe5Qz
akkPNQIyfuiZlt6j+l1MUD+VIvW5rBrgm8r8V1VevUP0c4zjvNk8FCVsL8fvL48b
MAHp2CjBMHvB8mJ3cQVO5Oeah/W+reDMO05NONNBQcdh7SItUx0oP0JzQRQgIsvb
OuJ7TVpSQNHC0wIm1rv97f7ZdtZnuxDioewvkvTwoqg14UN+Q55Fgl1tY/xfCUcR
oul+TnsC9UpEVvghm3Pi2V3h5Kl5810MV2+oLgaIFIzkB2t1FyVNZhSyO3d9oxPN
+85pGZSu5g9y0b3DMHraw0e0PGJKed9YMDQ9vNMY3KcYU4uInyg32UvgR5ZIQ+9R
2Fd+pjGLBuQs0UY6C/wEZthejjYntNBDFljLxsD6mnK2M8iJSPGQQl9lxn3oyK7e
0FwFafUyvja/bOy+b13ALLW2A/a71M3Ph7wg0aP9SCr+5Ril64xQHp3xJs3r6hFE
kp/+Heya6IIWbpMl2cyqyW0/F854/3N46hgZuyTDpB+LBgVn5vMMPqpAFgxXh/LK
cQFrk5vDCXf9CoSfQ5xPXT9GuAlanQnso1o0Ho46EWk5hIsACuHHBQVD2mFBFp0C
AUsBWvvxRds9KekewrCG9/1sltC0Oi4SY9hXz7679jVe1nwfVJ1Jb6lWhQxVEofr
QEmIUtU6V8rVmqQSV9dONZ8nQ6YqFngEu4A+f3uLkes5OCtAKz0/1r07NrN5Vz6P
dyUqOLoiYlNvDVnOhZoPcoyFG8YUqpvn741OXvP/Yuk225nZdTgGXOyn8YpyezB0
JJ/k0ly4eNBsaEtetbIwPyJyMST0NoYunaOp8fbQPtTcm8Z9pM+GbOpZ2U9zR1jr
z52BflJ0C64P1A8SyuAlQtLPF0TEneYRaoiT0zWf6ncgwc+j0K8eh2bDCNdeei/P
NbJA1QANc7Iy1Kt0ZSL+iaVRt6Lh4+INVpdaJFKkT6CXdVs7txW79wu5otOlFrIl
6ocoHLsi4GpHwvm3mJaHnKUqKvl0S5xOeYi6EwZXzKGD1yh3NxMadRGzj35T1/cv
T+KG0htFKnTHA0gzDiKFA5zzAEujsh5cxpH+PNbEj4HDkenIvMsTDHsTBVQ/MqT0
Wh0NzyXCrLTFWtHlwXldXV23iMOGv+ZXkd/yNgPeMtrd72N2OFI8YTGx5Ic8Npsx
GKwPlevZMRQzJ1sRF2uDuKn0UBviKRuudJ0jHmc4t3CIgYb0Q3gcN9btnS4FZ/4U
r/ObMoBRYVwKwR0Bw9ABkbW090FSnm192+EBVRio96ab0hRtLB/S/4uM+0SbtGsB
ArRVp7s0li7uwwkDK+k542o/GsSTRffUSjZ5VeDtO30pDx/sxLcnYLK5u1i0hc/V
A8FPSsNWm9fQupJUFbDpqZSGeBVGR5jCuBq6fkW4FhNP59hXfJMJnvZFkCmlqCEZ
fCGoriLes2R4TW3k+fVwQvKOjbBi6zboNFzZnN8PCqTi/ds0KIPkCb8OJns+8ajS
LUAqQQjlUsE1mvrS3T6Wf0VYFrlUOUtfTEPazjpff8dNueB586v4/bbB2dmip/1l
yDwat1cHTULl4ShLwB8wQ0D4xzXyEvb+RzwwtAX8JTkkspQp/wqC0jCoDBLI14ic
GAS0Ar2JWrJq0enpTvsbmVRMydyOY13/ALuxSMwpDsCMY0OE5o4tiMuaUAjt4ewd
i2E5SRmeF4mrd88PJ7j87l6+oWoEkrAchWxjIrfjTuw8fbQ7c6hXAuRnFkcDheYD
WpMevF+ubTSYChJPW0wmx/DHIil2sngdrSAyDBpW46yPbv3taOFhQ7gklhg+HL20
Y/ad2X9DMnEKZrcNvxJl7iUyBDqvgAn5OSlkce6wx4Nc5FEowOjXo+Yv4CWKlbus
V91ynoY77gEjlb07Q7DX9jnl4YGT3+blNqXA8zVzd+ag8mmGswekGhdh8Em1DLK1
5Mj66Xt9SfLlQItb8n1YwtfdvPgPzy26qGVVZJ8Kzlg3F6k2zvErk8B29GvhylQq
445QHWxnUfn/l4BluCK1QHn7nYNlhrca+Gizs+Me/fAPZ2XQ1vCHqiW3GmvazPLg
e7OOUkexC/88fL2pNFJNi7/GMjHAvWkSFNL7XgeaMM0acywqhNwmQUY5tZ4qczpi
flie1I2rTB0UuedMarIcBtEjUEqNgWs1MYqUXBGHKn8l4AWvA5y+TC+fR6Fu2biQ
B+t3DjvoIvjxdZPYEMSdMJwTYW3iv9uFM+m2XI+sDKOLbwyWrp3ZyPMF4+BKNwcN
c96r0uZ5XNXrpB82eiO27pfZ00FtdphDLXNyc5wSyUiM16Jl9p8BNa9GjsXns/HV
4bP/izIG5aUmhppLfWgzZqKyITMturHmiPYph6Av0Fs++Xs/Maol1sulclDQkgFR
nhoIHp4re17/tB4WzfpQ7AV4Dl57kMS5LZwF1IbY0Lw4a4RuAIKM7atU1zS3U6fo
GHrVb+0/qtolwlQnuhqBY0PQCDNqe+4JdDJ1dTGzdilIcRWvMcQ7miNnRVM/3vKG
9oYVO/1M0lJhVnGSclpIj+ztilyeqYbo68ih90pHaFujIhT/xlh2TBMa7tJsDto/
8za9u3kA4uINz4eiRExvqEX+3Xw4AhPahVC43wx1VQmRvsusftvOIWPp7bNE/gXk
cRtMUlo6EEuOhrw/Obopoa7nGnMzRJQQkqdxd6ZTWEKCklf3Ql9gAdPZQZdPk4V6
y8MsTHb57qa5KEk/cw3r66QSMcng7tkq4AG78aNqRGHcfTGTgcMueOuQtxx1vCof
N7cR5B7FyYdR1A8B+VeXybkwX8+Z6OIAk4iXbExjP+yGbXbrMiQYIxBZ+v05ZwF5
JpXUzchy2wZwM/Ti33NtEyPhtEoce7mWmNgY77hX6QjG3cqQeecWrTDH9eyvsZA1
egnjShGKxKUzo3K+I4J0dfgjIHQV+G2b0z08r6cZNcVtFLexfVpN0z2gcSbcR1hn
3zyXFXWD5bOAg57ophIoFBtBxROgvevWeO+vJjRjfH5DeDDwePRusLiATWMyZ181
pW+hpPr16RW/l/8s7mBLt5W62yfWCtDAkAZMSE1pX59sOC884QAViqgUXOrw5ub4
fBhX1rQ/wLxiKiCv7ypzLamy8vS/qPXu5bN8yucPFd0esjkvlkRauUgKMhkb2puF
h99L6pZlVOifl0d8FpaoxceKG2DdRMrod6BGBuBn9RkJlZvPm9fG5tCntQCcZEVo
u1AHATseGD4qQjeRIPDNlOBVHcg+HNGgRFV/ESspx7mNivrxfy0siyPfJPyHdU7G
lDIllsFM9SjHTsT8orzHtwXDgvmEas8jeyKL7QV5PMy69HVoK7kAoCDYL5FbdLoN
jSCmuBhM2Fn5T03N2VHhr8r5UbcVzTkxlVCuDZBc/0epVqcF+OuCkVQ9J4crhgJu
oJe2J7UkxGZRK9sLrwoI7tdq1HfurrYW9wswiM0is0gUqGjoWo1ynaRTh+/Zq6L8
QuNZeTaNy80qdTMT1T5rIPt71SKMyuqR0Tjh4z5bIyZmfB4ay7I4BhAuJQQ0nBz/
KtElFnS4W+T1XA/okiQwlwloZKvvG2UMChDxNHCYCAVOG9f3Zx7YOweVjStNKqMl
Z2LHXTX3JCdeH+S6f/v2G2mM35ZDposxY++IS0Dq/Ej6QTR9S3M9l8XuL+a+eCHW
Nvz1h2HRQ+mVeFhneM5AEVMFUTZKA0aY4kFY+s2/MsG7wqZSKHDBnerZSApgd+gc
/d0Ff/SH4FSj7TKAAKvBxBJS6wPa+luWZlk45l8dw+bKcdEMhRMEn0ldLR1vVl1j
mP3iUqVqDX9vumrotcvE45ysRZ7kzqiNnBWabiTL1aaGDlTscJsbWS9f7ONquzov
gC4IxpiEWbSXGLhvn/1kWNdwR06De7KnYp6fq5shqezWIubUfbA7dzfdwi+q0vwL
TraN6VUHELajZHdQbmnKs6PuGos7c7U8Iol+E16p21HRhQRo4AWfgylHU7EAlOte
aFXiRgBhCU4hpy5tXIN9mnKlBUe28k+c2ZAr8GzmGq7Bhk1ywnxo7SnbvEqj5HOn
pH4l5veRaVAdq1SWSCZX5+KYEZpufOKLK+y7sESRF7eitrxx+Q2nsyBxBAK2GHJg
CgLOvhGJBkqNe2OiHKqBEBziWtCQC0dgsSD9OT/8NKv3onGFlzboVNHyOux4x5Sh
/9lSTzqpWuF01FoNJLFZ8IuRqJ0voVz7kj/ixVm/y2z2dqmBjnlE8X4390+3dq0Z
AOOtMR0PQU2T7PaN0BJrfT1NdvBhit4VTwJUgQpdI9Fv+hk27O/RpBuj4tZrN9h2
tMZAqR1Qh3+sc3BOFAEpfAEyMdL6MoY1mgAXMUWyH7463MAGJu/zQP8H7I3rfzak
uapflwhls6tv53NIqKbiweFm3+8yXObXQCZJedP/RjVkeHBRAVxka2tJbSJ5MKBc
lszeLpqWFNhgFklj3b9f/JSt80olmwI84tB6OSuIKZHFeEF0CMYUgCnOpUIeox25
vEwY/Ut0B/z+m3aYwfGzUezk2IgA0YLZGxEAoTYxZOaKC2yDtAakkOPpoqSWD9UF
hCgkeEwMfPU+/yr1ImwVKnaSCvIzGd50H1qpsq7YYhRNldDj7oTcDFVPDETU4mhc
Ado1pENoh1N7O+H0jPFRg9/oUr/8SOdUy9ImFt7xvlGZ/nWdL/0xSzq2t1Nqvvtq
KG2AwxkovjzG9wEOIwrxtJQuZ5eNJz826lU2kEOnKiPo3bRddYdrXRwU8zU23g63
t8a3CfvwMxIhb5ILky05V2v9BlJzz94qQtL8Sgi//m3WyZt/fLZMWPhlQOljsVMA
APaxE4Sj58h5CSZlqHImIVNBDESh8P1xSDjgWKfJVysOrTVt858SbeYFFW3XoLhO
WVy7AGRWG/haxbiNpXrgLxCPKMTvo0TNXGKtAXJPDuu8sESdO87hIO1yDyvcYGz9
/kAvFe7awC56r+kDtZUBApqB8JC5w7nEKjU9ifCYAGXZzKcy3O/gDugr+Y3iCeF4
4llMHMSYG2VBs9QbEZ/gS/uZZpIB3Vbu/RVor6YYDkAW3P8UqBu7h0aBZQGDG6vr
5zAJPKMsyqtLcfqkUXBE2IfF5i00Jvw4Qovr9zg2im9bu13Ti5gKvHjlPwVDiMut
6BQ2Q0BNLmo9j8Mh5HvTnAqxZoM48J9eV1M/oYZZAGm2Bz2aXODra5su8UREJc3B
StegOAka3zEymkhnlQ7ZmcoZaxENvDK3AB61F8vH+luciR3HUykFx4LYAI/HoBFS
ZIIoo/+anwaEJPQbsUYMjR2kBNcxxGoiIRWp/sLc2KwzBUtR34HGeY6K2YA9yh/M
EOP4eXDqfPMQFW60o/CUOiGaP8WSLbMg5q51TvQqr0rHoyu5W07g2BNKWKul1na/
kOujQTpJoFYvP0CKkPuYEuL0zywQFpNJ33Z6rmqB5ncHTkBSSBEJKaNaNq66cc1z
RCixKrM+ZgmHIVM1QXu8+xLq0wND+TZqstTZ+aoEOJMAjC0BF4eAir/Tk8OUDx//
otKeTsle++hsal+ei78k3Unpj5CjWioT9meRWaqx6JJtWDpi+jpblVgQmlWOrwt7
n3u1Epvj3rotGT0GJZgORjypcPJIg+sgiFre29M2y7Bs7KDQwmLegyAxkgZbKtaz
AGptL8/kSIFgyEp+CmqtH4cedmeBxuDhg2d3xuDOzvzGG7VGLpLkG+dfjsifFIGm
ldhFLbfDsMiA/6xj9Y+pnZwQkyTBsstsRV2wI5RveSbBDIGP+Qi5+281r44TS0AG
o5uUuXyvY31tV7q7/dGbkXdLH+aiEID35kG1tnkgCK+0KeZozr6dpT4dhlcKmcQS
Z2Ev6lBL0fHnhbYmu2jD/LJsbYcO6S/VD9Yz8O/zDv8BCKOVrTf80UrbqOB9hgjE
Bv+sZV6iagB584Byv0O1nW4pnJo2r4RytDLTNVsnhAkmUno8jer+Smy9eZ6LfpgZ
pZzI09YRQKBow9W4CbJpktnc3TbvZiKV/6llJ6aRJ7kjRIeniAF2+9UQNek9pIg7
rqSJSZoYMpnyHkZyY00eopJkjIjx+39nkdFvPogZdbr/xbTIl/znV43xXJShjk8+
j58t/P4CQq7+4K9IOdfntbeXYqr2AM66yTa30LF7yHa4yzMBIszlR0pzkbcidRdF
IdXZWpegvupaYTTg6LWw+A==
`protect END_PROTECTED
