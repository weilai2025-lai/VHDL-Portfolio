`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4boMG76MR8BMPDgqIummGogDGVEeezg6gCG1IbWVOVKNL7w2m5ARGcv06sxAsK4M
v28nXbKJx432Hg0YfhVU5okeBVsqURpHll8N3AhnbZQBkzaf+WVz+vCFZSZGtHQj
4wo2NKZjhS/2qqFl1VdQUaxsfI9a4p9FaS0Iecs+cPIBOUTE5gd2RMF1kIIl5Nd/
8ZH25BOBl9CeLnYdyOUWBGA8P12F2pw6gP8wbNpYyTjUmbkOoxKb37u1IJpBEBet
5+jK9ug1tiEFkPtCrpaH99ZU3b6+hq/guR+4XdwnVHDJiTMqyrma1AauAEMCeIqr
QFv8t56PuaGfyCI5fsPIZNJUOIUaPbn5S8K759SXCLpgnjfZIbGcc0MJTy3p37wo
fTvxpCQJ18OoCRkjmIwvikc62qOxxyY9ObakwIrxSSkv+JE3mUodMNQu2vv570NQ
wPsjDMe3WJCAh5mfFYNNNFCu3hfnjnl3Q2Msnvd1ySbgutfQMNJzeicbVfbj+5pQ
I+kLUaA5o4wiZiZOiOsfLBFbHYunJusVslPAZ5vY2D9ac1aYHbYqSRJcXw9p7j8H
ZA1Ia6awLSWiyX2ObgpET881ENns+lJ9AKGZQV1KVsb1XiFz6Ya2Lqqkdk47dEDL
5Pmgp7PSOPUngJCBDRa8uitLTHPKIxMPHgNA8C6yiaDNAhLIX2XAcn0NHgDCYVNY
l5AXPj+DPfKn0ffJkGGxP9xr6SJ+RqX+zrmjwIo5fh48zVr2Fn4jdV8C+TRaXdcc
86YKgdfxZAAcIMFBOgk1wBbTbtmrImDiqiNxN2bn0U0attV/ErKe3AZHIOy124ZE
j7LlYt+j4+8gQcwSaGfOnMMDxM1zGFozWP5U2Urc9vEXxVeLpGzZbDGXmrQ/E6VV
cPi4ZJD13kwUdX2WcWU9xWLaOZXGQAaPMl4KG0pzjt5qk/C6bZb/zmUY98LaAnRX
V53j8DnclcaRMAEqlVZ05JVgQzi74ixdl7ZbATqlBymCqGc5/paG1MyP52ZEYgV1
T1DYa+21M3l7nWXvqDWY/M4aR6JzDLz1+TI1i4Ri7//6MZ6iSqgB8xcyoslouksD
sP6SD4D11Nt/6Tj0jb7hrTykFZhWE6FuAbUpYb895iUtREx6FAPbfUirQiIFbLol
nIp0VFQ7tG5MdpOdmUQvmeYOa73Y/nvjxFaeWdVuSnCB+aFxazn06S6AQe/P8TTM
N/hNtmSjN8B055lwlsq0kmAZHP3IEZwSgQCAuaPFsJ/BbqtTMtC1u6dGRh5lHC/f
x4Re+vujUjhrghpz292nt4k/yldb3vZ80F8VwbpJKsaV8K7yvsaOQzigpifg8Fog
qFj/sDQwZBOhWKGY54VlMShm4DpAA+Rg1sdDNtaaWCOhEkw9h7S61hDnmrRIKt+O
2VB1JN94bZczBQA9TvzLPNyboZHAWwK8PSgxr8c84WaPseAAtESywyDxEXDSHmNR
snnHVCRZtd9NM/CKthisyKv7ooGWAV/X9iyz5aXDbzdxjdTB+TX3452MUH7R4ZdM
CLWfrtN3GXPHASPC2q/XRGYdsUV9/Lq/ML3OZVl88DVNo6XmMCbeTS0UczJqJ1B6
LnQ5uTd62PoHfWFeLXuoa32AaUlRpnvQ0y93oeJLxl0aZLu18HNsBUcUw2pdcLTZ
m0oSvDw3Btj5b4TxTPxT6zNEo/zWcJYdWwQJDjukyTMGFaEisdt/uR9LI3Rc0srz
505ORDNnEvLrMKmEhPBvnVKv6xhwhK5AutYxFYM2+OT4FMmkwx5qRO0p91w95Gu6
T/yJAzwbhP60FByXM7+LjsSSaYyNpcxfcUyiivzseu+qe2GQGfSbaVpccaE2vIVn
KHaEYXo3GM78yUHfgSUJtFF1buIYkAlzN4FxGTGZXRVWNvikI8Gi6bbIz96jgwJs
6mcQRBLQvT3aQ4fJPIZP+3uQ8fueqM/9OMEKRGlLZSsn/3F+tlat4Qos2FaInpmc
Hqi+I1G5A//NmxiqUK0NZ69JveoUfqaRfHPWpG0VVOWvY3KTL05BeLfLVVKSfTXQ
wSmx5T14CFVZrLWHfeU4xYQZyw2TqnEXtMm6n4UoTVyKRhxhlW9PLyW5poYwwR/w
o9aa91QNZ3U4S79LIFiTLqk6AlGBIRF+SD+WBxk6ybIT8qOxd1YhaOdxRYRfjOUy
F+a8ybDKREPubTQZu6bkcr4LCG2RYj7NhAtvflCDG2y6YhyBUPQSvjr7ZAklwHQd
Ub7z9PiFDxijteH0oL0rHeU8C0L/uUIdSlz3vBkIrk2ztFsG+Dd7kgfxECS70DKV
arhUobGoyW2ifA+KHvXx48CDG0MXtiGGyaopr2lo8YLBM1JD41K9GMElGY8XAYC+
Zf8eTtr1YcPozskKySkIkPM7ODrZd+P4bnni9GtSZHirR6Jas761w2gUo4WvE3Hq
GlRoYzxXjMOPsiy0Bpc6jPGcMsR1a00SPJtkHOoRb4ksL+0riammxCM2G2BjSIda
Bb1h7/cS/4KGZa80SArYwmNcHkCYJn5xfRP4P/g4FWB5bLZJnZQdODp2MFDOE4io
`protect END_PROTECTED
