`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aIGyqAqG+djySQb6wwnEg0JchPEF3eMcCJhfS/lh8z/LTh/1CG0LV/7Y20iN32D
bduQu4fAleGeptKK2RR+hHiTbcdJutHSqFF8FZbrVgSRFraDori8+7yfvKCWvREd
BAhMB2A/5ciucqb0HqqtonHoWSgof4l/BiEyufyqSRgUqyvUHa93QEfenaASKNHm
GZtfL+lC5hPiZOGC3Dpsw4MocbTw+DzKZx0ZXH0qYMk5PiIdwiqgABSvpjLAT2mi
CyWY4PiVYEktkKPW764yxYczufpP/HTvk+L/m96vPHK2Vu3c5sn1qEC47koelI/b
gS6p9ChpwMbUGM1caHfPkdn52Jen2oIKXq6HBNtteIpMfxNJViBQF5QudlfMxY1E
yRR+HY97Fyl1EJITbUj/n2VzPFhCrWzowcDBHD0mKXoZ09pebYFl5HNo/jhedr9a
+FQGH7D9nfjn1UvUFhl8Ctc9tj2HD2BkrxmMqPpmT238sqUHqFr9NANd+n+3UlcS
7NLPHl0bDuA8+ASp4hrniRB3Ccb7HwDgDhiM6IWExOw2lCEmUjE7ngb52uRROQQt
ZPGG8fcKGstJqDVtkHo18Xwb6vXEd4M4tubjgVQMZopePRmTIsSCrzvWjvwzPqVE
YB7RVHSG1yuPc1pUiDGKdXARrBsRA88yJ6cE2sPj1nz7jxp8OXnOmw7hvjV6PfGG
sR1WR7Y9jy7lEyrHFZN/VrrX1I/SANEe034qTDbegIGvmCTOgrVD/gPU+A9cbdS7
/yr0UkfhQeY0KyofMApwfG8LqEpF+qjhBzHWHGmafWSh9E9YLXZAMkzTkgGCbzxZ
xT0SC1lBJhXtwgTa3vulbxUyJcoxilPQs4BhsWEW7J8vYPohublPBf07Dv2kCeqB
rBIErU0kkzuoE9XAt8w6keXAv60U2V2IxrODjofgG3/rVFEvHW+bu+2HJe5SziFY
pxRyv8o+2DeCE2+GHn2oaUlvTRH6fN5xtR6WCojx57YzrFabTTMpaiYTASZRuM5m
d+yaT/GNnVhvdFT2DcyNtA3CjLjXzA0b0DjlNZ6zzcY+/ciYewR/FWc10V71uQlG
Sr+OiFYeknJAWGt7qhnWy30x4v6dN725bJIIjN6rlLhHrZ+xqkk9A9wmzOc1mPSr
V4s79TXOFcaKZhHrJe4cjOhCPmn6ja9/vRa4/TE5WI84Ju+jLIHwch1iJBWna4OQ
LuSWvUn6CUs1mPGMzuvAiRxJkDgm+7TAbRJJc3UxqfAqQgFXGbLwCZiAlJgngM7n
prQCWR7vcMkLdU7MfpiWTdrzdIKfNuc42L2WgAFyqMS2DsrxqwWQYJaY07gHT4Wp
dEQJ/tjSJdanDTAwDxJw5/C+wnmJsMDwpe/5nMM+5BtE5KgJ8l9/VgbaQXy8/4UI
0fY8LDuks0rhtsXJRG1mmodxFiB970FneP4Hpdw13bSV0tgvZN0UnTldickVEsOD
Uh02fMvE4tkrT8D2IEJ4GsOmw7ear5I3wcI01Ac2qOZeyqTAxofjTfa1AEZz1ROM
RR2eAjX3Jo6/Wf+0P8+ftgYt7FRe5s70grFv79Qn5PCZnvq9i2UrSoPWNuFiL+CW
SxDOOpnrDwPJeyl3KcG+xbaAXnOIubG2hhtvpoFNlhfpEMyTpLt/P0FC80Ibr8gB
HMPJ7rtR7oOOD/ZGeemtb7jaxTR/ik38qAUO30dRU25Zb7XZ5E4/rV5e7zU3gD8u
OQt26h8S/3Ju3L+GJbA1Q5vJJTn00EuB0vyJsBY7/iVotHavmoBQnYVR/+8N6R2g
rPoov8glg3UgRd/FOvQCjs0vkaqnr6rD+QMBLXRM7JdFvucSqehJCwSkDFVKDnlW
tgqBFTm5frIM9rGGrP/y4syH4ItkuI4af+mb0fMJkC55XaGZDXzDfbOy46QhsX98
WBUD3JQCaZn66VHZJPuUNyMx27qUySRaHn8cPQ23E11ll/wAc9F+ZUsz/PinXGHL
/qLJpmnWz9GpYEKXCQQWCbcYvWkmTI2Ilb6KIZzlRC8PpFx5IHoLknJSdYwJqgqq
AqmtEAkQeNfKg+pMfpM2JQNyBvUMSJ+EYcDcGfKimmj5Y8V8KiujvmW/c8Ic7zYL
ZJVMpR320yI3+mhj33x2ECfYScSwvSpNPOFXvxdzpTRpo54Bb2imC43YPQwGFYRj
eUtZ/im2LdVKi4ppmV4b4OzCqRvz/DnErdvZsXNRfUqTjfegyOiptZyUN9L38Pnr
3HaQH/j++p4KaqmUdrokdGpsRr9JQmrnqn2sytKLXgaw+nJpCl2zLNqBOdSeMPaF
iNjYpS4DFRvcFAMVw+FlPzKYDw12Ub5oC84Bezo1g8GoUCSKWDcnSOM7CcdhCxth
bfALLPDMljpwdSyOCpZCwKwsHB3KEOJQBFK2E7leLLtkso3zUpGngqetcXbAM+dZ
HNTielK/Vgm0N37EnnWuUDp6mQjgxCJqQiyVj4WQCjoFvRAT7Q3LYSFSVVBeX92X
7vkQPA8/s921JpJeCJ892OvisUT5kvZ9Rxfxh44WDzQ3pdPRa3+2jKQoCKBoVcUE
UPXm9JyQCwYB6iMyLSUgWY0pjeBa/Fi97NnMfQ5U9+7Q5jlR7yrL6BXfToomVI0t
8NZPuJEgEs9nWcGc8n6PXaJrOm+r0tkoi1K5sCLNFo3p9X+zbOtH1FxO7jrx34Vl
1qcSkT8LoC7I9Gyrfh6q1FF8lEjTKEmAuCY6n3Jk5wH897QL/ArJ3NoEUrhDBAVy
v8DfcRYc7VnOchEfYtNJS6MWfE/zr9H16rMghdqZo5h0mHzgF4e5IUw3LGvycht/
CKzkvle6yoMt7N81RjPhWiaHaBhUSIEk199vrWrbyyrhQmQeaU29JFg/GRIuVVue
+wTC86MPnQn1WFHS+wVeBfIgNK3O2he1KJfSwRLxAEF9a5dDCpsJsRG4yzW7Pnws
F8P6BXPS69jeZkQ9HuB8GaOATRH4jeMINOYaExYm/rHIsS7yOVU0fdhrD6WveXD5
yfGZDWDyt+uVzAa/8HkjRF1nw6jlIhB7KzcxWNPP8+2SCOf5KadU73o5/aMJvdDP
8EThmCOYISJrjpJ9JsJTaqRwy1bWP0jLeT33fOnAEceLQTaTwJJkGqvTr0A2op9S
+XKaT8iCZoh1pRPIMA2bgX+fd3EtlUn9MgOxR++bXQ18VlH7ma5TGwaI7mC1Wvdu
Q9pygo66KFBFRtTkoy0IpKNQ3tthHIaXUFTWOhOfnMhldCeE0/9+VwAb0Q/CB8nt
Me1/A+tZCcB2v7urEcs7xTIzBtOVAd9a70ibSq9ztbk/OXIhLp9XAyIfJL7b09Zw
GW80VQ/uKAeOw5L+QEa9d1wVELJ9D5A7nq5agUPB+4QKVLKtMkXsYqQjMXAsQzU5
RrzWODfTlvCing3lzEYkVjUFtF49S501/xMkWenJiq/LWqlxLe7OpFxn0FO3sv/v
CFiRcb7rouIRmKuPOdkErnq2N6v2xAf51NaqnTad9IaQetBnEwj7itfPUztMga8v
/JYEzR4kci5Wv/J2ZfZqjIJAlTsn9Eaz1a2pXhVa0nJXfYlcK2DdF2UWOssAuSAw
3mpgFwbImPxIQyRzuO36ek2EB66z81nIL7M9z+K/YgVA9BdO22A8T8RHdx6tD01R
oTgM/48dra5so+85glYgW67cF0m+wIHsMxtdrGIb01idHZnAOuvkeE7t7KRXK4Vr
ma2VbazSNx1La0CmbNnNGRlgF9YOw2ZC43oR/bCxxmGa8gWiwojPUQ0FgbkFl4Zg
uGXMyQ0SAz6vfUUmcP6f90kC6XaAWAwbqpUz+pdRZST63ZjJ9J+/2vBKDKxUOWUj
9FmOTGQnkGzXkLM7V2o72/KOc62RE8vg+M7xfO5Kn/gzBWQZiATNzEBvluXsLlFs
gnrD9431WisS+qT1uJc9WvyFwr3Nocq5HXGqSrSF8AtW3iQmp8DJwBjyq/Dwu02z
A8FudTPdMxKg5MV/m3/cdzA510nQ+8P4ZI++BOoJJ+on10+mP1ZuI4tij261b3u4
0C+KoWkvT2q81pN7Ya+MAiQZ2d0kj7LuCkCwxJHADGP/XiMOxlBaJKbBMhUZDAUy
5sc5BvrHacP9ftA7R/c/NnStfFtS0NaXUdD52u9iXmmkQxLPEmDeWuq64FRyjDs8
aR24ugxQnurFhMd17ZXf/LII/IY3e6gr+7X2rL/IaV8ufzShFL0em1OuU3jxUkGG
kich0aMSEXpHjekeOrMBLpEgFEYnaACZflPnH9E4a/seUkPsAWFiSJ9CecmTnhA+
JZvChzSwHr55uyknCheYely/WwON9azxPROEalGpKpCvwoeiguSayjmoM37sZ2sI
hL+evPLWA4ufAaI/BUJ9GM5vZ9T95n1P7APs76UCZlFKqRG5SXuu6Yh5G57p9w2m
MsT27DY6U4XPLj7lADz5/LwSCLp1ggO1QVkO/TBqmc9So9r2PwFkg6gPA61DufO5
Jsj1LXJNHH4OFDapIiBqTD6Q0FNNasGuS7yV3lQ7f+Sx/5SvpPZhgNp8nP7ZibmE
kRyLCo2vfhd6uyeTMniEn51hJFLWoU8nUnHRt0nHX5ieJeQNXnjYzfkJAXgzutiE
AndWbWbWOM3nz2HHCQVV2KvtpUcC06U5iQjWdI9JpT8p4jPM30DkWPwmR+7LDUmz
GhOTcuVWqfG4y9WJh5UhBj770QTrj1y2cXg+SZKGFLcmVR5yOeyuQcGyLdw8if2r
s3WMJs8LBxVu5SRD1iS0Ug6nO2ByH+uW9AXMrJRad2BHVn0Nh4sNbReG6OYPOYJg
cr8RMQv6FAN8QIsKbLUtm77zHMfINsjyfXpKKNqN6QDjuVqANRCuVA3WdmRGarPp
sPlrQTHr7PX842zY6OO8KHLw4zEZDs8mBMbngcZxJR/F8q5y5TA2z7nMdmrBAaif
Asf8gR9cIfKfNqE50yjwWdG5h45DfXLc5SNuc+qO+zcW+AfACY7Uc7UatsqO1fPj
YvuLHIlQI4qvG/bVnot1/5ySRynflJPXbyES5isf60ORtshFFqICdbNC0FO3EMsu
Qu3wFKot5jziNHcMxkHy+41xk4Q5Csw3uSrEgu2HTce/f2mx1L2dSbF9iIKKWVFL
ENm06iucBiAJJRdEgrgxpJCkxhnQ6UuyV3bo9bWGj3yv/vYdovVZCv1on7Wp6YVj
m2Ft0R5S3y5pzvtGTA7fLIhI7ddDiHe8DhiSgucbMYOkk6iHhyWvP4VeRv0NkOsa
02gKAAWjD3ggKgncqYL99X2IX0XcnHdP7li1zMIUcDWK+UpMfk//13woQ4eij7ym
uiWUMNGrcnQNXHV1ZNCpr5Frum4z5v+qzisT44JXV9CBMDj0x85R91LhB147849N
71ZAiszmGmRri+2GfFGAwEyyuHuR/FhW7NrvfNuxSECbrl0HCAbni4Xdav0EEN+4
RmQBbMHIM6JpG4I2D26GMBUOUaUtRqc6TvJPeT+EYt/OSwGGPYeSRJp9ddGtqJOP
/2NLK+lXHt+f8RAzwrlj6hGEi17pQTe9+/+5CLQgQls+2QKWmV/XhRrSbw7izmGc
L/UbHIY0RFYnQb9Yx1dzgeNxRaX6eoDKCYljw9pro70dH3/SHsGWl4vp9d8D7B5Y
eon4KgD1pWSqnqn2g3dES7lkvi209qJAmRQ5h1vNDAgdC7qWoUpWEXgQcwkcTa14
RQsy5IFYXnL1nydYujOlsUlkkoU7Yu+mu/VtfTC11J+CN1m071wPbS4j7eN12oR6
m4JDEE2HdBucuD8csOi9OUQ474JVKxdSjC8/+pPhVSsjEOPUi+X68N5MfaBAOFBX
w6OR+UmD5Wrz1EVkDfIVQvMJtA+eKN/sOSDSpKwlQP748EKrDhukhd56Cd5ehSQ3
OBY1/Gsi/JQd899x97w9pW54cUbjIf8iNrsP54YVtbmWVlVrNoHHDJsD8UPNAnqu
pkPuQ9HOPYzN8rLU3I3XeQ7eaTw6SWjpGlo4Sb36Cdy0KI6FsUKfYBtnkw4cAcG3
fKZTuwLXTzpK86amhRLYXLu9cxQZZFKI0Ywb4y6jcfE8wCyCkF7jxtqxSECFk/to
g2BowxKiQxPt2051kWLhfLKPhEGqwbt6HvVl/LjpRjk491Y99rLkVZCiBHAHFV8C
SwcsucGETUz4W7kFJGYIMOQrCOHSvi92fadWOT69xkuXF0Xxr95Bm1Qo9cdfUuG0
k6hjTsks46GHqUfSKms/aXEsT1DbCySVuGpatjw3/KehasXb2HXQNlGafUZmXA9s
LbYzxKJNfQGJo9p2YVrfhmb/FVKD5T0fxrVZ7ucAzooxvA9y8fwDKWXC0x1jfhoX
HNO5yqff/vkmBNRMeg0xi8EUhL/F8d3rI13Iy706ASS80slu5ecGCfRAcdqebvci
wjXlqIKkns3pJ7olUtTTcKwWEYNNhNCBb2ZZPUsqAdlzpcA8ZxosvwnP8gCzDJf7
7+80mx1bOStiNKoZfy/qxKPK6gNM6ZMNJ0eqfTuvXhRVSV3AyGTSyDvH4gSPL4PI
DSpmBdRU7O3rLmykwBUcLgGeSjv4n0QCVd3SYfy+UHSE0ziQW19pI4aGgmfCuuwu
JLhIyYPBxXqsa0PjTjilMjm0TRPCcR0eXecIc8pHc96jRuZZdW533hBaNKyIk7Qt
v4sNYCBx7B5LqQcBXL7dWL4UrAgNKFpuGLbe4Wo83VVa/BSmGrdSlWuBj29jw8k9
0hmqM6ImfK1HoIp9OHRGLn8klrKW3qppawYwaObv7GhpTFKmTxbzH05qnAwi1BBa
xoYk/7a4WLxqTajk2Qy/hCvjTDC/ogf3ZCLCK5kpvlcP8794i1vGZNNOLtqclUn8
vajBb3rZjjkb8hhLisJwF6bgxzgAdrl19xx2pKXFd30R5gwlxBuQHMgbzln6mArK
XnbC1hjJRbV9uEkqeLeCjI+2zDoLYW2ELMvz5hqw8wTq33wrE61GrhV86/Yk/s17
y5mwMiOO8xCRmNIHAlCPhuQpggDKXv02r8Kby57A1yPbz4nUElHjlLuX38cExz6t
/97ojdyrN1OZcQqEDwNqVcU7KsWWLXLSCp9PvLW6R3NpBcMNb/Zt3S/X/oaXFCdH
wRm1y5NvO3ymJuVoIO9J5oVyZ7fkxDC6WjgGWyYi+6Voa4V7+j9bwhZXRiWOuyRM
adyXBCmxRMlMMfcvJn9ZS/Y7EVmP+4gSC5njvW67wAnU4eXqP/qNuG+/kvT7gsqp
jeA9YsFr5lMJy5RyADmwRa/PJZ65XnluaFsR5I0rfd2+SZ5S9B0jTsx3IOG2RhMw
f1kEMhm2m3LWRARrVMGebemawequAZwiJgGX5r78L54da+XSAPh9tEbjBShMA7Rw
66RaHL8r6twknnmt7iaM+5mvUKCSoIQVgyIItc2i+F4lvLLhL3ldLLptBzaEAu7J
x9aLEa/tFK7q26/uSukLRdCGlGcslnKymqsZQFJkn6inFDzqoCqf0pmclJt2++1Y
AvWIMqA9VSFNF0iqUmPyXO9KecRX7pNc13r6MjYo51xw3NO3S6I/idNVLQlQODVD
vt9WltaupOsH4I2u+lGCepyNRNuJOCWt7zABOBKPRoKE7JyMlpklu7PuzmxDqxrY
HGVpbIIJOqM1A06rKwpGmS/8CjOFYaRwsLvGw8ahkWOPIa2WCbAr6Eb3m7TERpx8
28oOTQ8SBeasx74yb4NGNk+GnnBU2wrQaT0y6TmwXoNZ22XUjrHvlvLp7aB1OyAA
VCTVUuxd8XxcXP0b8XAZfw20M93yM0+lsV5s69UFacTHBfCghlQp8w4InNCbxSbP
6uvFf5NitMNhaaI4M3NGzRRKf4MdM1ihHK53UQSCdPdV96NMv6ZZme4MJx24BVNw
H1wwq4qcksVwAAI4+axD4T1ya5mu+Y6AnLVJXbplGDGivXtjO8Ap0zvwShNdpcOo
SLHZm+XsHKuztO1Dn+YhZHaPxdM4CvrL0GUDXQAYJrRtm5ckvo8+m3n2ljYoOZeP
psdP+Pan4r97KRfhWyNYImCUlvqBRQ1Qp1m19vRoHUmjEDT6ESpJTmOzUrmbJpV7
PYuiYqUKhTO6bnSDv3R/ZabyiU8OTLa6yKrezFJVoUWl0SuR97ZFJc4r/Fzwg7pn
zXFo0smA82z3X5/WpqPVU8evDr4q8Ew98QA/hhlpTHRaDSDaeojBNKFWdNYeN4+g
HI0E3DbTU2XCngckqG1N+B1ymcl02I7kY7HJzozLcIW0t5dH4LqeNo5lx6SvFgR4
IhNfc2UM3+RlEdwBwFXJhvKZfo5pn0YBJTKej8rD+62+Es4oQ2p0eQuANS+iJycr
flEzcDf+IkHeCbn/38+vITiEUowoIRAMjB11ABVPLVvj1hjKNLNUbX6BtP+Lwqha
2djQPORLRhPgL0pgMb2uPwQKV+bVelaOBcWGc6pIXOqHcgUQLIWlFYSXwZDo7FPd
/TKB9J4NZ3cqrwSA2g+prmeLoZPk05AJiW4TfxPZlmziROaGcGr+ly4n8AeeUt2W
j7Nwda0ktlctqZT9Ywxc2f17oSODUMQPDNQ0jVjlweJsWtqE9CX2H4ZxJbirxMxB
mafIm32LlR/dofvOZUEgfhk+pxpkIr3LDILunHk5LaTyT0qb+cGQXOMVEs660vte
X9Xa+BbBwMpt47pVed8E2wsMvYGylen13NSmtAhRzRDqf8uoDGBYk4bG1S7No1ko
1LcAM0GngEkgU3xqL4TZXAEPPEr03QmGQnjJll67UXvmn4CT5UF5DEYRBGjlp9GA
013qvyoWkm71ei+HHwJjzFli495eeKfW6yLkG57eit3ST+IALoFsvSwkj7UXKAJg
f+bAUjElBF/niMBuKJKfa7t4qnJrmv5RRsDcwVwEjv8l/9pj+6kfI9gsrLL0hHkz
BKtNN6XZO9xbgz53byYGWb+vLGM2FCRV39134fqwJOoYz758kVWGeYYof05s+EHT
j1JQQx4YqH6slfu942NGpP6om7qYpRsu09cQcitusHAatAhmZS9rM3oT/NxfzZZC
BBi7CaiM5meXUIUOroNsuhrvdbj7x55xa1hhzgDxiye8xdIl7ybK9DL2HP9O/1s/
wz1nFbc3nc4QLvMpKKaYIEEzfF4yXT0xUyiC+womYCSr1wOrYy7R7XI5aSEUA7JD
b78uJspPh1Px6QRRXpD3ZXvOcW2+Bycnl/riDyZ5XN8Kc4LCo3FvQwXL7cyrrePe
mECS7iIpoNlcmmqfytszAIZNHNSqQ+CpK1HG+7qHk3SeObiuCb5LHEdteXRSC+g1
TykIqJYhUc7zuY9S6SSjbdw4nvaEWrFwWEnPH6TKSN/22kApD0hiW1IANu9l93rj
PnyrDLFrJLdUmFXoduOP+HAJxjBavNIqngN7qfKPkccs8HHfkdvsqnvEYG5VqU1w
WLs06LSgJ3qc/6hDVjH/Hmnk6MHzo58x8et5h/laf5AmCi9PXvqs0hPT2opdOCpR
sr1LrJpkTOr22KHB5MIBpC3pu/uFGli51PcSAWwP0bSUmI5+vIp67NpcbErZ9rCe
0ZNOGMv5S4AE9lCuJES7FrLmAQC37yqtNshcVc9RQv1e3dGVJlmEcm3E3bAyxCdh
IkYrdPP0cqXbfCcvRCZ6tvBBhEhR2fT1IUG45yLKEFqtvTMU4ch+yjg9NKCd9zFy
OCETvrEMrwkUV0qkR0cPb4m3ITl5FIRUiRkKXK28xtWNWl9O79snxhAiB4neHC8A
xrf2y4lQIaMfEe3UbjOGNrReCdwS+9WxtyOg5SbVjQWon2XbLCpfgMU3X9Iobkdh
ETZyeYC9yBnl9C6ivoZPmkypLu+bdOLyX/rfJU1VsoU=
`protect END_PROTECTED
