`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tX45Lo+hK6LWF34V8z7tC97cPU9oL0/KN+pU0BESjf+iVwj2V3MQBt7BPuwky2cY
ok5AASaehP6x+Vu0hCUfvot9u3l2C5yskP78QQMc0J+27ATfuiBK+Qlx/VOBiE9L
PdDEWhX5PXDhJSfrHUWrZ8XRDST+LDJe2nMhfp5nFze86J2P4y0rd72/5JF7ahed
6bwkHNZv8o+KkJcg/vRWUkNRwYfBF+elINUDWckFWwqmqqj5PaW/46La80xtFAkg
s+8yRXWpL7n5DpOxn7Wewm1axbyHO2QmDvHUl009vHQnou89+8Vawwjt9sHhHZBF
mTvezSFbXWKgeepj+np6LBSI3D/BHsCgnfF6kYLqG2WYyTSux0OHkz0buIcOJvxj
aSg4jRA1YoLnj1dYdoz2DoTfG3/Xu17squXc6gOm3RohvvmWF46ag0vwPvDmwAGH
Hs5UVex6dE9WL2sLvX3jH4SWrHdO5u/2DXZyTJM2HfvvQ1jV9lU1z3P8siyeLIEu
eoAua/Fiv70vXWZWhVaR/5Aq0pr8bGWFMF9THhiTtXTmNIcVoIh2ACeJ/U9KXfKu
73EhADX9r+vprv7iWb5Zs4xMX1FFZ+yH5StYXtW6NmFAzoTiuzJhJUH3qblWxKXt
0VEIfSL/0r40zbrrDFsoOHy31P2wAPC0tvJfNr2dL3SxzHmuq9VcVe0OzuJI9qp1
n1/6godhu7YaEMqHo9MOTgGUX8n6R43NVQvgGsIV9ZB3+NoKJEMaTwPAL7/lMZ8L
76Q9CQJamg+qBedFDBVqgFF2dxj6wUjvg3OpCOlcC+mc/ytUjvUUQe+0Tth8IgU/
gS0urmANJxL+dMJkjLDOdIEUr6ddZKXBBnfkY88GHANlLjUSsCO4fpTarspTHYjQ
D/YfUxVNR0eaJxY/laMFtzSHdR3+SDanLokU/jNb+CDiLfB+hgFu1dkHKb8lt9G2
zI6c0CE51lhnsIMZ2nuWFGVceXg5+w+0gR9KH5q/1XIe6Um7fRhuMu8a7tyBqqdT
rhDG3IMqRqjWZ/Ow512xSrvtvTr4jKFGI/Fruh2atOUs0Cqon5lCyi0HfUWsoJ8u
SnMagEpqS1bH1X2ZoQ3K6jCd7t/dbhOJkb5ovqh9XYWNKrsphm1WNXGT1nEb6oRc
XUw0L4tLF77eft0UFfuq+eziMNX6Id++zrVEggr0MMUpSqQMv58OQygGVsMBtX1p
Bby7fu9nAmSNOIHtGV1qbvzAoljPtOAdIR/VLKWxR24nMlDNlkyqO8UeEziB+KxC
9iAEc86y6u3IQnVYSEBWwUZU8B0b7lqcR+5IEyOB+oIksrih8JZk4tQEd3eNdlfx
dvqUj328eFyiavRnI547HCZ9hptgh/KXDh/O2C7gDqAJmi2WwbBDEhuxukTZBDQW
cdWWTcMuMkEwtzVYVCuBWvrICi0yYJxUZ1mtgtncLMPrIawOhJEdnSNL/t0GInn8
mY5myUoCeFWuoVZikb1BVAutIEuBE8zaUkEjdyYRIP4x6vHbHmcZS/R9JcTfKCQh
LsPbmNsWXwTwgeakWzkBGeYfGdMwPzxO+zuyII8j3p+n2vZpe+Y2fwiQ9iz9N7Mv
/6z+JFruLBIyI5a6xk4Bhd9DPPr1NU5wXyizBy2sRJK297vonDoTFXoLka4UiM3u
vcJlO5qyttChIu99pcqN6YYaVDQkN1hyYgUQkJuK6XzjTA3EYqyXlvX/0EUsuQbe
JDxL6XTDMvPklsEY6+kheo8XAbDdXjC8wypi9l3QEusXmoAGTEhkSxBPcn3aYTlU
P5X0BIzJrN/BJj4Vu9PNeuM5EwyF8F/SqoNxhZSM/QJUL3H6b1oGHF+UgqQ/QTcX
iqfS9xGjQd4f9s8SpeXIx89M9NoeWSetFChG0WMtN8Z/zMAn6AIeX0SAJK3FNDMU
NVhOxlAdLWUI8PVcH+5HQEs/VC+PWqSrq7JpG3+7eQzS7T4MBpRKmiAhs1qP/CSY
4QlcbO0hyM0YzKaLkfiL3M4baNKeKuxRfkD+UPxXM+YbLGqc+DsDln0E/c3Cus5g
2ifRTNXrM2tJu0NJiTp1XZX2LhV+FmT5XOXVu57oqLr6rWpIrOY/5znure9SQspn
nO1+sSertUiR7K3r3o8pBqRQTu6PepVYVRTynMT20/0UeMIl0dWr6MZ31b0ihnQY
7vXLbg+5WGM7BDWQxZGBwRmlBVS2K6q8OASWkEajkFHic5yDP/9iVLFLkCLRXZV8
7tf5tzj0DIO30eLM9hsmhTNa23BbsFwjbs2+En07/KB/TAeJjwQhDEZlWQ0+UA6T
Gcaz0wd0OqCEq6XnyBh7orHMpbRkEtj//nD2KW+h74V3ba4koIqR7hTEMhFW3btL
uy44L8NsmLKmNUC5Xt19JoCZBsLObgww0gjMgiOnwwbNOK1+CtHo5vQ8ISM5L5hu
+ahv3c643esBGt4j+xEgl8McxVIVQsEfXnKocQ6W3Nots9YCwBiM+mpNeZdD6+zZ
jK49bhZyMxf+AK3clVmuWD2R2YA1husyh4djjHSpICT+dFeB9H6o321paHaQxV4I
mXMZ8bi/gorzUBTXvWa5amDtE2Ym5IXcpKQ/myAqZhJT/Ujcz5h7OUQew1s5uZIy
yTp4yUt8eAelCcw2o69Ts2iyyHwVU/TBNTisa5lqvgklLMXM05uoiP+jnGB+XvLI
klo78P+p/mQ9VLVk2ZZpVAXt2DGI73l3ZVVC7/13QkJj9CNWXEeJurrr1YEhMMOh
fh70GcBEPPGKefKPtPk/JAzqNEeQ1dLv3FYJFEKGIDeKrxBSIeftG6tsEb4AQms4
HipupOMru8DdS1fWh2ifkgBhDvLf5W+kpKPDjd843Ly3AwRQ+3cHoOVU6qqNz4+R
wzwkKWW63z0j5yK4Om5THDAnOedJAXMFxlce2D5vBQ6/bqzwyaNVNEXDCwxfSC6Z
J/wFOuNHnyRrWcDRdwWX/JkPaWX2t/OBH3mDCtcvogSSz9GNhrzLCM5061W2rYY8
65CWcft8MXL5+qc2yGM9THJkKzvcmmNxuIkGJ9wLMTxVGKW+LgosIx/jf+2ftcbQ
XqrI6umdEB/izPDwIF5zDVj566idWfloOehOT/med7KKdJ4uTnqBDFnrws38MFgw
xzVlhqtP23BhYi8axAG8vRFfawPiT2CuKKLaFuh/6r5XweOKsYlIYcF6gAwoIsKZ
DS8koMYsKK5g/z9MVFLlTciNgOtFI0NUc27meTMd16/7F6JpkKImORrryr+4aFA5
BTMiNC00mXu8IVH7V5jsJgnCpvS4SzA0vcQGHIOTJbkfvFURSLrP6Uui2hjTkGc+
72pEd4+N3gDx8PAHJ6XJ36FKTUM2J0yOQsEmaOEwgnwoXUiOQq42VCNQ20aQzmLb
lCkTUyLGb2OrFUUgs7PBV/BvWAHiG0lRY0aKUKA5f2QSz+9tIMoPcV1IePpUupqH
FJ1mN2xCLNOvqOL9pFwj6N7sn0hKBHvqoDxLQhnsBQ6qKeYfu2zBSZ1J7yd4lwqM
tLmFmnzEYRIDid1dqBAVrTMJ2PX7EYwzR8AzdWkJH/kaarHi8qIdpdO0/VN9HeTL
oNeUPUnKP05qM1ph5rbeR6ha/siKMUBdZEjJyz0K6rElBZOsTA5V4DhF8+P0IQga
rw/ieYWedapEt8nQOGOIRl5LpWKCiY4DiPTebW8vnFP9izxzxVg5DCq1+unMTtaj
DbrZWjISAvRqhmcGitf/Rm6R6Dx8XEwXD+xv5/+JMW4gNFRlDm5S4yLvgqvmomQY
EedKi0b464zlM6tuFP9YMpSftBHI33DMH6siBrt3bbaZr+0gA1aMUynIWYkqwceb
o051E7rddOEotmQJIYnk45nq4l71Abg3e8ytY9dNEV6n+L1+CI94nyLpvis0e0YW
T9djomS99VXPJxdV8YcQWfSm3xnrfDTF/EOw2gBXU8TEBI5+lK8wfdMy+t7dkkZ4
8yPL1NMr+XrWKqQh1J6OeoftHhDOkbYY8RLh9w2Z+CBGuEAbNojAkwxVcI2PArt0
ZqmVTOF5iUhaTdoPfwUXr8lGkot42kQyuOwhTU6Ud15MODNtch619VtgKLr749Vx
`protect END_PROTECTED
