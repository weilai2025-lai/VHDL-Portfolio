`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDl9yx8PO+cc46YEgzHRECYANmq/rY8kaTrKle/xXLkA6nOCWtTOU7M70qaAg3jy
2YI+NvWI6am4eZtFOXESjnn7fvo2kfSPAwP5zaTjbuKf4VN4W/9o1jfzzFVHwXP+
yJ58jJoVbLxDaxVfKYqKNdiV85Fxn9nUAgsXTVShIGCSqTAIe1Tg6IN1a5dZOUXk
JWMRg+je4pZfSiUm43KJnbSFZnaE0siU0ePps2q0aGFYgUcru+fiNutHTtgXunHR
5iQ0rh2ABK3dqH7916O7+j3fIaFpOimVTS9rjAYRwQo6FZ465QIXJfAPc0C5jZf8
DN+yq4bX98ylNGDSmPFOkbADMnhgHjo6Cw9ERXnRYgcbcGVUmNatSmg7SYtJCpDY
E4JcuiclM8gC3TEbWmfGgD9bX0eSBa2KYmiTv20swKmCm4IzIxtjkO8x01wcr2sk
fKjPrWU7YYuKbwcBhxR/TSn4+sqm+A4KuVX9clZfki+l3CfUJanRSxwTxWEeS16E
4A0BDLtfgXAgrmqH73FlX4CmDmqW6Pep9Frjzl70V4WptG0RqwCkXASed/IaEV9u
J4950FJNmO6qwatOfWpmsLQi/bfh537qi34dVlax+/XjM/fjGY6ATTmSvZtRXUXc
L3exmNGKrArfT4Kt5T6VxXzc6BQd39awonkvEANhOMdu1Cuvg51EanY5AXpgJCOK
muoDYjMrSTDXCm8uSuv9mcpYWzM+iaCdk4/Y94/clkCp5t39oDX5wwiplevoU3db
NmIAiaq9wLok8CbrjrBmf9e56lOYY+FKlCCEdaje+kZK8KSKt0qPl5eHcXhheRi/
BcwbJ8PWdRfFXWt6JK5oAzF1WTzB/GaaWEdq7pjgSrR9aQJAbwT4Eravw7td1thc
ZgkT15QdmeQAPqpIWrZ19NaJMSdJJjuye18KIJhXrmU175N7tfhUVSCu/IwWJsu7
NbVPqu3nIavD3AQqvwMEnLoSNzP4w55DGTVFYjV5GTGnKi7ui+I1krpBifpdvMIl
vZa8/ajpkU1/v8N3iKFhrlURh30bWutNzFiEWSxcNqOwZ4wmyr71zYH4lF5Wyf74
PY9RuHe4Z21zOjcuLQhEYGvxVG/+uIJBWePWYojInJmOSnjKh7Hw8SFveoTZrRMB
+N2/i88v1e83qfqp95551Ed7YCx9O9CGxQHI5YDjaatn5LT1SqvMGkERwI+YeSG7
+3e/3H8fADoz1x5/GuPMr1afcwy1/ymgbhvI6bchd2lkoWNCCPI+WOk3U5djKucf
Nw5YDGxeECrd0G726mKHkMiWdIhg1TOKHIBSp3JuJMex4bXeQ+jbvxhJeRR8BHzT
4GUQ/10Ul/uwnI9+X3yj4/LZyXwU/N2oM5cxevBTGfmPWEp0p0AskWQ9oP0yD890
zRcKxVhvqicHVaK6RAEpebYhfPsPxnmsyfKIoLLNXKqwsMLywGsyd22iMv8iRv2B
tqljx1kf8C/3eO763PuQ3N1bRWZUcn2+OqYaFIqRpyvZ1+B8ZlfKkTi0c1tqPQtw
`protect END_PROTECTED
