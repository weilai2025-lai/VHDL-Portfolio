`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pwX2cSliKGcubD29QZ5tcPQpkmf+lnLQJRpkQCB/GlQL8SfDOjjnBUowZ2gAvh1D
No9p43idcLVfLeI7oDkQP9H/afCaMJv4aNysiJXQpRJ+wO+PUhLW3mBsod6JU66F
lm5sTDgChyLIBZ8VkybZL/w8OKQ2IEMoE1EbMSzvnnJLDzQl9rIaBftp4+EYpucK
aJlnEzvFS1KpUYdEIQOxx0OTlI4z+jwT4Ie5C5RP2xODSMY6h7tW2SLi/uxmpL06
Naw0wWnpfG/7DLSMIOuD+khoR1Vjob4GVDPNwVspr9yB5CKKba/SXJSuScpsWQCB
RvCimxCP/DGuAygYFlOickBu44+NFbx4Ax3YYUQ7p3TKnZBdDZ6UQFvn0jZmvhlg
AiJnIvirSLGllyUFAbvf2OQMerT1I2TR+LfYS8SsW8vCiOQun3jFkKGcc/B6DSaA
g7zMeDJvlKhQ5WxRV2l6o8M32a1tdTnMTQYJLOKTRn8J8EXYvN8GGRutGy3ACOcl
2xpNk+DxY69xFLy4X+byXdOKDod3mM0RlMeJWNE2fBiOtWzmbM2sme3ZyxE5/7lM
bX9FTbFH1qo4yCDUt2EUVhR/npMOca8T0+iJ3+LwkxRki0jetTQa3W59hxB0n5BF
MTl9EWYuj8+VXh3FOLu6vD4bMt3VCZLVgcWDBE93KC7bCiNeImvbknuZIfUrF3hR
k9aY9Trl9snWAttjm6FtdGZo7lE/NTHWR49DMRh+oUneq09ujQx97Jx5+I64UI/4
aPowrsZzNNaTz4rJsci+ge5ioHevn2K10kAytCPeQB+PR5W9R4vp9eHcy6dgGUGH
BczBhEPa5bRat4hf9a7k7QWPAGaCh7FU9negy+ypi36vBXZ0xcNp9m5c/dIBsO8Y
n41SXs7lDM9pR1FhZxK2YRdJYl3OH+ONlVvX8a5p8fngqFv5mqCdP4hada62Kz/t
3Uvt/2N9wbOzUk/6hDN4Fq9StfJWa2rsACgqpVvjYRH5g3XYl8VmMavHE4uM444H
CSJkiG+1+SKkYNZu5x0ZbGA00Pah03WwYNvGaLkf7PBv/2pG3DDqNn7d7+5+jWtN
`protect END_PROTECTED
