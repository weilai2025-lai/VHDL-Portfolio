`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYNmT8uYP1bgSsGtlBfiAASY7W2+ba7+bM/qo2R9auBop+ysHPJfd4G+A/Iemv5T
1HUVmKGiLAo8FdKl8HBYOswqeleEIJHQK9UpWRHDlmjWLGH6O1WexO6KS9ycsFXp
lzwdZ3Y7ZS5Ek/RkOekgwcq78FA1kDaOurr4A2cJzAGWllsXckVeKvCM9oKevFM1
OCSd07mOoXdArxfo/leWrDI56x7rmGlfzkdfyw0ZM6XHNcoXcgmcDGe26FkfdkAE
8SqXAjq4P8/N9g2f8/QvsTexVB5UmAohG9q6Vyb+G1TGpN2YV0cjUenMU4e6TpZV
3ZSm/azzQ4x2dRKWRwxDED9gNZw9R03ELO4swjrjErjhoyJQEdcFylwh49ojjugC
IFiO8v0rGa5uXdZHFMaT6PECdvX/Zit0QkQsyOzW5GFDMtRTvgNHzW+IPTHB0B+a
DDp9wvM5D26gMnK9Ej4JMite/iUV9pOMNYA/K12UogUkU3+oOOVnIEgaa7fZfOC6
mY+C35mO/iSF5OjaI510sIKvgzZF2kc5CGfaX/QRzxJcSgjmN9J4wIZZ9lXXPXlp
Gw9C1JSYCncWFp/jKJxgwn1O4Dfd54dL2GnxCAn/PnGS/xNPm0IdxR1quG3I9Apd
Leykjya8/lhGYcxWRJm1QGSR0ECCNKcUNJxdFCg0in2e9mKcIbyrNBFjCb1oBxQ7
vMmYQu99h2SbJsV05DQxZrsidhlRxWHZnBhVTEXkeQZywiyNrd5zSHjQQYXHt1Ep
IFymDMVUWGGLjsLwgWvkyJxpEw/Vo1NeeWMhV+ckpgPlwwUUK070TdjU5mRP4Xl5
WaUbW26ZgLO7R116eAazx/twDSq8ibhCPGiNCbSZJ+x38T/0NXlYh0w213MPV3sb
S4AiNeqex1sRiEFtglEFZi8N80wupKoCRcjj0VtqUbxhlwd+LaCFdDYey7uTCbHf
a9TUl+/qxztHK1Pg7OlNe7OH4OeyJ14TNbcur4TP1Yg4NGnul8iMu+deXu2XrY7M
eLvacB6E/PNvhVKdsN5uQGCdYKffub72l7fOCksykv27Pj4AxaIkmSSl0mgGwsdq
hzizwX6w58B876sJ2Ib5DDkb58efE0aOZNreJNSgDTWoMISuTKfmUzGmKAKY5jB9
xSkxK4IWrrLY31XN/ZDeTBzrfermSFYTrZ7eGwc2GSgliE7VD0/q4jSdiDB8OxVI
VD1B25jUwGeHwqPjffpbLITk3/7ztijHOmsq3cAcLYDAD60Kjgk60GeUBW6AoQiW
7N7XKTlDifw5IdaWAgRUqZQuc8OClf4q2ql93YmCpGw7QrTscwVoS38c/poJ64x7
0UtaTDyfPrKc7ZMXVHW9BIEh0KCXLcW34viwBHojfpSKfLAT2US38NTnT1S5gzGn
du99PYXgsBz3wTsq3TrmY33tynSm8aa1cd8qwlIIN3dpntmtZH/t43TYRBkiRZUy
OaJkxssIMQeXbtAFEKQwXG8Ita2vjEPl6uaq7b9Z8vCNGsqrm9WEQxSAjapOllCw
v2dHrwUvL4t9aQMEjvo7Ds4sKguSLxVD9zni4u4Hemyw0ftZyt0PHEZXST/WRcQ4
DTwrvo/qWHH8U/m7sbpDw7uHcldhreXfTMIehGkiXBGC2Gj/IyRuurbZrMHGLvno
/kx5gDLATanfa4csJzsMvOXg29uv1zlsOwge8yp3w61Gw8LkI7Y4wtAOGB1HAXen
P+d7qdO8FqENJ/EL/o4rSHqGlqvIO8qjgIzw5RTk5J8kGoam4e9gXgoOTJcSmVsd
J2BiIZP5OJBScGjGjIRsOAEI6LeHZh3AeeZVmIx6djOMRv8a7sNWRerXWTpdYUQ6
YoRsP4kwxjT+uZNONT2rghYnAd1Rz5jpn61x/ocJwBF0cqeYdaqDMQYGPWKrKZh9
az+MEc8edENkItl6V6UYRS/UNt9pH5KsjeIV8s89CEHZAY1aD0KGz0yzZSoZnGh7
4ey87wveL8izrHgYq/28MIBAvl/jiBAUvGI3HGdx2Y3RdHGwCqngqBnSLtysNwaT
XKH7GSFtdAbITcpNV3+gWbok6BUu/5j8XQotBKaE0nPAGR7KYGI7EoLf3FzGkYkh
hmoMa1mksQbwEzJDfNtU2jXTnjgfwztiV1Y91CCYHEgWOG4/GN4TT8YHMLyIN+8E
FtQsYHiWFYyNzzK85Sb2KFjOkO9i6MbWG0DQUuR1dDRKVPQX107sLNFO3yiZXvd8
xd+sScU6HbnlK4BSTxqy1+M1KsiVoPfmQ9VsoYpvvOO8WMLZwm5SQq0NPjJWyqaS
tOYlm2327gjdKPRHEzFJHRjtLlTzj6nZszZG4zBwbGjxcCb1oNRJ859ZsXQDhk56
CfUdwsxqcD2yiJNhfkHZ89EEIUTUWpYU0LbbqLe2QOqBqoEsdQ8o2IomgGzlnB32
C4QISBegIycnwS8tmJHittzl1hH8uXIaoJ2wRVTspq8Dp+QHCXrYvDRltP2pNis0
r7+GinvPO66bFx/fA5YNxUNHREKRZ77Ho7jVf1zM9ZEN72ObYmObnVi3f4Z1X9ip
yUtQ68QIFV48y0vRhpEH/JDh7Wut45D/Q1n4ShEwjDbJMeQCC12e/ZEYBX3YAbza
VEsO4eD86bhQO45iq9FzaVGQm2xnKT0qxO2UtZOVDz8snIiTJijeinl1UKxyopwQ
NaVlIGtnk4jE/uXkk0tDthnBPDcRdlDCK+LihrMCQtTwbr+75+Mva4AeHXknqCdo
KnxB948DkcIJpPOuO93rrAbTETpPyaw4dJT72odhaM+CSPeRwrVS5/h0OgNtJUcv
dURVrxqYYany1gqQihnu54Jy426PLT0D3zuSi1oRL4zCVue3S67Ot9Dd6tmYS3K6
E2HFDZCSevPk0hXJo31DQzPfMjVpLb8sHCr7YgyzKhPlmo2HzHxTgv2Ns4WSfBie
p8j/B9P85cUfSVoGXJ4/M/bx5dISqnu+xvzz4Y/zJMVBIEis4XFF8H3Xu4Hq9roR
GrA9zJml39QN72rtejWlTIGfLccMHw4p7QdYabRenc5JcVJjTnOPBKrgm1wGhIzx
MqDvyyU7AMdKYZIphXE4gd2RDccr5vFd09oGlHtOPbWCP2a0rp1oa0jsqOH9glo2
LNS9U682QOZTVpBqkcNJtTpYroFR99VvvDjo5D5AAw8YzuRvK+sGGDaglAoLfzIy
ylc8PrBF0IwI9aVHVdh/mtioKhIS/2YiMQyGmnHBnJ19wlLyzYmxFtQEZXTOA9th
7JzWdcHQQ4VtPyvGUAEKtUKbtUlFvcouVFtrYAfJVPrklSh/tL+GB+Q53mZWXNQq
xyim6C7nA5Yp4l7Cz1ZJafUr14L89zcwnOCaO4h6RxThr679utAzr5Y5xDPCC1qu
ZI5SdTOgWtifaIUsJNr7lkK1BqXe+7p5U70ZIMT4UWHd/cdMmthpF7WQZTAPiY0M
O0lsAOhJ4P1WnmF9u1PkTiDRrX/nScyhu14pv1Uj8E0CFgt3YGBkEyIf1l0JAra0
TLP+c8ANvIggStgWC9HiFlnNEOG51QZGpQfhpYhEvS6E9l1/HtTwkJRfFrcY9ly9
rhPaI/GpJJDyhGJVKC6gLz90LqXlG05OCcdoKJIqPT6R+/QubVJKzN4aVmAnfGlI
ML5udLOkpL5c+gIo4DdLM5LZVpnvMSdVv0zqu5vWZ+eK5bEEOtMvHkywOLOKP0HW
22St+Ynvl/OL8TC3TKZSpwnflHx+X2fOm6fKw33bioZTII/kl8+bW27LE64svdAq
4q3UVCPjszckYAoBuSumoKv9agjpIuQY8QL07DCw6WIzaC79sIvYiz7awKHNAoOb
0VNG1Ruge8ZaeB7To09jBYg6Rvs5+xxHHIoUvGG2dM03JQpLKyoIQe76OwZnMsOY
ZvCiJysnJxerElDKNivfaUcTf8+a/IVeullgH14JSZtZW+0aPOuXI1H9EVG3zCFl
+sAd3NX6Fm3IH1yPjMZkvQJN4pS56QslkWjMQgzILYKd4NiUvXQT/2BreKUN1yR4
qOB8XTIWxhZFlapJopkar+eXaCOY8QspqWCpNDZ6/tax8U5gdZKEArikIFSiu1V9
nlaECCUBiktEBOWSesZtQzys0Ua6yGkF8ZLYWDRqiBV2vnk0lqvJovP+0MVhw/TR
NQViQoU0Gjp0jgDkoP9U4VudNamXsZqiRyYy0uJvdhn1tYIyo1K5P4MdjzhWZ0e0
ZbuqIctnDsYspuuzMsk5NPxQGYDofD3uP8RgfNzagQgs25YJlwL0WalhehWKnl/E
e0HShD1iSHMbAsJ/pQxhaO0qM4savvDOvJeNgBmqy4y5pZdu0bzG92zaQNwiHZYV
A/x01s0X/IqYypTAzea4AgY1nYBeMDGL7Pk0Qt60N5rXlQh9s9RHFD8am54qkDfj
DZCUcYMTm0CV0sqLKBXyPPP3Mfl1+Wqx2iFOqX4ZCXl6iFaJQsPx9hCWOx3A/hn2
hRmWHwmDOgeRaZBIe9qcDBDi07++BAlJgtXUT7Uc10R+B/wlK6u6V+9Dwls/Vc0G
C75N/Cj866QcmDRnpCiwTQYdjNNIlwFBfeyHj1PlVhVHeaasowK3Oy4w6fwCXt4R
63pOz4SMX80aLu6zmPt0IGboGAJwtLQIa+u/zsDds93/QWGH94jfk1cNElJ2ZtBB
x5GHil35h31fXh2dAXsAWzmfd7C9PLPj/mYn0ArRkjjjlW7RuAbI8JGwIiaRo61v
ytvp7PxKd4MqCVH++q0vJzHRFNhirhwtERdwpGAaVNEnht4BrupGY4PEpokjlOml
pAxhDneXSbQLAnIHzs49Mxe4weJZ8U7E+HXbvu3DXna/Buwuke1lmi7i+Sa5h2fo
z8foZftJc8CQNGck3oJmsGnUGYYMBAo6gR0cxIrRzzA2E2PZoefa2g7G5mxAqsiK
DlgjF9gSRNMUxhTvrBbU5gKJVsetzbWS55Ynp0DHBJDAs0JRYVC6tsM0zIBv3gXV
qJVIStuOYW/+UYuW05g/SDOfNy1ClzbwshDGYLj5jdjReEi3QJnu/Wpy3befWerk
uY1FzZtzHjmmsPsJEcLg99HwRhLlj+nku0esX2MTwu+nu+5FhO2quUzSWSLGJiNm
2s2nU5gOOaneDpKlcNfhobSIvbsINpJYzoWcXfrZgT4kUVexDACVJs4HsY6PNIgt
Ea1OePRzUZ/f2Cn/VkiA2wUIRKs2d+pFDBd3pU9A3E9oAf2WWJ9STLnVrGvT2kTt
nEJealNcGFHz949IW1gwq0I1yLUKGV7KzYISvzW1syVXgSpba4JWoerlXpA1F3za
n8U8lXg5HQ4x8ElanU6uxLsqIcmVDUC36dh3NHhtEvqLrCVmQS7cVcWj2D0ehYjd
X6nhL+lyIARsrm90xonahLWgxQoHtH5UccZkVociC5VDhA4/KSFBLsjrgn89JIoz
9icZ8ljR8aZnHPpSEp1/ZhhvrNOAYOwxNlwp9a/FDzgCO4UmFvZkrz08RYNNfj9F
iN4hHrN66/iu5xJ5GG60aQ0AJWk/iHvWwPbrW1/80Hcie8+2SwL0vwMMWB2yw5MI
/YwM4pX2eGKFMzPKzRM9/1H8+4JX2mPjYWmJ3Z5URCB3MBD+673LJTSfxww98LnA
EypevcVkYmtr/3VWdX4+Iv2op9epq/GcB/Xd038+2G2WzqBkhjmu7GyrF2sTw/jy
piT6JJXXtLTGK2+vluNIpcJG+Y8R6HHqdSRU9q4/WLGDcDJa07RFMBFGyg1VzFrM
nyQaJ/zdeMEpNQrnOyZOuQN16DZza28DPpfDmEe92pK2iVwM1b0sSM8YkTiuYmsQ
svwiHiprIrlPQXRlGUR9lcADm2Oc15gpz+SJiD3YbeTu0k7FLTaYxhhWMYATxCmu
+PQbswEyLCoAAoYu/c6+GXA/MxkdpmVAkNXeqRJioQcU/Iyux2nVI4Rb3cuvlYYP
Y3bnL8ghOfReQKyQ3kaZabb7bkqA4YRqQA7uDFZD5liGEE9dFMFgS/lT2EhAEIq1
eliVXlWlMi9OQ4Pgeoqhh9acpYdZ/hhPxjeptuy8zvg=
`protect END_PROTECTED
