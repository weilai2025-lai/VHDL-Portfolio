`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErhhYWmJlwg8lyX68zifg7FnwnLmk7svu5ccqMvp0YtsIjZnTFN2DckLSeENfm+d
tDXFO14/VVljcJdZqD3TkeADqK/BRAuDXs/TCPSzaWPOmcso4Hy/aKqnksIuBSOC
yh7ZaCW/CCiayo/M7jQcMHwlWB2LJFrjW/heeHC9lfQpLSSAEgcIyGAUqs8qt3Z5
v5g5SdkPttY3uSojpx0TzgjXkV0mNRp1Ypyulw7oXOjU9oW/t1x9IBtPhrqdbgkS
k+DeHa1MkOAlZvLjnI91Wob0+PbhV+5Ya+9W6PmS4ZU2kWdCjw8ukkSi0y8esb41
MODC9VFa/+2FFLUuigUKEz8yZFree7wEmV1TYJ364M9S05jUbE6cMarUpcWRbuo5
51aNGVANBJq4zwtG2jRUMzCvrUBjGD616oAN4nGUbWJdMwlgwMSs3v0Fn8jGewHE
YDDPpnDe3bPTccalUpPIbwdbJWcj0t8YtlrLsi89MhFF84XFe4z0JdosKkQwa9Ot
sltOaShbuAsyqQqow3ZIZPG9/8cuIV/novrtObiriXLFGIyKoxBaVfhplsYi+apg
5UBQNejMdG63A/ObHAQG1qGLzTicSu4z7C7kR5C9gATerviNE7dc837kqUwm4c4I
nw2ScgPeXKpXtTmyqCg5w9+npFLkRcGa9I8HlsPVlbYHo6naCOvOhRbJ9PcGDLnn
KAUqy098FAbGaSnA5TnPMbzemnWIP7BQFbzG2qWY0dLbRPl3EPZh0TgZsQ4z/aoB
n92ScsePxO7pk5X+1GfrzcG52moviSvJPU3p3Al0ejTDRZOCTbW6pr1QsZCN3VCw
i5JPpREGD8v98beezFlolnz0UxSBBPqKHodjBBjdiSF09xHoYg3Ky7nfVbqImmea
vqkyE0CoBcPOXk3DvrTeWGh+Wng/JHfODnTfnFXReGLWOSuQNAObec7kSAbuGKhU
+toVyrswmPqD1W5p3o/SbkG45HtXEdAAL2aUosz/h6y7sg2lNTos3I7GbbZNGorV
lbXYT1a+WJr0Td4jwk2Y0OKYHiVVTDxdmxUPZJl263vMJ6DPt/JJhSxyZTs/kDck
kE/bE3TR0wyuCPxHbdtjLxu0pwO+f5QSWXyLdYIE39MGSuEVS7rICwT8tzJG/MYa
z7hxr/4WodRnS0txm64q01Xz4pDbuoIIRXQ8UuvnpAh4BQo8a5itPLrXIfKPpo7+
dmN+H8S131DkhBZNxpuHFS19YZP8M/kIM4PaFJNpcepBGqNZgRfgzkBFKodPbKNS
Rhxphu6We7XYOtMeNzG9PdIsaw9NNwiClvS3uuquQm5dHDAgfGn81rq/VXP1bL1j
wOuFUwbFZvVpqsfaB+dUpthp2njNnpgWER41RofVp46jDgtnxvc3Lts072Pr5AK8
2+/p1M3ssoJYCY1ixw4MGBZ2ixni2ImvwVLGHwEvksWiFknZLgtDq9LzPztqURC8
5498+EVjiwCjwrtwarJ6/Oy2gVZEPlCbXwSkT/S3PYFbaJU4vz9g/5vVIVqCqHdG
wloLMmZ8vuN/w9FHs+S/ANtKpcMW6gNsL0itkPXeEgVRh/4aBRa5XWfi2KuzLboB
R0maVQ7CS2ftnYufIP3C+DblSPYin2VQMZudgq8rvWWvGXzB9kMPZPn0mb83ImRZ
68RtpPhseA1IAeoOouJVyq0dIXEsOlW8iccDifI54RdPnDbee4SE2rQapIbybc3e
+Mrhd1zs1C0FGb7h9QSppUq7H9eiqtmN/6qpxL+W0yVrtWbhi5uFexRycAKkprhH
OzliWEb2tN6hYiagvy8R7WzX7JFgRoBGjFZNvlPZAIc+IZ2AyecO1gJbIaA2sKsw
+8ALXaz+UC9ZiBVprki6Pb0ueVtfkCd9xQYT4mzfEWutPtwzgj9GUEvpQVO/T3OK
ZW5UNK9NqbB/6VAbskpAhwe6Awr4TCFzfENHTnVL1w6q8Rq2kO7HrP5g2ZP41iiR
7ZqkNTCS0BoQndhuYanHhLsg26Ae2xxc1Pv6vo3PZFBXNeBH64mayF0kFACfyjvn
VokwRowWr1HYG3qNSl99U+jzavFAkdBBj70tcWiL/rrH3D1gUzkmUWwrfnDdaFN+
zYUBOeWGXEg//PMzXLlYDch453qXBmfdkUTt96IceEgh0foYydHpyMSpaeJPs2Cd
QClNvVaFGRphrLjBCnrSsDQUthYTvC1uvNc2thQh0NnwiuXCa59v4bkgzYTPoLGo
+zsyLn2lrtW7AEHM0S5kNlSNqpc6OIJZHXeLlVIcM+Ko2CKZ97QQHRkf2OgQxje0
lyBgYDP1cOKVkGYMwOnXQfSNLuSJ0dkbwY2N6yxpvg8NXgP9RtsPhrwy3AjP6PTL
Ssh0E8M08Eg4SVL1Qyfuk/k0q62XP7CtQff37R16u5vwtonkt01bHIYbCryyMG2Q
2IOprI+x4mC9GSm2zTjl+QKa1Z0uXonchrQyt/JSTVh6XUyHeUPCITIO9CuxxBHP
OYy9bOX5eUp/kVbNkkCL9T8KyxUsDY1SnG0h4qWH2BPybpTl09qVKupFN+XsKv1z
bPRiegLZK+ZYtSMN6ryWIy9AwAEZtjR0lKgPuxBRpQ1xEwb8WwgevG012X66+y6y
95LBTNWmsKSQ4YL3eNfR3EmT6kHN3kpFOubBIBMCQMQ+CXeaxPn0Op3F5KmNzJ6C
AneaVaDmLgPUOP63kA6wIUQQ6XqjhkrL0MuxQoYtHoQ/oitNyTKpd55/5yHVc2EC
RD479ikDdTDmoB2k0qRtSgoDMhXeKureHlkuU7iveVGW4GeOCU9vYyQFIzjpnJZ7
mxl7gBDVVHY6QTQw7f+namydyVw3eJEoYTn6iGfr+s+7qLjual54iweQhRre6JBv
yx8gs5T7qTXoJ3V5NnmUiW+1SSEkh9mMGgzIAbV10bTfkxQ7FeIKivJanr4IONYq
lBXY1Y5pNiQ0YID2Xh2A2FxLr/AeX9xDWT8Y0BhDEWAnXwp8Yoi8gJW4bUA63GoH
E4rfOQExcYmnr//JaichQG4oIYkmyU+vLM6ye7rVWep2Duc18s/MkP2m6hDZ77Bl
YF/HJ0E5Y5C3iYtuXuHSkY/hRuiB7zpgX1hBKTXpLUBu+o+M0CzYmhrqlcOA4TEG
JBxesoLlJ9z8Sh3CR0xftq2BVltsyhEEjF9ibri7x9+pl360sdcn9hR7mxifdo+G
81fuOgu/Lo1MveakFHdq85zHalytnb/H4E1GP1Gywiy5myjxs7i5DTX58BuZzu9M
xYf6d/vRtbax+Dx2hz27vrcDAAFqrc6QgU8fv47u8wbMm0wYP8N/kiWSyotkqWZE
hvLiU2BN42aTZ5BYHG3+uxAlmidS/fHY9/AmiVscY8H+IIHURIDfZ1jvv/z3U7/O
anAGNo1T++4hJNp7xv4O7YeiWrO9ipj2RErZpyHZLQJtJnZubn3tTGvkIcftfgjk
inAcZicoFG+iB/0lNuNNXhzGC7+v2sSs2NNxFKHVACSy+EPF737fHe3LHZZlR1zD
8rw7Pcp0d4IRNN1RhMM4EmtD7jm50cXMbqzcrCO8WoOA9DFYGbwwz9Vjpp0hUigg
TJBvWs9i/xB0YaSd2HfRv6H/PqlJ1K4YnMS7N603ekJr5SwC3L0oz7/5yWNXZpQb
jQOBufAP5m+wfFcbicpy8M/HoKZAVr/YEW9BPmZ6ntZswmNc2CZYVy6r6mFRODfk
Uc3686icqCdcomKZLiD+9/5hM5M/8rK9QlWpzlQdir+KnQODgB4AZQ9oLjmDDJ9N
u5vNTA4NUEpiwJf23sv6jXrrOD2IwDEzQHifV4Q1WQVswZiW1HXIUrIMk0Copxrd
KGQUBmhLDUdOWdWhFmIGGW070II/zgwSmtJ2tx3oYuDvrbSvjvofPE81/4MzfxT3
7BFjE72doIa69p9D23kiL7y/74YoWSIwWXS7MJw6shSe3DML58kDsr/v45h9mJ40
CTQ1vvCkvLf5CodW3Wf9lyGWYMIgMUeNpr61BIb6wYFnY/4fT5FrNQb8tJuNg+8d
roDHwbeADEViXjPDCKBZRz2UhVAQxP8oYx1puNd2bLpcIZpy1EssdN6TEn7dzSOy
WCSQSMfs/C7EGuyyu21M74LdD7LbsgPOfB9TKlsV5QXtSykTUPxumOv960tSIl0f
sRk+XE8txO/eJowY8rTwIhqn7tta4CvsRV+xaNQHWYyzHoF1gqsymNi+dSaTm8i2
fn/EcaYVvIZjSZoYP75zzUjodXHFN3aAv4lWOC1L1c7JI9nZ0xZZO2mqQ3uZmCu3
h3JePcNeTWlgcQBOZCFITnnYUykIe2bNqK7FOpa1yuAkQsxYGuHG8VC5GOAi0y+E
4ZuTabrB2PyYy23WlJJoMNOCCCSr5LkRnQAGUOLcQEqab11+DtNYC96KNe2B/RkD
IOGjnpvKJB6Ck82s1JOS0pXZ1uFxOsI007fTl1aA9g6nUomVgXHIZVQT5QI8pgJL
obnnd88+ohgWVe7BtSQbZ6pPrcP5nupqH0SzjHoKJCWIkdBW4H6bjDESVQh4Zhmg
ZoyY4z/O3H8qwIWMStXPvKTc8M5f+SJDKzM2x8kD1cmrOqPUHxwnFgnwQcr8Xr3+
Ntw68bGZpFY1DVKFDAOLq9Fe+LTb1qgdSE+jP5IKsub3f8b57z8BddNjYhJNWhsu
stHAgDahs09HX+Qhrv0j7+uFKt7SeJhjlchC05OrMJ5hbz8aFrjWymsDeyOEhVn0
c8x6jPNlvKlkiCCvbvnPmzDZnxfROzNpxRponly9tmrMzLHky9dUQNB3aVLFbdLR
e2S2OSu/XQB8lTYf9p3G1GuWFiComlh85ZerBKRXFSfkBqY54InAJorDvF96dyaL
WlZ5yE0sZ3JXCXIvQW+qyUl/U/QQqdEd+qMJwSl+YM+cBnOGxDOUTClVxtaqJgCx
Yeer4WcKK70pJVa2PW+EdsDKguKUEGoXwV9kE8IjDM1JayIiEQXOxLdSjP5lf7ot
nzMoPm7cvvUXd8DJX5TvGZXxKgao+8loyQZmMywWReks14vx+wjsmE7IZJQCLNxx
F/TjOyKOZfGk2jcVQM7jUEHltofwauDdTABpUe7xuVtWs1aamO3NIRm8bOCsipuT
iTzcdrZ/n9Yk9fn6dlfEQNt/i8i+TuN7UteXosVwVwvwfzsHYhz/TqhWmAvqgR5e
YWRhKw2Gwrtz/xt8qU4ZjiLc07BmRthF74oMjhXP/PWrKAPZUWJZwAToCPi2vBhn
yzbHEc13rPzu9r8AYTslZueKzLQoySHCJZADYEqgidGldLJ0AHUdrd04qrlpPU2o
CjZ7Nd2iD5kM3/7KOWk0jWMmgaVvjOGzKhmeTIHbN4wS4Bg1Pp7zjiBqcXsZp9eS
X+toOCQLKIhPGeVKbk6AcgCmuRmPx1kPnRBh/3LqKAD/YkXX6OGTE1cq22XGopdo
ofP5guAriny1II7wDM2WvkPZiUc1K2KL/7o16Zk7M9ZKXGXmRvkouvO0fqi8gkMQ
MNNJsb9WmO4DlMG+WsIq4QA1qKPU+YrmwPaiHQJmC/aGswA8TgZC0gtkBD1s+OYU
u1i1pbepJdYNDoxgGxfptk8F4+DkwZSL+wX+NlL0uhu4q/W1bmOJqZ0WO0JJ7cPC
LEFdZpLkwyoid/Vcy6eH2EzlmQLdyGKOqVumEiRy8O96qfyj/XpOsv2ZYrSRkl/G
sInDjFSxAP0m3qhFL+sIgG+PR4hJaTtxMkSoJ6/UaH97W0jgEcy08rOxuJhnDu6e
PfAnBxFnRpwqZ7NTv9EhwURWShiy9Bgh8I/zRfj2bjugw1In8G1qTyXQnVdrlfWm
SpdqMLK3p+bYkKuhNLpWDpp1zkVL4kkT9h1RfM1unDJ/bXv5D7pFooYbeKA2WJ4Q
1lzU3ybNFFvnFinWnK57Wg2X4FPrAIdPtbfh1nEsSNdpf5YDsdQ14hv23m764l2R
Ruegy4D4B2ELatBAvx3aUVnJvTOY2sDkOX25KXC5cH24UH707J4zPSaWd74ZrVr5
UNccQjambKKh1jCrkIMHCP11ecjhF2tYQDVeLRn+0h59Q0b8pzn2O0uCm/ZM61Vc
apw3e4CmRBBq+z4qw8ohD3CLRXdtCpMVMChq5P/MFobkTCsP8aSp5Xw1SZENqhnp
4ocuS7gkvGtlTS8Xkxq1Fwi1mGx7KnJt05C35WJ/TO8sHetHWtqU3yQdR805G/YW
DWF8W95j1bO1FEJ9bZo9/fzGQSbRv0sKKrWO9bbO2BmMTQpinovJwmtLwgwSyKPk
n1lRHNNWDy+z58gYHgoclpUmmcogzfR6Ld85dd/auCTRPvPohEJ7V4NdNDbtq78V
dROdGS0hIms3oZtRDDQpXGY46jbfZajFmcucgK7XAX/t6PDlDrb7J/f0eDnXS5YV
QSaiSR/eAwXFNXZrgHUEwIpdJnyovtHMi81P7j19sqwo4eFtldZtm6J+FZ4R1dHl
0NnF4kJHqwPkmXCAmEEOdN27YqXiU8mI8j8LDtBzcZYlyoJE9oS9s9a4/CgO11zW
G5pTDPMaO2l4SaL/VjFZ7I93KMD6f7weYVhb5BzxhnQ0dtX+OFdo+qcQeaR9a/mP
pClNthJD4VVaez80Yb8a1hM9Trh38ABBJeoiLNoHshgWTSVe+VLlxDr7/GVScsLX
ydimpXn3oKpmB4nNaE5Ttv9C8IALYUcwoEkLRuiRwXMayQeazhE3DQyDwMO92cMl
GkMgv/mUmyg7DO2Kwe81r08kNpUxRZ8RLBeHypcZXgk28s9wNofq3DqkyCumC/Y2
hY/lDdLmUscg6SFZqZxEELQ2yQVge/Kc26HVxxnhi32sHdV7s6a8y58YmpDTGOaS
yfFPwZIMWs0oJxyxoM0OmuNnJ76yrKq2Sw7XCoShOdQYzC/p0hwKxBOGHOOxVHHh
KP5qeKd78qIvQ4x6Ma7/Gg80d2COQwiiYyh8nqiXAbBgYG9Oa3jEdMLBqHiVBXmm
DvxHFLG3mBIxdsp1aDEYub5SjkxFlsgv/64BaaQmilIofujvN/8SEgpy6rh1AZPs
ysEMAwBIimcR8mA1iFdQrnRxjvTLT5ABnnk+WyXSrfu400hS0nQh2jcn8OVZRc1j
Rylx+pPxxAAoozWwnWywQXFgCWutIBKWM8OgdqeemYZwJpLnizb67Z+pmfJ4isZe
wtIOPz6Brc/lb6dRdfF8NJoWBBNB9f1bjy7r+VhCToZEc2qNpMPduRzf06uRHsA7
PqQMFCN4PUCeyXYNveQngVq8aucL6GJpkLlPPyAUVrfDeqdP0nOfz0ai1F1EvhY4
KwLYOYAIrxsoA/58lRFILme8CvrEpmk2GX4RS2q0/Nu/eEqGasRJDFZfPx+9TwoM
/W82OgCyU2CcpFJJWzimgfoa+d0EOLQLhmjIBQKaWJpoJYXGzxtOE0Y32nAG9Rjt
CPMlrpT/aMWVcxZcaSg44hRG6hW3cAlQhhU6piC58/AHVlmEL/RHsOIEeoBxNK7m
JeVEPyafJ28nCqfMb1hWzL3iCNKojf0cDgZhSO/mv/ksvHQlKegtCnQOQMxtDz/W
AvDT7QIpDpEvz0eZnGe5v4yFxDjwWmdSRRZCh4IqDwiOYmaZdPCYF+YksI5kjetz
pNAyR0N/o2JU2hP/+KQ35bZ10irtIgQYFjEmAn9z1TgNBjhECfepN2Q/fPm+RJ2Y
ux+N8hFpqe54xOdKtJamva+mnN6JFAm49KINSgapN4KnrEEDv+lOApVCpmI+DE2D
CbfpFs1OxXBwFySrhJgZE0ofBU0FQYOpERVGXLL47zU3XzgUL/Hc+mV1CXHyXXDr
lURg05M+kGu34aK19DrNoUXrTe3XBbrZj6fEGEBMzbrtcmkoTMwX+YBiGAdBI1nQ
wJyIpIWhqUtrQ7GSO1l7MFxIQlb6a9ej92LWeFMiMzOBKea/zhWcpjt72P06EJw5
9ubvMVVnDvKmsiXd16hfUTvBQRfbpEcjCR3hbz6Dtn8R/ugjC9IH/Rb5c075Dqs5
44sEp3OJHeGVelE/WXCJ2Rp7ZYsXh4JiDDJz8xG+m3ysiW6HuxM1u3L3ZgiYnABO
GAMpiIWRPLSJeD2THsVGDQk50V+ajhH2ztCwS0tR2RAuSS/blF5th16n53O6ZVqg
zvqhfhocaGAWIJkzlMyWBm95pyU1VXz/87U4rTA83N/FgAtHsmSIKBiufcjcnbQ3
svh+/6FPq+2AH6dNNDRsPdVHDg9XeKn9NwgouxgZfGLSBsYElx+QjommPyKGy3SE
Uuu3vtN4AmOdPaaSyuUzUbamOy2835B+MYiFaP3ZcE/sGcmoBgs+aAGgNxxw6PU2
bApHDUIJ5Y1kcpEaIAsbEEBS/SNG1uaJGbH8JrARiLayBsgbffyyXsVgP7Di7LuU
gX+2nrsV+Dt6EjmM/LLWZOLwwYPSf1uU9TvtmKhL9NPEEHIsee5vpQxMinfXvh0+
MRkcmLkql3p3oFqXOIxxN94Mj0L0//4IhOZOiZfwVJBJQhRF0ah192X2wYR0e1Cg
ZspDlrpiQkAvA5QwUyOdvmZAp/7uUyHtz20tGCFElqJOHV+b8WUMYYNwgNbdZO/h
lOBdV5tYjn0zS6BEY0wLElMdXvvVXGrkJX6QOQ9sLtFo97Y3rG4Lquz2/B4nslgS
NyEch7In3hHm7YEH98d+bAA+khgvbc2OLKwhez4G9xaOMmANM01UMXPA//1Q1boo
o15L+f42sLKvMpUswuwTKx5l5MbL3apY73oPxfkxn2QaOyEf3iLiclW9fD+yRLiS
1yFN5FFm/7rDllfC6kGjyewALhWwM2/c4iOSKf/rOLunXLKbVdeXaYPbpuw50xTD
nQfsgwyVfBVzatvUfiR4d3QNm/uLKAQYXA2dzOy7wtzZvbPILrFWy7LkuR+vgaTM
CLZpU4KGMZcTu7h/f9OzcFUDFoP8uioCe80qe+jZB8KninoIjK0BT12ZGFN+8vRr
8rg1LZf6OgfYN3jZg2XxjXwvlkVZbxlfLkShEqVyMllVf3St261zhC40NnFZzbhF
/Y1YASR4Yshh47adUFKeX69KCS6r36KpW/eQE3SUjDYVL9xM8HyTqkv2bwv2g+aQ
CztCQVGytidpPx+m2beTeEJphDn5FoH8J2ZLeie+eypb5tBwtf/OLXYhRTJNCyx3
D9LWOEyAdgdhHmBpAXKp45Wc97aTV0W1gjeGJbKAVuHecxIy7rGKncnoG+Jjswxy
lu4bN1YIowhlMKZ620s4frGcjyK3AcPuJX+YgAdgN4P/XDknmea/gvy7jDEUHWEr
xvvUrgEAruBVX8yhhCsTF9GUY+Jw/wabGsDWJiDTLkDgFR3epz4DSQfnYim943s3
qTYxYPREalv3lkTkXLloDQM2ZbkBtXKSFnIOqivFocv/A5B3Z+oig/pHYWkaHfUC
tMmXYXFa/wwxCT6MiFlRG40EPuoOeJfgVPuThkvqnTbbbopn33FH/thTb+vXm5Oa
RcghSQKCFUHP5Mwi+wXGrA==
`protect END_PROTECTED
