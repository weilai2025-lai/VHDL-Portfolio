`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N3EndyIVniN1tY2cy1xdY2RV4JCRdQRsTf1CAijdBolpzlOF2qB9X3pjcoo703RE
5v+xbC+rw1xvEGhFpkYu5Lct+pyJgQkGPxnzFItU+NL5NDjhiVN3F+fc/Eb6uWMU
mFHg6XQKN9se6biWBxjA/hYui6pDShyIQBNlU9AvxmPquaoMlJ8l5zhxbXsRHntv
20nvLnoQWoBWZ4JMu0yn2d7NLcWuMgbM7nagUSsTp906l+3k0utCPu9yvXH5zvk1
xYBYT02Ih42alH2DUkFCGD/pgUkkl3M/AxKAad5h4E4bIWDB9JtLtuueEbe09w5w
m0MPP10m38B93a9vSRCg1NVrZaKlsO/QvMKmAWtSrhaDGfmrq98ahxRyEE00fHHK
VC4L1yVYk5wcaqwwvyX5im20KiW0/CLryYGzcGUoq19P7ppLXF4MRkbtncqaDFMn
NoLvvlvT4rtcs71XrlqobewFSInIS0DrEfjtsv8KmLRA+Hbq9cIYDdkBQlMRa7Pn
3z2w53+zJG50c+DqW9eYTA==
`protect END_PROTECTED
