`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kroMQFvi6vcodaAA+sC3socghjWP2c1eloFCuWV/EUb/ptdLffGmJROzcYM3F8IG
/DM25YeTQDQMzgZrdZHy66efM/lR7IDzsp5PpbKpIXbj9AQaR4y1mX3n16WgSJAp
0e1Zh7Yr3RC/gMKhTBe1Y9Ciqe9URBkZc7SnddXUQ4RDO6BfVw8of3tTE/ydXznI
OZzJkxgeEdrWACZBGgk6qigVzJhK5AwD4fLiBdHS9MUhl87T0l9P2ISfwWnxdyU4
aFlFZkCYcMdX/po/Fp5sASw9NnC6ebzdk0UFrfGLJi51M98RJxIKgIiqPm7R8RZr
zMginN5QK5kyjYPMWYuTd3xi1kFCfOvTISjB1wSKk4chx4+VbFj3SPywLHmGr5QQ
5jtVTd8Z/k9+9N/7RN+LlQg8Nw/libRCJ+2Av8EF4BVC/k6/vqRAwMkxVK0Kvr9g
rIt29SZ1dHjuqNhyYK88mqiRTGOkVFqVXIB1V+rLOfX2nGI3UfZDjUA5rkm/81Kf
u7xIsF02ujTqulUZJ7Ks5QEEEQO+w2wLXu2QaVrhwFMYi2Y5wkrOODV3Nhg+oCZU
ww2YU4lmzqNZ29ZVcDmEKB76EhHoEqFiJolZQ9O9ycqqEv9aQj+61BMh9g4zlDij
m1y0RR3apRmM5roocQYO1zgSbkFPHsouZ7Fhqype5AP/l8ieStzXvzfvLDAR54KP
m860fmIpiBvTtle6WIKjpIyQi2Ye2FOq0Dg79GKLxoLS85ULhVVEE3Xw/cDjkTdu
J6C08cWoLV/evLsNnREFi94H7JOBOf93J3PvQv+09ZjIxp8FYzYIsmk+HwDKhGgb
qry88Gez1E7fKADlXBpF08Bz4A1nQ7WipMnrD2nFSkRNRs91PHdAA7cVCZhq5uUV
CJegyQMZHTQy9aR71OzOQqXc/OJthwBI6BCOs9qEWiOqusRpq92YX8JmOLyy0uW2
3ib2lmWytto5satqRxvGvMVIFgJXnQGW3ES7v9MrGoxQj7fDoz85lPpJarXpe0jb
hT9BQV8K+AbWuI7ST1et+iJMCViE4wMTqPbL4sVpx91PQzCgUnZOX+d1sBD8OYqK
+Rb4CdqAZQxU1x2r609+qicg6Y2QxQlLi5peilg8chnyrqu8soxz6ql0WBGCAsbj
bUopY/Dj2edpd22IaTROlCpdkyK4g2JLgNY1edN7QD1/aKzQc+1LZrkcE3Wso38r
NVMfZMedXgwpGLvXgyDcVpgOJZhvc+oOQ4Ac3EOud1ASvOLqfIzffpLi4rTgrD5f
Wzo3l8LuwzN4curktelLmSb0V7VRXaGQptUNeFkQkHwFP7vUEx+jdj4rWIxXMMLu
spxxy6vjT6JcPEpa4MjWgGfyRxBkXl/aJFsDDqitxXDFPBKfVNkz3UcSgt3ahY/L
iB5i/tUtvbytDutMnJueoOQnHiRXabJBZ/68vDRc5g+IvTk9ubZPilazfXuQGEvz
X/yjryqLP3WZUBjdAkJmvttFD3amj4uaz61QQi0p/QMruQybGGHwmraFKSCViyAV
d38P8q1oSZckgBYuJR7T1gkV98fpACH1V2E/fQpZA+HCwto6DSgEOVEc1Mv6yjkb
fNsd/SVoib2YNdUwjJkU/TqV6lU+U6oVBL9aQym10Ld1toUlebYi3LdOd5wFhVmp
ZJms+147+F70qo8bsbYcLE6H+rBpxg45bXk989s6RyL7Q5Y7n6TuMfTeD4MwEY+Z
ZS4sViDHtlOHprwx+rknj76wnc50Cmv2naWoOkKIvaOAiBdZfPtlkOoExcK8HWK+
`protect END_PROTECTED
