`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+334YU4/7cYsl5JkfjMvT96t39CK8rQ4FYhbyn5QzmdE/MZa1bvUoHDiaSMO/wCt
aab7h1GUGHRVkxw+AKwfRQiwUtDZX6iE+T8QD/J33826+EC71eph4EjNgoLOaRwB
BguwEO/DtNSbgsNiYJ2pZV8XwVSqIxC0aJ7dlL1YbTdoxdmXV4KcnJROIQBLv4bR
CGEnVXvShlRLYLOvtKFCBaVjUhaeUd4MB3FDiJhMwqc2ORCiL5IFKSXa7QSkZweO
psFNXJPe9t9RxzkG5ebtPlK4aOlT5rC10ogKXLl8ZUw30ELR8nq7FDX9+xuOPX5l
WJ/xkNK2IKWYDohoaHpXbA1CQ8Tf9KMcO8EL+/4fisuykDHRN9AfWtQ94gQJSWad
djuZx+FEYQaoCGyGEDYA4HX28mKDJet0/7m5qiaB5400oDMCpmsiDw2AbgebmQ70
jmmoV5DahNw9kXh/mIEdzfAE8yVxCMD9YHgPgHbNDGOLYL8wBN8ttc2zGAw54J9D
50sPl/+5uoTUnjqX4ttOh/VWIJ3yKRuWTDbu48cymbEU+y+zFR7LuWO2emnmg4TI
kYlJGJHL176yZyIXHFg2RWmyM2jJGptdoUwEUwBIHMkZacnd/lLq4JCeKZVgQbvn
X9shqu8OHUHA8vR72wGUf5DVNwnJMPwXLh8NzmILKu4VL/IYhgdDgzjtXYjrmiEk
N7Fk0P6J52PpZCBPDVrCkD0A/uuA30j6xE5R216gaGHGhD+aWbhbRA7DyXCJV1IA
TABUut2pFtDBc2Xv598hTNlWxoTx6fuk7ixG0XXPUv6kLvIVtbRYrIZz3MZjWEWF
bVCxIgXyqq7aJgj6a8SyGO7iN0U6eFqK1ZFSP533TIGiPFlnBei3kyuCeavOUB6V
aXDnoAcGRJV53xL1j5DgnlSL8Z9uqwJaKBMfycusEe12Tn1i5qrro+ubgqXy5E8h
cORBn2Be/sgxRO/kderazW5KGxGxz3ryhKf3WRQklwvg+hJb02GFCTWqYOn1Bzsh
RBn/ZI2MZ9CdddDCVugWTx/fOv42XkpmmhB9JsmGiY1JIHpjdpbqTGvSOdfDv+ab
DSvzw1bHrK2B5UiSgrone75TaT2VBj1waVQDdm8ezJAheXLj2lZqvZkFJ6VafP+8
PHWTP3T6IdqysmF0e6/ENXaugXmHRWCC9X7oLerGfAKGCaZpwO/AMzA09S6TLSPi
0VjR+H6+Xi591rFbrYgqTTxxaVeRKhmKN6bfEW5/Vl7RnhMj7ekjzCmFDoM+fNKn
Aqk6x2ObJmU5butfviUEtJSmX80EYUC1F8POTifgGCmBOf/nG9TFgRBf4tAvF4iw
U9gmXgls2TKwYIJELu2c/clbXxjYBAMNmJF96cdOzbw2oDkUY6X4ofVJDoTZnVr1
CyuGMgEt3SrXFmQxhdl+nbc6+an8I5MedcJeWo2zorkx2HqzRZYzLkchnRlsWs0k
zTP6+dKskfjeoDfFBoKRC62Mo3jt7Er3l0JCiKtVJwxQTpkPuZHBj404d3T7voTI
+TfmQurvLY6+An6NgZj+x4ILBFVcaVaObUNyl8xqQQb+f50mQt2LlyBGDV7jeOTN
cQTtReN9G/iOW/+3mrs8MBeCDwSTznZvmM8aLPMiIWaXy/ljV5/4G5HNFnl0fzLN
`protect END_PROTECTED
