`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UqjOn7pqrig4/4DMfKnCfaNRHOjG8J/LxV/XJm/PjOot5H+gKyeVkJSPYKwmTCB0
8mCerEGLb9UBKSp6NsSoq3oAULdVV19OHdN0iusA/Ple4//KsHtwuPXSLhjVJhPo
zThzcU2sj2OGsc8rKBPt/fwS3Nis0khEHchOyquhEz4UHdjBzVzfMZmVuDvhyewV
i96aPVQdDyri5oGf1SC+j2jALi8bhxBBSBnKwnlW7E00es/gx3cSsCxrbUbPYtqL
V+n3wCoLdKdDDyWv0rlb1CZKpe4FoOOaDAuash7gbbHVFvZNTHFQv2oS/zx0JD7t
qpRhBbIB7Rah3IWJ714RCA2vpdk7uST8x2HWpkYlnPSB5uCdHsdcISzoC0WLnm2x
ilFizK+f1k4jGLvfJFrzKMTCtHkFRzwXKk0M+v95Q9IVeEhWPfWyhHnwqmNu8jXX
szUtGYTHVluQ4vsnQXezLy2/hrGgG2dxz+S0h6kcioVaDK2OaqAn4bhaagaeghEs
TbrYbfXZeZR29C+B0U9eZwiIH1c0p0cW9zMbYpRagN8HZmOkZ1r4lt7tgN9065zn
VHYAInpvRXEnMgh92GOWXdIuXvFyQsWpAT1wcwUPa3Rrx5sCmbD6C1Sk+kyF4CvH
fBgEGkS4S2LQ7NT5rQAm2dkfyaOURWEc5EurN7BLFtnlJ0SLdjlD+41v3yfE21wk
1kTAnerbH7oV0Zw3h2+6LiQplHydwvYKHlTSUMBJ1qb7znK/cn0wcrFfC8szzICY
osUJxPYiaADuqTcvu42igVJJsnNcZX+np26mNuJRnDS6sko+J/UgHCUAtK5ZOQAk
eyA5eoRLD1irjj7373WnnQ/vmK8j8AuSLvzM7IPtFehAEr91MCNAeuK+18Y65Pma
RS9I5nTMuEOCl0tVipylJ7DwUSaW8yF1D8rGXC9eJxgkeATuFPAI7LL5jQsFV9IL
/P6Yaq1KIyR7CSpiQkfrKeiW08VOO9/EZupdhDAjcotT+rzDU9HYf7x3ZBtXfg5g
d585EHxiSzXaGBDplTiG1IeQuq34RLzRXt6oS8kf/JvkRPAIFoqJ/V7YN2v7LGdw
FHM+rQIlkSSPNMqYokugcOaAOqtLjQvtPf0+6LtZe5XnVBtXconetwltebWRosaZ
Ylyqnkibz/EwQgoOzEhPtay201oQFPa3QaqOIC9RRUkoemrLtWsjg6eSVIOciRo+
9HM8LJ8aWygWdhobJQs9tf+n/u677jvVrWnnc/s1qj9UAlZqXLLCY98d/LHuPwsu
dGVsmjcPvhkvqikC93466UhNro3Kp7I5NpaATTprJRu91CQbv3EYajJEjYK+nzLp
b5ySqmwDLxvDmsb/dxrJKEcLBsQHlZffi0RInFN5KMfOPVLK1vCFRrUmWY2+av4Q
H6PGCFqw5q35sDgMYZ4KqAPMPy62o8c/DHjKT+Ci2wNJQLn2sRv9LaVOtc9UjD9v
MWZs5m+emuKIVekhIwWXOiUAAJYSIp2BMy59Fd3XWxHFdobxOste1sARDWS7d1Wf
WqPOygpzmGGSZXcIgyPXqhpXe/5Jg1TdvlRpLK+FFfuBGdtHObZ7pOZyAldwjJjp
FBKRHDs9Pi16p4Qe7GpoiQ3BKtWDPm4BVkKfMdasG1Y5wNojb7Oo/u9TctV1mfCw
zhUFK87nXXK7Q5RytjiqxcYkHsT3+iflcAJZjs0pZQbEAkluzQ//s2tzj6baBO4U
QkY8ZwLkdWHKV0nzUQg8X1P+V+eJOAeTvJd8NC7xk80LYVQaehRrTV7H5mpaRmdL
YZHndcQpLEt+1obaRLN+BVnVX7b+atnXAIopJcQW5OARafs0bocmM3gyIzA6VdKx
zDV1+Lo2OPTeWZYJKkbXj/bHmRublHyVu5kFINLI2D68yP29F7VBYvMti3SxI7g0
ia3RqKUK6JPjoQDDEyDL/DEhDS0vwbPfxVPJhnmaEwBIwmJTum3z4pMyy/2dtq34
qRbFycYE0Nw3OeMVX93vqhsUMHxfGFdleRgsVKpxcEpaFYbyjDK4l62jMHv4Z99I
b7MVbBP18fywAdWFw+YnYNrt7H0AyPUTQ59oCmFX9l6IF+r39P8i663W6MRD6gjG
c5AjL2SmJI7S6lZF+t+Pkx2C1GRAZbcigJDnoxXDmtvIDWJTwDEAbMvMpLlDvF8J
c1C32/YabnalXF/NKgHDEu6UVRK307bXuBbXCjy0nXieBsTB2SOA//fpkca/4NqD
6ZYkNNfVYZ/2HjgJpl5YBozSf5D+aOYVL3Pv7Ez0phj0BF/8rFROSfd1UR3n3xtF
5fEmg5q6TkgVDICqZnRXIjHm1o4Zdch2ICcGUurEeDCSuMN/c9v+muuhoS3sojiv
jPOgS0cdrmpTiBPCAto6G2Q+cAXc9XzLiSFog/KKA30Oe0bOeHt0keNjxctNIX/2
O0vJJFuE4BtinUWidPNynLh3H4Mp0mHaTQ3mm9KBjyBVptx2f67ef5/5RTI4QWq4
YV2VVlmUQWRuB2BLw69touBG4ppcA4tqMn0s7qVhmkxQ94rub1N4uqJyMo8oq6Ml
+s5ZWKheswJR2BziT9bUS9jhAVSnnqYMK7AKg734l2rWXqD11qN1LBN33kF3TelL
DfQEq5CSVhoRboO6PGZmuex7EUuh5tSx+4aRxNDnTbNY5YBsAJooZilpuguMB4H5
sz0hEMOLY+qLEJQKpx6ooygSNUWX2Lq3CRLeoWK1IlXT15zLyE0luMG7CESlna54
AV2yVeFEVIz0a+gSXgJExUSauxAaP657OhTp2Xd7skK5QhobeRIYo4SqxM8mIF7t
9zxHgYWJ9balG+if3FNHY3kfNTLJfhTfsWjSaCWs60f3z1GHU+uoYT/BEIhXdTU8
pyGO+/+bVRvrCI8s0ckMZHvG2Cs4ioB4McmhKu/tnOdLHrEbsdOljyduEgS6pbqL
J/UhJICt92tlYWCtPXeHN1/1e5fpAoFaB/IpS25nKgSxrE/Sej5L6DQ3VWJHeScs
dT8yMFYYzBluyDihoGP7BJtxYiK0X6Ri5tS+45ndvYZJLW4ZcjDo/+iFzRjHNBlp
D3ArahJ4x0R/53CpYHbvXjTiWK/E5VmSTGhmE/fFf/Mj6483mFAgHj2HdDjdWlBv
7RixgVdLO5HUpeetARaEf1ofcwtKsJmVZbkY9dPKYYAqS7VgJdh5hodXlUDYMxkZ
ChYl59a+UAL5auDu6xVHjuZRQpcsQ13rbNQGE4y8BBDKFCxYWyK59DRi9mmL/CgP
0nuPsIrR86gXhK+lPDciUZWsAx1zLj1D4NQedCsX7QQWrihl5JeNTmPQv3+ontOX
u1i+PmaEqLS3/94yA4wx0e5BKVW3S0ohJtk8b+5LDBhcU9Q8BcnIXp0jsfWlrdLL
c99FRpOifooWxF1LTK9+Kd1U4vI5hroNmrxB+AGbXGS4rxOlntyWULBk9kGGjs0+
KPVQ144j038dJbXxuHGXAiXNnmuP/jfeoI50LD01ei7QIjLivoouz3nH6s1xZL1w
`protect END_PROTECTED
