`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28SIN9VeiZ7g7tFkluoiAvd2/3ABe0WWgH0f3NNPWy5uMiKV3OHUZTy/S2/Btvh0
sYgyvqahGBZsGdcn6QKLJDFLn8bqtBh71hk1kExzQYp8KkMn3jOt6QWeMFSU2oOU
OwghVm4n1bpZPqsPzQIyl3uJkyPz/YoxGiwJhuJtvBrB/dCSnlXo3c1vDzkKQ1kw
UrpsMOvgk62TZqbvHWvqN6+aBNKYCyW6p1mlRAD/Ovzte7X/X/8HYyaF+/MFYG90
QcvTLgBTFrgaBSUH6v+nRVqmT3QiTmBTjGpCLGshFaZupNLydiMd74Cf4fOeu61s
XQIROkObIJinZ/vIUmlmfzLExWAZXyrLaXzJv9trx+979b7NyeD4k6G0joY0PmRD
F1ghyOp/BrvNgW/p/qG7yK5GoOKgXWGOGT2NVpt7Pq4J5Dz9j/mCqZ9UugQ5yGH1
rUa8IAbc3QWNUW1zuIuWTrvdwHzFcn6cIayhCEZqAjrpkvjLzJQzBgO/WX6RuIUH
Qm0xLvJyP1UCGWeNZeqaqXTYCzHmDiZc59i5oJEK06B8FAWXwRBvpz26BACobcRx
doJrC8mtDY3Zim2qdy90dx5U8j3ov/M+jzxpj3jWiIxWuGGJSGu8xNI4hCzusxXH
paDxLBMSZczfFPRxBgViMXEWbBKSpnGCcYqSyiQ3u5fTnoHaMESHL3kkZraeu1c0
cPsFl7f/qQaozfpfULHZgVPT+1tTfzJ2mZiPyhhyCIHnI/rGvTUT+aOzYHb4FkvS
N3gek5ENgdZm/DisoixkBWZ9wktqcuhovyyeQxyzQDAsXpnuoid+6RKxKjddkHl9
5qPEOAeBDHpQ5LQgPWEJZ/dtsGQxxOmtJ9QD2yFqXWfKBarR0Uw56QWskUCi81nt
mPwJnp43Md+zch5SbleaDe/TEIMRiz66UW5gcX7spLaA5nI2hov5a8xGkksxkIhc
n4yY7Om0kl528VhCEzjQak7vBFBQyNlvSH8qwA1Q+7V5G/DyF2mlBFP3mTi9tSx4
z/zY90XjG+mf67nNE1JlOSV1qsyAlqunVZIpcjLcPilhK42wXfvlKXdBfEEQe1Q7
eTC4nDsxafz0oJ1+y+qiRYqXxyJQ+EOK8KyMEoxRC92Ey4K5ChW3QTc0g/fneVFo
VqY7olxWT97S8Zg9+h+yYrbtJBhxGwdc1t9/xR3A5p9IcuJ6HMOza+z+JkhhuieJ
TfOWVI9CdNR81u8RTBacWOs3cAqNxm8olNfyk2cdjJvyq4hxOxgOOmYNPZzoqakp
ChUzLZ22tm0Z0lmVJ+1nB+AcSrO/dHSpllC7JCzWyYReImoG9GiT58DtR+V3LnAa
V3b8T/qRjsrDQkjWTfa1ZMhm/D/lNe2RBnxpNtW1citz3cBagUuxvT5rj3+wsp+G
OLgbOetBQKitYu9OlB5yYqTAFN1AHenTV0hjVYnXOdlWkWtFy1+dPhyQe1D2MZ/X
fjGBXpukXaahH8wfjKfpAUZYL80Wwp5XHHfVkRNHJckpFBaCZ34tI3Z1Fjer7BwM
xicznxVXKHrQ2WsxCxlnuWnkIC4C7hRfJBOlZEINh917y6fC4MAeru69LwkprEQd
U1Gh0VXjDJi1DlGzBpTBCtLgxyOhEk1EfwYzG0UWclR2ID/GMc8hXQv4ur+qUulY
1nLtuoFwZ0sZnLmdmfGip3f6bDLhmSIB9Q3mzFkEOSAyAjDWZ6kXSIR437ZU/r3H
7gN8aTFHj5XvTWPJtfadaNn/R2DOfjC7HQ+9UAkvbCUQ2HiWKHs27q7TwJN8e5ym
DuLGyfVFLVFRSI4GYnwSzQoAQBPHJgnFogNyJwvZPR6IBEl28Nh9ejXX4DT5nVTQ
g1SlfCbMm6600PQMKtIyAYUTXKq0AKqfYD7tYTGoH/BltctUoekZR2e/rm6E0c1f
UzC0ecjphCDixEst3yZyYYpjOHAcdh6Pi0QVzbw9zYniqH237GjtetDI1dzFSvGC
l4dQqRf4pgf4tu/dnSm/uYtRmW0x5mESyO7lVDZjRpFrSQMrOPwVCm5TETg4avPW
2WO8oMZm2SYK2QvOaTrCvXdunIYwyz42ajQ5WEFoRmbHK5bDz4Vd30Ic27Qbq2dm
sZa4y2lyq1sZDdCx17uuKQDzMWQTbO2lEgkPpiowTj3zqYcQt+QUzMB8RrCNdnqO
UzFalNGS3AQ6QnL8M4grYfbHxhcQJ/6Z/qcoCjt55//oUlP4hi4C6UW5RSref4G4
2/dQhuBLcqQUxYUjo6ihGDUOx5m40IK8UBKV32reg8UwnB3ebpPQnJJzMwJdqFYK
TyOt5umAKdQOliw5LC6P9EV0bQuNzs3SL2YXC6dcCIzpYQEaeHOPjavNjYgxugOA
IFF8d5UAoW0X8mmtWvAbPhnxPez0VcUIXNvWDg87D8ZoThTkEDisprw2PgQ4OKTB
jfUb2lDgIpE7/+86RT0/LI0dNkuBYILMPbGv/yZ9tOC5VSeqHaFhoBN3VYlDrNxk
WO4FauwpuMhGLdQfQMNkz/oZv2nb9rkTspTS9EnrX624BmMLIZ1Kmk1PEeUN7vzD
D3FsMokg4JGdnK2LFqk/+VkO0Cww6AV3BVCrY0kx419DK8NSrUohDcnZN3qMyiah
BbUXUNfyo69uCgrP1/LhiGt1tghTOnDZUbvJGm4Gf+A9psZFFyBg2xhMy74O0A7a
5gs97PqkB87Ff8HwgqQyTloh69Hdu6pFGniyOlMY1ONhrgTuuHqHm/m2NMKuMC7l
sXJwI1wu6clqYVrBfNHBjrfmEdmFpw+bfGe+hn2mc59PCCcNaHqiJBTeOrx3xenY
Un6F+99G/QPghVUEsyrElhF3S8fAySY4mVDduEjzhbL2THCflxn0atfwkeIHOs1+
2U4jjkyG2IX6R8osa0tRlcxLiejuiouo5sKvJVhHcBVB9StbEp85AwREX294J6/W
in3KuvUeJV0S9oGqf1OTRk1uh9u350vKq43FM/nHH9oUSbvmgjxWMf1Mqo9JNgDK
ZNrTkFzIjZqSsKJG4vaQbWsRU+THYaKWAZYfq9FKrlYsr/zBiCeTzX+bOvGi3umS
KlqelrYT0lt04bCFMlPg167LnxFcZH31AgvyRg7S9FIPt0pah5Oi9k2U0EGluUui
dGUBYFQT4bnIVtTjO6AoOTYF2qgULVmMhCxFePPMmkCmKFlGnNnuYtumhZKwi+eX
wyX+2BXxkQgAZQmxYIaOxBEOXOe0MUItYEk1u2PHvKt9mjhOSfiWncdENG9gGGTD
P2roUVlh6Aogl+sWetIGmX58HBxr1nxur5XRE0zGtik7x6W6SMAbZr5AHXpXG/qm
MZAiW5lZaZ9AImwqdx1f27ef56LYneEOqv4f57Ck29cnQoNeBq2NJu3ueI9HakiC
7EdbCn+TmuBT2JiSapzfV4mznyp1kr4MZgGDWVmHZK8poXE/wiLNGUuinmMLjfzv
DUkc2OvR1jMmucgXym6vGK+CzdsRC9/zVAk1YsjoGGRUJgpMmyRSI4YOqgJNqoBX
YXyJLWeXT9Px4sRCh+R+NwYRNT6qUW+aeV3Ua/MB2bJKu5ngoTkYe3U1jDyZUASA
/1nlcRXlkIXgjO+khSTGyaLfHMjGl40G5xjv4JvJPollHlyi04BpizjYx2EdK9TK
iO/R/5ZPWVmFjmrah6HK8KPq5VngASIxjvjcnNlsGcggxYFbvSkEzcAXYT5ByX+C
VeWxRbXdUxyDMI0VtpTclw==
`protect END_PROTECTED
