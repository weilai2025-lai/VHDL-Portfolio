`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ru+Uy1D8cpjS/K+NQeLbGtkNO3WV++KJVDCcCa0YU/bypZngRxTHkxgj5aANEpag
J8GVefyyZpHv4meKUxLKCyuqIBDOiPEgUG98LIZEon9m8DsxXEPFjoYyzoLd/A6Y
F5bpzJ/utHYIz1mo5kU75yWP9GDUWECYpF5mdnyxHYtL/yrOSK+leDTRAUvaPMWF
GoRHxOQtvcs1GAGp5CBZ8kaLUJWCtsustq7RxtlmL+MVrP1Qurocul4ZHKBXWauZ
g85o2ubfkzZrnVKP7YBQjoXXjEGDXL4NugK3DDDLepxVCmy5Hl7dw+6vDZrsVhzc
6uvGAroL6SM1ehh5Nk7IFxuk4AQYJfgJADrnO5L2hermbG6seSMxnedkDgtS0Tg4
hxucFLUX7IYvmLUZ873nAZqN8MGg50krdFQSAMyLFD+VaZvON5Jzsw9TjEzEX4Np
kFVTeChzyq38vyY3VaBN8J+Hx12nHDk5194L79LQlC9fu2181vHvgEycyefgQExb
X28cOVanCn8HOUNlMNnvoCnTdIcM9Q72PdnBGmPzmwzctg3j9PQegKpugFGFINcd
jS78h+VXdPz1g9tfmuwfSPURZMe7nidhFUMAEr6hE0uOwIoQRd6qjCaiR5Hny729
eEFpFTuKSXTNLSZW4pAIMlo0Jj9Br5V03Kij7SuqIiiJsShGRMEk9OaQ5o1GbB9z
3OFhfhbL8PsVzAYX6zWzmy6QznJawqVYl1sSpaHphc6uO4emUoG5I+/9XBzX1lie
mFhIpCvo/zWsbVHXLbq+KrqyljXhQsZiTAHlRnEAaj6Cs9+nUSvaxCjTR8gY+Dsj
0J2KcD3xLfoCRiJ/TZUvCFiyi/zrfxAkHdEtPA0eN95nNma3vvpboPYxsUutgxyE
0EDFcw/uwrW72tl7G4ZX1g56SoG0glfNUTUBcCiXxsr95kvKDhxehUwnHyme7hjg
dA5qBq8Ds4Q7mc7BixscboxLepSkZ6RR5yKVZo6EF8pV5mPPQfp+agxOq7ukgWHd
yWALDz0Pl1brMjgKGv8O9m7rvVfrK73DlR+/3P0sAlBgMeePOvIZODeV6EK2hn7N
EdQqUJLjZW0r4rcYed83Hddzzbz2XqvLMMuj3WZxJVmwGg2fFVNOgOZk+7t34ayt
4P+dDpNDmblgjNz0/ua6xDutAzYIJgqeaVpyJHhakfXntdGYQkjOmbVTOmyHb2qg
RDA2nWHUfpdGwI0odcLswJj/ZeieFkFxF8MdWvicaNhIlxzRMLWGAIC0VkG8HNUh
K7gOGwH7VPprv2TJkDzzpEKRdVEeT183gHv77INFcYaloJ1fykOF1O1wmvkFeNLn
F6fg4PYHgL+/XuUjp0TE/n4h8DhxlRmkR4y/xGDcC/GkpWfvgInO2NODG6r7Mn3x
ph6kEb+R2t+ItyBGND6Pqy4iw9ta5oL/zWZhcHvOgkFe1RPWHndxBJ0c368HV6gS
xqRwjeUNN1+TWEkNqJMBkccImqVogSn90ibQboERp6aN/kcFSvjkDjSgldXAOmUP
zLVn+F7QtGbSKPuyTq2HjWa2ssfRXDdgKyxI/zTitds2UJA0jDLKgmhhSMLNTGX4
HQ1ByDneftWACz55ijYvSIxbYqdY8/piTK2Su81KK+ITFUuZtl4r4XU21v3TxjeD
1WoW+qXSlJ6U+PfFE2rGVaD8WoCpScKn2+HwzBk2+EqsNJB8dvf8uBeIj165T3k5
eNjfgo1CyAb/KdQGu1R34s/pf/bG9Vf2Dn4DI7hooHwAbNlTrq5V5p/6n6i/59wi
uOhkDWMExp5dITaee58eZiZAcVGdJaIG3OziwLnAVi25oh0l9pbsPIAi5N35cCFv
xNCH4QRdlskTlS46hILEogrCtQxowrHtaTp533vlWbNzIh6MLdT9MeZhZekjqTgn
waM3EbAuHRKgt3x5X8hk8lyfU2AgCVf2+/LX4DpQu3IW9j7Kig3MQoDpLkF3jvI/
0MLGIBgsKZjZfjwSzLZJo7ltEFX7kdCqxTDsqjrCHixKMkVzxXpoY6Q3sNePx5M7
+mCnifguj4+Au2AQcnuy2R46N6q+yZ3oZUzed9vspRjrWwpObuDtUFIkp4pCaWym
ZomyFWj7zfRKi1sASxF7DuGKHOXbbyDdQScycMOD/+IQaBuG3X4kH+8wOXUT86HX
1YtR4sm2K+R/5uFGWxfP20Wk2Y9XDD6WZpkhhLlWNIHVZB8U/oa9f1yDZp3JJCk4
7V17KhOcDjDppvzt/pHQgphVTgyldzYEFFW52Rsgw6zznK4EsF+QQCd2BN40Tiir
b2YlfosQNkwKQv4jhKPm4Ps+WlNSq4om+TWDxjgH2S8PPtQATBd/TdhCkAJXkJgp
rKboUpgrljj1lOwMwGN5qYTX38/YYSpTWgEQ6W+ecKU4iEoXPrVLkYu/yVcdEs2a
BHLcbAHhqL4KhdyA41np6wfnukPh14B+QqkcsjO+ukpXFfv6DZxKikm7lR9wAjgG
2SqTi1ygk9/u2YTMi1SOaGBklTYhSYrwjAKnrA+SbeJJMBJqehpjmE/9KPOuodOO
SBwcLNlxYvjTnRZhBPumbxM/MFMuXU0ZdsxrKHSxQOFjmCoTQ6Z1nEJuwL9QtTjk
u47FgxIkktpUtd5MSHfXz6BsdkolJdFaRl7pvexMWYkv98eQMS7O5MaUrnTpaZ7c
hq8eUc56n9aEkkuCQNVhJtlzN9VQlBlUG3kw5JwpOvJv+wMsIUNGJVqlGtWSKfJo
KKW52MNeeWWZRGXazBiMgArmcRVLOdFrFxkqWkHORpqrnkW/FnMuX2VVRNh/tREG
ErY8otTjjv/QOzz0AjfwyYMZpdrZamKj4oBkMEyQrBeKS3I44tIDgxQ9YyFpkJEJ
GVNXD7mn2cAmSbwc1+ltKeRRbvWYVp3uFQzQ4TQbRYF1kfj3oYTEYpEpRXzuXhjj
ZrJ0M23ESxL/DpybiIjCFXgQYBeCy6Ol2cXvW/nNpTrZI9y37ia/BYM5lERYFtU/
+I1t6Bu4sOkQSrteUlv0t21mYLAc76zKLi6d72UnhR7gdkyZ2W/YCOmeXUcE/Op/
krusKiAJjRQuwI8boyhoe5QHzmPT6wpjevKU5SaHaM0j8W15xT2+6cjuNrgkldO7
0a0WHf+ukoxYtk+obHI1rs4aKUUrEe7sE63XVYdGu577eb+lwtPyL1uFz5LFSDjg
MQMEU7TwJPj9jXyhR4SPvfV5KaCdNDiLK9+B+fVqbQERxklWDfw7A+kEbFGk5lpv
+R9iCHXW+h/5mddJ+O/BxDDDkgU3NTnlpzmLpODjuKyKSrrNS9lgK7L8aHG2/ENP
ucSfSOumgL1i3UyTDvR8HJvDwNxZOtnKYQHvwl5lxdFtOLBL8b1b3hdAw0YhCZHf
3xjtgFkdK8agmUelwxKkmt4x2i3HyssHpJIqINQtGll7XAC9DDpb3yd2bHKcvSdv
SpxNloPTb6AkZ5dff0zo/P95ZWZJfLivy44vc+WCVvee3LK0Ygq3kVLap825yHMI
Mw/OUxaG/z8JXhBAXyP77IhHNWkPsLHsa+2vkmKZrPYzZuuA9yYyje7g78BJbP2A
RyMYXBgGcb23pz/LREE19Qg/msnVqcFXMMfZhh/BvyJXFXSgQtc1aXMF6HtnpH+2
6ofd+Yn4qROX7CjJcbmQcrVK9qInA3Z4H3VLDCZaCmgjkqT++5jXqO5cIcvwf3Jy
8ZDYuUociCB35uAe786Ts4WwknamIrZHNPSBvDi1VhyLU3T+Y7Tz38kC4URI7EdR
scY2C/mKYL4DPWQjEfi0J29kH/hAODOxBqR0L+XlSg+ybNtVVtmHIWLw28yyeUiU
3uwqe4U5mXaOkfZ3yucAVN153bQ/5VlaMmNHz5zN4MHQxwPxvxq1Hw1f/M+ksbyL
JnzouHvTV4VVPaJny8oJQj5jycxJufuOd0KnPP3cQreBF8YO8se5EOyoFMXvF+ub
X59PUx9MHQOeQA60m2iqm/wt3nv1VBslH28HYJ8j2+hW1uCj+w2wHgXA05tjyTzS
3QPog7rfRCGwKxuKx6Mv+zNOpITe1kMqa3gsxNgJGNKZumtdrelDRhB0P+LoyFsU
AEfeRzgDdhH8QSPOESzDfBodhEFm29J4LSFTuVoCXLXmmtibtYQrwHoDBqSxXAmQ
LckTSRvmKTRFoJrAiiiaOER7mBs6Nb1RxxTuJL3i2CqTP9BtV+BF+wb0HO4nZf1a
nq78uLQN8H0S+8dOaX4W8jIxVzZk4AZO8DhpOKzvIED4g7ypQullthotYOsjVUsl
C/pb6RLKEfq5Qh4DJ7Zw+2fN8UX/CWmv7qBOduZaTxUKBqk0qdURIMB+LNV4UtsR
uI7cVTbV6V4vbw+urL9zbU/1K9nCz9UJsAAIfwoAD4I+O7TU4fOcNmnjvVjA3f9X
61M0/ErrzJ+BlQQwWXz+T9GVO47N9H8LYiOXzRioBU5S1H0Z5thqJ8A4ok+3vHqP
G0zSkaZRhBxm/CKjrKZ6h3SxKmgxCUT9pfJDp1sQ1nKO8y8CW4YA7BmHu5Q1NH2+
jEDVm8NbIfRJmMQt/OjD5tli5WCYi1jYW7m6QbiV3NfLmllfST0/z5tmRWcQOIKT
1EmT5I6ycOENeLtkRu1Qs/Do9zz1YUviHpZba6YwtM13jRdmQrzIShE7zn0kSkc1
DJyk2l4ZiX029jqBPCnaGHIm0gwRYoeuXadil6bJR1F6uvWLYUlFCJfoPirLygm2
awQIBox2bcTeOcAdnYDaADeZ+A6CNBjghfRNxjv7OBrnpptJ/PaFyx/QzG1xr/SY
DC0LtWEQI9eYJ9hKBOntlcuVAFJUrNFII89FwkZOuo0S1rhJd8YHsPzPvwmHF2e4
t8h1fUUoYPhrWEvf3JRun2AfF4TO6UCtbm8iqCF5IJfqnRa4onWJdrTspA2LQH4U
avurM4opj8FFXWSMzGl+53Su88JDGEUazt1Z93a2FB5iU3K+9RwOdnc0eJ/l9yPH
NVxHv2m2t85mjS6IvGFT4315C/hrt+gCdZzkRkzKDcUCZXBOH9Y1MprrTWR2NRVc
vvMYFkimqBs464y23aRA8nrXXo0tqR5X5o1QdYLwPThSUO3PD4lU9+IlXZ754LTN
An/jsMU50QoYkM0f8QVrTydnEX8jZsn+qetQV4jCufrU+2tED2pJj03RXaRNLBdh
qodJyQHgubKAwR1yRz6PUGhWyjhWMuAHInoHgA1gFGs7LtyuTTl+fQUj4dJdKDL8
S1leHm/kDusoqU/BkAp+oKKcaPxSDEPTtxqOZJlCb7rW1KgfJmrSEXmpVqMOylE4
nJ39FJ3Dsms5AoLm2VDQPeZG/QJz4OzwrviuWCrmnOoa87DACzDLnNhHhOB/NtrA
tzKCl0jJLg6+QIdkONQZiNdxzdPmNKlpM3jyufzW6H0f+E19vHFTwtl3TKmZOQIG
IW9Z+pVNcxJ2OemPG0gtYL/Iqyzkw5ZGCwVQM6m6xNw8L8E7AbMaqBedo/3IRM/L
4BUX+FzeUOdboXUXr5CkJPZEb3iqIb8JAYkcrr8haxj15Vex8izNnQXJ7JbDj2bs
KAQMIuCNQyiE9xfqabJ61MbvUzSxYl7b4N92JinSaocLz0/viSGoE8oKbFo6mVWp
xe/WIxmzom2BWQjWIKYBHtezmpHp17awEuxUtdyX5YcOSXQpKqUfOzTjpItVST/S
FeXIBv319iAnz2MKWbI1BRTJ72Ps4rEozf+NgkNQp4p66hKoXTNfX/tuWyLIB0nC
ZvHSvVwi6ksgYGV5llMe8HN+3LnuE8+LEcw7zVMQRCq76MMPEZ9rGif3c7+w3l5o
lyFVlh0ipwFi7n/rZoE2dqkIum9X6zWIWqoSiJV2s8zNCu8Ci4ntuXQ4wyQBSIsM
RLHdhyp83pIfoAGOlg1t+PvBkYNTmaaEZfgJdKRmhAGyA8RSrjIWBWZ5DJ7UWAbT
NaFkEcgyc3l/j3d7K/zZE6FXZEv3A9tZO6yP7I+BZ70aFrJ1PWzr1YW2Q1m2tmW6
eYeU/kHi2bR0VxZ2O+1GYXoz1cXUTFfv9kGIGN1ROMLQ8tVNzVXozYh0lgc/6Bhh
pwKCtaVWH9ahCI6UAzP0xMxSpreKglkn7WPPOEkrFLudMq+SWHYMFjYNCycXxjtZ
jQbqMNA3UDLRw7jW+x5AUAAFAuNPBx44HXlIPbW8Q688hMihATa9MERBXmEHtDJn
OZLAsOLW5LVUJ+MNQVThwBkow/YdX2Wt+9DM6nhA/vVUt7Rncun2fHDw3M5VRMNU
QrIgAiVcTTW8VrCkx7y76U2M7cWDF2OvVGrT1tBKwG7b7VRoFArtrVPs0gd5roO0
eyW6YIEfBg43w7lOur7kk/5gYwkq0+su/60CNUkIhjqU4Xhh1bPeuhYXO2hrLC3/
vidN3QSBmxZto9eqg4VqBgCnnBSN1c8aDb1JYzWNChO5qR8WieJlTsPxTYMe9/NL
F5XXtPIP8RGFlwjqdoaUYZxTFaeO50+bCqi9+Umf0SKRT0SIshyfVQjsMIfMuV4l
R4IGfQngvsKaHHpf6XQ3TfhGjc39T3GB58YJo+keXfmZqTls3lIwflMGDHreIdmt
/YrRh6rVJyRPUeq2pBKIB5C6ZuuOIk2Qpq9C/xTA4NLeJzN1gCPUBclhI520A/Ky
4xdLb21V/PQf5TLu+MLz6tqXUtathTrwJTPAUpcRZWP5mobgnIVSfRp5k1wPa53B
+2/T8rrdxMZKaremHhlw9c26mVEa44OFPxFsGEwLwZW0DDOGqd6R0SjLTcpd/ZHB
l+pWM6mHgI1evdykGehd7SIyXTW3CI1sHd8EdZXxrr2O7BQsQTo/ClX04XF9dhYQ
p1p6KH7jgZ1YtnVq9pthOBUtySyZbiCXGbTXMcTtXOJmi6SXYo2mWJkVKkQZVA/S
nRwgxBxp5HoV7eGoE2xdZ/czFkD19keuIXtbw+N/w8ZO9hcC5ruzrtZnCuQEFCcs
z7Tlgzci+LRXh+Qy9fdh4WH0O8wcWPktNejbRIcAOq3eiruaFKVXmtljRxUurZEF
aHgk8HhWGqyxLrAggq4T0bceSqGwzW51YDA2VxuyAvZb57eJfaxPJspgp1wEwWPo
w16DR1Qqf/cC1DhJcrpq973cwF2yrRg2uF8K48zrclIXoOUTsxMKjvzoks0OUBow
wEVOy+u+Y4yS0rYmuI1dOnJtv5kwI9PHEQo5cF1XPZ/ldCRdUx1zBAcxS18u5yco
9USoLK/UlHZlv73vvUJR7Qst3kH+Ynp7+x3MPBoXVGTQeTFhjHsbBRRXYB8QN9CL
KYrYWcCYfvgNs6/GcCMKIg==
`protect END_PROTECTED
