`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KPbfGXj+jHHCyNoueIDJ6Zkip3bqkSVOqVklUCCzUCTbrC7JOoAcwLOedSqQZp6v
rV77xZxz8gqPf+tSMLUwzTv0bGZ11mHW+mKkmk3v9LfnzYaH2DqmGo3+ujWtu2iq
DbPxiwC9bKPPseoMG7uDxY2MEmcJiFeWpBeE95Z0XDLIrgUCbUGOHsTg6UkD+wNS
SbeOKO8YyH5cA6eobPbbbzQQHqeF/rEDYD2JXLXOY3lELrv9vnsdJbsf/4BeaLkr
K1ADFUW84zL24Fe/ftiP1v+avZ2mYpF73bozpBs3LlCSCVoj2cijRfa57KZ/VxYC
v2kYa75KhxLQomkLxdYwRV9Gjcj/GNkdTeaKszSMcxDzz8bypKIQANOPWZBVMzjo
GUxLpQCjjehWn0N23Nzszdkm7goPhzkdQEDK/HlOjogj/E5EHVWI7HnwBmun9ltL
VExa7lWPgWNqBNCo5/UujifwBraqRsrzfSCSJCW0CB2YLf6beKssJ20GfCturUlL
3MJRtInPWy736I0C14kaLiGyhZ72e6tVoxxOwsN5TltmAZ/d8wKrhLvI7YzWM3uw
0FYm4fbnlM1TehucEBuYDibC/5Hq5cAbeVJqdYy7oWwHO2I2Ri/g/kO6QM4+z7dt
fyYebxTglMtMmZ9Ilt3om6bLbno0hQUADHoNqUaup+mY+cgb5d6w2ur7zqjQujO4
AqrCaL37UbZxmyzduQkLBQPBBfW+HSWmFEuIbTsxMIUPJMS7/tB4LB6Bh7p6cfnc
LfsOTjIlzkeoQVIpPSlqpGY6Ea/nbLZgDthJeoYb6cGH+3p2ALKgs42hPksLgz4c
T5JyElerQCySJjWQPQowsdEHN7l96Ih7BNCDtOBMYZMf7zDw1GsmmdhWuPbMWhsE
w442+rhWkltLNLXtQbyRLWKpiMJgYzkRj4K2VgAe+HJz6eDIBWWBlu7zfyCJDh6Y
HAol5wYQ4r4LuHy0dmo6plz2FOXqef4d0XOkTuQByue1aFusfcMeTLYRcO98gLzA
Cr6y9LvWi34tcg58apWtagvtBmvZn1WdCnqr1P7j/jKoiiuW7wtIcN6aP7XPrP/Q
PdeZ5162y0XuiKgLbSiUkucUUWrksJ28MaET4niZfhfNVc/1yv/eNR0SURsepFgZ
L6NZ7rtmZDPhyNrXfsZJm4zAxSAOWmzvGtmt1gYsS8OoFcdDRMxtwKpwl4JDkJ4x
sv0IqkD4DBEpCgJUazYZx6OCoCEpqh7bilccPsvD165fiB3HxtDUtENnXHlOLrP8
MzRQ/kdRpVDMZV7JyxazDmeygGCGb7fnsrXNIycqBabbalxNKfelYvh5KBr56rUC
dgza84rEiQeOo9OXj2FMeouYeiAzuPuYPJoQCTIijED90fuOiMMTX5ESeQIijDwp
x9d4G33ddkE5YtzF1Rtkk6nwfBTWwJFIZ64R6E2x1oemvDa3wVB89xarPFVmJRxZ
l3JzbC1cp4l2OFKe7ICkT1y4i+SnpfUN2I4RhNfC3RriHhK7elibXMi16tTBI+th
sP697vQFHL8l/IAJn5sF2VJ9nAe7D7oyIs0YkM+srTWJp1Gd4CXQRKJpYEK2MGLi
5TtyprakBdJTieu6mSG3sxYXXEhlFtmEcKZ3kFkeG8X0nkI/LnrlRBW1De2beqBN
AOFeQKTR0k8u586mp4TcstcoGo31Ux9ik0fgp5Ac2puIjFUIg7LxVkUxWW486c7c
MsRjp3L93MAheKDrWudKGXnbWfhXOJ4NPYHYBiQ2YKw=
`protect END_PROTECTED
