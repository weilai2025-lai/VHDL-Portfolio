`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQEFQ4IeUe9FRa57ejkmiyfJhh0g4g9OPjiNBLN4VBgVJ9Mlw/61VUfb46fw7up9
65KTy3lqN37HA09e/6CWVZsWy7euVBGDN3q842Be73Il7s7VSJ4l2dU1SYNdkPGm
pbEzypG8iLUAMic7FzY4lxSXh2J63I2KA7Fs5tAxno67n9m0rssZAMiPyr0JwVKQ
JLJtSOzORyMCIvwkPvcn1wxLmjpo8cw20ugFjsCv4iiY5nIngiSIjRYR1PuSbr3R
54dR9D91m+DenUyQGseL5d848Q6n9Ly+UB26ZHUbhj4BdY3DGm4sX2QrG7b8KFng
wx/gAA5qkvWUWpAPUlx/m+ln+rcmWJqsklkr5bb3Bb4=
`protect END_PROTECTED
