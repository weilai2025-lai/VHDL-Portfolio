`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
si5m46fLgM6BoZx6A2mpPWt/r7z3vtAiIJoeW7yN58wPKazRbAZdOF3LV7fFdE/2
l53BTTaykgg19VYrBM4MFHkzlpfsaqEK65mMPG7SK4SMpcReA+/JJMq+oL1R1TmJ
oa+jsry40eaqR6L9iN45ppKI6/aPway2LvStT7ZTzZ9cpuu0dDRWWH+WR4It7+G+
G7qKkYW0qByh7fCidx7q6rltk59GMNGsKkUvuofk2IlzaV6J2HcScvMsccWN3y9r
6yldAEaCSfnLmi771VLYsJY6a2ahmAnHo7utFnQDgeNxiqa0UvxFaBNu6LYNlvyR
kpW18c2ecuj0nNWRp3HYcnV2usWKstGxOXu+bJumW5A7CLPHYD9dFjXFF+m17Swo
+lvxbnARk5/KbWKxc2b9e9MWh/s7n0c3n+OiMSN7rK0KuOHKgBXkJwgaGqLh9WC/
zwdpEcON2zTEqcsDEdTIj8UF770Kqk/3kzOb0CNLyEihDQ709CwQ5fmXf4q3QGMR
rVWJnR8oMQ3b+GlyGvhh28yZW6f1mIznZe3arGb87Y/ZtZ8Yi9PgQdneabC3f1Z5
pjwGL6zKAtrjGYhu+lKbQM14pB65+uijPG90RlVsxdnC/VL2gROYRTWIaz0QkPne
+19pm1ip8A36heeFQqJ+nDUo5Q35PXSLw+xy/NGbbr5HxM1Ue4N2CT5RqssIr0W4
iZkXyGfzshtahLbaI3VsBI8RuuAgZjAjaNc9lESwaug1LuZ66tfR9PN+Pp48Xcnf
w4pOvkwEf9pPwy4hyI5HwN04WIjPDS8zTk4aSDx2j2QZGNNhAsYNN2HWZ5G0sr7C
MxgVFeiS7nUuuXB2YfnPFQCcQLeBanb4L+MJ9J1kX4ZTcFtLbHj5UFBrjNEVMaRV
dIkmEanCEfSsKKBdTpGGk6IzOLdcBC0X3qih078VHZf/ulZKd0oCc08+LKUPdJou
kssuAdrbyO7e7nyHWPIvZknKGM2Yge0+oSoXyDNKhTkllLjkyxU/IzZpILoXAIH3
CI4Iupx77ILTEUNzRjM9fZuPBPqQzNa/yI/XaBYYTFq1Yvh0adZ3T+Z+bOnE68aK
Ro3FhKKzWycCm77UhXcqjYqiXhQ/l/zoGpFOXHh4KJtYoCVa+30jzC11Xd7Q184T
IRfPE8SjI44ws5FDdB8Wcw==
`protect END_PROTECTED
