`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKxTltLYvt5gnH1t0jnlYQv1+aK+hdHOO70wa7voHybGjodT4x2mqp/cZcaqplUg
qkY7qvGG3q8UcTZTrJJxVPjFC3hSn0Uo4O4Yu4xLPHCRRSflqc7PYmHU5/40xn+d
IpYHvVedYu80FO9StW0JUtU/xvIuvl9Cbh0+Lq/AMe5R59MGjGQ3aGqsCyVoHfn9
7hRL8AIkhPIAxj1Cq6blgXWh6jtIXSg4LA/gLEenQwBZ7SmnMcGaEh6qMHyz8/mm
bCP2zUhnCc5V7MZYS19AFp3y+mouXJHrrsNVI1EIZG4a9FkICkjpkUtCSJt7Ep8w
dDD/QYMilLelIx8wb83c2dZAP3Pkj7HtExrrzape4kbkgEGuWgQmL9oHFuOIsJnM
C+xNVUFyyDxpQebuCwhSt6Q5dm8jrwDaMN1ZBbnTCgUaNwKjVPVA/VnsS+TRvQa+
oT6M7IAbAj/5zRZmlgEl2aeDat/WVMmKuQUG2dctK6Mn33EqzsIC7EJlgMUrL82g
/OgTlBszTlzvtXadZnAihw==
`protect END_PROTECTED
