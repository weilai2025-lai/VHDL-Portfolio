`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7FUI7Qt84Ahy2TQrMTDxJNNamVEGuVuE40eqCQBZlR4SOipT7gFil5YrbWLM6KR
5x9ImTRd8mNoAAntLguc2ypM5y7dMbhU1Dg/sRwmSbApNNeEMXb+liWxd1o3Y8Ca
Ux06B+lcoYI0Q0YXUgfKBB0vnHEY3gdTbSOSniDCcE4qgNaDh9O/+wr6hdRAqsay
oZzy54tfmo9gw7NspbOIu9E2lZshebwZUYvOppLklhAQZnIbd20GVpswJUoKgqtI
AQhHPgKJDhd3HpPyjJk/DQmHkwpLU8FjsIiappX3/JrtF4PM++7EWR+lW9cFtd+I
mGiASG5aoYVv1G26RfH/oOA7+eBxmOYBvrpBm1xxUvqhc5y+oj/kb6qgbux5hoHq
BELLCLx/8Cc8ZLR3SsclNwndcR9hG9BnJOLY3oz4fAcuMnwkxGrK4xMHTd0KcdI8
7XHv17jOoELYuS8djK9xmNSe5TsfsYcgJ3JoQKccF6Jeno+sPmt5l6N/sL4VZ+/4
tWVSSSpSAiCG5WRov1oGJfmWlbOck+2+FhwvR6dUcHu4419k6El7fOhbRwSyDqLV
DrPszIspyKuyIdtqjFFT2qhr5ZufW+am0bRvTtnMFznL6rpyi6M9Cu5aYJrxbJk7
1zMyPOUeunDUEChDajP/Ryd+Ix2d86NoWbY5hn08aGuKJZfyHlinZ3V0cFtR0uPx
p7XwlQiKjTWD5Yf4By+iMQq/FXghZZEUGEXnXFKXGe/Aibsk51TAOEucdy7P15zY
t3DOE8g/RWd36gv17SFzHx8YtXJwcLDfXBtHXk+vol6Zzb98zR6iNbZG4wBJTV5V
um/F/Xs/IwLSziSMduXG3Zab03fCmq2VZ3+AT4WIiEimNCv2dfq4E1yxKmWoQNea
CVFagqG6jjEsep8yTS4WfGo5gWY42OoSKsLckqLyd9Fzwnsa1dI3Z9o6Tcz8SIky
Gc2FLiQxc+3S/l6aeLSTxb32ue24ZmdXKlX2i6trW3QgzSK3HXPIbcoXBDDEvCZp
pXJ2HjKqtSpt91uqXgfbB+GLoUWVXDIpju0YB46d3YsaIqJaGH/8KPG6UGV5mWBc
NL9X/4skDSRY30iufCCeS0onM1L26XGsOMXJeW+nG6nR3GiHNKfyiWtaOCIDLJgL
HpAnZgxzy72j5TKLby3OXuxbys7Y1zozPQTJbCSP0obtMOMzP1qfUfrJMF1AY6aB
9OVM3W0KKf80dT9L+K57wCaxuznNzfMpQQyypZV+OqS1bEtrJ00oC2OMDhlS3vDP
YjVFjzmTaXJVnUV7hpcQ6oZ5CVqz6lEtkmfe9jT0TZ+lfPPYsWG4Zsep6Mt3kTST
HZ0DE6hTDo0sOYblc7C/g1YA5lXxRL4sMcmjKLea2EEF7PTaVpraJD4F3AfKxn1W
oCICcqCgEEnRbGlezHp+dj8NDGqbR8RHu/UGAatRj9KXNPw+4U4m1BOdfRbYoAJ9
7PNYE4gqdbJn2xLidDbh1Tjg7qbVyLmHijEfXpdfXh4p7Nmrvgi9qrHbRuRFbX1P
oeg9ODEQoHY11FBug5be8SxClYSa4WPn/mk9seR5+m87wmBqn9t3Y2s6oIP5gOg8
NGDF53qjluBgo+ct4xFOGcI9xYxnzMpKfTl3XScxKi+sZwMh2g9EyFxlzp8/PZ8N
INd9V1xmMM2t3AUvU5qSDQtmyg64DsXJFrj7l9alEjvUtSXYJC3IPBCoXPkfQYm6
Si2LWpQUmq+MyQW8ayb+ICBs1RFJ0a8pia5oysASjc3umbCM9EZHaaA773gBwuxe
XNuyYeDXjo+kiOw3USzBcPI7Iyo2gS/NEmAPjcSHFIkuwN9OhbZmJLwL+7WeXwAU
cHDp7FIy0emcNKVir2fBqKLfQ1kU1qVy8hOAtwzjGwjj+oWbGbCqELkAUyY9V7+q
E3cZZKFMyQu/Ie8h0IWFP84PRXIKHLgrTKwIiwgbgOu3XRCvXdbOYrSsLw9FCeJA
XKHECDNjVRHFUC/AI3ju1Y6yczER/eaOZjgnADX6KtSTkERzI6uuXP9zoTQFfpR7
UkbddTGyzIsUSQhHwA3f7c+hYgahjBLfErgDgiTxpKeFTTE66p5+nrOIKcs03bHW
99D+WOOecGUpkq6+fI88hHCIbGaF5tEWLrY5dtzSlHZ1TgtbYeetSl4pe9H1v5PJ
pscVg5JZ2SPWRlxLu9V7b7ZQMymGx1M8vfJ/8NNxVIqEZCtUSioVTJEJyNv2dNrK
/1pv9ZTwauzChTg54v9puOmS67TOYcPdnOnI6gpEsEr8doj7Wyu9Zoj2bOuYxSE5
scaOxY1TBL7W+ijL8/8dYFPQJPs6WovsuPiM5Ki4N5ei+mo71rVoMb1Wv2NQDwE0
RdmBChWRnfdSrlmf9kVUWUG2dksjCWgbZfSSBdMEInAP66y2ZNa+cCdosdeYqp/O
`protect END_PROTECTED
