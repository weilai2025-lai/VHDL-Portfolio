`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZuPHQnJ9rGEPgH0XFIOypCL/jtiOHpHrt6WzaKyCGTdlgMq1I7mybJV/kPZDtbp
LtO8NOOOJHCnmjD9pUUD2RNmJStrD5W4rVgL+IbFTKk3kxonmR4vgQzPqI9e+2xk
bnI9dadP8UQooden1UPTje9ncbjCALaHwYGw8juSCw80t8jA2bn/MWZlXhWrTaiD
D3DkZ0wS9L/VvSqRcAsCW84Qiop8ZMoxDcQDv+N4ZAKHyK342Hmfj/86bOqEZfYc
sugckco1u0fX9zqwu37Mg3lwriMpc9Jvr4GSSsMaOpJ7Yxt4hqVtwQ5lT14GtW64
wyl+5Va4CkjkCCPE/xl4q+b2SfAiixzPPoAVUZUCdiNsamveWBtyU8ATlS8wKOXo
+7QWWTpNaE7gFzVL32Y4+/JYF5zVryTIu2bx4STURo+zOHlqACDFG7QDRiwwJNVw
OOephnFVVCCAPvQMCe/JjvEB/isKobjFPtgaS/xgqJ6rQ6hJpG8QcYBhA2Iah4V0
YidCiHb5DEd2379yx7Zcb5r6ch3HDIMQZfarDBPWd3hkBE6+4yqDBmHgZxCJL8Uu
/l0IsloaGTKTichCMSp+hOx/8ggDE9GR0lroK4DL3aOvJctPPdvidKaLHMwa+vYG
osSSljxC8SodikgVLSoDXYFk1Xmt0y6l0RWrMCBnaBv1PJN7BytiwL2qRGFEN2Z5
YHK6mGdEvsmrbqyv2cHyYYrXrIXrATx3xkM4PpY98zicFY914X/7uoqWX66es2Kn
QLZKWRXQ4Ty8Vku9KYQY5X1SYuGMHctulyWUg/fo0v76H3uPd9HL5RXrKxGiwucg
nVbtQQ+QXTI2fIsxwaGZHdnFqZ6DkGvYG/YmNOrz1LwLQ1Q8vP8ay/jNlyAbISeg
MP/uziJMkHl4M8TqHRJVGGtzt4rxTl7XgaESiRLL1jygniyZr1i/7GeMmaEW8vhS
rLjwtcOwH9nZKJLSlNkt5y48wR15ntxuxzXNBFgwEskteVyb4WzFEv6il6zs5y+G
GgzyhDjneA/iWEn8QPeozeL5aKJUehMY+lE9zlnEPsMIdIpOnIT0hQf1iL/k6FM+
KNOg5455BaI+H1km2q0xWroEUGPWVSMgvk8T+R5xaBg1xxjamKMcyq9X1fJb4DxB
FfcYwsHbH1ZtjBg0UUVHXkJsLFql6KnVta5ipMQCANbIYBZNTWaSEXr5+SQmhQBV
yiB6Rg8mz6TnWQiLuUQKq2FUd9EaaTSMtknbeEYkEONa612GHGBKTBtv03ZWGr8h
SIBDTIu8hugiqmYlraozYDHJ6lHjYYTPcC4yebN0T1ZpNhgDWXwREUKW4u9ZOFgU
qpbvO6KWxKso/7Mo+JiqrqTX71ricChx8lPf5d5O5cJGliJMX4TZsnCHsiZMJ3c3
EG5i8MCe+WsSruw74QyUuP5vKAdpE9xcA0QfBlQj5PWheazjGQDLgQscSC5HeqRR
dm0Pyoqi1YAdN3ONKX01qc2ZhxMNIkmyXE0BwJIRdNWusuecYrtnGBvOzQkJLFEj
B5lTT4vL9+1fk/woe5VQPi1eCWfhYHFhEklPvviCHCS6rbgJIlF+MuZC2xLlnjhd
kczJ1jZBBOa8w7UDSYB1xwskgU6fzdBknc1aOtp0i69xo3/UxTx+c7qTuoUyWFpf
OcrS6eAUVgKvYstv01VZq+eCse5zNcsyc6T56ME8YsgI9973n7hZnS3dwxv12d/B
wjApwnyeZxr35KEh5yQXgfXeg861OdqsezHcW8bXMoEk1Bdw+YhlNfYhA8cmqXmE
i24qEOgs+s7M0ZUSK4L7e5udU7AhzfQefyfbUu0bYjeg/7/c+jTKqNIPqKbtarBw
riBDhZuNiUBwPbOlN7RjG3Ws7zIAMcp0IZihzPjZ6GUvw1qMU7KvXTxt+G3lB3XI
cy0pZIANdJlrqDtStIpSBh0r9+GlEH3yK4c7azU45dNroNZgV6jEYXMk/EcC8kJx
cZNWNHVCEPogsuUP+dTIrRGpaoDssGufvmo5qx+i3OlfMexOJia4AyUMhSEXq/mY
5+7KRJKLNUAoQfHWZIxZsLEonygrAHNhlPYhMBT2YOucDmoWrw5k8saaRqKW2BtF
VA0MbSutmfQfgYOc2doj5w4bgBKI4nHLMyKOlERK7CCWqVOV0EIdtyTLVlXj07PD
nAWAU+6KUTsOgYMFLC9tP7AepeCmX+GfAHVig4UMDyQKZV2bAUJ/62PY0b8zu9Af
PCIjEpKXpCmqR1qCBvu+Sa/IyBr4xvQBIxnDR+2iQjwwgZuoQu7SW49y4CUhgAl7
NBE4z62c92J/PPMy6UxnzzAk1krQBy9yt1Pbk8ABklC202dEu3+lb3XsOi0XNir6
/fnRtTYsMsCh3RJw98pVoWFBHlVpXs7nYwWnl7hFW3+SwvGWLxE8LqhsmotYsBgA
/MOHgSRL/Xoqp7RicjAwwrMfEjjhDaCXOmjfaa5td2ciC6uYW30Hejpe7jyDyjdf
eMdEugGSUPIkXRG4WI4xifP3sIoqRWqVZ8Qftd9ZjsumUd0OJyZl3Sqg9PBKNk/Y
BvkF1nJwGSpnRedFdgU4tm5LNw5puKfirHc3JIkNG81dQGFWJgy+nSxOOUowVY9m
NCzhb7FNNw1+alUfspKVevgrGBFvxWFtvj4DWlCE8ZUX8sxkAqZkgrriKCOtJ4i9
QSqaNTiGn5950vHKhOYfWI++7sE6/sq1SAO2mMF/goY7ZS6Baai/KnF2HxUkUOFE
9VllHhSf2RBU5QvmV0kjYHqT//SGJJojsJ3hyM9juS/IIBsxRysWjU7JMDZCZuZT
yfPdLzriIArS0Um/YN7NgloWeu8M5jcrayOdiUo36nOp6Sq3mJ3G7RUZRezOwBuc
V1wDWI6LBn1hoIfBCsaUJoXM5jlSMRVXiKrDurjt1WyxJ1vWFC0nzeK6IUOULpd8
fjZW4esjMzH2dgLu4Q4i92vN7w2fzWWH5xYk1AtNRTGcrlb5wsHE/bLDjOPqORim
Ihyf7lMfTawRd9RC3V8c6fdy6LvBbICmo0kYDceSuGge8xf4zrgWOpm8oaWNmXh9
kpGsDB+fnuLo52GMyyNxnSnFaO3Fm9bS3qjEpqa4B1Ap7fpZf8BcSP2X/Y8Fhufg
E6EJUxmYyrtIzz3/S+0J7YVZlqtuwYTSkHVTM8/JworoSx31A9Acm/QPwc2hFSIq
7+1tuWMyBuTLBiBVuzlwtlAEHiIRSWPTpRh+LfJTAptlT25n9CzvX+V0Q9mbLvR8
XwpoYzOf66MWJq16annf4yAPVZTitPcX76POwkBfuuXvfDgMlrItQowM/TKu9Y3E
CHiQZRsx6Vu5jf7+OfTjQ6HUG14RJHDAmHpdxHo1YfuMuf7ZvQwFWuL2LhxQovJy
UTP9oCKXukJBYUTt4ovRIXSBXc9072g5z+/kbO18BKk1OJohIpLIEoHj3d4hxOcV
jEh1d06fjxu93KK/1WQwvjJFmQJG/HjFnSXpeHbsP8MzBqaEb5Tgia9Jn8E2YGVO
2XxAHsVHUv5Z5dfdmtZv9s5hmtNmTxQkAisgOZ6DsLpDEyXrviy9zBugRRAWrrmE
WwWdV22wGTq73rChK25TE9EGBLd1qX08EQmkfo+rQNcwl3ARBBddnD9GsXzet3Sx
YZh7IKUPvIetRbNrb4DYNriMI4ztz9YN5/2uoydSVAJ/0hYlhQISvmkB0FtfBwir
i+xFpZDMCFTvEYYbgBiiPqjSDMUcTJQumhdC7hUSGCFkWhNWexNmx2jdOZfcD8UQ
zIC6eaQMn9T96TDjNYYk0Hu7mOb6w/5mSR56ejnzSgXygPsFM1rayBSV8xueYVV+
QKesSXrfwk3epJ+9ZwEGK+SlvdF+fiWU+jBYZaT7KouWhX++0Jw+qlpp66ZCiy6r
VF4ytcNWqJfjsWYi+IZKHfrfCwJ5t2/QhqOReKDK0LZ2mEZjwpNy7qAsVmZenLYo
Esus1F9o3ZeLdi3exV6yRa+SR7YVehkTm3bMRrjqgm+ClQ2YoYcWb3fIDF8DBiNY
XqYgwodSOUK0oQQbZZeB5BNi85vflQDeNLKorSNgjpK36HMntK6kb0hAzNoBogLy
UfLk3Z/vL4uelYCS7rP0ffOgwh3j8aCyWnQ3rBbATaD9GJttfRGKV45bekxSo0NJ
Dyh48hoNr5Ya9EJ0MPbCYshloa5CdZfAkiyB275NAhWTYbTSh55FxtGVdiV4vlLr
SQ/VHAJq1CjgAzMz7xrSjnWmNhy8DmOGc8EXD3rLcIiSLWHLsLgxi4M1ldSSRdzn
cVHFw3qXfb+HsSCCy7Zjrq4BuJ/+6LS5vmB2KDiUPAuOZQAJZxYgxTt9Pyvix60y
OuNP9EgqK1dMmDF3VVY90MT1hBQLS7D2DLcJQTpyhMhalcduGVcg1HhMC5R9Cbqz
VCFSIjgQT+cawnkgRkcrIYlgxI+/N5hEzI4iFlUcsKnSE2uV6qvWSRyO8aaKb5ws
N0m3rhblz/lf+kcEUl5SR1W2Q4ghH1BIS5YGjtn0VWQ9T7HrkNt0P96Oq2eRgxSp
5DUqqC+Xkj1VC9c5hsW3Wqq63q7N+8rzdcb8WhTK0DjUkScNc6dJ4yyrkUyafjLd
ig+TckTjFRA99EwnhCLjLpMz9D5ENOQ1Shw8pZEnx6kwGjUNa85Uyej231XgQm+V
gLuQx/ZHNa200twTAa0Ih2UDDmvUffw424dnmytcMCWiZzBrg/sRRvp5u2rOQN+s
lO8EqD5smqy3OrpAzthe5eLVZOfWJHajl7nk2NjLj9ZlDk06w7oeZ6gKQKb9gPEb
fBrPoZJwWU3Pyl0dt88GG7Qtnaww9scwvtPvjGDJ8IsQZLmCqnC4uickA6ZWBa33
f5Ik85Rx3yS0W7+tDatiRKhMpazVJ+WnGu5pOe9mP6/DU8FCClgjD515Uoa7dAyT
z7OAvtZ7xyIwUV8/Y/UO/XD/48npvG3AXr1dwFKv+zSCgIx9Hfx0YRKwEZI27gTV
WO/w5DXwS5SOlhJXxGYZ1nQHJdPbXS9hbF4uSAHuFfXsv8JmTXiDVqIVWowmmOJ8
lt735/Fd7/DSPVKdKPqOcw==
`protect END_PROTECTED
