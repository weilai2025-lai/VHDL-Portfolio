`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OMbaGiaC/VlJ/RYPzmEP5j3S8zFlWpUhqaLEE4aOL1VVHnGwztYBYbCD+njKo8DD
cE/1uSVtvPw7VZYiejtIUQTLo52DIrcsGpOsFtFF/mpYg1T0qvStIOINfY/l1cku
5op9MEJrRWefl6ATAoQ45r8WVW5kdNuDEmDO5+dL3wrT/5QIPra808Hngy8cVXzf
ou74YteBi2xkr3YatcJxAX6EVCaZvQuIMv1LeuwDYBtQ/1kHHQuYoD9EP7V9ywBW
cpRd7Q9Vs7uoT4bK2K+Cr5nS60xO8d6SML5K5XKqrt60jve0mNW1OBcooUQmgT4t
2KP866FbMTJq/Vg8UZjnj5qVxGqF+XCKwKGV2yztP5eoZg74fNGef5MK8DZIZZxy
eJlonRTHlJJXMxymCwoj0lz01GpNjc7MROe080jMnDKBwaLvXVe/58YVooovK4sF
HvMuAKzEsfpyoicLLqdY3cw5nriyN1df0irflgOzkpULzD5lRIekNxU7rOcJ69Y1
jz7gCody3C4VK2fboULpsLMD1DkbvJ6wrXCYsRJCcJk=
`protect END_PROTECTED
