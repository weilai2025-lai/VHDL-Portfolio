`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rcvv46++ZymS6dNLdaUCehWF2gLN3wBk+6uN5b2unWZ19D/WIEnDawF+NSih9gcG
ECa6ECYhf9wRi9gnu65gR9KMYbCGV9Lh9vigUbUDxk1LKvhkZ4Y3D3xdup3SATMk
NRzCTbcTb9jhrTDibp0gSJIHOfFK+JYxTg8Eun06nOOzujDbnlK8PTa1uSDepvF7
mta6GKlsAC0rw4xU5DIiEzqUqYdOndTmof5massBmdL+TbJlhYgEQxkTyI3ILNb8
9yzZz1ANWH+ZyMlmxkEJFVBmJfyvqaoKhuv/jJsOrZTCW6BnPiFVcoz8zn1uXskC
dLSBBY4IlPRdnCtHmvYpLm3X9itPGKlUs+I3cKBAFEB0i/yhwdN2bGrA1sd2BBWr
Z6Upr1rO/Xp/6PMv0AKfAQZqOputl6ZxScNmXRrMoXqyZcCgtegxKzPMeQgndzuK
HNq5OIxvQL7mRJCcVPnyak1YIURyCD+eQytGsqvOA42+ROza4dmij/ZQREZpKPCr
Mh/mQw3RAr6e80qLMBYo1pqW7jYimHG5i+QvMncAoRhD3VfvJdWac5dug490lqSY
v6u023ij4VZLs5E1oclvG8Mlm3xSfkd7SU9Tvf7poFB4eqcBs7U1Fqqt+SVVZREU
U35kgT+TKdGbn+bhVUsv/XD8xYAhZH6MjW1qERO9y/zB/Z9vb6aDKK45MdCl4PQH
gpeXNXhw3H1kSNchv7TtOhc8qSFtMxb7KkH3gKyeM9Swx3ypeHGuDYOCBZsgjooJ
nwjwSpb+K4ibs8Gv0C1P3fCQ0bXjtwx2F0YIrdl4uVfdbPcpIAa3c+0CrJj/4pLe
nAd0jjomSQU1/4/mZGMpwEU1rHhcEL7Ji4P3/tM4vN/ZEFXKYbb/CF086GKTTpVu
1uAcc481OfXMczfZvLbkZBPt/yJsVXd+2GuYZnPBo8OCv6IctassQrRu76wmYVzy
nToDRoZyguj535ZRW+y9mArbgrbjJID85M10h41ft7tw0V1w4iR5u6rfvvweVoXC
iFj3GiXIzMjX9b9r0lEwJX3qVdzYLxj6pRuh5AHZ/vu2MmLkzjkcBushzQaGzA+3
8Y6oYZDOyFwnSSrXqlSUz82NkU5t8oI2DfLjdrbIjIR2/VHCM4Tc0FtZXmZZFMXQ
DiGM0odnLNK46PQUd13Rx69z5nLztfLXfH1dacvkCaNcEuzlG2LEBRMxcOV7ieV5
eGme8ykA56YDCdAcvwngHQM6gn5LlqCLj89rHEKy+6SFdwvDJAhVKhezLRkjqUub
Gffoh7TqreO4lLiXMj/mF8cMZpTXH9jzkvP4W3qwJWtfOJ5aJGnchbshAmWDhVNG
iD3w0HweiCvZvpYzRQdDZze3ZTtsO1pEefmXwKGu9NzUfl8GBHZgpVOS19GjoeAw
NrL1EEKFsXUB4q8F1I5Ggw==
`protect END_PROTECTED
