`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afQLGlB6kJgDDNMGKtjEoeYdX80VAO2gAGvAJ5XcnAE57K8w+p/ynPQeWIhPh+u9
0H3gO8TuXYabMRX+UKki2hwYKyjvBAbDByH35P7VJLDMfdhXhWO5smMt+DnU2gp+
Yc+zkDvZmvq5jvztzniHK8gxhJRb46AKZpbAIQkDAIb32aDkuzKObiddqxqBcWDU
fjgkn+WIj26PMVajcPXTNnWIdNltsfFFA7exePGm7NLdyIAm0kLMRQ4N+Q0pV/w/
OyEJdE/Tsy+HMCUkwOI0NEkZ7SdZMqe/vWYSfWlMfHy4Fawom4HGj4GBMGiypuas
fkdVkEjObLhzfDoBrbDWAemKcuvRSErXpjhA69f3QdpmEyTdATFGIYydFO3pAVef
kF0H0eKJOnTG5j/fJiNcfE4U5zYcACdHFbeRFawPXdgQOO5+AB2sDRcKSMRWBIzR
REu/z57saRcHAwLtr90ykPBmS1oGPzNlkSLR9LqAZ3xpZ+4mFdDKNjLJTdokdWXG
/1n26nMLbDLRdxOWZGSrSLPUxnKvblFTCSoewSXrzut230qj720FLrQWGSH6qf/r
fWH6l08QK0xbAzbdhq3dF+3Pm0XZ+D5uEGT7mTuI3BT4dOE7+2fDvDSX4Rhu54Cz
bzzHTKeRuKrq3IRZ3L1SmRlQX+8EJx/aj3WnHkR6MJBFA0+wnvkGNTmdBpXC9i7n
QNJ4X76fLIxOnL0x2dN4Ov3qwFPKHb9ibSZ8VIcoEI4N2+vfm/A481xGHr/tztcK
RoSWoY7wWx7mMq/ptpmGKPiqbkmDfqZDZdVdAETBuhh7RGOCYIHmriZ5iFTLSHvE
DnT7qHzxQoDLsWiZZz6kHuQxjdxFXvOazE94fYMfOg14TEbhi7ttrDE4K04xt0la
tzm9PM022skST1WYQFpbPUDFgc99SMhbMrCDvaD08S1jwdF+GctV+MgFDECW/y+Q
dL9OULvYK9n+8Yz7TlRtol/l0lsUjbe32VFViW8MmdIalcgiKGE/EeG+jfZIoLO0
MePjehBQ2cbliEZGgmsF9bu+ZzNj9UHkkY2t/rroclKJXyqvduWZG16yjokY4c5U
8rESSva5g8HqYI6yX8YNsJ1fvfQPe3QJzw9ugHs1b+khAurvYhmdrP8eLDXD35T+
LS9Arjlvujr8/wPpy2qYY9ids4tR3Lebr0WGi3Qv5GJJhr6vrI9CkGNt7InCI2s/
t2q1yMA0p7dEnOl4mHtsGFq7KRkMwzUrRIxbDu4pHhN9+dMNypji8AImmOIrHtCc
ynwWBeifOgLOjWToFmyvAPkjxKMyoIYs/mfXePsRBBF6thBzmh20hJDYTD+gLCY9
UbwoUZ75ojPatUYEOoFkmVQEuKvRQ4OYgbuubYlB/VqF8FUYadRez2kAHhdNzdPO
UaxdX41tv8sl2g7chaVaBHWYpTHvPh+DKwhNWR5V/Ze3KaV9ybWS6IQhaYErWv27
bj3z+0/FdXD7scEjNF27m+NdgXOSGuzb5qKDNjzQWs+8LRaarj8uAIoiU8UZ2EY/
lUYoPa8UOMsTnYLFrNlyTu9I8E7yi/0f0DugwNF7lst9u03md2pDJZsIRmR2b2UG
iAiXUWVtqQsH4aXJe0fYpMX98SkMHlvPfVJkjPJ4EFom9lXuJtsQe4HIaxaLXZrp
3dMBwhXSM4feARDvYU4/NhpXyJf3BkD2GxZOsHXwbgiMo5IFq2tpxGhfhD9qBT9f
b0jxTHk+/hyVbfWLC9JSFBqZR+a7uzfMFjBUmrPQvUS8cb8fL9Bgpy978s73dU/E
AibIp6Q1FoAeVKKmbS2WAPy1FCdXqWc5jzEDFXWG2sKaLLmwqElqUid7Tm04rKxn
vCfs5eqiU9J6wsch3GJtpVNW43QszgK8ApHbbZJ8R+mD8buDiMfZfvZ9T4/HyfSc
4qRZIcWPFh9UDBmVefRh53zxA2CxuE8d7gtRLtwXGLyA07Ut+x+04vEgzFtECiZ0
+l6ilsWOB868nwUCTBkwrX7IUPb6SnlrwHNbhHP99178P2EZ/5sYxB/PEPnPhq9L
+lS+xdb4WqFe1iwUy68xqhfzvHP2kV/M2xr2wZX84djoLemaFDEq1OlUZmRfMUJb
mMNN71rGohVr0Z3QzguHNm70DwO2BgoMz/dVO/FmINdNQjzm1zYKoEXY5pReoD6b
300bCzy38/WWbHwxFYsN/j9WS/ZUP7ZkIsibunO4KXmGj1oyTedQVnLfSCI1wW/9
ndEBg6cac264CVj0hESdqA2DOQq1awK0SbrY7bF5ZWjYdhFx78/8xd4Nmj/vgfdk
Vg1MHzZUoB+JPzry6hV3j89uoazj4h6RmXGvvvIe5jEB/vnRHNrednXkhctzRBRb
ypHrmCGeha7brrAZ8CHF4xMWiYleL+3pQH6NjvOhAFiXuRfauS/XH/b7F61XTHjo
hq5kuW8mlyHrdsmkJ706p1pw2Cup/mWqhw+pGD+x2z1j5mqs85I+RwCqA0Gpxts1
zoDzPt/jKjCoVpcPRw9ks4YJTG2wq/AXr3gZ3emRoIFs7uqKS/ZMJ9Y3Et+Mii1g
o3pjxYE7xYiHzLACOr9zqWwEH3ZtmSmjKN33PqAR3EgAx0e7tOcsDnYkYfDu5Tna
zJOws5dFqGbjrV8kF8M+Vazvc203Yx6h+TVvhc2/Bp98gG6loWWI3qcSBatV/+Ru
oueoXXlixfovo023UeA2+6mkFSXbeLYy30Lb/O3qZUXthkGdjeIeJB4a623kB/LF
6hJpu1lm5R6Q2mEOUZJ3h5IPZrxALPSTPTFE5cY1PHSx2+EGkiVLSKmq5LyVhrvF
N0iywTCGGuxInjA/Zz9/6dJ9gr2jiwRDhKRNXOZAq1VDR1Yn9fVPHIvsvbgZxUU4
v8ksr4ph9lcnnPFI9PRQLC4zMDYat1Pr65p8hFuPPknF3PNvGuJaQZe5aZdA9Duq
HJRvlCMmKdKYIqdLHwo0LFOkt+juhaRqOC6JmcmdfafYzPBneAtvxd1HMLnq8ukg
cbgpd/lrKHuT/uHj96iwp3MpDtAnjOHYrAhKAyYQ2/b0mG1VFjRQOcdRk1Q9BXRO
XdPOG2ge6vnCwM33xnv/yABkIuHPMwXfvVCXleWAbwO7S+EOtuncuQHkvdpJ/AFD
pw3K29ExXVvfp0P/J3ePblOg4Y8eYl1fhGLHXbpzZJGQk13uPJe3x5oYkqBiFn6W
pmYk7Cl5WCKsUTSGVYikrqyATopZNcvge0L7mmRY5+FoVJRfhaqlYNOFFUO2xn+g
e5xkFJHOX5p31jHcovXatY4ZIyBo2UOwPtRh72Z++RXmVvciURH+fBDiNqe9JOEh
CAQAQK/6saxB7BLiGoB4PMLUP3lc7dMEondR5lc3jzlyv1FjLx4OkgL/uqHw2dh8
Fmgd0YBzzbwtD+W0WrLiROPnrxlwxKGC0JQlxJN/YLvUStgrFSLA+ehsj/mgdVNY
4SVYMFIsaB1F9zGv2L5jNKee2mBWMhw/bYTfizc3rXVR9AThq8SuOn41rIEBcYM8
imeMaM5PD77FV8uDvfJYdXFv+bCMGc11Jf+7X4LIYndbxXDMXTkQqS8owd1oq55+
Rww+cQrNfeQznCuGjFznD9xaee1sdhIP1GgJS3Cgojyndqto/vG4+OPj0GJUl3Wi
enbrTqwhncRVc3Ry9fzEeQ==
`protect END_PROTECTED
