`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
huNmu3IOLspBLwBAja13+Os13K3xpshjug2D/RUY49HwYs9AkO/B1Bzlcq4wZKgW
8AHlucvg6tk2dHRCHM/RhDdBZtCWAE7O/K49gNbw3s2NXqv7SCQst4zCmTQpl0xt
vNQjXAgE5KXCX8pErrbgBJfY3sXcAMAoBI1rbszLbPGoaDQ3TRZnWLppJNmOC3z3
5jgk2GhSCT5avdglWyKd2GNFbwDZ88FsZv41IGLoR3w3J82ohd8PR9SyzLv5Dm5o
IrcINx/bPFZaixbAuCZX7xe1aB65WtD8EDxs6UsL5KTxaYGLZL6c/aWohixtJs/b
cRH/TtbZWcsFXz0PEge5ohLMmzuaccW+aKUIC48xXwKSMqM3TFu21/8jRozrKIcd
LEp3wCqk9we670q1DynIdwUCEEt73Q5rqT485W7YBFJr0/csFwbU6L9nkh0gebH5
fmEITpNeTNkqW98lqSc24eLTAmClFbCbQ52KaEqYAtneQpQndNBpfPaYYPNr4vID
GU0DVVxBSQEObJPUbv5+6eyr+V+fb9F9zb6NBTsTrqf4L/XFRFVnycv7Hzi0CsUN
Bk/3jCw2/cmD2Oyx+4fAE78RzqHzh9afW5HEqlo1q3jbt/mJiC5bRJ4BE9K9haDk
6eDJ+5xri3Yo+oWPGWKsYFDXJpc6wc7xyBpFgWK7khCwIUd/Q1z9P3caXmJmJpxt
zgOib9j5zB2FO6yNmr3J9RsUESsVbfH2a5IlNohOW2l2h+BpBT3uCH7RWbir+YTL
Y2JpUN2v+jyD6iC6ItKHpZspd2EWqYATMLnsG5c5wf2iZ+04gCO4tQVmnSqKSmID
gQEdKiCLbMn8Q+rD6hlfVeQZ7Mdqxjbl7gDhiiVXEiFeJbJslMf48x41Va9nEOqE
6tBwDdiLsi+mNM7BUetjrfv+Jx96eZcogRBcrxzc4ZIacsIYfScHYy5J+XvsDH/p
MFEfcw33vQC1xk7qA6Vw5i81U2FKbNqQ60SA8eotOkqtpwPjoDDjL+kQiR5vik3g
oE+fU4J7qtPDWUEZSK+EXLbZDsEyEoQ8UCYKWluaWW6+AWJ8nXIRaQYO+bY4AIBc
iAPofb5dWSzheUJAQag9MQxg8mqR9WhK8bEgXXncBZ/E8UaexPlniRDWPk1yC8W4
wFn4zVA52WV7j1/iasAhLjiLGcRXy3FSuz9PaHrImA7If/djgESPzkbhyBCr/hct
/MVa6M1nDOdW/jOeuUVIigaV/yLRpuYy7KEJxD3M/YWjwdYtIORra3M+lH2F6wWe
gKQx5T7nm3Hc/mfmxk11bKFDgXHoGhe26PNlbbp6AjQJA5soP5CiJ8EC72jOK94e
c3qCcj1iNGq/tfyzTe0iNscQKY4NdY/kBBtRs82aldv6Kvn2xT0UsxiZKtAIRJQQ
G1ef50xmyFTf33CZXExLagIBPLjcj3yEJuQuZu85/Ol35FSeL6lFcjMZ1vpSFM0w
`protect END_PROTECTED
