`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0oM37WF1bB1VVlUz1qZ9VQi5b4zcTYP26iqfanFAM0G0PqeDtypls6ZaIBfI0Nfg
Vb8dWnDx4kRAYqQNVOgSQRMvIBGZGe2lQwiXSY/Ch2IuraTLT5So3cMg5MH5QmOH
doB1iewink/mkyYiDtCrNZnYnS3RcOcimjwr1imYnmHQTS53obQdqGtVF2CoKyM/
2jRNy+f9NBTtOXsN6hFHwwlpIGUKZxfVogMS6IT5Ze6ASHb2czDEW636D6fyNRHE
ue1fVKWhwkckMiFlBg9YYf2e38c0HppaX+35ZZTCD8QcrOTKXhyWxdgncKGtngSa
Q7WOK7qD7d6Kh3hvkEyLtiIqYS8t3f8udb2Nk+jJaZaieP5befIYvCLKA5nxyX6t
Q/bMsUl465XteCT/yi/62ars6+Jiw2iag5ryRhz8LYa55EM9H3mwX3S8IsEEhb71
hJAobM8tNGB4ywMsZ+nWl7h/cfdyzaTMTFDpkY8rTC7dDdHcuCkMFsyYtgrHuIvU
rjYaOtpkNyPVJaaurV0nJir5uypZyY1yb+nfZWzwWn9yhEGwM9xi0mhuh2k/owGc
`protect END_PROTECTED
