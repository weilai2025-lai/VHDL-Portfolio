`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UO23E/sPRvagwmnLCDPljgAQAbSZ+mVXgffmooVXPoh2f8dJRSLpEciOW6IF83O2
rVpp30a6po677W+TeZhEBVJCw44iSeo6RKb7bkPxDzhiJEjoCdkJAhsGkyohwQ3M
tG4lbe5ZIknaK7l9XYThW9nZK8GJRMo+RmCt/o3DKXZguROCnNfYYJILQkV5U9kt
dJ5YyU8c03XgwHb/+ot3InSeSTzmE1N+aFXRzgpUfQaNMlGMsdGgpyLBlQKzP+64
22jt2YXGGCn1F88K1hWdzFI2fiGZE6Zp4bjGaad0DECv6OqyIH9Ucb+V/nnqnxWt
7i3VATVnKFLwXBC6oAJ67KIvBM+vd3gTpttL2fUTbq5DpAneiMS0EbK9lRkhjk4E
iZTUusYyqsouxQnfoALjUMk4bvT68p2p5A1Rzf0zJ3HewW/4rDCgaegWi8DUoAwr
OMis2cWo7c77wsae5+fEjxlEmbOg6L/s6Fw3yrZ9UPNWnJZyBGRdxlXk7xwp2onz
HT2OCToLTn79Y34qJD7d4u3/Z+KTMblOEl//53nEWZsB5TRVIBWSg+WMjORN5gof
JPFpSDkxa1/OwHggpwnmYqmO1ujpRZKiH2J1Q2JL0yPpqfG5X9Lc91358N7uxIwr
6wmshLisSQX16CHDtfJv2w==
`protect END_PROTECTED
