`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XhfjPek5cszy/zW3KO9uVqgx1+XJgsAdgI7KpYAOBJVt2fLaz//9ctmzqLz43uDd
iN8y7kuIpFpziZCkgeHaqER5OQWoDqjFId6dNxeadctwiNmtvqPtWLaU9cWcH+Ka
9vRJmbeSItCemPxXki31QqxVZu4cKwt/eJGxeuyL9aTajR7r3rh9oeu3O6uuLFgT
g9FNol0AaouW2xbGhJ3GjPv/jpEwqE9lHYs8Qn9bi6H6elxkGeyfCYP5JvAeN2cT
JloQ3Unuczp3yBjCS6oEjiqDH0qKKtjFV8UuvwrOPiHIUcdxjAAoKZAV76DRyuQJ
0Auz8daUrPY5UjtwJgNXh7eKHMuCUvu/DaSuBnNn38ezq4EnZX4bLF4p7MsUQtFG
XTJF2RIWWYqHC5jS11Mqg0QeYvadw8vUP8EfI2hBzdvOohgU5pep7GHUqBoDmLkh
mw583bQ5jdlQbX2ntMeyaae34UXxsUEXrGwqr0Lewpc=
`protect END_PROTECTED
