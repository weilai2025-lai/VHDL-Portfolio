`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7woddbsBUaBolW8of7if8BdM5KrBSHPDCfsUQKAdF/FXF+SXRtOvAEhkZK032SVE
5btei3CeFG8aAxmyw6lhScg8MB3En7zJtLmrxqSCEV045DMuN01ajIKz+zY+4erJ
EDRS1fVYQv95cHCLD13464MvL71JxxkPGun3LdlPdHQ9M+JmkoYzG9moMMEPIiEb
OKL+icF0IUUAHBpENtEibD6GPSdfuJl+IXTOBogSJmNuFFv40hZdQ2RKTkHuOzyp
1Ek048SUulUnmak86cEnupaBMznbCMD92Y2fJHGutARw2nsdNvjgcloVQH/y/+Co
l+i038Wg/urR35C5G2noWkTE1SW4xT5IQ8FzxUyd+kcznpzibcBbOeQ6g1W2rTqK
/VorQmDcRhfXAtiZl9iuzQSPXk58Ff+3PgcNTSNha8TIXV9A05SjlKKdFXwDLZM+
aExrq6LTDF4oes4iXGaitJoKtctJ97S0tyr+qkc0fJT/3LmdoYUF2u/UEULpL/Ye
Q2VFYnCO+idhzq5SiQ0kuvJAsPqa8lQSYNeBpLKT4+HdvCpLFSKVxq9bCLzBb7xl
cVl1ZU2tPlBnxQm60o+xWMIHNqBWP9Di+6sB41dpEnjVErDyjOL6/XpUOJj3W5XB
uVy97XPADTdSHRV+bwxSYoYRFuE186ypiTn0d3KGxfeJiyHhXgSL8iJunFET7CWH
8qtBfBA6GFjNPtGfb230psXbD7NnSdPa6bmmnevfI5ksLfT+t9Uz/Gc1JndUDpcZ
RI5uW5+87uFCnMMlVYrV81ZfXC1YO+UeOnBmTSHgpZokI5uee5Gld4qiap8KJTiQ
TmDtLPDPEhNooMloC2tgs8BEgzM1nzgbHi8sE4lraQS2PCAelI7/P8rDoguXwu1V
j32v212EgxDpCcqtzSete8eotd75I6UKsgPVxfgTVrbjUqkMvVt5MoCokE5pisFO
2xtpBxXgivaO0aO4ph4z59Qv1CcluJeAA73mlk5YMDVD0LiarBOAaDVzmqRg732K
ucatkldrpT8spXM7SFejWcqF1/iAAt0dw+VPBJPPirPdMrMNFZTVy/MUhWodY+pQ
ylMh45zNtpXOfvi37lH8JBvn1TiDPzRQkVTI0zQ9abp1GEbVsV0Mrt+pOPDBW4KA
aBUA4/v+ZC3MSY8P8W9SQAY1EpzDOVc736dupF/JbomXKjX6VDztAknP020tMQwf
mtmxNf5t3HG7Y/3OPTOWOee7755IIiKmlDM8jV1k+XcXoTvGRDRpZQVjYEKfLLHr
FmoSkdMQNNLl3aga771BwGMttd1DnEU4JHGhGXwmYxxWdJ6uxYFpVI1oZ4XJX2az
IXb1SbLZ4I4Yj/7JIt0UbiM7u6k91KbB5A/TT99RqQeqLQKhZXcorW+nBxKxAuOA
S6KYhlq5Qhq9qr3diiVlalOrlotFM6lCFVBqolsOB/ehZLmlBXD2MfU4xZrw1FKi
M0SzOUByNFZXXQPkHGE7NsGQGIpBQJtSqP2yEra5xu9GZjaIm13EqlAxCuTNJErG
LvdJsq1a279lY+wkP5kxpnpvtksjtNKGuDRhDABw5M3NsF0NNyaH4DiQlU7s7hnv
rF8eWh3hvRDSGg3eK012kGtfITlWsFckqyrMPO59pi5TVFKLtmTZyY+OZzDEawHX
NygfdvjXe+u3gEaFu3LSLnaQXJeFkKVe+yL+4YVAAL2I+3RjvqdajP453UfA8g9N
xzHJ4i1P3DfOgRVyQF8zJm+kymfEWC/92VPMo/NE8wHGRhWwqbQriEojbuEj7Z7R
5svWcoehZXUJRUSJYMHGwFa8oITy3i5n5X8P0OkZR3jQDDoppC0oB+D9KvE4u3Pk
tOwZqrgMyDpSxtLCXOQsT5MScoIy7tGJni0OhnUFaVYqenp8uzw13j06MBqhkDDC
7QxJoYYPrGpK+gJkdRB2FV/LBrW+JLCFN8DFJZDeRWoB5WPGGXtjDHXTeA0WfbOt
JzSk4XvkcVSVbUZtyrQLROvwKvmNJoRdLBRoOF8OXpuFvhCy/mAYXzGqy46P4yKT
QL/KctswppwHPf3xQHvycjLUwvBqVs1uxPiBr2lbweLIsvQw51pcAKL2Ah0ndMrZ
uhkaPxYEjG8FE+lbm5Yax+bKUDfNtHfqeSa2NBVppWRRmouxa1QVucH2nS2SaBbX
/HUBD2phNgpqQ2JAIIr+863TXVtkiC2O5oO5erNzYlQl+VaLMFuzFkex6iuZfUPW
Cg3I60G+UYIuT9GmuY9uZmb89A4daEjYQCquP4QlvIQ6GbqF6wCC6Yxs3ZV1Hw/E
nVEzj6qBXSmTWOLssOX/Zn1MEnRNt08mDjdtRrA0lq13pWZQD29TC1uxsb1jG74F
3gNynRBjgF66chZRiOkmVMky7Yqk29Ir9gXOGQtBw+X4Cq5g8WYCuqjjQUuwV+MG
pB2kHldfAZuCr8F9E0NSrlJQIkrdCJIfhR73dUKhS1s9INCoaQYc495TMxBahoGn
myWO4nKUOD6wvwDbDR/D6jxQwcXS2rfvphjPmnit3VGWOtO/b3SgO8TqqIkNCpfu
bn03i4qVJ0GFF4DJzLHF7glVKohi15VGs9VcOrIoPZ7NX/UhK4q8uiTNig2dAvbx
R5XAKc4TmcIeA3j4IcHgBFymoQbUsC5gubf7cpYNuT/I39/DLpqR2sh4oKqxaKwL
IFrhCPOJTCY8DLSreK4UHCfQb/7FB/IVJjelwlDACf8Tsn7BJQ3FTX6sHmXNdBg6
5l46WO9EqhTzyhUNn1p6fh5zKxDKJo4P9lI8lypuUSYJU5fq9+qqKcJeYN/rvyB5
wYFBHzIF2lP/zb3jrMgKqr2OU6e/7Zij6uKhzNFCbUADo/Rs043cEP/8w55m+C6p
2btu96yJfyLEgn2obSfu5ujK1e1TTz2R8wCudUeYwZVAyBAOOe4J8xU8xukmrNAT
UgDY/DtyXqhxU+SPp+3n+kyooInw7A2MBfTba2ks4s40Ipf3mOOWmYt+1yqabsiV
Z/59JVHVlUBp54j/UukKvMTBo4CgzOo2NIMexAUIbI3wsI/hPFaWss4YbPzl2ndY
/CRXU6ZMiPqJqWOzXpfbn09QKkpJW70qTKwzRLHqpnlwWveTKUdi0k/O09zmXxDO
76DWlNcmnR//9NoENfm/afZBIwoWS/WKwsbMElYMb0JM9PAZrfCZ9CuFewM63V2k
9GQCxnstxzTum/5p3j9o7Rc0UZAKoFslPITMhK+YBqqSGeVzzqCflzOUAq8gsyxe
uNfKboTmxcLTVFgEVFqqvK6rkU5oe71xXfHlMPEHiKnTVGgpG3ZAUG5T1NNhWY3R
bhvt5nLQSNkAbMGvVbcmSYWLcoRCEeaU26ppbJNe2HWDiTYFB/jXAHmLZ2H8CzYv
f3M8FM7AScKgWmY7oYHSJPWChmjj3BoIsU8TTY13+d0PJhKoEJ7UWyyeLGSZzl1h
QIm+CkErz8gFTL6wq2SDtDvjRvhbKj1bilkvrHqEIg1DqvCEItf9mE0p3p6Le5hk
OpGyV2ELrAdvA9n0W8xlOc4eTeAkzRb3iAF3LQyTfq4aLcDt+e+t0/hKIRFjg3A0
szE7FvqNXcbE/vhiTw3lSCStgo8055wG5szUnoG1OQDMrFGE7o6GOIp1/urf+Igj
G0sFhJhtscozDgCPtWiHMXxKEJMeigTOIGRuQRj+oRSQZzTvz/EvW9bYU3I8CtZN
CBniT0RIMyGPFkGgG03Ff51U9sPK1aYHwVBcZa1Xgj7XLYkeBXOfxJBTCr4z5T4x
tHFxGfyJkSAgi4bEyp9XyzgChhVMl+3vV2DXd4SwYGQXHQb6iq8i0YQnsX++N3jc
AOlPdz56upYF1VMaO7X029fizFu5qrVbavkBPnrWxy4MnYVakNeqQD5LHBZtp+iR
8poQIfQSrEguk7+FJYU/+8hY1epcDOUvWckOf6mVX7KEIEHMcNUJ6a/cEpnVhkW0
5Cb7GS9waM3WDIOjsfJAZ9eJTNdLV1kGppdsjEKCSNQXvrtJkBKCXc42LvNbEmx2
BlNAmnL7OiY146FGxOWiiwvIP9TdeSqTGXd69bWZFA/Q9TbJa3260KqRLTJpQ9JX
IaQOp06XSIafhaM8ye9vuOhWBHxlUfISjj7dRO70fLZ9w3Qmr/+EsbB9kX9ucb6d
SChzGnhwecA0IgM9JhJBQVdPLU+PXKSaVoKpuxV0lx7Ise6Hi/k54UJL4afyvnwW
8TMM5Jez/GkFjcxrZ8cMgScZiCXmK0sH0Cabs7mz7NnMtTtSAjHJls4MvXOxJIf3
y3kwZd7YE1tMopvEAo7L1x5Q0qFofuj1EAhMRy5y+24iYzN/heGjn6coVbMPgLVh
ukTJ8x4JMc+9/1ZHSMpo4xcPcKinN8lAe9LXS/Fy2PED85k4J4NRCnWnFK9qcfNn
2Bg2WEd+pMmIIzZNlo+AQyKGcjG74ZxQ7FWjDsMI+jgk3yYkfsc7mR9/IRAjt5iX
waxxlpB7d1zkya4r+iPgT9aUUiHBwzJZuooDF3I0ZFpK/tmd04eDWR82VcNXkWrf
au/akHlM9WDPcf0CIIkz8ObKVS2SGaxj8jjRQJ+X3rI+jsRKx5nCyqMaCPBTe+A2
lBsvqSaMXYzRrp7XIzjS1zQ0aHZcuZJpF6wkcgM09Hf5GbYHWigNn1BD7rjZl27Y
LnzOnnCOv3+2tnb4TMUEYzE7SiUjsZ2eC/5/i9DDQCnXuJb5Y6UCGwue9WpIZxQl
B8Bou7nvI/6Mhsh3/qhPZkbmA+fFrk0KAjyjYjb1IsEIaVLrBmtMGbz0HFytnl7J
CGgq9WxrQrEsYYOrL0vltC+CBXDAoHoUnMJaMArLbg7ehOwKAlf+ig8Ablb27tvM
2kkNMvB6N9/MFx0srnOPEpVoVMQCCTaMmWM6FXwAmUpAxfKSA2696ufqaL/rJp4o
b2Hpd1gOlJHcktZVqkRVFz9HuPtf4fouA4RwWdgoP+7mz9DJeKyrG06TIhQP41qf
IR1JbdmhcCY1OtV3mR6mDz6f4PGSu1HzCrwECfUIrtRoTwfmbWwnuIJfmJrJuYaU
WPCQEeWuVL9duXeXDFk3mJd6y1qPnHNepCrsCaBRjAXDUL12MGo+kFJZsKYIotPN
52Hu1bDVEYhfBQArHZi0PzTlYsCeXEE9UhB9+ASdbH8DMLXzP7XwPX++ptM2icOc
naHojni+tvapqVcl4lxgPwmiXH+2NBkrxCKcRLQsqArZxeSbrI1oja7bRsC32Yn9
gL0ovHYVnT0rogmvVgAdXKiyk1r1lvKa4WaxZAyT5dbLkGNGyzJqjE19dWYxJZxY
xdVt8Ux7vR8qiv+OaYV7kkmg9a/0eJsg/NDPwQOK+ggIfo1uGXdDLlaeICIKQcvU
9ytF8fW8T2X6JuMPpXwiUGrFV5fAirkzjJoaBya+4QkTxHVMKtNV6S9Un21M7MyE
93FgIIpLivTpJcqACFnZbx1OMzOWvAUT8icQSSOmt4WMoIYdf+1twJl3UKn9P6nx
NdLrPHXAJzDMDotnudP/jI+byerNK6aNgv8aQ+ZsjI0+4Ph/V8WDcLSdLE773pXm
/lxjGO8dSRBU90HH95+ZII7n0n5kpEl2DDzyV4NSPns+U85VDuB/gtd33DWOhzUC
q8JdNXhh12mrn7D3GL4siYyDo82P3pDSzWSel3vTe40wlrpVX9WZtXgEZ5+h4knL
9nRASZ99AY70z6Ub/mQNPRfVR8RmO4lREt0zf/NrXSjBklThmTWcAi4UwbegvncP
Z6l46G7mje3AegkvDYy9V79SiN7y/5M9r7KnojUQznJCTBB7XsKehhKHtAglV7tX
5uzs2uy1zZ0JWflrJPIbVhPNToHffZ+3WtW3dqTHXGopUIjZPRacyj5Y11nrHHnq
7qRVhPCarRKe5sX6jByfkYYUuXe7aAuUMhtM74jhtLP5k14UWJdnhFGhkxNFbdDo
9JJCsDQrw4VC+Bj4rcQBuu6LnhwmT3u4Jeoc319qPFICGxG2P5/4p7RD588M7wYs
I4tBkpqhVkpokCcPNhe+uTfg6Yh85GCunCyRWqk81CthnV277hN8uRmrWpCdhOQm
bXbBhNHK5AT/nQHzSEEMHopNMClmJFHo3CFP/s9Vtift86JDcCU13BVyPOb88TYY
xxgfD+TrF+MZMALPrhK6CqNWUIyp0Y0oBr79DoavUdpjNC9FCag55SauS9BQcrfx
0i1OUMiBYHvg21jv1TiVr2pzrMBZoGxVWCNYKRQDH7RbCn98nHQV2AwfI9fgx8Sh
R1qk3ae8939+h0J8tn1B+7GBjAqU81URxRwxqOwConOrSM2Ttw4k3WwadbMs1fce
FFuMWisQ7RFnVKtj0jvFGh3JR+v3W6MdOI1UBp5rcqKOTYDA3019ZKEuRiCrPmbP
c0Nsr9BhKnrRLnWTVmYviczCvLq6dhDLTXmJceUmNqROonI0ahkiumu8e4+x5x5+
cm7opK7ToryDzE85kRLCEPSKSb9sXjfvzbrNNlTQfr2yTwK4JcVnwCvpZEX6qx+4
k3qHo61+4aaxxjWFWzKPM+IAs4Qp0lWkjck19HKM3SU7v8CFJHxKdPCjEcfh4Dy9
ShrziNEpok8uL5sLXhvJzps7AAw7t1aKGpdk8Jse7J4ZBZEEfLpSc+A/b3CCHgip
SGV5ZC1eIVhWbm8Eb08e7U4t55a/LQm3X4aLV91mSlKiTWZCBsboDskotN/xwaIf
id+4rBnSaB6VHYBh768nHwKgnCN+4ci1bgkKyzW7CbavUu7yMovQOLGLEwVsbpVh
2cGvF3dYVSDqnv6cEtGkSaXi/FHdVp5pOh39M6IJCrtxOJ1H3ioacSF7GF4KyzNR
bTTZUCw7PjHCS1j9FQ0kojmlYsBxykjR6fp4Wnm7orSFAsL6GpfZKV7zxqB3k46E
dI28ojbRppALKU4bfBsIxQ+pqpm0Y9QUAW8WNtt/sZRlzyHyyJ5LAQP7tvD2/p3O
1qgvZ6WMqRNsnwTdMxzlFpWtt1N2dvZrpx7RjtjiPEyN17QrmEQAMw4tRKsVE8yd
9rQ48dLCwEMI0/7rWmkvCpxXYrCzoLZpX0dFc6VZtKlBqPKGiRcXeD0G1buuOPV9
oYc2nal8D9Md3cRaBmuRrrR2SuuCTW7dWKWvzDL3jppuKSkdvdeupU0aSB3ZepXM
w4gDvbx5ZUmhIWATUCAM1LXZqMWEV6RsXb/I25g4l1v5VnDTDeBRLS84XDj0b56K
Fo0VwigdpXbzF/MXsyalU4JJVCjl5sRYamFJf9Gx2HiHO4T97yMsl26EAJvVXBNc
jwYhwri48rRGJyhYi5o0RXKW5a8NfcZ16w97Ff7JfPFuQAmJEdtKysNYFFXQQPNx
iTtN8HcUlshiZKUBrFrciz0MPhGhz2ex2wrDucxH+hUU8ZdvG9BLgGI2DlHuy8jI
uOKjLnnJdk3pvsFeq731sv9qgrBLD2NXwyEWa0NIEUxcQS6Tn3uZ80FSxfS0hYP7
thl2Jd8CdFUmENffiqW9tdxlNaC8AdrVvyAkmgiagGsZnc2PgHM9ZhkGUd3aF5qU
yGifxQKwEDjR4qz6V6OlYPeG+VxTTKvT0NiF0fXuzceuDwiAKHojdq4dY7BeEtJH
FD+oAoVOL2ZqXRMowmuYa/VhvtoiSJjXcBvcU7aMpm79FobJ6TLN+fbjiE/TUFn/
JCeriFjwY+VWK21HRE0ATAy5skAunRSDOUDPtPBwmz/PCdXgWBCsRLjeOEeKVUiu
JoGvL/0e8rEVAJ1uZgl6Vm6bwOrDZnFkNcROfCL5MCe0yXV7ENyyHsWk706oP7XQ
uP6L+Uo36WOfU3PUQ3hImoBjpxEQb6Wk6Q7Xc2ql6BwdsEmvmLdwQyJaT3SjGTcO
QwAWtxfP+8yjoS88t6HvVkvCe9NBluyfM2EkRJ4AvN83hBskk6HGQsTsMbe2k5+i
YPILPvM1j85TzY8ZrV9qCN5gU47muW4CP3HLQfWE7KfRXl95MEFFAG0a1eU5bs+E
odZGpnIy8ZSWXUzMj2vLKxpqf5n/2aS4rHTT/de5x3eRWI31excC9tFiO80PeO00
MiCo9aNul6L6Mn5eyXxpztDFW5W2moopS2EqKnPQ6l6+RC2MNA4pUjePMdkgkEO2
gkhxZ2WosCN5VBZ09r8hvLzO4phUSSVBcRcn0oWbnY9iExWHysPujKu7uzCQVQMf
xf5hWI8Kv3N4JlFHMl4/XnxAvXDfbVYnty6UU9pVR0TTVvKDfj3IQ8XQMofDL05n
toPEq/RJoQsh5CSC4tRE6NBbF2RSgaBkSR3FLOQl33RvhUVZM6iodmgiX2Mj8A1V
ZMbMvNcZqzU+vgOHWyskJ/mQfKjThm9P/14PqRYoE03QBp9cG9ZVemItDkyNQWlB
0pGiV91xLl1t/C4yo8ugfZ42RLZd+2QgjV4iuaXPQD/2f+3nqF2uUfLo6YNuXIva
PH1yX9PJLsgNhmGaWlAPPgtslWB2eV2sZwfl6nqCohy/XMpxQYbeAUdMtPUz3fdu
PQKq4uklTCgOLPLHWKxk5eT0Zanr7A3+C+CE9x7FGD9LjFScw0OhGmQNOMsJpgHI
+HBhpQIAp3rtr9iPgyrIijfiO4RL/oLHpLRf4/ytFpj7L1HJmfjqbu8ikgzYsweg
OyBTGuwUXOtK/qNcg5uzPw0hdyQMFahNhZyhzedbwGpEApnk1mI8wqa2GvwZbM9T
NKeoXOG55oMTBb3xnEANAfaLvCPg4+luHxN0/V+kM3GBDvfp7U12WUNBgdcai9ze
utAgKSSaW8T8Ez6otGmthL0HDLq6I4S4KW3saX+MYwXn6I1fxhpBdyBMhjGgbEIP
BJgtHAKzMyVquD/dFOHPWA+NMsLM5RMSDnW6HTz9fqNsWyVVS08vCFwGvm3BWSjx
YD+Pa8GXakQ1QVk5nwAl0rOgIWs+4Gd7xksjh/NRt4lMiDSqOv07tNE2u7J/HHPa
WojO5P1l69pDRn++ZknZ+G5GKY9o7Xp48sWra65BRmt4zt6iiSZ4Q9012taycFOm
nmTBvuycP74MYNp2AhEnnU03jnnJTeYbI0wrhUBY18+dU8FVCPJLekbe2LEjvwv9
4AiN1bXq3H/vjlraK3biX8vmcWGWAI69TG/l+7QYr3RkvB9wwy2jtAfT4UU2ihId
oLMDbWcBMqu1vl3vW6avFBZ0s4HXJO/yjiB39eOJsd1V+PGh+F5ADd4Kj659LVm4
hoMYLee1AeriXXrSO+K8s0GXzBny60Z+kze7O3TyPg3gIpwJ86/LJHjd5pdmf6F6
wgcNmdctyQQ970K29Rdw4s+Yi1Vs9Ye2Po5Gxo1fh59OUqKj3AnY5k3siulR6EjI
BcoTQbrVF58UHnObSLvtprOmrt+jfYlXuBVD5srNoxZpBbH4rZYpBVwClG2433fk
+GIPXdh09g6EENH47r0jp5U5SKIvJSHeA2Pp7zhXcPXGCS17YUAF+o8EvYC7Du4d
/hvkP3Ko5TMnguEdijiWa/eI6PTltcidwltfhiEWpIDpsqst3tmm2JnRlWjhPJjS
NNGu93dEx40tVmIvrhmAsxOdXNqyx5jqoZ0wCy0NDLzbF/lVwhcdvNck6AD7r3gq
vlNLfztyEImeDYu/EoHLdZpTXPtCBI2joAdYACKlVa6RLtUl0c/xW7DsgXzAQ16g
9ajVSzrINCBksNdPsZzQxUubwFjLbUxaoJJCYtB4sNGd2eUF16MaGP7RJERiZZCt
0gwVha6Okl/UE8LQBMbADhuMEDjJfME4aBEWNk9qg0IDfW3a2wiSuPXxdIfZ2CwS
UJddc3D1Eaeg5hZUegurraPunuQywVDHHmEaOaeoHrPEpMQctrBgGRaqndL1s9tB
bRTnv+1hkYCDg/OqkxJiU12ov5Np1W3MsdCT/zYigItWke47Ql4wbGLbNwT+Iaxk
o7NBArFBxgCiDDUDzOH+IjH0MSKH5Nx9My8XVi+CpQv723kREsJVDTD/kROvGKMf
pvXOAThhhHadgBDTfVHhXwwMHeVMLNUyUzhO3mGVS0kK5VFkwSbpFnF0bY9I/VdF
Fg/eK0CAAWzafACvQS12IZc6Oxo2oNUALcU7HspZ0gUsaUHreLjte6ajDr5ClCTb
ItL/Nkzkpki7J3T1B1G9wxz9qAItbAzK+YTVKmXSxNdIzrNEAX+NodKCvQEq5eWG
KqQhdc5Mq9Ud3EqEl5I7328TRftQec0MrmBQtC7A2NA5nx9rak9ArXXkTieb+ah6
WR0u0siWZvvEdbpav7ctfsgaYDbGWlqebt4RR0qrLsNy1iSmGvT3xxMnZHCxTwuj
hOzLcydE1Gr958dtr/1pR5sbf7wNvEXFuWvnEQI3Lqx9b1uQwVQXXuvbHNAOAQ2t
h4H5JSXcsjTI8DCsxqpSIH5dXrwmtzdJFTRCLshfEKVl9YbH1LLHhUhp8K74pTJa
zhgpqxdE4DVkZWO9AeXqto8vAWt5apFH/fjnybrSedNJUJYieA5KH58B/5t7b5jq
TKFRLDD4/3XehWV1lBsmK/vucJqNsauS+3z4jL2/u43BZWJK2Z7k5t2Z4gsanDw+
RUkuxR4HmlyAZeFxShpfCLd5DmEaOiCjI6HYdQfCfNbPUEkMDvTynr88/p5R/pp6
WmO3ta/nmGH6zkNGCXSMeKDNCIVHFKiRyPAhGW9nvOQJXArbQp2TkpqgEiQEy3tq
EZ03oFeIrXqdELDXJkibX1dST6ZqnwTynLcpdfx8LoYUCEJVgKQ/ce6ORWO2iMaX
mJvAInoaRiAZ8P2PlmlhY12zFUVRT5Ljdyg0jpimWLdsXKWotTyVR05EIyOlnuUk
pmTZXbnm/C9vy0EN78K2Z5rqFytELh5wkmeSekxAHevSIrI/Mr0FJWhtDe8+Zxiu
Olhj5ktzzR7c5oomuDYrYFnXu9uYQDTesMSxINSLr6SQfVkG6WQyhWUCtyUUtAp4
E7yXpAAVCB8PdDsobFo9pfA2HaYilJ31AvCSB4pS/FKIxA/bldeHKSY0NGJTZyeI
sH0Vz8qCTyxRFRMBlymKoNNtEt6GqkEEvbTAy0PmXOkXsBKKWIWqYxSI4ftp0q80
xfGj+O8v0C+TP7ZPd5mVAB7q45D0YiuO/GXL6VGUlHHY+qP9baKVS5g11uOg0p97
g9YyaCU8oSp8E9t+M+t/mvSZ1iv/EaO8PX+1r1QC7ZFugPhiDffd47702O3pEMiJ
DnXJ3AuW4ZLKjG62mZG6GRFOj5LJZKDRHU4xO/C1nMuBnui39LPCREsxzmi1ocQy
wvpZiit5MXkpUWkjeiXnMWRzTUHLt4M4y1ZNKO9KzWdeXATiM+uCPhKz6/S1cLO4
O0Tw1Z9aXofhEoVHr2WsojVVhONefeZSPRvdpkiSPBfNklypI9eYH5bfWntqujs4
9tMDYoBcDmyRHCpiUFl+HRPOCjoryTiK59CG8zn4X+Xigxn5E7P4sz5Yq0dXi/E4
TkymOuehXWXeROP7FmtRnPMuKRWrqOTcnnyUZX1MiP5tennBua7Psh+OA360h3ZI
bGGFZp3yTrjOQprcG4pG/tE//L2JdL16Y+aB2MFbghSTp+mA0dRluovOVAxiy9tt
g0CSV9IlwqK2iV9uu/dWKlGPgjD6valdIk8cEVWinGHuYgiYnYFA83D/OZkUOz9i
epB7ThxVqjFhzjNCt9ANu43Z0LPW77gETb81j7l7eTBhryotXvNF8xqiEwVFXBVS
brKVk9dkQeVcW3zL9yYsshv/bN4x79KIbu1whMKncI0B90ZvERxXVpxxHOSq6BKj
2blSBE2LYhHNMrtwtQhx7jvEcpKW7pQnv1d7YCWhNXcnStJ9HMZe7aVqyIK66ah0
WHg6IqIoh7mR6oqIhN7f25GcgXRJECKkQ1rsZE/XwTLJ1DutTDxTH1JgN+Z0dfKa
fkvyLHAAHTkC6YJNcQt0zYu3Yxn2AwWp371I/FsgSu408m8+la5/8sc4H55LYtix
tp+phV/CajTHfBm0iajlDwYBWAHGQSxBKQvK9E0haYwDC0lN3dXMeSPXFx1i5MgR
ZSX0z9mJLqBg2vUqlttRE0GypmunHExfI2dnjZj2iMd7cM+cxjHDyxY+BlO7bMPq
pIBfviKbjia9yObzsrwzZGVgnmdXTrZZdAmshtMN8ZQmrqy7VgW345UHwmTys4wO
+ijDwx0xqbJxAOmy/U7IzPQ8xIIkxrAkHaKJk8zteiOXRu3uSIJ8fQ9M0rInc+c2
XMjipNGRlwPB40LBbLOFGtOiCuZQKzaryRvz2aLRzOYpiZfidYNjG6lm2Bd8isFH
2NGiiQLPVtQVNVviaJFbuIuRMO1Ree6z6ra59yAyl//JpiZRMxtyn8m9kqxNbXzp
tlVOsWWPCDkg3NPMcTx1wDQBNfF6s8iI/9Mxj1nx2Z+oFBe8tWt8eQhJCZzsXMRn
StdXVJfjtX1pBZISUuhLXNjN621uOmKkpIr2yxjesZaNzeGZDadZDDmsgQn1aQar
e8E381BgtZ/K3Kp3OD+OfK9+7bzfFL4a+Ij9ivvE/D2QU9t1YuzDGG+b+CmSxgPa
Zp2YrLmqxk7AltLKjh9t9rnS01YMwNl83VGnBgdVO0wmSbD3KxJIY9j/IbsELm3W
tD0Vs4Q9YtD7Kd2eLXKo2XQkt4hLAAEpGgInOoIYVSnMXDoCpnCwKf1OzcHiN/E7
gEde9uI+zFg4seDG0B4GLK6cR+ZBI8e/e9evfKLyUCZX2A/GOBl5bvr0zFv4T2T1
y0GpI7u4G7h0fyh1YwXpdwTJpazpRHCzRmOIrW7U88EtZV+xPaCq7XFJWKwZmytj
u05wX+5kPet2xHNOQ46tz+xHN4XT9FyOwMnSE1uTJbM2DravF1vxiRyHEy7VvPgK
zchb6u/aOn6ATmJf0G31oUEKAnv5nco4gZsLtn0AqsTsKaVGP+pbcaazNjyLyZ0V
utELxsOEH5GDXqOItshM9rG1Y+RdM/wuzZhLbOEbQeNFd41dLuICqmNSLv7shg6Q
bhzO/VZuctL1hEpPQeNAZlmbEA25qc0wU+LCcIHSuByVteb0VPRy2gZy4M8E66xg
6c0JBEJxes5U2xE/DwCYUxN3i+92VqK9edAd2HYL+JbMmM1lPym7YsiL3D90c90R
ttl91Fb8fviZwI6mwbScuGnKrzozEwbf91FkH3Um3GCDZ7YUqE5+unfHCXWoPj58
pc1GliYlxTzT0fzoTwTtqLuybZikPOGnN2ftvFVyH6mCnSq/H4MAikRD+nVdyDXW
xEnv7MLTRfZBK6YEreKfyUR15mCtkQc19/paaVtQPG4I+NjdW3P5o/q/Y2Hw2GGu
EToZVwdjqi4S779n+hAufs91VhHAZK3TXwMisaTOXmtvTD6GRoBsKmQzUHxkwHGf
88WoVqI88y24UjUVkfnFSt+lN3i9OLc29VW9caGzetZK6e9LBCGz3RIyUUzfqilF
TtDIAuX5wDnzbhKmtlObjZanrpzXkxEA53KiPOmfCkTd8bryASCS/mVEEKMpIyqW
dKHN9x9pQPb88eWkC3918rioC6JWCqGlYlHx9Dfv7AmE25Fm3hLDdH2JktAdlgEB
Y2eCKNblA8eWSWyoigD5kQvquYh8UWMN+5P0BEkN6F1q+ylOh5oVFZu6ooDgOVJ4
coBRN2j2CEG6vABkD6D+gZ2vzHgkQRKLZOTyi8g3yIiL7XDV9RShv9AD6CFzSSMo
kaa6beoEEOik/aKQr3xN3vQHjKwJ/C0375V65ztKSMqgWsJgWPpu4UkYLJzLFSBe
ZjSEUI2MPEGNr9zHh1IuklwiIyoZnJRBPrRJSEIk792y51PPUIJ9FeNS7lWseNbL
t5yNLwAKsKwe4v0KnJTcmxxgQ1hmZJA24MUXsuwNayPFM0q3KqDeBSTvuIE50wTR
leqNYhXNBvWFeJVplFGP5nZ9+BC0gmqU6ZmFT16wZ9utOjnUC1qNipOqfk///oPi
VNy3PWnitzNaeIly493zL5Pyrf5GcLTGlOCRRASuvt09z9VRKt2oqfNV9syEKmgG
KeXXjniJhKlt5dzhB0SHiqPHAI3nZ9pX34rlZFIeHhbZuPB2hiP0Qq4B0t7qa7eh
myeQxFxptd/4+TeafwMks4JzwpBWNa3O/YrQbp9K3ckWN7GCUHBg8VvdZxpMFIME
o3/QEQKuntt7UgwvoB51Is6465Yh66FOHrfYT/u9RsyR1Oq5Bd0zUElpguG445BP
5OwR/zqISJ98aqQvUoXsWcFnK5gw9feuNAfIJo+QdNuwf48F4NaVGt33t4wnhW0v
qk+ja6IBqrTe1/L98W7CEMjh8FSU4vqdimJE4rWceqT8NFITyEFFtZxkNaXzkwJd
vAfCALAhl6pXL1arz/StEmY7dgp0Dre99G0BJxH/u5VGe/jo2LdHSyoJOxoxUhe1
DjsE+LN/zCifiyzRNLflVmCcaro9ap6hdTcK/3NZkx0b15vMBCEUMBSBjietv1ie
WTXrK8qHjdBw+nW91LcTAI1HTSbXeJ5j+Bf0QXFW5h9/hO3GDSh2S0N1RxvRuv9R
JRpN7hxUtEM2WWt+Z74WEpB4f4deONcZ1DOdAwCd02XIuQnbUsojLh5m3all0HuP
zswe3rbrcwTgpT0PLZTauT2eRzjChmFcoJ0kYVtYlqwcXLxCBawCbEgeGWb7cvE+
hjEpSatTRNoVNnEb7GF/0SemA/f7mdmC6pr/njava0hvORBh2NN0Bo3fnWPuvtxy
AUkSgo7n9dBJxP5uHghdXIfK+l7b1SDm+Sa6i5X0V0h7F86exEkwAayojdbsQads
bgtzJFbhhMXyr6xdx4EXy10p38Kd1X0Hiz082QYLh5VcNUbXLYL7VBfSQRhkScjC
j9+R0qTcJU1JtqpMnJLUQF3UbI1B4Sl8yXoFzPlovH+aW/UFO+Gzw9efww3u0czp
04WeT130wBF3MrsgZn/5qkmmsr8gMYaLFxApJi18UskpRRaBzGHN2gUI4hvKoA9S
Ywk9LFjXHE96ybexV38WaFXSGGd+BH4c3vyaZOJVcciRvni5q9BUNZl6j029QjJc
ec7+/6NXDcwpH44NTcOHkiohwJXea/RwSZaGKR2USmrmWZqyjJKWoRvuLfCO4q+V
1/qP6KkMCMgEhrItA+8EIZ8WCh472T/ZhHm4Y2kH1RxQ1DrkcRqoNsNJqkVIF2tk
2dzaMrtdvEh6SwLQ/l4TDxOjy7caCLNrl24QEdmQ9I6B9sz7WqVZ69J4S7TKW8DU
fDFIE2hAiiRoV6qGEp80PgOyMDktVDNW6sD4WeJ5KLlFofY5VD+k0+BimpajZ7dh
rVfqQrBFo/P/R0JbYopLK8XmaOSG2CqNxQiM88vfe9UeJZYhkRA+pZI/PNMbpQbv
m9A09QUrOKzkRdHw9vNKSY4bqfc9Jq+BrXw1Fze7Fd4jNSrCYZLOKCpafX6vr5xu
lyVWG6I02ALiApF5jdS58mBkYMgcjyuXJ0r8uc1xVI3unnDOr/PjG8PaDf+wuoNT
0Sg7YMBWkCrCoeuE8GMsZMGRtcIQ3RSI9VQ90unSBINR5K/zbFPpRQH+PsCTmaY8
jvqaO+YYp6XsiTd93luAcXZOKiWJ+ibUYJCfAjzRTu4T6xTgFq6pZUizhWMlItkr
HJRQ9fIZSS371S9+JQwxzWC0KhBBXt80nuPJsXmFZdkqArCKwYDRjWcgW0g8uh7h
3rklvr/Oixgj5K57ZwsziT+47wa3J17bhxQtvblNLv8ZigcD2e5COf0ooem2U1ok
6KG4pQxX3WzX7Mc3aQwRve7BYPFY6ARA4srDV9HlH5ezEI9dkeDhbIZNsSirKmSR
cDg/6KgJ+xAIB9BGXWgaKlyBrqaz5Usyw3c+U+MS0DI1jdIl152QmCaIzIAdh54e
24eRPp2AhjPFV/otLpKuPiwDC7cAtpNGA/4FZTVSDxLcMnnugu6tBQIUOjaDTLhu
6Ps5VwR4wI4PistGikZ1YFZTt+VLYgdjwaMxN3Gavpqd6/aqDiP8A7vAxnf6EjBp
bPA7GySEVIPM9nCILlTUVB9r//lPiu2ao9GC2aE0XpwAkZdw/yXSgzrY4Dn4eDSL
qob7/GEGt5mnLX4AS1IeyE/9u7Wo8vk7x0XRDKCK6bW7+dUSST13ITXqFGRGbYEm
XnS5R7QpeRH4fA/2tRUz/Hd0gIDFfoyI3kPHQUbB7R/Oncf9Pq1mT+0E0ehZKkC3
P3LcqnRukrAztchU3xwiJ+pYZvZ9sNwaI4CC5l7La0PMZ9rEkP2G9XO3/E7trsow
ntJmTgnlf0JQP5h078qdeC0ERVOMevH0XkIsjvc5+m/jLayTmYYLI0/d9JXGeswn
mCIgc9eBAA/mo1KGVgWoRir2daDY7j65gqRcTgorF/mYBJsD+fcqkTJ0vhI/4DTs
aNVpRtN4nZfuoIcQVgrDILO2iS6/WmUguRBSdr/aJ2YvDkOPkbA8hy7hdiVxi/EI
718WxxORUjnsD6JaItp7nLj3p00NUcBEVnOK+/R85aPlau7clWgJa+lKxaVBg9x8
Kc2xPOpx3lC+KYVBWsOZi98BdqEhpO1xWdgs/7Gs9A+LDQw55TqRBBEK/TaPJe70
MvUKsz3H8+rvFzUN5XIa5E9Xi7HWXRy705tx6V8mb9c7nMyKhu6YjXxaFhe/Lihw
5bKOHYqqWv/EWMeHe6VNDQq5X4JCIt36+c5sXAuL2NO9Fg0f+MevyVy858yM6HaD
xElzL0w19sCIR9JI/tKpVbi15d52CD9idUwzNZCxfUbEyNdFiVozDFq5LHdF6Etz
ZCvH0aEHe7R89ShITx0wlEiagxVm4l8hUyh/7IGapkIgJ6OjkKuI1VnF1bbjTxS0
qsImzqCbNV8QQYqYI5hXSj4jfmoCcRJe4g8Z7sY5WOnwgYnUS7ykdWaWGENhfdNs
mB5DAiRfImY+4Ba057U8Ld+SS/fFmVg0dNK/WTSJ+fTSPfQXh4FHupXQdGYzTcYw
Teiv000g1Y8Xa58eNF4h4WCA//pyCnns00PTLden6LaTosPpsvF6RKlYFeXr5NPd
+4J4++R/480EwX1kiDYwbnuMqwlRrZbp+UtNc5Fw8jFuDqcXkxZ4B6QggLqpObaS
rNrtML8P82Pd4G3tMxOu7s13xmi3rRKt78lAWKkM0vwsY0rVbUyNIvf1QJfymdP1
ssZbK0xt+18Q2yCjK9PLTELhaHnH/osU6NiDfLYQdktq8tU2q+ENdP0zVUfVxLXU
mhT3++0hQPpOYF3ZtQVVACOE5GkBAsMY+vdbe+iPrqqGfMYefxArdRBqacnxAhvY
b+mvQ+QngLhAP04du2XnjKC7i5reO91esAB3oFxaO+AHJKqNmx6+4gntKmwx6es8
FEdPfyzop5x91GXnKah0dxqXIrYeaQQP6bgxjn4+dweGM6pkCPUURkokK2MZmEQx
IfmHby9Xz9Ldg98QCH0GyBFGiydV1Dq3hi/S3GmZLCkjlBwGcDQ5Vy8o4dnZumbR
Zkq37pjmTdmC+EK9pdEx9dGw33lRB3z8f0LGFX19nNtQNAXVNetP2xl+kEUZamuS
5woFrVB9m9Eiqkr4daAwq5G3kDHBZQjwu7oKb6KjHd17oZ7ZkM5U4psHF511hA2X
DZTyl+n4NSovj3m3kSrDcEAGwMVGCGpCjZREZfzBhHBXlKbikTo9mC7z6ajyG4r8
fN1HwPMVYtJ9nC3bo6nOIHpROrWr8p64XWzOJRN8x+K0pHqG0ZQfOHpCQgX9pAti
mkyiEYjNvOGlcGFV805KCZhcL3SiFa9oONCK7VjmsAvlLN0LRS7JjziE+Wdblshq
gE1uLaVIqIKsWfs/vSNTgd3fPc+/lb3FHtwtdAm72uMtPdmbI9giXIpINiPXvgTK
GdPyQDOGObjutUI0bg6fWYe17Ff3t0PNbAzeyXQ9MTDKvfDFAIXu7J+3myYmby2x
vF2kobLl26tk0BueJeT9ecNdh3fd3BQZq+L5vy68BUN2YsBj2XaWsffnXJN5G6l/
amVkc526EXQI+noUnVz7w8ga4j+Jk0+cpfWjEIdjeq/qNhq3Y4hJPL8UAb7oyZWI
HyksA3rIjuy+fovSXlfQHj2FCC2rm25QWfbp/Gjw2C09yBll+NXa9xwSThfCAJ8/
1n002l3DXfpdia+1klJ0tWmhKn5wEt8QLPEVfed1Ua2E6fjhmhNUlgtIXu+a/1KD
zPuRqe/1I3G0g2HniaMWJ2oL+rAkRClL94daPSTU0rSSY7KGkSHnZm8yKQkhFb6v
j3vf+G4ijJnBySq9YWDplfh+fQ8ZJn+MIR4yCJhNdBRMcbajr03rKzrX4JIE8xsh
c0+UiHyVMsv7kvNfMZp7K/fgKq7v2bkafYHfXAeLyyNRyASeQfF7Vu1fMZMGaqgz
aCGfOhFFsJRMXqc2G+A0Dz0eWiOyevVQoMklO+lt01YvDiWdpDB07k+tIrHLmGfw
IU1jS0wyGkidjJ25qnHeB4H0AGkCF2oyDxeY8/Shr5Zl4H1ifc6GUxFCsVA6WESf
PPQVoFZ377zVXHusefkFReW/pLeBAeu3BjWt2P5vXGd02tHKVZBybRB6gK0aAjAk
c5O5kU+1JVFgiA0y+/V08Ukxx0Vbn/nC4Y+bIsYRl9XqtI4ywVqAF7gbTHRIlast
2v93xegF/NrJUGX6mSTLFTJ2DsV4/OW+rUxBcalUwCl5eU2MQhTyT5v60JRnnvVe
PJ62UszT9NYENkVEiBU5jAPG3ZYyMn06oHqvofdz9awNfaItmKYNJfEU6sPm1VFz
7OLJe5tRvvXNYaxeTM6vFVftxlwo57V4gzT7GC8QrjrHmq+59qnVmVW2zkaFiE9h
fJ1s3RW0PZ0XidI10jQ8fgct2nap9WRl3HL0jLZRwhFCDRHqjzWNqoLbfOOZnl+2
ZIrMi1evi2QsdM/UqJK68hwZZkuU2/qFVPZIX/4sB7u4CIHkUgwQPrlhvhcWIpqe
VCQT7zkuee90ae//TNjIfEM+zt6hlGyjfIk+svkXlJI6PZUSLNFKgil5SYhRZ9jI
b4n/3fc0Rh1tM7DcPPtDOQ7xEcurFgfQrkJesVC+DyWRedu3O9q5HyKu6K31+hRs
em/W5DFCtyWQjfuulQx9PcinDOCx3QDsxeLQUdGJ7e4PoFw4Z6wUOcHSGCofyXUY
jtkAPRb3FBwaYQVbFUMa6Epmsvoi06vQXAt04o5U/Kc6AD5ssqsPfyVKBpex5OJa
1OxQjw88UtC5JuCTiN5WkSFEzUmNG0VvFEXTh4kgrguY+wUJSLHZbLoJVJjwuGuL
6RaQ4U7Z9Kjz5ADMS5MtuDbS+Qs5D7+/5gcByeyWusbDR1uupKb6uCh7FyqQF6kP
Bytqxh4WRg0MKFdQhMq7dFKVB8CcDeUSBBUzO9lDaxsIlS2504o1V3ma4SZS5ib7
GKryaqIMgxaPdoXvHLRpCMuBXhObNM88Rlf2qFzDOmeE1JJe7TeCyVsqQe8rfb+W
0rfbbSlv80WgTBYE7ki7fDpgSadTEptQ8b53LMFZTfxdLVD8DX1ecMQ8XS70cdTJ
RBwowxPb67asWydPGZb07+UazYdBBjhHbjna3+hRszq70vS/UbwKxMHh0OE0LvHx
2hNVQ5zR3JaKAucu9xzJGYGiwFiIOBCr1FbBitJ/abbU7W12rNy+xTsskBEAkjtu
Y3/zm6qiJQka9LN8drjbBqvpgdo7QnKOjrxucIDCh7x+b5CGYOiMsoFLlvOn28AL
ykZuEcA9a1xDBITHmqarom/OM8Q/US42NK0e8fCkY/Jbn05A5a0NsqyV7GcHWJ7u
L7vkspdu2KmYB5fwxfwcXGG/4jPVJQs++/3I4KFTtWpn9nptZQjd+5XsrtTGhkB7
YxwxXxzMf3FV0Wqqd44dQLeRAcElxMZTKYzQuE16Qcp1/tphZP18wu770+6aLzww
cwTgR2TkelOFEKkzsKoK/vYdL+Og5g4Wl9pRqcTKQls9PaU35dbQJPksJjYmuzEZ
Au9xWa0LHv3OLqt+Pj6+ex/ne81WGmUzvPKnxB6Oks9Rf2hxn3GsCSTZDyJLgyVs
wbHaEakTfWpuTKcWeqFDSecJ2M3fRsCM+Jn+lacqrsZ43CcD68Oh+BxNL+mH74HJ
0ft2AwsnsE13MzEJiFSbsk3tde3RlK05npBJCaOIAdje6IJL4QfPH2jKnOB2/P/j
LfwGplf218G0tsq0KISt33NkGse6IaWxCb/4Q2wFj9U9mDiS7ZA2r5eVYwQ0ZBWq
2QlRnkp0nrkNVgcAT1MnUbAeBJ/nwfV2tyanJNx/6xDOeVl84y/jScL38YY37oJp
XFKsTU03QwCYviiejbNFabsMBoEoReAu/5cDNQAeN5weXE+IS9XhuFlHRY8DgqTL
kRXTKkm589j7zLgHVqTYKHkXP9QhReAAZ5aQJ+RIzL7dkfMYq/YmyL4LtngNNeLi
KoFJr0vVQ/ilUgWMMWAQIR1qSDnomK5AWDwtmB6wY6eBA1yXkn2bmIvoyzJa0iZZ
eDopseovc+jNIpKxgcHqF4BDTGGPANPUYBIqwJJzmYFvLQa/ScnO2toejfUElXHo
qu1Nk7cOtDg6Zn7n+RirIipmTX6f8it4xbEnh3xFojdFoMmJizD+fQjMd6xJAWvX
rBk+c9KhTzlu9ui1y5iBq2fgRsyoCDe+DCZX7C5GPUchgwGUOAQgSxRsJRdloISj
Wa+7W7TKjW1wsLcmSYE0GNpk2Kyb1nAKqCL1h6OH4QUx7+jmOjzkXz6p28gs58TE
V6nvHhyqpjg9td3LStcil1zsoSYDCCyuzuybRuWb2bOJFJ51ICnXZwkLFKo9CzVx
qt8gq+/KtR9anwoHtVu3jAk9hXyAvdHUH+Eze6U666yo9+wqqmGe5R7j5LeJDAs/
m1FbL/ToErjmjtCbIYf6S5+9rtnrwTSjBb1CCjrcUJlsQFbOigGJ7QoegLq8TM8+
Wvyh+qix4JPkGf9EsFNF/oVfu+3061M919jg1qQCz8pr4uCMTSh9cXrSwd2lHGiM
5WvHQhOEpsb5Ptc0j+oBZ2zFXU12aMNOj71qLnhfWKzoc1tzQDyXZD5cuQynA+uY
dvCPq4gqylMp6vsc4PRlpgpo5ZuENFvut+PEyXQWVSs9ZARUrfZ4tOS6K4TeEwFV
yvceWI57MVRaghdmDxFS1WzGXrAns7x80qDNc728wXbSD7gdMNltlL+EJJvUl7rP
boPG9xXUqsTXnZfsmDQKyTpg9AABrS0oQlILrf9+pbvqFK6d168S/5Ga0DbYv/Qr
mFiIK8Fnz9IZnRiGiDLJ1pMlzhmhd95T+3n+wmzn/0hYPr14vDTG7EF5cJKLyOxZ
WlV/yJLtxJT3brl38p48KS00WSpDzwQQeH2XGZ4xr3Ijy9dmIvfO4ZN7g0DVrCJx
iqn2FXKm+oELfycgLl4oh7sPOR3BDoEuRpIhztf0dgFwPs1s4ZvGpCLM77S88nd/
+xbAf6wAQZ99T9s/WURMA/RlxTWI3w7Io484RM/kA2g+yWL8RXumqjAhXGBJmx/P
i771anHtKLD1gT9dh6JF03dHtmKjKX2X7Sw2ADC09C/nF++Gbg46l0Ctom6sri7i
gDGQZMT8l3Lg/iIFi98NIlUjmQNPwOw0WiW+kUF512a4GmJhdoqoWcBPRtzTm796
ZQB1Ab6lBEP+YvxH4kT8nhG+cmnhSGGkBIPaIAJpkr5epU8PLv8srM1CpGTmvJVA
/NFstlIvB3PBEMiyc/7PDbNRH9wmgXTAbc2rhsFF3q473D6WNVU+9fHA7rQCpALK
Be58OIyK8GZtN9MDRJw13VZsMhFuYzDSmR9BW+Crr2LvFG6DiOhDxpIr+7vBBX1W
032jynWY4XDL7ra8Vj4yQnXWnTIcDamxma/M18h+IfbUCZNi9ZGo55R6dxNq9rEh
ckE/ALSU9+/p9FPkESC/hYAuHHtqCV1Jjvt5MvBG6Cq1qO+c+HW5TCMKxq6+CEr9
5Al1E75fgDwLKcBW/SEXBvEg1S10cb2EqB/n92QcJPcagekAtHTSM4dGI6gt+yCG
GIo3LpJ78h4k8ohNSzDJbnw5c4M54NxI1uhunoYc7dKCzuy+DIQ4NNv11EDfkK9w
tRo9Ho5k46rHrXsAgTS2Y7eM7dPB/ylrPCQb4KnQ8yDAclheKi55xeXLKEe3fphP
k8k6KAnHv0TZ8Pzsk+8x+1lpsjif2HcebX+vJTMeQ7CBJ4hiKKHGZ24DOTIvKkia
rAhYarKj0swzPqtteYuNpw39mUCQWFXr8vWZoTf9SFfFSfXDAhfLIVwE4tiu+Hvz
hEim25Y9V+d+OZZuowRotvQO1WfBtIzPMLUuglhRGQ+qnm0NfI+4czNbYkCUh/8A
bmcAKqy2eFJGwAKmeBFSfhQrEm6NFyzNiMihY/0dK4tAFzajweU0JHjpj0rZj2U8
V2bjocwvb04vgTlrmlq7x0DMG7Q3V2bOH/3xOcKQ2bRCjmq/xGBgi55MudHKGq0R
JooZuN7iDue0Q12dC74KqdBfDoauG+zudjaCKYyKfOKvhmqYupZ81kQaKBN/cHxA
kQQ4YDzA3qXDqasUAdprxGC9ZUQVOopv1oqJx/SlWpSLm04fDHN1gWUhVzoVRzXD
7gKMm2XQ3hpEwIx+giWtpp00ucleiflvel3KcmAg/SfkLpmQgmRzEyu2ThaikoF8
yrzK93MKWN8nzoxOzSE6ly2YVpBomADGmvIZBZn6ns0ZA3S94IYgxeKV6ZX9nHIe
sAoffPXB+d2NXie1LD5tWkpgQHWbVqlRH+KERTxmtxsM5BH9A7hl1L0lwBGs85fo
hw92n+V0kkHQCJQsbk223Zkab8fbqn4XDk18r/buHSvuDlSIcMcUf6m7ceq7ywZa
SglggFmOxpBfCZ+6GNomgEGhrbolp0nlOs3Jk3uNZQyqqIxfXqWU4gddl9dasrh7
MuBdTGTkuAHyaHA/mD6y+1Mn5FJ/TAbcLOWpb7B69DQbXvYzbKUCMstw+HXcLc6/
9YHYXRgFFHP5WpwBwDjbrNaIsu/5sXPE5rFYnaOraEsNhoh/8VISoRuoI1n6X76c
j3zwq/jHUcE5Z+0egTZgzyq4J3m2MG26lZbZfAZYlIux/0MVqBMnLrZbrG2GTyjv
Bj/Jnxi3WXpO1XzGLInwpFGjxePcibCEC5sRuTKFOfJVE+wNxDZuWxmQD2jHjvIz
UaHkKFS4WneNcfO3bq8j5++zHEYH06mrykuauICRDR5MjYr/zkGipkrS7O9JZbOQ
wKIRfYiaTrw+nmPTWUORVA8vnlQOkeWREJFVPKH+hJbNZxXbJf4eP8qUPcdr2yQO
Ds9sDsHs/sdPyQJo45mxEE/KVJ4A6nnVjhAHnpBn5LYK+SsnHUAdPN1A6cSi70lR
4R5FbjbP61zpS9IlueOrtCZWogDq+sWzFuXCzHHIc/w5Ru/66WsXuP2v3y1ygUIu
NSF5p3Bsp4REs9SB/tv/8sHdQuqvdt/5fGF1Sw0BP4RR8VTJZocaBCELb5QI2jYh
zz9Xlh3Yf0cnLEt/UF1uzl4Ynm9Eip1e7FMwh/tRIbre2Nx26E6fMVRhP738gMeI
v5CitD7axdRFiz56tF8wVVqjv0QbHdfxSwOU1ZqFrJhe3h4SZIcwrwiTarZhCTY2
X463bw7VB53Dlkpuy2P6qKZIpHNnnad3fT/gVFKg64jcgKwfmp9CWjQUvZeL7MKf
48F1ovIMIOmKqtsycJMy9D4X8maJfXfMtiI74MOhhb8UMG0Jm8sH5FIV6lLJjhfZ
jJgGENQ372Jxp4/gxIIYd07k1hB1T8uZpYILN1tEzPXa0ZkCN2KKht8B/MthKXUT
LOvlf2pW2OB0yrG0D+g7bkn0aB08uG3sLtskF3kTz3ejCc0fiZQSBSXwpCZE+q/9
w+Pcw1alPPAsobOCsgaQeEnSpBgphRwT7uwlEL1H9nhsxs2gT/0v+H0prFlvaWOG
KrVxGWDW9giBq2FsM1lywXc4SSyMlo7bRxUgSwhc5njPaLfJFqU2a9z4rK4eoNx6
hLqS9Ue6OWqAx225QEQ17OUVkanB/3oF988DuPRAdKNy0k1+TZ0q7YcUD32+22D8
o4XmvsBeoxH35UUWvOjFA2+nC95xatC4qKvwzSMskbcn8TBDX1J8RPC+1cmH81DA
sGHRuKCI0QpS1FDdNa9dPQCpTsATDDNDRrvVWMpARZyWC6qDKnxYfuTlHWN20VZI
rkw+oq+AQ8uouE4FqB1puZCGR8afyBMBdCWqhdqCVqlOswRTg1Oq9ePLR0B/rgim
PZVkjwooBaCHOA+wNQD89Q7cJl0T7osOT2oNPay4S8AUf1m1iq69H1+rzix3NQfq
+gLlQZJiSX7JQF1NsunyBiTlXhfJo5tD6Y+XaF6zkLQL25MI/8F3GKR5FuxO2ryh
eyz7DNW16QlaTeqG7F8/rtdxotbIy4uWJiV3dHa0c2r0kTgKdg5NLyeqAPW3irMv
nkU/2XCbk7NBDpHiK+dVLQJgMp8xjV3zohNrcjY6csTpM5eds1MKAAkIC+mDNY8g
RV28Bmp6B5QvRbf7F3HdRFPSW6PHlqsP0IbSNrZ+LJMK7s4WkVRwXYl3XNC2NpNt
q6MA3gc/4AGKu0bOsK6vVue0Au1bnmfumkUJC9nibQehxSalqbW7OB37hkPRWalO
iWlEUd6dBvpaFV8gfcyzAwwRrpo3hgqIIF5LSN5N19H9RHGNTZMB0ToRV2ujt6jH
vUvIKR+LhjP84ijUFIkQriw25biSrfi3Z+TFy4C8pxtJD/WO4gagVR03sE6Y364s
fErRlcj6SuuOoQJ1y4T6oOllMLpp22w8fS8cs3XtC/kp6CtE646qWcg/4gVpjrKh
Ofzg8tEle9OZxIAA+mXvOuW9a7efCULdtbXO1+tsVJJRq15dnTtTsWNO2rSsGyhb
m/BbSSnFgtF3BtpmSbhEot7S6z2GUxjnJvspuUf57OxsJyr5izvQkCQrhK6rRN0h
M0mLGZV9YSvt4kpH9/zZTh97Bvvqb//RVWoRTZE5tjxFJJ1fF5RWexRAw3WQhoyq
GaJYelwr+qrjYmR6qLBnFY0JjJWS7rT0gflJcQiaiOmYWUi28q5mcySg1QIVuHWt
Tcu35O0NtGLdf9neEX3s8OrfmuAORiUxTSbn/wF8W6C9HQzUx8oWF9CaCNAFA5iQ
nuPCU9iuKVSdwc/ydiOfYDjVRajs1K7IU24Ke/8R4zFXYNkIgmaJvSvLODIf0qwU
N5Jg+QirTTOK3G+iKRoAUiPoLJpP33TyHF6+TAibs02cTWm/AN84C6MZzkeNdWaV
MeYfb5hGQnHPRCmcyeiQNtBYJyayMQ0rGoc7U7KFqZF+tl+RQeqDCAIRjg+5zjK+
M0uwff546FFm18yjsZVx2frx+L3yElTpkFlUH/tYQjk9JtstHqD1fAmqxOilviQH
NiMHHTM9CtmtTMoG9wgyKSzTHV0/hjGSife0p0bIx0hRtrDO9kE5BSewbimwayFz
y0QMIJWqxYhjvrz5EhBsLSLsmAoTAj6yaWfchxjMynxBaLeLXeOAPmDUc6D/sq++
Fy/yjiVHddoUUxmFs6ANf/XUyTypgDVab/qOiEmOzAPl0d6y4riVIeJlM5KsvLsV
nnyRIF/GIq1WW0jCnXNGH9bZVU9ojAMcKjOkR0NFFMNfEpBnWhSabDJLe8YZdMO1
Hq3kYTm9XpZ7Savr9qlAhEGvaiFO3OvRwi4Z8DA7FS1ddva/tgPcHv+R7e7koinA
kqG7tSY8xENa4bG1PluGGjFj+1fZQbQdGB+2fQtm8QMPMQKcuqsOZQtyPo9NAiLw
nF1Oh7ayOVkAUm+165tqAU3GEu0353L2qARAYoZZJlfJch/H/1YiQYxKVc+dJBx2
BwoJJTOBOTRMDG6UHznQygKkShCmgHzaF76sptSJO9iz81OTkSl1BiuU3cG0AevQ
kyRe1cmetiZw0tP1amNS6r9IZg3UWh6K3zMO1kjOeV3K3kUoK/mQ3n5oSd9S12re
35xDu29QxDX0IjjibgTNw+7wbcZ2nxs+T/vJDELVlIeputjBkYx1cbckTodnFjDm
mDOcmv/zhF3UO96zeus1WNSJkqmrLlaWujgwkBOqEtikwPP2xOEGHUZKeTNvkqm/
zNQywS5zAZ5VNy7rk4ohiDVedZG60jL9t+lzVhX86XipOipX+idyHG//OXf18H4L
WQhqKtitLAENWpMAO+5dau1ic7EFPTNhim08fimFEV5iEh+XRUYN+OXPrDrQxE6m
PgjIeFfiBom+Hze3SB5f9TaFB/BZYFE7I42o08JEAvWK1Ko8nXaZwcyi1NFbZbQ7
wpYfUcJ+gfVO+7r3PhYHX2QijlTioISGvRbz15HdK8RyhfFLltLRjE/RCzhldEAY
Fjz/y2KxR27jiJEHd5z67ZNUsxIA2O/fKRJQyM117zyJxAXFxdEOH1Bp8R9UToZA
ysJEy18d669SvKoFf/etwpXIUBczH+ZLaju1BqYEPEdOusHfAQRu/ygXl6UJLqLI
mdoS5+fO8A4n32j6kX9p9yh80XNY+wEXKIiR6GIWLiNqi1PHkL8/Qd/yP3kXC89/
+EQoZ8l5/kYSGEaj1u7jLFW15Zi/nc6Gj6kQNKQA+Gtwaov/mdSDKqeCg3c+BEPQ
NzqD8VoRzD7QIYi1A5GU1FfgxtLQK38sivCt2KTiV/cxoRFRyMBklHZegmVNijqP
oZRg8wD1PKYjgUlSdp2Z70NkhTqXK0TrEu9kjfzIxOUSwiahwtf9U/gJPMHke0e0
pxc0lAE2JAPVHzgc7SJSSj7Er7KV7FKIeqbo0TF3Z8OPfi31bMPaQiPcOE9n3J0x
EPxBbjhqLHa02ceCrBOjtDF3NK6+EUziHre/8CrAzWXeC387HcaDYVepeHBboKpV
ox8E9OHcWXj1oRraorMF/cK61hRdTmgAUjJIAJ0ZL4xtIORt16qnG9JHzTzv675k
A/d58Et+8PyLyBNo8nyezcSQPNlq0p2toVaBb67dFx1HAP9uC3fPu1rBsjWXzvIx
5ql6RUIRGkDhrBBU4lU4nGsqm2o5kRXMgERwvoFAVnucPdCYPsWCecWERSy1Gk+F
4EzlQjclkVbmDv9v/pgFIQmgPiaAtHnvx6EMK18SwmOgLQaFArc4feGHJVjflfS7
KoRH9f/vgV1JQuk5BxPlSZxiEf6yUHNqcWnjJdeFKANvFIaFLvGwVq1YkxSgNIxM
yJeu31MjWWExJU2wdi+dGOaRebL/RRT2/9ng9qGQx+L94re8nfUt85s0Cv6M4AE3
XxB/388xdTIHN8itXlhsMWOU2m+qk6ZUjFGV2fEb1dLy7UuFf6iEGRzagvRhVMuF
GaiQDyZfgOzO9E7d0+NVAq86KxS4mzmy3V0Ovuddo5EPvGkv/7bphEzcLRuzGZ/n
koqHinx/G0EPeA3YryKSmNd+ui+g195oJNy2/Hzj68LY9JnMd/vg9S/uVvrr0EkC
6B9yq7fhstzYUIWL+pVg7lTdYMnU7A741OitBjVvjlwM2ZAfE6pZzzXPLfgYuIYx
MCIdVJICxLa8ZPsLv5jzekyZNW3jKCeKLMJa6z84XHVKIwVQvEFRzTsok/Fl/T7j
ELbWGlIZ1edGTNJ6oyqQg/KcVfhgaEddYZobTlxBdmUBks+6CQq5+PfSGr02QLeV
YF/qHWwMQE/rnxCWtJEAVsAfuYxqx4e0IHxIJ9QsRUkKprpOQalJiqq8FCFQGNMQ
kZ4LvKsIf0PjPnPs5FmuNdLrOsm8ysKx6rThQpFKeGpPD1O3U0G771giHN6tjJdI
USyoD0Tu1/LzZBXgYJZPivntRcF8VA8tEcF2FPUnB2hOzDZP9I8ZPQljgVFzjuJO
8xUrqcIhVFYPr+wMaAMt/wJFtM/O4Hvpn6sZR0NkZwsy07dzvOC4DElxNA/25aYH
EI6rl3TryyVLjb2uQwSGlVg9WR4FnAnQ+6m49U5c3GQxXphGL6ewt+C3+h57Op/z
EZwmQtgIUiOxRnzUYSxCMM2W1W+rbUp8foyZwwTKjq/YimvBY+XB2qJ0FtKAD9Oo
iLvvn6lBxsI4BEaQsx218KusD1L5Hlf4u46w7QpAVTu61RbeSHeXFfMpPuXruv5l
7Qy777odX1A0ImZ8T+0i7LocZWtLVXGWxs3Me5gFJECRnSV+ntwa567jOm7/PyJ/
hTcIZAzbyhlyIbRRWD3W+7uTl+tejU8V3jhz4Hs8YEZjPBHCDHCCSNVn2sF3BR7k
qrErr7UBDJQigWzQxJPASkfUH70R+iBGzkPXtrpoTbgQKavKaCFcZa1KVuh0puO1
chSBkJ6U16HiLLaxUU5blNYItPCgD1XFkdUZJz8OJ0ZE/LD3mrZkzX4yonOVsWB9
7pZkrTfevEbLbMGizRX2vBc/60jWgz4I08RoRbHSVCdnYA7St1OombceEximACTJ
P20qM27RVdXdBAwgaJ8qz3O1Am9gKa9w7RHBvJBXpF8ZiE+3TolAuuqe+89dLlN0
h4eTEKZD0dugVnCOtXMDlFL2gynlHU55VeISOgCsMq9AFSWa6S/DJKlJyh5ZdjhU
K7E1A9Fdbhl7JPrAdhNgwdwjqERnN/GjMOe9hSIezv73TnYixo8WjHQ+Rtgfsrmi
njbSDICQOBp3cNbIi3dJfBjBLQ4QqsTvP27FUgC6Kq7Z+Xt4bbhbXCXJdTyO9tBP
ihATKgtd5hyJRufcpVOR03ZzB4tS8JhoQUvj8Y2D6KOq52jWxVc7aUyt78RMU+t/
tn4CHdpYLCezgEdGhOyJ8MM+M0WNH4IqtEMXX9O/L05lyBRN7hvd2XsA5lGmp7Yl
fXWBOD53V4O9yRDww+gnp1446pM9yPjj3Yii5MUuUc/LHN/tvprI4rybS7RPk/Lc
ymROI+PCMhvLJdMREerbvksV48ZeE093vOeRIe2tKdERNm3c5mVRWuraL+LOiTyN
Vo4ZR9mo2+0GZEfSGBionzfwmtAoC/j7F4peH7gSigV6mbL88Qwma0rJVUWrbgc5
IXy3lGN87sZInA+kew28Zknq3tUsH3r7HSEeqo0eimJ1asFXr2Q1Hx22HvVDCBNZ
KC7yzdcuA1pZ6NpRgrswBY5fXXtyL+Zm1+5Dn7mtBu1wR5HfsYiNBiG3nXh5SNt1
pWJNFDiqYv3msOoBd6dn0OzJEf5qZbhpu+fWXt7xGF2Nn1Q4+VzRESh4/zRBFdO6
OromL2yC2MhUGcCj91Ky0MBmoz6ONqpoDmYRhuq8n4P6tWJ8Xw4839ii5aCwtkzo
KzTDSr4/gT0TclzmMl3aZZ0cp1r69TjgeN8/3sGOsW74CZIv6EjbRYeLXUqeOs+R
Bu5LQjUQH+dwcY9mOOD1jILflg7/QDN79Wcz4P8KJNQzVpzSVWIhjXdRD60XyLCl
odGC+6l02c8G6JfsEegNXIFK2Bv5/n48LkGl1GwdN4NuRAan9NnYyARBZdQS4+jo
PImDdvSTJ3i1sW4KUYgH8SADGmsXfq6wHeB6171rxFpdpUIVvVLBUe7I5xySZ4UB
f8ym8RYVGtvVXuTf1IrCcoNb3jxIxBKxAJ69tsEC/MzI/Cob6kgS5ne3MGjBPOiU
q7+5r+65mqF3/ZAS0Y3/yNQElK4LezkmteDQgCjN5L1IPoD/ydWJ9/jTEs4/X32H
bYoeBBiZksu7TkRMwhfVgA3HMLDLYHBU2fTptz0VbUD1ptGu32VDEI2Je9oFVAQK
Y0lpRcsiXOKhNmiSeCmMvO262CwN6BtEP2/AeAAgl8qhQUrWDO+wA8LLizFQ1NJd
R0/+DZoadqOJPf5HquMpGoRHor/OPSBl+l89kCkpT+KvdmAcykv0wUoHn0VCMoB2
eyF8K7GDblDldd0JI41Rl9F40M9nyIMhmCspzNEryKJlCdxSKhLAs957dnSJF2ss
IJrKC7UVx6Y65K2rH9IKjIXsJgceRFpMWLE1qmvzH5cBY5hKW1ThaKYK7lLS6vLb
izd/pIq+1IfkM9JPPxkzTi2rxEWmHXozPizMuVJRZ0q9COUhQl7t/f8xd/+/oN61
H4GD4xy6vejWif0t2g8lbm/z8zDHCmr+amSKV0WNzXEZxhp7EOMg8dc4XV1acIL7
YsHwo0SToWdJGfuqvESB9Rw0hO+M2rkHEEz51tA2Wh0wB8/dtw5rnl9RraArQkRX
MA1j2v6++OEuD6j/mopy9W4J+XapS1lc6/kj13aS8ZqGdHyRL70E+xESSsUvCeIv
pgvUyy+mmqeQyAmd8HLM7zTsM69naVtF9Ur77YKID2DZTlQ84wngZMag8/60ePQ3
PSGa4SnhNzFmMK6UC4Ceib8Hz7maRnrpvVE9cWBozWclxvG5j+AsYYu1a0aagq+J
2c8zAx4lSOFA7BoyhCc36aLTQeHWPvNFu+V2jGE3JE0WSVlQnXi/4ZpxSu1ewW31
33H1geiDeE+o9QxGG/AW8YF3VMJOWQ3qEEaC0lFoTxIvPBYVTZ0+a3/qZQ1eKl1U
LcOHVBHuSJ/GBzQYbNdlCL9NkPgCC7zst+ClsARO9J0B9QBfU8glLl7i9AIi7dXA
LipKMUqxi48y0CeIoniHLOHVATXTuYzPIKxQjvePB7mrsnzkxWF1WL29/Vkgq3sM
t/qgOI3DaJ5ybE6zJBtLmGzp1Jbj7PWyiY35hx1jvujMTxzWGhFGqe4CdKXa7luW
WQCxYPZJjq3a2G42f2ggTH0ONJzTYF22hlT9x8EOlZ+Ux7YUUCIX4zfQu4zdpym+
Yxnx3y4SamKo109T4bHD/ONlqTO6V/h385+xb1vI2pKNa7hz1T3Ep8zO6iENY+5Z
8ygcCFKZ/k/N3XtoHcYgp+LIN9ZEyPSULmKC3Abd3VLBj4YXJQn4hEYorm5BBjjG
uf6O/lMbd7yMnzcxFlLr2lSaNkvyayy4DTqGrdgRnSeW8lV892uvwkw6Nfl6jwmU
dANL8K2ArfyjVABXtpykloaxVfU9NeGglHBHSOJX8husYIGEwmyrft+AOLi0nCUG
9PlqL8D80RvZCQpslsSxOSZ5x94uAqNPvoBhcG8I388d+0QyCwVGBXYCslWvdKnm
ZU69kjq0cSaMqo9BnbUSGFG5HkKrDbKHewLtzsFC5h++n6bqp1A5BMtUuTi9gNLw
vHQynRvpqROjrTMEd+97SJLAtEVhV2o6Fgg4A1RPcApJ6tqH1B5JdHIQM3NnvyVu
eZJGBOycpGVOrgTa3NQzS5kWOfI/Nd/r1J7JeXxv1+eUa6RJqUotWYaDHPGNFNO6
lnRpD7ER5bwFip7XzjyDrrVKAqLHL8xyr/kqJri1QM5foZ0M7xVa6FalPdh3VetK
lVkxiQ2fq62QGG4Qm6zWFgAwjeiUksTaMuQ2vGgVS0fv7azQ2uAeHB7dm6qlUaTw
UaQWCW2UMkg1HDtUX0Bw8PvtckWB26sQRdNtx7Fo6UYXgqclehggT8M45X1gsYJf
okiulxwSZ6swJjF+iBgt3d5R3gxZkAmjK7UilErv7kU/wmDCn2SW4OfRRgusbvm6
j6Tt6HvkSXRN5ubFTGKiDI66+rSl0Shuwg6mUnUeyO1a6Sx9VbNyTWtyciTWsFiK
nloVWCneTvBwErwIUIF1iN4xr9Sv/RDyCPYyYJGmoZGT1GC89oW2LLyAwkXphFOi
iZNiKOH9sflnsHmUqvCTyuIOoJVtAuEJAqPkYrv2MuqQH+H18C1J4uRuQEdT4v5m
H1AEvSU/MpNe4E+c+PpvVGEjIYzk6mvT/+zftTCUjeUxPHN3sTP68NlqNWUaCFSh
Re/kUupHc0gG0p4CS2kfqM1tJM/AMKi+u8+/yVwp1z8Xa3Mnys3eK7g1cxbSVYwu
ccj5HeygiuCLoPgrCBGNLcfywZGXOJBlYJYN5rH/hpgG42IG3Qz9tkW60k6mdhan
iFvnebDw3dyKJ3yswi7xr37Lfeud5o6DPRTPVQb3z4A0OAq8KNKjXZfs7lc4+/zV
gYlWALcm1bYCxm3Iq6w1lycRTcBezqRzDhB/SwVFV3MhdjomvLZeEFZclYDKKHlF
CCmcAnBeaw540mg6/YURWZvuISnuQGhgQOY3yNLaZkirbAz0vQdQS9nl3s10hiuE
I4I0YvWIH6HCHgyjQv5oo2oMU9oVFc5GMptMBW6LNNs+FCXbqYohVEpkDld3vbOT
KuRtdKHpI52EKamo7uZJLyeSDYOfn0s2Y7Tn9BHwEoClwcyiqr4DtqFaelhW/z0t
xaym3I4MuZP5UtizAfv61dQtMTvMae2Xuu8eQFT8o9Ey9x72wapa09LhOFoQsVjc
MjYGPAgSF25FaNbJtGPkiiJMJlzsrtZRNYnmZ282+Q+jilwTjmZQPRXgdfKQUykf
4spYZrrvKoMTETgkVGuU+PIhhFvKX+uetQPK1EXFoNKAxZm/OfbRH2bYoPoqK2DF
3UIi6f5wSa0qYlC1tusD6Tr74oGTDiBJGs3+KEI+2DAXu2HOZgj9pQBds0o1Vm1B
vQgaNYMOxScWVOpEvLxJH1HSi0IPQ6ziU/U7JUd3MfGcV2yX7JDFp+TC3QH6t7iB
CBmkjcMLvQV5GIAFulX2L0qiBpVesljy+7PrZ3qLgoem0RiB2q+oc/DeeN/2btpe
/2fqF6fsp178AuaKg/kRGw+r3jMapMzN7FhhQL8VADZRpTywqwjwTjHCxLH2HIX+
+yajFhsPhxXhgnPu347qotrT/7RbnnIgktBfF4F3Ld8xuMMfEHR4DyGAcbObJjJX
B9fqBUC/5BdnUo/dC7RKJ4fmSLw6vNmDJ9S7ZtpT3MD02EPUopbwri1Tj/Pj/gMT
pkDOh0bQBJC/3BXuznOFUrjGYQkMq2+G1JMzHs16yw29lMD3BETZNpbyFJuc1mqY
EJlt8Abu9cnN4Wdkd7Mr15P2vQMprxEKNlULds/ZTtu7wKc3i82O58vLm2sGCASc
LMcpIeUHUdAnypW0TjYDTbNDYD7IOLRzazp9TFUqj+72tvb91b98F5WgrB/aZXGf
Qw071x2iE3RixEcAv+mfbML4ET1E/m4hdlh8lN32FYYfvEooGEPi2dGZn5+R4vB+
Le7lyCPDrwOKhUw0OjO7d3z0rb1ZDPQkysKebQn2/eBSPJ+PE+hpQgGDV6+QJOl0
/244OYusezRLH88l+CgKCRNk5hhi7N6F5AJJ26cXfpbaF2f6yY9uuGigJHvz8sg1
9beTp4e5a7WbdoiCucdVEwFhqfV2yuA7iM/BiOlzja3eFF73n+c3n1U0/d3KbmDv
kgCkLz/lni6tGjFbsGezk7URJjCOSNYeutmxrC8CTiMr4DeCwY08wi2fba3tjOnw
i1tzBLKZzJ6MvDZDgEbqa+h67RzVNZriwnhGB0ICbGbQAOkd3BfnZbXLMRPXmllO
0zRPf5q2uA3ew29CZ5eG2xjhnICmFWwIt+W+RNthJw4Ia/qvS/SmDGK35mOvTl09
M0a8uachb5PILp8Wr3DealB/a1fQaqPJvxH0KkGPaOMQRyV4pMslvLFi3L+wi4Eg
cs31fgN1nNR5ZEku25ZqtOFUHQ4fti8Ax9THgZ6h23+NGMwfPGHjNKercAqeQX3r
zNwLPCsKJPKdx2G0gzEdaJ+j74N1k64PvmF/GCB2Gcr8Tvglbnrs+m8KTVJw00/1
jLCWPCBD7JVUWkeXbWdKWsM/Vrn6wFfePUTsTyhYO0Gjuh/wc8hmM/RAmPhl0o9h
lexqmRbJ4qRgdSWGUJrXhTaaB3qz57uZOfQcdtJBtljxZJVCN8b7LaWQ869elxw5
YmHeLBNAsQ7jeVkDp9fKI9JLmQ3olrfF5yDwlpCYwXTcMLxIUM3Q3EcUd3MfskQz
LfTt2qOasTTEuW9++GcLbgMiFBDr7mgETDCFK84cRO65JGH6B4wPUhPWeyAUhUGP
50MpSbj/beT/7rEtUwHLoH+rFFqmPcusq/eaK4M07qsHNxH8H//5ZasT31wlC4/L
4xkVTzA+YTIzPA5xFTUopFYEjKBRYjijmSSyG+t6GgOPD5X8tGU2GKsLm6ybl0aN
c1Xn1zPYT2IFJOXiMGWzhHAlyRKi4M3y2mQDeryLxMsuIoaMESHaJjXTJFa9CJuJ
cwcjGrYMWayP/Ho8J46JVWbwXfjLtB7N+YLil5utBh7A0D+iWJfHCRY+YWr4iv85
UDi7ncd7Eppg7Ti3iitWeWqtPKaZ4PMjUwINbbKFAIi8qr4AJPMrgFO1ZbihWJgA
pykfVr5FM7+T2W0G+CRZkRHr/EfguCMYRjyQJ6z7q7TXFUgw2IshNzYZvw2UbZ6W
lnuNhBumXFtdTZjpKjkpXuKznow3XELYKkavMvxmzs0U8TuZFcT8ovwYZFgUh+GB
7HZjfSRcWe1Yr6Zv6996Kt6bSAvohPShuWE1KBJRNHOOb5d7MyApbEQtqvDp4bVv
F0eo3Vg7i8oorluZcHeaT726ONKQGeDgNNjGNsoy24WlYcOMLlq67zpPCCSVGFN5
c7R5LIugEWlOLR3L/g8czcVg7ygkVcszYBrp1NzCxoiRHDx8GdhAY5EHs1A2c+v+
oIIDsuVgRPjOcbnRYWx9AsILY55k9cHVWbhqni+J57Fpn6okiR+retFNoQaQcuNs
Zft6xQNl75dAKQJIVLDIPz+mFLkfOawyv0gwvzRQr9m/qlZ+6a5dGrPX2KtyCCEA
5SNMTZMKSHJbPFL16IczXCE53dE7A/AsoO42NSlWCPwCJxvbfTLzxTVJnBWU/xDz
GYGY8TZwqvrqAslCE+nNTA7LqhW5DIfiMBfyzC9jCWwnhVfMLiyYKMIUl3mMx1pt
3teo88GJoQ+HmN6hllyRKoUmLiw2f9lGFHVpEIjs2cmsvXLsTCxcBPjXuDfJqPoV
ur6qx2J0KSqFlB0U19UZWsc+zU2ESLUBCIuwTZncaeG1naX1Jh3qW2GZe8gvdjb/
lQs8C1Pzt1UkGIcjxm9oYzqz4F4pDtGAcBrl+bViaLbcJaFpx8v1/DNmgJFvvDe9
klxxe+B/QwA3gO6Xb8RQcDt3c2fU2xoRU1oKarMPp+m9wCqzsMLjTDEqwyROSMfW
GryUySg0I2IMsYXMImWXQatv5XGoM53ylzBk2QjTs4ggLz1PVEdDd4ditGqdlpfG
Z6OyBFIjPI8WF0v3YIcxJr9RfsttnT5R66Oi7/KtV0cCy9x37l+J8cpZtLmbTNYF
DdepjGndYs4L8O9/fOtVX1PBDPxcW0kgM/U4vKGm0WJ/Iw7oDMTNVnAR5aLu2edc
WSan74PqIfTKJ3c+Q4VTYtbyFQ4DH31yQHipAnmJCU6QNfduV8/Y57SgSzRZVgc+
QSuot456AoWS1ec6M87z46AWvScOVDBCuHhekSVPx0dOrV16tWN5QI+5gclmv4+y
3Vqyv/nulUEe2WN5ZJVv/jzb/ShzdmLrCiug5KLjnQIIvQKNFnQ2+cZabMANDeEW
tJD4qkDHrz2tVVGXhZrDfVQ8W5BJkM0nMcb4oYqDrKYpibW899zB9fjkxCmNo+Mb
udEb4xMqmXgyirpHk/peqhecSQz+akNKxQ1W/AHkHDUxZQCAQuq8+cyHcu7P+l81
f1JU8T/+5b5KGG5FivUHmeBdlxIizRk0aDsua24m4n7T1++rrkcRBjHvH2TgkI2c
03xuV4UJJOcV+LYIXRuGC8TZYwa02ie8nhCAqNjKX7JSyeChAE3MHlQMl5/9gfZ0
KtlSdnV30Td494+ZjSDNWj7d7B2zUpan912QuZNOPr4c7SveIO9A+2RR0zS0acw5
mPTtpRuyILIueJ9xDWhCSXsX154UFfyx73SwJlSYthHyoasjCXqfEOEn0EZs64ZV
X1o/kec241UbKCt8AHoHZ1naGWjq5EGbeUHr8lWSt388YjITN4bKaGRFCa1Zx86g
n3zxY/9w5Zci66ytCQCtfeYAflGV+HiiEi8lhakciWkAKYSxhwFoxs/pF7ivoJW8
TlyDu4Oo9BoYPAQiYh/GLUUPLKeUUSrwx5whIzNsEpFQ0QHbld729I8zMLmjEHBw
NY616SwKln+SkGthT94h67IvmUZYsiU2rw1viY/4nrI8tdDJVYNiw+Be+JfUljPw
YGSJWJkS0lheoUHUc8HPbim9Vbz00fEBH0WQA+MsFnyHwMFy6IRz+ZmxvsGtyavt
zcSMr6S9Pe7r41vY36+cM8N3YvnL8d47LgDwju7/4K0r/XMHdyzvteMH+YQPuSjn
uNqs2GVbkgAZdddCbXMCeWx+jIgiFqo7QX3o0ahS7E7PUyCYbGVRYx0PciAmmjth
5fX1LL40Wmm0QIimOCStMdfhvLF3o3tNYwqkxfLjLTZh3EpG6XbvdvHWMI3jrwSg
9dxpgg0+KfQvXJbxRzBbqgN3glCYgnsVFATGk0oi0yapBT0bJLqhruR6tM3o3VSF
HF1e/bVFcKElDmwSMq8TrsnyNlJEQF1NClsBknc2jsFNC5sEVXrrNJJnko5dSKBI
eQ7ymmDEHNJJ24iX9nJqSw5E7rfkKG+Pw2p1BlIOPzzhnAkxHwu65SXSDNGuLcNp
4cBY6MMPEpqmyO4NVQkXIFw0vojn6aDZBW8ZWq8KBt5kfT8WCYP9FAQYRZh/R1+C
wuU9g+AINghDhM5uJP/NDk3QAyC+Hvop1GJnfugrOUXU36/qWzw8Ik7JBpDeeViY
tFrLy/Sn0yXHi6Q76c7ddjdNq06Of6My4AJQYpXXvD9ETMexTS2kyJoCXBwhBXht
coEyPfVyfi0dmE3MCWA2kIe90do/3pAKjYzFJzuYpPN7KHJYx2/VcaJsXqBj9PI4
UOtfhuiKg7HDJwi3odwhQw0VyekJmVgmiq1tBOlfsCuD6tape2HhSXhK1fhMC5Bo
qOCh1RAkRmDVQzcKxDKyYyfZ4IDSzGW2Q86pGFGiq00H2KuHj1+F4FB6jD7me9xN
WKv4EmOtXHPFuT9CdZ6J8lo7TSEQ+lDqvkdEVwM4JeOpjWJoNJAdw14IlTuEB50l
e/ac6JClzESwohUJE89JhNaR05dgjtyiJ9Y+N5Sosatx/c/NvPjKDEzGQDqQrvK8
N3yw1QtHnciqN6rE2EVAQGCpZO3FQ5jwQch9Nsi7kycXfQ3Bavn6tVwUzcU5q/ro
gQQ22saQVQLxRw7/ACAVO/d8zXcN4fgiTXT6G4MQe7Y29Qw4qvO5DbnPaD1BKhgg
aUPHX3y188WKwoepxffeAOZmbC0P7qqkU6fkmwEa7kEGbU/8HveDnCh+fIeBYu+L
S9fv/hLzMIfqKRG+73dKIb6NQ+Slug8mkA1MecZvjwGLsYgf46xVlSWqRKWUMmXn
FQuqiL3Oh7ESkh4Txzed1gVokfEsTUzmuNZgYswnQ868emjcfVX87NsKC3sSf0hJ
qN6/NPw3WYbo/L1cCdH4OgKlMw2H6j3SWgAsFWJEbPF4nsZxbW0UJGkq5eumsBK9
gj7l+lJFQrMTcRVyQCWNAdEDr3gt14dkS4V1vUjmItlxYpxIaYfqF6WB6rm5BuKF
Qnz2kRBfTL2V6VfnpT24i0d4c0QuqeU8W+GaKcBHAAyPpu2yoMHqS6BMgtTPCwSF
+j9YK6R35KQt1KiLd2q6Lw4Eve5xuTQQEPmaYLjDoW9Qzp+I2FfaEN80981y5VM/
XoonCtcVeKiY1Y0boJyGkQqm3UvKapbAZS2qNnskY39k2fgGYLC3ijX9NQbGNGDQ
eLbA2NdNlJiat7P34l5CFI7vgWJBAQOTaOM69yGsmGaf9RPx51XMV0q+cxgImmqY
S5Zf+Cspp1mONzc9tqqoTGpqkuCjEEK6JR9+8Ab4RmAg9EA8fzJwR/vG9nqVTVEt
zrJ5I95TaCpRiQ1GjTrpIGsW6zIPUqDXbxYTLVCwI/u7m95fKnynR5fu8M+VqQOi
Ow9zcxCkz0VDOKn0Rm3ba2vUJa9ef50x7YVvbIByTrf5b0rabGme6ClkGaTrh14g
ny+tXaNMRkovF+6LO0gX3JaMzNYAs7da8DBy6t91fvzzJJNK5I9hakqkxYvVMZtO
JmJZBoI4/kGBHFv9/ZrsfTqKWOQtOVBOM1NHubDioydIjhW3QJhC+0m6XqK8oKOn
F4n2iLC2Kd7rZMkj7zF4v/zbgdzkix/X66+KYu/LBH/tUre7rditCD4KcNwhfVXz
HXsZfEioecMSBEroJfWob6lP1PB7MTkGIyJi9gy0hifFeglHljlVuIlLUrQc5fgL
SoVNTMsNHfJXkgoJ4U4niSq73rT/gxC/BTZhSCTUdufaShC5LFck4aQiD5lUtUrA
fICNM87qtazLUS+bVqD9k5iaMkFXGvh0VoBY6WMayJbjyqXMG9hJIjR+4xpMJR10
/8hKOVLXE/vAFoPYNeMatPp/4BfGgpxNuNCnIhnzNrddCXdMmuBJqhqDo2OZbmIz
pvw+PqGSSUatP2De/mSAwYblQfOTNTeF7Pfei1DKXPDCbgsKGE2KURZSDiwwyLQw
/i/AEZ4KHdRbbaphoXIsQluYBpZQy3A4xLP7bX9XTux1VHo/XDFPd7ylpVRuiL+Q
8yoKOkDi8rS9KiTBt63BsCsnWelYLoBlUUC3jNv/ldhCVy4eWOE3CWEDtnWEV8gr
i17urLvOMdA3jpp/NqpS7tkE+4sGVJuZeqplGnJ+QjLpDIR0FY+KRONsyeuDq5VN
iY7xNb8EQSeVk474tI7qvIbEKKHkS/0WQEeuEUTSsIAMDeFxsrGE4s4SbZG3AuRr
JJfwvEyE5L5eooleAdaq45UOLEv99PmK37DLLpVi+e3pilV+LeoWiBQG09nF5PZt
J5atqaiigWUuVRmzuw4wOZvdaYAC6EVXfWTtYgsLezhYO91r045TIFQlqK7bhXvy
gs6VOZEUy4eAuhorrNLNPc7Q46DiNOBQ0tzLA4miszp7qMQb1JRERMRI3hQrneMk
NJh5/gzb4jgmN7KeGt8d2kmTE1d6Tx3Y2nN9iHMmOkiQTMeBff7D56KMNucuiHl0
MfRnNpVkfErCEGc7x1ccOLSBATkgIDED3LpHPBOiGU/0A4uCZvz9iToOhPPFIZDS
ocr7si5vH7qrPEHO+IMNKPX9yvRrooK2CJlwCNxarFb18RzJKQRWcbKuhKZCbgQc
iwAzAKdnodzLfQS5LCTWb24krL5CtMvd9I3BAfUkRwtU2YhXz2E5KG8EwNxTKUkd
gMtxrtx4HdOllWwnsVN1CiKrW4ViahDew+xi7WZiUoOx86uRZiejcvjzHlxXaQ/1
HagRB4pxYcUM7P/LNRfKVZPtwWMx7WZEnHSnDFOHr7m8knEmnPmeMwNrMFH5QcPd
DeqzgihOWzG/wi9V1+OpIIS8TLn0E5Dz3e4xnpXZ+0fIVvkzBruHMf4id0zQWwxf
r0g2dyeIWkPZhDUW+THn2h4urhGMnxjKaKPOnIGCwnzH7SFLbNzwOUOjxu18019p
KyrIAv8yePJLGKfOHhLsMO4kkhueAUlMvHVwnPHlpseDsaXJ5S7v3jh3zjhIzql0
GWsKILEfvYovIc9CsUGsGwcWLCyQTbypX5YZhJI/cUDfLLVvNUVt5t7jrJuBPkhp
VESyBm1rcP+VrxMFG+Y8QNlvzFihR4y12etABlxkIc1W80EO7Sh3BekHnkJVnXV7
LUQgPD8epNL7b+8W/e/BmhxdWkyC+0oDZq8rFoLBz4tC0fK26nEhwEsJAUT+M7Yg
4NDMBwe962kZzJfJtMBm1uy4o+wFh2/wKw5zrw6VFLw4D2NiGCISX+22oHGX9dPe
eIVtzgWP8wHg00sGUdLRU2YOsHX11k56TxHUGFwjFhGBOVDdhl6vpOV9XjtVMpPs
p0Sojwy2JMq9BrEL2tQEC7Eq5TrPI2p7FqTy43cNQj2Fk8ym5thS8hh0xV7t7P/S
KuZcuQR0gUJW8r8SzmFEOzsYsDQkVok0JNkIzPbJmXGmGm3sPqD/x0I0Mv8oeyWs
5vziYi9//2wXNcyvaRuudsF4GEHxtC/nD/7NCLK2DaSLs8jMuCuKxx0fvdy9fbUL
jKqbRzC6spnKTONTqauOzK6aox75rtcZ5dG8VWI59qyId2FxhEBQfg9fDxS+W/id
/S6UHyNnvwe1Cs0o2o5TT9LlilFOcKsG4VxXSgLZRAmgV8xcIYangDfJuNxhRQL+
vOTJUP/yC9NMX3P81V68wT/JnN/8FJrju424jfht4FvaR6ZqwkuC6FkWg75GAw7d
sDVE4eKUvU5FbcSn74QUQaFx6hz+4HoLJQ7ZR5GEcvjMZCUP/X4jD1IPiKDGSIks
w6bLnB0wxZM6x1CbHm93wF/72tsqEuGFHpJ76G4OWGfJLpm+aY8UV8LEj4+wniPL
yCr7pRxoTZY5a2iGHzvOpvLe46BV3p06tmxAUmROpkas4AbQgh6MGaJdpD7icEDW
wm1InvbWejGv8SCB38YwZGqEYWc24y5UFGv+qkQy3p4yzpO5aIbD9vZc788XWH2G
yQ+ccLJIN/Uvl1IigVUxUWi3PQeqZs8LbDVaiSzUYoDSExmmGMvftq/f2bUvbXUL
BlrM1WlZaZsDavKxtYWSzJs+286F4S8dgB8UjY20M4a5zdZTAjxhFWVuO2HctEp8
/hERuFSjwDr/IWU5twH43x0v22363BhPN7nvPRI3eMC9IBXM0+QIpqhk0fkARDQX
BFIw/uughWxk78+fQNxfi93YP/n03SXphclz5K7pWgQ2zsCsO2j2Q4mKMkxdDhb0
WfNq+Nuo7ER3oPyhzJ21ADiE8cgJGRv/VNxNVHM5SDzgbd7TKPvcpAJhZFtoXvL5
49KwKQojyUJTrPTq6zcv+FnBM/Xpyb2RHrJecGonTnm7FlWUE5yvYHTfUazwMB1e
dNrOJAv5niqjwbtTN7o+giJQHceYYmyWX6lCSeP23pPIssHZDlQGGMsClXIlSeCz
NahyGThMjeW4YcN9O+XPLvNoOJeRJLb/Yt9sxTGfnuw6dOiQ1tRbMO48Gl9cQbaV
u4rhOnDnkZIs1A4B9zjxAa9BJByaGwaoMLCkuLBlhzCUvWVnrGy3zEJw2PJ5rHMD
whS2XlEwe98p7y3iAGo8XThRuDcCfYAVDOItQz9vItl2YWBVCFyvw5lXG0LbilZS
Msb7CL6OHzGFCsr0Ze+BqX/SVHV8hbnvr8tMBpBmF3BH7kQdxqp1sXNKH2Dgc9zM
PX2qC/E2vebf4rYvAT7OzkYsMJs3RFO+kC1K1AVpKTt98ww42XTaV8UPC2YSI0ks
1oB4NfnX749bSzrOHTXhXLK0U2XFLaNsXrhW9lPbF8TX9vG0IJ1WZ6qmdGctppzv
vgyLOHs4x/aVkH1sU0rIBGQNKmMWjtP0E3wRu6FpIrRB+cFGq0Gr1Ai5pd5iKMAG
pyXkBUf9wAF5Np21oFQ58FF3FXV4oxXK5iNxOEp9xrsyHFHKMFxYe59TjcB5oKBu
u70mrwhCvr5Rh+HlXfwqMuJDEVFj7/7Vb4/nUl43JxKjqA6KjSFRIyNRNP+XfFMQ
wVaZzX5YN7R5Q+ihGTRK+d7PHOqYZ4ziNeQNMk1Op683bYgJr4QtsRJ8EFa8pRj6
SgrOC6KtvCTilvqOv7DSfK95X+JDSMRQFkKotG1RPscQL0JP9VTUrxgGvpeAa6Fx
gOIQDUzE+gyho1JxwhlvcRUalldyfxtwYJQDhx3sPIeXKdxr3h6V6K9ATFliR6Gf
WwRLBC6C5JdmVc1qychQUDGJfbuLU5KVZ+F7o+BEVNm//IA7TvF0QTeq7uhxYguS
h3E51kaUHKMFAbhcjtNcUzkgIOKYCTpJOVkecWjMbFL4Wic5N6WkYBozNE/BPwqj
DUwUpBtkp1KatRlVYAzgT8SLw3VeoPdNDu8B+eZ/gcO7UKoW/b6hxnYuRDrG3qT8
McYNOdO2M9ld/bPgrelvPn/7DnXe9TkFtNrVkYEL20sOvvXII0AaRMuPOLGCHVFq
8l4MG6B3hu93ib/Z5MMzz6JKrm8tVoj9bUmajPXEgjrts78pfYyrBGgQqqaDshzV
eMMpsAVm7rxXyAFl6lD/1hVwL4kcB7pZPmegdAbp5bwpOcQ2zm7ShC4CNK9m0eSZ
VRoxGLBomDkM+1IenzxiVKuuUxcgiLb8HPX/gW8QOSAKKeV7RZj1tTdLOFvXg2RA
cTqbSmcPCPAB0+EGhHZNRYgFV2i/wU06tbhN6jcU52wMePBIwTSc07E4/f+uXf51
l7tKmXbaXDb44642YqPOPXAEeLQirPEdysUuRddvclzmV7R/unJ+kB1VhhCRa7v3
hrYJh7QZIfLythDKbcQi/TbrReKFJYdpVpoTJda0N6PaYY2qkv+zHwQfREjK0QKK
Grd85vrIo9QXY6kc8dJNoUrBUxhMDgJv/TNJyH4g1tNWaZSEVM8lYXXnd63C7/qa
6m5ldwuhQQc290U54DGVwTB2MrF+jjoHtCVAgPvrI9iWOB+6ezyv9+kt87hilvga
cUDpidXMGFa/pIymZdWEzQuMBu5I4HQuGloXHgxEStAcrU1Hi+yVbAtqwDBWaUww
HAepvLcQCeE1wpyuFWSv9eowsPuMj7NLx+Vhw6BA4O4QKrlLHAt1075+3Z7+2sCU
K0e5y2WLzM0Pq8w+Cef/e8UgOtnxaRqe6TV66SXhi65t6eyf5cKRjznY3+PLh+6z
ZYlb05JDrBrn1gnvb85ibN+syodzbnd2rjzFH8igYRxEzoby2ROktB32I5oQ0fPf
8ZOGkFSpXn851rT0ODSUKzzEHNLaxSQOlN/Kbe141DfAd6gxvUOdhiexB22h2pGz
v5LJ94lTqWFrk3UMPLtgAYTXEfuCQe0CIeu/7MO06Jo3u5Sz8LWJgkPfI+/wPUP/
k/vyDwfF/EfARCpA3XXSTQWq5c9ki+HLQhvx2/Hh7+ucrNRcbDwqyWtiGwFWic1A
pw/7EPunnsYJDpgRw/4ksGhKw6M108QOfhpZF8N/FGyZEw55fqhV8mTYVAHtK/qa
jW6Yl8XmDVMod2yGMCAiLPfDnkJ62oG8P4ZNIT92rI+DvH4zNHKX8IX6HID5NMym
1YuvQ1b8daaSoqbQbhC+cywIV6++CK0Hh0Eeey/XSYEWJc5Tnvc//6NFDrcLBdSl
3qVtvgllNOcgYMk0JNNcFfRs6STOccKX/Wc86QsoHWYc2u1toOM2qhoWO+iufelq
R2m/nTyUQ+O9MLVlgwi5gb5Bo6QQKsF6b3AaThv6PvtO8dwdTYYRFEtQYMj+ZB4J
vvlzxDdHtucQJ0n7fUZatos9yA2XlYCEF6FFGBZgOoH9jqxZFtQajFu7E1RW4AH8
uxI45fr1laoGI6BzDA2R8I0Iu1zuLuc/EmyxCOKRl7sD9wtPRKZk/tUNLVrsmoAS
Fj6KljxfV8sLBsn3ok0A3pXvqctVL8axEvTkn0KkrZGkoFJpNAPzLceWShzUPea/
oDTpqp0QGC/nRwEHmU2F30F5O55bQH3HVsn9kwykP5HjFXB7GvHNuzlHQF1dPNWa
ma6e0wskK3au0L7DbmN3GQudi47hRyFxqNaXPV9yXwSKqoOhqJ7WcSZSbWDlzqgf
+DJFk7HAUlUj8IZvn+3PDwi1CB7ZVROnVOjmyCoIMV45dFdOXRk53t+3mymQpFkO
DUymY3SQM3Yjb2ij8N6fsNeK+UIMIAR8bsQx5ZKn3gOsix62bfRe/Jz5GvY5Jgyh
CV53Nzme/FmDRcTBV2JXi1qarLDXtEsT3iIuvW1negUx3v4MQi3+aqZjWi3CwFXV
PwoB3UOR1LAtZk0Tbtv3iWwchQgyvURadg0y8CNRW4Mi0N0+HXxQEraohNtVaJ1s
CXnfafW1cZM1ANibbol00zldg0toypzZZAi+AP5nqgq3sP4EGhxxJmWlUoDvskDy
vSG3jDgfLk0LhKbaaj3zVdVmRpmgrc/lrp4H1OZ8HSkfVBUkEJR+QLdJnxvRUZ4S
cFdT3NQRSUtBjLkgUjoPOo+jPGJA9G4zUMtP146kNX5DRkP1ORrumZxQbw61RgvJ
pkU8u22woP7tYKOUZDvAhuu7hRJsBJYSFcPSNZFa1qkUYoQ+Xemq6IgN0WX/lAM5
vj56H6RV0L954C8BpQAaCA68/+d8Fy4oS29nqBABEC0pUXZSmZG/wrxgERPUMu/f
+YXdI3H69dPdyZs9vpSqSMSd2xm5Jngef6cYygTvX8KvBY+ucxBBuUhAg5MMOCse
u/hpqIAVYrbs1dxx/hTUllriks4DSciDH8M0omn+CEhQ4ozXKBcCxFgmOvDDKHun
4CGsSjzjwt38/M1oXXUtB3dwNbGfRKDRF7lv8d2VFItlSWWUqLm8ECfJsMliXgmU
A9aoLki2FlaCX0o8gkIsz3ib9rXXw2YfsKw+4ZPNS6F8K1oe/U9CWH0JzjYi6V4n
yTJpt4fBNCpWlXV8dQyZ2KuMt/ms0iZ04Q09RuB7vpvarhS35BwpNvtcZAeWx+Ds
UMRxGl8BoWUEj+MXeKlXaScdY7nRjrNKB+fMAIls621ryVseZg+dGkr4PWxLqX1z
/EJuj12rZtU9bC7WmKzINihmitliyefyrjv0inUyzHsrXBTqKIWdoTCn4J1MNKPA
tto9OBHkCFkIwl8Pin8dOWedwtgQp8FauKcpOtqq765wQ5Cu8B0wqnV0E5r9fZP7
KyEgGRjYeW/RXpmX/wzfECtOdSa3YSGrKQrVRA+ZR8yaCqrx2FtAzBRLWH9eXeDc
rpMvt9Gs+HnEH0BlHQUqRLYs8m/X+AKoUf9whL2g9G2SCRjPlGAYZU5rTdeKi2v+
0dlFIUjU38+XIWbvehYdELUFscMUeoWpvHyYrO1EO3/OrkohKmoS+gMAGd2AmKnR
8PstqmkBjOnRD+AetO/XQ+vK4kjPEhnCtNPFtxL/MzuP7CIuuJg03gB1u3hYlwjW
ksBDcqclBI+fV1JTiLncgE99PmKJ47G1pvzimjsR1sPeWKGj48vxKr4ueiP++NEh
eaOTIkvVp9ezH+k/AIGZJc7M56LYXRVWCxrmomY3f9sh91F0MGjdxtlNf0GtuIl0
iaO8Bk9Ppx4xrPyYKyPnoPrk+qqe3Fr2TI1UGfv+Vj67SIRouYm8LmuJkBUV8VF4
akmd3BMlm29lrXhY84J83P1IbC4krpNhvT6x+5q3I7gFMywPp0FfegvNUHPkH8Ic
E3CztTlURIHfNiZMJjQueCcfG2OeiaRm4AFCkIoRI1p6rntO3VU22jFRkn3lJyUm
JwCO+XKoe7b1mB5S6RU+tlxZHKgsDui4aa2od+wv8g9pVMIbFM54BB0wGnUI2Vcd
mX6VTTUz1s8tclvKHChxptjAdsSU3Th1qXv91xpY3q7N754C62uZ8UInWuWRVamH
xi1odCQvi6ZBz5B9NSr/jD6vBrqFfRAUDYFgbdAcEvMIzGlgBVccKH+9ZNEmEty2
TeXVbsFHZYPoPjXUnv6jg8p3xnBv8ZF85+lv1FuVTVAMtlRkTZtoWEszux3tgUWq
dyIFRemlIVJXJenZvxAL4A9LtpmDr94KT2aim103ztDQkV4Flsj2NkGnxigyvcVv
wRypKqIsZ4QuaWTPRw/qdwUGsAxu4jHLxk/1BYThdHE4HidCuxpJ3GbcC1bVDVDA
kAiGiOW8kOFGOQ8EC67547yC6d12hYB0BYedVyGh/M0u/duQ9d1cCDhsQXgxUPVO
mzGjiIVIYIl7ttX6cnDw7ATeRfj/5eQoywIkgED0z7zJaPGqMmnpheIoJPcueJbk
ej4XXNyEctNDt+g3fTrBqMkqhS51qCU5XUCX+Lry/OGDz3MKQp2G6HDjNI970LUV
fc2panOvjole0cVjyrmgW6VVQmufOJSBW5kTnAU7pP1q+XEfdBAzLJD8RL2Qoapt
HpcHH+XAWwv33CfjEJZ/che86JAZhVEmn+oitVIFGLtTHRtjY39SMDPMFuttR2dT
nOy+11fu3zQ87Y1iTYQ/JpfkiIDmMBbOSjzoXLrPvMGQjKdKAnLL/3e9HYCyq1Zu
cNz2+ZWsnt/RP67jZiKV9gT0YI+91yaiLfXmK9nomv/6YwxPk+ITKcqcj4Qg+PuR
eP52MJBj+s1zMnGUgg4W12DvyNllg8g3Ca+py0HM+gRx4/73vR+kXutpyHV8j9VL
QiwX4QHvSrdgJfWOuuVvTtiIqV6FDNNLwu10I714wO1hn2GAU2gSpEWJXDs8Mtd9
bM1jpCGkhc0S0sIVOpzeOYkzBCAPcOnMMoXrYVM2kdL88p12CVGkmccn+SmZS+ON
G7Y6OlcPGTdaIBQ1/HlV9Q3X5Iz7W/QUv2aY15DF8am4nG+bcTEYRb60GmmRfSeB
uRcGNV6LK3aL4JM913hQ0jMmQ3MdeXYU3u7kq5L6c4ZZLDEGn6lNYEibYpDG27kf
gNKWj2Xg/+kfi9yec/mifzW0rIDkpkT8DRXOtxKhN0+ENoddgEVsFAWkH67AfS77
wsGppU7ZjPfV0EiEB4nde3ba4tCmQ4GvHNR1uXm7jFAiPzo+7mkkpE9hG3yudZut
MQcmrd6Ju/qfHIBL8nAVbq1NW6VkJF0aduwnGNOp5W6+ToY9qwXR52j0wJ4T4rT5
56IbE9WylvY+WdtP1uzH5fTNaMFQbbAiBK+R39U+Gaa5W3vl8Q/iuUvMghCU9Gy7
d2Bynay/zktIhaNSH6mmor4vR7fQxapEb894CKdTAvImbLosbsvhuUKJq+UWeaKz
Nuhf+SErTzE2V9yXkCRXI9WgYtYQmvKQMFpWnPgcWKvqnMXJwXM7MFORKdtczNpo
uWNmrcuoi5+AeDFuotFxcOeGX3e+gHspUUfyjd784dPv3b2oo2Fhqnd8eweWZyaL
ZfRWjvzSa0S2J2q53HN5TPTfhRoPBd0bnhAnJ52gZbBVY8pRQRhncUR1cmJIiENu
BWid9bjcaLmJVZ70S+zY4wMCC1MGZ206ofXRTG4FiNh5t9RCP4nIw9tDtZJiy1Lo
r7wNFiU7mKmVkbkhc8l4d4b0GBSgSxQjEK3l4wiMpTA24vI4tE7U+jn6QGcrZDYU
KV7hnGovOo8zpukIOTsuQ6GRJd6cJ13NUHJBnyL8/os8NtKybkWFR/CBDZc8k7t9
LZu/WZPGfOkEt0tHpMW6VPf1YDHC4dVG/8egxkc+V3aWGCcMLOyo5GkEItIYVYJF
aVVI6aD9TSbgK1yBNNQF4o2V6Xinp4npqF2LtY7TUvrGUriukx4TwP5Tzo7ItVab
QhQ2o6/8VWx2cPdfCkJ/uFonXXyU9/T6JzOm+5M9I2dTBIIqOnijAP3yLstDlT5c
AQYIMCTwl39BAWCGx6tyoHxlc0vuvXc0pLPbyYMuyyQXPgQUpkXJ6XKO5lTKtXDP
4dGTKrTHu2AyTG33r80//JEEjL7aodClN/Rcl6PPqQ3FBu1C3jUrhEobmhzTWB1c
RftGrYdJtz3Iur1riuDqM7/AC8jPrCg54JMUTiVbgpXsRVQJKhVespl/LcgdSVf3
F+N0+HZ+GFMOWYlwfrRDaMME+4wBTkWrpwtz4Dw4GIV+1r8xdR/SRdXOiV4EPbqR
ffxkcodnkiZc/YWhet//M5jn7vgW5M2WkFj/e0rpi6h2+esCncjArOGQ2FxeXehq
au24HIizb6vEwO0qwolOhW2vV4QorfCV+gmP3pO7utAVzFG6sZKpyeUeMLC3Ii5+
yYHj+Cv4Js19g7xeCuoD5yOUQAOgMzn8uR7APbPMfFJ5Yq2iNRxsNGzJj27wA6ED
VQCV+UDok6uSn8Ver+mIkpX9VWhFBmvLhm/1zzt483J5xLkeY+0tBEXt3WErjUGV
DGkuhPIx5ow2KyshDKwVBwAwbcBJTCS71VIFOQC268L9FYIanEykMiv2VWW0gVdD
eInB/XXvETeNcsyBZy7/8WTWum8heB7KMtP/tjPTEwYPBcg3XYnWionOLNK0Rb/g
QAKtDFPQP15UAaQ85zu1sj91v6a4oDTGKwQq0YOelbLu6X5GARNc4eQF9D9Y4yZr
xib/HlQYbwBb0/ycAbG81qFGFx7C5Hda7fjjunjJrtm79NkZ/QCA9l2jWl9qF/3f
pliT8j4UNGQntxlIJNN1YutBbKBMujSUs6WBQZPzbgiqwnC62mRtVWDfY4hE2tRT
xKocjczG1OT5pk0T08Y3KhTrJCxX7pYexCymkoaN7RwSh3Tlej3GcQNMfSwVC6y9
3GTaO4A88+9pRgd0+sNtyh1gD0z+2q2k2xIydv45FvRo8+DAsf6OjA0LKewePm7t
Ze3Ys6eSYJzZ0hkbsA/EOcK6tEubE+fl9lvkZTeo9KrPpwDa6MAFeXvSVKCM0RXk
yHsm8GMcfIQxEkvbthcHWC2woOpJFgrfPdKR0mSL9iHhiWZYH9PR7GOfsD5vVibK
D6TtsmqjS7EInOnwMiNeREjtOhbz4cNyT6tQOSP25ejYp+Ha0wTvLq/LASXbOJBB
CNYe8gQR7zm2vSaFnUUDlkDXMdYBAwNyOcxj2IeVJ4OdP7qyg3DnjQYYfCuhK62J
95bsGEEwh/eQbph80cb42xU1uzSJTTOAb5Hg4pXjDXTdxhqIcNbeVuR/JZb/kcgA
WzD+8d7UWJvDSWD4TYSiivUfxeCkEv1g05O2k9wh/ilWRx1htBeGxf0/uochsTjG
K6n2u6iYSticEt8KNENKEnxL8m8Dy0aOQ8URZ761uruUtv49z1UBEIkXnfH6FQ/7
aJulLGm3RMornVn1xtxfvKa37aTZSzOptalibg11W/XyFDxwenGMNv7ma7MaBkN5
IAmai7A18niOHmbW59yCt/ZGIixFs70XsfDMXtQ40ZCJ0Z6Qt2XuVtMe93aN4XOR
uLT71+HG8DWT3L1LqBnQqZV7ev42fPZ6IxOoj3NO5+pte/89vdM3ZL9+U8wTvH1s
sON9RyZKhI+49ak+qmNpN7FqxdtkyllIslMGaHo+svY8mH6T9I0VbJ69uF40gxMz
MnAvuTgsOImmpELoYj2iVXnEhhtTFoDoMzH28mSA7iVs3XG4lPjOw1WK6X1HxIXp
B1RHY1mHaz1zqr673/Rn6m7FbJCnq/phP80RfF59Z3nsKm6fAOfLsvBgDomNZZpH
StpUBfcBXGl0hQi1BP91B4SJ9fLraZ3PZ4MqWa3BGkywMdO79xVUEiYjb++SlAbd
HlI8odW2gK8OC8nF7Ugf3AV8+ZbDzpWZvxWPX1a0hctXjWVB6Wa6Dn+pPdV0jEHK
5Ng2uAAC1YNoo+fhHXNXyObRYMlJWEPKD0wjSQ/NJYARvB8+9LTfrAIh/gPxQ4sq
Pwa0Jdwqc2L+8hsECN4JTg6tAX4HDhrNFC0q6OErXyIZFd5NEHK8plOtSZlXl575
/68ggKouO3ciSsr2OBwBsVHtsHkp/Z3qNMmtHssdfjD5/+r4QVPMbMOTzyCHqMlk
e0T1mC4++aWxiJEwTGFrI8uE3fEtYwAf/nCQqKhtzSUe0NhzUGy3AatOQE/veL83
8vRexNoJOyYwwbIyM4RlJoLvJ2CXQUqQ2d7VOvJxsctVPLUSkk5wGcQ/SonQ/zC5
2oJs92+Jp2aQvmCAAl2EaOsSRabNHSVvIbps7sYW5UWcKX4yERK8Ej7xI+Tc+vv6
oF34eWdk79mFuYr2YkjtSN8Yi7AEcd4+RLx46x2VyfXtRaz6XjSz4bLcsp7t92Vw
bHjtv56NFcwTolOT2lUdTehAH5O1sbUWf8bRmE4LAPjgDYxVv6Q+RztRtKnYjTQ2
SoRs9EdJmr7Gv+fmJIo8OPKOBXEhfgARsr7KPP/vDD+ph85VvXu1W0q/H9cAoHkv
tCqEwnlxfLT8Dp1E7oyr5sfBRv7ZQaR/y7tXl8iFRcxgxpBgMSLBXLh9UXKl6qMe
OcRpWeZl6QoxO5t0IvQ8nDgsLqGs0odA81tMo676m5gPoPYtujbAmvh4+/PlMC9Y
/YjIkqv6vmaifoCepy6iNasRblB/qKWTKzcG3N05wy0OTYuVossHiPub8c22xjMD
niVdeX/DwF9Ox8PSuEyZzdshulYILWCG5WT0QlzoId4Hy/Vu+sg8wOpbflRp3JKc
euf5iXNZdzccJtt1VnXFvD8CRvbFBo7ulXHUr87mTkPbJn8hkiFRWkO8pWwXpvfN
P6wi3DjPwvJqjkPeDRCyLU7uZUCxfG7f8wcOViYgCzEegsV8D+b1RI9epvyb9hgm
Xow35vxGei6LlPbqtr3/2TX10RoYhxfMbe02VVEpXyRDrX7gzoyrJV0w/5Llj8Q5
iqFXUsVkJnthyXTiJsAmdZXjak7yw6wQdUdtR0Ixxw8W99zk/V33WXEiF7y2giVj
Mlw4kqyPIhVPf2NmG9ffuhr1DCQ0szEKFUR/OMIQjHETKVOi3haCp+zD/gOv6Sc6
hQHTNeb4gdTTd/zmHnY4sr1E6H4mDkrWmChPCFHANXnbgTsfajKncMgNyCs0MMiT
SorQhMBon0te8UgRU0jvc2qQqZ6/KYeuPGKASwbOzo2NHIyk0o9+q4COyYBAf22W
RUMg0GtGdL90ocxhwgX0xQFdBZcowfr+qCkSGNwx3Z8s7/pRJkK3+RLmlBxizD+M
wPZQe50llE5ZEFBTjNO4Z48jqFKM4mzdr+QoJWa0zWBZfCfjQAbtJgLOKy+B1ZC1
uxdmkrqhsalxwFcHPDJtQ9khvoNKOxBA/SGhgYq9TpncHzZmilp6Wh7V5D5cSjtT
gIDihkKckgX/gYE+343TbSwFlPO33AgeUvy/yhx0ep1odnpWTuVSq5tXEiaeNL7M
d4wTXvTj/lsY2K0kmpnpURhsbm2eeeapDdLTuKVD8WhYapJV1rK7k8Usx6z7T8Sp
zULXgbsCe0DLyUH5wirpL56QaIp1KjIOCa4DfNo5iK/wHo3PtqUYQtxz24KS26H1
nzzeZ2wuOvGSlUmPefGpEhvQnVxq/PwVGOZKxgfsVgb3v/UUgxJrRgoMtqswFqta
SlP2VNjkL2cRQTVCbRz7sT51u8JHGaTyLz5RzFQlwE0cYlNgHxMJIM5w3yH77Pcu
O+PK3PFCLPP2bnnF5rS2O48FSyTe8xy2DEwl6djRnuFJAazH7y1bGgh1iovTqokF
3nW7ogvp4v2M97NShhcvyd6bz9hH51eexRAtZx+11WXUkNa6CVIQfao+Zw9pcbWG
HrkH5N9ZrEHFHL9YOrtOQOQf3D9QmE/EKL+s9EWuUIGf0qeGOTjUqeX+P074lRYG
AneNHZ6On9/F5KpDoXdtfynbkC9lgj0pRZTU/d/+VgQn30FXXyC74HlFzEf6sisF
IAd+zjt8n7uQVDGD8i5jSfallK+6Aig2AYb+QUcFdVI1oktmDJ6KydaO3MwZsxAN
7wPJhjI+QHBHHJg/J2hxO84/01e19jtdVo96+fjH1DtqbIwiHO69oWr7+bClGiQK
SWWPkUbmM5In3STVjUwPGTK9JKAXG/GvPoH1ZPgbWEVZRWTnpi7and33S6jO4End
DnOPf/ZuZMXBgiE/fKfut8LVQWc3+RuOrxrJaEG0NV3Rc5dqSFCCGArt4wGltN3n
A+ojaLAkYRqCtHcL5lE0ROSN0J4QzRWwWbYfQS1y/mt6PZcQdIGOLULlTbJRjfNU
4FjFTZ5izvMZVm7gvl3ryywJUE20HYCelYYgtjYcZc2q3y/7OsLZLIhRqHM3xpTP
usdzuafw5n2PqpBTa6ZNceo7K9MzRkiWalxk5c/R0MiWEF5GhvT67N21blOgPbmL
C5c4ocbYdHgc8xZOLG+Da/DrSaTmLcVanAxHcL2hxp7Di3y1s3Xtv6L7slQOn8Uj
qxULR3dfQByruUOd7X2iz3HpCmqiC58fsmGTkzvieuNxtc9AEBhxSb62I1KVSmuj
X4gtehNlREt46B83ifyjrqkmYzHsdhWxGorHARu5wo9XGb5NzD2ggjGWyR1jhsEp
9SybTHVvZV2Z4Ym6MV7dwb6e+jGvWLf248gPD1ZkbS0gqgpR12be7G3iETOonX73
8eaYUt1Np+g2areNTYPpZTauaUQJMj3Sm7917uev6AHs3fybwFwq3DLPwVycsHBo
uuGNorpHbqLD2u0OtyYCRnEgWol2HMHzmjDlxgHRCwhoUgSyGoAlHocrPYco/p4Q
kI7/Qb/gjtHb4kWIstNiDVbBoZygvALG4HtWjBBkQeNHh/pkRcm9O2QBya3SjomK
vWbIxuCwP2WupXFBYtQCqicQ3rE8v2RxASveytfuU55BquJNPGciMZwq2NlZX/JS
ro4zoBxX2/6JWtVIGoIiJjsu80+XGo9mDCEdl+gev9jLSymWJStZUbTm5GQH1DOY
AS8v3AKeTfOfH59VS60+ZaQ97QIyAyy92PUsPVyTfCiRmmgIEDmmVhdMPQtQIF6b
099klEn6JWn98eXQ3G56UPgwkXNtHnLt6OUKfQJjyvvVBGT+gqKCooefSrS4qGJK
4hRy9owoCMFxL7y6UMsv0VkZprB5BBrqX1Xyglk4pDM2I1uOg2sw9Aw2yixlt6uH
OG/dlc4TDgSV3V55gznY3rRcKy7ILNfOewzmUidkAvz77zlrJ0kWz8HUjC5xypfO
zw0fsAbijngif4RVTBlaSjBqOHVPNuDGGk5fHvbP7ykHNS7uRJDjZ7uZG/XkvI/l
PCOgmn4As4vg+B13cfaKRLwid1YFueNUXZBqx2/9AEQgHvzTZhr3eSC+PrZAzqBL
UY/FcomO66RKwd04FPxbesYtJRJAqDrBgcrGVB50sRZYxa3wx+qwEIo3VhZCK7g3
JZZjUFpiaxkqutWwz+ZFnia9RXqXbiMn0Qrhe3ir9gKQa5hJbbj+58eVOqVJIgBa
ltnsO3XStVsSELNMVSi+vCUNur8stNe++SSJY9oYy8RnqT8TMQcIQXvjIZVUta6D
n3UX5CvMRXRisNqD2MRHk463PwPwx4sGFKCdU/1Yc+HCyscMTFOg4aoMSbihKfEg
zO9fiL8CS52GDUBmusHsvPkZWr+XwhFK1PNloSTuRsQTrTFoRbNHwl9zK5VHV8i+
nBv19oRa5Fu2yQPWBfN14hCK9mPayFpT2gOPB+4An2wspuVbNcVwVQzGQ8a9mSFe
PkINi+yGBA7FTMDOV/GcgPv/4HBvN6dIsPSSr5L2xupZL53YnsQKrFmnKLF9F4eY
xQ7Ij4/H/pVKeqrM0UVHU5627blVZLOYm8V9oltUuJOIGkaMIN69fXHvW7VmGTH/
4Qu5DC2T87bl8g7JMVaHYTjfmsMk4A17EaXQVkaYX8TzQ1ygeBXkdnzqEHgb01pF
nTXPekzEF2itGFzdOuFJ7n7SzaZFzKOQNL3+nsMA3nGbSSOxF/BFLlDIMcJfdarm
C2YFvWGsVQJK1L+MyH6FzWwVTMnf1XI3Ar+ivQZt1eZuy4GrwY8PODBah+NoDOju
BQVB3ttK0HqdvI4kReXvKE6VV4OABZ8XmzknvflYDQy8kdgMwX0Ps9iaTzlga0Iq
NV6rAF0X1Qu0nVABNdb3SJYHFT5WsRrkP/Sulljf895SNGIiiJJswCwD/bZVQHCX
2zaNUcJN7MvQjNLCBHdf74djP3pSaCq/RpEaJbhI44SRKK3Avly8wH99T+FOp2RM
PCiYbpxF1+gbUkDOIsSnuM+ayFJMLoxHF/aX3cbWJZOv8PbDlPP3yrTzFkve20aV
ykfN/Tih8dfbziXWJAFbmbRGK3OA6UA5DjlOHrOCc1VFD4colgR77Iqty5MRJPAC
q7HDswiISzusRIbO0tgNoP+gtgNB+WuLkhHBWC3hHS0B0gu0tbMGC2hLIcZIokEb
96wM5EA0+f7nBcYs8rT67B5SXvpcnfzkqWoelUX22VBPujOKqCJh8tRkloIE1GS0
mZkqAy4z2JHwmoYGrhYFAzreGrHNJZ37yvacxAE5+UY64y4FfXwMVaZYpVZENQcy
atijthjusdLpaTsnpfMYXSoKRnWKESlruVK8ySFokjMhngCG464RPTrq+SHqc2yG
tV9pqnWTQ9uV3XC00deyw0H1DgQ9i4c8XqlPLBzHlX3uCxAkU7Gom5uNNYlfUx8P
2MU1YWiPc/OSe4hV6bgV34l+e1CymIx4K/KowsMg9GYKZcQbGE5ymL/ISPIQCraa
KcRnYEhd//C2yqg8Azo39ltwnbmeZwBReOBtTbYZuhUcuN2zV7/iiNwnLKqjXKqg
vADb4s2G5wY0EMvDf/Re1sUguiLe6Ch9wqGk/sZoDEiSb3rZqeWLC5zAjczDcQ4A
ucDpYLa+dVeW9tKE7fW3HkMpBnuhyTL83/A1VsLw0bJVwRH/iIY1VQqVytshQlno
jPTMCH49iC4dfnKpiin2S0eWI0Eiue541PSvVHKMwa+M1wptFOvrE67Js6hRYM/j
wswjKKAeXFg42Y7qiEMqccEdm5ujHnc9ULJK5r4bpzy3XLxf7we2b1kH4YBXMyvo
bN9KP6bs3agPJoCmKmTYfMxMWYCufC592goPf+ixbJnrykc6M2Ny0TlSgMR4xBOS
9+KhWguY/8cGtKYj1Jm5oxLbKga1/7f1xLOKhx2336EjNto2pbkBJwP+kuhLu6xw
yOy6CwzO6stInRjty47M1YcIGgTFzYpzKOZiLmIwQX8jNLYAsetxWE0px9ABSE5J
Ky7+QzxtveERcMpFHJ0DbYiMZ90+S2KodiuUnj/pxc62q5qygfjkLHRJImPK9E3U
Ks8/n1bxZjTVbxGMPTRpT2NpAGogcZWSrujKxSjl1xekMKOFdoM4SJZqt6MWe9Hm
rpSxOTgOI+FPWzGUwjouUGNbDhCxnDYy9R5nv60ExU5aCCBXVrzEwouYbcPwsXp0
LNWcXno7OG5ZPGDKUwZIDBLKjaUdXTAHVTD/SkBCD3+QPitIcgs3kHM2C3V1/UCU
Gb+GmmjbHB6I+RqNxptmykVA31KbiKF9pZlPhw8yiiHJP/zWvyQOo2qUefaaeZKC
WOLIq/acbQBZQDGlj1j0Y3Izvew6KqSke+a0gJdLO6enYUQCPc/V/IVIPbgoVZ82
R+NNJdaT0g1WlaYH4ZZ/MpLdXEUfd8Qm4A4myllsRNJjtv/qXq9Mo25d5cGjNQFO
XQCKuUeVCnZ9vkinpZV/SJ24iP2AVTJQftVmswMBVHDikcpA3jeKRoljzsxmcqVo
2IgYZ2+lTf1FQDUshQUjePWtBQxvKRd8scw0fWPg8ZuKQVu0IuwQO1nRFsCNPG3y
wzSIZPSTY1n2z8OsvEXs0pSfzX+xEExnpbNU7SA7MU9pt9QG6be6DA0/NSGz4H8o
U4BTKUVID4b52BZAjNdtWYxj1V6d4/mkdApayLpCsxVOJwd/BrgBrHtGZdagkoPz
VGX0C1Q2vOZ54vxAnuONY2BYdz1FcmbJHEGB7SRkRBRLjGYTYV2O3SH+/1eXsSxZ
jDmvmrmtia0UF+VbHtwbFAWqP+jCiXgYYuQnhEYv1njyA+dV/8+L9X4xuo+o3/A8
HUvcIBfsxBGCOs515/yn/1UmeuvBK0inqvT7Sd45xxj9yOWDbFwl20rRQqcMm+bR
Y1nhnKJt2Hy7a1YbCHUXfwQ2zHtLtfVidG2YflncozpOG956xO9qaWSTw1B+oDG+
PldzeVHmvXTGpxbjc1Y8lRFW9fQodNUJjsY1lxGXIhuqCmcZTDsXljllHVvaBxMY
Hw4IhSrk8+ktz5AeHksyEi0BVdVj9PHqLengJFoPcSmRTxSp9q/mFN9PhSaP8neM
dg5Z6tuzFCTm3LEZG29GDONzo9rmRlk0eZKjBhbrm84uj7iLtzW4H2tq/tedh9/s
0eYqUjtnYdZiboAIiZH2b56c9dU75QjJkWVHfuoHltgBzAGgOX+9jmqiacH4CdWB
EZwi4HeazN4Kz8h1761gEZNOuCY1UD1ZDjmIEdg+Oxb61AgCsfbEN8CpMTaOIutd
45SsWIAKMpxaIlTFgUowc4S6DzBmF2mliBdyann+i6/UBouSgs3UN84fVe/FcK1J
CvrBssGdNjHLP/4/7TkxCHNTq9M+3k8mEmP0816mBz9yZfbLarfBwjomPbxhK/AH
m3a0Yj6jVNEfwHmRn7s6eoYF1uoBi+FnYgvR/khPxkLLsMRtTkCkTy5RUSVCSj0C
JKZYUCPbsAJG2S8aGqLQnkAgm6fDZnYU5rwN5BRkshjAn+1J7IlaYc8eAqQ/kWNR
xz68YTxCxwikYQA12EN16tNmJp99VquUrJL1XV6hHynv2ibEdeMfTK4E11xhaU+z
LK6THX8C51OLAPTfGlR+/JRA1cbYxrXvy3vc4kciyddl/DD2env7M0+NC76RJ0i+
9++iMVh/X0E66pAM1CYODFM1xAPhrc3VN9tA5s4WDgn2vGUNWCx7CW1czFFNrsA0
1CsKCCOyqRT9gDwHCyiDmCS5Zb8xKNGIxzHp2JW53Z7XmxtD3SFqooUH1sLB7FRg
yOW4+rEB30aCIC5uZXUKgUqh93mNDPfxlyCajBQZPm2LPm82mGFI9FfacywGsBIO
XAD32HdPsAN5ICmklMAL8XKPao1kWq3y/ReU/aXLvuGZmZCzveEgk0MFCmtw/UHE
aNb8zo1dyTkfc5apkBo0SpDYGN+YrORKLcqInU6/40fQoLKYqOdQJV/ZKsk1Mvfl
6GpTU0vTf+/2OuIVMiAwMECSrpiAxWj3pcm665sUI4D+wS1Xs4JKPYkTBZmUf3GS
Jgvs6/Y7b2L66RnAZTwmHmq0/Xu0SITZD8QZiAO+x+NdAXS/ONtPCQXwYgqm4+GB
r34OcGYfplmUttDHBpQxGGgdu8JiN2SAzQyiDhoQanqAEDAM8h2VR2jwrYWTAKWO
MI0QNNBbcSUcl8MP4SCl12AIhUb3S+08ozFjhhX6oD5mkZgN35janQsBK0pkGYId
T+0iGiCBGA8V9ZGJd37+NmsszdULAS2ejdr5A++czVZQy7SZouEnD5uC9w1fTKmv
o1lygiOT3My1NHPqWehW6pS6Pbv5pnhwDncGR0SGqGRdS90quMdbyLlXgj7dJZFF
PlT5gN67KyWfk3CcLef0RemZNwzALPcmM2eVBMMmG6GLUpHX6PCrF2lAugNoFJIj
A7KGYj9oKWr+CYKaDAHPqxRNbnhIVHWXApjsgOLRUjQMsv1yqfm2hbpCiOJJNJwe
SJ3JHWTGwQhd3WeUV+wsLciYDcK9hBe9FwGxcnkTb8wihXFAPct4D0QOWzNONKca
YgOM+FQGNlqZcmcKG+S9jgMbIzgOgGwMePIQXEMFASFrXrPc80sXN9+A/FTuZYgQ
mQSrDDJzXLdtfINR1350R2ZtbMBwoqa9EGoBL+pRH5Ac/RJi9G6mQXi1r/zA8V25
jYjr17XlMEuASrILB59M8F3jfaZiRKHZNVrFIjm0snA9aL1eO3PLuY9BUwnztspq
ie1UOi2OJFOrOyDv7IM6FlBspgg6m4gPnH2kc5q7up8OiUUJotiXz6y+ICaIhXDL
3YjfE1A57nkRF3AqBKqh8M7SiFPtShBuqSFQK8bDLvty67rG5nP90bZfnIBpFdZV
D+7GUZ1xvS63euYmtgMlb+tKLpwvNh3+3+o5FJmRTu4n+il5Y5HwMD2U27iF8wDx
Bd3K+kM0y89G7dvRXdwf7MsRZKUR9l2i/nWrjeTENnZwouBMeg3BeOifPNtH/WCb
sTK58+NnfyGezVXlwjkxH2v1oAtWXsi2k9/oRMLHI/1ua6VYB27nyY+bY+2JETQQ
XdjJ5Z/k2M84ukV3r5I4T0F7TltbRk9cqoFhxmy2XvtHNrDdfU4ACyZak2g2qWsc
36qW2TnYroPK8WgMTog3qKFojJ3r5kB0hrqGZtcp/8PTT6SL49XYQ6K9nxZoRxk7
XoiTQGViU7g/H71j/+dpHv8LvCIzSNwu/aYDd/G3nrkbdGefYXVAiJUIjT6iYExW
p7Bd6tjs59U0pJAmHktUKyX534ZuM2Oa1q9RTvo/6PnI+1CTnua3IgCbV5uUyUQy
LHj4ERVDfhSpz3E0GSeduB1n0cIzEKALR/QucOiKjR0bFo/JC0jZmaeFIeRdwjfu
Il6Ve8596/DEOsc83ARJutwyZeoF/g+dD2g1DGpltEOl/pjA6I9/iAVqtdH2L+li
n6SfE2u0QvpsFWseYstNkSBFq0pDFMXB2pUatrg+gzWNCmKRoFRjbDGdf2xX5KEd
pT9vng1pChW1t5c1aZGQFFN8rGn/IryhwbKiUr7Oqsam4kLdlKvjrJ1IMqUf1VeD
Eak6tMaVORUScohZrd9JfynMg5ANZhVcvSWuwFMz58Ttpa6d4kRZfKKKgU8vgNMi
bB0FXsZLE2aD2b0CSoh5mdVtNhmUwMAjMQm+DgLCVaKPn4WTdX/DRHrK6PiwZ5o7
NQH9fFCMZ/z0cyFWIYI5c7eDQHRRaO7Eb7FYG5WWdN15bcSdGc4tbxeU8+58T7jJ
4pk0f+/3ZpNPH/ZhNJndnX7i7OnVpgRZDu7ZF8ml6WsvA6Gzcy0QwOKgYm4zOXmy
32sppEBFF+4OfMN1ZvjJ8wh+VyaD4Hh8vwuS191H6cUQ2mxeHF4UR60CO2TlvFop
3EjpO2fO7Xsy0/1V4QYi/0zVqzTfhcyqEe+pH92n0jxogGMg6JdeikY8dY8Cg8hR
ELo9zhE1GjVvKsXGNcBdfZ41UNNlXka/9iestWvxyzQ8oYG1clVbI6PKHocl0Ij9
dl6y6XvgVMYFKp/lcaIGo9pZKaL+qUrZySxbvngXn1d6TYGaOutV/Ns4Bzm6uQuY
vDo2X6XYguAlOM6SQuj6FhIWr7QMSew4VvB3syuUC0Gi/0JAgUCv6MXZE+TeHioE
KyUG8LC9TIofP9j8j6OjwyHGd/5drV/4s2spFRnzoWga39vypow6FaJszX7edZ3X
kzZGKecmlpAK8CAkQJoM4sIMSpXwzNnPfgwWib7Vtd5oTKkW7mfF1PtJPffsScrx
TRxl9tewETSqWY42pTtFZlNOYtJvKQKznqgNPikDeV+5nenHTaEDpz20WPOdiXXh
2WoqCH8S8N/LbtI5noeax3nk0QSOrbuqH1vlaeW0itR/p+Y+avVhElY+8dNO0iUB
KynbRtQHxcS9h7tqZHmder3Uhp5HsDOEp1mMdLiAkCZilHxLYRpTaPRiJWOKJ395
fFMMJ45Ev+Q0GQdCcCyLo1E0wr/ghhOP/SBR12avO4JAxjMaOnrGkechoe6PU34Y
p6/L7Iy7ctJz5CvHimdqUnfD/qFVbeqgGww3oDn2Rw9tSA35QB+VxTEmpbdynTqP
x+XPgs3U9bjpLllcEqyHB3cI6V9AToqjm+9o7vhzmqXbLC4+wGH43p9FUpwHwonB
BIaU2A7eeBJeUppIdz6lE211WwCnldbAkTjnXsetc2tHyDxedfsjFto6Mv6xWCix
Uvo8EY5j5gY43Pk6SzrkdGje53kCS81cXUOulbH6B2dbYdNWrJT/jNf5gaZzZUK2
JCgUVywD0He3imw2rKQ4U2mZ1RMDahAHFiUdBCuB4DglbfoEPkxL/42K3/YAvUpf
OJJhOhb69sTN2LxHkDmIfOopswFutlFI+rh5Q5Tsryi7jwG3QIfXXqrxVXtPsHbn
pXMaQgiuXwVzIwwzRWpwuop+ebnSeLaJ/cT6hEeGk51rsOne9J7bf8vbNfnrJMx7
I2jDpWNNH/+tZefY0xC2kDVCUvsBMt45O3pKHN4gUAzuYW/BzHFsJuzsLaEx+aE8
sgrzKUjvXexozr9sIaB7yucUyUm1yrTgMErOULeItKBzV/Y6Cny+sQ5/v86lKixA
2a31lvraB/qQwBfW/JT1AM05YmcsGOUC5qlGH6vPd0kB2IIAd2v25/8gQpBj/XVo
46krfmYL7G0dabAabFz3vcVthaBFHSd7g18TuwQrAK9zFh5b2JM27SbXktM7odPe
2yvAY4NphdXde+BJxzbPSKXLm5Er/b7CTmPoufHtW9+ND0nO3D2gga5+nIMKnVjK
i8BKiih7cVbt5iSFw7JY8cYo2TCl4XH0EBfPIFHtPjn/C+M8VEY/qi40HObnIFGq
wjrfUs6FmQb03DqJs6YHXoa/J61GPezgF3AfDCEZAIoI7OsNciD+VPpbmT5dRA4K
EnVwxBxI+KlOmfUsQwC+o9tiNkLxpHQDce6lcq+FWBrAF3CrUz9VZ/L29XLzBXGg
zNd666IclOipFJgT3WO+EC02OoStFJnEirE2tcTLWkVQniNMT3qzXA9sUhpvtADp
iTvNbCSYRA7OenrZRcI4llDsD780eFb/85PXbsGeglWKE8EMXXPpk9UvYDU3byGq
X4t9izVTW5+1b8BCLHcHgcPx40FIo3TMlHyqQ0n1gQxbYIuTqwadezCawuaucx6Z
J6Sicz5Y3SFos8hUzujYU7WJa7no/gBBXPHuV4F1EbvLyrVARKc3wGxAjOLdfTOe
W+qwyCHsrxRmfYU3VV08Eb+p/zTrjfGzHVsat8awRztLm/6w3Tz28MLCQC2ElH+O
o7faeviktmX/OUhdhKMj/D4SDxPVR4k87L0iMtyasatJNZM+RwB2ncB8OSiKKW1n
CMBE6isY692xBjwQKr/5pAXPksL9M1iznQbh6qo3lr3Frzc1Fqhzyd27hr5+ADYA
50/Pf6bE7dYRjBVN0J2U5B0zL+r0uawOL0zpzFR2ikbzKahcyuf73GLVPbyr+4Tt
ejy3UdyPMj1vWK2aO9tsjvT+L7xgAzH7+PEtIm48NMgGO2qZkf/2NcSuLVb4RCoc
v+Oz6m8bbPsOG775rjl0JW69j6RlrJxEWr5YqMgZ8cie36j4sLIexRSiyUekqoy/
fcQJMbhM6B2EzIrjXrkt1RDFE83f+pttNtFKv4+1G124RmoMFfkNjKKAeEr/KoBt
7X+oUIcfByK0/kf8bKuEx9ky8mb7i5Jm4lHgduDYj6cxepXpmD8txollnYZE12tp
zfAcB1UJ2OLuSd8bIWqMqllSyrNVC7ysD9kcSbRMix8uffnyO+r74elzB68xg8T9
eHAbwHH4LJvFAMnxpU43neihdfUlKaH9wYN7AkESdc9nI8wrN9wZntnmsYDIqtK0
Rp3HyJn4ipYnVbkowFPq6KQnLr7aGRYyQ8Pg1kWzbCzRKG2kZps/18Rf+hipuRnE
uw6t3WPcRH7B4CMpeqmz1XUBTLid28iM+g8+SGXxoZVXPtsBtZkyKTWKv0iikHfo
iWDPoqOgNP5sk3ZZL2fw9ELLjUHTqHT+iIs9/yBMNiTJt1cggBiFWlE47boZOGmj
E/lfS8LO7hOsjUTYHlcMAfGJ1UW31EQbmbpYogmIrYd+nQB2NVmueEjXzv2EP8S1
filHX0avzU+wZV3fyhvf1WbcXKnhiZDhHJl84/XBS+3768xYxGRDNYZGzeIhsz5V
El8dhlPhlkCVQwXR+yfN7IHxB9jjZ+wAQfpc6I4d0KlR9vKyxX98HmbvNKqC/Lwt
WVLWR61Df//U1yJttFO4erkNNOQMBAvSslEtb+4JMDhUZjqfJSDkYNf9XFQonajO
JBDeyERZfXz2rB7t9T4zdqGAGN2ca9IaXdd2QQLFACq3tn34oKT7nbEhRS1vmGUO
DCID48kovfm5HtbPj+VszsP5ZT4R+bbYTf0lMFK3HmoqtkaTLiGC0p4yqumCPLNW
MCqpsgeV1GzbqIejO2V1mguXqQmInt6f3+MFwuglrN6t3AuFqQ5PmeBIExm2n4QT
O95W308GbM9hh+ZJ+QcLSMp77+5wN9dXZWIK/ufmbe7dGHnP11sd7UdMc5M0NQPt
QurnUeQejyK5IGt+vAUv4F6zHFbE6PyZszy+M1XisQnzoFR3TCWcwziYPZaClLY9
OXRFDUq7iQOsdIPT/6jyKuUVQ33kV58bhfgtFT0Bi5G3NwhWtBnZT9/SkHtC2i+S
sdXemiNpcNEbhBuBWeYIDaI2wtkF67dUER0Y/NGzSMr37SsvVBF1vzZ3lMAy7L9q
tDRFCx7yH+FX6lCtgQaEuKaxLsE1tQEMzir2LcWCusVWMXihG8EcJaTlLhh7TghT
eJC8dR3RqTafdW4+0HjLuZwuIRPzazSkPVuL1deNt0AZvUTh0SHACd+n4gFPPX9M
NDzYTiVA0UZgthOsko+e52maxy1DNZZBRgSyoZmI/xU/zu1SEJWN1gKRFd56MYlg
AcJPIhqlZsxMWl85dP0Y1jZLYxMQaTVY63ec5PwjHZ68/nODsy3TyMfsf2hu1bKr
LGtc0kLhiWh9PE2/mMVgliZ91AUcAOL10GcX3PTLXQQ1xS7vLydv4mAZKsFC8rr4
kIxDQcZuedIgdT9FB/aK7dYJjaRY+vy7KWhQ1xnV/dCFIc+A7Jaa0lIExv3/0tic
+hQ7nVrIFOjtCMerfWeU1tLP4bQHHT1vlUdDJ2V2GS3foX/oQbpDXkwAatdv1PQf
Px1uruUjtYCAtFi/WsxfzfIZbTb9ZpCSLZox0pK05W1Kkgsqz7LfsGyPffi5PqXq
Y5+OJhJuoJCcT2lpiXtPBCnsAsaodMwa7evpnfPbBkzqWLElp2RqWnnilCFm5bZJ
Y3/CiP7AQX6zitbQ6MIFNLXDpzSgEUbPdrFiW92vHbqPMAv5R36vUNG+NxFlam1P
eE5QMuK/YMEVb2fjRPRZXniiSpRXIWcH/fDmHX4HET9AQ3lBrxYhjkBH7jfPd8zl
2Zr3es3lD656a76HPXcw+Inqp6hSKau5bv1ZA2OFV+z8CUhM96xHT4kWwxRQX4iQ
ihzjdVtqF7zz7jZVNUozlxOBamDylStEOPbjN9HHyyk5T+XdRIeV0k0U5SYbqmLJ
iyknHH0cNqa/zvoju1Ul6PfAqUEywPRyR5GCGTmSC/spuWqokgKG1DXPV8IiLTzk
p/28J0faqjcXkFhTWHcy98iJaYfP93Ozsmxx7iC2Xcx5z0ViujrnP1eW5xgrBl6g
Td6g1wDlNnQmN12sSuaAwm3cfhdfr/C0MQbAb4AzxZQUnpfAzDTuuoASrIqqxvT1
TdM7WDLiOQp9izdLrPUotN2FPklQHG0UA1K0evguNbtJYEzLVw39NXu0v5veve6/
yo/8Gd33dQZ+qJc4WXnLazoLJ3plue3JQtPPtJA96AQBkj3besD/PLaqAzxlqLB9
Um6VuvSROLuq00egqg/Rhx1h6LjaSceLfRviACsZtQ14OM5H88pbEEajpXPowyUL
blf8XQr4t2u5SZ5ixyYhX3LPDRdxd10q2ZURtkSKp29vIGEQHgCdmgZJZjm3JLnP
XiQ2DDwPbcjz3O01JzV7tcMMX+v/1AVJE59WwWDmt31oCe51RZ7h7/F/vfiJfksX
jvfvt8Pzz77QRdip0/tzxBCC01rDgXR55O2yEhLfWlIgTb/jND1twoNKAdAoWkm2
KGSxiv3eeiu7fLCyLA+mkb49Aw/6ni2MXOTDmpzQghoWe2adat1A8xuBIQvMGWtH
W4pDGS+uz373Wy/uClhm0xsDZn3vY1b1Q+DpTYHEXc1pQAY6k6xj7aUTO5uG8ps8
Xgu0qfzK+6hHBlc8I7uIVofHBbzYaq+xXzjP6+WZwDnneFDtGgetXXxDdbLF4bPp
NlpqEQcSG61HQ1/kpw4bWg+PeqHZGjVDDEGuOVoUFu8mFsgQEw7wwJbUatbRm3Q7
lb4DygwK0gMA94yFeyHGP0KoGSq/aJY/YCDSueg+a5Yu00jZOU9ITtObBelvbAXt
9XMGRLKKtO6WJse/ba68ZAhej8IFQBXtV62cuufAyU2vUxqbtdL6K7erjM32q7o3
Aj8efSN7vY0QLzC71aoJ8oPXPOblH3q4Uspl28cqwIKTvJh0E0sakG67sICXN+br
JjtGpF5OJhjlHN5hq/b/Ix0DfodquhKZtpP0zXnymdwAUG8xp64BjoO2VIEfjo1M
uk+d22IdYqpeiB3RWX50Mm4GfN5rrBCB/NgcmcuDtJ4ET6X1tpq131/wqAIDYH5I
S6dm/noa6PcSVrhqQimbh8YXzXnZ+Gs+8PSvEB2BwdwMoGkiqz9ipTjZDMpxV5uB
/ovHECOU61IQ6YyuXJfKP+4TXPNpDs1unb8iRXPEPNbisTjFmjQ13DaUeerrKdeR
07yntjzyAVUuUYBBa0gKhkDaleAWSi8IjDPPxuUYjtP34uFUf0yi2qmTR0svN/hu
pFYCFBDsZn/Ao5KVMM8HfadtGjzmpx11NmgyNF4Bpl/BLEuF/B1KEFnp6BQeMMnO
O+G7+2Jlk5eGSHrUFCL0sWlSC3u4u+DjJVwUxX1dTn/omQhOQ0Zqtgpe/3FPrMki
nL2PjlLK9pxVmm8gR0UxeOqj26R5pFTxCJGGMrBRi71qaYhdy1Ea1VRJVDk3MT5R
mCEB0GBJJeT7wlce4ZHPWfnHRDaou9Bwv/nUmFQ9Y/9c5mBptmxNmNCa5IwGhOMH
QK3Kz0ibYK6vVxoyiFyt7eFvHv3ugUe+xMW+PRZSoVbRMzD4Jw+I33zxZKiTQhml
gQcclfa8gCEVb5c9YUs2TkRz8C+3f3LfZJf1o905vxMzrBCUd0L2+JIkDh+shVpd
1lUaP97SrpUWuYiqY3Lf9WICFUrFsbzWQnQw6HGTNhEbBw9HsBJPghg7hToIRIjf
JwlC7IW6L12ENa+BNTHEq/l41mPKci0ABBk5ca/V+XCAdD1Q8GWHaWtpKVEr/APR
GL1kfewyNDAC9RZTtJrJDh4OfLLFYZ2P3BRsOpETNk3QIRbrHcpEqdvcZblsNRpV
yykNP/ApClvoOUn1zA5PsSKJPQggFoTgxeJmhY4pWsX69FwGLC3WS815MMlAGOch
0tZPewyuw5+NaoJYE5fc7sI98IxKQkAosq7cTg2MI2lCz94sd7gyhOMAVL/VaWiR
CfpClcr8sd0cd2X64feKEjdBuZw6nh4QoSq7m33w21QQH83QdTZ/roJOGRB7Pggz
+z7FYXhSzctDT2eT9svloHF7OPw13i+8FWtctUuXjcPvuQtg1hrMFqfRNQLreI/O
erfpUG80OtOg1gN7IB+LJXmSp1/f/HTUroBPiaPtCxjGDPX8NJT9epI4lpShnxUg
bzPtMeikoX4qcGwcs57sv+H9sO8aq0tZ2iV4ZNTotVFLKQ+uYRaPMMPi6c/kZ0Zb
x3NwNdxCEKd/eLelqLI/DgxgY+QxbTOQ0jYHcMb7vI6+Fl+GWuGWA7dfJaZn1OiP
uEGWw/1uBeHO7fs4iMo2PHzxP1xv/uMAOt7ulfLS/L8pq39ZhX7zipUHL5VxD+PS
aoXBkjevNyVkqw4rT0FgUoY+014qhgwqWQfi3yojwVqd+EhdrLeFnMrSnZ6rcj+V
7b+oiwj5hyCuRfRtpY+37wqhKDRC54ml/nR6JTffraMr+Gw8t5gqNdGSWu4+pfh5
LZFRoNwkELnvwgT6K0OEg82QvX69VTE5O7QOhTDZJXXSBFVqmouh9CUtQ3INyZ5h
pidbn9iL+8+1pj74dMTQ1++qKkDB9/oR7R2XeuNF0aoRy++xrWr4lFp11e7yy9Rn
3E2ZdBhjbH0aL66kEL4jt9uFPfviOpokKI77gN+0r9FlY7fmTWXqrIDZff0fiOE5
pdsz0JC6BQYPUAsV16KJWuLqCHGfD+5KxBgn7izEq9LAA3pa4U0nefG4xbcfCNS+
boeuJaMoqVrLH7twvaD94U+67Mxus4ZtWFP61Wg3UQYqMZ1cAr3UCI1sTzGCjCUN
L04qICKrik9NE85o6bJ6ChfrHvV6bSZAsiugwHoKktF76xkRVU52itZvEjALTbkU
ETcS7eyywp/dBIuKcLf5UaJgKYSiFApbYqhLb7JXdJEae3Li4xuRsucZq6ZeL2wE
/aCtb/5jWrIHEfhYZpjqkZFhW1+7XPixpKiSAFjlwdNCLNEGgkscuwR/YaaJsRYE
TQTZpga9zCeQWEGpKLnPowfYVVCcdZCqdMqd6C3Zf4HzWYUMdHVh8Asyn9Z/aTxm
GJ1b3dPZWJJozegs4ixDotnxcViwQIxiOV9oJ+KZqDv82ewY3pq1MJFmuXAJYa/p
RZPnSItmDmSVAjCzwklMYLnub2+XZijKrImli2z6vT6I1gekLT85fgpSFTPxsGuI
3uI+JI4Cmmr4T5Kbt/xyYOGQ44gHOAO7qsz1daNbyIlSULcJ32PzF0+++eqC2YeK
miUi3I+QgfAM7dUn5NdYzZMiDkBUozRRlAphzILAPa6AiFKVkdtjb4AsF/rtK/Do
/7Fpow2xjnKZ+VHfC3vS+M6NQODio+7gUYWIu5CRQa2YgrA90VLCiP5PZczPh0/n
bg88rcNofi65RQgBOj4eK8WB6iAt3+bB0ofGl33tK0pQpWbFMrUie/80z+m2TWaM
0vBnITiUwxFdNNmX0qif/0J9BYUxsyMc4DnerOxDmOZAtPIjU2iPCuA8basW0GPN
UIJYX1r+1vlq8rKiJ4p5n6ruroCwnZO8vPBY+SJX2JcYZa0mr6rYoExWMEWbK3hd
nors1IqUlImGkTeUTfN8OugITLRWyJyT9yCZzyZK5yiTwNdRdicarbciJkkS0YVY
/Xu0qLqnLAK5467/buQPAdvrdu3sUeLuyq5dRq6NMWidFt/DKxErROmntk8LvNFM
ZSOCbuB1+o44A3yTraprERwdiVKGD3Qb1n16oUgGvCHS77YAV1A1NDuSoSfVcx2E
1OHhe1BCp8kRVHfeK/nf6Zd3xGybUM7+CiG402jOlsoP4jiCIX6EXWUai2uy/UMu
JzbjsnxwEgtj6kOGmnz/89FayPxiN/TmaBT3yB8rs4JTV5DjbHvgezj8vXKcoiGo
0nh0ZVA7w4U0SzBo6xkKASpBsp+1jofCQZszPkqiGnU9+6NJS1y+mVTZohr+QXzm
4uy0nhovPIJGG81hXZwoiPZ7yG8Bmj8gSBqLNzytajdN7MZxWhkZakhrZCJWjJbR
Os0KzFsJaWAou3L9XmC50BGd+59kJsAQJsTWfa6jSYCNmvtnZCfWllgjcAerkRWD
8YjSnlKU4Ph7R/M7AwSgrC66yC+BdubycskNDOEHWLoOSHtORaC5NugkCEODwM0V
lgSL5fx9yUAKHwausHuhMVTE30EAsM4SQwzWGuHPtZ8pQ05yWUhBKt9ycRuEd4WX
vTwGmDK0doTTW7PsBkt42rBGs70iipZPKMb6igd0cjDwqB6m0iq571GzaIuH8eQF
dwjNiR5HTH3CYahwGnGitXAh90wK93q9QUjD5IBD14NbBcn1rkm9t6ZMma0DMiRR
33DPegk1ICudnJtRcr/vLV/9vNBkKepTgSPBFmP9IgBkth0dnrrxzAsqWJL3zSas
dfnD5CIPXyPZbnIRvWzQs7tzNHc9QCtTmYhLNNFslEKrzB1Lh/OsyVlrUvKCJPEd
FlK3jgZqItZHreXg0UrwdaHuMNravtd3fzEer9ItN9O5JsZJXhDQtrYKa1vCRv9+
UYl7NueTi0x0W/LoopOQBamZP2Mk97Zx/CgbqKKvJIko36ULPhBi/vdCj0Fo0fEh
4drnNjxcIvj/3fdXkQXyMvYrgoxvia52ZACGfGAzedF3YOxd8xHUT6jtfnm4z4al
qe4SwPIIMj7GsXg77unoC5zYm/jR/cWlQaICouLTgl9Jw8Qx6SEm6hm3ZtZwvbZq
iiZrL1bjKxgkbqeB1Sz/9aEuiHONzwJIeAGR6EydhxZ1GVuhyZIF2mdpEEXkBNhn
Z/bfSXF9Vssp7bnMvKlLolG5VDABcdkfOEulrhShZkMSJVRHEf/e7uOeZRtkGVDn
VS43SJm/G2HfJcOS1jwz0YCjz10hrt53++O7P7qsas4xf/Aef8M6COZ9CaG/B09+
Moct4cQ32Fv80QuJIX4rG/nJ1UKaG0twxsx+DMaFABCGNdOUNJnXE4MTYMN+c/d6
YZrPowWBkpouDb5B8gtT7G7pSCDytIrC9Ju9a16iNKZFhigenMmIiJpUls8Sbu1b
IsJlHMvKgLzILzeVsNBH0/lJXWLt/mLBxjV/vREOSWSWl9t/Sg4MgTd2byznAcST
sA60ebNaoQaDLAVNRpK9SwWflrxH1JLCEmpB8OdZLgS2UgK3XXjtA1njQfAXDyBt
AsKJsnxrzkB0A8UCxmNDM1Oo4s4IxJSGo9nsBV0eIn0nt+HMok8BL+vkK27X5fmn
jHvUIY0kr1MEcOmCF35gTZ0ikzlviD6TCC0zLVo79yz68QUZiz/kxVF3wWwZfJ6i
6Tah0S0r10CRV3uEjA6492OwLwbnWQowWj2yaQFAPv2oIhU2MVe++qzGzFp1bP63
n4TJH5LOErXIsSSR07W+szYIXfG+/DN1H0R2SBlLKWXPZCH+8vegvCSFDsk0yrfU
Zm0GwpL5cnKy1gsSdz8jwcG3oA331Y5OjqhaTV+KhHYo/zpbWzUY2VSOFTC4jBut
o6/N7r+Oxx9ttfiu9BF5pzJZIcugHee0bf2jfOfqlYEJVWmYhe4EeMJ7uPHNmNdy
CcLNA0t/IN7xQRC2rUJnerB4cMZ+h/cSSq5PvTE4uDDNS037J7GGIZhu2pmYYqt7
VvUwPqLhUYVrUB9zCGXPNrebiUOAPf9JEf4vmM+wcBTr2c4x/qzFZTTXwXnaDaHO
tzY7Zz+xEGKB2xzttrCk9+CUyFuiBKiHIHeuYH88ApbwdPMnTIJNHImEAoUIP3cW
DsnteMBUMVKxaBB8R8E2PiRM/CanyAd0cped8pzbKfQPn//ehPTOLu+Jkcxcfh2s
NNDo5mP3KZOhmiB9ZTh4fkKeBi1nEYu1xj6E8bCYfAbHhSsX452GKRgpFoC1yb1F
f2HNyMb/yCRdcSvuVz5H+tuNZB434QOxV95uQRSV3JvpvWnLTi+6Iz1p6xg8MvNk
gL3ZRCsinohB6NZpLVVVVeqGKDbGaemM72RT/LOVgPeUYk55ZOerTDH94fAOnIA5
Sx1PbhCeqXPPsldol0l9+tyBEm8wBTlQfeQ0LNPBPezzNw0+5ei80pxDi00Wg++o
rkhy44BAzZomxn2BPtqGlgOj8wVkul8tA8lsliM3hdOhk87shiToAeZliS3Xvw6P
OBFzAaqpnXJ8Zh1VkHcsnfDayBOutiRweQjdMdSKot0zirVLICS82YPNrBAJ1L+b
5EAALAxrPuWFq9todRhPEgRebcQ3JmI7E4I51VK7FCRvsDplyWXtvrUD5Cx0zdtc
j+hR9BQvHydQ/GDzi1SUcXSnyHo28MlHUPr2PUf4bhj0R+wUp3qXEkKBcwQv0qVY
xUlxKYzYVo2CXJRpa3uWbKxbKQSsuRx8QKNsx1KKhlL6+PGtgC+VF7Lak1SLPfNc
oDPp/UxQePBEzcyUNFeYgCJqMb4G3Z6d5t6kGWkK7tVuuw9yYqymvvHbECtOCI5v
m+Wi2wdx4Ju8OFOBW3UIgQ5/VCiI/XuA+ssFdD9b2imQtQwtZdbfS5CkBs/jRlE+
6KAU0KN1fOpZLqPxuUxUW0TvEHVhE4Qrl/CbUDQtiHCBkKxwlFEPDKTWmex9k9wa
0MHsL0BWPl3+X2vp8PpQ9a+wdTaAJ4gKLs99S3jYP0S/1iGKvNMWtt9MaQwMPlsr
3OuHr+7+j9o224pC2YWdHWUm0nokqF2nyWAQwBDgqZkz5KY/fjXI+3GT5UEO0Oob
Y72ytEYOpDIBTc3aJiR608TfDS5zI74rX5JDFyZ3oUBhRDGfP4diwFuYZG/WqFyp
s2tLd8mLEnV4aWECPwnTbFg8VX01iI6Pz5BwuUeGNx47BZ9Z6C1VwIvqPprFFFVw
d2d6Z84uIGgf4qWAMf60yH6uc+i3usM2j7HK8VqKNHvAn2lDCzbY1tpZ8Kcav6od
TST3dj26rZ6k0eM48dwVnc/JsNbBDb9voRZEJ6hPIf1Gu/2VKf25Hr1U2v+ZPBUq
eHzMACQDwci+8ia7ojJYRnkLiS49cwy0s44yWeSeS7BeJhXsJGKmdaPeT2fLml8n
08pYzt+SXWbC+BmM6Bh2qvyH10T5/2/w75xdu6im03jf2W489QpoCE573fVgmkrp
iPkT/w3QaIACFm1gf9bMMNCpmVMxCoasCdC/broiUuUHLeNtmwETDDNnxt1Zj/kT
wULcunQ1Pq7+Wp+Cr8fXYViiMgwIICyoH7HkR3OmZ+cXz5aWZGEOAVpljltO2C2b
gpboWvQrHiGry7sE6E0Ay6gVGfhJRG8Jq6puNNNQgSyZfKd4HxqqNT0osuoEklXD
dpdxYB29JfsSNuslfICVKuR/K7XFIvTZXEVAXpFcjguCx4hERrR68fqtDwt3UV0e
PnzG52YGuCDC9e9ug6SAE1NX3HVZq88o+2jMn77TkXjSt2c00S7ZKmMIfrhJF2bv
jBfMJXPXkzzrH0rOq7hcLmxcbWCu34rtwhtWRjorrxzOsNYNWR0LuiepMHxzXSXV
nUewPjES4UPKID4Byh0E3eaF8zrfJiGKlbg2ROeiyihk8DHwphxDyMbiA9OZKP6a
fsFMnT4P6zFDXv7Y+2WLaODUTiUAyyK0D/3LTc0Iu9R6xHLP7IYRa3nZ1mrGZMJq
xtNGdE6p/3DLkkjuezt/44qSeMVpE1kOs17NV0Th5Q3MM64xYfJZ1e+UjsZEYd/h
2/rvvhzxMxjkoS2JmsvOCb7JHkq5WqmgyjeI/rsgOHnlC8IchcfDPBshVBLTiobm
JsxLtGlEIszplBKcTfVLIiIGbZvy+ZkGsTL9O1Su7D6kuygUUqXGp8/PEtMopE9A
ifAdG56zKmE3SnrRXwZnG9nAhdCLxXSfHH0DeiBjNNc3f1YgxDYSCpl1QFNLteTu
+VKiUL9GXjnN0PFpHW6lVD7tjvv7arHLAMpftE+3rM5m+utnA+ziW6ZkiLQ8LCK0
S5A62icNeIVa+qkuspMzdyOms0Dthnk1x1BSgVHNmozJ6kIMFb4HizyIQ6oD6nHx
yUckzfoBPrYRGEbFkYwJywCOg3OoEfP1wqsAo8rctJ66snNIT8A2Tfh0/sy6CvBV
9G/iA/+u2I45+Jfz2D3yXidPV/EE9uhRx4PwOMERBT4cZTzyLcYuv8TDrNdaMf/C
JrvNZGhumeBIBR1puKokHIrhh/yPkPvTW/wwvcgGlsKPSq4Cv9w4sW7qGxNUQZjt
3AScumTsXncShZMZkmJVxuLEDZajk+bMkqvEqY0yOpazXJVT4nKGkfqu/mwPIzS6
4YZ33hlFppkTjkXXSAeRen5+R49wK3NMU3idVau2HCbAOLRqktKmvuHmvpSg6H/O
YHtPxPEhnyIoYvfVtYD8z4zVWX9H60OlW+GQIMicrk/LZI62Nm3V3CUkb3cMCVGs
1R6oZpOhEGWh0Jx5qEQASaF7+uGZMWcyNNDEhgi/cOM4yef25iCoSWYfV7rIyOPI
vukb+qA2wwF+zUdFXf4s4mVEzBySWvASRoOQm9lK6UioNp6jWK66HjYQqV+PSAu2
7CyS0iUVfvlVlIKtiZpPVahfjFN+sOYZDBJd++Y8h7AN3PoiV4o6lOpy2aSXzxK4
qn2hB5Uq8MEinrsQXXye7MTJn04mDWHRAKQe6M9oNI4bl6f/ZZp29jQkuyjjdAIn
aNKZIpfwf4BOCg8FbA5onhOoSrz0vVJge3PmlUYgh/UUc3TR3ytT8macHduvmPS/
xJe8xuCGySik74Acj0Q1siggWK89fziyCmRB84gOd2+1WxvT8v/RwSiTJ/wVKdXv
xHhZqhNZVOZdc2pTi1+sSu0t4t5dmtERrWQtYyVt/nNalJ3uaaUdVW+LcdmmY3WC
/aKNNeAcjcFBrREOCdcyNGxrgk6WolKTTMP4r74OOgYVxFYWs1MicVnIyCyNaSTS
7jrmcvoXiSExv9m2PzcgBlCmsAL7pzGmRVsQgqqBHj7SibiL3eLP8Xxlb7f9LEgf
ps5lHlveyVFtnSKwPmPuScV8sLzksvkKpTCi0QIuTUOAf13WU/HMRPJjc3tuAKoh
GMaBSmpG0DZFikfAL/gdcVAQ4wRTCcva3rCSjobRHgnLu0t2F8ekr71irePGqa86
vQcIvDTrFei9YynpHQfJTJbQLlcKJS+XOWi0BzGBp3AkWOIi1cIfBxjF3LGFJKro
jBJ8ZCT4cyprYrkWvfkMNJ4YR0WOfzvnM/nYNX74euEAu7jiF6+Dxt6UWiE5lLoT
cg+9vSRYrOJGuidRmjGqrxEjRHg2ku1mrD0DaU1rvna7YVy6n8cR7UtLXmHy5UfH
7U10J8RVO4s12MfMlk/c7mDcqVlArd4+zssVHjtD/l7l3hdLAPj1c5wNRuhE9JwA
/eCpJ8N4hBOuFqjff8JRLOguypbm8IpNbihabMqPZwKbCcki1RYp4ykayYlhtq0f
hfTNqPxsbuE96P+bMtHhuFumsyWb12UuyAhc30aF5byDPI4phM5CuDPNJbzSFoAA
WuCmCmbv/Q8Cy43dumsDkJQjDwwG5lg9ENgA5rE1SE57kIVYoqAZRzW/hXOFqonn
Dyr7kmDlGqw1rP4JN5q+4xQM3r28S8cjlesn0z8lk+WU3GuNpqeGzhnMTQpPO5T0
yyBX2rsaUlXZqFF+ijF4Eam9Y+AgURtrOcAvwsvkHbIySNzzNcXlxZo2K8OVXFmq
baGyeW/5xrwMQSF7m/jHHfKe3Z+Ko4q7ybxDfh+ciVTW5A+kQG587K2TIM4ZqZb9
7gB4JwlW+EztDIGbZzPC3yR507vN25rZjtwRz8DTQqN/rLDaM2dAFHV1+Vq97uEr
W77TTMxKSHOyS0DZxGKHyiQIL0Wt7MjLQUiGcs9i4dNknak2H16z6bKxDqLJUBzn
hU1AYSaUhRgkgoLsnqgdw81ehLecWbmts22D3ddwMQASHQItSZ1KJ0AynOaXHS0x
iJqNOSieZRr9rEknuGKwFR+0M1TIHc2OS7c1/Ut3vfpn5YhVf+TDfGqDoMYtYC2R
z3Z7b0RLswg7FqRQO2ve8TMS7sck6HjTKFRUztN6Kk51DjLFIopuZLuzaETjaYTS
1Y9EA2HHbK4ZcY1Ztzwa5cVyHUCPW5c5da4BT3kk6oVTCZQlOF1tcT4CjFAahFGw
YbHqzN5CxsX2QN0c6RAO1FI/Sy7AUviH6oFChNUkvdraeuVcJwEhYMBxck0DFD1w
EA1OyFiVhz6lH6c2sJEBUYjM2EzVO/0dYlE6vP4xVagEHAtuF2srv29AsKYbi37+
7Yg436ZwtYUZCCVpb4c2qnssnS6/kKqknmAWLM6dkUL6dk0lW+h9yhLimE7Pwz8L
000nG557BHQ3m7LhXB2d+cqsj+hG0wUBAXc4HlSS+n1UXPW3z8yy2oXugd2DOHS7
8MhxsF55FHzqCtDab7uWR366+BqjzQ6MG2VJBMSIoItfNkSFzs0WYk5L+5AxMLJr
10ojYnNqy7qa1vAETnFIus+qvj/neLZMPgad7rwUpDql4rnjgf/ywfo0I2qzjhFq
1bxBIzghs8vMvbM+zYCMOJTfBsw6lHVkDefAGcfW9phEKYSkm8aA9Cjy+rqwA3vh
ESi0wQYV2yzQXufLRLai8MgR0jaPFI2ZqfmHWofTHMLb1m9qtin1hoFQf7vw5VVv
TRundhew37XLFCeKxVzZLL3xIcuVSFj917W2rd44Egts65zb3XgztVNr/XmoPlh+
6q4pwZeEMvbex7NKyFrPpYz/5PKa0bZjE2KKLd+Rv1kqNiUNrg5O1y0Xv4FlRjmY
TTztJmneXMbfQ+cL0Ebe0sNq0ayLRwrkr0uoj/Bxb4Hez1j6yl5rQtbavZHgKurV
HaGAzGNrSkWZX7wuL/8c3L6vaV4ze2oMm0xuxtJ+HAw0EJ/Xx3HJJCt3f0p6q2Zd
AnAliSAMBYTDLIOb5fPPS6PVLtCQUJ85R2kLJMadS5aN3l5lq6daFBkkkISC8ymI
Lo8t8bBXNCqu45u/hSfn2K4mqdQ6H90dtKE+drYG4PGWBKUI4UtWzPZzCBLdat/O
BhN7UlwhBpIx1c/Dt58Ta654bPXaoKxQmxBks8cUF0FlD6rItkB5fu07ODUIMAP/
zna9FWarieh3G8p3MUpDPp6LcycjZvBMKIdtJD+URp+Ol4cjQJZBykBZPSkBMIQP
J2orypkv0Cj2y7LzT+V3jRrL3NEXX4fJxAMA+KzKHYx9j/2qIoZm+qKK9QACjJZM
FLdVrKLOOdA9og+xscYAhh60CmJwk6vUEmTFwnLFxIjwNQmkJPkb53e5NkwoU+jT
WyuTvGVVWtBR4LrYt83JG/pXi32oFFKFuyGt9FD0k17CrAtB6nfGyD+s/Z7JkbYV
qYDat7WJTf5oAvZZR5eAK9rUsoCbMNW7/0qS4pbODU30YbIJZ1RUHE4++97XYOEg
OYa074GWPSVRI3eRx0neFJVLizak4maUr8tFazotmbiSsEf3zmJsVSQ0fwAkm1uR
6RNg92N8TaEkOq1o9ZO18ADqxG7ypV/EUYyY/wAEulcHP9sP095k7JjziF8BgzPR
XavMJFyQbANh86wvH5vGnDb0EBu/14mlRD/5qiDEnLSmVyFXWQVwvW4yA5KI9Em0
LGYEplPyitYZQFbHUkMphWldA7cTWYHhUMVK265WaqlgPCyP56+YwgqVS3TbvAnu
7aH6P76V4z2Ge9LSYKyGhXdOAxM/ndtmJBw5Fodu5jeIvilLDgKMc/PVqgDdqmpy
fDxb/gAcQxBNeafW3HiHL3BMoCl7yWm1rWo5XEtwpxzE81oI0qgbyLNjqsYuHDP7
cdnroTiqTlL6JvophsxY6aYxSZ+suoZFONtTM5CoQYePIsuoprKEKh4dcxG0eyw2
sZdhzrWCAuPs1WqqHtKzN0inIjJU4WEwrc2Li6glNqzlMr3MhvuXtxEjCmYryquU
zd23hxi9PBFmpS0s2dJn2sQjYkDRt6JMMgJjbOx28j0DKa9N39oEzD7GhHl8NjkH
VrU2DbEZ4hu6lEWDApgso77XBGKYo0Q37mvnAzxLmsCI/INP7k2H75FLTn4pDCrU
0FLa994qvZRUNyKHU91R8Vp/Xz49RXP3OGZExBrmY81q/HW1sp0Xkhrm+NhR0JKr
YX/FYbfQIdPn4mto6mYBUMzEn9wolr0FDE0IOR87JtLshK725aVnvEJRVazl1JoH
ff953zix67kxZ2b9dMlZaSLZJswtbhnQz2SmJnOMX/SP4ncKEP64N8xgQoWYLauR
WOQ2a+uVh5k52dWqNhR6qI243c7REVaY191WmgUs9lf+CwxFs+tXfx7HG+5VLofp
V1tO9rEjHDFcydbqLz9W6Mv/r10TLvRgpuQc8EHTxzFmVbbLu28swvDWeTdyJsb2
cR3qefFItu3CBhD5fukHA1WL6bkbInzfy2rE+5hLgtdTRcwv5AJe3I1X949kjSbl
yt8horZ376tpur2ay5o4tMQNA2KxtC0Yju0szqryeXHc+WxS5pcRseMXf5fZVk/h
bh5g+N7TcbDBvTbuOpYIZ8qOh5OWqEoQzJvYOQlBj61Gbz1EVs9/mOpBEV1eix5P
UswYdTH0UIo6JNfh36FtS+eWfw/3Ebi+MnFAttpI69YYrVsDAR5XxOe/wl/tDI6x
z5hmO0nhlIsV9BQNt3yJavfbUL+QxA7r1aOsKqMHCuFJyBVjDHZwzsCOkWkZ1ILq
3Z7NWwFnvo90fO9PyQ1QBX2hU2QGK3pWLQnX1GDjzR1ydIp1s2SeMPkvHzk7/rPc
bBfjOafvvZ2QNmUSm/drbf9f/uzrs6d3NQ2QmVK5z0pyHoot7XBebx0MJgKypDlX
qGcyDjyzoXcx354yJZozo4Fa1GEY0FxDtnuyj2z9FkV5qE8B4buOqiNW/MTGiS71
SeNoXLa7tVSS98wGJqk84sUwEtdLya67vCNntx7oQ1ZWnf2fMhQ3bzg7VAmoCT32
m+GBFlJupJfobCz/yB5N7SZUJGhytom1Jay9gYrh60ZoTCpS+C2AJxpNChCN9ngJ
xwofB2APT9Lb2/VFHXOuxrEsZyolJ9fz66RaDsrbqPTqVONlDKfwuI4r0ejU+TFG
rHraUKdVijOCPgjjzhu2+gx5SvL8r+mvKTLOoIZDHd/BD7kXEhf0S5YJUCwnZyun
+Ty5WqynCmHHrdHO4mNz8KFGpqhs4xW36M1ju5Zmrt1utifPAkcX5bGeFnsn2OEe
x21LfqFsHu3fiOp8emZ0N+fXUegYGdfZMWrTBZ0RURlSfcKxrqIJ79SiivpK6IXK
66dHWA5b0xts07rogMPbATu6lwyt3JqSits8W7JFeu51ZOBZuHFJDQdi6FmeWwNk
rJr+LTrqGnB4DTzh/NHpZPXDRvnlaKG/W77pxfiXLG0eWA3+66xtUbaajpWB+8On
L4tPLzBMK0DJFWjvNV/GyDMifToHNXDnub2pQcxTK/V8HG0Tfw+5IcbfCpBjczDT
FGapUJag5RNPaXkguBJfpfYIj7CIgA6RXCc/EaRRvLpaziLs4DiSBjrIVD6rimW8
nXPk0luGic1zA4OpaUCLy2wQHIQ5p1fv4ZlJzOrMoq/xVUu+yPh8kC+q7/T+Vj1S
UzI86rOtX4R8i41Dvd8sCAsrap7U7j536iaVGPxZTzV8JGs8ml4FjVwF8u1VRAZ0
gtPii6S3kxU5FJ+/qWuhbL3ZyR1ja2N8/ibymUPmM0F7hTxweY3nqxscnPuj3QEy
iwIlp4zdvEysR99D/2qZRj53qyeNdBsxX4OiL6S3vV+AFXRYZX4BzyihhnxTeOaU
S9rgMB0YHuZD0mmqsNnDPJUQgZ4fsVdWkAAbGVqm/LdT8T3HeVGGOQ53NgcPw3QH
2vJYbNapL0g9VKT6EuqQDw9y+AmW2TYOiswKbbqf8AZdGJwyUJOchVgImdd8yaxT
RZ534hlTfRd3ew+IhZoWP4nA5Hz0qJDl37aAvUOcfMCmVPHACqu+QFrufD124hQs
PkfqxIpsGWH8ef7WFLQAXFwLTsu2DR/I+gCB1jApDyP9NL++LrCiO/yPOxo6rJnV
HvUkbuzhHHcMt/fVC7y/B+L3ss/nPdqqPDe0jMzbEy7V2JoPLSMDQYDrqjTmZ6RO
ceBCq0ijBtUUFgUolINkPSVdKF0WNDdMbfF355oi4Gw94xxp62rApqf5f+JlIIls
gXTznp9yAV1veoNiTALjnkpSPoVCpM3WSykQiEl+URYpsKaz02RipLLH6lTF9lH9
nTarfW3vG1LDanNg0JHaw0+xrD3KZOrBJ2W7fTFOwpSwE+uy1yt19sgTHm54tZJY
1Ms5JJo4Xq8El5bnymtD901PwPxZLnqfrvpFweU3QkK29meNwThEQPF9gB0Bszan
Dfsz6vueLoK3DWvy9Vfen1T0aq/OZG2kRTIwIGzPRlMTlwOM8BHwU3exb2B1SXm1
VO/HDwXcgQ4+jSu5SkndnnIzNSH7rPnvqa1A6WZFMkfGozsfwDp1QuJhREB0mxwB
hfWzmuSb1ZXwUs9zYQmuAEI05HgIGt4zQOeXSCkBy++H0NS+DIKgYnqGEHKdY09J
bsaAr8Lc5s9wpEqbd4lyyndZX3zpjm3Z1A3w+KxQnImvOyUMFYQt7dy2KISPIBEj
PGZ4cBaazxvlzb0AQQahuSh9H27oN/ni/XpWZa0RWF1ZHBsreBkcAnlm7gw8pHJr
dr7UZcYIaGkzQnz9PJ6IC5fLdDS2ZnuxYhv2zX6xoO6GE9o6o0ChD6+fPSf6VdZM
Ll5DtdN3d/X/RPdStRjeI/Oc83LU0q22FcUDV5uqhLMMpmPVr4XIoM9RCP5CO3pA
2UsVWMC6ZoFfHLdJcush6gzsDG0+kPnBr7rMOkz+Ej8W6orMV39O5VffumoHqFIA
k39FpShUdyzu35g4zPZxcuEhfoG5vSAQQy40r8oJ8Kfx1JP7YSeAYXRKYLQjVnBo
geB78ls8GSxZC2x4hQFmJ3l9ZEXTuV0G1MckFWOTZHmIxQpahxtdduOsdtHnySSI
E9qCbDPTQXz7P39rf5sU11LyiBin4SxPTB5krykYC+HN1kaXScYqJNuT+l5JJ3hc
AJV+crQi+VmVwtEOZZVW87c8Is/9Uwow6Wjyh7vmzxJS49HvvyVl/+dBxhSOmEls
S2bAmeJTNIHHzQMfacE8rvrAfVJJBeDBldKuSHWKgUsC8/c7nwj46ev157OAt7VU
BJUX4Y6jw5epVn0Xx+1u+NpCqQwOnjFtXo0pcED/xz1VzEsdWXgdX+PyDdzsxXx0
znzsVjWxXCBXyrqlTX9YC3iDKxLiywxxTCuFeSr07UVAGuGOp1rnKG2NJdpZw+ak
KD8tBQTFgTT/pKt85sLggumLHsdOlPRFLbYqeQEfDOeX1ru900so7UvNRq5ooVWL
SKdRUfn3d6AeTTHO55R5eg6+pCyCFvJsHYsbiGzNlA1HDKd7HlsoOytmSATvYK/p
UlqC7PtxYkVXkqRWD/dgXtsRrFlGrGBY3CogI20DlaBiSHsT+fU4Mv1pLVjuflV8
/ZjW1j4MfpiL2GHy7fMj9bs01kZXDCHJQ0IWQ6m/N0kTCVQOPsLs5aU6ajzQ8zSZ
hlG741gUJFBtUWg9v4/qUjG3EM+RVLAAYTFYkoc/52/EaWV8BBiab8cE1JdChSxa
xvhRyrBRowcLxyafS+8RoAZvqhgUL6bEh0TS6BfybDXU7ThbmOw2oWR99rd5JaWJ
kc4/c2FpCZSbdPNNcSIX4SPYckJSY1D7Bz82hphRxsblPG/TolHnBBWa6NzmVSv2
OyaFYRMcTMsYhNysLyLZjZZy/d6t4lw2m9HcJhkik2k80f5ReYuFFmkf8HbPKjAb
iWOYBBov53s8xlQb48he9zgLM9wckUvKC7fM6dDSAB6xogXbw6CL4xEcYuhtaiy2
BCogxs7c7+nOckcwOjZosq/xwQI9ua09tLQwfsc335h0kR+nZdv4b2dugQpQFY18
N62+/IRrvnXpVDnVtBgG+oFOxhvV6DpNhuWrU5c+fWoBZqbqRwLjR5iiXWHt4nNm
4KSVDH8T1gx98TEfgeJA+WUC8eR2Xb++OfT3+kZg8P1s2EFx7EJnaLztL4lXVqGY
9LQQKqMMPLoU+lnJ8Dt+Pq8LpxUurRsNPceQak685szTRH7Gbn4ZQkVB7QxIRrsK
CDK3EnClGjeP1MythxgoElYCrfpLz7VrW5sFp7WEnQd98KOyE28/HgL8wHtA6tTR
i3lxpJ7LiOjAQSFpADgZAUxQg9IGfIVF+40QQlKvz8T2jyCv4BWCiIBSLLTGowel
cpxL/dh3cQzgH7cJmVxjkHPfB2SPV0+FWnVY+S2nOBe25dDcFvyLRH58Iz7TOF4Y
4pSvNontUge16eD9FADeAIrOC/8r/dgd7mQgeyOpt7av3OqUAuXhfA6PIx88Omrq
2hezOfT78WWgRT8fzBqnoNNThh+rc6hA6p/BKg8UfWHbIIPmgBqTumYDCT9PzdSb
e2rB6To13SWB3veKEiy0dYgZdSlHhy1NmKHaZAoV6i3YITT8od6Ge9m+1nBdZXvy
TS4CP2hJ6TW7633zt+X1EdPgAru1yfUf73UMAOhiZtOfwSnbjC2He9W8zR3yHGav
Ms5dPZRGn0yh+wJ8B45G4bySQnaDmo3DXSkqP0qWemZoezLK6wnaL5q8ZaXqoRrt
JJBkfwSJfpW1O8RvE8bI/hI0vv5jIKNvVaRv6qg8PRaJu1hpS60ZpD6SuDqvgn/c
SeRuOeQFIYobSeQMjK3tl6AVLnBnCJCrsPa7+4YB30wTC0JjyAPkermEKWPY4X6y
7EMveyiw1XdAZehL73gYSenybw0W1HgPEWAd9+7XZ3A5aCA2ETX3qz8mxsu9WTm6
FT/X7FDpZ45EonUT9RH9lL5sKDLyd03Hil9JI16yWxqbXhIKhW0ReaLyi9kBKjtL
gu3ySA2BEz54B7PXqUpj9cxWxW1X/DymkqcTR/Ja6fTi/jEtAfxWZYazg7U98koc
URfH718/+spmdyX7YatKqYIo2Apt3Xovlu3t8ZKBoB/XYo7ywWL4R0hlCT/T7SDJ
w/THww928f+eZ0qteTQyKSNVIhlN0LGTVluAb/DcBu4FrYfEkBl4nf1Kmskw7d7P
WbRkHXSk5sSQ9XpWjBEixrS1WXcRkBRcTmu/zv8ADuI0PDMHOLEN17kK7yY3Ex51
zlgsfpdNQ+CiJjgdfgnh83uf2O0KBdjOyHVTLbaj/S9aLaZt/Dr+V+sMyhf0W7p2
00+8JmtU50o0OTSU6AuHDEEmRtcTZzBtE70HkT9P1LpC225qvR+fY2zcND1m5nOB
cvZ7PyHBG2AZeABZesk4sDyiiuw/STDaQeAatpsaKkBw2dHpLPkfO5AKo2MI9yII
ALEH0mITI+rwTl8d77QCUGLIP2QchqBqBCNAq3NJmGfrr8rFZcwh8CabKMeRJo3o
Jcol4YF7/0FwUKayZSsIqmM1ABBfMFSJv5d9KKnBleNiBPkGzP6S1xuq/ouiwYZx
P8JeLNxL6rj7+DcQH1wMrICM9i7kCR6uxbID98E1g2dsuJjOXW/K6AJ2TDuoJKmq
sZCp2T0MPGivvcOfseYgCD/laZurnCZ2SmSNYRkHzWpcu7h9B94WstP3gTUpR+Af
M4OZeiZ2ePmUx6Yf/1eRI82BMMbJeaSwlgPAVXQ9dNVuMksVDocAIZLbZLEvLbOt
S5Up181HbHSEODcWIFxo7Ur62c8Moy3Gt2/y01WgjF0mcUzUgeuP5piXwLnGmUsH
32jHiu59WYdR7Q/h0ti5MOzI9dRHIRo1CZp+CMOw5fml9h3jnBHwICot9ORIYhD8
CNvGLhKBRSi3Nvs2CE5GYZ8x59SYkb3IHmeRQnF6OYS5le1Vlp4oabE72z3BaNKP
HWQqoJG34ouiLf9Vos0fEPo4q+XVGnHVL+qbGCeFDkU7jmOmOH0Upn6Wi61Svbmt
E+X6ShmnKLPH975TtVJq+pRoyn8g/hUbyMm9Sl+PtVLOu1Bs3IxV7eO1pAkWtnrZ
VbGVHBOZ6Rj4jLMcxW5N5jl8bPzizFWYSoSrhHvKIcxKusM7HDP1/twIAvCe9Dfh
x1s3yNckZV46CGka07QugFaSTm7jVKspZJYiiGPhH7uIN4IKQN/YgNgj3QqmJwmo
aN89Dn6TL8uGoAu1O8MbTDP5pZdc6PHP2EO+QZW7gdSubrgURp54Qr2C5PiAQTGy
ZtUW79Y6IRUWa8MjK4WOAu4ZWRuu/t+fd0GKgDGGZ1Kn6rMY3kIXcKe1h1f9Nqv0
QLwzh4eWW3BobBpGzfyUdemNDSNDq21FG0LnIUU671IH/XCoPHiNhiXXuQHDpH5o
ho54+GdBbPcZSt+wh5RwovKKfRFeSMI610rK884jbT+Z68rVl0nnhLGDFDbMITfb
jxgCc7/4IfjwpPXJT7cfJvj/Jovn9uY3smBPlcWF0G/astg120Ne0pRRMp/xEKI6
0KHBW6W3h04scmmY6FutYgO6Z8/rLMbEzD3K7u+sQBelKrhiDVaKdoY+XZUCnD/C
WqYgD+rdAg8J9yHL6EDjokc5JLxXTjD2+4+u4w5cKQulRbQp6B0nhgegDruXJaiC
knYDfgzbKWqoxW0M0nv2g1TILT+ByF2EP1lxU5OzNcUZmulHhdjvUPjKnmJKPdFa
gA0+NdHjLABKXbbNSqDvec2sm2P9E6506jl7CKBY24iGh5ky4Bc/K+R6eN61ag/Z
SJOdi3Y3Xmfu3ReROgIUNFhUAB+Zc6Oe1ixMk46ce+T6F0eRlQCvBG5Yx6YMOVR3
DW6FUgPPZaiZNMbRv6A9uWeIvf32HD/uf81hbXORzLrwQbkPL7iA0HEjyTp43MR9
O1gA1RphNqQz5SmBPxoT67h8365SK4488KsL1nGxFiNGQ0faGUqP43szMwMUR0kX
QzrCfCKwYNCioRNHzWYbUxMBf2QlHo3ZpVR8tjDlYjNus/72kurn+O21rQPK0L3s
O+BX9kLyswunhKnX/Lelz3NrkQkFEeqIG2palfN0LspnCU39glHesNOkYfeLO16D
EPiOGwAKlIAHfMeUFCO5pfcn4yHhIGwRYnwxw3D8LHkvUOZEylTC6J9f6VhhmAz0
gSI2dkm2cSr+Zyy2jcTjTkMPmO8TtRIApfV3g/lk/s+H7vtbfMAb4v+zN4I/wP2Q
bzlUlqMan3DWWv+IDLcuhnaV/6XqjD9KCxJuaIJ2sKv2iI2PXtvpvfd4DZhkEoNL
IHWsHQS2a9QC1tVjnR+KpojSLmtAyYyC7jjQ6oWMMIR7jqSdh+ex6Eaex1R40X/K
n2uCYQf5cFvsdknIUdogC0V5LMtjW22xCkY7aryLB6LWklW0lWEzlEKm4ejmRlqn
skYvBb63LAR9WulsrJcFQal2P+a5Sht1yxk0OdkyQVLg3Hm7StVMBVYjHgCBGTBF
sjZCZTNFb4SQ+TL/Sj5Tz9PWtPkF9c+5gMUh8lmiCjuTjdXI2RKApI0aN+oqBOEr
x1Qj2Lw9xHBTzjpBM/43DpoayZm8VKKs0WaRsmkiZw5LyYkY/VE23CpH7KUt6FPT
kzOKdQgW0mxh3ThsKeSFzjkrrG32a6KoVp0MA3/8KaUElC4ZyuIQm5OiDPtxkFNG
L9vSg4i3cTurWYoOKXju5E4N/u159NSXz5DOmzFGZZBAMJsFMUzej0Z5gy1T2x4r
rPg70EgTxWAKGjNi22dwCcIbHnuExxZwY75dG8nkBpFOM0/CwGembWteqOjq3+rS
vFmMhJwZkVhVIe3uxpcX4QEgVB/GWhnpR4yXbzUGSKZv1mDQfjm+NP5CzhjlzWAh
FzNTjNyP5LnhiuMZCTAP+P0VFGIj/Fl+9ofemCnB5GWLpu6nnhfdYo36ddRMpm2B
072dbW93fCdjCR14sG1zvSaLiit4fE3CZjzRG7L5vJ3v1erEyKRD3RWcALpUWhmS
J41FAnyVdrqvb6oL1A6QplnSrea7br7Xb0g08NOrNjOHpoJqeYxyg7DlFJBN4lxZ
wDwG7+w58gOIrJVlABOYN3dTOjmA6mNVIwX/V+4rVgoSpEO58Lp6cvZP4rceA0kG
1MXG2eEhosEGRxsLvepO8DU9N8lVwV7nEQHqU+2qVThH64KqeusG71sACoshzgUq
fIFqM9DhGS8IvkoTU4lLt/tEbv0lsgGzuqeqRJtdew4XjWQ04C4JcQyP2gyO+8cr
kqHa4+rhbHz/WFu3NM6fpyQq3+KRimZhVWn81J74kcMEoYoXLXVkcP3E3T7KoPKw
53PTA2T/2FTGoRwAtHDs++MeaiC/U6fcfWHjPJT6W/SB5zKu6WvsIZZUsFIRwjx5
KcAhEO7UqBZkMt6LdANddI74Hq7SP69vHCxfp5sxiEleGnPiO3xli/1iYUOUh2+h
R/NeprDBH/6rpa0ZCtfuT59jD7E/rJTNCeK2Zco9lFjZfn1TXBV+k0tVnEZDPqvL
ac4AciosGTzN/oMixnZ+wZBBl0B9qi56K8i+ei+q91Tj68cjX/rH3MJEhIj+T8Ws
hxRI7ewGQaLT2UUtNukHdWA8dhqzWX/XSapAKT5+qREhsY+Ut0s2h1EpH3obpvLV
/+37irFyZr9gpxAmDeBbMWJiRMw98asBbP3vR5fCI9i01XmsRU9NepZ8XSMuSdC8
GMWKeMoH8QZMbSduTRBeZFj1Em+7JXjy2tOi/OYBKHVs7sknRNLVA3rujtvO6U2s
h3QBjFJu7RT4gS8LdfHEaDhoL954Yc4WwBus5WJQ9d1zChHJn2Gv5caZhySc176r
Y6a5c67NLlX2zXuewyA7Jy06IbzwPLTK1BZw90Tt0XIzXIoDSua9hsHDb8aWKkMQ
0is1OExvMluCUREpZzKs/ao5hwrq/QdWtzeT41AovaeyTXyo4Djv0hzKjeFSgLW6
Fy0Orx3ZMZkqBOjx2Swl8eFyhfW/x3OS8n0MaEKGdYJ0tKn8mek58WQXKUjiXSvS
0ZZvOxhBl7mPGqifYD6lVQlJ3rUN2oFjlqaoMyCExxhD0AuTR3pOXDsh3XmVdBrF
PhXjzMzXbLa1c+YePKctPfWO69/5NrxnVgHXujgsTAlcvep1R5Su/WLZ6oqTJQZW
HUcmVZ90ChEOzoeWyP6CEKe0S1Lodyo7tgzG9TjQ/oKY5RYpoDvfObkXJMQlU5J/
d+9eNRkZpeu8kQCFxxEqhsrb254FWpG7FXdUlkf45+ZA3AIfUdsrCVlH8uvCAhhV
WCtvhDpcZ8k0JbACmDd4GsgbI2DDDjT4NMRw23rym4Q2MWLFOaFJnkmmGrbsKb0I
JqTD6hC4WnYz2XJghX2W0WD6sDWBXlNzf1Wjf41Ll8IJI29SJKr51kUEQ61wpDm9
9QnLeoPXRYMZ3KQZRlVva3hJl6r9PSYbH9jPH9hJSIDZYuXYGtks8hKDtmma9s5j
fXei7h5MyZIfhQLmgp74DQ3wCfDEr+SKicOx2GkBoXQsdIzkEJji48ALRh7mNlLX
RJzwX1VSeIk8CjDH3jXLgJthTaYNEMK7uW/rnNH0rpc8MpnJvmXP81SvoPNTAClt
9n634W3wx6HanXYjEza72wBW3RpWrYX7k7Q0hBTuLZsAx3cdFXXkc7OLNYfPv9iZ
5JJfvIzfLu8wJbCRielvc6wPEfSIwgD9ORUomWCiP+ZV89OcdvmpdVGca50yCk+R
IE1tn1hQUn5EaMSH8G4DSMZj863hroeOFOXMAGq5v257XuxHDtgVctKUR8ibaxTL
q6c6TomZkdIBM/DVwIpcPDPAvbBSn2DokBDQO9Y48ww3xIx4PcRn8KufBGnoYpnu
WxUBL+4Lw88vdoI37x3G/1yzNF67UWDtT/mR4FygKPReOVoLgqdMK8S2Ukd4C8a8
lg5pbvOXeJ+ZQgHy1VgunrAQ4XotKKEOa/zvWTRqPbqx41omIj8YtAJ7FpVeH+J1
mBTb8sZxdcPlabiDSBJnEYZgsmD+3wK9MJdVlj/lGwq/DQS4+/TNTJQ4nvrHb38o
AY/itTpRj+5QNKawVJqHTGWNq1TcVPyf892ji9F+WBWowH9gEEOhYC8Fo+UApZln
Wv93zkVhZP94nAkU/VnmOnuHRffluVU6OPkkfORc4Svz5LLqLwYaQvyWxR7QM6Dl
/wnUp4A8CgF49XmyTnLQeBoIGYEo/An4OfZ5Dh0iHCJIHCCMCOaxmOMmnU520L2L
sc/YHhyPruH/zWzCdGMK7WR/Y+4EBoA2nVel3tAIhwPqWUTI+ORj12bVmgY/nCuG
pck3LfgSv1toFpDX4E77zvWg1k/foCz5J68RTVv+8M7jwFVnSZAss5sh23WP44GQ
T4IAugZbQ5bsq7OQJ/0//vfsQDlGjnkD4w2qggvsSbfySK65qjixmNxIK4EagKKv
YL5PHh00cXNftRsPLfaMbaBuz+C9B6Jg3xvFkh1GeWsBSofQDr5getUaOzDyrPG3
e12deKykjwhgTG3TTLdpWchH0f/UH4nZd+kjNat+a2O+RZVS/1/b6mYwybleKs0m
ZjZ7s4k5eqVVixd02LqzE9NTlorHTLHeWvQIw7INSbWP1csA6jp+EpioaGNLfELQ
1vtLdpM82kaWn3XJ1PBp1LGsvrdX0BW2rQQjIXVkcqw3VpFSyve6CdJnyGiRmhf4
aa5ADQ7C2lMzqMkuZgjYYnhNO8dgFl2hjC5X5rKZb5Sr8Dn41wjPXkhiyQroXkOr
ZPUXWJHgxR19r5nnPb4Wa0mj9J7E/sCa5w2qhv2Eud7x1tZxsw+yopW4H91kDVrF
zrIN0Ido8tVqlPP/QbyUEEeZdbHTbyVnRsG37BrMGY12WIN7Xah3xxMNfZNhRvUj
NZQqxRjUZCAz+t0eDxlrkw7YSn9Xxt6CBpjsW8GOiKM6/OxKINyQhjmw4SthTAdr
F4pgJo6b91SYPGUg1DDxlYcB9Y/nkQC31Lm7LltExih0oPfKvVJvWRPu5UBCetj+
90vLgf6Ce86GUnm/I/qXZdtGaAfBgQhw87wfEOdQmbTvqa9XpBwe2kqvF2Tspipg
N6T0+hkEp1nopCfd3g04NX6QE2utwacAYksb81/FOMPVGu1QYzzDnf9ps2DOX93Y
b/ue7zwMnmW86b/lebqrK+wNozSxYP4AzbX7RFyob/AmnYv+MTDXrOtUPbsZhhTp
2Es4lANhq/KBbjFoMyvIzmbvL+Swwb/nmF2b0F6TZ2N7iO6iqHW/D5q9IrInS939
60sz1Ymu2Xh5TfsXDZQZ30vqDVlDjWkJ/IwHOGA0cOyYlqfU0VXqLH/UsqeZ/wOO
0vE0iBmIsI9z6x9CkwHdOZ1YXIBGqckQtkv1O0zpg86ur7ti7fnzDNDS+uNgQoSw
Gzodn2EThjlFhSQorscDl9izoDkii7H0lk/oevTRuhphnsHUVNaD7dxYu3TtqXvp
SmoYwhX4Qq/EAyKjxfDpOMJJG0TFqj/hywV2PCaRm7o0ZWz/b6AQcMfIdqay3gHT
UuIIQhtKcG61PwrQQBrQH5Ox0tzWLLOLwcwo2u0I+4JWKQqYUy6QEq/U61mrhEW4
geh73VvfRb2swL/vr/sessVNviP/IeQT3SKG4Z/S35D70f4ODu1x1dSfeP+BUR/F
4tKQetWDxugnGNQ4BNW8i1Jj6D0Flxr6NLcdb5N4iITC2jlsc9NJnhDtp1pEKsen
jAeO5J3nY2nKDVBPGUzsoQ2sVt/4A74plsoUphWhKeOeeCvde4cx+l00McVHEiKK
mz5pn/0RDL6kltqqzV566zLcaEG0l/6JUKQD9e5jXmW9QSbdJSg9Quo46KbQtjf/
K6CFcIl+ynHcBcXred/Mhg8rvuVjlhRADh0tpAic3YyfPXd20lX/5jjeNJcDBGhj
QrKDR46hWHJvxKpuH3ZV9nn5zN2hvmJL45klwP4W1yBaldcuRLI+maAQOqAQwbwX
wqrmg21OpraIJRWx6motGi9VQ7j2UcJQl7YY/+UJ6CBmEdPC81R4jKtSBbGiebwv
/ohsxh33Q/I2bh4VGPGfd+hmpI8u62EVXutqiM0e9ukV1D2jXw/IwFrK2hfwF7Ee
1JAYIg6avtUdFcZACOPIMdsmt8nkwiYTO+H/M8iko6kB0sn6SG3fan+IM/f0R7jn
rCyxRMQQZ1T83Y+rTdaepU9CJhRq7WNQkt0PiHsqffpRKbtndya0IpZc3bWzBEEp
KqQ9z5yqu4iOo+hGOhPGWvf0CEbINdFnbTW5R87VuUSU09ZzsISM4VUh3/CODmI2
ihxYGL5lWed9mFSp2asgy3apzCAQOa8gVKkAShEXJnU9BI3TOXDJ/kjPn3mKoK07
4yrRgWLkngK/YEtXZkATeTEKho7phQ418T0y1y3E30+Mqw/KQBYLTRjJxvyI1tap
82sjfi6HFgDcasqPH+n99syUdp5H5LzV8+wnSFAl5GKY+f7nYAq38GQG9NLCXOpU
40tlTrF4/uOyvLCw2XEiTrItodeJdIiFUNg1SptPa5Y0Oy3sTOqb8miQoh2lQz/5
X+GhOrPnzSAQ14TbbigYGu8BI6na9b5zGHjbg0anhDI4gepC4+O00IrtXNpaabB4
C9XKk5cY5edA8Npnkvayefc5LiXqL+iygROEyDivxMhB7emkiqmti7V/doAg9Iyj
GNAp2W5oummUKI+ysJt/Bu1DAGlNm0Ei22PGI3FUXC0piMOykXLpZ72o2N/dh/kl
1gkxmDglnwM9qXROS0MOucvvSAPNX6g7rHKNco6GMPt0k239RYn/nbJfOJxBD4+P
yDElhh0IS4J21sElS8im07RmE1ig93Cd0KMMf5PJoRVzRWL/N//35c5dwx1rl1Ft
NDp/6a5kde4xxpwIOD4V/wXXrL0b0quwMMN9pMXqEivRNa79hRvOTB+HkP8lV+ge
W4NxNSz+PeAMgCozb29tTezHsrfMl4qNCzfMRfCkxCwQt3OjbxsX+oNqRF5fqktK
hQAtJgBz0TPhmIVxowasoXpF2+AWAqUGp2k7KoTyev3jn4ZxbC4/dY5ClReCzpVm
/qohhR3YqFTqAH62wvI9qQkbJC+EI6flNPl5TEf/MPjxvgDMH7JRfMvMsUOjeUg2
2+q1N0juUgU5syRj9A4XaQljX1/67756nkrJvbiPjGmFQCxEB4k2UBP4WHBpvIUG
7yq9XzKHcU8vknJwCkMy6mHw/RORokpYOl4M/yCLspZR4EaM69asaJ4VZCzAaq34
hacFiidIu1ggl3DJ1bsdNkEcRLlNWCIiGZSANVl+sePW+Tb7rugIK00LpdC5w09r
8EIjNdwTqyplu4VoJD2nGNwzWw0wzW3CxybkJdXde4ohrjIadgrSO8hCrv0TSLsJ
9VBdssBdDcs+JusAky0p9h446ouL1aau/JKiLEEB6m8z3KFxq6Jp/kkzVSoWKWRR
BSZja/wQh7ecyaZdwG4bbzBUxp/UWX8EONdVVmsk+wMFcylXMqr7IZfhVg5zghDJ
dYxRdIsJEAgSCQhiIyj70FwF2BEUxAYzFKuTKyhmEOqquZ6sO1N0FdGtLbSGJM/g
5lnpg4TjMEmKa32lODF9qkNoQJgH6USxlebt2ccMjO4p8LwiR9TaoJM3dxprV8kv
4fO6CBYGUEzvpv0ZLWaDnklAGNqfEuoBMfkwIHXCAKO93yiEGtrcOcvhUvhSCOlP
4pRjXUHj6Z++MB1TaoQJ+IOq7+sdyPxQdo23CR7FulSh0yrLNZkoc97q5Nu0DqfS
hZYdH00Y80iio/ZEWALmi8XcM4Z8L2E7UA5DwORsysyDmjYW91LEHPQKvK9yoSfC
KdZ2XBz7EH+10BSFG6qaBBRz97Kvrs2qZvBYAOzZZC8c44A5lTBqeIpKfBy7UJ/e
RUozUxwyQ7XKMNTZ8a0tYPIsGCmnY+4/xCRjKcX737exe4Ee1La/Ss9ACeFoM5PI
oURxnAARm6v91Zfkx2K8dy6YbSUyeZIHobe8PDe/p6B965vP5Xox+Xf3zXLXp+29
r8MuJ82RC209AZoWo7rdvokon0FGwcPCQVciXnKKrLmX7Djp3oKvvMIRaU82IAVh
Kqgo5DNHWR0f1PuQG1bzQzykLGE/DiCjDdSeqG9+d3KPeb0WrKQD3oBT2jtGKqiS
8kLFfRFQxVO7rp6a3iEeoR5HB2ZNG1k9K8ec+5fHWFSgqoLujzCvTJxkMFdru65j
/7T5DWBOgOtbaG4bVG7YGpHBMKEo0FxkllF7pWV0pdXMWn+GOm+h2kSyl7pJMDOp
h0noBW9EkxvRFK7xuvFBqo9S+dkooErcrxvRTIyS3Im9Z8A6niegq0fmrVlW72b9
o/tbJPiI3c81IRLVU31pz6aDfKAJ9Xe7bdr7VmN92B0aQcXrb2PEoMFRmpPO5YlZ
dVxkYHzYwenIHMXF+Xs/X4j5GpM1StCzUv0H92r601KhmqdAgx4zQMDq4AFsiSfB
OGIyumGMWxPGv8p/jXGvPhoTHIcbQEZUbKKNU1exfAHJWODEuqXtmL+iolTWzGV1
ykuZYYUwbyS2FV7lm2IFNBMpG37ZYVyl0QwAXjCnNYaAWJMGNXF1sMOhQHOKbOeG
Bn0ATyEbz+zMAUwHaXrXiDeJrTsSoC3TJPnO/vbcnXlQdpDjz2r7NHJVhmaYc3zx
TzRwlACnCTfidSLLtEVS/TZ2tDjYmKHQ5/yr9hbQA3low1jUNdamIXyIE4vGfXeA
dM+vxLd7qHa5yume9+XcvxFdfjaDSkPjsmyFeajxP7A4JvABr3bzWndl+EqkoIbl
8Fst3FiA6jaBlYXRX2+ZpJWRWh17QnlsKMJ1xZa5ozc1XF/CPmz5j/ydiH7FmyU5
XhOCO0tlHQjqnKsTIzVm0Te4RToBrlO9as9QTyO9w3vKFAv6h9LqQPoetesd/4Yq
0Sx5vPZOGRQ1yeVWC50OZ3XUv+/swPi75ycqj6EiTSoVMZ+pTm8hX/dE6mb0oVWP
pxfx/GdBCr+WuyQegRYW+wA60/RO5zUurCD62U97q+mnqXH1l7U/NQUqfwcaKt5x
m9C57IzB3GSyFM3DfVKVJEjqIbTGfIEpQho79/aQDOOA5V2y7ayQerd4UAXIP/oY
RpZLft7jm+E0XqmVeALYQ8Z+pyc+PTTsKjFYO64e/DCO3nTFl5O6xIW3vsJKrJHo
FNR277dfYRxBNRa7yauHev/c8BH84kZvT0sKd/m7R4bxPQlnqfzXz2Ox2h74m6t6
YDU6II2vG4H4/xrgdUu7RFTu6X7Cr4k3mfso/7ozmJc1LYr74Gg1QhFUZkamu5Td
mUdXenFWg70TRZtfGaRQcyt3/wMarnc5VuoJqlCbiNkn9F3ePJUGI2yuOhNsJduS
GZqEPa2SmLA+omeqgTOlthJzS4gd9qdPZOVsoZuMfuG2CiFkTGmSj6Oe2dSdgOS3
6uX0/QJFLvmXVG86Q6DyjA5wm4mnTKMP7xTlSwrgFDeYrAyd65IqA8iVEYSOnpE8
3L7ZK+ih8ysXSKP37ogWvH4AZRh39eJ7JcPq2D4BeLZjRqryzlu/d7rSPAg1Ko80
vYCTW/zVq+IX1u7ezpu+d4X3N+yEmUJtAB0LO1636h6ZqRIsSlIg69oCLV7X6753
l4Tfc12zraKL24G+fhkfuEZwBLnE1pnDioK2i+1TC08ADN81MzBEN+oae1tODZqh
bDIfpEdb0qQZpb6k5ChqvnjQHmcGmTwxBXgbN0SXdNBVKtnZIbhYEKWxjLICrVqA
I2ptUDJphpYDB2K2zH8ZA6i4uo21HTy21Twdz2XyuZyBCWZ2ETWgZIFEGr2yxnpx
CzF/0yFhDzUr9CfQmyVmnZAcl36eWTz3NCdFMcPjKgdRxY60ED362vCcpfgiIYzp
Aj4sUD9pGTt0944QILB6ZuYnD7j78tmoie+dmtxsXFaRT4uGuAfVpqvznKVU09z7
6gPDIwvq5QJHfpseD3DHcFGVam9OrCai5kIfo+ZgheYp85eEUjn5NQ3iJASZqghX
CIRnXo3mPUuq2MGUmGWWR7pk7j761bAJ233lglxA+yQqd0jrtx1YiJw4ZkQEzyYj
ak83dhXlKPZBMM5PGgBlnZEJZj5OIMGQdLPbIc6a/1XeVA2HVc7o0xd5gL25zk4z
lYEYlHcZiIxUq3xecoTzwnZoNv2NyGOY0kspG3e6+9kw/Q6dE40IpPjlu+RsYUXG
m0N6DGKVb81NJzKj4U83lYon+P54nWu99KWl0An3qwsskeiwnna1i/1VyGhVSCgy
RBpQuJ62D5IEq3XeowbJPcIC/BHV3Zy5Zm+RnQFKYzb2hapLMpwkXUXNDCkQ5drY
sn2YF5ZdH+3c0khuJtpScQnn8KGeawoGUC+iieVWRj40z8mNp9ys+dEZZ+06u4hf
FGTN3sdZF9aVo99Fa7i/Q0AfgvJZroMn+pI+3sE3cP+UqtylRSUGIWVDr0h5QxVo
um2GSKKl1Jv1nEG5C8ZlGx8/VmqCJ5Q3lCUwPs+HyBPp3FTDAx3UaMZsZFgvcdrC
T0E8NvuTuHiofkElk72I8aHOCy88r/pPhnq5A2XZ2Osjx1EEF2sYeFo1bdURtl7F
/db/6zOrc0VEXUm4MMjCAOKDugOPqsZKksZ2+Kh5u/E50xUKqqE+2le7eRps6rgY
CWa4VfbSVwU0niz5kzTFERr8UXlM78PqsBXzxW5GDAmml5wcH3EDsBy74Ph5LA1U
rhKsW/Dzri6kSuaD+7E3+ImDLoXas41l+4RhwHZTf8bFl1ugmysNseVdCYJAhJdg
Wecd3ddf8Le6z7Ye/5aWCSXH+nYB+Baa3wMa9sl2EujV6NMMGn0PVfMnhCF6VzFB
wP9BTXRjUbFTShGAed6ZPZD7lLNS4yDq/f/wJw/+JlL7XTXARXDHUWc0+rMhmEmf
F5KfL0ArsMQ8fp2i/pVpWS46Hi/f3//e/ikQFkKnSnDzZfuYO+q1Fb728lN8VoEY
KsfpX7maXW4CQzuMXExw735JOq7+IQ2xRUOYBrFRlO8VwsvMdOBlZX4zr/dIc8ZK
XnR2XO3/33Em6HiFnz0d9UkYNXRnnYLiZzkShb4IqkEtdaHx6k6W9l7TYuOfRE4K
XS3HGM6iUlRWR6/li+WMJetGZ9ilaAdtzWL5JURiJck7GZd909ELfxSqQRYPnQcI
nRzSn/8MRkFVo8Vu8RccMo1MXNPnyIMbxrsA/rrz0DFFcgVOZezYJRZ3+0h21K0X
TfpIskDP4N4emLiWbMxW9S2XL9xY0usAjL45lrNSNBsRz8rwvJeJoDqskMAR5URV
IF1hjUxFFnWQrTWf9WnTkGd5N9oqVk9ZTwDdAYk3vcKPEBkvcG0lUxxZ8LxLFQ8L
jViR9D2pFeLROtZkLScpT8YKTAUA/R8I95kO4UMp1UryT1eu6WElFrBvsH4syrU4
O5jaX4gtxE6/Zcuy3dfvPEeyuyaU9eOKfQ/ezuKqtKxRSheoXUkbB+K00nlqy4kt
GToFbdfkZTEXv89ATh1S8xz6qbjBtzP72LrLCewN1/w7EluOkPqn6psXslkYJF8e
UPhoBF8tnQP9YBN+zImOx5RU3Vice8ewxXfeHkTVN/XPqlOWjClz3ViVVKYrhb7x
bCc1dMfXTz+fktM8aA/CRGamkU8KBi1Khwyj5jlaaQ51gq2IJCUBtcVREDLo7b1G
WASrOlEURtbD/NDydBknI6TPK3K7AfHi/lxJr3+y29m4H3bhbeN6IeyXROzo9lay
dgYUKXpqpYbarGuwmcQGcOdmu2z35bTtNAKlCIc+T6if33E3i7wBPxvA7L0rLTi9
7uKbA8hVCfqgp7DfhrD5aobBKMk2qoM8Pk/g+LqE2je+D8QiinKEW/M9mbZwBhoN
ay+XTiaJrMnmkZqZiZDlQRS1dDZEIsHB9heIYdtgNVXvFa84crbu9vpcKa7lsBu4
nvByf41HU6iYdb9MKenE1zBCBTp7wUtb1rvXL8k+k7/m3jJaIonTDddu/YJ3b+an
huIGFvGQTDIlyJk1/a3WFUcrum6saxoG//ZviQXgNHBempoR5/uKPJquvAH3fRg0
f+HNL4IviIcV040qi8o1nDWiS2bZb2o+Cn/z3gR2G/UgkTjtM8bV3AHpOLNcLBJb
QOWJ1d5aLXxkuAzeHYMVE45mJZWYOjIAzHQLkwl58nCvCslbJyCCdi9PhiNibg40
LV+bfJt7+U1cTiBJ9t1ACgCS2efDRg4gCnBdXcR1v9ZYL3hu/8piRqHuKWHRlTno
pQQXsKoHlIPm32WM2Rjje9pLnaBiY01FFvvU527Kw1Pp4AY0ok+q4eIO2W/bOQAQ
PnRNcVfMrpal813CvnU8Il8ZgeLb7nj/BGf0GJixQQfsDRAd4G9aKwTY0fuiMEgw
EWr3ArH2L2zkkeKC9R/OQoEB0P5wTR5f5MZOVUyonDvzLD/cOM63ABXE97Hku//5
Ois6hPLp3bUYDLZjnLFr1UNuNQlZ8ClLpG+c7/y4yw7YMGwo6m1a1ZDeS26FITcL
Zfu+p3LoJsFjU8pqB4U2XTv1TwOpP94f5FaHTNRmMsu0wQ6lSsZJW0EQQVdDl2HM
DJp2kpZzB4mmDtCKi4zkzpsZzQnOJgY2yc+E3D+p85xfdCK7nVl1vv195EQbtKhJ
N/D29/2BsKchZpWp1G9c3vseVjT3io2v3U3ZlNIJbRm8uZxzX2RBs9hlFvex3bTE
l3STPhsCHRsV+4ulWdSW4Cf6a5FPnZzkqtXokpk6X/3961kWLrMZixU0rpc7cREK
hYH6Q2m0Ae4xKLABInXmEJV2lhJ17r12kDEPYNR491dDJUArGY+5HzuLJhwt4r06
kR9ZEG/YxaK/jqcjMucbJS7OIgIle50tZjtYFnnMIwNpl1VadPywPQmY5mkJeP5V
KkxIw2muhJrPecuuN0w8oewjJybZV4ZTjn2Qkq9p2lWkGXC8zfCdMPRepMO6zf8V
7l+TcH95QvFyQvnpQNEKmPFX+AmHnAoQBM4WbCD9K74OannGDcsJaPBKqFMLP93+
D9j0Kon3xtBxfCZH+mWk2C1Ez+XGpI0zc6bykK6m/lmNKZIFooCypP9Lr5F+5d4p
4xTaRGyxqmFijMksI4t5YHCU8q8I9U1fFPBO8pOMvb49cvj7HY4R6OHPrHQ5+sQK
w1VMW293qLMJME+JNjVAG0klvsL60xzsw0bfwNUVovV/X5BNlPiedaeqRCsbe21E
`protect END_PROTECTED
