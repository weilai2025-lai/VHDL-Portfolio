`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVG6h0593SzAZXMcVVnVofDJk4+4ldfp2zQ0kEDq7Lk13pX7ZMGMRRrAUAsOjls3
Xitm3MBm2jHJbk+VPcNBr+nlKAwzSmLoSu+JKeIWTQ9Zj5jeCZ80v4DQemLxc37u
Bv5kkjKlZn+0h6fVoGiag/k2qwnBJ/Dd8aV0hOVEk/cefDsKIaes2zJ8bJK3SrSe
gXDvDczeArv0T2kh6yBKhySSPi5rmDDSoLu+MOWrIgfKGc4abJhnihURJAizxtQe
J3eDN7CLG6unvApKLi01KZgdJObX94OARsryaEf1aTgjvVry1uhfBHKy6l7IlHFH
rZYVR/ulRHGqeR75n+iaXCvN0RZcYyQ+ZQy9MrjknksYvWiulxzp1r3K04ixF4+8
FWmI6eINpz2B84sCnYevdPbpHSzq83yeRNhMpALfNxTcO7yeLKD/2c43IsJM1x5I
KRbDZ376pvDuLDNYpzbvA4MX5uVo5biJQcR9GH+FeH834/rOOsEyiT6WaaEfPlq7
FkFAQQ2bDGzSioMMe78wG1gIDJuAepfdXfh8PxZKt7s7Qy2K5P+ulxOMppP3f+HC
sXSK5bB40tkil1AfhFhhc0hR2NvEiWBCY/sDge8yfY/wTQvzhgDbPy8RFNdu4e0y
gVhf/9tcCWILsWKtTFXv7csb5Y3MwaHh8seJP9MRz8B8/rvkEY0N2zV30FXKgLjD
LwcOxQnpMqQNxrV3MgxRXk5zludK5uL4307iNRUiJkIaA23vZ+MVUhdRAZZsNAgw
p4JLaAOIl03A85Aan/AFl59kZvKOVybfx+wd7JZkr7Z1C3Hv8kTuS9lHYvbH2YA2
uzYWYu8hquof52RfSUNCDjuZ5QMsUF5TBwQ9q8puf/Mg4sYW5SPqNw5+yNIQlHP3
5Tjz8/QzSdgFXPU03uo5smyCD6hryzGINKQdV8YjEgtbCDMHZGcT8TbNqAj/Wn0s
/9vVlG2DvTDbyhpGjyTo8z2VV8f3IIOXADrEXVA3iJFU0jvmFRxq8kkzYFfmWgqh
XxBC+kRsva8n4RwpVQ08W9RJq3MjqWQz1ovbxv7SMQ8pewVPEiyJ3mGtm6KZdCrs
fkuAlx+lZuA/oU2el4ltw/y9DOUQFB00bX36S9cTWit7Mtz4weqd1GU9oMacTgIc
8RMn9qkRR0o6i7CHhCQqYSeZ1HuAaK+clcX5QEGdWDM3uue1RYVKIATXvsbY79Os
PQCZ9bStEOKF1np5+NquTNs5+8PiGFSYzJFP6bRj4ZltFkpw9FgkNZWYmm3+TWmz
euIF30Ny8WbtFyaTEkFvKgDSKmmKuCSwP63IkpJlSEv1QkO7cafyBkq/HvPgztNZ
QK2/dTwoV1pYOqAaTjwZaC9maTbyDqq9kgxk34HyvpA8Gf3boJrZ9VBqtOQUOXoI
TdNvPwRYuEdULOC+Fi/DmVT9dZYD46mAofjFSIMKUruLPmPpvkINAqi6rqVUEl7B
CGOdG7M1gvyCGWao2pQvI32DUYr+3Os0KZBHPURdNpSjmMcf7DEX0TlI18ToiJU/
/H39z/nDw5QxqqqnEBn8TvzWIK+RA4CpN+HXjc8ffMDD6aegkEEbSlaqXaME2TmH
lgLhJ50413Ywdyzs9tJZGZPUgmiVl+IriyI7eHQxUsW0klMnuqxHelDbURzNmD42
NcZr4Ex7bcKzQ2P57P1X7CDI5u2CrymYnReaLppl6K07L81ZQ83+DdKJznJ4I3q5
RUkCBPQMTLqok7GBxwM6UEyhYTLuNYKv+hNr8DQ/WDjCZB/tGIDlr2RK/u+QQQ9+
FAjO06L3lgoRNVxs0dOvRSjF10V/MzVKF0IkQcOyKeiKP0LxPtDi2PhhfPWDSOwj
oi39yl8ZiSsRSQLdHQ28h/A5sb4ExjHvJ+ju1gwFx4dU7SXFZQmkwRl8Ye2zccaB
jGMFn7XHWT/JUlJak2jsx85zq+QO5E8veRtILz0asGy+vTbHlBuwJCoHS1e1pqbE
FLL596r68Zr1VuyvynxGasmdzU5a4rWiL70VWxsZ/YLDWL9AQBzaC10hzF+h5plz
F29KUfxr2qvtC4lGoAnDihrbAbNTdfn42F9cMPtx9J1mSNsDN1TqdLNwX0/pyw2A
7wqKtad3LGh44bSoU1sCPXLc5zdSkInznb3A9fpkH7ZwllsEhjKifPvkjrVEvKAM
sEcjlLaoIgncu0K4lpI4tQt7VMLhpkCg/AM4RShdB1L8IvuXAfy+0n6+RddOdTk4
5fkoYk0UQr1KV1f0U9pg/uotPX5eOuYfSmcn7bHGvA2+UTbrmLa2wPMXPb3N9qWy
B6YGfpCLfnbisagPG5SGPcRScpydtspH+k0QCNH0N0YnO4/04U7B6TqrEykBBXcg
vnrJl5FazQZnKe0+aOQDkNusHJ0oGdf4J7oEoHvrDYQgVacY/2J5WffygGoeGL1A
cm8UAbw32PD4WuSrk0UblrHil+PUF89R84TZU2ciVMjGReP+MrdtFYgrU6tRCO2g
agI4XCbXeu5PQSuY9CKHokFYcCnSWlE0m7fgExNa9DZmEnkKxAz8m2cvmSI3ncxv
Jpc+t5GuEJw/Is0jYCik0TwoDDzdGwRKOBvgFi9V3aQOt44CLNUZ+Feu2TLmm/xj
2NU+rvZ2XKlj0/KEsxM8gb/NkvLYPsHnmdf2nEM5imKrx9//FwPRGPCyq0CK6EBe
VLEAhf/8WFEJPbPw5nTFR2lg6jx35mjp1+Gg69PKgiqr2tVO6FMjExDv/hMEu4N5
QpNq6cIkcxFZBxlTBk63wWHjISOPC1piSJLPxa6Q1sDWz5rmynjepbLELQbvDY9L
NNpjfRbgjk8ao8HKSvhr2xEpugbqL0Jgyf4lHndUrgSFb6HTxM0RSf2YSKY5NHgI
dgzfsa/g7AhKX2xcJPS/XOMlFSEKk46lKWTo7Z7s0tLpPaF/u+k+0Goafde9cG3D
FEPdFIvlm6qt9fB7NOJxneGx6VCviSGsiuRwDFO82Uj8wn/VslxOpw2cSF2gN2Vo
gtUxNfRiWihnvw8dY8Wo6J05wfZWq9GxqnW/zowLVRu37ImKtE3mtWzXpFWZJsKZ
L8rpcwGVV0qNgAiZ5xlWqfzKeWGpchyldnzwchlQ+uL+27k+E2YgFoO+vSPws0dH
XzTHHunub+nlKQeu+WNOUgu8M3m8TFeGOUZkN3liF07TLYo9LxDe0/HOeiF+qz6M
hwZeLWsh3zY98ofRtqVqZpRxrg0tjof/Ovi2Ke+74OV8mhKX3wziNG36E+1wAgpP
5MspyhZA7n8pH8opfdwe0pCROC25y2dkts88ErbaLFw7K0BHx6T2MfZDoIv4aoRa
xvN5V0a1V3wi5zeT1FEX0MJzk3UmPNEbAD+sj69Bsj3Zh2oM1bdQS8wnZRWVf4ZR
TI8uOx2OzmF8Okw8q0RHzssqlyWGrLpXD/4Ik2WPzdlepB+w3fkcJxsoWuBkhPS2
Uq95cQd2o4rWpZQxOYfMfA==
`protect END_PROTECTED
