`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHHeuCfQRTINfDDO+LrdctpXNM0XiOe+Ydk3zXFElZME32ZO7Nsw/jlryRQiaV1d
g2P4J+cuazjZ/U5LPE4n7Me/4tR/uscY5E8H/Kws20J3V2PQ6xdY3hMf6T3AE1Av
4z+vcAYC8FJmxjYJg+mWBs7MAR1V+ygn1wy6ChX/Y3cd7s/Bm1geynhlY0qPfXRE
bHxY9j4IYiG7REeTuJlcDe3kRJ5BTcxHt10fStp7oSz5UYitFLsn9tq77k69zrRc
huOrEcAQn8pGXsoo+g5e17JYCecc93wSzfe2P4bkV3ez1PWBSP+3pFEGIBVcVT9/
cT6aiaR5WQ8iBAZw8Iiir39DZJiwEzFvfgWpPen3NyN3Nuwfbmz8qG+P8UxXVt86
DH2HLY5oGIamd5SHooy3hG/vxRQbAVxZGkf8h/2t4JVBekPkWUKYpmelgAEHgArt
Omvdr6HjhLB2GqF9cEc0ngMSAvbZnHXITsvTAXwNEygvzCo/VBgwvXCKS8aqtSo4
9RMHTnNr3UCzZjzEf+IDkqhXUlEUZP4rDa0L0mu/GMJ5r4MGyGsUJZElra0M2QAr
8F9BiLQo2N7Mg6FxfluAC0dIlzgUSX4ZC1/M10ToZCsIMxInfw6C9j3ibB08/zmh
UE0p/g04dWas2GVFfpX2sNc8lLRzHmD2qm7A2U8i/l0ul/DKkVrmbYoX4R/owrcz
rqjHjse4OxZ0oxha4QMibGyMxR+ZG8y5bK9kGjT7BiZnngg/5oiPxEZdlDYOGGp/
124cAmwUwmCaE4xMUhTmKytRzDLEBMzNwB3we+5OpIhOd71q8/YzVVbTIWEaidPx
1D530aQ3xx5fxP9eW+dJ9T7B/R3mIw3iQ93KgDo/a+jaYPXgJkyaeRzEuIfE2PN0
IcZRVwBl0eRNrP6FtNvNHFuahAG+NPf0maZfLkaas1P0T6MSt10EFr6yDRlqa3MY
2khytRfffvLp3Dsks9/4YBq7fhErKMpI4AE3B8IoMQquTycf54lYnFtYKXEWwsCz
ov1GshOA75v9X1iifhl9Rujre1hESM1r/3+ZTt+Z8JIglCU+pR63Bm07Oe2YNoes
VHKtyODFzVbGAQ33VCpFGpao93f0l5Vcad8OzExwS8LMPMQGEcKI4Ute1U3HViO7
esljIksID9E6xS0/VaMYrRY3BwUR1ap+LlOvl1iIbadzEW5wNZDzzNSQmWNdrDQR
UibXOMVvBzss1oNKayw0dqyq2aUBe8iMK1wUHmNbVtGspvUjyhemz3CROLHMq3ia
wEKKJMcCRcT3Pafxhx40lXHlqN09fieizKnF6hXKcL94jgcTG0+HFzATM864ykMy
Lj6Ha55APhxprRwAs3WvcYg8h8oCgfGNxdseQtHpu5zNarVREpPW/mbnDSsqA60O
QkA+VlShMd7HwOyPGIXGt0LSDlaMwxupIbzGul4BDSt8V/dzIpnwK0tAtwdcqbRB
yBDDX8nkUDxglGvg3o0WmYYztWUfUhjhnMRpKmFYoAiFTitzvy2H6WCceb0TgVzg
+V+GSn8M1HSKwctaynKgN/MOAllvwf8LDKrQIGHrVoApoEuAehItRnzGM3mpxVQR
vgCMw/24wLgVtLkclkugGkUc5z+Svy5wkpEUh4kIL+gs9A7ki+ba2RcuxoyUPYZ+
Biqz2HVR5kQLGh7HZtkifj+lkY2KJSWyZJAH+lcKAj6u7V2jy9LOyk+Bf0DppakP
Aj61BHRbfk2xv/WhTTsC1y3UTmQ1zotoz+de/YigethQ0ojQHZKT05ghEfsjiosv
zmQ/4O8Br8VT1rgB8hn8+gq+L3Ge2NxrNqD69ibSLjUix1WgUEc/LRJDHlB0aiBx
kPRMjSYvBWyMH8BaHfrQMiTfhai+Oi7Whlrcs4ASJVnT/SiDBb0wG2On9M6ECPGX
saFJY1sVdfT3tIwDqG/EqMXV1djk7eoV6PwgT9XSFQdK8kmlA5inVNbd3HwpOYv8
lIAXDcYfdHJfe3KBVCuunAM9BM7kCyXq4uemgCi1s4V4v2wSnqwXcsvj+P1jk6cX
nmOgAJuXldy1s96c0LoUv5k5s8pT3TGZn9gXz2vw36bIPP0AohMMRaHdqB9tslyp
5yW6Lqm5KiR9X4NE33fQN5Z4TsuNq6kDqd/SA7lQ2mcwV32vYmGfLu+87zPBKnjS
xCYArjOeE2Qx7JmF0eBYz7TqTPOuxyqX5EwVstSUeZnWyS22+MzAEkweNuqxrnyP
9lJbfTNQMVCUVSbBKr5qxrdAXEnmlnw48LwuFvvSruw1np24K3hprvBXCFUidY7M
kXf1wMrik2/j1NbPkdcjGGaOn0EO+ZRXaz6UkFFn8YnVvE08lQ8PiUinsXkdrFYc
JZ5z6hXbRPE0HCHChcLjjqYUkXKNcJNKr1BHho84X5WdNcXHX1AdweCQY6NHYGBn
TvUkYzRnx2qqgB7xLpIVcr/85cHLDRTXcq8Fqb6DCreJ+f6roU8g2IjykOgnwvPg
6r22eTpef2t8CRavcPvDMsGR/qUnB4vjs3+YdMSpD/huohgBAXCCvIi0RIsEQ63K
wldWMrqhZY52z3sMoPoTqkc+LewFde/AAkbueS/wV4bi1CyFMuSjnF/JJ663JgT7
NMT6uh6aak/ih8zDVqFUG0QzLf+OeUYFAK97HNwQHFO5NMmjL/rK/SgkMLqozZ2x
v20M8KRlPn5SUTSa0l11QFR2qjVSUIrTQOqiGKNP8VnP+FYxHeL08j6aSUAuXuog
JzW/zVMXFnviwkLOl8sELza0QN+KvGhnCz6zlU6/7arfM0tnLKf2b5exvvuBkRmO
FFADTrBC4q6dYLXhsSOZf6cIIBbil6rcw7LrdfEulT9WeySGirOB3700e8v7Qi7v
323GAyq4LinJPe+V7w9LORuCjzKl94JqbR+boFmsaKqbKlMTi+bmrTsbSAFBRWMi
7TFqX7sVbjH/PplWcAHMC8NkBDXHomYHkLvCMDLRCN8u+5KZp53l+BIV4l65HCQJ
KTVMBeTGmgJPsPCjs/cEv8L+999YFsOJ0NyyIWS8/vMjOfaLdYxDajqLvRc1uMwH
3hl4zOfSEKAziH7A0rno6SNlAhDbtc8TEaqpYgHleuYR2jYaDXDgmeqGqE0l1qsy
lTU8LthUqiEc04AGecmkMLm3Ra7Z2hkUGnI8brVtpbzwg7QVGm66sLEv/T4rYMGH
sBtebTF4pcXnZnyFipCqeWfWW8JUvK8FQSVmplWjcG4/qUiJpHYFboj6gqhmSUU5
Y3K4iDTOVXBPhBi03jB30PmFzgGpuYI4/gnv6GLcyqfOMXcBOObseqJ71fCNxLqJ
feEYExORNFL+wxFnlijzDSlNXkMjA330rKBZGtpY4fgfZeRiIcKyF1Z8CBD+l5kZ
1ZK2yL5pkERTu417djRmguPH3VLpUJHLoJ3gjH2T2xDpGDv7baKXVzRWZzpxbMmi
//IP/iejPiIvV4JQjWRj5tTI2hsYXf6ba2OqJVxWxylnS86od+vI5M5EQ6KyTKzh
KnFIAm+7qGdB8qUsHqu7fp0zpbTYc7rKcyb+I/Xk1PIbw6syI9bP6exQoJdrq2cU
8pNFak0in73sxlOM4dWDzMvXGL7Uv6P9JEHr5HN2CvApP1HYWuVsmCjMNLfR8xog
2DukKjD33zY9yqE4OTFGSJMhrqTLcGrf5oZGYr1WoS/Ra1nYq9Qt65tGLVmMY01T
Ek6gGp48Q8my8K0F0LJ9ZhTkeNJ6ltCXnQzBh4gTdW6iy6D0R3QxKTfXqOyVGyDL
CO91E7DP5H7Gur6m/fTen3F4xdp2iiAdUZKlE87kt6ACG3zlLCBhStpMA3eE+AVx
/BBGKvWxyFcF9q4NY+31zbgHOIFuAm5+43Gn1WC6YYS4XSUezRiifFS+rvCLrl3F
YtTVumKgD6vp0otpoN2KzAmozE00bMzjDetq9zaZNnTLdgkENnbcqsI+Yv1sTJpF
itlCMtQCujUO8A0zMGYj9tzHDGfeJzoQg2Ck2tvuN7pRgLVe0xQjcwyorzcRLLil
izANEw81ZzrXMSZl06JS8e2FE8H57nzfvutPpswjLJjRuCE7bvy2xq0sAnhGCU+j
AONhgjqM5CQ7L8vViTN7yFZSFMySuPT9Atae2vLdR7PJzbhCynBpwZImKU1ScTXW
5KyIBrPsmZW0gStfgIOAQaAeA9aFjRRzmkgicUObLAoWao5L2p3+y8b+/m/Ynnkr
enkg+omPPbKzemzlrABbL1BxEgJepwJMRTqnGt8/MH/QB6Qt7InbnQbwdbkLdLMX
i/65ArDPzWdkoe95+juxS6yyMxFocJe7sGE5poLgEinCH00EAXzuS3nMx1fyeHDj
oNm8R4JWD8DuXsBVYO3ukfIPmH4PYfpNGuEztZAxII+mjlWuWCTuPbOB+01uyI/4
xgl60og5Cig56Qlao3+3e4YYZPRUj/VanaZv4bNiTEQCRku+2ZmqwEVGoWUrstUK
9Rh5DxkFZ+FRSN9H/r4nw21OeabcU62KMUPP8JJd7LAudYpZd5XOrv13tZ2AQCnx
3ySF5nRS9EanmWYgYlK46sXLboxdRYDZCZL3b8EZw283y3OUAj0qKd8VpvfUNkaZ
uXm8FrEfGRa9ci0v2j3AOAIY5xjGGMbX2wmWixFFgWzJGvZEeR7TvKcrlTwBaRqn
5yvcnNXWylYBA3cS041rVBc4KTv6fvka+oIiYfZg4kbWuEBGJztNJuXnECHVzW5y
5bmyjob9EO2FXY2CHMH8NAeYw9k2L3ewck9JiXFW0JNsFfC+QJXgILyp7y4CXDML
1OkuCnjeFs7i+oBmJ1TkhuTFbRp6XXrYdQAhCzLaAohKAAdS5Pcg5kX83GZru7yp
zbq3bEq4wUAw+yKsvuuo1nWUdxYU9Um1bxm+sjPWOlHOgPgM0Qz0j239dju4jHnc
BEPxHjnP6vfe8WPPGIdJOoyLua76JYM37lNrqN6iuSoAGc5vb8X3PKC3nxgeSOuv
Q3kdVckLaf6SEHlzSV38FLk6dheeydlgTaBtysMwtvmrSbZZ7kzptiyAnKz92wAK
73+I8TIqrt0AVuHCqBJn1Gk4Z0bRSckqMvM3PuLmWRCC2J5pM9v14koQ3cZ9hdXU
n2SZd9isPQ/U8UOnbCNAaQ/qV7xN6zbeiOuGnKT+DJobTuO0E1xP3wvPXWbLSlIu
xpgAWPby/2GQEZN9YHdqwNlhXX3qAm0XB1pm4mDBHavBG7jynh4mbiFMvkm8xS7D
VCMI1vMuyQ4A3j5Rh7ZmYCvE8cCPbwtSKwUTZUCFm0/zb5wPvUUKCgjSvy5xaB/w
vaLtxjEq9Fw8C20moiF/+TVlwLMcMLzJd3/fD8oVEukZixwR8gpfXMwPtoB2HNxk
CvzBhy50rlEiHcckCejoHS/Ho3mrtsu1edQhTxZs76U0oNJl71MeGmY9QW9r+ZM+
4l6YhzTw0cVVEQHvuBnyStk52eTbb0kN392CCx/MbWBgMKZEUCaOVDYY4q7RzV33
TXH/NzBCvi5TRfuRZZmEPx+KPgUcZxRu+cVqOogPWHK9nadCnqNGH+B7VaXqTBz0
v/BK9sGOJLOeK6i6k2UV6lMjhkhiUplnVWIYnnC36c7dj6MBcKocBKT6mwvqf9r6
IuxZMjsG08Um5elZjh0bMf3JeUiofUQwn7S50YAYY2nKMWlkHFONXxxToe9hOYIB
/H7def6+lGamugy+rA7PrFZPs5cAvAi3KkrCFg5ndSHdiWxw3aI1OrQSK8s3Xwci
B6n2V518tqd8KdA4IzVmGA/qy18TrGmu5RCNMRNdCwI194+zDzf1Gu5ou2pXq06m
8RPamBiVD3cFVB4H7NTgQxMBA1tbEgBPNntj3L150Gme4QVG7GIBuQCNcic6u9wu
6E/Czbv+9BqtjjyZiV0kmLruJhOXL5UGmLGppjTIAPFpzYOtexs9IQLefPJ4eaI+
vep+XaBwLlMFoe2exfgWWc82cThcGPSHXN1WbLZ7ZOCkP7yc/VjdDM8nEshs12FU
6XXmSXKUGwRLuCvPvUQgjE0tvv8XdZ9GibL4vWGH24uFV7wu3d7tCyRl2wEqh0U+
QHXfV+Vfo9B67ZW8lstOWfPvi5qA35yr/3SE2kGXtf5CSUssZYNf/DieRGQawBPI
j8Y6CbgHaRa8eTdfSiwVKgc/fzCUeaxAjrkgKM39mlOC7MlwRfP6WnioQwfIkgV6
oNe+UE3OViVYXqFMXhCRO9q7bft2x/ZL0q/MY09TJ5YhnLBaPMmHo/BMCP70tfsC
JoMWnECyu5aznhxDb1XFTv6SD3XLVi7Df54lwYpQgahYjilRh5TEFUXtt3NkHPd/
JWD/2T+YqId20yA2G6lx3g9Wxhsbm2AT9KadZ5WRDG8DkXpomuhtx+DAbh7FCZbN
ihaeX5xoG+hUu3A3vVNZKVApjLX+6tZXsVcA2NDshl3YDeXgnUlCjD8CaIRYEafL
Pdx6OUVCA1SpatSNyDsyjey5XiyqcAlmUpb2ok1ee2/SjDoWtktrDkkU2yMFejza
P8TC0RwjYuGra4mAN8hy3pF/gF1LWxz7wV3VNFly7Mi1nAXJmepV8I4a5WHtF3Yo
SQgapyo/F5BydF7bAlTKPV3m9cNmk6ntQ8+zD2J/QW2ZOv2jyUKZSb0l7ctMtLEF
T8ahK2xyPd09aVKh/Pkc+Tz/NmcXbrn//vbvfRpWgKkYQ8mbefPw/W4uBKxCMEdZ
eaz2i6JkGQEC4+EGWsBl2YeVuIETH3tBvMU6LaWGwkqpp2q+rZ9joMFlkibUahfP
Hsviz9uPXhYrmAWqrNjWChdOkRQ3IChmwVzqKdnLd8WiKCqzVTUAfUP/U+cKoFLr
uAC3mvVrTFNO+EiqxmMG4OnIUOBcsHanj/KyMb5Znp1lKcXD+TilptqL11qgKf5I
r+i8zOj4v5tBn7P1FscY8pbMwKKcqx+AvEvDupUIK6yCRn9UD+RnpKoWvXoqAE+/
ZAssaxDJUCvCr1V9xF3DVrdAiIo0Tr7GuW2I6199b4yUmyQqlky4RiG8k2fk1z7r
eCdrZPw9fTrjwNstlHAc2UaOGwAmwz/yM8x8RPd/ipMrm8Ncig574BgX0Q8CII1U
sNiYJ8ThxOVasbqjbleKKfdDaOLqH5vdDTLyTUC0jkzJF0IhiaZZRbrP4GpA1X34
n4qRqAxynZd+ouScMMjy78iaqhQ1DyTnnNjUeT9DMoRY5VUXS2C8aLd6W2aaMGOo
IRqwN1fpPqXqv7lGurVxN8lpe6UGSMoW8F2yq5QzLVkwUX0Suf38SI4Pgpgde3qa
DZ+Ty4F6xijogAhdC0Tr/UMchmaIT8Wxr9CPuUA+05Hp08LEoJNKCgfEgDpirgQN
vE53/0Jgtggva3RXe6YpXNyigTB6wWXjtQYy+dPgXUPZGay/w3OqQU7rG6JwEYkE
32Ks/xvAs6vy9YYKsZnOX07UFr9sl+UnOgaOHYlbF3Prv+rHTgkGooP+CqKW1t0o
mGHDSCjuMZeXrEAY+/+Au/H93KnOmkr7l3Ve0WjcD4evig1D4C+oKLM+RUMqzF76
fJrPiwQqWnVbvyi1JDaBgGi3BK0CHk4lEXHriWmZsFKJB7KSJdHSBLP5X7q95N+Z
Q+FuDxqzahVSp8LdukRy0TQArD19QOUB7Sk9Mr+za5v+SAaI/yaOoNOFhYU7ixuV
DzIJfKs1ZZOcxTL7IV+2gfeDKzptgmYysU/t4Qi04Ap1HiNV91/1YT5067RKNDly
nX0muy0lToZo+vaJnY0y82F+8A1sqoo6k72YLeTG25RgfFwNsJvG9jllGAqB7JxW
mbSFxtGGsAO5bQ5CIa4KWmV2avyism+hf011eWTvb54niYZgXoTHz14lfGqBFF5b
wOFJgTe3jn8ZSehVymKFly4ZDkqUnpy7EnYhmFNdv8U3YDcna5MR84mPlJXT3wQ7
JRbh/0y7xU1Ng+wUA+pcqq2yp+sDZUr7EOTkB7eU0oKQkW+wtqjbI2I8v9sUPc9F
ukRcBzz7Gjg3NyjD+K5EtSiELQj1BAmcIqeiCsvI+fRRVtiSnsQ4CR/fea1CfcOH
/6musLGCjQHxho1KkQKz493vJ3zcRuQBoi1c+8EYlkylgPwyaRjoKwPIFJzj5PXW
3K0Ugn32+7HZVz82IFZDio9UfhgNEm+Kq8u9JRmiSbEO6yPEKem03Rc5tEm1h79f
PPRvGX+yQOTAps+l58UWZ4Z820mFjDZwdQwD6+zNmUzl3f5SmGG8vFzVTSM48hcv
7S7of2k1WDuBFhlWYYE5J4pL+/jc5xHyjbk97TiHAB5wriNDwX7Y5TjdJQDJycED
E9gqECD/z24ecE2NGYewCefWx9xeS6DA93afOCAjPuSzVQtyO+NPVQH9cfBTTJCL
Sns47VixLzwRlh9684YKgjvPnqcreFDKEe3us7GotZXDGDcEwh+yjKs85uZpabXM
HEl/mxXSMZfIiLtWghTKHz6udTEIMUqy6iDg2bv6JDB3L806oe7sWSpuJ818fllY
vlxJApOzQWog2VaIGIOEPwEICW/VzC2O3PEmruUIW3snYEEvZf0BFXhSL+ez488U
+hKx6SQQ3bLR8FJlcFeqPICIj+rK2RsxSHINxqYLDYqjekZrIiiDhegg5FnaPIG0
eeTMdTrARsamwzMwoFqNkcMyzu1lXFCWaWJH2hT1ShU4tOnfy019CZvKuc53bKBx
njEd2NS/28NKjjFN+Din7wTApvxYT/OB3hxQ9Uz/Xhb0z2mSdgsbFuKx8fr79m/D
7J4y9JrsOQgud+6PhWgCUgwPRQ1MBOUsXf5oHzhj+WRbZbkm2IQo798DNQ8ZWC/+
0eaxOjCJihtjXBI4jgONsAGPWxkjpdr5B81JrOEmRHK1MnbrLCd431L3FqrRjwof
knaGzvTiqRz9m0c8NV8ORCbYg5Bt0k0+dglTjAm/04kKKSnTwbSj3x08HGxuAT+1
e+osLkBuhJn3l0XnhCyWdFK4g+un6qzDy/JzPtK2XLeRlW8PPjBXE10Bosre98Nx
WRAUp3fC+r8v7CgJzX9TCuxwY+wUskFa74K5jkDziNCNGWdrtJ6d2ASDFjqRZCRk
Njs6Eb0IAwxP7JgwSD9g4pk0mztxPyI9q++VK14TMupPwzu3LrVGTHJeiW+MfrKD
9q65uyLY8EmwLwEa7YHnhRBdenZqYQsSeLrseqbzj0c/5bT4yTNO4S6pKMtYljuP
527XRkDHYjjY/vNyD7mMekCYdzrme9UVp8KMtRj45oj/aSXWDKCveo2aSj0Yr5+U
eOyx0KsoJG8kpbqzWczP9m+GQeUTDZCPk41gNDJj31cfWyj+vu85O/ydrYyzAc70
Ov5Ak2bTXkMMrZaNOyLOu7r+3az6i8cLpBRDxvYfO3BNzUQVRetES81WwxIGpFlK
7oDfnT933p2Ugo3CBbVFPUy8J9lmdzqBLvwHI8O6AtKRvFq+72Q+/hbxEXscUA5o
L/+zM2g1bv+5g5TFp5I7p8M85axllFY/L12ARMpaHhnYdYJwlW8EiDyHRuVzN0Ca
1/b2vpH+EWyyGNMsMFHPQzfoHN2O1rPvOo4pkWm+kl3juthOFyiAMZO0YGzXsADE
PHVb+OgDibOtkfvKIUhKd5tJ6XuQUAV1nq4Ghxeg88F+niG652um7sDqDlh/Wv3D
2E/N9gc+hIERK958BonwD6KKneqQ7eU8M7kwJJTzSYyQ0Qx/+LnvvGWWKL0xYr+X
D02AzTeq79eucrRIsdfoGAWFQpGNhOdKksbwoeTIG52x11U0AKnElHiMYfppYIQ+
JvvtNa5H9J/nWsMxh47lvO5TRFLv31TGn0BFlyuMcpm8YoE/jDJ6paGs2EXNVsPv
UI+KFvEUBuXCXZEKET5rgF4z8q8IfwedSiWUB6W0f9FS5KdsJcXQ7z5zk5V3KTEZ
gx7N1L7Sx6saSF2RKI5yh3JmUr7R3/gocxOGDqmCGMbtgM3wyTYXvmJRrMgMPDvG
E+3rIJBzvAVBpW2ORZgRh+Q/gFDWayrZTaKROGJv/lJdL95yUuFXX4Z1nOYjbLeF
Vrc9wM301rG2VnJu2SYjkhrq0HmIQblBAmJUj5YchJRWYDgqKtG2GKIhLPGxT1Cq
OAOTwJy43SR5xG8DZUUMKKay/e2B0dfsL1SttAxbq7kLohT3ZTFES/e8L7C3LU5c
NvrovxCN+7ddkZ/qLsDFlRFAsHB5K1eRKkdvWh/Savt73p1rkaF7Iemq+EtPgQKM
dVuO1+OiZiQThIi9c/Cw9NQELCCWFlIvbgnit9vMN5BNydK0mhbuEN8Np6/xmPfo
A1or6irLARgVHyXpIPbLUpInzFyfxdBV9HBtqPk78nZ6tstiyJx070nOraBmjUnI
tBUh3+3alwam2uDPKeLnMnFOptFqnoOdvDvwumoFtZVZgZtVmfEwqX2Q5cV80ITk
QfFBxMgIAB6F4Rsz1jNi8+CDTlfvE6z58HwJJ1RiGyqTDCh6iY/ulS+kpD8RapCk
I+wfyIFMKt0zH/YEs8Q/8sinWsEpnDMpFnahhC7edoNlhd08QrEZZ/KRzhqayzqD
6WkWVA5itdczeJakeZDSE5VJSfWfqhaOX/uUpfJQpHsWKYv96CoUy2BAszKvVuDG
lnmbDfvYq5TvzXa11izC9mHlFFb0s3VKkNo918PE5qGoxBdHOJ1P8dio3AMxc/Yk
hYo/fn1dtnzztzATiQcuPpwEEVvvumQq8+pLeggBRkhSdVVE7YadWEr85iocZuKZ
6wVugf7YK4gfLb6Y+Wo6qcXrr61/gL5ROPOWdzgXYJw5aPdHIQU0dGXIt6Y1kV3R
FQ3D2eF9Mf9j21/KuuJ0zoEIrlHyFE4IFFQYLd0kOBqB1hbSyJPqIFCS+TXTgHqN
QVDOjLXuxoo1HUaB0CFE8i5HFDyzA053bc9HsqX3hUzQwRIRCM/bvbNzPWt/sION
HBLYWXTGK/8Y4SxVdvdlXjRDdK90hwqEFafbTrJPuzk02m3lgmVO3e3inSMInIw7
u9jE1dqLZdTW5kqrhY3c+e7LiV/HxVq2SXOOkY4YSxQNVg0YRQPOuHQMWA8KIkpg
0IWnr8vch6fj3vsz9nQVr130HnHm5sKyic962jwaTRhVpSkjRfyJSs0Zt7Yf7Jhu
bv/8cG40IuowUcgqlRvxZ7I67S9gqk7PTtKm8SJvjQOE+PeINvMVmnaZSOEkiiDx
bQYJLLC4EXRBYI1DHAQOfl65AmJ8N79u8qi5RKvF/69M5qgrUZcvQmQmFlkkF0rt
vuIUaqitJ6rG8X64WTk5VBplLfMF5zeTOYLL6t4q9PiwQ2zkLdfizIpKVJQD4Q8W
YrWKmuwfc0DgfwNBkPekXHValxwya1RN/3+04RRLn1H444xl+zlHJakTMIMPPF4C
ytdlPncV/3EWciZNgUcutnfDmoiXgbAprtscoFUHgdyBRFGkRyK0f5G/0ydUTVp3
zlUGU3+EZD4zWLjYig+vIr3mmRroMCmCTEoXgorm24q1yJbKwv1TS+4viYUOANvu
Xdhj5/Q/+Y9CMSvEAcMC0NJzUrr2YczJtCxWyjZDUIxcQINNdjv5nd9Vu4H3f7K+
hZAhgdnrCCw/OTo3vLTakg83p20Pl9Vxg8zcWAQL6YyGed5PlmVLRE418rw6dT+x
HfwAd95DJIoS0h97SSs9S/+WS/rBqlHKOdiKdwD8E/hMQB/Syy2KExHvzwekiDse
yDmhniJuSNmvEtvVNwvmXUvG2fGtAMeUak4G+HBGcTits+V/GvFwGvBf7sYEdHVm
OON1HpVe8pcFajwCo3dMsk0yBvCE2G1D+9VinmU8tjIrH8Ukx73jIxU4ZDvLmSaG
DlnyL6uFduduQyYtzJCZZ3eQ9xrUJrmGj/FxiykKmhvcfN+DnqPMpyRyoOir7xW4
9aR0VQt/BeVPY6FeHBTAKUSBBVjExAvpu5DUL5mVg8UhtrcepV9o5G+UlFeZ6VYB
iMRrpAPc9NyejS3t7PbQcYCZ0DmKlAUtsTIL+lBZxA3CWVVXByW5LzcPnw10YEho
hgptC12dzYGcYeWBUD0bZ+srDUYue8FBF9bxIhheHDjQ8tWAD4NRE6f6MyomtEy6
+0NuQpahtBnoBuLjXIQMUlsb1vdNHKFDtZ9DKIeSMNVJGrBVfGvk5V9dGHuWJ0nf
Fw+ZZa8SR+8BpJn+fBUQvbQHhnOziZuZx5j3IOnsNIyCqeNCVovxHYdJaCHjJ64C
cpr1rbwEJZ7HUzHL9wwt5AdWIwxmQBStQcJORH0YRk6xjGDzfyvRVxyBnC4VCJJ5
NmT69s5oD8QjhTNZGcC3Fx09VpZoJnPf8DRwrx+yGZI9W5nrQ0W4M4YDfGIcQXGO
9exxcpHRlatsmuwo71oJ8uiKp9aNRvEVdcQzBwMiqWsgGgLkFUC1I1/KT8K8HwRI
FrePXXabz3n97pG0LRw4JWm4ERIJZ4mpGCP8MWxTlR8c504DqA+/AQQvfZ0gag9j
G1kkpfwJk7lcmP5ywTonbMbUVOmi4qQpK43rzQh84jFm7evtC/RU+beStP1E5d1Y
OQ6FInFuShcFO0oRHt56QErKh4WhXIn/faLj5f7k1ZHGWiL8P3FvH6xhkVi+u3YE
MZzIcVYcLJ8o0QcRVC1cF8Ro5m9j2MPkrnzQ9XCZ9H2Vo3E601c5w3TFKNoiYDd8
2Mq5Fab9OqhbqlQNwn+aDHe0Rce7sua0OZg9HCFa67Y0MV8B1dQqV3VZnkXBU1HC
THETWg/kS6zlzyksyLPlX6jU1+3ikMbIAymh3Ed7msiiaATNzoY56Wx2SMxbZ5zQ
wdc+HR/vyKJvw6tEyge6fMa1C4D92Ovgf5wEIDhSCxTmH5XAUlOE/JYip7CUBGxO
KPI3Q7kqqSvvZNCWgOci+6jw5ajhPM6Ak67e5olNO2WvTc5HMvop81ub+Ummd+h4
+cMhbn4sm+BReyZ6mBZX49BS+gX0Nhd+41qSxQJdPKPvrJHXTgcUFXQNTcqzKyhl
KgadIMg0Apf0NS7GKJWBgkjuMRnFUDNMYeb9ksT846DCd5GcsMjLyW60NrNIqLO6
QGIFjsMGJDwoMIww6om2OcDGwpzsMhZrW5R0ZAVITymvBcvQ3y6e67I0uu4AXCFb
g2YJdt3QaqdF2pBMQUENI4ahZPnMhNC+EStQSAfIxgGUWZOBk/MV4Pg3DQXvox2h
dwrQLXZuvva4cTLjmS+XmVjTDJczJRo4gbgYdXALz/gpstfa70ty4Pp31IHbYAa5
EDLoveCfmxjIkipYV1YDrqu7ci4XRXVNFvy0KCAGFviOtI4dmFI4ksVUG/+Iepez
MlE00YeKQWyIZksq72EloZDds5Q+ouAmXm9FXu9Pe2t5IDXR0Iw67Jp12PHHz17m
FqvdgOuBySRT3G7hrCJtM5rgvXDjy/eMQ7cRxJir+kOrVpTSb81vXij+xT9ED20s
GkWun159OU+vUTu3Vv8MJOYTBagi44k/SLpBCtuuuCAQCjm9qfoM+f3lPzKsJVFP
JRdePgsFhOX1FJQOeWzL+hwUCBggILziuZSGHEDNd9W3hB56pS3mTgSGlkEMwuUv
bEXY/3DbSOnWY2mni6RNSMvCC09JKBiOE4LkgVNW/xCMWKvV5uEI3zLaTqeYF7rc
7KNB3Y6ylt6lOQsGWMpSJnZY7l8GWNzBJO39AT42Mrp0uHa7KSf6a0QQdpywtB4A
Gd97YQxKQoRW06P5UVIFA0l8x6zHfa6ffu5FqPHU1IHaEwivK6QITdLi4JPhI47f
p81KOuJjIWg0W0Ssm4zVYz4vni0XtK5ZJEoCuZNrqnUQ2LyzXIHY/sqeo4BN2tp0
DukLqGcVvtox5Q7Hi/PXfn60+X9JjLE2+RSID0tYtK9/t0X0xxGpayUTf7BYzQ6E
0u5XazptCt1gvcdQly6OfZTYO7iDJY/EsVI2ShnUePeamcXj5iaJMicOv0ktcOIi
EEU+ohXZeYEMSXRCfuTF9fiqhc/hSaP8kl2TKLgwPiI/8P1cHjVqchK7m8JEkZ8h
XMrRxE+C7cSCN37pXLzxTDaa62zscEAUAtVnF32Wc427GKWykljherFlllqFcPFP
d7gQLMLtQoeoeOVQWW2rIj1M235h8l8HvcqOSHha5YMlzBsoyq8ykSKXUaKTTiMs
8jy3kjiRb0GOpthBlJkY/hWNVUF2NsBXBMAo7PVhdtusTgY4aw9eC5zCPv7E8uKE
Ec41QHGtb8gTlJRDt1tBsnR7Kg1rsb4gLdAs3lp1VF5cFAgtPezdShand4RD5uHz
A4/GIm8oVySgtrY6XtrdL3+/uJtjTMB04PSFyMn4/1PpxRrAQYsGTHFIw1yy1s4/
SvH0f0N8Ll3czrjGLSCoVK3Y9ul72/5rKY4TxCYGktnJJn4zpYORILIPOULAQgeA
7cNE9Y6Vxs2Q3jNWNobD9t5w8GwbkU8ZyiHlRM0P+yemRK2Y2Szc/WryIzfBSZ2d
vO9x+OLU/TXivlte6zCuvlXTxeq6DcYn9DtBwiN1b8E/DT6Ci7fRYiBTbUwcp1+c
Smzf3Qx0dwF4YKOxindBW0R+IofrhpjqM00SCpc0rTfW5GynFmK4PuBD8rM2TZKX
Srw29Wd4y5GnmsP3XCiIARk5DoyAnh/UpfMqS9H42Y5cwDV0Jiyq1Q2GhqxuRUX8
cH8cHXSwXAcOCwWTwuoDo3Lv5y1AujOXsMSamipZoQkvaEMqn2x8eBlYBi0CR8rz
TKrJovIeX7L4KwukPqIPFJX6kDU80+vIEES9cBL0XCr3rzKfr5VWjtwjEN8YaXEr
gaALumKmoxGiJB2fA5PmYSTaVAsXOgjwhhaspEjWnDLNlujXJ7aUS6eZVSFJevvW
tFYczdaSElm/FIc+hWsZ/SU273B2fqbN+fYl2NlyMm2k0duHp63+v3DrlnMHeFpd
Rdbspz1vzTDFXNudTvcssu3R3RQpYeRKpv/f41Wb6BcfXOOEX0xTP3tHeH2NfXOG
j5/wWLAlspSvjQ1POC3EagO0OGQRWlgwrcSsHGTN7v6Khl0KJUai6pf4acdL50vx
TQnkjOWpGg9gMvDlPYh75Txz+tWe7DBtcAVuGyJ9yjb93Yv37i96jDGcVmynVpxk
0Hfghdykmeds1O3sJTxDLjkOp5BdQvTlAvmFLMsnPq8Or6gyqUa2LdFzrPsgQd7t
OjtbtUZRccYgWg6KCfJ2U7au9S9ujoSKMOhCcodfJVGFWqjSPdwywssrkNBzRpez
RTJ7NgK0OGycyuMRLvNaRQW5eBSArwblWJVsG2100+NxpHtZDhn8xw7KdZ/OOwwb
TcgwYHYt9dzOhUxcY5buKuvI0zCn2/X66Zqc+FAnZqrdRG45sEe4a86FUWsvKUit
YwOcEHZoJ3PC6AufSOXXJs+diim0qZHtDU6yO+3qdXpvF/XgMBEkYxzDNkYxBqIu
zSZQiXc6pNzaZvrWefKMFJwbFqxDjW2tN+lX5KMOqmqNMEUuNxBFGgjzzeVJpeY8
4Y0dQ68HHcMeaWW2xMl0i4BlGd51zM4G5yEPolu9owj8hMSOdXWNS+6W8M2ZPS+k
7DMukYMkTqDPMUfNFkENrzOMHa9j++Ml5cA0/bUj02QDIJnFTYEfbqf4OPT8gqB9
fvs95lTHddLn0vHW99KNxkAulOsskgomykQgZ266oxrNmFB7o2TCJXTZIyZUP7RM
5IAhUdVeCEgKQlVKuur7EAs6Vzl7ekOsozxpZCTzfKIOq/nKe+iNog8GY7vIaiFW
rXwiP8N1LMnxrdGQNkenNwejGSOY2zGcgFKetQkAThG+Q8Mg1oF88I/5fzhhTlzA
axuZsDoe6p0q7Ma/J1mAZbxvXnyxXQlbYV+4XbFwcdedGQlufp3g4cKH8msgDUCn
GDXuc5TdXIxz5y7Eax5H+gIYRucUBspqzFwbYi4poA82dVeezGNIXfNgNQj5NPKB
vT9Qrz8eaF6kefyKTxvEWijW4lSF/CNk6wCh536oBSJQ1mVoa5u32BzsD2OryMQ1
jpcxJTbVvHdYYYjQOzQHcY6/vjgmCk+L3ESkYEIyhhk3sOXSXxhzBzF0TurhfYwX
srT+5gUO4m1wACaUrJO5WoOqXrVhQuzeC4mU1QFGpS/hKbtiM0G9FFhzKUi1eez+
WNxIF5InqAadP9GS8b6fXqH6gdnpCUQdH448roSQUKgSJsp5P9685UteJFIeZAFF
GeSKTd5ecN0miOzl9ribbr7k00TGw/omWGV0oNu41S9c2xHE7AKrz9X/t/uLBH7A
Np+mf4w/Wf2xx+fdTOBYJtIzU0VBWs36XA3GeBuFhac0UBi7E3Ykd2rd/oZQmy1l
V242Pw/KIVwktJb1Wt2FLJ1HLyzNiwlnYE/tmGD65YUXOnedtXTKhG8yQWTB8Dg1
T2JP7aQKr82bOyHvxtGzvLjgE4n5dsFj1yO8jCX03DAaNMBdSbxGz6M3/0ltDVqi
fuuBQPqBORHB0vdvLQurW6LFWaM+olpYvwUubcTqLF/9YdYBwJ3B+xtAjJjNxQLp
03TkBnZvHRIJ3GZNv++CtRtqL0CA8VktaUjlaExQPVawaKQCwzGzwTbDs15etmZG
LBZCoATCM1IB7Tb7iElx+rMIfC31txP1Wt5zA3RZXaJ7EDi0AhP4lmkIjjV4TszV
ppU3QuPgY5mKeHhwhPetPFzf0Z5xv512GvOyTA2u2bLbnJdkcORIPKdlKH3IL8+3
Ry07VQ9THr0CSBv4BfmU//mmBkVqp6wrwYjcKnzzs3/2EtAsE3qEG3HJ+1j7n4Jg
8BHrv37R3V7t6k5KU4sY5pSNCHPtVuAVTgzzyYPEBw+jnNqybX1qEvQxxAI/0BLZ
9+XebFDdCkAPphnU+AnZpDWhJ2gBvjR2WfHcoCI9UXbihODUCb62djNwacByjyk1
B8rJovaIyTr1g+ACnaNOMmlhw+6A3xG/AOy2LQc+YNUrYCwvqZh7zg7FFNRMddW2
9zuMY0ygYRSTiIbL65ARRork1aKBuAYcXK0n3WU58QLQvUJLNEFeVIxctaavmbMx
1hJWYAPOVLLetdMaRmT6sy15VMaLgfdVbe/ppbpMwVVslkADW1kHK/mcdFtIL0yo
XRFT2p9q++WDKnX6SVJHFqJTd5y4uM+iP7vxTg178P2sUKjS34eZGvs+UG5VIk/Q
2MRZU9QByx5+z4xEu4mbEPfyB1ZnKmhj8hqQgnVDIw6Dzzo0DN9ey6XnqU0fGDG+
K8U/a1UJLsTImjTKq6Bap7R2/SNjYUd93Ir+y5iEaxXJRhCX8Kd5ss+g9LHw+mar
m9aD2neEyVXqejrZSZQMshOKw9NePa4TucwNQhzmq8Fz7Q/JeZ8Tcl+G3Snij4ti
1d6ZpSbcsOPc4REANnMGatzgNHeLs/mIarkCL+ZGvFAmZObJxsgRzdVK7BIDROP4
y3aDxvtcbzQ5uuBlkATL9r3+llnVK5xqbO8dwAvo55pzqWX0u1V9IIxQqah8rsmk
ErB7KVXB319iPGjAEcv5WwRb0uMSaIgz0XE3wUE54GrAcm1TdKaJcmmToYVDyfzt
JxZk1cIug2zwbcHxNzZRxAfTzRnad56zcYYTyrZiQlQGbH7Ixnq25DnZZBUreXkz
hc/AqNPjKGHGaFkVA7RuHWl8wXq+zxEyH25BCEe9hmyQNmXZgmHiaGKm3++1saG9
GpL12HKSS8rTwNB9p/3UeVIIDLkhSxUf44+Rt3W8rsNrkxRWxem8Z3L5a5kO0wgD
gkujB/nNEV01jfL60I3tMyxkvI2HZEPAQpDoX7T1h3W5H3m8oeBFGXDITPy9wgp9
ttuZxf+pXTQzggbal8NBMMfW38F6k9XyQgtdZAItUo5QofIDE4IyBL1x9/Fzng6X
18jKMHbvd3irU0GWUbGWlcCsUzr+Y89SQzt0mp+Qc1Uh0Cfm8fhlDIovFB0O9VNH
iP9Hhu6vuJIHwApX5MO7QmZ+F9dJ2uTuMcrbEVI0nZdTU58/GFrd6/RLE3ahZlyQ
SUQgInGjvKvblBkMuAk1tSDml461irkfnc7pyrCm1prrR+TP+XgV9KUxKxWDOnQ0
vMLplJVIqbbvyfOL/d9I8765/Hj19aIZupLlJSSRpA3Pgo4VhSvaK9AT0aet16EA
ClfI48/FIKEdpTjtmuoMpGxfzGH1FuQ82f4zsdi2knn14nb+QIoCawb9BV6NrFbY
618FCFEFG+Qw0bp5jm+uwFEJBMupPSdoHW1AdR8q2B7IXK0idTSuinkgtis4ug9M
HNPHFsaCipaL/ppzQHCjdygv/UkppjmmQrY3vxEcomXkLuU/WKxQCl7OiDLWi0Hg
+Fe1NH6tZRKPY8dwt4jcy1IcCFN8slLTUPr3n7tljIuckCIeCNs0D+hmCV6uhWkx
1nP+CaQw/E3km4hvrJamao9vusGn8MwZnzLwFr+mYAQUVlZI7/dMA0M9RY9Dho3a
8x3ccFy0W1p0bkG3CWS/2AmToGjNdby/mB1mjHd8Wgn0PzlIoIS5Qfdcl3gZQTyg
wa8bTZ1k+PL1rRR7WByt//ouNf0l12liDTXfJ+b0z/tLGsIlbowjdKa8PJAfES4e
Pq91hroRWszb5bc/jbnZaFsMwIXdkkjvw/kOCraNSKHcyFqH/h23H0S9jcfEkYiU
gwewhlFDSNjGX6KNovdgVA85QVSAVL1yTHiksXnGNzkH5HjzsSK8WT6khZV1z864
lcTd9xnKZmYuzb3DQWmVtcaQeCUQu06mcd9/m8iC8j1WjUv3Gj1ohKzkQ2vgEb4C
yPzCcmwY6DJpsAvKQ8B8WMqQdGvV6BJyPQgLiBsFfexRMfVSEBuqr88pMK/6idzZ
lpHKIXGfI65xtfeermjuujUDMsdiRK/fkb9cAfzBHO7Q0IFRe4qEJRq29nMGr8vs
P+w8Zw1q0jWoCMP9/1w5UAluWencu+hYo/NbvRHNP4++5525iXIvIBkOw2MNpB9V
4QQ53HcvBTsxIwTgMcPdaQz0pp+Kt7fghymB3rfxXugXEpTWZMfPxwEfVKZBm+b6
2A3fbhPCeBqQir0Rsdt1ZOErP2VLl2KEHrH/nTOFuO1bUhyrFNviB6p+RO/PuGZI
0aZOE7parDRTDG/AkDlZuHDbcMkUSqtWoZ4WSgyIcW25DOcErIWRCBVX434l5tn1
zpgbi3sDFzwFV/CbakbtoA2WAd0AdC9XFPEw7cobB8cGbwSdbbG4eX1NQmC1TuXr
LkjSw+OjB4EfAJSqgDtS/gEoyyACWr4gVBOXIbCom59snkrDqwh7EQFTVuu14UAA
OPEuxeTymkRya43KNnxxmNjxIwHjBdghqVzqGAIYr8IstOHjQ8t7aoa83yOLpf8x
sa7eUXgHN4NrRCgrPUM5BWKPSYHRGGKcUYRelfGqz/gTvuNA1O+SUMdq6Hn95Xf5
lOg1MYxgLJegHLavk2gOoR9N/xGlJxINcGBRZMeHpiTdpxvy2jVtp0EQbEHpUq7m
oWeSLQiD5SaFM+QHSYQvnFjXyr45g1iyc8bnHP1ZM/HwsISKRaB9Hp3obLzRQUAp
FNzsbCCIXGjuWs3tTLFkaNwgBID+Xa1K/AHe0PKwnhkmf4Oqi482K3aZXDA1IQdi
2nKIUYmnou2GdV1cPVtSWvuHzP+WYQxQOKTWbbeCAtJBHVf9oBES0AF9u1VXdq/0
WpvxUT6A5fKSWMjWCUwlkOE+etxRgJq+uJRAd9/TTwgg5rTSJsohTKY3hEJbacP9
1owQC7Zuxfu3tMbV7Up7uU+8w0YuwkuN9yZyduh6v1Q+Ab073ZuBLqmJz8qeorMo
9NPfnIWt3ojNJaA1zLet4JmM2Yw7LU666rvD7/mIhghcVdKmz6nnj76ra+9cLxTI
+8jBzSJVwjK2jiTNvQovig==
`protect END_PROTECTED
