`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MGOo5iF9y1VKH2Zh3KFPPW0ooelBg8Sn4cwGtO50uKKlLxParpjIEG2Tb5WFAs3a
IgYR/DKmbg9is2cT7HxQNyN8eK8ZQQzZ7EOjhXebD3Pxwb08RvLErC04FS4DRtAg
KaFZilcabCZRm1QB3IhokQGL9kNsnh5QL5cmi0r1iq78FVbjddVwoDc6VMD6jsJ0
OrLdekJG6yCZfoZAc7iVRMeesLsrurGtFlm35unmPy1D6aCTsBgiesLA27kBL4Dm
lN0oA4R+JZcV0I+ZEO50VAYr/OPhPYoSNAeTn2TwiftswiVZh5Hh7BEC085sJgrv
uxBtlEvA+A/oOK6O0dX3upMJLkrMcj1K+cmT1dixLpHvzAnbTLRXFqtCNH5EQT7Z
gLaQFAzAKf8wTK6f7jppqJ+xj/OauUj2AKl2/ocO0IojNzxU39npLKIMpcqXEmB4
XneeO6aK5rYKtJr5Ty5u3LkN53iGAtdlyJ1eGd36XO+u+b4KbyBYLyRcne4ROxkr
R+plz7m6z0unVr7CZlFXl92WrBZSJUezfSBCtw87pvK2izlxBtZH+UjsWBKgY03K
+E4t2GExvvSzhqc8+dSCbA==
`protect END_PROTECTED
