`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W4aKJdBhAF/fHq1pQqUaGWS5cemm0BV223urwyd/rtrx00esGjxLyixkMWEgfios
S+mOH8Il7UnIMV44HVwHhpAUL59BmxUfXzevnLPUn4fbLUn9vlEU+IZzyVGfJVwW
QoZXFzEp1MJD9WBgx0ArLp549Nn1MQMXy9quINrDSzCKb8E5EnzZVVdyoJ/xTtEu
iOO8S5JOcLnGktd9HjRWlZXx8rIwI9MSSltVJGuusgOZPbJADguTDX0tiblQNkRI
q/ejIiy4blv1A7fua+JOP/4HwBsdxoCyIzSeX8B6FOANg2cTZ6HNutA1fwdQEHH2
NLZm+mds9jpvbs0JqfONHncSB6Y6wVqKNFn46qgyrWEPJAXU+e+yoJESRRrUWZhk
T1CQj5NKqWf4qHUET9kaoUhuAFV5Ht3o5Rd5+CDbueFAED3hjXMNxxU6POyg9SR5
iS7uytdVPTWyPhXxk+2VZHEmvfaC3V+SMnEPxIzSmc4Fzf+tDpj9t+J4z9IfnlAC
hRlasehKUe2ywp6qraCu4IH88FUSRUrH50MF7LyXoTvsNS6e54mRpGpM443j7+fo
6vJzhhijH4sIoqq/QmbEAW9nocTMbsUcJktHKIENu1ya99XwssJBbcOOQTjWtwb/
+UhyGNU7TCmom2a0edTTDtpmD2j/Oa0Yxr1/o0/j+lpNFK7OQqUC39ndVqjy73Lq
lpbog+bFMRy0O7EBfWVUyp2Hf0T7+B/Zya1M/siTPpshtCL+aGaBPM5WRG4VypP2
UnFE+Bb67jF3awEo+cw3Wsg87LCb1n5OS5dns5SFdAPIjSGWXJa7DKwHW6lpSgJc
e53DKLB4dW72tsKHxEwHYqfRGfBFo+7RpMcYFvjdBUKJ7pZWm3rhEm4gwBMldfre
0iLIBWB0CCz9VKjD1hOaXC80Eri1+m9giq56qmepA99RwND4fGRCFElxa9CpHV2O
Htw2a1wB0qiuh7sKKg26D1GLwpNc6t6xsHRiYjIAWd2Ni0DNh0l/ZF4gJsTps8r2
A4K7MpnPcZkOwvPv9q/WzCIhY4r9eQr59Lgo3mYlIAg5rk+TUwQCoEbx4aqXwtmv
g21JQ2m5Y5c+AP64pR2ZZPxWPdELlvFVbuI9Fhr+9kEwu0LyBkPhZE/coWuWOkL+
lrtIV8AQbEOnMeA8v7a2Aoatn96ErAwDrndJEaZGV8uhu6VOUy23aZU5cunkcU+Q
bPpBR/f2x1VZMDYcx+0SZ0svzvOc1/0R5KRQBQNrsVEz1D+9txDqTiFzTbxab50s
UTSwyq6bjLdqlOYK0DB8Mw5wKrD+8mwtnNw/81Wwv7By63S5ZT6fhjiYdRfT4/jg
F8Z1yGWUhAxxxhSyP8GXwYTWrWDiWKMc722xumYheIs5QHoRV1KkMYdcVOLQgaCP
GoQ/Bjoeh9tPX3VFZ8BhKfZPbiUliWigPdD/tJr/NQ23R70ZlpMErXElralGO2X1
ximaWEDGkV9jyjW+ZfWo9j2XJC8WIh4BYqmcmKcnxx1hp53lTK8xpsh8acNUUOgp
Ciyy/kJIy4CUjBw0OmY6FvDFXLyQHZZaX0SbHKEsPPVf2YdQg+byeF14cXnOJO7X
2VxJdPeVIiiRzPKhgfyW5QC6Gon35mQjQzBID8oOfav/OpVBoixvm9fYDKq/td8U
jBFk7sNvsjj9F769KVnfgqsAquFKzknqUwYzYOBgvinY7k2FuApzB6F7LALA9tJp
k1k8CeDkakBgi50WuAWU4I/5A03Wvg+DSunNHaWy+lzsvK+fC4onYCoUGWVR2tEq
SMbmXSeZtr7cnxWn4JCN9xHEs7DCYTKofyHSafZl3xNvyC4lKJMHMZpkkpSZTuWt
smhWPavUpcWzhyKQH4wx5EwxMjAVTpfJHHKAubtJuahshkgdQih71kaRpmAKkU6B
tvT17j0jiS5EOC1F2MJJ+RpkzmULjxtEs3KvCgIWibq2shRuYSfdWmqjKHMoVzI1
rpdKsBgTpCIBXO9a/SL+Y4snk7GXK+iV/WpKoTD8Q6nVKCdYIYiOMwLr/WTDrUCK
HTE98D8VilfbgDJuWrZuBjp0SR1nrTAuwfeOOOCdNnZL6JrY8tY7K59fjQO1aSfA
MCDnDTNs4KoAbnAcwKL5CDqTKyu+APsv9CHPizUA5HlYnmLrjOklRXAnWoJvSrp7
pRfaTPhXzqkl8QZdNKubktxfM7Hhj05KBTpk1b3YOmYr8dX4ePMcBlUdCSMIuPEy
qn6wKVVRykvWXWzp6s5xgbPl2fi7XI3EFmf7uNMvoXFbDf7mGyhKtZeP5KDCx+Qt
Wh9EvhB/sdHlBfTQcxBhoM5lI3Qt5I6KGroEAHVhPRhWhNZ9G8m+CLEwZJ1wefGA
TOc6JgrALdjSrdeeNFDc2smwakJnmHb7FnlkBNfvuV0BWvsYEVtA4iDi1TJelaFX
2/C8ixYxSxuB8DNCesoS6nQ9l5MpzLdSct4xK3q0WzFT2x39qUwD762jQCLRug09
EfduNlChlIACvez2yIZe8IPnBNjXefdM6c0owm4YzOaB6rj5X80QfOu0MkXIGV+w
0dFthFxFVyt7rpZeFUzNulaTg1A3DHk4z4GhwssiI0u1MYungwGf2+MmfcdkIYFA
b2wyGTWj1d5JXfxcx+Te+rLabhG0C7A/4GnCfotv3Px1A0cmzl2vxyQGKVXoCMIN
pz6Z5GM9tzCRST0pJgldNmvHVpSSoVL4cBLk3fHlGFRwH8yTUhyXljielYtj9xdp
HSrJAi+jzx7egyTh9fK34Md/UqxBaVX6NgxXER1H1gwGTJH8C89tkErpIxuxg9Is
2473IRKq3aK81CI6pqY2vyFMCrGzyo48YYCEXINmdUzFUVdPOM6A68QNPph3M3iN
v2dxXad6YRNPGI3XFUfeQRfDADW8pNHbg4b7JTJYgdvJspzOoQf9yxmO5grEuekF
LRUYWep9a1J+jsfU6rCEs106MoTUDG6bX95nSfZwWgMKDesGdDiV02xxke9X05CD
2otGHfKnwzhhADnNZ/m3OEEUjLQWf80oc7Ml3BIuPbBtrWmRQcHdqZA3JopaYrZ/
AEqeDPzDqX8DFARRon3+Nktio9erXFHrh6+oNqzJPnt+q04Xr1xNz/eWE4Dni2vi
SmAuzRGCGS47UI5yr44/BzXW10lqfSbdgk2DiIr5aMzfwHsoVIUdqCSOfcKCso5w
Ttz09C5r9ksyXc/d9FD5y2pCHtdtt1RphJ4EdfcZT7O4PvKY4yK+7ySM7rTANvkr
wAQEXXGgwoxCEngsNOtWZ2IxMfYwQZuTwnAmBZ/miSwKMSUqqawnWHsGflaZGxGE
VZRN5LKkmgMM3WswAekEVxGFQlfzvEOMK48d7UChbqI5LchNCUohtI4LPqYHEsly
PebRkYTGvdKusezBwALxcZ82xlF+Kh3fqyVUnLivxiiQaOt74u1BWlnVmzghySyV
BjOQrC+VpckpnLGQGnhg3p0+PkzzJQ8BZaJTGU8Dw7WKvQAHljY4bsm6+FQmRm3k
7WRuebvm+Mx5ksfPl2iZkLPPLyT/jAYjK5nb9cxpmZJYGNeZyHFCMlc30Kta1PUA
CplPdIfUGK5stLrNS/nqFqYe6zlHql+pNI7xasLC/h688wpyGTVR4hpqvWTos1Fz
dyT8OoD3mQ3A+o8lQN4aiiLW9izv98WFE1gTE9hE9q3GTMmNBxCYB9vyNNl5QRp7
IbgVfzPnTDp6OREeWLMCnL+C5bb5VF3iY+piyjPIugmJNxElvp+6xGLPH7fzRRDx
RqhUSF1RzfPg2PqAs+bDwM+WBH4J2jDovsLDarq4ivEUasThqQExnguD27IPLzW0
a5ZVFU+Pl3ZaqbOc3EOjnMQaABQd79+qdWO/enBK3nvSJ/pivcn++S0X7BkqAqrD
8T+3cCH2Nrb/t/CcnqzeZWE18MIWZXJPK2HgGEHEauur+OoupwCYxIhy6rKf4J5p
UWeZbzono6p03oZmyQTRZZFvPePsJK6VLLr1/ryKoaGxuqeXPQU3MONfRQ6V1f4h
ROMGQPbYOXYEoUnFAR4Ng+SHZXFzZEAKDW9GHzOhpyXS1RpYiO7EzQpjsI4BW5KQ
dI3SCrGlZ6nsuYjRh11WI7hqHdRHOGwswzT69xoaax8K7E9mNtgWfjQrS4pUcEjj
lJATaQdpZu3CwCYxt5pnr/rzcQ/E/nG/IVoeP9BQJt0tzawQzbfkaXDCc9CUKNl6
VuxmVTKHEwZoOpldbqF/JL1PIuUkspGnjFl2WV/zw9VAjSCti0RovomTBWBi35/b
eCOw/+we0MbWfZ8ItMpjUS02Ubn14EKrjw9zEXcRP2fVl50jbcoru7MHBYmmqG48
lNrqJs3blEbdlUBl88GIWM/FOr+VoOUDeD2T4GJn+dtK63Diy/6MN0CTZnr7uRRw
iie/4uNbEq8D+jx/RWixVCs8lZ49LPvgnJyCoRmNReAWIzqO46g1UHWuF+ervt2j
xCRHwXPMOie8s2q1gUHJZ+yS7D+IJu/dziPnQ9xPYvopWvvAnmZEHdR6WVdE8tgY
dcnNu8ZP8IAwfQkwZJbEg2EN0gtCUlde5s1sTpsASvF5q1n/3BFPGLVd8C2lSwNS
bj0RH31Ed93bYbphCHYGIhh3UE1V5HRIC3NEx+WH5edTK+h37vNfS/13Ah7kJyHy
+jcmeQgJ3xOVnTYcrcrRxh2a0az4JrkgahkW3jW7JtgLgUs3A071mXSNmTstOLYT
0SsXQ9aobLj2LQqJ6IekmmrE7AiIQ84ejUsVkMhyEV4eHeg/oRxwiUgZi0hLAfWq
osJCVHndqbWMfxtzmCveErQrLtokRrGwnam/Sw9uxijbN4+7IoSgL7ZDXPvl++ed
hOK+2CcQ06YVphqfml68ZgxZ85fD0kapagIvIjWZ87l8vEW6LqwS7ZjYcjAcoNDx
FG4O1j+/NwsBBKUnLNzBorJAiAuLcKCJN9pulyaqpJPzo1kkTtkVLmMM6QLWmLIV
6ST//6miIPFmr2T+8/+Rv08fGBM/C+yRscXr6Ls5rdxJmoxqdNHR8Ha5zoa3jRNe
HSTnDHWhnYh+0VE0pbrZEgNk7K28shd8giCAHV4NezkJRT1zGrVCDCdr7701W703
HBAeYwkmDNmZJL1XoAVOhjCTLQGiuxVgAfH7l43arvG4FyOXmqvBdQD6apgNdMTG
/7NmqgYLTTiHRo7FNp18+aMHhsnLilre0FBcNQS3hwToCNpRNK1B3YYEkhgkqqA4
H1tIHT77zN0/9hvKJilyYCB1SBev81i+3/jHfHrgvJqVa1wNoQ4/0YIyK/i+f+tI
CMn/nLs/KVNvA2FfeL2scN1z3zLGO3ht6XEbepP0jK6uVZJI0agcnbzWVDhYL1Sf
4X9KIPSy+1r5LiadIV3wO5XBq1NbOkepgDdIyr57+kqRZKQftyuhwaWn5z/eLV5s
rFUg5MLtEG1R0llONfbjRDZMcNsXTV5vzbv7F2K/QE3q4A/u+HDqVHNmZmBQJUEr
nwwMjdkwMG8sdeCGdt3I+iAiGW+Q12VvOa7L7t43iptOPsDe8aU9sSQsfLih517s
RO2sZCOgSaDfTywn5mR9XGUTrIBsdP2z8gq7DBkmPYiPj3KYI1qSK4zHYInkd54y
QCCuEIxPK7Ud6hr63bf5uHCLEeEyxwhYmQOj2b1VdrxpX/DIdKiSpe7tSk/7z6V4
aWnjDIjOoZ2pbjLFOvM0MNDxAkce+CwR/op3+G/AxKYBiUaP37hTtKvkw/cbXz/7
M+N5W4BB2BAUfIQ/CyWRIh+9tQbMKy8QkKaiOvaX+YkkddBEC3gWCcGO2cpRmlM/
d36hk8tYeaKSbwpmLRe9v7udTVqQaTD0l4Mwen912OAVfeBTTpcPaQ/tqZdTw9u0
cUM2lfUKRpHKtJghf1c7qUksFzMdcooAEMn2AOCYSB5t/S8G7oftbB6brfrH09z4
Nfypv72+KxS2G5p+wZw6gKfDsrBfuEH5Nv5/CzhbAdz5cZcJQ5oPu3uUND6WdTFc
pSrIcnJuJyDS8aaoUz7RvX3ZFXzRSESAgEV/cvTu5Zux5KtGsWryjPG74wxj+WSa
LVfTbbwF4K5/2htroK+vbXHoykLTEd4uZss5ZA1pPGm2+N3nkJ81F0jw5rQ2AIiM
TtdijlKpZ31r6f+sUV3Z36S8iX7c3xwVr9ZkHfCtklhJsb/lb4xFmajxiGsm/57t
eVbX7iGf3IU9W4GW7cnRfzcYk8BamYadF07kLxUH8R9lbbXfN9nQhZqDatp+/zr3
vI+fe7NdREG0J6/V2Bm0WMFXLvF3I16TfqF2rues94H7mtBYMYp5aHxNCY35HRn0
oPQuHFC8kXDkZgCbjHFUUbIv1atLvqRIP0nIz4wdX5E3jCXtSCEPciP7fyfPNrWo
FNh1e0dlFqY1BA19E0Fx3W+y+3f68pFQSi0zt86oyeoRAQcNvB71w7dJL5I46HVz
4vkZMLsilkop17KP3C/vbL1LxtS8Pwqd1uNDLwUryofzIocuxsBWy5Igx6A+DFUL
nY0eesQR0dRGEgbN+pXZaJFfU86rqBYSYNo9+R/4EjYvyhTp8LFX/e2FaC9CUx8D
ombSKSwsmkJ9PMM0Z5c3igPGsYK5pop8WboVB3dAiFkmO13oL6jtSHj4UvUyFZ2y
2Yk7pume+qwm7Zfr5nrdLG2D/o7hG4a+n3WleyytgbTMCAqTw99znlKEhR2hML53
I+F8S96c65wq6Jd/TL/fIY2WjLtpcEbRNTbLrUy/5AnXmr8Q5Mw2BPr2zYocFErt
s2c52f5Qt29N+dWgx+HzwJrp0XRTyuwWLzSBBJUnC9aUuo8Li3WVFElNEJc+Z1hZ
3T/EtgmVpgLYxjgX/lxli7RFLD31g9LPlge98jiM5qlmIsUybzuAzZaXABxLMqyJ
KIHlK3863jU40C4r+Y9cWwKOKCy+3MD0D28MnbBiQzPNil8yb+/n0d12twA8R/0Q
ncITN1uPISGQPjxXeJ+zkFT6GNsvZcHn4fpEQLivPbOTysxPBZ9oyPiUFVqgC1mn
DUYbV5/wK1MQFIsOHip3AA1QmYJ4+zGl53MhSpATo6lmFk7w/MywhiwwBQKyEhvN
eFknp+IlWfsL+Fbv13mgoPX+kuu5flFY0zSnK+BB+LVlYtFstpnniwAxuWYxBKic
Cl0jgIjEERxV0NYUqXOkMuGO5pBfe8HR7K0x+6zMnSaLsQE/tj/dOVnJB0T21vS5
S7HkrfygO33KrRbdEp0z2Y6sT3nQ556+yjRb+uXiFYDSxc+h+/LMhf0MLmnp+XqR
Lhu2hJ4EraiTInq6pAgHuIJhLuhT1XAXHdiQMLnXZ6tVt5zEyeXTxGUF+0VPhxc8
5PtbYmeKZHpBmJfU+uaOZCeW/Yk+DVwWyhS+T/pDlf+OsGXMFri5X4OElkfJ67Pj
At5jisX2u5sxY8HYV/K6vG+DQLynXDRZBcAQUTEpOqrfBq8dZ69fEo45SqJykeaI
of25aqejHWf+HZ0j9EArC+giK7S7AHTyEnlTCEbfd3Dtj7Cl+NL8pagjTMcgOUXL
SEvfNs+P+UEtuDREHVxJ11OZ/cD3AnWSNpt99u7E4eQ1Ol2rnESG4/bzwci/W30X
viekqZK26S3XsyK44itlOF4y8dzp6Fufe5nYBmK54bC4NzkOfFeWKyK9TJqdo3fh
xEAaQOS9QLE926YbQruRezxDQmW9e3WeslRT4tPtt/5OLZNYYVxoLKV16VfJ7BXO
+lBJa1w+XGQNaHb9jYRZ6CVOI+r0BV1RS7/fNyjfyNzkjwmbSLSYL6JfMhogW2Nt
+mAcHlEQlOBVRBqG3jX8thKQYBn5MtuQjhzgB7+boUaSvAieTUKlQHPWRPMWqs2J
Pq8X4hZvzUNub4aWzyT5TlCrRkntH2ZLSPKdLXQzCQaa+EUavuXbJWnjiUp4VGgl
bPcU3R9zswS+D5MUl/l3e0LLF9dzWhdc3mC8Im7CP1BcPCWbwQzEocrDhG59jQRu
tEWsopJgG5P9gsPwGEx1RIgMXBTZLq70VDhx36EJEH3njGDl+nd/uJQ0LypBdovd
Y6CsChxNFBJsGln5WttZ2eam98mTCE75yf7/sFoDHukHcCKCVWvAU9iZQI4rNT+Y
/PVoTdOYN3xu3AD4T6KDJaj0PIJim9byzV3clJ28HACcLVTIyAEuAKGAKSjuWjBK
Lp6O5nJs8wAPvyYz4aCQECI1IL6x4NGpLElOpM28nGPzQETdR8NDBpF6U3mH1r9X
QGEG+dCz8D0rinFZB2a0uMoAYbUa68YcAk9jdxHw8FnP/t+uuklJUAmpnS95TlPf
vLuA1o2+wLoXdp02NicnWOmw/zQdDIy5W90farxiEiKSJJaF5nernAF96CUP/5FZ
7Fv4UQr13lDIG1DIJfKE7BaYAqC5W2Oaj+vJKm5/aOa5u3RN/Nkce0OfMJFnqf/t
vB+E1tEgSfyq8sCx1b63VZTc59pXAJisvfSppvjkB1NQsx3M6mSlqE7PcZJp6am/
A9is7I/XLYdVGa5m4v/FiJOk5KHjhJwvFfoi6+meT+Y1OLHs2mmhoQsIcxsXtwcY
9VkJhpwTnpqL0Df6eiO9Ytm7ngBeAWiWIL7MWYUuygxYNN8T9RO8QCfXzKZ3cAar
+xQLB5VYuwIS6ns1DsJZEffjQpo30/WSzYVLX1nk6oJE0u8l18Q3iNwbnS64X5fW
QgDHAiPCuxobyC85DMSQYv+OjQXlsvdKc2OW569AGwfT6FnL5OZqO4nYd/vejCFZ
eXsw0+svFr2JNpmXiycACtU6AVSPe+TFpDACCVUciAECATsSZtYjMhOv9L2LljGZ
FcA249gmPOwEsuKZs92lQUlrx8GP+2hy+B456NRBE5H1pWyKNVhsnG2CszMVXHOt
5oYZ3yoewbBEC1/n6feBJ+GPAY+4o7w2x0DmF9gmP93p/9T+jBJ/zwBlkJAJbfTW
+6F/h7cNJmmDTUTwD+LYG4bs3cNwV3oDYqcIIqXYRD/0ZtrgroEruSzDLLRXEvEE
HiUsFUYMVqf+Ftk0hKnWrk2ySAed4uxy4vZkaoza8PlCnW8ZFQD/0Dp3Vwg3qFrR
AtbTnYiHY2/HAPYGEt+KZbIn4kaUlsvPJAlKSWW7sCB0ZcKL4e8Hbpnz+PU1Dlli
r93iIgKczEzLPm0UoizVc5ojqLMp19LR31gAnLyCtFaaRv4ITdaicMohrTr8Cc+x
yUMGO8QFU6XVZs7LX7zI7cmvGWt8ZAS4tbKspLJfdwNvGzhVjHR8bxU/XWPBu0ad
rFQVHig/WiHR2T3LMXYKzj4RCuNWk/WvJJxWIeZ0gYDZSyflS06TSQawmQH+QgnE
1P1Fb8PIO8mVAF08mBSyAK80irb6IkcEg/9BfeJGRLb2kiuSFO4WY4R/GS1C8FGv
SVZkuz24deazjaxU8pV723GBnoj0A42Lwk3RmLkNGY3QbE/8/UiiZQMM5dfVh5Sn
fDfDgx3BA5wQFMBQ0sZ4DpoED6EqkHJ+ov0pPcUO1I9kRdh85ssGoaMFx6i3CwkB
xcz2upmyoZv+tACPMLJULjmu+BStxoVGcKgnu9NYj5C2D1tDXSgNzKWx5RGvcoAI
sHXAz3rQkwmbgAz5vnJAenNrVnz+QNzULp/TIpKTCwgfQTH5n9KAIkSj9convFgs
`protect END_PROTECTED
