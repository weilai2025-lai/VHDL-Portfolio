`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifZckHCk1784ekK4gD6kqS/8Y9jKpNg9nryww1fHP89mQT4d9xlh7N4tSktt3IdO
eJb0KmXmqgYp0bLGlOLDlmExiMkv/yqsxK0z9Uezh9Zicsk4lagtrUjeNXkdgwXB
p+M8DIoHG9IE+oc001jfzdl3Q6H5vp72/BGgf6sFjpfUyQBzf7gJ/VC79JwTBaAA
9tC2s/BZ3ozKI3TW0R6N4I9TY6JpJVDbhvrADQ1xZDkUjNg9F4KacPOzBnR8pqn0
dNFYo1EKDDSgC6rn4aU82K3pSip6opg3UV8XkzGVAYIO06N29ILLoJBZ0amjBeAa
VylKF+bcUC2u8gJKWMQ477a5ofCBH5uSeCoetRQ2fKAVh5Qa++yn+0vJW5MEot5I
zHwJECoucZmuRArYGjPYjrkisDF0ExXUm7m0WMeoDEXzGOr8sO/KnWInJj0U55XD
aPk6Cf38RwwDjPKNDk79Epni/HRlill0E8wQHtFK68QvSgCo/5C/hQr67nvaEQP9
9qX1QDt8jCcpSzsUx7BX1zii9vkXEf7gPuZofei5HEDYcnoHK9Oi3R9DoludvIg+
FBEk6+97UE4uou3+yh3sphIb4xOWJD5j9t/J8U+qtJPizTOhqnPNBdk5mV0pOM4S
+vRELWLXxVOoQ/k2OwrKZlCaVmU95cnkaXTHJPG5/HyqiTzD1EkIILevW6nQ4+m+
6DUDDwGQI3GhF5EsZGb/yp3jn6OTNPmy3Tzh42Bqr4PLkIb7wYu6eO5m6cDyHVeo
oFr2CLntXBqUu+qcjVvLmMxJ9vPOILJoOmclsOgKw3YUGdjLOC+fPs7aI2FVHe45
DYHsM9RALTnF4cf49rsBYJxuXaqnZlUdwb1bJKdD3NNuSYaScjd0tWfJyd4VeNbH
4OOJyUCYKt9DcbFfL4S0EJRXgxoeFiP9wIE4iC8hu5h35U8YLfOP0iairMNbJr7r
xEFmpV0LWD5tC6sPrvvixCupihibW/cN9Kbuv8u0sDwDm1gV8KmxzBBectXrMu1P
pZP5TRah8HEAg8r6pzN0i+YSwhbOis1Su5hB5HWLS3wIm1oRmeZUA+bYGOe7E/w+
Pxkl33FSHmzyy2RN1Sbz8l6eKwLDw16tjAzuTTtExzMyxVX2v2fRM1STmFkmyxrn
9kfJafDrwBC7GsefPvPjtGzcthh+1ge+9BLf/QUjQsIIpK1RkntA1BzXw4EteyxT
JDgDcBTyitVBEihQO74pK+3mRYiqyEi0FVHgU4J6Px4yVbv/hgaxC8/9ucA+bVE9
6SghV1GpqF6ErQdxoTh3XH4XLoLqi/usj36vmasc7kZuMJEbsBcYnVPtAIHtBf6u
OCZQeu1fhpbN4g8lalQxiAdLXtANCXoKg64oYyJ04+ZNmjeQxjeLDkLI36DQe4ET
paknfLCCY0bYPOTTY3ymGxMCRRe+IeLBdrZGLO6Hs448A4xqXCJeOxBbWxuGlI9h
7JdryKDLX2AiLl9E0Ik3ABcQjw+2A3t3btK2x+LDwCgM6SNUX5EX9tKXo6pRBrcu
mmiVtly7ZGtKtK0L1q4GmotSALffzozyvLgm0Mx691+CPwzjYDuzPRaHXv/JJMWL
XJrIcL5Qy4SMQyjdhvw7ER/jhMzo+rvVPVxon7dHk0hlrWg4zH7uZWeky9HTnEJu
BNl+iRQq9i1mxLMUZKs6JYMGqZyIXH1tMGF0mmoYgjZEqtPEMu8tZkiCAC2HtGbx
+CGLtDj6gQwjsczylAlJCYSZFg3mp59kSoORF+xx4sOL0D3z9EFujuIFmnaQwmKw
hnBOHyfNMrWIWVRRE2l97OM8HodwIJw0YBD4LvDhQ+pnj1n0pXPde+ragB7NLfDP
FLRxVUNEEtmzVUrt28toHJ6j9FT7QaoEroCiHuQtGupRwSgOAohCKeEFUHpWPOxW
Ib0+dXM8bPz9TaQqMK0LpWGiPEOHiNNKsL7eIiC688BfsCxqo7iq/SY+pdqM9sPC
n3dbmeayKSvDOB8CEK2iUbTyvDZMlpJX7C/wWygeNbjYS8sgW9ZmFDnCnceJbNsx
redqwykyvY0hXmE+uX3PK6NxLMs4qQGEuqb+QwPUBfd9Y3gXhozjsYXTLV+UZyRJ
XgCeHRUTdO6MMsngtUTm1Xq2Wtbmo/aCfBjrznBcO0BSywn+bTpFOzx+oZiI0SR3
WaDDvM7Q8Fds7k4eiR6Vfrn86pgsF6xdN8BBDJkUDcjoGuzcQush6VBSxzZNA4ZH
ws3RW1/mCV22GJb452F6sI00JQhu3+rHwTq+5Fa5vGgW7KAjZBonOltygDB703FX
cQGYXK0U6iYBNDhvnOjN+IqZZ/oa4C6sgDwacBp3AhpNCMqZnVr0c2SzfWVadYWJ
7+bNcNBvE6EElXu6P2gW3Z+y05fCKs2Z/WSnem4bWyQae18NGPxE7CGqFYrZCBle
ciD3IHiyn12MQmtGrHnX9qMrEzrcupye6y1cJwLy1CBECf+OB49LQgde9193HzWJ
IBCyXoSY9q5DVmCoEGYbLcqVvl0LyAPkIZ9pq88sEThBQoi/HdkgjpuIzqUoc6qT
vdrwgfBoAQhbSRGuZqbKUILJHoiwqRp6PiAsiwKidQO9huZ4xQLApSq1eMNmo//q
vnfSkOWxfKOWMWK8lMcAXZnczgsV7k+Wyc78U11BOjq+DpFVEHPO7Z6PyW2dz//M
4JwN2IsYeUBooQDld5YaecbPZ5pl5UhfQCSyhs+v7TvZvzmgRu4dy7RlWDzfMnx8
+iiAMLNgFMEyjjL/dX0l3in7eWQZ8YAbem8XoyO+A8+KL+JKwraEsJaUQ/4dVqzS
P+20KQxHRzuYgE+gJOj+k9qGv0uHxLKcd3aP1+w62xzBs1PZjMo8KOuXoWE/u4lp
XL71gWH1ofluULF7YTZCCsT340aXuDXlBWfUbVC9mszvuYY88Xp2ObDqPWNK6Sxg
EYR5O2PD6LDeCSLE1R/BL7DDg8oRMj/gd2gwSPbhLz4XdHmf19S67qxLaiRGTFJ6
kymWLG5tZd45XnYQ3sB3+b5MUBmxDUPP2MPvqpoSfy2YLnOmRPHK0qXfJ755dcH4
OswVxrIr2EBhxCq0ZsTftTQseXucWsgJRYifnyIZvR9qnxeoKwpXFB0tSmYxJtPD
THQxjbUrO9SeaQL635+Da1Yp7uf8ybWxGTYLnfKmUFSgr/ooNLLdLNW1eqLBa6/0
oeYKFQyqA0APBpFeJGtYTTEaeJzc/O433gW8CLl4z/Qy9H7GAVxuhJAdzHwvMfT7
68EFgd2YFX9meKCFkkH2cGX0OII4z6DWiEjWwN0hdetz0k/XefVWJEeE1h4wk+K1
FKmzKZE9b8GdXDSDHSnXT5VimOxNfhsvlQrAI0GLxChijdBH6mk1h62YwFghuIvG
+srC9s5Jni0tRaWPbCla4x7w7EUa/TGEB3R5S3VhVcxrCRjBQDTmQhNQfUYNhkeL
Z9PHp+lNMv5Krlt0aFbM5jt9ll/yDwS6rp8mXvCfhA/Wm2mT0H9xl4dcGqifaEER
uLCCkMENpYWH8LZGjko4MfnBPtPKDTQJTGOOTMqAZIRA2nTsGeDBoWVtxrCbs1ZB
AfsGUbL2UBfNC+q6MOrB0OksYLau5isnaql3Fnf7CM1RdhRmlKOJ6RGAhwgW4t4+
pfsBErjCV5pfy6gyBNd3sb9swdJOuzHj0H2a4rYSgX4RHu0ge+MVfZTuv6wlRZrX
ZipjxrD3d9+aio3+mSRZ4ht62DQL6e8QlKKgcGQh7zbxVroKwqAo1uslp2xI3+cr
LYNZq2+c2PeO1szy8rcLRF76x0+A50DKWB2deh28MdnkRwByiiVmrby4kC/gPZk8
NxyC36e0FI6uM89G5Pow0NvcCDUMKhlgIj1PRpOZWfg7l+50gOki7LekJ1ahtG2l
pFIiDjsTgWR/BTVkkuuoi5/BAtnLSyl6rSQOhjw3oFEIgG3Z3Los1QNLQUOzIn3B
9p9GFmDgdOZ86Txzqg8t4TLvb/9ce/cw9Fk60cXGmjb9WEKASqh/1KOsBORCZ37y
CmGs9OhJYAFjLNBZGGevKTCs/YGkBYxhFW/kXolg+6BzBRMVF6gqiKI1zn2jmXr1
4Xn9muqyEXIl6Nz1LPn1UkNSmjht7rID2Ki6gogCeuaxcglixy7q51mH2DoDPsWz
356ltHuKZwUYP7RX74Fto/4qn+AVpEg3o7c8ZCSdn8G0egyra8m35a/mVo9tcNOu
DRXsybEbfWzB4mbQBfNHGmDW1wJT+tnKb7NezGGIonUSehjYcmf6rn7vfl+vxhg4
z2YIkNWLCmczuDDeLXP+djbv9ELLOLrJOHCdKZIEXVuIkubNGzJxxkF4zfpIUpAE
5sOqXeOJrzygANJgSlwhFEx7IIZNEmFiUeQX9w/MrqgpKK2ZZOaVxGCFmAWBwNGj
Zs9e6rwr/nnPikkeqCJBbG1oSRQJ6/tLLDRd8Q2iKso0jlAdEOHTeiO1N20WYqxB
gbzKhUW3+v3ZYwpUuiJZ+0Ck5zONF4o3+MMglkyjNE5X24roC2poOJ+N8JYhtskz
Vp/C6pUkXKQjxe4oAEKJt3MvLXuZF6JKt8vz2UyE0MlRp02fPPahQv3+0YyxyqpV
tZVu0B4WgKAHvKedll/3PSJNuXsjb6BAhoApCbpBF1Er2coRV2hjC6unUDNzg3sN
6eRHHYzZFVVFvbhbeyldvVlFy98tLZ3Jf3G7NqMQUb/7LUjuGogC4FOKhYK7gtQC
Gut9BcFV9bp/59qMYvFvepbstOukuW8FVM+AGKHfreQdbYnMmAIxnqNF6S4jahaW
LFAEd/u8jR0uvZWCGTScz/cm5vcqlyM8FWCQqtYRJI1J5a4eAzsoNnSBa5V/4nIN
lgv0nCwBrygcPVhObv1BGFAW92iO4Eeo/CbHH5LSrn2Nr31YyNtUbgjdyfNfUvEh
HcDYJECV7XiGJnH6Jx5hDBwLKyYd2Wa0aA02AMMzUSD97Qaf6kJ2LRiYcRxPBGLc
Y8HxHuoRIlomxM8OYus1xy2/BFabXEcL7sMtiEU/8LwM/G76Y7iAjOQ5vhKTiWqd
XUENrG8yUsSSy3c6WmOoZhP/v5NJWmSh0Vj4ZUS2lzvYuY8RV+JikZUe1WZ9ShvP
dQN+jGP4sDZObSmxwXFZ7Gcxq7V4HPVCTq1VphjEzau8F4u1jBVJ2dtg3VKAJVYm
Ti4T52dS4pic1Vt+jLnduPDJ2CLnap8d0Db8Qxa0SUmDSfnK0o0HszGkLjjl8lPV
2GasMhd1y+2EIqUAOKW0FRYvQf/xhJzhymUsHE0LMmTyJMOeDRn/hYQUZDTH8Ljk
xwamcFKjySeg1pAc9fONP2MjaZv6gJliC/9RrKrARxmdIEgblGy9pkkPX5lK3qyP
Gyo3EfZKdnwrzYw8jGGmELz5APkO+DlzOJFT9p4HJerY0zrkO2QfC77Z0Z6p+22A
R73CtEWisZryr88nBYKnuZS1kodCp5fWonmab8S8k5Te/b0pGUG12td1DxJxpesk
ehRSZsDrcdN+1MNPQy8FvcVF7Nh1VGExeFfbrI/UW8isbi2Tg2NNyCujfDApklUh
qPQrqEcWCuOf3v/vg8v4iGhMD2CLubqsgZzmKMQKSO3RHsYvF1ypkauYbP25lqWZ
wrRNyX25g+yXtZ06uEvGjQ==
`protect END_PROTECTED
