`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFsAlulEkpZdcK7juJAXKvY2Nmx7IxFxN6Ta0r50GaEp/m92IYeOvfMKglOArAJQ
+uH2ghPXbq0sca+9J+Jb4fLAZklZVe/yaa5R/CX9JiDzUzHjuNCMLdZBY+QT3DbH
YhNNxC2Nm6OWVffqQQgzQd5eYPXwW+WTxh42USMnCTCXlTEYQjiu1Z8MItCXdNDo
0E3mdV95mbQvq5N5skFAE3E4JzSzpLkbK7J93K6Z7Q9eayBfH+0aOLWA2MR3xUmF
qQlMtLRdJ1Qck0YGUabaFHHa2Cgl8nzfAenRtzqtAklHKfHjXb9sKzsCIutjYH3N
3lkFCiOZoNEuexrIe0dR86oEgsNuMLpgRrp0aZkPqqgMrDYdE8Z9W9sqKNTE0wdk
pEde1/9DIA93hflQ6CehSLH8j3QL/+Zhj//bU8+e/7uzGMjV6UZBMyfLa+3seNJ/
y6Gt7rF9zor5J4p6IpErHQpUCzf28PSDJ8PlYl2lNys=
`protect END_PROTECTED
