`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dOuJyHW1gWxTDF8QlROw50iyV3I3DeOEQorHPQJdonX4FfHUv4eGS8vFdzb0HMY
piGhs/qpUQLsc6lOH8USgmD4j4rc9SEKud/TCPxrsclHG94KsLsegORmWSq0EY04
qF1Z8Qrl3r79OzAZk5PEFuwx3EJ4KThqCijBSo8nYxQhfvuJJqyCJobBAJ0/nlfl
pGLNQxmLkJEKC+wdMYJD/GnLMihvrYpcm1u+Turj6sHR4JvEF5KHF0eEtKCTTDsz
hwfIMfJg+aTk4jKqHBEo2Ql7s1dKwCDnlqll9qG3HwGaNdLfm/42xqrjZBicrmaO
LpODV9/V8c4lDJ9wNpUfqrnTrqFvoGHrHW08/oK7/0F2eAatuK2eAFfu+at6qIVc
YaTH4rMB+Yt6pYqI0fGe0FVp3PFuYvQzGKDYnwk1omnUs+zjDSB0dbdr+ai3/dPf
DBzljcxEaEKkpPmZq5g3MpFRgHZ8W1dpe3SB8QTtYIk/sCGD/wR+5GRm9QkTYSZh
EyYjUgp6cG+effhIoO8J2BwvZL6OYYkJ0xiiCxLpuJlWjUk4fdf3z0IudJUY45ne
lLm5+j26p/ya8/V7OErw0ky+kprWYRrKZ17/8tNJzbc0uFCYz/5B6wMC1sAYFx2H
57aFi/O2O4grrbFVg/i1O3z8mjPAPeCgglJjEGxssANviDOLyEXUIMUuA7POeq1X
OCn0C3DAQAJL/OABr5XqqMntieGqYrg5SP9aK76muXfKVAmt/3X1k+ferOlG6YrM
v04I0YDiEzrj60lVI4xS9GokJXOLN9TeiKdBJfoUSKG02YiqIMN3zbBuKLJnahxO
AhvmoTz1sElyjilfTAZ7SkchGBe194P9DXejQNkOoAxjfINtq+LkuDn6X5h0JpXH
Wo37mCJumM8J6cXsNSM5Hyv8K5oH44fKsRyY38TtGirrqTwAnajZNIij8I0JzaW4
S1770FHjBfdYWPc3ruzGFyRThaJZuQqCNXJ9qBFhAunWS6mWBdaZpv5J6jeNHL63
shxI0+T7Hu7enNr4RRXSBPnthcvTIycv4otCvGRyirdZh2FFf3APbaFazeHjxFAW
7gqB//C6SgIT1sxp0iuFnyKAOjruImdZ8c5yJSYTFP2IX4/M7oEjtqAAbK4XAE2o
LGaD+GL/AKpNvJGpReGpSgjN5ufG61wRn4QT87khgi5unq5FP6W/+yZJqb5wQeQ6
/SYdAJ3qEhqv7dUR+OhYczqTsTasfxds6klp875qGHMsNXkemlktIKGUC83XvgWz
fDEtFA+grb3y5KhiUADc7ME3tBPrPzYRawDL/961hZ++CTRXnGYsSOesyq+C+O8z
ICulE1CbLbXF/BjqwXdeFcgABWISmO5+Mcg2N6NC3LNu6s42TE3wwCRMU97//Im7
eM3MrkxD1O0ZaPjk2BL/e+vdJO8PXbosWoEkiNuUzIxOWvJ0ytCZCOzk0jh6vhGt
WfGWBuWDn2kJJJV74dq+pom1V69CEbzkVg1pRiUD0CVnb9UbKf7FkfLvJ/y4FuWS
QCVIjcV2oYl6fAqu4YVA5oqJigCx+t92Mqxvab8Cib9k6n3HjZ70GG3J8OU41vaD
zimi2GWGzCoblrga/De+k2yCI03JMx3OZgDb6RuspSd7yLcVbw8BrfKuNulJwatl
75wzcmu41UDEpn5FBJhkdePJ04ukqhxIpIw6Arz9er47LT4OwI4GXBopUpLlp2iD
ZPrkDid3ze+iuJBgFBrVNWEkFhELP6Kj58cjRDhGu+RgeRD+DcSiFEBk8GIIAaJO
G5CNtVzlWuv3aGKObNsHjrhMiLUAvJ013xdrfaKGzTQA6sxEpFBAnzQQVLGHNJbT
dQTvQp7LfAq4Cn8V0HUj5RfPS5/xIkrASVnPAYJQPxlCRUDi0qjV6X+TzkVlXGHW
XggVagkAlhft6WPAE5wqYA==
`protect END_PROTECTED
