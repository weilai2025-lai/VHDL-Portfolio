`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMv7arHcETid4rCJRS6Z+uHcdqw/rND3Y/6chEjvCjm3xiraIPFL7E553yJtBLqO
TwSuqOZ6d7Pe0PnlEWA8mnuSmtHp6eticVMoFgRlNdrzVa4yIlX3aJE6jl1ovNdJ
D25x71M84kKm5CAjdyLzxhbd2SfPcZ0goRFqvtmiybDpb9bGclDzGnVBEi6sUtXh
FP0l3EDaALHF9CEfr4dgR4+JqckV5g47tQAAa3d2trk8yyFmJpUH0805ppGRe93f
NxBL6a36UqCRwA3O6+ImEJ9h1HR/2qzQOOffdYxua2h6Zok3TAbUa0eiXFXI4ZbQ
k/w+kEWNj79mnAoxARrB7V6ZOkjY1JiRTGQipy0XbMO7PTrlWCBa6ESfKpfdhofc
8iNfqnw2c2Ko0TJ0ZnJX68/GZdOhW3Zn5+aiGd4Nnh98TzQcapJ0uSxJOsxLeNGF
FKZDglzRuUEptvJD7cSa2ieuyYKvqiSi1icZU931XNIbYAM+DgAibNfrQCkiN0NL
NT7gEH/6Ie/LibpLyMHogWI/DqhZ5EXReEY17OGfzRUzDalitA8Pjq26p81weqCG
x2EKpad/0jNB3GHFu6S0N8rkXWJlFq/yHrTv1dPz4Ca/s2Ko749QhAAltb9CcP8z
PiqPN7jXgDeKMTLSEx66xRQacYgoU5++pfSFpBnOFp9Magw9oszwThsvBbJ2hqXX
Y9xqQmY6IZIEt8Rl3XW1zdBrl+NLPXuPWTSaYiqAYgUODTC1ZmI9cmD896XATQ5X
o6YxFB15cz3AjWGG8hFPplGtTBEW7snzBGmjF6Z0pk37msgL9/1b9jGak5E0n4yQ
fRKcmQNZ2QDyXdABw6R5Ec7PhOsSgccIalL5NUYeUdhZ2gdb667xh5IprA/3/fkX
2gIaamRIVArbIHef6Vf+kZ4lIwhd2ZhZxzD61EGfOXm7bP6l0laMPJbR/BrMOJn4
lQNDWszLUPsHrjkz8lwyW3qXZ2svulRoMEQeynz4bhhPMroiZBIVahw8z2qZMypp
ypM787VknIqaF/G+L3H0RCCMSLRdO3bPtQrrhOpU1E3lKzc1z46yHD43xzSBco4e
OpGpZ8rYdEbxuYUb9PCR4pKUpcHaC6lBYqlwuVGZhO4fibk/ZtqbzBsIcBZGSdRR
oLGtrtvVWFDgVdrVwPR7D72gXDQVh9QRs7yFJO83WTl3pPDlKxwAP9Mb/3+Lgw/K
Ts1kDJBGOgT6AJz3rLc+1vJf7/Vwp6ChWAFOnoNiq6+z5VF/MYDusFNlO6pe/Jgd
MD5lOqrUAzRe7Mo/WupDoo+KntoKAdjv+we/vEjfw+t2GM27Rcvuzb1QI3vQyGdT
xlMiQZlr3xucooLM9G+TTykwM5Bnb1qUPOdi6slJFJpzsZ/oqGiFULo9jJTIdsNP
ZGtkD9Cqbu/zupWP08WkvPNxOXvKFrhkBMq2X5t9hYPPJ3d/a03+BgDX07hwT5ak
JYo6ykQgnv6NP0QofNYn116OsEnIl3pktfE/eYJ916I88hx3RGZNjPUuQuHUxOw7
lEMxag07sjF9+IotoFSkzFuo2o7sZdt5nELY6uLvtVT/r4gRmQ+ToqCiyTBx9u80
EDg0d8+vcY2GY54NFr9HW9O1WT4w865zVEqZrPaeobwE4azKwFOXHZXnYYOIMiZi
vfreh2totJZh71ya+lEI2leb1LvgnV8KNl22CjBFreuxJz50TUC7F6S6OEBGbopS
r7oWV6GQswBz12mUKHrHKMSIKe9YIxYOaHcWU4NQkOxDmi9wyqrfzfuXaGdT8Zai
nBosaHadUFegzft1o196BWU2k9CTzty0+AaTUlTnf+io7alw1XOAlQ96KOrkzQca
N4wKCaWcYJX07kSnDXc3JZNMM86asA21i228K3j9r5pzwv9jIJMmX4W0sBjGeKJI
fWb1mA4ZrZ4KymFELI3WuvYn7tEsLaotnmjIirYOlR3eTLilZ2WtU1P0iNV280qK
Fyx+97ktJ4mg6+TkTBB4G+zFeGQsmpbaeDjNUP/eqheqM9BfV+PC4uyLDzY8M9PE
zyJrJFo+TAx2f3tD6PnS4DsX9b87BW9GK6+Pvrcs3f3Mu7XE7HrwlYizwKr36rKx
LAJh0ImFwEnUlKqC6jy98oMpl9lTZPCDITTA8H6mhl85w2kEPYdEXEEcAiqhKqaP
n0Mo6qbN4K6Xwsi6byqp4Y73RfMZEc58OBJvW3VSIS4CZZ1Omw6hAjYHoVDSOIHD
8NBdg4pUGWvF7L9Y2balT/8nvIohUZ3L10Uhn9dRkWhrifvo2MujovGTGTzONGIv
yM8EhZYu7z27QqLQihYwwV6De7qnGlUjJfIWDNpSJEsc+Wta7qkoykyUeb842qZ8
SbC24b9kZJmjjHonF8fYZQ==
`protect END_PROTECTED
