`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jpNqmMKtKAnwlYYh6LWX267t1K4amb9i/B20Kp/bjmvpw3mRz/MKE2QpIr34n/f
74OaE4GovSDA3S+SunC0AIDPPkkF19Uonb9KWn3u2+fFJrx7c2Vcq687MTflgmTY
D2Xv7Xdi5Wbv6sO8zpsQWJG3BMr1GuzOZ7jJiWZz4cLkJWanCR9hTThpyFbffNe8
fXkh6a+eUXvdVRurq1gU6qJIDNsvmDuDiqo5dgxSS5KQ24BfBe509b0yE//6AJG/
nguHHAtLZqJxr3fD7IGbu3V8aDFr03QUg3Fy6cr4gC6tsiix7zvKFndFvL6/md6M
1poTpnhh7wdDPVrbn1ErOx3o4gmQ5kSK7CQHsKBG76loR4l+zxAYpazG11RZu9qe
+gfU0exmD336jndHuf7y5xJ+LJnV5rlnpwtikEH4J5HcYHesVZwKUyQJt7T0+POp
vebcgLgxA1t25svXhX8buH2QcsMFUm1xcxbCrLpUuxoJGCT1yIeP8YMtIg3Ee612
84JLgp9SmR3sFjMXgXvHZbXQm0wcEKA7VoY7Jmcz+ljwU4zgxLD84Gevr+RMT/A+
rDlYvhm6onv43HK7J/GsxBV+EkAPpN7RQRPdcWKpFO5Of7M71yxprzB7ggHFwogT
ac7SrlXfDmk9uiw+7LmqDvPOilhFLFT+pPayqwEIH/38R1IdBWqiBp4XED3GRyi7
SQvJ0LmStHOlM9R8D9cPR/UaxKQ0xbkKiw12E6JYcUYLM05MeiEZJSVGQo9T7mk/
eunmK2i/u+cjX/nRvtok5+N0oSXEBXresIq8iNvSRChPJAxIaQzgn3IwPQjDNL1N
kTWEIo82mqqNDqh1AGai4vleE7LUr++LTarWwOt0I82pj51Ijx0CNMWYG+rtBPKa
LrPeh0Qq3QZzSAU291mKd8zEjcenkyYsq4Jz+KaJNHizjVnzpGC5wtR464ROmHjf
dDMn3L73G+ho4JufkGsIezt8wpcVkrsuIYNn0eoyZiazXUZZo98UBbNmwKguD39s
/4e8BgLQOsEZWElStMtdUgYTzaJN/X6lOIR6yjMbDcTi947RVICSwT0NWoxvHeGK
PtGDlwyXQiojxBCypn9hXauWcNIMJhxZ9yZ/OeMZLSsmnoYVwQwcFxa6faR9fgiQ
R2zknvPV5qn9kXFZQgzTJY44ka41MUfYm5c1wctxJpUfI9p4URC+KsWrnlTYfogA
6mxjQfQiX/SbNFrDodr1/+gM+N4Zj7aMELjqlI3eAfA6npl6F3Pr48wZ2CEv8M33
JpOmkRHWan73VPltpkLK4V7Z7Muo6Qyv6efPHfBFWmfrPkXDoLup+efeNe6kBoVN
neqQTW6E1m/yAG7Q9rD/Tv6F4Y/PKIg8tIMnp5wHW2NXPeDDC8Ikcf0ZXXnCtq6t
erZaa4Fuy3G0qGk7QLkr++/imVdaPa92v3yNVR+J38JYVaOZi2P9xObM48mexVH4
TMVoTSnTmdclFrJ2c4HeZ1emDbos/glBOB88yM9ZdkAngh5SQ7QdDzOZ3j50wErl
ekXr6tA8MDuQKoz/jD+lrwegm2tEXTFQqD8XGqZug+Yp7LkUTjF7bS6SATm5x439
rAWHab9VjCPNMvh4mVOgAODTJqQCW8qW09OMrij22cnfvwbCxsbOL3s2tqPeKAYm
G1RMO0ycwaiYDMb418xQgDwwprQieaQWHSrCfsZULbbPbbg+U/8DHl4Hrb7GZJU5
gOcOeRdqFSvretD8txxfz2hgn9BVyygJG9F7jDhwpZ73VOVasV2obS/1AsagcN9d
bQ6sP2joqu1LuC+MUwq1k4DtxcfiHxZC71nHU6OmmeVKVRWNRutSP7/RqfYXOeSN
afBoHBQMqts5SEoewv1aV0iTYw6J8uGe/C0DyxlgycLPRywocyIpNPZkclEimpHh
argfWTAeAQl4fMQGv+HVmKgDZ7QtD17crouiHCIa3oDB1mgoVJv31GmpZVuYzb4/
WJS2Lw0Yl49y+JUAY88zbF5JIju8f5KgmuejSf9qivQMNcquayTRkyNcwicDw9zp
wQf9NHozdqon7abcGWZ9Cm9IXdZNgdh9QQvezqmK6JkUrj5fS2iW8VKeGwOntrK9
q4OX4Mpf+oOdZaL4eN6GSyAX7LViEBHkGEsYp2I411CBqX87pSw73TeEjWCWvhOq
JaL77c3iYuqVuFs5OcG6ont21ZbeLl4gb90bUnWX3KgPqFVD+kq7km8Z7bR+sR5g
pbfUaMgrEImnQGOsnuy1u6yDR/TFr1PqTvzSCUbsKeAJlCuwQ3694KozBbw6z4QH
/pDCE+fdE/w8P967QALq5hx4QdMpzgiT1b7OJHW9CsBxSj2Jl5xSvT1tld5dKTsn
Bu+7UeGDM7JTpSmtSGRJpEpvgHl5K1DNEPOYqYWnxdG0SZQv0TDIJUfkderua2z2
`protect END_PROTECTED
