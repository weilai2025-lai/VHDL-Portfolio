`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csh289FwrDHxawT5ishr3Z8ulLd5+Aw0h6tqEhXJ6ohLZZsawdhtFDFmozLJMLGv
ZCQ4c3ck/ZOz7pH4w4K9xfn3bK7RtymsXO6KQSkI9rlAiOSihsPigtpxjdrmc5iC
PBHUkksCwoAROvI2cPSSK4BItx1Df5/qmXYK+eDoFyG/88yaWxwQ0jm5ViurYy9T
gLs/waVY69/nn9jR4vapwG8Cl472bfF2BXbK7ZGqaXfbgRuh+RqC26e3GnqcZo1C
30/+fHjeyoKb2/x4gD5r0t+Lu7pQjN6+EjSfaq4yZdLB5ipMVCTmx1OKjNby4re3
77oAgzeNyipwyqZXUOjOlwwKuTprgfTYfICMg5iLcztPDs2o3GS6wHBUhaJE5JpK
`protect END_PROTECTED
