`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vOLRhV2xgl/OIvfTEiR6JeBNVrDF6h1amPBXLbfQfab2+/OEjQMJcgdNYxQ3nZk
D4qKy3H/LgVFYPQKToiIP+cizboJfSG6FH0OFxJEuRW9vrLenXqp5HG2NxUZzOcg
aLAKPUjRiQ9gnVgdyd4pekkWGpMLWuRjXcICXm68w6Uqp1eVoL2+eDTL46AR1Co5
l8dRLOzjeFhTHVoI4EAp5m7a0AhcxWh1dQn/lXLZ2Mw+relQqp1NWh/tr+DqfHjX
sDnhFqySOE4CIK/pewrcLY92e8vEFrcYBs8n91zIParvJn+zdwBSGS2i9tjBNM4Y
chrXvql26k1knnMd4kGNxTZRbhlRTPTIjI36/CaP8KyyQZnOqr9zP9PVbJvVM8PH
0nVTWmu/AOH6iF32MZxD82Gy+aleEimKIfARj5dEsmfmLEh9gpGH0VGjnhmX83Tx
fuaJrg/eyQLpbk2af3PVfy1T1wW2RvlGZn487GNqZKW+WAIhA6oPFvwscNyQZEn4
eiE2FkhP+bl0eF6PsFh2MSpeSDcSvn3tTbp/MwtiuZxYs70NuKspyA7LeuSDwSRW
H1YaUbrBvAAf8AwKpzKO/Dth47oxPXRXxRsjgveA4O2yfpZ6eikfOR/Ps6WY/tmm
vUAvKkqIjT1kXYL0jFKR8NbywmcLtS6amDEI1AAcJX0oOAiHsbi+MzVbc6+9O/4Q
GVWRqeFXpEqLlXz+3WrGZO86ADPuGFENaDz8gvBdIdiDErCJN5kVVac1UyqmFQh0
R17cr0gZAa8ypeg7s8J+GmAr+n1enGPaVYeLN1cY7CsCtAkFkIHxDm7vPInqwgZ+
ZV9lZEORc35n/X3kr8ykxUQnL4vc2rZM42nsBX8TTe4jCixA0IN5c8ZSwVlS+5Rb
W4FWzlbmWehN3xmu2/FfB/GZ6lR7Qa+OAchl7CJu+9Vff7EAg71uljaXVEBLzZAA
te9+Rxq9suZoRd1kA+fGxpAsZa0F1Fu+iC3JqEIoZGxDXmUfSVrkMolkwHn/qHn8
x4R+csqPRjgKorrB4p5pSvYAT1jKaauo42i48xUOyMB1pAnRUPVNY+/OkWvGO5ia
yXc1uB+pGs8GuX3OIX7QY8LgffkImoKm4RwSI8EqxqIArTzhRzNs1PmhTqOe9GPW
A/GwhOEwQIvzHWectAcELzx8+x5QIPN126azAeJu1NrpQ11D6ZKMIka+bo66fKXB
ZIa/uqRMDBZJU9WuLV+YDs9kJVt7+kyqIRk+rqY1+I/6WM5PJ9GXGJEMe2HECRtP
PQNqqp5+oWDFIEWywwJszXaxX351m/xmF83HdeKunwbX7yBWHp7rw0wuYsgFKAWU
uP+yvq9GMgVPoqTGwk4P+zSnSyol1jzi0m8poyH4xgP+XSUFdlT3dRCUPlSdgXzj
dl8F0fb2oIXCgQJJ76bVGCzG6LMcIke79npJ6Ibo3bmdrzpU8ypMXBAlhNqFlv/5
4akc6ryF1FlPJghXQ8XRAadJO59xjKupqO8u9s0Y2tmjIi4Fz6Rco8nrm/yp//u5
FR6An2LPY6jjw8dvrac4hlmQYFcxOcXZOkGfi6UwDCMBiuNnH9CBAd1SqSmeH6Ep
EVxCVOoBTLp2KDiSOJOnftlQzTNr31o/fTjttJ4q/IE33iDJMdliRg0IkyLoscKO
70Cb6NELevmEzLCXxz8BgZszipWB5q5kzPXB3sfzZ1Af48kBy4gFRN7n2hnrwHk1
Ik5J/k9beVkOTSY4SLByYR1uW/qrGzcvt4V0pCblYg6gZ8OH3IKgSqeGuLT1Q9P+
9FGEvf1m5x4YZkKm/mnVEZ8YtGUhcCe1sS4J45f+03ORAI+5yKXlvmZ4U2z9llFE
KuWOu8I3XYcbgGfAFE2/Y9KL4kp6F0d6nQOyvb9IYFX58LxE35G0dgv/Np9+4Pdl
8oiSXB1uIklg3nZuixGlmKZuNWHcOoj8Th3QWqdmPybouvdgJZOHSnEvO7qtnknP
V4HdhGF6xabqhUwYk/VogVf7+F51tHvOTm3Wre5PvFImqmjkwGHtAI8sJHvGJ1Jh
drgTKrLJSsrPZ+PWdbIHkZe/2dPl89j6oJ9lW/Vgfnm8Ve2MCT8v9zuJ1IOiRz9t
hnx025qHFbV+IZuqSLevkpuFUt5JtaeBA9DMtVPIzTsqDjbud7zJDTSDIWb4DlO8
DJPRj0LSqveCZ3YNXsFgpRhzmLOwd3ZnXp4qIDloqldaP/hUoraS1tLkMlGnIaVx
t76uE3HBbd/j0QhVb/aMDQG09og/VsPaHIpbg+5MQZJi7TXCzzxs8jX0dzpx2v7V
Y74a4sQ+vYwV8rz25TKLhc1nZ1/X/z5QMQVwHpVLGCWWL+yRWt0A3x+edm4FmCKd
85jbHHIVzlPByrqcYgWxzSYvFPIgHc1uASn7qa2BnRXbueM1xFqd/nof4yN9YCmL
ilW5Xx0TyIlgQCbn//nr/zbdV07Y2WdIFCnIBpf0lEy2siOGjvtIq8wIvuzotsJ8
6GOBRxANVwi9E+KQr67QdH3P9xs/h1dOAuvtWv55ufxM8KKlNv2O6NG4NJJ8bnSP
DT/Tsq6f2tOm4+nypiqskBT75aPJO9r5P/lwGcUDoImQp+V7h7wzRnu2uLm2h/GM
elH2cOQGTqzw5wwvXnxywoBUDkpmQSmQAsa6C3JnaL1YJoclmMwY16BQoFyzL5Gc
CUoWcw4TiR7hByfhQRWZDmdAmhbI7actTR51WJUCLOXVMpGnrtoVGwVq/Xv5UmJ+
xuN+FNqo7uomj3pDYMRHqYmiXUh53E0hm2mW1pAw66hrZCACeHCnalouq5fW48qk
sPf9YGviyTVw623utNF1N5K1n1JTxVyH9Z3KxFVcGdgKUgNAVeac4sqlJ8S+z088
chme8VxGfEVO4tGh5Jy2r2PkAq8oEoLFrX+sd3DG8lBaWEUYRz8EhNQOh7JUfAg2
saCl/KC+njPZW4P1VXwcQL1e5/mjAt2gk7XD3s4N0t+h0lnUKbQdTAJXg6dZD6n6
U93C0p3Q7RV+r6IuBNWKVsTQTSwtEkrecrOcfpXFmafXCtrGytP1fREJIaQNo0a1
uzVv7AhCKbyYrohza+9FqVTYNRefKARJtfEbkwXsxvr9SgmlOmxqxGSF/ctBFpVo
M/eJYTpvtneM+J/JHwBrozYrSA/9lnWAMeo4tLJvoEQkOdNIb1Oj1hvxwfxnCiUc
0d2LMdCdDPs7HtQ70OxpN3YyavbZcYIKtMrKY3Ujf/6JCk4H8HLiWSm77Zo9iDJG
IQkYZ1fxJHH4LYGUQ4SlpbxMdzCC1+PYzLrZmLO9LGHg+iAM1zzQemOPVKgyhmti
TyOQBrldHIfGsxQ7mQ8Xih3MO0XaHzHvaEbx9Cxmzxs8APqQrBzbmOYabTO0CZec
NKFL1c87a57JKsR5hj6lmTI/4Ydl6pEeRkKNHVWvU3y/wd8VOkdwDbj74oANNBUQ
xrTO93KsPnxC5pACxWrGRTNsBDff2UQzsF/FEwkuBRapnJClU0x5UbiN/ZBp8ZkC
suc/EgtOilELvoSs9V/8GAGxxHHMk2d97mKvueHaCgUJ3DYVZrpyFNLk8UeS0Dpi
zDhfmSZ5audjT8f+tOIUJwZMD/BSN8xnZiUAaIoUp4jQrjSop+3ZwmlFAw3TTJbz
mSgs3rdY2fe+SAQDkenrULQTO3log2iMMOZOeAi3/F0aujM3lcdyZgWUph2i6/zx
X/Kquz4D+SyU45n744tufIjAnjpR7tDQZDCZz+5/tdyOBVrvwRQPZiZPuJMovByX
iE50RoqHk6AHprxPl2pw8+OWSuDRLIseEhFqRf7QR1qpSSwHS2/YfTocAb+CRw6L
D/5nlY6pZKs5duwcMYhCBuPUpC0bsbFHVL9W7zmxQo8K2WIbSMyEK3Yf9Q/Iuc2A
ZdIYoJyqYi+6s6VwTpqp5D2jjeM4g+LBYi5r8juNXs+HN3KWSJz9gaSBSjrtYXcG
8ZdztwigMFHPqfNDYeC+y8HVFYacb+I4Ti3Lfo+etLiVFYbwFV+0IO3VKx5EQN1/
568lmhEcdSXRMVWKZtDxOo1+s/u26nyI9AU9QwxldNi3SUjIEGRnlMUaJiiL4jh8
ODR9pVxPunGmtvq+t4zVt3f2QOsSy5eUjAGuJjGVF8wiTbJy2CPDLyWpcCh4lhZi
h0bFV2Z0HarW0lnThDoNY6/DCgOd3ORoBGcPDiJl+mzFGdK18QIg3W+4yLoR2//m
`protect END_PROTECTED
