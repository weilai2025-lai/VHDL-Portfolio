`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rsAfhnMOjCX9VCkDXr73XtJmL0i7QyutHvptPugBHjgNrwalEqRG4IEAHYhHK0ec
TzFfGlIPnFUeJCF956+gUPLhBwGrkbP0UuiE0IzWnm1n0f7UvwcbHWvTOWss9ob3
8GaLCyOjagW/vW2dJ4nkE8pL8aOrm7/taXsPayLtPN3gT+3YhHF1Y5loqSDQLyxl
memN8TxDuzt3sJkK1/a7brShv017mAbPztzepzKJj3uj5WR2ivLoqvBucu1ETHNQ
WL041YhmSmZacl2B/R0oerw9xtgxm3Jw1orizNHpfppNxtd+9SgpEF3vIq7kJycE
1pktyCgzIfbYI53FMeu5cnKxS7mLl2t2qgQPRsPUXge6nwjrIAj8VgIyQurSXgM9
jRw6zVg9KgFrECk+XAt4fwnHRUYYKFSQtV1Pe/1fEih209m6oGLfvfdY/Q4BHHru
YGnwBZONesgXMJbZ+t481jiJ7+9lvirZVBcdcKJLmMgd7apo7ZQyNsz6XLVmL1gV
sx+E1vTa34BPV1cFWEuGeGrFlDcpVpq0Ba8eE1swBVPOAMW4kljL1Me7ppGZgKf4
gVryOFG58/+7MYRKMFBn13ePyNmE5FBxqgOabZKuW8Mjm8s008P+B3+XmXTMMvh3
MshPbHnZLQ6xQw+E6MHudKw/1XbwhY+3UtZcZJQHfsltDHZXnEX8X3u4VEzZ1J9Q
xSEOsZ6Oz5DCwzznN2gKbLPt+HuqTEnJJ8d0ZyoWewtRQhtunWqp+axAcAdBk/ac
qORYqKmr3MX+avT0zU+9Rit8E5bC+XhPjGSa+hr6Lg+19tI0MHPrb889UtspIFjo
yjrY+nSoIwR2wCxbKoanfmzASaZRnlKAPWg69lqJxIYKMhP2GE9X9/IxJfaFslyB
XnhuLMEj+FHR4eMlWHJzlSQzpl96Bre21j0XKaX6K+EFCitHu+hXycsAax35jgr7
8WVnghLi5+OHvkLzQEIO5fJbtOsGtR2Jqk/d/o45XjRltYX/UFr0BZ4RR7NYgL+Y
0nPHWCcKSWJmyyLVSdz/CjOTv5eoe9UI0kLeBOcUVuPQc6tW0CAOKKKbMFR+zgJD
QTgvgPzo4uj/eGrCxTOkxhMw6zM1LxY8rawyaZBNf2shC0B8nxpCqIVBTf7YQvgK
S/IvLDKZiKpP6+09JLwUUJdHcJ+QR2scSUjkviPy5iRjLLEzLU0M6GLsxaBUONbY
HTbVC/y2VNGAgfKpE1yFtLg7lkdccLfymhGUB1jFvglLvsqwzKYCf4qhlDiYrqRM
Bq8a2AW9NyzyDQGFjxk74pLM6KV+uE7kjOgWKoEKNnwOfIwupAj4lzhF2iY/Rnz9
9fOKPprMqkV8Qfxw5rhzDNuROuSS+6adUTU0YnGVuObSp0uGHFm6ATTqyvJrsy50
tyrmNr+aoxSxZ0NfxWWn5z0mtzEUzKyLcJfYOB7/MfaW981a35Zm6yVRAStvh0/e
V4mvw7sdQI3KT28d5ytx1guFY/5N+U3kqmLNpa1m+sEeBp+IyfN/O4qucrYToIj7
R3S3fLOT43lQIlxjhYKxoVv+KtJjHWf4hGtijfhk/jakAU9T2m2gyHtHXB1yCcOo
/cnl24pluguaIqhD2B/kymqSG38ELYOK+Ea2HsGaf72dwRcZYbbZKaeSxuodZjI+
OJWueq517WQP3kdY3mAaGmT+iD2SfWM2qt20/Nh3+DssJAiUJtWuTDFJpSdH4IM7
DDetmAPMbtdgtrXNh6EpQYwJ9jeUWZCx98BI5vnGo+q+6uo7UNB5pjkYTon8nkmU
vQskCjXvrcH7enkPE0mWqS6NbJuwvG2QS3BevackgeutIM6dSRSlxwPlcQyniv8f
CQVT+cxgIaBvJ6yGuk+9GuMa7++eQ8QnkO061UxpZwKUL+wfZvP/dTIyPXhL1+f+
JHf5LGUwNSjvNjlYOjo0K7IzvTXE0+3pkKOszH7ecZRL6V7YU+BYO7ks7ZQmY8F5
V4pxwsVbhQc9Klm0owVJ+RE5t3yklglLhnxu/WUtkTWv3Lq4y4fZeemVTRLbPn22
fTYCRFnz6GEA2Fso269I07qfpNbBa82fjzl1sd9JCTIKkgm8F6eeAT23hb/3ynb6
Pg3CiBmmzyi7PWw5YJYSHXJe3Ew32VSmiIyFBKlCIpMg6ewA5n9z1NydmXKD8R51
D+WQE2aGE9TMbsdYfZ2wEFMBcRIl3T0Kah800iNMfMB8t/yKku/+HgWmqiyAQSzC
s5BJ/T5evrjUVeV7E3+A037Ua/aq3wfV2hYhggmjzloTgP2MnOFiHjrAyyScyi1+
x/o7iBm+HTYjOJY9fI893zIm0Cgcb0EVRKjP7V3hyt4IkgEDfDk8jo3t1irT/LMC
FZnBNkzoMXPZqtmfC2Iscxe3jlAfaOnOhmEYyD2jvMZIMQRlbABl1+WucGNtsH8o
911MMDpCcQ1LoaQIP62unkfdZjAIeVv4ls2lVoFoLSttTWu0NDHDjY5h8lwv5Cid
OVwbqjff7Krl1/GvB8gXlIwjb3FX8Yw/OWde9BkQJCuBOVB13+NTxJ8NfiDmv5t2
gtxgr3QCYHpo+UczUJU8DySrBe9vnlDdMUhIH/sY3bQ=
`protect END_PROTECTED
