`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHPdIDD0CNqtc7skAL70P+HxDIiglwVHuI+i747kE5HI5zOJvLEkRVwUt/SXAqVD
t/s8T+jzUrwPfZm1dXiQ/49w8JvL1aYq9tUxzEWapd7R31IZs2Wp9iosNKtQopmj
rfwdE6anISl9xxDKHHITTyZcTQsX2Sc+5QJFNq7pO7U4nGgxTuLo46E27I2AZ2+m
Kxc7r5Bfctzj11IlAEM2j+DcqpkfrmJOSq9kmod6IPTbFifaHQtSq3U5ERM6YlS2
JmqmVsm8K676dbVq+ZoXtVolsQnV+sKRZq8nlEFobQv8K5z3gt8kh0bT/elMMmE/
cEFMtPFJ7uGNp/0e8bHyIZsFUIZ0e5Ge+E4kfeH3kyKR/VOfwTdlnatvFwMre5S8
r+pqJ+adGLFykaH8eV3cqafU6Qjiyh0FMgnkJ2lZ9Hi90886odN3KtNY9HGTANoG
USmL/pVTsoJjR3JOwF1KxaXkkTPaiYMxkeoc1ORYoe4CJYJl4v7j5Ub+4z1yARiZ
VpREAugBnp/oS4rCHbtHI9xH+ptoaG3res2FghumicMm+Wy31YgN2CEvPR7FxlVe
9/Rdnc35857EoL5Kp3FORyTNTw0TQsTh7swX72NHVGJgdD3O7Avb0kLF94p77vSn
KHB/AHpYyjA7pdWYRZjdVJoSkeRUdAbn/g43plkGTd+o5Z9tHqqgzzVau87ziSHA
L9nb9tx7RW/gT8WmW5uMchc4uuioXQ+3t6qAgxHiq+3ClL5BeAvto0vYgl63FcOJ
CVfJWwnOsfpwfThIbo/YiV9dflc5x20M2gfZWX1RYQQt8XAEVtWEiIUHtXiYVmn/
E6LYoNiVZoB7IUU5SBIZC6Z6lGraCFPalr838HBTFhYDUjaKGdHv6UgLW36d5vgi
8eo+nMIgr+SPBmJuOSHJBH+nbe2QVYIvp1bkhh69O9ppnWIUNR7nR6fQGJstJdOm
ayYTbS5gRnriT5tWr0IzIVzk65fNopISKNiZVTPY/2YOE1GLaFy9AvgKTjaTXHeE
4yY1W79uRSr5ivEq6VJtZg0Tg9nAlmHY9ePtwca0O3ntuMVD6RL+pWtKH8s2kekt
2fgbIwIjH2tyU66J7d1vdRFFU1iYkFFqHhT5L5ACdXVqdGITpPmNumaahwXjBbcu
xW0HOrAwwlN3sBmbv70I3E8Hngk0wNLR/wM0hqaP2dE37QLIRYfUuXbTotGUkRnu
iGxiewZH/0OnfWX8fiAsaD2Vn+48LqToYlmlMhMNUfI=
`protect END_PROTECTED
