`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N6duhOfosZGb41cSr5tqQuIehvIDLUDWxy7G1/m86jHWlX2q9i5LgMaThwaI+hOD
DLw44mcHF49cUcSqL3RKs2Oc4J18Gef46+NBkxS3hD+saddiSusQFWLdzs1G5Onz
614a/G3EvsSanVN/QVDmSteeU5RxervyD7lb3Koh4pr3xCDwyjIAJh/8ublRHEDS
9WWx2pqp50c/LvZdqw3q9QMSU9gEOA2SozQwNohgycNU81Pdu8LUIOjK5wig8Cbn
PHICp5FIrq47mxT7s74ELYAuUR3tS6Qxi8yTvS/db0tJeAP0H9XWkYIHML7mOJBm
1LM17TWqkOCeyltvw1XUdjQwOICr6X9p6d+Vo/DeBEQjqSFMVvMkLLL8bdQajazV
Cn9/c5Pc/IHW9xzbY1OKBQaEE75GDTws3XJIF7+ZngYpgrF6j0MRM2FOBuJj/zEm
tnItgoR/y9hj6Q7Eo2sCwTVtitsfsc8rPN1Z4ipszFlxX7MwRgyrMst5r+X4vylj
EXm7hoGog2zwKyKWhveg7z/dP7ghfCUF3keTx+B/fK/3O92a8vTvEr7EGBuU7BXw
GPpgIE2jHprSbEPLgwECYE+uMCdriYHEETze99idz4fhzwX3I5Zu9pC86xpRXr8H
W7SqGzY1EnbQWqF4OGE6ZwB7d2NwZHBZEkp4g3O/p59J/nqklXIeRGEPjEpXfk5V
S7mZpENJzrgdHBsN/Y6BJqtN8EuUHbUklyyAMVnl1h/YTm1MC/ZOjlHoPElebLAA
nIPWqn4Ux0c4ypf3NRF+YiPWQATa5oJCEjDJVV8/LXowBUwiVnVMl2ay+q+2c3wt
irKS9760r6/qZ8da2ved4NJ/fk1T4ELZl2v1iGZ1Y89vkRnWpRoq4LQEmAcMCr7q
0TPAhTDOt6WlaYauvBDg69Qh8Tp3PZn6u31Rf/3cNltTlXfsq8/TH2uX3E/0q7pb
TtuMYNzOH9IKFckYiShUIjuHwS2PpEU9KMwQervdDTwwq79K8SP8nlKztWu/YyyI
TneJu9sqmuVHIJ6jrvGoQQ0JYY/HFmpkQ6oxaD2g36PnzgHg4+3NrCCyOasgtSu4
rujAKLscqxCh7rc5RalV0wVni2LQWkbKJPD8snRLDDLVG19/pygeI02v7g9+YLyA
2mhclgs21eXFc/y7gHhrIun5nSaNg8yTnbC9sUOSbX1Y16iHbZMEllwTJ2MXt7LM
v3GsybTwBPgWEEjP3YBRISo81FOBr2RRaNsjMnvCudIDJcCn1EwzbiPm18mfQMku
HO4IwAUUy/7QtdMTyRBl46s2RYA8ARbpDTouAnuQRFYQ3V0Na+70egcDt5qfrB8z
PT8Em5DB0abmJjxOx2tosxtVb/8jROWoSKOsDUeXa7le0h1NilbUCs0OkxeP7Vo3
hszJYjQgBjkczYPxZCmJvYkBxmd7SR0taMhdedOdJezRSmJU9ZAls4FTbcKh0P2d
13LMfD8ikZwYAzIzmSTRoWd2xwFrbc9Ms67lCFfmVGJIWD5WocoiK5fKsQQrmjFS
aIwQ/Z4D0l51jXTtv6Ov9e0iYlNn1O+UCC6YV4QVkguHERlFGPLRCfBMUHDqRBa2
qDQkqQFLaOA9tABTmFb0oBoDIakIZRsXwkchG1n7nj8JefB0rqIvIVlyFil8lX1P
fjyE+laHj7Ff+Cngph4yOzQmfgL7zRinqMHUA/PCi6PBKKVgDHKvC4Kv5WJ70eQU
zBNzKZjbTNlFiBcu1ChcIry5tPbfymy5YiDSbl6ic86pmoDhoGQnE8jy8y+FNi98
/++JTeRQ0GImOf2hkUJ6uNXFmxrHrxbVMJPWIdJkY11dR75pSPp0TR26TNjOTSFu
95xkxOp0ygVUaYELzJWOjersi5RODPPtaWZ+P7V2OOCkjZry+zfieWYXWhbeuvHJ
qZ5fcG0HwEl46qiX+hGQ22GAWzVvrFslZbljZwAxJa06uPvnptLzBIivT7mfoTGv
mGY8ywyWn5o70RUEg0UetUxipkX9i3HJGQ/mOcb3M7m5tmsB1qQTBpxDDQGjwiFr
bbmQKYxRbERUNJptca0oAxxb/NfmEbp66sh3fgHQsP/8w1X/VvIZ+URvX2ckxkFb
voOn803l/ZQc0ODLwIF7+5S0wHdmKU6I8bxx0L5hVSuL9gLKFvvAYTcGGACyaocF
5sI0WRNx6ED7JiXj/EZ+v2CcJQzBGq0VFWSLe8mTwLU=
`protect END_PROTECTED
