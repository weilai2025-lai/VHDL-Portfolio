`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l646OyV8h66ZUZao5OkrL/hrXaajhMjYN64kk65PT05QMEgH1q4UmivTvNFYAHiB
sCFxcuOsbRZnj6ZKFcgJlR5eMibxlSwuSrZJJvtKlif2ua5xVFm0l6066rmVdiUS
4cu/jkCi8Qx0ZE47EDYPXH/CYQI8jH1XOfOb3V5ChcunAneJQ+DczTT7W6O6dkQe
X0UaYyovq+M5OqzlftS0atxqTdj20DJl+LzKjA3n7TL/GAWGkSho3LMPA7IFC7wW
fvkoYJ1yOLZ5fvw3ayWAHAFB7VvVV3F3fQgHzlknRItvmKnHOeDVi8G4gTFH1E9+
2pBcMHW6ZAYCdZUC1ufKnSuC/nI3lajCZFs3GeRliY7fLc2O828JHzmcPOK5MKKV
KzxvJr91zTohRwFJvYcW3Wr+RIK2I/3Lf0ZeruzvwrvjU0sQ1zxdWXbf2FfM9KJU
4oRXG5d8V9+iL56vmHaBGNeEqXWYBNBiSgFc4EWG68DUJmgUufsGhAYb6WLREjoF
qrYLkMJLeNrFgd2DXJUs05Y+yBIzs+wQ47j+3OiW60MfSPGzHONVLGGQ/yzsut4G
JlgRZdNa/HN2eUeIbMbNoYvrcPV9HH0ipcTYewIP1Do68z+nfP6WAPC/mmNrHvHh
24YY31GRPcxQ/sZQjzqDYP/gxFW4F3BEmpjR7igtSPtrawe/AdClvcIbLzwj4M2Q
rIYV5qovcg5kEE8KPNKgVRkzuREnWGiG6LAKNxqfmHKX6PqfoU4n59zboXBC0klZ
n2cCU/H7w8NAYnLPyzzEgF1eINJJhk5C3dL375oYrx5omh5z4IgVie9IVdy5LK0t
gaTsEnAYQ6noFoMnJe+eXw==
`protect END_PROTECTED
