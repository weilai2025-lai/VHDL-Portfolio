`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mLEDs6MpItWI6/jvrisTee/tefRRtS3Q9Yq7CEH4Bb2ID0eLWMAN0TgLGYHu8LF
nuyIt4bYARetNmzuDrPq70/tlnjZRO6c+nzOpYJgfrZ83kNaIk5J6kCL6iYF6DWE
a7rslb7yARKEKRoFwQ9P3DQTpFD9xQierNX+0IGg8+pFKTKKTDq0h+3Nt5ffB7cp
/SJgMZrAa2ecr/WaUwP7LCcbqTlzZ5J9BDvMWQ/s7n2BOSG+GJgO8z/JnBqx2nX/
STwc8xQR+GaEwbMNoPxnHgDzHM036shNYlNPUnv6Kw4wSEZftrLhjIQOFUuHsawi
pkyOqHWnO8NcbV/Z3luiuXh7po0kfqF8PZPQgFch8it4uKVZ+5dptrlws2vBa6rE
kAgBxEzXKY7frjlqrj3mZ1SahLY6LEFpQVTkRsLPwFkspuoakPEXfpguK+kDgE5K
HHLL2vcQcj6h1SJ51gB60Q30PpJ616Uqr4zRIn0Lv6M13b59oUct9lg+uoPbg0Sb
Tkaz8emKwy5jtnQ4cqWkEJ7q0DtwS50KHZyvB2gMgLXDmCnPab4put2er4fKTtW8
iGsnygV/glojcAiK9bQPnLoDmZugmrtUyT4t/nVg80moXzyJRUVk6HuT4CKIhPGV
ewFg8AWiGVm6dB+fJWlob7k3lGoZB0GXXgyvY3VGlLoXqZyS5Wr0B1z9DZ4dGvgT
SGgHna88qeqvhYqTwlizr++R8RkbSZq890WLvn/HhPu6QnBf4iwp3gb22uTxhMpJ
D2/zH24KpfeoICk/Z649t8GhqCksKN2nvE1zErZI7QQNzqgH4Y7/ciiQ+0LUet9H
+RDoNQG7+00n2thyz5aoWTXnglf/iY2NYMRTCi/2Yzw=
`protect END_PROTECTED
