`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5BcZnrhIXyS8s3+4VObwZ2bomm9kqRCc/GM57uYIbrdT5/Ij/6N/eVeBzT0oxF8
qCVkfS318aQp0kT5KK9WjT1wzrnii+g5Q/zFykD8dLiZRoqsuTfN4O4FEkT6qZBq
kbW9xPA4yNoiYiHwLvQNAdMHpXzj/b7eYADtgfJrT/0JheJMs0YHI7EfRYMwq51V
iT81CeBmecH6dBKUh/BN3qBIqiblcrY/HNeR0v9Fkt2KGuPq0RpwyiLfSbQ4oVVJ
kmNVMz9GJxBZ9GHBrXHe7+5oCEvKcR4kS21d/oO1NjieTDaFYcfZnppW06g1X1MJ
DcHeo5GI7qdEGJwjDuv491Cf4pJb5Mim5QVqTl53HTXMCC9tDXqqsUvPd6wJvOSQ
8vdKYCLAYlIkA8QuNavonTBIcAjJvsDUpYEfq2BMOt4b7d3PTarxvdgGUfl5KZ4Y
3ZVizOqwnEfOw+ppFmeTO8i4NDB5B2Z1UJP2TPFdUIGcuAyITE6w4w8lA7fsyUQ/
WDZ7ynP9zEJft3p5kZdNKo2OgjC9QmSCldPfdz6vu+RmCUNlCBd3TJHl4bARgq+c
vssecIxki+41A40O5Y1NM/O00bU00I9rQAdZNZpOKSo=
`protect END_PROTECTED
