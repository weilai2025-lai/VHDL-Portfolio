`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cC735x3RIZnTW2Iq5ZyhDUuKwZ6h4DRmroNBwjwlMeR9V0AMdkQwI54qxEYSyG3i
Qwq8ayct2JdkZeHcEm9uAqZBWxQLlmue9KJwutn0/ENGY9HfoeEHpD2pEPlEZIQW
5Q3w9OSpK+eruRef1mLwCUU2130iAyem6ueQ/g04On3dl5Rq2HNjPK35ph+/eW2y
nQqo8aNmvqzp+9QRfoW1K30reNcvmWStB2qixX7hHEVxSAn/1/Il6aspuRvO3gKR
0wYPnzRJhIvBiNf7eKxgIfCALugL0phj6FAOuJ7uB0KENg+1EPDctsOTal5UDtoU
nxIrTf79zurIaf7Jq2xqSRO37Fsm+BEIk3isbbf4foNbGARCI2fhjojFSVRs2WJb
E4HHZbw9Z3BQCH8DVNB9I7YV8B35K9zwp6tiCI4GDZF6Zb80CSJL68indQrz6Zp7
+ewBMR11CT485DApOrS5ujGbE4wj9TUjDYaSESggiFUi8kWhwSxLiow7WRa5KNi2
dTnmHiwGUcB+KWpTIbiFB/Ibk8M08E3pf2ZCdTC17RQiCErKAhFQaZmMa2yJLU23
jOWxXBpW2TBrZ43ywrL6Bx1qHjfdU5ot61XXFR9H7K9ZT/jjY2K9wPp8RVHQuWoT
kAgYKflCBzW1sJkW1MpcZfK+PTuZ9OGlkx5DodTfIZBHUafYi2zS/iiVY0DN2cFK
qc0fssw8kCNCupGGMLRT6Ux2BspycjqC2nagBsJZoAWpOrjvGt12j6iZgWqzNv9S
O4LrzfHRGdD+aCyabqQExOf/G9Ccofc2SuTKumJSlenx02D3hMvluEYyTMfacjNQ
IkBglPEZBOdNY3LQrEvjp2rXd8FPbu/1Qb4qtaDPmQ5d0+0H3teBeWOVLrlej1oa
GubxmckdTRBnwrqnx0fdScE0a67zOO5fZrLjFTtlCJ7N1eRgzwqmJD6czHWrkhq2
hpx7cuj4TAUVfGzGsI3IqdlBJh//qgYoHCE2HV07GfknqibZ0psJB/v4aekW2VTB
5LVePpTVuVnLnWww6iFxV922N3BBJN2KF3SEvDMjv+Yu/C9aSCvNSW2V7hUlo3hz
XX4XG+LbQCkrtbCmrSnkwr/8vsrd7fyPC/R95euGt8KNkTj3c3ZrpuvTCu5V4x6N
K7M3OZFxP/Yi/unXs3IdKVonL/UCePEjJepf+Nl+qpLTmCNQzce19/Pc6/mIxQkY
Ok00GNySyLdKAQbDXjeaieZEKQdFqLdKvlwKVG3HxxZUoGvQrg5n9ZDhbrtA5De8
xqI6wwrD62a8MjyEFytUNPrv2QuumXxDLfRByubPyoF9y0d0RJBJUK1+0ZRmEBG2
YS3IE1hpyvG/kzzc0+5RI9p4g1QDn5E0nc/F2XVZ/kMgx019qdx1zshKpupp5SQQ
p+oH1SLW/kur8aOq1PDCWxOpo4ZdC6VfvbbxlHW2/izXle6Jtcj9IicVnbZvDYCe
d2hDaQT/AUjrVPHLG4Xy1ngKxMeei8Z6pO4TVd7zFb44hEI2KVs+jl/6izhoBcvg
fYFH/uegg5Dm+fTLs/nrkGtk7VS8LJu286DKbEiIHtqccpyH2Cl1UvAXt0zr2hy+
8fxJx/d6O4mDSORh05C1TGZMlgRTS+1BLJsiZmJYJGi9lpnMnkZH/OlVOAzM9WH0
3ZER+W5k2nNLVD64+Y+9lvvsnvdj3Ogup9djGjuT6h2vMeyPCHQhe9oTBVi2I6PX
lt3yFJtezP+G3t/85b88TobvftyZNBifvqjuhA0PUjJUW+KKG8bbouLbzdg6nlJW
VBHot/ZKl9BRKY4sd0tcZrfpBZ/+CUmHdiL06Wx0NiDWMqAftl35xFrkteIOyRUn
gRgokHgY4nxny4Ej1/Zt1h+IXDS3fWzuVBWFWdcAifGsz46Orb+erezqP0QPR/7M
A7y4jKwA7jA4wT1EXZYGIQ9gju03UjX+0ghdfHbN90dZEfHgYwdIjjujY4QOUzz7
26RMGjwfSEFEYnFfxfnsE43DJkPsHHFIMaf61b+MWPFH4H5vo3r3soVqDlyiEDMe
3Fm2Ut9XLL0RTxo5bzJyJXsqMoLf75VZrCkiYpVeq1jMLt95lQ6kQ0ug6NNTF827
vm2c/45AdcZ0Bwg4YmRZBIk4efsUmTNXPYT9yUt3pdAl8t48inyG993ZZ/modAy3
lGGDKfY/iHCHWNfMh3sVg1IzCCqKe7eDiI5fFteOpM/tMgaDglH6tJangiv4w3KF
s7CLg9u8ixQmsmjVN9yAaDEDVvWHDKNB/JOjhsvH3lVHcZap8UOQx6OHza/hBCku
sila8YKY3B6HhB97kM++G4IexYANIXuo5tnpoEELSnDT5/m8NkXS9QDi40NX0Ko0
HpgbQ4o3DqW+5RvVBuvmIiiQewStmpnltY/9XsbEU3fnub01AvV/RPrVNLy/8waw
wW6XxUlTos6Sb2xGTCuluJAgTwtY6Q3P3aC0EqouYRNa6OaiN9h0EaHZMKjG14sT
Nj51u6rPDj+CGfbuuKoWU8wxtvcncTJjnfHWINDNDIBvoxjsO56TLielF0Wad85U
/4Pe2HeJnutsyzSkpXoGHDWG6McTm7n22WaTY9CE7UkDRXc/e1cTYQZa9aKMjF8j
BZHLAOUte5ag4T0Fs4sw3V3V+R0c+bFDnbY01nk6Cpe5PwBDWW1Vv2NSrWo6rDXU
G/ZOlNE0/sv1j+PvqhlKqRVd4Vcvcf2vbcHRQ9hqWv0HfzTO6koyeSfssQod+lHN
6GsAT8VVU6iMFyYW2ihSifkl+uzJjaj/B9ju5qi7haKOhmnN/Zc7HyLa78PMTbRH
la9Vnp+mFhE4ieS2HxJgPdXfElxTP9SpMa7XpRftTM/wuE8fYXPLDSX12tMdc0A/
OIxZWWonLQ9Igw2jE0Q6aeJNllyMa/k5Th592UGA4dI7yzn+CVp0g93eRAwUeAse
aR2DDXKcnNN62y7U/ioN3i22/yDqfG+86kOqKyu1VYjMx2t4X4jSdLemQcEhTogQ
z9xURd8kbbB6Hq/q8VP2X+abmJb+rxIbLl3mnDv1HKwAF9vb7hh/EIHMbMLKwb4c
ijrQWJr2LNzGRMBqhhN7r6Ew29REGIUKP+XGSljTcIRxcg5noDzmm69U9cJMOOgu
idjqY6UlU/lya2QGmUoN5DLOJKyQ7DSscqVeHQ32r8wZKRhe+WbYKKYy3FU5cgLi
9l+zuEH3zrWXE0aOoL0wMkQmhgggmqVZE+qTghoYu8TdNumbanzOywzeV2am+KZa
gCul5j4cx1KEYS85DB0n+FpmnW92j4Sa7I+HuhDw31LpkvXP/pZFWJDSx1QXu4dx
t7mTT+jtIp2Tfwhq/qfLECKW0rKq2uRCZIusaoxiP3sb59MBWLTsTcgvzrOQnWKy
s6kIghsePZgz5ttsoU2qoEdr7hHX/XVRawPNa+pKML4G4Xt4u6BPkiXYWAZ3rv8c
mvorDYMb9VWo1ZGKUUDY/XxCXBFWEcIcetjYeaFsrJx5lgyxvx/39o4FOMwLXB3L
wi6mU+XjfxroWvaGA4FRRhTiXoxUyPB3KIhlP1yHyO/D2iocoyKrMsV27tNBLHZG
OVVyBtEN2jRxVEIMNQHf1TFCxikN82ShNAsV+n49tSh8IebWnXIXRibZ0ASJ1mbl
PSU87l/WfXp1SRWj/1D19S3NFMtR8F9W5S/2sRdS2/ciC4A+c/B8J7Oj8lGTvHcX
n92BkudJmPNbIEJXzOnJmLhBK7uflgE4WEaqzhmLlWna9nXdRHeMgGs4Iccl9HPl
RzdhNnuNqwN0b+q12rtnssjOglWYUQqNAi9bPHwqMfUlKv3nLyJ4hDlo+fO+gVS7
NeJH4Z1cLaUtZArrllwhRcw4Ai+zDmjIYHi5pQsEgUtmM064ruFCeo4FM9as7zOE
43h2CGqS2FURaqUfLKbcOUKai56v4hG4nGxM0zPenL3oPaafDgtC1Hr0MwCd7m+X
ElJHD+dMBTvTNNOE1omIDmtWodvjA9sdLCqmcH+0OdkD+rA4c8slafFggST0z+rL
bEsP9QiJmoOAPqNIoqpI3wHRjHCQ6uWlk7rEo8kimjM7XW4QKq0gjrMhyD/lLrGL
RVnw1sSPcNYTUSdTgIJgfA6bVEn1DupvcwEN0XkBX6DJdnIjIvIQpUoLwgmSz3dX
2z8rBsoKtCr+d90vYewRfRJevrVVbNnitY6Szvf8JmEteJluS/2Rxk83CJLjNXE1
qay5fhdRHgVmdkXF4KEf9rTdoaGMacpRVZdPvtzrqgxeOSb0AiKdhBmdgRBLSH9A
X4VvMpKO5RfDuvmd/p8/4fji0xh+Jr4CvzuExQvtBn1O1YVecuGZJPYu5UjCDgU0
S6L7bzzbeYh9KMHRt1MizCScqysG/gXViWtMx06n+k8Jrp22Moqmsv2EnoxxxXlM
c7tgT6Okh3velLlWTaoyfhXbdeSserm2YCySgEDvGiArTRa3Y3s9NYpiPbKHrqOC
YOxvEyiVyGjyEe2nEiTyC2CPRuiEVf7/n75p7l6LIZEFVH/iBNdam24JNjGy/gUN
I2eCWaropLIfMPN3tnls5xJm4jpcRZsX7Dn8HWw5AVfYzC0NhPfzNJ94BXymNjM8
8cgc7TaQVrSlVDLwyOH/W4GE1+saucPZbFr2alCdNy6Yq60SE7gWb6ASj1x2/Eli
RPmbHVrQu7nHt3vN26Yl7YdU886FXCSWjnT+lRjOZsytTOHKxVu3AV5S5iE8D4H8
Pa7XDI36ZGMAvWeJrlm/IcbUl/BH/pynxp70ThqQ9i/Yp9kmvAW+YcZXUTsse8s5
/KODBLc1jtgoDpJQbYIjOEtb21PF3Gg9PEs13+AALdUp0kBzZ5Mgz3DOy56Qrhhb
kz6w/okOc9pO0KGmL/Bt2vUr9Cxbp+basCGTMSMc5OIyHBXGFCKxVMve7j8xbDpj
n3jDCA0HBG8+gHguTi+uxfLVvHDwhDEY9pXwK3DPz0GixRKDORDPCSpD3ebuErlO
C/FmsIKf1kGGwj+dPKS9oRFvhdLsR9AJ5/ZyjMWmNXeppnXc+unzx/Dj1lRvQ2AT
w+V2sqkbAnYsWARf5bia/AHq5K7AeQpZTvZrj72iI6l9uUnuDEEARJx9tC5SP8gx
sjV3QqOpVMwmZfUqlpk2dMK+1kIl1yhcBlnH/XX2NmL3otxX3wMe8EHZAKbMwNjc
Qrt4iL+Za7y3J/wAUDiLJZg8jH4XK1f0+71+sxP+no7SNWuwbC9Fh54G3ON4IXbO
fFpcTjH6mF5EU2Atg5hJaP98tDLION/e9FuFmw9LmRuhdxcjiat1pk+fqPigdfxx
ZF/soZnLqEUzTkdo/ksArlaKbT1bDihG8/aBpSbXGr5ezGxNw8KlRui7IQX2WwRL
H91uEKB31hJ1Yvrf+Aky3w/TSFHA+JMN28jV5g0oDFBGcHJ2l2a/Ey27ygruHhzz
nt12HLAxxF3j1MQlG7nE6o2eMIpsC5XXIJCiSxl1E7mgmSlFo4+nkMScZR4+Y74A
3OrxO8iycwoHuRQiTU/2Tavq0wkh+gxVWCtc0jt9JR8Dh3orWWWbMs4Uo5y63MK1
lJ/rbKcUardOatEl9p+eBzcIVCjsxt2Bs/JbudjUYVR5JlRILksBCvQSI4r+JqdN
rnLevTIW3tM9yqGl9bmgJ2vLtfhEJkVF/GgzuFS5Afd9Pxj9/GHTzdmzZTEnAssQ
MSMR1w4jlpWh8AnvTiDpHsA76x6glNu8Uq22q59bhjiv377UTwTYmb9No7E8mTQn
yzlq/RR+telfFYFVCx7v0SdtGM/RiW0g2Eiy7Cmi1BEODTpNywDxHlpThuT+1NxZ
OlDFALWNBjSR901XtEgd3iOyWIfhqkQYRvVbLDbFcHj3jbWKMDAmWFybKJ7vn2IV
hDzb77TAC6cgAuUOPPHmzoD989dvQ3yZerNe8kvFAy3UWAN3IFw/zP6ZueHufkma
CJr4sabRoru8Id91SZMluSRY3W4ba0UqCNkD9cI7P20z17biaWchlwJ6CNR6Hjaq
nSVpJyXYCo+pl+Yl/jRpghN3aEO+CW6jNozeb1dKtxaBD0m7BrZ8kaS/95cMEFfc
Z64wLsMrSrgn6YKp+zAuNcsO6pba2EKM+QzDyxLEuseBd4Yq4tNCl3DR+BZ9Msu3
AYBuThXRdB7Y/g3tD/1QQZiwtHqjoSTeKM7dpf+jZ8av/87x0ZBMRuUaBYgzkhXY
NBcHviyZ9bB3KJyBkv6Z9WQZ3owL0dnEmpfnpjC55kPWtnZoDjvaOkJhZCD6DhG+
MKcGpP8CXihF/lFGSLv4C818GBXtkgmNDzNlk2WvhjDZLGWxJByvLd1jJy7Tocb+
nAbpiOfX+ftO/e5lGqzr/+Sq7OsRypE6u0FFRIThkN4juPwaTn6a9kR6yp2TxRrP
TcS4cSPfgOT9aJ94yiMt3ZsfnX678y+8vfLwnCM7QT/mNyGXf7bbNA7sDXrR64Sn
vF/9aOZbDyOnxKuHzFCbMF0OJWnwgIp36avcrnwQNELGTcgAPhFOo9O5yo+7ZyUh
poBw/9e2t8uPK0Y8rn4uj8XnLiZfDqVDax38t/JxQI4ZLidMtPW46duq3uQqIIXP
Xfzh8cRejPRAmZKewxTBnVF1qmMYNEQbdcpqFVm546qEw7zaqGWDtN4Nim818X/A
csRpTq7bHsa5PaYVwIUidnTl/OSl/qV4bNkJSHjVuKR1H5pccFLhZnW8br3axpwk
hEIzDpWK3xL40RPOnF5us25L8fH7XwmDpc423p7DomiXLikORpZB5ojOBLx8FPmp
x3wQpzcMQNcOLbtiXEbwfGPwi/k4aHzyPCZ5el1oJ7XKRF8kNxHQ/3pHXyJXqt06
m0P8fi1X21yz5+ozx8HDfZw3U8UjDGQBVlHhvIg3/Yy/TKCJK//8aZQu+GATH9Kz
mDzr7CiEtv8U6gPZdhd0pC/cJ5yJZxI4otpaUx2bqR34RWJb/ocedqtfRrjWsRZ9
erZZZPl2IfQ1sUaw8vS/ZX+uRcxDqDdAz2Rm1J7y1G71PcYrvKP64I0yKmKV+MqY
IMK6Gu3GBRGcKk2/BCys1C4Lk3wq38+r9JRqrrtiJZFampg9L335SOKrvDPpqLOu
UCI3GhoNqOelcmpQleNZBzkNnNigBjGW4/6niWiv06Ly0oxYs3T/H2teohZviAwr
FndAzPHKCH3goOyPvg9Li8896tCdal7m3wXQCvNdxME4SUSxLejEAg2epHWZMWM5
2K765VgrxIIlAJKiGeajjHQp7sXp/Gdel5+4N3Mb8eJZr9CQ383EYGEucWmBX3nT
/73u1f4Mk3ERmzhwHhchegx3c4qP8W6LZmP3HcQwp8MS90Ht2K/wPiiKvMmUpsPe
zwQqKUKSaaEcsOyz9gqX1vZs/zB3WkCxtQiiX9VKHihVEz8YoRk1rBUCpm2ppFZ8
gqN5F6tS8FBMcnyiyO5W5SGTiMRx5VksJBITOcFabS/oIKsGAp2tMEK5XX9apB9W
dWmM/Xc7oh6lorvD+YfsQlPKsx+hR02c2cyyRxEtW49l/nUCjoVis8vMlMumhgiw
kVVlbrORW1IbjQxUlK8/anOGjh/A6riIeaIrPbRT6qYWI2efasFXQWgg2eAbTlZT
FyrSB4mRmqObNz/1hYfiZaoq75yswPeOGX34YbJWKg9DapLL0Pm2Hn1oN0Xd79T9
I3CULh5vN/6YYrsqAL3UVuzL513/Qhxxrcnie/if3B2qog7EBrRBwhTq8yCbwXjN
iN10qndvhHP3+ZOd/zMp12UHewL+LLocsxw6LLpSYlPUdi3BBjs6SjTMcpb0Ioxi
oal64c0N1vJLmsjwXgoZci3QWFdnobXWeq81u7i/bqq3SXkZIXatW32cLUb7dkfG
kpGp5yYYsjzE6U3X00ZQjBJ6TvG0BnKpIKN7o0Y4KCQriIkecOFdRb7CqgWr8YdN
RF/6MzYB1Kh68H7tsHybMmFRDFTi4zt32JQaqV+9FuAO4+stIvEJn6iPFJk1JGry
mPqf9wcGQWZA//n02G7CUaCA84xzrR2hWVT2sgR4TErdfXXlBlnYp44Hy9cmGzZV
KoK8gpgIQqlNrzlKzSf8tTjBM7o/7ciQLq3AMVemHuR/qoiSUs812ygDuOYmY8L6
iq5A7TZOKBK+CeSAyC7dOm0JbLcCXUJaBsRhxaSIR4Mf038xrLSy7AOc2n2U0Das
aLsT35jEm7NdkjO8osq616NLO+UB2Iptm8mnmW9d0pe+KTI776ZT/043UuooosNA
T8Fo7cF5/cUmsSoxiFWt8/npmiAQmFw30ZyNKC0uAgdTrkf7P1HPm52anhs0zcSv
JhV9JU5zP3LMfI44Udre1NyWB9oobacO5bCL8ydbfwJ+xQGKk+wB0IlW19Kuu2ps
B/w89rFeSuwIq2OLR5BlIFyHaDca5tJlUUUvlSt21l6cVcFaF2DDSn/MsyTIdrmO
I1JRtaXPlaU7HExkilqtYZrUSd7xZRAUD0Z9VDGKws4zF8xNqB5wuEeKqjZe8B3H
7n+vTY2sTqoNlfQIebMYab2vnCMgOx0vc36r6Afk6MedjUm0M9vcnxye5byc4u+t
cCz/An2IXXQvXD0+9y/WCmmjZTXxeJzPj62skX3wQtEF3hGRMeUvYP2y6bDmdTF0
SKrLkAKNmx4+DDumby5sLdf4K1hJqAqN+qs3vaqBFi3k2mJbBXB2k9rwrTiAVrs/
UjXd07ZAHehUYR2HcYbWclnKxVDBWZQUJ1l1GInV5b0PyQzemm8YOyjQ1OWajBep
kBxPpi936NRdggAQIY2Sg6lVTwxp3qeScUQBpUmrK0BoL4G9YrxiSbmI9mZFWMV9
Uj6sjni5sqYl+siDxJ9OTCUQKaIO/PAkHYrLP/q6jMKwjrB/7Bi+01H13hYNwH0Z
KdNbhT/7Ij1n0Mn3og6D68n8DmHIVdOHDuLt3Uu/drPd65+dKY9XBaGm/YG+BWkY
TjxJ6O7E6lv+D+WAyh+Jv7nFphbP4yZi1Dj50eRokTXbkmlWaH4mOtNnUzJO+OEY
kP/YCIbloYMTxptBw8bwxDwOwW/KLGWQi2L4RzIlplBxGjkxwf/RO72WhJ0dls7d
G3rergP7uuJxyHesHJQi73uli89pT27HjOGoZgW7gSTIxvy1Mj8VSDiaAL5PoNzH
rjuspnzZyFqdzXjZgp+rLv++MySqGBrq5KpHV7gGSEteFdUadBnWLv9YdR+ym3vi
bdHQtQ879qzDKBHlAogIPqJalqSMfk95hESRU2DiEz+eZa7YjK25PXtfMtFQKFV5
traKjBoW+Mf6wfbMKs50zWJx3ajXUZOj8sC7zmrd1LyCDL+TiV6MamyrXLCaO/HX
tHc7F5OK5B2DrmgCXnRlCRmZmjjJwsEpInjlQnLJeE4Zo1yhhR6NgTIRErMsHcXU
YzdqlzkTQLn+DnmMiGeJ+tNA6qZfD6V6RS+uixBvPg3rszs6NOZDgJhYrpm1U6QK
8t1LtMHUsWY0V6IY9UxTrOuO2iCKjco9pEkc+y236htgQ8YdFy+ydz7/uC64wR7h
3oR45bylzST6fTLW3cLiJV2Y8uW1pnVplTDCXqslHVO0ToVbwxVeEVcnzxiCCOuy
FGwiv2tJ6di8gDNSxUDyuP5X8xLcone6/x4RHNiVIqWd+0F8laIzrLUI4LbzPX8O
rx5nc9WMIhG0nOmuQVIkU1BJq76MFziLLfIPJfvw+xZg67TghRwnLIl3J2fDi2H7
9KURWjGYKGjiQGh0LsovMKY97yLVVlPskqI+wPCb/2wqgdwm2A8wPCPRovEsO+cM
hHHVf4WCZLf3SsIh/iwnC0/Y/dZX6MmwURmFKPeBLyxDjpZQ3Abe47ExKn2bE+h7
gcKzMtk+jZIcUmGpUd869ScUif5k1TtUu2MKfG0XLsT/fruw1PBjsi8NSbWNLv4T
7LQr4z5LZGnRHX5AlW8y6VLLMnjdkDRf/VEUt1k3Q7xw8lBStk3fjXCpM7a7xMfe
LLZtawJ3vxWt1dioePaSBChfqa9L0Uehg9E+kCPuAUpKKWQGJFx6L9fThBByd/Kp
CkKsrFfbL5Adz00mMji2oTcAjF3cQeRoUKr+53sL0PZBPz2B5+84EYYMVJZB/PAl
Wuv/EKIaxmZHXqLikLI9kemB0FauhTqNyiiRVHY4iqQYiwxnBzeq41ytlxDPYPWw
P9e/frhoXqNWGjYtToKP72WvNenxmFKu3EL6hv+rUQh4QjLGZR3QfDfR7ioolR2D
JrUEtwopgy9DItYj7PhFZzPQilvaok0QQaqs40WG0gn3CEJd1h4Ftc36jUZahvKc
przVc0GF2oet52dzympA9BrjeBbJ6TP6+XM98kPVvSUt35285dsGXIR3G59KquH6
Nd7807v1cLXKbZLoXRR+lQ0/d06VM1644x8tz09NSiVMVjdzA0okYiVdjmK6SULU
QRcYrFfQ0MXye4fXHpBErDaw7I/f3xDGqSfS8IW9X7VZYWKVUys9FxpqDJQwlBdG
GA/amBLQugjzgHuVKDjbw7/QoDlBXi6KiCkfP7Zg5TQDJeg7Jupz+2qg4yOR4mAR
g46RXoRolsr0zj0dJT2/v6mR3/JVa7LvZYwV5BiGGuNakF9kV4s7+CK5ORtiDwag
NzanuP2Ht5DWeYn8ehsfP4gt7HDhJv20jjZDHpk8NuWOQnd+ps6AKE30SMqUfkK2
nkVp8rA8c/T+XOPAjAsnH832NvETq1fH3CXH2IFLDwVlmZ3eLaSEo3upwB+5RXCs
IfKFyxJofuDaTwf5Lj5y/kpAWc4oNRcIfWuIBEWbeWk7aEnyb3SjlUq1S87skeol
AdPB49yt1A/R2pVt4x/aYCAWlyqZ2EmZA1rV09E1xvPNcYdY48RJrf9a+D9JonYo
TKDB755hCDLNVYEcOy5cvI3zH6Frtdi6MlNuo0usQs0QrAALR39tyhYufl3xCi0r
1NXfYsjb9o2dxobzjsSQEg1tOmXB+ZSpU8dzA1ArMCuWn/CTmU2oTLWc/YFw4XRM
PbRpGf7bSv4ILL941Rt+DBUJ3TZfooGuKIuugKWziK8tOpkjekAtwpS1HkVbzDs4
/dC02SwlHfNtjJFITMoqsDLGQRo9PPUKhCrRaA/nYQI2SxIMU+Qnh3UhLXDdO0Xs
W8r2LlKnHEwVzHjmn4dS1APHzO18aQVSaiVD9m5OdOSpmzk2cx1Up+6bVYYcn4ZY
0C8OMaB2uiXegLdyYR0OiA7PKEui8CQpBGDfW9IjK8038LCBoe8tg9ehYhbTKr/u
5sAuqHUnvUUR7iQZ1pevCi3TLBjH54PPBmAUyGACwF/tRno7tdZt1z9yj+4r4M2w
gX9ZQIRZuM7aM/dNbsEwe2UrwFRvQPKraKEoZim6A1SETJxYZGnHFMnUnkp0WxcI
Hmp7U6j8YZXnJ4FgaS4i5UIZbD4XcRjd9FhM7cUgGRWsiVOAxfLJNTU6oJQWlw3i
O1763XlzlYLHmHfcO7iAP3bzSfPJ9vha+MYx887ZXCm/wipwFSsekzn+lu3XG6eL
I1F+GqgQOtT5U9FCgN2r9niJQ20eD6GDgIuBlGcoBOufC6RiKC/dpBqPh5gGulrD
eRkVcGE9i1X5v1RB4q4cIgMNInveAsvaa8n0RjNIPBlpkaTbfc1E0Q37o7++0pGt
UEXJo0zAtIIwRupgtgB7POxwfupu6U3u2N/45BP4bDyO5RWuRZq+DLJiREJHZr/k
cSvJRwnPgIGx1oF+pX2kP8yR9xNf1xngKLW1Ibj/tx9BZNmrbN5nXPBeZxYptUri
vUI3uvW5+HsCwMUYmdgR5aKdynbGm1tbLfhNhTy38qBs9P780jhNG4GOtDMBPqXd
UbI9++fHhRBIhhK4PKIQuuDbI5m0m/6ub7v6jbMSDRX8yFd+4szE3njKEp6ycpcg
JrxOhRA3zzJjJjFMLh3VqU2UPCXS0J4YEKr2yFlbX1F8D3epHCgLeCf7gzgVyUOP
b7ybYmjeI8mwfOs4sch5bX7Wn1GfRiDyU6IhKD0MS7GtT+i+X2dXmBxEwCU/0OzN
oUcbUGU1SYN/ICZn2awwOBci5jzfIRA3/r4MgZZLodZQIY1fi5qBhXTq/WkA9Gwm
OdYZkTUD9ecjsvYNQL3RESdmeWKBfNFZT3b8WZmLgMC6rvdBQii8sCul+Fnjreed
Bi+5NIXD++1A2Rtgd8AM6r5QshWxjnCP82ecPXxfcts4YsmJr2/KAC3Pt3nKsnlY
fcCFfWGaRTgKpqOHY7fFIMER8ULfI4bmWbUiBMWo/KPdPn/xv0Mx2cy4iv+40Ram
BvEvH7Q8fsiM4NZNVQtGlX+X49SJVg56Qm+T7tEALylI3VL1yI7lInefM8EkEWqy
mbjr5s4pbQXtHcWopKHAX1G8kS5lMG3corfHuCnJ0ECGyw/ZFrdPDFPkwzQlRz2h
l4eT8J2EQQzNHQAQCXT3WBYGLr+z1C96CsJPUEuLpek1124XugbnN8Oeq8pEoFG4
S6sV+hCvpZMdC9WxQl07GPLov9BUX+WfwAY8o+aepuOKuNnNkXU+NcOWXsRmv0jx
aEa6Ca1hNW6pW+HWgxYu4XAEA8E65QdJDKghV2HGUIqzdc2+ikyKs/6Vj1dSeE+U
ab8GjvEXZxqIoRuINUbOQR/9mRXrQe+1y4U3/8h7hq47yw0DtwmMtnvlG61QkS3b
Rh2Wn/kKOPsocYR0mdbn7yAJ3NaeLuGyeVZ8sMHVxTma/U2aJeKURXfKn9TlIzne
u/QW0gEGfzEzbCQLLgtCiF9hBieGSf++iZmGoFJo8IcoNfh9+SQdnIaPifDNFy3P
LDc9sID/l0i25TYO5DeyOLMYkHq4IxKiNrHr7ioUrI0km+Rm6gbjEYY50aknCsEE
1M9ZYfdTdcUpopYr3yCjy6n4AKn+tf4KNbJYqNtEsOpgdfnaYCyJfYFA9+lgWr66
qnRGsgW+SvRsdIkd4EwMKnsNsjihBchnU/FJP8QxDICSdX3UEYY5PG7QfgCjZJuq
tjkKENw+J9iqzKFVOq4gb7CrC3ekMXQV2IdNENYbStI9klmTowgXLCP6ZWIfI7a9
ATvWOj4nkas4wSr2J+U4tMqZg75jTXswXV2qUVh5N2tsB++nul3F7qJxFMqrAxx/
Q06buYj4cte3QoxngWUCsnzL27CClSMeVEeVx8Cvyw6D/VFwUM/yOgUOCp2OcEf2
eDrp7GCfRhu/OLqF/wGzRGVGncQdEpxcSiobrVANT0QcZWRkg8JxDEvRsZ9whTNy
d+AaG3hy7/3JhZXs3BK/FBPfNcezPqCnd7lsVlFCgOoK4iiiEfft6TfPAKHcDLfl
GSwYHXpRttupGiwQvzd6D2lIjDJRRoxvyrRw9OP0cfqqzGohfVvDPgNZYYGq1+ZL
CFB3HbIthnSxYgeOdmMDQbPxBpJZbtohOSscLiRiGRTsaDkSlA9wGqK5qDnXfFE/
klWGY0L6gRoA31cpKAu8X8PDcvbTxhSJbhoiMXkcCxozuhGkdgsTXZ4QnShwx8HG
dJDBgsTx/eosoFoNBdUtvA9lzc2M2PnpqcrfMrREtm2rCNSnfVYUYocMe1jrueMz
L9xUGAo6ubSot5oFDqq5XC4jOw3XRu6RjDwbHas21ezrj+UJI48a5RaqhX1kFbDo
tXUtxG2CnTfLozldhtFlIAO0f7pEAP4yW0/wgoSRZ4LIpiytvFeHu1dmDLCSDEK7
jq5k8lflp8yRZmUPa6rRGzWGgAyn4KQ+46eq3K2FdwuaJIrmh0ufaYZNigoSrYv+
fbyfVKruOfQKk7R1/2y0lM6S7pjpPK7R2ZqLW29GKq52dckHOcbX/RWcAE8uLK+E
uQ1NO2Tsh26vV/8XZELioEoCStJ/GrLFarMVSHNsvr+YLwIswyGWH4zcpLsxAeWn
teScqz9rJgpi9ebNMKghjxSVAAvYQ3maWE6UggkVwwL2hZMd9+hZb5zubhQQ2QUG
hjwH5nfNW/U8eGlPh8Oxqiyycy5fGnD3hpB0jNSXGcbK7QxZsFAEMMOHQ8w5Xhg6
bhxB53SDrlizEoyDWGptu6MnTSQRdwJlLDckyTUSuxKz2DJf3J2IOssc2mjdusxU
W4ObLge6L/FRfJKgNpTzInu+gm6nUqgM3yBoNwze2vSWXtxCP8l7XthuuQGIzf/O
ZaOUD1Q/kwQMF0Tg88FENvlMa0BSIS4BSODbay6Iis4r3QFiGYJ5+zmb0M8PfSVK
9quhCzbYCtF9VajZqTOZkbS8k1UCLJnVpGPtytfHLq1dxVgfX4K88I8pJD1+pIVD
OvLFtXoFyVLBFu6nzVmmSeXxGmS11JFVKtdK+wOFNkwQHKHGs+CnWTrVO4phO39B
JvzvhFUAyX3GrGoKGMCqFgJNRl2UCiX+BxuZXNYvN4Yg/LYRJvNA8s2PKiV3dcRO
kiMucfE6fC7LL6Wn5w9fpyw1RqqQa2qQvYnD6momtRpR5toSn0xnTeYySYmDB7jP
aL0dgVkEo3MiG+QzUdyw/Np6vvNpyozlpj7wGDDBTu/UiQO2gNaE20stQnLSPNG/
xGTaXDSxDp0rIx7GHTVkkFQ5xPbBIR+V6fUeTzrCaVWLobkU54fMBBzUfWmT59GW
SX+u/sjq+sZQfh+PfoDUNa5uItUbqBLWWHJKSct+ppfciBMlLXVe3qNjGddmMgnk
kqWZS2QVeBypbEAkVaqbzCHOhJMyvzBnlpD/lWB1J3Gpl2DzDqdMwKG8XvXHj+ji
2QDL6UEtZ9t2X52Z9vPL5Oj6gD3E17/p/h5DEkRAwAr6mrlJen3JmAWDez+xajif
QhJLpA6tGUjrPwnYJDuphX7XS4poV7pPykQ1aAs2AzIAldXL62815b3CUoj4ZSfk
Gf3ViX4JHvuZ2YxjrmmQZTJDdVmXmXqsUmF9ZRzl3xWXImTTchRTWz9ldMVSC3f/
nVOsvtl9s2jAV/fBQ5m8gfaNtZ1crkh9Vin8h0dFkGNX9Yv0rtsiTX66FhJhxDhd
nDWOkopuBzEM5VbL3SdA1p4mmkp5fxMR1cj/mxuD17QEySeeGTRMGxzn+hh61VsP
/3AOWs5TSzpd91VXMCaQjpj7YdrTFI7ixEnaNfJvrPqhh7/dsGJmihlhZtdy5/7A
5yQJF8mKTVeLDCmN94C2aBbJxu+9RXMqBkq7ikXQ/40OJg8lLsN9gIWSyFPrvWtq
OYqTZSdNvYpnDBwjaZs3WRuDVkPETgxIZiCm51YLKcOxVmJyg/Jr7/7onj9txjFx
NT0TIydNn1jPq2iHalvwaaqhUj+H8ZW2yDthrQF/P1CipxDYPuhcZ++20M0uU7i9
gcB2YthdhucKiO1/5W4kXlQ+uuydHK80EXxowLvCs8f9ovpfaBpTtMpMelgCaI7H
/Is4RfkAKl75O/HH6JVEzESBsEpZezLvtszoPeEPNdhUeA55bG+E/Jkl+mkRn3yH
HWtmmuPhbMMy2At6NqyoFWOTM/7naU+yGEl+5+xRtGYrgeB+fDM/1YK7S/PhhbDv
wtBf9h1PBJARi7Az0HfHg6htVqAqKsECyEjv3EvCdNBFxVmbUYrM3pOZ+1XEaS3w
Ah3Cy6yri+xVsTq2s9tzbzfZUccDeawhqkFZpfJy8TswjP33uD9BA5cKhacS37Ek
mhkK8t9crbQ/7GK2bp8qxUBCEakiRdXj/baREoP9aNCHrcPp1Y7mTcb5NOdOPQOr
RC616RTKFcFw5/4kn/RYi0/ahyF1+gdPkQCJmLnhbJOYXbtgLe9+szBkcRzB5bm/
mBIj/sg+MAF3XjEwFKrXeub+UxYV7DM7UYrwtrQOiuSPUlfuXdxaHrLwooaoixLD
RjbiZLqfL/qjutMl2fGO+Cpts4mtGSTGcfCFfLS+rqfWSvzg9dOiT7aY/6Bhh9ae
8iO93omu06shs/8fz0G7CY+qGtKG12x1JYOCzC1ipLA6lUuyA5bbwmAoO2msDLzv
1ljPcXDv+cbRMFedRS6rEtODQ+TiMahD17xfuVfRax4PMZP/OM/opWk0A954JixJ
EodP36+ifMQjm55pNLxt24IKWTXTI9gYZB4Rs/xZD1uCMktvtkQTyp4nZZw+71jP
zCm6361jsyWKJ3xNlP78rojpgva84ohESUKlm985miS2Cjf+schk8g0Z6pJ2F9jG
Uaw+T0OUeT8WVCAVgC3UnZpnPVx4QVPsfRsCyiDMNOeqR3jANAqWlClsEBQmDjcj
P8SDs2AXqDlFsZqntdlaKJ40n6hdqTZWWuhRGKiRmw4W1gL6Lv2H5uzPwoXW3AfQ
SLy5SdhJZET9Go1z8MqvzPRZjJlNn8+xJc0jWa0eY7g1sWQz16iLIV6o9aI109wz
abVpo44D+b5SsqCBgufOwmT0JgTuOZyPe/RLKcssKSK0T+urNkC/lkPfjTeN89QK
JXL2XFLJSVQLAiCJdZoGQscboKnwKdyUgBBk47L4Yjk4cHLLCfP1M54AtE/5Cvpw
F1wmYM4ByK+DoEHYbrhyPZzjOxOJDTFhP7HnirPLbZexcYoRalJy1IbhRksDqhW4
iCzm5cVy1EF1Uro/C4kmd94hEWNMUn9RwuvCUh/nKWxZp6ph4Q2E3SPoQY3WJPvn
w4e1QwcNhnUp/HyqG68XqAWDfl7HNOV8eImL8i7JfizuEd91q5ats+YJ6CuIpkyH
JKP9rMq9eta4+24VVLjGPQ/H4w7G4sxhI0onZmt/XdobEbOmO/QZkzzoRtYk2DIb
x11+V8i3jDv8zaHNEbmLT77ZHNy+RFG+ZY+DxHAJcKdDKRs6CFnQtc+CMxBxxIA7
Jg5PpkjEmJBunOnxu2lYp5H2nhMah2SSgbFCHDkshDsGFUG4ho0wT07Sj0g8/cU6
qlZccFGi/KHYnc47NCXNIs1SORRIjdKNKIAe5eOT7d4QU39qjIyCKo2ZlkPgPg+3
2vbkTp/UE0jtZKLJqbaHhU8+aNTwE8oP2N2VDDaVCeEF17Kmd7/OOV8iTDyrgqB0
VkRvssP/Er/iXaLAaCeO6hDdZG/y1ImZzBAg2qcr4XvYCuDdQc8op8VAGbTLOrak
/fPyG79X4REOkhK27nLE6BmSC6pBUVobKnaDf0YtREx5M+QoebpJkDixlaJxg3oY
PUSZJc/lOs8JdZ3+mANAUGKYrCfD/NCuCZU7UjKZQi5zh0FfK8tW9mWgcVfknQLV
zGS6ZjteqTb3TGtGfAxCrvFRaurlQ+5GHlifRYRMOk7AA1CH4Un2foYfNtkK1z5Y
9ow4TPCgyxiSNOxjc8afaK/Dp/LscASV606scYVDXbxJs7XY9/Ll5QBXutjzZCnh
z36MXOqzR62RiJJF+o5aBUQJ0CtJVA7CKLkxkAXvCdbB89fV0spX2G1t1hYq0KBH
ZkAQAzQx0RVcd1baWpIguT9GIHqgdNT0besKx/AjerphtNz+kXc5si1Og88zTd44
anS6PJiPNYvxVyRJaX+hWEUyfumZTSSrs6o+NICmvWuTn6VQOoP2imaG1pD/dpXb
Fme4WSX/e8schypof7l9vVqEa+K6EhTqu2HpER1xROksJYclAch0g+72extWqai8
HLdGByfnlKxYl2N/5bqzY/ufEe5tmywL5jrJ96cY167x1QnRLB9HbdTjHnukRVvT
K3c33BuPYgz5pRWzJCfUUnxbm2TsDPmIHEI4hn1bWYxZ6mMuklO7Gr9nU07+RIPS
Cugxx+mnZSqovrJ9STOw8ITsUWG3YSMwt9mzpK5DLOFigfHW3Wi5yTTFa0DKBeRJ
wtFeCPmuY3B3zYiEBreDnty8y0XV76+8eZq+p85ZvfU7GthyQ3GtpRc3JLxrvAlk
4tB7IZOI1DKPIN/rcW6mhQuKX3DKtxoNbCWtSgLNy8/re2iQUPAo3ZoyLv16XQBs
Ao1t0HrJFwuWGm8hCYPi+m0W5gp7krn7HIqN209Wghq5v4lscNzyjHzbIzhWLEUy
hfJpjr12J7cFqyN6RlJ03pGqHTIzV9ljck8+hX7JJDrYYRHEA95YW4sfHfLWK4cO
Gcq96ORuwtryzpOBgzcN7kk6OJ2aJBtA/eEejpoRdMCdy8iMdEcZe0vEFdgFlM2s
bmLey9+97Btl+zawJOm7jfVTvqIgug9MzDUsyOUQd+4zDgKw+AdcPaKBP1R5jf6o
6dSmelRawoTG3+iiq15z6fr5yVFghlvj6lWMKj6JOABD1mGAyzyjuTLOJ2ulGjG4
cpVSn3icgy23Eoi8sG2pWaAzLHwDvaZhmX/OWiunoIxQ7cpFkdCYaB90e8ZKICNM
yGhb7qUCO9Q+FPLRqikfsAQNn1uU3cPfb5dyN8cG/9KzD1O6r8PRiPnK3hK/xK4u
je7X5AkOOs57iS68f6zCGfAAAbXxHNl5ojP8DJfkKBSwwuSHoTw3olrjtRer4tBF
rVqI2OBio+VqZ1I+U22U6Jd50Zgweh+ViRK3DHWsuYFnljG5qMSrSYi1GxHvnbkp
IUh7sM3kikdq04FPTZkfrKp2ft7+fCfwNaPtgGcgauQBq8acqWtaBBdEIe1SC3fm
/Lpt942pk55NSw25Ej1/FK7E1KbW34OUvNviN0xB01wPryFLF/dnaupo8Q3/1WAB
OAeaN9Qyq0nNJNqQgCHN+aRtQdhcIwEWY5ZpN9NpTRe7vMOy0DZpVNpLSx9Kg3yD
3c+beB2g2de4gMoska2zy0EjS7e1Ag6dkjqIA2odVKhfKs/bJV4l/ifzp5srSQ3f
dMZCMu4LliZBvKOEFwtgI5ONlambgGUvB5IVBvKcLn5rGLvWKfcACOBicG3VAUAJ
mE+piKUXw8Sg1shKR+C+HfRSbmkb/Tt5QVrLRuQ8ou58kOosZL9/t6xWwYUHlBob
QCpcz2Z53oxEJQeabdqS9tvo4hemS45A9IOXP4aCClwRvtyOSjDYr9z3mncFjbKo
nhyglw14iPDov/L6BmGUMtJU2VCmDlEHEhy0VaeoV+ccWNVgoUpzixkbrmL90+SS
pjJWQ93EEMQD8znWoZbvZ70HBcIx59U6Qyq/M88ebBSdNIGnYbaoBBxRAVFtfbUX
7/NIYmXm27qyh8K15NX5l+deuWgkaXTNmYz5vyl/nXnWdBPTcqrpRjpE/6VvV1yb
yeBWYZDaRzYj4ImyiK8NR8hDAmtp9unjEiWb9pw7F+dSFbTzgBvNIY2W4/9TWhPB
BKRFiH2Arp/XsCU/gOS3+owwjm99HFj14IHnUMmmXoHK9U8y2Wq0TrFpiJpV51nj
KTPnO4TCg8XLfL1Vc9i27v7zxfv+KVfqCU+bBrvAGgWtDlm5ebgBTQO1stIa+O2f
CDRIXZuDoMnVXz07S218I1z6kpWZRdXcPTUbX/13KmO/FHry+61+6LX54vJ2ieqh
TJOXr8hHxvgqHFjuce/6QAsbQTsyaSOyUGFyIbN2X+x+BFdxzi9Vn0I0QHjpBgIa
dGN0Sk2cbCk17vWy/vJoakpy5O4LOwsPYVIrcH4MBhNVA/GRDKw9bueEepKZpEdV
IWtqQraBFuJJMtjTdmTy88jGK8oKMHQl25wKLcK1KJnwB7GkqKf8tnssQXo61DKQ
kqZIJtm7KeqRPEiXvzf9GLQp0iqsW68T5j/Vr0hXMssRq12AI8dyqts4cXu1pnWN
CWgsId8x5fl/fckG6vxm0baXzeXE+2ie2qzBx9UAP51LqQgedmBye1UNbogcYycp
wjVNGcoaxlrrYmFlQsi3uP/1KhuWfXq21/ywljbFifUzhxoW0RiLoqEB46tosMF1
H9N5xGBG/G6dmTdbEEMZJKaxSY8A6GbLJfPdfXXWkso8OG5DSsTPDpv2GdiuwYL1
r8V/VJN0vAMF9qWiWGedFE84fASX5TTeXkh9Gwl8zQG44PFEq6CIekn65bAKCm8z
y6xqo95hVfg7yK8VeW2pLfAni0Hb6HIJRJX0qSho5WZyBMb8tJjdlKqC+5UV6bXX
CaPtiEX7Ts5SEZio7rmWL8C5zuWkIK5PFJsU5NUDyk3BQy68zdKwuc05wFxHmC/G
dHXIm6so/HU39kuqcAoRRpo9Ps7OAGvHVt8PYHrjltRbL1P6YU+MsUi1TMZjn8AP
W88Vw2MdGvBZPS+yMglKrNYLQA6D9ki1RjAc0swQgV9g27F/JzPXwHGnrE2A/E9d
K8LWGkkmI2BB/eCbJQBEmt/Hke4Mmahp2rNVjden4VYDsN+zNJXcNOyiBmfkegY7
T/dlN6XO9REhPd/wKvsIvqkNEL8bA6z+eKgA6EU6U13Pgr4Sfu3t5FSQOmx3vMAG
4jm2DCE09qWr5cfK3VEQBxm+Ul5uYDuVp8pRAZYcm2AR6KG89HK/6tEyfAzVp5br
ewIxft8GjKQ1PHwyvpW7B7H8Lqvyzia9EQTnFRzF9ZRLexN75eY6IbCvuA3u1Xlo
U7DJQEEPSOxP4Ymn3kLzS2olMp0TDwVmPxTIrx7ky3E7nNZNjKrSLP/71z3dwCFO
uk2MJb5/pSJ/eXBYdr9LZGsdq2JKQ/5AHvdWs2MBBKOdbg0oaOgOJeEzEb/+pOfV
/8tM4jWB9C4m4I16qyrm20W1kTBCeU/LIpA/S1pn3TWmXeLJOQ8AGeGdabgp7xUY
I8ZUnsdK1a6qi1S3IMzvGo6fZ8HtZ+uNyVy/Vmts72HiRprR9Ifrx9B/UX8c4HNu
X4Mw0r7lxgKK6rgydviRDs/po0ZHN7gJnXUSxoWzmimLN5y76oNfCCaOroWPF7EF
Kp/51OV6+ienOs8Ce0KUIJgscVvcwRhMOGCstUm3Wbwd4tB4M2TZ+QLisEqfCPpY
Cf1HGNuYheIA/e+a2oThYlPZgwMeh45afNAAa7oTKlDsFkRXGYYSqa7VuvFRFaJQ
W5jo5f+A6Kznv8Ea7PyFZYXddPGTEiTd/MTa7DoNaMSg1Ej3ygHInL3ml+kMDcX3
WeokyPV3Tyzn335FaEulMhd24dbks/UHUnk7K9T0zTfiR5YkAZVRjeCBnRq6ye8s
Ijp1dKZzk3ArthpgLbeVxrv+sdBQyL7QSoWZpN3D2co8KWnrqNbr0VtbVQIW6yXW
S9t2bg9y6daAyQ5/1p52kQuBg8MCUEREj1PHK0fxoeAoELQbcW+PHU0OgrdFH3Z1
0vrIVzDv3B0R9LjiXbvy2Qcp1jGF0m9e6l5ef595eQZuKWpWwtadblV4w+JB0qOn
jCkfkmKZZ99pXls8/sZ7HTWeszEyvWycbCehd0Q5Oa1XtL6ybpDUpAuBdtNGS5ka
XALtI5xZjTJnO0acCrAwcZmznyLchDBDBLpXt+067cQ1EvgmGIgr3clfFQx6tcy0
SneSXLL7YUnhjWkQVtxDkDGXPocJiObzmaYsF7ZHy9I0r+Vo5+1qTwmZVzAEtXd7
+InPOj1jm+hu8vAcTm7go35/F5TVWNvnqAvUc46w5u+jaX47q8lzDMdfSeJJgZoT
VvMtRlQlMBv2q3AC3wEuqjG0AMo1/s1IbwVpJmIbFUTkqguG5JwjSvd15IRb2tCM
NfCwCfq+x7CeLbAnXBbFmyNujrKk9h4FXtxswbcNYnWC1yitIuCkMu5TPekxluyS
qXGgEp0DGo+r2VlVlMtyncWHeRVucqC6eRsYc0PB0pCr4emyggYRn0S1qVHPK6SS
oxXoENpyW/eLyrWb5BcNCnrYVfW7AJMbcI+QudHdC/JMqQUflpAPnR3xc53n1IDJ
lUU5nNJenkXi9SHTJuETWXhi5Qlr5s885OvusmYK7G/B9i2oR0UhdEoLlKQQ//AY
MGhLJ7S4jM9fSteKFV3S5vU+eJ00yD2lVN6Pr8BPfmwtDl0J6DAA4XjHuVHJaNfi
wxwwcVjiX6vET+0vxH9Dzy7sNXRXU+pACvfNeV+JQMt8ahLw1wR+VBRJaBWgn2vl
MABSKOnk7TmmaAZPW+yVhvcw34uKxwZcwv9oUERUFRik6asIHQvVUoBGfL66qj0A
aqHbaqbcPOfidePlIDDuovJYuuWjDP0+gfI1IXDta4DVUscxlPDIDZoqVA0w4xAb
SxJYM17IdfxMs1ho0Gax8KIgv3Ngs0tvz+qsyckyvOp0961Cj6teNjYQxO39AT4R
RSx4QAJ/6EwamI2XzUwwFWKVtiNwwaePbOkbZwkxC0O0DxQcUBnel7Hna81Qnw40
9rppVsL4bNyKVPx5XVOOrQ9dGGA7/X+TMDDpfFxAxrE9pykvoaXjs2tsK3Z/MUzN
Zn1BmlxAm0Z6jvWBwPz2d5H31u/8vKDZ6ilQZU++cED3KQorjGx6mVBUBFveI001
EB0JOy6fzHBSvmvi5Lbw0A8/I09u2x3EQO+c2NKFGEQe1rW7EXBdN+lQXQRazwju
U1Qza4238k4TmAofhE4q3GpR54OtTzf2Ev736CZuTwk8zFQLTF822c0D9ir6jq02
qSizCDiL0mT81Pq44WF+4rLw1TqMlsHbDqmHFFPr0oHei5r1iEJbzd174g2aUXjm
WBktqWZq2VHzOZO9p/1NOHlKbt5UN3rwT7L+xH3loHNdKrr9GO0pseHBZHC2lYRI
IFnxiRf3y1Fw0aJxhNfv3HP3Tn45R5tzcyY3C0ieJpyANheLFkKv++VfKT1rGcmY
TruVF4NMGbDMAuEmspFwGopAjQBqtZUABOijBK1xVwXPK64fmnt3r/9Fq0ShWbe/
mHeJerCSxYqo/iZNhd+NPDwR2Nil1S7lUf4xSjF5RMxjQyYrMCp8MHwSVnSz34Rl
CqJ2UfHt4qfx1pHsYxnFz2CMjdShaWYLWOq5HzfgIjBpQbAGnhxKWYRYkKdR+ItD
JYhjU4DcwaWRR9R9er3BAClHgpzYb6HiAyBuXJ6LX0Y7SbnIAljCPeNXYZC11PhE
8wxCFG66pqWHOjFhzwimOho+wRs5rR3z4+qjLZEOo7QBqALIHGHH+aIJyGfOurvf
+iZxlvabf6pchPygRYmU3O0EChAj1QXRse34jEMblSRgs5JBgSnT48BqT01GQYpL
YJyx+WmMlZ7o6UMA1NEWLQRrsKN/22gFIQJU2m9PMwNG3p4CgoZTjqyWbamDFoDx
tCaISGWByY3NRP8P92Vnpu0qCRrXOeahu0d6MVv/TYvTRR9TA0vSr3pehuGQI/z4
jUmnisUq+cpmBji2tM4VZ8Z0b+m53pVEVXPLGb/7TBsJ/xhf3wRGIDKihyl9Kn1N
8mr+vNBGgwa8xtYU1av1TgrjgGRqwzcWPPLrNehzJNcM9qKFAYpXWgI2TimLqucV
w7sC0pP9e5nFwJbviqFmWYg6sbB2deteXu13xTPI6MNfzimxuO3c1N6sPSTQ3tIi
ORhPfPwog9oY9UhA5QQk5jFXeMhN2CuCqLBthIQZ2h1Cf+V0sOejDI47ZuGaT+Ve
U0rb739TmxIo9KkrrTHqLCTBinZmCExrU9Qxxw0wpdPcySf0PIS/sohwdAV3Rg1Z
c73j8m9l6Qx76l4z4u7bjp+qjcZyCSVezoasv4+CUEipaUwiYeb2B+naf6GxdKOV
ntr4cpITI+2AgUa6MwE10vrSmQVrgxERk5atGTkCursWuj2mxreUmtq5gbMmxnod
xlYHzYdWTFEfssWpL2F6yUe3YFcG8ogm5UdRD3pAOU5w2tO+dua75eNGBfxE+jye
YhA/I1UxIkEmad6MhFAQ5T8YAnY3vkqTPlxM1t3U6tmW5SLJlnzxjp9YOkGOlo0X
msOyoL/0tzVOFreHr1yZGZor3cJihT87F8f1nXnbgd+kxNUQM5b7JHL1rXDWfM+R
GG3I13Po3fyLXI98yoX5WxN2Htj3XAQAetf2tLRUAjX1oAGo2ZJ3zGRkMszri68o
tbHva9GGQhvcmX3C8uMFITVPLDehVHJXgFOLP/SIsSOuxufIIjvXVDOzvdIO8sUo
pfsAW4rc6a9yx6Xsg7g5iqPH547XAUDCnKdjhf+aVX5w9WV0Pb0s6LzLCci1xuuB
qLKMguduv8E6tcT6BSTVMfh++4uWVSwCQk9dkKCyjT9VptMUl9jokeGvEtUXPETu
jvH9yndtMc3lHwblsUwFBidmdjom6lvExx2Q61m+4q8EISkjUbhJFASTThlnkiW/
qRtqcJf+yXpJzzhevkjyVoiSu8rlH7VYVM7piBDj6Z/32Ht/YrSPtmdd/sbBzD3s
lWnfYX8rMSDYxg8KtTxFnD1SeKFqHH/lae2n18bPgpbfyJ9NxBJLtw9W57B2aFM5
HN+mJ569k1bJ6WHYdWMvl6bFddYQEJe78ES2LvKhXduSJbmbdg1ips/Lhe1vqCUK
V20+W3jElRFBXTiKDXl6jl4reYjNYImUr3YXAm3z9R3MMvx938ciE1wNZ5xZR3M8
O5nkqBqCkR6Vt8jx2gsaPzckDWjJPcFFyZrxPj+BT/5i5ukA+f5B0nl3P+YsiyBo
hd+5xwV6yDEkdkItTSOWDYr3Kkb3YHjdNuGDOf9ZX3boQp1yWlrbroJCpJrcIypN
Hm4v0wVk/FNvplVeKSRYGRLsNzqgzKPb8qh8Lj97DtDqYbrDCJOtTfVnI8MDJY9t
BJ/2MguEBJf7cKoTp3pktCnQcbIaeXqnEzJKOyeEuhbWv4GVrn8eC16y2+Az+xSo
MTQfY5xPJjs7l/t0oT5W9ZJ9JpAmrMTPhSZ/cZvU5mzhNal2Xgn8PHoJnjwkSLGW
Lm3UpaubECBEbwhXszEJICLXYb70gZArbzNRXW4ZBFgARUcAJ7kqfLVM1xoijL1i
QtUM6BlbLXijy+eYlKuR7AOWb0l2dzXmV3gngoCOY/m2slNJlSgoDbS9ZV1ul6Jw
SOoeKjZIrq/WsgRZN/pse+NXmulXeD5SSxY5NoxsLf7Z5jzQxVQ1C3B8Qg/mhVxl
nnSGqMRfzoTBplMZ4+uSBHyGo0PG/ms7hKdriRMGPcHpcdPJwiDZAmYj/ZgRKODB
p7GJeT7P/SvPxz27UyDBZQwF5kj7cF86hGOPGDA64MawOv3MDzEMAYwo0krGH4Y7
hjM8751psZEaSjXh8sUmTsiIlKtzpltsRhgZLHCzpCvQRvlQQTqlX7SmkMCzX93t
2wOCGVFU1OVOGeXTOdq3oDuzcl/lMIr7k8Qr3z9FiiUq7ZT12cEA4yN4tK9HLfzC
S0w/1OSvoqzbTYsDnjE2rObNxLuk2qB9RUuGD9ZEaWx9/bALZQuJMdpJNwExFsjz
iTBO5bHHU9vGUGgXPrumQ2f3SYaWsawTti9N9Kk+szplhsPvOJJ9sDnmID4tl0yY
4ML4Q/CXSUjJ1VYMOS3W7lGeNZ/MQreJoBmO/xT6mn7ph0MnsUfDaR7DP+qT/H6N
FE9yJkB23C0tCAiCZkT9UKN7WrIZJl9bMPyrvPylHcBV6axosr3hWHRrA3+LvjvP
ibvKdWKj6vh5xX85/5iyFDKmjMc4wv+veJNrAB12Ght+MQUgllQWlEUmaqijnVop
yge0YLPyTWrWfiTwQq5QaMm8q40+7rGb5nBjCHwnjwvLzQMAFqg8AZDeKmc2xCYp
UC+DcBuNbX4pjeG1s8hirS+xlKScJledhP3Of2p7f/S0zi0QvoWArgV/UOVq+xod
ZVe1Dr71HJ1lrsZ4FIgrw8gqoTqVHLqRrjLvl3y38bS+/qNgxsm9/9FHJoOSDlsk
RelBObqe99ElJAVyGkoSDT2HQtMzmeVNY040FUZdN4UoF9b8dMZ+Ke1DIYl5isII
GuzIcS99gSWpefNk1GnRkcQOPHL8BlfhIaNuM71+TR6T7sWnlBXwURhtBAsnfkw9
lApTTnThjj8Bk2tnDs+R1tI/PoQIxmDvd/XA7Vl//IE0HV1oiOzsS5n2lqUDfJxz
9lsx20i4gMI7iDySKU42eGICAQJrHfg1LFrKmoCZ0Fli8X6NDlbP5e6nKi3uBjUm
6D0KO9zVQjZIXRNN0EmOlo19leQzYgblyUWl8c618bz0wUkz5APurpCRGAYQgtOw
nsGXAG1pJ5yGMa053NWqhgEjKdNDpkXH/SAgTkKCGGuS0g7Q/qR6XmvfcRaSI2C0
9V5LuFeRWLfEqe8ZOjSypXriX4Hy1uoadVGki56zE/19LQHqVcqgkxJf/KNKGxMc
Ak0f2c42EwdzbM3aI4V2dal+CiM0Om+xVSKfHgW2XBUUHs0gXj61wCdN1R9k+sj2
X3/Ovrg8wnmagbp740cwDLLWSA8Qhjqv1yfsIUqJ8RylguRtuAtRNs7e+WnTMXaX
KpLm1LKy3icI2EpWM6e9FCreO25r8bNc8X2qcDrNp2yZb8KfWGPns5W+19hDmOUg
1zOHliDnSXktoWS+mZ3Zv3xavbThmgk0PB9PJnzx81S8OHWmMr1RU4ahstyySvhw
kG23II0mADXFh/7cWBuHHqIo1TAzt6d8c3Z1/DuuACMw+SeLtHFD8xbT2Jm2gtr1
G5Fk8+sb1ahG9CUh/XFiiGrAoP+GyLCFsemiZNvkTaX0D+9sErv7nLghrI28Lwl7
cMcC8DkZz4wxtSxl8f9Ef8Yzv4X7CkKqltYIjY0CtKFiX6jF+ZxyHGNMmOmWWXPL
2bHPrukepUldjdFvkRHiwasJewnFCWF66ONvHzIHDx5aixEyMKlqoN9DBOPAaUn3
930i6ztU2kEXcj9p4rNZxJYW33GZK43SIoWduhQnQsaws2EVaWHg2+Wvycnw688w
fPGRhRmTlGnFQO27F9FQZhlGWosImZgfiR0rjhWzeQfV6D7Sp5ed1l3HgJ6+dZF2
gyfLzESPV9/Ipm0DtdFh+et0GOzLJ5ukJgKIt/Zi9xT7MxH41uYpVYGyeCkqpHLE
ayP+00xCQ35nr6OnOs8i87+/DgP2ga/nya1kb6ZcD4MPVpzWkqSe2zjlXlNXERyb
0kBgzzn58k4JnDM4vhGoT+n9U7lG08kZvHkgHZc0DVMAa1Z8TXfIWLPKR03FkpU6
M6IPtWQi034fBtabnek9IVTvoxzboLjx3tU3mfvOGPxpdIulS4c6ztz5Kj7G5BhM
C2euzaLpL/CIe6Yr6Xll91I6om4KElmVFEkLUdJzF2pW5vWFEYt/wqZNlEIx7fcW
PDM2mZpXBvl9Tjdqbv5noNxzqUUsPSOzHXQoPD5MShiHu7o9X570e3G9grtIAnAv
ZKxAkXnDfxKQkXCA8IdLvMApwvTYR6k0Tkj7sxQpDylHTQYW93QzGJkjA22Ov6Z3
XBUBnQ2/E1aSxuzo0D8ppkyoKhO+MEpQxMhG0HWBTtN81dZSDC4nQ02OYWRUadvq
IjWbwAH8cAcExE9L19drhGv/17tKhSksgkpgi6IH9To3VT+3jJsvZjfpdsu6eliA
I3co+tPLiKXlZ2Fwg7zAbYz6T6+t9/lBsBFeYU/u7+4pcSLmf+ok7HdhIqYQFO29
a5bTiG43AXau79lwBxEWP8xPU0PHyc4qrRPraeI2Vc9iLoVO+sWvbupImYEm2cyK
NX2yXG3JhPMaO+E8faayzHrT2dxN9GSzgLqOBhyuQq+PElrfRJehrWFCaSvNp9Be
zZQYL1CuaceEhnEZmchtP3Mgp8EHm9gtdfKNhG4oR4fz1OMPrkFOnMc3vIuJBciO
d13tdO3M36f+VGuJEDSoOnWbMVkHijKAcZfgzWkyl++4Dsr922zvJFVzxf34B3GD
1ZVWYDe6WRg3FfPgygyqmSR1zLsoH0t/1tRBIXnUQsNmHsFEK1jQEfcN3VS9t2wW
GxXAogoxoYxk0W0kRjuIg2i8Cgy3Q2/sYUH7qxgXjc1jzjWGxTbblT0PHNV7Jcok
szEKGO/zk/oKQPVrWGjegeE1R0GG6G2jtXcL/BvxgKNbpgpKQWKGlwuLwVTR6F/6
2Vx05HlB/6zuD5yfiUvPxAvV+KX8QRjdCbL8cirw0JXzjleofo5/Dw5L3oS8yh3w
Q8E2i0i3Nva8DpZJoSfsnsJW5wW6ucwA+oTZRRED8MVAk+BeV2OkKiOfSQRWcvvZ
QFC5NJQGxeL7Qg3GN2H7V934tbcychV7PgHdwR6NbI6n5lTyqBfgJXOLPNYok8JS
YGaUMVm508BpmGuweiaROwkLZfJenNThvFPlnP6Z3llkhirQrkENkHCMkA9Ox4ZU
TxztDXmEN9BQIYQA1mJuOKoDo4HDoplr1UexGr9sfMbZzGzfgF1kPD0mk4ifhiYh
5VkkR0n9wQGo507CEnFhtxkfAzR1s+xD4V1G19WWaolmLVHhRZ/q5FFnBdYiKqDv
T92iEaq7em9zq6ZJC6uV1TKd3Jd4+3YOYfr1dxLJF9or8+ijx5moajZcbI+0BnZJ
xGOiu+bAxZCKbduovjpxS+tDOBdqQcwXi01B9yWKPw0D6UqSAFpPu8M+x/Q38ikO
2cIsfpVF3nMBLL9zvJye95wwsbaF7xJ8up4HLCu+4j6mHfC2+cj5/h6WJ6ZSOFam
YX/jcmo2HWI9WMpiJU0qu6+LEmnMZqEGNUMzCgpDHSqLVDh54QCzIBcu5/qWw+sQ
pgkn/mZkKrkLFqs/lfT7W9deEZcsxyNttHCs6gINF1+AB30a3YGX1ehz9gvxqjWp
tbUW3UMfcX/U7GiOAsUdEHvBehtEdG1Cc10hdwEsTeRcmal2U5mRX2I+gYeHywsX
peouLSpcEcQ6vqVxATfgd1BLke66S9p5M1ViSLLMixfcUJ3Co+AkebAfYiQV2DUC
1TbrtpUckQRxJ8W5D0UV8FfmV3nkJ0Pq4JmgoTWpJcmtlloEFNQUHUDo7tsSmUDD
IxMKppsRgmMoJ1Jn7UjRv6egUyNHdo4r3SBloj1QiyEJWzKyZA9ZxBHjd0Qu1gFZ
hT3n4OmZ5E3sBT6bZT0JsWBgcm3zCLaYHA5mVtOl2AD20tp8AY1jRQhM3kFALdAG
Ny+17ffrnCxIn+XXiMlYfOxsCXOpKP1zmjGP+bK36+wGP2Bueea0CiDN85B1RyX8
1khTLx1ZWW80pM7J3Hcp5vc6a7HD/iAjez7/v/nWu8EeXz/dIYrH7WIeepPEX7Pg
Co9olD+PeWstv8ekVsibAyJFfDhP/s+Oev202zGE18IRncfTb3/+hkIH7xFRbX+i
C3O65UNvL1BR8EyQLpHNj7xdOw5nHs448b1Yr6yzK5ClsE0evKDa/Na0+dzBnU5J
DdDVcTmI4vdNY4z3tCbTXUMDJuaSEx6wE2PIna7F1joVnktlR3c3BM1Nle94I18L
d+4I1wMn7D2Yt/vX3HpmioE587ryW/uj7OQUWxlVbG4v/IqTEk0O5+/wbvltgXYa
Q1IBZsKsvGddOhMtV6Yji0SDyE7wCIV9bMuM4cITHSjbDgjU9GkTZuLLfi0svcsm
MT8FSvAtkqSEDsTPNF+wWi/vlhrRsxGoi+nc0Z5eT4SwqSPEKV3eqrFq/7ICPtMd
KhHviw/C5vLbhUMBkqb5mYNuROUr6MZRdHEm5Dd9J+kuDeDoyHxofmKH7IqkOiwe
9pbpXQRs1fix7Wdr2Y74OuKi/zdcroigH5tnLDWvlFbbbf7PiXIdUQGCcD64jTNZ
FDiFaR9Hkx0inCl8ldGlPrUK0SlFka5mI1KGjlPoF+M0WH0BSP/bUNJrIv8DOj++
XLYz8rGQUjPYkt30kWt0B5QyS0/vPiI0tLe2dMQJdt6Ctt/WcfyFK27LqwaLjSlP
DIjDW3jfgoNALRKDkHmYth5HHg6W/urlsaEsaMgb7n1Bcb273I0SmgvWZDLNlj4G
+NLB3PaLYxCUhkrlhnxT21NH49TP8/PTAB4ttvihsdYljTKNOt12rt2qCIECKs3i
bMz2CYV1KtYShHgkOTgrTJOe6GZikFWIq9eD0EfPVTVSkriAGD2M2NWt9qfmhjgM
lDlE7sykBunAQm1dpLevIeiJUBLgjwsGFuYEoVZxPH+oIxgNj44/ghZGpD5IlgkH
oFeEUkOF2XCS4lCwxGXht/rwTOxI2q2WZKk2gDs2n4t5ezldHiiO8EAsbNiVg+kS
4MiV/jnXvsOW2eQgpiUahBFjo+W1+XV6Y9zzcffTIOVHPa+M9eNrZ0IBgVwOjhae
zagqqll1E0YPWZCFY2VVcYkxTs+05dSirtnfgGgNoyWxqEVP5v5/q+2HjZj3pvyi
fbLYlEG983b1jY1K4zLk39VOGoO4zVfScoO4NiukLc2a/ewEMLRELugv47lJfPcd
YyacDraZ4+qdPtZhEEza4jCfS6KLorsXkyXh0ODj5biw3NjOxkqzjOqzJpsgyWjy
mNVQttOWLVyiC6rgMpGW10SU8GOo1nmdPnAnJCk1DOjq/PZHhoqg7hzDG5wbDbXs
1FoTAoZ/1CzxKIw0ysrqVnd7eeAF2PXn5/KLgPhkLztNLrEaJScNgesq0KK5Rjjp
Omv4etEZy7YumrQ6sJSTnxFwhbw4LhoWhB+7xz8wVCoASAMwV5w0mYgcbGP7rNTz
ERxdJiLLJc8USujxTF4IsHMb/PfOQEhZ1vSjpgCZLSNB3NdYitadGN6BrIScxT6b
YLX4xbI3162wdNfSF0SkUbh9qiql7OeqGFH3F/oO6yoX9Hou6x+FvVuHf6lrf1iC
RRGzpoJq2nSEnb2WxWWYmsCa//YlWMhwPMQgDqtcEWdNdJa7myVuTunQKVrPycnA
Vls4EYYYJG3mywxi6RmzrsNuTXP109DS3taHMd9a9jCXWpzhKUlBMFJRwsE7Cxyd
5P4kfi+AFT8Vmdc5/HgczwdfOfjM2twVMFeng8HT2yPf0lyJURis4QFdZFazJXpb
MiFI0PoApV3/HUidLZJ2S0kNBhBixbFeLmYLIIA/ZdQvRUwpxAChX81ivUbP7bIh
9kIC7o8c+zR74Kjj0mxUpEG9dKX3iCWom9hmXZmOATp4K3ea15HilU4iRRoR8DoQ
JZfrghuX/pEf8lmGmySub8MtDsGpVW/GhDxursiXQHvijWR99ZMZJ/z3iAScM/53
Wiya0uSUtJScQ2nwkMApCgOUl8yso0SNxwP9QT3L5vMbqm57lY1NWjz9UCSowF42
nzu2oGQ7gQ2lmeFxP+cBJA6B2R+HGu25PX5H565qbrIAidY1D2sSiZySC04tPJ86
lgaUbxWNspeEqQH92Yn68JmhV7jB6pZ4sEHrbgLdAsC9uXLMykWIsqDaySk1bd8y
iseqCh8My2WyswQH6yuTaFOjbeiwF3W+W+LyF/mnDlAM6bgaYDh3JNnmudfCEgJa
DmLp8tvq/k5yu0Ccilz/NdHZWcrXIyjWbXNx5YhOdxEK0pjkNugQC4Gx0Fm9DpbT
sJ4goLsEh3h7HtqYqNW4jB3DzYilPOWrQnNGJNStfs/kfNw+YPJCG2Ai7fOyW3O0
sFI0q9o8Vcq617xExugxVKhAUveA8fQYXD5tAIAFRz8hUOhDCgkv7SN89Jw7gafu
clvQE4xgVhQu9kXHasbt4cdkcqWUEHsk4M9/cXRR/r0iXwvVlDnVaqEIKUzZ4BqB
8aXCOLZ8PyYnTuiShcD3Cp/0UcJWKIXkOL7+aJVsc06VLf06UL3djmWGC1XryUyO
R0TojMU9oMoo3ygU3OE5GapU635O6lajxx0WfRF3M6Box5+p0xu4wH7mpOUx6trU
MgYr9vtukf2wxRsQ+tkAJWTcmS3BxNjHf6uwOX66Ml99S+awk0AZ4/O/UTXrJZlh
QjPIEUuUpaUjlCMHS/GV9eh1WX5n0i2H+2t0odf/rQheZik23++/s/95eL3B7IAZ
v0QN8cBTF5S0d/PaB0hR2kaG554XZMu3DJPCpyEyHs5EXiFmymP3u/7mhQd9wee6
qwwWTSPFf8c9vWVGcwb8bGaQl0Yjjc2hYDrN11RVGO4Rz/sJ7lysmW1IvWv5Oodr
nQadaunSQFXnY478NyfikU2gOz5yhS5fF4FvhTXwaFlJV0oxQbOYSRZ7aAOtdHCm
U60URlEslzL29n4Af3OJDsprsghpfgQY0Xxyl3VzgxOs3V6KOajTS5EbgknQvx9E
mwADpEzD375JN9wlTeLHGN4B1FKSwuxGSpdMBD4DH5G5mkL/wCTcxGGhgPZeMlx7
k6x0vP1B0uJfsE7TaJiFpBk3w4GQ2Z7chpfkPRCrZyHwB/OgF7kDtnJ8wHp7I3so
qmGIPevX/JKoK4yoUWMYpMpeR8ePpEEhYmhYEruGZ65nc/+i1Aip/z/DiCUI8/h+
4p0BH/7fiOcMXPdfSWL0+OxNpqyef0UvZQ75sMk+CdpCDMkd2fxtKMh5a8YYo6ai
LrO5w0LI5yhGysNlJiSBiRloFBJNK9qkUV5Yq3sU9Wxe19hEzhSvQr1TI0BexotN
UOF8nxy+0QpDo284vs47GwYPT6qA1q4FGlKlHTjpk+PPpxt9HX2yxNQiQDhYCUbn
e/66NvUYoUOFP1gcpN9xWXY3iAN1yvV4EtB5WuKymcuQd9NiyZ6ha/5ihRSq//Mq
FTbzCyGDavXHyl90f1fshOxN8R6zsfTd3Cno4delkJDHtkm+xEyxmLuyeL7QtnN7
GlINYYyieGXIA9OxI2MWsXMn2grHzbrLh9RWk3Cxljsh71Z6vgydTKgSQLAc8Q0e
O7Wh7n91uhBqJi7raVcrzWe6Y6CBnvN4CM9gcYfM0CwXsboIQJnA+GWRiuSH82ID
W0bI2E8nbpAB7QCkeEtrtGAstYwZQtCnsUVc9J/tRJ0lBgFhU42Go0KfKDq5qfaE
/Dmkbl6lpgOklzA2WD9nFSiutlprJYWcpXs2xUFUpkvqq6IozIuWHzTgLIZxzQz0
VJ6OMNxxz7IoDr5bn1B12ULQe/qQO2WZPk6hLMU53TBAZPWNu1cNBxBgkUl3yJ9+
AW/hY1334ikmY2SYojok/rcyEccQo5IHAB3lVBfXKRTKyX5VK0Hzevtdxl3xZJ+E
SKl/vCi7EEGX2QtzuzmEqhuTDZYT9mH1JBU7X/T66n9ITM/N/n3Z62MHe+gy10Ux
LoZ7dkpPdEsn++Q2ErbMRF6ny5LabJ9Qx0yeC6Am5d7AYdC6NNM7kTEZCfJM5TN0
SOgYtgen2IWFu1+RpnM9OXT9E7UdR+6aUkeB/vmTO/28LUTqVokrYSHhkN9UCOk1
QjVW1aI4jSR0lx0AVLKgTbbk4P0MHDHVNjQ0Pjo5YNoCWNkftmaOV0vieO0vLlMj
j1YDPWvhmLDtakgp5XvtVJzDHDgiQ6SObfNfqeHXh0mKDUwAS4qikoH8dQUqDskG
aJ9kY74Ugm7ReyibjM18GMBZclFuhUNUk9jTD6nI5D5FEgWKP/wMK9DVT8wcP7UD
Zua7OUiVK4P742D9wnRobE/bMhidy8aKs9yiMOfZHKXWMpLRzcefo0Qx14b4PZqT
h4F8iWqF3gCTe2ARA9Jy0ZAo3djlf2IFQb6758hoNyBbwjOspmLkVL166iShkAmB
JRBUOzAdoQQgal+gcAmKuw8daX3WT/+rDGGTRuE5MsClMv4SU7mbfsuzRIqYpVjt
nZ9ISq9enZUnK7QNmHLULIjtPA1PE9upt2ZpGzPIerzhnQycdbZXNsGJC4kpEfS4
fK55/VCl2TcQ4fr53GWFJmiqvzXYr1SPonUmH44zqmrxY0z+8zB32oKFVKFuqti+
13yHO4RLRfDEHQ20rl2srKzfSVb8JDHrnmgACvhoPN9PCrfH0N3RBH8FbxZQw2zQ
9omSCekhuyx1VHlszu8/ZIm6W7MmKzp8dQ9KrBd9GT91OiruMumaKrXWduPhu2NE
DnPYcDgC8dRGH5qrpp24Vfxveu+JZDeENBZMP9xDsavkUL0tWahD1ohdv/bSGSPS
WtgW+eVK+bpRVO4fSnhA5Eclx14vEgLCJ80FV3MZbiOPj3wouD1TZV2YHJB+Wat4
dHDJwqZv4B6joKaBfTdbRhZSrYLklp8Og6AdwwK4gLByzTx+FP4yYT2k7TpyXy0W
EXy4AOgyRgSLVjI15AWzT/oYDWfOF2swHRU1lbik99XztJRvL+B7FuqVOCJW4V2j
5WqjVrusFGwskPy2mjOkniv6+aKyR1/g6FQTkk1rrb4UEqVq0aBZL/L3kRiNZn8i
XtfrlbDctYa4u8/V492X6jybxlocX2ePu8iXWHu1KF+3i2qLOxVnbkgKSqIYVu6e
DXspUqT05HGYB72oa8C62snKw4sWZw3ulB6GgwDijzOl09wGaec4puGVCm3TeEgl
x3BbdGlxwNN7LTncqqOzSV4/jpY4eNYybW1xzYa5gdh7zLmf38yPYFCzHGpdOqvS
PaTL3rILQTTCtd3Lk9n0c2wZ3KhpqUtv6gA2LaKPqD8V50u9QrYeaxwJi2CZIMY5
mycERxAvSEyW1UToBrelXtPEh6fc39uVIAPPh6u9ejoK6Tab7+FDWtDLtLPrKauT
4Qqj9GisJnc7aL7SEuufyaztIBGP40mMeTRDLXgD+OUdxppUk6F8NRvWsrJh0d+1
bLR3Qj/Z5L5D3S8gD6Js+7Rm1LgfPIZqWt1veJaVcF63VJfiL+AmGQAmmic7yz+A
+2NQ3vRlRORIWH12sMcBsNLgokCrUEVCW8LJXWcwfS2Drzf76PimVfKGjxwhBkVk
Acp09hNLK4Cuv3D1nLf7gfdnnInVQXYd+4y72TG8qIFN0FiZzmehe+Fxfg0LjqLP
4qivXXXPqwdI/tig4QgrbFOqXv/F3dD5m0my9mqQuzPy1J5iakxTeoyvvJDM6Gim
aGobd1pBSE8MGUVTlp1nuk5UajpjDIIYz13+GYXkTXXaUrY9pYCZjWyy4H41t7rz
+wWaQ47BEj5Ird14M8nmLrKuICTamU7eJw6sp/ziTgjYskl3InGCKfzB8U+n5FBf
V3JWE8mmXXiFnVHGPR0+YF3DjA3hpV+Q/QtZERQPSgK3W/KlXUnW80OMbxBfg/rO
8/Ujq/IECYUQdCwgWGL2wjK7il9U63D2lCPuEkzkHNqRXcSeRBTtN1grG5dBnf18
H/yC2WwrERe2DzpqLL/060KpgS9Av7to95EIdZILI9ZVEbr7iek9t84snUAlO6DU
wigDwdDVXOnHlnwEKDna7qJcUZUjjoLgUZxvAAfFkZT8mnkGYawjSxRq1pkwtORV
4yDRnQHvz8HbWpdeAUGFhFTY326/4VwB7gaVMEHTKWWsjoz07fmODjgVnvGLnWrG
BCSHAa7ng0Z2uVPORvd7er40AesA25NhSHARxw/SBaUx+Q2jK2cv/Y7XJN2DknqY
qrE8hUNF8ZaJMrC1mMtMYCc+UcRILkZhjtXlDU68eJGhynxCf7AnKT5KAx2O+pYE
7xYUX/OS1GRUCCdLMks0fjxtV3wqaqlpBxiQLzOKoFWhvWsq0pKZzUABT0b+4Lne
ruAZ0ceYBydyybTbsG+ZsugXC4Q1wVw3cUpG81JtrUAZx3LwUo4DnqbqTQGSwtUu
W6Tgl7Tb35AiZPSPavjR+ySKlaue4zc/YJDtwxvMljTyoLfa84ebVbyq4h6Z33Pp
FMu9UvgBgNVICowxLzHNcpB4BSD3Vhsdshi/z2akIBbIlX52ogutW1EZL8H4tst0
YSa3V1iAO5xlNhL5iGWHw0GZA6Le0Mt8GG4s17zcpOZ5ZsBY1emfcQCmkZ87s5I2
5lLQ23shv6w2axTetzTEDWdIdzWlBwU6vFGq9c5d8qIC+coUo302D/791tEQnjvf
+ecdJ4nH8USOhjzvKcGorYNR0ep1BtmbDOBUcJMvfB6AHjEI7hm7AZrfwRqxEfm3
xzrHhxJuljVpF6GZn+vVdN98ySdPfPadcxiY/nYJFcMv9ja7DxAqHXuzwGtHEh2w
YOk8o2yQ8L1mV3yVaLDs6t9Tpx7YdUIbyZFOIry7GlAR8zGbZipIKwzO2zEkVZK+
ymAxCcTwJ3ZHFA2gTb9E+X+W7+bpFaSFNtRqrxo65ISAN4SEbUWwjK97NDPafZ+c
qfocWnBaqE+jHFY0Rc6wDSX7KoSQkr2fRKrr/baRZzJxqSNGXinSRn9cQVzeM+w5
Sb1KJTxhGaRD6yV5QNP8fE78FSiRvmN7TsMHR0sPruWJRaRcz/f+x/V1Fz9RaUck
PEYnVEvxAhNbPev3MNGA071H6bDi4Z0OXYaX3Q448CoXvZzWVfMbE2XkDZegV5yC
/lFVmOsn6kUtlbUdC/TPKH4CxzCY7p6yLWHfeYLbHhHfSrNEqvZsNypfFAtROrn2
xz2gdI2+TQ6uAsP3f3/3yEP1DvyErc6QNsmvb+OcbVtSKNNt9Wpg+nzzJKKkSsK4
M/SVmTzCGoIGmYYuZahY3ZqW8/fnmIDr5us5Isq8IIC3YAHxm1g+zFIEDU8YBKzx
y93P9tNX/Zf2D6WN3+suxMDQAi4RWb8DKMTVdKXJHRWlK7+0qV/t1xywLKfppy0D
X5/PB9BFnCbfStY+57JLaFUQrFXJCObjDKm+JRILpxHCpayj8DZ2mC+wWjvny+Kh
8U1XfHtlCHGjSc0Q0wDl2mTpnTzJKjHRp4ZDXp9Nh4jcxFqdSMPQLlMCL3UKTZdK
fRhcqf1lJx1h0J8oLhpupV7nmfesOV97dvXk8OWP6msyadPGKwH6F4UT7HB7fdU/
4RPPflFxtMHBqNcDpTffXylOp3lWemV34KckijNPlxxnFFBa201oqrmgAXJS2KRC
7b++p4urMez5unX1VuQXgHeJk4hIEz39Oj9I1R8rGuvjp59DPW3EDP5yScVDdzEX
OBQOeoHJoVbdLaHfHWJRlFAvKek4PVSheM+BqDTEpRX7KrJbIt929YnPjHd40nu5
2+0eOSXKIVGNNRso30UrUMefcV5aZSkcM+gw4XpoM7Rs6VlX1P6YMwnJEGr+bzI5
2d8FF4QUH0RylrtVDaqaZDJEvOfYBbaNAVwWmhds+Wb4G3vFrfTudHLEpEmKbQbc
MAyLsImPnCrdvRDEHffh6DsMd9so8VsGKRZbQF//JqgJgvfzbgWJkXWSUE0oijG6
YoSvW0x7pL7jJZp2POSPcp5hrgvYdizjelHz1y09A/bMGnAUx5COtvUQg2jO7UgL
ZO0roeDsqg8XcpgdqFMJcmkZOYPacjMuEWHnbYoId7HXaZCN8UHinXFQtuUm1eX3
hcS9eNCdLpqTEyNLzcDOo4/WdPBiCvJ63R1RQQKlRZnwsd1T2SzwmWjVikDKdjbK
K3Q95zCwkT+V+hxXxOWxVKKFZQnYzR1vEhpmrait9WjBoBx4RdglQpQFBVTwKurT
kt/ERwTF/nEG7p1c9MDPNyJQLyqRlJysfu/Qwpz2lddJU/7P6oDSDvRqtqqyRupj
Gzv8cIPWXP7CxnDGb1p1rhzL3e9OSPSwRxt/10FpV5uhT4634z9OuC8l7PMak2Eo
hXLGlRozAcjfUvbT5rFoTGmoPnmvMa0dxc1QfxshUXccQW8RofWO8Xwylnlb54Wx
LW5I0/BVjRgdccXMF808BC2pn7HuAeETnE9c7MPDS6bc3WC865FIBeVMOurmrLMK
kB2lBxjmRKiLBqv1b9QY0BnD+xji3z/SvnOS0hGADcMQ/abABTr7WqlqTU9ebTN4
qv6WNm5E+CeaQLhtEl0tVGbsG6/YHl6UWPJxk9Hu7qv2a5HeFSrkq4sPB5NvGdoR
AjOP/0XUICH5+V0cxVmRL7CBEp0vXodqjTxoSogavyONjuf0F7J1WHr8JvkBP/4B
7nPbv2TmKjX2yuEsX1qPwAQvs4jIsEX/TLoZyAx+rVGoDwrzbuZ4AKkkw3ZYKPLx
w4UL/yMuMan1VaVLSfTFabJ097LiDsNGUIpxFQlsloyd9apAo8iQTKEdYgUgXOSo
JyEckixZ94KRQlda5sfxUoFp8glD+PV7eaEh/beclD8DJVMd7ciYrNcPeVhN7RXY
sDuxbjsU6X5j0GneHU3r3w9DyIrias02tl/d9hW+EZSEDVgMKI+joiLXdW8gyUt6
OqNvuwCUUNsurREGh7wJgbb4H1DbT1wq+8vnFb3c8qoUc7dQ75TN1mZk1Ct5rdSt
NblIg+IlB/img8zQ+JcCCa/BhKw0WOzaY36Qw4Dd3cT3nikbeQxTyiSmOHD/yOcV
f++nePFEpSTxEIKqKG/3u3BYTnQDskyNNKzKy37vNcxdO4w7jH7gL6NOxp1+uSuP
75+VNcNrWKSNJTHl4CpfPMSr8xHufvrQmhvWqeu77NttxZiMVSVrKswZpotjIAv9
ZHE3gWRMxDEyIjp+7ik2iTg5NmnsCEaFnWi4HsMh/qBeqHwMvJSXYDKJUvmRfjUn
KQw54MQGsGxvBm/nKD/coBp4JpLwksZIH+p/VDY9ZsQ3Hyr7PSrU3KQZyZCU9hYz
bDnpg7SF5NOFRHPdCCiFPGRFgJllTpHnA4YkrgMULu3xspoPv90t3nOCOOcYaQ4K
Owg+VYrOrMgkPJBJSKG9BSQGWwBkRvIbgfZPtrdDY1YMSZCaW72vK/KfMFk24Dwf
XHUWs873iNjazMsEogei6l3WglomWPTGIU17ZteQRFlJh/Lq4TkCms0rKV5bZl9I
jl/vf1ttt8IlPXo7s7Gkva1jfGcEKGp0G7e6eDD9+RbAx2tlz3iKvp8dSwHhhvDz
tniFSnJBbuC9+dIGbQEvHJt/hrtWRgmYDI90Q0FnxqTbz9Jax22G1KOBg/fIHvAG
ANO0SLyrAAqMDSJpWchPsrVfzf+TEHKABCgkgtFeXuADhT/tNej0jwdZHjfWC+Wq
12AkxMPvlxWhmc6pRVDIVa+KhygSwxOHeDS7sJT0IHjXADFU8YL+HXCCeboK7S06
ez8H94v8kYEYNVkQiEFlSYxnz4Snc+BffceVzs09FYTnHXKOEP2Q302MrJ+2N6g0
qpg9NPgnCAaHggG81oAgF9cmIjIZ1d5r2lA3W0zzPyR+sU+9yakOWJ8MACZg5eFA
27gY5XvXm+qtH2il1yEmuGtoeKLgtBLdjR3TeNN0Nxcf9D8vw7kD9uoB64FdG8xO
iDPT+MT5Bbwjo8Ln31zZYgVrClS6eyd2+uLGSxcjhdhq/+AWlK9Q4Gl6AZfXca//
WlPAomwV99LwS8z/wKzxvwcbSrRrvU5B/0oO2HWPSxgVmJfpFllJ2D7dWmCr1Yfo
CIUwZIFRAoxmSZwkmoSyvF9b0QVszwn3VYDGuUC8hnpxp29FOqrezIzfqQ/0YgYT
yirY3PSodLRW9+dCEdowee6AuetFewvl5ojx5Ry9KhDZ2BG7zCoaIZVikMoBhLEq
a9sLnCxYNppcnpBVyNCB6uwlxc0K/soLeiz7q9xgp4q308M3lMQIuWQjs+wvUcLE
I0cK3fNl/S/jDLaKYEr4Vif2CoFIumbMBLaV7AjU/AgHENHN4PciiMMa54JBoWnu
usmJeVTjIgKJDmMfhVhCr5v4a6iViDp5gW97Jf5IO6WL+nOWQhP3RUOhs4Pt2nfw
lESxR6dI4RMJSkgtcBVV4cjrGpZv56aZjUR1401cKV/wUOCpMSNucF9VOASO1b/K
UXJmpbQO+333qsK1+v2b7dHozzZMpyUDfSk5mcOZbnbN1Y+cq0bSpvGdpoXEDoa+
E6oeJbaVEB8saR39MGywtWm8lViFy8rJV/T2gla6CSJenx0UOuERkrFocJZ/DpEc
GX1KvTl4QOYqUWAM+iXQBeUt6CNhI+5at8oPCCyxIY1jNIn7rYLCZWrB1bLq9QlD
1SvTFGiQrHbLVEpdFP0kqVYYCkvvvly4kJxt/oFsuwD8LMDh450sTYNkJxla7hdR
XE+3KXcbytbBqeFMgWoMPq0a7k21ONb3i5ZJFaRaK3Z+QNliJ4Qsq01X4R2pfbfl
OfVD8E8kgdBVH0yH0D10cnNVDFq8wA/qjSu+GiDM/pYN43Y1DnFX8zxmY01CKby9
+2a2EwxtDqRLPNU2H7+NMdS5KsA3x4V61NrXoYQ3SeYD0JgxD3gEPXAIzohoUidq
ztgIwqPNHzniyIYS+rtC3w0xBI1ZmHlkNRDqBwBAr8wFyUGlLKNbIq77BN3O0dKf
ndV2aGUctIsLImywv23yncpxGmuxUCh2qPPsFkrE9JHYVoBsni2uy/4IYJCYg5Qy
XVZO68hmoLUPk0J1xbyqo4lOFESuuaErIh+J/dGzZLUBj9WpJUrioL7ZfQCuqPW0
anSwmokdH3Kr1kZPeVqhikR34HlNg3ElbtZTu3MZqRRYMrTxj2OLhBbPNQJJsvPh
9tUBPaAA+fIDNZbh3OQKi2kRjcpG3W05zKTQU3Ye8Tjvdg73sHZuYpoqqWBq2j76
E5V/HMQv3Q9Xt8nSjYBU1cMyJudc4JINE6nNHcv2q8gHkzSLmbA1Y1kxAn/5yN5r
qVfrScyGE4lvwtowtf5r3z1eOs0HTFZrIfAQRSAHXdosBGV6v0OWgwzMiZsfOATL
50fC0Ew3ciH7aq+e0Rn9UlWZCbUza2y4BYxBkksU+QcFcYSPMpMOlg5ig7BZomrO
auIL3xwBhKTkqmUjrb7Wq+HJ8f8Yg/dupHyOOFx8qIvc75mj7gSA7bCPQiLrele6
K+hoV5wC0ZVyUaNP+/AVZ0ALesmVBuO7s5c0VfaWZJk+bNARHykNm/LQc0MKEv4K
hgEsHXpXxLDA84eG7wqibysIsT91TY6gwmM/lKDbSm4xOcKC+CKooWBCVSUwoUZn
jLOyH8LD/f0ek/ttrC8wQNKwfWYCUt2FkUAuMHbXZ2bLB6m0nBlTd36aLpOyNw0n
+DfudbOdhHxJQaskMZfqpxpGYW3kglpG2nkb5o5WFummTXylRgy8t8UqGXxnhkOI
a4sVPJC4h7nRJYcHn2pNpqMIOAyFc7dx8lMjGKsvDZ78UtbY0eRKP9gLrPG3qgan
gUZuXaxtjoLaLll5c/0lPu0TLb7DTqzA994qkJ1TE/ZjICF0PxVEWRBJOJDiPixq
cnK5VkxV6pZB7nvc79yD8oadrPLuP6gUZa1NN8DAjdTTCC2TjgobVTqpXqW17R0x
HCFzrbuWLYxInNZEHc/2i4EqDWK1DVtal1S6X6eOtmXQ2RsPLBg2UeN0QUat0thC
UBFfxVR6CDHDFNqEYWtD7jvbR2theacFAGcjme9W0LYOJtiQW4jbe/KYUTYFgLIf
WBS71JJVt4H/DYF3ja6F5r7+ks6gSqrh7gav3o9EX7oaZD0alW1137vJhADHh2pp
htzlVtLNjKZ8+oL+kmUL3jf3wbUENDxyNsadWijmRdG4eLYGJy2vJn9X7kfdCm01
nOFIeAJGhYk7PnH2Xa+cYY5KU394n9Yg6z2MMQgAFUDE+4PI04SVIo3pkNWX68bU
mjEyQJ4NAgKZRb00AVRC8m/8D8Sn6I2+zT/xIXQhZYw+Eo97XrffTy2nX+6MLnFa
ibH2nZN/UtMWKSAUsZ4GIuPei3EtnpL3tjsZje0EbVxSxcdil54o1xobUmELIP4s
6FsD/H71lzEEhZdtKB7/S45KFgRLDUdSMJOAaN+AqAZJxpsgVmB3yQPot8AGusSR
n1k2AFpWu+hZI3pKIem7bUHR6AA+rfCJV60TOOEEFFNQr3o8Kuj+6I3Ou27tLBOP
GUl2WFqLmEjCy58AmbO78Kr6tsQEoupBwh3n2kYFNzhiuRi0Obgk4VxeLFX3A059
3pqTZ1sEC2PvckKvKNGtz3vCzsSq8+cqEast04Wj4lcEEnh2Dv/5mR5Xt96NmOtb
3cuXElBf+zwbMc0CtHmu+OKGK2ANdJqQJWicghH689xdQmjH9UyIJ8l2YdvCc4kj
DkldNbSdw9EIJsnyqVAzgJDt3l76Y2WOrPU3JUVxf6tiyssEyM+5fxU0j95I4CDh
5H6L+kMTNS6VJjMLES+D6/n0Ose9dJEtu5nzf4xGRHGnoupGBfhOdwkxqjbIiNn3
QfFh8CNicKc8z1BdhmoLpUnkNnVDcOmZn7sOvOM1R5t0MBffxUjtMiBlbbWM8Gl2
6nRtnvpb0aknKpKxAFRa8pOeKCHTe1wgz1l53HblETqP6oRr/4Wan8aNPgVby5GS
c1Ut3TT+PYm/BRmA1Dla0FLKo11EIJpWG7vDEos3bxqN74KORJmZfIhagkbmPwk9
2TVtfF9P4DL95ZmEqOno4YhArFkmYcNOqdD3VWeIzV5H4MCilRMqxTXOgfsSIB0/
T1e8PVuJUomgSX8yPrsbwAnh+V2ItvR+Jho+YbkejiJxtGEQZdbs27piIjYwtabq
j24jSotZzoH03d6chPoMT9AZD393xkqMoSlkIZmm7+ELXb7jpDw5wp32//LPYoQG
DHmPiwuKJ9RNZLoJa7BEQ/eaVHmsF0oxfWy4kIiwbtPkQNOkib5L7svZlpsvWkI0
/j8CjMEUDmjNQ7rThNpFT+XsJa3R1WdSiIXlNJAg5zN9QNHN2cXHslGsKLoEDjZY
RCEvMb3qSNLFmndR11gbVEjWiniEa30k3K5NkbPaI9vClkkQEHabK58wJzli3GoC
dN47H2O4Q5ourA14ozWvc24TKP7IDTukNNDCXSvlDCRM7Jnz8LHJQqd1wEuPrEkU
SGuCU5M21tELRaUSvvzqfUX+SGAZwPigrdQmGiq5eOlUM3+p5e+Qcem1ZRe5eWzJ
DGGNDl+rKRQbA+6Pqe6V7N+4jWJXnPLC+vwdZ5FTB8EwIA8SAAIT7kV9eywGSdfe
e7TDsKQCnKGMivd/I4ym+6GjpeX8YcqsJH9S1WHuUKveR9xbI3DgYPkPOGoUibZw
u76z0k/dqpmtOIMBLWLiNOxZgNOjuW11MQZyL3MIb7vPysdnxrcoDEgNNRYYYY1t
71ExkExLqq9iVvsBt6nIj2FfJ2pInydYE/oPpk57ZsXXGYYsg+gXmda49sjxP+tJ
bF9CYlS7rHO44uZYJPkfnTsntoZ4N/WJX1K/OsQ3nt/XNDXGkOSGuYUE4P++hJkm
P6nwA2XSclwzYM1rEkG5pPCzutVfkplI5cXAawO9T+sh/gzXpsM2pXjf/kSIuk20
F6kPLXU3wlN2JN9I6YnDFU44ZW9Cp2gqeE7tqWtDvhQLUwiU/3gaxnUhgCZe+lJ0
6kCF9l4i/wKuoEhJkY+4X4wyiUZ2sMvMsn1zbjpulk6Nh5+JUatIRntdP3y+yfjb
Zzc0Df+BlGeKynm8cLKiQxZfLfWTlvoGHrD2OsHDIJpLd3hLlwFp9sVCMfeiO7Ol
r9XnCg9hmEiuu/dqyclgTBNfjt3GpGktprpjGTw9rOgyjF2SVYGPV1EMo2jTA8yl
yOmfsia7UyEPc0sZ7Xbd1PDsQLwWXRhQcu67xZD4uVP6SwsLC9HQKoX0LcuZdvVI
EJ8aQBzhdvxSoR0vd/qgDIjc9fpPUvc8NvOveygBNAtWn2/Rm0skfwCNUeLst+0W
yYc4sfaTBrafUJXLoyTfL5AlR5y7zH6MnN7bKtNjrAFmgtpQKW1/DZUy6BpMO7Nk
xQZh5rW1dSORXsS5qN0JBUjq82UE9hK0KGNKPGIdSx8WdyK09OaNav4/4dm5FWC8
Q796ztLNVnX8MWEuWaTST3eEKe6WEY4HQRUqEdCqRLPqF011R67fXgRo9TcDx6eH
FI4gKavddhWY2sadKuEZGQAW/MwOEUarBeKUqe/Vlq3rl/i+kzSs/YFr3FZF+Lqc
1/PEIRx959dLh7S+RO/pz5isA0POw79U86N1OTMeOewFnVbD/w5ujtEZ0uHNVh8w
+kJOJ0o6A8F2sNY1PFgKxav54rrx++1ncF4VdlgcAj9e4g4x/BsXwkqTBbtpLlVN
UbOzDgN4N104r5AWJO4ymyG0uRA3htKNSUdowDvpavzUJxeoYsAnRWVjWQv6IS/9
Ni9HoD6MD1LNNV5qzOOjthmNO52Sm+3J6DfI84gYvG7rOacmE5MJOTgRuCitYvU5
pSxks0ddGtuT+fiLXccgGHYJ3nMgkYMyAyigXQ6rr8o3lRcgG/yx9CbTbCRXaODx
oq+XpLSoe6LnHGZbkuJr6C8+W3ygNrpAuzlKn0DlBgWzducnEvsfcaIbRbYi7/Fw
LRiI0affI5Xl55m4GdobQ1xpdNoHaKcoty8u6FANMAfW0Vu+UvufrbDTUwmpTt98
jULhVGu2NOVDzhZeeM+5+lFU/gS2xmdNx+/Jcao8k6MGaMv3KSbsBMMuouY+66BB
GrdqvQarxP0ZBl8BTQv7BjlJ8JxxeS4jJ+vs+hcz35L2kVIset0XxTpHwQXga+11
SbzQun8Hm9khMtZL+ejx/j+qGQwQxu84oYznzORn9K4TVRDPMlbkYbaR53Ipqh8/
Jd3L+9yz8L+VdQYRbGL8nzg2pakS63CFZtuCMqXT/ZL3nJH5Mlgb5Y9av8uyjjtu
iyX8VWZJAC/yX//z1cIlSTcrXhZ8ScooMH0T7Ls6VWz6xRRs6790vbjhVC/XoLrs
JNmIi+fKjYomtlcWeDeKQjBc7YuC3IOP/uZDKkjHIrhrxRSqoZoy9GpeB5Wb+jfY
U9GliEB+CaswU0zrnU1kWvrr7Co95gPnIgHD9F43EGdT4JxivhqedrDaXJymIV5o
6GR28ptvtj/cKeEP18+pWlIjDAqafvJ47cQ+pLBngOl6RaI1MLQ0TZ/vTdKAtukb
XlWcwAFOSkgvhAuDvxBiEFlg3tmqoM4mYR7YkbiOQ1rH8b48oUw1REQGlzXkpJHQ
Nn5DjqV6RTlAZYXWzRThke+8zpYmSc56PiMrf2lkulVSJPco7AjJQyOmTXgO/cuV
6NSFKWMnQsOOQ0dEBxwKYky1rEo6wbbbefR5XNbiwddvroiO8RyDzBXdl1Pk+xs6
TxnzqCuRQk7ngPMCX0jAF/rlpTknDgUCrTZVQWQDv43TbdOF6alBRar9pa4T8MxC
dpZuy8Xyfl6znqtsDl5FpLNrxolypZ6aymF3c+E8oPoWrm5XQtSwdRAb3yDjdjVx
XqroSIdqNBHyRhYqAYoBn+IeEcunCNLpR0N9w7qJzvU9BEnjj8Q1Fqy2JUPDr3cI
7wpQKYel7YB410jPs6Tk/q88kdBaHNG+nxm5HVn5Zoi2BdsvPBoPhBzvawNvnQkb
yzgBqZTIe09Y8SkCQha75IQ3MPvr9PgANby4OdwQ/lkr4rfWI1E85dc/mZHgqnE+
PkNML5ciPvEucNP3ya+U3AkrKGOzAlYGoZokA9rmq9/Yb/1DYxUaCxIi6tTfejrB
h+EqW2QA1qNK3rvkrs7cXn4/mVjf3yma8NYdWVw5IU2RWeVqBlrW4t9gLPP2RnKR
69lAXpPo193bVsCA3TEb5njOqKW3yYl2MJ8zMFxZRDApexOjqtRaXpsvozwjTBkU
OyYsuJyiy/7Mrejb5hZydr51eFmEnEJhIRtycvyfrPKb+T7Yo505ydnJ9yxM2UlC
9yXRMAUZmhLfMHJh0r0fGTn+jCs3SUEbNnXI3ZRbJXP60D9HMB9Qbm2VomHXg4o8
hntSWUS6DJ2c4IWcpf+FwRhSLH1isHOBXfc2Bgzidhm38fEAt4SLqfnmGAGd5i9r
+OuDMXbkLI1peG7pcSWq94DwQCVAogZueY42qt0YfLRdRLeiElI1M/p5bu0zU96E
hU2XEXFYhAjxUckdQG6T0X5C9kX9XPfIfGrrkWFJ+LA4MMWqTFUqJrZNEIgSH8KV
u9yiaphyCYyfO4AkUj9Sq79iQ9rOqiZmuVZWeD+Cz3A6fDzNtELmQHDc6Urep8pV
xnvc9Dlo0mEkzpNatcsjfV8VP4D75f4lOS0RYpn02/PIE3dCslbKnaeuI0k7x+8v
o/mnSzdWEoSlwrMLowiEqCwXeWPeha7rRUNeBD4daIuS6VFUR1Rd5HNzHuWeK1aN
3hkkGz966zSz7wgnzXX6+4hs1VSDL3NT5lI8DQFnqewdHS1ZLlXYQcEn9pEr7YBP
fi/orcZqsCUM6xE/QI6hg1GNv0ku0D9gO5NRIXPcvRwdAV6mDAXpxkUXXVHSvsgV
eXDjP5nBI3JZWHVBHWOposLN1pakWErEGQj28rpkonZPGjlE1tynOSpSRtXV/1Wj
IM/HzuCxoPFmqLixPG1OCI9szSmayc/irv7jA3icNnKRapx3p7gLFNmlCCulSCFs
k5BqMVYEZ/7kmQyasfeFzVNCJxMIj6U68LcC1GxSm8LxqDBp+mqSzcHl+/QcjZfY
w+hmO7lBGaxbPe6DhJEIKXJnJ8zXdsctnCLbOYcm89gDsibnnyd21zfqWHWnl1Z8
D04FiHsrsUW1KtoRMRuhNNdUkPUuuG8aqFv3PfgGJQkK0bPzP5JC0QWbD83BJIJp
VE3KOiowPmjcJbxC250qmMr3QXGujXvnxFy8sBq0FPNCMOVvyHWGfAoBW09/jn52
LDqKGsI/U35MTvusWzIcrlxtyrr3IylO1YA9rDPELoKGVxQKHE4yg5PL9wJSMP9F
9xjmTsfmhx1TCWdc8GzlfulyVYuEQvqmIUdrYNFhrqRKAMYZWC6kiEXxeh9zZ96L
7nS+YeqItFoD0uqzYs4b1y08aXyL4/9T+g0k3X0VVkVERg3qZqU0Xi3E6xwenaVf
rRyCsZfWYVcySuxAP8xaYl4ByoJwISx6YsfcCPYBRT3oS/kpjB8DrYyce4JPaNTD
J2q3X251dz7bTKqXYgZETtNzf5oStGmACZrE4lrNHye9JHb6MhqtjnRQp5r3uL9N
5tENuJMMv0yTTQyOh+a/oOPKiNBFe3N1HNmboh3sydwHPJYNcD7XCJKoyXJL3BNi
Yb9NYSsY5Qn2n633RZE4BAFQoUSxemT3Z3QuFHHX7KZXwTkDpaJLlCb2Wdxygmxe
v+p2EtQ+hT0tHzR4d+bFUFV09yyUZ1SBmzaY53H2PmdH8BUSalQgL/efdvK3jgQ2
LclAd1IWBKU4eMo0PxqgCP6b6184lmKqNG371gb3rwTtS6L5+Ll4dgblvoYPnsLE
FVYbFJ834r7tLYUpXWkfAXv5u79hQBhRgGP0H8qHGiSWZdnr0H+R88+/s9oCsKoP
ndVdndurmfr7pOaKcdEmTd1q/2Sp7pcdlaxWcg6FPfycQ7Opnetd2KOyqAckuMmY
LmuX3EmthLap+Sv2/2+xvalq+qUiy03khIQ3SgWxcAB0bniMXHGWEep2IP9PFJzv
rNptchqG6D/6MB6lEOaX7oSGF7aa+alUFm6/nyocrgbiAtnJolwOFbwdrPfvcWhC
avWGjoz9gtqKg9+03/vi4SQMbXB/1iMEsD1Pzch57p3bvaqkLwWm8BNTDcJp5Zdd
+7m+bquO8BvH/yR/SgP0I/lVZe2k7TPn6ucWMsFxdJf0gtLz3SB9D3tI4JnZ+ZVj
m+U4FDGN+Y76iaJ0Wx+8U8FW9t7Cx0ENYPue3mMwVyNNRdfK7C5rZb1WQpCeazaq
9nUrQwvAH/RY2PMjjXTnt1icoLnKnhpwwV7DBV8dBtiwMswaN9appmm1vsq8Sa0a
FbbyuW3MPGFE/dycB0/5qhg2sK5cQR3gWxic1EZOMNEwjWgFFwd2TP1IjzBrGr4S
CHApcXRNAd7y/myf0ShYXM5SWh8KFV67z3s1VOwTtXo60hAXdmwzh952qsyCbpXP
WL6JMJwQEsfceOjDVYKDXZquezJIQqYmi0nvPTOhQlwbsCXuJ5ZcEcmFXmPhBg1S
b9TbXiPqMs5qUsZzRt9ApG4DYaSXKltayS50G3blEVUiP64ECEkxTnuThz/BO4UC
0UqjXhtpccX2ShAQ/mcvGM/cH0kyDr6hp6Xwz5GglK9XggPcdBAtl14ttaCpZq6I
TH8RHxDvkCpTV6ts7C9TyaNlRKccisntqHx0zPiJA7Th/t2GYdT+1a+1yUyhsas8
BNO3WT2wQONU0qbnzGQgU69fv0r8MtmObd3M2/TfL+fjfIiDsLHRLKVAe8IsSLpa
ek+6+30eZhsegXSju1d9QMQpqX4LcyXv5+oyDdeZQKSEThRv9hRsP6/+czoIwiRG
8RdalW3tQSXlZC9qmCnr9Ub2iBpe6sYv1y9Uifp4wQ8gQfWt9/t8fLi9ja7vgEah
es9h3IHJBmBrmHKZ7lkinvGpEie0dfqhV7JSYg0Mn+xq75Xi/c8YUo9ciBJkbLbc
U6oO3n+NFuil7r0BdNLc6AClJGssmE8UbRvWcXg2v4QuMwxdAjTPgP2Uz+fpn1Hl
vlI67EhCkX4/hhnRJFkqg3pwP5a+IjIoGTvHLJMeMsJJY9EaMJj08eCokr3IMIE6
NHXoC4Uyw/a+g7bwmyRbqP/HxeEqVJhRd/HkaiBO3DgF1pS8P1VQ92o+9ylN2Uwb
1s8vWq8jrKaz+OlWNwm2UKNNFH59aVH4MU3P6kHpgLulHvSy1alMsMO1vWQAGQeN
ak2KSC5sutorH1J2lzuEmy0h/5QYEFG1INki+n3z0orbJ5o3b4qZSQP/7fy+vKyu
W6T4a9m3HSirAoKkpnl0mumR6vIUfIdF4Fmtqmrmy4GWQsIm/v+PMpuqfQGLwLe/
ZTpZhZwGGEAI1XDEMOUXYVE7wLobSZMq+0AEOp92d+cuepWYtG8FvnZSDU1OIWCy
ow+qbJFHWdW9LEssGWGrP8ysvPlEYDREv3tIx1ymbG83tSI2OXhAjKKZV+Qw2lnf
41PLJXy3OA+Cmo3MIq3fAnOQ8/2Lqk3vhEHL5mEXJsfdAsznxtFDqUEd4tnCq5vv
qXpGkWbqQa9Q0HQMLzCcbm45YkjyWPqObVlmHqXxo/Hy/QMeBI2C1gwUA0C6tvwo
G7CN9//Iff1qrNO8rXVrpYdYSpAo0gh4R2rePJP7uoUDaEQ3axEUbie92Zwlxmxv
VW1bkilUb0FRyygNnH7qTe3BbseLYXaATssIhKAA8bI6sYQmHJSQff46iJuYCnWx
OSvk/2lHo4SrVEsdZgUX+pLyunWtvUkCphtupZEZl1mRajhEFLSq9F+TTiPdAdRN
2aEx/YTmmBpFf2f2hQLZmHWdq0ucu2dIYc1yOxJDtxBU6G9Jdkedna/7SheSvH8h
VGiyHkTmSUV/RsZ0SQfvQwXcG2fp1BaIye/RQi9EeN1uwBJpYvTPOXa3Xr1+HaKk
omGAVIPGyyUY4He70fP2UEUQ7jqtlXdAZGUVhzld0jdhUDqkuCDKMU3Xikm0vaIH
G/WiBHK5L5akyf/iRqmTYgHHhPDrOXmRVqckaiwxkJGFFFruUWFOwf/Ilyw9hq1H
hy6ISYUgtQdEBnXhEUBZv7Pkrdk88VmYrizWmhQT8w9KucfH6rkzpZ5dvu5oLY+V
Sd+OWKMLnFrg8mm+/itDj5RawcQ/LutivN5H0UvvhXJhAPXh9rhclSVbQgkHniLC
Cth14PZy1EuI04C9YxiXbOcXhTdXj+EB9L7qVkmxsEtEWXGXCXVcWsWraqycaFFI
T6y51kzVs141a5q57eYIaxJtyMrW2hl/Pw0GBZni0lUwJSnZJYI7PPan1dDVY5Ee
6nhJ+X/MteVZ76yB/fsm5uy5GvookoPs5Q2diKjXfy7l3KMxXVkha3oQ9no9fMp9
RlkelVN39EkYwIUWsfE+ZmJsnSdTKQHAFnxMuwbXw8rmO39zsPSCt+Y1npNyatsA
U50PSKYrKhxEB3XsAoZIy4L+kzg5rlxdF05ziQYfwUNmcAiBB+dt7zCXopEcCevq
2lja85j57z/liw8lcewuhbdrbU7P3xfVyeepm67ydaQbOhuln14uB6XLb9HSzAp8
HjzCy2/SmUa0XtnK2GsGadK2a16zP9nT688JFaZgikt97pDJSkO46f7NR7ie23Hg
OHXa3jn4KllTcYnTsgmi81JBS3xioyfTrplinykOd1k0E0DJ1VWEZjZnjvYGBogb
OCiOHxhaDVOjnKOWy6efuK62WbCV+hxN7nXrlrMl0SYv3cI03B7jxTYvapSr53TD
3TdBAuDNch5lsO+r4h6IB/gVdNFTX37xLFhQIxYOEVOqK35UdRpcshBJrT86TOWd
t/0qPagSS2AzMqu1J6UMhLE0haNcf5s3yzJ6hufziBJvQDkXLr/Xu/dYBd4M3T0F
WRbkEwn8Q3uTlxClixTZ+dQ+lzQ9t7o3WSQ/ptmd0Vds1zp5mPixA/cyrRPhZ8JH
7n6rjyWniE84ee14rP+ZaJPwAmdpdh3ezsd1ogvAh4QoNtW8KHjMdBFvOfhybrKX
3/jUHnAUyJRRwCNpr/LbePePZBYww+dBfAdqQKAmwyVDGNG83O2HkYKxEHwwQe2D
pRA/8Po9wrd5CA1Sl1+dXYkCvFSLzlswFO9kWiyFAzcDqzdIM/gUhSGBijM5ElUC
ROmu32BC7FL1W9OVwqMjben71hsFhDhpLd+2C9WiiuBG7cHVKOD1qUiCmbvYAcA5
gra95gk9ITpMoKiXA9aA8OOuJQ4m+PcRnNEyDZN3a5SsecI4jzUL5j7DI/ty6tVD
Jy6YHd/BVorrTC5Ig1Z+/dhSPM+HUJFVp7yvPCQKuPrZ0AXJU2AluTAR7M/0wkLC
CBq6iTYOdGnMMV28YWf/Alaw/dqe9wbv9ATiXPWS4kpIbGZUnMMKlU31k2fAfD2b
uu96tyWFgB+amoRQcWVPD6qLPgAdh9n7qOwO18iveXmo+V11xVQWk+xL+9uF9gxU
kgXzp3XmdG4ETO6kxV9h27danaqmtNNPM5Pny8dS02MAcA74aGFybMDCYcQzpyC6
CB83Y12sqpW/yRy9txyd541ulIX2wB0wsvxezB8L9X8xEV1b3nBOFGa2qKqj9qgg
YDYkv/SuV/elNLklfGRA9oRFwQejfanWOEFFmS5VaUwu3D9B/4scAwaU4i+V9Qya
nloOP+bqBWi0bYmw/gl6iGiXxB/7eSKAe3b3ZkZGWM8+mz1QofdZvc6vjjeG7SWJ
MH2s30+Uq5PJg2GOhNuSFUoentlD5TWVMisvE6eqHa0mWHaQNXXfm147ThC/aijj
HDvLMo9OstfIi/YXXJwa1zldRp8bn7fWVo1eB9qilMLXE/nvEJf8/hKCCkSY7HnJ
fS4Dz0yOYLin83qjpzGljh3cHNK0/F8ifRsoawzBE1drGxFX0l+RqPx2IS6mzs9i
E+stKSwH02qNp0P5arJZpCWf0QgfvNgFNuz1qJshHv5VXcsakSUtu1Pz+Ni6+4zm
MJrBDJlaL0qE6VDb/jXKECWRjg4cY/oq1vyNRcEoWQZu4+hxxV/BXMP11o3iqQQD
GUq81MIewexywMBDs6GakZbFbsSlysXy/V2eeqHW//mRuLSdcVx8dVzzXUeMWQ8a
Dz/Im8pq3RWn0f1rgCSbXAl1swVkqa56mtCGVYm7cHSqXgCfvdH4EExv+p4FrYBo
hDAt6YRohcZvck6bJ7j8As32nI6KfmAt5D16qxBH20qAYTzFzALxhfp/fguteS0m
tjOijnVBj1AJBlzSXo+Hfu5sMUxO04MoUGVieyOy46p9W/XtoKjmUSKs0zUtCLQ2
r54EiCZhme5v9CueVFLiDmLXc/jkt35Xfp092K88A5V7lBrNFs9Gv40vsDc/K/YS
si1UABGm1gPy93Opt4TcCnDUXTGK/IqgPXFfvHTrxhuBhT+75+CUBe9fTnJhly+C
o8j3fLFHeupnqmj8+BTDhYa9vDKDwOBoVWZRnp15WqqxtAvOngskDomkDjyhv2sZ
vN94jPxCv5HeO43nt0cQScjd5YqfRSUUmH4ID7d3VmP5pnYLBBPu2ney2nVaHebF
gb8ext9/hLTxD2/mbG/XNUyyPEwPjVMmmEFXn9sSqYA3fPT9tCu8zojwGJZzMBIq
RZ6LCrRMoRP9MHYzmPYyI5tnlEg6Wo8vQdv9GRosUP+XNAfFO1/1a+iAGfWNtq4V
ymit4hDZJHOx3wE5iSPfNZvOhCURNI+STqxC2pxHnGkBdIzr7/5v8/JWKBJy1ADN
zFiEQ8nO/Jc4NUBfaD+I7m+QhRTeyjz9Wydc3mhPHJM47ZGNXNTPUonLn7+UC4lb
2mBaH5P9RMA5o1yeRqS2JBtI25NUJ8waQhRADSBYS/4wWDeq1vh0EN5V/J9qWY/c
2LJAGrPl+8ReYGH9Swp/294iSwXKp1i4LFA8ZXz0YVx7AAlGzaS07XcqEAWrAQuz
P+zAns5hhmIPiwBxc/PgZJqkWjcjm9RWZrRBSMMdSVcv/WMvDV0FoXCd3vajWcMH
lv1MNylDqJCKyysaATDzzuZaXOo9czw5uepXMnQ4qVILDazVFMda0zputIG+nwnL
fCIQlw1NahTQmc1HGxzj+ttZfTDpATDv7UAXu2SHMEsgSNWMXARKlXPPvy51jGfC
HKXYMDWdQGIf9QdTLw7RamLaVoHI2X7cZ+SMKeihHlwalDfCOdtY3LMAAZUKCceW
UMApLPAeKnALHthArSgrvdOKdb1AiQCKxMsK96b3yJrSgOoyKUsTJ0Ihzr+4FW2c
Zt3KwWZ/pGsZ647Bf/rz12k1QBpHvRrdkC3uu8KZO0w+9qyc7/liK4GjHJvwywq/
nJDEB1cBBBZDmCmuWEXOgOD/nb+pMJBqdyIrO+g0nqOEElNOFjpSm+XZ9xewgLxL
jaSCMrtxBFwfKVLPndlW+IqIviazDtK0RBFarcB7opoZ4WEkiytfcFC2huyhbZ/3
d6BIRQjkk01zklMhr2HDlp41v0s7oa9hOlC12AwH0BGKWzXVUpJczetEt6wgxZ05
ms6NH9Xr1LRPGnTmdryC8TLEG0h+guiZ95qVh4Ao8qxPlDGFA6R8hWfB0lz4InOS
0/dPlXDB9ABURyZ6x7RkuaSUn0i30ja90RlS6XuAxEOmUJmFZlhOWWoi347cNKTh
wwX1M91BRKHn8LEyOUI5Tcc11O7fvYX4bBhE2zEHoTw+Q2KedIJuOc8pW3kJNrYI
PcKJnAvjhfSPRqoH64Scl06Xb9QKaL83jeDn8RGPIGvLaeJySqq7sscnMYb9uNkm
N7qS4Z00Y46Qs9NQi0N2Hmt2lWiWTWk2o1cSe6V4Vcv6aif9Vnnv3ZhVb+GaH5Tw
jzMgqVgCFwvc7HlNghFCgW/L8x4qlploW4UW7ndyCBPdEtGCaLzXQHozEldYeBcG
dPLeQJLn15CJxNkZFm65/nE2AjDcNrDbUd71IM/iBMPDthpP2ODGu027ni0nvBYG
A6qGtTrCEXEIKwx7Bo886vAb67r1c7RiQz81l9eqJqR850mmhH8BOVRHnYk4OoLF
2o1k5n6cMkUh2KU90Ho3IASlvmWx+mZmtOF0pZpmtZ4XIJss4ZlalvYl0cWCBFaD
b5LftcVYMHAmRz1KxBQpIf5pWsNMffmH0v6GEUKouMrm5EYNt6STlhM/oTmdU8CB
5bImKBlAya7bEyGrqSBvcQ3MO97PxOhlq+L0xM6TvR25txphe1bjQNn/ae41A3E6
trKuO0El9XsiFLS8Le1A09WOuqNIyM2PYMzvuTbTN3c9jsqBi/9cLFM+T79oNwpC
feHq8w2BJof77XSTAdCIWigKsz24qepLNUA5klc8Rj/V7J1wIYvUJR2nHgrp9ygS
mPCalwNqPvIFdTJCWFgX0rQlF5YaboahhdFYQd1vGPP3Oo8N5Hm34hLpuqQ5z8sp
xRVg9cbd/BqLn1z4JS0mpRVIKvyWP/aLBw+7jSCLhdt3v0peoLQx5uDHZhbv+mMN
Sd/G+vhn9lzt2VF+S7t9PyW1GCzOWPHFWCi/i6L5ubohDrHywc4w+h+hsU2c/68z
SAW1A+ptyVWW6TPnZnVbiePeJN28FwplpzYj/atJpS/InClSh8LQOgbC0uMCqtSP
LnkNp0htn0qcudIu/k8loVl53uuDTFRwitooxIXGaBjlyzf/7YHjnzV3qoni/QqA
WVlmjlTyp3rRLVQg4HNpenTxvePa6ELDunIGO45Xc+3Jd61Vwt2XaGgdfsKQnIye
puMBtZt0CaeJidNO02o6meY98v1en5mBvZm2X+rQsCZOaVB51ghqn8iy/1VctEY3
WRZGlOCQZR7M5yb0pMRMZiNToObSNV0F9BDFXRrUKeIaFVM+eIrBCMaopFhhvdNg
ucDhQ1KDMOaPtOpTVcL7hqoSUdHCSWDZsKiT2fG7Bvk9dimHHc1ow5ewR//Vnc9T
VK0w8v/M26HGTIVDeXI59hGXwYtQAtj0VHSz4iLQC/F9Mb4crmiZwaZlGW6vDNt5
/+ew66c3HoedTvRTz1sMYMSJ8IHgdqjTVM4m36wpigUt+PD/gxcn1bv/zKMUV0il
A4unstwjna4dejXEcFQh/8jiqxcwb7oDde5xM73r0l5FJQdHpuk6pBUKsgz5Kmwi
5x7ibT9q96z0GYLOyhe9J2c2oFqLF7D+5mPyxdcQCG+faIokhcXAB7N3TyHeENx/
DYWKqr6QqSyFx4iW1h9wY4pP+y3RiOo4rJVTSAX3EjMVtjLPv75w6Mjy3JjOX9PJ
gBA6S/Oz+ukVY+ztvOCkwlQXhL4i715Wneigh7PhgCuROaspm1ryiKdhfvKkLave
rLeTWdSCPwJvPV4+L27vMbDnYUJIXWoXw0KNpsuFBKX+TJBZk3v+qn9wX6M5OE1x
Vl+uKSW/jHoqguvDhjahOfjmHf/sMS2DJPg/WjJQPkhBR1VU11zV5u5PjfNFnkBN
Yggess/iy3HWg1ZHlAaAKuuVbsQmtn7CgXQIIrYPCn7Car7ywoIoJPGrx1h6Z/4R
/huesdLeobEPDSzetx3DRXEPIBDJTcsUOX86sn1Qm/5yJzFcMvaeAfLjUMwxgC1d
pbnLPoEYj1X0JlFCSZWm65ZYMP3vCtQrmEq6u6o6c6ZrKaOrzqw55FRn+aIaaPOe
C/dDAH9W+Pv0AY5H+tIF0fP3X0rWhBt05+ZTqM9Uf8poQEHaSbVOaL6Oa7iSgiOe
oZ5kMGZI3lSaBEA9H753BWIH1XQr/nzHdsKWyf+tE8oexzTGfM8S5suOKAHCHKmn
EUTvFERZwN7nQwO3qpnDkn6YkN90Inb88J3f0bKeb5bjmiJ5tN/0RzfWKmdI2SNS
7Mb4NCZAF8t5KZnM39N0Jg+22IEqVFV7hmMOkM/qwe9xXuzHlkGDAfz6D0xvPO7E
cD4iw/mrJdP65xFqCdqzaJW0bTSi7/RW9E+W4rm4eKVztDUiuc2Ax7KSSqARf2BV
CGsjYU9hBky3iCNw0koOOeXdCCBoWyQNoyfnjaaTK29yxEU5SHHM0n0/KLb3+Kcl
p7PoI9gY+M31Dlbzva2+HTr2MWnjfT/4Jh+fQM2BUXT+CwGCJKmmOta6hiXeQtuN
xVX4/REDZmEha3qLiEiP/hV/Rt1jIngbuT2xaoq5incW9XCm1fRCPbZZG4JNW4ky
VZ0cF5nOI5BeNZ37znC19ZW+uldQurw1Lg5wePqpIuwPMD4ShPm/JddEC1kn/dbi
EkE0XaNpV8xVj90WW5oaxeagAEqJ37VxiqG2xWqlWZjkXUGDNS++KGqto7/u7/6p
iniKWVPjbNZKZNtLynIHQjimCuwojozXRPr6gus7Fr7IyXvhK9Ggb1V4Tw81rjz1
wJXo0+wrGy9TG0nR20utQf/SjpohSS0ETEaZFF5WgchRFr8xA2Xl8cGseT5bawqc
Xp2CJdGFw66rSRG50vCvkgW7xNAbkIVXkxNjXxAhFXXiGdxggcqempEXLv4b479k
8424omWM232rncLVw/MfEgG3RpzqGWaKJB97p14TE5fMEesxNpsFPEQuwe/8/7th
TjSuNofLuZMgWWKribiuHHqnHoi5fvDkw/Lt3XoEfQGpJ4qzkewhNfA5WdUtczXJ
tqC+1mCj7kXdcm27fu8SwLbQ+dfNA4S6spgsi1mF4kPGX2wqB94im+1SPd03Yfyf
URU/Hhhm0MyHefZa5ALLrHiGUZWAtr8YUJzH9O3sXIGr9PUDusn4fUBzdad5c/vq
aqxGjHXSbuvEP6eaKmfkLSphubZuEVuaSKojqKZhKkqrfXJAfrQOuP7HCy+7P2zB
t5dB9WWTY1qS/dtYXsVFCQiPuIfI2YfLfyGE4PBKvMhD5eThOQhVPEjjSToS1zZS
BQ4EtFh8lQsqzcYKwTcID23/TpqA+7NZ3R//2IZnzK0TmC7LtiSqGwsNlUrT5Kxf
6ITPhwDabyG9I8HINDsYwVRHcDLSDvLcKgClhY9f/iuxTUqzNfIIamQy/V9PDw1f
KEzGw+osIByeBn+8N5u+dtvTsuaNXR2LZq3vgWYc9y1sIzZ2lt7c6QFRfwE87ZHs
6EGvRZSM4Phqa4MD6rcOI3aIOPpuC7g4Rae7AGORRIyTcEoYZdLM1EfweNGY45V/
R1H+L+LIwXQqo/PY/Sia0XW5zMqNITvE1hI5etGbJORtViyIcIaxz9EeYKA9r3Ot
6gTxExVsotHkFs5zMch3A+RjWgKuAcvhgtFDGQ3kjs2l+PGVTUn8kv09+BaoKWqg
7/8yP2RJmKXXEkBUVeXMNerks7aabE8R0Mur9t/DZD2Nb+hQKy1ID2HYpHyyJdml
kW5kaoER+cxs1iThhjca7B9CdypD3Lie5eJNZ3/L4pqkxbCpOq8W741mbg2lu+h0
xnxI5ZEqY4+UK9jmZ/nlGE4/4s3BZtB76b4nKe9c/H36grDfjTnHjK7l+GWsVRtD
40Q6qqNeUgukHMmvn7fomSa1GcGznkWBefmuGJMY/PoZwTSyv8NZOlCQ0tm2//1b
EzJvhnIMp5Ulq6EGCGSJpfBQQbBmmIsKAlSHfVsS9W06NgrmbFJPpKBLsxenGGSs
ztQDLAYrH4N4kCMDzVSer8KPGRPArJnsBC6CNyhCFPsEv2rG1PCrE61nekBTmgeB
Mvze2Lr4GoBXsYPsA/m6LRlHx9nXs77al6o6fynpnx93rEgljxrc6zhrCV8XYJ0Q
fmdUxQ0ISABLk7xdIj7JLvxrzAPZjN/Ei2h0eS+qjZgRjvrukZHV8aMRlBRg2x7P
Dk31e/O0LqhQaR2rnNafCCVL4DSO8VLl9YqAySpzJgovDbIered5eqPKx1Vk2w8h
vgtvtmIfdtpAhRBZFpFsdnti9QNcizhT6OOp+DqZnRR0WfuaeLZtlyJ5vfVquW7S
Edmx6JuRzYj/rHlJScRsmMqqAEP336w84y7r9wJtcJ+1xCqE1+vyjAI2UDTpTF2l
t4a66QBsrqjd9SoC8PMm789jztEIF9wOtPM4UMpJrJcEjo1/ducXoC9qR5lz0+ye
XT3IQMec51QACvRsY4WT1ezy9/UR49e8rWw6bGirOqBBLAetntii86l2fY4+ZlvY
CKEX+NkOykVF0fywuqKsso10iciR95fUx+A7u6atneNdvOeul6vuc6P6cJssjJuX
U1Q79ofS+ZoC5CcKBilbDBQPecGKgUsg1qLDiA2MJBT6w4l4BLMB2T5+ymQipH1a
YDoNXWcrLYngc+gXbgpPwgg2IbGx5I1JrbggjS2RjWsX3mLB5GHCxbR5I0VgBNSm
vPmALhHF0kuicYt55gdxuu4fdWprIHzIvsqNMLGLUUt59ecNJVvsYj4rLGIX4PK2
peJAYdgP4RXILab5ZLtlINkgfzAM/mB/A4NB4lHE2rsLtCxS5+TBbRTxLYe2jhB/
nFbY4iLEbtK8fShGxkkBsEE0lE9XLjkFhC6NEl406DLN8nuGeuX/M9AdSIhc/KTW
0q6Uh2EYXJZZ2xDD2YoNCPrKnZqM9PbWeUbFpAp3QU+xjhBrUtD3odMc+si9aad2
xY9mGMvOntCWbx9s1BiRUilWwEoZaekJQHUZIc/J+BEnjY4zTgJrq2YxBjzL21Ri
/wkLe9vDC2Bbusugl07ruB1BB5oN10VBqNIAI0Ycff8UZAWcM+CsNPDPa0obX1ub
7LGYuZe7gqnbxNZMJigrlEAqREdRi+yPzKURe9HaoxsQRF4dZJMBB55sUipNmhBH
K5laEyyHU3C0ufJWFf0sfx5tSZnDGA/LqLRRAGbXknoFS+UqXBw09hO1npWW091o
ilq9MnvUw5U8xNbRhpbwW+4K09CY6Bb44bvymPmCvWaqjnGKn3+vD37yIsmF2lSD
Jeulh890xEhwjNBA8RU/s6QBHEABIg7L86IXE8StHyRFu2rp87/i/m8lesFiasgz
65XTGYfKWkvaI37GBsY9qUUam4KvqdXBu7tIbot3aeszJYVKbCFF6yOfR7jq8H/4
NgrhlTPJioecK/7+lQpwSRvqqmb2x/nfdNr8SS/+/1gzOMHPv/uFeGm9V1fAF2ug
aGQS2LBOxGfOPfua+6Wi+u7y/jN01CABaK26Oxo1/L9pjo3gIwUJhUflMT+qD0cW
y5xWfU3cHiNRD46j3LbkZV7z3StEzgy/BLHD6wQO/dLg1tq31ZTkhkFWoqyDPLJE
SgC4SDLNTW3qC5L7AuVKqXz1u2vQKqdFL0A13G5dgWtEsOtVxm5yj4SFmrRkYPXj
ekUZaHtvxnua0q7Y3q2/DPQL7Xp2BwbaOch2QhAtvzOrrFhtSSURLc72EbnbaxGY
LJ/8VhTs7kqLDk5Mio/zdAdL5cHh/KhYR5PiLGqK1Tf/P3cwf8YHL76t0I9kkbIo
3GgeBmEtw1kvg6Xck6bPmxrNKzu/7fgUMnCuXQCu09PUcEHHvYyVkbWPBLRHXUfe
LdeibkXMREPrvhX7F+5jNPYZinHPF0ZDygai7fwAuYEMpt3i9F/R1AKpNnhpJAj/
y/b8PQmXYHuc3GRy+afz9wyU74yf/GvJomnuTvOSUVw/CGPv3UAbFTwkl94Zu81e
fholWTK2AVmBxp6aySmEo/AcE9J61RRFRSAf3RLe2U36qdlvbqYCbpSyCSxBYM/z
KgqPxfGfvHLePYBJvWkPJgeNr36nSCrNaQ7OFW0NTODYhhdX/gqKtPGB1b+H0Cqf
43AS6ZxMayqgxmvXug7Az3GIhIpvISyd2IL8VL0ZugHyY9a4MMsJADCNnXTTLpgU
HU+3Dh8zkaAxQOs+ntrTnjGSBvtNN/cCGysEy6r1R9y2DEobkB+nQzf3WldyXMIW
t+k2FziZxkB723XV6A23hcxCfB93bFGP9JpDAp6Ef9WehUE0G/bQladet/zy1Vi7
cGn2x2v5m2f2v2GJ54rUZOpDC+qRo8rmq+N1t6D5nIEbRylYa1VjIcXjl8PtNPfR
BJRUx6yKCKPMKOW82UNtz/x1k5q4Wv6h+OkBuLcLb8fV4Cc47rpqwLTjKLBYS0HK
HmA4+eDHYV2Q2yXWzoolLPfUVC7GjHyHoxXH3uIGyG+448M/CEsc2yKqyDP+xzW3
PXaQHD7E2a511eNSOwW5K+65OC4vNelZWtmFH/qHQr/5xzRH3PdvF4pnX0YHcLqY
fWjzADEaVy0iTGNAaxXJeuSOs6eMVjVGPBPvhcaL9vReqJIW12119FwWpXv1TDk4
Csfx3J0SfNt6Zhm5aK0HhaammnGnHPYWlJYVWphr72wmQ1s/E7SjibhkFipZjmrB
52sFR7Jh+IWFhCXNGMV9AEcWeOCa1dH2UbZhMdN+0dAeKCXQfidDC8R/4cm4V3zr
QqIopLhzn7r1Zh3dHHjWY79BTzT/OuZFSxB4QQfsNppUzT3TbGNjM+9lcFZncoYG
70ZutyY9J8eknj0+iN9SbSy+gpFGbYO/Wjmj/vZhhqMII5DzjKcQC+s6KWhx7ZaN
Bsavh/Rg7oDMFrl5VBpj/Zq0bLSlrLgQvRzbyJ88Lrro0nekJt+zLBaeB15NqY3E
sib96P68ZkFwA4ImH0WZP/sMMfzPRZHJ62N9YWHLAqmJ9ig1rwj/LFgfw5JloDi0
YEf3uNjomwvtVOzyUMUo5ySHQZFQi0lrsK+qaeT3Oka60zz8r2p/YXFjswrxjXwb
l4GNaHb7sadQEt9FCONOq/IE0aTlO3pneHvB3BSue65vYV6GYvi6E1snuFZlI6Wk
2eoMKPvgoc6JcN0qFYEvBv/Ueh6Pl0HMLXa1gkMPTD3YbkfnOfhSfIUZA17QiG26
kZpUqIAqXk91yRFFAdqW6oLgrMyUm3NeHey7s7f5iJegShdAzmy2V5Wf/nqRZ/87
C4F2uJB6ijXbyg6pvZ+nJxO9jB6uxM/dBayJ7sOf6tOtHU3rR4x2smG6dGZ1ttMY
/rvfUgMwjEB3cnjg7Pg5rYnxqFOTAa2SHxhGX0zoO6ONgiG8jr3zEVJjSBycBtGY
TIBTsQ/Cv9nWPkNzMpb0DnBpolL67sktxP3HiavM8YZ+Nm8JwgXwE7k4lVrN07b3
d4WHj07QJXzS7SKjKjRh07ujBf45AvEgT8X32k5gAPaxR6MfXSSE9DzBmwHeAlZr
lTrxz72gHJvgK68elKnLTNp7+L/aosp5X1WLYiN/M7Hkr4rRY4D4yEdPEldEJEWl
hLvtAJlH57MNEyAG6xKwvmoqdzIDkS4h/uxOWU1FZ+ymgiS6J7L4Y64soO5S7oAW
FO65TjAL31o40ax3yAYzgcujU+0d34xHQQliASLI14cOTXvmU+29RZ5j+znKSfNo
T7IoAydeyZN3rLWaU4pb0Wzpb0q+M5k3TsOCzUNDTUS98W3RdDAgT01wOTzwzLpR
X+bYG9SRTkYv0s4SZHFZdYxGsVaYFum7gK2N+6pH5gWFlN7RT4pxjgD4YQ00rmvA
so8vvuUAXFG2crFb6kSc09Ne90Reg5bjW3vmAjCfc7c9NS7ZgdswU7sdZtPTefPo
+dNtnKi4eD6eoSQVkF96lQBnA4D0U9am7tDdeDi8UoRAyvBHCgO/g9bZiMjVg3lU
oRGcYTPDVsJoeduWCUkBpvBa6W+ly186DlCEhVYB7QHfEeYn/LOrKTS4OeFmPzaR
+/Qhikw5UtG58D8ooMw0IYwcI6z/Pf0QuoHxUaX2wRHTYVwrkvFwFNqokOG4CQLJ
xeLj0uhJa0LVeqQ/Q/DGmnkwrPtc2RwZH5iX7MKixHrTql8v8eUzaFrxI+0A98zI
H1mnGwG8YMlPS9ZIJfGycWjuyWMQCRII6JxLg61f/qA1+9ddZhU6hf2VUApE3/J9
U8IKYUxSlHtaiIbFGqoGq63tb21OrvRs3bVMgH5nhUBagyAx1+AxJqwCHfIxe+E/
lByyyS0qdc+xMsI43uKjvwGDYlPrHXyxELszh/qBPSlJlM0gJATkxQLGxJM+8sEY
Eqa8zrbsf2tjuY3HgxrRd3mBfJf+l+M7xjhihIn7h2Cum9Mt2qbp7Ts2YqIf5TI+
LD0KELSY6AFHrylGU9s1JctwPV3m4CKPbP5BiUIdREJn/pwaXznZ4QpXNDRAdY7X
jt39X1h2eElJ+zQMpxJYTfsHjYuBn5WBiT7KmnaMrGOmowBAtjwDiEq9GpMnXcPi
EBMiYdamoHjPC8P3no4L9ReOVhwd0xpdJH0tnkIFbAghDt0clcUl6O8rKiLXbk4U
XbJeee0Cyeky/QUoY7plyZ++5SMtddW1NjMrb7v7vU3W9QbDuhMJoN88oIG6Xq/n
76p5op/B09FZJAGeNajwxnmf8DmXoSt8NyvDK45qx5xm2MbQsl8bVy5zQKSIsZrd
b7KfGytK9cOrIb+HIWxZ0rXQgMrDpx0dbIcmVc1cU2DePlOQKIz1WHMkAw7h7eFz
8kluL+3S9Py0Us+cksFkJtVcCNlJ4v2zS3E/IfLSOrlcLmBkO1nrecxLdSNUbyra
nVq5tc8ZovEGlPdzjVKNUJnFbdtLOABjBvBM6t+exwXTz2w+FqrfIMSliKGUT/u0
xUgXDLJcg1hvqWiuWmG7T54HQkZ6wK8CpEpGw+fJPT7RdYDa6+zwJ+9usxL+g8Vv
d0D7ws8e7RJj2vW5EaEqv5wGVVHMcrooGNaN4vZgrOd62yfAgPcXksYeftcLOy/y
yQ6qOhtB+k9C2XI2sUX6JWy5SM8aLDjnoPNXhdJrRFnT8X6hH+WN6sxGKyaXfwU6
oAXXuIfgPly1VCnakULYfBVQwQ6Cy4bY/Ufpe3RIcsw3JHLMJpgpCUy/9kSL0QK8
YbIUvJ8nCLbYEIZpKQpo/zuIit5u1SH8N655cimVBdRNRZlFvWvQK6TZkv9fgbVf
mw41CTqoSCyz8e9x4zx4L5037BTnFOGxjfl00Yr1Oqw6qBFQsnUeylVGreTkZN+e
YRDwutbW0mcFmjuD9LxNYk4LKzQrHVwRjjrK3k9pqYBtziEzD/P3lpoeB/ZBCpta
dbvYjXT5jk5TAgSwsCvys2j28O7NSt17/Tp5tA9K/cMETKpbtS6/pR7BaIaZCcs3
Qt0qZdlVrpADl5nYMNJKwfVUUHmmbJp9943pWhyqR1kL9b8mLXYarOVYoy/QckpG
azzCkIbhAcu/wTrL8ikMQZpZTWOhn9pO7ilxnDtE3xmnTpoBaxbtCDe9TE7XYwXJ
pFLqMgMYGc3nx1M8m0yo1WFTotNNNHFkc7pnPT/vEUodQUHQqritrKHp3ZeuiWvP
1t4HfnJ+UG8J0yLfFSoDJ1ogwJN4OxLhDITceZjMSrJJAaDM7InVIXgtbJ+uIhud
GspIPVYzI6unbsUT4aD/NJxHI95MiFfevyCvpNdzPXOWGJ8nQXEuhVc/gKxtDgcl
pB/jVeDJlvTXz8ORX4tCwSUfVV90R3ret+5egp/9GzJt1yANwOPmiCtcI3H+t5ao
wAMWGg1uiHOmSwTDIU7QLolqOOxaAwlxqeG+SfFUGeMiaRVdMJP5FRp+2bt+B/tf
lhchgs8+AavsKq0fmwIE6Buaaha8r2I9VK4IReVOiPB4drlddXREQYnZDXv8puJF
t6RUgt07MGxBiszOLsYX08qjKBbqjd+UIcEqEu9RF2F9DcBDcdTBrKB19GfLFre0
bjagjBvD+USEDdMeaMr02l5UsE0Zde3TmluIeywD72qHTYjOwM5or1ZJvZIaW+EL
KPCTd3V/soJQg8AT9m7hhXlnRoXhzYCFU9ojaMt+/gOS3aKhrlhe1XND7QvGst7r
jQ6ReXs1VSOcxIETdkdiAJKviEzWRX7hSscBYfQO0AZ+mxRzhs9q9OsdFAkXi5wv
yImv7uGdvjbycR8uF5A+2FuvWhXsaignYvAZCKtz9Pfk+lPFKG0wO9WL5pFFYxOC
h+gn5Y/gdlCmkC1tns3eIzSyd7SwHO0g/rjZTUnXffDIxSZwq9wfim9ssQ0f1CSU
fXLoS0DtkTCtO+/DKjvPIz9eKHgiLsQfcKUQ264AYfWIUx3xN209ySxgMwJRcl9o
zlo3gUhBBwz30vEYWjopxEIs9dHlaYwhFRiEQbySxMnE+/Q1RBbRyFUrMKMwmFvz
cOmK1HBD2K86FpgOm8s7GiePAnYaNid20LqG+djHQ7qcvNPass483wXUJ6RKD/oE
aymgaLI+b87I2KeMkzeDaWVhAnCFDrSHoPt6k4ichUtdhBMpArG7hSxbJ+z7k5uU
2vrf2ibjXW5Y0wrc8B8GL496sAbVeSOAwYy79MBm+Y7VV16qaxrN7jI6dxG2KxKv
BuviRGJYusghvFP3LdfDxK8VxYhqjrIvzp8Ov2CvxelTBrWrN/L0kcBl4KGC67sr
BXXe0XGfNKoTBu9bxPShq5paM0KgSawCNO5rDgYY+3Z8xKezv/wdZ17MXQkwkW9F
ILVXPDixEYVEkzE5d49oOzY3pSOrlw7Pj5VwOe3dlK44b61WJqUIWm58sScZNB1X
vUOsUudWQLvMPRxXLiONzImuLEsTZfDSYUHr1YknBmWkl90yXZ0K4XcbKCbisjnZ
Cx22UgmSxDGCSgEDN+FzPf1UynRXbA/6e3/6Dh/WoLeSzq3lCeXGNJntMrP8ojh6
ND8+n42dMYm8XJJ8U3Oy5l/dmQFCImbVqUy4zOp0KuW6lhS7Qdlk68VA04V0q92y
n2bJQW3rt5hMrN6VP2LkWS3j/dVOr/qIapiHpzmC7XQLtzKavg5ZC4ymPkahez65
A0CDX6r5iC8DpndFRZqD8sf2L8s3Om4j8eL5T7PJbgObLs8r16yyudvn2OjeQaVJ
lj4NkRphD3q08zJ+YN98rfHlyTdNY9s4YtY9g8pmiCPGM577tq4e/pcAOIBt6J19
9TJsZrhQpy2shzRUJFRTg2Soni7fidjWz4pbrND0r0iM6h+CoIkPK9pUhdd9w3X2
rd7669i/C//xS56VWtERnnbSd3op3+6RmWo+h+sGT/2x31whu/qxFcDsuAtmxzId
94DOOVAxOb1YmHotihHiOdcrlA5Y9ZVqzQ4GmE6+gDH5z738g0ZY/VzmVpHvVrub
bQEPM0TxYSHLy//ITc+bobYuzoSHNapteEPuORv61nH48wxmsvKLoROOeqxsTy0r
0EPR5eP1B1LCX5s8DLIgLUx4rMpsbrJkiX/UaZ0MHqYejijPFWbxLqp3D89q0hhu
YEdohlCx5Tb8xoSpqVx0kkQtMFFSNSPhTc/psju004v+hFAxPKxhEcHJhAjufJjY
LT/AszztO4bsGeUnRpSWWbyb6A9/Sn0R9SxQt1BXKb5ovVB4FdI1R8+7eBSamFGJ
m2cDnMa8SbMl4dD0XSBBQKj10Vvl4m7oHqSr3D4VPhgf6hsJq+NnvzYj04c/so2F
oEep3vb6ZQUAbr3617WEI0hni0xD5jWKcZUh30rg8GNLSBxI7qmUP5ohGAPJZW7D
2zIPCyScaePBuWVyDDvtu+H8WiZgnECEDw7SOLiemCZveRPZcYVXb6FTuqtsRlOJ
G/uvluTfHowS0OZmqu1ayE6sYc8uW+bSYJKL/dAlQW9EwntZ7Z/B62ZJ1C1933gO
goVTKmN+xvmtfuO2rFsygTeigyOuL9O4g8cIYbYGicLRU4tX4tQfn18uGnft3vAZ
FIwWduQ+2708Y9BAd50oRJfEP22qfvgmJjt8EC+jZoTO/iQTKnrO1KMtHeaNlUX2
+kZvXOVDP6ezSR3BFTDz20hZYc9XNE2HPFb9iOJLPZtLMSJcnQgZDQxl00/ncA/y
VxSPVef+Yf8iIernuCDWRANifJ0NoKcsaVtSz5Dv/ycL/DMbYaTSTyncsbetGQ9B
Ub7SDbvQnDks/fJUTcHCHmXjF8nf8b2Gp01/L7AWt5w+AqSG4kzC6r6WzmEoWsRA
hwkuVFpHH+gZOLVi9wLsGpAohnrQ/2babYadFc3I7uMnvT5WE2Bwsf3QM+lx3jW5
c8NQskJ9hBsxMsZgipucrYiIBFDyyPNmxd+4a7vaPXS2GgLP0F9CyNhvzAh13aoK
evfnfaBMCEMi/bi+icUxdzX1nM1ifuDX7GrKErlzgvJKbCNM+F94tUxxTIWH7eqN
u6P/JkxBOLfRhleRDjlenrDuMER86pd+x+EjR4WbLmiNCr6kH4iJlBb6TFBr3p1f
g4VN1iAj1bSmkVZRMyMCVX/3BuA+8aDBktRDlwkJ6Kk4VnGafRannDeyCgCojhvl
h50CsRqSoOkFUM7kTkZhjFMNpcOf8tHEnJh5fDGNsYU7FK+JIwGc9FZkKXGoK5pM
siU4Bby2P3dX/1GhUoNWLif+H9XVoBgK/tO/sVbvbc6NDib3tBGCgS8FZTqEdSQs
QsT9zLiP3VQ7+QS7Y1oJmohyHCAXD6ZUq/ZGlSNuP1vLoeiMS5OOuiT71N5GB+9R
oKFQgkCj0zRm+3I6HxhQxq5e0N+BJSSpr4awUG+dTdr8mHaMBZtpyu+HO1bSHyUZ
M5SJH1pX3dSOIChA4FJtnm2JbPdD3GnSnbyThc7H+tvsMq5URgpDylV2gRc2sjDS
Ys3ZlDEd0D1F1JcKyRPKkToIz9c5e9kfmzUaVKd3w1lbD0692kVh8echV1hj5c7X
7K22RtZdfhiQJdB5qcYjO0hOFNqef/9mYOKJnMPcK/zKdcx0f7TXx4VUJCxE5aOO
s7PQxU/U6/sjD/3s/X5d5FMqcEzrmep7toDvBubvcHM4GWiE/WIrrRUzZvZ8XrwW
69eMJ5FRPhiiyWJpZB8gccXVJmqLQvd+bO1j/cXLXY4yIPf2QWBshU0I6RSc6oPb
sIP4T8PJ4EL9llmbZNEsOyYnHGJv4W3K5ovFz1DRzwKbDV5tINPqGL9fuJNVJkxc
M5EufTEwrFDGXbZF01tHVTngTR8JJxt0t8JZN2ZuEsxwvGAXNAm/tWrmWKJ17T4L
NVkaeV3mFYk/1H890/opfGJo2l3wvxgdtpwf1cYDiSqSWThi/g0i9eljfd19rNZc
zeH0sbt8eVF55ojjHhV/v9ysr7SHuOoRH6RPlH8ccgtAU5ZYt4Tvtm8zGCsQo2Nd
qOqjw94aHVzuqOCaVSUQMTKIXUMlxY9ZU6YnpSCjWUNkH+a1ejs7cK4yiozu1NQr
MZvZadHhfPo8WRE8R1HWMItb2ELpsLm7NoRx8/s9BJ7d79dcDc4Z+F5FG0hfZCyS
Wjfy4/7EbS+PsrIzwBF7MzwoHTBtvi5JuUPe0hAZEKKGEcOUcRKbQ0WTxxdDpzo3
7B1kuC/e5KzBPx+4BrK0jCXiblDWYCrdJAjZgt0x/HHbQCVtn2WoY55shyuhf9gW
scYJmr46PHQYOdt/gRzx7kkiBjL1KQwRNkI9Os/HRtC4utb228R8apt5hsl9fr7J
U2oYb6IHK++cuqCb0R5sb5GsnOy1XKnW89+bcFr6MKTAQJ1Yu/ua3jAxmCSkL1El
WaPiOSI91awjpMXkCo08TjEhf7EReH7QKt+wLuV/+O3prmzvGB7NjnFNU+9/Qu45
ORya52ZktHR09Pop4+s3s/pC3vJQUGJrTHN0b7CvH4Dd7swGkAUmAxaIv644hnw3
F+y2BJWZmEl0Dau7uKMLnt7/TzuoUkpgL+RFjyIl2vEt3Gaic+CWfH9i80/M9hVF
+T04GpuVfYW876UAeXEzilB3yrO2GZ8oFhuXklq8L4yCLSc9lf1ag57bZL9SVr88
ofHVb7k8P3Te3dLlEyAmgKWRDzvZiIUQRGjJF6INnCDXeUiXRr4Dlv/GGusZ+1tc
wzA8SDfk6HETWMHWRrWHBd52K1Ctw1hSsWl7uB0uxUkTPTLToF3r2RO1PvLS4l6H
0Mj4WRT2IK3YT7BQsCtKMx5NRPemTMMbd7Y36gq64xUtbgil0evFAQiW4hes7vCb
aBsWlHZs+GywI6bO54Xl940A8ymxWso3m2xupDVy4hktjkBAn6HbZQUqj3Nf+Pyf
DCeeyVIo1TwGj6HK01XbrxAjmMfXkHK8JSgHQ8mfPRb8KIqpErYW1IZOL2Lk60o0
dXRHg3avc7cAbUc+VEVvar5PvekR6ggpTwOiyfXSYetGovsw6xPHklnwgXKckIrL
7zUx+B7NGjbGv13413IrF5d58mFzrRZ7oYLnVGs9HfD9nuc6MR7I5T1Ru9KDqw80
P2K8S6X8CsgMQz3m778HskeDicitccEVWnC/xPHKEEJJoeX7DZMHxnyUwSQrPW4G
AldpsOdk80r5p7VlTHGq3YVxvMBwjuFXyrCTyojvS3eOlr8HrjnXx4PqYTXK3Bpv
b723bLwgmhj5+KQzJWO02/OjHw9sViX3TrafVO7HJy8MCHwMZ+CVcueINHx5B6/s
riKy82dVWXHxmCX4ikbqj4ycEQB/fftp7beHKHzdPVjstsOspu4oyzH91Lq3nbXG
qLuSb+SIEMxKKhMTzA74QunJv4d2fzdDWGEHailTv31Rap555oRxRvg2umGiDMvY
ciXYvW+lfbXOHSWhYYd/jUl2KUvHBdtAxYS3jhtI4T++EZFAJ/2IiUU/77CskPlL
O2fEuK6fILsenPHRbqgq8DwHmgV+1QOwETxDQJA4UYOrwVulWtqJtn8S96R+T4tw
qGMiIwRevWA9d3CONdHfDAL4Y98eSA03/HRs8U6G5lFiUGWQHwtK3AVvoHieplRh
NsGhYr9Ndn/xZj1BvWoNfV04zGA1mAKEZgfWWLxXtF1qf2SE2gcamwrFBm42GCzZ
AEhPjUqt+8SEYuujvvOTC+Lp6dYq7kyeVuSvo6otqMqw479JITkTSNfTZX2VyIS2
xs1EexWR+lsPH/SfbERnO+i24xikOrFXOnjynXl5K+5SPvCMLVlAaweX+MV1CZv6
gd0IgF/LXPCMxINLKARcG8sT6+hN/7XD6NkZAytXENAQ6GiF/H1yzH7zYUNeJzjk
UOw0fO0i4zMw//JZPYxgppd9tO532sppYnaswgnwUUyflE/gOHurg0z2Mwf+tuaA
pxtr2zKjw15bwYwQdm0MjePHe0SPqCQQVttEdtxOH2xkDPH3etLo9nIXIHnbXwmm
xnKOQqCghxoK2s9s9jlDmYMjJeFPB5MoCOFezlbQk17BJv7Sjk1oX/Bul4XRWEXd
4rvkhLrAFQMw6+GrHeViCQ66zo3pZJoOYSp/08nky7bwRPXyGhh+ngbR9NvkWJpN
K1e08GuVMXNiyOywLzNW2eLCd1q0YdwZUVvG0wk3pnbEzeMnf0dqE79QRRLY8saB
cONpA4mhAR11QhdCsqfOD9LlkhmwfkcqBmAQ+DGA8LQBmFBsVCT+sF/DlI5oZQnF
cNVcSOBXekeXED9T2uEZuYGWVoLznwrYv4ZXZ/HbfOVlwCaMxUFLOb3Cb9iTGdES
quYweHEWCXkWqy3s0TjLIUt+3szK9xCQzg3DmISVJVblWP1wGspbIQLRfqGz2nuE
3+gu9FT6cbbuzxTkdF3zCH+rSiktMn7sWW3mp6lNz1hiMlHKpCxgq6c9rDDYUYU0
12xZdbUayHe325Uzrmca4jG76p5cxJ1f7CMZAwtVFsnVIk6aaPPRxqp4vYlhn9JO
LvnMjGos4HQyjYwterWIcsJG0YRUWEQxbMM/29BJ2FtAC2KwwTzv/FTVeL9rFGt+
s3zcNqnb/C2JegoLH/yom/E9jQQv0EDx2C9cUuO2JuQRdDLrjhOjeop2LZh9cYoJ
KVthUdrb0Fhx1eDnl8wbR/1qxyHpYqJB6d0iZZX0pxVgIw9xqhGoh8V0DSAU2rxS
aH2Y9WlZr2VQhHH/0lXSGmFZVIaq6qNWfBhgbq6tm0upm4s0BJKJOZdUYMbLQuL2
TMD0jy++bRUAwOboMwi0mJT+W+0IKnwAg2BPLGVzrmP9dFD5I/Z4THHfUB+zm8bt
9hTZ886dbSAixdJwDV3LciMhrY/z7jVs83pFjrClOhc/sBNcTnjj8bUW16hgNNYa
2HVAW2Ky+BaUNOm3NMnpIgG/WEX1sCwptK5fXJ3MTysOFe81Kbm515tcMXZUska+
OiY8BTqWfuf51L2xhB6vFFi93chtQZP8mW/uoqC62i1t3mI/FWCmz5phANWXHJop
fC/RLfKVjblYTU0z8Aj++T/NDsEzuacjJ56Nfc/65DKyhZM+MQIEtbiX/fIUmwpX
p/2Gk1yoLqeWd6YKZx6DIsqh5RAqil6FCaFUXrsksitiVGhdfjwDmilKKZZD5EmY
kKa7IPr8ECNDi0HysAgTfqFO7+4gIU88W4hrNwGRTbhf/hP1VWN2wYP2s9QYrpKZ
uitBhbAIOTQKjQ5ylNQJRlPvOtuIxj73+AvZb7gXblc7bnxtJ3VjyEIedgldLI2q
4+dHTXr7iuIdxjmnxm2Dti5nVmG49P23t+zHv4VfZjeFUIrqBcnCFR55bZ2tvcDj
vqJR7E+yVYAdAc8kb6P7UkjuPOPBgrgw+wP8+dqPobAnE/WS9NNFimDP513325yx
5IXIDinxHbRgxFmtI7gCezalsFNxb+KPEQi7zelkbUN0+QPZyQAbrfyVrUNBba6j
6GRhh8+V3s2+NeB1R73RHFrBfCaxj50a9dWb2S24ssT4Qp4O/znxYndBQHoZTs51
LEcFrd0M5YWSs4S9RzEuhLLyfzHp4FgkDxKECtmpyr1eDd6jZmkKL+V/SkKr/Buw
g2oMAUQigxk/PffV+8ILKtZbCDiGuDXX930GzVqgq/Tpu1giGd8WW+w2pS51Dxyz
D06I+/7amubdoPflrF0qzhgresuzcUFEMjkYM9di4jJmS8cqD6RL/+qL7ILzWQ7k
FvF/g1BCE6XM1u+HvlrgdfU4AriYCC1lGm7GcZ3QGzSrKotivh3OnJnGSqXGg5B8
XHarDTDSKp4ICZfNJf+RJq6h6yyFK/zH4UFI7HFFq8w8EQUsqJjmhJPMneg/dIGY
mL+EwVbEQoq+dv1FaFF3UEDABSgdh1mwDyN3pmJY1lWpOJQm8aFgF4q54/lo8GWC
URv+GszDzXKjW0fnb4nSofkT+g/9tEt6Xqlnv6Y6Se+BYm6p2WCk5H3fSPMSTBpH
Q0lTEe/7bQ2qRvlu2hnpVJb5eGifEfOvR29t01pT4neuXDnJPfGOF2BJW0NfoaJS
eW+hfldkeiaBmV5xw4rmazpRt7OmxHIog6kcAM3jRW9KlCvYEjQtM9IzZR0yCBM7
kdcK97F2bk7tRhwYGVBs1LTZ9sh91MCARUeHEEY2Qqin08g6aQ5W7QFvVmyb2aYx
iDN2ocAWcVsE2hgF2sNg6WeUh81rgZAH0jeRTQBfRKioDLwBhY6DQNJsGf8wVkEX
gRYTAtclpwtXWRZFOfjgA0Pe1wP4Ddy5g0w4ftUdlTQGZRiVVZ6jaajWES6D3sP2
4cOOA4PluzqhdI7OruBsrFPbJ0jtSC6e7Bx8kMk6Kukubg3V2k6T0XyiDFoPvRIb
i2Zs0vdGpAQqKai91fKxz6tqxXfZTQEL9xrcNcckrpaKHVvxn/JT+OGFHEZ+S3/c
IAjtlCLJHK+/jVS1ueL5GGhv6pK/lvGCxjIcOtJmoA/Y0LYw7dbOUiWd4xq93jhR
EaKVK7I6SgTvRFqPV3Y51A//BHqnVa026WuBEJIe4stRcn7mWxoNP2t9e+pEUmxZ
w1zmgB2rMO0GzfVxPCXRF52X0l08VchKuP3ZO6flRDBJcPJY4UflFbJeWp8bEtKD
+ir/QH/yJVrPlshJ/yKs/Rx8Fb2JFL0MnmY5y1GFQQGxr48sbnYrCJokv7s8Mmm4
o8gpZqlHJuIBvMxgbGqWozu8qJZa06llwcmlmi4D4gK/jXEyKs1v96zHaSm/RESW
G1xCA2A1Eo+kC1efvlaoF7WfC86tuOQeQG8mXb9KLHyqG0DxCbY1OnRdxj0IZGc/
L7QGrnu/iNE1MSH0lbjz9wWZfMUHVgVHfNPsWz3mY7oXkY5WVVrpfZq+IpMzgOPP
ghUK8k3ETPS72mA8PZL2qKHpaRNTdefFojXOGZ3ZecVBeLGtPIZ7fWlBeDg4SZSr
SGbm7ty3h/2i0HEien00xlc8MFlOP9GdibTOSrlE51VOwCgh2XHiBNtt8xDtWoob
de29n3KAoc0BViiPpuF4msyU4+MH+VF/ISRHG+ymj+uMuPtQUOXJv6xCwaqE8q+j
AcnURTOVgXcYPNBYNvKX7F/1YOEJ9odl4t/iYdANue2Y1Ltt3sZGDYwPYE+hAC7J
f5NFgYNDDsG++wupe1Hg1tWhLC9iBUB5hY72wKYEPzx+sR+asvqkqTCpvkK088qd
UTniiBaz4FevuoM68OwHQnI3OtZVnjqwA3ua291gPQVyt3GaDlA6zVUp7hK0c7qe
iD0BVvUL+bFN50hsPXaBpJtDLTkF3YbmbqPz+Y/EW6gIm5/+f8TT2sbCqr0lcauT
jfO2ShVMkcdJR+PSpFN3p+i3CPx4b6ozWM2X1XS1plTyX6ax0ce9nWH2uGAoDuVK
XRsBOuxeOcUUeJ4gZUF0xKv/8wVReJL3m3EipclBrtQir6KkZN15EphqcfpIdogs
CzXSgfQ+vUR5fbDerhEfC0lTEWWjS1SNb8Lkfq4xmn6LS+I5NzavKZzE/32Cj+HP
LCAscwyJoEsol9mcbfSNwCiTRE73bvW5FxKb3pkaeMjS3VWGeW+V9MekEbo3TIcc
J+fBw+VGAbC2Yvx/ToibwjzsLW3K4Zl8DLNuqE/3q+w1a1YwoHrpbyjHojOB6bE7
xEoKGWsGcVttlh4Qiqpn112Vmivk+ObglfbWAKnePykKGUuPx31CDVCCteKpRqTy
bU2alV+zWYXpaY9nv7MpEZW1kYcidRR13cJaOcNrO868zt0LOJlyp2tJHkXoExQU
sRlBvIP1l2f10QkQrNXle1n8THAM3pBBdzoGYIl0bYag0pDISyerT+RGZRzzdTZx
NGgKVOEHBjXrctzaXP6w/xG7u5tSKtb5tsgzMuoApaJPbxZmSiqZkk9n0ighsENt
kVKVFQ2JLnUnKcPSA29DTUAewqd6wamTHtaWkkC3xeCY9wU9cKkBDQVRJJF0jZtF
PYM9Q3IcU4FcyQCZX+w244kCoBocnnaVniqAbLdIQMwSZq1xkv0rIyJcw6Tpoxry
xM2wuNEu4rMktTZMsOkwtf8JyQu6S09SYm94X9LO3QcH3ctjAtaVBRct7GcNZJg+
dxWcajuL7NkJRcOd41WVw10pSDu6okmz43gtWlUE1R3XxRhgMNU+omyIwlhIdz52
V/RJv9KKqxz863kafMNHO9JY91u0CUfvPsCt6LP5t+ADjyw8Gg80D10XkZwMneBh
eZpuyaYv2usbcWvSNBT5xvKxdIRiAwpwq0GGj78wUNXM1ZWP2DQ8oQZ/XJT2jlmW
FfnyMsClY5+P4wYAxWkhUu29bP76kk8GrJVr2l3S62QigRwTksK8xVddN0apftki
OhfxYpOH2K50KsnhqzdSs5O6NheWLo4qxA11B5IxH+YeIRBX4l/RYnHSibtARlT5
Ri/YQwrWxe5Lc26prQrWiOkKz0jV7Z/diA+7u+sx0VQot3nvASrUSf7C8B/KqZPT
SDPayl5WTt84Cgr3dTPKVY2O17Jq1IWO9BN9KKEVOItHtdil8YtTP/T/Q9P7SAqx
onC0YA4ja7kMg0TsNyyjMsZH/0/iSuCcyYnWCSbmF8f/7T0aXQc6ZB5vh8Xp4NH3
qLsnnT7UIqESfaBTuK2T4smIoABgQW1X8zgncY0P3ogbSlp2Y6fk3E+WgqJKKr9Z
cS5Bh0gSyA4pveZucyo1RGZLfv3MThHWcVfXH/ud5FRewT3YnyXpiuRBE2E0ajEF
+rMcIW0H0fjwcQqbC8zwHHo+R1uQZuq7DvLiXfSaomm44CHHvAPn50zHYkPHIWd7
Ygh59Ie12XP9w2WnjxkAMzLp1jxY8DGVfIaSiazfz5+DOtcGh+UK6UwZKYb8pMHT
8qLVPQgjSlNsfA8F14dqMYbrTCP1X1nZQEN44nEYAYaGDx6xGCI/c86ClRNuPfvM
fTn69MbOUm1OZfrVcfSU7iTEdritsLcNc+nVOh28ZsFbRN8vOJmHW7g+OK8rRN0n
L6/+fNLQJ9mPOoUSxPNafQO6AFdin+xK6cveb8svePjp6Rocdwd5vxHWX8/26KaZ
M0rwXghQonFpsw7cCkrRqc0o/FwhNbuLAxLuiekueNI+ZCgUMlFEem1iYa9JK/F6
PWoGQhKm6UMdL2k2tgdZMB0i9WlKv0jQQnd0qDkUDmAUI3EDsVE1amjp8qrlLUYT
tDPPtNJkrgSB9vYgtV65x5sFeO+vAfGUVEWEjGxN1zm7zC/BuCUbmyp07aHQg6Kz
p6SxP2ku7u2CfHnGmjaCu+sYw7yQlJUSfdDzFjQWPgnh8ytyXIFZkbR7ZhCmGH7f
wLRUVrf1X8cGDdeAjdlve85KtQMML81+TucQ1IO45Hv0F1ow715ooJEoA1T0pSfs
rXarU9/SLWvglOLCL65XDGc3Tl4Bgcbk54Wj98yBec6ntq684BnChX+cWbuA5UZk
I3hoC3FmfiLeHYiqNps7EwMpD4fTJjdy/THbKOZk6Tzfhoifybn9Ih8o2YInDpr7
1kPCMw9OOO3vkm1R3VYhS5hkfZ6LeAV5Ts74id2HlRgTy7Ny738KGW8TS8sdl+GX
F3GdiQw4+Mk/FkTYgPbeJSo5fAMy3aJ/MSxGxoxMlgHsCEsda1PMb+aWOXoBLVfO
RoipttxJHTufvKxR5YUwekw5csfhGnrloxEoYecvULRAttt+xkZmDisjVVgl8TMl
NsGKBNKUG8re89sxoHEuKnwr1pHyPTam9Av/iRujC6XjyGCtd7j64Ch/zbw92oh8
7s/zZhopXmSux6msEXNT8UHLibuwbdUJpW1XqgKf5q08sQpxe8jAgwv/nJJwwOWm
MUyPjSeykIb0QdG06jqrFcMLv3IJztY6awzP4isU4AGUMh6TpclfsTcpt36kGnXE
dfOgbQITb2YMbq+L+ACMzFcDRPZZYADdYfal31jkFG+7iw/VqJFFKZx6vOr83rQL
5jcZ2WBpHWzyiO97re4+CChsbjKzBoLJjdSZYB7ewtY7aTUiWJx7FikZcuYFOzb2
N7/csKj5L/eNLkgNVCqV2ysuyXEkxYL/00XU4LZjdt1tZ8/CrsAXt22Y8OC9BIPK
oihuKCloibhmI/AwKB+vp+Nl9+1eC5TbJIvvBliexy71KarlMdLvr+s7lNeMKE+K
C50ePY7NoA6X2mcnHnsS9aImbhVAWjUzDJGxsH6xL1aUpT8Rv/HgjTzKPYILtIoO
bqLAP1p0BTq/Iba07S3bhk45Q83BXZFvPWjnNt+gtF+ip89fFJ9Igksk6/t1Ilga
NAluYjGMm1BbNA7EiORd+Q+QdqSQY8yQi4c0q+fal2HmeJIwC3Io1DQHpPfjDan/
fbV5TBQFCrDArFtj7Yq8wuml4W1W4NnZ63WsokhE8CQocuoTjAD06GPZPOkwt+/6
CBx8G0ri7jC7OTcLemLZ2GYzbXcvIii9SsSE+PDu9D75jaFUIa6Z1ihdGGnfsduB
iSCJRYPVNy++LCX1JrAkqHh8ShpI8qA2xRE5py9eaz81JiqhlYUY+zWIB2PMwGWn
zmuZsDcAa+xdC9jcQQaj6TwuAdrvthDi0t4HoMveFIoaZdGl5gGrPLBPn7Qr/22T
67RsZuh/WciVz7kEZegqItsMuNE3ZZ2YpMA9a+geAQh2Oz1kwgaBJFJVoMf8Q5J9
tkFvsnBJ1JCZdDFcytc/1bDbwN6SKrC9DEtGdrcr/44dS4jie9AvyY7E8h5UGuUJ
GUqTa4BEo8fZKr6mFPOzy9jM4dZO1YLKkLwb8n5gSPaqrJFbg71fR+IhOxqS18mz
lMCh674HHkgf5Sgup1lTuglCspqtxWqC5cWbRrBSTAyYn0o7qIj0pj/A5yq1kbX4
TA09tJDD/Yj/x/7QzYbMmzGGsbuYRcm55uvzweSUHF6Q/gDq0mlfNqBHXBVFEOsN
sJoMXTBN2T1LglaQk4roiZ7GRmYHYMCsEV5n2v++JNZVvwm9JWlwRD97imZmOVR4
IuTN96aXTd2mEmQNF045GaZ62kTNn3d+dk7m1qi/AOMZsrgwciUMgHdyyRrUXi/v
i1Um/lS+QKysxAaoG42xMJZkmVGpWviXExdiGKStfKveQb5YWJlJsu0yw/M3m8U6
lErCzyaEkR8oFUuF9LVWnLzALGYhtJix7poxOUS/5iX3tTG9s6w7y4rJiuUdijoG
E25guFTpjtJlBP4r+dDtHRC2b6M5m8XY8XgQFIW2km7zgJmjMW7OQSJXEGsZ1ckp
Da2dmCS0KSyY7IODOwLMWqLhPmvCI/Td8p4g5Sn5W+qUFElSovXP4rpDUfjLZOxX
FgMq5vYbD0UV5SNxbOyqAJby0gwKDwJgsqQOaR4d3yXjPHmQyx8bb9O9aQrHAjDE
q1eTRcwkLDgHsWoULR0ZXmSffb3YXulRfSjFGmBXiIe3f0L4fQrN2G5WuMC8Uath
lQirIzhNZZktcgOVaIB4dwMMA69PNMZ/8cHNHHlQVXdbSbeRzCUZy3XpuLvVOZuz
mlR3YFagM7qN1SSk9TqFgKdaivQKWj8BpZfxoUVSXc4PYKdP9qJ47j7e0LkXkEgH
zBFeEvA2vznzxT4Od4kK+4sRdEbsCuHuCwy1JW5SkEd+DYI8DRHByQafXXPgDfM+
2bdaLeNPEV/K64uA+L5QGBxc2JowFTvth31H5FgsBptWPxeUucxp7FuhUmaQbbi9
W47XeSatG7bRToFZIObyRAqD9b3smHtnn87KN411YC605MlJXGEIT9+vMq04JT8U
M0677SiCS3myuVhsnQ5lhNnq7zIPm57uWCrs1WZufbNOrec538rseBopeVR82Ps6
JRGVgindy2Lt6TgVbxJ6dGeX9PAflY4F7rxlH+tX8tcO3RSbkiMd1FapHkve6OVR
CH+381Xt7WvG6M4eJsQfHHY9DoX7ib8d+0HOIdAyQZLJanRepdhjPruTp5XdERq0
1eoizf4YDGUJDsV5XXO6G1beDgp7rMczAp3dV06KKdiRcdEta9nbXoe8tA0sHI0h
dsz9IgM6D+JybZyDeNMWUwWQOJL9pzauN+o0a7QgcwlY1r64r1JswTUxXMKXb+yK
avZoJe6NCplTpJ6N8UpZuXb8kdCCgaTWsqoALz9e+by37C/snF0WhgSy/MVyonv6
Rzv5L25Ed4CV94vsDh4e2xEOHmmnDFEYi4FHa11FAa2CpqgDHfWOyQ9/P3BFZpRv
qfpBU1ro8v0aY2rieUd+xCZLuUNKlR3jdH/CALuE5jwEhzAruNnyYDI7ug2h+yrS
F/ideIZGJnjJQUZG4iWU0D/+YjjaKWZi47qoAwC2JL2QtBPmvy62OGsttWu6BMB3
pikvW8O96olKKDHoFKKENVHohw6DJU+Z84qbidyykLXiv9YS+Z2d8IIHcCnMjA4t
T/P432ZuonRCs4C3thwEOi189fwZ3csrMutGtIMl9cSAAlBSgm1aEi+z27FefVxZ
t9EVeK6LQ51DXpsS2ioZ0ThqmLcNI7M5yV6qSsYsZjFgjcjBidR7+JtU5XM+dFnG
3pP32ay+1zM1zxa1XayPbiDetdguuF/6u/Gv2+6St3Bwf1Mfc4DO8at6pMsPtzv8
aWgUWVk02lIw+qEdH1oK8uTlf+0NltfQv2yuJoNziglw3uz/tEmivPY+jtIoQyG0
y3M9l4ED9/ITVKLBXbaOWl3YBHFwbiTmdBTCPfp8yGNFw0DFKRa4Zn6qj38vmbUh
GeY/G26UT1BcuXjjdnPOMnVtXoQ/l0h5K4rTxLeCQ+4FTzLwU1WKxXn7wPBYZ50D
TFJ9lXooxGOldh0bFc5qoSBANfyRxS3RXxUdBfHjee6nNPF1qxy5EnF1q0qbM2Nz
6wLybDSxSOBvuswP+0bZ0C9Jc68bdIg+VPh+G2JYQuLbwWhrb9gtMU+U7pBnRJsx
1claZ+pkiLxSL/ETiG74s55yHF08ORIC4GlI++4cMGNYxVGDCoewFcWuTOk/ZMj7
R+hbQnihINMvD5W9Itv/gLeAS64ho0uw4RxG3PK9BT0RgaJBTjbR/nkj5C2porbF
7A9cr4jDjLlRzn+3A3S4hL4xuVSFetYcd21AFI2PkN50mFMi4xWZB/LK1AVJdIZT
OzBRC9AcV5Q4y1CH288qStcixZeKIQR7F+ungGSt3g8g4eJRSr/l8Va0SpwlCyt8
Ts/snWPC6L3YVlqpBBQig2LLRrsEEGXbzyGNViJTAdJTyWJ67yPWJuSsipN9Ji6e
NeO5nI0m6lLnXi/XTRUzxkt9QcktuvMT2xg1kUJ6GpwU2snRSJcldAIzAQivCtdZ
B5+EcmKNLjXFXUYfeAoBg2RpWTkkFJPZ/IzTzm0GQYz5y3U0jGVULaj1Zy6VPCDJ
JmXi/JT2MFaVQb7rEBuVE9guPtjq7VLYDTQGPGtnf6/PGpmWAa8k1aDEhrfYwPR2
gUEAajBaF2rb/PoM2UMqINyw4Lp4t9/LhZJwKqOdlU1UmhNhLKNLfeC89ZrNlzdg
b0ZI8IiS7pIum2awDzFev5JYRB7GsvIn6vGdJJnr157gVdtOyMVtF3MynMmoeBza
kL2QUQnhFFrI4kkHe9hGSXqa1Rlij39y3GwxbriPSw6K/08C1mK56Yi5zLRh9O+Y
mRn7wBXWGW6Iyv1owW/NnaV4LqboU78HyrbKcWdj3oSJPXCkMqIniB4ZvAbxKndq
YrekFFgvk0BamgyTI41Yf+cYSu1eqMOnmX5AMMp+/O2yEmN7pRIFh6bFlLzN4gMV
/MYWT1oimTmH85nhm0OojJivZPkdVSxrnXRSFlB1RDNhuSTyQeYvHJggKOnpFRjw
+m5sihOSWj3uM5z4+JBDJXY/y8+T1g0Tdz24vP8sR6QpXu/0gZjqeoQYcyFuc6iT
aW/afqgNxPmzr38hNxtZVz6GK/gI1ffN0JxgZuB3XvWAlG2sRU7/mFdzL8mKslql
+sduKqO6GldLnD0CMRkVQfC8DnTt/8KW8CFkgX5Hplw0nammGvMvztrmryQPHeyX
uiRmJ2Jcoc7hRSEBl3IJpcpZiHMh8UwXvAbAD2S7Lm4V98cyVcYE+QNguThH7rSV
ObhM2LRmN/faxdPHvrkDs/dvYX2U/8ZSk68OG6HqUcd/noped+2aDvw61SDCJhRz
aUrXXNQgNtL5932nwVDaUdqaKEMpZIAQw4nvD+/oYkWOlSXZ83NK99M/TJJ6FU41
dvks+VyLbptC9+4dnXdFba0DTdsE7VwiLhP8lIgMFr73VeTEDPc0T3zd2kgE3jDg
yYkNJni8Y5sWwqsK5qonVOURjq17mQGQeRjJX7EajHs9EQIQjXfkkqO3Dffmpke4
0pBBh+X11v28N/8eGrpLr3h9luP5kJGQXaAFAO0rXs4kBVEVe4JpEypB7TB7jl5A
n1HKro8KJtpS/Pe5nb8IuTQO+cnWZSEcz4imSQ14xnAlGdgFObfYC7it/zXWLLnK
Ze+VoXZbgqU8/+0LvTwKh/nZyaJkj8j30uwyTnfHrw0z2mCkgjPrkS1pt2C0w+A/
t9x4+ZQglscblz6KRKfi7PMcF4jpZ54n/A9Mmyi8oOcV+k5XpRvqPwYEAunqGN4N
UocpfI6kdf0R/rDhpVml7Yr397c5bdy5ro45Vbcl5tfRPYe4M+8ZoDOqH2KXF0IM
cpxExb38sjvHSe6VR6k5GZQG6SNwSNdYESYgQG0GbpCnNcY0i8Q3VqNZMfidguEu
ivsz9XeFTwr9WMLVTZGAaQ9N+k7fexLqo6DgzeRkumQW7PcCAZmTzYx1aYHDvE++
LZWAreRXNkEsog/8X15p+zsWRtHHx3rFhInkRvKcBt55VN8AylF/9pLoe1nK+s99
UdsHYS/eUR2aqC1oA7UN5bXAtosbnLu/pEiQpbxHJjnQFYmjYk9e2RCMugB/bKAA
6gt7Ex1oql0YlZl7k8tV6HVa/ckjQLQTVBFFIvCGhJ8Vc4a8ZoKrEryoFbPhFM+o
W9gli4+lXojMgpGh+OSHDoyRd5NGOlBv/RI7NgW0ISME012yALGfOtzTtWkDn0LR
yydJI1fJGGc5Nj/CVneoNJ9LTvHM8DjLpqUsQXWVj/aBaWM1VBWV8ig6UMl7svIr
7Io0h2WLqI/NUwmoJdpFMdiX9+TOnnbtIqAwgmA1Zopykb+4x/2r+wqXCT4rFJ9C
1+n9ktNZyOtoUwpWH3LJZ0dCbndLd4WLJ7jcYhEVg749zMmDJkLW91Lx4pPPn5VK
sw4qD+MGQLMVh5l3wakQshiHshqSw7CPnPlm87ul46/2fg83/GfRfZ8EZKrER48/
mTnz/IODLl+9hzsZDVBsdIUpYZ5LTFroswFoFcazUBi1wVp3Mc7Z/RK54JS4uUXZ
zxk5z2tp0z7aoz0+KX1o+O67UJpZx4qbzgdElWGFp7CQW8H2CuZyLXzfekyLxsCP
SSCdxbc8aBwmdb3PcRyJ9LQhFLUv9jDroiXRf5TCUr6zPfgUUjaXbKSafPgSrHzS
xxCvvoDoDRtpXOHWHyJWBUIf5rC7UyrnqcXP3wUV0cHyBGpXMUNmXPNk3xq/3Yu7
YbQuEUwHDl1cNiSY3gC9vCk4Im0jDNnKSX2vdOf5Tz509PPCLI9yDG1UbVrfiurB
qf0x9iSGg/mOVm6+wDFgvgCl5B8wFQai2Ax/KvvJjdW1t8/pXmlnysENNjKx7Ykt
aZwwvwDLD2KXB1rf4zCBw0ls6I+FeJeRGRrM2O/DE9yUXHhqjRahQwBvLZGGjsCn
32v5DAPzFqgLEw7jNATCBY4J1ZAPIUsJXgn6ZqOo5wcfZTAM9gTQSGrryeh8Nwfi
Kqo/zjAZ90qQSbnWnreBcWPOgQOGYO3JzsnajOBZMmZqqjubGwKsYpr+AW09EHIa
kRV0F+snMTz9hbmIDwClBJh9zuf2yD1xLb2hKELnxHj7O8HWGTG4I/hV00GSnSEF
ga8ksAwHDULn7zdWJ8pdKYU0t4mOdfNDNlTpbGgKmamUQMlJbK4Tz8u0fU7Bdk86
rQZ7TlyfcOuoQE+KXv8zb96SzXNC7ea1N79kpHNyTgbNR/HtT6l8PAHVM+HfYwed
uUL0g5DkYRYAMfcvgBvcTj+JVxaNKUOBUeDJ3eYLSlIm1qQynJFJuBQaTOcO3RwE
XjYEKe76fW8UhIFUXZVhuwSV/CNQSdgoMsuVnIEE3LBMTL9IxnpN6v4vaoDr7e+A
Iz3widz+AxvXFih1wmLRKAZ7CrExDdxkqtONZ7MzeRmQ4aX4EqlGefZv7/ilcpyr
mP2gUj9U/XbiMtgZiEjjn8EKtDSzugGDnkJEeZnZLFnKm+R+HgkHie7xC52lxmZV
IgH0yN9k46F9CyCBiYXdt5hkLRz2yQrBIT1VQrY1v2+9CgcoOr5pnxz7FyyLsSbQ
j6pH5drH3yqh357RDmUjBjDm+TCZ17SzcjecrRoN3M/zIXx74+vHDoqU/axnZnXP
Cirm8ZM4/mZP8fp51/7KWH/4anOi87xSvAdBB3wS5HGtD6FWzJjv0kY6VSujcj0v
ibFy8hDSFCBHaRZ9zFYWiCv9Lhh9WpmhhRZjrtpHeY4eaqL+jCBfzHEAW5o60ikr
UUJ2nGm2RSQLQ404RdIBQdv/MgTItPEaZkTJ9wD+T6qmx2HD9KdeiQ/nTDniA+bH
CVjK4Bb1VSxsnK1EuoX/55PjDuANBL/E8iry93tjsU33hi5ZZ1xYNfPjAsHhpLm7
P59aRvCjCT+Ol1O5hUR+PSrjwkxheBUBpKNFb+huysJJIPuezChF2zF90GjXhwNk
uCyCCWXZvS7aZ95eD9P59TI0IMjtR/g5IuSG5+cdpXOn351aTXX8pgmRh0ViZmvW
r8ZgwFfU+/uZbH1HzFXe+MrL9kZK6/7AxI8Hk0gF8Ap+HUCi0ulZd8vT3QAyNu4N
gIf8OgWR3A7qTtJt3ehyYMRgX7Hy1uBG6FLf5riLZJSJBAiY5fsAS1rT8ApPRJNG
fTellmeeLX5fAdjdakF2Lbb2yD5w8V+VXXoG3z3FJits18MeeHl4pZ6WOFbNsVnp
wOGGUjAwe6eN+qmcS5LtLleiB6wJagRwc3+hTPF3Q/onUiyh7bWkThDESDBkO9wS
z67S1/KjDpULVYSxZZWu2wQKsHJrJrFsWQv4Fgk/b92p2mJP9JxAVH65w36W7c35
d+oYPb/B1dwLDJ9vr7yf1UpBtXebGrIINxqhBRm4yn0qzJDbHbh88wewcKzI8rzK
yFchMzGermZIm5FNw3TJ58JQm5i0w9n5nADnAUPrGt78Nvyg255rCuzWk//8EuIr
34bS6pgx4pT186E9qUqqtUeic2cv2Jq2HxBdydbD81eipYKj4ClY3d0Y9tBWmKYV
if84m1viv5CNuGIMSQ2Bf4t4qzwP3Y55K/SGztsTOkM9QubmwcArzT6KZfNxCP1a
mHXXSMP/53Iv83DTHHL4MxnY5XgYv8zsomI3OBEAMmeTumb2xu1/z6HWWEwDQYZO
Utw42lzind5XSjtM1YIagP6qG+SNSwcKT9UTd3o/z4ECs5wTN8ztiGF82yXTRbPA
yTU6VrW7GIZ6dns5/RWPwj4Cj81/6c2eZ21uvRw701EPFobPbHsSQOvhtQHYkDvc
5KDNrSQuTSNvqiPjx10Uc3bTgoZMk1fAV1gNMWCpkUSyrHqw/P/xi47REo7ITS6b
9ZkWiQeOUF2Nw8jSLkoE5F575fnuT/VBJbfuUws1xQjZRE3uXtsRzxYAqaMzAS00
SSmrG+sZbEFi5Tzzh6KbzW58UIfIHoex8NgV+3otDd82rZ5o3hBr+ExOPK2anSaK
CLQca0tdxXB6v4QoEOm5JGZZSTfOy0uArcwsnIhF4DS3IH5QHU3r+jMy0bl43Aa8
Myl7Y6kGYUH+y+wOCkFmu0zEhJvlCyd695hBdaVu1zAl61jGbzWqG0WSCLt3RhVc
niwST1XbQGt/4mDiqEzBUzNpid3Fjlq752mKya/Xvi3+cxDteP+Cibz0eYv+wRd2
Y/E3B4UrS0fPKmp2y2XXxTByyhtQqy6kTq/T7J8zxddDGErVK2iuOXmwoLOkJD2f
twwUvs7sQM21ng8coJKlIBNwft66KV6vaBq7wqLrRKdk9woHDfxyo+3UuDvG6Mgy
F82sjj+XcibYnEx5TXQoYXTl5YVMSQPbHEYqIJ6CFyWbLtjlTwHfV2nweG7KbC9o
ldaxudUwJejYEhy6cR0tFXBb20x/WNmnYN7+1UK0EoITtTa+phaFu5GRuLb6gvL7
CH/LKJI17Nb5n8aFTsfRvmRgdKSxgVZbBXp8NVkmcXiq4L/PquqHvGAqYGsU7zqv
//gIN8F3I0ua/pOjQ8TYEhcXCca+0CWnZNhZWkvT7km73K9dEc24dbvjSHYBR6wt
yCwPmUpxhuGkKBqbpkowhy05K6zSXIeLv/qy64kdyzR9dluVVZmqC2Hbtr6ltY/2
Tf+9jthucBeEgqWN1g82k8PLNa+NnbobdgrN2I8PiBX6Bc0cq8Ix+I8/WAVpkLno
bSk80cTX8qK9cxfTa5zhjLxbr8fSP8QLQSZhlT9Hhya5NA4ysvXEVm+Jng03Gpzc
jSvPDmpha7FWbOkPkPKRC7F5GyhxjVj+Mrs3FpjBCHi2onlvTIWnghi5yJtihaL8
s1hWyT4Vo4W95iu9tfOJyTXLOuaArn3+iz72AzzbbxZmhKcQ9qu1D3fVeeRChZVG
viVrPgrDRU5kLDE9zzpq40NwFA71WShBUDPBTbh0Are9fTxFB/jfRrKJPtvdYHEM
yN9MDWkZQUaleVHK9XJXdDgAZC3CLj+u8+0UsdfRLsEKgvUmf0gqRFIOih1UKfFa
MBeJto+LW4uj9YLupFFiSPGHc4m8kwh72teKkOmrS0z/O9p5P+IuWY60zcGRfvTM
28lFVZEhvCnp2g7TrvyGcfFP8Kn90sZSgOQ2HTP/1E9KZgUg1NiYEXjhhX7TsMDG
cLy+bD0TXqaDe0EQ8+OkuE4UbDRw3CKEtn9Lqb1ZOi+NE0DRk6QSW9rQxV1pgCki
s9eY5oVd4++4NQLkDN7tXM4q5NRWaXVjXaKiy9Q8M4tzJg+CfWrd39tYQl2PmtXn
CIQBU7sPHwVl6OrFEjVlm0sqCV+awAELBRYvEsLFDlTriNyKD+AUFKVmEfyUG/95
m1mw8k0djcpVuv/4fdSnlCEFNWfJ8ROZZdwgse7F4dORBirrJqzkp4W+NroxMVNj
LusuD/n06ie3bJbt6JF6BY+G6YX53tl7I3s09OnTfMAegRnZo0G104oPHBZ87pj6
vl6pNP+/1Vy3qbAPU2G8ORKzI1+rtkKSq5UpWhSZsafxvnBKQU5hvHCnj/nkuv0Y
puhKQ2T5hHO9KTGTS1jO4s6LJWFFbW4tyPO4XF4YJbbqFvKrfTmqdWRMSl8UyQD9
91PgK8EkBtxDJI9+xegwqi+YR4VXU9tjrKDeFekN6+A7eyFb1EQmxAkNQgom1IxS
6eL/Ui2/TcAKIdhTvWd3rz5euHOyCZL1/jDompACs3bgbvU+eb67dsJ+zs/xJpPV
zn3aq9ezoeDe48zsf9e9Y6mCyyioW52KVwrgIPP0ES4nHvfyQou/Tlgi71TZDZgw
0TBU32dN7b2D2c5z6U7rVToaHGbF9DWrqm91kATQ5TRMteVoteCHBXYKk5OFWbHr
vdJXfvQHOB1mRJh4DzxH4NV2WY/3ynIdODCGN9xttLeTuH7LQ9FU86LHYOYNkJJ3
hQQa9CdEE5j/1irpoThrKxRFHNRpSGQJ2ZgMHq6ndFzomnnsnJcqjwW1vVYvQXua
t8Ysn4VHe5NunT6VXspATl2QjBKrIoJnvsHfGiSY/MyUAYR9uIL/lcAQTxYr2Ckf
z6MN1o0aa0upjrTrmqd08+Tv9VrzSzZX9EWQXAZFXOmAgMF4gJy0tqLj9vRss33r
At/7kGzfVoGQ+GZzqH9JugYQv1L2NjyvsYNFYi2B1v4xfgOLnjAnYjzNFRebymQh
UtmmbzOjugIviOorgG6CSI+PxmA29dF/1wID6HTkCYwudA4PrCz15TkrTsS1sZJm
WN9L461dpuYWcYwOTb2Q4ZRln7Wu5MIoiltn23ulzkOLNeAkLlLy8ZBmKmVJK9RO
V5ky/M0bjYXeplri0IBpHqd9SSGWQZnrQ0MpFkbhW3n11UpAr9xyJoWbAVI9YdLF
nJjBkj8eb+Hvb3ZtiB7fZL0qihVdybBFgVnmUUTIIho3OMESHmXoTcGwmq4oHkSZ
bSUosY/wfegzo53OsmghbDE1pcVsYXQtXDx1tnMKwthhpJS+16GuT/lEkkKjqdLc
DxP9YM805z8aeVP1yz1wnnucOnd+VB2qxRyZBf3XBje+FqDnK3ECLGBgHjo1CsNI
vjqVcFy0af64uW2bIwYzNmjY8LUjJSEmvBsklLndGFzYvZZH2LI/ylall3uUD5nM
yNAro0+rLZPReY+Y7a2LXPhIIXd8qQ1iSRod9w0GRC7ND8ijGW+JayYn4qF1JQV3
IaVZgBvrl4vg7c8nE7dGqwwS9IPcT84fSj3AITFFlFuKYjr2I38ZWHSBn/t7e0zE
MgmD+utFCUrzbY+9qWT6C2P5Rm4lnMWhrtRXzrjt8mPTlrET/OPAMirexQeAwIss
lQ2qrKcOceJ01Dt88ZWeGVo9LRShcQAUHPl1uIf5La4X6k+serQ6SqFofQnkxJVa
SuCzMBsII2CDPUxR1XA1+rvGHtKvlptDTbWFlVYI3IUJIfeb+CNNQx7pBjvi5mUC
Zf5jlpRh2F5y0B9jBF798/bWsgRHE8ZS6B+vQgBBMkm3SKD4k7FM0PPqAeawSUOG
f9UhMPjs5/7V1ApCXeJSnSLXdriP7uMRzL4XJctmYuBAwROs+NnZU2kuMu/3IzsH
zgcDfhUOhrOxNuk7Gvqmw5ZnGw4x6oNC5T8HhahRFe7i5aVlE1DA3xh1bgwkuDvq
f3Ynju7e28qJv7m1ES5/HfiKps5K88A9FDszqMasjh9sILXFjuw3qmvnMBadwFDl
rfwxFMV2RbhLIav2h3ku7CYMUxGQOEf9aAXtEUxEbdat0ZoS1tDEx18Ef9UT/SI7
golLrBiEMh1y9MmdJ5z0S9ZiTjXzJIIwKAnENA8b3Wb2azFXsGSxzQi83/jUxaTf
68zXqEgnwCet39CsGVmrL6HDPZ/mTw9puu7hX0OO95+hVuVe+Hd+G6uQ+uzuvbcJ
ThE+Qat1oVlsMMlKvH8lcSnscT8v1VWS08vA4OF3ziGN3dSEHQ4DTNjxlYwXgbNb
u0WuhSM/G6Hx4MCTqbC4lQPCTUNVpQUvIL4OK7PgN4eof0wOWE678UCFkw6hV8/f
4uDPRlm7/gzHw5yIhTy9sNNMO42sPc/DtSVxdoqFXosdrivbhEJX9LLHZ5u0Rv3P
rxXvsPBpEC+vme/KziEFz2syduU+LWAqMpZU3StvtfW3kuX4azLc8E6aMWWg7uVn
yy03rHgP3VxJ4/+XRCAZnJxydE4jLN8GNErf2vv6K7cVFC+/73wMXqqpFrNmD2sW
h1vcIDs+roc8tMK8g00kKCuCminRFIQAO6kPxqTNZg6bHCqfIC8M1T2pESDw2B9q
kSo4eOSng/uyZMcX3XcoHgTFdSGmdSIzH4aL37KqAgZP7FSgMNaWB3JwDCDStLBG
JCIo98oHJTPpP+ct/6SLbzDqyfh0Hl5XYMt+6UzEBvfk+ByC9tUQ+psnYLIRIaCS
GktUpzaghp8Ogp8unjLxS5+IvInNYEzaPES2qrn/wcUie8m3pr5SBGf+b2T33qdf
mw+q+0KqM+vkKqLgAqvJBVcQgzI0g5a+s1uZfYEJ5sW1M/6vKT4hCeRLFtDwvesu
Hu5bmc88WwgpdWOuZAckZYTFzbHSOGSCJE9JxVsgjpQOtezyLRBXxizEkCKwDApo
s3dWjkqrOWkH5dejMRr2q8D44WzQ8x0PEIN3C1xUQ/7zbxHDL7kmLMN/w1M6Kx/g
yI7DitoDlj+uXp/tH23Ii+cdrn6q1hDyLB18Nzgit1iLw2oT9q9kpHE15quPRLs1
nGdF1qiLEe5A+FruJMFYQsl486Yru6nE6hTd6BrZrvOg2Pblb3gwTsi1oeTcv2Bb
LAi0Zg7D7doxYjoQR7A1+8FK60ST07o4dl0Ngd+mwHuni0EV2cLphWyXmWeQy3kV
m8ByOTDIiYoxe1arm3fkZ+TLMr28KlXPvyGOgMo3zOd0Nt7VWRkCfB/30dR8S/OY
ImzC8R+4dtDCYNNg+au92G9COzva0mK2H76W+H8Uhcmi5eR+GxpEkkYAob9E7um1
U0BqToao+QNoWhB4eRMxXp+a6czKsvXlQb32fz5CCzKLRa0y4fU0pMTZY+mjwKLM
tyryXb7MoTfnPUreEXWRJwPW/hX6P3zm3vyNSqnfe6alPXQv4kLns9cG4YnSDJs+
Ofru0jOI1/Y89qWWZVWkwm1vgVBzFprttATADjmAaa8mSUgENzh7MaeZ+dDJgAlF
Y44rplz3r+XjJBTUg32GNc9UBzuuYpuEkGal8jiaqv8BxjRDh2H4SAEUiCGFyBqI
EKMrY8rOke5BJdUBgyiWODNW3VyfC++Nx7a39PxLNA2FSksa2fc7QTsX1f2uAWwx
8rNfA4y76KWxwMvu8tvpJftuFV1DfstA/tbqYHyRCNQnX4oWb3ZJc0VUkyh9B3ee
w48rfNAY0UdUwjcbL+P/sJ4M252h12E9iBw5joHBFc7p7v0chgODxXxz3YRbAKNf
ySXQcUVRe89mCWLBCqXEs0v+js0jeVa8R++ZzG+hqSbqRt5czMAgadwsAXJ2z7v5
lzdbCPOVprHTCUaXsrXumjPV6H3dd/SrtmIOk8sTRj97GeisCvAwieOcDj55kPhP
ycvPoK71FgE9PQsNBl9LswtZwWR2yFx0HQKORycrEf3rLkhpLli9fJeJ0Vlg/R4O
YqQaIxQWCfjvQ3xkOTYPnW+dZDw7iG/Hphg/aXeMG/u40YUgs+sG+SuUpKD5xeRS
RKJBpzsd0wiRoDKtS5/HbGuz2XKL2ctxhaOhrgyj21PBOm+1yNI2wBywQlfhObab
L9F6+tfPLwTq1Gm1y2o/X9UFH5CLRROEa1owxU2Z3X+IswIECh8W6b5/KF3APeDL
9pq5MLBXN/VF6iiRbjepxciMmrNNXZlLRNCYM84QrOEwSN4gTg/Gt7sKWacNEH2r
hnk9tQWGK/zwrrWAOi7Zk5MUPJZvNfROjiLmt42rBMH5XIYqAXC/qYPhQI97KGHA
7TWpzMBVny32AkkA0jrjlUWoPNG/3SmkWPw9a+k32eDN+9OLhZbnIfFsxdz9p1CP
fzfibC3qQt9UVuqZqoasTzHV3qJpjDTlKQUBL6MLfwI9x6V6146lOP+ne4F5pBiv
D0hcHjQRE3qhkxJ7GYV4j5ekyXGX/+8oVXiLxmjk7qyyHL9RQC1tcwXhl07PA3Bi
XBb7BdWWJnClyDDgsBfGMVfZY3GKfReXL7VrF3R2zqnW20x7L6BSkG6XWschbz6u
Y0qbcMmgTBbym/wtc0AKtlfJPAUONEU/1n/sebQmqdAfToajhQLgWIoF2/8bgFOU
SuCsqgDwOqFpGw8z5HqYElopiJ0yBEGGA+6P1HfoOb+ncSHjGM5nOm/gJ07JyLwA
MnAt5rUyCHPA6Bhc/6A46oIEInlgkJQTg3aX7tAa8FTp2qSzd1sGmiB5h3OKIvvN
ObkHUq69Vr3hSTnvaaLUaColOCnL+J1dGIgXFuRz9Yo7rze/2A/trT+iQ813LrBT
nJAGmUL/lor+ViR+OxcqPrUZYwJPwPsQELZtIm+CmmDFFwByHWx/PAXRTVnLmnCL
Oek4CuiSygjYkYBTmu9EEV0R0eQ8mRqQJAvX+G3WcaawAlaKKxHwrqogzV9wRWhP
INRqNnI35+RGhJ20SCbMr+nBVUYVrID0KndghyaLQMLrW989FXBTKg6SuGCew7Nh
//2WgAS019vOO5+NkTufBBmu8T7f0s9BaIps3p+XsIV8cdSxrmCdEUh+p89bt55z
t7n1Q4BX4+v49+SSF9Ei9lkHAWac3/u9mUh4AVz7o+2okVuUahC9kfT098wOQeE7
ryymd04jIcVHOuJdvggMp1k6filWrtCmFYNlUOFuOUgXW/9ss/t10kfiLMJFEuLh
yhpSCau0HIYaBVyOY/Nm7R9XS/woN6F4dxsdBGycayyMTWowNEhIrUQCgCybwl4p
n0IeUJ6EpvnXM9Skft1HosU+zvEZB/YSdu5QcYb1HiFmS5cGBzCj9DLi1cVR2P2s
rKhtPyHgGDIki+CxdcdGt4+dQZirepTIRnpwmn2lZP6RvkxlvGB30DHJ8Mxwo86D
pMAbG/RZQD7VYAEbivQj57FRJe8l4O9K+K4oUxrG0J+vKcND0PLr+Ar1EiPOO1/W
m5S849rQv3lyytgXN1aq6Gcaf3rqRFcVgK+O3XrEfm8nj1gtO1Quc5/RcdiTuWEl
9U37+EXfS9IvPslff+90ZoI+iOqkSKj8iLUJyd8IarUsO1hvQcCnZJXcJ1cZn3Pf
kDtp/F98uGEExf5dEkgDyovJSRXS5SB/I9xz7Cka/ZWbVatoGRpsWfdFdRa6BR9V
/0oZWiV6SO2YDMUgrxeYByP66B13gLbvwfMxlwlrvH0JZvQyVN1RdLpaYX3hLZrX
GjESG5I3AiOrsHMqgVg62sj/J6ce5Mb+CNLkgwylLbqq8yUu66MywtclHbcv1ppL
YRN7XYnr0rK4fUDvZbGmQkORELye12GpSoFgmYqN29zx58eFTt0w8Ik7y9dDjYXx
iQpTXru21lKiEhqZVhZ2TncnvlPYiAfQMecf058ShuKGhDW6efcdRcqNKhMt7Mzt
j7DjPi5xs4eEvsZYEzCxL90Y9E7EDiqXF5EGfL3+8Zjjgz0tjp2jWQmCOqaJIMMs
IroPgjCx17tDTYjHkh9QrmOTZsHOF6wPhZm4oA+NElSMuaDxzTgJZOW/AN2zdy+K
TOJFrgK8x1SuOk0nznZQFdK9kU5TQ3BDRlswBOW1CcIXLar7q4H7zR6++yz5a4Lg
EWMxxJRC2hKHO2KvBXMxVpDhwednakyMxD3u+vSA9SDhyZ49yvv8bque3O4BuRpf
xf9q6LUjyUoMVfG1iFFwFIX/RAud3Yp5wZYiec5UlEQzpmsj1H0JNojZsDaMaj9u
uVTIYeWnNTuuKK+VaZBqR0UrkomV11Nmf2tgDwJE52TABSghNno8AXr/okAj8APa
aJxQ8wkwywUaXTNaN+SoHEs/3B07lEXBLjHwNaGplXYb90CZxItkFOYcaCt34Mx/
HMrZhKrczWR0FCxyUTkAOhXqimdtHR3gRh3mKyFiS4Ml6j2wTfGD3pDY+NIx3CNa
Xn4yhBeFdbfObqOiV7BMPnGwMys8qUyel+e6Y4Gt/h2Bj7F/OVHim3GahJEJl209
m1VS4yu2/y318aYwHkHHz4lzxKnzBveVIt0X2gJjeMc1+iIB1s57yGiu/BYdpump
P47TcAIyml8I28uWjzpoDELaVjBi9b7dSGvYDcFln7ytcS0183gos1GpxeXkPgu7
DY9J4HuSpG+F7z+4qFk2Kxw9GFupMUcoEIOUUCyKBde8mdpN68SwnnmFYDXl9EpZ
y/Xj7dH41YPMSAQ+w0IkjB8L7nJWh0URF7wZbglHvAdCQ7+1o3aLnqOZukP94fI7
auRSCu2+062vCSLrwXTFRw0xLpKJn92RoKyM02fO+cfeoo3aTW6aKe4Pk4DiR//j
DlZVosn1WCRTYI5U2KbxrptZDz4d0MJs+rtoqPbGFDtgmhbxxoFIy9IfunUhRNUR
d8LVEpJxkNKlG2lEuJFBd7LQ2FX/qR5sAb/nC41CB56iMljFF1+HvLIICiLoZtrg
n4e5Nxlv0SU1kmS+UfnVPD90vxk1sS3K81x2/BRo+cIymQmYgpp6I9A9wUql1qXZ
K+x4NI2l95QXRm34I70TcRQWK3kizPOp1FpDU3qExTchn5QyyVOSidwGikNueU3O
JVpvfS1mwJErrCuqKcHVGqaFa1o2gnFhCHM5MyfBD5dkqWP9Cfye51tIS+5GM6xT
EuIrZFQQDPnbmO3NsjkXTnVEqseCaAW7G66Nifkzld/nzf8Fj/aun7YZBDkroG6X
HsHzc+J2jspCCRPbUhfhOyzwrAONCgzuswI96+MNkVPr9GOBdLOVV95KaYiCXuNc
cqTB2XNQMelVyPxz44towDUU3zHdpU9EQNQshhwdpTspCum61TjXPRKS1cyDns9u
4TFVagXqrJNyXzR5rKsaMVIHXMp4WZ9xABvAhJNVIJNNFZCsKawP91bS/Eb0IA8i
jX5OMepYQS174qujmU3s9MNDiXzgiMKIlmvXQUZJ6S6T4Hplgv7I4OVEywkOPhb/
tx7stQg5N/ss1RPNs25Ugn5GKMGote9JS3Q9MLSV0jn9rVEdWxDCE5Ss0Sf68aKa
fpX03KaY4zfl7p/fmJ5GMxqrAwnYkgXu3ojC5bd+aqy6DoBYAW8eDmwaQmbTPfPS
YokGMGYXVQQH1RsNAHZhhThy1uPJrKvGVlpPptztJ21n2uJbaeXo4G2wyvm0+U+k
9I+z0Xoq1AZsYZbT07a56+1s0C/00hm1qQ7vSibE4vRArhH0bBjTAP+2ntJKt4N5
M3pv+sNA0pe7F+85/F9itg6/T2pwdSFIEbkUQEEST1lxGL8ErY94C2nqv6jpmtb2
LsCFM+UbCeJMS7Xt7ByDRxBD5R7K+168IUFvEGrnLWvJkIo5yuUVH1jjDTKay6X4
M8bPwuBO5aeozc1ACm2zwm10FRrnZQSu9msOvADqP2AFH1H4V8tA2YeLkMexi4mv
vZ/JWdJSIwwW9C4T6BQ0SrgKhlx49BE/TfrB38IlvA0zcuNTt0/MnBe8j1HJe1EP
YN+cidM4LETgXNNXG4bZbE81rcjs5T/4BldZitIKnYeW8h3dE3xlSvv9o6CluZPC
a4rphtA5cpSyMZOO4yGBxr8jSRBghueNxhrp8RLt+PxnFl7ONhxehdwX8cpPFdCK
m85uFQPPPhY7+EH6GWqFJWReUZ19J0yBTvdaVgsK/ce9GneP9+SHCPpGiRSxua9q
Ic9DxlyjZskn4aGlmo2MZS6v9C4Gwh9Bb0EqOrBHg44CL2G3Yk8Tl51chBEgzRTZ
YK80+/P59ZJYOsjHVsnp79ltjq02vpY16mfkRJ9X4bhvb1OBdUfAqxoiDwolwjAh
UUOj9Y99FZhUPMo+iNECowcrjWr3KQxiu0JH7UlOS85gmAP6y03RuldlAwu6fdne
RoM7qX67RezD9qV5LBi7AR4SLoK2BT3415NdUyvDBThyKSjHkwPMLaWIB14rtl0c
izDnBBFDypKlzvdQSHLX7X310k9OXq2QnlAIe0l9hHwbFc2aUZ0PvkBPtf2yNt12
/mapDNwgUXXw8faUZLqFmIoLyRgYLb3003jD+YfJHcjvjyV92BRphXvugxL6OiK/
5p3cKh6YCLSyNyVHldNwN378CdZbgAMCCBNutqE4///Yd8simVYemg3HwSJWi+of
w7Xhd8SV0DLxUjlnWt3JcNNNkKzJmid9XKKLdzBqcWztb9dNWburcrGXdKuZ4Ih9
gCw25G+GXLcH09SKiU8ZJ28K+arlPSAg2Jx2UsLWs19pzQtOeHI4498LygcIjnQY
lstEiLmh38+xt95fUejJavwZ4IBxAHOQlzsJWJKotAf0Km0bwQKgw4Vqy91Anan6
TO3BSh3dpTBhSZqWpAehx+cypl0wH2SoO20lqmFpU9RqEs5NWBOtzKla+gcIkivv
eJhWc5X/slWnLTHcqHIugnEgrjzQAY+Va2FWt/JG1NocWMWO+/S9q0ZJHiIvRm8G
LwBvXf2M0PN9FKHiGfAE1uNCFINSIP9/4HXJlAaagDIsntccB2n8idey3QmOw7oL
fd0+KWo762+ybFebcG6HS4BA/FHK/kSZBoxhwY5F9ue2OZGvMsqBQXhorBA3VgGC
4XMidJIfnejK40SdkTQAX1hdrS/fWMHkcdysAXYMv4SXsQcowBLVIAG+9U50ksYq
adNJvHlIdV1lHKI2OoYFHXZmjJR8E+Ug2JFUl7w9pWlOqg7NsQMwKpaQbRjoGYFr
9R9xJDlxUoTAC2BOMnLdFqzTQK5F3wrVfSKjBZ8E6sbnAoig0iob3khH9zrixjgo
CMo0ZHkprB9e52VlFp0xJmMWBTPIfUDdWbpZJtrRa7Zf2nbR3Iu1L7UhmMgofNW+
7nZtv0bDpga6lk86vHotOeo7dd5QluKjcyfkW2iCbVRVYHTPjYvbJic4sZ8DVN6C
08wBJgbV/7n7qlJHeKiPnkmj9qqXHxNsLEcXwuT2dnKptpIVn3tfxVgaiBRKxEGl
qE/8gCJVtVC9TTP29x9MRdFz8Z8N1yTVR1bWnaiTtTC1SQ8XdJgEnOXxf7D1DYDu
vERs3H37Wo60L2cDnsTu4J+IxY8Eklq8nUuF6G+WR6vxqL97TdH2BHvo8h/TJZ2H
4FQiNyN3b15wtKZeWE2AEQsx7bRjbufZJHTijcD0S84/zpTdHSya5mKJTlQh7tDO
KOgCR7CjJYfyTCzzqJx4bjtseTERkmwilUjvxWkalEUnU9f9l2LmzYHSO3Umllti
4qPN6OPczBgIr+HaTulXAxZeXU50R88MDikTNNryCqX9pPyjh3eYw+tQMEFmgEHG
tSSNbs2Zd5LtF/8qi4DNYN+1wl95UKDF903Rj0RJPkwrRW4i2okXUz/bIeKCr4Cz
8NWm/zOuqoxDhULRmRJ58h3jydyEDnU7O0S8I/NomfMw12XaxgPN1T4dsRkZLgAq
KkbMt8nVsrK5/awEZ0/ovb9qUm7JwKJ5l3tVsjv+PDRS0m7H0exym+P7smyS84Ga
cAcCDlY97N1YMPc5LTQBZEHF0rGj1CZxu7qzMR2rt7wxL/1+uX5jOFjPJT21sgCt
0rEPbQkFA0JKiMZLGsGXh3mjMbOO4YFNiewaTHcpanOrfJDw0CB90c5Z07LXRnNH
tyJ7crgCWgAkXtnPd6hiFBHELrlyBfvAhRHSpNWeZKaE2uHulI2YD0vgDEheE2RJ
ozbT9eUksmjjmHisgCJpSo568uKYycj1uo4ve8vsMCKJ/uEIq3CBAdI0qr/Pmm1z
fMZ+LZXCaPE78Ad7/mTRof0F2ZItG+L81CIF6yKvj63/MWKn7I+/77hzPXmggygt
cjMkXMQpXy2NbuL9fyCi3EthkZAjb8Wwurgk8SpD8GdshOwmwYKFcaj9S82U2yJZ
S5tYFlT8Rz5q6YIkdKy61ctFdUq4NAYV/UpXFAtPtlOGKNRKdBgMCySb54BNERQF
+Cq/+vamSjXDJikrgTqvXa0/DNOJEVSUipqoCQuDyLz9PzCcJRTNyQIWWFGrxSfg
5fc/D4i5i1E2khdYXvPusOSsuanzI3pUoU77CShC5x6SntAkyTCEPTakURD5YJD6
yaWtrDdNxxn9Rfym8fQiWf+SoE00DVQtwGjoswDuBfOGm1wOwYmid2Rfcsw892oP
TL5j5tS8ntxYNLzXMGJF9nV36i7XGtDcHNHqunJnt5by3mOOBZlSp9VirAbXIkSK
N+zi49Zcd4ykYtpJ5D2mx7NYGWpDlARS6yQ1ZC7hCkUlRdMDpTJuJ9KhpIJ7JIT8
CbYaAu/2YEqx6xPfRHtR+MASKmEqv8n906xbPahyMzCev0ckEnUHxjB5iqb8s3Eb
qo+TfvWA4H4j/aCOMnL7eLWvTTigeNIN8kZW22EVUm3wgDZkOgrV7zFxDEZ6mQ8f
DcUUDYJmIwqdZXisk82fDuhInZWtZu18pcNJcCbwEJYpsYLpIUdpz9l8UGCDowGR
7Rmb1N38ZlzKZx69QQIp6F5npgX6x/ATSIx94aIJC5kzv3tuapQp3Nr6tViveHSb
r6RW1IvKKFdU4c4BNxB8sb/VQAxhAYPHpT8wcHDu9fmbEsTGpv+nPgtmWFj48jOz
jsiwiGQfvR5SW62HCTQm8eOlFvSpgfefGR5lmVg/Xxz+lTpM0fKp7cANbhKfWeKx
gOx56Hlibl7HrNnHL/piBRpR4kfGAcMeuiCWokWXS4+nJJoIqrqZBmGgR17u7Ppf
`protect END_PROTECTED
