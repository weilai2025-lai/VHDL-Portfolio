`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIRzSWTct/lFGn+6IdTGf1pLchW5K9a8z99CxNf43Kn5qDc+Jpg55tJxB7WKn7Ci
smHecv3fZl8FyqRIn6rr2PprQ1cjpGvJpWUViD6bHDWvWnEHTSepiT64e3yawwDz
Ib3EhuJDCwN8gcVbf27kPdZRBZRTiPUyUbsS7BWH8pkp5vWpurkKsAMWH7VEyZz7
V6SSEDHjMgem6q+TznsiUsIUdjVgteislfpeyc4h5i7En/THiJbENEt6seJiVaOH
Gn3LghfW6/c8ocBrn0owQsnQQw2d9H3otyoR4bpa0WHySNjsArXWJsHPhFt1O6be
GF4Fj1pFpvY76cwr5b9EC8tBsS5IcwkML6WsXMuUSMcH38G90kOz6WpB7NAQsIqN
f3uFAJiOB9Kq3IQMUtyphp9EIH/x/BWkN2wJ7AQw5LpVl5iG6Kdq1aQOqypyoAW1
r24BcP3vxAJiQ62HPa9gLg5WewV0u4pzNLMXA9+cuT1tL+/z/dJUYfE8vqh67APC
uYUFJisNIDQWbzjJpct9nDEtbELafnGK0W1yBcKF51fJpx+uMOb4p99MZUqDdLao
w7PRn55sE2e/DZftr7CX9eDxCaoSEoArTEOknIkeO5DAkf3bx8FFtKvNZvjdI1wn
CsPdD3yEw9rctPfOMjW7Rdghf6hdeSrzgfeXKk1Q8xaUij1gR6hikeXifXfAOPD2
UXZCPTACG/layQ+J79mQZq3mUasWEIkatzictMSGvdQ=
`protect END_PROTECTED
