`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bi8auP6hgbNJwrnXsReTxLYdYTcclksN4oxO88wurcV440EJ8uW03sdPc5weIBF
i2Zl3UkmU7d4rmLEI6LIfb788PsgUGrB6JBKw6MhfJocsGHXez6gxtw0UR1BlriW
qmKayFexFUuZpJbjB9lmJNm429kiF30aq5elv4zdIUd/65478oI2e1tutWDr0rzn
9X9bslJdkwQzIScsyfA/gdwTmN6Vp0KZ3vcLnIVgRWhnnwSCcAjHDR2IMJ71/FET
RCW3ulA4HkQFxE5qQvOuRx0LWghoSg/GpSemsYQC0+aVNYxe+q6pn2rbLXHZTf7H
3HxcC7hG0nRoHAS0bRU0nvv4pABIstU0YKxhgUrHtvoT2hK8E+2QmPXuyjqMk7L4
aUQHLpWajNcZeVVsmVmCRupvN2HZkfXUL7QmAD6TOkFXCZUq8L9Jcxgz7ZYvZLLr
cDtalHCxHdiT0us6l9/4GAFjgNe2hTB8eX5xll4jkApl2t7bsgW4mqYOaJ4NjsCp
phxOdhKEUOvvhsmjoobg0rdo2RdHaWd0wmnRo3OefVb4A4gIQQ1Z1uf+p73at25f
6ONDUT9winpx6d9Y75Gek/bCNXb6IBc0tiKa4CB69UNf0jKXH4g0Ao+9chsTPp02
D88KF4S/LIAsEo1bzKN38gKWD0FlnPISbxNz9zv4BtBXCfxoIiOlDgjZ79MppSvw
yQP808/tt2x3LAQQ0Mk2/NkYsqGbwkujV04dGQx6v6NLWDm/37IILGjx+zE+gTuR
ZAu4MKe205HrLhUGBLtLobKRwqaPS2e3Ptl1PIKgYs4wBYnUxTgjKfHCKVYuA1+f
55lBRqGbGYvRPdPsiLFdga27JcWJGY5g9e3Q5CeNx7a6WyAbz+09BanthvKeGa6E
0pzOhcHwsx0v22mwr6bnHEI22NQdHsV/lp1HnNbSnGmUG93HwnAOR5kO+xIYuRzC
9KX7JUVBcJddp/V1xvy1iqDQB/AHBv9aJGbcRuSiV99iCw9KR0HRmGLoe6yyi5pZ
10ivieHq3O+2GItUwMVwVoZZxJPp9bN3RdgxFZJ3RcA9iE2Ql5DcGPWPji7n9lXS
lTYWRluV4KSts2MzaowXIQnhzHbbpQKXWV6r1ELLcxkAUStmwaeek41oDhWPbtX1
J6OG5fsE/TGYenDEU5WFfXNDWl+bzi+TguC0pYWTzDZk+KTIPYqv2OS/chzX6jKW
hP/Jt85UNRG2nNpBkL397oSjqw+0c/FGjbWRPbdGtx4orYadHFWFJZuIGICZ+Czx
N7RyyLawShCbf+Rmc9D6X5fLk0hK8pepEzaBf599AtStMdFQQu86p03Sz3ZfAdXL
/kvwYhWRMcZoOLlFG4ouqHQ1y4OQL70Hw072LhQs4kYg3NwB6efM9/Av5aStlPUz
x0/djWApu28uwZYSvpjgHM/RB5rbTMDjPr2tgbgR41L2MS5t06sp/jc6Tg4bBfoT
nhYHXN+lnsyfVfLcHt/DVodrBBAkz/oY1+/O4a+XR0FHXmswZK8ZzRQ0qQ5WUoLY
FoJspEyOkptrHjl7jgFjcC+MbvDTgRrdL5dO8M5U0DPQwoF3Q2i00nRzFhWjf+8B
JWig9P0tM4FmohZAyUxJ1oSkvVkTta5vbOT+oGEDK2pBZqi7NRZPDU6AW6llOPOI
g585yV07XjILI/iOajaLY5xyINSY9MDbLaNYdisP6ZLo1ZwDdN+RTGrJtc9jN9Mj
ql/5/SkY4WVSGBUppuclXl1jtvkAgzIYbiAWzTvimWKhQz9YcHAI9JLAPG3FxXuz
h25AaqCTb/BmR/K+jJ7NbTKj/DDYSENUn7cjxeFdb/SkIri9hY8xShZ0Ra6dC9oM
hEWxnXPvYaeqJlHKOe4IZb9ZQ/vFMvmYYNdAzQFM24+IY4GETOz0Pn/rKDkxazq8
e9+xCETwuNOFpPeP+F2V1RoDU2HPpNFVqLi3EK9qiE9OgkTTC1FhBJkJk7tINEOA
v4XKJHbP/tp3A1KAgEFUe8DF30iF2BRZCokiTGOD5i4+q8Iu5iPml7PhQll+FS5l
Z9TC9eom/bx3+PPU6Vh/BC3u0T/fTYz6EbNDvhroi6sx8T6KRGlin/8KLNVcxKhe
bY/AIzMPD+Rdl0IPEfnwd8/tjRgpRQQR5dO1nfC9y7Yid9EJxANsLZyAG+U2NYof
tDTwbxlp5NvgeE3cCLxpxTdFGuRXsFoGnCuV3wjJv6wHsl3QeDEjhFuyjncxiMzv
0SCZ2QHLJgm7MIEqfiCts+zU1HK3lAdUb8zbOttllDxKRwDi6h583sjbGm4p2aJF
8y2262pV3cV1ZKMz6TeBvc6kxqXmwetWdyY+TtM13Valaqj8sHswGVDi6Gph2WjI
3SEDxiPCsTOZkDAYa73g4ZE9LRzbxD5fHs3RSFgy2+XtHXTiyVrm6GHJfNUSGqdw
x3oXW9KtY6BaCXZUl+/gIKv7L8r8BIcZM9YcN83ubo382OgL0/yZsOX5ncQn/9RT
ysv0sw6eV2AHmTb9tBmdEJ299GnasrpuO0lxbr1IFOALFAynJnW71CQPAhml6rvZ
Alvq586t5yvKgeL+Dd1oUmPH2WJ9JMW6PxF52oSy7zEP26a5jhyrKn0NORzh2Tpp
PWv15Gu7y8cGmfNuyFTJ+uZIPnKVRq6lXifSKV/oerfT+D5o0JCzHgqQUwHTFGcK
R+Ls3YdKvaJ89QibfJZ68ym6odL+GlVK8HwTtLmDktJPW7ft4A22V3PyPiIG5mxy
AnNinzT8v0Mihl36gEWO1RtRVthoHQ4Uo3H8796E9BdP9nAOc4iR8IythJ/pRgWp
2qGBWMB1PvkKbhtIdCABbzEuGMuNNQvZhZGYXKQVDA69Fd7jecOInna/15hPer4p
5UfcIcGyKrLgKrEa67MFuNkFIUqjnZE9/FpQ5ItXXtN7YJxnkeZXkQ9tBWVzCfW/
BYtKGAeUiCGv/xwJaB0/vnl3F51aPQEQOHwPIEYEY8Ad5Q67igCYwDaEnxjAw5pz
tRmqqWb1ZO6p16pegchD8iDNg1SIeLDzn/Lz/HH1+SUf077403gb2mET0Bqlt0Xz
uCJ6G0reJPshDhTPI9LiHct7rAYuxtb0rnVhBM9xPzlkHjKG4g7zvSUS03Djf0sm
XVNOvOsLfTL1MdK0Xr4BO91yl554vHY1vWKa/yyXbxaIrAV/k/axLkRswuaP/xl0
X5DqroVTKvR4BPu8Pb6rlPIA1z38AcYuJQlw8EFADDnsiK7qVbn/Ye+ebpFyl8kG
fZiZ/HJNfVqW2yJRqUncuF/7pqlpxyKcljuQPgYtAoRrmEYX27fo/csp6w22V7Z/
vkWx9sYalf7Kki7zx7Gfd9lytEZOrGHjlghhPGAGP6jlbk9haAdPrfj9sx9hCmn+
ahw+MYsVbtyBv+dFZDv5P73I8toGx6ey4NyiTIOtlTqz2INyvbSapmXzVB1PqN27
jybtHhz8K/N39WLdF9bm7sOacKZKFiDNk39GiEpI60iu3FNZp7zBf9Fb1rNyb5DW
ofS4/MdehD6dgfJweo5ZCqUa5mf6H2V74ghEd89NoWleVk0lFyUXRRjQg56qk/8w
irs8nPUcKrLNLqZS3n2UO146bkvRd7wPLNuIdVkItVhaepoc5oosJS0CF2DuJW1R
Dhci8/Ou/0R8mthJ3+d3kLGaVuX7KhwCpKt/KY7u76ce9Qz61fuJjK7D8fjOc45S
J/w525Yu20uZGTwlKPADOLGLvXk/GQtcsQtPtSa0Qg3fExox2rDnM8jhSPgiJNuT
WO1M3KiIBXRBkWUnOTl8NfJC8ieEEMJyFJG2bhDp7FG44Bgj2w1QXPnqCAZxSTRz
fVCdeXgzWr10V0aemajtru7VwNbCEQ9THDwMti3UZE52JoacWK1ThavYS0YKOE9j
q6qXPXNZDlrh6Pbjjv7Um6nM4md/BQMH0cDN3cUaJxCYhiJ3H9jGsETsltES9Y/g
+QQJL/XwzIkahSlk3h2QIXAkKPYS14a4bMHrlz7hrY7RLMtsBYpD/Ch1aFxEo4Ns
OMYMeClpLf8V7SORxhs3doBdirqbTJWQfOQy4f4HwYNssHH5C+Wje+rdSoZmW2oB
6lyWxs+WFyGkeEX/ShO7dpbRpt3cwgkHj5Oa0nsSAlefNZh8PQs8XKLfQk9/ZCYD
YvK2QYwLNlFIo1NCZS4rTJjgEqDy5y2NHykw+VsJolv+YxywGlranASYnGPx3Tnn
LjH3Av3eKwSezGHaqsNLgdR41GvcIxWtOTA5Fz26mEVwUTJcKpcnvWHufQ86Zuj1
HCwMfvGP7u/bc52UVm00DMWGN4jXQZ9ybD76atoUB4Kev1YhsdhQrjvGIxlrAZvP
eTIvrDWAUSiSCvhbPTPqk9yUFCf4DJDRJFIFBQ6mkB/pvI7eyhDEm/cWKVmMNvQc
ngoMFSAmTIZMaHwD1x2mS38HXSVHeG+Q574HGqGqtkyujSMyNTifp/ersWBa9G96
CF7GPwYsgnvHffTmtRTb5HHk4VumMMkH4b/BwEBfMHgW6cmI5KNsSHY7fo3Uo9Qx
/VD20VfCV6PZYUTWMntwTPPu44/1SsCyEBIRDie3DbH2iYLgvkwQ4W+WuuQfPfn4
LDmtNPa7Qd/nXrro6+aupZMkak6j6r5mwOi4XOmUNlRDP8x2eXC5gs++Fkn2Mu0G
PBrhoWXnHebiy818hjFCs7SXKZS6+o8X0m9itHqCJG8f104IHnxPEKkiq3zfoGTM
8AhdQ0/KjjKGWTS/QaO5zNGfo8bR2zBA9vYVla189Mt98Z7Wtaazv7kvjZvLPcT0
s/wzkpTqVu8tOYQBlbdLwqD9xmeGK5E+t7Y32k4KhwtOh4XPqSvRg0L9A9QAoizy
uJfsh+A2wsqjcAQ1MfX+CsXxIbUOGrYa3UQT2F0wwlH6QYIVnIk+fWAM5QIWH3XK
KLallzQBnwpjpZGdHPGuD+qIFA//K15/Bfu3XpgFBdiQWCLUzYK67cOM85ASYqPQ
9AJX9htHkooWUehWbXHWuNFTkxvby8OWgDp2pw95ROEc/+pdFhW0R5srVwHb53h8
347BYUacdk4nDlrWe3Ai3PySON8XfaTOPN/CtlttOXUY09JEGjzLYpvdzyyn3VkX
gUVOY/NhVB4QMnmAcxzUqW+UP1P00DjyhOjs4yjUP2Tm0jb+/2wZyf7a/QYU4Wu7
YkSN5o4HhEbxdDnpS2dL+wEFE4ct4YxNf7ueM0+gZrVrNNRrus17Wb12fP07oM9i
/QFVJW/IgMolo4SA3K2cGhw/481TfNjBVQo6xQxUIeFZIiL1Yqk0aypZ1m6wK6d1
9KMuK/Xyv+qH5ktGHa2Er3Ozn3KrsZOJUmOJCMahX0i6eXvQEQtjEQcg7mcHxB+W
q5u0ZKN1mIIvX6otkYsRN7uPFLwCVPFgOyse+VMEugpqvhqukjVym8YzsaxyK+mc
BZHsVBxaB3H9Sqonryr0+ManHBf8Kc54IiZ6Ytmer8max0SZlPJvH4qvYPDrjmvJ
lz4ujWqBuray8IRyxolQtmEnm+lf78w4B+kyKGFWdDnwrAPa5oMtaWBhnZ3YMZRm
e12/kcn0Tw3qc3VEhf7s27e0FKfzZdZPzcII8Wqk3zgccpZ8ygwHY5l86azOKY3h
TNi2fDM8nW3ll8AKNA7z5J0w6PWBlkDEKSHN+hcMAiyF7mV8RT/GqS7xagwDcVHw
PK3kCE+wuXFqdw2pqigB/r4dKrCqwqxZwTrvjK1rEYGvEGjRkSsXXJPpq2YDNTEt
7sd2ikApp68eDENMk4tYewgNTlRB1CrFR9yO4FTDRLef9Ne3W8g4lm/fd90MzQQF
XJnAn/YQ25bm9CF1balcUYeCekWSUz2lKcMbvml7hCQs2gP+M/KjS/h3Mr0/KQv7
IXLlSKz8dUceGdLAtg5AD9jlHp+DpYuJslf0pMz8/Z96dl0GLA0yY3kmHaa/W3ua
SLcaoRmS1JkMiO5YRU+VYlyKcIApuUJUm/4TKbcd8zegR8Kpow3w2XFb4isi6a42
pA7HAoy7BnLkjMCurpmhdXOELZDMuFeqhabOisrS8EtoGyJzWcQ42HwZ7xXgdwxc
rjOONEFYxjeGzNERhyejce4sksMNGTKM/AOWsaHR9tbhPMwDWBmyoOnmpgoQx5/r
Q6woqzfXCilxGa2UH196wXxrnPZ9YglgLDKGWYOpak8fMMlsaaq4bmGjli19Jtjj
4MIo7Bj2xVLpcDx+9lZCRPfLK2SP3jfWaqrdb7PWq2Vp7B8ykcOpohse4/6HI+Um
bOlPO0JEdlNBJ2pIU8l3bFEtakI9XEVs/9mj68kkdR2AcJ9ExOyLGA5d1OE+VsD9
y84KFRKhj+9PBfsSLdkS93nn4j1pS9fB6iD1CLpBHOys27J/dfCEhdKmf2sK13I8
Ht+WOYdaNNQV2OS1woy9D9IdLCJQiWukiSp+jieJ/mxETOLz7cTmqKq/lqqnbKqZ
KKMlwq94Opf8I7O+q7f6tzgrbqODwS6hxJADKMzOjln++FpC88C1Ps3Y16z7XePK
y/+9E1ANuLueGvAIFzwleOa9hOAnunO6di8fl5vvcTqXc/cSFWQTf4T126oEoSZS
OZjiJuB4Gg15QV+Px1syizsoPF+aOaAqWLYXalExPxDkZ5hVkoSsENDFI4BEa3du
EvtHaUQvnJQd1iUmtS4nT92oxWTP19NloqTC11SaVDooNPvQATHhV1pVTKRCsbvY
sGd+J8PchmrnlbiEbtNcnwGju76nNIngCjUn78KKAlcBCd+3dHQaUdtUsObiptOE
yoMxFduWnQji/PqVVLqhXGX/HWFE5ldzlDaGNxrw6cVnBKhF21X2ufLFJNa9aE83
qGJBbcn1q+4sIqGJowTeHaNoAjJ8yHMYXZQc3JW6sa6qW8wdoYCb/lPJSF9qlhyD
yGR2vrm3W6gB9HIlYwKSubRzErh6ZbfVEYG3/UogZlqZnAH6gNETio+WKQgaeoTY
EgWx7J6IhN0g1aKDgw1jVU2pc+EiQ/+vniO9P0hB2+9YnL6+x5OOQyFp7O4/IAfE
jjbRLJfnti2ZaX2tPATkPc4BAPEhlgA5qQTQy6kxo+sVCI8TlUE7+apiHZwuaoOW
40SrBzc0SSjYWJ6sSOu9iv1GlFz/0HCJOQvhwRSjnkZWWPkvgGaerI0Q/Qcm3OVi
WIEUnAuD16wxWO8ClgIbrALdB4temvg1m3xBLQGYLbWboQGOxPnPut/ud2gyHbig
yAwl8CZxZ4C2eAPNfvghTpX39XXyfPqHPl0EVh2ycZgXBCdxlqbs0+aPJAH/k5Pv
1S2MWy68TKpcc9lL+q6Wy5uJ6+DLKDrtnhpeczmm53IpxI7t0M/eN6GZufe0MVbs
lrRTw/eDuII0vVaT421sZH9DAQWYp1bNx64cNCvXEPvaZUpfHBmAdfL0aKn0/Ory
6Q11W0f1AJ/uIoIU0vORVRW2dvUWX8BnFmlGGZUdJ1SmGfDqEDhS2746g95YRbrd
t0/ZRLIGDgpFC8lN7jOmtXqmF9qF9WFRzBe/o6O6ABm6Er1WagqFMukdZ8IGPoZz
xyDdDR99wkhvx2w5cLijy6hioYPTAA5BgM7tug571PHkWnBG28LZWC1+zJbg/yI/
zEAdkR27OJ3ygD4T9kZqyNVPDbC7OYyy9AUDSzhP+3ep27xxsDe5DtPN2Km25Tos
zVVJsBctBrj4ePOG0iU03nheClniUfB4OVb+SeMXAUnoffT0EC2LKi3XDoaucXK8
4w1RR+1l1zzS8wC9kZUJfxiDv0kr0FDNCRr8sOIbCSqoM4kHMY81XqX0U7ksLk6X
kuXVvhDcAh9t3053FIg2BaSITvLWYGxib3vxsFzxNg3/6E00ZrenXvjR1PlBtuej
6pTce2RxB4LAQTuLKUa2GDoFKDd6K7c2BButlzVvAEIcY4W9mw9RBpodgj2H3mOQ
dDgNGV6WbVJcKcny7jptSVuk9owZtyCgQ4uOTbQwzWETa20QV+VFczBWyEz1qyOU
q+4+Fy4tH2c9HhavOrr6YXVhO0iOfjIVtL/OHAdA2x7LDt5y8hpPY4A1rvSaWYRg
rmb288LCN16lFW+9Km3XjMCF3gJBNExhR/YRUyhs7xZgzIOAMveGR3ztkynyAiS7
TreyzpUuZIkgEyok1+oQAy7XHpqJPfKLrXl8L5HR93YIyhp27kky5Ltm/lN0YhP/
BVY3rCrddPupsa7bH2HZuNdNunHhCUX9EktEH7zkbn4jDzN7HT/inAPsPsrdeLT1
40r22cikSiVBhYYqdIUvSBJrHykEk4XJWVBzf/fFi72WGH59FVQNIRMzEg2etqk6
dFwhyE0ptOLi9EE/hzcQ8GAZsqK/JKWaDLvwRIGqMwnSRfvQIhSTsWGGEIEOxTSQ
gztLcuNjYSt9HdIUCnI+GTx8z9FpNurA1g3Me077HVM4nIBRCH7hSfsDvJoDHuw0
mIRVtI9TD2vwNXUIZzTkFiRpcmFjTK4k/I7ypFmDYucJl2ODIZQ6X9Djq5AsIRug
rXBLoNk54Y6UbVBegkAhgqzVg0X7vQjSSbcCMAdpB0ak3UmyCLzYWX1RGyNzFN64
jgL1iaIDw49wZcwhsJs8vxBHOR9089DtcLdzHPahvfpD2kWYgC3nGwA7WRu8LgP/
G6EQH2YAc0nER2ENmIChFjlmZ+/Uox9uCZx3yEMkJ1EPGOLHVo85VWed2jGGDvMP
f5h+IsgPaoltYPaa5HuxcadP9Q6tJnbAQNOOaB8kkPgT1ePW4yVpuiPjbvwGDvB4
IvwgtGrxrOYS/LpAwaNIa0UzReiFuHue8zmYKsQVtcD5uXry3If/1LgPKjTLGkUI
BVr0Yvw0WeQ/Bron4m8N9/RCsA65WTHuf+fTbcRnxwXvIVwSLD6imnSnU6Yrz60V
7oU/VBnIOfSgbhWRSnDQa4aN2wgxyfJbsuLmI1OvrLgnUk76TnHY9saQAKR+9Cb+
PWxRZz8JJUFmBMRegv+uhu1YBI+SBQ7cFR8dgQLgh+/rlqYFP4t/xIBO5Yo6AQBF
sINNj2OcmEHG7+5Dq5S+dVUxT5OMJo9DUwBWhCay39N+DTeu/+Z9olObdLpI2trj
ajLir696JgNmSB/UWpfmpySEiBb2GhWRfl8ecqwaDeiDlpOR4JPu0MFTyL05m0HR
mEzq33agNBgM51Sxgf75gg0dBEIWs0xTWCFvtHlNLx3ZHQrLhORcckxwEFaOx05A
EMPrqxLhZueOThXnq3OSopNIhwv8qNvsKNJWYot3H+P5E3f788G+8nrFj/TiUe7H
UhQXuPmJfbvbbI8pq+dhD4tyq0mUYWVfRTDw04xJy+AwT5chQhUcbkASUCOeYcAp
p+AykgsM0INC4itaVShl2I2oh0L0e3vGyrxMzr9CzN1ihJeIsdzNHm3rVrceMcPZ
0A10O2OQVcAh8WzCTKfeKnCkCELeeJPzr1x59knHzYzYoVIZxXObrnFsylMcjaXG
HdapFBm5yo8fis/Zjlfju5ez4mWUElcDHvsmCNlzmk/uAnrwJjX6D4Od/rVch4Nu
sqqj93WAAmLvepL483PhnLMSxMlK+jy94OhflS57AT3a+4Ucyvs2QNzuwkCufdTe
jA18sJ7E/n7K+jAJf4k6VARB6lrO9LkoRjHHyQgmG8arxkmioM6nFxLsSiJv58ZG
2LXNhbdxodrLqr1m6O3Qq4uv2q+7DZy6j9HVLoGyJ/BYPeHVpLdeLB1qhVY/1Ts/
IbcGW/4Q7cpg3qZi2b6RZiWGdq2hPCoHNKsngM+6uUIMyL1Fn4B+7JWfG4gLwGBo
UJtkVPm2QBfQS+0sDxjS4dJCJTEjzEEsubFWhbhYJVB5ImvzB3+axrneIctEGz2w
9u4CZZKFO2aujOvBlVVKoRQ7JkCQWaKsAmpRWmamlC34NlFp89hysHyAWfU6G3hx
bm0ARMD/7i7BHWd3YPDd9QPWSU4LhF2rOdMzJEZkvCz1usFbFxsv/gxmsTFOamRJ
KrOMEXOwdP6KaBv9LpLZT1hJoLSaIuRECr79BjQyuOQxPWaMqyp/j3uiVf2Fyf39
K5wbwzQUHrfDkUWAxtxn0GCyyf0ApGT3wZSd9f58Dw++2mnCe2FY24XqMAICer2k
BEKT3muEnqhL5Cm4cL21ylfEEPS5JhTPm1fkR8HBrul3R40UvBMicQ6Y93smism4
xvG7XIVglS/1lh6BSgvwXfh4K7vx1itszPLAVTI4CidLKRNaE8sKk5tF09qb3YHI
zcCm2BDIYEAD+kFS49GmTXfBQds3d2lUoXQUQD6bVCKyhxVYV0KKgp6zwa2s7Bbt
NCqgartXuHKh0uJ6npSEfWjsShccaQU6daj1Bv9W7aUcpto4CtwD2iDaUc8nzwQj
06WOWjyAIDZQF9vk/QGPGYWTXcUgS2tv1vVCkQcAwj2+R/1/PHWQ3pVzgeevEeoV
7GYk4Rj5Xr7lINRriKb+uqFsFMbLGr76SHgA12mC6SyqyHAqqXp23vTNHOkQURuA
qGXxbvSkh1BtKxs3BHgSQ2MXoQPuRYlCpJ3g1+FQP+LI7b9ISaeNldbj7ho+k/l5
hEQNEg8+Lk2XrMsT2Aj7gfHKJOpOp1Z/Z5QSEw8I2W1Z8GodJPEi5sXh3y5IaunA
hBV86/R6UO+B2E4DP5GeA5GSEuFhUKiR6KG87Yclh2Lx2ch/0VgEiBuA0Lqs6Vxd
ZsNK9QEjASDaPIgbTXCM03dppOJ0L1SjKsGLtvUtDRxCjKW/dgZpC2EvYbQ8EZSe
x01+xsltqmxnAWTnZFzjaY1ZClvcC0AokYodUDFJDUpZ9+h6F0rGi/vxULT4rsPJ
PmDsvcUyOg6weR8HySRW2B2mZsQMpvfJ7Y8KxJZfDiCECafv2ksR0+nuLxx9SYkn
uZBjmJMYzcqSZl3t9WxAom7Whc0VvR8Orq89fRXLXFi4GSSClPDg1hBYcEfN0VgB
JXgCXD3yPRGzgn1QK2/KB09nrTjz4LMrwVZvQak0ZyT3CJyet2WZxmPgiptXe90W
hZv1XUWMWP217Ih9CmNkqYuc98bdJgOa2iq4eaVpFLu+9F4D94OoECa1XFgFPzaG
hsMVubnTa5Y7LTtQilzCYowHycSbJd1vF+CB6TYuXewcarT677mC48wD03EhX+sU
3gCspvzcrDzhleQiV5PkVtVDW8Uayd6NxEUk0cumJQOWHkjfT5Ggdq1QTzgnPKwr
vArEdacMXJuRc2I5xL1I9e4gVAY3PkDe/8P53jihDHB66UOrIqVYb8FZf6yhl+ly
WlhBGZ2Lxstbus1NUcfr0SdDDwqx6o9CbhJ8h0x2keIxZC5oDAGausV6QS/vTMYu
emBWkx/4BYHVv4DpPc4PQcrrxGrFo0aYl2fZBEGHJFZ/FHypeuNB+Lpw9e1Xo6QK
e+yQwu/M4A2dRP9pdtOFhJX1SOaMrw5pbV7UlcdbVxkY8TVN/+RfE+44MesJQzu+
0SRusS0n9ISn3ddN8Krf6U4aC7N28t1s3Oo4V/9nCHPYxRugTlpX4qQN5nCx8H1q
F1Zeil9uacrBi5aRVoR5Vd7DvWxj2Q4BP4x2U15W/ldHL28K2SwprnPGFHZu2lJa
+g6u9tiE+J+gSS6C6w6AhINikr6fM9LqnWecT9/iymgzvhI3tjw/AoTa4IhBqMSF
vltTt+rSkQHfw+/TkZWaRxDj43/lgpQOiBJ4diBAeH2V6Z+dBI+ZbWE93g1JzWWx
jPzIEdJE8fYKQaDM4HuNsSssEwiTOasP/OtLFlVi4Ih/DBkCGo8Q6gWJn4MccL5w
oYjbGKE6rOtXq7IZkcMP/CoQ118wJV3YUWpnLYD4L+X8By848OjK+KKDkc020xKD
8G8vXMLFlZyljvLbR9AMwGNT7nkKLV6ijsasLdJongjXneqY4J+Kp1fcxLTD0H1v
QJB9TJ4PSQ1irw98PoLY9/C8mOaCNpn6MHqdWkvu+1r2fqD2AHkxDw4sUmBVc/su
iRqWzDtTO7qrBMxx1ow241cz8vM0fl1CXnapSPWWOBOj80AyImOJcKc7kuItScTK
JWFxWYS+A7E2RqJgRtG+A72Dgi0npsfVQH5eMbVvY/yf2fAEZv7nku2Spa5wmNoT
H4w6cl4Z9LwbVwDFGOG+1IHxB9wvuiBxI0waaWUK+4Y8L6naxZGhRRR2WvC4Un6I
k0Ni8Wq4YjklULDMi6Ho3V4+YcaTG39XH94DZMaRDSL9zvVcijxdPFbdwxwxFqL6
Zm7chAW+c9zU2clKc7Pl+lFGrg3YeL1V4Vgqo5Yh+R3rSxxHR0bYyrLw2k+G+9a0
Id3kDMBI6FvKeZteGj9ki0juPc+bxtzf5Pl0dXSGUp2oDQQjmyZygZrJ65uCO12w
89kcmHrTTvYyoi7psO9fhVacLo43mVG01Gz2iIuVB4O6JqFzNpSBh37TxbR3hN5O
P04/zylGE3wX0Ej8rbTMrWj67AQ4suNqRrqSfuL4WcYhmpYgirT3MtBKZnHgQ5Bv
dguJikJrH+DOPbRVoGvXNIyTWRVtvZ2egWrtsnzvak/AQRxyPhBdW9vb3IC2pGuC
D8W3lv+8Q+EJYLZ2FDSTPDiyD/9d0NwIZPrlnMT99g9gAtwEjFxmueLWkDjbiwf3
bOxat0WV2QKgPQ1DCv+ICOPjsZxPwHatLFIrULhBANlus+qdKKT+dP8nakokiYOU
YKnOoczv8Zm/JZpMwo9e07UirmebufRJF7V7KWJapGw05H8PTb6ISpuMvRpe/re2
NWQ/xytzO1gcvMCJG3muOzbmB0a+C3nhe/dUrxE0gcSQECMttg3Lf/grvHG6Kkdp
cEeQoEDrCGY6TfSKA4bU+sHZ9I1PMiUVbp9DGiaRQRTCVwZkewA5W51a/oA100lP
gKIEGlO3Rs25xVjuqOKh6dGaNbzJ9GWOPhXDz2pvmPCs4y3qXpXYT+n++Ec+Jk94
OC1B+dcHcznq++lw1Gzah8jgLHNghq8bQCGNr/HIvxJ+/tEA1M2NVFmGo+/5sQp5
SRC/E0cqz8gk+nrjpmcXGhYKm8rpojxj7d4emWuFczi3yWfKj/s8cY69MwYLoe6Q
zBn7TNuF9qPeH1m6jct0q2ZmCMW5r6ZRUHor5GPhcdCY0gU+Cc0Kd/c5TgWbgzFw
P6dzbGXygmY+bB2H1Qgh5oStpht659DHyzuUfeG+NUaz2rzwjsPfe6rF0Lqj1fZn
Wbdyba8K6CtY3aUUmCMOcqxPmQjOvXfj9jDReGF1J8anHBM+9y4HY6damq54K57M
oNY0DD1SY3z1bilkeFI1uTAKLGEEe5EDoVcVBIPMLrWJhFMB1q5JQPTmmqxJuGEr
f+zuHUypDOy+kX2prw/imr6jnlv01SX8/Wk4D67qg8gUe01JGV3/jrM8gyhpSy4j
P+/vIFhKBrGgZtm3Lkcxtgwith6QwyHdzVho6lDmOvSq8k5Cus6VfBbfD9Suci13
Y1Er32AX84X/2iCZH2gGEjLjcHxtL0pAe7EeD5F6S04atP5DfCz4zVoZPXNuIdwF
vw1WtZyEhC1Uh6VNMwyyVcDig/NAK51Cfiko3McBpys5LMoEHllA/D3zaliFOqq/
Cs2OF+ChyVCi+hDc0b+JDUbam3u9cbS70aro18NjaeOa1Lg600JV2VjU3E6ajcJ/
/gg6yhYtEV1pf4/DqQkgb8iF28mD7LQQ42D35p1H/yPB9YoNL6RPrmfuvW7zKief
PClxt68mCHyWZVz4+Dk47K5fjFAfeyvPqqnJPqyUGX37rBsrRRfPGO5bK+IWmKbU
CKp47GeDvq6j89TxCGYnmR825vdRYF7o3/iUbj8bjtzSkLOtAdUYf4nCktQ36n0B
mH4Q5lWblQf90Op2A7UADPTByGjJ5MGAIkiQ2mlZT/hi7vZshb8BKVPpTXDYVraG
sOGGnV08nUrjc13c19m0f86Nl71R9lNGzRwSxFwKfv+Gp6bepd7IFMcDemiEV7rS
XKaJPnedNaLECRZy0iAVgBFF6VVnLfxKnrLUBbqSJr1shhtFyypLcJN8A7M/YiQ4
r5rQHYLB7+TVy+jZyzxeJE46E535RhnnKrGPFnHdxYEO9HnbgpRxuYNIzS3lSEOR
qqo8COP0dogNsBmI8cX5YcBlvT5GXRD1pzl5k++8GA34S0XTTZrygmt2OwlYYwPh
MIcHCcefpSNGXJ2WL+vagmQOWeMXmptLVPAVfzJ4S0qmukBbbqKTgFeAJqCRa57w
VmSYWUKXhO4o72L6X8mkqa7JZyQ6t1EbVchfmM99kxyx5dUKOITGuqc9cXq1uLmV
KedatffHOBClEAmpw1GyuTVuFZNdiyoBlzlavYnl8Y6t3bHGZb6lCrf4K9gYLEKk
KUcYwcP040EI1ymCWS9/5LzKYyRFjkAxCJN22ZoLXHKmc0AD0C83+/gyr22pWRXA
+/+HPXhuiKk4Dnuivv6TGqvTh3gAuoXpVXzopCgB4zuZrRNfKKqWoyyfPmRE96qo
pZ8DDTNW7p7I5OfJ9rHComh06jpDnbP/o6Z8zYCP7YnVjYCFWJBVpPeIxJyJuQGv
jI56jwocs1aqSUT5Ne3anhSLvQAKsBXh7gdnz43CiZ99PITLmT8JamFMJ5i2KRHl
0rlMP6Zuihy+W8KqhuKptNSVrN0BXOG3hOzyooyGtagRuq9AO1plalTjHtzqQ7mu
WG/sy/yj3Wkvs3dP5jWcEHb9EJgd8bO20cXfwng5qeBy536Gj6shloHX2WremMJA
TzVahNj5lf4PthFZRjw/v+dNwa7Ignznmf93JnY1fdfBvC4XX3TxwqsdIWdOhRlP
U5M63TmkM+VdTtuyU58z1NOcvWpqwKx1rnnYUg9ZmzhmBTfEdoDluz9pE/dduYby
tggDzIrDkbZSEtrp1NS1BKeCAefFuvRzgKQ/dnsPhvtBXKfLBuYHdbThzpDl1vqx
Rw08CvX3HfsPGgHO3EfNEh1PmYsRZp+UnTY14nbJNu5vh3gO9veCjSY1Vqx6Y3J6
eW8bRnZyN9FxATgqUYRM5TkWcq0mKqglDqy6O0a6d/HTS7FdX2nRhYt34McPATpU
Iun7i6yAEU8RVOix5tCi1RBDQ7vQW2qgFsGpke3B0RaAX55dX5eKu+IZBp693+RN
uyLMjIYeQPv4AumMHitm1jO4WRwTYkSH1pfiBGwEXTBvqkfasmRHFKFUXQOFwIXu
anTPqqkWS6wpuvJCV8qAsQFQ7F1tyhBQOkvsF+miHP0cvYYlkmp0B0ua3+y7I9oy
G3eV9iLplL3er9KMGBWSXG+HkCYgFTBcAaEpPewQpfkcw4poIdQvjofsWyn259AO
FrIpQhhikBIECtH+bFq/ypuBvVJEa+TiibpAmQzfFQPg+SjAtboxTvbPP5ZHXt16
Yk+1P3JKN11yFweBki9TAxtr3BdtP8avpiZSlU4m4xb1FvIwlRHeUqVv4qzgu8kD
0+pc7zyHIy2leVfDPIWaPQQz/UzHERMhm2eMsuOdK+3UXA0oqzf8KAoa/tEEY2C1
haUrOxSnyDhUMc72hFdgyBMn91/aSam0X6tCnG4jxyFww5wX1/blpfRlxwg1T0kO
lR4mPIizRavJiwgiiq3UYUKy9VYYjYgztZmzyvxB+4+YxPFXBtLNHIRjxa1ieu6J
fdhxtRLcnrPqSJFeR7zO4N5V+pdLy3r475PvHYbM99uJ7+QycStcp3em2TkMRZXR
DXyJhoj+qXzRgotb/lWC6Qe6J9uZ6F6a+vFkRxEBdwHLaCsa4n/23xWkIZibQcgl
yKWnirbbI4CmIbvRHT/M0Un9ksrdOHwMx350AJIpaZRav0psbEauSpn8A+sv3UIo
yPyqOLMMj+0MKWMbAp72L22KP3+lilKpCvXjcmzWdet4PVaWevnJS5Zo4LNZqB50
MXDGj5sGTKefYI8EdDxkWH9+QpnCGn/Qb6EsUCJyYuhm8hKRHWEo8cqg/IssV1AN
6DUFd+itRLfGLA0qDD6rpv/Iti/Hoilekdg3lrqdG8SaF7WBpqVTpNdv76vXYHu7
ioNod5b8IOyNd+CkNYIhKp/YtR3lJVtilsU3F0Ql++A7/eYxECGrdarIJwyzarCb
YTGyjtiIBIq4frqs0WXACFTJhbAhx3HF/vTtYQcepVevYX68NycdoPle6f/Sk8iG
3Ez3u7qyjjWZD9i/v/7XZ9FVj5eXj+pYm0sp4Y5s3M7U2cBvLKqVxD6OIHoehmf6
MibKOzYfU8HL4MuhoFyJRB33Nin30lX+gLLvNTapuASiuLzzqLsaqWm7IaBX1/ve
o8uaRPuyi56k06vdKuWft9syr4TRAP0iuIR3CnCExHWV9hjSPAAEVh7L4HnpGI8q
1JWTwyrOFBsdaeZTacYQ0nyEk6z40WMcPtdQGklfuu2+5xsmxwakgrZsCk60gIAq
wEcbxVZkkvwuxXJXGliMMACxIjg4i4nmLvotubRWc+yVetyTWYrqQij55AqHdhOH
09yiRN5iUzWVi+ARxJzJLwKEtuztIdNL7r+y+D0hV4XfAramHM4EhEOdkb72f221
wLETbByDP4jjHWjhf4eIDnpWyllQpd9Esatfu5hq9LaVUWQbBTI9JiqpGsOTZQOO
KxsTTJXuEDJ/HGI3DkLvlyPAU6ak2Ii6mn5Y7Pex60Yp1YyWVU9GnhN4RTepEi2a
CKAkX266p5p60NEQGHloU6WZckRGjML2zHZZEOwNG+Om1EKk/snBcmtPtUac2vyF
bozOit4MczmbxoAsLgQVyeLNB5T7n32ngLVDteUP3MW1jMZ6fs8crq5K81M6CSaW
ZrHZvWaTlx73MOA61e1A4o6rpTCJ4yl6SQsH84fjjP2fZhjk7Kq8mzt1UtNggplJ
J71K8BgZg5yNwdZ+LWceOLoTNmpwsDUYOYELjisGeF3CRqHj3cs4iyIFIFERpRUD
RAjjWzJNPerMMY1htFactK1r3Nf9rNTPRsg8NNJjT8UksTJEmzwjRKVcPkdw00U6
QWESuTJGDPWliCFB/ScwyAOIs8YpZOCl5FsisxfFTlU8YdbaDg4GvC38tj/mpA1+
kv5L8t9WQnElqRFl4gjvkDTo60RjQHX+/l26cRF1JfRR8HmhfQrzk3oiMsgTwaXt
gNupv83+eQJhb/XNIbPbHWTozTS/sxG8cx9G0S1YCIeg02RRu6gT4k9MKYxTp5Mo
t+YRPKElJV2IT5YatAcnj/bqPAc5Kj3VS07AivS/t1WAKSVr2RmZTlrI99FIWkCS
i8FUGxHbZSk+BMPfb3m66SupWLcB5jbjb+uSvKjfh6A4le0dgYhiJ4ga6WUuV3mW
xA4GTXsSc6zwWD+v/0GRD/YaM59DxsZhonC7aP8rUXOfw0nfhwMakLZi10XNj+7v
Sf4kbe4mKYOWoBHOTn9gms725JynyNx5RvxkEv4967afShUom7c9S9xtPx10bAGw
VJfcNLvZ9npn2fNbCelVH09wbW3h+ONui488VtwrvMmvPxgo29gWXasIHbXmANEw
oLh4++8hw/uI9WxntfljWW0xtXvNYZIMuEr37ql5O1QYuw3+XPpFQW1f/twIua3/
zWs+rq3lg63HLUSGAikkze1nqGsOQaplJAi975aMaAg8siosia9lHUheBEP6lT0w
gJ7T6qYAN26tzC2vKlaVVEMT5Exlt5I0o2lERJ85zi9JlRR4o+jhHORXuOZW85Wz
5s7IGWW7sBaoikmmFXht420tZ+gEbLOQgUlhIN1KqB5BfP6xa2XYTe17v/0NNJvr
2itNfBdPKHw//h3Sili29eF7KTa4YuR6mYAgCtiaQhCZY24nglXUqny+r6XLjXgl
ouB+XG7e4PNo1gKQK3SyNfLQhpaDoTImn+blP1uUdMFRlOIDjaCrC3eWIQtb/Dbz
AQgbhhzHeIkXXdcjJyJPEiiyo99zPGYal7S/t69I25IrJCpWuEuxyRhEDT5UmodK
WEn5rgyeC+TGy4LX6qxmH0fus4kgkJp7VoT2bHz2mM0KhXz2Kc8cztV4fxcR9uI5
/108FyU7NXjU2O0P1oDRCSmRbiM4NwYwSLn2mQO977O7zI8YBawnS6bBsgPTooir
maAj0HNRLGbiNPC8+608NFPjEnBWnhEcReoDBbB0XM5Yokc1qMoW1uRj00xRNZSv
D7EB5pHiWbFFffgnfIFmXvCrv7nJSfwU+BH1/snA0Szudo10ncwbMMqCKxfJnHME
PQYZuf/T/c9VIiSxWDNNdn2ROClQwqLa248fYcvoOLlntVIK3bTZCrubXAeYI0Ag
6Ty5LrEZ2YRk2+Z2XdBUxy/x9CGpYUHUpqXdCZv+0BFso100b5JYOkU8Nqhj+34c
BCu3sqS3bBgR8tkbmtvxsKoT8lat5mV4+pcdWXUSzWx8c77fPdFWtIhEerMZNmPd
cMyPnhTn4XLJQl/UA0iV+AepVcgmH1dkegiM3S80ulPmGBrxuO7/FlE4owLaWQvz
2eEBL62ftY4DUQCPwe3qropYchpIJ/j+z5l23l7iJLWSpn6Q2/WqMfe2/iEdPNbk
pK2wGF/oLWmgcxiR/5fh17WwUSi9I8bmkhRIixk0jN4jXQIxhpWn/c16rxULWlpL
tzc9fqKXHBrMN2ObONXBoRFejj/WdnVkxa4vl4FfRKA+RE/oIsYVXfwt+rOJwkK/
gPk3//VuWTrEvXj53Pj9+Z7mTa5Kq0KEOtNWoX51TrL2iNSEsdfbdJOG7AGMtWC2
dyn6vPeZkgQRvwBxQ8JPZ3aGGR2ZaZ4lGW8QhLobbx7h69ypJjkvpkVbi0fz5jGW
I1zjpuXs0vlECpPVTmAV5Ur9uRakA4eXHjQXKCFa953T7WxSkw+9550FlkOCGjnh
zv0Tc+0XOgoBS5Vgrgo3rQH8JLL0FuABzh5EXZPupKzjaYDWA66QgzalxpQdgM/h
c8APGT6Bu1PUQKl92FpzYk9nXLzHv8Af9FFx6/rBIS13YS7anN0ZbwAGOwkOoPq0
w0AFMxwBzdAItXsveCQwnTgpzXuIKKQywHBbMm+A/avqbbtBGf1FyIG/Ig152Vl4
qXnQSdTWi0CgScru4jJ6URorvtGWPOB8FAmJbRgZnkZqjGcEJWv+5kHZjpDTxenG
Yq1DXGZT/E+LV4wg+qSTE8ZJPs5OMmfCWLWRIa/CZhxuMeZTSIlIrU+bEE4tzXrS
2Qm2v7erC3bJdGqHkw7Oo+Syr9+vdeCj25HCNlRuooGC63Z3NeWFsQvpWhLi4EJF
S0pbpTYt2xkqMaIi53riDrhVA6niE+vhHvez3EcaUY0VstEwKR7BCroK8OihqPVM
SNqDL5o9SsadrVCDPxufGvLn48BIAwJ2KVnsKJshUtOcLtDrMTz926NRI7HJeZsA
G3g0t4Ez894/RpK95oApulRZ2qjuo3D20wtYFGMxwBVxxan0Zy1Xa7bYTow0/+re
9ylXjHThEYV7mI4gzSLejZiFVvNlsDOxUgKKZNfmwDlQeeKmEh2RHjbinfsrVibT
O5dvtRCyjAJo5I6PGZ757LeXSi76+PQbJYCssnxSJ5yzBHvg00TwahU66K3B7nht
fSdYcLFLOAWlR8NB9+SykOZEXPaeMvs9i7TuIst6yLd4qxuVzNTifyVFEYtN6lS9
Gt7EiskR2yBLI6I19NN+iogP6NF14frDb2Gx5p/cKJUyEu0C654R+MkU4ERuodm1
lSC1daC65gN9HKHMUTZvTXiSIqw4kS5iakG2YIJOJTjcHc9W318Hstd7qTynOdfM
ItizVAzMIXTidMgZ24JfP5dFixjoAaeAgl225rLlheI0tcB9FWdng6dvaNbzWaQm
uyTsiGzHUBCA2DqO8kBzosSwcV3DtwYDyINa9e/8D1zg7C5H9UdbYC6Yl6Xx/dfO
4BdXARN3RYf9nqY1+lciP/Jlmknhf6PJaCs8NWjEecmXW1zxGLYAW9QJMP08xMG+
QuFb9vP3ulQNq41PocwMqd9NbgA2ICC95ZnxVc+1cqm1T6NzNXHIbVf468HpzC5K
KxZEG1DiweVP2nx/rTItUCuFDCUyhL+rnHacpwiW/dO7DkWxnUyToROWEs272n0H
y+mKgKUfs5sGsqtO18QDeQgTAx3wlD8+3yffdLsl0hcnzAb35+fkgCOhFrCZzEaL
PVM0B1y2BytKaczyP+S6HUL8PPEEAtVZKXDS7NUUW9U180jICUWhIoe1T+GoW3wW
Yun0n97+3HkRdntsRoHQVLfio7LJCFGDZ8PCW34mQZnJOfPF+AondmmVi9BHZhst
t8RA7vDnppSuHMWDpg+6tR6UoIB2gYtrK1RtrOldslBVsg6eYFAN7OSLMBftax+X
I9lki/fKdwPgNxmamkp0cEGm9LtBJeiFPFecruSmC7aFXlsiDV6yJQwNnrkxnFcO
O2v0Nu5Imv010JWLu58x2aAPLZzXihBSHcoeUY3fZq8Zr0ifFHwcUPYDGtNFa8q3
vYk5mgsbF76RciFzqmbunonH320oEB7bZUoisEOuu+WqFIj6P58Iz0eJ2WkixedZ
yYOs2VmcFEefbi8zjDAqC3Qbyjv2+M+eC8iHroQwsadbFPHmawn+uaIf6L85Euyn
2VfDMOWI1is0pKoeKI91dNSCmT3CqsVfctfQcV2JPGdBcw/itq0EW+3XhlxESL/y
DopVIOOGwiT2hJT+s1GkbRmMBlhHMo/+CuflHQUD7z55tonjfsewsNx7QGvl9YBW
hNwbzPk/7khj+Xe3p7ZVrDRTFgGpx6TMwItojZRgujgvkCgCc9sXY+iSirHnA1Te
5PWFyl+vMry46mR0UgSY+QKRBKxS/IzWidUsoojLsKAFsV6Nss6/Wj3Tur/U0DbS
sjsTbY/txUnJNydQQXu92U8f/b6HCKWQC5scz5WF01z8TqYsv4BG7cb6nBtWcBMV
rAyLFKKZkpcypUmZedMpfkPU+hzasfQfvnLdZs0kMOq1EqtkihAukSmMOverjfJu
jrMy5Hv6J+2IFPiq0dmINfbg4+JU0a5S+KRka6mtZwmzcQU+IU/H3IAGZJYT02JJ
3WDIfGitei14YMvRn+Ym+X+yujC2mhZXvfjlJ8+S9qNvkIOzhKkK5S5aMrBp53oB
jGJvi3PfutcUvYFyOwP830wOQ2bI4eqY7UnQ4pDQbLeOQwEdHVGL9ylyF2kiOMMv
EJoh9cZkUUIqpnWdaZkykqH/pp3RaKuqXneiKvOqQZHY+oEwCnss00geWI0yKgUa
fIjA5v0Ua97XUay1hR7ruYWXyXiFMMtlmLt6TJvFSrDhSsWqEcK8pkgybnJ3HYzI
g6ccbyN0u3esHp9CmAqinvqd1MZTF0xm1arWCDJK5WEkJk6jaWbESgs4MmIB3hlE
escaFvk7wu6GRC5+HMfxw2tlZfI6hTSsqd61B0ffFkM3I7littwJXeXdQ+RWRLAN
jqg7A10X68qAgsCkmIEV/4xvqGmOLWUJzTS8UQ9U2AwCN5DVodYapPseCS12ty6Q
uOlB2QqDmHQXeIlyQeQBkQcT+oYw9Mp/JUIiXUKEusM/VLrhGZuoksSut+TWsr0l
Qt9qMVxp4vhk+3RMUhTxBgktwbPyv953c/7pyCak0+frqRT8MBrFrs/3540VGFzm
fDGDvf14HzQSqiv7k25mIsj8D0raSwzptkYAhS2JeT8GuAJE5X0xyCeedKYCxYae
rQQieXUBs1Wt75k63s11zEbs0Xle//D4PGyRliBv4e/FO06n8B8ot/brGIBlSM0W
1kpspSPC2u8/PIHBXmNkdPot0X4tOLBM/z4GiKhx+3tiRXRZYgyC2qys1pOXQu0N
5kw7DUs60oV6Yg6ZVE0HfToZJ2FBNeWB6Nv+zTY3CJYAK3dKuK6TpHAWD6jc4qOr
GmCXzNGef4yhvec5Fb0hg1mCQqFtq6zjEoMKBfLoUUIhJV4k9GEd8rQ4eRoo1j+z
uiip+ImSnTIUZ8oOLrxF/jT+NV09mr4MQq6e++z+DxX//VClG6HPkvv+zOYQZtlq
0ZI5rFSP04XeHvem2pTFNBcykuyCfyMc5sFXnM0hoFmRz3G9PODC3ofwk6lwfOkp
TfjEfXmfe460jIziMrk/RRRlhsRQLXOI9VvORUwv7B8U+gG4j6OLfx3cadKN5hKS
zBIZlX4bVtuu3M6rzWX+4VN2h6x1n2ZxzFmz3Q9mOR2rzj1bI5IkcriJZimaxDri
eGYBjW4MPff2wPHieH34y9u6OeXnyA47VD/y6pfxKbpjECO0MM2TmQgFROif/3Mv
VyhJw00GzP/tRnuCg8UY6ZLERU92SisUprtNzR14LePkL1tjDP6ROoI9iU6ezijo
upsrbhhHyD99RA6ftfDBvYv58PxNyIqMq0w2JsCYj322PyqbOW9Y2FuW9yiDMAHp
g3qQVwAokXd2XkOHo1/zYnFUWhNzfQov3ozwrPI/H2NhYWSMeE+s9Zd8grsPPLvg
QOaI21iZWwJv/6lL20vyStme3uchOp2thbTA28zraJtBd6zVuoTP20Hy8yjAzzCR
Hou6cMaveMqecxSvfILHC9bWt3iD1Hi517vsaWLXu+90KrKBMhuOiTLaL1DIERl6
aiXJUHO0qRXKCio1oYB+xrE514HhD/mSt3SykIvD9xhpQpE/HD0bje2tEi96+BEk
788gt4TICUrKhbQDn8lJnRLlbHXiCY0D7OSX1ZnYCIJJPj9M7ZW88Xybwu8womEB
q4vBLVVeyKXhA3f6fgCGusqKs75v0X0prvgJ/tw+ityczBfsdegnsV4wPG8I6NbK
AQ90/yPRv9PffSl8iuepMa71GuA1V+3fd1VdygHCwBBj8jrPemdbkiQTRn6v1pm/
yer/E94T4PugVL8BddyaCW9OwIGExBB4iPO0vPwquGjGkDQ5lSxpB1sb46FmGf5b
Ry/kBh3a8u0sgDqWLlthzf0T9Se9gzHJ6tUw4OhoceiLxCIwPFptW+7HcsLTOe99
Od7qDw/1XqY2aLQk8ZDNvcT0DmPpophhxpxoY7J8TlCqO4SKcMAl0+rZSNt633dA
/Weu1kesjYPhbiyjUKLLjj5g+N6TmV5WtS/A5ajh63W88aVHZTDBe/XMtsJhMn9F
7r+YcRAx71iNQwPXZMu818LEbug6dubOvvW+T3e8oeRILaG/ALYC7WUzbv9iMphd
hQJ1Q99pKz/nv1xR3kwdqEeaYb/SgoxYcdvxXcu+Yrx9k/RZTvdIayK5RXdp31yq
QRPlPmEgcUEZRIu1wfwHr1Ngkg83YZLrG86HrzQRuOspjcpz8GsO4SSsPvcZA29q
EgU0Jko6jvSJDNSySKNCjeY9XdLBMdUx0kewU1wfvXOJIgQuXAzQM47Y2jBD3mqq
4PI9x01TBY2VAQSc7ZGYZFVIMfy1tiaYnU50lRJNO+1SKFIwXNsJTVgNz95M5Z+v
yi9B6v8jpUklXjh9/nZ0o4xKFHbIrOTd6aH1B791VkDDo36/j4jR7UYVaqubv3Gq
MfdczCk5+lHTXau9qwDHpdlSh57EmtC/rLTilx5WVUiQBvQRe8IoH7kyZmb+7Sdk
V+zZdTzuMqcllTKFeLqCMAjfU6m+AUJLfKvLasGpU2jFdCKfE3AIWdlpx5ZAA5Cc
l7r4y/3SqS8ruUpzdj/egU2P2Es/quhkp7ahk0M/GBAKQLer/UEsim41Kb3SC5g5
6dlw2RcsEsf/AtR33iGXAeUcNV5nZjjIyvu9OOfWesie1fFs7d5uE8HFzx8fgicQ
f3vqEPWapgEemQaO5BqU7IxsGZoJO5KRGn2tye+GrsSD/XiGgB984U6Ufj+9FOo6
ajiWOfDxtNElH190dvFeOGpKZsAykQdClwza0UXFTO+i8sfw2xVVNesAn3kIX3qf
K8tkzIakx1G0QqU61uaG0zo3uQs4FHc70m+S78iCWx9a0KDjGr+n2g/MRebUhmr9
vFYyFIZH0YZJ3crYHOi+t5SlCHrEggUHRapFoEbaFMJ9uEblC630ZxITck8GTHf7
pXSpqYHrWpa0cQakfLxYAS+wRy9y/gk1YNkzGNq1GZtsGGzP1t8+F1Qxe+4NnJ0V
e3InGIdbvtrxM9OnRpoIi749I0dp527mw6dNGa0+UPrq0v+1MNo7weB3xBdL6bhr
VUbk+ubbrAnLnxyFVZ++LECa2Rn+B/DSFJeX8qJKmbRoszwudOaLozsirdmHZCK8
QdwxUcqzBuHByqGN4gKaBQiAdM0u6xbyapNZWnEaKhcmkH1Au0qQVDhR3CKKUlnL
AzRTfnu47lc2yfnkFLoPD7uo2vlKIBTn9/kj4bT/SiE08J1jXMwj3vbXdCku/iK6
XkfYMsL0DGKckA4Rb6AvXXQFBlaZy7QmOsKDnqy0Qab1px0IhcadPJ5FN5xa/Hon
3ktuVKeE4WKGiQJuAOKzApRmjoLUQnA79jKrfO74qNQrtcN8YREdPmpgIzONv39L
up+GBoMDn8FJ5Ifrn1zHXPSepQIGVYkf9O2FxJdnYEww+NcddLkgweUjN2Z//o73
h1UMZMlIDqK/LVAnmWoLqW8QHmFPKeETJn9GyrEkSTZpnVlp3a+kCtzvXqwVKb81
8I64kbmWpsTHOdXViaQNmPwJdpFIWKCrLOUcOICNYDU=
`protect END_PROTECTED
