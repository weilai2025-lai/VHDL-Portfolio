`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vnfZTJY0TcKzLgE2ya/wLe+OZfCbIN0qdG8anvpnjBXscwpIGLBAxpBXIToOACXw
lHbDKy0XMy0VXmNjXxUTGkZTt561jTsy8StQefPqDX+ixdFBMnYSpZfOCOMFWTpU
8nzzDSfwbxSf4ztVAw9eIzHm2p0dRM54IUVGRCxiGlxbz1tUe18PrH+VtGX1Nezg
qhlr72wg2RImPR69KwyvAPNJ6+cXQ2yOCYy6HMRWon6arVk52xRJphahq4ZTQ9w1
KHsX8yNtkXmV4UJKYpy70+gpoiZVrUmG4PS5Xm2CVFEtJnYyf5v9PUhNlVWL3k9t
FZpqxVfOs9iFwHpMUpaoT1Yr2g/8Tgr93DlMKxVKqC70WdEjSLWQ9BGBOwPFVCZF
x4dRgtxy4oobOpqkEvNLqBE5yhSK8wU31w97QEs//3stER/8FyLoiAx4P1u11ttX
tISVqFYYnkzUui9obbtVmrmMC0N0aYk5GYfcDruEVbq7JQi9wXf+EquVRmrqTOii
brpNfuNWdRQQn5Yr/TglIeF9b0UNY/Isl7kbEXQ9QWbfB27C87AmwAjsiPXEm5mN
8DBK44b4uLNQZ+C6jV8dDnP8lLfSd+DEv6CgmPK+mpHDiM1r689nzp/3lu1jhG/8
M3+Ty1TgQ6Gbn+JDIldKsWbabYxi0lixNd8DwQwME/w7fIFRY8yoeLyN9O1/aLzT
aNBOCT4N3fow/xhQoxTFYOT5deGxADxd+St09jj74XSQrRYSEg2qaaL3hdI6ONlZ
fflknTK2W3Q/gEo7qTcb5mD7W4OMXRJ886y93VJa08ck8wExq52KsA92msl/X6Z0
Ff4jgf0wXeJGU4/fJEnltLrOSK6+rFMUgna0mM/JfSmPv2btbJcNl1REvrVI5D8O
bcqiV9JnWPopHOiUsH0Uctklv9TItAE39jGMPmWA19Pmeq5GELiRV+O3J+g1LaUj
Lipn/vRZDVwV+aBxJ23Vefexokp3k+0tUC4fGT1iSBAjkE2t3tSkxZjf4eIuo/qd
ndqzkwRQocwhF6s7ONeHfxG299IxKzyfy2dDaqGQSvEE+9mRv0zGnI+vILAosknC
9gheKEMaHj9swXLkj2e+nTCeKgfLLigMFXm2nkJ/ak4WAkxsX4rfxdbU6lZcA3OJ
JUl3fbHnI+9kQ9qBAFWQ/5m18bj9rGTJqVdAffvab3J0LsfhwUb2XSv0v7Uzx7Pd
AdNkWwiAK1s8xcQqdygcWJJ+CN06W2D2Xw/5X3io4Pe5KO8xg6tz2atArygca5cq
Oa8MKas4/TGXj2BMcNsfEj/ilPthrlOLZj0ARtDNH702JmpeVAuDQ6dCyZobsP1f
q+sT+XI8M4CSIc0qeCpqNSC+ixbhGWsHlDEBb2czGYVAu6FlufWtvTdGYzAhTfss
jnmfa4N04t8zpyqxm5QRUPrNRWjR3RiRNMq2YBJs4HOxgEHvb74+ynSwybadhPBv
qMnlaunTRRrxg+jBohp7C0yxeiGV6VxPXiT7fqynGzpRKoJNEyiGcTxW0hn+5HGl
D7a6u8P8uz6A2igrDy80fMfy3dwEzPShp3dmImiURgqgxAIH7+9A1tBjOXiu8j3e
kGGIGjTEzHRstFFKdMkWxLm5OR8Uh2KUARoHREV0bgh2Cv2juqhATtacFL7vQYIW
ryozJwt44CxpM3ajFo6SpfblpNsmhyittgkcAK8AMGuQGu06ofPhR56cSyWhEtNh
8R5jYwO+ZysfQnWeu24F5rBqdvPRIEep0z4ga+vPaPTJwMrJvKVrGpm8i6fCdLQ1
XEZPhKCHW1TThd5Z2lPJLK+QgkDJ2QdKr0b3C7XW1DAFNJv0g/Qi2WgCbTR8VUvT
s+YM3w72YX4uBaibN4n6ccl++PdcIWJZOAMgP/v7JVwdhHgPMbrIKXPfAKvv5+vF
WLbtnrNnoDX8EQcYEwXsUHTOZDn4zocvm+Fg8blPzY6QbOlnur68SJ8bo18QGAU7
TQqFmg1aH2RxlGMVDU/0Afj9YTr1YadF7/BH3xtoK8fOPvnyug3UWCUw5VEruAi9
aExLNdcda+gBeVGplVVSQhVwZ4FuhzHQQMjUHTWXPKlSpI4YGWh6SNaXFrHtkujW
CoY50pmyeR+oXS7TbV3nX4/uJQSobvfRMEb2NFl7I/QZnquszV3raXdrkJ5ToPUy
S3nQ1MnqpCfiKeTiJWUesB8yj5U009QJ6YFnsLKVqe+XDs+/LOQU+lEUpdx3+eyi
GKMMHchlj2IE1LiEnapQRs2ii3GbynPFCPrVVY9iDUv/SxA6ABLPMm7dVuR/Q8nc
wv9yGYQ+1eYSRRlsdCnVE19AwB63ded9g74erGKFJwl/Q7zkJrWksr4Bl2Dl5HDe
O4vE2ir6d9DnNzTYKXlN6lQ+ldtf/sqHJBu0/ZUWBPD+3yCnB9Av284ehfdau8pU
cs/S8m3uME2RzZbBqc2PeyKfAbAYx+ZFPS0cp6/qgPPdcVN1rbgrSfSKyijqnZoa
ktv2UozO+JieaJ3/t8kf4Utii4Un1YmkCH0fnJ7Ci0PieTgnBGIy5Rpe5I/O71dl
2gZPS1YeF9Q/xZVxO2GH6wbximWFlVSQ770xd6G0skJW+xr824DqL9AZzOTsNZi/
Osi+xxPhmgGVfe1vklveUV0NAusK7Us2pk1Q4uU63Tt+xw2fN3H5ibZdqAB4zR0m
95nDLc1dfE5rpFuhIP8/tP4ryskw7abrYXXJFns75ZbxEqvnBduhbPuTGcDeyEFD
f1219mGZtS9efsIDWcX2YH7rWIezf6T3v2RqOwFQBgDCypw6fpFpckVwlOdG2JZk
xEvpIP8VBraH+i9wMcGqk5Tm90107JhusAkb5mr0bqlTIoqBueU9tfjslRWO4QQi
519tKPgejLtPGqw04eKzqTkfrRiiis/HkCowMJvn0FQG2AaTcvG6O1jW/idfKuxr
FgRJrHV1zZ2bRvL/Xhn7yn9psfzmRrrfRphVx4mIr4fZRqVVLRqwpdhW3W8/98Kr
LZVOGeqx79CsG9dZW1/KXlhNkOYZr+PymTjaFYj99HtKbJmhGZrACTBwOwsQAqpM
PdUgDoOY7gHuh0Ec2vo31n8l0JkFGb5G5xckqreCMIsg9tcwKPBBqcV853+nbKZ+
3m+p4JszM5ySJYTJ1bUNZh6Wsct+HlcMm8JBuiz/2unUNt/ZF4VjzpBAQPlcCs5k
VfxjrT6TE1mNFZmZ8CuuN/mfRXtQlp6HQeBos+hizySJ3m5VcCv20FJdAnidpq+A
4MbTjZ4GZnjfsU7ulWe9v+M+FM6OQRvY8VmrjX7yGkOJ5t8ElyaCjW6yy3j6kPjM
tPzDsnTV4fi7dH1ziP0RUCqtVabGNV6kJBxvhpoHX+3RGnRp+4E5tofy43V39RLc
LaObIw2M4Nf3ePFUnSqfmKRSuAPmi3eKNtHPPVKLehMMApO4dTB9srf2WOTxv7LC
b+h87/5CySU0u5qExz+tFSJ0YYMZKXQpU4CnTP+vwpdZDr2H8ZlVSnAyV7pqPep7
9TD4QuRtNDjEfuuLh82xXayfZb76mhlfCBE6j0ZjnmXcBw5yVDJTd1jM2ICn8FW2
vR1OcJfcYjGHR4wV2gXtpinT4GAE6SwOEvD0e+v7/3WYZ+writ8nX0lbs9HSAVnh
SEDKPfERp5rI8I4vSOR60bbhya/BqER1cZqNQmsc8Y3z8jmAY26v+/oSGTCeB77W
76Pl9STjUayFoSIdYq/2bgypAOPAZXhgl3uCx1SQotoUuhW4TO7Hq6Km9IzraoDH
/i0edbj4B1lHw5ZMIHS7otlmSbV8qqt9wOgvMSZS2n7vUKvlY3teeryri+ZVF1se
ou+gLPQ2DEwTfP17Jv91c+Z7Lr+j58B9mVmNjZMNlUM=
`protect END_PROTECTED
