`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMQJt5U+rSFdHP1Nql8k7RoWxInmvmiRQEAH0dlgtUfaXbVg7rYw89bArtjVaYfj
LkpzKHJWfXMtPARwriaet6BhhvzfufHxOMjaxAwCcXyoIDMBZp+bcYbwHzYE5UeF
k+/4eX23wDpAo+jgg6MU2T9ob6zx7P+kiCyT/j5R0WrZST52lvGP5u7wUk3rXqTt
X8Yt2EFMvuHS/kd80yE5O3b99T1j85vXmnECLGrF0hnbpUnt3xAPFDuk8kjNg9uO
L+o2JO8FOwsFayNc9S8qCKdwXNl68VmPAVhZ0ReHkYT2rWTMyU9h2nBL/wzueKWc
Y5abWMSt3/TpmmwhzJq0GVf4Px4D8+96SzI8r4UokqhVaZa/w9tDYT3zpo0tEC/S
d2mcx0XBfUwgmuGvIBnN2u65Ow3K/l0ltAMD18zmNSQArFLwSWT7vFsudNQ9zouV
DGl6evI3XM+8j8JzTbA8SktASEqT4FM4ZP9CrcS7hXM=
`protect END_PROTECTED
