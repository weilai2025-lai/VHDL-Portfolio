`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNFGJts9v2md/ybpAXj2QRYdT0MYvp7I/HSRo/EcCoGXEnmw0S4SU+hfpnbyOha1
oa5uRMElCv7Y31iN9BOcxmQctqxcX2RiuekEWlHgJw+VB44SMPQdVmW1y+skLyJN
Vzfn/WO4l8+rA8kGqsOxChsj1FqN97AtE2aamOL28fjAeprDPERsJ3TiZ6f0IFZf
igPIx+4V+U1NGfnvaIV7j/3f/a5bsowYezDu4KJgzVDbPWeVc1/Sf8169o6d4jyZ
92M63WCZxWMyJyLnTtqlBf4YOypSKB8/1ZvvKdkyBZXFhU2buEhjlykJyZlS7KlI
cu/kfWp0XOgfkSyDSsi75B+U2o8oraqSWOkLSQ1iYEH0p+C9qi4XJburY4ppoWfA
/I3O4oSWkSF1pbuQ9aYGSQ0caM1H4o9Gk98kZ1pJzHVIeaeRXq4bRKFmAG2XwEAr
1EKFt1fit6ITUIrb/RmuL+4vi4e8gbbyV31SAZGtOHzNqeldComRAQYXDtdvaF49
jVztKB4I+IGRRbj4pSOoIMjOtmdvjcrZVZcCKcZlsTRFfpgkLw0NdG6DQMGXkcSv
xoY70yiaBvZRlW7RvXzqXNkJRr+4TTHscmI4wq54wtm7ElaDSZyvf2d3716BkPEm
4PGjPwtGJtbjkh1CWEwzeLnkT3w6gJ0Yw1Ck1SfrU4k84MWZ2+F7Pazxu/TQYrJh
QSIa7rZJWdLijFovAd/2Sl1gU1+9VCxL6LGPnvD71lQJNoLMmkUY8D/C4EXfHPI/
Xrhk4D0MvOr/e8nUBotjrOasaah4jY0b0d4KKuD/IWKUAfeC2JffNxt8zcfwsPVC
BE2sCEi/6cAfZ15ItCtNrcU1OQbi3kiC7mB4VaPndZ1NewO4297eCWyFUD8bhRbc
lX5fgioBywZsAt4G+J48173TgKn1hlKmRuLBg4Jj7KAEdrh7es33W2v9TXAY1Wpb
O+jsVEzCRForSogrWLucIYqxlSAmz7LbVV8ZnHnVv6JGhF1JyK9C1vduapCIU43m
ZqZ4kfO5e1f9WlDS8Z07A4QeLDB/q8mHiiY0IJIj8Vxuu61ac/89TtlwHq80cPgi
jub60PKLe86ejdEybXiWTmXagh72vVOCnnT7eR/x4EFBHx8lEOTrlkQXRrQhLd6M
`protect END_PROTECTED
