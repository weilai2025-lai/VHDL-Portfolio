`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YY4XblF9k2rJhCZjAGNViM8k1h1sdr1H8PvpgFYBaWq5Nh3/+ZIym4gQMUKinEb4
oU72Rb7N6gGc+VyY6T6RKvJZ/glhRDWflXqan+nXhHaosjDlXd41kSBgGdTFiEvv
EmKjEW4Y/xm8gXNBg1OA2tL7bbR7UsB6g5KOe1MVi1PVCA5CEYTSl9FrALZZnFrt
3zmOkAZneQP/S1BBTkeNlb4V3iY8tHV/Cy5kIRMnaZf2rsh3/0lnQm5u+xUp+BkY
W8SPnzwdafRgKznWsYDvYVaCPbafngZXHg7ZSQVVPhy2BGE4ks1+MDgExOiBEL9t
ax0N9HuPTnwwyyGfkfhlTtSN4E85xaOyRoI1KDbj+XE++igz0N0s0k43n9N5UcyT
KM6my7Qt4pooX8D7XcIW9rB9Mx9pL+a/f1X3K8a1ZkUfXwQDaY1/qCSZbks+9uiX
jsldyawHHirHLHlObx5ajSyJoKdN8euPdStnKWMAlZ9KcLbmNYR/jRuDmvNMp7Yo
`protect END_PROTECTED
