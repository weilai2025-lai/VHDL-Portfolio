`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WSvd8qMehKTFV5UdhjSUSNvU+TfQoJcGbofybzkupWo8NrhJIf6ECIdl28uL00Ez
blaDAjlCYWJxA59nOCG+j6lEi2NJ/EdrXyoIa8rd8ot1H4b1CImf4SQcyxxg+GVK
BEh4tr0iU3iFY3ixjn5WnsMHAWEigsWZZPoQlIiz+iEFbq5AEsiVFo0axq13o9Bt
HW84AssIU3c0bP/CYfN+jeMv+CZNRqGEu4JTSgMv/teRqc6JajqypesKIZ42Mgie
i5E+jQqMO9hBYeCo8fPXgDmYoQnnxray7iAMEl/3Lb+0/++nJ/rOQ0dqxpwKDcQD
bLt9loqmDItF5wDRjWncD4KvRnZtYpoy/uH0KfCjujxwdRypPXiRsMlnnMGYci6h
O8/y3QuNz+7HPDunWZpj8QaIHhOzac8A0P2dOFEdh1YuIP1TqV55K8CqZUFgDBrd
EsGRQ9cBi50mgDCKt4wx0y/tJTpoCTzAzIyg2FLTVCSWb1any3UCOoEA/dmPHq58
rOoNPMvh2w+gC612HbQxE2detwu5VD02BE+aRFMvFdg6WyP7CeJfeJ/O+HlidXZv
rdhyvVyHuO6xwCu78yWO+Z3jpCxrJdcIDXPLfIL3XMe0H5AN/a9R7zAaKrLDSiQr
NXkeHf34fyPDGaLiVw4OkIM1IMW+esGqnxYOiyCJWPqeEw0xcxv0pVr+AxdCEvTJ
loytZijUGBHM9h3jLoAMEyYD+NxeC+Jj4hOywg5JhgZ3/mHGFl/HK+Md/lw/Uukc
QydnSA6DwoDFkielrreFBEUwjJKg1H0AVO+xwCVX1kUP66f0n/HtxpQtzlEt7KV0
`protect END_PROTECTED
