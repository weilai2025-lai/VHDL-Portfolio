`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4hPihWGfSTbyKvJ58DYmkhGKBeJjNSqq8mXnnfBl+KHme7LuiCERuO+u5QBjhz4
29TbR5KnYguE3jZLS6yq2MxS7RvRy7CCynHJxFMS1I7ZU1VV6e8u1gzdhbwdhIGQ
kW4CM/5ypPY8qYJMfjv217wDTxyKok9Q8zVxNgX0PYBdTRN0SjA6t2Zpc3dBW57c
jfeperin1F8she60TFdIZSeyWohPj+MaAGXJFa+ffPTHVwSLBaI5FUnnnN6asrrJ
lRCjayIKNirb1MPJDwCVJICY63x+GHm/PowIGu2fr3sotZo4ByDvvyAz9f/EhPnw
aK9ZmlEqLAVU/ga0HA/3O6bum7RX4VP2NvTxA6Jfd4iu0aDYWhZ21qyoNJrIEyc9
dH2rF2Q9TBAyMFDDSh512CVInYXIxeWXpvZHxVGCVjnQzrxnfJ5Hq4LOBNjpt2Ob
OvHLMwJ0UAmdlvy5cllFXY1xuJgbivbaZZZLr7vDR2iCX05VS6ij3gzcoVp5HTPK
GZtRpP3y4bBgaKrDQ5DIPFiTZ5TUaSuq4ut/A7d5x0EUFYXoi4BHH6eBxmQy5maK
gvsNwBEh/EcxAIxkSr/W5S67q0S/rOQ6rUD69c0FEMlikLUubFBxPlS3DSNlhdio
q7lQx8iCq3OrVLytiNDBTmRoCFyG5ZG/7XPYqKovqVuTbechf2Gs/UpLsVrn4bON
JoFot5qXa3LnAQCDNy4kWsCuVeMl1reswRHBvdFa7vXrESKPJIgbvNgq2yw6xlE2
ckMYYhCTAqIKlfp4e6B8qpsQN1049/FB95bm9w7lyasu9jyOMXOvGz1bOfyGSPCz
dhkjYB2TyGXaemt0KUOwmC1PiYKT883e188eex3BqRRAhMVSAyCA6rdxS55ZGRTK
8VIYL7eXaxYMdHHv1M5MtBC5R3wjtFkIpbxGm1c5UfaRkD0+pUqlW4ICLH8LGUeE
A/tJ9MfIYDma0lFCPDdHb1arbjce6YtJNnhHFzJJAm/OOE3W0Mv7xvLfh1/VRL/+
Dry4dG8JQAkmpbrgWSiDuQtmbJcZ1gd9eXlncVqLuMPUW2XRru08rLYc4akHPWEq
GeU5weFJmSiw/l9RGxfHYUTU5xbUWjGVHgJCm+q+WouyS4mLJNdHqW3rmXS49O/a
Ub3SC8QY+0Gk23ozJ4aVPrGI03CtMdqWJjm5D27G/YtqsVJSSREbku16/UXxMCu2
+zlVAifVm+LSvhdUBgoU14L8wsXRCSWMNcTXiMudkF4qddtyrZfNvxTHZpsu7n+7
rhmmZscEOY23/MmOjalpenWn76DBog5qsdD2pxeQLP6wsIk0xYYT3Y+irIuy4c3g
G1BA4gvOwB5zNdyAljjJeT6n2XZ0jLHNbMaLhBDCPGmtWubkTuIv7DqCI4rE2VJi
u8IpfRZyErDO7weDMr9VoI3MkQMkskBFjah9k2VMeg964pFLN7bvZ1wmA4FxKVDm
oxi06giGvtnPDiJoc9aGMka69bFPEskRDE8LL15G/CvZjN1M2qoaSx00LYDG40bq
tPMhYwFJqTvIsZMb8OYiO907ZB5EnHNtMy/ea/0n3cnULs0ZAjFXF13m049aonMu
PdThAzAvh7YiGHPL2WQFERtL1/dkNvM11E3LwTviHwSWPCeK2ndswz3euGUB2kLS
NRJX8pfA5/gCCAN48H9GJ0t29Qx3npACguIiAPShGVU=
`protect END_PROTECTED
