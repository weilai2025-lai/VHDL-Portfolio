`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lq32T+fTiG0jZ3uNJTfiBgLhi4/zggqILm9xsRvxUgKBIAUayElLnW6usyjS/vOL
WvRlrvRLc79bZ574rTRKkuhmh8Nkgep/CEdC7JyuDNkUXsWzTR0K2l4I4tNlf3y3
iENZzghQ86mvynJN/955E4HNpwUQafLWKZS1/F6q3cWzQx4N+wcgcQBskONCHvCF
Ij2bfzRfjyg965LVjdsRZ8eA2LUALk38UZ/LMyFThx4aLcLXw0pbYkoN7egtHuyL
3yhHMVz46XsEYNucu+LwtffJA5GmKN0sTEnUT2DH6IgOucKySjkc/gd7SS5pmaQb
FHDbgAwiHoTTri/lBM0nCw6O2NpU4jwt5QkIt7AALOeN2HAJYFprr9KQsashjh/L
4pEceWqfGafzR5zydzlkol4+BNnTx6fuQIkWOGNCaHir2/3BBLE82MNw9nKEd+4g
NpU+QN7XqZ9ZEcQqBZb6RrtfKxZ1mNnWeESe0BLwXlZkkMmp+EMimb5XYPmMq2vR
kgS8DUeOdevXE45LEuY/IKmuYnespNCYV8On24DjeD6MWXrI58vDX4B8S+NLShId
76sfAVwp2e6URgXO22dvbfo/oNb/NAA8NB/9IzrMZ0qhU/OVuDpfOy4Kj0aE+j0H
5Cm6FKfSwfU1H5mIb1PBGO2BT3lTxjASp04CPYr8ce6gKu/QwSPiG3Bg+WEX2R1q
hztouSgeoY9mKVjdLp6+2eBvdjp/NY/Y79eBtCT8Qmj4hx1AGYW54/dAGN65U/8L
UcZFTwqJoyrtxxQCvnSKOYIfz2OQJlflXdEOwKhOZHSIzMwm59FzKhgse1AzyrXY
r/hC7xr/RjtPCBrhupDqPGYBS6IybOkVB/YTau2303bGaOn1mt5VNNq+4t3c0IWk
QgsVBgiWkjVBfb3A/qh6iAx0i39qEintkdsiC+hwQHxmrBMBGxCVVqCgXEWoBgGy
0mytOCQoqHSqLhMwhvcrSbUDmXOvNMor9UG8rU4UyhFt6UQf8hPSZ3XU/2zb017M
T+s1CoAygnWHaXTYCUCK0Y1hQC+dz8TtTweHz9NXpL1JoJ7MlsKmMFm8WyXps3NI
JuXyRw9SV3wrP9uhFRdWR/SUkxlKXG+OVOLCQKJvmvefWJk1RrpVUWoJF2TvtxGf
FMg1cNB8A7Er56yeSNewGHOU5rApgVmEPEcqLNC1aZyMc1k/NjebZFD/p48KpTeT
Nmgw0BGzFAyoRk2ZW5ggDd5B7QicMY+mT17pQPNYf6g=
`protect END_PROTECTED
