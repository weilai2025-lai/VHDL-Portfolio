`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzkDZZswxv1db+UxVoyOteo5JyQ0U6nt3q1NvE7wT2/WwUKqTI0QsUfqmHmZ+R0s
GtcJFqSVx7euNEHJIFlzfwFBiaJjUxOGdJYA15IXEi4/5p4Ks/aQFT0ZdXT8CIyv
5RU3+6VN4hXNF3BCiHKNhOfQZTUlz4TY0DDutWNrdeqqhNEWuB174fLt80mNw0nK
faVX+IHodN0HMfIuTd3o3effp5Wq5rGG5PvVFXqqYzFVZx+wuoi6xR3EAzpmi5Hf
bEtt85eJ9cobkW4UIz/ETg2l7Rva3yxqsnc3VbrLOQLD4PTfUxzgPQ5hbtZ+b7Ky
LAXo2/eO1vesUJ3jTtSfHTq5jIum4WLEHFoUJzAQrTsC/M/WwVb9lAMgiqXJap7K
B767u89bLqa4UNLWVcD2qYcvEBL82iTLJY0gBe869mkzycpa2JxHAARj5pNP17OQ
sX3+doSMkmV+OrkHLO3dy3CNvnrDesJgF8dqmTkg7PPpzTjoOoZiGs7+4eBYJZDe
WZUcvTYyoL6930BovLUyY2WKZ/V7t6yVESbT+UIQIeBCWy5jifDsK6txUOQQpR7i
pSzVWOSesX0y56lr/RYoa6hbl6UUMBQR/xqSPBQ9Lz/HiocmyR7nbwi7fdIjUOCl
miuY3edTNnZtvzkfEhVe0ix7R1wLUo7uUPHk6GiKhpb5XQo9D5sJcTIMiWyORl4t
2hMh5BsWoJ3ONgWlNa7CEeX/JK/eEKo7x3nrwnKo0Z7vPWz9WFkDy7ICGR0d77OE
ZG/BDhHW4Jux2DSSwcB388YgMT0nEIPkhVjKUrVW5D3E4D40pZkjQUGnvBsfMlqE
yE0/ggVZbn9PixH5sU6dhEtspMNDsq8706647Dl0hixLt9d8PGYwFZByq15vAvdO
Zr3qOWMmZTJLXinVUHJrPdAiSG0bY2nMewI/wvCFiWEfAAjq+C6Z7XEXOfURUI+h
uR1b0uI7/36HbFOqMnU2wpnoK0Z9fJYS3f6fIt9/JQ8hq04ddrOLAk+FO6m56XJB
/+mM5eqzrJa2JISJRIHfIsWpD05L53U1Rqqu68CmYWgH8M+MsHxSw5oMool0/MWz
9opnd9Tquxg9zXge3gIshEI09Wz7hdU1c8YBrC90wsGQ2+UQ+6vH6brcytrvdHtH
oJivrSzlDEEQvGDOF4BL20ajOWgCdVXf8PG/3Q4WDHKPX+U//zOUCSNZxGocMtb3
fcFF8kkxGuNkKU5y9vHMHagqNOBRaRh/yZMpFQIa398UFXssXt5k7KqvcRCffMiV
pM3kKAOriuoepFRIJZYx1AgNNxJA/g6Vl8f6VjVUJJy9gNvp6dktRjQH9HpSQp3A
yJiQeg5vk5v5zcwLMuGcob2Z/sMDVYd7T6iQ1/O/0rqdpNj9KOXr3PpPOCgmsdmG
vghA/8J7HcinmdmPLqShp1FuyHRJN9GA6Wn91o5G3yhk1tVR+epHG1giMoAlax8D
`protect END_PROTECTED
