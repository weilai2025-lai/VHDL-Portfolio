`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3yLJ7PD/9mjZbQa5AV4grE3l2YVdAiDi+E6AMg26OzQVlbQ5xWt+eYqUfK+bs9WU
Whbv4zBQnMY7Z8LdvBm7bTfnTOG6wLUdiYzHPUP4z04ZXTlg7bwyUBQlJvB0OW0B
KxP8bta/82ZUxs0hz547/AfAOcWZaWioNNefQXLSKjwsxBWFf11hgKr8la9mDtLK
qGV/VYB8DGCrvnMN2ov+wrDFxgbV77kH82/2TptfUHCUpdhBlEl6R7OC/d0m2/D6
nroIVfO0njhp2OQIOhHKs126V211619zwztfOXRoP+TEO7Y3jCWxpKZfg9CGbQec
UNnq0sYfu+cZPfXmGn8n5TeckfMVe2MchXihPjDUGxhTEGoSgfj+fqmQwp0RRYtp
SSYdVudu0zAEPnnCw4iJfDkInCqH6aW7baCLo0CRq57VIxiczXAlFhBdIWfeVOlI
xdktxEpSh79n9/5dQ5qubIMeLpllFBDlc1tL3BH9lbMYQz6LOWcCGMt4+n5mxsR4
+jJT3LPe7/fXdqR2tlgs+UuJ9dszOQ6c8cb0MOvUj3Q+C8W10LkIv4VsbL9hd7hB
TPx1aW73z9J+de6NMgfUPP+2wTcayN2u7yMVQeVtcdUpuADPSiIAFncUIuIWC4Ff
Kj+oSJ3zqMb1NCxjRc9jSnoybLB21YAhy+yA1fzBwylcDlwA4sz0LGfjSWBcdv2k
QR3TiytGzk+28Vfd3dx/d4g2djsdlk1eqbByVs1auIHY9e92ho0HWZ2cXTgadc2O
9ab9plYqIQT8F7kby8agBQozo0hlQl6T4dZunE7W4FkVibmpNDBX/U6JuzBc/85l
2TIMySlnb6r0gpST9lj84Zl9MrAl4Fox2azLRPzPtigkkNbPSsP9JmwVChDAgl7i
jsE2NBLeefRvlMVtR8vMqd6xns8BW3kNm7gAGaoFT3qjaFnnjg4WYTNLVW8XIFNB
ZVdh8AGIFr3Zgn9ykshscd+DSXwH/sJNv3Oj9QKp/3IK2cEjWH7sVADZZx9QzFiD
8ZCktHGY0aKfCrsRIeFCD1KlfgoVQb965d/hHyO6OPRH426O27WwMs8eUQHeiXNJ
AUMpwJrPRfgKqOaXFzhERoGsQdNF0M8T21kYHckTdAWMSgS7A3ZdcRvMx+x8MCkJ
pPohrahiBdrHCt/aqpt1rMyEbWujmTpoM3dDSrj2DfENnC+8c7BXpSXPeqtGFKrj
IyaeVcD671aAnhqAX7uKaPpV395ae73jD9x9+vSlDs/ntYf0+O6IBMw0SG0bKFEU
ahVcSPcW01WbtG3v3FUH3HDKyRJUwclRGiT0qwDrxcqSatZ+4L7oxniw3pftELNc
q4NQ1lpmRpLKIqqYNZQO4FcktvsRR6NjATn7wycVKClETppi2WMQhxX8tNtLUm8D
/leUTknrpJnCegmptNfUPYeBnyFUuQel9rK0tn13k/+sPciuXt7Vemy9AGczG3L9
gCsmxy6QpKdREXxYdaqvRpAZqbAjByyJFacGQEurko/4Niyi9I7UkutFbXSL2DZy
vn6bgjvZ6z3sBrxLx5RuuM5kUWA7TN8zKRwuCIMTZJq0o2NizR09b9xOd2GwueJE
i248n4jv8S2H+dh3JyWNbBnmoC0Ovu3HYkZ1tXtGwQc6G4mPVhUrcJs3P3Pwj6S+
O/WBWKdBv0TpftyCxpmb2f4YLSCLJDlzrT8lQucsSfRCm+RQmEk7JePHHj/3R1c5
NvYF/a2wkxf0CYnOI/Kz0kzYybxiJNRGVUIsYxyoo7APB58i9HOy+XVVHTIFkjGY
Or9go5pSVJb0uzS4EPWip6tkVNa7Q0XAZIb/nfqlLeSsFwYbTlX9G7m37/aE4oew
+YvQYjkcqDT7+rd//CK4uj8Ve9TrPE394N4tch8gD4t7EFQ2KOLgD0Y5JyjwTNaE
RKTXfgZvtdvo/pbk+15ljtXE2f7WVNeLJYlAzmZw+I6ivCJNmj/8xKkW9ZSgMLbM
4fowyIGfYrvYrr56WUYRa01WlVURgcvIlGrjU8e2yKiFqwZjZPyYUs4wsx+lxtHG
uDtT9x0X9/40vigP9XaJ2D+vTFA6g95lZTMIhl7vPmWgsRjoPtlR7xqobj1aQHl4
o73k6k163aBndpcusB7Xa1zOwhN6IYY6k7I0S0PnYUz96n/xaLzp7OnykFs9pB/w
Bji4DIk/3LGKxz6/iyJ+JYYcN/oDa+poas04f0cC3qfUOpyFMJVjbyBf49ndvnBw
05moU2qQZa5W+pfc4d3en/oofT/vqRe1CnYxKlOCumog2UthjW+7rc77AznMCm6A
bm0nk6TCkFZT3UeC8mqS77RH5HVq/sZP9C1zpYw6b7Mc2PPsSnAHLg4ThAEPMWET
POfMM3EPCYPu0BxptE8GMRjs/39rKckisqDPDeT+VCWLXkFDvjnm4ZBPtdm+xxow
NYTY0YXiXjvfsibyCdY62OgxlpbDMbhiU6z0BQWfzpIY8YaO9ZzbLx+0KXp3H3B8
K2awVvnygCjS2G8IWRf1anhwekbQRKN+32vzu+O4dffXsVVDlfVoPhsQhuxgfmtn
pu2oR+BxP0JrQSWxt9GZoeTXya801vI/VUpqkJfylPbsSPoKywrtdvJrl84F98Op
+Fe6TskBXNmE/POE7s74pyzbLmfjMoa1xLi3Ffp13bpedz9Gy7Zv+qlpemC/arCf
eEE0bmLh+uETm+B5iQ7eumfErgTV/cMPy0dmHHvuqk0DSnHfQamRlgesTndl8sga
H+oB4vC2Tjr12lbJQnt/SUY8jJvVGR4W0iUJ45cCOcpjBJNhSNSHDt2MKiqivmBF
y5rV3SDjI6ZGUeBADZOgeP1nnhKaoRltjLBVFF1i7ZNZgf2BSfBsqGodlXdrkcfD
lagtQmxO2kaHStVScZgpKF46tbjBpxjzjgS5WnKjg9pYgFbtsvNhnF1VZ4LPpKFW
7Xw6Ts82m/V+psqK/ElInaQ9WwA1fFjDD2iuCqQ06g/EnwUfNrGKY7FXz0UJRdMF
+8mNssAQSMqiChTGDUCJ+WmnY7cCyvz8GFvu+7GKVFg5wxF3fNIhf3gIDjuVGnYs
k81lMIdkIpxyj9u/Fls9p0rHRwy6Tw+3kC6izD3IFGPvcWxsl8mXTXL20c/3cqNz
HHQdTouK9Nw61LE7KU0pWnbMjlOf2BH3NcYq9dmozvj9DPg0TcuoNzULSP7EqJMH
KZ9kd5IHdPEB8tfJ60yXfPcL3buM7/qaK4lOdVecp+NeUKCAGAg3wZU87CXvNVjI
+opIrzun+e0MD9Oni91yFb4T/T8D7Fs0nJRL0abO+NHX0Yc5AEu9yl3C+V7vxaQF
9zcC2A0PlcL/5Zvkwws5NM5VmoaVNzD4G82mAnTqNQny2g84DyPPoL0C3fVLNB2L
0F1yhM4MfBNKDjUhn2dAEowi/GXBF0UWvwHCeEv03CiCgbtpw4R1g6UztEv5jHV8
qqV5B4p9Hu7gC07QfgMM0bsmmpnUoiu1qZlNNKv7JlY1b4Uf65zx39I7Sw1viMrG
V5X0id1ldHb2v5zok7Eif90EvYdA/rk0eEUQiw+JkNEkd+r+Io6mZIHbLw2Nzz11
thF0dZzUp8cBGs9KE8j01J7gf47RnAt6zeyO8k6eSDgnufq5UgiWRyE2m8Prgk/T
2Ueb6HqBUVpegnOCU5kHB895MpMpyvuj/3RR88i1f/bMDAYKgVM4sODhYwkpPsBG
rn2MjA7NkqNp+i2/zkvCzwVBBfhpVJ3BTrKkuynS3efaPHeEmSqnXkl/YaUZxLoZ
kRfykAaOpTlpkYMjF6YonUt2tCX5eJJYpIQ868cdXW0DdOkxvQq5FMSEjDvApJtE
u6GGacTAdPN9YXe3Tn9QiWecdnumJ5OCYyZpn+aONnqy77z+o14GIJ7EE6Ox68io
Gun2UsGYtTqOWVoPU8GxjYOBOrBYJd3BjNaKSMrtoBg83wd6G8Pd7CuZJKd5GAYr
Y726U8/NO6UTEeheuahFqkHpsXZnv8R/6VPHt9wDhdCxu6Cs0QkFAfrG6Nyl6lHr
XmeQRHSjskEQjlTvTKG1aPAy6Hnf2EpIV0GZ+bOvYqk1bXtM3DQSRmk5vYotbDpb
l1Puezj/PKbwMUKSP2EmsOh1n83nrKLpebJSyH2EV9wAnkQ/sJMCKP0FbEHOdndb
wvPMohQdlD/h0zy08BxkWeQ7A6eiz2QU22tHofVbU0lD9oKGMEYj/y4m35IJe2dN
txfQnLxv5MjThvSlFcouesQVUBRQVtP+RD5YPi/PCJvSeH9Xqu1sCJiXkZywbY9a
9et/RLFqt4RWxvJZ9JK9iItZ3vXxGzBKFnttvQXk8aUiPQLG6j+0UwsRwa5+X5TM
3GHpvpGMDEkTnML7IWYC7ts9mZsZgwsoAkdzjAbxR1W9OPT423omdcoRBfhxMBOA
mSsXMvGwBPCqAVG+Jor/8EJOBEnPXYxoiBuswG/nDKYLalXwWQQ2OhHuim3Gd5FR
+7bHDBQiwq8Bu1SVxRxxGQxPj+LTpetIHkpcuBXSiTkLRThAL7OEHXFwz1w3xQSx
C8Ta+qif4PJSriG9v5/qJ5xIsYuqDE7XgSaC6mruSOarVGCDc456OSbNLOzvDoXM
h5hoSrByPYicz8LktwBQ9L0nE9YMUf3ITkKQiEMk9Z1/AWs7KWJY69p3nq9rzw1W
Gu3J7We5zfWTDgvV0vSAjZanKTNIOFhpyf/ghblJWmFXqviZKIO2BxszO2o2c+s0
fM2A8ekvXU+Y9p8Mvd3WIymClMXsB+5+uV+/tWc8nGuSNvDtWXkNuq4e45495JIB
XU9cMmGidynHhTz9qhEcGUYi8bwpCRCgkIidahP2gL2T3IZx2mCo+mqdVNw4cmkI
7YjBlyVEkhhqhYKSdwFD0Ziy72itHKVwf2QZiQpmB1xxjvHiUvEzFWsoq+V3Q14J
cv5Osy9w7/vDz8IWi1DQgiUAbdGb/Wn97KPG5f8RqOC9raprEzCH7ZIdwSXJRxnK
3pITHypSRhtToiyw4VYWhu3KVG0732nUXIyLFQ0eEW6IJdKnW6ZdsWsxqQIjPd3D
W2tk6MOZBxPo+Bd4KsNTwWNVt4+aixO5HWZKY4BbAOo0pUwIm4vx6dt/flcAye1A
c/LsiVaZ7WDM4kfq6GBxQfDvesmbj3L+a42hjqBpnYeiHh/lelg7iddA47xu1YRY
1mtVleGp7aUhiywcWlyOc3DgoAv0pjrdkTdhchlEn7dtK7MDV7eGYF2W9LPOqEio
/QbG0Oct6v7EIdPKpB9CBBxgNbibADrSYpm4bbr7K1AoP0odO6xaFRJtFz1RPPeT
NYBiXtcBnVqiWuPq54Y+F/xIuQ/0/13SisaUAbHNeYchKEcu23H4pxFiUBHWeaaj
dosGWdLLBdZD1qPBv/nuCIjtHXPvhhCcFwdLS+lTHIHnW84Sb3CfZHDxk02CnfJ0
wiILHXSHsxlU6+It+gVoHgomOykrfbYhowkzywZD4uL67hKk1dUmTeF0YFX7fXO3
9J9A0wFu2CQ9d0IFryBOq6Y1NUU/FO1W69H4VqNXiolhj2t4iCZhcj0uzqW5LW3g
YcPOPXPKv6wN7OBh+tQo5pLZo4kFqf3UGNOjM7dAr2ya2FHVQ9odLJdulPrcVBMq
E/vnZ9E4iQP3K1o5HaHN6EMG0jA8SkPHqYhMtNxxcQFWuXNAmqaLUPF4b5RXJdhM
o1UkbKir+EO8FQAw9S6kOfXlTB6/0Avv5nX5Xh8/SAOSMANbQrBx80MxdWvL0yn2
v6O5gXYhGWABzFtogELlRRWMO1jBi47oJFpNCNU5jF+U7hncaLBHcWVrXBXyiqcT
fyJRqrMo+pgS6JQESheUzVuptcmC+01UTvt1G9AcrXvmELmILSzO09ey+VKBwuGm
Lfnt/8lou8ABrdWgNst99aX/If1jfsrMqXpAl9A6MYmFt7P4k/eFIwk00JxmQmK2
puAJwHpouC2voXBoHccXhNJMVuHETC2YX55AsblzaFMRzJqWYelyDBwx7ciLX8KP
6eOjbr9UvPOysyTV7yuAAs8QiHCds1QjWPF1Jf724gsaCZPNZC5gMpzAuF/qkLT+
NsD0r12h+Gj8hAY9d/sujjaG9muiu0FzC8ORvfB3BNokt3/73CotY8BawEE5bVB5
OZUXcyo4vmK/NfupZ7ViwUm7f0iKCQLSV7GCiV1HPb/dd1/5NwTwfxRcUIVKLoqt
AZG44iOEmcQy/oI5UjY22slXbvSHFcrRbl4GgUy1xDATF7+WbiIUnj0xvgPVxedC
qUY8f+sn1FPNEnjwZtHgbHOSre+CgsGi3sIDKeys5tIe90zEn5hRMmdgyF0nvYa9
5ZprkAy6ucwmttNl5btyVliK/Iv8WKXwa10CwanvSg1yuiI8ko+j9gWbXTH+qA0j
8rmPp8adVPVln95wQHnmiwBM31SdrGfU0/1p8iC6MYZzEXUbUfQS1pwhoNaZZqIz
H1KUuqCz8WZnqBr6yaa00QlWrWyEGfztn47mn/ql+P8xObcZl+CyAQrQvwKltbgm
PJghYZ81yaFKAUk6YyQ65CeMsTl1kQVXD3+T1e0VMIZ+aIZQneW9kWXbVFMdLgWp
jqZNZNp4SjHJjHPDbQ11tEG+Joy2fd9Asv83ywq9PiMuLx/5I8oJUts8hrZadOd8
RLAt5yoTgCzGAve+OFsfzCswVsSz7EBmwk+Z9BPsrahR4UI54NO5K7IWvCKWMVUp
BZcrkZ6nyvyzwrNA7yYSHC6zHgfTH+DDjyc1IJ9hzUbxQ9LkH1umFbQRLVgg79gW
HZolIcaP2nyPjQ7l2fThA71tj7yLzWMgLpvqxTgXyeyeflmmKgMmcVoiS1sQQaPs
qUJ5Bppf3q0Yb6yuYkMokvVew5xCXnvv1pWUb2+7q5Tiz/GiVo4wCxMKurj3AIB9
9bdABoDkqj/O138XWAG0GfFL+oS6ZDnomnRJ0NPNPL3ISQLcO4rjJtwffYJF73FZ
63qSLh12OGhs+ivi5mKMGoPEgFXXfGFpphOry6ci2SiVWMSZs2fklhFBXhAhIktW
v/Gfcpx4VS44xI1Jb2EtEn99dBes3ptt+hBMjCn7Um/bx20z/2AFbnlQvYlY4otj
oyRmnf9rk/4NNw8k0DXLkDoHDWgrMiPQLkoA6arVLXvXM3Diu4+EYEdcpGthZ4RG
0dszupRjIj+iF7OSsWeyrj97qnfGWHiiL58zvIslZ24ft8bdxCR0RFJn7b7XHvDd
SqpLl9PrIQClOYad8qQToDLgiTxM++LQIRxeW7FX2LYkcHll1Ub2QbzQgDFGI1ys
bIeP6UUBIhdrX3H4bqBgMY8QYKGsKxJCKTDYOg/QJ4tRg/JTiB2tMO4mLd+Fjj1T
wY3rjsqIVNe0L6yxhuJs6OZ3V6YPbkgZ8DfQuhIWjE+42lW3Ar2tAeB4Q5+uUJXr
KEZi7fEEVGkQwHnOiJPtvKrCN36ssNrqsJcj0i4egJROh8O4CEfJewS7+s1tphAX
zoqlu+bBGwzQ9fEKzEIRl+tBbLmxFoJXOsjjb2hFNMjrfyislUbJtxHjHwWqn2Vu
tOmNaTA6fPt3RZ/nXJouVTyowd8ysfi1tsljVt0x1hI47HV17L9wJel9GpuABVDx
95FlN6drAwAE/oKjoi48WJSZtOfHgHUWx9u2mRRxPsfmYYsO/qdRsf3bF4zwG5o1
FMpW9Pw8U0IH3GKrJa1a+PBEvUbVcfKRp16/CApvguw1fuAjjpvIIGGFMXxja4Nt
9BfOHcnEbdfwuQBJFvEkHhW0ydIgdQvrmDt9SQdOMYizRjLP0MW6CyWliQcUUF6e
8orfeFneot2MFb5GdE7q9EtTpxbtHTULxFueswyZM4pA1n783mpoz2lpPu9DxxvJ
cJeYVkDzX7xXr6DYAYA/VaGuBxClJRZOc7WL9MlMU8YZNNsjo3NqZ39rYX431BWw
vvBaWe2jdSAf6a5XB2fo7xKVZErUu4FsxnRUdr7R51eETBelEpj/vCD9jNh6/amq
ZNK0hm97QUTaFJI46JD61/g0W0r17BQuwb5YSVmJqcTCA0gUXkD9Pa+t7vr0jsky
gnzdzl3o9PQ5IKqPzMGEXGzBnDlwuVBrjeCJsDzy661VaxcLkXRJisG6dGEL9Pd1
Tlui38NVMBNf45xP3zM4AQQ8JGzVcS4964wguqjAfh154hhYG8Dh42E+X+ZpY56a
uJttrPz4dxSrWRrLOK7BVySkDfhVP8GBaZJrwqoRWZEZc3VKbChlVSB3H0CzzQUv
o8zJDC2hgd5//6hh83RQi/ScZK+H2Cr/6jXRS8C8W1v1+XynCiFKU4XZO8avwdPm
Unb5GD9CN++YqH8iw3hKZ5edOuitoZq/XU33r1N2gITEUjnHlMtmHIxmF6HEBmH9
opM8v1P2a52/8HTAyt+L9YOYkRo4i8Km3SJzJxwiL0WUAPRgqH2Hqk8fVI9/Umqa
9hGl25s5f34OxXUNcbDz4A06s++ql/OtixrLZxFJDFDE/G7b8xNhqHasrlqcpo9+
fgKqrxLfyuOcYIY/SHI0NO/UGaiKTwVBmZFkwsT/goivI0jmCsL9gTl0ix7GymD4
7ufXOppcZscMH2sAeuLiKqdI4qkvA4gq6NOd/Q/ZOu2s0scgFQ2mKNRSRsCfEs1T
1NTS8CRHn9PcaDHSiHbzVl4U4c5G1zeu9l1qpmrdhUAY/tDA8IJX4vbQEhm5YuJ4
gqWbDmZ2F4vWKG+fudA9nl84LgIqrkE7PXmo9bNTwZvBdH6DsJtFh6DTGE8kKTXK
TJkUiysDOv+2v4+DY0bElEsdxidDazzOgIDsyQ639TPW+CV8kPYD3nva0ddvVvLc
2Z94V0lLJoZOwMNBqnhYP9u6wZzJAIRa0kbn3yeMn9z2vX30BEBQhYEd4hRiHwnw
xyHQfwKmv33GaPl+1fsyykoGZFDNbqavM+3qmfkFVQVYXSzTMQuEDwd1B9ZRiooR
EHWEBO43b39C4oQlsiu1uPAR/GtTDQy8WB9qVpLDrlp9MEduCsu0vPJgtMyj34b+
07UVG/gHKTVmK+7jBxsp//ZBrk5hotfqh3e2eDmIq8CBP7vTJLglf1rdUwlQ9BCS
DX8TkimLmm7dxyoKyiZTK8NIva/Q7xhAJkrDIUF59d/L2+/DZ3ywT7jbNCoYESHg
qkI8bwGyJaQGN/jA7nXdQmwFKmjaxfcbm8m5kpNSXbUt3jECmChXt7HvZ7NKUeBY
za4bmHww8UEZ20LbCvGAlLZB4FtvPAm73xnlK+PVcgiiZV1Jvlcg8gRnEoyhoxZG
LsE+0zNafxRw7DkUbje+NNYiIIXXfXZTEho8/6BqjiJExzgRrAoLfJ1H3uNzF76n
Q43is5m9RIWve8t7uo8ZGChA3PLZCrV0kYyRqgl3f2Fqf0MCWAGZGfC7v3Gjcyj2
e4nIFOKA4w2liAMzr+VqiB4R6d6o6sG9mWHGpYbVMrdDJz3x2TYIb+rGYnjb+90L
YwHRJ1UTk2L7bKU0SkEeEZSujZ4RB7eRZ7Imb45nH4AktVB1M6TIadjUv0eHPelO
aDE2ZbHzaNqUXUHB3JWh/7ucmjwBlmeq/Qpd5HfOATN/3n/SQ39Z39FO4NA4fLmc
G1+vf+YPMb+vPIKVPuGDckd9UHfr/ge5ZfrMT/Fsjbn3G9kTOb0tU1dZyGwBKFB2
iKhmX0ymtVROZaryLPTsyQHWhsvckHHlKbwp3aTOVltgTgeRjFOXVSMIh3iQZytx
UcCvCa9IPgXPLuMXqJ4KwVqsRM6BTg11I8qvQng78zYFU0+jxR/VRATHP1UlUJdL
REEE4FM4fkulQ+cBSmcYNYJwULdZReLPhZkDHiuPsgZJQFsZG09P4vhkTRLTQqBG
4sVb/4Tt2bcJJWGiENbVkgIE2x9jZTAc2XehH45Fp8RwOIYjaG/JrxkP//y3oz8m
S6WGuuwtpZJNwkhXpuCuvzarciy2vSzBQdwo+qOy7f9MAfKk+DqdK3eQC8XQQlFu
CBJT3U5FcUZbMgyAllJRWmu4JX/AhPo7zpVR3k96oXU0YhlawtSs8+ZF8xq25Tbn
5/oCOVZdhMm4+b/uWcIXre4tAlWPalyKocbkpdgJ7JZlMTSSI+07fpLmYIq2qUx8
nEnIqoAi1SwKKchFPXjIWs9Zqkt7wrB7bMk0UvzcpCIPENzTD/V91wJu9d9b+oEr
4dhf+vUSkhmI/y6x0ywL2COBNfUvdswYwmV+GpbQ32eGw4BWThCjwdutXiSAKgAK
pIyVzww4HSoEJCODt8tZHvB4pLXD2qz8SnN7HOxB7yx4TvakM46T5qcx1udnPwe/
6SkhprGW88JmZFo2QA/dKWk3GajDOFiwUV9/CGABWmw5fArLjN/whA5SYoLhWONs
+skKLZ0+H26gIM4mQKneAc1EJwRBQXBTGjRjiCMjzRwBnoKG6NWY6fFWw27ApxJ7
lYw6sHazAIrKr15osYx1oGc3YoW9dekUVPx0KCBPfVKs4+ZlLHg5Tda8iyRK65hw
QEH4FWfqbybtzW4v7H2FMlkVnvVe4IrY94UX2jtMA74Q92332hqe/pin6QOVDnZ/
JC2j+lsKo4qO5KKTZHGnGl5ImdiKf36Yd7Sk/4UCrCQnV/gLn+PtAdiYva048E07
VzCjE5dyNQwKQmSAIxoxEdn5XRIQ4RVPDZ+xQZW63BOfRfzgVTJSUnYdGE2oDNyg
pGoGUItywMCejFxU9uieCo1VRNfB3roVC3FvFFy+WDcSQF3CQEK/6aUo1Y36P32L
5Xrx1JYWkVwZBUzu3RXl3UFbTAqUoHV4duEVPYD9p3E8dUBZDlshLe+P18BQSYFM
vt0C7fAA1Ii9Y/RsqeJROcsuSDmoLvafS7dtQDnhZSt2xjcFYsAuRumlk56IAgD1
InYdoCLnEXTBwOPnA5sWVo0u8MCwOFgHhOHqHT7xv3kgPKh14gWwSPql90iP762h
cQ3d166J1IMO2lerzXZq78ACDNGn3Umt2ec8+LKp/vfWu2qnHDHkcTXBjiFF0voF
LBNbLlixclvm84z8aLTSBhOYCvowQVOC9gxhfAiBRnNLf5PM2m12jxyjsPBfBs0r
0nBOl+vC17xcUqDBa7xbPytM/if5jivomY+2lwMeyPrcX44DElCS25CP0b/c4w1Y
JRgpsIACJ9fIJrbFtKsMJ9tx4O/p4QtqjADPWRimyrQvob//OiP+lF61Su2EG9os
cwiccOhp88QKjJ8jpPPRcqQaHomdu3LtifRw3DdcZDzqo3XypFbVsRgvE+1YrdpB
Q4qvmlTSeKMc7AXP4F0zOimq0R7IwtFoz8xintCEV07iJ0ktmp8EWkQ6GoPfB6JZ
mBBgePBCoTyU/gcJcgiwlIT+De7NPyfbL7Tij7VQaLToRI3narOM1DExnGFK4ySF
w0oDAhePQTQBLBbR1rEr+XwVM06ZH1A5gc3Y8RuWuPlE00//FiK4KS8IqrzjHl1N
gtarR9lCSCp3w98oKCubAzvSW7iN6zeS3aakKd9yHoYpYVE5eexws4qiy7+5kGzp
qDcg/s7u4YXZQiRkJG+ENgOSEpHq/jf29Vml/W/XhUqocr5pqrJ+vpixpShwNzTX
QSvU5hOGyta2N5xHqCKz767mD4VsODnThrCIbqGTBCunTiESt+cc8Nx0BD44qHml
2zT6bvDQzXjwt6XmzHPSzKkd/vFReIthxd0iJ8HVbz+/UCeEzULcHMeIhd2PZfdp
X3SDdHpFM7uADBpFcsAeYDQEkEnzL5V4ciN3zL6xPGv4hb6pXyumbm7YSuRT5jJ2
BbQtf/wh+M4Yw55xUlNqXC9tVsb8hkx5AF7j5PzSBZOJQaVgibK4wpPbNpaUOFGA
RLSDjFQ6k9lbYE05UucLNzJAHVrcDdEeSbDCjkp4htvvdaJkH2FboWUk2x37/+FJ
FVRNarRR8zvEavc+HvyaId/xIteDoWR2klJ5afaiCWf/smJUNijx376Z5UMkCpje
Lv63wzPCTEwBJ6t6infuugW6M+vc6kgb7SneFvNRk3SIZRMiDMvtGSkUbAUHaKI4
gxHPK/Sch4CYJsLdJBwDFvnSStBOYwlGeN50FWyy28DN2wmZ9KmZm7Qq4+Ltdrwy
yluyW2DS3I2flVIqma8M1tMygQnXtqnx27d8gahKxB/4iT4DwkL0/LeRBDlRttkT
w6PgXDA7bmWKEG1/txaysEu6MrViBEixttplj8bPxlQ5nP5xFmRHb6vZtIbCOfAb
WQjuyNs0WH+ta85l3m2o7wWI/c8XPyEULbSAm+LSGMEEW6kD7/+EixvCcVaDCyt4
DcLxIuHlBJyY6Iy2HjYUkzOJF7UMs4cviFitzDNafRDi35WJnM3Go3oS7h9CoPjn
yAtDS8zHfRVhyWoz00Ify6cBLGPxE9S6IAqNM/f/n2xta6TCWCQP692CVs29RPYa
gqXuDL2MyS2h4mdmEBXPZdD/XMUC3lNuuORTbDwH/h6GJRzlEnvakXpbyy8Mb9p8
MxG0vug5g+acU8Kx/ITnBzG/kRti1lFsUX8RqeTUWPnRKzc13Sv36EvZOlGv9MXy
F9hEq63uu3EBHI/de3KxKqUMYP2EDZlCmYbqVAUhNvfRkMfEyCX7iMxYLP9Bz0Zl
6BjfRCDk0M1aJ1jnjGZ5QoXiE0dhcrvd4wK54Nce3ffp5yRNzHrPLJYIi9hdW6R6
Wxa2w3QN3DJQATUDsjGxf3can/dqwfLjpn8e2Y7zEfwkEcbKaIDRWNQUGOBvWH0E
GnhKXlla8BIxFV30OXE4K9l/cx2xoG5pi3iiXTkjCOJGKG/SSBCn6sKfK21JcLNH
ptJGetSFibfpkRn420IM+qsZCEgaX3R87cE/b5lsGH0+dciDECB9mhec0jG3KcEs
Y0ZeAl7PuCW47qU5urXvFf210U2l84HuFWDGomTXomlt0Smz0silOx3CyWMsyzCL
O3LlCNvnMICjhgmExb8n3lHUJjtXIOeBWKvIWYGBxzyUrGYlHN+NBLk10CfKpRrk
4m/gv8usIyNgYq5Z3MHaPgBtyVLdjfMkTWKfbwadO+chRBmYZSLI41jpN68fHEN8
IwGt7jjPgkDm3hNKKBOqe+pwhTc0snpypNOXZguchg6aDRsm3CAcCX6U5EQ2kEXq
xmvZuhCW9EbMRacTKzbknb827TUAAgDMlBDjXnQNrmO/lhJsWuo7Qv2ZYYpVgw07
ssIN+XMDQRdhRQAYr65hh1tmyyX9MebpWzqYDPustwI=
`protect END_PROTECTED
