`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CwRiuNq3CWtqFr0hUm0W06jkRJT4X1WHQqy0NPVRAkBqDZ/98m8SoVaCOn9QEZh
hzJpKwmbhvWqbQsANuRCDojEbjRlbsXKdAhqNjw8AwfAYGbJO639ROXiMVUm3kWY
J+l6vXj0fIkvV2hvkQkp1UraHTIqxsxRr+ltQJP4z+KWlI+WlDkRmPoeyMEWFYhQ
Db0BgrOW8cx4W7/Nl+YJwrPDidJmWvkFZgqzl7tKz++s9C6dCidmBw525TKpZkzO
ojSq8bDk63GeB51USkHXAhpkXlyHtjsX99j5hHTGskhOKf59/3zeTG2JGKzvZjuB
WjPWjJTgnD+MxIsg8mk0mU8QgD7AAIJWJGmL4E1bb+XV4q1s1czjUARE8jA2VBv9
KgliTQLlAIOD/JcIOeJ9jnXlBcVh5XOsCf6ZWl2VxkhyxYPx5GvmEFcbdU9RHl2b
rHxCSAEEChOg2gv6BxkwpHTgrXJN66os6ts3oI18wCMh1PUkuZ7xMt72Xs9Snx2F
llbXCIzlEfjJXABSb9MsKs7pwQDteA5nYF+a7Zn8CnZR+NCstGMwClNKNDRpUwbW
s9b/3rGhzhpMnJEmTE2aid4MiclpGnGhcgNOj14phgeamlGsn/klesBXzWymGumu
Q5BcdIuL7zxDAoGSMLJWAYqghgbNcivs+DDvuFiA55/T0jjtmn2ZAjOJO8eXAime
88++7kDZLA9qP86/41J8M/rCaaAZbUshHsc0VZFzpvM+t1Z8Ns/M7h6GT8/Wcj1C
6OkN62MysjweC4bzBO19rXU5302lq5czv/vU/YWC+BEJElDKQY87Najf1bzGBIp/
MqiskzO60aBIfLDL1oGL3WWnji/LkPtEVAorJ+++A8nT/dWsIYstszGs6jDkxFSM
ZizGZGFJXbkKRn8uSeUhsD93WxQqlINa9u6DJoUHBeX8mqckdyLL/Mg5d+29jcOm
pVEf6GpGqLEN7F/L1KMXd/xEj9Lkdot7cR2a+t7yeYRuSFvw0YrQF7xO78OFUywv
JOeQtB7/dFSQzO0aOZxgpyDJuaFiAwVFhEcne42RXIKGXHi6kiZCoS7cWY70t0jS
rwzF2k5IiQutZhFfP3cynpS78x2dCY90ZmyMXO5+a9jy5uJHPQJvL4tSC2H93o6t
4ZVQuQHFf1Gx0f28ke88gzpe/lA04uVktLD2HXiBQ5YqDMX4q5fsHdjweVBqqo/w
BpdfO93Ae2qRG8QikSkC5q6MJ0tRcrcTOyl7EC/K/CKUBkL5r2/NGnVhftz2AzXv
q/8PrvMhzyI7wyPutBtI46kSMmY2p/vw2qS4f1Ja3CiUex7YnOybwsj+NG8K+R2m
rSjph8SGiQfZBfaBBEVFhgO73z6J0rsBBx7ibJJ4ISMeCYE2156LJHG7nHsgkW78
5rb36Fbcc4mUzcKvb66HtnjYEK3ZXOenWRFMiKLnWEJRy4/QHRvW4GFPZVhPxPUB
`protect END_PROTECTED
