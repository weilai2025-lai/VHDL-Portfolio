`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p07D4IML60Oe8VSTl7YPfMv9Xw3PgL1BttekRk5mblkRZZNV5+q9dyLvzLcafz5q
CY7QBav7K4t6D6P7UOucXuRJ1OvpPmb3BcoVS98OHKUsgpyh8xTXoSCPBxzTZbGA
wRq1oM6QNHcOcQjvgYOSTQiqdhmjd8AxncNSdg/oM7skybfVQyKCTLtY11aLLOJo
vg9F/t20Mg86hn2VocD8MXR9eu0riHznulGc70l1W9DfH7nyoZ3Bu5kFSrO2GnWt
PpUfWFzctIWXZj+goHtTiSuKLGR80AhZTiC1T2miiPQT7fkkUMTyNbhfzTAUIWh2
k9EQGDuz57hdvrCHDx1jBdGuZOI1rwjCIeP09xrKldCu3QYAPmeApeGsEQisXBQm
t3I07um/92Mik3NtGqQqAz/ZzGrCf5TcKbPkF7G32BReoG8kHrP0Tg/ZU93G1Gf3
fMhi38+N51A/Zp/lnKcQP49vfPJpYB5Kdh8pArdZjtGlUTkf3ZK7rMqewCSQnq/n
V0xmdHMsv3CpPkAlVeGsXZOU1zpBpWS2oJg7Ogi8QlATQ7bsMiU/jVDhwSo81lEb
Bpd5/2FNovTPrBB8j/5ngiC657v3zD/oi0gdQ5wimLwHkc5MBHHNlWzhEcTFHPGk
0OyK2L34tELTJClxZz84QtTd9wGeg+9MpFCeZNUh9pSwfbE4uqLygZrtjIhNmQ+R
LQU+aAH5sTYOqxVwh5W09W0r6gfBQ2Kf9UZCdUoRqxMBEcoMIc5LehrZqXm9UFtz
1uc8WxyoM+GsOnvkKAg74i1H2mb+MLGUyBQ6kN3jls70fFgZKMuJfbLVJ2m7Joaa
84qz/8jjc33jPT1RSSlOsoilpjQCe8mGENcnRRL4ZYSZ/a+grwCqKasL7kDO5esx
xkfY0X/pCaXV/aQ3dm+uBtpkDDYcaYTVxon7BqwasEUI3NToK9VPDF1hpqGrLOql
FVFK67NMaZ3z2wf/R9L3OlLoKKNY9n744ykIPN//X0maObOS78wjwx6ZeN6cYdSO
Nnaydw4mONDhZYyRf6RwFiwomcfxo+gs7HyZUXKWpx+6it06ZgFapM8M0wSaNhZq
eghP5qKGUcmXQOk7w20w1HA1tn1PUq4v9pTlw3qQ7CAfXzZ9rv9XCUc3TgpwJlQM
8i35ikM/qVGDDB1iK6dHlepryXTExUW678ViPMlJZqPLbJ1tLt/q4nTFmJePDuig
vJFJEAaYsdNM24eBu2US1QrMhysKUzbgthMM7W8eajR6EVNA3AKBRKgyqqm7bRhA
sYXD7ZVwpMdB8pkB1Udvo1tFTB8iyy3TidhBbuoEalNkid4UWb5Np4NeJBhjXb9n
+ez30OiHcwsWvM6Q/H904ruqMLhMOJDAsa/T4sxNoKwEK5rwqgkeSKinQdOu4dck
am6X4EiwuW+27sF30GTpPztbB+enn5INB42xupAihtlc+r1hn0ZacaVsJPmiggqm
EHo/6ZFNQvJ3MHyPPC8aF4Xag0gE24CqNmFrLZ08yvamJmC0dGcsdCa0PirmJ2AJ
fHkPbJ9wSSJDyhHPrbmGn49pq8xwTMDUXyFjsw5up3veiwXXvIsNRyd3dkQcxJjr
dbOzPj34H+pfVyJZ6CnacyiLgT3Azd5XpJ789I5XNoMjBAUJhXsT44C1OnTufVUG
GW7Dja2MNCU0nzwbWvyPs7/Z85EbEz3ZeGlHWh+5wgWxOjkmw+bwkWHhLkDQv9TO
OGol6FjXR35ENaJzKXbNHRy7DBGPR5H7bqOKhY8k591rxYVenJiVz1xqqHsMN6fx
QWqrm7sRJ7aTGhu+wVuH8ckMI5PhhWEb2MJYSPDg2uv8HCsklAWHnpbrCzysnIBi
DLpEQ0JmN4sC2PIodwE5PpWij9URVGBfUH+P/iANiinJ8+NsXyKSzkjF/gzOKAP8
HIJGMABYPxL6xPgVEFWKOw31lOtH8aUrGI0B6ucPQGc3xhlMKdkxcletdACwFKX2
RlOIRnEZLYyv6MdC7f2oRj/yDnPKhmLpNjV6yYNH+qHwR4xLmV7N9Hp2Key4/NA6
CwzI+8nMks6ersOtoxBl2FDo1NDmA5uVrU9nb3MhRLd+wn5G4qWX+CQDx4j/a2UY
U/gL+x10c7CKYQrA/APiOcGO9i1rYodzOJ2RIKx3/Rnq68+P72H8XLg6FlPLb8og
Mn9soBZtK8J2LlfjTk5qoi6FkhCTxJ7WUPYHouLNaQVawuc2tWj22ZFxza15+Sji
x+zQihGSG8oDq6jF+25Jee1yH74BZvDx1Zxqn9v0CourZekPfQ89uBFgW3F2+U8T
jukqmMkyMFb7ZV7ZerFNrdDqoyxGOzY6wCHcg0wvSkjhYmN4xEiCq+wuZWM183PE
eb+NDjIXcyoBT7b44kWrmdC8naBfnnZ3eDKDVlia/GMD260w0Ios2Mkqjh9xSSp/
7HMXziYr7bFX5JLRnhw1j7/2YWjfqNwekJXr5tWI8TqiFfsqZt6+AeYW2IHv9aJB
pIdiaWETeo+MMoBM8/Al098pvHT2XzS1MTkRoJxNnsBJUBTTF8GusdYVXc8tlTUL
H1b1z9Uc2teurcMf+jsMDWuaEBz8+xyvS2XGN5av5d6yUUzXieyGwMz7qg3Tf8e3
1cFBR0BJ9DBrhjmIlsCa3sFwjGCisHYDFzYNZlVLmgHl8swxWpeDPbULzDXyCmYK
kOtGK8/3s5PSrA+x9/iA3Agiz3iRYIbDhwMKTM2IWNAoh7blTw8y/swRyDFSUw79
gGdnhQS7M+6lD/qIlqQ+i7pLWYuvYEQrrmWA86XQGnrqsz1nhPErYKVBXZ0NA7Tp
+b8DSFqPKEYDIUPrycTfzLpyqQjApQ1Fk34RhYZPv+QhsLmZwTWCBdLTFJLzxlBO
PWWdW8QmIjQtQ6hBTfbFd7hMkylSAUYyCwCIuqnJCtPkVDRIdnAr8B7qc4aOmNvs
XGqEGzZg6yXaCEbK6OIUtNfJjMnCar1BZO6ic7toKqWC1cwf2F33q5988SGm3BbK
lw2O6cd+oovCnU5M3gVHrlyZv4lT3KhQwVnu9smTWJRHY6AI9FM1BxuS5B7RVvTq
2P1SUrmNesHEooU/XTkCXPqgMmK0GKn0IGxt7NVG4h9f9lxm6PtBbm6x3eBdOszL
QcdPcTaouyw/D5WxMVmDxAV41XeE2Dj/szg2QkpBHrFRqFbDMYEdOAQ2zBAQ7c+1
s4TKWj8fWWJHWNEWTtcjHoU40Wk9n/W3fInY03bCABao4Tdr+wNpJPt5JPxHdYW3
VpOGKKxgAOA/4oEB9X6XyTFBs5i0ksEHKgrAgyYQkTqHw2lgzVEPvQkIq1J7l7qH
3/V7L937vVyiUUEenM1OH/ipSRjFoJpWnNXlMVVjEw7qlAwkG7IbsTczps9z+ggV
bP/yCxKRHx1voPI6+Mh11wE1skMRUKKoBnQN1vZUpw/EIK8sYcQLrFnygu6l3elv
/yWJx8JZ8RfQSfG+m3mhiFxXoadeV0p7QFMeIf31x61+M0AcTn59pdV+BLAjFd7C
MlQW0ddNhM/rcvGadHUi9P2gIGq1TAxivegfaZupNtkv09mwbOLikhzvSEHIhha9
VUdhG/EwNSigJ80hYhiROSFvn7Q136Q7Z7NL12LU/easPX5QWsY2J/neq9uxFE25
q/BdqUbaKGTTw+R8GuxCRV+y96uD83Nxku29ec6LVEQy0NuljoA2vKqmTn7kMybU
AJRRKrmCI3KGAARh8dR0JzlVA7jXblWEpoF139T9/VnkuqvUIXpvJFUF7fmyK0G+
kRdFwOpSn7qzcJWFQvt5D8ctCviz2t2u4DZwrKZutb0snHz9TO0DhYsgib6Pp+wK
1+KVJMrblRuenTpz+saPBkKeo29x8+PhUqZbLq+4bHRZF/9PxKPJkOVgQ/emtsGv
GgLP7hH29c/uWCtFa0jipjAR6XLrV9CekOdSVi6fxAAHWAkb4XH3qfeO9Pqo7Wvh
dot26xoO7PBLVOA6847oGKUsgCq/ateBPu1Os7gA5fykZY1NKT/knrAOw9/t1Yvy
iSMfSItHzMOx2vg9R1tcgI58VWqlrPvOgQkPtLUFq2j2v67Aj532mSN6WqWIzckR
ZKKG4IxN6suGhxEuk3D+XZDt0TVSeLOXi4p//IhtUj3wz8upfT1rzB5cknP+e8R+
eUZjtn6rhE+bYwMvo+XzupsOe6hjShwWn2n2gCmCybksrRtu1wLHQZ0K+ITrXgpa
Wt30b6oxkh6cVurjLKBCK2mhsPBJ7rlS02QRJv3Xf4X9xggITP2nq2HSjeYiOpYA
OGCEsLcOzI8Z9fY5IhQvZiKCL06UqifN5K8L6h+e1Dl7iVKOHOX+cFFKyXjYwF6r
9qIFXjn46FIL7bO02Yu7jNQqqR6KZ0cOHNXXB59Xz1Rw9Cpc9mALB+qolL46Nr4g
F6G/VeO1LNv9U76/GAYMfTc7RqCBvMNAf4YDM4KTCk80UHUOEwSeZJa2qIyc5K7Z
5wAm2ir4P+aWzutBWpzDhO8PSAJW6hVrLkUu02hAEzjAkVn25G1fJ7U2RAZkQZO5
Kt/UhyHs/VlcBerisg6YTb+FIsB4KHQHYbLGXeOGAmHMchdpZtkqec17cx7DnmKi
F3/PGRuQhftfKCqLUSn82Q==
`protect END_PROTECTED
