`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
os49M3cgJCBWjtsDw9vBrr3CdZcrENplbsMZfJZtq95yZw/4V670kPEGyPH4lUug
9D2kKAsS1nED2CDmzZ69Vet3tGCFPNwmbC1htkTmIdtvDG3+HViT+1WIscoRntyv
vj7I4nsYYcbK9WMkZw85esFRth5vj6fIrc56GRCJ9ZwK2CD/Cf0Q3Jw6Xo3uzSYs
uDKTgzn4k5t2vQdEV+Qzfx04mZWikA8/qOlJMA0Eb9b4ms3G2JTVJ7u21sTSA9+q
8R0eyTda28d1OTalLd6eOiyF99102PMq6gfamD+fITQ88oGIx5QhWGf0P9QI/4tW
/Ns5rGmVxkECqOvdFV8jtu65Rx9SXgK4akNd4xjfLxX9FKBm319KgQ9IziCuL3Xz
riJWFtG9xcT67yaCsd4Oe3EuWgv4t9tbz7g2MYh9HmAOd1tl/b6G3eLhknuvfaQf
BdZESmOhqVl+ZMUMSPSAFKYTSKnsbXZku1nLajLh63kfjJsTT6+KeUctxZmXp2/f
M2pnsKHo0ClKFktj1GoZbYKSwh1VtgAQLNzeE33dMjNdx/vRc9gyesXto9EgdgyO
D5SHvll058zr9+ipRSOQ0RqOsloBmAkSKj7p0ryt+d9qIY/x9cnG4JI6kdk5uave
E9BefZm1zPjPK7EV0UEoVrk1l5UQ65gnZApw+qEy9rImZRyEPiAL/TkqzCZ6ToCh
mO89+0+D9p6nKm5odGyaubaueAHC7jqcC+qQi2kvOEkPYRCyem/Cn24BYbkZ4wW/
Vu1CCWYsiCGTZt9C8qjHS/Nh/5h1LUZ44fMH4R0papL1HcHGB8nvJk40L9J3krth
ljHcinbdwTbrc2he6hRf2xadt0Z3ze/aSPQcXwmeDySvUVAFpaDJTA2+wTfGZ4wq
3f04O+ki09A5/cD80wyaYrWsnbb2CnyiZU2ZDDb4HLFEz2Iv66mVn6J+mhd0Q78K
LqUCDKq2cQ3WO7FakJ2qK/CuOm5d/2Y12XyCAPZGqxSaXhdiUHmwmi34DNQVKZYL
Oep/O60vIIQFNoC0XtO+K72wUvy867syJVJhfoafI3b8mXGmN2ASv8V7vwRyPa8P
SyAgZowG98a8yMBN8XV2e/5sBcJicoqHKNCtrKcS4VM23NCr7XlhR4VN9sH2UOrf
RCZckuY4UFI61lcxGXiEPcpyiPqp4hEGPTXIAPYbpTfdW5H3LWjookJ2JZkK9bHg
YuTGkGw+jCSPgbHmWOf/P7Q9DLK/VaPDp1bVYZ2+yPeV2IB7arSfSAnJ725+z4QG
qxkDzgZbF2Q17V2bcQ0qWvABuYor5f1GSjB1YVwmrdjsPjE0HKQSaqmRM6h+1qeX
c8V/8TZ2+a1sb4CfiOPULJWvyqoHiUb2ZtbwA8+Sx06s3oNTj11TQdg1vM7uDABV
sKyCBf6fJQE8V9dJYMO95paMVg9z3a7bgpNbVUgVA3gCPTGZY3FxgWp4vgCwb8fO
mc1BFcOi8SitvnpLXuSz1QAcpCYwNWni81GSBkXtFfJcCgvFkSFnH9wewXtbmF5O
KmH1Zr597QHx4MwlW/QZ6CUhojREfgS+jWmpHbMiBFXFgpk92vdqJunUD85I1xRb
iolDhiX1EurRvCFj1CMYigRNpynfXI+fGtGxtvHOJ30J5Uji/e3W73EeFTASL8yn
uLoT+YdeX+J1uMU+iNKbb1getL2gyOjyM7c6HPnlEXlH2mLNnSVIHeq++3IGQV9m
dNtL8yd5Iw572jDg2SpodC91xMT7ovaij8WeX/GNdS/SiG2lpBBVovGOMo9XcAiX
FuadkbP2onu6A5wQ/q++tut4dVRR5an+9SpsR0vkcAW/CDNAfnOQEEyD6/iV5mmw
p7ttYWQPe6mwlru/SHl4W8bUCG7AfPNr63Oq8+puxE5V4rvSLnitXpxHAScCGSvs
nYTRNIxxLtt0/FvJBS8wrfMaax6fm5zpUUJnMWAXe19qb3MZEGBi++QWE4ZEcPyi
jN79yGJe/WI+1aGXxmTUoGRco0dpZhjefibr0pA29hnaBzIUiQjS3aG9bSZSrVxK
FkpE69NJYOqe8+FMwEzDe1IGIrI84DxevTtmtxpA7nJjVujTK1SPQwVy7QoWKUB0
HVrSpjiziuwSgT5w71VXAtqpd/nFHBvPpYcdwrEp3Au0VxeFaHnkUpqO/bWTMysz
oP+oE9ePObtN2qrN1zaxHM60w4qQPNJCx/OtSItyNRyU7aFVWMaAsxnVoWYd5ofK
kq6aH0uizBqMTCkWVIxX78axd1VM6lAE5axZ8gGhTFFNAMamMWD6DhZyOZiAxKAc
pKA+kqMeFV4s0Xhld/49Gr+sjJ9zAoou79MCBFb/JNjntAB15rTBRF2d8tnlf2/o
CUVcZKhMptKdURQz4tVfUW3IOyGD3oGZQtTwhBKok/tJdfm73awdVD5Ewn312eVy
yQYsjtf8mg2f/RxDpgG/iwYeqk0NAWwDSONOfwtk0SYFuewlRFtG942tKREmJ8C6
QHWtiJ+2w+qg/+bDU3aB4yUbO9di4p5jtC7DA/LxozEU9Fxd/b86JpvoJD47uUx8
XLmirL/X/hC/YLw2ti4EZKoMEmoki8THlS16DF/x/39QwDXHtAc2oJSYIdXxFXKS
Uq9sxjUVydh2bvg1o/i3og7obmDGj+5gpCb0wbs5Vi5wInsn/zikU3JJkzq2m+hK
YXQQ7sDs8b2ck5/gfK/mx0HTFbexB6hB1bHnPWPQpztb91hhCzwObV8jXYnIaAJ1
uOvZAX2gu+zH498XoSOTlZkVgh8xX3L0ke/DsXlU+W2Vi0f08QD88TcRVT9oWPKL
7xMsgaknNTMBDOD2nnHMbHV7rQFTNTZH8LAKlojDibydysdUoKJVqdIQUQ/70GHS
XXN0r8tab4AYlmbi55LGfr/f40H3QebKxidTCL597MIN17fGgPFKeU3pN9BNH2T2
4KE8u885hz04myyMKYRfipaGtNVJnA3IP+ICTGSMeW3fgkcvq8APdEBoPMiel0ay
o32qcKGVUDHHi3ZFjOUnvW+cf/HUVdUNDWRnpPiHAH3mk8v9d5K+yiazV8lfV/zq
3/+ufLiWG7kT1+CmSNrlgkPZhMKDjARHc9/SScOQF1HMY2Vsb7eEpLkYyhveJ2jb
b3OQGzgt1sRwpx2MyrvWoZNMINB+bkJKW7nIK87W/O0rEQQ5nIa9WZXnOjujLs4V
Ymjb43cPkVvaTUbCgtSLjJ/e31vn0X65plaviPN4rpQRsgMpHf1mK3H44s9jL0tr
6GcIGgG0FaYBnopWJ1mQ69kIUoRMOk4s7zjGP/Tde0IO2hcN9VD/VeKzy8bKjz5X
ikWYpPfmGRe2dP7HU9/pRDg/YIpQE8oAVXwNEMiMZmKanLP8b4nPfMPRIWSBzuhY
WUXk+fi4ZAlrbXpbkK7EaI2Am5rBCOOvy+ntNtWxX9Chqd5QWEcFEsY0HBgaOFIv
x/LJ2zilE2Gs0N87m69KYM8OCsw5eyORVv5IUtn0iwGgzfmpIaDtIwQONKSPlS/l
Qu1a61VAdOOH02Jye6yO1O1+D+W3wHINoj6xDYe954tDpWxzsTXogt0fDmOPVMvR
OOIO1UUyj1VgD3b/csYxfracTR+IF6G/1XFDK7UrY9ZdzD85Q/byBa9UfO/mRKT3
9nosnvtSHbQW9e4beBTcKjSC2Tx9UOVlK5A8puE2+6t/CSWg1kZVZ2HhJ7zuq7Fn
U0Eu1Oy5XhU/r673BeZlarXE01dSI9W2EBWun4PqqvlqHHa/OkEVxeREe3NbgogB
nwSBmaT8VF0zhLKgdPqy/YTP7o043tKaQxgXOD3sFMCv20KwVmh8RxBlmo44GDeE
m8slPxCG0Dt5EITEfAnMwF68mSnC/Ru8nEMlycB9zPle4jcAAEgQTiohfFSZXrfm
nZVb6y8ChbUueQF9RbO/wsqD/mdCyvxjDW2XpqFcJU81V5hCMf9iJ+VcgqBD5L79
618Ryp7n5om8UEu9h/iXwlob9V5BRG1FEu/eJb7+nQBLhAFa4/u/qpiQrBrrtTjE
tnpPrE+EbT8mIUhqDGTh8SzQuLOVXofQ1wq+Jb49KE0R+DeVWtzY5S/KJMhQzk2Q
qGgJ9SulG5fev58FtAnzvdQfOoEvALHh4BD4tCp4C3JC0Qj8BVuPEwXHCm4si131
ApB6rl4NbKco+LCNnydcN+QdtEcH6p17fh1N1yb9RBbwEfELWu7WIWz6wYiSt+fP
5FU/XspxrJKANV/3V+2jVRxxvsBpe3iR0JUD06XBr7KY8LTMp+na8KaY+F0uaXpq
N795yY43ii+nz3A/d6muYmBK0nk5uPKXvkjG1TuODnDHP4CXkUVEU7yWOsjxKJir
pjeUm1Qa0+kanVkHlOYk903r4tVqnuAi3/gsDUGgJ3Z2xwUYI0BP1r6LLOR0fNc6
Mtu8ZGDFnooO/KwJlAz26go4Fnt077ONnMCKTcMiw9VBMJBd8052J9Pi7KA0Gad+
Tb0emMD8SB92Rmio63Z1xL2Y7lNxZDVz9k0iuPq4+JwzyvwozeuULyB4BQi0YNV4
GrWKIZaIuaOKsIQeWJivWNj7SeqgywikhiaxQ/r9K1y6Uj7NDXlf6a5MHdMqSii8
6+ms2/iNQC0ZS9rFBdxgpPk7BhjecHryXo4XYJFLqplVC/hypRAHZeLSSgWKUWid
3F5RphTuXmq2081eP+sfXMNwCCUfxKFD4iVW+HdWCTLctwd2ybqxCYZ4ePH59XQ6
PPWFiCcORJX1dULP1l1or7/sfcgQCXasuV4JKFqgrD2FtXPYyEB2h5Z3jwPM0ndO
HE4zqsHHJfQ9wAxJ5Nej9VxETXugeHz2x8s28zcMBJwikX6WSDk/O+9Z4Y+9PzdD
D1dp5Tnd+k+BGffE4ki5ype3jfKDGSNdFJ+LZMRJCZLWeD2bqVIQKOZ2iepA12g+
rZaDAZfJZG0UXP+nyh1zvJq0O6BbcLdHF1topK9lijGn9xTpEYyQWaT9uSTtBj/Q
QN2DMSQ7AI9ThuAjUNGZH4q86DfqAmUNRlPG3cag8KDS1eg05EzCiC8C0OcpqhAJ
JMa+JzR5X+DUoNFoU8Wo7FVqN+6mtHWmBCyRYjrkv50KxspPw95OkooAZvqGc/da
b/dGjAGsMLmABPJKttd7DVaEWUfxOyD3BhX6yf005IffyeQWWxqmKpD4jQbWNRSv
AHUtn0w2bPGKJ746jq62ACsYJ3sJSqtz7apMNJMkRZOkyghBh6lW/9wM6hopKBFP
TJcVyPDvhBqwV8Ypyz69fRAjclVd4MckfwbdUrqx4Av47ZWtpngwrYWH2wyfubPe
c7T//jKR1UGn1l9wqu2LG2QWWJAUTeNExC4n0SKD1sarJsh9n6JFA1AI43xiSTHg
L9dgr2pNwhKpI0UHSjvaxwUK7KOoTDM7+wFGjkNl8qwehlKrFwWwR7yfJti5Vq9n
NVqzEpzQvX9K+ltgv83Sqq/VoevqOToKCHV4+46nNrRhISb5wIQeZYEdFE/cvANW
YUOn6CbwCiwpchLgwxYS9qhD1Y51Hbe3L58LccBgWriOUY6tk9XPpkZi3KVPErwh
drAC/CUC/XqBoGyYdUONmB810Tdjsd5TMaDv6AKRF4T0TpTApUEHHCMtGaneolNl
BMt1fAZ+Phm2BUPOrQWnWNAt7v+NEGgjGEYBkWk17JKzdQs/I8HQQyOrK1/FCAMd
LPSNgY5RAMl2LXdic0BZGfA2DY+sSYVit67qvwnTbnb4rIugqsRrLDu0PRBYo1kO
28oCsg6LwqAwHvWTqRWRL2+Sw8ohbtQybgKqlhRSc9sV+hUgGgNOru7J267+Va3x
Om0dPMMvXvvrx30QWWh/dVECOyeBlPA5QZo6HcDDGFaiNLYipgLU7MwD3VLcwdMO
M4h7doutK6COPiFvxhl5/sJ1A9QMPzcrJx7IZTJcMTyobGkdq4J2lL+QxX9lEj4Y
4I5RGSx+I/s1ihNyHIwiGmVB7FvT+JfBu8XJPmN6Fj78E17330avb4cQQWzmUuvJ
Ng9Rs6/MzuXw20PLDubTGl3UGJ6bUkXr8f6HqyfMVZdQG/UQV41GsD6avCCgWwv/
ERmAlnzeSYuFgvAuDCbVAtzgpQ9L+SvqK26Q/KjZ/ypGbUfIHFZ9fhUHfG/okkie
nCOgorJGR3T1R3lRviTumqnzaXDqgTwIToqGRCsrRr0gfDEgks4mL4J4gKUqRwxK
3/B0cE5QSMnQivuctYixBFv8X+9Olrx0r23c2iFqYSxQetvYMWC7pBCLeeEIS8i3
396lY1A38KymjOr3HoX0TkTQpAuryohG+8Jyti9pyG31F2MdsUlkgM1c7bTIA51D
BPH1iRS9qMLn/xjizg627Sjy7fjK4qPqB+rASo0Ktp1C1SguukYmGAHi9Fn2BuhR
axyvtAgB/Z4zBHKQqcszF4EkVVC4lOFmLIKjZFC5rIx0H8Ut1z7daykdxjYHOTDh
YaXMpiiWhNPVZESpv3bqQ4zFp5yA6XY6VwJcyXTJUfgR8njOWx9ZZqL1ROV/Coji
pjqSiAvw5KleUu3CrmPprQaV7U0grGKidMHWMkI50yWCCrrZjvtuDVkO8Fj6evmh
3ht5AJHefa6XACxmrl+buSQQMiMIhB28Lt+1u+6/sk6G9OMOLM0ViQipSplvat5Q
T52SNeHBlp7pFNXPRwiydVSlpLpO18sY7zt3GsBsMy7ax0aqWtSXCZ46pvnI834a
fM0tcdJvH0m6mPefTD1YybsCA5T8vENE9JuE6vQbUDayZfz/gOBzrMnBWn9Jb4rI
svLCsx6S+nPxERwMJ99bN6SbZnoh/wNfToT/YJl0fFYhsk2WUYZjJkm45QQ6wv3k
y3HnWBBJk9E02ZAL4NMo2t+aV5hZavwB9TkK4TgOBkEXTJiD8sRudNdet8Q3qkUJ
7KPc3OazxzqY7pknSgqcCvsa69ObMtSxTxxpGTuO4rFMXFSkZONaXQiSFk2VPksP
Tc4Ba+IwBAXnP6c3bnxpB2/eb9NH13KJWVFe9L49cBbXE46KPkIDZgfUzfLoxisJ
v2jo/WkKPbDGzpF9C2ZCHWYNWIhTP1jfo2kjH5COkNjpHQPFVmEoUEpMDQhzdkd7
VOegrt+E8Z/sp1ecuD36myxfXBBs0NiUwS5VxAynkl+X7F1DJhj1cOLvKfo1X00r
6i95VCc9dIZ8ttjR1Nx020FQgYrd+zLui6+6AnQMrW/hEiFB9U7VulRWW2sTdYE1
7FIl2onghSthOM8Bbrhdhhn5az9tZ0RAQeTrxZQYpN44qyZ0hDT5Iv9dA9DOg8BE
ThhbPp0BWLXiCwsNYZkLDLKIpd8xOa7N4+mgWcXv/RBwL/St60CF/BOuD1rYgzuq
Eth0tYHhPP/55D+6ooOMtArZWkcRipMZcTXTyWxluZ7X58NW/778lPyFgB2R+esL
+pIBWKFSoqJzMlN4E6Mp2pVxj/Bym6fXDiFnvWHN3dohWtm1P/oGQv4kRewZHGDI
mZ4oGIc5RRxHNq2B4/s36kNCDM8GaazsR78ulffELkw344HceMO61KAIchnMN9/R
Y2jUdQ2AgL74KqGQvvD/Tt+MpYLZRcC5kzzawqwT6dhA5ohHlfLVuXQyJzS0R7zQ
hhuOI8JwNYtwHgDgOFQmGkyBeG8wa9JqtkCNiJ3cPkVeERvvRgCvcVhFXOROh7Xy
WEisa00VEnqK1r12gFexrBMCM18IY9z3SvB3LvP5MqYVqO5FyFi8KbAGxI19PnLy
tSAecpJKoqfw6xcwIduPo0+4Se28KokJ0NVzWjaDPpRSMoSzk1+K/eLUASEYsSVR
cwD1VqUimCFBgHSnSV4KtNhVwYjLO/Db558j22K0IyQ5qmiK9Aag2dKCsPnY3Uz3
CDiXZJgXL9XKMIfPPKvXo48c8Pxe2CRTsKtfzOnpYywtvR+uOo33MqunO9AyyWQe
tyV95idbanZCuvCyotSp32o0w+kgMykut5pHDiUQWe3xBs/sqIv1qDj9QNgqtTZk
NIti1ol9F1NAuu9o3aY1gdnuvQwhrhIn7JQO3pckSaiTueQlrhFfV/lv4hooFkFD
YJ63DO1sHs7JxAJR9TXusXj2YW2MuaVZ+Fq3CYA+SGJqoBUxSRslFRXLw9Ti2hrc
ObijFZkNFvwfbuRbhRtpuueXPBAP44dpunlDOYtwcaXPakH++MJZXXlMhvOzrgxv
jPuypbjGwnWQ6SQD4ptCAuZ8VHEsIdRZC+9I5FVc0pHFPp2PbhZk1IPEoVIs4Umf
d96PIj1B44wa7OjAUxdgggzwf8Mk8HaFLDhysdL4fDpLC1uN9xevIdzM9VZIaBbF
VUKmUwTDnqhInaQyt6qtWP8jc+6AdZprkjTQtCElkVF0hVs5BeJ5Q0HzHODHshsO
lpEM6Qo1zDUD879OoSg3exBTvB6ixgqtt3GfSRThRZaGj2Av1REbiEvG2Q5MMyPW
s+5rUS++GmL8w9infGwKMGgAI/X7b5Aayt7/BdcO7bWjLtyCQ7JKbRDV4FO5dQiM
zHnngpuKTmHy/vFwV2pCkxg4bIJZv8m0cwCTHDd8ZwS1kGjcbjTYgvifZ08cdhS4
IwMaeUh4aS5fbLURlork9yOE5eJ78uZ0fKOq3m/4GMvUibeUrg54FC1yJCXJtWRt
N6XXfo6O/L2WHGQTfgtMFxVQvTyJxo2XLjKUs7q3/dvMjl1s6eLyuZsFEQgqYIo1
x50l45cmSILtN+kmu+8EfuYsU1MIdfjMvNJr0IJp8zKulV/RyTQtLxfADNPRK44n
7p5t0BvnJeT8NtQaZ/ppQM0c4qVm1VtqD1J9cQhLjkP96BiybdBu8mzzFJETOkYa
rI4pj7cPHTnNL2t7RiugAcLZlwkN0C+IFik0vJs0LolQJeV/Czti5qB6Yss8F8Ms
Hx+MPlCzC+QCveLfU3t27rZZ18X35DXiiIl0QPHHN6GY4prEUksRSaScEKTQK4aM
JD5jX/QOKE1fd7dLJ6GOB5DX/thRlnYirKZD0KyWA7rRcHWm41N9vHy9wv1cKNP0
DoANRUFQ5WAFXm491BxW9HlvesviJIzue39mmcAV77NZ//bKPMXBeqF9B/FKRP6A
bx6kUJ0ilQ56AZ7SmwxROnr69RoZa+Q5IW6biLTwFBOrTPgS0uMkZkHUYaD3cv+j
5UcqE8txAeirfPM89tZzQwQNUlzICPdurt6lHmB+nOg6J17KMoRH72mFbNyTuuot
F2Z9vjhxNk307mugM3Z2wKd25hr0Q3dXI6yBN6h867wmphB2qwRgK7OT6jzu4oie
rsAqtSWfFSoVXLSy2+35WMVMz6Q3u157qDDD5Tgha26I6E6F836Lg+43QyykQlP8
JdeQh207PhTMmvVjbBRl2MgnYTbbw5CQihAd4Ur1tFI7+ekip9xa87Id9/Vg4IH1
KlP5AbAORsFlAuvby/eKgKYkXfalc/f0lINsZdLNUWxsTAwdl8PO5BRtHaFEyecF
k+Z/6E+S7T1wRSurzf5s8TwoTuTqMKEwjUZJJ9HiiuAGhwgEwh/2YHYuyA28AfMC
hqj5WiuSGgFv50Znv0rmuDJ/Ae59K9f7/ncKFsXAXYH1vQKlAI+9CSXyQtwiusc+
HDwJRiwhabfvdY7gdJfzltPghnfvhzDtuC9NjyXuvW4edc/fnUWibCXp76i0r2lU
KYByJ1TAF7PHaaVNnaVR+G+eHhHfPRFDEEdj26Cx/ktlKTl9pJsdkHUrG3OAHG8b
FE7IWLmdyoqf3MKS0EOT9xeBnQzqXY7ijrFRqtxaITg4CVtOlEdzJsIDV1ozSbMb
Ly0ohLbI3BJY29fHuMsA+m7M9GC5Dkg153rpJx+qG7rEZHtAWzneVRR8tptrscnX
xvBCEN1eVWgO/8iaoEJYTd8umRHp7EDJb/reQ/Sv3D5pAYXzgl6rm2jSbASuxgVL
QE/YlnVoyVubjT7urpUEe+fOR4cIWLocRzAlXKZ7vDPDbfXrfGZAMsLfaIRRe8sm
eaTRZvCvbqCSwy01aUDee85tlUZ+xae2gT0EbSRtwX+rhMDSGagZBXlsaG6HtIVI
+rLeO1Mf0wdtG9lTv8VA1PihREmaWRJ/QNs1A9rjiiko2b1VkZ0ugtVFl8dlTKOj
XABjguSGqTyPPmkFrHdsfX7/P2LHU5pZ8A90JGl9AVXbM4lIli++4rNZBpbSBY+o
Yt/az8qdHvUvDVWSEe1W3u5qvoDgEKYwQyEZMl+dpi3pgT7ua/hmLBIiAghf5quF
ppOLzQGihCT3mO7nxwoyC+298wU2+E87sp2PHsdvetIkebHX0/5WktZKOLBGP6yI
jvg7sejNnf7qJ2jp8gUeUgBi1cKN6kNdIII9BVlcdI1le/uYHxk0z24W7oMepanP
gKcA2S+hnoPfTXqiw9u/Rmh74MbuUqJI9eQbd+uwxzQ/2w/12vqdsTNgDBuAqXiC
EJKRKaSIY4Pdmk0swqZwmBKv5G9ZMAf2k0eKGn/DMBN/61QkEuhqVxUQFbIwDYdA
bvaQOhsoP1mSh182wZIsqX/WQbgDO+E8fZnMybAu4MftAEkhZnHexsOitW1HEx48
1eCi4kupQ2wlv35qGaxrQIARmlrLGTSnKUzdUpZffjlz60ovJuwgLH/mrEx0RqOO
etemfVB40HsT7u3V2zteo5dTA87RmDTQ4Vc9NMJP2H8JdA4sra1VQn3kll/I7ctb
M/WV8/5YRhSEZDvt9Po31JWYDGhKiBKpkfktbnm6jSZQ6jmUDTd+t3ZQYtVXOy+F
9Ze1vbVqM00euV1zYigGP9U/mPZj7klMCZKrdvlfb0XR8YcZ1EgU4AWt0kAcDqTI
KpjGINqs31I9RjuKHLu6XZcvDrA3qoIjnlIy1D78D8HyboyDj1Hgv2memfXsHzt6
J1tnZ9LNRYjcrTwwaWwiELXBgtXFHY3cnNXZqrripFnANcwGtxN6SFyCl0x7RHOM
0yqVVkvj5kfFWP8quYLLDp7+SqtSKEg5qSyaJdpt/BlJGjtVThBLvN+6p9Q+8sg2
Ip1HjYfRyxXNuftZHLR0+h7nMsS0qSpHQY7npv7iWPHOzwx0ERsF1cbSpAuMjD7b
GexYJtWA/up4MBgZq+ybollDVt5TJs5laFnt6FtVGgz35gEVIQhDS9F9LfhAV7lv
gNE42Gvo2w76LBZdIFdKxCbHexgNg+gTMWaGUjpT6ZMXiJx8tSP/FjXnclBrkZcI
rlCj7pueZebpWstVTpHUmgquFhLWodTbGk0v6Hho/+MOaZOqT3bzu4558MuNXfU+
EdWeyjTl+wXU7Qv91OJl3IhIsE5DFfIFMmkuwPtwDLKXBO2JoJMq4TezUxs3dfBg
W5Os1Q0RR4XC4vsO0O4yHu4ob3sScajIWTL/XqdaonsYtyB5wSO9fBlycXptXSiO
+zcJAEXYnJEZy/THvUGVpbelJYnwjodmC+cdxWXAtrukg0TMHyChcWy+QHyNJ1wn
HzxfDTd9CxPg8It1eMAn+Znb58yd7arZ71wMblegrGj0IkrNat+PTYa/j6hMXMQU
TcHXE6SucM1gnJ50B+WskzeayQuozNavir1wykikzTo13EiaM1ykO1o5TSwm288x
iayI7XdaX1yS09AiW2kJrE5WARP7iQ1xXi+55TfVILY9UIdxnzbi0GBpL2HnPQ6b
dh59tjQPGmcJneKeW7PJycHTfTYQGJpG3wUxclLSw6a5eSjTEKWb5iEpV/HNxtI7
ZM3MXY1gRucyvboNSaGBzD60ixg9erl+nyQ/fGTYivsnKJQvNrbHFJxQl6vnlJc5
4wTeYMpslvNHcOCMS2pLt0f4kCARhihl/5L0OXyn9ePq4vH/yOWyg3Djt0qJaWIV
nBjTMc8yo6crNJ/2F46gxTt6ml/KmVrMCBhS9s1eI7lvEuoPuqZ+RgFSoF6Jz3AA
PXlAFD5MxLiOsBBjwqP3S3nOhdyrb6yxWrV1X5RWZUzOe0pWMjlgdlfCt3BQuDj4
f9CfkKrd14iI8uwZxSy8CW1rflbkDZcV9z/Va1Iufobkq4NGT0ES58jnPoHBv9P5
OWSX9LWdMMyvD59jLu8pFm+8XFPZVV925jeZ77BP47WNJ7x4wc8Y2p596NBDI+v1
3MSbZj4XfvTOWpmPtE+iNhTyG475mbX+q9VClWgVAqbTEfq/Am9yYORLMHaumch+
Vl32nakw6/F9hg4Nq1jU+vsH7B50cOEUCjNDF84cOhstEbVKoYS3kJlgQsapMZrz
/mqZophC0Oxsy8wESS83hIHmMkuXnIqshhD0i9UQd7isKfYTYUUvTshj/XzcnYAo
jGn0r8n8WywlrrEBrkpd0S9MamRNooB3isD6xy/LaYxe8kmq31h6SNKpaLiK4dCW
jBJIAA78gCSoxRctJ1g5dHf2PJBZkrjicXdWBmYNs/nMRG76jfnbf/V2N/7iIxt/
6GhJNRyC2cSkpw9cuYFMYPGrju92X4oho+nCvMGZjFdba3t4Y90ExuSIsmaILWs1
JRc1V8LHYupjgMYlDsJNz7tJ0MJ4xQixfEFWz+hdEjxHcMRAnmEXA6GplDBoBk2f
kvlJ9GJTNfUoK3KY8mWXKdMdGLeW4YuqRbHepWAvy+V9qtSPXQsE85ZKbUPi9sWS
N47x5HRnO8z6cjtqlGlWy++gkehnu0F+8N6QGHOrmfrLTcFkEQlZR/8Y/H9CCD2P
P/4H0kMIKqWVn77pfPKGLQjczlVWxUKnxaByQkXkFIKs8d87+6+yGxTUVwnQZV/a
qpkh8uxGulSKTU9xl+ttn6C4qlveZhJau6gOC4rq3sY6cGiphVm6tHym1rILbEsX
F7rUbMpEFvpoELxy7dExG1ATghXbVUmQL3WJvLD+9K68xY6DFaW3bk9N+5hZyRau
P5cgfXUcgyJxEf2m/usPxdoX9WIseKavs6WqMbxEV3+ZJkG5bK+QWI/z8iWPCDgr
ekNIp7uQ5MYnuWvIOA91JCkcNLSRKJRuZW9KML3g+7dJZZpsJwK3brWshSCLMS6a
Mzila4unNFdkL+4RcA8z9DpduBtlACF1OhT0ZWe34sESLLJlqNc1pFXxMxkKC8zH
6nUgMtH+uMO3OvxkeEqXgcKRn1qPSjKrqTlIhj4Aw2yk9yVxMuR5lNYauDnp4p6V
aFJJVPep6e44Bokbc0UwV5meqZJKgsASgUTfjLVNgXOlFfbeZTDRhXDlKn8B8IXy
PDoNhXNBOz+l90vQD6XPTGzetqgKolIaLoycnIIC5mVSQCx5Su6hV0d0mkykkeMi
xUCDoB7PyBJ9BA+mxdosXyisjBgV6RnNiLFCK8zvKvJOh1B7wbGWrqBdfFchU5Rv
`protect END_PROTECTED
