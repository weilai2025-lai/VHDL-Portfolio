`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oobzcUMM4J9LlC7axy0LxGSNEFPNzQwbrZrvdl3mfUWWp2xmwjviGr6CySlitO6B
qNxR+PAyA/QRZlzaVbF4XKNgmFj6krbsO90RGMRTcyrrXuuvm25iLDXL4bl1cLOI
i+GduWMBB8Zq9wM7srHSwYjvQCcE4X5WXC7BPtFDJEsTwycC0PJF8ckr8tT1NfpO
HN8soLsidVkc8fia20PNsXq8DoiBY/ee2QQvjCq9p9QKCGDnsEFraHmN2CnR98ok
HmEgDLuEoyhhj2BZHgzh9WaAynzyPR/LeXC0Kj/JFKNPDOcXfl3eAHYX6s26wg4D
VzGVtG3QRiLp7aq4gcq6TYuFQ57UINFHTzLD79YpJUkb3uVfDdtn60mCdMNoQ7eJ
gOGZJkIMQ331e0bGmh0IeQ==
`protect END_PROTECTED
