library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity fulladd_4bit_generate is 
	generic(width: integer:=4);
	port (a :in std_logic_vector(width-1 downto 0);
	      b :in std_logic_vector(width-1 downto 0);
			cin :in std_logic;
			s :out std_logic_vector(width-1 downto 0);
			cout :out std_logic);
end entity fulladd_4bit_generate;

architecture generate_structure of fulladd_4bit_generate is
	component fulladd is
	port(a :in std_logic;
	     b :in std_logic;
		  cin :in std_logic;
		  s :out std_logic;
		  cout :out std_logic);
	end component;
	signal carry_in :std_logic_vector(width downto 0);
begin
	carry_in(0) <= cin;
	cout <= carry_in(4);
	generate_adder: 
	for i in 0 to 3 generate
		u_fa: fulladd 
		port map(a => a(i), b=> b(i), cin => carry_in(i), s => s(i), cout => carry_in(i+1));
	end generate generate_adder;
end architecture generate_structure;	
	