`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eOceVVQG7nUvLtWQNf+XkSpxSNC7H1HMf3/yUX4DMRkostwFAxaTyvA6WIYddCl/
M9FNdTSvYWsHHBgHobDQLmCLBLArHT3GwwTfhfLzZNbKTotHTj+qnnJtsAJ/jDnN
Q+9KhNs2LMjb93iKVZtPDVeojk+NjCJTrQ1luu2C5Lk7UAV6IdedqyP3hUyUKevg
qcutnPVDu2WdG1S0BoStRhtGJxDQPCFl+z0usWPyZ3wj4EpSyJMxvFop0eAfGpPt
NcEnZJ9rIN2eFhD1Wu2aLc7ccd9feHxnCkxjL7vy8AQypesJM2hV4EVcX9XQFuYa
pHpSfE8V26QU7RVwPLyBk4Uwqbat6iVg5kTFLgPePCqGGuOe0Uq/LkXslSVARIH5
ctL4NsfEQgS1OVb5YFMJDS5GWlNQZpej26H9RnqhGtVhExkdKA2dazqhWQxpt+nP
I9oVohVtBvq1/V7jsEU/Wm3E4yDTYntAjfc/pUrD12c=
`protect END_PROTECTED
