`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmfDg0oztI9FtGQxKXjB2Z9ctMM6QsDwjWdbOs0Fg+TW+VXJE75FEywcUdr4xsz0
u6eDq+4mLNVl5QYJNSdjYyN8Aa8mA7yKHJFzJ5TRW2kpmPM3umVSop3zrLag32Mz
KlG/6NFrGYHP9/jd6oMpYGDP96ICVnfMarZ5n6TRH+1hbmN+HXv5NtRZbcnY7eQe
uBXct4BlPItVyGU8JKZFgMgeDB44QrNXsLB8xiaMOLyQLhCr/D0rp0VtdJPR7LjP
qmVPeEBMQsyoYAUxeW0VvURzNWmSbhmcx0nhvkVgkrK2SxeD3EQC5WBp3D/CgTgr
gyxX/CM3A9F0wz3j987kPf6OwOBc4B81oUHXkyEzXB149M3TUWF7JefLTN0H9phT
6XayGzeCH3ST9UlW/WCFBHBI/pPNoWJuKW1rUbE240fSQIw6WimejDxxols/RBFr
bckHGt83krRIoqP5DYJd8873xAd7FyO66Y0Vm6/ChGRi88jr4eUOvEDh4NouipHA
ht6mdfdYDUxqMv/0m/IIG7fGUyJAY0/A/jyAzDMSKWF4Gk3VMoU/JFAF+k6++3u9
ipJ8zC1djympEO35lyWqVdyGyIXDVRuToo7KFqCTJhXLdP1guDqp8QRJ0g7mkSih
ZEea5buTMKVgctAh3C8hsJINObFs+jd1FqQgrIptEdSmcOClE9PXj6CtPIezpYx7
l5j37O8yY11Bk1GbwDZADSVPZ04JqYJFxDNs+A7dPwZ76EMRVRTk77ijomSyNc33
bMnduvne4LsdLi8flr99QmPCK45Yhk5qPp5uvTmOh88IVmsLMxrOQN6ox/rC30Oh
pw/eoz0caBJLCA23pFWAHB+6VvS+xMq8R5SqXlz//nfWhuCTbz0Cbifn+Bx9TOlm
6e22m7ZWzv/6+ZH10mKmkOAdEEZ+LCPeMXrw6x2OW7j/iWO6vWQUru6xrzEk3O9x
mJNjE1z/q3h2gf0jwrakgCZAezP97O1wW6Wbe5TZ4QbxTIMfI8ospNJHAEjNaZWN
oN/4QYj7K6QiTljHadXgHFSbxz9VwvIVOu3GTQ1Kf0oc28ifo1tpS0UGsgNzB/tS
jPLjBzleiPrfmrm6KOX7OTHfz/9N4IiRhYcK9xXbS7NuipjDfoqLDpVNVTPC3vHS
i0bG9LBKKeGHv2LA3nz/2xceLhQoqvJULUIm6CrOCE5JgRp/BGY3LEGrLoqYxWME
0VJtfJQxIWUxYxiuvo6ykw==
`protect END_PROTECTED
