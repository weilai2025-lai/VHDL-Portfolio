`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7sc+abMFSZNMpyKC8LLMHBTEijQ/iNnPtDq0N4QVyXF3OnabHh4a0uvfeT9g/iz
Bb3+AdNuOBP91RkkdXdCL53AQq3ugyZd7fXIEjC1cCWh6p1HzSx7j9mpheOAGJP4
2ZH2rghNhmd6KJg27Fcn6rtz//DVuFkeUbp+VOgXoqUP9mTm/WAMT47akQ8AAsZX
D+h7MiRAy3UkzFRxqmXSUFGYQYprSug1nZCe5D3NL50CoE7n+C4jQ4P8ULgVGeSi
U9PvIcmm2ImOyiREZIuGEMAQu5xLD3jLmzsBeR1rPTmZ6Mq9C73VB7cr2nejncQS
fCVoduNr52c4EfENXdwZA8aXE5DafwjtEwa0PZABeN89fjy88RTAO4mhobInWvP2
tT2/KBTWmWTZniImyhbJsRlm5hKVci6FXcGxvcUuC9XSmbkHEx4tMEVnJbUpgbPa
BgDC787TGc+W6tQDJbdGPvPh+f42j1Q3GvZ23bo8FXTpFOZvtbj+wFC7dKlv0W3d
nQ6ds06Wm8iTNhMnZK68wyIx99A5I4aArqZ9Q2L5zssNs1O14dsXR2TC+YwSsYqW
/YZ2C4PjQzlS5qxIyBine6btJV5lpuonqkdo35xujgVvHftwdoPwMZUofLxKblTO
LbnBMJBenDkQmYXIExtfnA==
`protect END_PROTECTED
