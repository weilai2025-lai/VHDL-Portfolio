`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ozhY/XZEHSLssTgAQHq+KGDtLFCKgG+deFAOmvz8W6Gxy8ES/pAIwyO+I8BHlQG
Xf5MNO2KO3eaEOL6l5UZnWcjSy0tSv0i6y3bnkoQUDLC3y3xeUJBL0KtIOGfXNTB
UQVZGHOj7ZBS2fZz4zX0OdSBMdCj6R5bJRsaj+N80iv5u7bWRzBIqb7KsD28nv42
v5A1gzXiTWXeVzfeb2LPcOszUXo3yLjkEP/lzhCFU5XZ1dXgxHFqh2ApN5m0VxyK
e4euzgjTRC14PJPPTetTQ+p/7rkshGwA+Exhwn1rNWnSIRe9K3Zm2sPE2FDhjiAG
u7OINhzYfrhvWtJ7J22YTU6xqk55Ui350zPj+Yf8Jv6UXZiulkBK54XdOwesjJGM
gKmUIN5llH765QRtuxJV/6pJxozIdh4Sp32dZI9Bm71e2ad3FJsLuF0vSozomw08
er5X6qyUMuSIwDTNeQ2X45w9nqJwaE6J4gakeR4dO/IhGUQC3P5k5y/6uMfD47cu
jtqc7QyXhPxukJzcJ3pDKHppiRU2OguxwJg6Jo/B4HjkykVi2rjR04nAzGYsR/bC
mic8R7gEG/hZXxzle7gMNv0PRYKsveoBKmLmsb7p57OkDcsvzQjZ7/jihmNPrE1v
Npr9HpVdMZPpNHY5BtDiXyz+Evt1i9GEvkfwGP/OW/pxy1QH5DfM5xCIGQBKUCTb
UfoM7lIX6fm5C+9smFpHQxVe0KUG5hm43LG0xCQJnMdXdtLDRUS7k3HkYQJBAOCG
K2iSgbLUWR4JFVo+wPkxHcHnnANu61Zjyhsc02JS8X5kS2mjbHrhkAcJwrd2hr7U
RMiOeYbh8ZVKey3wIMnSO06cnutdaODuu3aVXKUMK3tYEh4oNzKK6l9dYO9nCctq
H2Tu52kwCt9o2hU/tRKRue0Umzx60fRGo99RFjSAKSurC7oXwrD7CtFk5Rhj1VwW
wzOYvlt2Ap02RuWVHHTlzJ44Kqg0qSJW8T6QTL9B/SQg2bJNZbR/j9kv7Cm0vgEl
LFUBmTRX5ZZ7CrxulcTXeKCssuPyGJz4AQoG/2u8xczGLznMzbL8xitt5J4OA2YM
yDV9yMtQEOWxMo5wsAtVqTK87K+ptztQ5oNATYGK1EgLsbZERys3Dptgxu4uyDMC
JQfWHKE7hsKl/Af4V7YQUUAttQPl64N3l8m1lpob0VuaPwf2LGKSoBdYVJNuJTDX
v8Qlv+MoI9UGAsfs2P/1uoYnG+wGN8wfHdeFHQuN7vTZMTWdhuHvCvsHxOEcP8et
LpMZh2JYENRWPN+fFxMx65vJTMH8uHIuFOWMYF99yGrCmss9pZJjlmBZ2VsaePaQ
rWZg6gUHjqx85H+7wy7jJigqg3R7qtwXLnJPLx6/79xob2ltahRGx+VeGFntC7Or
AIirWmt0xDpY/vOks6MdiZsvAv4ynV+bxx838enw7QVqwhJoP7KBJut8Z5r3Wplx
+7QrURlCGAglfOKCdyekvyGUOqUzQGh6uEo9VaZwoQbFSihepb9kiahYEKhXhxTS
i+6kBRMzysI8KW+argTylhlsOYvQLhMgY3yjmzwGtQzH38ro00ze4n13L5VNgXJV
fiIFqJs9lNuKnwcI2qFDblfxyW5DrvOP2G2sQjPD5UtUhYyfLCeQXAK2q/iN6sUP
8toEjMwhQGFRId4DiVJ5M9R8evXdfGCO9fQQYkGv+35AqORZp7fPnzhvOIFJ/Bum
sxHIidGkeIcEKC2lEahLTXWODgTfmGM/JWy0jA1UpBjGmU4GWBskXP6MEIzTqnv6
43n9vm55hNpfmsfzFy0zn3nsnJlW+XZJu4cM3JSGWalvdX5qngbNatA/5NTuLcNl
d/ktQNk75XO/rR4Yf3oTu7EJPSgEg/VEYfqBA+jGsmRlZ/9KdaPQApDIRBggH96v
jlNk9+XsqPaIWzf/RWXeHlJU78y1jUGEv0DrvIupZ4f6dSwmbOVwqGbB6t7wH18T
F4fdGdgLo3+tpt0+DZeu7dl0ONxlfs9Q93rmhLHFlEZwTHzcoYx3UB50+34D1YEP
TK/1VO+WV0MSM5zwZNKMjhBHzk7omz1p69S1hKUx2KMi87YQc2zfB4TDcHobqW12
YAiChkHCqet/B6OyLY82hWF+X9QA3E49acESVYAAR2+2umCSk0oCK31bqLN085tO
wapVAWNmIutxZeIuYwe9zMeR2TirJb/PZhPPW5dPGNs4aMfw0CKqMvLqTZX5nwCl
zSbsbzvh8P2B0oUAJxu631Xcim5smUw/rBTSMPQwxkdXZMoure+nBSz54QDNgrs9
HcClQG57XF+nRNvjWc+cWWYstQv/CtbJMbxeOOi9REaGE8pVWktQmS3ul2QrESv9
riSMwa0KBzA2unX0TmQeXIu8QT0EtQYFE6irWPRYJNG2O79zQ4Uf6HJzihIVfExj
7ovxWqhjp3P0goxqwjaw5ch7Hra8xmoglqzjCb24J07+mZPvUjQSKNai5cyzTa+R
6Ct3brcfPz0mIpQ8xtGtOatV+8Fuch2EhrtrYynXEf9kLnHfgH4qgQuRfCYY18fk
r7xH//DtWnzYHmCPsUylC+P3v2XvtogSe8nwjsNp4AJvCAESEWC2cAd6P16Knc/4
G22qQrZW+NAOycImU/w2a4pOts4XjJxwnrngVt+L5IwMXnsJ8mqTRdFLJ9EAkx3q
JY7F5zNQBJsXh27T7c6HKmAk9Bn1Q4gOBufJf/Id7sOF44JVtc3KRjmpMLMGnEGW
JLNOqArbvFNV/hWca/+xPEsvC/eqlObe7aNkYCBYyQymW66f8qtlgFQ2KetMrfhi
pVySTySrmP+NogOHn0csOqE86NFJjFnht8byWky2kog=
`protect END_PROTECTED
