`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNbd/+1wad6tONPfD8dZ5SXEV88MwP7QCZyVjWXuWj+BNKTunGuS0suC7VOD6zPz
59o9WCDLp03i66fz1TI9rFv0CKXgg9vlPTxeK8B51BvVHgPlKk7tVQe7A4/ZAM1o
eFsz7ZZBKIRN4nn5YAKr9bhN2nnzRZpYN4F2axaZR2rSaPbjuMKxroaHPtk7/KSy
CoyiRkbpCOLSB/vs3HbggN7Ms5pQ1Bjle1JEnn0PDYLRAAH9hxcXEyNCibwj61YZ
sLt9l7S/mZWfmO3K1jrQCtSISu62VMXcdhLb3hNr7P66QGby3uJtJFd6cGYfLLze
Pa+R/arKa2G9ZzMGRPZhpNcw5cBF8LkHXWlEAYQMO5hI5kTWLq2Q1qpnMmWziI8K
EIwxZdWiWT06fhj6EdqPBo9GNXX66uhSDqvznqzxZRp4N7ofsL1cabEiIiX9NRmV
Rr15UrnzvUFTRgH/bDoyyG7y4LtgoEtyafrGGnAqg/d8dfKXku+qcYbcv0SpHgUZ
94iW4wobNUdVo8TILO7z6Ty5Y7HXtlWgPH2oCDloLF+ZtulQXGeYL7J4j4UT8hvc
04JdC460OvSBOLV97/aolCxXIdqozsVBfz5QxyCCGF/VfUIEmbCpEQQeUjKEC/pw
cSYXb5ot/j+aicqamaJVftNtqHu7wW5aGEDwHhe9OIG6Xzr+5c3DhgTgQ4yYPZYf
yseB30Es3SPpz0eMITffulb9IEM/BMJpIW9KHtFdqYpFdCwTuSF5/+6bhyE9rdFE
CiZXPtI0BT4NZaiaXQC4TbPyAV986SFmZmDUP5euRgCxuupKn8WJFPZloTeTJtbt
WKtANLWK3OSfP76Zfj72KvMqd6MZXXDltLoQEd7MSCYIqANapkrJhx3Ye1wrvj7l
x4L4N9oVCmI9guXpNyPoFMjD0tS4n7UmTyVoZXsNHYDe41DxKuwx5RXcK5CUN6wO
X0DXorhdz2dWaa5Vnf/JhWvaUFvJ+AP+2G9WHbsrBkedCb+r/jfPBkWzEjvSGp3B
VshymC7Q8YnElNtbk35DBVoZIuWlSJ2Nb299PbWIK3MUveHxgUSs23TuR+FeSoEq
YjUIY7C/FdDgTegNXsmkWY2rY10cMPP/jYn4FK9imCcsHe2hczXOh4/k3okYxA7j
zj5tdqeg7u+Bu006X/F9j3mFcP47oZ09WSYUfasprrIs0/pRfR5IYSXyM4bwATgq
v2s0J4sMvnr/FsiAUuknwfV7Kq3SwJI2+93xUt8xm4FNZDWiOUcTIJIYOF/GHsYf
VU0U+QXz59CKRDEvDNgRyGr/rZQ445AZi80VG1hwJLq/ddzOrFpGdu8beMQSQ1Xt
P8ZWyzlKXLg+rolU8GpNJLkDU9mrQm28OXAlhnJxznSQZkJE1gS3U3jXZejS2zFv
susl1ak7zKjkEZ9l3s9Xk0xxyC2YFHAxgERG0udV7Vp+wOwWBTi9Wtp+H0qkJf2Q
rKk3t+co3UHC8EtSfGxZHWdf3Fvrbu+586UrAADLR1hXy/6Xcdwx4Ra1AP7yFhDP
RkQ+pjz4YJmm3TEhO5RzbSLhxNyAc7/ge99oqF6FboRW5RTLJRKl7ZX8k3PJmILC
`protect END_PROTECTED
