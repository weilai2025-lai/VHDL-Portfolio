`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NqP8JXnn1/HmBgSiyE6y+Ewf/vwmQ77bu4NamaPfWikkP8MKKseDAKmq4MjiZ+fb
1VkqaQ89XW5lhGUjiaCMXq6+cCmusPpxkq9VZfvkbN9RJlnlDuwp4w4CnIKdq0TN
FsZHHMQWXS64W6rg3gg+iK3gfk1jWIyuafXEk5johUmnzdj3VpezRYgae/auT8ED
wYtXi0DFmASg90NhoqSWWrQcZlFbHX73X87eLlryhGQrfnLbgXuAqR+jBuEwAhTv
aorypYq3qZh8lH3Xz4WzExehZ1PxmKpFGCgUOxU3FSApKaSLWz4qRUEUff6y4Hn6
IbqcjPIAP/iPmdeV7j2kQLpGW3K4nDr/f7C17vELUzpZTWxJF/17CyYlva3nlGPQ
z7AuiA6EcPkV6Nq22uQmNql/+E81PanVoafphXgab9W8QPtI/s/dgeIQgyJDxycB
gpHaS5+d8ISD8aTSU915x+D/mgJ+zugYAaom2nh59F+BrXz6vZu1EwCEHai22FLy
/OizY2eKXjn/QIQts1/4Qg34ZK4HORVGPZw+9/YC/9Vp45beD/D+xltv9xov8tUF
1MeZ1TOYpTJ8a+Zk2wdyywncULj7hnTnBDQiKeCZ4Fuy9yRFa9b5WooWYbq5h1kV
g8CWzyuKllV8bRa5lYxar3TgGbaRNWYVBiuFZNyljufHL9ZqWaRZXsnQ+nE17ju3
p3JGGUFcZXWddQvisS9/HOV6QAQmU661VlbhwlN2puOUk+TrTrA2gQF2CehsFCOS
RI7xBwf+Cn2go/FEBEXnqmNv3aSx/sQ0bdvYR5y+frM=
`protect END_PROTECTED
