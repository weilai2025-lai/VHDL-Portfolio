`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0ZFYoVAkCwumS3Ml8TP0n92VQaI6LI2LJOZ+r2oaLkxH1nxx9KybgY4/LFlhy9o
84JFiQJCJZfrDQNc1qMfpQ9k3UrZ0W3lDpA44DfNTtwUJtO5Z8iVD8AYNG4RGgWF
TXtkm5RC480E2kNm7e0Hi0319OrUw2XiagpuGtEkDaXg12FhRxhIAW42YjAOBnZh
CIjyTM1fkIBc4tpb2YrltOtpxCs8lBkA/Iw3G24LHf3Ss7SX3Q4bTwXhMpAjZta7
yv/cibRwzVDOprUCA7lq837Yiv05bZVUDVAh0SgGg7fT84QEX6xdDpUztGw1WJIb
QhCd3eAqeXEunq0DTpWctgSHknOYdfJ7g9PZSbf/DjOc101/m22BI3ScPKsFME4t
zkaoepWL9sXSjsBr4xVrBdbtoPZFn1+6evEzg/oSVlL9vkVz/AW1g157RUDS0gLF
LklRMFMae8iZvE0cA56pBn1NuAIekp1F38SJUEQG0jSoW29qiIg8DkZep+/8owgg
zZROybIBnqlXY9/OyxBphyxd9R5eS4LVnZgBlaRRyCgCXTOyKAbba/rUyJpRTvlT
tzmJGq+241++3uZTGXmnWqtEhth5WEsCdQP7ZKT3YL+9coeC+iuEoY3go7huhs7E
is0wrZc9Boz90iZlXCigXwOsUrKKr1lNvq2ZR7AM3edwVyDdhY+UuFJHdAWGO4+e
FCTfXPDdsE38s6lbHRm7dcCqKv0MCaWxuiwjJY6tWO0xQBqD8NHOYJ4mKlndHqQq
U6Fu6t4Wz8TErmk67xYCH99d+1oxWIQFqvMEKJXwtwdAvAFyQ3/zyP/tl2chiCpg
KwXpfw2NEQd0TZhC2JyzrAUX641cP+fgOzNEMkPffleaoTEw4vR1zngLjkUsJyJh
nlPMwcQ+5Nj0lZwa88PSSRCTw/qYc83vBT4TyTNxwkJh48xa6f+Gubvniuj2IATN
Zy1yfZcRlPZzpqth2rPOlsauYPQ9H9oSAwocVzoDghf3aVqbWiA+48IPzzX5v8HP
ieydheHWERXTpRq7K/gyLULSMvcOINOqzAM29JSe2Dc2A8uSD/U3MWupKu4HTXbJ
eVTp4M2ezfeuc+JoA4+YZEc67lSzkm5bX1hShiEpwws0GjH0T/7N3qGpc/b9WYPW
zQ5WsqaU/hYIgUjIbG2PU44TwpkvcLsJCnHPjJp5hxhIoDFBXcHmp0HY7/9JLuaP
7nR3Uswnb3hALPZELvUmXcVfwUO/XmhqgpyhWJ67cNY6e1Vt6Zkn5wvNiXKnfPlU
qOuFmohlfGhVS+reB2U1gFh7D1gEYnezmZydZcrlyHWeaTBo1WDckFRH4ZLDiHkA
QfgHiFAs8IlTHEmMVphFV4TnzrEON+Pj08IIpPcE7OkPl3sMyNXYAkHD+zWL2PkZ
ywhLfZ0vPAfkclsdx9cQW3NVXfqSbUHl1dPXgLTt9InSJSHOFAP37uBXbwfvhEB6
Kyw2GX/g8q8aPlPG/yhWV7EFOGllbjgPIEp8j8KjYjSpwmqFaXn0DJZasMQtYCTN
EXUr/IhPBHo//2QSSiG96PIVoLgPF/bpg65V+6Vu/GJvDEnQ4Y6raNm7UjFfBTbM
NSC6AhjL8JfHDgurkK4EIIvh5tjJBNf9zzZK5u7rB2zEZgumSWlePDuYK3St0BYU
p/On0Thzzpsx0SwIQmBWzfu9BJIHnPmoQxwKOeE6tv+A8WooquR0efdhSCNwQUkn
NcfwAia5orusCtC+/Ykeo5jDFcy5VDCkLgedMAjHVwma8ocHM3X7WhyQFozyy9M8
Yz8WOaVUPzIvTI0SoamL8HX1CefRQko8lihUMizPM9/KQjsAcm8B08Zy0fZSHkmG
wdrXknAz02dN0kA/vnaV2IsbRV5nHi5WXm92CdGoMX7f+P57x6qZ9/YKib2aZME+
AbxpifDwkwVP4hwoTWWegEGmG2b7wICi3Xn8obdoggodbmCUH1GquFL6c79xqOqc
2x1bUw2YSqfeXzo7dSrIZzZ10q2VHBPnw7y42OR51vr0kBUoHlbJHr4Vy/u/EPPb
F0DHGyibVrtqKvGkouTefoIHZhuUCCweOvfXl1TWj5gqgmRkTVNfsRkRvQGu2LlX
4PGkP1Hf4oQGoZcr/Wx68+ykaX0RMVQ5oVjaiGrNR/oZKfyPhx5im1tjKozm+7dg
hhAf2YuSGap8mgo68ZG7VTj8Ni8nj4U+Ih0U4RIa8MQ/j99m6WZNDEFNpPBQjeLu
iu8fkXQXV80O34nj/f+d5m6Mllj9tVuYDSQy8/UpnRSKK860wwpQrIddv5m7hAEt
YX/44LXXzKE7/M2jm+E8gpQgTTwxju6ubJSGKH0MLC7twA/Tz2ulVUWkrf98dg2J
EmXe2AursH2Ow2fdh3neVusQurGgVz1OxKqbvjPfMfwxwRhxV94z0iWLyErpxQOV
4zChZ2DOZCJvI0b1ic6PUH5PHxx0/Gcf/gDIpllu0VEck1OP5m0i610ClYII1m7b
c4M+ygxKoW+ZUwujqS/WBtx9XPEGglNHQrVu52ygyvsMq3HCfMmOLJldkWD/m1YV
WuPmuNkSON9dJ0mPGWYE2T7pKTHY3Dcn7o+fSLu8kZh78yLgpBxnyLtNXPaoiN/a
uLp09EzmEv/eLQW640679MabFOl0eDCg3t2Kvy7Dml3jHwAwF3eyiTwKNUymtxqr
aDRchG/UauIgMiDETYPwaOiD3YLDv6y8Bdn61nRFgrC7t5vRFwTZogfkO+fwrqPF
XS35/IOPHn2UDqrB8+D3h/hJihuyv3rDTNGTLYMiByaOVITFXXxr4nPvX8J5d2P4
hn/x5Wl5PM59NuG7viNQMkPvCZqBvPuTug9Ormle8h/mkUAD5EiJwPcDZpFrMV0A
oji762h8oj6GRbZ1kGQH63cXM8w0Crn0JIP3NxA/Vl8Amc9oFiiQsIUKIlPm3ZHW
xfbYYPYX470Uc7Dkbz2i/5zkeFuXEMLnpIRYKh7x/pkR6b3sYtzNrVFyEMNwPbPd
3vhAxRkaX2Irjiq14Z2pCFxbvvDbfn8uQ54wVVHQKhOnfcdb24+V8V7nI90ZO9V2
KeWgouZUWKTeNQq1X98HvO7bM7UqzXILu+r5tAeyRFCjVQGlbxBVxPKGp6jv3XlE
R4PuYHXn6ZmnEY2BFfgOKsvMGDS0C6PdRDwFjTrJoG9dFUVbwXqdNq61QwcmE4Jc
drV3/9wQ1mhRD3O+li0Fygrjuxa0P+owr5uPMg+eK2FLpFBLxteYj2nQF0q5W7sw
JQvYAvWqhU+dcV/yNlNjDjGJ5vE6kocYjNvfBzrrRYO8+f5a3wHFnxXax7z8nN7q
GDq1UZIhVRmhPSFhh+FirohxXR9fMPZZQ3zEznpK4TKkMNS2JMvslH1Y728m39f1
6qygzQv+ac2zEf4Oy1m28ve6k6rIt6p/xHSLJ1Ci9h4XdgXll03KnfvAiWLk7MHD
1z0vFuJs0A43aTEQMq+rDpvRx81ZYhse9mHnnld4mPxhVLi4Ho7x7/GgubagTsQ1
zOjxFR8WkUokZJ9W/I2iyUFlR/kbJ9ssJLwm87SznCbll+GY+1156yiEKu/F3PPu
n6HtMveHrDR4WuTebgEKoD1OCpbzT56rJi5bLAx2Z+BxBWTmSeXHe7OLW49AX3RU
5+UUwYjirqL1EjIsX/ic0kDITiIafXp7wRnfpvQswfwwWcKVuAcjsxWFu97M+BBE
B0aWwcXVixnkoLM2GovF6bu4+Gjtbk9Ih9+ok1vpydaNn7M+M6nMQgeUx7StE45O
lOqX/DZ8zMfDzm26u+3KOUyPR3HxKVidUGw4mOyFv1A4IEBhBhXFOkojvOY8yzgs
yv/rXwjB/hFdt5dT7yaFozIVsmMSAsAw16GfX9CM9+jnvjqnr+7g6WrK4wrLVaZ0
xrVdq2LxHwOHc7cp3LvDV4HdDAHFAlk4yF/6hLHhaayPIjr1Fsgz1NhXOpjwf0No
HWFbMUHGKIw23QU19sEgJcpuwg/mWo0VFa1Oplb2309oodaTvqgufFotlyAjHYmz
pL8CF1NDPMmoFyrOm08M6RWDSaWjfhwXn4NVGkFmrCYR05e+uk54GEJUT6MGsRUV
o/H/JKewYhMhF5bErpUD+0OT0qbvEtGuPioJBlwMs1Knkb0yLYO2He4O4O90z7bU
/GSbMlwpd9zL0ItojtSgZ3e4wt5SrkPAw0bvATVhN//lwXpvutjNJtwfjoqd85h0
1WYu5Ez4ChRf2WCfpKhkJqdEAGHKd0QaUErfXrvBeyHL1hYTdbgrohssqtafZiOC
px2Yzn28hUKFBEJMadBPOj9+exiWoavtobnojX8W115lubY5mqd/adHUALKiS1mx
xMQwS0nN5t4+KbNgYPCVIcjNE5JbvtEZ0XWJ9fLQ3f6J7b+VycBPicYIL6UzRIGE
YmmRJgl7KPnkSl3Z+XJVAVUSRRypRQq2iYzEhSTPr0Wo8d3mc3C8fNHACZPR+DGY
1CX8XS9FzBVREIQX2zioZkiDTGZSfgjv2RNCXvL/Q2esaN4V8aGqcCoPhYLUi6lQ
Xp8ewjIU3zcXFcgt7ULp5sG9KEJ+Y9X0Oe58U5XqZp+2zF110w/01ctyWt0r0TRR
NaK0c/44B6aGuBf4kOEkSQ==
`protect END_PROTECTED
