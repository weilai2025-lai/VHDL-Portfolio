`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2iqvyBEW0xV57GroahnchQGnWaVXpIjYI6nxH7Rq6wAHs98wEnJBA9NEbRIU09Gs
6llT7fvxYwdTzSHD6ZtMrPsgXo6jySuY0c+c/p2VIvn6tV3xqawPycLiDFHcLDom
E1oXwPMDiWTpur/k5Z/vHtd3weDw83ZTnmdRWg+i6fetg1Z8lYkb2+xnTyl90RZV
/+Cb3DBIu9/DH4eapQt7AhTuSQRjtq7U5JXYWeGGphlxLPOPKbO+X5Vat8bvbZ7u
gMc3bQB2yg8SCv0N5QiQd0JCAEKud9Cr6rV0yXCROlcPWge8KB2i9LSzCuL4pGnv
pAsJAtbXhei8LUKPz2QzPXRStI2JbMzKi+Gyhrc0KtyyrFOmAa95dr/TZa+PGtXu
22Ae+ePKtKxuHTKU8TL/NxQgC4sAGIP2PUKq6aTihC6lCYntaHFSy4ef/x9No2xE
n7RV1/kpTnWMf28W2z/SM9IU36sOi7+MJyKd1ajb/lUAD2qo7lh4TBUBp4vjZ9+p
ZTHqU9so+5+PXd+8ixGsMdSfEfEErlz7/aH7FrZ9TtvlwRDJWQI+jovxMW4TFy6o
iYayeuz0RpSQRfBxPBAsDYlIXHrgJihocY5gioYoTwKhXmi5zWaInU/u7tr9I1H5
CdD98bozPPW/auXBbvR89u4c8T0DRoON3aVnFEj4kxEYcxcWAUXoNuGxjP4z1EpJ
Bp+3wIsq4IGWSoXLZdrwDReWksAs6X9oKp21ngw/5IY=
`protect END_PROTECTED
