`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aj3GT1I5eUhr1qNnzI5O9N4OTf9xWgR+Odj8i676Anz0SODv723p44zZZ5sysMH+
I2M/zaXZiuOjvFFsDZyjvwG5zbzu83rK6dYmI8+Ck8Z8cqKLuQWO1T9ViA8F8VPx
g3ArHoCYALxEGXU8oGVbi6bXHvXVIaEuNHaYFYfDxnndYIJvrV5UVaEwa9Nv3dLP
2t4ctz0Scf61S89LaGEctcLjhuvhnK6KlfvorVYsBqrj97cQrVa8y6g7DEYHar3G
22YJu1iAWWKgvkmAdw5cLqkV4thOIP2xaK1DFsnn3MqDy2GdLzLyPasZbvp7CeYp
dhAYPmi3x28NhpHAbXpaA4BfLAmRzc3ua8DxGyNqS25KbMqfprlSNsiuFGFk5AeC
zNx++yP/h9a95uAqg9hAC5e6wD/b5PcvDknh/TNFKSEA1LQq6YfnYQ2ceCUgawGd
+f/yEQnTfYbtawmIDXonQpnzfz3KHh4OCu6OaGoimZTxAFaQnfoS98+dTCTLePiv
DAC10aXpB6xgiwp2zyHnP9EX7J9d4iBNSN4kdCr7pkgf5heXaxkO/qG+69S7RWE7
Et0aV20dqKrmKiMpEAdxlxilmzj/C8OybVRtAq8yjw963YT4eFg1zI3pQyaOKhQ6
aUTY26AbTuqFmXc1aptKq5JeQp38YWhPs/lYAEAtYfWE86zygxS0N5ytHu3aVsrf
VReg5wW6q3tmNUVfCRFljyXGEXNmksl9ptu20po0o4NJ1nQn9L1pBIaCAwgVp8N9
T5OXBRBxmKeN4aiKRa7K9N3CELYWio8Hov7YtGf0LcaXoJbwbJRt5aRTPMW03Wtp
8vxAP6L+1op5rRQEybhioDFN0aZyFHNqJAxan8dWko7gaixNGiZDr6YRXM0IJJYm
Ki+FDmdjUx9tiH4wE1AsswVtenOePmv8y2rCf/pwzYY7bLXeCJhe79OwOvEwBQxw
TtmbAESFJDzR160bs97/WpBBLRP7T9KOTMZ49SfO6+hr3thr+1CMoIx9oReghi1V
mhXQ2A9wN/mUF5LcgxeKelB2BL3DEZSApQfzDWR/YJB9EvOfCmWdi7AHaEhm5jzG
gj0+lJmQd3VIzfbwm4//XTjIdm20JwWGzWYlyPnIn31miiVCug7YmfUhPToOGP6S
KHHUWo4k4WTMy/9N7Cc9YCuQf+ruK2yae8u4M6sNTJ0FwhP6T/yXoBnMExL+J5DU
clYlRBqURSUqZLEw28adQvX83QqSFyzZe3wgoRqPiGAlMJUf7gqfPk5WUdUwKVkd
w03vnLQ5ViFjoZAzqE1QYGcsztNzlS/Ch7qmr/AtlW72BQOQBI89OjOFdPBelG1C
vrskeyd7qhIXHBPXkYI9OO9zHhaqMXEJrylABGRtDaO4e3eDxsi9gpPySv93CF1C
u8dB3DvBpyyXlSW2fWxzfxYIKy3Rz41DoyGSrKg2FZ4N39uH39jNxXmX65ZYiDcP
VSoDIyD7nmmU4Ql0z3jRsZjWq398JauVMVTQ8NFNGToDedFN0un6jduPfa28ETII
2XCLxgUcbC9Y1s85R494OIGfQdrUYDYlO125jbredY6pMBkhqa7+89Gd5XpeGpAC
iXi7IwVtB77rFYeQ+how92zGPBJ7zNQ/h85SMxWPwKZu90uifNm0Cn8+bhkB0GhQ
x6EYZI2xKRh4cuDfI4v/c/KPMrEUJvHxe+AJNKmw5Av9Pf2ilIUTg9JST4KI14Yq
dpxkT1PJaXkW+yGIbTjLiudHCOsUT2oKJawgBIoPuzQ=
`protect END_PROTECTED
