`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EOQrJ2bLIcwwOLlmukUAsagbCm64RDjvv/5dt4PIZDFni0zgCLaw38SB26Au77hm
0FB9VCI3q6PBgl4jyMc3ZAYjdFQRCUd46DAltH/kMzP1PohQj6UVtGCy3hm5w52C
rR418Vr5wxGEiVAKWTqaxGeuGQw0yGV3N2vPVNWt0UzBMXFSa0tPa6D8Slnhspub
PfFFXspj+Q37K2CKkjUKFccPZYh0ukyaR3K40JoomAoWKqYAy9OlD5ZF5K6fZPTZ
F7tE2TxtnvlToZYm6Xa2QPbyZkNOJtXGDU55wPYBxBgmGLFgX05kR65q9vZtSVed
PiqO8KZ4MNaVx+VMUUGo6sxa/bIWn3dNjGwwNCicIyToJwWJlnC4eEzBjyiFRD4G
Sx5e351IaTGAyfTS8LGvfXEU+7Y4areqeAPwpBKKWwqXc99M4a5vhiC6aUcvpTnT
/bHzB0DMwB4HWTpszOeM4dpz4VA9TD1/2rT/rCzdQ9ZA42kwwEgVq19CSkB8JC3Z
m1eAhxr+60P0NmHLWhGjxR4yb6Gr5f/kQYqxS6PINffxVHHMguKrJUhMh0MXF43E
E34moEbwIZYwuUYc45KjXg8q42ERBoSsIVHRR/0UhSg=
`protect END_PROTECTED
