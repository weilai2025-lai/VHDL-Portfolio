`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2fp7G8NCaVjBYK29FilrZelJms8pJJF9xHTldqXzuwHnCixZXsKwDXLwqWDRKWu
gCA7/x5sHoaUrSSen3vnIaAKsLhQ7U8gEbhuk7PeAxMAuFqDsH/UPrR+nL3mo+Gz
QMnSAXctwHlZJSBhfaG/nEUDBG82u8pRYPrBBNJ+T/HNMi9Lpe1BuDk4T9C2VC1q
Wcz1omjjEA1x0Twe+5GSzvSU7noAJbXCyfDsTANrK6pXOJ6bIGNmdxfpEXba40TV
LtQphgc4daKBQFpQyOOsGRA996njBpJM8CS+fxnTDhyutxY9DDuLO1Zp0f/Othwv
4Ar7Tu46P/TsXgDCIMcmjliMEebJ6ibYd6LHQEvs4aiTqfZ2s/4vJbEqizg9UN9J
pjaKSYEPok8XaunkAhEOgpdtgLXW1g6Am13ShacsKEPuyTSao5/bgSl15yQqllWt
LCKFRbrCF+2Oh/O0UV7f0h6ZRfpYFD47XgIMBlhgPRdc1Hpvh78VAQLg08bsRyod
JDSH6h1KsREZw6givndyJk80Z4l4iMWRjI7F8nwL/Cw4cufs8Jy7i7RlmzFF8f72
DtLFLrBoqtobeacZ9/KzlXIGyvRkDhWd0qOZdbuFdlfzvgAkW93PoCZI63dU1LZq
tO3bN8N5vsWDWgZB3Q1gQGDLr0AbWpEbvy2TxS4tV/MvkKwcX0r92EiY6fbNVv+S
6imLae8au1HkUvWxyVN1imb1zHqs5SooMNCnL0G2gJt7Rl1pPdZk/VFNhDaldmn6
etlSAehShQExBv/DdDOe5y8iTLXVZ16h2V6BXtsK/1KOr9yzTsyiQtejpyz+CLmn
vWli0H6sQ7D7UMwLWhQ4pZ1ScbilF6suYcBySPHkfR/4uV6es3YeXOFfPmeEixZP
2+bUI8pLgX+RcFBrr89yj0Dwzj0GsaNfpGWLe+5Nlx3euqtVbf9KOQNVlNuNNDl1
e2kl1B5+cS6QeNlLBsbT7t5H3PkvRXER2a32zLVR2zjlu8I+ECsuCYjl2awf0qTC
ISIMtqWaED5jBM72sdxx5LGtbIK4FFupH+r9Ay7RWX5fqeqyCcwX4LupkeOUBRPD
WxzdMKpul59SlCLledr5IjswOdtRQUzU3wt1pLPPgWZpem3Lqe1Vvu7nZbM5yPuY
eiELsycwzgkQ98WmFN0+3OIVCLLDIjIEJgBIj9udM/nSR6N7PGcPck+DoNyfYCAI
phnaxaRy0P4z2Xn/cYzkm7bkE9E3ubfeq+S7GNe/oakdmrVmxrTyfnwnbfIcCKs3
2OA3CxI3czgl8pqteTkdsruNV397qBtju7a9Zp57Lp81PnVI3m8bMuPlKFvpWp7X
32qrlKB/ymc8EsUDjFSIGRjgkGpmRp8WbBE0t4W2cKrs5ONIfLCCZl4k6zxoy5D5
kl5H0HUa5i7kGuYsfoDEomh03wzcsPnFxcuqNXQl5T3SVKmT7aA0Lsnf6oahRF01
ChTktYxMyJmDx88FBKxW5JeEsfbWw2kHtWRRyncncg0akPY+ldHR3vE8u0KJ25M3
yGQ8BRqfL0z/A4GKx9dqjDamy/Wb+TrmHr3QluJObmHVwduInbmqp/yuxeIrv0gK
t1J/+BnfTIIO8fpGXAsB3BtgbBRGH8Q73mjegswYlojY8FJKY82cDzLG8qviUcih
H6ICHVYFXSLnemDELGeR3MqKMYpw7us9SjQlOkZlZYqPQMUEdIaNaPaU2wGNU0pQ
oUmdm22iJIfVdli4HCXAzWZPTqufr2KJeSrMm0c3ef8JXHx2lb++zaDJJG+3aJPe
KTXKDWzoTmrVojiWskbnh7SDOYLlQMo1A2u94BozZMmVS5+izodTfdEtG5yg4U1+
ifqBWUJQVxUriPRuOqGubq+DlwzDhPa9M328B1rsVHlUoiJ6HguesdJ4qoy3HA7j
TDoPT7kN52ej+BexKj9ieglzU2MC8wq+v7QpoKu1V++vrYMWZ9HmEiIHmPUsvv41
D+ZWTGzqIPxN8h4qWgqA3LOyYfyqaMkyTJGuqg+WQrhAfYF501m5YYED7nHR8pQ2
8HmaSGmhQCCQz+YjNZFrTa53RjFH4bq+5KDTWz1yxGoCC+jy4pexpFWg/aVBw/jM
pFznZHYUspUEQHErFJcG4R5dLVQpdSyi6iwcT/NwmKN5DBbhfnALV3As1UDl5u+1
91K6TNJS9qNIRyDV7kNIEwkFkQnOL8FN+kweSXTFfYiZYRrtgl6UWueYCsRId2/c
un8uUBjUSDpRUyRij5p0qw1O0hUr7Rp3Q0Pz3nwuqSX2MLYd8a7m0nR3w3amFSds
Xhz8U/Hx7pqluXskjpzVob6v4Afbg6HTHvvz5x9tQ1kyPjzNuOg+MX8o/vBY5KQr
/mCzJ8uXrqKaJl/JjLTaxAgFk5f4dT3i7XmTGGlqIw+EuLWtQVe+t3loyh+ZebOg
11yAgzgDuyH/XGBi56NC5uOt6ejrilZw3d+gExAJNl8KF/5fuUXMZSv28AhVxbwp
Hd8T+hSFIppnzhObySgAi5B/07tanIN/gZrWHwPu9siUalT8WNeh+vWYLJzbH0Lz
Ia9YjvRcAdK3aDXE/RhTj4VD21mMZHPxW4RRi0/uCAwiXumzwLq/HW+K3ZnnvH8T
nv2Nl89yRLgzSXlKRj96ku+8UeX8xE7iQZ8MZCukBzMd6+fYRrsnB6fhlbuShkaN
bGQwFwCB5VJnqOQGoUcCZwHpRBqaEiwEKk/xQ3dWtmZbTDVQZY8Owsw85cZK/PMx
SS0FgMzCfKeVVHOPFH+3S2bU//mMI0BLZGNWyCm8Z5venpQ6HxpiWgaXZOtoNA3A
cul+QZV9Lsd6VVHilmdouVJjl3R0FBqiFASZ92xrzR7bjcSMYTkfdclQwOLn7pH0
wUtcy8CEbvox3G8aAdsx1wzgSYD4r5lMBdYEjbSerRdgqFV6dgfbKd1eL3ZDFxp8
ZP6WRm44G39GOd4zroy7r4cKmq2qxfOjuJPCFrkHrn8ad9ELNyJoiBSamWnN0oxH
wGLQ7NNMQ7D43+LeSdQ1oicBt0RmctnuWl2yr3GfqgCXPq4oDVOPsCZ6HQpjTs73
zgOhFjuSw1zc1g1SFRo7ieRjEt0zoTombc65YzqW7M7IdFbgTMDB+wwPVoha323c
IHE6kG7BZnloowpY1JK/CUxk7Dcz98m9XF2kGrgZHO0BERMQnYFZRrDV41cILLwl
E/3tsXau2wzPGsXxgLOs/ICEi6nOojOjA9Imixe2HNNm6n/QUA6lGCU3s6lxhqO8
gzS41uc9uYFnWyxY6Sk/oGsUVsKbXRDEYzf74w1I6yU/vL/j/8bKNEPh5QDQLnM/
yyRmZ9GYm0ED7hfAsUtG3nOJxgH0t4KCSyes95pdGnljR/30D06v8JxBAogslp+K
7HbIEJ6vk/sCmOLvBsyZ7Ue1M9F2YMnBuwuBeeDMSKN7YpJjzXgP5liJxcsjw30W
6HBdyC8rqj9pu2WueMt/JVxvUzHdkPPfV2FblQHUA3VWCFOmQs//odnYnh6xvoyo
xYGPwDbCN79wa+kRqZUu+PMIyd4qj3S/2tQ6d+cs9tpInWYlYNewc76wcu0GkBJk
PQtU+LidBZ/Sj2B9X+y3xgfxQJzfH6H48tU+SH1EpWiUFycmhpgfUcRf5KwMYPTM
IJOBrZ2uICIxYBsaWNPmelveLV2LXsO+aUtRb+o2enCLnnkW6u/SprfHFgxL0Qw7
d61WuBlYKlbqS3M5ztcRJyqRtx4JIFJWx56nyuSmqIRtEqfu8udWIvw8SlzLP0Dc
VLVs88VC/uPpmaxMBPSTCZ5Mc9d79IpT0yLZvIym6ee5AXIkM1BYf3SWTJdMr9AV
5yEk207OiU6UOPLEqZK3F/1Zw3XQSO32tQOilyVrRXrIhLV8adDhSrVRfx2TjPU5
pbC/cY1+CvdkO8BDKwdqNjWfPJUFDKqm9u8/S1L/P6NlTA8ltuEhV0H9yhXYkPAg
iVuvCqU1TqTy5CiVQObvHg41vfQc20kn4oHUnMGCgA+qH986XL8CxoWkSrFmf7AA
cf5lnom4mxPGIANFrtDGKcnlY39Pg9lREHmES1XfEqFRKOD+1HhMdysBhJXdcCjQ
mSf6iajlhvf1ZsPy65RRFJmLEfvxRXNrAHLdJfbe9UKvC9w1L5/BaQg6ffjerHWJ
ns2LoSfsVsEYu6gGN1bjjClox7hUHRH2rR005fruILty220H/O9nVx5lY3s0dncf
IY7eedyv7lGC+GF6qSCbH0IxzDktvDhA1uEL1eeJT5PWpZPLGulSKl0KbvefzF8j
xxK1Yk7WzExD/SANCPOP3H/U2DPEIXWI7n925qB9Nt2nVRlHVWf7nCBr7uXx5h6E
pXyFBjSl1Kttq6rQFipednmzvAXqFy+QtITO7+Q7vUdWGsW7cOQQrJ9g7mB8Az1B
e0hAmRTM7HBxz9z3roCIM1SRGjGWc7ZIoLKTWDJYayCwjSuz6vwNW4Hr9Wbz/6eQ
`protect END_PROTECTED
