`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wK8REnATevfgNe3hbK5N8QSdHVTEZqjIGKsTxjG/fI6L5uI6jkoCsbu5XSa8vlRY
zsY97AogUVS0Y1fftvKG4yJbM+viGenS1iKXm0Gxybe1Map1Ofst9fOlapeL0QVl
9U/H+ScHJCwGIiYweA4e508LnPheuiZh48O55HnZYD05MaiQQg/gnc1rcE8/6DSr
wqNVAF9Y3s+P/wCrfOydExmw9w6/XpEqmE847BlAjck5D0T7dnX3lH02x8q6TBD2
ILi345kAmAHfOqhTXLdwDhDTZvqXl1+//5skQMBhOwh7UbZO9Ww2TyivXKh4CJT0
h11GznGtu4C8IzXGwdHSKksO8JQf9GhWNF+Se6T9M/wfSMjajlAc2MBFJVdYmQiz
WvWQqWSZF50oXWN+stHulfV3ZNcD8x7B7dbIdYl1s1NTOnbySphEYU5bsdCLKWSP
noMwh/HAPgaxg0yu6+6akCtHW+PhLjpqEJE9mwuglRQbxGo/LbjbGk2AN8DVug3J
Iadb21Oc3kNpz07NfuJreDJN2LqSpp/bFDF6p1QdOOBcafJ7u8uIKW1HXaZLkItP
lXMvwJVaso7Emc+4LANHQMrYb1TDQgzBk6mg4H9sXhV8x940VgsCWTAZOKPld3eU
uwy+sFa8kluAi+sQ8gviTw==
`protect END_PROTECTED
