`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtjW1KW+ehlqqIDQ8wQtAerFpU49zHTOwv9/HA599S1+hPsiDgbNLoxnt0dahbuf
/819spnsCqPYiOpziiS2fSvee1cDYQ/a8Ig0QUoqGBYD3ckk3AyNwho26cVy2jVn
h66FN9VgtQKT+DZp72oCUBSeQ61UdBXa/0FGOTcw0CU7bvr74BAI41jppxb5NACl
kPxbJNbKLytZROekSg5cFmq8KtvefhFm85LxeMsyUDhe0OsdcxB/kHb+ILieNAGN
C4DDwlDNNX5Iw6hEDTVGq/ezJA3hXdG6X0YTbI0lnlnCYrjr53bb/KJdxsVFgbAw
ZJoHrG4Y5zEtxH8HMAa6yfbcAreinkOQH/LNsiZGJVMvu8Vy+3IRprwuDg8Rg7tv
c2iR8xoxOQTu/bkIaZ5Sg6D5aZNv3F84Ms2Or5qJ4XqD9+0E6A511m6bgh6D1006
Xm4DCcztx71di7lQT3B8Uar79p0M0rgaNH73Q3ysepf/cvZjk7KDD1YFSQflHbgx
y8aDXUXSr1QFft5Mvs8F7PNaYc2Cqjh2IFPr80UPnLdflMF4rsja8z+/cEqRi65C
EidVSJ1wjPR+UYBjTWMSTAosJ3ErxWI7UZeOFQNQjsm9FtU/A6yFgKqXxV8ynTZi
IN7xK29sY3clSDcGC/sVpimvkkyLbGP5auIHwAwTWr6GVtlousaqfg+R0Dtw3GYG
JJ1w5kpyvVKHFoliPeyCSt6fT9UlZdGyrb/GRgx/OMV0do5n/U3anmnJAhti+Eh5
N53GVJXBeLidG7Br7zO5JNIDcJxlvkAcF1t1X+tnopmwlGv2zV7BqJpt6KoSF+lV
urLbXaEQ1NZagKQbDMaJJWBet7huxevtHg6Ge8H3tUM0cnWVgF3NLQoObSOTBVbY
LaGJLePJsZ7GR2AVM7w1hMZJgRWF6OfViEQS7wffuEqAjSML0zU1f3ruDuzunIJB
/3311lhuch3zE5Fd6BKMSkQlICgWn1YYzWTB/7S4/yA80g+s0rN/t9v1RmMY5X57
BqMylAllzPvnX2PBiL7mBR2bpAFe5AInD+ZIjkzEtvZEDt4O7cR9AX8wbOeYv5Aj
SWPsEsmokn4MCrb1ds8YwTmFQemU9SJUZngPS53P21YdkDuyhglbby/1SLxAPU6A
Wy8buMUss6CzdF74CdtfqPlkVIohxmSB1ZmN+WvBATRnm6X1qfjRpdDflanbKY3H
s4+ui0IdENuPqg0vJ23oiSM2EsXCSiuRTqgfugKklM1jQPV2gR1ZCFpc2fhxJcCr
7NLGfPkeioTaKwyK73PJ98D+98o2qLoDoJtFRxf7F3XUhJyzyF0pitXlptSMOw1U
cmECHk5YZ+ci+0NDFGkQjYWh/V6pUFfJaZ0EbZzjmT2RfjkQv/MtniuqRfeoi2Au
nq+KpD8F44GwjAT70ZECLpqEtOCmxIvR/RV5qsJQH+3RxUbkU67tReX0hOm6wdKn
Tgk74xg4vd7Jsq0ka3sFAvQIMwiJTkwXy8Ks/zflSYRy1druM5prcdEus6Gt8anu
hU3zamz9Gs0DW5ir4uRdpleDa4l8qIWPDeW6y+Yueh8zeiO59+9hyAetPdti1Xdx
eAT/02Ubp+vsav4f83uEmY0rjoqu6XY9uZIpbjxuGHLmk9+MzAhrwATFxbsCA2KQ
c8Dn2aTIGGNErCzzchS4Wng6q58jH15tR3+kDE4MYjFmVPy0X6JTKi774Yi3G0qH
Zu4tRIccCXwhA2heRxnq7OtkrWrdLgyWxnfYM8xB9az4CpzknQ5fphp3tJk5NQuh
kz6T+YovNL9Q1w9ut73KfEQufZ0PNncZZS7jxJc8kFM8m5cJm+ZPGaPLv1dbpMQO
VRKjgmRIvKCR9nornLg0y8dVukhFF70R9Uce5dPz1cFhXL1/qf8pY67xpJdzVxsL
SiQPYj4KQs1n7PRPcj1PNozVlAdfRgxiktSMYg/p6aj3GMietZd7Y0heOxp0vC/b
8tvnpbs79sOUKvVke4nglMFok0P93MFk6zNxT8AK0I6PS2+9KvOGTzIo1BCq1wVy
Bjv1QS0HOoD2B9Hpr6lulbDsqwJ+rttfM2UHMs4+kj/phScdK+y9vP37Ee9MRiU5
iR/45mEtKNdPV0tp1L0O0YZYWLTEnJkNqCzF0Ve370coFLJYKQcjYupTNwtzEPeT
c3o69dNKIIc8qnWqkX4wmh5c08RiB+hN2cIpZCmaDZ7mHDVkUe9SsAwESsl0HLjV
6gjYgs61mzmEBoDD69fWWoo8Mn2FMPMsFryldTVzsy2/IjrEtNcFMfdsNZ+9+VEJ
bWhtHMo0tRuKyi9DZZXt/2AsG0BvguqyY7lzm9ZA7Yzq87mVaRr95jaL6l5FCwSg
paLaSTY2xsxpb8zZHgp41lwhNlA+/jWAPFnDo3QzSU9kgpfZHh88CgM9m+7/IGlH
lETL6ojQMoOaO3ALi7QCbPp7G6p1Uj4uAGetbJPfo5g2yfhXFluhK/heoJZ/NfvF
eOZKPs/lLJ2rjUP06WXUlmM9B7pxdLnaX8aNuGCm+hTgYEP//mhFgrsjqFAQispT
/XWA3O6zI+4EwSGvgxD+51OLx7AaEA8mg68BpCc1FxqMZ0IMTolRC00C+4LZ0zcx
D83qCBuyHNuGDZsvbw6hEwDC9KFpsDS3qp5Jff1AJ5F8wICDjrVlYvlFL23mq8t1
Uigy6sBKlI30NP4smyeNs7Jzr5WAaeVWcD3Kx+OR60siqWM01RxNvOcKgThNqB2R
KKDUiISIyjlgT24n37hBCbP8osGXD4jQ61sGUyX9VY1jfdX0OPwz7JbhtZLYZvUM
CpZAftLWwRkYkkKrcKdfwYNsOLXT2JjE6X9tyseTzntQrsjS8/pwLf3UTHGnpP15
PWUPzjjED57TejXZAaE5Y6sfVrlXX7+m8n3fWT3dWDhCmyKWzqXbR7k3w693kDrv
t8EUUwprGaX4qAsFJ/90YUVi2jQITFT1Y7A4R+j8bK1T86fEZfQ3skHEqowJS15j
u2GUolUncgSVx063YfTuOhsCajdeXZQ+nA8j+l/LTRX7zYmaqfmK0HSRXXytRDGl
XbywZhzwAtUle7gM5noH3yta1p6d+nLlnOfJnTkgM3T5mY827BQLJKZZmRt3hmid
PzD7YqTZ9MSfyEEWpITZVIFd3oGbeG9tub9Oi9lss/sqjScfGBDBrLnIO4y5lf6g
kVDlaC1Z5xkK3Sb88hKRinrzoRkdizKPis8WpDqS5BIWUcplgcZ3MH+AGmoEkPyl
V8rwahHZu4HvXATaolSW6GmBhM6c9jmLFaT376D4gOxETZ81ikW6JPrUk76AHHw/
a3pkk8XHMQgYm4KXGvc2Pc9vTM9CC2XBuCko3dfE5iLe0B+47wWoDe2rWe51GaEE
b5/JsWetKF+cQomAk1oStC0mAsDyrIQCOtXnSO7RW7pteQNfmqKaiWDWToFvb8va
YN1YY1EvVpfMmtuO2OEfoue/bWqsw/F1oyaynw/y5WF8Lfar4Kt0NhgBwNQKyFTX
ncf28sJdP0DMRJJtonu/n/f/n+q0UfnJ9BGvXGaWg1iGFaKGSs1ZvP1OKA39Ao38
+F+kI78U00BwLgeeQ9D2WFr/fBOKZO92ZTtbnDJxOMxuKuhJPE81h1zfP+WxAk8K
lit38GGHNqKYro6Xh4EdO5UJK+7TvSRqa37gRj8xWT1cb6SBohuOdlRhW6LJsmh7
di9buDKbVdpgwUf97Egjw/hbxC+a3jzNQ7AGR56NXZ+rcEvmXyyNc+lKwdPGpydi
OnZDLK4TidsRuIguXwQchO/YLL8rmwLlOlmn7bfnJtFWY32hzUPtNwRnUsBJq7wl
7iOMVQe3giXudq2oNqVkUDxrxNRGFCZgeYeh0alJiXPO0g8xzxLHbqDfZcepNWMB
Bo8gsfrxVlo9kDy11XCN0rdRyalB63JdgxyrgyTgVIWXlsDJAakZX89lpAS/GXmr
BSGskZ6igZslzZUd4UxEldGefae6HW6IpbRN6MmjwgsLo8S5wxObt8WlWinVyk1N
8n2fHxavJiCc7ynsfaHQaF1xtg8pgl17V0iypweH7x8BgIGdlf7iSEOJpJnvFYoR
a1u17gAY1PuSvxXBZx+ZnVDYyL4M8kDr1DAPGadBFJ1khvGEzCjM0oBoBW+jDrZy
xDqYKV3V5qn/BxGR2zwO4jkeTvyQdCz723+CN+0oWnAF458EarO2rrJgffljXRVE
XsVEXAqgvUMQeEUwHNlbvo3Vd8cH6aklmzY2l1t8uD6Da8zc1hiPKBaQPu5ZboAX
/nwZKSSVLKnhISi1HEI/j6+9EP4Ph2UQ8Z44fuDCHFiEog7LzrGjxF0hCqgPmmQX
NT6qKfX8OQiwKVcly3+gNdihnqLdr0sJ/eya5xIV9lOQHUvrWQRaOQ/4R2th8Rcs
JU41IvIi5D5Anme6q+AR5dNfy+O4jdiB6N48NoJhuXHiaYj9luWPTxUA6AabJOev
kgXgOxY/69xhPsuNJHDhKD6RDRuFns+YiWosDmCHyJDrA62LBjNnaF26Iz2sjx5Y
5WRvCFDCMn1PX7clRX49f9WbF15XbFm+kl9FL0YMYfQUk+UiSc2+6fimPr+IqtdT
z+af+0RTuDMkjuYJi50yeAFZhQis8FGROV0Mm1ycHul5v6ooq2DRFklf3COANY6j
+FLrWH29aTt9dgiQpX6JB0b9o6Od7vWU7EPrsKtPEw46SLcQHfKvUw3CHDoQ/0Bm
AvbQ4xKlupqUrf7Q52g64BZ9kMw/HnPB7Nu7aVGkv3b+wYd+99jq/+Leg+IcAmpS
briQVkMzgN5Pi7RV0g+jbkMeJBNAOqUmTunr+TDhqfYNMbeVaptd39aOEc3yXP+o
WqhXKJgxMbPnPXyVmRK0u4cbukD7jcRblO/19IYrTtPuUsfOl+I7j91yTyf8FCt3
IsQ5/vhM2E5Uiebqpq7JlPBsJtHHmOpimtEZW9kLNHGqgc7ya8/L2Ub5vi1FAIIq
`protect END_PROTECTED
