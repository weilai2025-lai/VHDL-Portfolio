`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzaD+uVpgFRzQWdoGdFQDHiNZz9v45LBYzflOnFjB2qlEP0UvES5V75Hdr1y5Mqf
WcjfTtFSGkizXgoD0pCj0JNPM6AMInTwkwcKTqZJBaqgrklFRax8KHxJVzOaqNOC
slKHkmbctjHlALZA6Vnd3d4wkXjMPN9l7lhRmiU7sUClNV4GRlvAsXD8cM3lSJGR
szGSFFJ7DepJxTUy5DbznoR8JZQ/Q7Y0IFSsRmrudCMGERvZrzbwhPqpsYEdgAvY
5J4Z8Stpc6qn26yPjcDrjc9IL1ScLPes/6z8wZVg7biUHhZ53WvFSWT0ZDCoLwVu
Hfrgq7uxN78is576sroyNW47CVUrsMZeWxEOU3+v3U5h/D0v2NwDU454AHMEUNoq
Qa+aBoLvVxNuIwHvEXe9+qlNUR6smKMC4qH6WPjUBMO+IDFloDDqXxWHwbmDMuzn
`protect END_PROTECTED
