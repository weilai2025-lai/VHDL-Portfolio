`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
huM2N5MiMl4cSrv/OmJSPWbTSJsxRwpMlM/zQMllsxeoFuG5sE72HeL9O7VM5CPO
UpmueUWkHAB0DCJ0GJCLwvD3OsqQ6FaHwKSW7ypJ4vMHMPhuRel9P7BddnWQ63OG
2mwsizhmEVviyTfrz97rcfCdP6MpLjNbBN4McTLXYyThQmpweQk7ZgpfzYbu8qm0
/ddl76MCLAQw/jpAwB8FliK7E2LnZa9WSE7sC0lZm3wU9Snd7FKARmRCzEcXwrNR
nVTdAZsc/eTW7kwaAMP87ioXUbLx7Rlvk/P2tOkld+6T4P5VXv8ETc0L+V9GHsjR
niVhLEjEvU81kJmr8JWGkCS3vSRf0j8uP11bpyEN4k5Q97/H2v3H2jU+n7Pzwae9
2gG++rN5wI2qZkq1SPEoUNESQIOOHOUL8izmOW+NFaTS+/Ws1lU963K4OLooKRqe
k7r9Kfttl0KGHWmIyrxk7kYHlPfG3Y6HL1UHbvhHs+9eN0Cx/Q517t2NKKU17SET
m5XSVjblNL2pXqSwV2D42gvMkqrOkZwdaM4Nv5ER+bVPdaPzVu+JY9dihP4Jv/3q
nn80fOSpItbL5wr0adYsj8W4EL6ciRnHeh/Xgmtr+xzX47lmMbhFqbEqzRf9NMec
MJw5M+zcLKzFeoqt6FfGybgep+1BJYfS+i/Xc+mXEtfhy7o2DVtWdYrm4tkBO4Xt
gpcPf8MLFLXyNK1vZdiQM1LbgG/0yG1ScAMoPD3gCjhJKNkYfrqGxra4q0rOPER7
rsv/RN6rFeLYUXNWTvKi9PwA/cWeHXwCl4SQsWboaxI1ystobMpTNLC1H3Fovj0r
`protect END_PROTECTED
