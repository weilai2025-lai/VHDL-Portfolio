`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8lhARAXiAZTD1YwqpMpIPLtxMlYuV+Y3ftlEmI4tWwLaSD5dLni+5k9jVdlfZwA
yjP+huQx5xHAIm8hYGIf0Ffr9egcKE0e0yPS3SKIDU7o0W7sIYvnarQzKQRUm30E
ENJdust8WSQY/bxQOUlUL80mfsDefWXThVkybMeXDna5ox/HEitsViRs+/S8w1k9
mIb8wS+CbovSKIUNynNjzetQtJBTvY3D7/VaX2Ognup9OX1HnJ+AHVS5iieuPxHj
mtoGXkxdxHbSuFvcw3Se2UBHlvO78zP8cv8KelXLhv+bPl8DV8+lFb4EyVFac46k
NG1GUTHk4Ojm7bAvD4T+08MN9O+fOvGaZyDIusYnRH+7zHqeh/Ur7GCPHmuQryFS
5SOqyLnX9yk8Zpu+inY+vAviCI9y7Rzc2dBmXmw+PTE7J38bnAcOkolB//N1DcLb
bblMxXLSHMLpFl3oXKVs9/zctYgNtb7rj2Zj2P6LHw3FfvdmG2Dh9gbKapa+WSHH
A3U5ia8EnRNwbrh7faLGS/oYffn9zK8XuKmwfKDRBPWzn/UKtkzRIWTdn/PHpZEa
+PbVkrIONTbYO9xX5wVrbPICli0Gaf4Oe+Ya7ee/yX7y+8x62qUEk7HP2vEEqU8G
C86q4qLB1jSLsV94lWUxIHVtHC/Jd2LjaPYi37xvgsPkZ9t1DHPzFJqHW+kOXhvk
GiuoDx1AlUSEfzLhxl35jFEjBHrY5l9EVNHO3wAaJ6bnaC3Zr0mxx4JQPblvm++q
O9Vqv9+ZYZjf4rBaT2PCNVdrYLcsgB2e6PD7jBgPIlKCqD7FKojdYskOIjwLVJs6
xfMjjdOQgatv1ok29KPRfPei5qQzjQ/GafUsuNgpK/Xkfii1OGt6KPx29aLATugH
bK58Cv20S3IrZi/waipoQhbBbDWH7yjqMD8fhVfWScw6ekde5UhBvV2UJu+B1MI+
4IPJm+WO1hKaaio1gcCisyCKolsYZesM1VpSADCbwwMYpPrYUH093DagKyMmq71R
RRBa2lr1GO8yvpXt+2gGE/9i2RvXsyWHSnVvqgAtTkjgHsfa6ZGbWcRovSargLqa
bXZJFT4VlB3ZBmHPN+yn/ig5kxxpAZHz++nVkdFrNg9S5aWcYSK+HwXE6XVl3my3
8gsLFlJZv+ksPmJv+LLbOOksbu6dk9z7kQupomJz1BRdK5uxIhX1Be+dBHfUoTG/
aohxqlfNh4tndxcSeopUZCMS9fIOqs74JP93a3XTYWpF+/gHJdqKnq90zRDD0vNu
`protect END_PROTECTED
