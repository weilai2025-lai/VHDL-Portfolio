`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K4B0dmcd1uv44zGLpvqPx80gGVB8ItEXQbZopX6/ynJtRQGJGdQPSO9feq9SMpMd
Yg/DCapaRr00iOLLXbmk1UAlOmAKnTz6S83faYCKN/JEzy2YM8VgfCrNCgZM2zCR
2qhuIED0mVGEQgj5sfz/XkN1v78JMxOPfFi5cvD+ShApofm72DFYMEi91j2o1SBc
wlcCe3bH+nQfpMIQTYxN866YUcff1WXbUjpRZ1nnup02rykddzO7vp39Xgh4dtp7
8Qnh9i+jM1lnKEVyW+ue11VW9gJJe6BSMYUZjZojTGT92NS76sSzQFe1RW1lb6Ck
VrAc0rjW/j3AtlA9P+EMDeBpjqi8i48gAZxKzAdbxvxYJeOVWJecOwzmG3a+JQ3n
CKP9Hi8L0pdoVCT+JnrqJhuYdncOZBukminrtRIeY8Jm4eXEZkNCb4obh3UG9kLY
UCOVjvzyqc2bX+27J0mAiMAlTgolaHzmmhTVnd+PEprSWvnu4ZJ062ij6qDl83U5
zuL43t2uDDqKeXUYZogWgn+RoyCNeanKe/ieUUM4weoMFh6O8AVMEbkYqbandkWm
+Hs5QVBSK6e2G22N+/VEdWZLjdLu09N/9ddUi5fbKEoimbph9w9O+gUN4n29+AA/
+VoR06M1I/vI4BsgY9MvtPxNOW+iI3590SSfzV7cyc8bnpx69Vh8euCwTQTmOHl5
WRUrH7s6zd5NUfbIzMtCPEWdw+9wc3U4j7fr917iXIZt6H0cnoRD97bD3IV2nfpo
ZoR4WCllKK6XRBLlW0cRtXmTptdg5yA7BLE4Rg2IAENtV3shJooRPMh7mV2Z9g4u
RcdZgtfrdhu9g8dG5hkuTVrN7/b35Quu15RLgI9hwCFhPOli4ZnIFu4cgG7LSm9j
dY0F1/51iNa/TvR6l6LNam2RDNTVj780ymoFhaqFsFQFFc5Blz3GyVWhP75xPFkr
nDYxMNA/9MjLkScYpdCtH5NfkIo7YGV8WsTxvjFPVPFAUv2hgfiJa7HWt1qcbA+B
KM8TX+V5qtgOIhMieTZjUzspTKq7Xwa7bwxBz8XhuykvtfLc946zDQfT5ZH1znE9
6jmWvpZPdAY582GaMVQI02PjNgV6uZtzd+bjePnO0r34NdOmiOE5AsH9jjLjrKb2
lhqoRo/P5gs/hiyu/3w63lhzUIf/iyN+Pa5bWUxhDkD1/SU5h94b8CqUwg9coDIM
T100iYZyG/QnIRIx6P+kgyUdoO4CGW4t53O5nQp8TzIOFLJdvhcDklO/DE7d8P69
Ahs+L+dmiPf2jBRr2vlNAJQqsoefvK9/zsWX1EaXcJG8GWY5xQXzXkMk3P42W/th
oWGy+jYaxcAo6H+Q83Wl6U8ZOUTCbqpy1CXtcLX/Idgou+5lLH67Yewm0QD3VT4F
8I90YuTxeOn0bKaYBUqwObDYE157XCNXTivvwyxBz5R4wnsH+B0LMQp6DLqiHyhi
XP+cE67deEcLoAi50kXiwbfUoKV9Amv7B7f3UGfKEWLknVWplZzdR7ftMZE6qjoR
vllhQ9N6O68Sn2pQuFjz/QdUEfQRbvwgxteQt6BiWv3UWs8Vtmg4JbqTk14lwmKB
0i5Wucj3YJJU0E7ljvjCVIS8i/2yytjIsB1HhBfhN5SDCoKuvSU8yISzgonMfN6I
DgTRhnVyUw8EMY1nY/cavH0OjH+Lomh2X6Ns9DFTtXHlxVInIbjW9wphUwxM7saj
K1sWaG/5zOBWZD136QHfuTFpKe69KdrIltfyaBZCK84bAkS09eTcTY4D2qyjx1ka
AmJhOzHlbVXP3AkPDNkufaf4EHTYxmeXMeiSlFtvEIbWSqsIgSP+lZ+Jrwe6DM6F
PBOn0/2ZvM6KB+nAEMLrcVsML/mEkUo7A4QJB6PeqfghTPaqcks9CWyCzIUPdktT
OLQhKiapPc1TENoAIRDI+5/Si0WGfqN4Gu0pHECQGbviIsJtsw5VO93Np6TvuXWV
q1wh1Di1X4UYEfWNlTDwA7GIlP8YNSzu8DwOjb1hy1G0UdFL6pFBAncqDEuoTJlC
nvC/DMYy3g4hTmFUmE7UWmI5HvcfeprUa+xXYdasTtVvYtVEgnNbKAjciOmufpsy
16To2wzLVL6xYWF1E4cUbTS1GfMn7XOpsiV1Tjwpbwd+gydibToGOInr6+ZEjVc+
s1l/2/PbYfk84sCc5mGH3hJioAQa7kGgLbSOFBPxe384bvxS0Jk+/EvjEoUpqYwq
R7zoaVKp/axnInsAFwNaYVWK4TwoCsHwg5OwLX/C1VMv1fNkrIfojiNQZ47NcvVW
k9o1p2WNdE18KqPMzbF9Y4Y1McHjdcwv8dDuBefAEUKjgzhnSPSjqvz58FoXjgdk
i6K0pXM3i/UDHzBekS0J6y4wT9co95W/10yxcq6vpHcU9kjwFtHtAKTCz9LvQUDD
90ZAn1ShLZavslmhTFQXix4yZzWegkACoZRZrMcGOWacKgGZx6bcudXj0mhQpKTc
BehPmj3Ts/105yEUMZvxV99LJEdMl21zkzjs0xgqfX1dBVMhIRue/qT2IZcfQwZx
y/c3/mPOSmRBW6oBWuopuCfWSNE8ubkmnpJbrmJtyLQNm69NL4NvtyYrdmcFBCVJ
c1FYuxBG1ZqZWiTj0AKtaj1RjckDPuQOCdKO54SFytFtLKTr4XqhHv/iy1ikMd/G
PGx9N4R554NWYwHFdc7Vz4jvRFLYST6aLiJzoYrWTihtUa/cdCwIQA1KjUqDdqEW
gM6uf9UbswcgFg7lV6rZ+xNOs6rG1uhMZD2PxrPrJDFpOGlUucMEI+w4LghsCo+O
rdIYw+lHDNFYVIS2M2Lv0oL3ooAtp/6aChTzsa4KxAo6IJsUICn6FUV9g59gWv+G
XqAN6ibM6tIO5dECbOCm0m00rZIa22Yo6rgPpzm5ogSWYhmYUcALx9Ei/wFpoFGG
+2Jvwlb/oRIVNYTEKyLzdjmR9LYJfUny+KJIIUlIlICRTW/Sdg9OCjUy/oIDPVSB
kUPMIhcd0XIPVqLimiNIt6bmdXiM47OVINWoo3+57ZGu8X4beYL6VTYnN/DqH+a5
/V2uK6VN49VxYbkfkU3YPSV+mYJR1TrSoj6fon1fFQGFwgVRNFuV2K03Gtyiy/h/
Dlkz9xSs5KoP6mYZNNVkqVDunHnKtsnwvKuM1h2U8T0eqkU1/1XXUcOPlTCaa67G
cpMadmznL3RZkAoPPqxNtKbBwIEB/iLEjy4rDprMZItT460XT6IPiZPcCPQp0YBP
X4yGQ2Jjm0HGKEXVTmTUg2CMWVqhyWZfwLCP2Kgy4WTm9Dw44tDOoC3VbC6QW5Da
FmSqG01NR7MGMQkx+bQE2UIUTTC9nN1ox7bX2jf3EaFudl1lusTAXrXQzzeEge3F
n+qJ8e+NOxIJlVAqACeV7mQMzkRG0plejGTYVqI12o4/wehssxCmNAnNETRitVP9
vn0PLodbCFfW6b+nRFRAr0lNPGiW7RS6DxzeBvtsQie2EsowvA3eU4ryJLJl0TJE
R/5twoPznynqJagohsIk1L+VJlz/jlwSjDCCmf1fJw1c2mv4mBDndnhQVkIVLPKY
A++AeuYT3HzLNTHZtOg/dFxzirgh44aMvatgq0DGU39jAxUEhaEHbNA8Ow7pxtX9
A5WPGDXLCJA+dDWM6dk4XkZyJE1XULW4Lu1ravwthHDr0vO0FOL1Z+823RUOXC2h
qEqcjUdYBMLzRw3fwjHapGSFsSbGvLEdqRhk5Rr4GJ/QMa2ROAHd99t+ZXboe5rA
rp0pzLzqoN29C9adfS5r9hpbmB66HXmlk6QFicnRU7LTyTt9DCgUY9rdK2Vv3s3N
JzFkHeSR+nCifWIa+w/cPMnF5iv0RlOFIAWYLu4fSiFI9JbbHS4dGQdRSt9Kfkdg
1nguiN32WZIr5gAp4W29qVojiuTuql89zMVIyXIdMg4UhDy2KsT2gjikCtu76fre
Rt+vBGR6VvCZKKhTlVUX89aZmmEcT3spbyI90G+lkZZ47TOHz595ksw2VKLejcmi
Nfe5bNAnTB5YqGPQPQn0f0VHr9yapr0fTWTKO4HkuuifBrbhMsx6zAJlwJDGdD2i
90TC2h/2IJNFm/Mpy4eLKXV0Kc2QLLD4Xm3xHPVKXxQev6YPIPIfi+MaMKRkAD5o
Q8YvST1/5lVnuZWfcmprX31uttAv9cZpuvKuZhrY5pF63YR7CkTrKBBIom9+l03s
b81skgoN95x+ylOweWpl4pR1UdOAAx02Y2uLa2ZES84NN+KnBnUFKAd9uNLqfyhR
KsN85iTKS6Zjrk806AEDXBx0Rggzyvr6I9IRwU8hAjh7Y4Ozgi06+8MhSFjSFhjj
YcacgA3Y8RXdn5DrWAWpDVeZFEyBEXh1GmCKQQ+ACGH7ZjhkjzsvoRsYh4XrRngv
naJ2kl5KCwYuP6RYfCT9ka5qU9AqbKSD69r3JfSyzOsvahVcTIaV7QfPa37B83Kh
hKSndUa0BSLUa3+BK1oxpLL64hffvsWE89gLSC6lMbECG0ZE6Y9SuNDuXwez8kHs
jvR/vDKt6NPWnsIxkDQ3bZcF3U/XSFRGmnxSVJ0yiIZlQSbTBvKkE3I1Zibc7/q2
tZUDAjQoLcfqP1L2EgY2l+hZlSpqbHiPJntDwbUvK3C+lPG6freqOre3n529+/6v
dJugz5q0zKvHtE7uEOxLFjMmRFeWrYp9MV2VfnmJCe4=
`protect END_PROTECTED
