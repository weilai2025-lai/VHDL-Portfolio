`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/VzVX2qiGv4Gvm8ILShMW5G/bM27U1ppy5EyxvqvLWyQyHo+hVpDqxXr0WdiJO7
ikot/d/ults8+Skl8fg7tDLnFE7wG5vy3jRko7T2lh6OB7Rou3+U7bMDixTvpUqC
f8nkfRX1ux08Jrewcl+fkyBia0Fw76xyW/LZRw7a5+8/CFGN0xpK9wdUMsrqsFuF
Xk42mBNWg7MkLLf6kMJ/e9k4+28778KYTRXaGF/YO6fxe2kycqAEdER2bqvfdgwF
H8TIphFc1fdKlCyQ4VFijRkfkSX4jArx91Ju1JYak+U4KnH+xgdFa76FYspROUrh
wXPd0kPc1QJwIksFsYM8tWliKJpXfF5UIjfgFoaBEk0nyYFgh+PsNAKFdboaqBSC
AUDt2aOh8r7UtVsvFjcROvzq6xMv3n6hRAmAWdPl/hnzo4DAvJ4F3wjLnGwc8/Q/
JKQ4lbY8lf0St2H/FB31OENidi3AxWuI7ME3AgTbhbN9HvadLM2Z76jPzsNq6/ps
9Xq0wUO6MUiqDOz4lhKkh/UA/Lj4sbkpIA+/HjzgQAgiFwRmI1CewZ9ZBo5+RT9+
xp57ZqOBvi5NjxDJLoKjJEB4rn0uN5q3Qt3WFp87MQWoZhsgEhdxRY5MMB+M2JYY
0dO1nl6kHkSy115QqopaFrcNp6poY1utiJWDR3c1Yghh57J0z0oWDDZHQ0DSXcTV
1UvvzFv1PF28j3/K/pdmcuE4assodTAK4VUbAe+GtuRazK1cueEdgxG0by+4P5vX
9+pz2pEpbXr4gPxLbF2Y0NOx1tYaY9fVlk+ANimj+h4AbbsWsZTPsqbbKLB0ty0c
AOzVxkUE3rni3FZZbA4BPceChkJLddLEssqX6C6xk1X//uFRIh+puHYOZ+Lnu7t5
1HE6bq1hHwy3EHeBwB2wqNG9rYqEU2LkjF6TizgOrBvDw0dtKAK3F9Kx4/WSUJJy
fDlY3+m7QttRVM1PLJNlMr1xo/oME1ks2521XYc7a2wrvgbxRPNbrHqfKw5SOAHt
K0debkAIKwkeYFGjb97ZZwtB6clFyZmRoqIz62otR9cN0YWjODcHIHIfo6jbiJLw
a5q0zVappp0hmpCZVQkfnOQsPLVjP723hmabcHmydTFJ78SRW21/nqN8pBO/zx8M
RWLpUCYrFmWRVPp4GKXhl03w1WVD/BsDR3E8Ejt0VGDyNaW/xqBAZKR4rZ5ktlbg
88j/B9SLXY6KuWF1ZNrACTpiigEvU18xP3ChrqqoXNkBps6HJvAXIsm/bTeGa3Dr
VFbMmHstt0PWWp+D1zhizc0V/gSKTVJ+7fXKkXpHft+vLz0HYirh/WyVGr6N9UKC
yNTKWXWsYBednGLHHrN1Yn+ExpjJpQaOqfrygIK/JX8xGdHPoc1hGbnVSsm7Ofct
/e03SubmKaHDtsGUq7sZb4n9glabbQGrbptBPyO7hRjeTqWqD5oEK1O0lev+2Ws3
497pEN6ORxbOar028g91YnlpRJAeihD/aNLR+HSC2CQ8rsiYsw3mgyARFz5fhfWH
7LWUvV1XJU/agfWUZ1ZK11z8CMcowmfW3bPUbNRgy0+fNni9q+fI4m9BR+rM6D5r
xBo8EYaknw27oaNy4hgHIjDdaKmWzMS+HsblCRm1xxiyayq4xwUQZYU1mF3HlFDv
321PRRo++ZEu/mP5aQ5RyWUuZL+WK9b1MpAERb2VmKMMFtCcxKAPZi7FFEY0a8mz
vxQ7ZoTmpcHVZvLW7LUCEJSwsugCkOVnPWvP7n0CDUA=
`protect END_PROTECTED
