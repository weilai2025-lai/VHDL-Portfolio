`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWFu9SR5qsHw+s+6C9GVuiARyV6ZMgV1umhQ/8YnkG8pcRYsdn5l2YPZG/lOLeby
IxX2Loqp4EDuSRMrW1jWHJSPuw8K0KPdSFDQqtyWOGJjhOEuglsp9pNmxq4owWM8
oG+3YV4u9FW25sBCoFA1QhBzQsVA0asRgE6bLXBp2sHy8KT9GR0sWYzkMiXUV8L+
qX843SKWw2/8fKCepRbAs+P9jDjUXwft9Ps2vKsFQCStdew6XGH40wzZUc+JpIO6
FHOETSZkrEsVKL8pLRvURXKwxqNTQy6G8At+8LNTwk7JYG0vaROmFfldcPqDVOnf
Pz8GdveDnaK1PdcoEDTXMeLUqv2V1YBEa0P2Zlcgk27Y/wJWH2p7DXSgS3QiILMr
yRuxDRWiXapsxx9kxxFnuwTzLjDHWJUmI/iiDg2RyKYptFGZ2OHGUpulZYjf9Ak3
ngGbjDGpUDt5nG3BB1d9ChvgP0c0aX41uhmoPlbDjzPb0xxYh3p9SRtITjrCok84
n5icIIMSVK2i1vphqnOQVTeKjLr+NB5mWziMgKGyr9ubEJZHX07z6KCu0skf3lbV
ugK0nt7vCR7kAVVsVteqzsLCyYjbHLdR2utC4uwhCnViq/8TEUhNKth7znMF2alo
JQfVUZygh7wf6LyRoBKMsMUG6n9GMXUY4hnvZCSIQS9vkz863uK6/U1Vk5NaMIQk
`protect END_PROTECTED
