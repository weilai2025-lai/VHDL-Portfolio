`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97z50P+wq1jOPgyBX9H4flv484bpUMp8QmzIq0rau8RGn/7v6BAv6dxj9WhZF03M
8cFwvObcBMz5Dy7r0nOJanuZG8GQoD92CzvBzULp6s/LLJ7QmkMqrj8RyQSmRGhe
rjPhfloc1MbvrJNDdMSfq01agLlWGvpN4Luz7zVbygTF2+wVqTLUEm28oDtP4p4D
3ZwFOAYOByw0N2PXZ/YPNhl2zDWMR0IbvCuycH2P3i6K3D3ZqDH/6qs918KdHatd
u3gKf1C5xSbieqpaaYeKkPEFwqtQLrDSf6XA2d9kUT3rBrvU42SB1bJxANakH2nI
DcJDd7+8qfhZtf+MNe/nowGqz0zsZBS5TFM0stSpo0ZVr12i8w1b/PXD+F9Fc39u
SO0iWg1sdDsgf57yFMMueX3UNg6gkdBc6za/dZrV3vrOg1Tg0Ekq92tFDMRD4By8
XvKCkDI+qz1YPejN3U3Ti5V2qge6I8AKWA1fKu+Uqfn9sDq4LY6t6RynVXDPQ71l
BMlIlR5d7deGm7g/9cgP923SGrcMEk7Rdg8Jsp/LyxIpDZssmoXaKSma+OduSDTD
t9kC5lL3sHkB8mhVhzy6+z2+w9Po/4SXM3ZfN01YDVhTFomRte6TwkyKgQ8Bzv5j
MsLtNhj/RiyhO5lU/FA1/+y2vVzcEQoIQ4NPaoTXl5zYkzf0OYMSAD5I69AmEYdV
ANeeRK6Azfc8QbXwZR/rPQzZ47gsOD+XpZ7vrrc4U3TruBRRrAASHvWh1WG3aJ33
wcOzdY3DkgyPTwyi5EdrVO7UkWF1aRpbdOVuZ9h9zk1a8kVfedPKp2EK4TRr2ajR
wwToDA6c4U6zLEsz6VPWt9GKgYzvndC7X0eWZlLSeu0R82IfJUqaXJotuNafVG5A
0BG+ECBVW1Cghez/3yvbmIYrNm3dOydsSZwL8M5VrOSoICyfTB0FkJjmz2gVxlQu
wtqwxT9l3X4bT1zAkXuYOVBt9mqPjfXSeQAOi88TyQ8AxkOSHOa/mQO5FLzy7/0V
7ZDsLGgh1V3kUJ1B1kmLI59tl5Hk0R9JxcchKjZlsE9iAzp813jSK1yrq7ZxaQS1
gg36AC06DbmZRYa0OOVwkBczfHvIJO3NeDL4E8nbRtWhjnNC0U4cqmn3vqIgXPTK
xnGAVQHYos9md2gFAenegkgfhgWe+GXykLVPNhzpOHjGHma9ff8hGK+WrVPr0sWA
YCTag/a/uOQre0y7rKSXL0tGk3R5qnZEHfI+fI4F0SnbU7EWSJox+gmFmI+GjyMz
eDZijbj3BM1I4rWoKPkUOMRw1DzNH/a6nkfudWp+SdrQ09swSkbRlthK5XPjKaP+
kS/ob8o6oQ7rrOisYjxMOueeoTgDSTW9HIoez7dRB7OQZWSoCetB/xtcAPnuQSKT
VjN7FdjUCeqQ6Wtp29fr6tKJ6+C66JnQ6gopGGewZCuNdrNC3MMZjWH725o8YulC
v+rWId2w5yscCQqHyNk4+gNNKT4DAUQ+iQJRJDiKD7QxeMQ2NNB+hkzh6W/mU2HA
WURB/NoqvM5gOXc2UwlT8evfu7jl1tPLWnj7g++ZpBPke6SqAzInzfuHZZjzN8q8
iEMrJVYUA7QkKytzxMEMtttrDXdsGE3xpe9ht7z8iNSLVRtQstMSctTajv/pZerc
OWYetma6Z5ZD33vhMls01jm1de2QwVvDPaj8wNuFMOq0/o/OJn85pNs9KX9hidzU
Vli6vErxvKYAfjayUKbyRFkAZPKzkVuXiXdjrxlY0OqBAYlJz7IWllpnZrgrThW+
XtBkRE45AzDgMfdCidZ52H1FLMfCHEGq7M942GhnXxqe+0TT4m+u6MZ+Gfso92pg
7aTgXTfFU4ahfpofWf95qBaWTkj+Lmvcl4MG2F0uZodX7C+E1LEQJK5IezoQsy4y
LzqsfKT0kZfuz3dxwWkQzFs7C9UxojPl1KN28MDwagKL1toTH5E3izNY9DW6V6x3
lTFgQkTPZcXbfIhXyF9AgA==
`protect END_PROTECTED
