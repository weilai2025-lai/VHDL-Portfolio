`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRFK0ghqqtHT1CYBslaFw80IY2IAT3fHZzuNccQWfUF6RtVOaLM1+O3k0xElP/+D
8yNnTR73/hu/BZ+LoEYDpCAkUoYTMZyXgoGqIu2CZet263Y6AqfAi47L98yLUzj3
HH06D/sB0rKKTq802wtsU6Yp19QELKhaVjudwrzzGcVb0WvVtEyQjQfqB5js6xvO
Ih6e/A06ysyYpDbFm6zuxX2TLaKtDXbuWM7qj6tfSPLQXfH/Sk8PhWjHMzTBd1Hy
6R4Fn7zYuGgfxPt1Jib5J/GPRb/+1QO5aLCWopPW3KX0NwVf26Ge9NkgFFBcHrD2
eKOpJwX+QHcexIYlSKiTKhxfuhigwNufBBA1Ns12UVh2Z08Ov1w6A7DNqp3Ey/hP
DZgWAjzHldSHDi0NDfZ1PxVWexnKL7TgNk0gANFXMP+qHI0/yvu55iPUVgnQVGoV
+Wf1qCiTsPc1HKCX4gfdfdiwCkBZeL2iCAwZ3zwB3qJSM0oy9vbjEMsAyJzIb/WW
h+HgeLoRVzRo8fjkYjz30YaDtai9Waz48typeoqDLV43ttxREt7oTxD7jwTDGam+
ccLiYrj+zku3aZWK45itAw4d7KsvLn057tS5WcIheCh80UAGfFaO9DdtBSQGKQB4
cvzbb2HFkve6B+rcqNyP7pbmQ1916cFsceOS5tpC0YTiyZQKYHeBz5IQYBdh9zeB
WieNSaZufSvKiDupCRFhXFWLiiPRDtbEnIM0M1AzqyHURN+ClTwONauUgFIsMP0F
xLX3lgDL47ILkIDG6GeiPg==
`protect END_PROTECTED
