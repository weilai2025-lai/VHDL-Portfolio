`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LfDyUFJykqXOD+bfeuUuTS3PQaC35SDJsFeNBvqLhXjaAQanS/Su7c4ovpubtSh8
jcOqA+m2xAgX+CniefPcP9NROYKX/qfUp/pLPNC6F/oVD4c2OF75N136xOIbmRTg
k13oKRGN0/SPTh4gG0qyKe5HiEdCV/zOqXK2ND7ZIZ4/ZDYrQw/Tz+V0KvjvYFaH
7lwWpgW/vWHUSqIE/+STQk0fxaW0SqXsgj7MlYDy343X10X6Ns0dzpbX6Cck30vK
R4aW3B0HPQzpLibsNJqGFPqYzDVhX/ZU7l9PuBCxJ8/gg95RL8dIIxJXa4MSS+sw
uXEHsHyE+TiyGr9GGIl4tqLYWfLs7EUahEOF99iMPgWnm7l0Cv8/ws0wChO83faV
hA50Ed5GLnOFvm01s9iUXyXc37kFB29vj6IXnZ24/zUlVr1KcF99mcSJvz1LwB0d
ZUpdkFE++QXamkGt6+l3Y4+GWIYLXJvpocDPIih8fYM6xdWjRLSRUmgJbXUCEx26
c50uQIgYK2cPgDaFxEUm4PcObrOdINWtKj2KXlhDjFM+onUrNX+6vLa7pCLo/l3T
LcVcCxJARwoaWJO/cAgjkqwcDQ7OPAOIC/DV/7/CBToBrRem4vxpj3rRt/LOao6F
zGk4HbwK1gQcQGHoJG2nrx/V1BCbN6mZcrcPe42hPascn4CtVsxGvRoGMEznHMMX
mSBq8NDNym2C6Wd30wT8Ta3tiBMj7jgq/7EDPRvxZRazFVsYO22lyHPSVBwpxbzc
IvYNrO6h4P10R/AWvDI3c04FVJbJnyl807vfs6JkhIpzPrprn2M1K6jCDB4nVdI7
ok1kDAT4fpBMKo1/lD/7KeqLL6vfx0543AqdFGCZrnNwIhEF55DiQ136YM0RLJGQ
R14LxeMv+pc36K/8hgB8jAxOqApc3K7gA6lsjxIaonM1S09MkTQ2Xzb5f1jQQeV2
T+59D0MxQBUjY1cvx4AMuM3fb9siBouwF94F6GFA47U/aZ3//TVjjDIUTg8eEKOw
B06Eo6641yBaJlINKkZrSm1UrGI0tdwevLBVlAQv+i4NS0CZ0oVtLvMKvQd004ED
/u36JMiXMcZd5TBuNSMaUas/rFO6OwjMciryCKFWvvDRKxILBWlNw+ThyzsKByXy
Y5SelFsOwv9M+zI27MVSQjz7ce+C1FGGEyWwNuinzmNeMEKj8A5sKgZdlKCP+6BM
iLfFj1Sa+HiaDMZQBf9BUnplJyelbSci2PWc0IGD1iroR3rkjdn+mcHX+wCExKvC
YaiVCWAAneL3b3IOtPI1Mg4BuKrQkTXI7vbN4lyiERQXoQmRugi8ZQwFmZ6kHPYC
DC1jo48pfSrfE7bmItY4giEXF8E+Cm+sJbhI/PZAXESLqNWuvRH7iXyDbUw0wu/B
oNpTUpF9u5ZVsZoR4liIz9k6rjWAYtCpSHF/svdB0e8iOIMiNAzo6OrK6ZhISMpH
t68P884yvGfUvkPtbMxEnw==
`protect END_PROTECTED
