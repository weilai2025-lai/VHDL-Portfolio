`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6yuE1KOr3TztYAtVbIzN2Q9S5NMTsAgRtq099OqsijOrtWveHDmeXif08mKsB/A
X6OXKXvjqa454h9KLq7u1LWmEI90YOAdIiMOt1ST6URbi6cX7dkhLCsrBn7IYV7W
TYFZ5id5C5sR48VeusXwnqLoHF/NVW6VEHzEKcxB6rtWlRAz+Cr4JwBb9lZaXZz2
jdO7h4I3vzb5O5MM2SpdoU64zPYVbgc+j6TNbn2xkTDNVqTsP+fQLFShWIU2PtOd
wdzYxGKpkGIqx372g+sOnOydXfU5lWHnBl+QbvZJYNp+eNOgF3mQOmVMJqK0HoNi
mYf2FSa7BEl8BpMRFmdmG9S9E3gNiiOeP96jDq0tOUGpc5H/ljVkKQLOWLEMBItM
jjSavnTWK3GR8GmOidVbkRq+6jIIqVbSEl0XhXV1q8AZF0uvn/P4+iNGPP8fr5qb
t+13lLjOY2zLbnltAALTKGnJ4oR9jd2NS8Ntd2DdiIa5WU6Ph+ghu0uKlRTUz6OC
eOMy/3cKNfIKPFN7DS92hvFwsJnM0arKYdsegVtRD2JnPguzwwlk+TzaiIEnwWXL
YleP6YJ4xyTkrTMzZKTJb7phdns5Pfh/dOe6kWaxJ4fN8fh5NJyLu+LHKa2L7n0J
rAJ/kpJ+U97QI+cox62s0n9Io62YVolN9i+KplmfyfYt6FLgzaTWEw5WFVIzzvx8
VXQCNdz7YO4xeGrLcSfWcD5qa6aJQ7fPEiYcSiPjvN5ekO7rq0WRxA718N32upXW
8KhFbBaU1R5dMYiTaDonXCLp4HAtHNLm49g8Zte4/WW5S1AzPjVkAcLha+imZTcB
yNHO89qOXAV96fVcyJCnQes6PC5vkyC9xTQYgS7S9nhvdplNu9qqICUe1cMaqU2T
J+XRMVCI1/3eYbJM4MzSQiuSzVWw7b+eiknd6gB/29GNLszzvqPyCHBtzQ57nIo9
JXZjTuBE0HCKan+sDHuAKuYaG6SjJSG8PYVUzk8ErlVesl4Xw/Nh2R0P6zPHGJDG
PgXszBKk/12fMAEXIU0U/bykZdUdeLSF8dB3AM3ksn1UHaam1sGwtlNI0ApBEvy/
lZJUrdxgkqAi+WAy4TOtxUb91hABgQcP7C/+8SOQeuo=
`protect END_PROTECTED
