`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUwwN6BdMDpVzu6U8yjYx7eVPIROHKi/f7x65HzPl3claLD1Hjhm0KKj7xiLbivp
T/aQ/oGNO3NHadaCYO726OdV71WzL1HJuLTaebp48Zbr7u9Inpq4mpgA/vwPhWw3
iO3l5ODjirpmMi/xPdpEXHdLAbWDUNkqPuzeTq7zkrNYEhn3oQ5kqIJe51HsaYaX
5Nmzq+0Ppg7PFcYCr2DD9mNZ6WDPHmYF0Qp9ohm3mssA3Xz1KtDCDZyZI8uP0xwn
db8QyvbzZMzMJ6fnF75lFDkDb0AIqYso5nvJtBeboTXFS0rgGP/yn8Q9kHEw1EG8
63eMI46HkiCN8IZvJmwxzNxw8ed59ottNMGd6D0v6fBA/WUnmSRf2SfwVmzRwTsI
LT7zz6QvcOzf/m6KZYJrmDEF+1X+lDrwUN6D2tKS7VyHL4PwDA7t/f823NAyI8ye
rXFBBpJWkYp3ZNbbHvZzXxPSCf5n/U4vYwlFAdslSN1pelvc7i9YEk8X0hrOU+Un
wY51JYIAqY1Sw3CDqOXUcCRAWw764mj1oV6SYdAfUI5F9BrY6ASNUZbxgng1g5+3
6svG6NLaUovKaN7NjyocfVbRerH7n4AB4HCZ/Aecj7oQuWdsu2uEPqheZUBnYdTF
kU8u3Yy3zAW3rwsnzBwJkUdXLHPMlNgy6EP6VzlN1PFLA9yMqi8ICdvrwipbJMcb
n7TiHij8GXOv3zW5ErlCmN/nSNdeHdKDMTLORnyzud7mPeWlIMZ7P1ZjDRgVRUaD
5/c9VDEUP1qnvAs+1YX9gd78AmvxWCuWlDkOpczLwcoNB7sVKEdXsBbzGYwmHcV4
SMnOy83EB3GlZl568mY9w2DqM/I6Dhd+48s9m4d9sxpndwzqWp6WVWl/8NkB+8di
M41U3sunEeRrTI2UPhC7fRJUo4+z/Ni19Q5hA5krQr5J5FkB9vwQaxssAGDWc30U
7VR3Muc0SeO5H5rTkY6nWv0fMaDXHUXQaWlsYhwKP/P7829VyqkufQja2kjBJtZ7
YgOwlfx3efshcUOz2atPFVfdYZNzfgXjtV1oSGXX5armxRuWdLy0Y/M3cA9H2Gtb
6IssYoRhR7VxXb3p91q11+H48TiLz3pCw2ohieCEfb9K/h997aOzBt0MJH+a5RKU
/fKm3S75ti4L0YRIQio7MeI+X1/pjgyAS9KXpXppsenK4GwHjhaDmYHd5sfqVLW4
5RaSO8iqaMxNN6xc+KXT2FJWcegpaRWGRNIGMjCPQELDDzH1aAxDtYD78g810GCN
5h4iB3rDB+jIxRwtShy0i9t1djfHdgSj24HbbG2pvrB5brmEQRD4IU9qf5MItWLp
fc8n8QaReP/uNY8q6AWOSvyw2XNB7X55AOHy9t3HJPWU1cY5dqrToSSZhX9waA4X
pXJC9wLkcrC3fhB7lcf0Vem6o0IY7hAqF93xnSlkhbFKIC5OqSVLnSzccgaWvk7j
gsczX6Ey0Dwk+i6HESCtDKKAngKCCpzqw/Sed1Q2cIK5hirpfMuUvTZsBoMTmRnw
qd5JJFg7lFKKBH1MNoiGHhYJGCr5WmQzp1KjMtYnrgAtldlIBBkSYsQn0t1dXKkU
YNwzFfHEZCq8pUm8Yk8US97WT2u4KTypDCCZe/nOlkRpDpQt1QrlKJAosLpa6zf3
nmmfUKBmqGLWBe3xVNIcUtyOFIQ/7zvsFI+Ke1n7PQJTV0nb3jXF8/Q0vDbrF2Xc
kDlL+vdrbrgF9xfw8jMkpANXrjHw8nlpfSaZwdYjLc2WpnxCtATeLuibPRraRsh+
bSTpXy0you/eu3VR35TGeVtgaq+paYWsnZmAA3k0ZXqM0R9vlb7fKAc/okUBh+x0
VDFwObNG6XugVUqrFU4LhwI7Qpnz+Z14TjoymfwTeQEmE2H80iYkQSa7nwdrq316
l1bFogCswX0v1KLuQKxD+BHTKNIAv+oWTBgW1nRxL8gje8DVImSYKHNGNn+1hh4d
fySBnYHbfJ7mvZwYyEQaTAIMPvVGQxTkN7in5jekmDjmIrIBMfc8XENa4RoyRIcc
gdhN7N3WXPbENrHRaIXey71eyRG8e3DmcE1V3gZ1wFFVbiG1ieCL0ASwBzRHv9OS
M41e7WLQr0hCmA9wH7nmPZVJ5tZSS5uBzleEShmK8tTHzTKEsgmKP4yNMNOZA65U
yc4j6OhevF72BqqQGn6BDtXORmNA7jJDsCldWDMgjrf46EYCWde1PjLxcY3KnD5U
jSx0YbTisLiztMwBTW4yepNs9waTbjm6lL+HMLBdWjuo3jZ+CEwrUZqkQZiRJmD9
gyqnA8CgYTN3Tt1ywM2k59FKtbLtQO8s46I2BbWDJPF/QU4Bp5YK44UuOGslqhPX
S4z2JrAsK3Xi7KeU8okLgDqaQW6RDHAFDE/cypje2pA1CMBYycgaohAE3JXqtRfG
nL3II68cdh9lxxBxOTXNJJ6TvRlapvUWHQuKtU90d1pxpX5aQxiagYKNJyrSQg56
Lkn/tJkUV8PeUlbW8jKdRe42ms7RVUoZw+ql7RudwFgSwPkwPorcTGpODIahC8hi
ur+9uOdTEY/obL8vWLwGBQS0/JPBrtC1aWQE/BG8zS7JSpNaFhZ73Lx6p7t+EE4R
aUI2JvJtFFTdG6QP526cTlI1x5Q4rHsCvzUTbIjZ9JzKW3EWadwX/OxsxK3+1Q9h
ojluu3x+Tvmq2evtiPARttmUDpoRowNCMCHr3P8b6qmFHT/aapxv4igiPqy4Xc40
VFBllZ1Qt58RrmQlxRkbVxuk/yR4jEjn3cCjutp9/Rs82ldXH8779Gzu/H1SDZHu
UCmSsZvB+ZL/0VUTOitjB3c8YEFwnlFxtFNzqcZZdXf6x6XeXOtvIb4iBlMsSRw1
tHlvXLq04vcmB0J9PwWj6BSQbiGL3Wp+uDlZZEVP3y2dkOOYNjmjv4h2q9WKYJF+
caAoZEar2N8CpVDaLaCmMy+LWTuv+AfwTAoo2pCMW9B8CnvheTSZB2vpriYKBbei
0odzYteNLTbAHoxQUyOOFTLGtEP3ltaiqwNDnt1vXNnf4G2T8fgOpMJ3pVoK7dIj
uvUGWZOA/K6A8Ji25NNrDS0eBGT/mu9079TDPfDF0lricgAcY4XjMup6wBwx0eoT
912NC9dfddixUmKRmi8xHXNfWQ3J7i/4tulTCTfGLdnNGht6P2IMlXB1jgGRmxe/
YSHnCeTBM1iqr1W+87opu4QHeP2Osf+CNYnsqj4tmCV94UDdCSBbVlAq7LfhuCht
QdYRKqonUCusIAAMSWDtBRh9Va+eq+fxLRBl+ob99jUyVe7Zzl622QEaoqsUuy4q
Cd7AMM2pwZKMnCDOpShK4p49b4QYHDLM3pc9s9i0e0C+ZELjpcMKm8jRYH/b5lGv
/KH0JI+uKjS+2e73ukMrXEBIydj5IpS4xtqktKqity2XuOmmbPYlVO+2XGxqCFxb
RQBez0HHcV6BGxPhlx2j1ud0Ee5bzBP14m1BauFAomItN8dMOkcfA7y8x7IMIuuG
dJ31/axNsF8Y1zG8tnon7CFfUr59ZYlRAx+GtGZ3MASIyiR9+T43Y2IG7Hbjovp3
nrloZ9raU9+qMrmEpiUtmsPbZFRnlddvrRW2elAxn2IL6CrC3tx4M5npZU6SRdCL
qAygDNa0vN0F+1iOPywOiQa4vUuDfDibGCpDUg1ZTVBkPDsyQqLcgGnWIGDSOFhf
1v58MuDuYFiwppwhqAcAyhYOeN9CFXM7wmnYr8FM4Iq6HaJ70wgI6YGiB4LZNONc
Io1q7L2+yilahgL1Usv+sOzWxpKAkQGAaI2PYJ5+Tv0AOBaRxUMJ93zlux2pJis6
9V4zsG7CxkXcPYIGNye6RFBY8e5KGWfVkKPdo8FnWP5Apcbx1GoxkLsXVuq4mLyN
fWCBbZnbbMDZZPL0OUOWMAkbM5HDx8ylx01C33mr0MhBW94xqnDGbda2qsbORLlk
vzi76UIutkMLHEg0Rmw4KA6u4c64ZblPBtktSu5PLHLb66/X/5j/zAEdrNUbnshK
HTDfWYNST00Uj3Ybk/iUcMFISvOzT0NfAkFKdJYuJ3ry6ORmfw2FDG9OzYS8ZSCO
7P0pp3wrzpGc/7+/DcFZQY9BNBd/XEr8t9agXWdExu/tuMv2nY0IlOAKzrKWA/Yy
NwSva+QZ9aS2BJdAtlSEy/TCWJx95RB93T8jDKpWRwxqg7eOgPBRevgiC4wFAKuY
btMPWFSPComY0aiwmpuB609+OpkFELDujXh+F1B7NbfvftAFCY6F99Z+rMB+nSaH
B9A7g3bz0zi3/+QFgBV39k5u7PodRiiwU0zSdZ/QC2Hiz4ITORtqeMorm6vCAGyJ
mauEWmDNBe3QDtmbImFQwWW6kiY2WeZ/Yl1LlKc1luZHIJ8vk0k2GgfNjH4uzSAS
Itoa0KTjxSR79aN+nlIdZc0pKWUWf1A5O1X4LjkrOkpkPWboMqsGMxQk3kHCOd/4
aquUcv1kWShkY55SO5CkChyvnOp/nz5QuJycgK9o0VXtevQD1ePtMcxpGZ9oVrIG
btGGsshMlNjUjqyPUQNaXuPNUsosyDEwPhGQTBQoQRASQumjMQaVsgkA6WeOeRDU
PbKDsRcTmVrlUAylUc+tQoazCgqAcQ0kqUvIv44kA4iChyriSWBoLbc3ZeYdYUZC
QkhHhyXUpkVl1UKlcik7wVXWcSDwiSdENOe8fHUZCX05ctbCOEww+/SDtldaRLU1
r94lEIgUfszXe4SsTpEhzoqfXEmxG2kpnWtEoN2db9JgRArtfTn07ModyRVx/0Lu
7RB8P916ytULOtdpGDNDV0V/K4QXWBCmLQ6XfFBD4ogOKJJyGOewgaqyfp8Ydq+d
kGL3qKZX/ARgFVIJ4suqzv6Cf4rQ9TwgxtzF5cSfsqY7bV+N/UVNbudkrl+ScmTQ
oM5DkPpKSTp0bTpJwCCO9/UI/lKujGIF3232dakQl0IU7lm4C1zaJMSxuwpSnzx5
AWK0j5aU7ijj6WOFtlL1O9FDXkLjZx1dLqOkiwzp3KCxhBI5z61ChcXFZsKX65Oe
D8XOSETxkDgpeb2xBCQ22oIAwlON81+fhKFcaS95+54h36tKuBJp8ipkE1HFrPoq
n29TJFqJ+w2v9SsgCvacqORcKwIGLJ8LNgqV9zttWDytYq5WYngtTfoh4WkXEEO2
YpVOgUt9+fvvFiN5tbuJgDC2OIRiWFJOq6iRPITGwYHp9nQupbfAQf96pTjJ1i9M
5pS1koU+pwL+V6i5SwCZkfTWl87w1qj9C4OvEHrVNM5TnWbMcijNGBgGLgN7PGb3
RCyS9eGPSkzCiVlac1+vjXqFPXzdvrBLBcQs166ulpS4AtGJcoLCGgzp8A14xv3Q
UQqHentIHHwxfeeblIgyzCsS1hVzGpXKE+4r4AnnTf8RA9jZprQ15MYWfOBRKba+
F3ZhaMC4vxx5uhQfX9miTjWt0iTPvoUSZIj9+T32FmKYUrg4v5NEcjdd682ncwpJ
xdmFV/OXQTPV1Zr+e8gos6qoB73cmcen0CO38/TZGZ9999vxht1E4/h2A2PVW2dq
/EZlMzav+XOtqygPA0OWIj5YsPI5c39UKjmGuDtecrnk8cbEMflf//OKmbQjkLK7
sYx8NM3uDM0hxu+aGuX4pNX4AuF94qr97kGvUNGUfk3K7gxQyq0o6Yc+bKYtuXdA
WH3hSlcEOZ7sbjZIG0/j7/ijYqbt2YBjVn0k0BD5BCvmHHb8rmg55H9qE3WSkCIR
ly5yjvzrBkhfV4fQ6C0Zp+S3PtKHQiNOFNguO6WixCQSY2z7ABlCqzwgtde0jVa4
HjRyt+hyfHAAG9cGP8k6mxFDvUhDeiW7bF5b1jeMsd+5rHDD0Qcnjv9h2BLUh0OY
FNp2XOW6W/sCxs72KuUu3v+DI+sQDZDZbYYv2qwdjvoRkC/sOvyw1VDf1N+fVsQe
aNpMYd+XD5YlKLL3sveA5Z8VHvond9vxA0PVnsQMYGpDJXN9jThXjE6WtFLtNcnD
q+z/x37dOneRCPmAEXPfHQnjxxFVm8bdNlaZeDT9Zg35Dfb4S6/UXJ2N0FDOny9B
3+Py/rGaoyJ/Xv7+LR9HJeik2f+Yuu2IRojPD0ZV/WHlIZwYbObsZ5NASUELHEgf
gt5oCA5DuuQ2UrwGSin7yQIL18tpmrtaKQ2P8HyLDc9Kz/t+HoO4zAqf3IshA9eN
ubIn0oOwSoiWmtKSmfsw1CAH/xHGicUhmWqmwq3qgD4kXE95g3Sy10DMi1X55J+L
KCGmyYIkHfaPlQjO635TE30Fk/vnAZ/QCj0A6dV44MBpZk/jP3Ur+sAK52NExmVg
JeIEARyBsvlcotCncb2xR2HXDQ/hYSC1qePj+4eNTbAIOD1ApKfmVFLpF49MnYid
gEQti8IvvyBYCnyB1cWKFLt+S3uU9kDNCeQ6TF2QU15sQCz59hzZBeCw8fsPZ7IE
v3o7QekBqLVfQpVbECozV6BX8m2X53O4x/HspwDB2mEZINqgg5k6XCFLFEF6Egfr
qqEMCZ/HuyCRmxQFRNy06mrT7+qUUAoymAm5AuFtLd+NYIu/Tzs+hzEhnG2GZRWy
G3JyVDyWe5AVc3wT8ZWY7Oh1IAnDIycIn5ICJEc1tTBOo5JX5Hk7srtELJvONjMP
CA64RPb8sVqEF6M4bHV6lGmg6SWKQjgKm+l3+5NVTFFxf2HDF4+rDUE8Azp5Bv6f
lJZcqZ9VZdVBJzv66XBKlkzneC6vARNklqyNBCcy3vSqpBEHhpDfQX2pAQDBwcOS
cIIoS4uWjh9y093iAh2sgVlhbH0JNQsIsAiA1LUJd0gX+k8qN7KGn+WfCkmSrFhZ
q79GaPT+K0soC/5HgePfIji0Q0pxLR2M/YApyovrQHDrn7Vl8NSqC7la6Fx8DqAo
n2hM+kGbw/IY6Djm+F3PLUye+P++FhxJgw45mIxkuMx4m61M/ssr4vp9490Jd14T
wctLJ84Dss9fqqRIa5Owht1AjokgXUMlTaqYb5s7XbYULU4ouA1hayWPKQQVhYQa
EWynd3XWE2V23jw5ProKei2ed8IIc+mGt2PkUJIkdU8Fp0rNdzVhvaSrj6gkqn4L
KLk4SvvETAwsIbTePU5uI451ungP5j2JTCd22Cn5LqvfozjDh8XPNEqMy/qfLAQd
wcw17vcteK+WnYjVXOzgxc87UjwoxwVPsJTQ2gi11c3rlczq5mkYkslbpicGrsD/
3IB/q/+O76MjXPrFwEI3zEsXS83f06OLskkHlUV3IUB2Ct8vZlnTTUkHdj5bttkD
8IjacCNN/q7StacehWRzJ1BaI8OLZ8ti7vXSheiPw2CVNGhWR0yVIo2u4G74kaO5
BFnabnj9qYchuH8JgI+ojF3TFvz+2b4Wu3IsfeG/QepU1DXayTfrr14xfIrmU2dh
Jl+PplQsjsqMH4hkWs2ssUQa3tSrknW5g3ZnEa6ZR1GLNDvG2XW6IXzRItFkGHcU
r5zCrgUOwbRxo6OD8GanGw2YYkK0jnXWm+V6IAvPSWA1ZhCwQjojFtW7421M0nCx
wjXZJ8+CPYe/BxglyW9x9SSB97JDqMv+1981ib/vGFyKnHFNN3WLBtKj+Sf5Knos
eY+GycsQmzh7+W35H1tn7wrbzXBTd+scHC6zHkXKuUHA3FGpRq2Fc/RGmlyxC4Cg
3mYw1ZNr+flsYb479G+X8ktIlebtseFSyu+Y7K07ZrhVirSuDZZRLgXGnesRGRjo
cc9fqY1wazutxcO0gnYDXyD00bVIFtdX4XTSy80LFZbwYIt2s68T0+UUM8k7+mgL
PWZeNpNnREsO20h/6FI8NkKioibUM/MB9qNzLAPhIWKOrO4qw6xqjE0gCy/RBvmt
gfKISRZX5zZtM/U4SdwBrlihuIOKmfhBPBboNYogEi+/3eZX5C0EZg/4/CYzdsdn
RJaNTWjwk/BtF+9CmYea2Yfk2sD1qCltUXpU8w1NYZsFtCI18z5a1/TXQOspv95M
TXRMci4CNrppRvqY/f4T/keB+lG5GLtg4d6ulUhWRowJkVUkqP9DVe6eS8tII/2Y
Fw5vIRQ3Cif/cSJpoWKvYYUHlwwSMOL5DlG1BKGv5/mifNRrf0E2otn+Fcnle/3n
KKX4LD6IX/ehuHCR+r2PW1FdcSshm23BGEYwFRGK7t1nyiIqkxumr4tEn/UOnCnb
SEwp0P5UiMWgbX/61Jvqiam8+f6ndvNk9q+4gI3LSK+hcCf0EbRLrF8CKTJwfmCr
zPBI/yr4EPPOXEcLdIGVuneA1wN5x/baSUFMNpJY/lwpBX7d5sBJFm2PM7kpdtwb
Lft+sbIjCF5BHHHMXlJHy74NzMjUukVId8IkaxQsU27KAcp+ttLkWlbgdbht1npI
5shH9GG5SlnbzK/4uOSWs8OncNtqioACrqpFb/E35Hw0Rt8ihjrfL7Om8j4lsSWn
Rpfi5awTqoVlwhaNagkETSxEs1ppoX30j4i27xPsGhPvRvdWn8Nc9BhPmNHICfRx
gh8NIEEMArU61GUdU2+eTxOF7w7ACZCzjBC/gza+UIyTa2tlHWSRjkz7NA5wI+aD
xMNm89Xmk+CKqsnuoSVxJ7+qwTvYespWUpWMotFY7PUFLWFhC4MgixrVZt472F9T
a7UHECc/wh/B7uKI2duHdN2UNYPRLuguwNao9dTYJmF5CBrOsbyEm4MQbyHbQNFF
BrekRsrBQ2KhBdD3A5qiEqPpBYEaRlF3xC57vKW35/JR5IhtNFByvfu8Fi+1D9LY
P7qxnWGOuWg5BX6z3NUM3o2J+z0U6ioQTHbucF8cUU+xMQ1Sa9u5tT4jG/BPSMfn
uj11EwRxCUeTftvf7D+cD7zsC+1uXK0n00UPXXzsJ/ROzRFtWHEny/RnzVHk6Ru5
Dc6izMI1m5jYfQP54QCcxvx/w84sqUpI1QSCRfW7gHgT2wAe+tbDiyS7d+jbXTx2
A+x3poDCZX0be7BUodEK81Q4sB8hej0OYh2LJcfS+NWu3sxZ/ZidURTDVpR7EVyg
HIF9YEDkEMhw54UdDBmfJo49e3eQb7rZZ7TWPPhNUWIGnNaQZrOEvp2zqvcezJut
LiQxOCf6mu6qk4C80CFP1DDznN3Yvpz89l2UsRW6/LIFkTS31PmAk4uONiN/cPPE
DVRlXVcT3+PE1Ucywgb7WI9DM7OxLROBuXuAdC5ew52V8MY0eZaP+ljtThv2i2H3
CPQIJbYvDVL42EHA79macFxsveGxxI9xzdc6a0hwKuiB5FAj6JK0IFiUKizb/XA7
vBI36yp2CN/Im9QNmPXw7wbystKwdZVQhYzOv/JJIkT7sqoIHHPzDhh5mdTldHSL
4sATwxUYlFflopI1oEPCavOEeJaUxBByUa0QPdlrrgt48GylVxXc4XhQ0vPpKO3O
tXpUCg2I+lxZXWTqrONyzLcPKeIb3WMaP6r3a8wj4Qw/hhrBIHC4CC1RyxGNk8n5
RcX2RAwzcf0UYmdAVI51GcoizQvRkUpURlvbUOEQR6hfIZTS9R+PMIF+Lamu46Ob
Z6okYViB/+gy21S/OHBHus5ljtYjohaJL7Bi2MbLOYWmk8tvYKKjv9T0nDwlCSTV
WFQL6AW8DYLHVnalCWs4vr9c/HttzwIA5bwSTyJ6tMbyAkUnypM7nydy/PW5Ngtk
sBi33d+35JzD67cK6zz+Jd8rXw7lmFiSm9KlDnX0KYWQ7p0OTn8/ilpmg0Lx+Gsh
2jAnRn5k9uSxhesgSunT89iNiMkO5W29atfy5Cu9V1wE997nw8vyffe0+MqMLoRs
X0q9AMGDnHVpYsa0Vv9XzL8oKA3jh4RlpVXW0ovami1K78tmdHvEHHtNAn8ESV0A
bkWMcOx1NQJKJPHp3v7jaJvvFtt3HC1FOf3Z9dGD4/VAsDeL/cUvb7nMkse/LpCJ
rUpnjty7ygDcIZsToEJfJpaN2LREXm4epaQGnI257vPURIBmqpJ3kqDqkrfXLQM2
UUX09IpjeWxecc/idpl4a3V1pvnmWoPsFxF0HolXy7n9/VBoxfSMngH4xrlYwuHk
+BqR/fYHzLR6iVjI+jtKalplMenK9NjTPh37L5sp/NT1x6oo+adGhaqS+48mGeMW
A4AR0U40LFlVoO6OQWpCTTqSmW5IZd0nS/OuezhQdEW6t1TZ5dlBbeLSsbAHEyvs
IVUmdqWOCkS8ZwCwKSFsmET5dBuRha3i4HY888wZF10mSmoMkuWVeHyUelfUg8bO
M6tCSAlnhmEfokaA0XOq2Kk5sAaOGubFGvEOF/peIMY3k92JsV8O/It5HMZiaiRt
lFne7Q3vdX0Et09mp400VR5YudnB/jlPXPYYazkothK+2NfvTKSxaOrX52iE9/RB
wgZmJsDDnMa7UTh/q47CvIq++H09KDl+BtNdpJPgTEUuTlwwNv958d3iKnwZfsH8
Rpr62WKZ66YAJEbNIMk3ZSosubqU/vffiQ34gisAmNKH0zvikyamGWZWyyaVlFr6
Yq44QoldvI0RMp2bM0lhEr4/QIJFYbb2Fpwy5WiC1u9xUtE4y1Pj2Q4qOHrrvWsO
Daj1QT+MsqmIpdNPhp0PUI3c095paeaVi0h6362kAIIafuKZvUh7nHRouBYR5ME0
sFeOUAhsDLK6OfVYWtujpZ3++i6HaSeE+ImWDtUL8X/TpoQvb9rD7sPDYcE/+qgV
E/HvZHRzTaTEMiJPWB3TDCe3GB1J+IAC7Dz7SHeqpHi679xPB1ZkGyBl6di2HDTF
Azm36hbkMLZqsNAmoH53tAATf+qNONm01wI+Y7Tu34VqPrEG9xDdQfZ4i2H+jDeD
mHW34IDn1HbRvtAMSvgiIrA1tmQaTrnw++tbB4imxtAl+29Ycx0SIs6H24kezCaX
bWcfJaM3lqiLI5ASEnrZWndJvAtc2GIQXqa/JUkoWCVJM7lpYleGue+Ky1XtNGAj
xKaOVxSdc9mDhcUmSStH4mNCAGTUYQ/P6BPTtBByArgG4EM643qkDQCHSF6OLGVK
9lUmU/1ZV4RMzK09wFxaa0BmN5NlaGAOpPpxwFI83RlspMohtQ3Z+WgN+NA3RWHz
Efhz6dtTNs1ika4XvDXyyD8zM5sDUD15hUJmvZdxHEAifuFcFU5vPsXQi1l4v/Ea
CVfSqqHcSgsfylbHRfi7nP9KSjdECMpGq4lvmyulLlNXyTUvr2vigYOqAqCaft01
35lRpwddYD9VV/d11/Fzf7/OD1kA3pkV2RMK3jgn3AT81mX3pFLNvIx2byBSEq+R
xRH0pZapYHT77fZChVu98pTMr8WBIZ5LMpk6Kx1Vra2RSaVHmdTxtn93a81H1kuy
bexosjOG4GkUwWTnMNHXJsuQYub/FJrf7IcoihQ23uHQHahM8ZI5olbkpn/8BW7j
8oacQ0TMmLG6tfREDzNkj0oR8uspTvQ4ZqzALCsgGOQEd0IIm34f3Yq2jsqPfU+w
SHxReoERLpD/lfX7E6STFAi88f20kUQY4iF5GoMZLZ+gNTq0TSVxDl7pWRTUNS2S
1jJIZokSrArpwKRmcQDdOZFbV/5vsVCdsb1vespUnmzY+/wBH0ONyFQpPJWjT8dy
jIL5f2wgISjZIzk8ELzDOAmQf1FKa5ha2I7SRTnVqZAT953JpWbstdHPu6jPPq59
W2MfJpdHEWyR3HZ5teY5eL4ydFIHWt0vmVCc4t7Oc+oGsk0D/BHE8rJ9KuRhdBRl
HKa6hvBTnSCONUDAGVAOdgUbKoHJPXFkYQDoCxLq53sjZK9E15ULfxG/F0gjl2Fl
Rh+HDP2Nwqi908osjED/XCv63yMtDeQ54bKmzxnHVFVH4bnhVGH2Fe0f5fBE/TTl
1aD+PyydJiZ6fTKRUVkj3S85yfZAikfKLxmnSqxKXGxqo9oJDTGE5r3znOzJ2CNx
G0qQH8b1Q7SHm7lU5BCMLrCXUa45Gawwy6puWFOhz2tcq+JBS94fqxNktcWr596O
GgKddTfKANLan7j9Rayylt7TjmF888arIOVCE6q1Cy27OYM3u3SIJyIL9td36FBv
rYL08tdzZmO5anT1iktDnM1hbWlL1gAUFDcPbXBPgEmZKbrCNSsuRvJz9BEhL8Cg
jG2Y4J78KGCvoly4zcDg8s3u0dT2PM6rlvXO8pxdYTAJkGbMEFj6nVEO4eSDDgXC
fdxIyb3MPA+2PgxwUvMJISiIr5l3ao8ZTWceDgzB0Fpt2D07uiYkkx6r2i8bSLjy
FLuh4g2LwnM/hMaqav3Ua4QwFWi+Rjow4cCSkBhYGGIOkiWPj/xLxQkY2OzGmeKr
aMYsI3HVjp6g4zoS7+BiUqp4Zuxfzp0/i+AgkJwSDeXFQcCBJ1DPawOLcF6C9cDh
JR0WcNn2XvbaBbOSjZ90vHQYIPmfOfeJruiJbkkrvKogp/rd+uhLtLDNLXoV8xmX
aWcwcbcgOZ/Wopl2300uWs1B1ptPicTkp/Lg9nQq2/w8WQSt6FP0GE0tsjVyJv1f
acfHwDw78F+1wB8VGjr+6P7RLADkJljdjyriNw7NGjaZ5kKgCAEaZZjxHwQr/0CH
QbgY1k+ZwIF4ss8h/fbXi5ForeLS/xxUJicCZ45crVcY1ItvGetExRKIFUAOgeU+
BbAxw4xxSw3I5wpo/mMCJ5TNZw8jFI/XMZ5t5FuYOii9JPCyHUMShWsgHcijB07w
JXDz68CNxGkEgRcFAKhfWuY8FcBEKFZdyCLLM1p0wM9RMbHZ2Y+65yzN7WedYwtT
htGhCElVX20tbLXMrtEmezXthtmZElvp89Kkw+O4okjcDpcvgSgvZalbw8+qkyOc
N3RbDBKcrrd9sRxeDRehJbrnEgKwmW0CdaRPl/wisFd8AlKXGZdjMD68M2zYPDbc
Qxz4C2xcm6Oj/wXGI1hcMPOIjhOknCRmWaQzlHcyk38O7MASEjvPjcru+SUpfZxH
Ir1+fqxoBURyETEQo2PPUh/ICvPwHuRkEF1UTz6d7WZmcwHsGhqips8P3id2TbUT
J5918rhXhssdeEwqiBFwEoE3p482d1D3tIPVM942KoUSMzZGYJ1tmNAyayXFbrrL
GDWz0x4V073iPBkDr5R9mn0n+d9hKI3zc2LXW4r95XFBTJq4vBtaaWQzwPDd3ukm
GchmaxV7gTvT/VarajMGG26O/cnMbgBEEi7onKZ7SkkGOZ43ocwnojT/8k7F2LxP
RrLUkGM8ck9OvkImfVZbTPNDcbBFjyHHhyr/stwe9yzGdkv+cErMCvAVFTkX6Gzx
ATv4pa2tdn/iEQq9RttvQQTmaR/vOnAO9br9Spj92NDPZr7Rcg/xr78uyNMcfB9i
+S4f+6KslXqUJcjyTyxM0UR0UqlDmbdRAJbg40ogXkLM+SrpRdhCd3sQiHZDiTtE
LimqTNa0BRgah+qi/w/FzTmI0yyS9p+cel3Em7hwL3p8R+9xLbxqrsTmMsBbSfF1
gOxiL/Pl1xbhrkOHg4wTCd+7I1dBQxzDcL18ENAVxoTxl1n5KB1VwQNwSOprVh4i
jtv5sbiBsQWdGBe8d2aeIH2eGZmXVPUxZQI3OlDsS8CPMgoNcZ4aaU62r2hMeGgd
+/0U9RvP1oeRfVGcpJTLn+G84EYtLotzJnw4l4sgivSONPZh9EdCgUYh1iHybrI3
QBV3dqISwH5ugBMhgc8mhK4JTWgA7ebSEYswxQzXF6umZ67kqcwQZXf7rx6HWCvS
5GtYGOo5PoRIVe9iygcwHnnoxdHXmFVhuhaoc2KTT3CP7dTM+QpTU3/0fuNaeI40
YoGKx7XqobICCx91+YmEnJwQQP0roghF+JpZ0+XE34h3ISZCEOoLIwFACG4r1/t4
zIvg7POtoFBBy8IhRAlKwrL5nQuvtnpL84xtJXSw+CQc2Wyj9guE+zw0l6q6rKU6
s23D8L1O6aY1XOjGfcGMKKMdVYeknThDuWXAFjCCoJVlCOQkbuoNV/jYnIUxmXKE
xvgIoW60z4HQTFv4CHDvKpKDx5VnNp+/BJ5ehtL3zoMrREU0eMy0wHEZjqhlbvyQ
q12p2YDfla+xq1pCuMqTLPCeDR4Rmmmu5T6nEf2S7Lr56wB0q2rKBGrTRzVMgxh2
xZ9uyvWdZLRzdtFpff7TdOOe406Zhj3rfX2G6jjHA9UmaXOi5d2mHp0/e7QIW2Yz
VvC7JrswT1DVxkZ8Jmz6sPaNmv0lCvboJlkWZHtN8jJHvypFHNuD3UDHqUZpdqae
ZEoMR0mZkO5gtSxwTrK7QVurckTVVDylzzqp7POYLI6On4OIJJyoTheviL8L4cSb
6R/AEegkQuiHGOk6N5ZXdDvxXS2xalRxMnBBREJkmAmICznp+giQsNxr5cH+ccb7
c0VGzWVBs86LhthDtk+ptX3SX+bvq3NeiIqZembSvPfsTfFDOD5TAvZQ0LhIYUkU
BXTnDZiBYNBWfjaLT9spB4y2FDM+Tr3qAbjofiSMUFrK79BNq98jGpzvez4QbqVn
3MHOIN8YLa6Q38ovRXmu73yuru9h0BRzGkpwy482BQstKG6kPchzYOT/oUkSrBV6
ZES7maTv5Qwij3jqTSEZDKAZoqUD2DoRgv+Syx4vkSKPlqbMIAT2dGCOh6Sq3R/E
MWXO1SH1goQEXpyDqeDCOEptE29GWjsTv7Qqp9/g6GMxz1YBD6Jk6Ylvn3Mw0imC
5cCsgPNWt/XL280q6qBYXRV9ak9TIt5+t26XLCcwEjVVhtzoc2MStQmB21Lux0M4
fJuzfHPc1a102V7qy11Oq4LhaV2h70QRNcbbphN/AqruCTskuMBqaj9wKLJ9Kf8e
DuRyYBoIG0V+gY4zwCAZJclgBMZ4a0C0xDawFux9f7zC/gBssKN1hui18ZximXAA
tZ5xsmX2SE+I5+bj7/5EPyy4y5PfSCNLBMR4hppMYoyc+fL3jlfR2rn5numE/be/
6+Osgc6CCcBs2ciB8RUfiYAAG27garxB5Li5yC0ZTbxc7YJ4VxsmfPpcGBUw1u1I
+UQuCMVW8wt9MtHZPqqbj5v2TXLOekOeoJkn6sZak/t9191Og3TPfKF46XnKeCYo
7FI/jTfi6kGvbeOI5I5ekDA5vCxQm1pwrMWpfzX60xqtLnBw0icCYnp41vlX7iWW
4E2xwWPQEzxE36F5L7CP9k2czeEO4LzKUNhapAy/dA1+RCRyK1Qp47DW8Um66sGJ
vpKDLfCb4bhoeVW7BJJlgLzKW2YN0kTr1DMzgGhoYyJQqSjYdZ5PrLhscg/HAoWg
lPItM9scMHrDCRFj9UaId+SqyJI7X0uX7IQoyiqRclZ0DEXpK9cKnWapmHXevFZw
ueXxXtsgiz+hqNi6fd1Ls5YDkhpKffYfmlP1x+sFVNGKKWnjAgajqG5PTpaubUly
ff2V4eX74HkcPJ31ucLwMSqxoZ4bSLw7U9LX85xOWks8ePocdai+3Sji9RU6RUvc
42rsNaYIBe8f+RgtU/GcDbfF08kfVMskmjhawUJ00hvbvjMG9yaUa9OzS1BHWx4z
h23rgk2hgIqZetpKQ+6HREgytDSyDhfUR0KaP+yCexozoHd9HrJnlvGNDu0WPSSA
mx5tfIoRJEcQuGcIKddO1j6a2XdQLTnYSD37EAaSPrKPKd4MWqnqfB4psPeyCHrL
WXMVLa0GyBKNpjYSU6Q6cMKSKXi+KBjRslMotm92w/pYWTmy4pzuDoUOvl2SbSw4
TgqJECLSDOpLLpEHyLJR7ChU3S2MexP9eCm/X/5/lbOIRI5i0B6F0T81OnlHFkEc
+JO4ZCjUe5BKPSd7sEr6Lt13kweTBHKKVESgWMwi0CZsvzrhRWHDgnemFp47JWF8
+p7l2uT2w/BIzPuT33S3sdggSDmS0BEnpGbvJdFkjUW7Wp+W8qf8XoqV2Fce+37X
1csdEOSSssq3fbLUCYfM8gsFCz8phnvVrXp0hoYru6EnCgFr++ZwSEDf9I7qBcun
kqsgKkMU7xA40PKWeApyVTMixasQvr8PMaN4DxG+wKg0fnwjxo4bECdS0lCFSs+A
Ca/UcR6I8K1ZN2J0R1V7wZzx84iEiXx0uhiTSzwhHM/AK25E7CfFZzYtwveaGXnT
zbZVLSG4smOvn+PTtzIBfkH3EwpPQ+Vaoc9G2d6FYRbAWKfnfN5I87Y65ooCbXwk
wirM737rDGhEHflH54gI1lGQgsjZJEo1meynnpgffh93vayqfXjtwV+MoVch9VFh
KVvQkHTgoEhRoRd42cyl3hjmmlghR4ikBpspp9+/usXrEfznqm0zxsw3/V5d7jyA
GTE4AYOI+sJXKxqCsK1EL71oCpOkmfN7A/raI1Ygvxf5pUmuJKP6FSpg7SnyZiBc
LCGOKi7CgFcmnU+d8IG6DPvaMMY7JaOn4Rvdij4gEy3e1q/fnjZjcoIET4aa4S7m
wy3bkSha6J0p5Rrpfx2a/4S7iypna0KUOvD9OJQJjceTn0b6mVNFQyoQ/Ges0Pnc
Au2PVe2949rdsClOxlLIncNT888q+4JeWysOlFVEuVdAm++gcS5+9ItTp7lbqZ79
e5I0Zxr91285SjtISjIYW8aWVvYQk+lNX030H32fLx5cRMV83zp8VKRZIcBiv4mr
l+c3epIs+gMXG9y9UCpTpUA7hvS7mHORX0QKbjW6vXCYOmcwTt2fiGX7HjnRcjJa
lTDMFvye5pB6+tjF/Z5PXfFB6MWt/kp3wCK8FtlSuNjODNQXeSBzSXemCY6ZyCKn
oO3ZCorZJwtxIf7fthRSaE59FhFOFxQ6xHjpb889E8d+jET5vmMQ8rAkNqdet7qh
Umvpb6C9ad4OeZyDAq3xnIuay+dL7C5kAaJzFOZ6XMK0B9ZvJg/FfT23SnPMf4NH
Z1581fuVT2DZpuEgem4o7OgZUlc2CEJTQB8BPqDGJRIGQVZLQVOWKfeqAH+ONnOH
eXpqkEnXgwipIFLqbJJflQk0DA0tZb/W+7jw3VwCUAvfYQPr0OpP8AphXTo9qZk4
82hs1c2itJOnaFTnYulZuzzl2kYxALuFJDLh18NZCTFbKtrW5isUU2N7AHY3vKXR
bjRl2L826vwEb4kzdc+0ibaqESOVRkvEHlRHsXU6A3pcztINUwMUzfmNKLMPSmv4
sbxh6HXrSCadV7mwGlA9VQp6Mc3jcMgbZn4DoR/i9kr2L/kHeuWQIV20cOZH72Qj
7ngv3kgEOPhTf4omn2c6aTH6VOHxT20iMF+8dPd7dj+igYbroSMLuq3S4mAxa189
8Zxs7R9c7Yz59lDNBZ/3I2ef72WM78agAT/kTbsY/tfzorKZoAAO03iLka/kbJfM
KduBYsrhcohKhZFxNGd2gvpdnYpi3PsFB6GtVTJChSp/V2db5nqpfH0G5o8IKr1N
SQKsr9FDFgwujVSybf335miphPaTdCAinEONsZUbabzvyV5/tYcqCkMBRkXRbP6f
IE7kzkNnsHZm9wdH65/8Rmezq06FVQKkpbRlJ6jkU+fTj5CpdcnBiNj4QgdwDRur
D66AXKzRCJR+za+5EyI84/kZFZ67sJ9BMi9v0HXirB23vGUnNZnAawVmg7UjldXf
bvfQ2pyjDF9Qsr0nFzIv5fVm9uQeUt+DZe/vWwDTs+VC8523z7STYJH7a4u5VnAs
YgNDS1T9/xoapjPg3DNXntQ1BsTw82bMHzOo/uFpHTJaLqBuj7WChOEedFmB3zMe
PSX/9uL8kDHy5T8FfEyfPh+RABsaa6JkZjJ9Us/ChamKHi3KGn/HboXBqLDCj2dE
vo7PJrneHrCktG/IvPE0m85l+m5CxWhz81dX1qGKNthxb1/egvsjMV83mUycL/At
ZTiBXxEMcELya9QGFsQAoHXaTtDmMbbf4YXhcjwxeheh9KaLUmNQDcpjaMQ0zcdY
1sKor8ip6xZv5D4nHD40H+lBfQDc7FkpJhNcUVdNkPrrvuWQ/mOlvFPCauPul2Tc
Ucan1tEOraFcq6evQRzhbJloV6s+lZ9KTnYGvcBmwLqY6tvsT9zQ4ig/jGlAVJwO
P40puSDI8Sv6a6wgAJA2DdqU+EyCy+lkFltonSApr/Tl5GPcADeXdnSaC/pISYZu
P0VXHu3SgPUBnh4SxlQUhOrUjwOQSGrxgtaAzLq+Tu3fFzk+42L/mw+RMV1KGiNd
HK3oEgkOywOFca7YRNOGMpAGvf1TtTsi4UacKfJj47i0ByU+/qoAJ6RGwC1PYae+
tcwY4+Y4k80rj+fVD4/cZCdpXTq+1yp8smTGcBLF0zLbzH2AGy7oeSMzkuL7xh54
q7szwenNsKSLvAUpSYXPDsWRgicz2oPVJWsFdxgnMQf9fVZjscg0P7u26dy1Ob1J
Lp++UYjhJg2X47OeP/b7KsjZ4nbjsRbEuo2dtWPrt8klQ2PMsaF4PnYJ+gi/ERPi
Z+O3TOx8/oUR9m/QVBi2cHAQGGKmKSPN1PPpuU/Xt+LMC2QBAggThI1ifkVOoLKi
cGf4YaR/lABIAkq63aokMNZofZHTMiHl1SSPWm3q/F8O5VsblQIrr8GLiuPHrlqh
UyBN7P2pTjmYlFA1e69DCCSRq13gDOTnYuDuMUQysIdIr2T9B3EfI9kbalhaAOVb
YlGGdEY08f8BrCDSBEbiXRXYck/fY/COyp+0PFrsY3HqfprkIymdHxrLRXiKsJAq
fzB68OY2ogzJ4UxEXownfNKBmIty+cczk4U5JUM6fbzI3lRK7mesqMVA2Css6lmS
5wNML/xQwuLIzFKvFZm6rLCh0Sp4o4LYPPMIYHYO69OZIGAyefHcg+K1Xi6tSG+S
F1OGLy+J/auZPBBc153cnMe/Gz5iVlmBujn/kTagBWY/Mziw5k6/YiggHP7yt+KS
ghs7v2GIo5qVa/HiwWUCAl9BS88KXJuNwDtkUYQldZctLcVZJbpgG2bHq5LfxS/T
640bw4JvBcd5b8eJocFAGX5hOzH+BekHrc6sdyW319WiPtzrBqk3ig+0fEZRW+kr
L277Rc8np85CnXvlhYVS1MqoIlZ0qlJzOaBUi5WHAaPOqSbuVLbeBky7aKOW87D0
xzOzI2g4glVfBfWZ957m2YVeKIMDwpm67W23lmEK1Ql1XfYFb0i0qYEXnO0NCn4J
0HTURqkvl9bsKbsJN3fZhyh9a//87hDX3mFfa14UVEeepW3OVEfP9Qp3jThDIrE7
wMb96w/c/YsuKp2r2MeEAkkUisKKTkEvNvLMK+88f0gS9z65O1fF2nxxw5gbJIzx
2B1DJoO4yZFXkFGhuo1+EC6etwb0VpobzZ96kIMwhcCQLuQaaNGqIqQb9zp39dOT
bEKanqgk1kmkU5jOtW8LCDS1F84fOEwdUaQ4zaUYf3LlFR1oCOxhbq3Jsj77BzGY
Up9Ap4Wfdj5gZXd0gVNtbnFfB/b3WGEhFDt4UJO7qqevgMVE4u06/4shLreUjQi2
IT6Fn2pjjb3dota+gyYQN60jz1vEW0G2Dw6IBlNuM9NGIRG/mbLhWJa3mNCkm72w
aFZCNI/hFVyJYhmFMs939R/4hPNfoZd2sEq9J8RcAtiuY4PcMPqxR9MtyTLHuz0Z
+L8qTmVwyhHBc/H+UPCdyK5DBxsPwIFJcvx3eK039BF9TzV/HLTYTJ9c2tsTTdUt
gygugqLd48ZQXPXct8+GB4lzONmhN8yj44MZDpcPg5kiguCmZZW9a14sLIVyA3jP
8fLxpVJyNeXqfkFVoYN0wMj+jbQK2hl1dpCa9LKBs1IqNdMRs9FjJxGklZDMTL+k
orryP2Um+PNr/dStH2vWOrwckAOKjF0L9HT5IRvy8UC8J+tC0snFA62ygnQfGAnj
/MqoghU9aRY+q/OcJOYbVxzHrE0DNHzbOUzG9qfkP8eqzeLeqGMeJck2U3h73YtM
IDbeP1l7aVYYJZzTwsm+IANQj+DeMb15cKr70jyAISfEGQkpSwa7MCEYryiU6oPV
+NHQuANGNYsHc31sdUuuJ71zwHRL3IBpIg3iazUfDMo3vGiiKvevQuBLOWnlsRDy
KMJe3DdRLroJBTduGU5UzdZS/tjq1NBknsXrFA8ZuoliZiIAVTka02p96684b8VR
M8ooB7HPzGFTjWqXAJIpJ2sK0YkAlgKY7JU8WUdxW+AsE7rmkoz8O+gllWfrUu+c
3Ogm8N/4RsWHF6R4OwZa7WBVp732PQZdz+fMXxhh4XCYTxxISkwDhAYNtl3hiZku
IYYmtJHZnS9eaJECSWT8D+ufQDsxPZ4dQBeWByQRZhuG9G7+3awQQcKmRJSprafn
mL6BWp43FQ8hOSjmWlNAjO0Fog4j/7Q6xAHM6QfO4NiQSIFaKQObZaooVZKKAiQ1
yeQco+O82pUyTy2AOeprFD4jZBBWUUxojeUCLKmfChyVVHlsd/wBwsss6sO1VUth
6DtRE8LFrD7my0st632ZA+nMge5wQajFgZn04HVZ8VrtyioFxpSmRNraSCu0MYoH
hkizpXz7e0W2Jj1/hNKw5eQL+8UG4Fsn3TqYXXNUqcwSLm6OG4UkVPM5eZtQw4X+
r5WWAPZK1cm4Kfy3I9sU+ZACLzza1uvxqEBgQS1Ofzge8Ftis0jvBuOmKtxFm5Fq
F0+kXLlNgLLbh1xIwD13rPdcJSr5sqMNp8A4vxyjXfhqQinIH8IlmVoUh75jGz90
AD590MJrTbISkoOLhkkh+ldxCwhWKIU0ZAKYVzrdiakEV4eKPW5nlWL1PFuVw0VR
Yl4ZQmPcNIshZflMgvo6qUqO59zI+l+nfZTK/rj/xkk1iC8oBKxwpRQZ3vMheS7t
/16hPRhSll3dzMldrCuLPlCvP9J0l3FpcXtmMHaLwls+hiuYBumwj++oAFw37mQh
BgP7UHYYOKDpoqiV5NusyHTi7w9B+qCaSpycKK2LaSU+7HePaXGltWI89/ZI8Uct
DX9EVFrNkKsPHVPHpJvOk/IIFffiIhLVUWZVExRj7OgVdxoYctdbgklzRQqjGUBK
xWTQa2hj594ng1KRF+tmNM1q307q66gV8i2B/27mgmZ6ntXihsFgruwXx59dRziA
xA75FpfuW77DdojFfE++m/PQ/e5hUpkeIT+ALYjwB/RidxRfq17annz3h9tHSrFC
Di2ffWrq3e8Buct4lk1YrrkGWDtxS5BaXq+xSFAYMlc9YDzPLE48NAwb3aDJuwMX
UUAkP+fr0j2XWeMmL1CygpXg0/MT46bB97ZA+4fYsghv4WZa2VfPtpK7micobNAb
9kmk41lX4NKTfSrn84oz4p5eVQXZkL2WFmEWIf3KBg7SSiSP8W+uAc/ZUEe7Oi3N
g/WxmwGSfJIqr1duAxxC0H/7ofyM3HGc8ofOsOUgjgr6Dd0WDyZ10eSktmWRxSUP
LhaI/CtaSdzLB1Vd33Y4bU188//4ZKtd7l73VclrogpkI7LaB/pBsPErgpAfQDOb
k2opHBp+SAvMAHpWvFSnYPzOhoG9gWk+SS+qXT8/cIRoIYYVFXe+XJ/SFrWqODBW
yCrsdwsY+RovWPvHIZgW3bixLy2hSlslmllwZBTUbIVd2jr0UtQtDJMJ1g+zovse
1p7ztg69r2YlE6VGux/9UZcxltCUL96scYjA/0109qiYyR/ooyzzdmdGt14LPXod
NsdH8IvUi0FR6XJKMS/KBg6xuU0QuCnP5kLlFjN8eLFtkl9ccex9rosMsOlAonKb
HzvWWy6EYFs9/2OJji/L9zxRbnGZG3L6GdCciK2i1fJshHaQw+4WKd0pkbrN5COE
B97Z0lElU/Jl32seVjGL6MY6NJk8LJeG1qmZ+fASaTubXbNUUgc1zbebvuLnbrHM
fH7qy/ntxxFHFM15arK27fdchPnfugoKYHQz5UeH7nQ8HnkJKXGXFiviinT07hWO
C6Zf7ZqQ7GwXadcRTjMR5qMBs8T96I1I/0A5QHHaj5M9hhR7zuC6gM+bWn7KTcAc
kLS8lx/TaxrVgGAlQDisU+Ul+AJRzrqnDsry6VSTkKI98mUiltSgXr1np+/enVfl
IgPu8twWJKhNyaW34Q51en7QMwDMJSetGsPs6E+gOb0hjIDt9uqWJWarBzoRtwx+
ZLGFKKZBLZKN3pF7CE1IOm0/NIYTAVY5EUK2n1zrHIsy4SRsVi+l9J0Epy/BPC5k
r/UHOB+kqH07Po4ypvTZktsMLmGBI1PGOhstoHlVJLYBFj8t3pBlhwciS2nOlBlu
RDIS3d9MgaTC6MTfQ890wsJI1lok2I8s7L5qPd4miToiyB/N5ILbesBhmjvPf3jT
Wj1R6sBgtB88Trs0zo9lU6mMvx+Yksn2p7EvjldWye/UWmuhxIq4py84Cwqx1Fxd
x1J7TlwLIG7QShrqIUtxlNZOU1SA4ov5oDCG2IzZxFTuHfsX62K6n4TwWE+vUDqw
kgJarN/DBIqOcscY66LvaWzhDoss6UIvhMEdtLrhm70zswh0uJiVg4Hz6tO2W8Cl
m7dArOfLCMM2hj470jApOosbXA96jSQFZWLHwhivR2Zu/016MV6OpvEaEq6Rp0un
jPXlkTUE5nSQ3t1B8Nn5iv9d3ByagCnj+/tacOwDuZvLdOxM0ZYuAy84HRsWPPMx
mr3/4kX+yOt9uQbPgd9RTdaY0LOVyqWmH8usrNpIyc0IenKTCDCtlAeFQYy3mUku
4adQ3lKvkDb4NUxd4g8QV2s9RWlx95oBa7V1MKMzRRVzFPzB1A/GZIzzXKfzzFs1
u9Qeep7dqDxI4hasFnsIu8/22kxsQHwo9DYdgYVz+Rn9qSlBBH417vJ87NGpR5z9
2Bv48Ui++zCcgEDF6aTaBV0U5wdFfKYa+UbMR/AJM2jOmKFKYrKYmvRQqGwYfNOK
+iqKm/0zcfMIJ/cxVAKHgayLmRyEvCW0gn8rNWNTO6C6ApcvHkiltNzV/tbjZgvl
CkM1/l8DaxoIGA5RWPSjM99bjUA1ScSKdZ6PVczWONoLrBq+L31HOqq5upQ+pFaQ
Bi0jKTi3wXnlQIXmFKluU7cQ8Vy2fQaWPsIy0c11sCvGNt4YrKVdBrAx1rrrH4LH
VT4GRUUO0UB1T8VMlU5IiHfZGidDBg/MicS+HvCTS2huyX1R3BqbllHqycriOKaA
HgJ0JMmn7sVwBPXi5oqOAoNS7DuegLtgMcIinJMtDeRDGWCZs1Tb6QJjF5D3nkNf
VgiJAKcqtKcBEiNLqPJpYnOI86t753zjcNqGpaPKEH6b6pb7Lbp1BJv/YJkoZoPk
cDH1L6DyPgoYjNJDCGSVCPwTaHzPRpsS7gJXhbfGivluvKF3YHkVbMHP7H7TldES
QUbmwjPxrEnlA7qIl2IZSpUmY2HXbptM0Qy+R9MIO+6IrRoE3WwZxqn6K0Kv+mxi
ZIHVpxBpQjQ6Fe0BBxPwivyw5Bz6qhVLFuJLBaIdnjnJRs0TUxoOUXgG6YhHJx0q
VFuaw2NRBc/mfTRZpkD6zTVPv+e0vvzhAJCWW3tvNn440RDk6QWvb0f1MVQ8i2dD
H8BR83rxm/SZm4pSdFe86cOmDvf5SuVj+Lhp2ZGuckwcEebU8ROOvfnI6RtPVOFW
e8SjgGeKZ15hwlM6T19i4C+y92tI/OssREgAj5BtN368V/TKBnNeD76Ph7odhAhP
IUmNth1mxFvIOZ+ooCPAnHQ/6AleBQZjg0MGPxezeacHJxB+7htNFc5wUVGsAjws
FurPLQK+LQLrXrJVW5EtvHrr3Gf8DA7FRpTnyYPmAoJYeZr9IEtGnJVJ9oDGCDBH
Wz/Ne8q7YLBF8Qvmge5Yh6t0hu3/L5AaaQ7xF8ao6xi8kkel5sJVQ4M+ndS9tOxZ
8OHHZ7JSBG5uxYat3o/781OdlqFZh7VTh4v4tyM1YVn0HhdfRGPxqlDHhOhFhPKN
bttQZvP+ojkPHV6rNe7WFVCb5OdLxd3BNveCpVZVn2Z7t0bMzQ+WSKJiBykX2ktB
o3PxUjRChX+9rmLzN+5RvrES3k79BNeFn2gMgDjIQTGSWppbj+gLvVsO8mVMWLUs
1/xTM660ROVHu7NhDLwoxojX9vHcFNtGbWSXLeDgXkUOgLfmdmIz5QLNEpfaFqSe
Dm6y/2xQQL7SNd6+Yfdds6kR88tSZSwR0fPqCdueUR78DnxasgNco59v3CdQ/xm1
wZ/+hwJQrnytMmw0HZIDblNRA7F4SQ49CrJGVNsBwf1zdaeYIsWIJoyU3MA8J3PQ
TulK1oz54TiDaLtN4x095+gahBwS1cd7ZK2j2236qPotp1T3HpW7oh4Py0KSh873
3TY+0HdajW4nJotPFW/AnaVG7vj42pWodAwxcavA6Dmrn3LAD67uFnHI6GUsGQLg
TZSP99jdolKzKiwjT0lijG3jwJE77BNLj0W9XnmWZpsLgYyMcG6rhm6gEHy7zD15
POivcsqVxH0y6GzdjZPDPPEGnl1netgGDrsLr94EqY5CVJl6UruX/EZCWB7F1pLf
0Z2jpZYZHki6j1FSfqLyxSbZZMXx5RnGAc0rGaUEk8GdrWWobVgjsggFmTQACmUl
9CKoTF0V9m+6/AbZIVX7ptV/xth5vPiSFlMnygGH0nbdH2BJhaNBmaWC5aeLFocT
cujqr09M/uWcurzuaqKfhalekzy0FNUwlbBie8jK3ntVjeT2TgfiMUK1vm+Pr9cW
t/Ox43UhgXL488eAXs5msc4V7XIf99P4yDkdkBEpUgAprY6bb9ZciIOAUgiDKvHV
0p9QC4HkYpOcNGvrLSoGvUzo627yGsSuTZ752xT3bG9vh570hjZsI20K1ypONlxF
YIC5ElPWL86DVO57sJh2ds4zPdOsdBvGOgQ09cFqezV1aiiaKJQii+Qc8vDkVF2X
QDoYe6jGQ8FVUrfGKj6tKI9K34KBwsXzHZCCtxIF0aPmj2H11PJ70cPwEijpnVi7
xtwpO5tEyK/x0dwVk/Gs4yD/RY8HAs7g3RcZRH6GpMcrkxtk362mIL2vM7FNtHq9
WBfIcjmVp17STYhQtvUqdrC4GnHgMXABT8WYnhf45HJUWearCQ4PZhjsCxpn18uV
Z0YGSrDE+zuqoqGFMFJexHVSu/zBhKLBclW6g7ezB1EAjQ0/8lqJWhS9GCstahgz
awV+9H1uYqdDaqzjLSQrYmqU99r5drO/qNSb17flrUy8ZT9Kztrz1L5rgb1ULS1V
2PErBfqHsCMPjN20KqzZ4ScV/MAEGquX/WBuYXtr7HnYGk1B5naydF9ZLqrZxeER
NbvtkK65g1E/1r9aAprNN4+VgTlx1+B4o8croZ8CWQQhf251PjQU7buYWYV6/Wrt
5DoICPjW9FlnB3d9oLUjULyxsa25C/ZubtK+8EIPG402l9NPz5ETr1QwF7w4xPdM
hGUWTltQs3wiB0xG4fz4TDu95bP9iLrPWTh/HAO4c8nhQX0ekjxa5jgJBLaZDrlI
KrYauelGurMvJm5KoEtFBcYrxaSGvLArgv6KiROoeYcLkm98tDL8TzvQJLdxVUMN
QT21/XBKCL7vM3LXZAUxjDU3FG/pztdVT12q0lVCuiFn9CArOr2e9HsRsBLbCHl0
OfQ/hPzLCbpso0hIZjpg8/OgydQyJVW4v+Okwyj7Nv8Z5+2400oFC0LJOXHpHlAm
52B+cC7pahHUJ6EqOneOybH1vbs74NlN52FI5KN/twJyRawWaEdSfKhfkpVjIHMp
SZGSU/iImxj2j2W3sNcIlEuNWm6MYzLllPVbyK/l8Gs5s2qLniv++lHBcGBdh2kA
juBwrm8zpChN5qcV163obhKdN0G9EvKnwol8gmsSMzLMjIt4yesXFJhtPyf97Sj4
qyE6R9SaiTo983RGtytg9jb3T3Z9Svmgri6iE9qOusA1f12Y1munuorcagIdXCkw
Og0UPEAEfdiNMwqPkM40x7URa4EoKokgAHmNm6H1eSa+fz19jPmgdgtI4nmxuj2C
OOTrR4LzXnOZRv2r68N9RFdabhTH+cg72m8bSSxcvWOIeTeYcmU+e9wWBAgWVlNy
OhI37rX9O0g+vLuY1lUV8IFN7+iGj3aSARfSAEt+alt+jrS64hfer4ehnieFdIK8
+Cr0y/n9P8QZqk7q2cW1lc98u9zti7AwOqaz8RAIZTQYc+JRFZMO23hZ2hF0v7gi
n9R5qzzkvZsRMbf1MYQxzy1epOtM+mxZ5Qn9/1GQ8q/LXJZhwd4FW5Y3eDD34oPT
ghpKWFeBhvdB7ViUK77fDphkYjSrocWwJkGL5Sc6ATrvJDLwbdo4Khpvw+KzF0lJ
KQC9PP7/zENyI+YhIWQL10nQXUX8UV9yOOoQ6xmZv+8nEYf3odfQCggJfckkELzB
xa4iOtEyTsCLL5G6MbPowsfhinCaf+567qZQSMVnaMlhF5pNtrSv2A6OnbKOtL5u
Q711sy1KZ6owym3LJXB/qT+taAmeP3ioHkrKASjtje5eZJmf0vj2Jd95HOzpbKel
vG74ypWJXZVGLnv0F0nVw50RVjRnvMVAeU/uEzcW2QX9LVDLuxHJHsBOl2wbTYAr
jirC0tipDtjSwOIATAPxBDLkBPyjJTjo3F6Am/AWeluw6Nfl0iY79hR5SyYbreq7
PtYVuezVvFCCu+uZqApTkWtHUTjyFqeIQKVLqgfz+fKwPqx1pGSgRECMfB82ZsDi
ZlUc/msaSK2wEIIinTN5nMsawWYge7MPsarnMFU+GLCqfDD9rbV3h5YkcJjhUxKL
vd07D4uXZ0B5eUD1o2d4OQ==
`protect END_PROTECTED
