`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4ixgqcvJSBxYHekuQP6CAHi2bmX2Ir1DMHAcAvlwdSNlI2KsXkNXTmiZtuqepDk
e4ihm/rW9XWj8yPqe6TofkZ317PdsOsPK8pL6Mth2z0JdhhC+QJZnmgnaCX2RZOx
1pODxe+sw/b4gyJV7oaKBBRjx+vtuk0WhOR+SN2f5KH3CP7CHOzeX759i3RGEAId
Abm8bZ4wI6AW4/CthAX9XpThcR6doAcpApWlyHnWT6ashoKVguh+Z6tKpDtR09Hg
9R155KYnLRyEnZH8RdY32d9+6CtsJnjMP7jIuJPwjkeXFeO0twGgUgcbs14qyQVF
FcMeBjc0s9BRAKYv/ZbfSRm0ld7dccGfABnW52sqVt3dDUGfk3W6PhpN9Db6R5DN
CDImDP/vUr1mguvH2SsULj8aYsUqpYwGPkB+aMDc6Fz4i3O6DK0pb0Rd05u6deqz
HjUUWQObOSQO1agId0I+oKAPVITo3Ert7Uf5ScFmh+7+ghnm8YJhXq8yvjuYRDIw
qblxr97QVg+FsKofppasO6sqOxRDORDB4ueBK7ox1g7rvHgGhMfUsUqWwQV9LVYW
jOG5l2P4GPkPY1Xy4OgFlUkNSAmUctKYD1/Iaqfj2JenQu6qYvjI9kHaqdglQW1N
PacwpAOALpHOwUIkSK6q3AMIjXQ/KDVF9Gi0qXhbKmUEkNEAqYUQzkUTBNOcp/T6
aacMGc8/0P1fGmYg3MlntCWAr9e3eCRX2SVq1GPRonHaIi14hLF3MlheF445biLf
dvNNnMCULqoTTf1m1uUdGWqwkLfJU7EGxh+8f/UUH0VA05f0bHS0fqBrLlD49YrF
8IQeBbH/rO74iI5pKPFxgU4qWvCclEdpSXZpRcVG+D+eG/a88WOcLoT9gZBiJA68
7R6rMnQFJSYO9dW+AS+RqvJ86r9+qqn4vTBvDi7UkFGgg2ddtIH4XwM4hm8zHrWx
hsztzB30mriAsysDjpfv9iLhN3h7GxeDMGaJNRoO2A8ylGduoi2Z6m/CO2dfVTD+
b/3VpEgnN/lec24iapnbJ+qOg8psXRQFyjstAa7HblZQQeMGFuKkFlDdOxevcut7
QaF0ISOJYtEClLkj8Fpfy2egBv8dZPCkcyVvnZBxed6jXRURneGYSUUnzUEl0FCS
M0YusptP9S+OPG4hBAPwSQujoScS0UPV1hi+lC3ERvKHbStL7WxyfrQVjj4eQHDm
P3HzBhFqRggRVXua0uFpWGxcLFM2OVKreTYI5oI5hnE5vnGtIxoZp0LVP3F4eiVb
TGc+e49tJxAlF+Y8thR747i9FT940TkSiVUZOgOVssj6Xin5fEAI6MVE/tJNzHXs
70zWbaW4DuJER6eUBfbp+WzvglroeZYW8c7/+CsKuHu84JIUOVvkZGcD54XFhhlS
p5QNcpi87lzSR1eUf78obN90ojV3EjdxBrrZ1XeF5SNOL3psb1c5sl8oezQ0ptEJ
BupMAn7ebe2LW1WC9smeaxVaNGFj6mZtfOsN6nuVBiCa2QHDuBL12Ci7XOniZyd+
pUFWMpr9xROF3VP7P8lZaBVvtU8r920VfcO1/LTy/ucOzlHRJUphm4izoXzqlTzg
tWDI1Ac5yQlbgihbxeGxgbU3tefC6qHMPyVPn0fr/kz16uMrO7ioxpmb4hghypik
9ecoR4roaR+mJdDTOTeO93gKPhqH0OlkIk0OakICBMfVUgmuFgKmJQm1Tau7hm8B
XHZoTmvZwDzYvNSPCoVYmjPF9ZZrhnlO8sV9jCzbhxpPfbI1bIYdhXfWF096Z49g
81aaF7lla3Cs7EzP5jNSRlvNCdLSTqbiPdjXj1eFz9PTximE4NJEtgby94Beko57
n4Ol41Pms0WpjEE1Ssh3MPcw93k+Y5y/+Crhse374bBADGaE8cPKCNZG/QYsWQQ5
X8rXanFEIfJqpcf3vYBMs8b9P2uilvRXE9x7UpudISbZOxCur6WHlBr9iGVMOder
MOIsjxXPokQRy6trs7ZvzLGHC42sr5NYHvo7VaPCWMeuMtZ7tqCxERBqKZ0F8BmW
67oTd1djgT6NcChPFsp+ZwZdg3b2rD2efqddzUn6wmw1Q+eNNaLSXAhiXIfvlPgc
XjJo7aY6/gFeZ2FFQygvZkQPgPmTB7Y4Ti5cXTrgKg37j7btoJCLRTMJGYb8R+4F
rBvflRj5/Tn1252zkn8NVREOxGDRbQu8VVfHxoXgbjan3uJdrY47XpO/gpz65/HD
gp0UCVG4lGSEVTnvmlKZj+/RmBLq6+03Y/8oAMWsfh2G1JypffkxvpYZeR4J6egn
qvTd0eKPSE1NsyvI4Awrlc250dXqxcWHn7FwXk5eqeHJYKyYFJsQgwoD+EzGU2qw
XXyA0GT+6/2PF3V1LpAgJwMznYdqfG90eqfy//NOZf5eafxLmA/BeKCMNv+CfN4j
BH1vtG3WzIU1ma+0SpsXO3DqLEx3FOSxe2oeTeV0vjU/tC1us4g7Tq5p0OxZyuSP
92W8LRiaJSK6NMbtbRp4Xfwp8nNr8Ig6pAm89ywOXvgnap3yMaOPVFabYOYac455
HQiNcyY+Bcw93683fbyNcwa9jozavwWg9EVKBccApTqmsdlNqLpa8fzkZYfkz30s
Kf3gUWyrwIb1vrItymKa4JpjlLMyD5tPWYQheEOG+VwYUo8wlUaeNZYpTdVdp3KE
xPfjQoQr7bJukmOSgJmASs2JKhetIMjQoYnwGX8szj9LjuGhTs8dLi+Y/AXHLSoB
1HugJOkWhOiQ7OR5A2+fQRnK5V42qEBKUU8yF+0rljwmR1mdK4Tsj3A3pHCW37pR
qDZVbQ/Y1kJKAh0Z+frPm+nW+RkflqASKXxwXJGwBOvPjog+7DdUEQHVemECa0OK
wYHN1+CKka5vfIDdDT6YNh4TbvvCxxYIPP1j2RHImTHS8m5pVb2pUHxaW7C2Fb9g
FLDd7pxF5IwbYiYtgWJ8wt4gAu88U1c9FUB0e1PLGqASfP0Dhj4Ig7OndfVEhWtm
q6Sg/54WKO/5OYrRfd8mz7o6cAWsixcjlBcz/FX9J3pm4V+F7p+1NvjPY1RCRlQz
BNEY+rZRDmPDk9wpXWyJj08bkxJzQxmf13fwR0GMnZbdAe1F7UPfpZCxfjDxGeU5
ThtTGubztMoxADofKZTsboWRZvlAYGp9HYrnqbloFlSWV0GZJHeRD8b78r+1OfMa
k851U5oKeZIKfxlnss9H9h4eiuR1UtqqEgHP1Yiq7tY5XmPxq++c2M8WpRF3cvm4
CQ34A4izpuC5/nL/GE9K94xCyurNJUKFjyAxILI0bwdxMkWlfwK4YWd+Fxovj2BV
eu6WYRadUherW5mg+DsFNXHE/djCUmvZJdh5aF2pquqbG87qv4wuSv/Yir4vit/4
WdpImGRLxe8Jms5hIzltYDr53GGpNn5E+/kOXxBExCN4IISqEzKZ/NYycZGyW8bV
bMPdSXn8DA/+xWn+px5B7bWobpbxNtcfLjiXEvTrqZcoTYB1ETjhR1yTZqdMCn0s
EnePTl3aPyfU79luKC01wkAVo4CvjkdXVYiU3su35b9CluId+F9zftrELySf/ZfK
htEKpqCGigPvCtzJQETiJLNhuA5FHG1DvoNP8TLyOpk7hPmYbWHL6dA5X0g79rZa
ARNAVXcoFL6Pz34Tsc9PjBge0C23if0Mb0ZFak2DfNKM6OK4QBJElgLXOUo/GJLl
iUAmhJqA4qLI9bwyLzsyp2ip7CgjOqGxY8CKguZ9Kn1qYMT2E1UZJJpPi/vQhOSM
J+Cdo8IcAIxb2w/4nTKFS2KRfZp0mMexEPMZ8xpfzjj0HrSsC5jXH3qFy3+uiQ/l
ckyboPnf/kQMqNNMrQY9Yw6HP6a+1rSxWzVsT8SF2W+x1IFCpcx9t5e/6Qag4Rs2
ZF3JLSFYJRsvCQE5+oY3UrDBEWBAw1dEKglxrb2U3voi/01dXnjAYuAc1PFg4jqq
uFX3UK3y83MhYy44CXHlUQgWA60D/LnVHoQedSD2agOigeVHk4s3QhWlT9hEAvRt
xmSLZ6l2UWL1CjUsgQ5UJg22wo/NgPvrExTjEDluZ/UTzAY5PnrqP3Fj/zJHbahh
qy3jHQupMjfxx53uY2WzZPcNnkm42Whxingxdlx2PKGV2Hxk1n5NunwhoVd6BT+Q
qDI3BCh/I8IfJhyMEGkNE1UUNXekKuoU1Gru8kmrmI7bSuZptQA0Kek1z5ibAOls
eFMt9gTIEy188mtvewcK69inTZkUDzwgu4eVuXVouF4tl1nEeMaAcnPcluvhatyp
66QHbPCnpF3ZCByFYtIurypHiqUn7LtDCzqYjSZ6ZWhnxUP2bE2K8VICEdhGopwh
tidHYfDFD79g1gbvzEfwxojGVbAhfqXdSbYvBX47Jkwo/ZXQ8OTAYqTx0l7ywvZf
wxt80s1bHAxW888VYhQjH7m9i1RTj8/YZVhivi7H0+5ScdF4j5PFeCCFH69yVbBl
`protect END_PROTECTED
