`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bdr4Bg5KUZt4OglrgaxfntePEAN1RMMNrHn+fykbCPpBC7nSDwcqAVtFHge74aoD
AgyctrpfkgnS5Kb6Rc57sMjZtDk/DZWK87O/hUR7EXiwfGbwY6Qu2SXK/okWqPPM
LNb90iIvlioNSW4FyLefGAYGrXFcNZh2dJmklibIAmg0p+fqAnouB5IUUijfEF8b
q4uSHk6OT/BUs3+CA37k0fHiwhQzJmdSr4rjiQvZ1WgOX11VtQse/TyCX2GTlbRS
RwGNF7PA14JewSoiWRZvRsQ5LcuiaLHk0t539pFPP9Ji0OCDCWXBHHFbnkhsK0o4
DNvF6ZwJ+deb2FJYLQx6dS6NfxucVFmrkuL1eEWHobP9Lb1PZ2wfjWPrH5o5dGbs
uORZwWGhOjhi/pskBwYNfwT0z9Cl/3mGItuC1PiseHDxzdBjN8bOyIPBhDzq2Lsh
i/0j+I22yqJDx2+8zRsGrllf87abrwtFpndPzfShTySgsuuT1c5gKdG98USJRXQC
3aRqTMX0VClP8pJhDhuw1K5LnjCGlDmwUI3DMbvA6edUnuGr3V72vfq03pcatIEs
0s3Mm7+8rkYDNSXdYMdWQI2yw6vq0U+P2t4AoBk5nnnFF22QeWwbybvRjJxIsByl
hbhh7KXrkMYTq2NbViuXxF8AcVYbRCyIkel+lgw3nBW+8VAFkO+/Qalw75yQr8/S
XEhzXgkAL4jjFiF4uJYWhhoO17TTbukbZCsDjYsQrakykEGZ9syhw0UIOM24zyjJ
jW6Ci4oJPkWZZ5mRdgvIuPVAK4gvRI8X7Xac57XSTG+1iCx0/HUxzB04YpoELOmo
BCd/7pHIUwu9k5M206HsAKYZDZg9c0wN0UXF6ZnkFLH0eEvngbNHdgA8i0u+T/EZ
1fNPOTJ4znBJqVARYp4biLB+B6ew1UsPVZOtIvhpUXnLvR4Z84G0jfk175H0QaiB
uAidortYJ/eF+fzUGSKlqySTWYliHPa+2MiGlWM0BD+Y6qZuup7XiBdJjTutisHs
+HF+sWy6IpmLd6CxfoC4dWneNLe1Rfp+9MzwobsK48JkxW+al/kcpAYatwyo+tNQ
3atOkB+IifXmLgD8FcmW8GnZEh6F4x4RxNI2Kpm3mgMdvl5gLpk63tmAm82X2vAz
OjrTzYoLLm59kafMnmIm807FT+8tcC/Wtd3CPEmwc/es6OfEcSGOTpWLj6qGDXkX
Atisl07012QqV1SsmGUVrOtOIiSWVxonE5N6xXMjKhSEkvKBXuwQu2fIm9YqvM6k
P1Ynhm2hn6ethnpgvsqdwSCQZOMrp933kBWJvo/7EbpytjNSR9iMiGUEIQJT7UKi
NP/I8MkZaHSjWvR9FYoTdyXBips7QDk1PIgB5/vthks+pOx3+WmxUT6RJc24nvw0
76ddrNqJKL67c/El2ogLzqCFTwMk830FdtNkXwI7+ftIo3Q5tf4L5viCS2Ubqaer
X5rI6lVjPWD1Wpd/FXU2NI5MfHTQv2jk65v8kGb/LfXogk1qXdUoSQoRDUjNGbVI
GhI9eUzLohDlkCfBAq/Mo+59+56ai4V1lmiobixWKt2vdx2ey3Gjwvun/w1uxaSH
WaH5XdJS/6Z6A6RyWwa31jGt/uY6Q+SU5aCPqFoav9ILK9T4oV1Ki8p/1wu8mJWB
sMrxnM/xv1piTWpiXBz0wosQ+QvSaMBJ/czdNb+TPq1F3/lKc2+6VTnb1SuXShOV
L6f+SDYJjZjzd0zOlvFkjzw9RK76uvEQXjpVMDp43KKGRNBCqzz0FZOz6ZaxF9vs
xW8KvjbSfvbH0syNPK3rzQmfaiqxU1XfTVgG0u5pcZPLiAXk+8lROiBArFivBvvR
`protect END_PROTECTED
