`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qHd45h+QYsb3axtsuQjlK5LQMSny1IoxJBdR8M/3AI7Dc01giFjhW39sXEfxImy
op2f9bdBEo/QzY4JcW3kuL5myUJQkLFPXyepRDrTa19Ar83BOBiChBDE3OPheGE7
KGi4CbaTxACunz+WDMLwMuZ/HBjHuhpL3TXjva5PG1qjqNqUMjENWS6TEDAHNrMH
b6hipwt+c0TdwcTmD/ZMl3iH8RYnh3TRRzx2atKTq0yTgAtMMARBjXWxL8blHzw0
zfLmsH00Mou1XJUHcSbTE3ncVtAdXu6ML6AFF68jOfkowplO/RUcF6K2B4Xrl217
nRHoHiSjIRBHt7dnCV7QJcKenBX6cglWbq4C2NYupnV+jq50KGJJ66Zf1zsinpmS
dinkdde2OvvHRQR29PGg7zViFj6qwmuijwuj4AtdsqLkXB4PMnbxisJSfb7sdVSH
m7Dr1rSR0kxg1Wv+kTWEpwnjcncMyJy/ek3ryyEaDo7/m6KhACCXcbyQVf86kKNs
rf7GDzHrRezGfqpxRWK49GMt1rjQ2ZwYlcDdUX9XBynbKbZQym6bYkI67GFfMmSD
qs4iTh8KwMi1VLqrt5zPMXljkDH9ntMCF8E0BQUgnzCPCS3LkwP/8uabEXlCwrgR
H5haliq5ps6XL/r1qMKki3cDXulmYwqQ1A3cKpTBrB9IDk/6TOAfCznr9Ug1oTuk
WQeLcGXRNQ+sr4B147t2j6kzo5HD1HKRy9UB2GX1ummqV8S6gWbYyr0Er6hWiDv+
4m7ptYvCF7UAWCxsPilUiJTOg0G51VQ2Os2/zzQycQaqEcpBPhtMt4PULotMOUPA
Ycw38f6klBTtIWfSoZZhtckFGS27YrDb949iRGytM7nvS6sfzSxBTs155eJmzkmp
/ArrM5WU6gpsspI8PIjKYMyaGBNsqYyUQzSyyu4/bG9QWyfNh124JvyjN+TcRuDN
WkZqksTbvNre8deyHbdGnObDQ+1uoX+eXl//rQ1qJNc49CS9N0apNoA5yyuCknL6
`protect END_PROTECTED
