`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZ+QWlnfS5qnGHVlYxrnZ55vKme2cJv8bjluomA25T6h9o4qgDwQBKZTyAOp4e07
Y2gk0YH2y5Qa+ZpvCB0YaxjAhm9l0s8XjXYkDpanUu7oOydmER1FRCYfFvqwXTlo
SAJo8glxFyEp9MT1yjlFG7PJF90Mu2RSoSz70KfrT5+T7vEMT0jcadf5Kl4Y9v2O
UGjJSWvU+1yJCYDkiFDL4t2aKZU+0x73LFCnpT1YNitQyvt+Gc0hogJ1ktOtMh/R
mArK83toC9QsHXHQHjQiyLueNxxsK/PlvFmzLDfaW4k9Yx39qNqGC4wWMzgoUb4Y
H4C3WvomTqdbtS/cedXtVxwAQle7Z6nBT/SmKzvWTXKfetSbIn3ECm3LK1ufi2pF
aYHRWxn1vca9efcoNWSpSaRHURbxb38Ol1TrR8V0ej0jhmNMsKWD642hFIlrCXjm
OAk/JTXxsQISe8PDqwoWwqwl/GklEdtye+kYtAv1B4903LSQo8iJHjkLjEMSOQWL
ywCxKGRkuA1DKYAbOrqA+Vj08cYpHG7Zk+cPepouB5TPl0B4gLJpyAcI61kKqaxi
x9L68+5t8sMNaUINUZ7sC4KqX3KO9CbSfvH8flxRpv+h69ej52K7iBOMt9peTgEX
4OvBnMhG/CVviCBKgnT5B05ic4o4/0Y6nxaflMSS5RmvQ6KR5xCh695fo/7+XfVD
z+UYDtX/gtBbmPrfg2sniYiFsUtrDQfU1APXc3/b4m891XcE0LXceZfNCOw1NQDN
K1TpL3Z3x3ijXeIa4P/H56Frdtvth1nFUuuOJ0zbCCSZDRk8xm5zUoBjRZUMOreH
i7SGoT73hV1xM9bVfVf5YecxL4BnF4ETjCOXr0Ljpo39uIiJF2uI20V6L36vJ1Mp
AG6idVNvWkePli/cah8ar7FKyhvRggMfiCwnF0lHdzqoJ+7Stt2PdTEO8tMV9lnf
rp1TYyDeIxn3yqZek9C0+8NRWvV/b34w/CM9jxatZQt6IqqV1Nfa5udhcOKjWj5h
qntzZoLe9WmnZ8m/iuV+/4FY8pMPHI07HcpLaCnpE/twYHpyTuRgAHpAe+BcZSpv
YYy1v2ps+ewNA05fSsEeTaqrfyouesjcVBJnVi6IErzvOdiysNw/ZgtpZgUtZZlc
0/dYbFO0hV3ETNKnKCZ0tUOZt+BTURZGYb/kmTo+8/LGqG1TlDl75G0LS+BNtGpz
J8a18tLwMiHKw6DJZZ69ZgjFyJ47WPGU1MhyJOxYkgj4NSfJ8brCcptzjZRvGQv8
F6r40b1p0/QQdjBToZRPpMj9naYOJF37JcQd6NQzAcN5XaTLQWww56QgsbUAhpR5
XW6CoOgDzUeN23owhGCoNKbmtclVKne0yaisi+6hLdiUhrpGgcKLhrW9wvrdJVj0
fnhBCGyjSRsvVDEHTF0jhOyhQG4R/p3oiZCM1siW+GOxEerN+0JpaHtsNAYHVg23
P0M6cepBZM9k8KVsGEBZ2H/T79Inq+Bd6hCSMSjHev4cgbgPNiNSGhY1QlUcWnaa
xsZHN/SgHgJ0S/A56qtSLOgZVmUwMeRKqrNkh9fZpMGTCoF8ph/P7AO9QK8SLdLL
iRScZN3NVb8Amqjq/LYHHq7TOxU+V47JfzTz0KNMA+E=
`protect END_PROTECTED
