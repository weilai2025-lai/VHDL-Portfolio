`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipXr6uiKPvYwxpCdl1/MNrf2nsPDPKz94852Qk75Qc+hBcN/PDJltd7UHXVb1uCp
sHnz6ii1VTaEqpSqMxJWES13XvmiDaIrseKQ8n417lkmOJ+ZJmK8k+BdDbyXDHxl
8uEryQLexGRSnlSJLuhCeMqNzNqUHfUVOaUor2Fg5Bku08VEU6aKdVZABQS7gPci
e6VZh+ZFBFimzcaEne7uHR26CihWpO/VdMLl8By1XlcnaAiSDfM9DWr6NesIHZgP
yMiTTHBvOd1groJu/jFDD79zlN3YGJTeyMopsxT+CQRuuTpkQPt5wAvfRPou8v6C
KPNFG35aZxzq6lKb1T2+erm5r538PZ6t6bsQPrpC+RC+JjKyboxX939ZiyYil57u
LXubUn6hPb9k91svV0PE8ltjJEA6FiW4ywStxbzL78wAPuCpjtfLYQa2IV5dcNnd
kenZP7dWbc1Qkoy9Epr/nXumpF+TBDbPm803C30VdctEDWg18hs/DvfW/kYygYlO
i+dawkIh9ItqBIgyzV2OIZuPdgBR8bze7ULJrlbf7fzx96tZw9Xr4e0rRjVP4pqx
pklfuU6PMJae2tyF4tWUZfMRfC7HsdhWCVPxp8dlVY878nUtqHXn3orV0E93KoL5
oy8lSp3tT8nG/QqFIWbFFy5KKAx2lg6hnD9hfvioLH6/2X8xXKCYPpF8XsEbLo33
W/5o8Dmom694aYGybXabIDrjnyRx9XoznP9YF4nqFJBC3miTkLo4wuFdfdnbJkzx
s6OCdTI2FXL65KUH1IAm80dT5QsCRRwkmh/fAhZ59T4K4jTvP4A2Uw+sbm6LwVVc
4m5k1JNIreU6McF8AA/nkdql+2kxRAPPFTPVp1A9DDcjnoZZFjhs9F/snNNu1BrM
H7A8gfKmhEcSHR/Cp1uA7WiGoxa95IfKGL2mfpowRDI3eRXhb1VWKxwOuqBHjwSH
jamM/fzo33hRi+Y/DtQ8l5mFuwieayfbXE/vqCVDCstTlI6rUcv5bIJ2IAcfBbFV
CmgQuULYpWBqP/nv2fqq3P5WGEtB6U4+DIpzGDHUS8Vw1opO6p8WOz7WlXLqm4Kg
daNQ8fujohg+U7VqPEoDWMBBlpoWGwHZrT6Cqot6OfJSOS7ju3S7habIKdG8Qshf
J/cc1IagsE+q8R1ZSrNoIQ==
`protect END_PROTECTED
