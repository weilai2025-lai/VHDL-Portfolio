`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gGSJsM2BotTQ39BquTkN89NQYzJxq9v6E7Znnj0pnPLVywFWlWfqpOo2FYr0CdJT
P73+aq81OwppTI8IjnXJ/sSRKhx3/+U6VDrKAMik1J4VLP9OgjMuhuawSvR30d7Y
U9Yn2J6G1zIWUtycW40BRVpw2eoBwcOd4UyoPdEebzemPVFQq6YWiR32SlnKT1o3
t0nCQuH/y8V1a3iJnijbtNBn2vrceAEv7UF03WENXdE6iJlXzgTasj3tEBub8irn
szS39ZSevHZtIBIyygHbJ2l+CAfVaYtd8AT1ehChbZZtgLcSrb5PZm44/nZAnBI2
dtE5aKEL/FWNkauZ7e+0ND6jqo5dj80IHx7oVOYYcbPF0Bzgrlb7LcNoGdM7ksB0
mHYNzGKqOUTo0HlKXyR2tfCIqHZIM9eXoiCBKJd/UnQ2IHFbmBH9aSt7mkf+rGNc
7Hr0DgFWNTXAVS0qw4s86+Buac41y3K2jd6ZtliG0vghuYy4tyuGVlc6Gm55OEQV
I1Sx/UvMpW7cs5OAQGaNGZ2DhfGx6rGWGmVO8TdtxxN1URIGCsXm81xdK2uTC5Rg
fyQTL3RUclswoE5e70dJImnhZFbg00nc0QefMkIyAEgJp6WkGK/12rqbJIK09pn/
NNp5aqVC+lzwjPXF0XAOfPajkE5YuQ/jAmckG4Doj1kwpCgEL9X/aDq9JhOTP0UT
0x54b89OvNmvSfQMq5pO1wIkHWnyRl2TbJF14LB03Fpi2jRDQMUHNSZPe6KO23A7
rThWN0W2OBpcYaMTaEdS55Bm+DYH3XxGoU0Xd30SAcBobwSKCELM1CFKWlffpbKJ
7liSQX6GNVNUdif05qbgpMxoh734+4J0Asc2iKbTqDSlaobcz+cdboRQ50WzkuhZ
KFXzdyPQ2NR9wmF+24WoKGhkuAsAo6C9BoJB9b9KBkp+zqimhiXWCGoUSHUBLcwE
rHTKrh/MmPNMq/MdD2JyYiFfCn/4ptrunf3YqHa76x6bDFNfdYJv4EUOGYmJ085W
Wu0V6jNDAKpubwuU9OeHubD19DNXk4ny7UOdvU1rjUVrJ8iolEiqsJYsYhUdX/cL
QJakTliHIqnp6yCLl/JmU3LE6irWkcHHi3vMbU1d97MccRXTP53dnXMt1uzA6B87
hZKxpNW2N3jfjpw3b484uLnnoxNsUOHZ4KzTPSoNKBPueOAedkdi7U+EBlw3iZXJ
SObB5aZHPrb9lar2nSSzxiYofz2DfkgTf4wFxO2EqSkA/4o08jkPq1GDDsZvnA1/
9URv3j5fXae0IiDMDJsQ2cXaJ+nX6Cprt3cN4qwAfpQAoTgDsFUTNyh3ZsTi4CQQ
0lkg8n5SuBKhQaXMf1bEOzFGltHgL+mLCzhMF/VUreMAkO1z2THsSsOI5+KDCz20
hyz+IneC3jxg3TdZDbQECFATLtWBO/++mkwabxcH/eZrDkpjxv/EbKj4+MZs+o+J
6fLqyiWSaeB1chd6ReDfJMOg/ve8aF/7gGhJfRUg3VRHKvvpzExrjzhB7eTNP9QU
RoaL4WdKVOtTwVi0M1pHeg==
`protect END_PROTECTED
