`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fk+PhKK2dhHzYZTue1ORc95AkuR77kD3gWbltRQVyWrxM77ExT2Jy+fvA5kJmxH
7XR8BO+bEvPib5s8uATITZN+BAOlewXpsFauXqErBYc0NgGWAq7WWCjCVaOaK5PJ
Q2tqRP99rFyrLDuiw+NbFOsYOw28VgnFaZf50jWnGxMRObG//yj/EtK7Gd11mrB3
FAIy9bBE+ki7ShtCRPkmblxnpBo0GWVJHYcST7co4kveyGGRJ409GMEnTsv4VcNp
TyBBgX7dL1h+73NyRQQo5R4743Hc4DOhrvuOPAma5ipIjAeNl2/4r7h9VFbCHmte
V0bMGK6YIYVFse109/qTMQGcLdOtENYM1xaftrcc1XXzHFlI/nk+jKAB5uK/Da5n
+XvgG1D662tvYvgQuDH+wih8R3NkNcYODSwi2VbYwUQHPJa9xEyfb6TTYY/HgsUZ
k1xviVPGlGaw3XiW4rmMsDmXsAUtQsXRgrAUXRfi+8G0VtsU2QvfHqKqR7q5cAKB
UnXlZxptHgFLEaX6BBWvNawUz4hAl7+SvPyzzN3Y6Y4w48/vQivnhKCJrGAg0vUH
2Gf2S18SH5You22gvefIZhDW8hOmpaOaZxgsGVkcvWAU8iK/xICNP7P8jHjim8BZ
LF7R9HNhtGFVXj4rkA0o/3P+dV7T7oxd8e+dIFRr8tURWzDX7t8EfuYgxEqixMO9
hxAberes38KGactQDMez/lPASEMxZGs3wnR40DDDt3GbNTCcNqO5oqYHENV8KsB1
teTzCKB82IHzzPB6+pyex6Co+GnislMCG/ViZpM5jVJOFRmx81P32pVJ79f+cldx
kYLB8oDRFDMMma97w7wuamBGCpIZIOnPxKEJumBUIh+yHYbBCAEnp+jpTEXgv4D2
IAK2YsQnouO4W475NQaxDeXO8iyQDCh0dTxyDV8WX28jui0y09cGMe1epsIADGQN
y1dHl9xphqF2H3//q0IrTu4liIL/Ua6GCo1qeRBY7WKl2R9l1kG4UDEN8GoAOwvF
zvJVTAzk6JWmDs+p7qy7PGikZ3M7J7kV/8IGaC13ZLoFu8YDrs7BwLSDKzYj/UpL
tqNspuf2s/nT1mJXoNX3Y1L2ASUTLErgdoZr/AzTgJFufAYtTyAet0YEAsu5WI4x
nrteZ9t/5QgQAjhX2sh8JapcSExuwqbOMrM93vcNS1Xz3hojh+s+qOsLoWkuq687
5xmtw7gz/bAlK5FdXy6pJK6RldGZnozVtrsANUFFmyaYpsWM80f6rUUT3ShhxJFq
Rq68tDCXsM+KXS6rDHgAiP+P/2Fzz9eQC1i9NmclvLXYdChByZHvh5/TxMY4rzzx
zGosDokHdC9DHa4A6Ovyj6tdKzxn8nESzK8SouUJOxK/sZtRLfxy4/o8GuAC7PNO
k9CJlFrBzYzsmrbBGKHZsSBKOY6wrkQMQneEl/N5otkXUC6cQuOEl8qoXANUlQLn
5+rRphS023TSml4vYyy/xdlcE378BPMdUcR0FxL/5nxYb0wM+weaJumQ6mfRkkhN
YxEwK4xMwBUV4WQGDCjVyA==
`protect END_PROTECTED
