`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcSZUIEWsCFbtED4gQeSpjqcP9FXTuVINGOVa3wUnMtweInDTthUox0+Q9/OrJhb
I8q3mHcle2LWibOKYX4CT0BbF0hS3mDLCJCh3pavea5LdZB883VhGq1lcKvuCxa2
ttNa5ml/dj0yR0TNuI0CzoZty/3odn423DY10cH4k0NZOdqMFALKvl9N/6oVJOC7
IYDzRJSDHQywNNgVfkLPbr18d36622r36U8DRvMJN4NNMWbBC8BSwh2+ZX+KWuO9
5ovLvy9ERsNffoQZX0HY5uoXLFfG0oHYFQjkfYzXBZWhDt4TlIVBu5hLD9HAYIRo
m/ytqtpSSzqdJM+z2scCUyaiExl0OYHgsgzo9kdO7RtnkoXRaXoyvVmdaJ73AjGS
7kHmTYkYyJvUNetK0S9DtOyFv/4KTHNr53JV3Gi3LIfrJW4SSfRgF3eauKYrkI+G
kr82QyHWgiK+O75XjTzD/uDv+ApK7U78yhxSLFXh9mjRL2gOjeYVCfXSEMqSZvEk
D58wPWyW9/K/lc14Fzbx+Ov0rpcQ3Z7FyszvtoO4y/++arvNk6ZIRUiyhJrRnJzx
YO41pttpgQ4ZdMk5igjsrv1oqu/obkbtRvHY3wooofztAWnbG3+JGK2K6RkQizAC
N3WUIekjGECc7kPftCJus1KWMRojBTa6Jgff/m6LqIO/B/zboz5QS6RiNgustCaE
DxlMcUebEZXtbUdlFQeXs+KItxcEP1a23SYy4gSiKBVwpCMtgnWG4Fa/JQxFBqUG
JR5y4eGB6VPb+/Vwk0dZw2W4M2m811zFBixrh5wVmrc+lqruMjJXDV8NRLrFL0EI
fUekNKJoHtvTpojh+owO+HfI3D4SC3JnWwEFe8Y02tLSVr9dSww+bsVVjtmCznW6
9jHARCZjBwV3g9NqBqwyrX+dHsE1zF/6zX78h9u2o6by+vKtAbLqPoxLtd9bwbsI
4hr4Ll/XM4mlW9NLeHEnHiy6pxuEZj3y+wRkfbq8sYwhY9ro4rTSQbwtBrKVTMiq
36WYBQl2e5LhBdj5YBg6NQdxb2fnV4vYR0VX58DQC9xbO17reW4w1sy5CdV0Y1q3
nGABBmFNK9f47P+6+xK7EXJlV7tgyaz2KwFhtFMWms51oE/5HZQs1c4QQZ0/H/n8
/ggTZsEV7YOQEyB0SSjUf857X9wnzbc1Rac8/kNQIzClh71+kMSViqWBFM8DGL9j
vGlzl+IpndQD3hUPt/BccpNY3r1sWvb2PoCmowWnrkJDb4zxMnCzAD0kNfc9Nd7x
v84V9JuHzh6EZSyerhKNR19mHDV/7wacznfTqx7bgWBOktG+6byfeGBB7r1vW1AF
HhUTnZtljgT+kYR3KVA0I0RTIqNYwUavCOB6o0MWNeIslQCfMR6lsABZD7l1YWqe
Oi/rf2cILosheIaZtxPOjVFmazz0UW2/EbbtE9PsQ/53+NAVfeL/PJfz6VROcNFe
o0mwe7iMXkkjLm0Lgw1a+09MYDEjBsWqRC70xNM9daJ7di9AI4yEdCVa+TwsNS0O
bdZsX+XhIKaRbtQYUn+gKKdFtx+5rzWv1lsbzdbZBNYKSNUHwXs8VAqHkiBqoRlQ
bWKqBGGmtwxnCwbM3Nk8Wa16d2tmnd+SRzoYSrapcyFtBBzOtzPae9Rym6Na73uK
zs5OWxzDrLila3LKreGwbzpAFq9lJ+oKJ4wibHlLq/KZPnHaOTbRdARg/Y1EzlMj
eGXCVRLmVjbIN34aFKsHKlqtMALCx3cO9C7HtHdJtzsrBEx6A6BDZnCcnDm3PpA0
cMPn9dPUE4PZk4gsohZsu/82kCfT1R5J8USm9HQtPcuvxEULEKf9YolfvSKEf8Vc
B50aH5RUKRinLV9t+BYuMdGX3egFopr36FZ+kuYuqzgW+KbM1/BTKQnjHQ9vEur3
hpw9Bs0eQBcTz237chaaDb9bsJdBaCYJs6Bw9DFjrSgGma2zdwsM+dA4zJKJRxgd
3zScN4EQVVl/sbc/d87FLgryVhFscyDpB0ua1sL0tWcY9U+XmJZJnMRq4mdrB7qS
8P0V8HA/Xov/0aNBZFR8WL9ouGg318XTRSJ4rBsRZdUh0EyIeH173Uu8/v9F0AJQ
WPDGEZOwfeHCkHK194eM3MHtd6/dkOFmIW09ILML6hxW60yPsWdSpNKi23fDwhH5
dwm5+XXRi8ngDHtMEtTysFNRjIgqA9CPzFqA+dCrA549QXEOLNyJCxseJ3ekX/NF
IjjFMYd0QiQJyVZniV/7q0ag9S1fhKjtBlsZNi9QgxyAtdSfFJjSMg432FmY1BA2
k3fnnN9FFln92HCvZqPz8YFvhKKqx5e6GdUdCJMvLgUyawLSWQot/fe2eueoPzgR
TLAfRGgmBo/xroNu5XClB0DAQ3gOPxLxH3Xa7HC5LK+cDCp+XNW7mx/eO0yiWIuJ
FE9WRQ+BkNulFFNPngE+2ciLmiL+QW5Z8bdkurROzbOosOg5W/cT0aqsgtYwUGsq
ci4ebbk5gmiCLDmniVKh3F6sjWPXskgghgwCTMGqaMauQGxj3aMRk0eyHJJM5lOb
OAWdiBMV4bCJB3sm1+Ybkfa/KHfdRmO9Ynh/26dPpKnnqBeA7/mdgytnxJT8SgeB
EwsDNFGDM8SxqvFPbZMBxhLe8bMZBJkZ0ZdlMJVrc3VBlF+pFk+z4U6P8U3/6pAd
xzLnwYwQp8HKHpPWWZkyuw9J7uIAhPuFfJc/kYXP6eI/4rKJ8/RHTCjevlED87X2
elE+fqCTbVgh57/YZs9r7LS1z9WFSBLIp1fF6SrWSsxLfX5rcj1IoJqT7D+xNH6V
odGdLmr6j95ftfeQ4zYjmaR9CFd6tUV0Xy8h2lwuaTkVwSU4ViNMVYzs0p6S0dFN
o2fm35Dg4oVEG9Dc01lRJyaxb/qx9t7sOtYIvVLaLIr0Pn65sMCqLbZQpN1S65A3
85CtyobJbro/a1ao3Q1qSah6jOc5Am3DP/Ty7NtqprWoXFujUWjMthrXrfp9u56a
eXAkxvHINyXGrBFaIghl2VUO4h1HFVqjTKn8vpme5IfSnyDp4uNkZnTi5tb6ar/1
hp1wJ/SJQmus8dMDMq5zPhv5nWGko7zfuOUHwy3kR0GxCT+eRBRjJy4swvoq6rW0
cQZzp5hgVecSRX+deiRC9ZdD6Pgx0wa84Ex7puN+XM5vOk14wZt/SxEK7StwhjyT
ybj+3AWC/HMpw2VwNT9FGwhNO73KH0B/x5yNncHItdz9et8NPnSEtBpZ3iyf0Haz
xOonI2CQEH6aO/EdIqIHgug6lwqhrG1XyhyHnOYVtVCjJvVBv/EHyNV8nHrgZoPa
vDOc/sQq0Pl/ePc2TjKG7CR/cFHNV7sVbf0pYDaqaJ7ofJyiQadPGw/3oTKk1Yw2
1bxYED6unIEXLVEzlhcMNKtjx7HjkaOtdN8bZDgLTP0LhOYxIDRA57g5VoR6xaQo
9lNVnGBDNvkvM+SSI2GmlkglQX+/G6Nw+yaD6xzc12RSIdDFvDGRKuz6CIkDhL8l
6JYcinX0WG498B4Q7icIz8F/KR/7+NOMYEzOwjRWhij15szEnMMianZd9uVGOukF
BxOzDDpvM/hF2j6Pr6PQkTlwyPIPvqNK0HXWPzFs+7ZazBp7JZEWbaTo4w6M8ZzN
eaWw1Ye1zO8ksBx+lMFp55aPvorlVqytW/6C47lEwu9+NG/YXDU/4flqRtrRueyR
ZaL1A2MU1DgjJN4+TdoWLeeojdlXgOmOi1XM+NElrwcfujO64PgheMHkpn0nhpG9
pvV2VkcsgpGyg8d3z5tKj+QGubQgqS/G/1xI7blqgaH7U04BbDCyLf61tcwxMNeh
4Dgn8U0KgJoDeFfW443aNfCSF3xSrEAV45P+ULPYrNXzN8VSyaMN2cV2atJPQCUO
YeXUTd7ud+LUH+uCtXUMWI/0tD9b37ySJzVZ8WT7vql6+XPAMWD+CLe+KUqwRytA
JbGiSaHSRl8e+2H37PDm+QVa1cf9KUxvRYvuECOZMK4JFZCECIpohSLGU3ftuy4g
hIdWNzVg1+uudV2Kf7zwAmMkX7gfAKnwV7ALu3b7bGFsvfGDkyww5MkgN9V6mMHi
HwDKN/nXbPuG8I+lPTN/s2d1dtQ7XQ/xdPO1q47SKJTwUAvMrwBfFhZ2EO9J8Jt/
GGDGPSSCrromGTejDYMJqNZ0Nc0aX5PviKe7mdsLvOl1s4E6ZqoSsEUB4tCP9xvV
b+RSVv9e4OzV773NB8176owNwWxV5fgAy15enIn2DQnDZdvfocMh9Xy8kc0TdME8
VocXGGEMDXW737YbRX6jHiZ+/msUin9+xwYP+tnWe15RKnZv0+/MQpIKAzxZ83yR
30IkrJDVO80BQusd/5SItoJ4lbchYIxjYMNusRDT/9jgNiHXMqsfrpivomTnruz3
pahF+5Mk9AR12o2AelMFubpZ5uDRPilqkHeBAlZZLRH1QUbNZDU5WiAd0lSEYohB
QZMmxOpEtSNcKNcpdTVJm2mUqZAYoBIJF+F85xeqbm+FjDphUYDuwWIk2WKK6m6A
1ciPsiVZPJ2zQmznu3QIVe7dbU3Oo2wLs1/n8EUyIpNQQoBurgd92x1X0mRSflgl
FYILoOwa7ASp2BtxxzmXYPtDPjVu9l5IKJhm2jxprUBc+USH0Z0Pya6I5/Qb7g9W
hI4uE5ahSAvMD+oAFE1VF0+I3ct5mgGdkmwLa13ZwX/Zl12/3J5KPT+Il89Vtx8F
uvpRs/ajGn2KsPqr3z4/0Y9K0TENdVb6QD5LGcSpueTsWJ+1kAC74eKSAF7kYdnO
EXbxFPny2+Wd9uomm5BG+bxzNCoX9W2rymqtBi9KVG3dWjZe7TdGG7NSex8xKk1I
7wEGgxI82eQz2u0ojSCczSwXwI9iQidwcOGqBTTnagIPzciFGpZqNJYxRzqqQoTf
TdaRIkBTzWY7Y6egPlLa1a+M4DQ4D9pTzDX1DVBCbIt6DWRhZC3j0NwvBdMLsFuz
HOJe3rgvCfXKPn/jwl9EmbLKj8fJfeGBA+/qRl3DCv2BD/n23iWjYCm9gGepdPxj
hRSeZLLXk+03UdIZEI3Eu2zLN4GYRD56sS812xIogrG33shAWkHfzaIre7KBsxAs
izKzxt6Z0VtP+g1BWyZAhLRUHn/UEQK6Bz5uXGi+ET/y0Caj+kiZGXG0RzQsf1i3
Te9hGhHVpcLJ/vcRyfWPH9rrFndJg13mbrtMzKEZuTU5ngWOqRCAOhz2Z5IjjDVV
b4E733FHP++t2sfwqXOL/OXxnfjJLz7qFVt4gWSIXBB+Fhp8OgIk/667ZLStxigb
0iZomCJX/xtYMIhis4Ww9YWiVj67gbiC7yTHH/sugembq+wQZOpKYQ53d2KluPUq
PwxmkGzXCaUpKcQcckUPx08F3H6CiPYEoKusDoonUZyMHAzXJkaa0I4NgHq7d1ky
bMXEuO8eXLtZLkNIDl+/szTv5vObZLuuRIsU/0a9GNF6LUWuBXpo0VeJzkM9BCx7
R6Otd3wXERGcg9mjGnsBq2MSPuSbD0YHV9L2i4sEARPQ2AJCZlLyIwYlNuGSEn5w
2SZft1Gg+EhhVpYotUXfggQ3+cZTpTeAE+fhUw6iSLZRGHs8onbuDGnpDgCxMU0A
h1cbe3RDkAbpZp6LiOn1iwaBSRb/4DFnh0NkCRpZwEweZCs7HcYfnkCcNaSGCzSZ
3XI483LfpSIF8S05t4Du2Tjp6dM9fYEMBF/aSTekfNkB/TiAmYb65r9iO0NKoVnG
PfclOJXaLOjbcx39oDpeemhX4lJZiLsZc47Skee2EzQ23FVQrp5rlpnoFln3U7vo
typVBVXtZjXDQb/YAiRhof1OMgbx2EB1v1/FyhKdPjs=
`protect END_PROTECTED
