`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8U/Hd/wKWUtKcJHnilzHT9GolqFFmMt550q/aUjxiafl5qnQINyAkiGyrTpItlH8
AS5pGUydE51UP8lZ8V4iwBfIZYc//9m43UmVU1DPNDk4z7bPaKxOOq6GrFtRD7hQ
mXAmuq7nIpDXJGL8GiDJLvOqGGfBCkoHZRjJ+RlXqwcbdmUy8L9dJgPr5NbzDyVO
7HoOjdPxj5DnlNJj8GmRfAbfElSqdeuVTtXqTMV6REK3LAACitRw3ho6f7TOytxy
f+oeBNlQJyln9VW8PrW5T79fVPr2DI4SXOh5Cm3g1HIxIILT/KZI5cGqcHv6kVFH
q7E5wcf0+/ZYJU3tVqesGg3pI8FhN09ExDdUZF1zE4XC5iqDYAZuy/XSvxzhSuEO
Sa/4XtdJ4SWdx9c+/bw9kFNMmfQdPtWHHzpbzzMdojXJAFx2OmAjJgOs1w/FnDub
VXW+9JtM/C02P//CmrNeMT9FGuxPmmuUzgO+q9xR9xx2qOcpxDKq9O9Z0ZYvBAiw
fLi5AAewkzNo37FDnyJL6rKQc9R2JjMqdpfnZUL1/0YdyTKxV+5ibMF7yvr8SCr1
QCqtByqfy243XT1HodyC9g==
`protect END_PROTECTED
