`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMjJzs8m85KVAlywp4WqVBzzM8voVtCFXC03hc3OyCHbh2HI8/7BldDd4Bfi0hmg
od+DzLUBbt23aFCnMStet7ixGbCjfEJpoZY2/LG+vphiaVcRKdknzFgsWR832fkZ
mzhvgrfKzIX7o0PEZddp8BcT4I3y0Hl0HUBi1SFV4Ds=
`protect END_PROTECTED
