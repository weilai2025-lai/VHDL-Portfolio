`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSwhKhlFIdwqalG9Ket0IfQDP+bZ1Qwa5VT0kVcyeACTYNfjYWaPQJdCIMFolPJk
fG1HCWrXs7n8qH8Xwdrfu0zdYjXWz8XjU6qTo36HHTw8jytbYgV1dJc0YcFPOFoJ
08WOpF77EvCVwl5OTJ5cggvEN2xNC2z4YovCpWoPOVUZGJWcPZHp6EvEKAUuG9BU
13vyuW7Kc7uJSc3pVb0ZJpSGxc0xPujtj5anpy5rIJxQkUwDFbSj98TMXipx7LHJ
m8E5J5C9jIwXmz6sM0I9hflRte6tNWd2hV6U2KEl/vUdJR3b2OIMB+TYhRPzN286
p/hZSqo69nJ1MJ6Qtc3SQkBdkFdqnU6bh3Gb+hFbBr3YOh+pcXvbJOw6BqiZzC0D
LDdkA9/5pD/+k1K0pkaC5DZcPjE3dzs0wX8k63F3Miu7oSqIWIyVykPD6n0OPoGz
sKU7xHhukJR85tBOLmwjjUZjfNAZy5QTFqLOSR3xFjJfY8KgbBnTC+nyvKq8n8Ri
F93H/3Zxm9W+00V0zqP4ll64NxoVyF/kw1ypmGRRxtFXHBXL6L30JstAzCGdwd/T
VLt/rBVTUhQZNmIBp3x4VL6xWKpCXVEFwp5JRPDH6LjeEhEwETR0mhfWWBuwkUnM
HIFHL1zbYZDZXKcfiochZ3qzLHNmMDuRLAU2LgE/IlvFmGyvXAWn7zXpW/Mk9rYW
sU5O8E/BTE5XOrHqG0g6CiZk2XP7BOthaWnZRnGry+ygaHvs5T1nth/4D6B6vb9+
RaWNcep9QQ25Z+mhnJBftQ5mi+Nsf4FoshaQAmoCU4uNH9DnbNJqBakyqFcKxk5S
3Eg40P3BssMrkOKLR5T+6YEkGGoec16VlMA+bQxynxDu6BpbPRRPuochCrFFadii
nVWtGBrg4aEh8LA59BZJwuKXqn0kth1PJBWY7Mxv5nC+J0iDbzkznh5Zguj7EvfG
upIhKF9G0aSVIhShpYEv5ZncUJK8wV/8FNqq2pgmn471UYP684exdf4IKL+CdcwM
7vNZKXLsPCM2j90v0I9aE84S1E2DG4pm6B0ACtVcUJhzImEsXy9Hm/R7LiW03FEd
HMCjJt6pVD4bOz4Qbwk6VrjjR/V56d7sY0MOeVbMU3dy4/D8eT4fddLZA8HO+jsA
WKGUhv3HBRFIGI7IucGs6U8CM4usUSNmYSjkSm/N2jRNidVkqjbL+OXcHdyW7UXe
XgejACyTLLdpAK3EMWqZvQOoxNy0qFmXI/83tOP4mXY5LRMdvtc8eFWgu5iXPnZ8
BiPVwYAqb9SAaczHq7X7Zp28gasDNouSdr5eFghKYqXmsEmQF23MWx7nnsk0mwFt
p0D+TVqoL/D2j82sIt9jirqmLzGJt311reOD3X6bPci68AIzZ6y4Aa8HCVPP2G8d
N2AJN6g78+NpEFLT2pJnvgE3t4KiEX8eTb/NRFhwW3hSE599dk8fVqUEfdNZY1e0
KYvW28u806/8ry7iFfKBaTkqWE0+qRpfn3dumKQt3NTojMXaybmVVOszG7fB+uoH
xO8PBWmp2E6pkJn0Elrl/Cxa945NuBDWx78dgLtqvxrLfUP7P/4wiwCNnnNJLyq/
O7yU6LPcCNZ3kcD9gTUX/RItHIXX9oecWo9TKTYs5Xaa4p+fzRp4NtLnh8jADjnz
XgI0IxYhjJNDsyioXSI8stsN+ieRvBMTXDX7jsGd2UeCgeSjl8UZ/5hAuQdP6R/J
tHX+NvD/7CGrL2aFYMcJlbn1ABxTvsUCXbUOrvdonRtzm3IUd/m0o6J5kRLWLKHf
f17gnJwLUJdoOdk0RhQV+w3SKiOzK83mAgM1+NU0rIGQv9CVLubHO/pfQErhGkAF
jz769f1XfjAUgFt41BXjiK2TM6VMGiyASjGqtJEDupO5jVK3orGwKyP1Cykck4BH
7302dtjNzjk6ueCQMnM+73VpqWDrAOGyGoNFBADNZi9K/c4OzFvltUZlVGgz3fg6
t+ahZGKfoto2pawcZsoWGL9gOaH82f8eSy4yPAAXWHDW5qwngBZi9AQwF0NDiEnl
jnL1Sno0MShyF1odhjA6NiFpNu3WnCbbT3avTeVKk9cv4bwC2xRqj1kIgaJwf9v4
9C00qjDPYfslFg8Wg+EbgdlwUZp7TSBpSf2rKF6r4z1n9Rw2fntaPAj5tCLxyIso
t/oBjHzMbqw4nQay4RwLryVbaDq02chiZfX1buNosVmlbVl4TACVggS+D6VqmMo2
tYulzMFs4MwB4gsslmpAsPWdTieRKp4tDp0wA/lIrDOrEFjfZJ1pR8prfWSkOBkX
82xxp+50b7HHJ805ASJC6uUtRsS9Y+qyG8MaHWx1ZzOS8s1ma/O9ebY21oQCZWcT
/rrkszxdosmQtNJROuiEPj3qTiQiEoF76tlK55D9nc/cMN/Wg8CjYeYUoOg96JHK
vucdP4M/rPTI2JQpMRIUJonOR31/CKyxQTeeO7aaSa6aMQ1Pgod9fMviquf+kzBg
2VKyRgpCtXe4FT9h4ERaYqNfvzPeEzBYeBvfx3Aruz8l8xncvhZ+NEZPtRDByEu1
SMT/APnAifOecSh4WgV+Dd3/YBvMSJfYqc+c0hHBsKzHVdDJ7W6GlRm63Tlt5d6W
7V1fo7L0dE6prxjJ3ws3gsfEWzjyPBeCR1uwHI0idWE07dLnP4SVTroSupRD0ugq
i9Onwr0nI4Gekcze2fzON3dilmnF3KZgUO8+fWzQRKtmBu9KgocmMrX3Wn0M/i9q
u3w4UoG/Gq8HImtoRNiaIaynClKxz+11lEcnU2Y6tPXJNj+J4uSdpzD6aHNSp5tT
+3c4/SbpuovXF2EzWldovjoineic0VN5JoyFKD3Y3ZuQYlk/++TnbMyeJC/UC8QN
nIkSDwP0z1qwHB4rR5bkvWvHiyZSquXOrXWUXWxGzQwkUNhCISW6odGsNA1eDJ1w
DhrIOg8CN5etErmnfGBBW0BNchpt/1QyW4YMQZ+MxaULyc66qIJ8EoHlHr+wq204
OLdNuhLV5BDbseENcTbddLOqPxLu6X2WGS09Caac7jG7sK+KtCLSLluFyd+Rq+wF
Wwqd7zvenyOZY5XVYHaxywI5dCxcG7XJgecbdrtcwWY6CpFc0XyDqFM4YLEz/cMA
Tf42TMHyaNbTfhcED0Ergza1Fcd+BWu62PRvSRYAUbKThEDad2U+KpHgAVDEzbgo
ZhBHlUW0GZ+UXYhMU98AVLDbFvof1k6fA4cDoeOvYSsdjwncEkNe4Cd4gSP3PH7r
BEl0yaDd37t7ng10LnSH9rWY+RkHVuOEzfOh7kBwz/ign+fhocEJXCGzuHVsWGlC
OckrEKoYxJfF8leDbDsAFJNMhT9ip579wFxpwLLLNmIiK9F8nDoaqwk9U6Qvoi5X
IBdjjG7J2XQSDgCChRfZ6aLYzTF7646fLNWH88fOhJCkqIrb8K7NRYj+fJ+Tpqx0
OzrrWg5P1710p6q7G8WaDCaCgzR9OnZk6GUxfcMmChC14A3/YlZ4tqdJqSmPDPac
FIS7cag/OWhJOleyozjfBF/vCW2zlyN1QDhKb+0yNN8KPQew7C4I/9MRE8Wg8Gqv
vd4v3+UPFOH42j0yAi8/MkYtrMMyon7VkeCfHDdwNMEVbeGsHdpGBLL5dcfj4ISD
m/JnpmK42OvbyNKTRbxSamiZVAiEctyIO9cNmz1FuYjK32JjxsMrlwhPbgJGN8Qn
/vPxKXgbKuTGtaxS4BAQQf7A15omrhaas3jbEUzh3zXS18+GYxnJ1UHAgVoz4NE7
Rgue1l0+SgpA80E8Uj9PwkKXtwHWb6jG7TCWNLEgUd4R5vzWWgY+C4LN4SllA8m8
Ud3+sIyXQPT0/YSmpuTumWKG4FJYTNqd4gjRuUgf2clkZesNeHL91eJc7RDLpYPV
+gFY5z+8N9zsYkuCgwvu1wqsyP/fnTyT14MJ0pUdqVsWOVtuPOTTDU1gG40OG0YD
3+GNsSK4RHY5JnXsHE9fpKCPKaWb3fOxDPUEwgHP2u/liuh4xnlJcCozBNqB051h
ZjZs01Y1t9fpPnsQFQh6QNeBcsOW2QNq32DxbC67ODluLn7PLp02EexgZYY0Dns+
apz4g4Q2Kq4tulEU2NOoYZDmw5G7MJknREGHEqSCgSqJiHWV0iHx0nhdh9ciSeY/
yLFQnfwk5wDqASwlTSuV0N5Gi+wUbkMKDGhYoPLKAPimtnN97e5IN6R01V5vjeAZ
16XZf3sjBoDHx2F8Ylc3oCz680+5h1pp3/PJsOAYBoyC7vcCdZOJsMJ46BjAzZbe
+V6bSPh8llAFnGH4F7D5Y3h/blpaax4RhRl0+rnCMcgLaF4ESWWTG7XTJKQLAET6
WLG3ru31s3xiHwh32H/7uRh445ir4bxxNoeGJeZH53YPDT2wkAnK3eO6M2eM7Rv4
jFJkUqHeraBgM2tE4Lew+7djT23qBQBq1+RrNYkw1Y06jdtJmVWoOKMVs/gWCwZI
pt6brDrm/BHREIhFrA+mukxXneRiD2h7Uu+DpHKlm9XydoC5pRdmkpy48Pz/fvGb
ZqWggQqyF6IWlVv6zDwaAhuYh6OJ/dlIlDhRQn5sUQB8c0s90q6LSnmitcMn797A
29okbyHElkAXS4zAIWh92V6DfF+wkd79gpqA1d85ra8d4XqEz4LDsQODCyDtbwtX
wBVCUd0aqQOlI7shKND4oX0EUyoSNeNVS3rE3Y5aqDHa/JmibWuHyLcYgPysHBAa
GhFuCbM9lRiHnuPQ3rNx6y9suJIKcyjWC6f0/IA/qfRfOJcHz6A+3zK+C+aoL+nn
bUmke4Q0I34AZKcaWexnMLUFVe2suCHWrawBM+scG6eLksJ8d+MV9H/jJl55f7UD
mHVUrTUWe6du3MqY8OSPadzXtOJoPpZ0RNGbW5mzsqYlr2o9ePyEbiKrqvvMGW8N
e2KECtYbVA5n/orQi7b6ntgr+RvMOD83QqOpCTCFUhbzoDiR7d0yG2JsoOOsE3kz
zZMfo1lljVFkQ5jvTSs5lk77PBXS0pEZ9jZXw4VzAwlk6lxMYhbDdGQNPq4PCC+3
Om83ICuW7rO1I131jvVEALX+PG71q92W7Q+MTVUsn1zzZEz8tb0h6egOirSzWfcB
ZiArlCkgM4eMy7wx2v7qUXRSWM4e2cL4ubme8FTrn5aBrbuhT/+aBQvAjDaq/F1I
mNDyVnOmz3802nulrZ3fQ3Ep2ke1L9IeBjWiOy3y9OTukBNj2a2wekrPDytFSmi0
6z9F07taREUzaWjv0UpSTKS+hWH+X86lb60ZSEgopCH2rpOoMsBnFsSQxbiCBYHP
kIzIboIgB9aYVT5/E2kP8hHfvb09MRD00ZgIRUl0pAo1nHoLLJ1OUqoFSfDRsIcs
BKm7HXBhyVXey3lSASc/OH0XpFb1Maszc9IJD3gQvAJGH3H9Zj+7VIULEQ+mOFHO
kwqnunCL+PE80YmjUj8iIj/5/60uE5wdcPEcUUHgK/IxRLF/s1ATFnqcD5wB+iNB
0YQpS6Qsr0o0S9ya+gbwY68pW01l5Y9LkuNuuAWEaEXZ5YlfbiHVK1BjeRmoCPsz
1YzxVPVwR9wotZq7dWhCZRjvzk7ktqdD43k9/FyUiP2X3sCzY8X8vFhmbRWZxbvW
ZXQ53PXwX5G3R1UJXLj1CxKzIQmOmbSXg5v54pNkYPXVLUfA15B4ZFKz7DzMImQj
mU46/2XfBszQFbqEnTvIhdwCJZwvYTrpm0ASvQwSu/VHXXM9rECnb/B2nMHPyd7R
aIUjzkOOO+6SWjncr/lx3rAmUAKJjgORsIw0QlkRubbSDHSepmuKhObZUDT66DXh
EdGMGQhG/C+/GG0UCfFIx+Ak1GuXYediDNWeUHr9J1uu9v9MPDnYPcWZR83db+Uq
U++nBZRzmswy1vEWQ8dm3IO1ObdX+fxB9X3La4/UeTsFs5nhx/0DzucvIrS/JElx
fJ8CLVx3T4nEdfosUaP9o7u3Ho5kFZelofOz7ApF/W4VqvrTI4kiOXXk26ThOtiF
kXwpYW5Wktgizd/TAq4n3X8RPZTpGD8YRBruyj9nPvM0YeZrB11MFRe9VYPqMKei
LY7uOcq1C4oZMHXREtDSyMYSECt9DpIxOL6OsjD+/cc7NBGT/kgFZC5/EGTAjgOu
LUJck9joHS0uza1tCeFzqEfh7hcaBrng/JaE3ZYgT2mxqRiYp1Qdoeqx6FGcECHW
8Ks3PCaUWKdv2lyVDgBSOzuA+UMSg/rjXFwaAymgsq5Jm0RyvR9XVfhJ4swIj3KU
ZU6AMZ5QH2ztFt/f2AvNSAwVp88ZunTeDF7RQKMPPmApO18ESAz4zQnciVvmGRoA
10+/ucr43G95ds3Lk8U3wuJ9ffsYRNSJMXHFlcfCvoTiP7X/nGKVl+1KAtfchxQH
ohKwG8Yl1GfQDPnL7aEf+kjXP3xHWulAopUAVWGp/Vck+Ie7JK/pA5AaKpLB7U1c
okEmYpFx6+b8Xx9moK30FtGhoZLG2TUjUGL0ceTsSDmx+9moUfXGJwykVV6ZCkTE
ijKdoT0uOHshcCV/gGoISe1CpfKRB6k2Ko3KMC1+mKl5anaM6qNcqpWA2npLFbRN
KUSk5XfajpStklHGBYL5Tg2Kv0G1+ggx4OMQhvhXZ92ZNU0MYpuhjLHZbxv9IbFt
IRrAsxN+vD1YaSxPwYhrBjfohqj5hs7M9WleqOoeDjmc9scQzE8cOcVOByfLYFgE
7hXXtA8i9uWOqsdm0yxYQQPfWSnbu9jo1bnkeXVD7M25Q1L+NbqbJVs1l9Nqu+J1
Wan3AvRe/wQy/hzMIChbz1JzCHoxUB4dSn1pdAAspbD/M46ac3fWF5a2nFQMrgQL
1CbE405kFQod9gerXOKUONrqMoeWy1lZBQcMuDbJuHUSQbeV8Y2nrTbmLDAQERW6
T11W0nJG6MxMOY7fTXK7yLSZgzIEvqbB6B441HBkAUUzyBnhXotPj0BM+kKDt8U5
OvZd/oB5o1ku0ShKtYfHdyDA/QBd2qddT/ooWPfGcpJlwp5liFETuILtkvd+8Is3
vVnLH4UgSK0zYWitIAyja3vinwKcpqjBALNGlU+qSN13vS1c5JMYKVV29pdvIvU8
IL10kBTAswPPnGnP5pl64o/4g+yOqEbuTX/PnegqtryIZrixbJan2nhCSwbCfus5
dXmUbMYNMp84u+JwRzGnrI91BV9u7b2F4k5xqtizxOvLvVVfm5bj+7nUp1oonuAr
PZxmzlIwv+BN1zbexxvrFrgqY0RDXfFEbUHr5sBjSUr2xliOxJOgbLLT0yYP7YMC
KmvBi7RZ0S4TKBA9avljGgASi7hFJfka24DtMm40A7Bx41DqWu/ZO85fcNFcJx0q
GxKfItH5xHgRDL+48W6iwubhNKHf4Fzj2YOeBfmXS3q/XUfr7fEsb87ujPgSl4r8
7OdVx+GiyLrdM8ENIrwLHO7101OCmC38G9bMz8QPnUyDnECQ+okdfYRuNTgk5nHL
CX2GdzZZdhrEODCiUaNyL1C2R9B4sxenpY2E75rkKP13fIbvel0joTWlkHAxcBZW
H/+numumCDrCAer+pMrJ7bLqEQ2mo89mMD1/nNkVbv/v2y6kDrIzTtdhhg2klJiD
duJPe0tN8eTO8jnd930WLi0hHOoVSyxa6jjCIO8xYS7zwseqkLMvtyM8B2dpi78r
0Ti8UdEWzTwRLT/PgXZNahOMnc9EqFAMZekTwpkV+R1i1uhZzqzFBBW8vhtz3TrB
u1QwZsGJLMrL5PjlEGHDXo+KXHXRs040zeNVY0L0nAvzcthxSG6PjbcOGKc/pi7Q
rG+MCc/0u65ExZZsIXHfETPTLVmObBdWESad2yYtuHhMmxmCbbx4yJW3Lt7tpKGS
dVIvx4zySXtwe+X5c4/jiR/54Rjwwtj8qlmmuMz6wZPVijuYjTdMkTCtG+xQpGV/
oGykuHgGcQZBR9nBrBbpMVQ9nKUkuSKxJRisFt3T3/CYvFq/R00T49P0l6niKc6m
QbTJjFC+zPRPKm5EhPRh3a+LHeS75VSQifMP1MdRhLXgBuOeN2W+rmvyCyPTBj0m
pKRTM2/s35FVLQtHuJMvMouMCQocoiJwD8ZGlbLmRJiWWa5n/x8fujBUOhanGkA0
uEyXUsSqfg3zcPibNHa3/8GExrDvw7AYTpEmbE+pYmVv0gNEWJocT1p300u8JY7l
o/8sJkTRpEWsT3W9t3YM0dClcHaW6dZ3TICfUCTNbWe2Z2D3HGzjKka/tiLJ/EdZ
oJzZ3+f5rm/1IWpt6izbI8xTe7YEhFewvyBKIrgea/Pvn+IqGjcsStBp/BknlMw9
96rSJrWpa0cvsG8qILMK+xdqeXb8TPO9AAg1gwoD0DhyfKoocoRtChGigNyfnfi5
dyDO6MPNdSz90qsM08zk0J+jb050ThE8UH0PLLxHl2pm2BvT2Hf4fIcTRM9QO5w7
JfaigtAMa70hp9zsrtwoZvvad4ptoLD01S7430mKEP+ubLcXabwx4RhkAsZ6ILx3
j/sfq/HRb0XVXaByYUWwVPHaICGq57/XUEYUOHIQR8HVgcfxiywvNMaVPLhMp8ue
+OQpE+e+H5i2EQbEvTvimmBSc9GFXX1TYrD1DcTcK4ZDRDPdgReLeD/VOQG1qrmh
1wjMyp6P779m+I0kQRVnI7HAMaHRMjYt8ImvQIduDhpCYY9xRhZsgSDFfBPXRntl
gyuKHCiDKAZnPW5xuPNWf1Rz1g8mUr8gXK8DVeY9AqrQ/mfc4PYckoqkF3Gh5Um2
MWZaiYBaXR8PK2sYGmEL/dFkZyc7EyIbehKoZ8kmfvj+l2nr+9xCI13N+eCHfEgi
4oms4NzDnnOo0B9d87BLVdArUeCqaLh7t1PjI8deTLn8axBwFZxQ1n6FfsXhJ2U4
gXfMXShrWIg17Wi/i2V65IZrbEzNKg1wVFxzI0SZ7VsK/1vL84E1gZ7YeBJgu/gx
nKbTDnDGQ6vQpFlw9CwgQoIqhX70K9dFG491HTYqy2u7FTTWjww8HuS08cPnjVTX
coPPSTyxjn+lzbiCiAof02vPs6/8AQXu7Ba1EsFfagPqVeJGxIQpprizwci1SoJS
UyqAl6JlUPMfDok7+ruvOWz2mzUk3xA51R1aoXAjHTpWvEW14ySW8vv/B0/9XnNJ
e7L/c3kyuYFG/Jh8OrusWwTMDe4Sc0082cR1mpyPfRqpWbfrff8LrpaJ7Z5P2prj
7xE5TEqy5x5Rz0QwhAf/DAHMAQhEZRJPTHjhlBuUT/skQ6bWtnXen7bji4Atrx0R
NEcRwkzOqRrUZgLc26TJiTo8jrl9l27h7CoMUmEsJDPA78VgCNdASnvMKgs0GNV6
/BQeZezV5i/WdCOcTir8ZskSzjnicxLH2wsvsoR+Ewam/j6XuhFnjnj/A282EFmA
nZauYP+zim89whAIhDwofxYHDiAl1MaMypLUtnMxm5wm1FMCJvDkPXTR1HAHJJlC
woJu02OsmMALChjhcESJTVS6qso2WnDKtFQy/+iZi8Wcj3sprt1y5DErkFi8eOTL
HppiGmECkX5VPS4VP7aGG4J3OGBqZ16p6067tGLZ/RAooX+21HCLRHaG5Yw9SBDN
NL3DXeQgQXxIQ9OaNzQwCULt5ogXkt3IOV5IWLw4+ndZr0/I85CyEsMIcO8hGwDM
L5a09XxLw3Tk5IrZ4gf6JOHLtQ7eW0t8iM0ritfP4N/JFgfxwuE/DeciL+dKBwlB
RlWsEaSjP76k8SPAP+mG8DjB44q8/PjkGXQIwRF/HpIin653XsOeIYPat6DOoyRV
VkNwr4+rXMaXiXEatcxzJO8Y+0EbRFtZIlDRCdP04Y7Rv0a2Rfmiejnba06k/Rmz
T2pCWXp5k7iGaVRtLossaTPNxVeXXVkYkAde/loQHWZ0dQpAVZ/RONhdVhRqjoS/
xAfRE4ApVeoT2zdDDpT4PV4ZbPiohmYXIAGscQM4cHjVSjnqvDKtqvh+aeykZS45
BWMF5pEp6HJ1z+ZxLVeL9377mq2rWkwLv3WflJ199zD9G0Zfjvjh30T6ubtw1Tnu
ccLFhoH8feWu4cuYmG7xKrUGXQbaKWySjWPrQ8C0y5FEkqqkBSNQtyVndB3NeoAi
pN9u/aXmnpv1zVPbEG6kmvGPZrutYS7Ogm7XitBD/Yq5D8G00tDb0c0oAgUyxfBx
EiJfUJ9kYWkfi0x3GF4HnTerwy0WG8VhRaXy/ayngtkNTfMO34j6hVnEtHrF0Ter
h8uBJiUJ+z2NqsMxrkf1VbGntM9+MDy8Nu3XhtF/AaZJplfWlJJh2xCw5CYZ13re
Oe31ZWEMe8MJUmP1ZVxsR8pfCHdWTSzTOQPg/kx8dQesbZJ/vDdoZLSXUHbJ2nXz
0X2ArzAEX78+OWgzCygovLEP1LMzpJP5z42fzV3RBvyiZ8+0uW2i1Ka1S/g3TI4D
2dUEdIFZataqIb3XlA52Sk1sP2YIoyPYlD5QmLlmG0ezr5bnKAzAVHnnktbnBhuC
Ss4rq/x0pNA22BD32q8g/du8jNWwKly4uum0/+bmvO05+FI9r3twS/I8zyY8Tek+
4h0eI+KC6EazuSue7VYO5av3T0NlL5Yke3q56Q+UgimSYkDASa1GPxVFW5/Dqd1+
N5O0Wo4ZXxGrv6phMWO+enyDsm5kMLFCvm66RU6YTM1Jj9ywJjAa+z1X2wvMT5D9
SrDu5XpaZKRtDrSKjUHW3S2+yzm4QMgAFylRPtfO5n298KUeu4nmIvQJWrHBh0GL
/5NQO8Y9K60QULWSXlILTSQEqXyu5VhyvMxgc5oI1zsALqFPK5O2/h6VXkd8n5zs
1YDk4hy5nQtJFSXlCk601Wm5sL830whuZDYOnnIASNRIKr1zmJA18jc2J7wEpyL+
f78HXdDYPLHxVrls3YrUaCm/7qqa39HVT6lQRhUtjUoy5qDWlVf1IYtWjhak/HEI
B7bPRjSd7fYmfonMRkxSRyqoiQgsEAhb9mMw0YZniLQBOEiHl34vZAfz/rYIKVw8
Q3EIdGeam9uirH6ABWYCs7Tl0Lw2KtnRM0Qe05u3zM3rKksprk9NCEaLq54f3BoQ
GSJnRfu6Jt8uoB0jcqJ8Hdz/U14zp3YhS/AmQyj+nuZhdOEWEQzJ279Ws1qLlmkh
+Ow8F6k6DLYi45WRxdmNcfTz/wfQRCJWwA9/16OjBQ5n1FGrPXybKIyX+HsRJYly
IkWMwVwvabpi8La9gT+tB0hqCSqKodppGFmCYcNpp0kvvBptjv7MIy5I24qpmihB
2mkZJb5xB+gk1eDI9wgPDx2SWseVnvEjd2wx05q3NA++Ys8/NaHQ8mpt6wMRf40+
3baroNdUkwKsV39DNT8YTnupIQslt+NS2TdWi7KBvNK+5hcTCHEtd+Ck55J1hwF3
ELzwZZKQxfxmlZLMpZNXWa+KP0P7S1ihLij8GzYFwmw7RqPNW47zbE9Noh46qmvd
+zFtyFaGkfHhHV6MEqj7J9ncJnInS/xUcI7nbocp+Nvffdq8tKhDvlWhbtoJA/ZK
7z+KsT7ocud9kSTkpLgkF19HAiCQOwpNCAiYFg/VGHwuV1kolAA0x/pYT2zXpAha
5H+tMZz0oqJn2B5Sfplyd3PAayk1JOZb1xy/fnu5IrLh57czNGHKUetaz6EBw9Mh
Q8FjL5XogEo7GjKYm+Zer1okreTgjLHuK2pq2KIN2SlO9E81OTXI/qk1yfarT1xg
Iz6594PdaaT1FOVLD4rmPgbBKgtu7sA4mVWJ3xNDFwUEl1SkfWKAcAEq99t4lYmH
YRFfkxBzDNug1Y5nln4XCEtMqoWinL5mE3sJtEjiRxyS+mIfjU0YVYW7ocVOYYgW
W2y0IOPrMxgeq5s5+xXLcBCB8MecXBAuGpb1e8Wwjq+GoFKcOD/n8cnlZc6B3FPj
j3d92uwrGzaq0N0TXJh5G+BJSZ9o0d6Fr6VeSxwqtHq2vVibrEZ0V3lZtE1r1EvK
0fVtNFu3oc8EP+QMu3ejKlb0B+Frwigv99cliJRYZbm/By5jD4VGECzHkOubGmbm
nomaCia2bnNInCRsMCH0PZ/IC5nTDElLykvNVdX0Wd2AtuKNQZmwOVJMlqhFAbhq
yTCjM4mAkzuRK1PIsSVuesBAuraFoPtgK7Gy9eEqQqJHsv/J6xdVaum+nwaor0qc
8/694SdFX7eHCJJrt40HWurvFQEodk1r61eG7nk3FIpC+/HWmXYIXqFffIjNq23Y
Fo0iJfkla3iRx+N3VG42AuvvKb76+Scp5FHUC6oRjtqqC2H79Dn0/P+VUybjI9ep
GIehIS5nbsgipfjNGciX7+0FuIej5s6RBvptZPDJt6CNK4B4gFb6EXWlhjEUr60t
/rT/Di+lspniFiatTXtcVinPN+14sZzF3CGCcEJH2OEDf4xmFn6MrQR/dTWZbIqy
lFvm19AGpTN7jd6taIrlZBpjmhch0FCmQpXvhp0HMaF7nCBz0YD43jS6/AN6bC0F
/JO6WgnjfeSZ0IIYiwfAqmQrvLnAWhOrbn5J4Tpy7THShQewb1L1+8vwrZn7VZtq
9tPga36O0sHAQr/o+UiN3Haq9kgiPAMVq2cRVHT1zrjlp87oN8Urj9R6+nqJtUrO
XrHoa+CXWeKodErP2YxsFg3Kp93f9DLFEKmZiUeeC9TehVESju2cy9LYnDvJ6Bfa
yvILooumxZjJiFGD9t+qmmY3U4LlGBB1LT2RCjw4XMvxtezYWBpIyGCqQ3DYMZ9D
b2w+zdFlgRLudbHd0OyKYucquQOvPQuYJq4HUYLVQCBL3PuwP517S662ztxhAPcN
anNSKVkdgUYKqDcAjpaibiTokQCJ+51d+UcIOu8pomIZzplEBmflK08nwx/NlEcW
d9vZD241JEQPFF4rUkT1XweC3ZSETBlcvpsMVN7hENcfWUjpTTFZfgogSEyCzE5/
Wh+CzCEFL7JTHp/qH8p+EQwetR08GZnMADPFDgjbTpj+/oe4MmivZSA9gzNgezRQ
iBDszaH9qi/iPOg0fAU28zDx+nihU88vgWL7jw/20xQUDydl+DLKmRQtMOTFY6gk
94ENmOGQtHmfg67LgjJ4mh4KXnu/Wia22xhPgvXtWuD5dvhXN5GpS7lyEMxQh2YG
hnELHJAIr6q60xYEjqBPInUkooOfYDISyynzrATyhuMMWyqxilPmCaIZUKbZLgO0
gKoAA7WSeDHoTOEu+OSn6nLQ5r7lJGqQZ3BmIChuPd/DrWcfiPJLL36OeUpitBt0
zzEBnhYSWkaj88da0pvD7MUSXVX9AMJhpM4AQ3MZI4RCZjOMX03x5pFfU7e3Tdbk
x4F/Plfh4enPDU9pAxEIHvU1uE+EoFg9bq5DusX39kAA9w0i++t8ZoNs00cg2VBT
AbEPQt3FpvVOT2PR0ijDcOxX36liSiABje6R5OkO2SqA7+06MfJ6EgUxLhIdidxo
dfFTe/7N+LSdWV2dmqLl/g7xjKRGQGGxMDM95sVRw3HPmk3xgr6HwX+rjWJMqOCQ
5EBCnAkRY/0V2B1z1tOuQ1lYSDInJpWfKKnwiLuYu2YvX4KZ66CegvTCUi7DszEu
Q2Gt0AGYL07JeV48DYlTF9lhibNoXHLkejKwMZkbM0NKAME3iWIUj+HlavKXy1ke
YpjS8HY9pobRofq1vNt1kjc4j+0r5c6flHR4Ga7dKB4B0HfHvUYKJqf/iYXjNIlK
wBy8wGss5H7DOEDC37AdKcd4xKETADReSSDy18AlkbAlsedsMlJwEg64PbHRlKY1
ijRhiiSph/7mn6lWclthbZkn+fT5glqtda1FdqQZxvlXadk4sJ1Vce9sC8rrwD2h
zLFKs4UxmIf6+1p0Y90Fn6S6xtqQMl2gAK+fxSewgzZ+Oux7mVUlxPSfAKfMKEYm
AA0XWQoSwDGRFUEiq4RcanodpD+QvXT4NxkJxZEVMSLnDAkJStKVx/4tUm3XQjfK
xkG7zqtDtktsf4Ojhv5DXWUVG/PhLTxfJnnnWSlKqf0z/tja2RdIyu9dB9dQK7kG
TQKYjptN76cWLo6ryrIkOTgxPGhvNhjGEuwuacx2/iwoVF1LtJMY71Zcd6Mpkpe/
J4QZgUmUVp6lVFS4ATadl2UQkQ3439oXNf9FQRaTTqbsnF1i3eVOJM5wn2GrI8SD
UjcTVU9KW/9LT+DQDGV+obTa1TtHCtlcElLCgnf/PYLzIbrlfcBnihPYvOmbgjY/
8JAwkB1Sw728Nj/hH63Yep091RxxnGyKNdRZQrue3Bl07xmE7/LOlFmvCO5ucc6O
fMtwhRx1VeDwND0c/bV/FuzmbrAIRwqGR4aoenfJtux0sHQvJ7afKggx8ok+Hp4p
jMxuBLmjK4dE/8D7JScT4paqj6HFOEbrgjLEOCAzkvt7ywWjv1vH0XriYwZCGWvi
ZEhw0kmN9Lhu+5TN5zKn1md3O3bbwSO2s1x6XFbmxpAp5gCh98Ej62lgov952ofy
PPQkG/Mvf//r/V6klkjYsSZ6oGsUIuzLEuBxO7SKrTU+uMwpN4ye2aT7r7tm3wwH
XuDQ23SUQsThwyYQM/26ucDlrzPB698HKVsJf9I4YaRIT7YhPB8yPgQtiu2hgMxm
5s1dw4pAUHTn8M/WmM2qBgcC4WUb/rSeZSTFltNMy7Ji9AtFvmjuXywj7EBj6A5F
rGZTI/+CtMOc/RgGcyC4hksrxAAp0MB1SJgKgBGOE3Mwp1Ae82JaGl8bp4Fr1VQo
nrnY35o8adFrZ/SWlpU/hcLtHbQLD4pXxziyKw22r29Yw9W5sDpYInw3rZDkWshq
7hzXAaUW7+q1DLx5HyB5b+Yi1Lh2RpqMcD2mt7mja5fTm1N5z2mOWTH30EYJn4Mb
VK3zY+1EEAEhn4W8u3IcubL5lyZIj06JdAikD5Nu6xqYPdjTAVsUUzNRbeElM+uh
P4E2CjG4HUas6qFrioJM9Sul6NDcHIgFVtjnrFneLEG+UdS7VK0JPyXbu361XKvi
TFRGi/Ot6CXV6eRDxIDD+HpvIQMIS5JNfEYZxUKlP2JrwRnwts+Etq+dwrVEjH8R
qlLWNfvKe06g/yuX28IseXQekxeC45XsC8jCuUNDI7xZ1BnRqVSOZlyZGqPOAyHo
u2svmfAvZb1qvk5l3pJpQf2Z9PRdR/T1erO4rBrM3SEMizSqO+0gE65k6dO9QYQj
ESCPrIjy1YWVUyMEPHI9XlkpOqAnYErkIi+LL/6ONpqRAILJjd486sOl15slImZY
zGL31nZyezgD/+ZyUZJmekUxTxCjT46MGdHVu+Kmmhslq2kgT+Vx/DJPi2w5e+8/
halUIF65AootBvXpTJy8jfs6C7SdevfTcDVJUqTBHurI5B2Azvt+ly4l8onm819n
L0h+fYo3FGlVP69/4xRR4AF1Q1S4YqDuR4g53GiRAMmOBOtWbNWc22udoUuQ5Ilw
5ccvBP80gXhIdyVmW1Sgzg0EDBqR1HewsQoge0Hjk9plUW8qFraWlrDnWeIlLFS5
fh0nBi81TDtfXpKG6CBYCXyRZ96szxkcYQe9WKAvDgN4i+wJRVC7BzDhPJjX7Wsl
rrx29bPKu6D/lQrdSWQJ+Yt7KqRscvPKZi/fG8EGAaaaNq85BMrvE47SDLSv640v
DJy8AzztOATv1RQ/RqRJeqXp0isrDorHKKufl2Q1ee5MnvWP2kvxo0V5MDrtnA8c
7vHUzLd1NtJbHBgq4YKYTaqjerbSMvPaw2VXn3s8W3jiGkpg8gWwmtisq47wa1Yh
lk1d/nH1MFmcWpSdb5zwIR9NtY2dlS91IzNVpN/lv9vgX3N/7kvwc0Johs8F7dvU
AD7jDrKhMfrTF5ATEjjnGKMcZJE4Q6IME+TV0PcMKsBVxeTPCsbDKrEksvNKkd4a
N/u4VavH7TM3ax0lv3oYHT+3Cx2wKuGYyIIa9kIRjCGgLBgwmAo7FDNriBsfvtXG
0/jP+JpFnH+6mXxcECRJ9r9ReyEZuvWYUArrkdOyBcSSZVPfluYclaapoXjZiGa3
EDgmMH3QQePb5POqv2Iflk+a9Fu4EVYs/2gzAhhiqPhBO8Z3Ot/zHgxgM2E/xyin
7Edr57kyml2Ibb8okQ83X791/CwsDKJAS+utMDdhjhT7FJZJrF7OpRJbSFpa0m21
9ovvpSRHXj3ZlvyHFPMJgTc03KF+KGsvmpxEeZdqYAOLi9hfW+udtQfjYA3UUY5f
Rgk7jYfPA1B9JzkJGq38dPYx7eIY+CAeiDXEvj5ZP3+7pF+NGH3U67v/wvX51OXA
IL0oEG3MljqaiMB2IiILDucOCtTCi+mUusAyLnByyctE7MFqtDvIljwh1krQ4xWo
QOvw7FwxlohTFCgjHXNgJHUkPMTDIq1fwwNlJCuqQ6JbEkBCXNCXwBNC49izWP9J
FQPyWvl7xOKJDhaEGBEGidGVBclMNlHuNxzjBdAxu/ddQrW8MVZksg8RkiXHS7pA
XPY0sI+w1i/G6RxI1MD0bQYuNM3EI4JN72re33Eyho5sH3cYaxjuFZ9tBUQlshgu
r7QnH7xGFepLzsXkGBVtkzSzWTTvvHqF5oMS5LC8c1sOkufDPUmOeqNdYeo04Fxx
4FUq6EsCbViZp1KZz9Bh6yLzeFLV03STGiUjgEVafAuLAv+pm2uVFMZo5/JyfCqy
vToZnY5ZdNMZSg0QoVKS2qG6Vw8ovITTjLIMdgIFtwfcg+S3WUiyVEN4m0TECfe7
ouyasDOXAStwDFs7aZj/EI0ri7zJNSkBJE1vzM/SoRhIfxL/KKl3q/pJU3NWGARO
gxF/rgXdyL6Sm7xCo0iR45c8mWMSiyJXc9EXwIF1lWTH6eFiWs6BLVNvynPGm1dy
QlalrkRjJPI1p8b1OQWNIZqj2ps7TbQ/Jq9YsQuk4Qo7nzmLyL1wkeCinF/oIM1d
IEXJiJyvCoxzjjBUR4bffvIE2N6iH6CNqISYsYMxbFMwLfLXtGbh83cGJZEd3ZVK
AUOV1O6acOXo1NRqRm7vKqeHutyZCxwTckGxH9zM+0BhB46YbAVxZuOwqkI6M14w
lCYk1rX82U5IyDzNucNXT4+8WLqStxBquAvq/CY9t8hg8DGRAFt5XfuvbKtJsQV3
zWKt3XrKhvANg/6o2cEal9NK543y/RyeICGzdatbSDEi0iHY5yyUtZ+2OTgeoBWB
8nT1GSko0d3WFsJhtWkKyuGUB8MPTOdV6ijvQfR8GceEtW4fCK/A6Dw3KkRdZqcS
QXCV5aObqm5Dix3EZXie7xh2Zq36zMxPgpsTRzLsZlhYHCCED/Bzg3Ad02nxI1OG
4dMcSxuGv8dQKpaR2cvrpa0lKEUPPsrEqgslZGZPgtd0IK1deW5zqogeFvGy8bOV
G9qM/V1OgNnVIZb8BVHANvzB4BcfXb3TYcFnkqZaB95OxKSFowPtcw8q/fj3aTLP
iXg3fDgY4ycT3RdplH9xUwIJzStZcOlybRrar1KdNqDxGf6XN4BIaGYW/UymfK6y
PAYJQ7LUh3+ddv+iTEUcpVZ08atVmRUxC6NgbsQVnNxMsNiEpraiE+Zf8YOlhqhV
VXKrmfGMzsCm9Q65cgz2ztvqL0K1bmnwee/meBH1OavENIHuZvftKdIROXrujsVJ
KPZABYqf6jAOUC7AG7vpaBLAry3/Ad17OlbyNWRRUlyT66a4Ghifv0z/L3UN4Mi8
5k4Fmzp4LOt+bbuQWoyaO+YLpYz7fRB9AU3f1Yf9DP/YuvnhgToGrg+nvfibM5bZ
83chIFvfGLbAhulFKiSegxuHJdmFPoeAMXAqfEMJnIHKg7uBTOz89tpySXd3fqGy
k8iK1ulF9vI4y5Bvg1lFBJH+WrOiFduwKCslXD4+ydqIJpimlYpUGdwJpoDZ3U6c
hZAQ4vXeOJgoYWhOXNInkGUkicFfhd86PHPTqukhukwjH0jp9gODSnTYFyjnJTXI
SzV+bnJtXeOT3xNZ5NN9pTtW/cLMz8I8MsH4tLSFNcXdo7FJAuwS4n1gff6VX2kt
a3nuF6V90gFCWDZwaFXW1ii24BpuOvFxa4V2meHIv4L/c9fb/HyoRWSA67E55NFw
VfABOT7caA+oXOZMBSnwkqF19NLeKRg+E/ALtKz04ySqvyVKnTMOTEy5ieWj5EEn
fgPjfpOxZ7Ev4XeXRBIqJxRWNQ/WrRqZkgB1V0qSSIr5MPvO5m588lQ1ZP9DvOEr
0glAf2Gh1FhwH90QuVvj74PoRY68e/iY8ZI9qX9yHi5VcAbaNbPD40dl4dLI/qJY
+SjyQBL1t9WW4AQ7FKupNwNWsZWaoX8EuCJxzknQDh2PkSgVyocxCe744GQGYPbv
xGYOMvyUt/OzImKKa01ElrkVKILOvDtPMixrjmonNGKtoYhxOgfWUTFS7BHD0qQv
2yQITZRsjj+KV0j8lFeW7PIgvPsEBEiH9eUhRnAWkMOPzTDgzkloGL6ziTE3A1h4
1rieWWkiIWdTgZC8F6txbuBB5pUFTmEvzbY/6NP/7aPqF9QhEmoZc0M1eEKp1nve
kUeDD5AKA6V2ANbU9Arj830BdA67BrezJKLUYqrOLWPzOidZkmhDsopKZZesoc6q
8RzsuVuN99gd0inc7KuVaizaa2H62OUfOis0usRKTsOK919Stc6FeYnxftBQhOTB
r0op6O8y+zrKlwsDQv94z8UU/i3Aikp9YVhl1OstYRngOD10o3SBRbXOhfjwe2UU
iFPES5bT92DPV5qWso/0f6HIZRSfXi6d7l5J9mOyySPNEO1/CGHBqfxWo2NubPoy
QAl70Lu5yopBtFc3zfv2ko7oG7iwq4/DcDGIE3gyPLO19oxsIe4YoROqLydFypQ1
eXInxiBkIP1cr91rXPBSXv5I3K/f3pXGE3MOcH6eNbvK4ytsZpdZcp7nq8f5OLbE
Geksah/rzBd6JGZSxC4psQV8fRN7Ql3u9BTT/TF10LC9gueyZFoJy8grFbmKCqzJ
BSA+rKkv1MLDL8vgw3xk2hvzbO1o0RUCKpGl7uKAmstNe0lQNJcEpiUBts82grE8
XXl96dRmlwdhPxF4ccOyvfX1mcBMaiQMGWOIDmG+ATuM+jhaaj+56utTTlr/2e4f
6mxkHGHVfbIm0iPts02Y6PRpNWpZ9i1luM1Ni7AyOCgGiCuC7YUJ9Xyub2iXHpZJ
jMMdsEBK4rcmH1+IY78/eWJu9y7IXPu8Jywy0Nf34OYXtY8wVNjcId4gBqSompwB
3KCE7Yx1Cm+lcK3fiegskblc60zvnmDkveDG16fMCYfXWstAsVUkFnOdV9QUPUVB
T71bvG6H2IWyZvZ6Q9JC8mD9LfuMLhzlwm5Fscbp+/w4FW1U75ZLyHHicbeIml8B
Fqhk4xZZerFTl0PiI7hKQEgFG6TwAXyryduwsYgT/QzzuFM/v2r2j9kbt89yBSvC
E2jdu5BhCm7xyQJBOmvbCY7zi7cAa0EJ33C/8NdQQxUmhfs7R8yyIZy4uOmLNUlz
/cHL5JJlTxdQ2J6I9HZdgzCvQAqA1iYLppEXb+3MgGcDBX0895wg4GaChCnI2mxl
b0cGGuK6YG6mh2SaJivQIttNNUT0w5rQs9VSgSg3aYhh2Am2oupnftzN4Mjy0dzE
08AbGcrgNGYKEYSIrw5kqn6lRgRg9iXlcN0dlyMqC9/KWPHeIr7VEL5C9UjKoS/j
LvqbHiW/5143jawGIid344ocOj1S6ftl8+6tIoEAscd2YXt7D3nDTloKcsWqKFHt
8j0Ly6UKx8Hxin9/EeihoRWEgzrmyQpnz5IItZ1yuNGY0cUFdi5CTMB+lftmcz1M
7ryOuMvVqjKhTERmwJ5tiWuHoXXajIFdOi6jNsOWpSiDaltZ4e2839gLXKNon2eG
hxWiRh8fzpFwTzbt/tmmbK2aueXGGks/4Io/wk3vP3i6B8acG3xn55esyyRLDGhA
/v127sQQcTSwMWmhZLFti4JEqm0iMyUkpF3TkJX2RX5CTkzkcpIceKfp4my53MlD
O4KtNXgpFQRvv8rqBJ3HY8vjVIlqy6BzUeZGKLNZE/e6QPN7WfV9rksDrLozDcop
dC5o/ouI1xLWwpfV5cHZetLv59Hm6n8dI1UrNSfrMg6du+uWoZCsNR0Bia/chjy9
gxXEjLY0LsL/d5gKEtnBEnBuoU5ZJdwcR9Vo5VVmx83NtGhWtF3QO8ULz87cHaUU
/+gqWq1CV1N4HFbRPEOssps0DsKm8fmhVdTYv8UfBpU0+N0VR7Y4+SbtiodTSRfC
9+WPwdtTWUy0H2KWqrW9WjX1k5al8Nd+Lcf4jWQCgsV07Uvo/xEA+JkyYkEx1ze/
sF0l7INQYCEFIsL78OSpP3iPXt7WuG/4vfyL6sT2byyWt51AUsc/kwN7f/cLa/In
ansODfu9rIWnopMavqZLBsjzJ8vtgsdhg7uQkItWCoeBQ1p+uS5gzM0rwM0Lou6G
BoNCAYlvSaheRBWCoceN25NLmAxa3RRkHKUl7dgFOPiaNPupmC0yxLZR7r3viJFQ
/yEaM+p98tBqb5ILUU+ibq3euSYQBDQ0PVep9iid5GMyf+foStPAAadr5E5DHsSS
HVMBlxuODLNmxMn2OOgX223exmHBFBaSsmDdSFlgZBpiG6cKqvtpVsb8ZMVZmGuu
88fQFF8rNx8PnkXaw3hca2zdC5qFLaeasY45ZHANyn8J9uP+sPZm4VE2/fwnIEGK
Tp7sUh6xRvAdPRi71TLjVec2thdPrAT3YZRvw5xLMlgcBzeWlia/KYjkA9wImEhO
veUoO4HuhU+g3g9lR8Vo+7P9hlFEOgYE4xNGGCw65ONhQA54s54i/lrUR+biDez3
SDaHnTrySy8xsAhVjwMZTR4T8NR6CVm0rNw1fn5bQNgsSp3zwrk97/cnlf91vu6t
+6MYQJj/zxizSwb7tYkN2+XTYoeiitWDUHalk4IGfiuKiTyfzXyTT33HJeZ8REbS
6MG3WEBFM64t1sdrPOAcZuq1FIZZ2ZQBtsJSNtzOpBNg7B8QF8j27d60D6QqQHGm
sTYDw45WdBtHmNPGF7Owag7lgN2svK+ElgWzAa8x8RtP9askgsoRB1g/BGRzBw01
xZAiOhMechYsWhqnMUFj3zLYCOAbKhveflbnQ/Fy9VV5kqJ3Rj/FmUtlO6ktw9ML
U0fW7wcQlq6cKM0DB8TGs5VIk67VE7DC2LK/kmK4pW6DEJYWHxzpZAPqwIRv2r2j
U+zBkB6tLqL3OpitaTiplaAj1Og5lE62vqEIvH/VYqxKHLR14b/mErTRNGBv/JtU
kQhkSF1BK8zJXpKUYPpWXo+rEZCG9AWAIwqhU0PgnA7yjd29uH7Q6u9ssJX+9CzG
psFU6IzoTeRMiBj20G9dloJkjXEVXP5KARGD9M0EfoFHFSaWgMq5AqjvXI1v+yrK
4mpsTxzXDV0hcbxMxZQw03cuRY7KOaLI+LQYrHjvDKekBc5USZPKJMibcP2fQbmF
TrFZtx7KUYMSSxswJFbfrk4o9CGBUn1If5+H8BTSibL/ks5/R4s8TQvYLVOhGwRa
t15pLar89Hol/UtKlAV3ksLWl8DxGj6rjNOlrZtC7uz02LWC5nUpFzKMZD6e3ZAx
Jn50UjnTlmy6N+g1C/A1NtjA329pwS/mRwAb/pg/xmMlZRcXzSbOERZuXt8bt/e+
khxGSBqMiGxzXcKgC9iTO3zwF6Zq+gREfkuz5ruh32Vm11Q8Yyleo8Weg441J9li
cKp2YqnXu346G6v2sJnR6XYw5Bx1R8EcZfA+v6A35xwhfULHPFWyaY0vMtAaWKIs
IWTEQSBlcHCug2aQ1HLNsePtRI7qU9LnF5pF+NwQatrUO7wkifbhYZ4+5MO2e1nh
fQuR0HILaDDw/cDJHviB+Nx8CdXn1LwWzzXlNpv4Oa8tb8MYH8bw3MOxk4C9ExIG
GDK2iqN4Bmc/StWhGRgNThR6pXwt3ijgDASfJJspapOQZbNIDSfoDTJASmbs+KBL
+YD3ZsJpHCLspD9VLu/UzzWNdXS5O3GuftEy45vbCFS6JZTeLvTcDnOF/j297dUp
rpXSDPhg6QEnoGNWg8aKyY3fm/WnKATJiy8UhefeV7mRAtnW9qM3n9jfXpBEGh+x
WShMue1iqHG7IpoGX31iimi6W1ABjgsKIqz3xl/ZlG11fiHEC8TVuExA4lvQtusZ
PvmJOIdws/TeMs/DhieFj/GbFXvn7B1cm2wdbmK/x1dlGSE5okX/FIeI58BtAk3X
33vfX9Fj5nW3b9qGM01y+jA1jpCmYuCROOf8hSEjVUpn8j55IU5PurjZ/HB4I5Ec
hxxzHjd6tO/IvmyJSZZcjTRlvOWuGvIq665McRsiiUG4KbkPYM0p/4T2kNo6dB8h
0vNo3RZLXrIWOzkuBitjUiS7AOZbEsWEFeZLtefFwdndYtGMgDvzOyEcND4CPeWO
JbpjnO1T85JLADpUMWjn3wq7aZBWVVp/e/qBcMH82wgk0RQ8Q84Acg1ZH8FOE0HX
WqXoSC3bRmKR5KGatng6FvmNs2Qjba7B8F99P6W5hT06FvPcMBytNR4nn30dIszJ
il5TpPcL6b+tiBOGFGYCZNKmjR1X8LugUMJzHYKfC/t+iCjQwn4LCxsIvlZWwRuX
SFNh9lY5rZq0eB0cxXk7QrtHqC2FRlkPrEiu2ahQ6hliOsTdbIprVPj64eBujRYf
pOTiquzqO3WyDpS9YrM1ivuWIMHOPf4D7SC96oKT3BkeDtWhK0QTX7XAT4Kg6YXt
n0gP+s521Fs2/3aOU5KiTOcsBIgsfEYt2cHOzL38MvXqjSTx/dMPqJ4Vk4q4ARsA
I8PUqOMVMADtqSjKyw/zess+Ol4dWFjaGppC+bFT5W90p/Q05lrCbdfOBoNiSMOZ
g9Rt6uETC+i7x1GALHL02idU/6HyYpd674/4/CNOjNPwYPhecxuUg8sA4GrvN+mJ
bMZ754pQpauf0jzfPWNwb7DVLJ5EHmTLy7sVGohewI/KJg/90s4m2SK+f6XY2BVH
tyP1eN3xhUYAG3w24rp1AOVgmZYm7YLh0UKCdl7ao6XmzH0U/lGukz0yOLhkm61j
2tmUruUmn4TsBB1zgpxaMygiLJZtm3YumRiabEbVdVepbFgl2Eu0sovr7V5vdvfA
YzxEkK2Tdh+FF5Ln5KHt0wbjNyHTEbZDxH33H1xZJvJ4gww6/Nq1ylAJpC86L5b1
F8g4DBWYnS1NQKM6rHBVUcEDKwofzXd485rFZ2mdczEUT+2Jd0UexWNBQU6w63Vc
DaAod9kk5I1fbW8HC7xF4a4vrRr00++R4IewaI8m7q+ztWHVJIzW0AOSDrtPtfEc
OZmVib8kjCohFDtdTBKKztic2NX48BN+W5U8bxoBuuGreyD9KM6pu5XshnfT2T7O
Qcswdc13OKPdYIo0Yb3PDqlTFmT30ZhB6ca5tpR5cP25nLPWmW8GgqbU7BcpKjjb
MCdMzgWn5lp6/ZQM7EJgLQwoPTcewr1HcKgRXd4E3fsU4KtWBxH5bmGzqkMcb0k+
L2uKzairBHB6hKiDed6j+tLElvMBTykEaqO/KcZSU5Qc3pVdQ3U0B9qz44hlouED
b+KNCY+M7a/HbnyhZa4kB+gSrcO2deEdcTEzjUNsLUji+Ddzc288BIQcaOpRKEZe
2oHtWvRKjZ1nPLJEBDDWz3zSQaHzZcQlu17X1v3ASHlUDswAp+XqZMYX7GkE+TPV
lOq2tTfPkokx0hyuBh9qgrp9qHviFNGaPzR/1ZOeHlllG/zyaQA0E2OSInALUz6a
Nin4QUeqFAEx7pbnY94reWssoJ8N24BwMoUa2acc05Nxw1fJeKk04iOCJ5eiC1Ci
ro5B8qr/hJgDcpw8r4j9cFxU7k3ME0sHUwseoQfRQtDWZojn/MVJk3GFuyhOyz2O
XWaJATQX4Ln+CqOCSW0J+HPFcwYjRj+ww3FRHzgTIi7hlQaCpBx0JWJf+zyIqXMA
ni9XKg/bpQFjsKjJwqCI0+RfhMqV+TZxKOmZ+1QqXySp6JPunnF21nfkbr+FvP3p
WFDUcLnh7g5hgN5bWXBxyzXkwJwFCeKkzOEVRsDK/s0OchFcWNuJ8Egzz2Gqv97+
Uxgt7AQUGdJChbsHUtboYIPdjpLQQjbxE8IA0Iq7uagA6Z/UDyWwDigo70kRbH+F
k6h+DmWwAWqAAKYy4Vra8pUbT3dOHL7u2fXvC0R1AtoYztrt/0/zgPY2fBPJD4xq
zjkgWtWcth1tNnyQwK445FyCKYpWRNSNvggt4M+OT6MzmTOMYKaTcvbwAAY2y7Xl
knaTXRMJ00ym+ow9P9m+z5K+GxiORTificmftrssNQ9h5U27B8iKn7w2u89amzbE
wCCgznqbR4J4AiknDNQncHkWo11tyT7Gu+aDe0dCvTAyAlLy7mSxQYSdJ1oNZ5QW
cQRmJiGr6NWtuOspnVavmd7zySRVYYQ2g6W2qwV/R9++ZknMOepgIJbbsZBjIHm3
v8ojWG9syxSwqEy71DhfgOjMsqmM079UjrFJeZHUxgpxJpCON/UPOBuyI4PK7w6X
mAHR80s+4dODb1bvQJcJhOzC16Es4YmTBwLMP6MaOhxQv93nAjpKy8S6BM5yTjHM
ZgAaT3sLlZjDyp2YDnyBI5qEB+VUEHEu3nnbOsyt2iALG06JVtMTsEPo9nJO1MvO
d8bOLWtFccnV59hmghcMksFLu89U64x94iVPiGk2eaObp7d0Pz9IxhKYqMGx/Q6x
Z3zhnzeJI6gM2z/6I6ORd828p37TvYKNgkPIi6pf/WGM0qdZgz+l2MHB470vvdJw
QEzwm9lJSzgqwhJByTrBf8rN5OGN1R/H5BHunE/lYXKRC7NtE7vzTM6rmu63ne5b
Lm34l/i33/q9osWmPCWDCL2QAB0IfjKQaEy/54lymaqXfhIgYiDk2aHlqcRBuE+C
MZjD3uOIJXWoFB+u9P3e+mePlMCNBzuSweVyef35PlZK+IUJ8AOhd6MMLOh4Vluk
nl+ibyg6YXNQ5NTHWt359LduflyU/+HLu61eOohmUq2b5sCeBiz7LAyqPytxAoLI
a7v4ac7dNw0yr4z5A/TOmvZYo7kXaEfBz+qpvKoiJV6JDXIh4d93nd+7HNYp/nC7
jKIm32ncjJh4whheblfHssny1rArBWC+rLEJ8zrGHXQyscRb8gM1YS8b1jY7AcsK
Z1hWnCTFrvccHUK7MKF6Nq8UNdp1DPYVboL1O87q22dwVFlRUIKYEgPCPJ7B0pu0
6yLimt48S6CyWBWViPW9qfzWSKjrVSbARhnU4rx7Qb+MYygWMz5DWyKtATAeOK4V
PV4fbi9Fmqj+VYwg4ZpiB16BbiNe6v6pn0DruBPL2qmNb1/wH6qcgr13Lf25UZUK
OvHkR/g2F5iXNP9HeYG1pI8nujf9PmYV1PzQDIwq9jSTasAV166lCEj1J72sqKuw
0iI/GXjsb/ZMHhp/lkQfK0Qejx75q2+Pg5kwHyzTvc2nKrYP5cVXDyuIIQM2dfOI
hZ/hfjAD+GPPgcIEyv8ZDAklkKLIu4VTHd1DLMq8Ye8qjfvdtxS14DsraD0FaFlA
9uPjAUwOZsl4dckgaN0oJ1TOq5y+tLkVxdJm+/oD3CC6PWJQU/ZSy7o+1IQltnbb
p2wMDBCl2VHu3kOsRcatsuVxDjkGzH5Rng+0J5klAEIDWmjrgezVjzDV3WZWOV9r
WqBQLrlULXv3n3p2hozOO5duAQLGdunME/gSPk/8c3dP9ZElbfIy30rv09fp1o0F
mx12Ih5s0kFck79Kz9oV8GTQUP9xwQCGoKxNOdacGWg2h/ukdwFAGXCaYOp0Cwx+
+7+aQhcpdiO7BrTGqnOUOdTegOAH4XYbAL7aYb1Fbnw88NXlIFhjZQl6pnFjeE6t
6aijC+my240RcWMw3Kqmvo9PfskCQQ3vgWJpDJfWa/fjFix0vamNkmO6P7rw4Gkr
hdEEfUvPSCOx/gtL7bFXe0foMyxmz75UjARkeVhSp7UMv42xcN5t8ZDg6AYN1d5f
6aDolDKrtlw1boTIKJoMWplbfkX1Ni3KRfyrMDMzuxjflrkg2a5rUWNtpGw0JF1u
uZYsW7+K6SYwoAhpp6WKlFPbtTs+PrfLdyNK/ijSBrLfxfsZT4BCMC8KpmF2B7+f
IaaBSEDHkfy9leKKKGKrW7ub8QsDYpcvkayO1G9u3evEsruO+vv8hpMh0k6Nv9aG
XGNvkY2ktj8DgopTXZJrt7dfjJoCXewOU1y/nYnE203z0s9FekZ+F5IXpYyGXHJZ
u9Yv94hYVQPftiOkXjHR7mFXxGbbjvZNFQK7E0AelCYGnga4+29X4svjxX4CmUoJ
4JZsvPrIvQgKmZKBGZtZdysR2+rQY0SjrhJwxi2ZU9LfKx2AsdMhFOi//iQnp5Tf
NyGwYSiiYMMucovVXHjhzrQyT99F/PL1SOOkFsCKWJdbd+uR2XNudvtabnVIbfez
Iv8m6tXfmVGp4ksnbuy/AQWsbnJ1g+Bc7HMxDrKxVCK48NbtDX6XgNIdh9iynzff
AHCi5Q5WlPj4jttkDT3vjhud0YVIbHsHJ/kIKtI4yfri9akaiSiEE4hCLfxNjbqg
YTwy7PApe/6y1aq2axdThx4kW4LX/O+0t9CAu5eMPsjM6XrTztBn3b+G2R424vQX
8YoETyGus4gqz/S5SjS4lZy5PQ41lRD0lFzVyWsBOpEqvN+uX1k/WEeVqf0jIytJ
ISXOM/oOfWJ1Try9EsNlYD7NWI8R2Xgu8gxeKVh7ZJ3yW+Bimz6AO/yFgaWhZ0kP
cJkQ9kUkK39otmEmG88MsHvw8rswgOy8UnqSQzZv2acU6LAKTvtq6jsW61jf1TJJ
2vHluQeXbQTti8dEFv304DjxUUVMpDyaMgK2p7XItn/KHxJenAFdkY8YQotwIDa4
sq/xwj7GRaI6dGllOOcgNx7xrWmogpMDNMOozFalsqEvjQrehoWL0dufTxbLF0oh
OHas3goTyMqOj7GtZdFeAf4390ocmz3s4lW6fMg3mBRFIUE8zP197p7f73cA4mnL
sh+0yVsfGt6LGfGglOlZEa3H/DSZO14kMg1J5U/LxenEB+PrDnhL7sa90j/Hi9ef
vDTpXspchZvkMhOPPiMPmIARuZn3u9CA0DV6USBeZhVCgk6EO6Bs/Xsot/JUIz+K
VB1F/vvcGk0xGRGgkoizNygxEXyBbJ0CQ6dvRa67VKcw5Ls/DepjmydyanT4MeM3
f+ntRoBnE+dMrjYHINwwLXbeWowpyKRKLk6TvR+TsLGpuxn20HnQS+Z0B7f3w0n4
4SijQXn8zguHesmzAzx7mq9bBBQ+yVj+Etwu/CogWQeWZNKSyAzmP+K9WY/wqZkj
riPD4Z8hXiuGji40UtjMyxMWiFO6Bvy4DWGRw0WJrn5BMGhzfLk2DUHBrN6dX6NB
WDrSLyU/vPml26ikshWAG9gO8HeRcwk/h3RhE6nNiXGJHK/CCstztie7OngHXA78
7nBe98cmf33knZ8HMCMGm0//3x97dWA2IP2WVcoLayFDHyzAgD+5t9ySWr45Q4wB
lBJR10y3nU742saaCI6IN2SViewmWVbQ4n1CSQ8tqTqodPgOoQkNo6H5CV+cSYJi
beN/g2eyYy5RE28wIDBj7C5ryX1bjRcgUJGvdXzPWabe71BC0ISyPrCGQZnvVurN
X2Qt6KEclsjXZAYg/2C1/1H2Qp6pAUxMWfWDcP7OsQH2o4iazcI55sZo70Mk2j3B
82MdNvmLoz1pXP4ZEByu/uKn+zzhuHc0GZj0hx9Ht87K6Co3pMIFdmANrGPTUFXr
YQOd9biBVP13s/g8P3uRfRHeuY+/T7D7oBnNCObIEux5lME6bl1ep4epQtxSyT+7
gNnwmfSrfyCwmyx6eiuq19mIJX7oQoq2PckLXG+rf1Rp9x/1Lwkbbz1qyH0EVY+Z
uD2mepOZbQ+KhQ/KVQiOhJCszsFpQKY6OTu1FpD/KKckIwBSHcmZzo81FeAlc/FD
WzLdEf80pS7W8NzSe1eokMhkSyMLnagbNcncyN6K4vZWmxt880z4WzDpC4ERxl0B
WCc9cQNbDJ4OLRg6zary9xkOjgnJf/IDtAEuVfZ1e49AQZsBWQEVjXBjNZFuuZHK
0GY9MCTWkpbIaNoldv8UXIHYlHhwNrxNUccQjdgNRGt8mDV3MuuTNoIqvHYvMIY1
ErUQiWIWqIdtVe6qLbQe+gH/AbXY69fJSq5+astNsU2g9nAVZfx7dwt3jRqdX/qA
T40dx1qca6nwychAAoGnw5lDCPQM3vOKVYjqwsAoQG3FQyBVznci5SDuo2CKxBo5
eARIXSc6kR3zLgu3Ugtgf0yWpqW6AZAyAqNDo9vZ1qL6CI5ZO9rHA/9jQ7Ek61Lq
tfLU2Xy1VTKY661fZo+771kZm7pjMZ2/0zZV5xM8maUQgQGQaX1xPsHNpNK3CzHt
U4fL8xMfiAXvBXxNSqG7AYhhN/qGWv84sbpovYvLk+jLG27zZdepYHfoIuOfoOOa
cttaZ3ISPx6WvlxUI4eMD2VhE5uFRE5j2mjoDhjq5vMg+vcyEE5pkdzcpAOIwaBo
0Yt5MikHYEl2JRm6fyaHdnIjshGfah85bb3F2pHKn+ryfUANVxYqntyRNoDB/oiO
Fi+n5JcRrm/ZD7zsqoE+CXEgpW3ySRVtdxQ5ZhKyOFN25KwIrqfbJGUkOWAt2l1i
Jyamyqpce1SgmgmNQErJBwuv7UpsEMIs7fmyOKcLMiamcyj3PviMP0iXwFKH5DjX
gWJuir39v1vhxYemlSOvvfn/4bMx76fGq7LGAb/qYFFS/yi8HigTM4yETg6jeVll
ezPB+cz9tDIHXaYjuf4lFQu42gEIQ1PfcJkqzyJBpHQg6uqbCNPL16VYbPllXmMU
iUeVfrBHx1DFzedEpYC8k0Fy1fUCjWkoROBeix8t3qLrTBcBhEROxZk5DtHGC8pG
jM8LX1XSDigVDfYJkx2/RblxP8ZLoZ/RnKf4cIr6y/D/wMJA+6lcwAs5K0A/2LKt
4PcNcr4ojgJexa69HipYACM84fqtPiBRp8fmHbpGwACYIJFuL7+KAqZTUqokPiAY
NDCEaqjY3xAyWGJVfegxeN5cc76tOjm0T+g+sjWcmHhchhq9Bzl4qoK6exnPlnp2
zrx5KhuJPVuDaORczc6SOBHfzPumoaCBtEVyEwwt/MDyDqC8KJtBxfTMih9e3wKh
TQiqutV8eqprlRAuQBEcRFq9N+GUS1oZO53zBqLtXW1W6IxN1nU+oUx5cIODlc3u
2fwnk93XDCcNHr14P4Sh5F9Cyo1l2wvzzCdcThiGqV+ysOTPtVGnC5DcdJX9H17E
QseweGuMJDVIIPYzfU5GbK2jv4x2TNMTcHC3ECLdCGs7+ujRjfe0zK2tFaUZA2sH
bomWGgi/ss23EPqgTx4kqLZyG2NMMfuAFQRyzxPOF5cDDwGcoKyHlD7xDisZFn3C
bvWZ+ItN942u+8AhQmGUFLQa0HjLM4exWaHWQgZlNXPa60k+raEeS+zo5SUt+t8g
z/GFXqVTD7nMEax/rb8wMB0LvG12lx8UAEgDTGUEaZSyt1v8+Cy5rsx/ey3KcQsI
lOxITG9Cw6F6idBs5rZd2KSh/4u56AWib83Z+19oPr2Pp/5ypWOpSodi+AyzsV4+
HLUNd4YZcNr3W4ZHulkbxDYHmXLDPHfTvij9vcL1WnlFnWfDzpQ1SYSGPeaCHAxH
93kDxKtACZhSwNs+0qj4u0vM2xKPOwx3L/lJVw/zsrw2H499Jh3TbIGAK+wi/Jr4
1deNMvPkAhrwBNrQdJxnwPZQ55k3RlSWgzZDwmI4aVt1Og5fgaDPYazdyfLSHsS3
hhambF2Vu+g1x8vKSGrvcD/R4AM2VHGfGbxJ+36CMv6+fIkMvnIMsElIzudQfxUe
DeC3MjC/J5kHpSjg6t9hVljPmryJ6ms7AtPY3XqgdigogG4Kjb1yNBtQH1Ug9bI3
h+V1B+9888nsVJ+bDS4cXUsfN1ZCmNYkfaHXTuu3sJ2sETovkn7TIXvne8Lj+DfS
zbKC6utG1XeTK70u0uGDciFJ//5nRJHuWeCOyutXppjIDWTbzXG5pHK1bwqoryZq
V1TXDfd2PkCpj7ya6J95FDw94pfM47GgQtkhBwgdJuwOvfEWSQrmEDs40I57LNqY
MAvZsTuCJu3D8AtFPA1qsGXhSbpLZLt2l9YhIga12GD23Vj6HDRvjCPE593Fj44S
pTavjgsj3lmhiOn/x8htMZQBTt9kXjP4aiGn4kE2J7B/ZbrzFF7Vk6K6nKNAYPYw
mlJoqWT09i33xpK4Rkk7QgRbpujLlABuFLGbuFxen9vTTPWA+4b9Gt3nkiwvSPEj
WkC0uT+tDdpk+eCrbrR2iYgexxxUjZl+2vB77mOHJXFD/TJljGXhU/d4N+rYdIiW
DSeYFZQle2uim6+n6KP9fLrt1vjhsX66N0YCgJsgGvaS6VzLpU5f29Xr227FeBql
Jtlkoan7FLYvycHCqTawKUDTjAYPFQ8W1CUjD4qMQxjbMVH3WFNicnJbiW7znTOg
yOVcajqGP3gneCU1hWwTU9H+4RL8lz9zEFpgg72/W6fjseICkUGDMnuXnI3HAK5w
eVqxEex25dDK3OPprHEkTiuyr2++BGVKfDA7n42k8/mQ2CwIckbK1i+zNwz9dmWq
Jit2Uov8dfohuvgrrj6kQ+mThdhr5CrgqqQH6e6v2MQ4O8imvCZrLi0/JpuxIqOB
JMSm3HGD8+r+IxeDERG6yRwE1FeAZAKb4mVsghFVlEd9bx1zO2M88c6HtF0i4Ntm
pijXfLc7XVDSZ2pUJ3KRixQeUNPQrPlToMDzFyInLt0sRKuqOXuHI2L5GI/XM8z4
rATuoRA6K+LcTh7cThBU7K5GIT63dNo6XXsiw8HYPyWbHH4sBMvWK0jP3q1Vmhfa
j3QDJq4kqQFGssm6+0v/G7nMth9AYfzxtclMlk/2KQXddRrWySj7uwieS9eM5Qm9
IC0IbH+76MuOe475Yv7XHp9o2ef4yzCICQ3bQVt3lLHNM7pYPgRe6XB6Rf4CBack
HeHzolPpJ7K9QIiD3b+YCuNch0c8JvXtnfmftF5X7LAfXy+GLWtAFpnHOsK0fzeI
d6cm4n8kgeHbmw/9tW4PNW7GYWOT5u+fnGPuuS/CH3Xu52c+lfsA8gD8AuSZLT4d
Jt3n48XyLaA8RTq6RdNlD4K9I1HTzTk0wKdh75on3xTkRMDQMSLnE8Axuorqq6/B
aKsK/UZ479BMGpxwJcnGYErztopEFXoD4C6G0c1auMv9gdR/hxzxhUMY21rpa5Fd
8/FKsvA6uoe4ixhjg4MRuXi5FOd7Gqubq0gBZ3C8qHTQjggIOKnf2aH+sBo0As4k
6nsyzqUq3nkgAQKwjaPZnVJJYI/Wp3msfBBJJ7OKxzVSlEfQp3U5DTc27hJYXYc6
q7325RA6MtxTpGHJB2J4m55owUfW4P1MABmXPyYlZQUXzVvqLjm9hhtz5x8fWTiE
NW+TshsmHZxLmJJJ9WazPGo/w/7vxwUWNaGC430Yj1ZoM3hSAdE4CL29WE/JYJN4
rq4XrgZPKyN7psIADmvaUzsKmwMgHvU6yoHZzvROQ2sXUvkn80YzD8z7prd/pO33
tl6WIi/yRLZVbU0jD0Fr+OeXPocLJnACxnsorx5BFLqP5EpznP0Ij28GVALJEPn7
f9vZF142fCyWd4hitH1GBMWJDg2nUWBiyJGqGgJe3hfMTAcEEVVZ5F6wWlD0l/AD
2g5HZnPzO5z7fpHNByD7XpHTA4NG01svzfNO1UquEJ4Ww7uC/F2f7ZR2OxhiEwHi
3ju/1TjhX58/FufYzvQrpywyEl3uiuItEYJBnjfUX0imzKVMTEmPbktpzmHradUr
b6oelYfT5vN/NBq+mw+M+BFahMfB/V4/re/F5B6GSgf73WG4fA8/X3watTzU1AJS
kiLg/FS2CenL8iHtWBvoGQBddqBBBDBAk7KKmSLIf91ipEluJ3PdtW0U/x880AWY
yWg/lplk3iaGT0pcacN0CKWcrdZNqxpSBZ/ZHmNn37dpAodldd8A1awldXkfcTE6
sP4az1IydXPmZlJCS2XewcF63ZDV1h/kO5wFj2EBpxYi+QFGqLyz9bCF+Bigl8FJ
3n1hPZA3Il94P2ISE+oCll/BtSqzMG9qWhE05/08qXnNt9LkM9YHF7qfmh8LLRbl
95u6eZF+REiRPZeP7ONyhA53kIaUZnRLuhHzh4CYbjT2wp25M/tlOuhmDTvtcGWk
TpdLJeKaN8IpJ7BFiwyuLMGozo/I91EAC6fgMg0g/BKsQQd6M/8goX0FwUtjY7Ht
HrM0c+MOt2MNnGCkl+MyO+80vGbylKufDC2fyYVbFLH3DM94giK1r5BOYnNjDVrB
r2PAIStIhL1HOm+JCzqUwnrqSaHqh2wEJzODj4wvSYY13DxVcopM9mjtK5orQJWQ
ud3oPjvFXLJmNKswqyDiTNqUkbCCwcG/DFed3oe6uoorebML8w7w9IA9qkosdZyj
xWeSAFdoVRMlUO5+W7YV136nYJ5EUF6RA31Q476Lbnjrc9aKsunS1bZY/eocROHp
8iXCNhQLfvKURpGEUGshHvEHZz7FSflAOveAm8fAk0gQN5m/CDJNP0QVz67Wusfy
QnSDiOW3ZDZPwLzhP7E4iQKqI6T6X/nS912lagqUX+RNcLStHgHRbWlNrhc+T86v
W+0fVYYCvIeUb/ZqmLt24hSmyazmX2DhVSRE62tkavC3d8etBmloLeDMZ9BtwxPU
aA5EVszQ7w295b8kF/y5r4J0ulHThEyurjmIAQEW8diQbmHZwM3F/djKiIoKrNbs
UOspa+SZzMl3nllHMFUPZpjVgkQzvh0ATg/ZOL8kPSFifYEjwN6Y2p+PPB8zy9no
LMxs2jYdm6AWixYbXwJWVER/ATQGEmVrG5i1xMMkR6oaCT9ITT+txs3jWUL6hwWb
a3u0ZA11neh1oGiNjv2OVc+rm/+Fj7RD/oFOmhIQBaBtxJqkVBUCtAP8NWeW2fO2
usTmnrep0Y8jnU7FlPNoWEnv2LFXSQX5NhfKGtsPmE2fDYlGgtlI/rzX9xNOnF01
3mUbcv+0VcEZiiXqzAeIS70VbUeTGdVnySclyZk5S/95cAbqhhuVHoqrcOErvDOy
XWFHQzRbEWyCgQC1R7vrhFnNa2nz20n2sYwiM4Bl2awKtPqBJ0BYHPHIMhCCVZe2
TF8Ygc2j2itJvX9q2C040pbqfSeP0zD3GRRc1C5hUB+OdctZ7Viw7ZZjc6VDJunL
yAEP8NGlFWdvXnPpqbsr2pIrmHjqgAoCyH77SfZsSPuSB6QQIruwmjabrYwVuJ87
6QGMyZfdCEzp4SsTeZBnRp0pGrMnnlyyNJF/ebDnMAbOkhL7xbqz02g41jdHzYZt
6oyDtHJ1ofhvB4SKkmfZJDcyjIf0uwx4QPc59lYgDUNaJSr58q8kruw3QOz+PZVI
pFJyBSJgoWYKYymHtoLN/AfAlI1FnFy919CZiDI9KtAzWAMo5jKS5IJYUyH9QtoZ
UIUQl/mkNB1MyHAqK1a0vue3l+ElciZ7N6p9mPmhSFQSf0oC0mGLHK2RM9ssUgIV
0Y423d0anNb5pUqSfReRaygtimuRjocsVnZO07s5io1VXo6GJoe6qXxhMCvarKC5
tiHz0P0yAWBpEFFPiYjphlMB3yGgCLUghPa9xplAgkNCiXVo5tBSJI2P5HqWVQOU
EL5COJmAjOEbnjuDVG13xc/oY7OsXgXrHhkAHwOsg5M2wxKzM7/xZdXkxT0E/f7h
lE7pYarcTQLe0M2hdwi5rG9wSYPtG3NmLKpTIYkEyPVZLcvG7geDyGGhm+tPKAta
m/q/3Eqpdlr3zVXnBqAgzvU7WEGMUMhAnQzqCDRzYpw1rl3Necvqvl5gdvbf6o7c
8mXq31RBwY1q6Ajo59Jw79D91r39eZNjYR9JPmby+S+SGaUib8ULQ/0PFE4UHdCJ
lNK42OzgVlGNRtd0TGk7owVo27A5aTVPAu92drexliGIwhzPm5Kv4NYzufUFBHik
+LdxWp8HvLfQok0AC2MUuCitpKQrKZX/md2W4/EmRD7snA4BSLMz0yZgzw0HZHHj
9cuizV+fxw8Yvt5Sf4IrV9BH19PEpIE1ev50AKz4yIlYio/FmqV/szbrnWPxKa27
Any4L8mbjXEIqpfb/OwydeWkAzv6k9Vd3N07eXJP1+M4kcnY+ThNEZfsQrtwCgRC
I4k3hoksVr7iKP+0t/sEfvwDj4uGdP8oNmVYmohTALj043kHDp+pjuHXgQ2TXbl3
zcmUV8cTZgVtzejVEbG2KaR4VwDQUR64mo5BgEChZbfbO00NZvrJKoiegxzFl0Pm
hlGNJWwcDfLQM5sUF1nY2PM6hfTOw5IoC5R6ygrTngZ4An72YHfVMYg+DsiX7SZt
mp2JvmprYh1o1tgnx8bL1hKhzH4JH9PAYmqrfIwwHsaQeXOkHXz7zepPx3RbE7Zp
/J+bM27ArQKbFSiGeHcYg1dsJ0GCkzHhV65qu9L3kW0cmuV68n1T17aLrNA3Dwza
9KX4ZMnRBS3+LhPwroJ6GMFZUFpxi12BlJW3rUwdKVdAySqMIB3L1RvB9ReGBNVx
8WM564tY/zci8KOo0THZrynY/lClLAGp7dc5YCapHHjfOJpUR4Z9iIiStOmVefm1
B4aNoQPhh+AVJqkYcTrVNwCo4NsAe0bcYtSNNj1hcDjqlQ/eloini0gqSsroVSNz
qVvsIkLczgr5Elh/7L1eIo4FmYWjVamlpIdfZHJYyLaxUc3BbnxvduNZH/JGjQE1
e2ciBYruYNMGtaIMjSQh1wDJznxUKuggvFOtF1Y51zu24hLZzcYAWvFbokARC7SM
i7HLJXHW+zT/A6ANGqy8eZFEnS5dMOBDcchW17iN8vlkAOEzBKFtx1497GYBxAlT
T4tyDvyuteMavL+V+V0Qol2GMjonVXtMkJeri0RxVtdcIpxGnbuoD0MGC7cqMJMZ
0efbJzwXtdhy0KT6m26pOTR5+B/Hip8C9OE3/xPL00eljsh7zGAP8D+gFKa6fw3r
dZnNlXkuJX0ADxGfmQZl26bn6qeI7MkoV+v/x0ThPteRzHeZANAVcX4DL6m90gi9
fRLErI9p+cVvkF+VaQRDRgk6O7rNREGqrn0byUb4UQFt4vuTfC/2BZA5NL1YkMJK
fPJScJPOqyZSXiZOXcvuvhz6vuEzgCnLe2cq5dJcZLRR775zXAPOA0/DB5oEgt9I
idwRtnsQFT3Ye6lwuyEf8KRlt6ih3dCq8kCm3OUkBhH+10LGBNgVePiAH0wsyAVT
4kmZohyIvmOACY/FassQ6mTxN5y0Cy0HFO1DF8SkJr8vlpULJYoiDjX2DWVndf0J
pUK4JQcgw7hC48gwUGiGn907L7AKvMAMACUhewCSnYpcOhnNIVP5ZcL6Evz7Mjjo
arQveCnvfrvcfYzeJd4jEJGrstnld8yGHTHtoM391b2NPO/8mwwvMWOZinSoL6YA
8LxUkvlvOl+NOLaXxok7TP7MdLXJqzwwOyLab4756uCtFoOnQcyB5ojCXQZCmPVw
2oRUq2NSkdpzhM0uLZr5kUEm8Xpy5w5jaf8Wh1p87/j1iON+fmAwNgi4J9SgbOAv
8fE83JqKPT6Wb4fhU62g/dXDcfKtIjvxBxwWE/koh2TL63SEFWggAYKN/R3xBJDM
CL5qdTq6xG6t+5PWYv2z2IuBAeQybRva8gMJvFLof9bilpG3esXG3MFdzSJ1usIr
oMnLFlao1w6nrjZGs+luWEQBvJN1CS80FICOAgLrVK6fk3a2Y/UxRxvEQRTsdj92
qHBZws3/zNxill9ulWPT1PVi4hT99cwI2ioEfYxSptG8SQGgt0AUrpUoQ4kONcUb
ibgAqrdJaOd5XNyfZNQHn4yp42xF15F0SU/rpSndmX33X3YoJWNts3uiPK6wH5KD
VHS7h1XuePUtkZCd6SbDbp9HIxN6cQ5qMmS2jRTZdxQNMWCYJjHGxz/MEjoRKbH3
xgRLwIRxQJINi1PI4Vzp01rK5KG8wMdcd3Qaj5PkD7z/dz2BbTu6Cd2Rb8s7P7Eu
xx8Ss2Rn/r84AgnMnO1pyu+5CSKmOOVVO/UCMtq5KWVgT4Ml7YTue8jML3FTcMLX
8DWm4y9q7Ir1W1xsPy0RRLgTLpsJepLMF7kcBpcC1hjG7IMarBmH/sMXI9SFKgSx
pEvPxtsu8YDKhLAidrNGYgUk0NOGKOLC5UhoM9VRpJmoC1vQll2SpLsH2KZAa2FY
ZtzJ4kjRbzk47gxrEsVed95vOQxcEUQOdrPY/pEZBl8rMNv5/ZDk1/YytZVtYpLE
/rIGAs+o1cxNf9z23kPc0L6zTn8Pg7Gf1jjTUPik7yTZ7m8fCG/CzMvaieTFwM93
nQJNvChcmY+4wP4u9DbO7aDr5MGTCPLQgMuR2y3puw31oaDQHJNwRbjS1n0hRJOX
2Pk+Ui7jVJ2O/vCnpPX4fc8A/+oE8Ifq5OsbrFnXXRmoCVjJwkZ65+RKDf/FaPBv
H+fet2tabGrvrFV1R2rL3gB774Sdx1Uk8GeQ3tRE9hKxWsgScC5J25nbgdE99gv5
fZ1i9btS0dI+YZ3Mrw3c0HlC7SZKYRvZaa1nsR1+qLMY+MLiqEK2U7BKYRLdfbGl
AJJb+tGcmmBpDVPf2afH0d6x6ZH+Ahaj2cMFbaUqqgVJOxBgD1lM38bhDl99RABD
QFnMgTs20chIIISWyaq5VdgWakQtYc0Z750OO/VDCOAIsPEgFn8Ik6839yyyD3Tx
7fUnwYDTA7S4ZpCqcwac7DjDJFzWX1Mp7LVzdSVHG/s7R+pMMCDIFxMPip0Eb5GZ
CU45DFbO2NLio913probOVITDeJbEqlvwoTm3ezOuA+EqKwuOTSk7PrRWUhiNrIk
ygUn5TPEv7j/P3gwWIX3L9wh0Z+LaEJEPlLSY0VM7InAMGANMiDt57dTaScIXcWq
HnpwI/Pk7K+YokTVhazi2W6moWIz8PuB9UgCh345p47xvUyhWdDmdEBEqKIEpk8/
G5CLBC+n8o7o6DM/7uy/PQztGIDds5sO6kHLDFC7qZYUkcLD2C2i/UoZ+eowV3me
2H8MAWwj519GW7VxA4/9ih8c765qeDzdkhJDHcQ27r3OeG3GZWzim1mkZPwkfxD3
wVuZ9SPChfjW9BMu5lhc46LU+JyvwyoKTU3h+4S/pD5ygTIXZPnPQCOo1jehy5HN
ffuKJDmpjdNWnnUu2mvnwNZsOtZwkYtynN5NsPEVOn5YaCe2/tIBDQO/W8cFDgLK
gtNuBEiYoe/8zCJKjCHWv3Pz7bYhPTW9eiM7ttMEublJclRReGdyi8p5Pt051ss2
+XRteyXUbUEk4FiIfW3x9cod0HX7bpUPVqay+tLDthAmXA4jt6VXXX3kD/iQJUsO
IBRTGK1r1Hp/9MX6daHQET7ZkJHUAm+w30ft4M9Znrxr9CsflcMMXjRGSziXbsA2
J/quIUH7E4DHxE5E/7kmtVjM6rND3oUXkE20JrnCyxwuqif2FhNEU/icTRrQeIDr
ABRbRgTZ2GSg2os0JRmUKnYT2ByFyQrBbPeM50DlnHCZ/CmM/e8RBYSt4jinzMY0
NkVZiDqy7cxEWWjtwrS2ty19G2u4cRuBFSeuLZj0iUtKQZe4IYDRW3l694Gv5Nu7
tBRXFp0qJBU+XXB2YXqzc3/p2p2cv2HhxXaHRTnmP/X2O9yd3UZp3zK/9I64eBJz
UlGXz+F658h53H8mQqPbN4w0lxaY3mPLF9aSpV0XTGf2i5XUqjeDD72m/dvgxgQX
vWbKYg4Oqxl8eamYClugUlgn9Hk2sNadct55b+Qoo8Z5Ey0cQFTDwBbYGYknXT0S
TFy+d3A5Jhs6vN8Dq55YdKVarT2+Iokrldose4XYRx8N1XEUdZdDQokH6Py571hC
oeN6eveoDsCIDpU5XDL+GwFU+Ti+XeKoAsmg0ogYxL3vas6U6eugEuXTg12Ayuoe
Om67NM+NtNJsUsvTqHpQBCCmkxFfVBRBvY1X2v2t2bg4frhDqdJ3tDsZgXQtIk7t
CabblJthwEJ62XSHQwEAPVBOgT/PSH6MubgM0qIIb1zPL95SZ1LS+gzAGaMgj4SS
iyxGK46YYbtfmOgWF2nXxr1wpZMRpjiUwhycQwiHmd996mB6vX5ZfnIwnwG8MA7m
2glqdiy7fio+p/BE441IEU9roqKziY2I9EdCiD8CeQqv2yr9Lqrr5s1y6IyucaT0
KY0BWJc2gcHjTn5iHJ6omjAjHd40mwxJFEnkvPMa34dgphfz23meTJQgYiQxziY+
fkqAFrWR0j21aIuLWnU1Tpc4EsgTl+YAocHhBQA7dc1oXVaxSLU6Qn5NXLtfxKKg
scRHlyL3AgpCV0xytsPeNf/KKgMCXkdgJaXYlKUy7N/0gfPBy9KJ5y88NcSQMOXK
5we/8wSlR7svanHwO0GcjWV3ll9VnV3fmHLBkaqnkFuZ7JqLrpXTbGSPdnWnjNz3
Bko7oRXCB9Pux7bsCHdhx/cCavcnQtBFEEwvwYNLBR1/4QIFY6zv0bjj9YsuWmnV
oVVET7JsscXe3zra2KlWgP9ATDbchxGswYrttl1pRaZtirsszEh8/tvPJT6JdXTU
0XQzErWOVJjTQhpcqdE5ll+jNmh5j4y6QZvHli6JWaKgmAyIf8bgc4u5MaI2gBw5
/kvw/csa1AK/heYHJ4/DdrgSld3B91IjwgnOzf01cLx7horvyUe+VT0apC7pKgCP
QxM+A7KDkBf8Ym7bMgDYXn0CBOwtwghGRnDrWA8Km96F5xMAFp1aFHGkwUua4eHC
dnBO4ts6vX4sNu7OU36s/7aTRPt2SRWoDdAlbmztE67dzhAmeToOR5zbuhCHaNyl
ZhrSlWMPum+RXjI1jdPRA9/oZSPPGNdxNDdhvB635Hd/6wBmi8Uox7qEQXx89z6p
X4+hZGqbVEk/qJor3zyW5WtCPz3j9xve/kHJo5LVjYzKeL22eQUlFwADSqIgmRHm
Jb9EknfriVPFlY9Z9cozzzrNe3I4To57v9IBR1gzd0qOotVTXNHJSBbCaO+maexA
mD/Fi1dCfHoTlsD3QCksIDmqLHZD0vWZNQynugjZewG1Nbn6WywPiFA4iW3RB3Z2
7Lko8+9+vD6N5p9Xqv9yqLS8wV9Vpv2kpMUsth5huVxwdjASJXrZE6jb7xRV3Clr
T6Lb451iaviAZ/x/tH+2BQhrlGT6+t4fcASWST0Nj14zTsS77kHy1dM8ggi+6PIs
3sdh4i3RcFQhkS0JDKBEdyRjuG1Us+i8xddUZaGGIsC4q7A/EsbdEY/Rpbk4wx0f
kxOUh9Ueu65JhbnsC6bacLhen5IoWIfTur17yxmnJoHlGu9nLWuHrygrtJTE4D8a
3GWC8V8DLtZa0p/ePQ7T1qa7cU/dgsENL23e5IPPyBU6TV+UAj842xwFfEjVyy7f
xnUgKLYntC7xJe95Odflm6oq1gILfC8qS6F+k8K8e81Unxj8n1jhyC4tuQyom9kU
uSyOj71H6pFdQLQY3KDHyWCb2iO24S6Ng6IsjXsEw0COqcid6OKVYB5ZueyE3XTt
BNsylt38tnm5E0YO9DGB65hIoRfOnlpBXWM25BbBIFNZnJyn5S9KUKI5gaY1xcUA
q5hFoI2W+Aw4NO+8YivEsGpLGPfoSDwCXvaKNKomaU4rvbqKaFmsWmdQt9NTJ5qm
7iKWqBSgL1Zp5V4auIWpnTMCXt4d/m/typ+Mm07ZZokDFpRgdUFudZpQO3JHKTGx
izyLAPOfF7PSdUNpZACOyxrrBjUg6ykO8BnBukcF9+xe3wCSbWKlixFS49bx3X6I
31Xx/G8HYEFBDn616f64p2YojUMOIYmT7b85N8caIWN7sLm60pQ9o+FXt0zBy5mQ
L7ryW7MkAitkJej+aPj8kwfGPkkQuGMMM0Ktc2F9rH0WDDkx6x/S+QbjZdpVT6wz
g9s1BSfcety5JpUmo7vH60HfmRCxlQn5/TbwkSwoshk0xbyIdWRboqSEq6/80czH
0xNn/sQEns5FwZ8PZsw0Xt34hnq/NHf5UGQ7JaHpuuzD7Uy7vMFcqs/ZMgsoPP61
MS9IF/YLgk8izCjw8MiV5enDqJYMrm/YgpHKux2iiw4jGpz1UYh14eE7pyW+VFFp
c+lVeQy72mqLU9Uq0kDZ2QIC+5ZN+9Palij3wE/EO1sj5Nbqjb56+b40umxOQnQ7
/cOxTHz5lcHlZAoffvNBIvgNDSCQMV4L1p99UuvYCoR+riLe7QK8ff7MeQiA0brY
JTEAk/EnzoOKZIHCs2UvNcj82cZzqpBXvZ2jNdRuHhRbKW4ttdOIbDYsObsN2C2e
HmEhv6SxaZIylRk+eehQyC6uxINQf2U9BVp2u5l2AkfksvNzPWCBgzL1t6Rqq7Xo
2/WD65Zh+D4Ghz1tbM2XXt2ZsCx1S8z/Y+oARkblbEo88fxFGXG6w9COvuN3mfbD
hVEMskgD4mIfwOvDdopRmwtxUnagWr/EFjx+lt5cwwMN1SsL/UXbDzmwsz5w4NV5
U7FTxJA8Ql1H/P4jcXuI2eefXz96oH5pibZvHOA9i/aZNVEblYR+JqOW1J0llnO/
+1lBsYq+77wNPkqAzkC+EOHehsuwmJp0rxKUto3c/2xbG/MXKtL4cxgfZIB5lF3/
VCSiQ1V4dIT7kaVu8pYu7oGAAiuCmaBAAghL4gCfvLvEK4mZoIe27RgHxDH8o8CU
3a6yIuvmRqarH5AHCba56frWK8Wmvax+ZpHXCKKiickufIJxZOn6bZb5SyW3TO0o
vHHote/Vs+uUDNKX6wvy1YqZEJ1M9zCz0YeJc3Vtw3kwpu8e06DCeybGufQ1QNng
cx5n6S3ENsqJDM6HPCYP6YWGpOQDYptWYo5ZtA56Q4eODiFBdjcoMYDjEuaut2b/
ycrk/Myt2u0ibbdL8EMrCjtHizD5IhVKVFKvU9en3LzJJGPdv7WMzLIuXDdR/K82
cg//Fx+9m8zyJCADJckc4SjKKWyZ3a7vAlZpiZOKMoCWzUjF14GFSu2G9GaCiqRK
hIMkq5tfmRMFet0mNq7sfCXNa6fwUARaSOe+5qN9oX3XPqOOpCE3FbMpmatJaj0x
U2B4Gfw9VMlAnYKBFstgC50MkpJboWTvXhq5ziHyKoKxdY4Hj8X6eoMSo7Mas8rs
JQCDVNXvZIfi5uZjac8rAqwXTaZOYmjoJKqSvt76f+FRfDteN4IdhCYAor9PvMz9
fhQCiLWvQ+R0ITIdLepSJZL9x+V7sS2wtx1seXAKz0xQ6MPyt6e8oFOZkhOB+9gT
b/3IVsLGn9Ucd46/3+VPxpHmLJQwC8D/P0X30vS6Ld1pJacuMKGtDvFaRMSTr38j
Yi1pNvHspRwBXyEHrBsZlhzzd3QHXk08BxHqy+M33AyGLyLqxpPnXl81SmGzAriY
rM7uJK1lg3HYnisLoR4OfV+yqTw56IuAh8y84BIqEbvQvrHM+PKZxkVh6r7ag1fy
PDe0j8GdZRRmWHvOm7HCeZBJscBe6G37el19sbZk1r6ZKwwKC7qH9ffpL/rVLxK4
wmWJh2BG9sRdmYlPCJrKj1EilxX6vDM7zr+OGEC1dI8krNdd9eu5eNgeWtfeMKNR
slzVvsm4AZuExctAYS69Zme5U+v0aVNc53oV3tDbdWm5xLXeIz57uoQLhqnqyFUo
VV7dDPqtfg0PEVBRhOIm+pXW03OI+CdyssGRRFIEtnlD2bdj6Ah5ezXq3muzOe1i
EziVkZ5nNGHPLBONtu7m1At89PStQwY7tSHYgzr/8o+8qjmOy2AhPAsUhF41t6Oe
vzXbpBn8z7BpjBNtEUtuGQLVHs7P4dlUoze3R+WuEaB2Fz6w1x3Be7Qm4zN+sIE+
6ugp82QXQp/VYTFBzHwRL5bbpWr14MBgdrBgE1O8uLLqmjdr2tmu2lQPQmuwiOC0
NShAJMy8jFZXPsXjr4zIRvM/86ysgMCxgUVEcx/00uxySCxH8hOkpFLXMUEe+poq
IoPyygK9axSERf3HOci06fQAnujUVPjc5cJV1+VCQ1YaYFm2bWhrPNmnDlMpk9bv
mxBxnsXmbLPvx2PWIlt5/RD60pD6R1L73T0SQlvjxazLeu2MsiJkXg25mmkyGFFb
tjHwJXwRXbzPaX4XjK2WtI4FjsqKihuVZJyP4AXXkuBFEqXL9izz1H73G/jJq91L
B7Ib7TrDEM7p0xTNM35aFzWjk+F/QvjcuhI+j5YKlMQWhGLR2TU6cNdxYen17zUk
BjNbMjLbZKzegsBmgV4CdA4xmKbVctgVNXS3Xpm6iTo8peF4unmlU41vCYc28sDq
69iWBibfKRCZk4OI9/CFgX5M8z1Wpb8oBg+twz29bfO7zL0pk5yDMmC8PxKEq7UO
ZbKMf9cgOlsDfzkuO0EsG49KQ9Rw1FEWJsu3HV8d+cC8S6Z7IMQQboQvsX9lf7oy
QKpVD5Sw7Lneh40iORE5kyM2JcZkd1qFtZUUkKhNnbOSh4OGmbm/dLcak0RP9mz0
X59+Ql5aBJHr1S5tLF9dkBo/aJwYt7WW0xrIG2MOC6cc4SRWIvd/U05sq5pGJWco
WsUQfj4mBWxp7pybvZOrdBofv1wQCp4PVtG3IMW5/j2R8uaSnJ4dt66yV9M7xfLc
RXl4Vi+V1mAD0BkeJa6k3iMMMN4uZngWAIreb1b4Qk4yYpALo2Npu9oBLfw2hNj8
y2OwSNzfb3s9Wj46qrKTy5nwK5h+aWqvbWplBFWOSRbmV9Wa+YjjPpF2jMaiKPDq
v5BuUnHK+pNb+G9D0v4OrkBzBc9mxi0BnGK/tYARI3XJolfuANuaTPYd32Sf0wau
nibZdiVBCoHLyAqb3n/MlrtD2BpguiakX07jvJ7ke+Guvyx3ixtDEcmUSac7ofcw
2egy5Uu/StR2ViajZH3PjYA7fbmDJ7hjo1lUse8OP0th7PRRfCLOQnnpiMG8Jm/8
jyS+ZW+D9N3YHCJhVaCQ+2O811Rw71ToBKqFyi3XveY2fSWmYunbhfnIQ4TOOWYw
ple8XUrNheRxuP9Us+kkOl4BKNfyVg1vx1BXexIP82HV6j7HpJ+uQcrV+AsEqOgL
219Y8H6UlzjKqGSlhGIp3tc48gv9nN9aS6kQ0WUHxl0LwnKv5QOZ+mIrwRc7Dv64
CTAyKwLnDBFP7YJjeUQKSvDWLd0GLilXaSkRx0fV26ALqzbKWcLyj5OSK/wzowV5
7eh//hYPLLVgYXC3u4ZN3MCb0E+0gWgv4urBOIIOYWJb7CvJWPeVcDx087WLGq/h
e/7GtZ4QITWwU3+wPZVQz5OIqV8ove0P5kpBpYcz/F60YCAyPgbr3/qUGcJxKU9Y
Uweyoo0LKcIoVpDToO59/Xa+7Oor4dHi2ylbRkg77lhLGxDvi8NGYcCzoPjCjwMy
kg656KtlLsrqJpa60Fa/znFMKuvcVWw+xOEYsSR3BbPrflKepsKlj8wlv30ulpI9
28xThdjOSAsFixBRUB3Fj1xt+4w3mTvHKZnACTGKS/1mSPh9MsP2ZeyfbsmgwqNr
xzUzAPNYTazEac8RpMh4D6w7AlCk8b0ulrr3PICYozTaWnkxdNRD1uePrF4h/t3o
Qw9F1kZc011HMzJA+10aSnEv9Op1pL+RsiXyPdbG7Wc37Y9tDWLv3WXqPiyiMyaG
5V04d8tzislnWsDX2nCJoYl4sR06Lh9SO3CTE/sck8znqdtzTyJo6PHi5qKTt5wv
QKkcAMHgl2B8ALYxzqm13GpivFDk8RPn0ROhom/n18qE46YhRuUDt3L1t7gzAoeE
s+8W0/STyyXD7o9FPnKF0gdm8zX8fa2Jx1n5RJck1z1Sg3XCQaXoEU9aiPe9zXh4
DiKijHqjLrlMegRsjlY8+mgH889ac4blXVeXOF0ex7sJ/Mxp8vjhwCV+F55b0IWt
UfKRKTAhHCmS5Ed1keIreWmELl31MYKlpU0dDUSrEs2NrHwpz3PgZclbGFxxY55z
no5mcFNLVZHg2TLNGN5lRFCEhTagjcyoO8s/ejuh4EocgGPAEcTslt2rRi/TmJEH
UiFCFEAPrbHI+S6gGbzeBCT0H50/0gijd/lQcIjw+fFzZv30Y81uRvvGCt7ektZ3
f3ZNs9b5JSi9KPHpiF0h3z2zT1rERJ02jtXQgbse+JHeHiyHbudpBa46zTYJRgGY
U2Cv17GfS9fPzCV34k2zcvi669h2b3RnUwpxR7Rqre82i+r2z/8zRu8xRBsbUBYV
HcRHjYQQYohw1Lh1kohnI8rgszy9bRnJozyMLIgUB4EJOGk2e/lcRTieTj4VfVV0
YZtxNhR/yQoyxPDTOWIJAUaZnQlL/RowiLJo6pQdokE8GXXNyokUpJSYtcR5diJz
p5sBwLV8DTHBOy0uhe6ZDL/M1wA9K/uSWD7ZwpoMOPMm4qOgEeVDYZunWnRkDSNu
WuCQA9wiihSMndYYgsG65+0RpledsmI2YxSYZWxyhFDzYAG+zUk+beaTcCC4KhIe
OHwNghLRx8eHq20I3HIYxxrfqgKl3BIqUkE6UFCPax5CH3ezGpqIswRT5cOLEg59
I3yOxq+bZ3lQbePJhJXhCOUp8JZyhQwJRE7y7rbReSX9RDoOa8kLyOOhmbTdyOS3
bN2NTXLzgYBpyJ30ojhV25VeiuHZCNCBu3BLmx/Wtvm/yxRSl2ZzJoUJr71sBnS/
h7qX7yAV3s3tXpvsSNWk2V/NDdqQsYtF2eLr9RZxe9Zp4KrgjHjWAOu5Tvr3kQJq
pRCWfVKI9vlcqoGv1HQ21CgnMjrky8UTXTC47TaaW2HZR0LBxkFiZ212R76tjfWl
QYql2K306L9ICfCQltHyo18xCUho+khhPP97zeNdZiHLe2BI+mfhSCtxxDN6LnOT
q9wmvI7Ao4GXaoHSQbdHB2ZVuJ+bcNT1nfzq4S4llZn4aWXmhKlmNVNLeUVmrcys
GGTOYlKvJ809uz/qHzd8rsiDix9rbb2kcqEntZQmdp17vEW/hRl6w5E87LtXQf2C
ZCXH1+N2GYDGx3yMmNoxWXSqa2EBsEzismoB7vTBSEQsba7V6r8KH2xp7yYtzMK4
stj5ZTVol36KVSC4VNr58ZW7Px/1mvd9pQms1GcUm0VV7PghNNygHkFsYVBb2o1b
wOC9cSelsVxWWse7f+MmIaLBYR9ksnii0RmAnb1cd9wqXuVrG+wGRSL1z2Tb0nLI
FiOnTHlqkac5iFYJoe0plAe8R80eCKNl1NmlFOrgCEWYIc/l8Ck/4hXLZYzuPQ5J
JrUH3yroaSBOTE+qDM1GyjVn5F9I0QydswJtIQlVFzdX4nAiCB83NjGcUhyaWknX
GaMH6TtSdWsk3CE0dolmY97psiXdkYnBBzMjJaznj4BpsnniMhgzQdXoRp6nTi3f
M6I5dwJv9WwDsX/BpbwG8Ipd+wm2cXATJRunZaQmlB/AV3xs8vqbDvERtj7GrVGe
+0mVas01MJRcNEgIvgWypZ7hYxcVj53wa0quLv9FqUCdr9cItdN2Qmgc0/TB7Ouc
L+2SjRcUbK3LNiiMhiWwyYkETiutphlssDtmOE0YdlbQmSP8akPVcDb/yVkA21Sf
gy9zAG2SjaO1BKKw6qJ8aqSLM6gBQ+yB133USzK8cQH4JYunfur6TY+A+d+ncJtY
h7zAlU3xmqi2wL1C8mokY9dwnfM2GgXTW2XLj7sTQLwND+Pcgl0izphb59ahpF5z
GucfBOWJdhNISmVHkgJmwRKSvLuIWurnp3sBawp/KNn5UU4xr9G0PsMaWTRtO13h
SOup9X117uavZDTemtcwa+3Xju4s0uIsWn5Y/h4avm+guexfp3arMAy5x/tk+TtL
GmHtEoFFVAaDNkjY5no4FAW+GRCmkTRTF3VHQkqGkTxDGXq4Senkq6bqNkKf8gqg
bR7/Zul8DlmsspRS5bcfQZTka97EffrkogyEe10aceAvuqm+4qQPsqjnh2XLXBAL
PscouGfpEvTRtDWXvy9Ymiyw1WMW0OKg8dngfngdFW5wBwFZTAkd7PbZX2+/Zy1Q
l+jyVQKkprvimt10MHF1Ns5c913Jeh9wmW1nUW2KmM6MgEuoi/k9ht8QiLO8bVY8
7sCc0OwScY+pWXaWboeyY1rLm2KFyhWm3beB+7QUbcAZ11Z8P7tSTkYAF6/uCU1u
M7ULAFEQtImHotL6QROqpwdLJnGMUelwjSDa0H4wUASKdKmZ1uOr5dTIGAm2cwk4
dDSwZolP74/mMEvucmXxtrpDLj0eeHphgtIqyFAiyPyg70kLHs1yYXfUB1wfkIyw
kppZtPn5JtGylPEVV2RMdqyAazBDE4KoRJq2kX6rDjUGasNH98bdgpZAP49qDkK8
+ovTGHWkP8xWYILGxXqZzI4xy989XBVYer5kohTTp+5uxo5wiZRhHojayU3/6QHH
XmE6VWiLJppTX3krbJQD4mw6KJohYn06N15kN4vJbfEWWJZbKAM7tT2+MY5j56+x
K9GCmF5RN8h5Nzce86Hfv4j4l5XXrGy2jhxqRbCX0fPyYm25qEzhOHRTaXbp+Nel
oDab4KsVVMn21jXOvSZ2b1vOXP8CJSTrl+eePXNxw4WhvTMlOjawO/fS3pLzf6g6
TCms4BoyAgz4RQvUVukkR32t51BB+XqEN2SsyiiHWevKP1YbzDmu3Yk4Y2kvi3Ib
LD6XBRyesdre2RBMaC5PNECytHqVDZ9xxnLzVDvOpAodCbjbY8QXHVfLRPpZXyh/
JenderA7deoB4CV+4O9+h02Y94pSOiMNBPIA5cylr6uw1uwaRfxPmd5joX1/nLue
cNSLyaQyKGhpP00NtSG5iJjLqRxP1z473P4LeJ5d8fgtvq/8ZZhx+tlvoQCh5Usa
NAWlPJRxQaxCwfFA2DIzDYY69ycM3mx8D0W4cEIuX38VAi41Vlu5E90Z0uMXHpTY
O1c5UYPXr6j26isXna/WhLTjRXC+DTIrjpPDxX+IWzeB4uJQOvCF/J14w0HEFqgs
r+DBEWAv4SaAka0B/3OTqz2un38JBwYinsjf8Xo8FpnBMLvJuVcK0wzuRAQaEtH1
Bko0o7z/rG1SU3C6BEPg8/lF3FtuyFox5YtuQR3FPzHt8AJPpn4DTWqBGPdBaok8
Nf6beJJpXR07FJXxcXqBIWSayAmD3+C5xNkeSl3iZN/ahnWW6Ea4kaQnbcFXfuT/
aUV4/0m7mqRk4T4/efPDwiusTuknNBIYBDjl4l0BmbnMJJi7a1BR3QcTqmF88de/
3z1285b7HATPyLd7Xhnf5V3l2uaybBorEiBHoQ/EL1CVMsEOUiuC3CrZz3aX3jV7
XBU5PSt2oGRXheRiFW0cKz8aFe+EB7APVhOSWucARHQSXsRFzzos7eMUV5kcwh2R
1PHaN4K2T8wQqSvuNmOd4axwLk+vwHjOwgC4oA4kitcqAwmcP/vNhiP8OHGOHKDo
H2disVM+84hfGhPmygWBtYUnSu8mx+DX/u/b4g69ElYVzoGPuq0BmasnoO3Pa0Ey
UhxowPtOsYaGfeTOez+1UPn+v5HEUOgjQlsiKWtM83p7Vff1zORnStK+BtRu8biz
K4xMA7pV8tBtMfiQLGoNPYHIkiAYwT/J+zTEnbBmYRhU/S4KKHcdAD9TeOCLk7j4
PAuCrjVWK6zPsp8I+pOwNZjdd3eB3J7NU+4T/iKW2LU7yAD935iVbDZSMDGdtY1F
DHtnzmOdcFpyA1K4M9Gw4MJ7loehVVeeR8jE/JSHy3MSg0WQXF1op8OIFt14OFjU
HpDvYgdmh3dlIWyWNcXFrNHaxy1WydiSDrFojxwoCGe4bxCbf4wJaG2L5xX7Vaqb
argpJAqhGihedn1LBnx9JJGuz368P2OuTK+01e1ml/6e9ApMV6i3xmC03iyKRokz
yg6Q8QALuVnWTUb47KNvp0aIVc3PwwTG34Ok5p85eSPtufimdmuTa6mXG3z6szR9
OugCNK72pUVNgNQ+JQtwcPsjEgZfXxpKX7bFg4L5ViR6HL55QgCHyA2Ypkr8YFMz
pSUDSPoNpq9BgMA0oprRzmpTBa3B2pKyLXTEqw8jCXY13XpYgxYzxbKEU22cZWBm
+fCf6hy317etTtO9j55KoxMDNhZlnPL/2GIz6d6yY5uDMvkuI55uxL3CfcWJGYgG
/vp0GFqg//cBEnCDwEvXrLBacbzV/uL9R+WpMQeQzM89tNLepLETu+6uxTIprU5V
9D3fIMPV3XDbaujA5KA6hsQrXarZBWFHAnrbM6CkJ3lheUtVh38owlGV/E6lDuwv
T2jRkSUlpwTx8FLdlnN3fwhVNrrrR76tJyT2Dh5B5kXC2UA/JBmAuy5o89RJVc8X
unqJp1tiRPfewSC2+4iVyZYZ8mAdwluOyY0D5YGiNN/gwJ+KWBvf+RESxYkaD91g
xb6lLFDdx81NTZP3MSiZ2xA+5KnZEElNkdi8xpmi1BayOvuRiOJY6Z9sVaboj2gQ
cr7tjnEVHyKuRsMOnYgYRjLjqYqiNpEfEKBMs5+TPLscVjOFHjRCTivt56c4W4CL
a1Pnx8dZvSF9kMEXqM5Txo9p3bl9cZi67FtaTPA/hNKNx1ahqQprhAG9Z3O+8glG
PQVJQOpoA0r1fEjDri/6Sedp0mPONSCFFTWrdxg6jEwzvFnPjf0al2PbIDLYct5u
q9tpY0QRnOIcFPtNSjFi0V7sRPr+sDD6hPen+N/jX2Rcj+ct5H39zLiXUEhbV3mI
AX5HFRrCkMdIdeh6kicHliaX2NIzjDKDFeSWIholCHmn0kADzR9j8OMoMh0oOSx6
PQfd2tOrqrPt8aIsdKa8qvJ9NZAKrzSlxdxNhBDKgodytYfkqQO9mafBcyRM2gDN
v5G6MEvH0uDfGuapZ24yq22KVI+jNwn5xcvjUd/KTzuv5fCuyU3ja4mT+inVn1EH
l7DBLUJdgyEidWXACLkTBfo92hd6J1mygVjt1vwT6n2a/n0kpzQfru4mG2XkAoe7
K2LY8ea6qVLJch+Ti/+r1xCodsT8tV6zLXVJREAn8BCMCx9p8USRWeJdoZDd13A4
+Wf/iTEU4V/Sr9slZ4CTRDHOR6HzbkRVA1bRhAd3F8u1zTuFbHja2Zkq/wbvkN2Y
Z6T03NUyl0cGfPCBHuuypgZY2SG76kAH2fgMfAv0uE8kK+K0Qw3y80mSfJ2e7+Ta
KfKZnSZl2ap6ro0mMk+2/Sk0p3/NwicDAS1VaFoOSWTk/PedgLt8D3KiMKUipjYC
A21N8xXUM4cFtfUlqh7xWM4Sq36R/TeJfwk0IOczOW95Sim/yS+8lEVpbdol5HN4
VimWNFgexRE+VuzoYzwPnb23zvCmzFmZJI+c+pCGarj0M1C+JB+RIjwgEVz3aJqX
1wpuVjftx7IXOMhdl/rdgQ7x0jPuQwOGojWehvo5OLn2KvLWHHty3m0YvtMX2AXb
pRrqy14j76VefJIX6+d/EpBvqlFmpWKH1vBPlz7+Lqasj+RmeXPnYhw97YOxjCYa
9MoLYeA6rnp9WveACGyKXi/pUYAb2/EJnPrcsvHQJ92RZkDULkcjhf18yMSORO5e
yj6d+DfZPVSG9jGzJ/xWcOZx7ndoXQCT86ebPWSKQ7eBDcFy1pHs5oftvPKKYQ/F
RpDXQ1nnn90J3ILkX4YqDHS5ScH1BZd17+8tswudPxsGRMUls7Sm6IpxhXCr0s/s
ofxpkOKsU3uorDApoddyWgKWPJoLcLdq6+xWkXu7U7OOxeYM9RJDv7di0uNnMKUp
MlNt0Du/VZ/hINw3URzt6sjtxqtkDby2fcnDdHLkL+5xNjlyMdWcmBOo5d8U+1gx
kTN/GMNIg2ab/wKPMzc+r9uQ+vhpxQTxdN1SeO/QK29nUc5kBomp+VdUtJwMXCa/
Ni4wwZNrytkxweA4rvLP2toz4iYB3sCI8Oqpluiz7NKfXOxGEqPavdrv/Brwhkgt
gKg+D5vBuO1kndheLut0XXsYqHYTfkKtkUEIvYUGRFOB9PP1rqq7JlBN1Fu2us9D
yF8iKqbPNPDkLhdvo8FU9y+3u9tKvDwgUj+rEBUdgeZJW0H98nkyt7Ut49DyupWp
AusW5xwYRTVYFZ4Gg3ANaBpEb1gVLGbyL8IGbR0CdiVpblwsdLkawudk7pVeRDIG
TxLujAndExNWF73zbBay+rY43IjAYbXjHe4zJyGoymDcnWUp8OTsZ8ygO4iZ7CuC
mKAvNZX3slsdS6+ECHkWVJndo2G15f8eDqLsNHSC2JIjIG26v9WkOTR6hS0Mtubk
Jo7vFWPln6DXaP7EJTR97mgYsanBvoi1Kv4QDGM8QLdrRM571+KWCG+nY3e3QvoY
+pSDIAvvFkapko2QEDIjRWX92tsGdgmhA0Q3xWmkV/Eg1Y6uaC6TpruIK4OCwvcE
YPT3Fddtw4agXzWjYALXEFGyZaEGVG5wAMts0BJhAcGu15F2H9ANpiHQ3qOjsC/l
bVXKURKrOvFm+y3tMM4V9zU3fovCwuf5Ifk22T7Sqt9lA3neE38hUEH9P7IA1YaD
SGowKo3eUSYezBlNb/ECpD9xeX1Po+2laSUWyg2CY3flIaBBVb9qkBKWvCTCkiSE
NmK4WPPidHx19zBeXwH9lI4DEP4xNbRaBt9wQZdGHocf8SbnS4flkU4WjeuyuzPT
kzHQbWEI01pQC0bzRytKmkzH/9YO1zKhgC+uCktySxyS/OZz6+rdaW9is4/DUzsi
ex6cxoZz8bc1+6Q4CiOvog0S/eW81SOFnpZ0fPLTdR2gUKKIKDag5zPaDtldGzqp
2xhAm+hoiMAPfZKQLrgD5EA2lJ4I8tJBOwQDVnbDXrnQSea+o7IZEYbdT9e5PD8y
c9WkVRN27gwFv+bdvG7U0myYc9zT2qHsMWTzYvl84mBAYJtYSRBm7/EBzyjt7AZK
UFvS91gqdqHi15aw9oQEfXCHAv0G9w6kr03ViLLMnS7UEp2DCU1hUGJcAWHhcOrg
Fo6vJc5U74L0lNnDzZbHS1da9EjXvbvdoV6yG2xAQp//taVXXfeuJAQsoqUjZ1s7
cgZy/Kja/4rbXsng6Vcsc5Jlr7xE0jV+kqL46LO9+lsZgMawIehTm3UBZeaTvz1O
eKCtDT61cHeEWJQpfboZ40apqzOFU/jAk7d31VKWLMbfEVkOVMBh6HFPk/MwAZ3+
Dkd5cDe7itMPJ80Heey5PCAnx202fr6rMAviA1eoFbMmeAevRDOPxXSOGrIjk2X0
CLtlFhQ8ZLBHuplTAr+Xh1OmfnHi5pmeKI9EnQxACu12X2BiezsFTBA1fGPKV76N
sBaWuPdZJXHynAfdmublGkPAnuhnPlNQhNenG4VLun8pEUKHyQ3baNLrCivVNrAw
6wT0KuN/7Hrqmfa3CvUviH1b2Hawz3OA3r5HnIg6CYh/mtCrzdi3vi0QW9j7K1H0
QqV55Zu7+Fy4o0KwJ1uU2cOlVXpD7oXuhrVpnaTXVPJKzcc+0tM6WIM/ofMkMseV
YwainLzT4Mp9F3yyxFkLdaxef+dPA1TRFjd48kgbMo6vspRDuUyz1+Pfb0YJMkyx
LtqUdi5B9eVQqjPWWu+4Qs5cO/kArjcH0sP4+hF9mPuaOtvXueIQuH4b8RUqEJJL
EO2T2+vhCt5vT/0Zn0T85MNZec8dNqpSP3aGhkbHyUuEnjVdUEM/g4t3FL4g5d6h
FoHdyp1g2x1ethoVnWNeALyeNpua0sOMq55kmuOUSA8sVGpBBhy4Et4e/ciRqPWk
+FYzTE3PDeVrlU7A/YWaikJqiKSGwpuQpG2EQnmcgOYvmeMpERIIqcKsgis/xRBQ
ZOfzMzEm8JvCpeZx+WRMkLkUEtPEwvfv1GbA/1ASI2T1c2WbkUA3RS0lg5RbTSSr
E1orcfC6IHwxf5d0L7mEFw8+svLhLaZFeQzXX5P9mKCQaXb/7tpn8UMrV4t6zFXw
CpmYC042iKQLGG5kMwR9x/lXlW2UXYJQ1TG4i80bWJPFNQew0QZRp7Q3XellPnNu
oq0KaT6HK5+QmN6Nn3dGXEnN9Zvfopu/4S7gkOB8LNzGarv56dFJvpdMkSR6iu7F
4KSggdaLEZ14nYKMQ9Mim1AUocEY5vdq2pW51qbqIQkGbD2qWos7vf6JMWsHHTPQ
NaC9dUL4OIfNHOX7PJot0GjXl2iG+3gjt289Hmqbkmj1xXnt4C9XoFU1xkcB0Nw+
2IgprBFmJHRPex/1nez18HCvitD6h7kv16ya1V51KQH5BgKUv7/LEjpJUMeu+0ri
Qgaa+h7I0OsCt2SUbk1xkQAJiQdCjAmcQ73N3cHdseob+D1o+PCIgXCxHm0nUes/
1XqEGCIl0e84Xa0LClTHdCiuVbSoAHcr+Em6NgO39d/cNDtyILHi7qc0XGnD8pxc
mvE23hvKkWETjjWUvzTZBsBklXGRb0yJkLtsY95kdBXKba5VLyVyXX18whCqooSy
ajDFC64ASRSVdKdKhYKX1BSfkiooq8jtxRiiklXrQWrVmG+FANDmVGWyGmLROGg6
pKawBTQww6j7GmnsYQPkQC8w/KjyuyhRm2eiPsv44P5l2dfdxyro8Ork9rWLVCJz
Icvm1tGm6vtyYG9iLA1qZJfubcDUQmYVP9VxWC9mo62X7H0c1XCPIizuCkKED8Su
3BAjYI9WE62/4jeItYYy22aVvyC7ZbsfGmRBoeL1OLtoQ73bRKcNH5fTwqwFolIB
1dD5H/NlEjN2G3i0eJP4pFHxnXbgGkOYNWriRnIJ5LUfR58+0T+GPFao0SKyHetB
eZ1APe/Hic2kLqxdJ7yQn2RN+/X0ZlN/2bojrtGTpsrWivpxfEF6w1xPnDRhezIm
gmuuyWmNvQf5y7I44qG5P3uouSkKnNet6fYAP1O+JMYfr3ds7G4QYB2VVZ5a50oW
vFmLgv4b3/4jnnMBb9cEBgd+NWUU09PXCT96Ow1qBQNsjDGxNLqz8iyRjtM8d1xp
/rMcBScf4tfj+0cZbSZiFiEySS5+51cIy2TwSvTx4/uq/dHwZDesLnMlc9ZtSFel
8GzuRsGpw7PgqKNMk/SpOmrO7twkYZOSDkpVv0bTYwepNtkh55iSswgNgNn1XWut
ypL7V8Uksg4a6XFo0LlEgCDbpx4VIb63o8f+uCS5U1lYOQ+BTimHrUiOGBY8+una
FUt8jogga+Vwy2u/e9JeO5AbtFkAMhTghBMhI9ggBZEINx7gXWRNtuGGN5y51tvx
MmP7ErMt7il1n7iax2gShUmbKgRGmGo8VWVMSm0g88tCFp7dFJ5HsSiqfES5rz82
GA7VLiBWiHpnfwv0dGteDZqgHDbCMu6+VtrrVgTZYlZu55MzhQEjEsCtrl7ZCRTN
K69j5GrYOzqWfA67XYY2y3OSR8VMqVb6UbEB4Qw5dT3LvVL7mlEILmRz47FQm9Nk
0RdXe9Ee0At05OaSY4Pg2/HdMw4++c/S/s/KutdFhhK25o0HqEMzqDa5WtBC8Lc7
CdhQCY3ueXl6Xu5BKy5RosttiZ3LH43J6dDiummoatuho6MwKEUDo2L36B1o8eS3
H99w0DSLQCzogHsTWboELc+UKiI7OJgvbfUBb9mojzU1RKk5lv1uYjnbdvuBrX6B
vbx0ff8jSeaQ4YogP+WVoP2t1PlHY4hS4Q3aV1mT30Z6+nfgj6rCHa9GU5DVzU7d
eVSXAI0itBRkK05UEEa21A2LdfZllUCOJ46JKd407BWVvEX90UMV1HKzUt5wH78l
n5HNEUP8FpOpbp7xekE+qkjCB5geyo8HevloYHljHxR+jv/FUqPg1fiPDt9CxZzr
f1L06/ReAArUWdN0QltfVFJ9NWDZTXr4J0Ef8hixQS68CIYSuwdL+Cdqp/JGsKqR
tzRt4rG+3ABYQLCJPiA6Nlv0kXY2uoOFozIBBifCaZ/zGBJDQGPYky+0MzLTGKs1
uKcJF7AnVaLa1dMM0i8tduU8wBbfCAiFhqY4uOb1atna1EVh7oqJal6xRy6+QyWG
DL55QlgpbhK+QCeb/p0lIxZU9GZ+mRdH8bchEVnHG5trUWU9WNIHqDNUMF6oXA4a
TqCE8RpF1bc8qbSvQVyDNz1BmdaN3IZkRTVhtb20IsoGab0WpGVDAgJnMwBx0GEu
i6tHZrBJKAu4iaJ73EU61lkf7dH5hvpEwqKJrmLTIt+XKMu3Tu4XxkENB7Ac7M0N
xTdc5msDGWnHA2lY4oDIV/jm32nv13A7vbkahBGFm0aECLTC9o9V6eJsFQG8h3Gy
FBbpoUzKItMz2hP8lxz4pBYO1uP+P1vx946t02I+hWMrqtLRFNiHM2KJ4oXpJemi
lIWu0YsKl0RVy9hZ+uFYZyIZ0aTj+Ri3hXjMte/Sp3cD1U23ANSbs97e3FNTohrG
lw3F/kDPqX/5kRdNyEuWn9ZRwIp0n07w5KZp5CNXE6spY1j/9QEXpKygR9XVSmSa
PFIk0/2DViPBwrwn6AKadB1J9OBKFcWS/N7hq5NR6zPDMcNNrsSiKQNndGIC1nnV
ZQ+CsUqjI/IYkmwE8pU/Xt9ljOssSTBlyZ8MLFBmn8GEOaZ5IwW+BxzclgwVMqtV
4SHYnyzCLGjKQbtNlZ4Do+zyZid0S+jTOohl+pjXPdocvp52jl+RfROmndaM1Y3h
W5Ja6h9fsJGjAWe5wxs32nctizPfgYyT9CFA8izKX6Gvayfp2RApIqNFwNmPc4rH
JnzRvtPlo5ikozWyb4AmafcgP8bgypn1LT+KrOV/qm6nS8V/yeZGQgkcIdbBWKQ3
FIgoa1dxqBbkhMPRNjGtzS9IRUJVf1Jzcs6lYwO/zAvh+a31eKeGNSC16rZrGZ8z
3rCR1zO7p8anjKhizC2TPt0FHsHqzw2tVU1SaOzTk6g5/iGT+0C2HuFfpr3gcg6y
Jvtml9M7rmEVzHNC4Qv65dnhKtvtG1lfUFbPkJoL5kv8r7TbT3XIkWu+EKr3Emmx
Jr7N5Malvm5PHgduSnBFOwq6KjvhZidzRwb4D67YpQVTIyuBPYbgWot0NqTGAHWM
KvsWsPcOTlFS7LB0PnjLLfvxVSJ7togYawWHUkJXrvgNdje3ugaqNfuCahG5EmLk
hgU8DDRkjivoysoa5XXD1/6QYPy/PNf+QKwKiWN7PWYDs2rt3YrxXkYJnYgT5EU9
oSyW7VJVVU1mMe3NgDjhSyRtA1eYCqncX8TexZbhrIysgzXxz42P4SDs8DbSAwaT
rlAsI4XKg5x6spT1XDr6u4IBpbnKJvlY+WOImDOMXGorU0zPqSpylSwNXoI4Z4Vq
jc/dPIBcscUR4DQ1R08ZF2bSLXzsR4JhfHgEXB793i6K7jJDdCFXIGUX2fu9A2uK
lzCA6A0tBtJsEjcTunFk2xbWuOLrl+D+Id84fdsEP05eyOqLSdiRVilDpd9VyQDR
UpWgxhOyqi+wMuJ2jSd/xajYhctcVh8pCGnK6OrxqAy+JL0TAett2n6dFoiVZ4EA
NDYupsrsinNvwjxWLEQCwISicoiJ/c1614NzWCM/3zst00tGB2NQw0KUqcq+SluJ
8+dCznFXLaDMfvEQlAMcvjL8p1RF3dqFL3W4X8FstOPb2VyAR4S+2+NAPL8u/2lH
c8cQOEDYmDFuijL2QZHewv+mZwHVBqRQcr7pw1b44rRFSrsV/so87+8zzfHN6/Ka
KS7F2Ag3X/GXsj3GVN82SGHjmrrzsorW8dspdx11P0c0WzJ9ijOiAi3GCfNnmGgV
97qkLyRFy+78VjnkfNlapeX1ZxO/G5lgq+IWtbKOUQCYLV2yYQmKbWJ2IxFn/BTO
/4aNzWr0x6dWGHvv3aim0q4hpyN3nwlF6tmZlFPW/zjwGvnSpdjkHvW2meyeACx0
FD9Ffbi4+aur9jnFZhjU9DuDxRWGYe9W1yubS5Q9/XJnodyOEBRfLQElfI47WsGa
R9rx6vP70fmaTH+ixh6Jxzwsox0HtUjfF8zLNlmd67grcfemwOL2Ci1WOKRJlsX3
Pn0p7ClBGrg1/RshCnmiG+h7jOTSEBtLJSKycP+ApdcUEtaJ7KHSMZY/zbYuBEFd
+luj0RF2Mz2Cc9vFxrtvXPhmx067sdgHhmed1paRdMJmYxfuY0qjYIgBc9LBmGXo
ZdMAsFAy3H1YrEmmwDaBu9ZMEIEEoNfNBPd/9yl50c6SDD54UEFfFUn1sKFujf/c
6mk0faB65mJXjV7zoqbXNbQTJWZOgv0cWD3IpVSll3ATyOfzNti5SgGmUhu2fpX0
lNb9m+zmfZ1rR/as7SLJtVbpOupHxi1KJBoCQ/xks26sfkSvrzHtu/STX15qpwhr
fpbrKsF+6E5QMRpIKaPwaEdvPEn1/3J4WnPzv59BZ1TtAyuuRC0jM2jofPvvTYqf
m13jIpcIhueowP7uNH8hqCAOOBNuIky1MXIODshp2eH2MappAc5hhSmlVRyUMvnt
qHuXO21DduYdjG6DTTNJajRppwgXPJ6BAX8MZmOP80NWV5tnp+cDzhA8KCfcjgpC
4z9jj308Oqr2UN2uNbyDqK5qsJ6ca7rO+Se8gdV+UR67GEXNAfHGvrPHW7d3p0nE
RnHZN2FPzcMOnFJjjsIsbqZT3ibJHfx3tfGXB5hDEUjQ6AIvoVNGWWgIvwiwlphA
viR12o/Uh5iH0R9+A/HcD0PJHy50HyeK2Z7lTdJgIGyIEBnWUtf4knVhmfznhcFL
ESAq9V0V3u8+Zt9BB9mlUHLeQ+OgFXzDquJ17oKa3ZgcOxJnIl36WfOxI/1HtovE
8WxobhaT6Gqr4gXcFnl6iCxL8g9Vqw5WWw+A5+3e+WvYGMIBi55WsJtf3zbSCVK6
nadoiOwiq5nxb57NpqYtExb3qIoIjQ/iG6tUcDhE/zSEU2ToyoGD/bhqmVFH8ZMX
97iAcoKc50HHDYxEkx9bkotMmBtVQIl8eyTDsPH9xmGEmlMTKe24J830WJyhT2c7
xvWiLndbUkI4ruFllMMdLYAG72K70m/ST8r2ZKVutj5vyPeTWXNc1qRIFsthw5uv
SWD3AAtiD1lVrliCQT3R2SBqqGwtD+sCjuBCe4QAirxGrB6nfi7bW8Z2V2GYBw0a
TTk//tTCe3bGXDPBzbm9gump3qRECduEPp88/iuiWIOwnIS6oesQibu6c5nRisIw
LMc6+4fbXzF7p+kqever5mznRXbKFeF+KqH6KTxmWBs0pc3K8yYZXZJJpR6BecLO
BYQk0oC6Ui8lIsM9KzX0EzsAbRTo/2zzhFouojcQD29xSMYx4Wkg7vYA/W/CrSZ9
6F6la71wToZpA+k6VI2SNODsY+EODPKBHBzPKDEi1P7Mhr9tsANuOz+cWeAIjkun
d+fwiF/MYqsGKhPe9FeW6/Q0ARX3Cd1T8Cgc+9E+RbXs1D+KQGNuwRbY5LGxqUi6
hscixws1He2NC8982t/bJbX2DDjuW215i0+BXmhcC3L+Ys6cM/FMdcs3fyEUaBhm
afQuvCImabfL4pWv2YuPhj1MdJPqkNOyjel6zvn6YETx534ouum1obRm9SvrhjaQ
YuH1h5QC3aFjbYxu1z35QwgXTHwcwCESFUnTeiBHj1Jvx4jgWJa6/E+hhTxnc49w
xdyhfKoFFA06lVnJEG3HivYO9ndReDMS1vQ4609a1Sba/68XKHHQyCbr/AuaC4s9
TRugL5EJSKFxfPOY1oZX4fLR3XXKWhvG1B1BJy1YT+O9m7xj2L6JrKGGyeFbkhg2
N5LExyYgPn58lkLeYsSI7HtoMNQCUH9sdvYq/SPO5anLHEpx0eNrhJ7FR4DB7k6j
H+WTpGycoOhuG7DftMwXdyfFtc7y6MF3BVI+OsvcN0jUiupORX5fzGGdvyXacVX+
a4MZWsHR6/q2mPze79FDm2u/0k+G2SqS/y31edc64QOSYf8T2o329W+4ns61051D
+KgSCY0OA/r3LPRcaLq863Ixczgalg2JBTQZ3O8qH/NuHDIXNek/5+H0xqBN+PJ3
+xkkhFsFJJcbzSi14a/4hfH+f6XSy0V10qi1KYeYSgJQHUdry2f1erPd/tgSPDUh
Wgg9y4X7R2dz/0QxadVB2vnr0Cngvr9JWXEI7v0L0Gdvb7ldYPJGGMHg0yCIObnA
suPs7uLH9uAdZIjjXAb57DCTAchiRJU1o+nHdFzD+hjzgb/t2PbqDyZP/3EPMHn0
W/j/7PWXcBtE56VwskmK5fuFi9D9k6dcUKbt9u7j9ISh1GRYy8ztonaEgc/AJTL5
d8JIxsMfjVC0ZT86cnLo7HDPUza4Aq8GJDbQE9G3ssq/34ls3GmgKTUqX/4NasD6
49CTTA6lk4XqGuUFs87acige2BfZQGZJlcQi8u1R1cd+7mpsQvgbKMbd9fN/5eFs
Nz/kPeOFriR1Z+P6LdO3fLvCVXCTIlCLzDCggCoWRtWCsaqOBXjsFCzfj8O0L5gN
Tj11fDq2NWUVotZmWM2+iRPnbXTW73JZ/wsEvAGANH6Ukn8ipEELvcZ8NsISdDwX
XEUao/eJKI/RVKX/A8aZwtQdEcJJ+NkZaDPP0BPkM7APr8+oBqXHFU6+dPf2flnM
T6poHn/aTPP9KGZnqfVwhEmuKyAjQ4V2hu/WKrrK96yTr2vpW3diSxynuM+l8GM2
enuINSVCBzUPN2wRoxhWDC6f4I+JLUMTu9mI+6GNsHQfiDjoJ03fDZMDtIxlR1xC
3/8J88yxV6U6WriXma5lGHdPrOU46Ld/iIGassdtHEQOG7zn4TtftPMrFHah9Zlk
cRmLw3RweYHEJkhsi9rsqeSNt4ZqSRQcBPlNFdmr06zICYyI0I1a4qyKoaVY56Ze
ueaKvPiHlAY5uUIh5COxSBtz0dMKVlrISJvZXjwFYto6LYRk18Xwcy8pwVsUzKEE
VFuKmGQG5ml/FzTrrK+WBpV/qeF51tBSmU98Nlo8qirDxs6ZNgO4LYuTKxIaeU1Q
IXJ+CKS8RKwoGZD+cO40uAlYEUtkYokSbJSYdasOkvlLaiWeLyqVc9+YYyhTvT17
kMb4JP+pQ1Ws4PnTjQRIXKhv+nesjHxWxCqKvmbqt1UETCXJqrN7jFpnovgLXDyA
z8r0eNWE/yidj6YMKn9yeG2Qv6V+hypH/PUaMZ3MIlU99zU5RW2wS0AHOYVbsD1v
isqysbOfIu8JxCTjb8sTlcKFWL8xAzJdRtijBOv3PmArTDe/WJ4Yncbn0BErlHrm
YGZ9dRWANydR25byrk3HnApGLQjP8iIyPtYIzwd9HABB10LBzj5m/iBSke6avElR
Df88Ub9uW47L8mO6w1a18moZwqTqd0RwupR2gXNzxFx8G0/gzDY0BCk65i4/rU30
4FKehXrN0MFxR4mspp2LkvtxECRGvaXR6SVWVg2fVtnhX60tEqc+BKhptmr3wDYF
+EcXZbotaXU2yMUCuGTTaszDM/WOwwZbNYIi6KFtTPozTETI0hgTpZFNQjhObyeD
H4FOyyEBaMUuaSXfdTTbMn3s7pjUaVsa8SUDvM3spUH3EhXbk8WpHV6GlzH4Yatv
xbq2VLnEEVRM62ZQSdad0BLs9OhqRw+9mvkvvnQYjfrfnmDifEzUuFcSZbUs/RcL
4GSq4zu/2YR83abFJAbFLgsKpjCr/VgyiRr3MXL0+ZheFat3C1KPp4y8QXaECjrp
1biHwVihXYepNJay/o4EUNjw7apWje682cvtHk4l8ojUoxK7hr2tZCbc2O0oJyp7
9LzyWsUsMKGFA3ctHp72SVF/nYZ5WwxEsYkYc6cs28Owv1D/kf2YW9kNCxcIRIwe
b89qvTb+icD8XwfSCYmXMeK3dOQ5KlsiojEHV/5/l7YLCqBdXPjDx+FNXgy+mEZ/
sy0R1ZvEqXpslAGpOG/PPIqcXtFxMf9BfubSvWcH2s/ViEn4fmLyEBO/QzMQaBYa
TOw6Aiis7jiwLzxpzUTsvRgHENmNYKfI+7Su7MUmYQjhG7+iUjMIvCa8egaD8IMu
q1Co2ObjU4+vk40Vn5gyDAq7jZWc6CctDikE04aJE6QEFxB0AHwWZRNOvDeEDALi
xfWfMsST4cHdE9dEWQAZwskKyXx3febArpAS+UMjIOCnY/K/rby1v8NOkVaG9fZ0
4/RwTATvpqQjuzXemosdbh3rbMlxBzZWdM87UEcqisOIB5tAOtAZlO/o/rz4PYgb
puP84nVwIhs7RUqdwTFoFnzluE8AyQkQnASVpod+vH7XvqI599Io9/d7monB63C5
b+8ibkUIoUwkxbNFoZe5yKKio/jf64pMYszuN8DjIjVovf+OcSRRSysOS3STAF0L
bigY5Z1RWfnoI+9Kp41ZtV+2n/4N9hdG8mhSnSlLnU1pzh0oiqzJc0W28oYMZTLE
MVaB/j2HRZBo9Eilp3y9iUZEXthX+GFGWhepzZDa+0y7xihE/ru8ByJ6PesfaZF9
Ukc3yzCRmXZwNX3EnCJ/yLbMTMOF9zmAh4Z8nuTPsNyULK1vrtRaT5/hVTtMrUbG
l67DObbDBNh8wRp1jzwuJ2FHR366EjVe2paMOdAsniPSdiR1v2837G7EeRqyZKcz
y4dEnQqXbX6LqCcIVzEJdgFycO+CahMEKkeEmxT6656wFjO5MGruuU2ljCVpzKZY
vEnxauX0s6STJP6BVpNQiqPoqv5KD2Z+zmv9MwXFj5zyKFV/Fgo/MHbpii1xLdLQ
BfLgJtl6t8MdzCKmIk6hR0/Cwpg6c5C9K9cbzAYMb58dm9glz3W0FwSTkdXdLGcF
pvUqB6dV7MjP6zzod9urK47MxH3fXTdwuCTeBKzCR3/CHlIklRBKFkHCKzmyIZHb
LMmnI4LvsAd/NIlO8u3r4136T0IOhErFItAoVF2BqPcYxHJRm3ooftVdiVJADsRS
wnbcrDakeB9ZE3zOK/2mS5a+4VyYHrZ3QvycLg1t/g0eAO2o0gYKMEedwyC9CMIa
Mj05JgcVllUlsk9or0DwpaH5AkPkGihslro0DA0AagBhZjmklqCwA2CKlNqsx6bK
9sWT/Azrv8J/GDb2sk8aV6P0WH8Xu8mKTYoKKd7iTZ8aw76I964G87C9tMK3Ly+J
iZV+oj3JU1RyRYj5J+/TbKFy89bywAajO1G30+zes1A0y8MA3dX9IIVAsDVIhzTM
q/pnNsXRkGuPzXDMndYAS3hDiIcF0FVK9OwWVTf30wN5+vcyvxZ7JVoulIFACn2R
JYNIAARVWYmtEtmci3zo5qrEWWuOV0rmFTn11Trqk0ZT5O6vr/QcYQeM6ck0NtyV
zBCvOzCaACG1J5Sb+HU+a6kd+GB5QVeqSmWvfoELzN/VsJ0ic1r/oDjrxEdhp5AG
/SnwaN5JZMJWfRWPWh749VvG7y7b2mviaTVR4hrosB9vRBTpoGtjbXXZcxeAUYRe
S7iz+0vE1B5N40Z+YwRFM+ua4nWHkC7SZSXFFp1GAzJHZFzTghsZzXPwrWTGGcRv
FUSoHZj064a6zWl+pHkfe2wj2zEhv38Fe7KW8IjXmiZigtAAmoSxNvcLo4Tm82Sj
njZxiBIDGXcNKvPIMs6aCQV9CTOBYYCJT20xLZO5hWGWkU8hi256eaEM9dQrZEu1
RHjUJQ5SkEKRlOnoJL8ckBfoJWMZZHwtkA+feszfD5waybw8ekGce3jWsVfHnTXy
gerhDAg3B+A8hQASCGN4UB/8I2eSGwzgncm8p2XaPKNqZxC4a+Gz11EIhjZQAbYR
AfHwIsXiduqRc/ucJG4YYXVuaGgN7A/L5UPY3zOtIcxE4JpRunYMvOAppgPbGzu6
LHY6++f1WeotoTCU1tA8dMYu8mnx5gPH35Zvbcu64SjLKPlHPpO9S7iUWe1tyOlO
VBnnyq/M3qWBIKhEK3HNuSbtDxcUJZ2jVv1RwECw90WW3NSIdjb0F3hfvCv/N1Y+
vjgRQWCXBY1rejjbpHvy5CvS/hKYiUmj3PDF9O4YkJDNkhofmzpcxksk+K7Unl50
QUy9kGWzQH9heq7khyXTrxyhtyvgyo4KupkquviT/0uQr4TCRDi88IpEUayku7Oj
EjAB830PYnv5USVSKTevbGZo8xyS1wWAM2/KWkDbDKiFbRF19LYEATxCwZSfF0Y0
nb4QzwyzEWy4fyvcgmBH2VtfY+tzfQ/xSiBmOMhw1hJUZREuiIFskoyYnBiAOIIq
nOnBEB6U86HxBaf7bVyrkf4jn9AX5DkSmHMFaOseYOCm/EBXOAE+U99EmFsmKBBl
f4+pG7l6AZxX1K0f3dbYiXIeCGROF0bRaM0NJrVc2KjWB7EEuOOXNnXekohHQ71d
t5gifbnfQYsI+UZvdI8ejwBRhhDfs0zpQErG6achXD2XFPTrQxHF2qHCoqj76yDA
6JoL05ELPXjYYEiT6xgiwSOaUTA+ianuukxYK1RNyPDmDO/l146y+/AE7pbrWWLc
GKT/gKd3MyB/1LfEdeGHsJhRaCToaLedJu2hCzXX2OYJVZBCyYvRsZOs1DCUol7p
CmHRGn0O4V3O2maXMNHO91xtWhbtGVAqBZw72TD4vi9PnKHJXZ0MNpshvHb4hw2X
qfrNbthLClruLnwqrjGf0Z14mXJMM91+YpTlMrCZtKgWV3gL3111rEiTuC1FLW/8
UFmJI/17HU34ZCBMAfgo9q7tXoCfhWTbo6rB9zXLqn/t9reNkbvC6kUnBQi3E8k9
EW920YjvobO2CIoCWTO5YIOE7+ZFvLywQSailm+i9P86WhMlXa52A+0oupM/2LHw
uUcbuuvCkpkSHXpRaFFwjgyjx/J9TLE8BPjY2TWfdTXBXgMI7TJn/U+7yefC3BBW
0Nm5PwA2FN9gsrzzrx+i6VhZasBJA/zK/qyTdep+2FcEcIfdrCA+GxZI1QIMEbAq
JNfavbbL6LxEnCw/KFcuY4jAriI0KH7cj/xLpcNSULJx5HkmeMhnhBI4EkjJMyZA
YMlYHNzzSekHmH3F/UPUihQEK89MIT9Edkvd3R3XZZzxzC/NEv9R0T0RXfFEFtsw
9TSeNG6C6kRlfCrcpLCoKdBAbDu0R8sUVPEyZju3g0CCBct5U5XGxnv3uWyQ3L2C
1hNEWE8g+sLwRqgvFaJ5LNLB0dXPW5ekwEWRtkny6t0DoIeni2mT8Lolo5BFQ5Io
buDv+YKWk4Rtp2UyfwzmyaxGSirDIge7LAaCBRuff98BoLSn3OXsV5G+HtsM2psM
M7xhnjnWLqlz+W+Anv7ZIUrq0XQRfNCWG/ycXJ9P61rUBKWMVRFm/XfSrqmQ8Zau
drADGduWl9/SGyjRprb+J/aa91Y84p7SRW+0GxH/r9cIAgEIlB1OTKYl+5XiO/vk
/T4pNqar3Pa28vO4Mvj/7rd+ZTB3ZflY6DytCNHRpRVbk9/Jy/7eZoUrN2KoxBPR
0B9wqyBzILKbacPKvmBoe6Qu0ZeCzj5IMANttM4cYcucALNe3OqqZjJu0hAYmRmU
3h7QQsmXKNLaVI4WdIZsCesoZWMiEMSf6e6UZ7SjwvZL2jOtIsUcClPr/J6XtPQw
FKn01b9AniRRppQyG5qKNGmNw026oHRQA2E29Oqkh1jA2UrIhyvTr9Fmti3J0Bws
2+5A3bmlp1bpCqQ6txJpxrYDtKP8hDEOp5zkGe96W1Xmji4Jy3QXL4EqK3tpYruT
TClT/pGiBtvPPi2f/HzRURkFb/D2HYqc84OZFxJfOkzano8VPm/Kp3G0kKaMk2ES
Hqtuqcf3/hlj9UcE5cY9AC0vGurKNMgg+hdDO2/iqmFc2siqJeHQjZFKoZaBNs3t
KA0MHenXq/1qgiT34CqHHoP5FjfKGMcZr9OowwIG/mhvuRDDzKcDv4+jgEZo2ikJ
fDcK+f4IS9NVTTgpWDhu3YbGDKnETXlqcZIBX1WJWbGPnZdcwXCrpbxzFKPkwNmx
WQem+jcX8SGJKNwCfnrdmQjP3Hukw6ui5l2ShVJAhUu6AZPnH0K48CaJimSky/+U
PmFp0UcXNSyRi15+c9kMUp4UQssebM3+lVlWa1M5uB1ur33c5iPqjEclCw58oHdF
tfWFnS7WmXV7IJVF5Og5OKcxraIqYKPn3L4KYnKVvm79TL9DxR6a/8dPey5N6jEU
/6uIKkYOSdfL49XQzw9BZVFy5I+Vj5GW/nbZNv63B/wnhtKLIQxRdVRw9fFXcCIm
G+oLnROCoM+AMKNRRlNME7rOMqSz2r7RZUG2B2BmnhTEUZmU2aeAlnjgNfTmrydw
vvDwccqp774kKFAz3vO7h/bpgyQmquIpTY4HjDeMbpamMV9dUWxe6g7Z4TJLqJtH
NBii+4TFR+jFusC/+yWnRSfYu9OaoY2RqIsZsz/j6V9tNyMi4DpyaMVz04WDwdKU
yQbW5K5gNcR7RdTQwpL55kkGlMyJmOflkM6YvWpbFZB3KEu2TAxNZzoH2xglDL95
uE5hBsFpoXdHQwlQbORj/JwGRIGtFRIdSQuw533VgdvXzuuYjKkh1lRfCQI8lw9Q
WLkRJ7MtTckiukv8qwOSfRnfrMwVEkw5JwPb1D9RwIBVHzWPw9rDyd3diQTKK8nV
V7ketVNB33BTdMzfVaPven9ZP1bZnyzSmm/3tjl3mw/sxGWlDNdLIvkIlfelvMal
aCm05niww0+mLk94O4DqMFGwZcs1wGlOab9X5mUjspa+xH6Lg22GT97YuuRIJZbS
3WEXURlII7nRuNY2CHMnYxKjrokO4l3cJTEev3lgvORQR7dB0yPZYGfexfm+rqn6
SV2CdblE4DW5PdY5h199OnHqy4n2woVjECTwvF5VEiCwcBSgZmY31CDM7Ajy7zXC
Xeo/SpMb6ketnIXBic3lle9Et6cte17B9EW0urFvGHjIx+hXKKLr7mVxnE7zZssg
+8g65ybXNGHjZW2le6s45/9PiIkjPhjqAlqdI9LXofZSVAqb9eJ3+CfZM55maZef
jJr3jj6fvMIpUpx3yoYAnwnD2ZgujpkUCTBl7xNcr1jZl3oE0X410DGJghyo/kTV
GR2PZP79eWvZwQZc5YS5RCLxo0LeHBp+8OgfeTILcI5yLVSkeo7ZsAItnkBJAgmX
Iz6kOf8w0W5WRwMQZjSQtujAHvEgulqlgwe3Pg7T/n0DriDsxa5dm1PGhU5ynP4E
7sbq65dqTR3TYsf7RwnRhUDDGSX/Jtp7CbZ4Ub3KRCkKk+ukOt8WAygxVvhz/BJD
Hyc6NJ2qR9fJDzYwWH/OSXGS1czP047KHURDg0IdCwk62TGvZwDgTPmmrWR3gSoM
R+C6tvP6u/tXxhhVrtdHpRGEAoShZeODd+LWvG2dyjLiFEHhIa1+2wh9ZqEDAkmA
ss5WHcbt30bo7fhEasOt6jyh2F5/BgbbP/M6FC8QFd4rNTSaC5yk7udcnybVY5uA
7d/saAGIqgikwtU18vqabSKNtQ8z++KNyL38rBghpirBHrVcdvT/kn6pBMMniRzs
KWcbanHrnoaoYj4lZ4THGeRg90MzhXGO7FhzVa/Sqn0wn0RGVDRTZYO1KCYHGxcD
Mh7xAWX6hJh/tqwl+HJWrHrOGeDLEleFiWkIBnzRbgeteq0PYVWQIwfsnIp56LOs
9joAlOMYRUQUH5r57cj8Qm+lLjr3E2YVDDPbMY0vHJUnZuJ9baVetQ0OJuEkMtw4
JWKmMK/isamW6al1mygzjlQsQUZtpAc3uenFCDapbZvtQbwC/kv4N0N8x9whiZFu
UlumqHVRO3XRCo4dPBy2cK+KhHvVjG0xlz15WfpGBq5EPfyDJnQQmOrvsCrj079X
Bt7u9X6vM/zadABXSeshomtvYFdAde7rclpGD1o6JP2XPJqnex9yV+SbzPZyHhJw
B1xtlSdNJXP+pPxtbhM2rtsOYCs/Ba6IvwrCRA+OUIClvuiLxTQHeJtkRBdSqprY
bwlQV5BpYawRzkZExdAto9SspJ12zygR95U9mhNBcYnwRDCNvWXQZ/XDo6yhaU+J
Y71/KGVeI1bv56yQ5Y+k9hxQlqIH0uRj+jxTv3qqJpqaWhT7H8rkDl51N7CAorht
NuX7wVPafh2D7P3+qY8UNY+h3qDT6Lvm4lXMGNVkNEf5RrLEAEl3jLwqnaLpIUsK
pLJ7LSDGqSbY+HcKdu2JllmlzuuIOwCXyd8+Qu1PHFrdybeUKr+5jbECmmP9mIBi
w8mqwo8jqftYuop38PZBTGAgTfKnfepA+Ag0+bMSPF+l4RkN8GeuR+w/PW5Z4uZw
ld2cJFgmfyCkXDk95Tc4Dd69hK6D2DIAuReYYFebqdM2Q0O/nSiU895KakE0nq/6
5AaBroiHvy33qFRKjmeqFIqjUo6k7A+bxz3Bzyc5x31XCySd6Cw2Qp/d6rAwUFQe
kXvDM35q6jlZdLyv3GEDEy422IMWi6FabYrCbstP8OyxNRITGjTLpkzcuhgo7LSu
1VM1DZPNVsMtU1eeYUh3pc2SlbpPE0X1PuPJXLFjXEEjFOdxI6SshJSGxEWnk1m4
2XF2Lhr7TmRnsKi0lO2YWdQ5Ix+a3GZhuT0DKo+s4Z+SPQFJN5azbMvIBJ48etzO
YYEUA4vo6zhjtH+YFNKWMFmW5giDL+2SqFr+jzwdWedwQwAU2G4+tT96DyS6d7s5
vFEDT5IPdjrHdebIuJt1QqV2ITT2oTmYvXSQU5rg9LlOyqecSn7mIajO4TE3pGMp
Ofr/nsrYDWH+XidHpTiQGtTe7cwYNXLEcPVxdzEyy+zH71f2YeSk5V8Npqp1eTK1
tt4UV0hNc7gahnbVmJPGLBkr0MgcEVJYNkadf6h3ExFaOOms9Gzjka3ZQeZ3Y3Sc
mZYt4PHyRBH8tSUZCUvEXJ0n7r6kd6hC3ApJSscquMYwMcXfXp+zlXDnnjhnP7jQ
LgiK4xaZ/J3KLdrNCiq/AEOi3gaoqU45mt00ijkFv1+RAVW1a7Pc4uNCiCsecwuq
AxmETlcuUbWQN5arTg3/HURNxhBkXZOkUlavK871tuxJXmrfGZgU6nbGBeit23/o
HPlhL6i5dfazaTrKCkDxy5+tuOP+Ch5TdkUc21MuL7gGMDeOIUuji5rwmdHHqa4Q
/1YqK3ujbZjOrfYLUV+eszwhxoerUndhsf1YOpQ8WrH7Hd0mElTy9tN8ADHi8KkN
76vRXquKDaZKfzbxdcMo5w1u06DEB4jIvhzQAyfdF3GeurjA8HJVgLaRvM6gEpGj
rZMOMBU6FxVQi7dXJwuKqTJu5RDm9B5BOyzF3scEi5ZpmLOg4Au1p8dClriDTgcn
5m3uasKYOkg5B8EBITqUx1sohuQ871OCVt+lEnwiHdrnwRCcTB8Pj3jABV29/UdU
8/aSgRaUnHN0DttM/gaW0ZrLjbmhLGjXqs/W17CMeNFp18hcdGAhOwSypRJwTeBs
fKgwgvXUcdv0A1SIeREPpK205nW5seZDeno2YlqDtupR7fB4O14LDL87I6NDkHUf
EGSeCbnRAzPDjCJtt4ZBzCHbBU9Xs65JJAHYSwTadlbQ22v9BE+jMxnQwjY10Nbu
KYjNqPyZ4RlHBa3rn9WvsNY08Y+PWJqTYOt5TitqZWesx5psKDzqQiwTe1q42Ckq
Catxqd97DiP+ghN1Kz/lX3ZY27wZnFDNaTZgI6egbPPZxego1t+ymMsMMv2fuxxt
zWrgPTpE13ZMP5Z+soyYSvhxk9NBiqOrEIXPll00ED8UF6txrTYuxHPZ6Q6rF+oP
8ZR4hgiRTochu+KPnmEOY6Kh1qMuePc+aAQPnCb+KmY7oJ17SnsK9U3195EE5Xyf
3gWgQkg5vnQNa39uyhJR1GS8MjdXBlBN+T8QR33XOYX9pkytRE1cTgUlnvwKaXNB
6emrzdU1ceSkQQj5mAMH7XvXLkhNXCABMt52UweSvHy5OKFsIxJK6p1Oq2wfPDlN
DteDHreuF/JRm5BLKG1BMeOciRq+2iJoi+ZWoZxg+1SBHTVhI+jvNlKgB/jvzq4L
JIkiqJuusR743EiKX7MOccSJWwChQ1rXaiUFhnq4D0NJ3MKrydRzWgKbqDxorDzP
HtKVMy63I+QIpIxMQLq3k6vJxaaFdb318cVCS8fiPYb00U/OY/Zeszq2S4M/GthW
CBsgZRG4jcPt47H3XktHSMHikhbMIbS2kKdp+9SlEN5Z9QIWHAALjKn8ECRLwmwu
WY/+eB/+rvGFOCv1ImeJhHFq+CQMkPqCiTxY7iETs9Lk5dRgLebU8vkLuasl/ObG
9C0ny3tEnPB65zZiYNBE7e03mGV9OjIzITmZ6vpeB/7TTGtxuKkGea/Wxoo41Chv
LS17vNT9jPT//wRUZTcFMM+E/tahw4BcpqnmDgSg9TVMif84ScWvIoE2e2SltlgU
+y0dxS9HPhaCk0/nw5vIlYHeJlmv+zgkgJtIycKQLc7GjfkUee19raat+9C+XGcO
nsdBQ7yY3IFcbWO3a68EmBHp6p4U0wHgBFPuBx4hWAVxAk3pQaEQEB36TWgDkZVC
NtvVfOzy/263T4cvzmsyHcLobu3nLkNe7Nxh4YbaZMjgyqnMV4N8uyUnwaV56SMe
62uZaoaBGZw+qEOEqQWo6xcynbYLGzHs04ZFRjROra96ZlFsUMhFAvn2fJA2Be40
DXraUKKQ/dLe3TuD78h/CzK6c856VI/cNVHTrrheOvnqrQxdi4NhAyNvYAgDTemJ
hYUFhvi8C5SXw9an1J/u5+Z5L3HpnM8CVl8wVWY/wGGLsHwF1PBsKgDYwQoCAQXc
xIL8DrikEnH0+L0J7mb4fusxATLIsIcsq6xVm/E9QqgICD8weDcUrohiqlKvh9cH
lJ2DzM0vdlXFwukQ1wj77p0jW3gSwX9+KDLIUCgFiFsuX0gFF4LkiVkCI1KTWVIN
gPEL5ZRMVx1JX4etviMECaHfkqaPHb+I02feXvLUxBZ8fwbwDeMJKo9o468BC9O6
x89nIi41ZynsO39BhKjCaVjF/dKTjNlAAhNAjjzw/T9VVttFcVjjfEi1+xvCo1qs
ztRDV15V8nF3xyB0kfK02qVOYHDhPHRnOkTYh7QQzTFBE6exY3rt4y1L/VuLsEqo
xykwq4ZPOitMMUJ7JvaOZLu4FotOjcx05sHcvbLUrtDTadB+w6XxTTT8CemPBuZf
MrEiQIdkjJfzzwd2qB4kvThZ/Bg0xgN/PC57chW8krYB9N5tPeEU7z/IzCl/2miS
BPxK9hJSSIFPchRphBqyFHMD6ryaCfP90o6jRCWNTWs6u2Dg9dnMNwTz20FuTfeT
tFRRm3A/I4UM9zFxijfDEBSyboD3aPKzjSf8w/xF3qI5risCmxU27N2MJHvFCkod
ZvNqQ1e6gt6ZfHMrWGCYjFBe9Z1TJtAmzCDMO+6gvrz16ylYKrzG4SqTOFF67xye
bGIc9HLJ4JBgCBXYNsR3p+ioOPFZ0Ubagt7xenvrDh/V+P973i3Wktm17iEBm/v6
hc0WQzgrnPulhq+8dauw3yJoHlTlcGQyI7P24F8eAP5fHNuw7IPTYB0XhwsEwbWV
g6DcyiK6lbmUtVY6yXxKGOEf7afXw2HQUnoRxBqIArx1RcFtn7Pi4FjVLbqvOMxY
tsXojn42xCg2Qi96buE26aznNnXXoxHJJqHX0fMRhFy5DvhmDy+XayiuxJH9KyRe
HVxe/ZcLq/XwEAlYlwDVoFa1FFNSS5DyeZtUuKJgbIVYTyR3zDsdoRP8DFHRKB4G
pLRUq/RKVf/2JIYqoDAjWsLGhbNoXILUHbjl4v7g/1Ysilg68IL2OUDcQs4L/A97
ZG/pV/JO43rWuDAGEsWx+6lIl4cSpHgPLxrw3SqwR9ZN5WeeNn2FWy61JRQQaMQQ
FvMvuZRBC64o75tCdBkLkV89uZS7b7bUNi3nhc5sabqsHvblkUjO/NER28zYmPJf
oMB+auzMkvxpzZH4oh4TNQQn0LJkBS/HjvclgdTv5TzFd/BhEgwrnBhnSlzbYCmw
ulQJiVs4o32XZQP7t6GCu10SooRx+KmUqjYXQ3L7HJQ2aNRh++hhXJFJ8rtzlTaC
oFaLgiuWZlkrtdes1CyzDB6g5udtzttkIHOZXhVryP8auiAE4l/J9QxfK7MyehyT
7Nwv3tU5ioYVTgQGlrzflkddfr1VpSxfj3fZ6Tf12TSIl6HHAvlGluaoFM1IQzcH
Xbq5V4FFPxRN933IGFqYW9kegsAqHKTdnwK55pemRtEmqxN6XGn2pUSe7zMb9I26
pW4iSTXdgDCDJb5W3FoSnIdo4p+nN/fWRAJnamIuezluwcBUYNvoX1Go/vXPJjhi
/WdNQK8lggmrNBD8S8b2ypN6e4pSq2lKiAaMYEAJBl/XAJbiPJgKVMoAaLUNTCa6
rLy3FndBIfn1qmnk7ZjatcNt3NJrdx/t8a3EvuiG1VFLKygE6ZilaJMGAYU8UENG
k2TPXwZL82UyoAJ7cSXmQsmLdkHy0C/gJbloSAhU8rPT+otPws8Itff1/iPQyR2w
QZGtpSDTNtBbMASINg0jHsfBFJd8HvFolDnP+SG9SU+RW9H29qRWVLwLCmP/HoBt
4OklX85SroImvvPC/UMBFncpb36l0AHb9X4tsfJzwOHdKcc2QeF69dKLlVmNHIWL
gX9nZYdGlBTlsy8a5XoGh7Hp2P2GGXZednRrR2XJQMHJtnTUyD178PrFkfb9QHUj
jn/J5ZGh+lvh+B3X5gJ6Y/UGMfZ6e/Q4nUakiTz9sMYCf5Yx6ppZDHv2H+xh2mZM
at34HwU8pPxO//RdfokhqSaRoNm2bRcB3mRor5GZ/2+6XjMI1/O7oN85eoSMu7mP
DGsnr/+OIvW+oEtvFEuNtWI8cBRpCkOGCPlQq/dcggW7QsASeaP7NoTdZcnj51vh
Q8qgpmJIRE7pjQuAGWfPn6J40q5MqypO44d2/cnrbrJWNCRbaAruYEtrRwaw3ek9
Bd9xys/1l1+wP3YpGK1ZvYgVoaVYXq5U8/MrF8pGm0lpq7ugiU4sRtnMo4RaESqu
O0cyuv1m40O2uoxTWohPHAJVS/CqxkTviKMKZBHN1Ds+MjcvWBsoRqUmw4smr9OH
t0DpaM8TnVhTMXbJJ05wJl+q3Im97zVBp4S1uW/SaleJ7f0T5gbCw8+HLj9Mppjk
mQjpFwgLq7pW4FfjjQPfrtj2nU0DdQrfAouFuH9G/X8XpVUFirkLBftdPJoVSX5L
IH6tvsg2lOmeCl1LnKIOQ+BHhAcDL/k9O5zrAtKsimmLifQZF90cLM5hUiqR/v1Y
N2jXDTKuRilvhA3Mm2/Ql0gpuzq965c2jgNZ4jgW2pccsULzkY3Ke9HqgwR+ymCe
iAWfQy6aVx9tNzGlx1fH16p+xmhlK7C2293IiNhh8e8MOCGWCLMjxqC4qb+mORVJ
TW+4mDz9r5ezymyZbgxs2sJZ8x5BzMmw1SIfAUfVHvD8Dxm8MmxQUiYan2yx/oSp
pdZ3VhziWuKado2CMWSE60bI+tPGY5CuFg3but/Uu/U/RkRSDxDPM/vHi80IpWy7
m7bdzcBlMVw6Lygr0kjA+bG7QqFZwiOC8H5BZef8Q6cajVSySBVBavEr4vYuU9oM
9Ki1kDilSkwWcovffaBHp8OwFk0AyTSnKFRjlcFvsozpAG6rXF9ZqBNDiYiUJSeq
hBaszFmjclEy9fcftYEEgQ6Uyan3XlvsGLvu6NxK2eVfTuHY3U5A3tA9QroAUC4A
hFsE080HciQsnvQoEtshF/sUAYDFQ5CpsL24MMw/Qa4bvFa+3KAexRZExdCwbXzG
7bfMykQf0vuv7RzAMYKE3phhQjDvBHgmFVhvFpBjoigigZuuT2aNiTD5Xg4LCWIF
w533jozrY4l3wmR11W1snMq90YCxHEUK4AM9cD9ro4SU8+OqqCWCA5L1svasJbgj
zciJf0IFKsB+Xt0fgVqtBPaGrseJpMgIgPIgeD8r7Qu+j1fcEcq90utPxysio+DH
vCswwIWMwIM9kwXTmm2C/Rclv3sXJNsmR+bTpUYTfNH51/2UTuhd68C6Jx+Xlr5S
aJseySjn8CSz58cmKNrFob0ZU7t9SJJjVqZV5iSs4wFTG2XoNmvf4m1/Y7gJ85li
MQPbOmQ+Ax8nnfBqhFWvRDi7iVHo97adR1ckMQomWEUZP/QSfjePoBTdG6JUsi+Q
jZmZBGSoCXQqhsNy/tS6uZwBi1aoqJ1oV2FwwP+n62qk+lEJ6XwM2jLclysWvAY2
1BSKWdpB11ys1BajUpkLGYpvSGx0HSGAfSHKISDGqVpC+NzZ+0It2GBnsaYBu6vJ
+Ew3H8OxDCKAZzv/kQr8AmuzcU2ySwrrSBzXahsiGjkUiI1vLBEwZ8Gh7dMfBvBD
rq3mcj56kTTfa/WxrJjLvjbnW6BBdqqp/ppSY41PEtLrhyC1NF0f2RpzsTkOtUwb
ZH+BKiYUcVESsfmLRfIcVDrnLv94gBkCvY2C6epHRGpCMMOZZtBQmvwyg0+wc5TQ
foPa1KcqIssZK8zP/stT+kbyS1Eyuk5d/9l8dK/vpksMLymrH5uEjD7Fh3i89Rhw
VOoiN56JkTDbjX0JIPXyP/zLzUq/+vSbtLUak2CY3AjZrzJHbX+/6lhnMR3FOcCH
cYb/+OgcxVosinJVKHq6hQ7B6+6mZz97qfF0W67YdlgKzDIjSJuGEsF0NzJdu7bm
JG3IOSs97n5nP3wFbEbakKGFnenzfzvmCKb6BptP8rwJNC/GOxOJN+v6spaMeBjn
y7qSh8uxIKTGoP6+LVu5BWPkL44kwfucW9ID9kD8Ld66bOydCjGoQ9jBUZL6E1Ew
A/yg0EpSLwRQHGMzYCcdm9pnu2Zh1OKEL0wnavtu7b+i4B9r0RLBNXYYr35gE0Sh
iiNwoub0NEFP9PKuR2rKLgL6S4nh8HKX4cjHHA2tkANNYrpdDkQ2A8ayPeTi6hN1
KYMjoW5AxNV+ZAto6tjiS0toZYvye1MFVuYUaJwoWA8QYGUswvVtnJ4T/qSf95k7
GerGwRsyMKR84eh8R2KoXR066HHt+jt4t5xJsnSp2iGR+j4RvF5D/M85ue8qvPZW
vCerzK0Fsy+PjEY520qTdzwJZwm41Y2g9WyLSucI8bwNJJkSoAdMykQFH1uZk3gw
Z6iN63rv58ECBcePn76/mfRKAl54lqO6W9iUdKK4mCZKIW62IG5T5FnGDSH3n781
EjuFFU+DS3wajGGVZA5zNKRjXYgYBkYDdouDC0YuLThvMQkYigsAEB6SzgNVtgD4
x6Np1yUoFTOf0ZchWKFZFv3+z83v2HmWZpAijBXJ8cfCkB5nwHWy4WScWe7+P8c9
Ao/ep90908ZiO6q5w1n2LvsOjnTcaEoD6sWEy6ogzZ16iPJXuDZqilqW+Ta6sMf7
czifzgZMlQdVAvCCi3bu7ChloaXqu+5IRe+EeOhZN8M2S+zr93KZo0OZINaQ5xgj
i2SORQnrSx/N6CSpn8aYuPnEPnO838B9sIDDIThzsQWVeQ6QbZH1eq2AR7c4kA98
chdzEkhbBOzM9N21Z/Wh9mMIB/gyf1plyH9OsoO+Fj9+K4s3N/mOUA/FLJ3EdOTi
fdSCTnFqSHy0eWED4MEQcy6802/pgILj/5NDdQwkesU=
`protect END_PROTECTED
