`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPzeO/n5+iXf3IimLgAoJuBiEL20bH+wki3AhA2KB2rcvqtpD9SEh97/xmB+LVVl
/AhEu8wTzQ7nkEEteVCkgsMkMQQRAB1YwoWc4oITxICKUiwz6qLVFH1fArShwK9p
9vuXJX2rER5MRuUn0jwzVwTvwKFddc6Ur8zJcNA4GgqOlwW/WZkr9S2rX5njpYUF
BXnqRTbmLh1Fs0XCvcQhAAa6m6bdVmv+brG2HmifrrNuE/ymhhHE6gj3BdHUSZhu
rMufPO7RYY9U9PCHPSAhR60FYKcNwchUlRrTG8sZmiz3l00fBXfeEnE5oeuZyNc/
c4WCad8Z8GqccUafvPjRGo4vFPzWDkRRpRHQA0mueh8cj+sYnrAxzTISSGBSNUtA
6STrDSWxm4AGJ8p6DGHCbGoInWAiJ01liId7496K/tB9z/QrMa8IezD1Od7vbHZC
Kh6LsRt0TGE/IQk7e5tIzxZDyvcIm8OZBOMSOuCRlI/iaUVvfZ1ErvPvcBtQjX5R
4u5UsXAvraoC/3LcYaRbMzwDegoIk1s1opVfLS0XB+efkp8gbBXGhyr6yxhCITgZ
SFHpYZFQyJut0WY0gXOW0u1WRaJQEhYySdjwz6f1HKwg1DvKcroLG8WTXH5EXk2Y
Mm16lFtYr0wM9y7PYlHTrVdG8VpAhJJ7br8pYW3lxWZ/LxcZ9PxskaKc2cpLsF2x
7b8TXrvDPFa18Z64H9JdqHQBVaxtFtndCZPuXLCQzqoqHjpl51eo+Ugez94XWP+i
yPytDrUJHRKecd8JKYWHP9zPc3Bx2s+mc+J4GXwDG3HHWk88yOs9jo94rU/HN0Tk
BZxJIdYNKG54j26CJM73jjSZpJ5AuMO+pTFgkK4UvjZZ2cNTQ4zzv4SmU9ZaSGYH
`protect END_PROTECTED
