`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCuH2krfNqxj0BNEvOyQWjeJTZ3Jwppj26aOIv5FfKn2CP5KmQa2p2dTY94l3MsZ
57XNA/WCRZkNojfdFxz4K8+gbyD6dARHnfXBJ5VrWXlf53xiTIgKwjXglUyMHjl+
u/fEclzDgVOrdeLIBxNmE6MQXJ0IIZDe2VaVac65HsSqql/hPWi9pvEe7Slmgdwr
QUmiK+20+Aq5gcrZc5q2s5m1xPfT9NSXk2otq5W4qy4R6VYqBuSctAb9Cyl91CAP
w9ccadhKlsNnIG3+7CZkjv9Syw+5LhepclIKcGivxWtdBk91XcbTF7CSMp4xZc9y
SBjLe69liGn21fdsD8D2I9nZ4vHpInXtj1yoApFkjx9H3bG6zLigsrveoGLd9gA8
jAwjeAzhul0jl9pFsm2ILTs5UMncOLjWQy1RthCbxdLxth+IhyBe77bnZ4COzjYw
r/JNTSwyU9JB3jvL70gqLoFLOhxW53KsQnWJFuZtpJPVMFho+Ru8vNNn/Wks/sZf
UUTPh55XEYIX/yO5+xTJ5vcVAEKVNLNsygdJF9080Zr64XCjHdzFi4h3JkBkqDy6
tyxNizKJzjjLomv+WHfwHazD7jJfQFrxYm0PYe99wH7xFYOageLAR7rMW0L1Z2Qw
hNKnNFJYCHjrscPLKvplnpeGj3HwUht84gYVHDS9nCGCGrvPL1shMn4rsPXyUyB1
y16hxiroOpFQVhbLPBv2INj5JHQLPO5VbOSnOMjUgaTLFzjSffl3GHlgzRpKJEcI
hOFM7l+CoGkYr6MjkmUcIl83DlhcqarSkloxgvpt5Qh0CYFMFy0FHacGlo3BOPl5
AI0olqQLkLt7+Jx/awhdam4jvrI31Qp4/xlOzkd6d0Z1LWmgNreuPq9ZOwlbaObv
rmAIWuBMOYoIxmo9XkajXkBpufnTHqjPwww67YdZy6eOaVd+Fwvzp8A8wyIuEg3B
nPzzxQZIfUUwRRjd2Z0FyAfAQuM0L+4aXCsC8U1nHRCLbzrVW+ciHYybhGA7Vk/i
WNmCy1jNYn7+zmiSWbnukgGkt59lAqDQYI4vH8ZVQjBeIhRQjryf2vleNzDy161V
X6/ObH/Mt483+DKVoP0oKNtAiMUiKDoiY0UQHPkhG9/fJs21OfwKl130NRM8c7x1
7MNtaKcVIb3vzfYpEVtxTIL1u/h3ftGvDfDvHYUvIOuGIzg6XpGfF0fT2JoBtQ6Y
RfGsaN620fmVn22zptiHpbG2Kbp5Nbqks5qvqwjUCi87cLtgBjCxby55C+4XXS+t
1bx2tzvI6vM/NVwSPUiCLlA0vZDWJi9wGWSxqMGUnIJeILF7UV2LKyuNdQCxzcBz
6OmP2whek8IEJeUiVpVVMfSh/d8j6NMHU7JMakSvkYDN77jcizUze3FVKKNHGCzo
lueCnggvBgsZGlNPX0nSsIxeCq0tIMPYH6O5qisdmuxHCroRP1DsgqZJi/jANQPZ
`protect END_PROTECTED
