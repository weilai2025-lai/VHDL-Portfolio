`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YXC+zJjTjotQ4KMPgY5BzWEZ068oMaGzXcdE87AWVIr7Iov1EeVC4BP6fzRKi1B
tHiIIoM5Nz5kFhFPfTnWMu4D37aYM/L3dOGk6wC8i9EhQz1Zie+bZX5RpZCfgqfC
SiREnQ8ssNgzreTkrdPplA2iaOkr9HD7CRgizM9T5f8U376q/TANewwTmwh+GiZ4
4WaOQg5dxMC2ODPuRJZprZCX1sSwIrQz+h75Yu9kDVtKQa3unC85811PPWlSzWC3
7JkHdaLgFDV4ywcx3YkcS81FEsqSl8mn6Q1xGDpVx4UOEOPSBZPweMSFT8YF7aon
CKbP+hxwqCsHup265q7JfsPuGMZZuFehkMT51NvIqAZWu118jDbZLHZ1ob3NYUVo
c7f+97lDmeN6vy8GD3Ua9rUO5mjzoR1mfVd/cxvgzanxAYkxoRYFg1+Wnmf338e9
3DdibCNdapzEPpJVpH4vKQ==
`protect END_PROTECTED
