`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zKc365vt0/Fb752NvhIQkPgwOrKtAJ090mOiuM2rxuKGbbjQuxNnKFyKAd3BJI7M
D0SleyKbzgsGqIJgrGQrkiWmFmpdk6ZlCV4Cu0JfJhfXUMrH0PfODnCDpxLI5jEA
RMrabYLjlNiR8+gbqJQQ/xKJXwOZbfrHnwb9nsqDkfBjA6+E/mr1nGvFtsTwuqLG
03xdGCUi7MchAMcaSBQH8gRUUg9y6tX4vy1V10b+YmpKPdol/NMAO6JF1MDc6U1+
z/33aq1TJT3ti4aRzZIEeAUCYx68CzYLtMUZ215i8YnwJLRtKeKF9rdXtr8d0z6l
7o4UMYZWtpuDR+E0r5EOxqJewZKFBkcnNL7twDgFpqdE1NHizEfoRGRQ0y1xguo7
YHMw9YkMMstn/U1Ixcc39VnlDJJ8H0WBAEW1p5WkDGJzqtvBGQjwuFGhdLE8kCZp
THSCobvwPEIZDEBpqvqnzOeNIsuisIsOImSra8PB7j+cXxBqD0g4cg7GAv0TpgDX
Gevi+mgUrNiayOllliHGEuA9BI00B8Gr6Ug29gqVR62F6NgtouQaiO9Tc2ffJN0N
7hGKChEYlHM/6IWPZAgI5sIy0dETqok8BUsEdwku6Bk9InCuUAPzzbnljPN4MFsu
B1eiIq+fO5xklZZ9aPxBM5a9pjtOd+jyqzBdwIy5gjql2Wc9N+UzcqIjD1G20+47
nNNWHoMWu/XnduRZa5iQ/e2i9TOHn0jmDMm+zfrxRaK26TC7/APcA0TQ91GF9ic3
6F+CjQ638VmDb9KZI3C1S0TLAB/JXCHkr0twpT7FsM21Nq+3dHgiBRgwiGZ/SoQs
i/R+vMe7TpiIHtj6ktNPcuiLTRKoBavkdbyV0g2KsKlMvYPEfw++2ixlXonkX1Bm
0Ec1W+OORWoCqTK/Lkmkaha3buaxW6t9P34NfdzxXjEZP6FeKUNfWbbGaxCz2qOM
P08EOOdT78/B58jWXnlNCsgxjXGyT/RVgHBWON790NT6hlxB2/xVRaKiX7Ev/MVv
lRXWR0mL0IltPQ6dPG3uyKNkFOsB12yj/7xFislzRtaccKw+VxWq6CN9OpSXN2Kr
EGRNPFilKIGQc7xWuFfcnojrJsQ7hpM98AHhDTyXUxH2NShTa3omzgVRR3/v3rDZ
e9XSgbhmq5kP76C+u1fdj7ABFM4YXOYJyZZJYWjw4Xj5MFr0u48N6vMeHwMyPpmj
d8+MUbEIbeq3RvQ7ooRj7u3vtlaXrt2ZeNVGqebidRFmCdICsr5WkI+E2LHHwtL/
1q5grA5FwOaDuC2JJ8nzPEVioa4BA9LfvgSSk64O1dyYDY0LOk6uKLnqWXYKrZWo
jOPCd6d5iI+vdWuYkLgiTX4S1BrbSgzOZ/hG4ulHVPuRvVLW7CskTVbBZX1PWqLM
0ipjtG+nTvyeNS/pCMqfMUAfy0j+AEgdwJIaqAkYE5UTk2DHiTMkTkeBoG9ZTecs
+j09BEP069fz6BSus8d+uUI+HqKamWGn9kg6zhDdsUmLtbQOfGfLzL1/1olVDgik
jbgDSwYKJDNseGLH5oJLtT+kNS3pr/gg1CvRhEoS7yrWRlT+lLuL9fqL4q7XJucG
WFF9AeV3oaqCdMRr7MElQC5Eu77KJOoLk1mwE12FP12fuQThPlvtUzx44zXSpRxx
2pJcyeNgSUN7hQIFD3hDzdFs9nyDximqYB7noDrFEbHeM7ULIisIhPhl044KRQuR
0zeEh6lS0IGPjp9L9O7AK6p7eX+3o2ZCJiQ57YwoAegodGoxLp6vf0KWFyVmfYoq
g4g1c/ftpWwGWUDGub9i2XYEQUQuDPqU90KcDRpRmhUuF+ccz3SUr4K9rBUd4EVv
RV49Pbeh17rVV7ybtKtW4Aa4D/VqDDjmSJWiiTA4HwUAXW07JVcxfyTvXMXYel0D
qxjU6wWVds0ZePzjrAENHGQwUvxmZg/BXC+O2yQcLq2FfdSXUEfdgiHJuRNOp66R
dQEmoJe2Vd82ZMA6G045m/48m0SP/mMgkFcXnu1iPM0tR9A02wVibyAt5Hi8vI5/
QWIWOLqy6d9VpM93nNcIBY6U7pfqbLOxeMcGFDq77LnG0ALzdVL8QyavSJOKJJHG
tutCTqDLvuZE8OR7E6/vSZUOGHWhIjpW71AGxOHFtk46v7d0z9mepuWZd+pYcgvL
fPRY48lysrEUCCxrXsR5ndePD9p4C4irq+weHVtWpLTltQGXfDj/zYt9b1LqaGUj
rIRVYm39M24I2/6TOgsfws16YHWbdIiADOXKm2pmWldlmTWh8DANtaC+qvZ1p/Xe
nWLSArA7ERqmLJDNXQmoDmtU410KuGz+pLsuORYh4aJODtXnv2HHlPpLr5G2D2q+
br4RHWhjmgEgQ5/Hc2TaX9tylRpEr4P/TSP+Ezn7zYJ24gZTaoYZVsVg5r4mWzEc
Pu0td8cS+cm/n/ffKApOLq5dHyyLlnW68tnyPSX/BJByymff3PUZNADgOUVHU0B9
OEHwaA5JpF7jd0G3H6Zqtldq8l3cz9b2Djrc3oNsLHdqPmrOenpRoum6be4Mbe8S
sNoKOTHq1TakGkdqVsYc5wRbHxTCKfjpEV97SdAb2fu0RMToktUKymHuFRw5qxcp
dJ2kGyb5+QTrXWrsK5EFYHpbmZaZ6sXgPej85PMfwubQt8RWEOrflnHZY1nEvfUw
ZecejaYTb9G216JOhxThp8uRGTKVMQTTw5IwbsDo0sObc2SaFoJBZqRsxtEkpH7I
1bk6HtgESbYVxSQzUsFnnLSqpk65J9xn6YCao3e9cyVaPDrm5T/+oDjxgufgGHYm
wj7AyE6LX1xUWWVhq+R4geOMpDdf8JG6G94bqxuwUQSWjKyCdoueZbRCGEywxN6n
vUnAAd5uS2hX2ljfAljRZZfv0prXgRCoA1ocAitwsaLwl/4bthrYqTpn67Od2BFd
ZSyo4q1XXkZequi2QSSJ1q5TSd1/g7MjFdRDk+NhhnVnM1S/ktW8ruVaj98JajnH
89CJfDodpZZ1WZPrFZGRItsK+ypaojqeEwV70TGQC+I1x1ItjvueLpJfSxzI4N5N
Y3dqEN75iU61YO+S5g9Ju8J59oOlwYKFZHa1XBLnacRyJU1s1ppYnPkSvKV3pppD
71ftlnDOfoqOgr0Go/I5s1G1MkRhCeYPAhpIvWIniUkw0M92cE1fqZulxsdpZj9V
oDiVjAMj/Jaqly6B+my9LoUlBdJ6VKiCw/poONJJSaqUpp20jPYkDxks7UGDglrJ
O5Q9y27oBN+7xtAo40om+DPIMcJKKkeHUdFpb3vazRnxXGiOfNx/lXrYZoxxt9ZG
FB1gmAlyQMeK1fktr8VOTM0jm7GSs0P4aJRDVqelJzacoWawD94AfoW6tPfvsCKc
UNAXN7idOuKybZaVxqnZ/O4rD3wQGh7sGc1YylAnqbMmKLSzqTl1EbNrInhvY9XR
q64qo4g5sFO3TCJIlYEPjZXBXH7CRtVfwTCqin6gakzcNpNuN8dMjxojRmoSMq1D
GWXEBsjlBFz/qn38mHrwAzaJs1weUnE82yLBB5mbkSi/3z0X9NjqbjjtPnXLWzni
vQ4edAI5VkTtYvdGRjaHBwi6y0Ffu4FRlLIJEyumAbpZPTHwhe4Gl4EK3EOWMWVz
xZnLDsAYNQVmn75wEaxtqVNhjmtApD9HaG73KWdM6YhvI6trC2D2LCgIokYNOEul
vyTirrYLD9rN4zqTOC2UcBG3hrWA3c4OUKArc7D86ij9h/ZaOcjUht/tEJKUZdEN
Hu/iSuPcPwDq303cHz3HWDEvO8TPyB0BrzTlPTvwBv3M2hpn+hIowaKap/uDkjbj
mZJ+rqBoVfLFhWx+u21Q/zKIlxMsWLSJZzz4YQUKh9TZNOXGe5WmWSMWszUjlF3K
uLlcGucdSgGWzw1gvZT5LnuZJFZds5q3GneL8/J5gj3dTVaJ0KVbcuUgSjaYpUlm
ATRQKDrFpAnIwq/Pqvd+aFoi+1yplUNiXUdVrwcbRxU24c111YPYCYNp49EKMk/q
0YkRYIy9Ogtu/wVzkfk0Hf0CSp5wT8xnU2Y3Ds7sBZ0=
`protect END_PROTECTED
