`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwkpWP1tTW/qMInrzrexB3Lk7nMSLKgDC2Kjdu9D2ICun9mXr67uemWeW1KO+7TS
n9k78IaQT/IVvW/ysM4FK4KLhPwD52fmqMWidqeILbzs6swPgTo9CCtOEqcmOc/w
EJ09FHQMSQhC0lbm3rYLbaTj5doNhe7CLwSNn+kuFGSgmVAHq8lQxjPeC83Pxnvv
2bfO+SvPbMqwjkjvSY7y7Hbctoz9cG2W8vEe0QCGpi+J/MjYjoHLA5wyooE2ALVN
FD841YHiTSSnML6n9+S2zIYDxihIiS+Kz9tu7Aku432GLVEs+8zXHkHyTqka/g5d
rxUnyEOA8dXodAz00jy7ZZC9znf6ZNTF0xHJMGodZAZR4Ui4vpbAtCI6wroM1wng
+cp/mtfKY1CGN6Q9FKgAbdEFRIUpHCTDjVHbuleloB9tv56I6wdX7pW87FbQieJI
s69Jer/c1bAbD6JyYEHWbv45psaM5mqf4WGWndgW+2JVpJZL3jw8nEcquORkkQSk
XOWlLkVnpUZxiFj1Qnu0sL32hBokUuF1YiwavbbTrFCoiMICRfVd6gmLi1bNIhVZ
WlgRjCoH7TOdSyT/8QDDhXKFWs9J8j+VuFErXpbU1JLbVADFyIohmDKTnEtnNhrL
PZgag0hcu7W81cnxAq34Q8NZzTn53x1sln+ezaIX+yJpQPq/js+SAou4Lv/N1YSU
Fcz8yBgKpkKr/MH/RONVCQuakpLJ3mC+tS+8PNRm8SYdG6G5JIdBLyQ5mCYcBQxw
a0UDS49fminjPNB/4wC29r1wIayRgQ4I86sagTRfTYiF5YVpqAiOpP0N8gkVcyxB
9+rHwZHKOkB/Ffgtb3snurFvkBpbC/c7wyfXLDZDA2/ksVUj/Mww1z3qgZtuwIw/
PX24kNr1LNJqGvBCCD7ksisDz9AwDrQjlUlQzyUdZibi2G56L2oRt1y8MAhZGi/q
3zy4bG48JrnkElEKQUWlEbvs07MhqDZ74EQ8zabedDoRYtCj+B2ZS4tH9kZZ2TZg
PNNNN9lRg8sR22aWUbaTATZrOk2WKkqx2b9Br60+ZODpT9pboXP2Z9UvfPGzTbWb
XrNzmG5Nnnw/faOf6UTPQkoSuR7x1qZrkl9xOd3JkdGKRmBEyzBUB94/lD+T7SPl
JbSloHDNelTMdRv+wOGm2MNlRy6HLAOIKdvnZNYJq8gGloIl74CPPi6G7JFEPx7Q
qUGSVvNes9etrvDOhxQ6BZ0ouvqhC1ukp859jZFPoBMC+7jY59njrXuBBQ5YKI3M
CBC4D2zD1lddD4E9+46Zen4zIsmfXqa5lLgpSAzsmGXGjiyTDzb+joBX5PQEVqIv
z24FlYxs8K/P6QOgNgtbbrqA7Lg+AJBd0U3xEiABfjuci3KrzBIx8ZrxM5YmdGXY
Hwh37ShSQIkjyW0ecorOIXTErei40Ls9GAcmiJJANFap4SG8qoEwrKZuP4f3V2ik
ZLNkgTVl0msnc4zfwf6ZvMdUTctTTASGccaTbVggWETIntXTPMwVSRiAYzCsUV5l
oLBUCmjfZWqqbqenxi1vtfvjd9SfuzEgVCZcqBvI/QtToTIIiHNxjVX651wRVFjN
Eo4JvaTuKrEnmqj7BobJniumH4tqEvV5Y3OrxVuLd3rKd82AEw2bht1IRLzwlwpR
iDOxiAJem7QajCOvHwCaOo7yZ81pLMYGfo+0lCSLx0r5rdo2kOSDtDfR9ynrpFmB
H5N22+ezHN9ktQ8AocR9mmGnLPd6pmeUf1uQybeBCda+9oehpFzoRkRGGmEhwSGO
APYB6t6Hs+j9nxrn7j32gdhY4JfB1+ecN4rg4iK6GZhvcULy+MzHMfIEKr3U2OQt
Y1CM8fM/aI4YIpe0BXGswTHGTuQ/ZwLz/Wyd8ksCpIO6xYyfWkC27P05qVrPCr2c
XyURgVewFClvXOk0FD490ePiyyTeW1jWJLhjqqZRqS/igJanw2p+W0UEfhA/fTaC
JqZMOYg8TRBs5Wn1nB676qOFq2b7tNCSiu83R4yZnvobtlnzqG1ewtJd7OVs1y3N
CUNJ2bGlaKErXNXsg54ncZ11RO3p8ONxLn9OlNmwYhUiUI2S2zRZM23CynQJzRpK
THFiBwmROZUnXrTFAGs2zVdq7OPM4D3UGOG5Zkf0mw+ho1JZ/KhTL5cYc2mjCQXF
9HL/612sMR4BP/rNXBxR2gNbQDIuowc+qrnJvBqVyHaHftcQxeUHdpa6pZaLKTYc
brTs+DkIVtZxVrtbXSnaCInZ7doz7fuGB0ylcT72kFkV+q33kdceThaKqgtnrpvV
TEvM/VOTGDS05kU+4r5bURc1IwV+xEqxHQ/79tsAQmlx318rmtHV+qJVTfs4ZJ99
R99hZmwAV6DkcGpEyuVFT1CTdvC+ndpcysJQgSGSF+430SPTsLBn08P8dkavpKKy
LJ+hNYU7OqAJjiWn7q50jVy2a3SRYLy+57UuZLMrTJ28V+ZO9RVHSzNyDMut9GoT
LyOH8OndWyzohPvfNdivfVcwXfnH7YkhLVjz4KRRkTa8+JQK7/CP0nBZ7X/SVNkJ
RErxu5iypH+fqLaK9L8UlkYIrJ8yCiBsKgRuwoK4VyhjIU5o7xFxeOqDv080rc16
v/Yrr+A7yUZ8rDvPYrgchE8JDpY1Mv6T8YOOR0cX8m+I9PKMFr2JtafwL6yeBmZi
V68qcpv8DsKbjVP9d25BBH1cvUnOxj+ri4S0xWCKg4YpSxnM7ZYGPymkQ6XNdix+
M0zGMKM8d+8MUmz8+m7F/WFge3cJcSJZ2dEzmLgT70pFUoqj9HjNQaul/7YgXEBh
TM9IwKb2pfcNzJJR2PfsgkCIdhhF+XJVyti1xqqCr7PAKr4jKzave9NJfifxZtN5
yN3Uxfn8/KqYAFiF7EIq/AZmATUQDfzuA80dlBzzKI5DPZ9Pw7CJ9MxW3zjYrVYd
/CrpmwSiSe+JrZdGRnPqJWculuzlnUDJlHbBzsi65y3SDQVC67rzJ+HNl/5N4Lfu
3LNje0sTC9wUd2ginunrm2u9e1++spncBzNwE6pdShEvmf3C3Ud+M6Teqr2K42PR
LXkT4Rzy5PhZMyKgS0fgocwos1Xl7sHP0wmdy0Gabxa7NFViNltr8cFDoh/N6Xtw
+oPKMMCB+Kbl+L2Bxx1+0/HBu51/x+8cUCMwdDYFwc6K+XkwcnuPtLCVwvUqhG2p
fX5xKYqtqh0P+aN84bk3OHIWFr5LIkYj6rO5WlwaQTCmNJcRUBQUzTHV3BJNyIS6
cpSTGb3SICCriRawA1CG55CVS/yF314Ss/auB6TI9yHsHKRW8GTOdJl232gbGTdj
IAi9/qbJm2sxSRNq263rS6mq/Ny7NXxCwI4Bp77Mb1XMHoPY7XSgcq864apWRzrh
8NfYZOrMSYFDgpTIEEqsPaBKYK/hZJvNU1Vp9mYPWOcjSH//7CfC7+12mcKcATMf
ECJCE4mRQmd3YdfN3WsK7AgteD2Ct7loQiJc0SFY8Yw1Fk+xFUHknbI6siMqFTXg
1Dww0SOhpgBA4NgWVlBpN8obKopdjEGX3Ccu9QVJ1rVvkewXrmApXX9OWFqbVLGx
Z244ovLJJ/SKhuCzUoxFOwpEE59nCcmigy/mIIPQ2LVybOXJz80MjE7+4T6Kvrdx
7mpxxL9oZ2aI4EDSCnw3/1273JsjD48Hbgp1izWgE5sTk+8cCu8QjB6CosSpESH7
pOX21yLdXsKdJdudYtuJpMO2YmIJkL7u7pw7EEH2UuYBau4cwq0IlIzsGWcGHDX/
x5aESrS7XONXCbxf/OvkxUmMvoX6WXz44RpF4uhBFuGQRrmdU/7wTLPCsCOKQhpQ
Lp0FPXSazBj5bkLVX0LCZRfho5zyRD0RIN6BdQCpam3Ir75+0uH6yI2DTQXsTtH5
4g/OAZ+5q2zSwxBO2cTUmY3TNcjo2hVCiHn+og84O5d6gStI9B5ZTb3PsdWdqgOH
W+47Zom8zoSGuRf7d5Ip30EqwYRD8pg6wS6bcyKlYz/uXETl+OiasFdXD2RqXsO6
VHs47rjJB9OANYzGLxcrNh3cmZwa434H3T9mwhpYjswhkXVmU/y4VDCOod7b2qiy
I3SCcYscRFul7Pev4Q0R3pXINqhaGwptMrbW6ph1wCg0/3QgeUABjwNFsiAm8s82
1/qafuMAICqbvoo0nCg0+sInorj9PiF2PAoi1zAeUHvI/HNwsTAqWYBdJwFRWFnK
7GDaWua3oAS3Ud26ERIjWzANAXQTuoUMkaAqc2n1tg5Jf47JUD4g+J16UQ8uvRVr
ydi9r10j2fFiLCWRzu+UIINttqBlUBWFfcctUWSosK6CQZYXuO3YBP3HkGnGVc80
HjsAwNQX5BSkJYGossJLQanJrCAuXaNIUkZ9OgHoSwR5nNoi8CpziHHeD9MuLYpV
7ktyudjawyauMmEb0ANgsvCW8fdYIYCUjImY2bnC5c/TOi2TEV6o7kFtMnl3T2JJ
wSjtI93GZGGiSHiJVB2IPHjhAeImgFVFtuRwJPX4iCbWpv3RIHErgDupjSSSZHEd
V5xtd88HvqxZ1CQMw27abAwCVQF+lWpfkmHtD8iLMF6RO/+eVNP9SSw4HrM3/nLX
NrGn6ExjNWYStWmuwYwN5D37TszXAKEJm1urqM6uIP2SfYHt6Crab9B5LAvXdn6M
gU+pNwyRauI/tKr0FcoWQVz8AK6j9kV9Cnbv245ed/6L3lAAlObfZ5ISMXCYQoZo
WzysqKYykfEUwAGRnJPwMcCdciCdIfCYPxCYJ1ZkCAcX/To+OI7PfPBGn/YV5x4e
9dx9MFEVO1Njhk2+xscBl0RrIVcexgGPsiGm59kMmU/hMKC8dCQC8PTrodu4KofG
pr/RqJRJVNidsQFalx/jHOL0Yoolsf0PcUTroTp8hsRl6t0vrGp0/Ck0eJPbpf+b
LwifQ3JtL8E8JPk3hmbH5uzxTXE95HLqEQAcB5q6aT2YaxMgLzMz/1NlcIS7NM/+
JAKsDcV/FXB7D19XH0JKChla9rxVanDINF76AMZN3txzHtu0AYiuLoxAZ03a2DsS
r6Ss/huF+d8xw9P6RSz54L8BWUHUJNIgEL+PjS/t5NySBg3f03ORJm6xOocSK8qv
O2OjLOqLKb3qtALn0FOxk3cUyzd+SU5RKS+JQUIaBJFenCQtHE/vyVAIdMe+UjqK
6lx/m8TChjhs2MrNKLl25yQ25Bz0z/pQMoV1oOe3LRofWOM/fIRPfaupnvAZLmKY
JSWuDLsreVCsrmdLygxxkrH6YxwJ6dZ1gr7zuzogIEknBGZGdrRVo1VTTx33A1HY
EpiePVDwCXXocxvU3B4iV7WX16EYF6YTEJJK4UOM7S2S/553OlHPh6+AbanMpSZm
oRIILidkzMlwW/LkcU76zEUWAcsGub/BA2SInFWlmW0qbcmuuhumZbZivSZGGFfQ
gP0KQZBNB2hBAYSYK7JdhSEDPX6q07BDFsrVvGRp3Rrzll8xlmsj5DYDtTzj6iZl
/wIetGPg6S+bYN3J1qy5eIA3Q/4LHRsc06E1vDLXPKQk3XBXDatXKf9WZUAIe3Tv
aliXxHVpufjApB4NrW/oTZEYr8TrCeIRUTSq+6UUMJMMfTwtN15/z0e8XxtI+YpJ
ehZ1SwMr08CZ/CzrbxaLZcN6fX0WSquk9KjoL6UrgH6idkBPYGeb6mIUbPO5Q8GU
gYFGADx6g9b9aH/3eHO91HAlZ/JTd2f4d9iKuha9hGdmibH/tEGUVriszDuM/Afq
2ZzeWP2JIKkyABn1YHoP9LGZiDtrAaeDaNWKg9dV4dWhR04iesMKC4Py3LFnUzAL
pZojKl9Q3QLzcE2KJAOkCM2YPyJCfNlwqvtjYux1PuSzfh6ed1ppvb9DNGBDRP63
EwiAlPdqVDiHy5dFRjvpbK5SBgjQgQ601fsMpub0uLIsMb0EZ6Otsfx94WauXl3k
/UiaPKCykWj/Td8Mg1zM3VliuFRgNRb2gDmi8CGO/uM=
`protect END_PROTECTED
