`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x54w0dH464CqnAfK/trQygiX3IQDVQYT5x01aGHnssdMZH8jOB/QrDNra2BNpPJI
zTQq6ACFwfnhDIVJk/U2kxxekzUk3hikYD9+Ow+nO+ln+GZ3bApDYSgLb76Ndp3M
C0FQiW9fEq9q/CxY0Y94IPGdyLQNkN5OiVvdgS7QggE4g3A5EDn18RDPgJuh+uET
C7hWAoYtp3RJCgUYLYGu5qGuMqfUIBAG96uXc1e0zLf6qv+7OGtfCcglI0171cBj
wED9TTkEF6Lom79snrNyfr2lCo5mEpzNeEq8ELf4G6RhnlqukVIjDLPGDZAqNbTb
A7m8L+L8QBamFNC5nTI1Yu2IY14MFRjKHF8cBbugG7yLun28HZNCZ2MluB6LWIDv
mSd8W7oXdWgQ1gsS+fe7ZHOJQhRdAiHPhgdraALdTpRTBxkREdHS+UdDUJn03U76
tLy00deUnY6Ptac0t0IKIiEcwPZmZhS4XGSEVKMEOanVNC8+vrsN9dgk2QqeZ8xp
y3j2skNi/CxW4vHLtkGwoWBARdwQCtKxqGbbGV9ltEaZYhq8wSO6HMyN2AvMYPJh
UepVF6kPPwe632OyZbtuibdzHo2VRRTRkmhbEynL28a8WQtxdHiEK94VSJXpWwiL
Rhf3W7SRPD220Yd1KhLnr6eFUf9FcWOvB8YViQVq+oifiUiV8vrLkMId8CJYWgG/
cGVgCTHA7BFKXuOk8m0AGGyCQVw9YVz8rmLDpegcspCnYyGmSg/XYnAbgFaweI9D
kYEmbHNxmk/p0W06Ev8klQ==
`protect END_PROTECTED
