`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIKU2IfVAkpppPhobtTUn5yK704jno8rpaJvi0GJFBjKPZPmfEejSREwnpHPVjVh
zSqmQi0QYqSbZV5vECtZcNQo4uRRS1uJSFtF+/o6in7q7qR45gDEFMWSYd6MQzYY
oDXEQysp84wXfooG+kbhNERnT8YIBL+HlXSfs5wpVv4cI0JSTO5FO/ds/9F5d62V
hhkYL2PQWuABjcNWXpl7YaNR+ncJs3Usp/TiGOxnb660LdXxhX7sB/71a6prC2wO
dLwU6NkVtwJCA+brMet0SwmFtW157nC+/Ug8wumIqaud/cwuCy3F782ptU7bcQCC
wsVkxhYRDoYbxoeSLNX1Pm58r4XVlKcRqHuYpqr0JKPfky6MK5XKOrkErcz9hQ25
lRYzSqiADkVBtY2jMg+RHcl7RljaOY3HVY5QAFdYW+OSJ4uH60Fs31tPlWp1JhrK
QZtWpSk3NmdN8KjKvt1yJ5e205PiRQBLZcITQIYNLhAA3AknA4Eu6i34LBNdSS3Q
t/fPiJ5vKzcD9VsaodArMtLtUSIPY8/Qsp7PkesH2jQLjGJH29CXrnFg6bgXdmC7
/HReb+hgOm2eVOLe2GujuiA96jwvzimR9XbnOZ7ZUy9Ry/N4n7ZiDIOCR/WAL+54
txjXPPqjU2eCXPhoYUZhbB+uhzYmSS4MITDCqMcSnekyqxHv2gwvoLDbYtG8hy/G
fvrW4G50xwZWojJ9xQlZ8Ab36GHoZ37aXvoo29oCXqFvIzUCMm8WCRcW4kvJ5BFd
DYxo2L0mJs/q7yRHCk6eL9kO9GsCZz3GXB6kMk6Qk9BFnu3uN2Rt/hRHbIvbgOw3
MftJ02FC6TRbqOz4yE1HMEDHuGfh7HT68miakXmQbSjEdVLtBwVjVBErWWYE1n+7
INy4aZ6UcBjNN/WTTCMRsxqSPERfTp+POtjsu22yzkVlha1ay4RrK24acjtArUPt
Sq2gvxzNRSqiGQ7xu5VnT87XZHNQ0FYqnBH2naj1gWLSARBpSCYDmWXRsde0gHdV
9maNarHwE2SjeVe+J+wfKELwfyVpKg2NHK0TUci27euky24tNDMBCttN8rz3lYgj
qfk4PxeiqO38NJiwFgINPUWOYZRMDC2dEJLMdiqE2vHewYi0TiScCGVgmDbT5go6
V7kzDICs9vedjR6lMl+yiN3Ci6wunBLB+LcGq3A0e+zyxEXunZkSZ1R3qD8rVXAx
XRwq+1GLrSklOgUq8XF6G0h4ITE7vhK+qTfwKfJFWdUCFx0mYYWRddzYWdgfwORf
FsQCWN9Nsgr9iULsJ4drkuo90mradu4j+0DV4i4BRwm+eCOgsU2+qg9UlrL9dxIA
6m1v1UrQF3CoU07Ru/KZSoa/VLgAusonQxSmWtMoTi6njkzCafO7uehpqMahIf6I
3yg05wBTKOqCfQ6BVP8ww0Quk+xHSVDT6NZQDsevEjaLstjryAhZ06HNewkkbVhb
00KL9XqsSvSsCxD/CDy/gFhlYItDx2gVuq22p6SYUKOTysZDmhEQqDUECJIOOE3h
Cj/jK2e304D66ML9omo5OZL9xNvAxG+QQ7IbtHd2XJmGWHhU7XnTK1GGh6RiJYiX
+hn/OX7avXXv4EBtpnKUPUjpX9FrgYPxJ5R9EsHJmldTuoTippmggh3GgihgexQ4
uLqAOUbsQ/DLPukUnbZPQDXoz2rMtZiMScjvJMUFzXuBJ8/Cxrd1PPEB91g1MeI3
uAkzqaGluzAJN9pblUtPG6SZ6SVVSVq41WLg9K5XIekGF48k58RFk1XwYvC0RHhw
KcYSxmPAcNElzwBKLyRhTcibJD04LC7eut/1joTBfEBVXlYrW+QVaah8siLVseWO
CqWTYeU06b6x8oRqJNVNsQSkTmRdA94+2zCbRm5vQOma20z4s3elEmLFwKi+VT9z
Enis9A9Idd22yhim7UybghvNRRQbDrnByGZsEFpVRUE3rI/ptOD0QBP5qaWqo3eP
UFGAh3B/AOkoAYM3mQOySwpzv6hH6PcRKYwbD2jNN15m+siOnjWn2YP9sPll/qxD
xTmAmadIv97Ij3nb3peGIJNnTVmUxPi+od8NFMQC3lJIDGLDhDd2UhjGkDUw/2O+
yJljMLygU6ubm2gu7Yk6b6Cn+oCv0H7RwAWHv0K+giDxR9L180NZ93SPkTiGWAWY
oXyRVq1RAZM5dbYVt/pwbfXALkAdYw6P45XVk6cqNdM2BMovnzJWgqzy3k0eLSCT
ujxQhgUsRB5l5pZseKBpCP1ReNpmuk15+5BpCVknphDYlHbWJ0r8T/Ie4A1IPgE6
hQHmB4eGC1zKjYYB1l6GeLhX5Yyhsie4qnTRysAHuHZJmUfWEWGHAuy+VfIUCfC0
0jE1x+6hY55rnqVE/1QQTnw6vpfVncYKO8QEZCwnE7lGcNYnSBwbBebCtn7uk5ld
ZghEy2VEono0L4c+JEo4Nki6alxI2oC1p4DK75CE9X9aIHAyz3QWWzNHPJVobnYS
qSh1v5y/PG66PfJSw25fL3zkx0r4zURj2suWip3GHOGu4cNrMdJZCdIrOHm8laH1
6WH8j5IDeml73Ys6wz82B3Y67VXCf9RsF6Me1WfbXEFQieVf/kJLzINI56apwF38
DX0iG+fVkeVqiGCpWkqYolDsnYQrYoZnhSYRgb0mm7a9Unm+5zXMYzEfRWZy8j5I
Nv81d4KtNk74Zb7EkBWRn3YL3hgrM+D20tAT2BnOBxt6GcGglIw+Ucf7gaG0ZAnK
xl1ol+ZlLSuZl2y5uo+gJboFbJ5bHVJGcJxRSfFLT6bV/jPDjbLyCrPS8OWX75HP
c5QqdYAqFI+hY37zbnF+0t1rIaEpUCXVuz0mccwb++yltGml1a6tJH11qkX2nkpL
glftOEjGDiWGwWvXU5FWgtHOJkIZBYnLBfimaC80qQbjv0E/PWoi+23yQIPdNlV5
ylC0KQFvNed7bi5ad8w+j/j5jordmrGN3FgdLmip8LEbFvjd4l7+1Mugq8B9Sa0e
s8jzFQXizJ8x6Vm6/G71ATV1jylAesdL+ahu21R4QJVNAirxv/6aBm+UW+Q+niEh
hCZiPALsSO1BCLlMI+HBEnfC3QvBln3zSZPcVdSMGihtU1DUMKywhrGSNbrUkTHH
kL+hS0SM4lwiS+cAkIT6uDfC1w74jQC1fKBXhNRsAix0uMcoJOSubljxEucKd8H/
GugCrQnlowJjL7fsHy1BN5ra4keAepHGbaTXTMkJd1ziASKGuncu9LI1WkMcybqY
5bMnf3qhdd6f3Ffo9V4gDVEEwq/u82VoE3n/HS/H5F5u+rx8ILibvBegxC1umXVk
ls6Tr1qoTsWJH6NZ+EXwjOeJurVoUXU2Qevua6cuAQrqTWLlxseIH1VEPZftZEon
pdK/2BBCB4ji1Nf0lxcHOQ3S+7H3+WvYTaZm8IYv+990PwYMI6gtZ4BINTH8SXX9
rFSAeIaz4gIfYsl8hSKZT8PU2JOJGrNn3xZj2DY4rZpjiT5Xcchm7l3Ug8Iqx8kU
vCSBQT9S5PcL9YoumZpIkx+ZfB5BFGkINPP8Ar2Cz8zehA3Nv0r84lIm0C+OUXVl
eRJu8p2KUSXYZ0iNeL7aNjHi40193MPYiLH7tknihV8UxCsJfZ296r6kGSdqjgKj
m5BqW3y7iO9DpzDvNEuk988cpq3+EOT770k0NHWEjXptGz9lQ+7SbBDOTGPOjSWD
EEeXIEqq6dr2X/yYkm1vht/HetxjkDqU2wFGvMfk02c4kUHRMmb3TszNz7FphQdg
HAwDN86DAfcbcOnXo1kdBuDi/SsdYBRcPnCxvpAgaaXN0tIsY0Gz+v/rrfNd2evj
kZ4ptjB7RRvHqlxdNHr3ohEzlquTZoBbmlWQVMZHCXI6nfxIiEBenezUBp+F3HeF
bpLmGPU3NiQ8YfD7y+xF6nGUsJLIMInrfbPFy50iHvToNEWv94OtlsSc3s/GTc6P
VQlNe6I9HMjd6iT9ND56DfSbJlRwpxPEIiZAHBMB0Cn7bkMLK+p9yisFe4kQBHqg
M8Fds8K8s11eBQ2ajR0HUbWAtmYfMzlVR8jUiPCHVDWpvKfeHtqSFLwrJBfXGANu
v9mU+fdfJOqJNMFpsnuzVT5LPGZfTuMCO6Sn+YoyKRFfW0j9Lg0Wh0r/B0bkASPN
Yk9OMWVsmfroKv36AW4iKHqL0sridXUqwy3jSBSrQRL7TZ54krr4NqWayoXe3r8w
Vtikn8Mb7JPQPQUj9Z99q3GvVL7/ucN3mapCUj8RYPAKVgtQAe6im/4UyAs3MEbR
Q8Wj9UDDUsujiipZXE/LYkgHBCAQY6AIvHQiFUIzLvdi0a8JNY4NRUb79usH7GQu
uepiXmFJYlwnzu5alMOa1mgdpxebADe+fvuj7fbsV1TYVWOVCmWRKxXd/cOhb6eo
QJlEQUCUO1t6TfcGlBOCpe99EPoUbjQDTrt1hIimAo/x2lUn+nssJhr1OlwggQHG
aj5alTPX+Z6qjZYoGG2zsR1LK26bdbx5Inr1mnbDDec81dNmDivyBuzH7XGJt50w
sWinotSn0xIiI3UhcnTuCbrQM4tH4waA0Gggb01vQ+gRmgZn34tt7Mp1zbuxsNx2
nXIzNbIXH6bntXpdBoKNfHnPnqy7rkrU21nJCoXiz1Fo4wQAHd1Q/zpXiK6dKrpL
CO6UcqolXDzkJDq11fLnz2WEfU3ad7nOAvFCHGrzQ6KI9Bm2KnleRpvGIjGswddK
jCmE/LBmmKtPbslROuzwKNfEyY1iMEnJx3yq+bw6IFI1SXWCGomJgee5mvRFvurX
YQcNnatrMLigVeIXogNiSfCKAlOhS/8X350T63Gy1lNRH5f+suZJ8kr0PLApy9YX
j5EvliRcvZPD6sH14RsQLLbG/iaF8VMTfEZKemAqzoEZfViKLRnAYSiaIJOGODGi
3fvIujA9N1f1jDj9h+qQ4VNQkC29Jb4mKb1ZIlyhFw/PihtGLzCvkVSBudfZ0/Tc
gC7cIdgAVOcGkPITdLudC/Qpd9/gXbDY4R7T5nzu8MIViKgfNfIJppQhPTUc0BMU
uSSyPPa7lfAec+Jhr2BydvnKErUgk7yqEhdoc7uxdiBTim5KPfZRQjfB59li1C8F
0DVHGe+wgL1FsjaaHe0eL4Hglx/G3aXu2tmznJq7q1Y8EhmMsbwp19Nxg+ntgqwP
kRvo0lbJz5yjfiTA1qF1jVhNFbl6xxHYGKUQ8/RShl4y2iP7BhGEJRfAWJVageLs
VeUP6bWZEgmWVQCAKVzOdvHzmJMjgAoCkh9IuPKgPA2GasXq+4hdiJylfeVjaqSk
jtCPtqdrS+uP2Ps2MJK8iAczxmhfSDSx1v6TZyWB99eT3W4Ho3R/aXCe4Zt6qsYx
2IutcTeE+ZnM9zKLBKxyjAwhvvyi4EyQak7DiZVNhA2qEX1v0vOwzJAMlKilyeuI
n9FnckQEOLibOYFlF5BLHxb38yVe8nx8hWnOyemV8F69SnijVxdgz4HaB86QFno7
x8xKLJB+i3gMNW0QuLXaZI3mCKXyBQH1rLfzg4cNoJf1UQjXXZOoQw9RxJBJMJjn
ixXBBZUdPRDtFoGgSyHmYTJ/E0ft4p8MvBp3qrzCsCZ10wEyjgpmJpx0etFDDu/V
iiUT7+ECISMfdpHwLF57xCw/kBovf3jDojtC0Pr/cd4LXXfiPW1KZSCci0DHg304
bET4GWllaIm+2MImvVqyVdv58YYgMba1uGI9Q94ZB82aze6j5miDfmb4Y2xPVjo8
3c0SxcLoWbsSadm7EBo2tmgnmxWSjcEIuUL8E4mgmV8r9vYuJK2KguCPm4pXI/P3
BXxECFIhudlVmq0UNUjv8I1ad1S6GfVSDL3znYXQ4+YDfFzA6G03vsaJrl0qQAV6
+94Wh87KKx0Y4c92HmTjjMS5ctYH2dssPhzgG1peB6CsHLdUkxy2Taw090wcmzjW
dgjLdM0mX5XIQTaKBZj6vgJc4X6xppfyiFjDmYiKVuuSHbXo/DJMT3J1zMugQKrg
O7BiyIK903jnH+UQYwheZ2FOiIGtlRSMKdc3ewRD24M8xvh1SiZCvpcTZvqfImPN
3zNT5tMlasnS8xF/4OuvLYb5fa8Tg8EjeBGZX4a9MS0AXRaWTbRH8YdFYiIHETGA
tiajjFOIlmapeJn+nxfKqD8lcMt1zGp9jbmzoAWQMeKEx72BWlm/HQX4rWh33Ipk
YqvPIjF0QK8TUxvRyRjcushSFFtfHi/HLORKm63AQGvHpnRBLAEm+CPtDZXEjXEl
bimqKfoYzPd7V3Gm6lIFeY9osOGAgvfRshZOiuvOYo119N1weMM9YDxxj6Vc34BF
wHe9+Q/8z1N8QGKs2wQF3cbSxMdi1A5EWP+MUvLpsGiuH0aMc1a1s04zHpcEJdsO
Q/xyyfjlZn58L0PYwP29Gn30zskwzJOwkt7HCtU9vNHtTdTzyhs/uADEqkWDOCwa
uugu0UECP1raoWfqNmTPSIpzvzKXq6Se0ZXz1opgxrn2iqz1s5d3zv/EBCQfWaNq
ApIGZkG5LI8ercR3OLe4tXa1xgxPD6V2vDmjpsqnWEZGnCLvWVN+sZDPWtcDHair
ujIX5mudEPB9Ggg7yAt2WHVh5CkgR/jVkXRpqPdMSt5i0iKTGk6L9jeC4w404G2q
6BiCDhz9oYMXYMYqMI9CinKyN3q1XnjS8m5Piuyoz9yJTpDE5phsU6IMM+1UWwPi
ayD1Ol9vQdOOj39noFdsjK3NyjTZKxal93rEkRXfZjev7nzuK8ca0ioahbYl2+QV
dGyJbjdak9vSn6XF5BupVg/OWq7quhJ0thpFRgeSJ++iG9T3o5/V6k6uP9Lva+Ux
sZs9HS4y0H5cO4Z7WhYUWOtNz5V1VyBlp89ou/dPrA/s/D2aoEbkRuHVynnbsHT4
AbCqZ4K5LsKHM30L/UnSxSfOgO2yj+WXcIiUKhyUd80i3Tu/p+TdxYGbwL3uH6dS
Axl2oTQ6KyOJztOJQ5gCBafN/8JEiGGr+IBWk9CUF2JHuM5YcfNUoYVu2nk6/B5j
fMSZTrg3Kam1Mhs4cwSjtnARRDU/PzOCAsRkSt4al/y1VgQuhFMrUr4NlL/IY0DD
GOXBimKZklNwhs3mahiqy2gQrqwSYTo7VhWHThFmv9yd/Mct70HmjyFifhpO9IgB
KGbq+9UBEAbi/sjC2ZPAs45LlYZoVESEQdTF0T+ddlpdNTL5xZy2aT2NcCr/O431
q9DIKjKwYh+V4URTEXc/185B3e7i/jLWCZfZZBqVRDCD9pxBGO4qldDCgvHFXQix
VB8+ep/wAQUJwKCc2jx7FeQBdMJ/+I1RWjQYwSgAHIfX4G+i7+PVDZca065S93LM
euTbu5Olv5AXp81dK7rtpHDLT6GrZSvCx2tlg6IzMM7F5tCIVWXXnrl6sQQth4aB
hn2eze2C7ddaZVpacUGzAVI3biRcLVB3JV1cN+zkU+ZFX05mZ3po1LGVhx/J3qAG
WP357u+L+KXUVLfHFmX9RHFE+oM4PfTO5JnBMxVK+94XhQwMilwnAMTLYV2gBsqi
wFywnMeg2ByHO0A2uMFaoBKulYVCwQk2MVEK0sdTy9XqTJrYcqoM6iL7N8FGuyPZ
myf3lPksVytHRP+gUpdAiFjU+9Ug1Cp+IW2M2djtgc9NaUzRt00h9P9I/ZP3SixN
/Fql68ynYKiH9Xbf+Ozqr3js1LCpMu3VLQZx5NlzwyTF2+RYV7xoBHFsAgO5DH36
UQuSVm1BCNqtxxS1OhJzdhO/+32vi4HakaDkwfpnAhs+v/VTwXbcV2AHqkmDokhD
JnbuMHGsjqydctFXLtcetFSvnfgVSvXMbv8/3i9AetMp6/cMzFw9VQ0mcDQzTfa0
G2QUx7WhUdYMR0h2pcFj9ALGsXANMD/64zoerufAxHXuwFlmzIBqYNmyJeLRwM8F
/FM0HJjIlnWesUOAuI7yM//veyRRoA8nMceAf3KhQyJfpdcgaJQNYadBwhmWMZDL
SMUODUD7mZoDDPy4lUvHW5QtxpMZlDyHWM/QKnSSxHanBhJ53FDbbBaMpmJeuDGL
K9sTmEDRoMXVZ2c3gdexFwkEiBSiq3MoUN456HaAERXJuJo1Pw335xiHQVXHveUq
hz9yktBaoMBdUJn5YYH98JfQTt5OKCogK7dyY4z0h3tByhYqH9bBzfNaVdRONSsZ
Ayn8VSR0G4CjVmcgnpJF1OpEO9qhPXywMoGqa4IR5xCEgSy5L4ohBuLeso7SgfgV
ABDjXPxCMVl4sQZvbfe3l/qQftZ5pIzRhbrvpm5W08TBT1jUmOfyg4L8sC4YS1FU
DusxJdcyTyX+clj800bczaeJHOU16WczlDWerdJWAESho91amEgIC5wwfuVf0Qhg
aCgJkMDw165a4cTClAJIgpFzp7B9ucY14NjsesEuzhphFj6AW95XU8gSKy62YmB/
e6dBJX0Vp+7uyq/OU/jReru7rGrj4E4japW+kFXgUw1IZHfSRjiVOWsd86GYzGZW
EcOdZUycUNA2gXDHdoeTttsWmBr3/pg+mDDCXY7nbHf3eZzFanUTfBddPfjB5BAR
7Uw8Lz09yxRsWl0DEljJiNKD5K7SHQkNm073gLQU599ovNnbTxESlU5eDGZba0Md
iJt/rNs3TUiGen+wHox54HueZDbvi85WNfQTex0A5kUF5UQgY5ceGqeCGY+yzlcl
tG0v7YNvFnqR/NI1SsuJ4Kp3XjYH/fEtQIGUn5dEcuzr3ecbfUBPnO1q2SipYRo+
R8CXerSPhQacmT2qzhPMU07zGgxZC/HBlK7VN/fS1SgQbTyNlFvfO17hTL/M9WCd
qrPhInP2MqAkSi8v0SqUyQqpqO+noxHApTn91/GZTTgFYYhyYc+gRbd7touiFuL1
Kny+WRN2TDrYdjUf6uowHPu9J3B2zoiyRN4ScyyZO1B/EeTVNPxPsWdxVd8qxLgS
fEkP7Uy6lZn53NUCyNQqzw1s+bJx2bqCmFgl2TAcm7U3c4Tz6b51nLxc4QiQBhLK
5WR8aqh7+Jti+zivqH9IY1V/nkny1f+hnmzaUiJyUgJQABhCpoA1VhfCTg6UYQ1h
J9YstbUXVrZB5S/9PWb0Vf4r8yABc17LLake3fleztHxyw4oV6s+sAIPYPyPMXOF
+jay6LsHqBjhcsKF3aZTRDAdMp+KU5JUpEONqdO0HS4/edE7uhxz38leY6LiHZi+
5Hmeoq60LjKN820nkJWs5N2nh4iH+/AZ8mf3g4iAv0bCBNHS31MxTF6uNzERTCZZ
Qo8RzMsWv2rPilST+l9blbMWzqQRfnYgABrwNip1EGSbX+Y9f1SxUACPOVEYieaw
G+Cq/OAyp1I4IGZEwhRY0FuhRvY1+k543PvFMizjFyUZizxEs3LmJohkLrxXt/Zx
rC98MqsFHyXGROXsVUZy+96wBx0O+zkfqqX9ZtHwDuwiSmHqfLC7PtDgCF3p0rCc
P+HLURjIyG/nby+CPDm3Rc5yenfN6caCeMfpgb+AGIntTgXGCc0YHxpA/5dGD6yg
cFoHxkL6JNXsYtCZhd1g/y6/0ZVFp3yGf6ATAtF5bk3DnCi2JKnC9YjhYPGcW75L
pIZK5Qb8V8HhgbSYdiB+85zXBR9XGgb4DFbMueTjo2gGxXnVsIM0xGn8RY1CKqWA
JqkCztlCjNe7Tni2q1lz6tvrYfVpdx+jBBE/aVfXNVxz1lBmVz2ogooHpbnsyhzz
cmLvJDs/EP7HJ6VSAzXu6mXpEJsJ0ghB2RDaaIsiyQ3yyx4CHSBIFI69TB9CFhut
8VATwCT+9fYRRfqNhwY/NNbGeNhlm+F8QegQd8cgsoteiypy6bhZvkfU/G4cfgWM
re8xfZvXYeRluzhrjzLOfPtEIsYevEVzX5HLl3QIMkZDka+j0st4aV5VAjqS34c5
fv9qoJz0yyR2MrKD/umk7npGkm/ecp9ZbIhQX5bxyJMOdi8kUcuwCY9S+RK8Wdk2
h+Z/tT5b9C16iVt/pVLfNJ/rAdWdftVqnKD0pSetFWLikBdjA37eRQB3YRCK1waj
1E/8NOE0kDlGLj8lslLeRJ4i535ukSYgqYQWEoIFmtRPYn0LtpjdwduygvNoKqSZ
mHMJm7p/K7IoA8sMBhjuOECPgZjhqSvk8RZo2KCG7rlRPXKWaJTng/0WOh7mq0Go
c/GqwmLNj8qW1J9187AQK3VMBlD0kWHZwcDXBomNYn1EwfEzkp3Bh2NnQgBkeYQA
f2DtSuMPlb8MFwQHwUzRrG46OKoJgtitfte+BpdZpMeuZcApgGArdFCMcwiCAbyt
1bBsWlr2UwczsDZe+KZ5oBGskyweEQt1LbphFvVDEUQ5gU2OQCOe0LO3LxBbOyYz
5hdoqQAVYTzQL9PTzct9WczvrS8BYqTzB39F9LroJpuzsgDt4/QVOekp0F4zfJQj
6JgBdtk1bITVWTiscD3j06udIR4WGWvfDGjglRlcYv6NoYjMTNTVA9sjb3e3HEtN
XEtjbvnklhewWfjC8Z0t/WnzK5vlWRyxSBlJZQDtYdasMdWsQnFuDz5hWQHdqqqb
f5FBJWSPyyIYZo5QEItk/MW2ccTnTaSXZzbUhRfUjn8V9WRLO4dFGj2vZg50DKHP
i1oAX4dv2eccRufZsB3Bd7uTDROfM0jZElR/aeKxyYkAW4Ew51lwpaKD7jOt9bVS
ZiT7ZDxCbuvVHCH1UlUgE+cF1SFOVM2P7DvItM78tm8cTGhc4FGFQ8SbyUHDtd4J
MlZspdsUeKSnilt6WM89FuOH5h6SSVkTlGOeDxf1gLB8EHMrqizFnwXq5KTIiLWn
7AslMJxQqrn41aLthkMvxAocgd2MDCxWVNS0FjeuWBPR+3oruqPTA/n7vMTpjJBN
Ya1tDVnKeU4eRkVGVWPx8Gu7s9uHh55CCrnTDULIwWgsQaC0GwVGybXqLytrfqtt
cQpa9NFk5pP4PEtnU8tbDUng6qUCvglZB1USC3ecJ+/4ffq8lEYkWIAY9BOcSsnv
dbFi/28fwYnnxvKmM6jYPEwEeRH+ZN5Vj6+r3BOHTFMDq+ysg+qikl0SMj/L4UIl
fPLqURr2iuqCzUwZDU5qYSvoVeHHh4Jz4zO3WBJUt4zZr5fJ556l8nJI9VpqhUtB
sOU37eD+TXA5OuO227vHKp4UuVakdLQJ/nAnNzUVsTP+wGnyimGg4sqlAU3BxHOZ
5ZUfFyiEs2RkatBG3Aw1mMo9PZT2XIN/hFMGGN3VKTOFvMxoAAVTKlMcEhAgDTbf
o8MR6nsBHZrmYMisMWrp88kCkP4OOzmBcPnIy8osaBssJWHz+KGh57KSZafSt/pJ
YoR+Klb0Vmj9HZ0GbT76ckCxWM/bvETvpgfeVNj1tcI1Wb+nRfz+JmG4TajnqKsq
szcIEEs2dUPMnJr9X+sozqv5nSTTqWg5Crkt3vdYKHUGFjUWPd+kXUMV1OitZJqk
ggzAsk6wM1EvkYdCs+Zzsb5DSmNY2m7GBhU1W0zzYeX+KyetBLHsrNhKtegjOq4B
csH8QO8DCGjenbY+5n/NIXXF10IJRrgsjw9X2bk/3qNYWY3EGLA/LZsCLF/I6Mbr
i2IkmvdmEC7T9HCwhUyJQRRh6AvVji+iRpkZVuz/sgq2EALDtGgtAHn0FcYujFc3
gcZK+RKE3KmoHB2hULtyqffZyKw9OhEAdFy3QkEreLtCyoiBM7lLKW8hgOFL9uPH
s4FaUsGLX4CGyuDoH43H3Y/aJjompX57fNPfAEG+3zP+b8O9Z64OGTBce5L+wJoM
ZQYYhIB/H9xe4ioAPQr/w7hd8weVVrJmwur8JYKG4KHBxjdFYPiUyVZNaY3mwgwi
2Gegfb5nyOUZl+2LX90jOT5JTJcTvaBjFsmnKnati229KmK/lIAGdKUrarf5uor0
7tsfqpeNz72dusBuHj9Ljvhm2hFrJ8QCw2Xh2ycQZwEnJG8wu+QRES8OCnLU9YFS
5WdiHMMZQhc9KUyNklUrB0fwraMYIS0ZM13zOs8V4hBLQPVmWJU7VRTuWoDzPdXR
3QrjkpVYFKJ0k8TbnXcrYiWMyE6zrwpWNGYUKA6KP211Ew70n23hwRq+JtGHLhR0
1TL48eDcdNPSIhGO4YZeVaOAeT0fwcuZEQ1hnslFhDWBFNAoThBf3/xajNPjf3OZ
eYIJ344Pvd8EgvB7u+kljVzRgXDL8Fhjxgvqq7oMgqD8DGitJsiKtZSdhVYyTYdS
6ojn3Zp11N5xSk0uiyKhJ8cAz+TNU0cZmTJAqXXKaR3Mi45wrKrRfHwM8Jv3N8Sh
XsZzk1SRre5Q+ODmzSxH2G6QlE3F7PRfMeMELjN2K+8rUynYBouQPq5hFfV0HzXg
5oFx83FCvS0ZIu+CBukvkJT3f+P56lmFcqFKc+tMsynqepJDwAMaFYPx7ThX17SP
3r1JcIVWGJbOc9LEFQf6W6Dmtr7LZ2tDr7bODzaeTH12g2584b1MXlbNefzlSe70
1sX1jgenFGSwfflVKujiZz7bZIMZNC5TIfMJCB7IjXJw8pk1E9opeVoK9adVhoam
JiQPpRcPBysHyQlSttDWMYEyGybB3jJKwqwp7KlzyE2uDj0aoDWzhLe8cgBi0tUF
97MbMGdnNg8VhJKycdGxMgpsAvJufYm2v1hwog98IorXeF/D5UfzcTRDbfESg7cU
4iYxB1X1YfWOqt5yI2JA8JzxRb+ZZcMuQple51w+SgmGgXb4D1UynPBg+RM1dFFg
Qdg1WWXI6nPGyevTyi/ehNkPtsswsD6XoIBO1NT5bx1MA7BRfL5HsUiobuYBR8bp
IfF9tEGPXEaHrYCgc7Sm1H8IbOnoPkBHjylctv24/7+2Sh6kHhc4G+LVJAbeRHPL
ENY9Yv+hLyTTOXm3orUVLGQ47UYaodQUF5TLON8mFpKjWECqVk4tz2bZfddM+ITd
x3xkhOmQhXi/gclEIUnJfhbGkCa8P1K3AcvbndzHA7t/nhO94TkMDYoZWYNmlrtE
0nuh2kkHspnvAcV8rDrT0M75A4pLGvhG1PPeMnLmri/fxVx24MdNtd17qe299Y8S
Tv8XQuhW+Zw/Jui+SeQB1MEf9HsvKWaOrMyRGNqXFpjH7aTbuF2W8y4JkAt1xWPK
t2YPmB+FFeQI83G0nb+w3lnibNZoRwjwAJcQKfndSNrqkXfmtlOAG+n/DRahfssW
xFWe6cfMPaDxfBgZZbJWLft4yH5t+UZaaRwW+/zbznzvP72ZomMYrOnV6FNnvI4m
`protect END_PROTECTED
