`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/MFMvZsJ09cI3AxUod3Pguxy8BkqS8GYL1wg07o+1m443lpjtcm1zR47VlZgyziE
sMJNLQrRRKw/7/oc1Hy4xUi12dC8gVGeWRqWHzTwTzZNDnf0EiKj4Z17x9kRShxQ
9MwyevmlvBUoEZONmdyIe5WckYBcmBtYvrdLnCCO5LnCpMpfEghKP/cJkT1F/1J5
RlkSXX7IDIRSqy5JXgQXNN5PEAmd9fabtW6+vAtR6IJs+I+d7gcipa2vBgtDOsr3
VevKy27OArLBjRw3uwyxQPyXRQ+enU2FaNmQufXlgoC+K6VU1IOfUlze0hjJOJVe
XZj6i8FsaPSAd6MVxsrL6J60ABQTFete2ERqnhoJl1AnoWCeJ+RPACDcrEuNE27W
buEkenoj8MvGEMH4aG4YZ1YWALAeYKNDOUHJ8633LMxTwiNAaEP4Fry5zeUNk+Ln
x2SR4OBQMkFPhkaSLAY+SHVASC11CFeYHBYGAJOn2HR85IRl9nnBQW+sm0paFL3h
/cm2aP3zxLiIdugwDpb8XEsB8yE3vMeGA2kkBixyqtxnhSp/1BuPG9A9nStLKhT7
bme4FG5NVbYlMp+JdRfanXJJIxHb42jtCGR8+/GX0tc5KU7Oce9cAQSSTDhr1qEK
Zw0pMnfUOQU04zhzvXdhl9hK2ztLJK/93xOoXe8uarCVEpLR43P2YgWmaB+Hfern
eCMEGd5sEHTDEg5QQdVTa/ch/LhCArEfyVpPpEc/mUJIl5obQ8BXEEulH/NN4FjO
a3Mtr1RDEmK37LxrB6MgMkiIsaeTQo+xDSkZWq12Va4eo/RZOEm1c9VgXSGETeUj
QaK5TOdWJt4bl4HNnlHGm8defKtpKWLUmUXlvDsegT+DpLpiSfs1e8sD8Z3E8O4T
+j6NOj6Vcz46p/BGGmrh1UZfqAecS3gFUqDFaowe0JuWINzm4PRbCOo3B0STsead
hgMA9Kr/BmjzqqHU/M5Yj74jBnLKWU9bTSNIO4NsKl5HfDW+BHWYYnGLwf4WRwfq
Q8gRf2isaYN6cV0vbfyyRZmdLXpi4Wi5nhIqUwJCXfX1ero34OdwVMGrsN0GIyMr
QQTlpdO3tLrh4Zakm5RRVC6htkDzUCXPknpIAA7OjS0OO5/1jQHWx8pDTaHQMsVv
jgyp6bWfW1Xyb4OZwIopD4qDj5pr/qS/wPZ8TtYcP1PHMqo1MgJIfAZjmLkq9utT
taZUdSfAgpk3mNiTicldqeEQ8mNrQ9wyQm2ibIJqfHvy0jJ/3iKP2z12n9HWm53i
HnOsXHTVrE6oIF8w2jjchHdrKirqMx/GkTKJkbLHzzCi5ydzQ6wi8cwPAd13NkVN
n7grC/ljjB5hz8s4nVdtzTraSPjkPPAQAOyJb3b8Z9RAi8oXkvBbXioQfrlpqKQ5
+u1HODCd8wn6EpeXCtf99BUxL0Kfc0T+4RIEfzFfHwiBYyo3EOb0EFidl9kdmT5z
WlGW6Is64KOmG/f8VFkM+j8gwSCnSG136sfxazetsJGwlTEoaCS1wJzWFP2pEImf
ymxmY6kK9MhxU0wfY/oHMkBkAG6y83AK442G+CJwNvSJhZ92iozlJ86DyuT09sDn
Nb6gvkkklmOVTyry7MXrUQaEhPXlG0cRUiG2UWpazJJq7JCl76uiB9zQ6pFdUa2t
WjwqrXcqVfs5O6AfiGgAcc28SnOpVDN37nd5Q4nX3RubhxAEsqmF43XkLntnlti+
U86Zheo8WROqg1kqOYN4qaEvR6ruooJ0DtW+fpIIAV7gj5ne6721hqomZ9X0FPhQ
qbZix//4X5/YCnxEfaDtCFJY58aHGYEVp0Fr7Pvm64UeSWC3Zisf2ODjh6XbWpkA
N3gjptZq/QaUspFZMmLO7Idy7jf/1+sxj5W8Vzf/T5g6APkua8GXM3G+tiy5O92w
JBzBQVzIhsiYEZXhVSeE5rR3tmuRhEkVnWgiKXvGyVFUjK5gFqXpYX729w53NkTJ
`protect END_PROTECTED
