`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuk7aoo4l0u2o8NgSD/cvSsj9+Hpaxy8Vf3+McwH1vRiJ0/G9BmOi5LyPNx6t1RP
7WJ6mmkHMl021bQQmTD+KzaejsubsXERYQVUEerNKXNi7miGawFHQjhJ5JrIuXjF
B1A2NP+2YPwOcme/XEEp6nMoPM597ywDod0np580FCQCoz2qP16R+Rk2xiBIyDJY
UE6HBOipBbMYnXhmhUi0CSV5G+qu+LMDVl26tQJyjfmHqiRyLoKv92xgAwrQs4UE
OwKXNMZw0a49bLxsA3T3vxfUE91WbRRyXPvffD7dOarVQ1wCL+rgKAK5LjVDxI1G
3LpccXx3TOia5C+4uZtH1Z3EVrKSgxYMzrABEIW7qEZU5PfGc/31IUh9McfPHfNB
YNFeqlY6ZpxeH0jotgqkPfsmEFXNSLecekLvN0J2vH5JF5TmWC2xZEkaqP/jAEgX
T3Em0+/fawcpHwGGITeRbNY+GXkeY4IwRIzS1ANEEpfQBzimT40/1IWToBRHZpGg
LwhaVjZVk1VYzy6cKcejPTYR3SB6+UHVMJDF5YUjM9f0VV2LqR+ZRFpnynBftrqy
vXCjRIxybiUiPjBL9mHsVHmtW4VZTnHuAO5kCHM/Ug8Z/Zhc1ThUIgWxaJfub8Pj
96e6oJvppA6/o7dnbDeoso1/mT+yQdDpIIkheDrkmEaNl9VkCQDfc+D1qyedBBEd
83u+jFjplfKmfseOseuADyvyhoLMYISIb/BiaNfalWjd3i3FhIxisKbIgf0QpzeH
mQtFY08D4rhuH77NcF1MmjOrIWzQsNLn0LUueJ2EZ3uM7ai2so6+4Zj/ZCzX+11F
FLivJ39n7a/2Oef6DFilbP4KnwMkIaEWuWrSPot2QrFGxrR6TA0RuYH4B22uI/9s
jz8p02uAX+PXtACFz4rm0R9yUWJ8+yr9Om9jY63QfV7/XfeuxMnpFoto1XNxaSvm
zT4yDZVaxwJuF1h8t+4z1WTPlq8+/KiXF7cbd5qYOaufzZWMpLxOHd/1xMtx5DrZ
1By/Gr4Vh299M4yXc6wZeq6cWXNTQUoeIMjuRi3BfmAQPcsEO9WkNJZ0vHDguXBa
4zUwmcxoCeKeMrZOXiy1AyOnI4FszmohF57vye3ruWKvSLMTeO4S6XkMkTDQ8DnF
vaKOby0a6RHB7IFo6tPZ8bb4Kr8xQOm97dyOzVgu0IUJ3FljfPK4OnrFUEN2/WXm
p9bEQtVEq45ZdLj8O48wS05lZKgUeO9BVVFyV8DvAhvQ+IJyVc9a7mQLVobEkxUO
jtCnVL3pudUB+CUJ0P6CTVCyYNWjo7CahceqxjJWAZhK4hg3L7xbgqyJKJtFQTc0
n8kSuIC29zyCEu2Ykmuh+hsidCA3+l78TNHh75ExUZTlx2+mCJ6fG2dPT1qMm5HN
ae+UceqR/tidDr6YOa9uPiWOqUr3dI6Wi9WWG88FXUZjZ2BBda+z1p7+Tf7Q4sjM
yfBy4bOMhnbiy36WtZTabNYeu1bNp888Ygy0Tk36yzY68jlJpoaOTkxHT6pdsNlN
1oXekyfrYa0FW76FNXFK3YKl7LLf6KIx89Z3B5uUmHhd70SwsD3A9QLDj6dy5aT/
JI7J6xPYepb/9EXFhbyV5wSWsMR+muGvuOY3eodF3/TtF3ra5+tjsV9AEW+u5G/1
`protect END_PROTECTED
