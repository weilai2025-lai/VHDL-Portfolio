`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YcnvyMQUJjnM4l8xJ5kZC3Jmwx58IMgnCzx8FO+u+c7SAzSzLeFWUTYgHTxGbc/L
zvY+RzuwpMi8brC91ovueOFvrYCP1UOU3DaeccYyAZYTCZVv+Hkg42uGuieCXU0N
D1Awdgx5Nl7kNLTkgIhb4IzFjskvMSkfSZTgosp/b3WgFVvd2TWunPQ6+NiFibGm
dcmnSGQTHqQapxj52MCE6W0XV6f5I3XocLqzHhQDj4x2UQosEFT6hPMZGYCkbmeg
l7+YUbhbrRNTyEj9s/1ecrtyVfMFZA+55QAt7845SmLp9dXQtx7k2d9QwrsgPJyM
sSl7WzQDwPni+QFzaIMlrW7IWC9nlun7AER5VMl/JeSmsHO4hYqx0atmxz86tqKD
kzMlwFXjuhaNYmi6X0oAKMI0CBru7ikbUtNVFmKVuG5szkUkSA3Jey5I6loV8Raj
JltmXhbDSiAWani25obRpA==
`protect END_PROTECTED
