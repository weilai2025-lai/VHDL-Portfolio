`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/We+6j1zE/YZOaWU4MgLrCz4WSyl6q7YwftjoDIwpyNjmfQ2qEGPKwY5vZrZxcQ
dfonHwAWefcviRFdQXpmbUbcVOJoVMZCgXhnB4lz7BnBkCoE4DzqHxtOQ2gc+h3T
Z6SUDjSzH6lE/Olc6LBlw7gniobaljJtZO1p8W8En/oQilhQwnfO01NwB3QVbccv
giRRuMU3UOTjCsZKb/WLqYe3yqR6AJsampwI9q11dO9DaQMDxuf2PB3OOihffsNx
LNUu2FE68T+boQXBqN7nYya0/jWct74ZV1DQ1OogJ606qEtukrxafmYOHOnpWPLB
bOmFn+BOJ2YyqnvbvS6r5GjS9znyEm7vFJizeaFsB6w46tl4V75FXreBLifBQCC/
qm4+7zmicwBhNbLZ+x6bCVxWFHWPvsFgzjaxVQaZufJdfsvzwnxMQjCu8jYGdBX6
isz2VPxlIgXtA45NSGJ+i5r3cYZrqlsG20D0ZnU16G6WzvkXMhofV4j9GyyIpzCi
3YyankAKBFVLw9/HUy7s6n77JIYWlmQVStt6sGiin+tzyjswXjHTprUOT4kQ4a6e
Ug+dkpDWdBTCZvEUIS8wkLKOLqWrbeySnQjOyEwOYBvx111HaYZCBojCkrvK+w2f
+NQJLIBN9akTtyOJ77JgDy4twIP3gboPh4CMJYah4QFy2mse+HZeWuwYi1OI962q
ZdNyRM8RLi4NMPnDAHFY5GUt+B0xE6AVM7cPIlGiftqIJxZntdOgrJ55/96qCT2R
QWdzSuYesSpxEz2e7VkKix6s1+8Xov4TKa3jcDvP0vR9s1mHFENWyYd5oKgqZ4CO
QLy4ForknZTjp7DyJF2QCGPJo8HUPp1+0/oLq3SlSgmR8QksiZCCvuSzltI5h3Bj
9mcJbUi/rb2JL5dZdIW2RXuARG4XqBIOBVIpjAI8tR7EIFOAExMPnkr8n97TL1Iw
n2Z+aBuFZav/OskaUDSOd66TpQBv5CD+5e4M4dFAnEG/PeC/FSnbObr06gNyfVew
L2Wzd1sRUigS2s3MAZ//QeKGgm7gqyCyWu/cOCH442uxl9r0/O776TNRQ/0KpuSl
MUq3MMKSbOzJ3olzBfViLRWCYcB6Fx7pdVEgC90CAtgERm2AqiLHFVsgoe0zO8Xs
WwTOnCzg51S6YhDNupPKiOhcrAGnqIfCiciNeEBtWRiRO9NR7b0/U7AVimX/ER5o
zxwB5pCQMiX/7D0eXPhINxGYZZvh+I28lncF8GyFxtFo0M5dYyNoqbuTGHe1rs5K
j/PZnMJIpvgyjxQ44JhiGpCGdRVnQFdqYaE070amXkSpVeMBPwMHQ+ib6DSZS0p3
2jAT+lzt62fKzrStez4t1lZx+AIRVfaBUhaDy6x+KA4djsOEcS6glwTteMKIjvmU
U1rqPzYPAyTKV6lcRnWfLQgVtTMg2mFFy72xjdtAAqLA78rdDYMcYw/M+f8je0C3
`protect END_PROTECTED
