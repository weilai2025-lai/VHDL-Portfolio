`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L8uneFswNtm5uKS35Zv9v0j1mSm7F2/y4ESzy+xB8g/Qi8zKQNlb5AMlGyDMGPeC
KW9TrKPAodn3djeyFNQzq9R4TJY+YoQmIG1yj2pxysqLxRIp7L8CslBEE7F1MW24
IAszLRwZW/tS8dQ8/LelBVbzuhuCXTkaTIrHzbG6dB/UbNoFbUJC4fMHjiY2nuw2
Sa7i14dEOb8gNqSHdIxK39M1zS+FUl68Rsuw9VENMXBKdiptR9Ppfw9HYfnq0Xcn
8DDIWgh66qA4HlWzVyu4aY30qRlOl41CoDqQj5vza17cp2G4WWlOfY4DeXGOQ3yx
otmCQq3/8nvd1BTIiFTy+ksOJpEbt28vgctz+RxhWiE5/BCF/zY9gP3yK2L6vhPs
Z7op9Qaigq8i3mCNedNejxlpeXw2X2QIB6xjEYVNIhVCySEWxn5XDfhNHNPKGxUM
SULOwkSDlXTiZvXvunywTJp1GHSSA5lWoPhJDCUnrglM+8X9e4GVvd8CQT04haQL
++Q+ejsBCtfFXQRuc0a6Ii6QsDvqg8EyeDp44CbLOC+nWpFTTC6FIqawkr77jQeU
VvWqyMi7nyQF3Qt7Ou59Llf+XgVn9u0JIIvzQQopwAWcT0HtSDkJB3fMMXpIn9MT
MQgH9ocBMSMqqKeP3epVhK2OIPk8e3WEheOruxqKASzoPiMsBg7kI8Y1TgSWPh+T
G82/17csANHEexi5crcXG1zIsv+lNhjRcuZctlrdqeaI1tBSRugCcAXeXqRUgXgK
zwt8Ih+h0ppvcRXbqgY+sSiyZn7Jav4krWkll98avFVE2OpqjNd4sJgPM0cIx0JR
3NbfALYnuUP/x+2RHvBjF7/+vT+rSBBqsZxP0i9Yi3gnsX7aNgwu1J8yQRtwD7KG
yHBpV8LuNo0yJ1DsfMTVlJWNdUsaRGCzqJQB8S+6Ha9Sx/W4LAdRkVyonZYEzji0
TYO0Dbqb3MxELwZYXUHJUJyfD8ekzVSUtN02l/PqaTjqPJq545UHznuCYiUQB9KA
s0luZrNZHEtkhtiAOZD07eui0DKHcbMER6Wo47+mmE4NMr61uAWiH5GIEQDFdpI0
SIMgMte/YiTrLXSd4BgC3EkIY51RQyeObIy5vl0xC8MNum5+hHFpKwtIHIWgsElM
N+e0y4WgfYadBh69+kuYioAbbII/1Ou8x9wcRNkQz8KOtKxhQEU1+0mDQOum0NlJ
ZQS3Y1kx+Rd6Br+G6yb1IIGxe/giVkXE9SzJC5mgfhtAj+4uDWFmX8EnUj0CRB1h
ifV+jbDREf+Lw1eRk646eYYa3IjnAnhc9RYf9grQo8E6Uam5qno4KmrV/jrK/AOt
W1whfb7dl1CAXPBff5Fms9MtcQNwtUo6DBqC4pLvBseC6X2dTf1iLCpOFO1krXYI
M33Dvx8W2OqPL+9V4VhbtHWzS44YaeVHljjdv5GtnDLGGecHXos7ObDY2fCTW/Hf
LmUwOogZGx0ePZKFKt11jq5slbX9GEVhZy3KRpiCymrU7jDfZUVTSOEK99kVwsj0
vfUHKzUyJ3HXnIPBASeK29pyQznVoU0+wvCTDnesPuFgYesAcLtQA8ijyxfdCNEZ
/+zMMR4jA/Evn9lmhp8fkD9dOyUGP0RwB7fgn4ZFpi+fEhclo9i6wWr0CXxBbTpg
PCX8dNFaqBG2MdfnJqIw7AnObpNJKb/AUV3W2t/aQOLXZsJKphBSCOMWKOqG1c5O
tPaYKAfEFmBb4nej7SfWiMPkyz4P6DDvT9xbkZwYwqovy6J7K34eB+Je2UrmTXk8
hDbgBby+JFjh6vNGqXkhEqgRLIEWDywBdfjOBLI2FRuucNGCfX1bRVN/n8zpHL4d
LbgjMgIoDT4SXNK3k+ajIcTOhIMDaMZ+LnDxFq2ayK/fXJy2QzRQcjJH9hy7G24O
lWkpa0rNKQWOOopp99su81uwNoT07dZicN7jXwg/GPKdrxXVV6LCO0CDhzww4XiE
aiYb9jRAn/goTgr3MG8t+cUmMuOSzlBGLBQLnNwE9uZUy5P9WY59FR8PyCxBEGWz
IY66rIXesr6vMubkTCUOAavrW4H5caPle/kun4bGu9j1DaPWhEdykeiKrxrS0KpI
5ipoRjU3VldpUNpvJncDk9SdhB+RiawpeOqYdUrjf4aDZYCrZavD8+pl675jZwbr
rs2tk7eswFq0AzkKHSAxYEO8sqlrsz/jYWSM9NJI2BSsoJVN7XMNxTn4NJjbwYoy
PN35jZdSn22Uup9vfKLK2QBmoZO3jQzaKAbi26iIvevpCQzrOQciWCr2yY79mKbd
0OxNNMEkt6IiGNguM9DwSFpmrPcMIOeRdiNy+HHopgBZy8DuYj0rkcqAkC2naTHj
WdIv7PPkp4Wxk4DOWEQd5HiRjl8BdyPkj4kBpO0+1KPqiwJiIskEtsASxne08Co4
tXiR6Q9ZkpbVh0mDKomYLesqD/F02L3US4Xd0Mp+TRFNpvHF639gagSLdWlOBXTE
+gNKphubbRgH2oOk5G29k/xLi4GWsMO1N2UrNrYBgWow439sX5LQ2oPq0boU4sie
gwwMtdUaPNc/aLZWurjf9+mNIImT8O6VT3192e275zOU0MQ8ZNat4lFTgKQr/sJC
y+YtdSYsmLKwwf+//jiXnEfRi0G+OWS37mAc5VSc4ua+qS1mszYMIACQH8m1KqED
pXxRi4vr2Jpjq1E1k7KV8DHbwsx/AVjP57RHPq/ZcL5MqqzuJWrpbATES2pkmoO0
qKPqdRk4uG9doYnr0U/MUpvvax1sPa5jhmKKD23WOKkhuC5rqXLcHXHoqoSLX9T8
bKkP+3b43SeRPot/59p7uxtB+OyPg6LknsFDAaZEH+z07a20QBTcjKhnxSlRcpFQ
eRuZ8/PeRjHPQX0ehir+EmxNe2ZKfpU0szca5P/gcihQpjeTiT+vmnBuZe3JKD7M
SSgjFnKDlqYoGxQI9dKO32uIwFfvhnGNPc9dkBC+Sivel2aUnnNdDhJcqs2XDh1g
PaaB3ccuC/3qctc+sx44A/Cjqtcp9huudhAvOU4BkJWDs49qXLpWmCjIOeY/fz0/
GYOriE+fKM55UzHYvXbv0C937skF17BNFyxKLhcpi3+noGoG/RiZzg585O3+OTBL
3TtevMMsJOL5MTzu/TuAUhG1TSa2QJVPjhqjcsE/4DxuHNRBJSzfik86DTai0u6d
Nwh6QA41rWGdUi3M5P4YT2z3GIaZCYVBPrOFMnZXLAxGGs3Cg4ktX7ucxz2Xz1cK
LVtbJOqPHNMJQS4qn/RSt7fEDcayoDDltPvvuMKoREN+7Y+RKo2T8AjyXATYUdUc
GxgcFGSu9LFH22CyE0RzdtMJwKYs4l/AheA5bdkdqkecejCE0j1rf4v4XKKJRxWj
0Cl26Z6iGKbBub57kHAksD93Pf+NmJtfX4HfbdYfa6atHN4Kx5tU83mrGZhquDD/
msCfi8R88bFvOckz6svcs88efU8oIXEi7uBeYKM+9i2ksZbR79yPYbYLKrQ8qyCb
AaYVwAojrbUK1J3iLEIxwcx2pTqQrxV18EFPkHaSHjJr1TYTpdvVmDey8stvS+3i
b/CyvUfN/8Yf7hdEJdgiS4aeHthzKsR+0YMLTCf4rC9V0ooQpK7uUdAjQqNboKbe
/LSclDPyAIVHVRiEmnfZoLAg56OqOpXXPv2AU/TfzvOajcqXsRP6UxzFtKykjsgJ
zG4s5HX8LuDCv0m1pLxDFnn2UXU64obC3Op5D4arp6lmEfpjjK6jdH/RZxnmtSdG
Ayvba/aEId1Lx/NmjiMN1kI3QVWu6faEwkppoT7Qhy/1peIPCVzJQd/NTflGJ+97
nFuZtS5fiE8GIqyHEZPP8Wsloq2fqnmI911R5mZ5vlQGFyxlaKioNXF9JYPWtEOM
ODeRoRlF+MOub/2cTSjy10cI4vdgXYeePNv+Aw7FG0b2e6PBrczgGg1VtzzxVEzP
kkq3+OKqqKNMB8KlMiuZJFRMOkIhPTVxAM0bTQDn4G8RXi8r85mHg9/hwvL0cf8G
MSQE6X2FCgMZlP4nPJ0oyyJOMI6wBB/tPJVNkj784GJApg9xex/E4/zcYOngGnih
gOba2YUaNwruY88Yqjdr85lDjxxIOg2V6LNshfCnuSuVXSt3qn4bFNi/uWk0tYHw
/XIqLRfQX1EyIISrgOgUr0WVPitH6krl7XAk+WkEKCoBeTYwrn4AKyNyTsqwJy0B
91o/9S79K4oXuK6UpCUws9g94KGxpCrzQRxK39QUGDEJ4Et2SVk2V94gqB0VzasG
b4ZvNf4rO6phFUTzLXKLBfTLAPR2tkRsxQrAKXj180s9+X5DUx8KoNYKnVQKVWXS
DEGY0GKGk4+fhtpXgrjiXjBrJM/8/xmQuaqM0j5n1fLjFTaxYbVC5mF+Xln2sjsc
cv04lgVE1usfG9fQXVbaVWcR3XdSzbE/XoQVG1oyuDWbLQx4dhskfO1lDdYyyVYZ
WcZR/aBsC8BVnu4nlEJETvfVKUZh3lkYK6fRIKyzE/boD6+9BXF42L6oqROYOsgk
uM3SME/Vh9m+KLnxFrCdl37snBjkrG+mUn8KJMhNj/htB7JqFhfG9WuEaeBoXukr
vpT9sPOvAoGE73mCI4fHx4ks3k07VdCxwlq+0YWuwhTvqBnAYjlalJGXIOozc+Eb
H816BAgNAPHdOnGSg6vuqoYRcI0Aa+kscrFARPqaEdDCD2J1+/jLWotyXtlXiLL7
4XTKrHRRQAieokrFc4SjugAByn/JAdQOQ7VO9lfzqBcjLhWa3I/gEuFH+HOx2lC+
/1WygCvAmlouovSFDArblRAwG3wGugTjseSlyUbacKlTdjEtRKvvKLFduMLSMlWC
VtQWEgTKLe8w+P0evUjtmOHjC+adZKDUPHMQkzmZzLz3T+H1ZWj/hP16CF8yNEce
6139KZs6f5YxBFBhHVNFEcg675rCk5auo2KjAu5XkYUDJxHzpu4PC6cNanN6ri9L
VHDLUsuA1gskNc5g/kMBfJym8/05PbdZVP88UXLBZ3aPngI1vT7OlaJbIi+nnCG5
4AZVFXFNFE1ekM4A+FG7F6FYCQc2Jp/+hAJqwKANOfH8nSGB+ufEFA1W0/H2iNFq
T04UYmAMhOa0yvMhnkzZBE15gBH4koJCT8XcwPWEeA43IFknVQVnmOZOtV8+At30
w06+O59nPLEJEq62Q4fzjFVPk5yfwQA9RwqXiwcG+ZH9CfvmG7AGyAy+nz2STlwp
zWHOkz0iJ6BimwsRqvpmbNJOwfwggf+XhID2loEq23V0lIpLgUqVN3hhpUwBg2mD
2rLEvcmDgucLajx+qnp+hN3FVeD/wy7JR5lteMl+bgXKHk2xANc6lgiq9yqtyTl6
5TsdvPvSzrXDdhR9XwLZuZC2+kZP/+3tnc6Qh87/Er0/cYPOsnUZHVLC1sLB0cP/
/9Qfef1R98v0e1T6uqoHuqd6FISyoB/dYCjFzPi/wF9BZMHYQQGUVMw7EwQ5+3GY
Hp4PqqbyDYpKhTdX3U/gmenPEOUt39qiIkQKdz1fhnIQ7V3siyMo2MSrMvi+5Rku
4Gghmg1/ZM4qjM4KpK6j6A4oYRU3xFFy/vQxNZyN7n2NcfnqDQX9T55Wm03NjPML
efWrdfHjz6ug0hxPivFFBUH9wUMDaeV5IoKqylNAtbbsAmKJw75HTO7aLUTTPwNt
0VAIhUDziHF4zSBzY3p/hN/ARVX5BR98H/tqxBE4xfAusgYuS7nzevoDw0y+EiIF
7hZ5UPdgckswxoOpwcNVgTLLgInbBIbXLnhpvq/Fb2oiNjnEIF1weV1Z1CndGdYl
hFf/S1QLtB3gV7/RTdfub39LXpf4QJWbh55hGBe+d53srQmgraTSmsuyBIg13Cw8
wX0K3LdL91mWfLO2fP6RvOgSeCemUvwRB+UTzm9cEAKRf52T8nexk8joZwQpug4+
7PrXh1F3+i5nwx58Ggaw1779C+x2waNwcywTx2DLeUA/qAOCDmPlYRRCcdSnSmgX
0PzWGFD6lVmN9P6TVr5MghvucHK+R6lztYVOw1Dmqx4SVD41gsHLkiMUBV+gwanb
9KFCea1VmtCcHAAdhTYYK+Xz/8kjAnDjmiOTqd8cesedVx6GsFz+vFjA0JYalQ6W
N9FA1wA4insrDdDOln0kYUwF4c+oOd21/FCLLbzBxi3ZbIGyOmmOiN08srnhxAhe
coH1R/KBx3O09U7BEddYmFGdDSdN0YpGbabLHNXZfZqA6R8V7MKeVy5A0BOLRtqe
dMPktGYQyLsCvc5zPyOPKgjSp4gc2iVIMBzoemewMRWmUiCyez9lld4zNALUUonJ
wFp27WLHl+9UQww4VA124I1fwd3qYhhVQTdAnUiAgsntW2ZUmODS/Oj/HxmyL10z
dxo/TDHPDjtOuKfSOqAqCd81mrl33v1HtqJccycBxDSV+EhxONUwvIcvduRx4ov/
eQjmqOZvABRjI/SrBihPiZR1fzrRaGMaAzq8mqwTgKlJGm22I8lwwkF0Sr757hXS
PUPB9rvSCMmSijaonfVLrzmEU1Kh1KiNu9tRWsWqUpzN+uJFof+qhoOt9pOb3QL+
j5FXIiokAAMhwRUgkc1GBH0HmOhpgumTgWn9hgG0OWKEc8DYQJ5CR3lktPczwnhy
OQPGnS7EIYmq2Z028ofRb3lVyBtaP1l8/5Vg8eDcyCpjgwcLEXx7ofRJ15UL2yGw
6NydFl9bPOGr/Rb74J21h/HTNyRl565kRugBpppwBz5O/d46Knvw0ebYak4anDT0
b5eopOCIc4zXDd556cgoYXZ31WMW8K3pBDnfmk45shuMP5gJCrGlav6GXs50pwNl
81YpKg1pe8Z6FSI99SrYslSnmBlAg/ziDwybIma4O68+o+RYe1bEK2+dgJ76M3Va
2FGFNqSxpaPbb4fprKUYq9r5iJWz23DtLSSrV8tfK3X/qQC708D6G2Gp8ZMK6915
DXoKz39bNUnTJZGAUZEcTVmYXu+lR6CUZ7KTA2snU4R3hBkAazJB6JdQfgumr9xW
HpoVGufgGNCrgY4lXWkLpyZNaYSXh5tmDRWhZGpo64rmb2q5r19SV+Rqn5lK87JH
yquctFF4XbSmzMfxpspRtSUEfnyvPK0/SRVVKUXAj3+bFC6Afo81LoLWgrVxdW+N
oQWWvVUMkoqxX4/t0nDb2HmhpPPm8Cly/UFM1zkgB5t/HieWBM7h811dWNW8gnuA
t5fEkdbivo5zyQVc49/6SHT1BWsjUPX9UpBuRjOEo4w=
`protect END_PROTECTED
