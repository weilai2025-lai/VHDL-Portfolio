`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRQLen38tDke0hiYee3UNyvvgBmPPYuWgiPeC+0wcE8UXObFYHsCrGXnj6+/lOvl
rGV0iv1j4l4npW42P7sE1wUArcvnC2pQIiKQJFR2gfh2fygohiHSWXxnBa8+vDPJ
GwP5LuM6lbZY2bZFcNXA7kvlXY4jY/cQIoaMAWEVzlRl2E9f0hAoS4/XBKQyuOMM
OrrS079hTKbwR86GGVw/mmIye5rWITA6mNcZ+ZRglA/ZdIoMgT1Iq51b0vsIINNO
4xFve2zPRaW23dm612U/5ZtQpjasaj17z+y+tlWdSfns1xYMg/+C10bF0NVcN6gH
vYOdKS6XGpa0w6qyg8hmWMBFphu0BKxvdcdDEi1pNFkffByzARxKccdHzFdVP/FC
poBY8Ti6yyDtukjPuwLdRdU7PsiLgCNXjBQEH2chIZQCixlxdnHIE4sH1KMFwtuD
hBGZi/DNuCGj2Ds7WeOUhlVTEhRoPSzNimpFSnjStT20nIrcEERaNq3Oq4re+9bA
9a0qigAYUZdMvxyVs/ELmI7kDXVfiyAhQeAq9Lw82Y/NTQYqhl4anVijBz6a1nRF
VzLMeRvxcIrQLy3u1zJzmVn71xLmZna86EH2XFLxeBGRaV2mOOI5WltGnpgNGKgM
HqIu2jGZdwv6qkQ57R4C389Zjfisx2CgGgdNL0ZinipHPIaOz9wZhKSQOr9H5hSf
RKxsoGwaItuCVMqrmol4f7n1xkvv2xk+J9uHOob/C/jGaO3ihqSSHApOcmXDs+6l
f10TFIRJp9sARHS7QzAiS36ZDSOgKOUi4p6BGWrrgl8b5FQ1SNX73FNJ2DH1Hs8K
Ggq+p7K51A7naXNPuwQUFlqrReQ7AYnDzJmWBMQuE77pnvom9+rSfXi05IRI8LUK
yuCS4/A/GS8BQ2gam8x0KOvXqGMXGNUn2wDzKnXcsuQqugoK/4vn3T2Pg6t9+2ke
Mk2ZeVyTsfoXMHaVPcsWLOfYVU/pWurMcuVfYhJkMTQHrwVOxmt1BKqJexENnd1d
nMiIBaP5ZnQrPp0CKeceDAkV5A1AAKI9+lM6Yoio1PyeKNuCMV8M536w61if4KBF
Un74hFdXMApxDD6cXHlocBTp8sKst7C92RrlnmL/YvYX2EG+ujnqNOT75Ma58qB/
aEoQc95I1eIUsUNJcFdfi/n187RXR5IyXcRBpKHyLI/4tXdKqfmdGqiJgrJnbBdg
5ZBrtYwaVn7UbqLQJU7tk5Oma+SMWJ6fvQvcXIeEDrWmHs7Cq1YO/6re17RUw2FS
qDvGqYLpj17vHYpFBEuv1q21goipYvc8Stg4BqZWxb36IEiFQwxsWzb9QJ9ppNA5
gue1PvZ0BULwxL8R6oHwjL6sYGwC1u7sQnPX0tq3DcsMBGt3Ys12ENTXN1u2CPjw
CIBptL9zCUMyFQwAAMDNwY9yVo7Q+inSfGoZauWGcDL+IQhsLqJ9j/IJ3WBf1OLh
84coIe4fper87JdKFbiq2PGEmfbG64lTnmgsOxxIUvPZVW7wbi2s3pjzIRZK10lN
vveTsVHdQNpH4614gNljJe3+e0259MTm8sQydiVk7RI8n8UdmN4+NFJhkFP5zhbL
x9uDaN9tRJ5sqS/3j21lzHD4vyOgxMNfEcQzmQFhCjo4LcGBTbtoScwZ469RgXu5
vYiZu/r751AfyhVM9667Q0Ewy5IbNhDxUh+iQl1TFFNYsxriSqTNxpU3vv+9kqBP
+s7FE9HqOA4i7Z9G2VdFvY4f88kZTIHLmL+o5W8Lt7J9TPzCd3dByp3Fif3NxOwA
JVRov7Bm3qAqHOcv3Bn+ToEiMHxu4uhYdx1NCavgm8BSkUQpnjc6OLOcyn93kVdq
J/tCkqR1oPbEsaSP5GhdvIxGML5lswkR28Dx2juaORjsaAVfHN4Q+K5oSzPN0FPK
2QUCT27dDcF1uvbxqQn4uONLM7iKcYZEB2r/DsD0iNOo3RgZjDdVqrQt/SxjzZRW
YPKx6HwaZfkFraWsHqaTqiRVuB2wwIDnmYJV84rpZw+IzxmLQWEPibHIL/PLsTi+
j/88RSILiD6L3cRTU7FdwaAMx0QOFfn5ROoR3i79RGUKaTck8+fdnl0FHaknNCOg
RzQ4+tywoIiaaCC7v5eZZzZzPfhTsUGBIV/u5Pakdg9o1DYliSzVH35YvnQH+kVt
puK34XqthCAe7D6RS8Ospsa+STP4oVdpTK+9u14B9GdF3iXLAc3BCrx37qecKTh+
caYdzRg1Ime9V/WbXi3x9g==
`protect END_PROTECTED
