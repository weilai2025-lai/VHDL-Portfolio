`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M20VIoaYWVMTbERgnMAvmI+48rrQp7JWR4S1qnd22XBZC8P7/ouCYf/ncuS7wYcJ
TMhS/PeVPQeFumEuk2U8vTe+46RYvjamUyfEYma253LyeifZtwMRD3JyIR5zdYSi
rtk9h9jMC0NRiYjbupATMnYJ3Tak2/EBhPkB4a5H8RuKyEdKwP+6K9SwnJK6vnM1
DGkWzdzMPtA9ss0RLtF/S3rxTKmJcUqWZmWkxqlCAnBAu1k1x9SmpOpuzZD+vI3C
DfSGiJfSWO12gsq5GjyNoLBn4RMQc3q41w6dBALCWsVFEnrA27YCwZUypj+N3jMT
WWCM4q17JVta6FrRswrmblZ6BEJTFPwieZu3+KkC0PdteVB1IKqFfDB0LFk90+/L
3/W34auDqLnIPDUPBbVSCd9FGjs1sNOe4wpOLfymRHCxbMPS335WfL0ZHQBJJerK
VN10ypgwrREjlL+6sk+1GSM5kLk9vAcgIqiZFgph9fQQG98geRF/g+bTdXnDF964
elWr15nKdmYPsqP6haXSI7rIB0+tJYftUyNRqzbZlsYf5nZ86WAhR5lEUQMSUijy
UOauDJVHFxFvGu+6t0G8MmBBIW+Msrv0gwLvJCCm5AR/3luTFKwfhr9QTPaNDpXv
89IyfPnZ54ho2iGoHW7OCB+y223dsLoQPAhXY8bgfDs3XKgtt/uyXV/RQmBahB3p
`protect END_PROTECTED
