`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4oQCfl2QOYFSwNKc8KDb0k8rDLDL7X7SsXeWl4rZZJ/3+stwutBosTh05x496es
r1Y+Hslg2vWSQOHUO8yGu4owFedKfGWtCerwHPIlvoXpAnMmlVVyP1BtlPianUWI
jp1AcnClpXgLKBh+YbgephFcSg16+L/3cqvNh72DMJXn0Mbinu2hoNyAWJVS1+y7
pvn8b/AiqkwwZDjocYPqgYT6tR47MRtsfeWoW7EhD5akA1a+S1AllWygIgt0NHGA
W5zezBctu+m8yU1VJ6IGAkfxqceVF9QJ1f46k8wJeLjAGsAE5dn3lklqDE2X/aJ0
N6y6jyZS6MSFXNr/7xwz+Ws7jVEvENQKQQQ6H88k4Ga9e8vUsSYxnWC1TjcSZiPi
b6tTlgYDReySCJvmQk41BAp81JXON3VTsicXz5bJYJbW3UR6CgOoX1vo/IGc1vZa
O5IlZarYnuWOU7eXmFh1Aeq7IVkv3a7jgzBNHYSenyDXEYlnWBw1fqku0bJLYu1y
fLxWisafAB+E5ywywN4Pjb52unsI5OKjV0yHnyq0sth0xUEqSfzygA3QVvvUrbrq
VLd20oTfkHPhau2bawbDRYGy8mcvTqyM7lrjyvh2a31erwZWVMt1sETVEOQ3y9jF
bMirxb0/SE9lUnP5vGypWtUVi5sWd7JeyanZcPQ3t2gXasC2pwVCY6p5Ywd6FoN6
ZV/Gnsl7x8l+s1r0am0catwen7LD0NY2SaKZM7BlaGuCGOueT4M25xxcfJ9bLDnl
xoiY6BP14Cr3NJH0KGXYZTrUQx2RDvEQQHMzuOlLKxZDZP+Up0MUo0F7RH0hDXYG
XlEUS0T4lAk7H6PkoYT65HDqeMH30AGvsr4/ZXXTMMQru7vSf6E/+OTruE7IkUOC
Ed7ew/Oz5DoESsp7hwE37iJRTUyt+k+5TIxtZuJgeVYD0lJjetwFR2XR3zr4GSam
iK3wgufriQaHBxQBzLwZhEZngXsmCgkYyw5lGYItgddjsfac+Ms6YzZyTOljFnYp
acqBPqHjTkZbc69F0h6sL3+1T0LjDhjbsvjYBMpR9lFNdHLwfbrlPyzZ3f5q37fa
+M3hfm3bY0/eHgbQajuYTyofxSV2FeoyO2YjA4tKfNy48WLaTOcAqlFzbxmKNLXE
RvJvFr4mVAP7UbrvUH4cc8r4ZslD2YS73ertvIcU21qdihKxWaEcXsEyFUoWOsSE
lACdkyR75So8PRdb4q4JZuWRZBsrOo9BJprEbxCbg84k6arnYQt/6jaNqExYNRNw
itCkWPJBGU+TDbxwrkcqUso+d4sLgNI6oyWgUrrRkEYR17ick494o5HkmZ8ZhzJY
/lvlYjbZG4ZmDYYWaJGSnkQbOyu+iNqg00BCzqLJ/Lj9ZnmBczI6K2ASx0kZYBy8
mNSPOqKVCocxDbGQAMjIm9CaHEV6S7t0B2Opo9NfAMCL+rYb9iSylIAsmPdsAxK8
MdePqTa5LUHw1KF2Et1SvniZVP02qB6fFFkys/T5hxTOn47rZcUa8qhwHzwT2icz
O40BiJNZe5ZEPVV6IL1khMkljy/KQ51Mv66lzCXnUDPFalCQmfSjS77P79J/ee0f
T2xqeehT/H2vXjQDWR5wupaKsxRRKEEKmY7hj50sihwHnen8eq5j4tGz5HuwqakJ
0VrH97A6bKmsGkO0Xnt3X7oy3sx4rty12KiDAdWaoXTkJToFL1oJjEIau9upk4k3
BPgyhTCm54/3/As5c115Aa1pWG262DYrn02Kd98aGhiNvTmtmyPODIQpIA3B+qca
qutPkGH2pECiaKadeTDMSWSTvyLVoMBrJVqLzdMsPzNxg4eXM0ouzF7NYNwBWi1x
JDkHqojPoC+LsIEDK3Jsw7ONu44TaPdeXSmSjeOIZgvfL1UmG/HZBjLtvrfm/cHE
cuu382R6IJE1UBS28WIsvOBLICdQVVAHh5DYEtnO9uvxM29157K+1lCpOcfy0l73
BFwegWiPMj08Fq+XjnctzEshHTtlnTx1pC7do+2FIzv568MITGkPJtae9FJ5lxye
6YS8I9Sr2Cmu19xXs/NL5+PxzbhHkzMOXq7ir5hoeaX8NG5gpfD5LAzgpjdr3sfy
bpiHC/AUUF+kBB7q0WJG2bWAbLXwiFQX5gig0NPIJPrFOwgwxdwHa9usOP4pAmrU
RM3ERduWOkce0BhITvgecAvOS19OjDUOZHXUk+Jp7q0NZvWyJiXfgk82y3BSJvMR
myMjxTRvBOrfMaQUAUvRTWViH3Y2FNeWT5JbFXauAVRPpq1M2MEEpBWTPn1WOmPx
aX+y2GvtYgG0+zJ8ZOzHnQ+97gamvI/sXszwXVbEiDnR2KQyQkJxT/huopezUDeb
AlCKV15uvu5wTr4gmVksdtZzI5zY84fpl5cOBwPXo9utac4l4LDnF/0Pezgdi8YS
om92oBV4fEePsZNDu49ZsGt5B3/ZF8MdKBCAyRWm0iXy/dlHscwE45I9S4qslRHo
I+gM6QFLtXkNAnBTVbzI9y3wmIryoTzu988/17+at3vmgJGNkEjqEIG6XUqPAtL5
CbmlBwTestx7Y3rTybv+4AWzOjcn8VgyuK0iz9bToYDZxmJGA3SN6gkYcktnFj/2
EYFiDdSoeKhhDgdG8fCfZyTrtBQ2yKK/IFOEr0eGKd5sk8KkOuzV0n+vf4s8FhJz
HkejF6AzuynIJP/LSogmcgj99DObLuMlbcGQ7aQ6EApVNOqPQLFQUT60yUlb3v7B
ejChB3d6iRYVcCODupYIEs3VgtHJ4SfqfA9j28e4syEdyH4L2gUUJSn1DHn9hvWE
opcOaWQbOffW6AThy59v6pg/Y+/BsbSKfRkhyzBkFbo=
`protect END_PROTECTED
