`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BhOrkaMs67P/enjREmSvAB347BDbHW6Gw4U9WWLTGP8S5d1IhUDmJSak0weg/qNo
6dyBWgoB0XOuF5FABivmsojpeVoUbG72wy8hxuke8YPMNbPre/s0GGhL7yis3Nl5
W8MsYBkloHMhAjv4cfGQJFMvpz0TLEu3ejbi16YsbLA7l/YUDxf0M0Z6jGUphf/a
kHZQNnYNJzH2WtQGxyxE/a/o59DoRHRw8ybx3GAyBYY/rYA2ZT0HO4bfZ3ho1ulz
ll0YRZBT3MFxUX2L5oAJ6NZ1e+oEMY1y56wnbydLQCHgQULNa4yprI8jZD0B2iMZ
Lww4r1vIW6rI/EUZSyBvoQQrTV0nwl/U7y4mw4LVzYW22CKF4dfadqLFW60Uuph5
1ldZehdP81z+qw6Bl7t9jxvr77YKuvw4nBSDach9TXbbws2Xe5GykVMoRJRAaPjm
FJ95jUfYyH+7D2SjnXcU/WYtGq1Vb15lOj4UwsqUBHeNyukNxeJkgF1vXeij2mNo
dCSMs+LL7bkbtjv+HBDkvN9zcCTe+c6TaYs54bbxFodzIND88NTIloMdgCAjtmT0
Hjjy6dA+DuWco//EOhbZPzQxvErDhPtIWMiIBJKRltgnLvVoQOVcqFeCjPR3Aa9C
nxs3/3IQDd7j5ffbAilSzr4rRuJbS2kQN2TQIWwLA5dwxAB/xQ8bR0GEOuruy802
`protect END_PROTECTED
