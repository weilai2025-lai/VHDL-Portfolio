`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cohRi9Np6xbbd5nb7X34S89X2W1a+mXb+XVy1mH2ID/SlaWUWP1ihdkm6Ap8UZ+
ObSGM9NNwrRBTkFXXeCCfnqNUzIdYy6tpO2O0FKTrvlgB3SVCCnpzfXcYxnOinAt
aAcJDj3TqiEfmRn+QcdO98KyQqa1yM2BOULpV+wb+bOmkYJClaVSsEyI59z3eP42
2CyDVJbt04FAD7vsG+Jp4ZoS2r4xqW8vzp5Asj3o+XCcsmi+NucB8/lV6YycQYTj
gSAEZonbIGrYcMvUXQjKG1sdCo6qxREfittdVkuUkLqs2NSzPhEHqpAhIRk/IW29
2itBNAw3wCbSYM9PZu1ks7zDNyv2w7dwQ+pSCmIs+BFXqcOXiQdX07dt5QgMgvvC
xq2pFrUDvRwmA0YaZ602kfXF4EkEGFiHG7lLHIjZ6beW1I59+M3bni/5H8Ex9/k0
iIhgYpUpwwpMrDRDPT2SU3PYdGXigfoEYuyKDmD1jD8uBnYZUu0XFKfLjssagqGx
OKQj0iBOjrShAMF1hMzEBssrA5XQS1+4J1QNNsxmoN000uY680Fb6I+OMMepQABo
/JHc96YHw8zfz7W4+h6v8uLJJqzZ6WsDFmRuUWoTMD3dMRZR+lyI1IDHGO4g7asS
Jhsaw1MB7dwJXrSYmSO3HxC6jnhhESGXPxrrDotat4nRCYKU8nS/L1mb0KCsE0Bg
pTgVAKY5tyIhLJ4Jd+7UBdIUabBS7IP5hQEe93tBCgcVJ7VrYXP6zuHNduW7JQUQ
tp/i3cQ328FAQSO/ScVh9IBn7SAhSA6VuNcL59M0Bhr53yqhR7Joqbc2rBw0Bvof
86rXOqKk5B5zoLfz42STYn5BIMgojOftRt2ZCWa4TeS8PyiuSCws2W8Qd6so5khz
wDwYu2gYwdf3muEoxDmuDyYsyzm34Hq+fuW+53a/NaJMzEiOHMCsxb9IfvwT51m8
zZ9HjiHvtUQHxy+1b1+BXPAqwduVHnO2WW3zm7SjrV1sOj7ecdwHcxE/ZA98b9DD
OvYEsQroOSVKEAez8MSzQ+et13xZoExAvFXrxzKRw7axqOA6b9KvEmrVEXe//wDU
UWt8omRBgHUtPlSgQiMrEB/ThOSMX0tz/RKG0cBlBgk+tzZuu4Xfy3mAU7sCQdsJ
C+sll9HmOCMsTVGkAzLBHM+G4VSWvfLwA6dMlBjz3UwUmdd3WWPLLCkUWTiXHdax
jlnJoJBjjohpSEiCSsD+aGgnBRrKzlcjfY8mvSvfaqhyWbk+zapur8GX3pL8E16O
vucPGx2yr1rvwVbmE3VzM4q45+Mz0I7NiNcZTrQqEAT8dMwaYQY9fLugEKvMOhzY
yCHAKTpfogc8Qvw/3aN/S7cMHyMsgi5O33tsOiHLiulf2sBS9gF7jT2HS5WZ1/rD
9ZGm7DG9VIgbcV28NxpIaDbVWmt2lwjdHjg/geSS1XaYdlqLY/Yl/I+fC/HEj3mk
3PhRIep1uL/fuVz2R05iBFXSF59HwPOxxDZbV1+1/DC3tvH/WWb9YGTWmSYNAfWo
3KU5yzN598JfjqExdzkZ8B50DGds61oTHm/IYx96n73giFB4dJsQvwga82s2mFwJ
XaMKvg2/QJ+zsGUrghgariinupAnyBYOl3qwpPPAZjL2svNtyRF/uGj/4FBloFzq
BT3BqjvYvgAWhREa+p9hG9lJOyb1OGOd4EFKu7si9zguroDGkWlzNR3fCFJqifYu
rIoZLQ9175+UpruZLdl7EZFrjEKtg/J7Zgyrs2ZhZp12C67ktGqNxupv7dxUsGwn
a4mgYUKdO2X27UwCtbuB8Eo0K87zFcEfpljzUxZ6UqQ=
`protect END_PROTECTED
