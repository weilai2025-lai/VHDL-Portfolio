`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bI1xekDX81/UlEUC4fpS0mZMWhfEbtv9+VKiAmtVVcQW5Wtuh8uN4vcglKLo4qxJ
6PbfUajF4WOuJNpRYu9CDkS4s+qZDONwQ/92erLwwWX6KYFjfTYSXTySelhzAiX9
ZgbjV41zC0kdsHhwCH3bj7bRqKiow1wqOB4HBYYqdfDoaIHMOMru2h9EYKJvx/LP
1SFRNQP5r/lJDzuBA2lgL7kJE/GNjiNqYN593vLNHEtgbhF+09zQn8XnyvbPVVY7
nE+JXVYQ5th4grl7nCwrSnOpiV6sSxxlIYCvpqUvkpwdz9sxrdM3eZXPFUM21EW7
jLnc1c4XgP5bYjYQhmTNplTwXGbGBZLNxKUgr2pYCIdpb7y+z/2cHLZBA+9qNwcx
7DoaRaPl3fLkNEpX/w2uGImi6Z8mnYTO2BGIZCn9rt20xnojz8XmPJ9aDYoodGks
sm7YG0Cz1J7wQq4RGY4dtANz0ayVCVZk5t+o8aCYs4e8inf1fp2qUBh6TJPurmyj
HW6VTkc95ZRAyjgbE1O480JyPbUdMoA+rw4iWpj7OF/AWka1Mq78ZiEmjNlrvV8e
n1n2RdsMwIV2cnSFacdtU7pF72GNRtMMytW0N6DfY3VSZQ5UOa/8GgjHAVQCNe74
bDr5CTE8C4zgqaSoroKLEd24eVKVPgyUfU6GjQfIuUl42VYKatGig6jJYD2l4axq
+C/bggJKzvGSFhDGr/kD4a++ZQIsz9y+mPZ45ReLkLFIL8YYUG23wlYXF/Gn898I
P3OerbgSUt2h0AWozOkGf8cYCnuO8DaCWeOMsY3HyuZqBDNrURda698fAdydMHto
PrbhsFSJMkXq+PBCeCK7pvC4kho9v+ZVk3mskmjeB98=
`protect END_PROTECTED
