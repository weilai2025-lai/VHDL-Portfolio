`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOS4sNHPg7lSb12GHvfXH2p7fdY42RBTRGuqiISj72/bk98sELs0M30eikaQMQ3G
sm2082dQlkuBYe/SDpAtNYqz7Gda8Fe+Y3hsZj/YfZR8waPdiRvo/iZbSOzMZi5W
EyCDxHd+ecoWC1gedyMkIlM08IeCZEGORYNv12Iy1rjOuvAbRw/gCyU6iZ1wOVnj
QiV9/9FJvI9W3UoUvyHh871S48TtEYxffHlpMwp+ub04guyVcE8wRGQT/+wMd2+6
JJGo2Y+hjZEVm9ZGLK0fSHinX7YJDD7txA7AY/5RNEX64XUzWV4B4lm101nFbclQ
rjxCQOOAta/qjzeev0zhuWOspbBkbbp77ZYAwrKNloUME3SuPcN7Wq1EJYNw6l+f
52DjLFk1gqfkoLf0/jypjfSFfkI69mkV6mIvlCgtTjuqLUWZH9As1Bf+Ljw1a1Vw
2l39khwacXe2Ak9k+tvx6GEFA9eArjxGZELU0eOh1AF/AQn7RIrfzYJGrekXsRta
fZahrlwc1tZZUDQvm0+4/zFknv9GCL/BgB1kqHUNeFztyoR6rMD6sq5SkLEkq23f
AiVV7JbRRYVab4pPU0y8X65N4UBL3npICrYJfQ8zLasgaCzRoZqzI+ToTpzSEwhw
0w44JIoZXkUJOos18wl9Y4ARykDSiZsGK+wL6AeWbWG7odPHMdpChpSN0z9u2p5R
uD95ruDSICA5vwSV+F0pPdD+hYyH5ZnLES/VdLWltoQ=
`protect END_PROTECTED
