`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35G7I3jSHUbuV2ReE4T0ig/xfhxDCTl//D6YWKZSEGo/hgnIhmn0voUbn37HgrER
1hPhUuIbR+MBF4XRH9R+M+58KwwUOsYOvRweLEkBieBWhkNG6WosUH72RmWa0dAb
m7M6CguKCSpFoIV3s1dqO6Gt/QCbAPh74W5ZTdRFCmwUFuas55qX6RUNbEcJHp0T
ceJFvJDwt00escr/hrZtfjUjs5QLP8eEpSz0GBaJgesmFA1W3kGU7SCyVlOllDCJ
Lgk942m9/VwmB9hnqel3sykHbR+8zV8EyROWr5+qnnkdneBFMf+b5Dk1oNDXcWec
cf/6+yjqwR7FukHiINfJ63TuZqaHpIwlFPEyRKpVzmdRVA38Xd4ut5OsYnsrskqb
wlJPm8CRmoVkN5FFxVN4Lpzy+e4T/khc3oSPk3GjkDAlf14b9VacqU7bOdcPIsVC
T9nLJI+x195sRWz1JQDkGEU4HZrHFALT8uNuxPc/pZ5lQuQQoNNOelIPeaOEslNs
EpsAvi/TcQWvbf6n9g4PhyvEuPZ+lBqRY1DJZr8TcwEomI4WchLDL9T19Pj8tLMo
/Ht2rEmMLTDbhfrJqCo19JnBTR3fZWgL5SZCFDQB1yDLNEu4mjpzyAYbtwE+jaWs
7oVCG0G8rWFDPay9m0etRJO3vtaHIxigkZtrvFWUGM4CNahWBTkyP9/PxcAHLXIq
XotwvraKJ6SdZ12e4ijqrFCVV9dTmpCuJe4GGa/y8MVS1Tq6YFvahmnT5uyYEi9p
JL0bk1d2njjOp/ExXDLZztAnXZVOgogrNVuYL8A+1iujqBSALOyTt4JPX3YVz2qq
4GeROZPTxp06sVWR57ozulG/SP3Qdzdkz+XmIP7cLcc5D9+axNjqSIdp5tpD9hQs
zzGirMkFnldmuiRPjTA7N6EF1iskcOv8gsHByzUmpwbjBM5+o/UOLiwtOslNxkQF
Nk2bS0OHLlQ2IbdlZv9o7euC5niQwAzjtN7IA9OHGLJulnmAZNHQQjhUihli7C85
PgEKs7bALVC1k6spUjcEuvcGjrV+CB71v6gqVtYEYtnXyfxHvTew0lcdXqq/HLXX
vho+jQEMTYOOPelTGR4tzFL4W0tpJTLgS0SgVCV+Hwk/IbAnykFXlyj6S/+PppTX
9n5Z7Fj8xumMuHM03BTlNzKuj8hpiBjgIm0wHFLXAbyPYzLpacLWa4Youa598E0n
/OBrrypfzpvJsFUfXWCrL9Ie/q4MSvexBT6M1+ijwjj0BstqvOIPcW9YH69Mdchm
vHe5QpapIjwoeIHWZuGM/oKBa+8Y/lpkES5he0VrZPdXfnO6em2ESpxLBvt/5vSu
eBaLuztvmgmruVaPBOIuEuSWmf4q+rIhnGH8fZrSM2fg3huoh66YTej4sW65KQap
3E4pH9fMku5DxfirQyubAcS1Hi7qsbJs82hMv4bZcHzWrq0RI8QmioAng/vOZuq9
BD7P/IM31xsLi8SxjfNI8aUHIrnmSGCKHRLw3fec0egSRzA+efQJbIGrkmolIr4K
ODhSu2bN4QPUUqZ/FM0zyPIsBt4aYPXTFBcGyEuJnkbMEBQcLVozVX+I2lsRjsky
+jypWsP+J/h+BZJyP0cgnX+py4B2+tbpDinrJScpoJL8u514t03ZV7OnNKp3aaPV
5Wr6XMQs2uvzli0O1EjsmKnfE4hiTqrGZvWKkKupb86azJ/aO+hBr8tePMoiResx
PMOfj0RhytYGM60BR2LkNP6H7rR7/D3HgUHJXR3bE4cdzrP/cagSNjLGEp2iAQTi
HC2HKwwehxTb7ph2NRDnD5AINz6mmhJfPvIYfACCm2m/Dr7xLSCK43Wz6354JrPN
LkTtjL9NgWabRtkgNWtYwcK7cabpw6FoLNsgsXwgx12df9XA3/Gm9b1gnzgmqmtW
fvRG9O8A7LkzqfnabENeOK85XNWbdBz0qjz+7b0aNu18K8ryFKsSeQLBTPiazGGR
xz6ZzLfcphCP91b6ZOjeICnA5Mqo36R5o/svr4YorgWunZgJ5uBkzXftioDdoztY
H/3T7A83gDk1s9uGpVBHks1LN3phYNaAwbi+pEn+RuKNWsT5Hz4/uUbgsd2KTbhO
tFmcqfkf2H3R40uLp1dZiLn0Av4QEP8j+rI8YM94b71d0t02ZZWlCpBn3jndIn67
VXV0Z/hbv+E/FrLe7qKSK9eXM1DI1iqeVf86tjQlVz+9smN8gOs1iO2OhjI72y4f
B1mWvKebk/9+YcyfvZyrB2DRSCBqEwpz9JvMvWZwmV80zP5jATagtJLX26jiLueg
zRnhDZ3Im+4zqwIlFd+uUxAr82+lCLQRjnQ/VDbqIFokZ6iE6VWhPY/8xcc7qZDM
Fsc7jt3xkrGQ2gUna24UU7m5Yi/I3S4BkbgTd7IWKbFu4O6aZwAjiI4P6vIvtkwc
CqcueTLb/J7Airs2FMDyqDYmDEEQ2sZGq2pAL6f1XwMo3URQSjgsDVFLPzolEgLe
WpDcq5o4HzofryfT3AXFIIj9OBHospl7m2buFbkW2xMyCovnnpdRBQgH0gufJbI7
BASexkTUKBAE7VlfOf+Zi5LFq1xxFsLqpgybFQdMB92v6+WXFf0owaco2CbnAtcL
yTwDBAv2vo4o2gv62nLPG4sCgxHsQ/1NCAUbIZ/0KYN1Q9j3gMrqalk1PFk6WJVj
eCj00eeVh7oH+D4iwE+WGrw9AX0XGYC3s8WRr7Tw2b7FQPK0ReMawo6btuWpN/Pf
tVCSDQIoe2zHhwb6SHSTMwBSTS3HACtSe2hlHQx7ZbXQhfA0ZfK/KQoO4QUdswLD
65bWbLlNQfr61k4cft1nGROGHjRg9IyCCkjOj7uRJ6yUjG2Mbdykd/eqd+gfCMnT
LSaG6KmxsPlTQeAt8Q4wi12Xbj4O1nuPWQ6ZiMm9DwS3Jn2nzbhDMNj4eJl6Aivk
EbNspvcjfhivKoZNzZnH8D5wxUAVezl9NQ8BrCm3QFTvla4HEkkP9yH7MDiO6jYE
gczkSOnt3P1wTKcn2SAwJNdWC1lLtygheGwPpULXKVKqjFdknU8PajKTy7vK7Mnu
wvK1z286V8vUs5GiGrGcdKu7yarltScF45a3kPh6YRr1yMYXC5Kj9zKxOLAFSL/J
jq01208vYT4gTxgpO7c/u81Uy5w1py2faNK3GbfoeQccYUA/bFn0ZElo6zPdp/YO
GGz1Epfr/yg6Z4R5Fk0EEOEKZWC4UId+IOFskxm1ZgL32xmIe2106pATf+yR06dE
hXUwiAyUwWWbWN50LGjFYlYz7XPk10kkDlKJs+nWbZKaGrxVtA0SIZW3xoCTc4pT
3X75s4Hbh+gZDtXBY1GYk92s7BZNwBaheMnjranAJjHZsqsvXJhwhG9gJDZ+Sm2a
J84u1sGw65jnN+3eYRF5O5X4Qa97kFJMlsg/+TsuM5ARl3/egHR0imVGNmgwpFrd
cY1yGIaVwtP+HMC+qCrpcWfBysUKMqlP/Eby4hYvMWQ5Sy5mmaXlxlsU/jsB4SYK
QtlN+qUxu5iXLz/6m65DKfwKgNe3xEhBYL97Kar5Gw6+gFCy4hMu+tkmOoDX5QRR
hNixyECzdhrLNKFAUYXeK5NVfwy6hB4CNmueZy0VGFr8E4a204aAgqkKeIpLrJ+k
SspHLw7tSXrd68qYNOAaYNpU2YFdbdNLx/S02XixEcluWMkCmSDSOBgNtMORsJq+
TmpbJFMrhyFQ7Xa9R9kSceUa9j7NwgYUA9VgsWZw8+AN0aPXTMEYYfSA3nGqqF9S
uF2mNQtcV0Tc10CuPuAQJr9bqOMjeaxvclXOBmNKjzvA/6HvGItPcHs0PQOSxZjW
dAd6PY8mz5qkIpVSzxwicTWyCd9ZFEI2fynHopybdGMaAynzY5IFIu5Au9AEtJPB
W59vqXBoUAsHuu3mYNBKRqdR2jBdkmHf4MWXjux778WfpsYzGLdYrsF3UaNqPWS1
GDAci2ZLn4BBJQSYJu0pZIP5HpCyy1nS2Ev2yuCpn1D06NWOs46jkskLpM+8NPDs
u8N/qYl52m7AzDL5uVIxFkJu315mdtIyZvM0jBV2wkGOZm2wlGvvZO8UG1lWhV2m
sAbhF9ONuTlmDGQAAim5bI+4szGpif9jM/QUUnGJnLVxqoiExqR5lO5LioSUOu76
JDMgAqq7ZcPMbHpjDMLjIl+P8OW8N6H7/Go2lvj+UqMdnrdKvFP3sZCP7XcBQqBv
YKFfKPCOHGyX/eCm73I99sAV+8PKGSmhWSvF2wnpYotssbYGQtPBsFtvDxPXBinR
f3/wEMDli+GmCsAEHMHwQztnCscDhnS4YoJUbH5cU7Wbdhej2GU3KuhmnHu5jwTv
YzPuoPZR4vtAzadq0UPWCVuFsqauSwHcmpn/yl+sU4m4dEIo35FXIEO7yI5hm1gk
aux3m5N++CzTHFIq6Vh7NdR10GcE4GeMavPr66HcNV4P+Zmx4qk40CdWYZKFOrb6
96A3n7QQAlGIU+gxJ+KJu6oeMGk6ayjIc0v6PutYJXT3ntgy6lZdcze8Re+1cALh
jBrtMuciz9sOLzgnvwxyo4u46/HGjb+W1Rt9doecNdRZUpaI7YjwSLx5NBS5pPur
vncsYex4IbgkntDaWUilJ8lA9cmTIQxMfJybHospt6+8QX7JTeMepuiFvk2Til/T
7aW6tZqkW4NtnqJYM4V8j2N753zDZZMMz8V/1ZXOLgTwHE78UtHLY0b87g8JwcZ4
/OPEl1UtOzHJRKuQm2DDuh4DH/aOoOil9iFAr0WYCZEpHvuQeTnE1U50fbdldT9y
NzK9Y20lWRYRiqXB7gygfEjMcX/zX5rqDcW2JSL163Vqq+suD2VS8zk47v16g4rW
FsKlAsVRmBceVfn0/34XIJr4vz9Rl1FYRN2Ap4Lk99IfaO2VsqqJGTNJ4KHqBE0n
vy5sySa+aRQZkptkgG8LPSM6pJMX6vsuNeXarfbN2slHj2MkFWkOGde9L6hba/N8
6jljb/TRsLMmW2rwj5H/TNDVx3keoDsmktOc9zMn8pFISvBFSPDWWFSoRXz2UEis
JlsnzDzhwuLEExiJ5NRwMY1QTN0Na5y+tkEYidS+FYok3J1+RkIyzTQy/nXRB+LF
etWFt11n0XyKpC5QDjDF8sH1z+BEhbCaIh5hImPKG54mAjxlY4sDpmciym/P1q5+
/n68snSvOoqc3swpS4Abiz5uVRUzU9wbgvlrWk8sLIVADBUhP7k39uFMDpvKFIeb
2c9pb7V+nHrnX4ylL4BvxDdzQMNEsRhcy7IhNTEvJ6WFUM6BanWy2X/Sqfo0N6t9
kSlbvM4pZzVA6Sc6aYabYtII+q8Qfg2eTx4au33fCzSt5339PSgDajXSbQ8aVIVw
mgqU55CQ8HatZD5kEmkdEP2VbGGX8vYs3cSOt4JC2wyWHYk3cs5POzek7+NSVZC1
rEjctxIYDN5evbS+Vdr5XZBo2QYpkIcS7W3RpPhH1qeE8m06cfEBnpP5dnjcmkjl
A0uwkK3Rz7myqEIiwlgFgF9oDsu4I1O80mP/S0bojORz0MkwhIJyiObizplmdJJs
a4iZKb3pK67hh2jXm054G4BnAeudFszlv8ESqF/+aONJS1DJQOw+5WFT9EbBfelE
imIKCJNsLDsBcl8ojJFkJ8I5DS5zGxzaDFN+r71lcQ+7i3CxpNn4brjvBsEXmsGg
PYJMoVH2FAdv/4nqrbJULbwjcyqjPpbEpA8uI+TGQ6guLWen/vmpz9qxT357iWeC
8lWAyYZDe2OnwFptAXZUguxCt43Ga94Cn4MpEiZ4qh/Ehh6NKgLCb8woC5bdhnY/
Q4iSXW/6oWNNdfgUOfUdmIN2RGo0dcCKHO8TvcE/rJziuxoSu8eWveULCW+8n1dy
7hpk7TIEQQD5Pso469aBzz2+kLPTVneGfBoStNwdq2LqVt2xaol72MkmDLbe/2E/
MKPyLZ6yLoX3zEzpTNeKJQrXE8Uy15CU/nTw6nzWoDRNTdmrZdE+LRfUptPjc+Bu
S0sUQ8xvOzlYnoPYDjJbyGxkKfV7zA21JHnkxy+zaaz1syPMeUfXhdUhS56r06Pt
wNn/IB5gekSIB3cC11iQqlaGICKcUe37QbTVSO7rAWG8vLNaDChiGRJZ8GXGblSw
7t29AkBuQVbeAahehaDE+69cjr8cLWBCmoZ+eOHV8e8qdgKO2VW47u897w33D20f
FxIYJVbf/0wbVW8Te4Ywn1+Cv3bT+M5xFYR5Ta4i0e4j5ZriEoyne6vTLZXcC0+y
uTVVNPm0YZSjcSE7E4NohkuEdNbbJvJCcJhWNFamIhUZPKdMmG2BZeGgACULJTbb
DN4p6X1UbVZUYnYJVQ6Fko2vojRoCjb11L5nrzglGkDdmSRVdV5AAd6arNNxBA1K
IYGQxvoAZjt3ui4ZNDqAbHr10JxErdZ+WVe+DGpgl+j+gZsHzPoXkhJjGpG5xpUN
d3ybuvADaUItFb60t7+H1xOgJ54CQJGqyC0VF74vDtkyBbZ8g1uZD9FpfoO1lfb2
guntdXODj2DbrqIY0zuDWPKP8vr95vDdUNlYA9zCWpdV/wdKPNr4RrAdtBBG+c+1
WQwT83OEql2azN6QP9ZPS8LfBOOn1IeeL//cxynTbazjVGkT2AxthYlBXg9PcaXM
spQ4b+8jAE56SrhcQcZO+kwZvm89QGvFC8IVjZpVECG74cvv5w7/atPrKr8wBlpQ
Y2adw5Y5DGlTWqH+gT98HWetN3/Ohxd82kVgHjiyhMK93PBCSAgCDaxbDCTUk5uj
cczX3NoHLlvHWkYk99bPAGj8cfi+LoJAABmbHdM1fb2yNkojzoacR/ZniCB7ohdq
V9+BGVB6DR2vpxFtqaSJrm1yjw5J8et54K1CcIo9uliU7FNjGEzQ8Y7TSD93sngR
B2orgGYMaeU8+nl73qCkT49RMTY6jcrQORXgAHKyn2ajSS26rjPFaJCj2zXH+8hb
Fz3xyJ1bphryxGpF6fmv8ot+b8KpLOQQ3CQsWEg6lIimVMkvcBy2sx8seSuHZeTx
MCxDmtB3uwAtLMF/egM+sXrSNJr+nQnokcpeK/QLhEpn48mPeKRSTDHKfyxOimum
T2ph+r7ANMf8DQXFZoL0CNycXssYAzWqU4Jk/8o8n3rjleBYJXqAMB4eunNBwlbp
h3sPnodGtGqTMH1cq99+wXAGjN3S3/jB0R8MDjpiSC+Lid7vgWay1LUOWwxgsT9+
aRU7WxwnaasTd2G5AeY6jcqMv+tuGzoNNlBJ2fpMWgaUlfzPzMIn+gkFLgCj8T+o
IFLtAh/7b2PLv9TR3hM1SBsM0nWbECgbBoZkKUqIuBPip1DCy+2C7+XSB9uAyxMc
oKEaJoNoVfyZHh52hAV4RFb6WAUqWzM27NMlhwViRklHFbqapXHGxSt1l5uGcl2x
ley00DTuJTygCY256cqLo5FSgkHXQxbw/2G8WN8FFMFar2f8jQWlY+7XgEzxe+5q
/+fpZvDypdFN3PQXf/XVIEoFfCMugWVpRYDadbVNk/p32iuUkbCMopy1RWlTTdlD
QRKYIIVHtZ3eNAz3oAdkTbZJYSUfuhdGf5QCbZo2Zvv3UkdkzSeWFWDu/aS4yaf6
sa4k5OI7icEzmL8llUli7bB0ZD5jlosqWbecaZ4mzZBy4jLOrBN3gCezEr6ofmfb
GmYQCZniP7BxXtuJQcqwOscMJIvjBff40dsjucnrfL+orjamV+T/6HJvIAVyx/da
LdrFRbPyIJGhR+frqVqB65MQbSfi2n28c5iabFywMZidKhL1yUuMXNSLh7a2Z8D8
/fo5lLZsyDKTvzJ4Zr2Gz0DPqlw5dod1SYTaLpHLvfZWBRGPMe3BscGm4ZZS7eba
axayLvz/eDl56nm9Rw0iLKGju7K9rkR4tSXqSu0bug5zFCF4EIdOGV+cvU8I0h5C
rMlvsFVCVLekLZyqY6l+LR8ZHUOx4LoJbyS9Gqo8s622i06s6Mp6G2/tblzsf6UW
jG0h7NCxiOAu8m/49wAayIUQYzcDti5BM9PxWSy068Jce/b8JZhBtdjLpE8J08IT
Vi/kkg0325jbylVEs3OHpExFZXDTK4xhhdqDPPSrlKiGreSV2b6pOB6uVP2DhZZ+
a9C2UxUNcE5Tz93O/1kcFA/3fUl9LE5eb+CYljO0iNEuq26EOy8FMK/Xc4phUQC0
sXxjApFNuLdxnX8lpAuCI+ZaYplQrXe/bin8iuJLNUEwfk4/F28Zs1yCk7JxMVv1
Q3aX+Nxo5VIKj/vy9tGDlUHlWSb1uSjmXgFahvn678+Zt2IcNz30HPa+tZF1YaId
osJ6OaY1nqaIMCm40n034IDXzHH/8W0I0jgDvCh+rODedtCfbtj0riYYIqN9x+8b
LuJJQ9MpNoxCBDiIjrq3rFveQO0l/ez9ZnE/JhkyCw8zdH4HlhUl217/pCwzh1vt
sKBhvVGQxmcj5670PYMeNhh8MsLVPzBV+oO+tIMSviIHP0DUDo94PSO19qJyxREe
+XEEH5e06F720cbI3eNBeprT7Z0JCpSHoemDp+YbWPYaZx8HryQAAZLgal5arsiH
xbURyMe0ZRBUWta6D96SBPfefj/HZFf7RojtvIlAdyrob8q7BOjPev53qZ8Un6A/
KqeDYD856qQxrHB3RlU+fyG/GIExibyiIGIeoZ9lCv2023Jz3CoQ92XD/Tyn5hHB
wdom8xlLYaXx+vacr0yaodoEvAQqFoJYMeAoPHTKJC+UWLBk3csTKH2DjHYIiK57
owuA9y8FB1GpI0aLNXNi6NHgBJky5Dz5zrBJegxTddrB/cmkhjZ2avTwNqghBrEl
58EIlnU/dnuKsRvVnE+yhMoeFMZIRAtyMjsk8v0GmeVlIQi5qW2UFH0LqR2fC6/b
tsPtaVtYxvyEvYg9sSQ5Zouzd/1uVOhVfbwG+cziCkVqDJWgg/pSwskNA8yBJ+/Q
phn0kcP+gV7EGrJe9UY8c1aUu1wacO4dgyNNIcSqmeaBSd87ZDF6x337JUaVLTkJ
52+ePeVHtKjf1AgVMZEs3uzuYl7kIMrju8mjUEBcUNZTfmj//KK47Iab9RigM2vC
k71EfJHMdVWJsgWP/069OwL5ENe2cP6XJ+HrOEzetulp6pVCLqaFERJH7/DFEceq
Yad9ig557KfT4Wa4Xgjz5t0N3B3Bh2A+f59dlpRAKpDrAfro/CpsWJUZ1pMKAdpC
6DEmM0+oc8yYtInsZGCY4nhLLl63hulGuCN4A3OTU6dOZuhDLWPHlrOuLHXc6yZB
xrhlyzALA435BW0W9+I+CbMU+qiOhLV1nJkwBLUszzlZQPYw6RfX/d6PEnr6QonX
j1BvWWXL20tVw8R9xLqb5uipyzh47EUu4QIvh/SCmsAx+uHCILpABCsy8DNLD97X
AEgLtCh+DArecXbYwAC/pFRkFMvm9ynljHZDTCvHZYLXqjVhp6oV+voASRShH8+o
C6V3+bYTlWvlP9uKBprQWxfZE8URvdDlrZxy/dna+LSe9du2t2gc3DhgQ/imlrYW
pw5R6oipjAExc+t6s+lct/+d6xpHoY3ajqJIStwJRmdaP0gqJSM2Oweo7I3tJjTC
DeYXMlbjTuj58fB6VrY6BFIl+xIA1JdBUgvnuuLOutBQIT/0EHEJ192kDdjX0/wg
FvT6ITk4V3mUPWfKvsUw/tzsr8lleX38H/fyvTM1THd06+lscD36YJGu5YM7kJ82
R626GtTQa6LNIM08NwkImsLNpNVevATAjGfyKtXP0stOPzxLvDFneR7pl4c7ECJ8
JNxSQYvfPTnvoXyZSFJkv8kTsEKqXXW36Ujd0OpSOwEs6e3RWKsEZp2gaU5P5pDZ
X6ibR4WLnf9SwFaPn5C0As7vaU1xrCQ7TTwsth03dpK6n3rJ0mF/5H1L2CatSYUu
PT7EcJVtZ3IBbtjuo+0Xlm221UlRwjm3MRkjN+YPNEnGi5vDhmODp7R7Xv2M/icE
CwxG5jLSjtOQBe8SCm7ooNmfjkMkkK1pe5SPV/QHm1cLE3ybZrcnoRTVmNvH3GFt
FVanpFbMFtQR1RsksZ1TYx8aAUVDPE99GY2+i9FKVOQbu8NUtyAN1GuDpy177v2S
X/ubXUmMU/sD82CFh8FIl5mRZ3AC1/Vn6jKwY2G3PhyvRpmEppiXUWyuKEKK8Ppa
vuus8PtcicO+q4tP9Ed1A2i5GEhS0RCJRcuOi8JVZuVIG6f1fiHxOf8n126299wU
iVmS4HrgUfxztB6zwT6N1UqQ97aKZNLIzyqoIWd8ZfLfz1LNLkAVhA4MUrfoNgS0
WAZha6bMDonC5+nLJw5G3IgSQ6Lp3FjRuiE5TBEstCI0LiuFhIewsIkPS1DcN20m
tD6MyawDNTovqcyj4XK8Gu/9/Ha9YiVlZRuHvFtBKunetd43a18504at5PD1/egK
KdFnuInynhmvjgm1dap8OCOYCO3mdVzRTaPuSOxSAqVADZ4VTAm2ZfAQLPXr2d5o
32PjyyV2vUT4IqEfj7p6+B5ALbYoa6YylYKKWrb7stVJY3KtIC9QWH+Tf8Z9/xIM
B8HgcIvFJnTWbQte2tSjc/5M3Sj9ChB0ebid9Pe5lP391y5w8AJ+V9apb+/wlrLC
u6b8+pNrCzM/jcrh4QEHGGz6QZx+xYqULGNqFDqpqip+1ETkuDWPRI8w7yYDN+JO
0lKj1S1OnrBncvThPXWIA8fm4bm6wE8qPrJSddIkmatlAMkIIzP1sRpCuZcMKXPJ
7ViZrBXh5xNNloH8vbq1jznr17N2Qe4zLVqjnpBHxpl/IdCGit+gb1E3xf+nHQaZ
JYYELjvkvWRfenWiYBLfrsOCDACUGpFAAXI5k3e6tGcSflceWcRI6aWJ2eViCeA7
sU3oSh2IwNh0jOyEVaejIZhPTlzYRU5lyGvzVPfSH6A8WdtdH+51PSCBabuazZuK
PzrceFAljfKotYg2rkoqW5Ke6Wum3Pa4kbJnFSn5TdSt4I+RSOXCj+yHu/tZT7co
OTH59F1zSFP/wmUdab8KWnCAVaFpW/ye5x5EoOAOHjIa0KrbSSC8S58LWioUddjd
onkLW6d+LuPP3H8MacvB7a576u8gYf5C8/UvC6YfXkH9h1rCVtpCu9U5H9hTP2lH
IWvSFlNuEDYqEwqcGGFA1GN28eAergWvnvxaeX1KISNVYsimzjwXrKOKQMtP8ZTO
kya53Nxb11pwHi0qBvrE2eGuvBV5P22PX+bPvidJE1mbEvCMbHX1IiSvSDdVScWq
CmIXUXzfY/2O8WNnR1RIe4jNv75JJ4FaI+caGAy+S7VobIhmTIdB2zl4e5mp1vbk
/Hlt9wpdTlYH5jl3u8VdZeXM6r/B6oN0n0RLfp+ATvPxdOnJnpGJJHuNw0f092nv
dqzZUjxjakd/LoDwFBvqvcJl1YEiimMCFFnY5864CZyzNMkbZHv3aKVYvc2AUXtP
pPtt3VJ0HpzfDEwRKMPn31doMrBy/46fctSeWWvyFTOCujfgKHfCremStxJSWYwb
5l+xGE+3jpNFaIAJAJdZKbE9W9tRILt5SghX0Rynd+3pORRoTEzISGXb1We/LeK4
1TQ6tRaIrAEAMkkmZRtJsbKhpkO0KmwbnymwyhkdpQbBbWo9XmGNmBcxTVlDQFu1
3iQUsbHk6Ga0rvIoV02gK78BsiexfscRd7gOaChtim176pIIIEIivu0zn/VmG3Tb
lOUZhDugcZPNAFpyIeVMK8B/zTqxAyQ5MsV4y2XrSxmIVoH/fYEa7hT+xuY9gxpC
tQ5+bM5y7FrhQe2iJFcOOnPm2Bkt7zGZDxb5F5Ds3O00yENEq5TewPmMxzNLa8K6
RSDXanOHjVJBIjh6fS1B2f3aDfl2bUA0ZG7wJajWOIAA4Vtmq15vvjMpl1a75z1X
U4xMGbZKx5wdl/VUWVFoCOOFtqhbPcyHILRUoY1olim/Cuz5WVvzuElIsnUMdA5u
RctAHFns2j63dCKCIS9hxmElQ+eEAcFtHOKgi2vL+YzfK7VrxndD65xtfnjwVJEv
O7UqjWWvbTCy6gUZmEVqkyRG8mM39BnJkuKY6xHbzScvgEa04PaeFe8lHiHi59N0
smUzPzNfARcGl2mcMaQFD+V5sbNGXiqqBbPrrtEyDvD6upvPGHCvNplOx67r7Agn
So9fqnc0+EgJ/VL5Orpwx3NIiB91RcR0W5JkzJ17ZhHgJCjW6YWgYwzRHkx3S7QO
iUub+Gnra8axJEVbg8BJxLZb8+5vRhngSghrGUBxdDZJTNJisSyAf9HwVDipHNRY
dSaUzrcwsKUKwglvFwP43PCie5tgXMvknS/JQEU65ogaJMDVo6BNVVXabjWZgeMb
MQP0iCwARlFztBl4qfPVB6DIuI1Cv+1ZENFbmpiqHmr2vSzLIELfrMwbso8qGDWp
mcrtetw0lMit+9VaaYEv8he9EPaqWOJJrH73E9/FmZXhB+YfUWtyG5WMTuqPYJ9M
dYgmVRtBv21N/8T/8OXBtr6CdkEYrL0ywqWsFGnK42lyV0VKd0wa4tzBsw/1BbdC
IO0eYVX1AxFLOE5ULD1LyvTY8sD5QWe/uen/tKw4rUBecMD94TJwH40k4U2hYdcp
CSrgHS+oEK+ERfXANG7mMB9sWAmSn5qVxpzOnEQBYRyR1deAg7TRrxjk7bjZ9mWp
wvOO1BV9DA5Tp3Hmlvd+SgOx1u7m8ikZCMoeb5J+9Szr9wt3hkbvQFREqO6XkkIe
FK8NhUZOeeWTbXq+GVBjyCbxYspeMB6fb3DVL+lWYXI1wC2zeBc/1rsFWuvQRD+Q
Fng4aZtRqEulxNDyTECmQGGWQOqsEPDOt+gbUfhrVGwqzi1wghVU6YiUD79kZ7dv
vQzunEt3U1o7jukuw8oC0ORCQdpbdqEdrjMDvaXZQ+DAkD5ZC0RxsxdD3/Ug6zoX
X0g0ennfT0L1KGrgFj9zXvOqo+G/3yjZYW2eAn549gkr8wB1gXrOpQPCKwShbLR8
oQPfgpDE9g5r8RfTxcFeQQLVdiV3UdwWXH3Vgug8p7Y3PNydpLKeETW2LtJtnM9+
NNB0ON3ho6L+0IJ3fHjIvaH4EU58sNcJ0cSZSVAuU/YfrmsbPzPsGg5T8YK1q897
7/PuQVQI5ttnfpBw1nduMJ8U5bE9JLZ1lc+Oyv6QJMoKFKy3zOBTWVJiXavECPy+
O/LNEy3UIMFTyBlsyWPoMe2YtiU+RZiXkgWqPR4Rxl1jvAvnNrDLeprhh/oPaYTH
6nwtSNuTeOJ3nIjhM8J+IOnI4YaddY253egm3VdgCmHQ+paB+qjJjJ9D6qNy+HR4
x5UYw/ZavLVWQKqQfXmCqaN9wlJPgmIz7O0vktff0IoQ2G2lvPhkKV8NXttB3P17
kuCCtJVKFdqht3A2Dg6k7oHLaqSpMfUugqDMw2/4srTQAcQ/pVqbWOelLZqtxBmG
cB0B3Mk3DwZZj+obJq/ZpMQUxfGZ9/WxE5xubJcMCEIfGYbuYiDH3oMFe1SMsjal
e2FZeV0i6pdCmYFboMeq8cgzWhmd3KcIPtkZTtCL+otfvbWrKcucTviP4Nlo8yHM
5nEXTH9+ZPeFuhStA7SvUADNL7uKTGouGh/KfXOwA9VtcYEgQGD9Ghul5dRZGa9F
C/hD4BWmTDzYsag2pFM42x5QJA2tD8f+6XRrVY6kKtwFiH1MzPdvN5+HvRj7WxbV
nbFqdkr6sNmuAL3tbyShjrVMvqSuRFl78Sc8RAItVarscCXPADih16Vh8S2I5Y8L
to62LgCuIxHzyi4HW+KG4LpGrA9IPraNKADHGfZeYAWdl0ZMzMJ+1K16b6cTcakV
lux2FEbFkOIE35uGFbzH+KwgCbklTPoqqS0aRPBAT45BAAFgUf1Cw+64SSPjhFnE
fzMQtpWOL/8Ai8l0QcBQL9Bpon44EFr7/nyODfo3+6ByCCsHXp6fQ3qx1JNkT8v+
wldpv6EztpIs3z5lpG6GWcBjPIYdNeO5qmfmMn6D/zxgNuuHOldoHl7BKAHKQ6n0
0+I3lilnXbU4PZKq52r9n94rLR70JQIVq6MmZ+DTSIcTuILnYVm61XlRIR09P1L/
Dhy0pf2WL/+CCy9FINvP7yTDQJouU4+1wLNTD34+tXNr6j3OUYjcbFIPxWjggdQW
P/fjP6n6s4CaeflML2MFcgTXIYoVdCT9ZRsDWV95IgvQUAdECyaPqK+zkHni1yXY
SyzUc+XyjnwgcRqqHm+ZB5ZaZIiOg6SX0n5TWvmjZoQFz1REg9G7ZbrqnXjgSmwz
wRWC21ykDH2HyW57Z2dGz9MZ/XjMhCnl98lRlVDmEccw4g9QIUAh+Fcdaa6DgRK0
Z7QM4Qz0jlgQ4QowlYzjXNFg3PGbDfVFe0JEfyL3aiza5LJfFB2E8pbNbS1fN58z
fj+G7PO1TwoGhkuC6Fw31sd1jBoxNeP2HUsaR71/dbBtSpxYT0Y1Whu+RThi07IW
x6gpexarxUUYCKKHHmTGjUUgTviuiWvKIANy91X7Edy63wk/9oYbBpTnLRIpFExK
21fu8gyoB/QQWkHOWHcrS6l3hdwODZcUEwmi3rPlMHm1Ii+PrvhuKKUZ3kXFwaux
o4i5chMQuu9VUeirpl3jcJzQVLEpJCHbQfBRU8gPheuB5NPSHklCUnnmKeUaQhEI
m/Ib7hwmn05X7yALMKz3oECcJT157oYVv/3GrathGAVDAmgeSOg/hXJpo4pukPt6
Ezqx2QoswXMc9R0iJXCM3WSeinZ8qQJaox5pdMLsFntwk0Mb/7x5Jhkpr5RLJzT5
45Y7dTvbUKt9qoi+sNVyPK7HAEBShnV82YfMfvj9TlbkDSea+QxxRfIsFsQpasoI
cJ65RrjUJhGeypobv4Y0T0kM+cn6LYeERHOvunjrF+35aODl8UuwGdSmsVipCfao
7wjP3P/GxItWb+TgcX4w9lUXQYJ+6bvJzsbF+9JX0LS/y42PrOOcwTOhKBIp0pRv
VVuwpE98kBmt7nsvguk8nUgRem1Cbb7uXqspG7GVu1zLIfkvIYr01UoBDlCAgZpI
02WNLJkHyWZBudbZMxrxfx7EmZZ9886w7upOvaIH4/7vVYeyuWQDvmvLEqU2LMQ/
gD+F//RD7gXM6DLTc/1EVQd8vUPz7AIaOGFzi5hzcLXGHcw5xeNIfdYFYokmg/CY
bEgIPJbWe+nmo58pWw6Q03e4UldSsPAHnTObmJJRbCDmos2HWSIPq9Dad6mQ3wgG
YYjnVk5XbaAFIqcimMwgBo0Sz/jD6z7ypl/Vc15ukoTGpjugkgUFdASPGDGr0Lew
94CawM07ujz3Z5Uaz50HcQAzAkH/y+3RZPPOmIPo1vKhKo/+hYBDoMi71gmtCGvg
3PzUorLZNlWcnXqnMN/H81FoOxR82/+accQUEyGRbLHfiWW6vHoBHDniwiBNMNNU
Sn9yI2AaAXfFW2Ybh7vYiwgGPO8WKeoHAErZNuoBPNOvJ1mn00HeJIxVET2zngLD
tLhvu+TBdEhUzqdMg48MxQ5D83htw0dF2hywgmOhrECXJOlgV25Zy9aS9K0czkzz
PYZk27GGXPexyWk/lPUK0Ap9HmlJ3oIFyEyxvntJr/1oM2hp90Rdr+9eL68ZZJst
ZjOUFKTYL9QEYocYLkXLl33pWwH9n2FwNMkfCicLf5tppjiq8GVVjPwMyH2uWDV7
PMAZUET5Ed80ojjpvVPtpvNxwseqTyfw3Zj2GHbK7Lxfz2s2tbdyF/cvG4F/swdF
9R244bDkzb+FezGqHOMPzUNu2XzJQFHySMSQGPkhvpCpQinHkV44HMPhMdpKS8iK
2AFIsPlei/EBBO/NU8bHJbxGrYodwUDp7qb/yH8Cp0aJRc/GkzC0caIU5dmWPr9+
cLljeSfUaXncKEzkKnQrksLEb813hLjcnmkJzZ/TIB0ntS7vU/7laOzCEGODNUha
2fVji3X1WadPayzvyPIBPZc+UZNdJnsce3mEwEedTADNUBBDd86QBGniubeI5Dtw
nDlx1aCvWeaR+mdjTdirO6+WCWknNiVvySwxA3b1KlxwdL/4fpYJKxatRBLvy/bn
SrL9xB8uMG5twLFuvHb8rwc8FX+k2ezA53piJ24YIifrkehEByTQJELDQRfWEsq8
rHLQRhbuGLlxuATBrcwJaYDeUwZ4Gpln/2rK6UWyiql+ycbYoFevLVIpXJYzk5Qq
W4FBOKCAeLCfBLRWa4qyZ49w4fL69Gsqmkm4pCj9G4njSO2qmXUFbB/FqZxkVB2X
FNSz818wPyNg3n3LrfOEh9AXX8mdacZKLWTgn4dvrJV7CQOKk/L8AmyDBNm4mBSu
eIftMzCqhbdUz+r8mTv/A7Q5SwVnnH/YKx8ep5jA398AHM3s+e+9CDAlVAZsmVCG
RAoX30tz/hSn87tJ/pYIT71icB7TVDjeta1OoDS8vRL8KIXh2Zs29I/BB12DCaI9
MkBXxUJGjHmLJBmlACJaeBe5/hYrSlqdop4u6RwdFE5M9JNmx6XxclkL2FRBQykZ
3OOFKSwjxR06FnDrMgmaL6ZkzFxkvywTu+so4igNyDDGFZajgtduS4O05sVZsO74
itrVxxkiwHn3iZl9WafWeYuGhFkJt7F2+FcmSL8St194YJaWa8dC2saCYfMPqw5O
UTXhZHsM1fI3vVKq6gCeWJwzaop8G6xxz3yA/QRFX4KeCWKY3y7au1kuj4YjIti9
AqL01/BZMlwxmBxaNG7u0MNN+HfiTmVc5ixcx/jX1zB0nSP6BswU4rCh6w2vlMJd
hx04IZRNIeBwR9dLRULqGhnl8Q8bDmzo8qHSMeWHwXmvdqX1sUGP+S4XljbQOm2Y
kz9y1EYUN8zqp3VLHAPsEe8NWFN1ud5TMgElAEQ/hgsnKC+DNZnLL1GksQOOHC9T
BREbaLkRMvGDBbfN6grRu/EHaUcNaoLzRKDTEnya5RJNmVI6j7d3D/llVbeamiBa
aQHnhvseClEZOQhE3UgsJVvTrtUfqjmuWGZYyggRJN+3920KYQj5xQKiGAA5rzMG
uJUEiYtMEl52Vny7fQlkUL4JamxcrqkKJny/4lPTiB/34YK/MWQh03bLXmJ0mpJm
pd7dUSra/p/pqUaQLS06WeYTTJGCC/5mC2JDE6ovBpnBBS6777su5+F1994JTLxU
YGK+QrpkGLws1Q6hWWi5chdZRhTprcgXXVMJ0GLpjdp8K9I2kcrnoPXZoJDVW5zR
f30EHk/Et8DNRPxIOsDi+rUYKWMh/WuavV7xQIDvuCAlqWyL7qFBomI4QQI8xOFy
+LIRR7gFEnSiIPFpN6J18TVZLX68/F5BxpwX5BthhuZwIzunCyhjO9chHYa/jeib
Mz9PADADmxmgNta+RkyRCp5DR34yoEQdDxGD4kpRcQVP2XMvxdiMF9kuacw0xpPV
7JKljN/MtQhDH6M4zN2KR7wiCGhwzLsBduLk7gR+1E47QHSVk8/I3FUM5s52bIhm
l0QQwSlCm5FKgIvZ5jVJyWqhCfjs+twCZeCQhp2Tvow0B9CoyHnTL0DFs1jouFe+
NDnAde7+eL4Wa3hpE/y6ugiYsyLOF6DN5xYfPOUySAhnPTDIYfKJ1C5ZD4fm84G3
P/qayC/UUuHaEiw5PJEqfp8pkdht21ZVV58FhjnsNX+23ki7tQwGJT48u8TeE82m
3KfK1RyC00jFD3zlhq3kVpeI6vIbI69qCHI4DZpnRRmdxypZ1LQSK9SXz4xQMEGg
AkBBXGDXTbZTxf+tr9uyRuV4SVGg62DEIyc4zQU7KH+gfu1dakFypYptCaHaVb6/
JiF0ORGdyJ4DRpHuh+Y5EU5SKxDXvJFx4Enhj326TMBbntk0XZnYipSS5F+72Ouu
opE3uD5zd4FixiU9W+MnqEGaMx4b/YIiKeO+2DZH4jqpajtkvvnZwSWffO47OvWl
UPUEZRwZJPW5hT5h5c5LYwugFb8/MeinzSqJQl6L95co6LaaHn5aAEJDq2Sz0Q22
pYNko9tSmK2KOUvBIk56NX099rRtme5SvnKkYDzlrSE5E1dCrp3HtpyFizGnEvQj
2VT7idFAipHXUzuY6u6UaUpHK5I6J42zpGebpOaYBgiZYug/kOL76GQPKLfjYDcC
mLNdu3m7Dobqlg//XmoKCoMyhOyMghol7znrvNHKy3Bh+jwD7ZgDGGI00zYx4EDR
a0YM/1BWrmDAnxLhCH+kaz07S1+Z+c2WwIaIdd8ry1z/w5gN0MsdwluKe/QPJNNr
gZPoYv/NdNI/jlg3qMkIvD3pctPs9+GkthkmfzqAAIpUVozv9SZP9A2DHyVXHXu7
qrZ5pvK7JZr8Z8OV0FOK/8PTCy3Z5/LizTwQ9GTPAudfTogU4jHpF/SJio5sFArO
dWH6MK8tzoV9qu3gdz40HAzSeocgJfEmlzVqOuVDu0uiWMNhLHjHBRzvMeeJAEiZ
PlIA9OUCXwECoGHs7qZo3JIhV14S8gJ8rMI2i8fv/a2gXXcpms7k31OjD9X9qN+7
4qNE+M/aW0sKtLOAPDGPUI8F4UlMatr0enZpFffZGpZ4dEhLaRl1cgyobpUFJVYx
QrYG6cSbvothfuH+4h08dajcb1JG6rsvaYQ6Q3jWJ52vv5pmWtEyH3sdec47KcId
dqIw9g7CL85y1vwj8HUqtVRoDkYz70Z577nOD2wUk6xQjk7FrZQPMpKpYJaNWg92
YFBZE6m9T4FPQVK7J5fuhQrLYR/9rRhj7JSQkdBc7cOo2nWzvrrqMND1SW6Qwvbb
+hwRj7AeRId+BkjfI93NLNuGN9eBFaSvyk+uY/BLC8c/rSeoJMyqFFZU0yXsf8Pj
VS13w4uH4YLZtnMRcu7VFUuQngLW2BBhavBM9Rg8iZ9WOlH98OqtE7554AR7IFhV
+vzt0tSmcB+qbaLgLpb7R7d5aLYOdfGcGoW4WO0SMVeMfSEhlxdsseHItuAOXAfM
2FqqrYfxfavH+T97V41LiScruHeRbFz/GXW9mCl2DniRMejT25Wy1O4QXE990AHE
hbPpoTntMt+60QS2WmVMprdF4fpTMtrqTfsG4EuaHRwrHRCQKxTPYTOak2KJdZ/N
+CHZXcuPgBjbwXVKMksnMv+m8lPTAdE3I0HZ+Tcjtl0SgZNx0cxF4XmDcxfGykyo
bcbWfiIuL78F7uQD7cZ2DJpVrruHI5M0QI9ZsGHN5HbROJWnvQa8Wz895f9bCJJr
PRR76fqWlvijvhzAsrIcXzuBWbz8ZZyraGB7lJ9y8AY+nacBMCrXsjQuiweEC94E
YIngvE95uyV5FMr+gTAOjrLjtHQ6UZybonpfWzpXsbv5AXU17BQgrDxgnrK1EYb2
3SBRtwGUC6nKblCw2h49pQD1peUHYXeeaI1GEDC25BtRCEEGSSTfUJ+2P04eTLJk
FFnJPMx8VYvryFdDK0JV0ldnD53zbcVpVPq5AuW2GoFBnPMjLOAQKoeLGeL+ljO2
LfQwF8l0/R51TxdRp+/kuyphrKyN4Oc50lc8f2WI881xyoZlH1CH2W50luIZLGxs
0oE2PGpTxRFQhhHNa6KiNRuxOKbEaOu7hvZb28ut889vFvAbnyJ84zPVX4bZ32HY
4DJDgS7WSY+7Favx/QDq6PZbaQImCTTqOFv1Myl4rjiGjrh2MXf3gn1IyuzIoFeh
ljpbQ3QoSkLiJEn2bRI/d2W8O/ToMTAik1psT37VLbKJ0n4MVAnrnd+SrIfEsfF3
LG9cAUjX38Wp+D/3sp02ioFFBM9VAHo6KCBXqKTE2KAytM89s714E2uSRX2mS0LP
dq1QXYk3NHoBPW68s67tx5ChkrRI+BzGztudg38x9O1aWL6sJILo3wI2teUgWUMt
XzMW0mWVsyLKVTYxbD0zl/SvsmiEDylNR926PwcVPPEyloEy3EEBFVaS3fsmBCU3
Tg3pnfF72aejw/PI9rObGhUogKpukqykOD9BmL0xmiLL9eX7WKGo2p8CJ0wn8tdc
UdqJuCyF33yV1FA6eMuItx8kX/DCwWVGP0mQ270zQ3epyEd8hOqoBSf4l+pkWWgU
4f6pDj8MMzi36WWvc4Y9spNFX8ihFofukrEBp8alnZ0l2kUavN3LduGSNzFs8I/j
ZaxmG9OC6b5VJNv1bZW5GUp/Vj3GoqdigUw7gnQfcv1WiQ6e/K97+8REBybcXwpA
isRUY++RIT2eC4f8HzXaF1BH4O8Byr5aYya7/0kmTXyM4TRmYJvAAXXpfW2DZc6P
rn1GuhMumzM6Wk8nmQKrOnesQkmZUKMDjTJryKRegMzWKDLRl5m6CZv3Z9A2loZn
j09vIwtgRGATzEQiWBOEjkqJl8K+hK4LlEcSd7KTDEg7TNfxWBgbq/bU1X2t6Ibl
sPVvqe5EvjnrOr73g5sQv6Xf0Rcp+j3vr8V3rTNmIDyHZK+hz8bbgmG2zjTWa7y/
gDaCH0PGhzlhfPBN7Lu9AeIczvLdJqVi8pjwv9ImVX7k0rb7Q3a2d+i7mFokGivV
ne4nZi0/m6gyrni8t9H6sfp3kbuBunKDFSMpuDmrA1IT7sAG1OCJYvjJZj5NHoj/
XzZHBVfwRibilaWjHjFDXYhfA9HXIe6f+zJ/xlLB1vu5EEVkhh2UIyZ8ITAWsUb0
LDHqzVl+xjQIF9TUev0wJd54zyq814hIQrnbwAT+YJeMZo8vyUeYjY1Tc6Lw6V42
1D6eZD1IwsoxWf7YJ74BGVkLnbSyJX/wxIiqnoTaVx7EkyQcbu1Ks9VWhOjnzNAF
ulLYkAkch4JrjYb5BDMI3QM7tLOJ109GFnhyhtxLUR3NYAwDD4zvqeSOT1hDHYaq
MEWuDIwrUKyQF5510PUI0D4ccHW9kUkc+Y64QClEoxrVp0xUfBdlIV7i1aGzxVPz
bDrIA0iKS7mignjggsqiC6SHD5pfORoJOH5JVePt/2sAPpAox3wZfqEbvSHXEta7
rBVdtbhk1DimJ95nTHStUBSCL9tRsSoD8DtgsaQ23XdddLUwzOLzlYEAh5ALmRcI
r+59cMRRurEP0q68Ph4gfJnJNNvpNp6ygQgGA3h8S5OWAl0teGUiU1NOs+Og5w8P
1COV+f0S7e668QRVrML7ql8/qoHWRidLHueJ4SemD4/yX6JMLKdoVTbcz1tFYAmk
WAaDbYMpdu0T0+H37k+uC6Ye+u8pwFVa43IKxulTN+d3awIpSQCqqfIZYuu9o/Tn
ps9lYuFu6We8GPJQyQAW46O3t2NhzaXrFHdQYETMMXoSxOABoAXHr4pB6FU07KiH
F7xDhrsafwGXw3PETOgzgkqs1hw/u6eBUvQ75R9cTFftIayHxh/0+dMdjOp+kJk4
Iigv7RWT6HF/mSlGhX5XePK7cIjR+PUXsHIhwEstZstd2pAruSdrPj+9mP5iK5WJ
DvwKa+L4mbyLHz0p4xImNsE1/7EklQBhUfdScDUZZhYkXiAnzUytQvPJlkoTT29y
wfU1TfyO+5TvD/JYDR2nwx9LY6PtJ7mQYOuDLdLajT7AgDCJb8xjhYznI5Uu6fS6
uok1RibX6CEKW0xkf9vdaYVdRmGHKUaulwK2Jx7a4Vx8ncuzUtbXNZiv2CBK3Kly
PT1VSxZO6mRonqp+y6OJfMUOhVaf8piDv9ti2yuARAYuGKgDx3SVGnV+poPNUl0K
VBVV2s6FhaAm5avrTCGd54UeHZRKRtI/trFTGorSac/hJxrbDpYZ513FtawpVt7K
VHtLXPEUUz1jvMrUd1g2BoDfbYx7UDF46V91byw0oWlM6a+aLnH8XiFjSwlLgrhb
TukbKkco0xqnQ6t04Tto/jHHGO/4oCw8xk1EN4cSXcGhcw5k3nkxmo7dyfOzYoHc
ABbV7+1um1mW4x6k//FdY9zvssJCkcmrm3ZjRQbe7nO6LkcnbFsIHIZ1+OxvWBiA
lb2/BMT37On0yTHgbum3APEdTgvgIJgSbn3/qIDiEhSkXW76h2QGbqRcB9K9lIve
kcKQ1PPPmYcup936nIBvxyo0LFk43LunJlxSVJORuYD3A8lOGV1lLove6+1ympqX
QCWgfGyn93pEA8fe0PogDYZNllemvUKIaTR7I2CZEglYKRC/4dA17C0MKiagDlIC
zD0SmWiFnRWycwxyaIxsrgErVl6UBf0rDRr4As4IRxCvY2cL7R6kafX97/jGUNjh
z6srsr/e3lx/JTriu8wiAAW2AGHcWB3SzhH4NzljYJnARtjXaEmlyEv/Hqxx9ny3
zmVOcK7ybSk2Os7gptM/5qVqxdN28TGhS4wTveN14I0V2theuMVC6PeZrSZUlZH+
iQ5970BasxaAyIcHPxsc9fTiQZW/uICHiKwK6IkKMyrQC/fGxXjV9aK+fbPqluEj
4Xil7eSAuFyDRnVE2LDCYTbeO4Mg+QoOnhQ8M5rDJsABOuAO3gZir9qbSpEI6xOx
tTw3WcZCSZPCh8mjzuVImZhowgpUx4akbQsTjXhL+D3wJ/NEq/bFRycWYcEIfQ1R
ENnwZAVukp8QwZiIA38FrLaxpVo/ED6XQaojtWEQdiJTOhvOGmhIHKySdVJmFSOu
KnittRUxGWNC6mLmGzLTs7NAbzMyk++TDP2NyCgOt8VjkyhJypeLolisy58j4k4h
Lg7o9TkKskyFmpXe7U7BDbTU8X55NGp4XUOG1jts28YUIrl5VfHuUgAkv75Jivos
fdKes3CtIlfE3Hy0OVPSMnXWqKXg2Wm+6thOwpGc5l8bDiaq68mSkS0Ia4AFoXW5
IZr+3Qd5kz+8fb2fl3BJGsiVc0r8frHfp3qj6IXKxNsuE3l/HSwdp14+70Qi09+4
DTbxw1USeqFrCE3cd6gSASXq8jzDBv40YJGUE9gYc0BmFGDkI2zORN+SI7C6JOUz
77VHhgPsSmZufL96O/Uo2FItkTgz8IPYpvbUtJCtjgYWS+z6BtoXdyDZCkoUlhh+
cPwIK0flrCMLvn1CBGCwHGZiIwTHLB91ghlR+ts7UwGeOQiCOgGR2CfM+5iwvmO+
ObWh6mmjxO/5+3ZevsR2sVoqCTd9tnqmMu7MD/KBQbYYevK8SIGcudJSoTFO5QAd
Zr68p/xxbMsvyPiIDoBZSr9Lujpbng0EekkwtgMD/x7lfDrx3a7e3iHrkbfMwKQ7
iohegNGRXtt1WuJJdcquRI3ALJkJEUIODddel82A/ixsN7s/TRFsw/2vWjSGU+iI
0c4W+W83wWsfUkFdBkU7XeOE/2mzOYFbYg4FO1mVRqpCGfikGvRiEWywUDuIlRhU
nc6DWFQR5CrLIHA0NkCrHlGIZc7wQ0Xlqa/1rV9rW/RT/fcczB+4WgUPUWJTJn5K
WRmEdeMb+H/kk8/qlqLQouUOzVUcfWQerB7Lj7JhG/sPf39F96KXrihNCclgxZ3e
oleqLBvp51/o/j9nqHGx4wEyemSUmicWF/feM25tQdxdT9Jv49voWVF/qi2brMST
TGIw8MdH+E/2poaw/lause8X6NaoR/QTH6Qu0kkyYRR+LdnRgeqp3hk5BLTni9YM
yf/1EDIzmfs/+3Zg7ZhcQa3jWbEYWYgBwCfGU2B9/XoXVj+M8DpKmTn6VuOd80mt
Uv4qzJJmxAWR9k14/zqR06FHb5oP56Wlj2vlFWbCAyi+AqAup5TUODVUWF2RG4+I
K5avvHRHmsXCEtSwi7XZTMKcJ31djprEqqlpLNwPMgY96ElRQBX/A3O1nSAJTsOt
J+PM3SnSKO+XWpclbB3bISrYrjUAghZM4KoE9hMnvks7IJDYrJWWW4CXjxUV2Uj/
xXZ/VCKey3qgCA+yPTGthVgkLUGy50VWphKq6ARdqY1JX+MKYe2i2Cf5wBDf9dQe
ltD2hw1M7emfJU4jQoMUAdkpAdSROGVC9S6HTyXa0hCP2DEdNvy91jK7NGrq7YfP
Lc2jQSRvFXc3kroIOjdBu/xEVwn+j/chPLOLLwvMsNqYoQUGsnuCJo8OCmytX5Dz
ODm5aBblW5WSvPgp5/I+erDMSI6beOQpx1CeaQmoonoRl0b5ItkHJmwtmljlBk4w
x75b7S7lkHdW1fRmnF84kbjNo1GihGGjpxSwxtv6SrXBRpbQcbNCcJYIInEi4aMx
/rroPkadP7MCc6+NmEdE01YDF683uG1la4aciJq/kILUq8zqWCSzs+W7Fl0OKq6c
QWvilZDEyjc/SvX97hA0KaxK7qTZa2TPTTJiDKeYn9mGsH4xW3d9i1KzjbImz8Ff
3UXcNyHd2Zx4ReUQ8492ikP5u4z1I6dWHj1spYAeelnznpA/LPll8yWxYBus1p3a
5vNhHcRouADc5n0lpk6MN6NMz83mbeo8hYa4MRKYNML+IcoxpGFniErm7iMKUajg
3iwnxp4C04N/nhrK2sN7xP8xXIFDOW2W/qEsilihqZAY++cXsAv9AA6WXR/WrYjx
oL7VKvxuyQRdiVKiNZ6h0mPXzaGTNili/RntHzqh4LiFwzo3JG3F6TgXiQFX8jZW
MMYTNiA+fZML45YF3nNwhLxhc1LvASUi+mU9HoYqEo2F2aSDoZVdGGVxS3hrcIBr
5UrPTbN/uH6lhVsd1MC6sX2z35BC+i6EBDNWyeEhnDLNLFxqaIggzOIf9XgMx+67
7WOXEd8tHyJm8Cn3tdkxJAmrnNP1SgVRadqmyeUlS3Cd+lg9PusDYtmZJDF8phaL
2TSBS6cmO5Z6QSDPGmZ/AgTXjbrsYuUqQ5zWdhyRxTJMciIKIdskRuI7sVPRW21u
n/kbvllH926km0NOCkcTOSnsRCSk8OwhG4UU4693ozxu0+f4ftyv1rXyncNhgir8
jb8WpKApt7P1tr91N48yhz2XzWQbfXP+RBJrC/hkizMY/nnojlRrGjnKyIFFT1jm
FI5MwU+Y2ip2h1Z8NpDr78Re9Uf4fcQufRcmPOzs7QX9Oa5Dca6luZ9pVD2xmVCO
vBX/yMuR04lf6LFtjpSP8PYSJZryDIlbnOdBRscILVDhJq4Jydgdb59dqNa9B49N
30fJtZAdcrS6eSjrwo5aP52NMVHkxGbuB9pymvsD7HR9Uwkf9mtXA7L0oF+Ge4zg
lvHnB036RkHrZKMS78qAPVHlP6JTu0rKWiDqUd2wxegN1Qzrhny6BBSCFvx4P4Hk
szld343xYXTg9W6tJlsjziClCzk3JgFD+zdMYHJEjBVbS7aUTNH7FBAvz/s3qzhw
Fio5u40jJ0UZmOxVydxg2nQJgQdTJDjnSp7mb4tEtEjOjDNGCuQpuriCvtfQKn9z
JbURDXCUgYnKMJH6ArmIoD/rWjWEyAxmrUEozPjI3tLoSTt6VgAKEjg7pR3H72p1
50Q4xAZgtU66D5XqV3A89rxLL/lA2BF4YCIguKcOpQZhEoRKS30E5LPmR/isQsB9
qLRsh6063PiZ6A3tdV86I8d7wVQQkn+LCQUKki8RvKcVAnNU+cOHEoFFl8s0fvQs
LxMJbgjq7ksJ/z6ERO6URwgVQD06vawkxP6we1I9SlVYM4ULhe9/eeskynt2zC4M
DxmM2qxOJUtiYv6hmAkk8duvudV8HqN2qguialjIsWrXGS5vktK6BQVUkLNF6vCM
D1NHXpPhCnsjFIAbgG6hR1tv6V1WH0ZUD4ZFYzeCWKc9lRsKp1Oa5EVNCjiV2UKg
1Yr0nLXlYP+KT9ADW+DpnlcYyXA64PnCB0lexzpslz4AwtQ/xbz679RB3SuaH6X9
b6iZcf5vqezJxoBcPr46oMdGZx+VgIi2mYl4ysqsqNM7wKpTBAoqA7+Xr/i+Sn+L
yi8rMFfQne/TKVczRNYrV0M2R68xOv35XpqTzBMJHqs9Qp0xo+yQmUOJ4OJo8qGW
RXRJ2mG/gtOa6qKty5G/T5i3A39i424CqV2lKysDQsXaldRpWgSyRzXKochXlQqF
YBScXxUGGr7aAKkTqWzM0wX/s1InXmhrbTrVPyNkCLz4oDDQs8F8wpLLl2D5Dwsf
GKoGMseMtjklc7LW+4wIAJLmu6qTG0BiCz/RWWnuASDiIEVrF9ZohItXtb6xoamk
Kg4D/Ij3SD2u7GsphPN1IvEH7DRxyl8WWm+QVOys9MPQJ1KDH9O1XQRQxzN7c6bi
hPs9tL4Pvptt/5xvd3ncVgFfnSfERqmyGtKrVF49Gtpjht8XJ+pSAgkOKkLq9ewF
5p85qyLVkIdUy+6UtWwQ/TkYTAFofSZWwHdCIBnTdRCKv44SVnlv2UvdbAzPAw1v
vfm0/xVwxz/0qfIBiVBafuL0X1GFrJLV9/T2saHisqKseVbpxX5eyN6ugswYhR7R
K4xd/4ruJZpu0nMg2yfib6BwWsRcQIegBq5cdmOSmnqENSMF1nlUoMnHPMfYIpE8
6OYNpMMw6oQfklyM6eEX2lZPpF0dsCTyFjHGFVt60bPo5hzy5qNFGcN9x3ULlZRm
Tf+Gz4DZMkxqZ15WVi7wJ8H4davQ/7M0dI5D7/kaH1QZcU+2bcG4HTPjjvH8Drn0
BLnhORvtoBPvLPEu6gtSNNpSUh8E1cEGXH12ODlNxyLBbNvpbT2YS3XnVKgrJ3Vu
WNAHZU6v+0Fsv2SKzvTy3JdjyIb7+dde4TE04O9k2wZMiHgX/eO1EsdZc110gSyj
wdpPdmyG36RABB4EzpgF3+Eb07GMG/hZJNY4Gth7rL2OLmHBQlpoNTWBM5vLSzrc
gCDTvMuZ5Pz6YdYTywA1yaParH6BPdc8zuflLESn84wtodia3wxvoQ25LspEHo+f
wnrwaIXlqXKqpF0m1Nv8xLGJ88xq6zU4Tw6MsramXHS89RIdLHlpidJ2G1QEMQvE
Ducv0QV2MuR09SxJAuERZ1GNS5ChL35PookYHwrksRgDVz+SmuKJP/jTa4rfKNOi
25eQtZbAY4gD/PQvzWe9pkIr09ulKUTRLTFDLfxay5S/8Z2iqpGxkmtQL02N1fsk
1NjR/EZ6QKZXHjX+xJOuE9IbW9Cl52G0g4+RRGBG1z5kDLNtXdoarMJBhxOWt3eI
DdVYys1s66b3ps0rNFkcN3PGUHAEUo4oDgdppT8cnaWAj5uuhrc2+ZEckSlBCqOD
yAjfS+PwDrcKAoYu7Xp947jvj8GocGXKgcXtZ2viZE2hdXlNC9XqtkiYpYFl/sbM
ZLvjiTiHRVz+W13lBdIpoBaTVR89FB6yXp4gxYiCH9pAsxwfSrjUyJ7sUP/5WBVa
EYlmdOXTpNEwHsdh6CrGdSOqyqBHzR5nxPHdfYUyEGWMZEhGRw+mp7tfC68+ejVB
sdSgR8UEZZM80WnaSBHT/kMxegMtSG8KrKWJ8Dtmh0R79fAiJ9Ly7jw9wtjZCvVv
l0buTrC/vewMHVne2NR+jeD/7vGcHB4r7ZI9F1TaKmHbC2n5MCTK91avq6Yi2cjb
Zq49riIvvXDvIhehBrmfqrF5lD3KUFR2S3ltm/otpOl5JRKHg/Bd9huZzlHunZW8
reqLuXBzFdR7F9K0aE9XowOk6jJPAr2rBMGpPGgRnB2flvb4sTQepgBkufzk7kNg
Uib+umvzXm1+Am8qMgBpXnsvOXpvx7qGxTjecb6PLo7XJhmJWnNJAR4IUiKG4JIN
pP1KI+d8XRqecIVJjYwYPGGVnNQECec8A28i8PDl7VUbojVi0WrQtb6izD2kAMru
TRpcsBPlfJNGwfKUoTMcoK2ubnJ5lkXHQqcpsm2Ns3JCHWvqeJdugXelMS5KBe1h
4NE+7y7SfsdVfdxIu0xFVy6ZJaMzMmHZWez03LD0I/HHoGghBvli+/od2KzKNxzB
0SLtRmcrt/cf+y9T1xlj7kiSSaQ9OxdUddgpoUCTwxCJTZQV17hT6VCWAkMP039J
73lVom6Bx6eEFF+1ugqppyIfMJ8dnxN7iGZlq0X9h1wTdxuxN9bVoZ92adk4tsz/
cDzy3OvUne4qRFzzP+nSL4f5CyszLonk8QJ/3Q/T7uQhx7DUx07fgTneNNfn/Z3x
rWvMgj+L1T3wex983AeV8NVM7nBjj0chT7Y910vTcXGvPNKfC9ZYQ/7ewsl7WeH9
PJoTIWdG6h8cunhHN4u5bypECKNH6vD4TedtbqebKK8wNYSCUka7jmjDz6kxhg32
RINyDXL5eoeQ1G+3MVsqq2UDB2xw0D++ixdgaQ1J8ga9xwRrz0rmNDeYYEJYmxfg
a0FLsNgJNcX3Y3KzaICZH+coJYdCu1J+xiDmdRVvYqzzi4AuurFlZjMuSpmHV5Nl
dI6PIh5t2sXazpLgJFI14dN4wyDukQj2DYVDtqKWWDTCDJtXpzYfbkN+OJ3KTIaG
xmZbGhZ90gW6ElPfGPo6WtbG2IyXT6uP9dlMMCAUqSdTGFXfAFMa9YVjktWBTN9X
h2/gZcTudH+W4ly+Ob7HdALCKGL1zKoBVbekyE6qlmaD3xDlNYQE2AZQXPQECrAY
SYAFn5Go7R1FQUtLA3qnfND5eP2DTkEcGeOwRiHEBsf/xO/FrNq7LeokiqkIU6VP
b6ehWRwlFNrsWTQ4rZDXNTgyv7oA884axUMzHU8jCy5qlzkd5XrVcl79lzyE0WWg
BesLz9mhol9/UALmpnzZe99f2lVtLyavPcBFDJ2J5NCHsrphU/LXM2n4kPaF+7jj
0ejPAfdryUN+32vnlv/veSqR1+L1QztzY5JyJWeM3AIrvAqpfYqH/yigKAHf3itZ
bVHUwyWhYKnLE55FkjYMTJ0EpCHRFeaDZsXC47mOZnIOs2ge+TcQbQvQ2+tgYR2l
fyPAexRj7fXSJacNZLwH9S23zaKl3hlRKtWe59JUyStcJ8KJTQuImydJLWV1Qgbq
h3gHJxn05XRIBpuAF4tsA227kTuDvcI0u3/EEm+R7WAxVIlzCK5+UF2QPVPKPvss
RN6zJEtrq3xtj70HtnBr1YClTXfk5XRQzed1CaUJParJmza2s6YsdcVAdWtAAWJb
cfn7Ifmy3xVNQwUA3mhe18JwG63L5duTmEbPQD58NXLICU6KeJeX4/iHf9Rp2v0A
wSO0OEmerRhBjs4eo0qehGfUAE9hYXzXdNpcsksTXV3PJ2uiIletUkxZU1LyB8sR
a0cChm201j7PenEwNp8Bzy9Pokp2HGSlizx8E1sPuxLl+cAv66d6dT3bwtI+sO5T
fQJrrTPOscE5YxQYjtLS8RHxl+tKKqv5sIfvgkdfwhrEwGi4/ZQStF2n+YGa30IY
P+3AdrhoUws4OPnPxkwlbP1bdJC0xkFe4NShI1ZOZ/bdnnh/pcNUgJUD6+6xvwH5
bOqItbcHnoMXQ5Q+jThpgfpft59CAKHwWp6IjRblMEdHt/rj+4zfdcLmvV1rvOyJ
qQOlbu9LPA8h3n5TmFqdjKczk+cRUOkzE2+FlpSZVHDQO2LyZtPNM87Mh8JvPELz
P5YMIzmZCe27FmXRb+LPb/Ya3WTU4OSmYkYBhaj1+eqAtpWwloDWVcodEURuq554
dUssP3/HSdgQ6hXN5reyJmmEo4sUPfFiXyg9rvEkUN2jluvK2ccJdS/EBvseMzkt
zCq/91cNG9+DoDGF9Ev8iGhP8606RfFCKpQU72R1yrC8tgjTgPYcqGmSOZW37U92
3cv78qMmSpd/ZqnD6mFZCAZCtK6YHpxDB5ugwNQCnzFAC75KcE03LtbsbSNlwhfq
JgVTFsaNMiC1yJBNZQwdHwnKjTJu5hhoTaZcVqJajlXxpFwOxlPv9p1/ctZoecPr
dduxolKGE3Djp8HrF2jKAY9A/esBeeE1c0F2U9Kj98UqjuOHcd+MYb5QGIgQxarm
Mxjb5NCs47f+kjPA9DuQS9bKRAMO37Jad8ilrRzZqLDlE5vZ1eYe1dOVGLVypJlb
x8Rx0qrOA4MtD3xkaqOtM8CpguN23g9T/5ev1pH3DK5FD63j90Jvbe8M6mvg6WwD
XM5toOpo05Pg5HhFw3NUbr/edsz2rfAT4oz+Wbb+rtn71X98TJoC2B4yHJh9C2qu
8jMYFI7kKDah8m9d7uFFW5W02cvrq+3EuZER7tNerb02YkhJv8ZZXXpVI5kKIZKo
RxH0Hdif4hb+uWr55tfsxtTHGeE00PkrRQ+vFoWoaJB+OKD3LvXCSImlZT6ryMaW
dMa/tvR0d895L8bfQbDgr6Iu6sWqLxQkxWwQcYvUkpF8rtn7HoFMxsldpFRElJQ1
iQ7plsQ/Fnv/Pn0nB3Fyneqw02Rdn5OT7A+hOnQ0fSmQBHIuB47ww7qfDPsm7lQ5
nvkL3JXHGm26TtMJZCzxUWLKfWcsDMxFacIGGT9n00iRkHs9NFrZUpEAo+cnrOEN
kqxzEnmhbMzgQYCvLtSOzM1qIlTUxfB/kNlcHoK+Qqv/PfOVLzCKXSqH1OqnCIjK
8eUwoePDVJ94hwxNTF8RTTLSijDeB6QmMgZ2aFtu1L0R4W647epf/5XZssgqWiA6
eojo2bh6TgR/R1W+Axr3gEcmDzQYSvWSbBnjdxCWx83QmdGTqkexegXdS9HKQo2x
EESPrFu5uUz1prqXqFShSM/Z8m2P8olBZqm2Lv9Bq8t7ebf6Y+pgKyLBjayIvqTO
AfQ2yWpPTLV9BcRmLVcM38A5mpSPFb3ATUISm3hcUJka4rdx22u1kvTp77KQFmFm
fbTDHovDBa2x9o7IbEHUYKAn8XZs/AC6hd85G9vblNSjbnfBc9et6SD8YrTfbDI+
iYbITc5qlpEiskHjPwAts6j8/f4daIvPhyYV066yPh6J6eL26gicNazCq6pCwq1a
+K9fB5ePup3iYcKVugAQXjOlK6WFHeCjWPuFWbNr/fd96WUFnB2681pbwiar9cuk
GBetaBBGaPq/w8u3ZZbxWJl+56CMHllXIjqNhc5YSIdnZbbJkpfWLALpm0WCFUDz
00CDDKjjvJhabVrGMRWo3tCbWzUvhgi/9L3X2gAeB+9H62uq61GjjMxbloZbl6bQ
QiY7b5QwCegk5w7NuRxAe+5Edt98xlZYBSTFkSP6tdQXYu5AawuweJpPGPPusvvV
ujoZpDSbltZrjanlkAeUNVY71A/IM3V9/6jM1vsn/wno1mWxq7fJDZrd2ZwfHBpQ
ccckQXiZVSk7u9Vozr72ihsC4uzUbTV1jAn9mFR+KyNijLLHp52idAGGxS1QOtPX
AbCSJf6Yv1pfszLlPLzW7m2m31EZVBoWddOktDROm2jGmdqhNsuvAEizL/sD6pMq
60wUUjq8mNzw7gDCxCyi0xNAZLpK0cvI9AhEXRKb/ylDLmCp4caRQvKvQnib1XEH
NdRfi1wRMNcd0gyYfCNgeYtHPuKYr69UOKlBF8zXmDbLZocl+iq46sZY4vLllk8G
QTSSXwprP6R11YDUvxcGx/6qfW//dmVGcp+jXK13w/5gPXPx3B1VTeRPFaHb/fg4
wnow6AwFVHNAtFgQ2lCQ8RBHGEhrp5enOKInPb2iDaczgxm0JCPqNKUJyQYWYUSq
IvDT7tGc/cyLVITQ/Mu8gF1ztqZgEjNAFQGpSi1aJrCSLuKM7eUmTYy1bYJVtyDe
tFNrkQDviJP/cCsuQZJnIl0wy1xX/apE1T+xjbLHSvdhhRty7LQLAYR/I5MskKSS
sf+TWKdAYzwkdvR0NlO9ksRzU/J5tj1iMSGiSGVefUavFO/R6DkZHEHkPzVLIXfn
+FxUJCtOkOz9w1MrJyUlEfaZZKhN5m0/7qpTrF8xpgx3z6WZa7Y5N3f2kzw2ie8G
UdH+AHIL02iNrMWv8LqZ8wXtmiCCBI9XM6yLv+zdYihil/P2sMpPDSLjLDA0x5Gj
jgZRDY8ZAJtjMMZxvbBSScfgRwjDV1WsxDUVAkLBMcl5oydnEXDgalDKUHG9ofp9
icwEt/0cnxMQzdg1sFJop7uiaf+rD+IjDiqp1JVwMsDorrk0nukqc9RE18wSQwfN
hmltlEiRqPC+0glbFjxamj+8ul1FY9Lb4dQ9VHJkN0rAvrrrNb/NxMccP3AsmouL
qN3QKG0y0L+ZS18dXsyXkOJrkq7guJ3fHXKuUcp8+xlmb238D4YB7JLSrD2sliLm
lnJinoFRd3VSzE/i40EphWWXi+xqLDRk9UV/L4rJFXpBZmt+LpuEseRd6L2msoIA
/mbb4oZDKUGEd4pvRqg074vYax1+Cp84awuEt9mmEDYSn/7nO+WOZM332yXRpW+A
alo/ch8AniqtN16ayvAiUPTS64PTj17Q9fJOE++npb3t572tqy8X7m7GJp07BdpA
ylYBPoS/Keq7cunWoe/KMzEqJC0t7QnnvXns2LVk1KRlD2G7c1OxiAnia7cr02Oo
pZ78ZOaexaU++zTsgOYQHzTnoqweShvEv3bbvcbCDDwaxDEYFG9F+5385Bqi2Xdo
w1QMGbrnzJMGo/YfHADt5sBR44ssYW9pz3XMcyCXEHlL4I9DeOIvE4DjGCJ2/RUw
FmgNautK2V78pD3VHM4dYbEBvm8Tc/sDZwWGO4Drr4YLc+n/LcEZdfjbUyAz/LCN
35cIepDPMKjh0VU+0Q4pW7lC2E1Hp5Fp0uVoitdej4CC6sj7jfHsEDhAz+XhdLnV
Oj4pHh+4AO068OFRqtKl0ZxgvwQvyNYAM3OOUvJr0oldJrqoa1rOtVxyibmZBFF/
kfZaeFeD7v/9o4P/XArJmC6Mp3dq+JAqASTowg7ffTLKllP8vh97etQIKwsg8V/y
TakVplpDHvpqBTgeQuvSaPCCRHl+CRfdiBK6Q7eIuIW5iEkwrun72An5n54WZSVJ
APrZMn+jN1TV7SZGcCyCi21FXN22kCB/f7vcFWB3srUPbygfhS6Tw0bY2WB/HhP/
s3zc2ZgsqLOMCUkJtABC7nNcfeSSzCPqou7/yBlk9R+aUWgtQCGX5iCGf2lYT0LP
r7ZbM34VnfiWpmd6I6u+QiP8VrF8qkS/B9oF0uKDQF/2bWQxtqkhSej2D00URg9k
fhmgEzhJIHzDDC2eFFBxM0L4zl/WaDnCQDTBxyxeDapMjacqY8/MutdDfQP0BSNl
qnz3W+iXL1RHo5DsFbz14pZK45PfcxowgO7ASKoIc5pqfveIqUEQIkPOjT/5Lz2k
CmnjI/Ur3FFQQkKoRyzVsNZRcYGLDi3eXXRGqIWXYMo9SO0pj6rIILw5H/4a9nzD
p8ioOGeDono7alQFN7zZxnBs7HrYCIO1tGprwAUUtuJvy3PxfBsiWacvTa5G5VKx
4Tll80WEq12gi/rHwJR71OI5O8aZrWH987OTn8MMv9wT3lqnrR7yDjJyM20HQUMT
SiYUBKLlLAcp23pMVhwDCC4g0odxQPeKdvYRzA0rmmCoNV/4a74L2TcCcbO5YRas
Wy9ZexlEpyQcw6EdhSJnAN03pevq2acFCcRecXeHzaOL7McMpcpdL1iGODq6aD/R
35HeAai1P1xGKwkuzX79yohAC0zQ/wPktl+ss/bBSWVDyAPikWLMtw1H5AqktlYu
xhBXYWrFn2pXTqCgRyTqXvIVNqkOej5sNXl6c+WisGVPbS41/Fff/qYcv8RBvgqS
/Aljrm25zUeWhWoaf4H/H3teeqTzd6lIhtMCw3kmqBvyp2Ej3dDx86kkMT9lOnx3
5/OQJ/ptCySSQhuX0IpahToaSKzsRB6YqvT+1I1w4XZ+74XfSa+YaBlF9Ac3fG0x
l9P4UNnAAmrl+rFDbvD+VlP47yOb/M5hsJoK8HirIJA+ZmjQfn94pT68K4q19w7O
u9XuA59OIYSutF/v+Rg1roYVmf6rUOa9WrCgJ/X3lhFjFFHFVdUwZbQfwg92ixhi
lKvKFl0TnIKmwMOEeAuU2jMTIXnTnLjRUBu5O1LNzN3S/aX3SrqjrxpBUuHsJ75/
d9Dge3R9GX1k7cC1owpQRz6gaOsaRFgd3cmoXdMeNcHCRwNfluF0ZtYSZfHQPJFn
MqQcEo2xhQzR3+LIOC/mwLBLoZFdjIYnrrI2IBlSGOjeEXgv7HWICDaxUgbATtHO
bYxP/+8JvZbzIShVbyyhrWV52mmotaPtJox3yPrE3K3k43AbExKj8AWPA2CgjN3u
h2+pMZvtaVFjt3F/BHSz0PobDpNDkYh/UGcTtxmMMViGEOfZwTwqnz0Cvwoykt3A
z5MW78dg+ae9TUVSAUHDhaWFX3VErMHGYjAX4EJm8Msu/hs+Y4B0U+0b3d5TbkE1
58PO4Esf4JWzv5fqanTifOGG4fRfBGa3YMrKR6Bidv3Gmym8SCA+Zq/KgzyLe3cL
NnKX9QWPJSxCsvs4kcTrKKoUmreL+LAPpBQWLUBiYborCPb81EHpUZmO5HCC+Bzm
L84VT1qbqcX8F/PmJWPQhZhCKTFe7usWvpCtHgP/BDy/Gi1PIVfRcZpuXcOhky0r
+s5H3sEFTRVy7jfgA/sODKgdsVUCk9Rnq3VEz6uM8dW01yn4aLQZ0fmnh1JTT2vw
S+l6uRoq3NHqHzo35c1lcbKLSX9UDVTgjr2Ivxg2UaVql63E2Y6JQD1cuccqr6WB
UsYWGkhlbDi2BsIDpmJVmjE13dUQNiF2FSBkVRhr9qp5DM8XGpHd3wO0kGYLutyF
j42xwMuY+viL0WMsWwKYaMbGoU1YPxYJjYo2BzolkPgBus1tUkV1z+wyCPHMG4yf
WHUucD5Wv8WrcVlp3y5L0jGlG0WvAh7djYXJdzDCXeTcZUs/AtmOca8qWBSNQiQB
YFpERGZTsXb3jzWd9DZJbOJ/Tk2Rf6W1tPkwF/Ow/O9QChDBwCG9bWKZC632m+/I
i02HHBbgL8gzUfvlRsg9zDGR4fjB9sagCCiw0SrP5h49e7MKrqf8/qhjxnUeVBp1
y05scQ473m4kqagGRJMsdWgADhSh3IVD+HMUJCn0TctN/N+MYWUTukRZ9FLhk3cI
142HbwwpBZEZrLFGjUkZaXh6p0bnB6w/3l7cxrNw35yRxYOo4GDa/XB1vP5ZFiwn
MsZq9ayguanmMrYXWla1r60WAHIwaIO8P74ZunJE/2OMtKluvlackc9Rwt3BTZhc
zEawQi4ft7ffyCUlmhamsg4mpSFcX97ggDwoSapMwvsuzZ0tk3R+v8lXXwwTYowY
5QtrBELfya7fXSrUjMQqxFjtFZoyxQTqWR9ECjveIjpQFCGu10zaxu0wz0gnUmUx
KBdog2K0ldt+FYE8pfdZ7XlEXJmyHTpOn9k0ba3txL5z83fqVr4cLUcbdIJMq3YJ
tJpdy4BG776dV4Knk8iBeGNQBtCEy5R2DR8uuQKMULq+qx2Qi+6q759ER8I2HYkd
kyyuRaIDL6/+Yg7EpzN5PFuUm/Pnzc7PQiniBsUm2znywC9iNRdG4YoRz1ONv03y
RbndyYYkeyB0l7QdIdWYujKZoczseleM3OBQSCKG5neRXLZvZkRYIl7knoJ8YIQd
I/0yVZZkuTISnWAqjY/wlMRvBkQA2C8Z5fWheEDg8m/FkBiv0zINKtuqDYH9bvUr
nBdjJcRZgSW7sKxqG83YvQ8vrF0yPfZ/yOJVEKLtBdfYgKayE8NG57eX4t2biyt7
L/ijMfFoJtICyQZZCG3DmfCuUNISX+5Sanf4zrlw/hSRZoZj6yXJ2Xqkr7Kh7olP
zYIEtpJjEr5FbvJPSxXyVFJpWR9qtzI+WuJmT8UF7k6ZH0iVVIBJP79pOL+4Wsih
mpiqfAYZSnUyYL+lB5yoI2xDB+YtZmwSaMJOTcOze+wsIzOPdc4KnPU0ZOiz5Pyn
iynhvWN93XwoAKQ/XkTCPT91Gx5db9iKnskUIXrkV2NqmDlRFUg6IHWj9nQBNO+D
LuTHttjed1RM9nrhtzomj6xEF1/1ee/5riUk67K5o+M4yFslaeSQp1iBojNc7yUS
vrJNnQQRrQqMq49UXzMgY0QWf//W2uw8NRnhv6Hi7apYR6H8IUcscIqKXQeP7yBI
GtccfksTaYsSOFnJULW9CDKj7tSO7t6KLmixFaAfVTtld9aUSoOjWcsxtbC1OipH
UCPHhu+ICSyNHmj0IEsb5+fNo/gwLyfIMoQBOY19WJh9PuyePI+aSoqsLjELS8u4
6PWK4h49UkTdU3uZ7KTe0pJdyIGxGHpxiCiCxsdxi9iLT5Yiamp+CTJ8L1ThFQSQ
yWpW1S5COIEF3+C2UopACXdj7vPIQdrnJQVKhK3jLG+bS5MoJudyJ3B+oe8MMnJI
G4OctCIMOf4N9+6Kzzl3JBfwEdFJSip5GurBanjpjoWMaXZVCEc7Ti8G5KaMFEnG
HNuxLSqfUOraKLw/MtHSKiWOjIpveOq6ij1/QFb4uH+TB68j5c7/GEuu4eNI2sGF
o4EGWroUtesGDZkF52NUO+nPnCLCD4Wg+ZschG9MD7ZcZu7ZBTVryZU+RZsezrGw
+675kEvCQnMjaRErIefcZ8/jsh4BQiGyudRkML/4k5IhMqZes94zz1XQedJ2Rb4r
kU1qptmDJ5VbJF3HN79lIGxS4vjXowkhlQ8MeY7dyjL/MWkQWhTvA/epMeGyT8WW
lpeizIKwOkoe11aBEeSIjYsPDSnS0XjIHvyffcQsJiNwRqYFE+rawTtc/stINC98
jogeRRScj5nnmR/QhOrY1tu69+XQWwrDbWRAFvMHtqcAtWBICndTVMkBDxsiVrsj
YTQ/9hjQ3l4y+tkeqyCK9SIkTEfAxCDSjC+KWnchvEBBN80H3MywR3cANHcir3gf
zpq6YNBIJ1PstlEjlPnwTNEjOnYY0zwVfNb6oNUnkqN8+z2gu8B3ONTegOHWBgM3
fMk/PURGZZTXfJlXynSYE1ibaN2KueyZ6xyJZjzPdmiWBIoQXYsvQ76xzhesy5WQ
NQUpHL/8Ete743jBDDZDRBpX0gSIs27Fm/v9CBGcDR36Ho47IVWDhh8Q+LXnAAfZ
DEiQhDp/MbWBbxwtalY3jgPW4+rKXC1dZe/d4MDEkC8896dnYeVbrzZInxKJol89
7smQ6rRQj5gwF7eX4/iAY+icv+c3e9TzQ384QwyPZlra6sww76xzDncp/M++K1YX
w3ldbW7eRV1y8NrQ75b+jHqgrYE/H1lzjyXRH4BNLwUjTLP+g9cOanEd9FoF0KUw
e7VLCN684Bf7KZMAlkJ0cmka3qAeidpAv3SCRzkCpAAOV/Y5xMVI325co8Vduw5l
mgJbqTRGWqlV39eEpHZQM5mbIMaXkIK7uZKoEXPKX1MzJiQrvx74XJ6K/RWor3le
d343NvOoAF/OAgOkH6KpVOGgoNh2ef2D6eo92q6FqGhFzuIekG69Ep7NAnatjjj/
YfnppXxA145wwvLsl7hKVXo48b8+zROc+QD5ULxNooe+6bz0Jv/B7iAlZYNjkHvi
ETTY/5Np2M+bxkTx1KyfPqttH8Qb/DJ+rL4YOcThq01r+P2Zl+fvQ+HdolQthozj
ZrqVsqd+VqzhQGcn2HG0ecEOkWqMpQp8/Jn1G8O8DwlU4J3oOd7o+y0FjInMlrsd
+FEJR3dg6e2OrH5fWzvGURNPEUJtHa9KN/aSkaDNJi998Nadm0ciuby2V8vZzIRd
rGDXRVWB1K9jnZpmmrNoZzOjS7lkFV365IIkaycund0MshQMszt6cf8881cq53ZM
Bk1g1EsSZ+C5YFUtMJMBfRsV20ZQC7sdbcpioFF4YPoosHVHnxWcydtZn+IEBr//
9ntYK2HaVDphYHO03tMGcRAYyIk3lsPl3oPgT2xacm9kwww7ldTv9SqX4TXHVqnb
0n5Ibp18phS5gBnuB/mS0FbQxY901RyvtwRfz9jjGjMyl16y2fU5cp2jbdmlO3eA
5BhbN9OONkYUsG12J9BsiunjGZyQs9JwpIthbpawjK2jbArGSHBoJfmvGR74uHEI
DHdg8jfhsTxYyzfOFDWnstmVeW2qWRprO4QDsUpRv3GKx6edSwkSGUn2wQMoZB1j
YB9DYpUAJ0RMVwYkGrwhPtXBGCU2jkt6B/rzJM8R48m8yf8/3RHdU30jQIv1QbN9
9wfpnnoThlHOxu3/LQ+w3axO/T2qDFEhX0h8nagUYU81HgdQ1hif/xGjnVgkNK1z
FCZ97+2IQe0Nb6V4/JjsQMTknotHXl5RGvOQHJdT/JAxkuyu7j+NYYu4RwjtKVuM
jptcfzHgmXW/jtjwUqxINNXrb+Je3NyNVa/0Yp4mLwaIat6AfVAAA5USMH4nASrv
Z4WvQlyhwi+2g+Uds3N8SyhyH4sgof5nR+5e/V3/K4+55oHhijXNonF9tsXKB19k
EhDnX1as9ipzSBbW6rIoZvaUWlrC+yKsZKvSA0EFJuPsYpdX8WuQwCMYwncKg6wA
CHjDQ4tzw1lsyCULfMEuGptAQ1prunMz72HoAwKarPXlhv3BBvdfOI/dsDt2S1rp
9pUSZxRToeMJvhSkMG2PRQL2wZwC6tThJNbLMAqtF3YxIkADFTjEoH3OMOHWKpjg
YQprPyoEbQcEdjKzxqM4o2sJf3e+/sXa8T6AqvM1Ufr23endjMSZTT76i7YWlYku
vrTkl//K8OB2StRNEy4lzyuwPDgjwfr1Aff5SiEAZfniBmqJUtUmD9jwhx3rzW2P
AqzTzjXWIFdRE/Q3z2i+63iOSMjbadnYBRAQe44S+V8EqHw1Aa1DkAEY4POCRPIK
gnPzRhfN9MOCNYQxRY/5TqVXTkyKB8ZGv0gxMFjQhUpgHHzMgCb0PZG51qZ1gp3W
W4IUC0rC+HAT3RLN9ynUN/lfW5aGLcl+y+6k6DpggZhTvCle5hDdvH4zjwtmg0MC
1JdzqZ69eu8SxPO2jdFGUQvZfhwuZbpHAkkvoNK0gA1i9Re5S2f3qypE6WksyE+s
cmiBEvWZ3rqon/q6BRhKmDERNidsknYLZJjCl0KPFWHpPImdCyk6NEsH9dahuJap
eWWyp0F/7WypeYoSpfNMse0KCiqoXaP5PbEg4QhHAf6YMPKMAaQ10f9/oAgeB/u+
usUxVXRrld3694HWC7P4gDM0Erj3AviM0hkJDYyaLEbxHWjEtLDMZWpxhY6p1FwA
4VP1tS8H5x+xGYpj2UuLwTSDwRpYuU/4AosvFJmxhPQuWHH7AzAu681fX8yjnWNr
ei8nonDeo8G6hfGvMJIsGRntYnXtfumTBCVBH9xAGriva7GbQz6gpgY+hFxPlyi8
iSP7ESWdSzM2pWslyyoPZ9BEFU/GDCXFFMWQXe2cRhi1/PkmfzggCcnwEUkmcLyU
iXJL5OAmBlMpP/H2uGsCgXyCU3ukr7yOoer178niZdOJi+pYCHc+XNe1V45e+oy3
+WFV17HsFcaJw1lF5kLY+0Cdw+g+5RLvg14cu3XgfYjLJlcv+v+rCV6pXJw3d/mR
JtfzI6siHyPzYQzWUlNyE4yzPW+VTP2eI5WkemgwIp1z3Zb60hhMTDxfivAI2HZW
9zggWicy+6AMCKJmTmF+Mng/S1osM93tmshIjc3N2uKMHyefYTTFmUZ5nXN7KyMq
g+7wsszOpiYUmDfK/4qJNopNUygEAxZsAP0i2L9XeQPu/eM8e70TZDGsIwbOVyaP
05DU3ucIyVt2GSyIGXL/ssrsMbxDV7aRx5an0q1hiBDvmX6Kvtbk5w/DPfrARmTo
je8BtX36DzrvRWjCBNytXveXYVCadjz8BBUBVV3Lv03FgQUWg7R9l8Amk4+BVl7W
ABeyUtHTPHdjPUdt1cLCmmAfpX74TGjtEuwHR1leDKCT0oU1TjtOPncTUzzCWaYf
xqNoMQ28cimRMFRL98jsgz2gYrBQwWQ7rhRxFhz8das1OVxsOae78cBzbr5dEp/c
nUlIu3yqDT/T+CLZLENU/zJcH7eMHpbcctvFVs2ZXkswMzRE0Wq5QyjT9Ah1nA5P
Qol8V+8Zetyyf2CvbfAXZVHUzn//GphEAJlN/VyQ6RkfJhJ+Vand+6/gH2W5IPTW
0BbPnmHzFXZelHH+vTDOO84xaf5fPdG1RnoO30RIjhE+ZlcKqD5o9Q4DvJoxmvIX
arkovEX7LjLfkV9jmE4mNzEMWIqc0vsNBlePlRrGyECVo/YamaoLeInzhPF8inBt
HhOJ5sAMPvMmPONzBdwBq2U1kHaW4Mg0kPHdUw8BZohNacbxZJKhAMANm/hMpMLo
IkdX6WB0dw3iS6iLGs2uMER+3og6w2g2T/rGjFzUdyQbQZyQdStIpfEfOeZ3yz7x
QQD3xlAkF6E1H2WZQxPshsnOpuzCMOExJ4cgIRJolth1a6OcQgU/RYlCd06a+UG9
uPWIl9cB4yRBeJYAD3XgeIJa0jhlxI9i2jil+NaracFkiU0I9HF266X7RbM2uPVb
dzv3YySQ4V8K4I+S5QLouvE71G3Sz+4dA5gyPV2a9si4m7gb0K02vPDUMchhk4zt
N5YoN5cP9uwg3sDnxBKGtVWZY2NjP3+IP2qX6nBcbNSDWtdb6jiNlX1Rf0Tcq+iJ
mH1eTOO+9735c5riU2T8IttUgKmSYk7SY1010Sa/nE1QL1WvnHdRGQ54e3gvHbIv
2IAY0oarS5Oj7pRlARkKB6DgFUCo0w8Qe4rUt6fB4hn19xSFXdRC6L1Sk+Z3GtZ3
/ljp4Jm6Xcwmeb+LfSAm6EIJvKEUct3r2inBaH36qfueAf7hZMx4aw4L7w8Vo02n
S20kMbdj7BexBhz7K/KkMa5infrOPnNJt4FVYf/G+46bNzFY6fEQQqDYLd9lKm9f
T3eVbL28L5E7F6MPmUm5TGlBdah0VdXGA+u2jNz+P2D9XBsQWWMDeG8t5Acqz0td
N6J98yOE2EfUUo/mUAkeJ905azRQcAptSNlWbJKitHujeuIYM9FnGzheIdjt/TBF
3rzWWdos9Uzl/XHIWFnTgjGQfGXdEbqdvR+wVq0xDovn++BWuQIC6agaoGNzzCM8
5yD8IFyfYe/w0D9Dqw51PeCba/dmx/qhL9dTVK4P9CWWuVCNB6E+iRSqpaaSpbfe
PWbxo/Dget8Ysj5kZzDW5hvNGOky7p6knp41jPbD9i7gt9fd1xSrvZzRHWmHh2yY
R26ob1o4sMf2PMg2VUdNH4t8ZxNMucSe878rki6+YMGmiF6OKqhergimyc+S1joc
Dw4JX2fyTk3knitdpPHU2hwOz5vok00YQHL2Ga4XN6kj5BqVRLdrZO3qmgsr0cLQ
9QR7/075WlZXPsm8qHPfwXKRISFHIJJafVyGNYNVJt6KjImScxIVi97rO7A0MDvV
ahB1taxDrGyzNUkO06TrWLvgo9X6/KVEUscbpUpD4jR/2jfd6op9PPlwhW+KoM7P
y34qYuN72G0THrZX+p6bmZX35/PSxJPayEDibJU10xeWdDCRmTdVzhCXFbVPIvlA
y0HojfSEcmiF030FtGJFvBMcIOqKzXUVVkDGOA3+8rFC1rykIeQRZBqp6Rw2ToQJ
B2QGcpiEQJATNXg23u2lE/U1bEm1aBQvKPn21Q14ImJiAZG3rxHQhmRmqvaZCm1x
n9+YRQ2MNNVDeRDJnZfoj7wkEE2jIfKuRqxcCzXOBUq/H7gP44D4i+n0QGUQmv36
Es6J9sEtjU1Skxw3mTh6zme50BgRz2LAaFVD8vEzF2la+aOF59ggU3NezyJaU8KR
yGTITScBFGvDpaTUSdkiqA98xeSAuDSa/nHkyL38QXmbAoGEXnUUdvqd/3P0sypd
i8tLn+2TCqYnO/msVAp5e3rPDbPUc5fCcQ6HjmJkRrY5xn9DAlStpYB2eEDVA8i5
YXFvlXdtPkus/v+tAb76qgKqENPDQtx36jLzuU08Q0HIs4nrbWQKFUfj5Ib7351e
/HGoEEREDvZPZ0y4Wu8DmMXr5kdnWANYiUOhCzXshK+bdcq+N9N++G9zVE5gCqnc
bU+kcCiA04SD8yqMovV4V7aAIouK1z7Pqr+ZV1QrLDflb2VPPjRrZWShllx66PnB
+W2sBL/G00qHVXSgVETQSqsmher0YvWq6Ejo0vyLEb00IpY0Mw5PVZVRQLlsAOin
YBlhl1Qq3dLKQ8L7sTh8zYoxPIDVxBCVVjak/ognl9ZRrJA4lI8OCoDCksVJX+Hf
RJXURWDROCMR+rftVjAbW+h5H6qjrMJuMIJUCgZ0hDcL8eCiaoPTEJoFW9awAPoo
rCqErogLhQNDE40d0nfXj3Am4sLPxkMD4nxehVAsAeTlJQEv/OuleBNnvdXKKLrM
6IPNZwSuMXYOPmerJk0tlELnuJbZSGH3UxBLk//Jrm8OjD0kNzf/9hPYhhqqNqnz
qaruZ9qhil20ahutiQ+sfsULDUrOpNO2kLtEVoZMh1Iu8/igoZUa4fzcaa98lHWz
a6XzNupkcm1+38AH4moJ4+qGCEdaintJGYSdeBPjKQKeZqY3E22mUkYs9lJmE/xR
wmL8I6UVOeQhMzcz3yvwx7LxoCL8JbcWOlibu5oGXlPu3u048XoUVwjxjFzL7y3A
tqR9o0go9s+twUIZ6yGzFVwHCgjsCJ6CjcaRmIzx4wEsSRsP1qStMOr++hwq9me5
AD59KHcRwD61fQ+s2/1denEDpJSgRgDirCVcntMbsGJrQ0c3jNJxn+NqLz1fm0ja
ynQSntdaPYBykdnCKjp+HmbRRZaUVH+jSSJBB7+KKs4sIjN27/L8knh3T6laKsAI
rcWPB0G7BSdgZmNZL/iGEbIN8Q3AwTSbqPKPSDs+15F7EHLvhOb8ZTnLZS57ztuD
hSbeWU8dAHrtjqp4EYwdXXczGdqG8bp0PBLjuyKbZ7K7mMWdzJAWKqK3V/Q/Ovu9
zbSp1QAveQyM34kVVzxYp81zysHD2ac9O0yJ3mHOe2BcsdNwGNdWVuwT7XAUCzmR
pfj91+tNSqZe41Dpp9RJWIlNMRspMrd0tzXbenvmnSS9Ol3W0glo/1d4V64jrgNV
NTWyxJlRwJ+2x1KGk7DyUwlt1/JTnKApNjOAq1yUKtzc6HhudRSlM67Ct5ia3jhi
+OAJY44do0uc3CrAL0YizKQwJuUbaWwJ+LcHlutuzCWDa00uwdqDRcsW8mwTrWie
1BZktDH1q3WWnc3vSTTi9WW7jtXGrO8d65ZMXO3dFJWslUottpMfH8mXNIjlsvCS
RKbmm5FsM10W0KTEaIIptrpP20daOHZwmF/9PVzux0WoqFuM51J/7wPKg0nBghGM
c2sHbHJc6kdfQq06Y6YBiwOSJxJDT2z37KxIyFZpnh2jjHdZnofKm3BViDIOJJIR
yWjshyQvSZFQKqprhvHS9eG4Dc0rr/f5fgnLN1NF7LQN+3nNAYg1DV1/oR040HNT
t3who4PFUGRU9l4krAf07T28no9J97+nz0I4rq7eYnW9aVDRYXDqduNXyBz0Nbz7
5g/mPAD2quFRuqXmmGhjk/dYxpSsjNVlYWdrvfFisGkwqqV9YCnWc/QxAnBRWfEI
S5+dQmleOof8zQ4fZTkADXUxgCWtLjDA1irARIA7uQhWRPDETnALd2Re6paR/5Cz
LbMU1IjjCAgeSRbeSjYxchTxccvc04zkxlmK2OILoG5DNVNy8AUkfSZKGnU+QZDG
QXA7OhNrQAfFEE+O1khlXVN0W3Oirx2RG8w5KyqZaNwpHGClq0kG3VXt0vu84wNe
0+7XV268qhHqQK88RmeP3uh8U4W7FBUPeWXVh9F5WiFyLaO1XTcpfrFkqjin4kNE
kGJRj0uTWfuxGs1RzL6Zd0Q+guHBn4+0nEvROPvMPBh4wAUlvyLYfi/GMGzJjiVv
uYI8mgsTae866xto9za1d7AKSUeTFJtY8ScpL93vDHBJZXzRX2OKBNH3XBDZftx+
q291ApIfFxM5s74jssz8PdKjYthF6VpaJB6i8YRxJUzchoR+VsROmiWBV7eQ/R1O
i4sHP0xDw3jtg7HOtgZRYLnrLOu/EY3NNQgs/bn9M3wWXbhCJZhmORc5gRP4C8Cu
ycuX5Hl8vIoLOyMDo4op4tVQ/CP2pDP87ZMNgFTeFPCMZhBtJ0rq++r9HMsMis35
1Fpn829pp/bbMCt9gT0NRvLHxq9prttNEA7LRBeAeZwenOMxHOMFhYyLBkK9ZMMc
7bkIKMYvIzUTrayLfMXGzejL8VyaLL1MUo0M59MzVTR0E5Ob7Ep5ob4mGYSChOLL
8d5xQ7nvTfs8MnJlfgQkLfzzZX0iXpAuWnlzUJk85Anh5ZpDELLynWNK9fyBjG7W
W9mcd+Ar6MvsUj4JTUqsB4ie6q69zEOfvWkna6FfhB0bFY2au7kG5PyGRWoEUutj
TGZcSGIYTfvjnlPa8W48VIArr3Z2fgXLktOq0egkYIWSiklpOlfiz2Ywkco65mSd
fHW/GlQNqIBoeyi/ruRXm4RnKfvSDcKHabRE3+bEy8tCsooHhC6IsoWAbedbsqtZ
oLtLdZ1HutG/g9P1BXZVog==
`protect END_PROTECTED
