`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opnx/HUaP71gl4gW4O8onu7tlPTZQkRdvXtS+u1AKSrrIRrfgZPDZULFahdUfuln
qPCxWB/u62CJPFDMzluSM4cNtpXKRtrxjgb/tY89BVvKU3nOiIYqTdPFAh58kBJp
bj6HQRPyd2J+JFb40tE/InQg4v92Yiv24GYLIEzGTop64K9Tp29ytE7gRUvf0fxK
xNUgPWgJO2BaxAKGpnVAGqIc1jy9WViA//mJ/O507FISarzxecU1S434IWK86Qhm
BPrHikPHTrLqd6Wxq1YVXZbUPwu22l0Mam4+fZDl/BvPxqNSRm3crWL/E5dTd9DC
oQ6u6ibmMGKShV+0u+5iSHUtMeVZ9uaV28BDu40AhsjUF4EEFcvCUrYKsyVVMVdW
LbHukYT4hzXIMchBm9qEKVuSmwtXL/VQorKisFZ1eXoqI4rO39UEfZmWwJBZ0FZr
lYOiTkukkR8F5HfkL32wuzR8/9kVrncdOSUNQsYFF+a0Uw+l990Kw2vSs8/ZnN22
QMD0sfoGEEwxiufxRLjV+4XLnIdVXG9P/3V8N4efXVo0Ri38Y56spCgeldgWH5CT
6gLKy5aA4kEGeEKxtTIKKmTG4Sy11xNVHHtg+LpzMNUvT2hbi17RY1FFdXR7gVVv
fmviODFa3tH1/nm0+wN9kbytExi3jPRGJ65E7S+jZJno9tnMSsG2WatlGUly1IjN
UHiVbTteZUnyVlSzqZJpWWdavGhzauSIoYC+9X8cIk8dxtINd6l6kK62bF03wRg8
K9PVE3NuLCk1p4rs/QAnosl2IAv/3qozwpZFRXtczRUkHUBW2tWduoGIXEXVobd+
a/rWFB/abH1Rt45WVb8SOJgeWcdWscgP9UhAZNfRRhUpjrt030hD9tGCv5dxrbpO
rodw9lsyweW89+ysj+17TRFYVwb9Wwcq8pycIbuuOtp6MPy4K0h71pA3t/rh85Dc
WaIoO1VmVomFFTIV+Hfp5mQIQCtj4j8Oyw+1PkEl87DovDmLIe0O4+7i6tWYLCBq
f/7LopLaLrcJbo8P9JwpNwt20DPgU3P5GKVmiKG6B6KQinPTRrlo1SlA3Smr8lvH
2EU0KbcwtqMyCySJHl5Qw9NYcyMnGSVDMbCLJSr5lBNVWQa5RtbI9gXP6KLRPEEO
Ef/5OyJTRaEYV5cgPGXSYQW8epfT/SbjDeyUAGSOJqB2tt7Es+4NkVPtgyoc4fg0
`protect END_PROTECTED
