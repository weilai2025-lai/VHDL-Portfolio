`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/8IF7hoPMFavFyOZ67UKzETs+sTr0ZZcrnVbfildUn5SzQIcReLbKCSYwyKONDj
AACVl5kVQ8cquG2CwGO8TbaOHXVAYa0bIa5wcbCCCz8ibBHSRcnXDyTr0yhZ5Jh0
gKh7hPytN12u0h8lHkaBQ8qB2Yw6iH/daqqUKssr3u+nlr8PpzU/5EfM8oKoH85W
o6HT/VqHzngACOuG21cyvJQH5wD3ziaH4pTuqTRni3FkOoF+THvkAf+IH4XyxrIT
5lk1f4FTCQ9OnnZXjgSEY7OLRVlDNO/sp1xmpbNxF1Dx2L4WZwFjHrA3GzaOCnOA
7HRsTsaaJjmXWayxE7dWQjqasDyg6m0iD4TVlTpcs3wEr3tjIZIk6/X7LY8jy010
YrIjO44ktvT7jBg13WIlOH6AhMZ6r5me98pYuyVDfvyXKCuZrHuw8AN/8s63kq1K
nnBYiE7MFSBpGb+KIIG907nXiSuQpdltiHR/Cojq+QMexBsTpNT2FwEzPRrtHDVa
K4IwrBmZKu4zFO5bs1eq1k+MEi/hyqIGBrqkIJGbMqknmPeY2aEfp6/NaP/Gqo7i
2xUEVtIeRWp8aYAWzEkM4cyz7JI0wl2PFEUUhpYdU2LS6jwZ47cKJZpKZwmtaiwM
kdffKE7Gzl8k/A8PV248Z44TI0jBU6x0SJ2L6xOnX2CnJn01auROY9nB8XLx/X9m
QAoIIg0rGJw71PNu5iSdCVYqi199R+L621HP96lpBGibIsFZhcwrr6xbjYMniURc
Jf/bBGXMw8VZ4kKsNoi+h2SO1ic56ucJIX9XQCI4n5ENu6V5AFZ5uDNNa3BKri1+
X33IRHa1AmsUdN+T3RKw+MuvfHFU3Lz/32hZAVm2nJ6EweCoGr475I1c+/c/X4y4
jdDa1voKSsBcWVtiK5a6qN0/Mu8LwdcT/2tBIqRmB6QaiBCYYO8NMidzDvsbnfpm
6BUKbzm8+/Zm5pgobZikKuC/qAxkRkE5oM/kY0JUS/Z892WnSxnR+j4C+fmKfSIr
xrUzThICnA5NujrrYDIBc0BsuWhvgVkF7w0miYwdbHxQ+dMfdG9QXyGEkjgw5Rp4
JOCDnKvR51mMjAB1VELmJA68Q/RBZrqboYO1hahM3ynGgHuu4PYH+0O0K0ad87zF
OHC9EK2ej637Ivhy+ZDy8NtHCiGnJXahU+Q/337lt9jdEO+eXAmadH9QnRS+/rFm
bvx4CZlBgkRG38yPD89FQHn+tzjzo9oG0MsD0ondRuiFjD6EFnPom7btHmo8NDvi
e2hZHkgvunvuo/2UqBkLlf1gNDQCA6GL7TnCBNVkf7HVfshlL0oLesmwt3dHU7zM
6o1ECPgSZbzeTDx2qjCBUNbxbX3dVa/uRsl2P7pXhPWiriuAYQh9cQr+xfMPthOC
Aeri0Ibj2f8hCcNO/iQ9RIFaGyN0SZzGkRFLzDINNCem9wEZwg5Mu+kq1MOK1cT8
enKNKdjRdkPkA0rcLwsga6+6F4SIMa9osRQFeYLNxRDxPp+rzIpOnc/3WqBDMI9H
kK50E4G1IXsuYpcTrEtI6FNU1sw5xMegEHmjdFeoKu5cehAZRLwQzqVgaEqyfkSE
N4TY+xg9JYecGp7Yrq5TQbQglRV3x389m07rwoxvotkNSo96Akdiy4vy7Vhzl6Xu
53Iw9wTGYRDppKkea8UzrLkUmbNvuCRED/Xn+9MnJUHd4bnbRO0bQWyRqgojPvMu
UPTPNr/n6nS3k4GQqg9xKpLCVydchdGD8GwB7uWtymXsIFJ/XdKyoJPA+BoSRY/v
dYNhpczgaOH/eVKCRYqkEPocMtS8Cc1XnCu1bB+5l3dSsIuN6p6YW6p/yG+cz7kr
aT04LVltpkPcRJ/LHrL92fzsgiq5iO6Sj7Iw5YO5vtpLwpfM5bABOYWCPJb/p4L7
2ub8q+dryLyoaAfGfMcgFHhAByUfBMv+5frsO244uDSdqEY6bikFg55j1ZlF0TDZ
TX1BYrxOdSspYdQ3oCfGfgfHAaH/KfT9auYIaH9s53k4pbXgU9CyDEnRkjS/nP7u
bB9auprrAdow5rkTqKKIkIhwjAIjmbD/9jI9Idh23CjKO3aloeCS92lis2OiZ2d0
zenXDXxD3CwUjmz1yvX3z+UdBSBsczavx2oxkQ3021WZHy9Q5I8+kets70hsL322
YofBxDTmFhfHM6SmACJ0FHf4CRJ4XVR2+WjiXyAeJP7nzS0mez+6y1Up4kOi5kb9
JeJwVQobTwEwIQwlDNQVOzAKXQBZKXDfgWEnybw/RGFNhVF3SX0H9gTLNVWTZA2s
rcQDHCkbkMR3r0oSt+ZBXVpoFM8W54tLM59rlWV9UjeqNTB64LNcMiS0AiICKc/j
VCdIwzmTQVBZeoeijat4y1RlG3BePR0BaBkuYMMRcpHCU86Hm+nmOwquUoBfyvUg
lgASmPdwSOZ5UXFauV7Owig0Op/fGdnh/EK1mE4mN3EAMA5eBusE6ev7SGKhQ1rr
ROjyFRe+/adE99Zfp++vUbviFHFtdGrOgAvIc9sjYquQBeO4ady073S9zbQW/Btn
eXzAmcR6oKkPSjnNnAm/yStovVhsg8e2JhsMjxrxvFfQW3HqxTWFCwgXRRcrK4yB
SNJ9WXgMg5eVrOzpKV/2NZU5AADpi0QNQ+ZT6ky6PRTQv+w5E8VsdTOclik8EJLI
GSPRDk+FdaSauThXv+2LJu0NNDKyw0V5WNLzJ/GALicGd4iyFqFCNSMmt1ssKfd0
gXHCyDu5vgNkSetsO4JMtswzNCYucO71Y2axNU9Uv/SVclDPSMGF3F0d8xxCQ4y8
ybQbcxfJYqcUxw/clc98YWfCow4d4svzH41OWiQOKdOSgEaN7rxpz0Sd4UjSkXuF
kyWTCk7Zxexq/f0IyI6hpkIcYW9TkxSy0OVZhCUOLIK7Qz9NNfJ1ieSrpDJ0aLTZ
q7ZhRa5xAaSzPu8uDNWs12nzuPiD9bn7dJ8gDHIVokFoiQfak98gy4rgefR3Syyw
KuB/O+41I+pv4jgcvBXaHiRgh7Jc/7ca8wpP19pRRwQ0134tqRchog6vJEvWoYXx
DDx1laQt3gxmcm900OpARAT5FIxgGtbO9uu+X/IQJ7dJ+U+INHY/QkE51DN4q9rF
kPQcyqeL6r+SbK/KvKpA+d/aqIz2WFYJE8lp54cWy2VttW0fhTIBD1TGQFKRpHoA
5aOqouYGVTsyn69+3fVRoUuBD2hJCXpjX9wtwf7hN4QwriQhHKpNH+IC0VOzjY1H
KCnjvRGJQgOA5Ta2K64rLxLVPc3yQly+XzYx4xhxGha4F96oOY9G8XMUesdh7ULu
49WczyIEefhJgqmO41IP3rP3DK6U6T9WdPOG1hpWgRpCMNdPsbH6ox/SawHGsov2
MfQ7zzE2w17konkgU/9eXwwFYvCP+kI9b1/qNaByFHryKzwAJwSvKCBuUFV9k+Fz
jPz6pLAvCk+YKbGy24NhOWEqL0qNQBU6KgpFyFG9A++0x8LYUKd03+kyNnzWW7p5
DsZwfnGrBeV7OixzHLZVltmQCVO2n0IlD/CLmxF8Olun5ga7+bkyd8Rt0u263RX8
zaHG2EYH+HZ8nR7P/yKnF0p5P5ujw3UjPRUIG4uUC2m301ZK+CKm6Zqx/x0Cti0/
K0DuijRiqihU5h1YGG4Tsdl5yH9e0gdjFs3P7smiGV73shGdoVMhH903/1WkiiaZ
echWJtIAJY2wzdOKa930fDhg41mjP8svx3yLJ/aSEZpOBM8Ktxn/6TxZL2sEzTcx
/RFstyVX9Q9F+sa1PZSWjM0c7/REvfk9npZ0LKhNBKICtCPYrjp4eteqe8hJLTxI
DOIa8VYFMkR68H5wpcz1T56un2jIQfpqxLgNu3mjKzn6aCcnRMSuES33Mh2PCSZ3
AFtrnTY5PTfi2KRTuW0Z6hn1Fsc4qhH1+VLulLkDNAtLq8IepHuBx0qRqiGlHCQJ
Ir5i1JVFxi8Ge5fwGXSANXQde0hM4DSU5SWtAXM9NVr7A4pcKXnQcymdBLwzNMDP
Tj65CYKDAqWNvZbIhNI+YDUa7OynUOzBZwgOdiWcnD5M9IZvUb1D63CQE5sEhG/F
8zQUL4w/ABjNazcCV8IxUofoeHhIf9PqepeubaN16NpLUar6XUT1Wb36vuwHBgiA
57L8sl/5pDedudoV6p0pvhucE6qBhZUQ6WVcwBPCyVT/UQCuBI/uU03XG5Xms2I8
WS4lHCc1W19srXORqxhIJPiyo7bt8UT6g3xhLWCPl2yH+bePu5kauVTPmPCCrNMB
/xQFvnvHtk6IoGKn3jbLyrTXZ7nCUgwU9vdnui3mzUHg2lU4yAAFNw5aGjqydWqp
Tq5a0KenGJhN0Olen4o3Uy9WglIt7mI9raw2r1DvDVK2xUjmZ1O3mEQ/bbUJkais
b9gfF/F6VX5G5mAMwYQtSMe9Sudz3XGrWIsbnhm/l3CND5+GEcB/TtgeBZCtVB8P
R7lrBGltf2RGygzM/nuMRgX2yjNXGB1LtZ+KpIbrbT+0cP77SRt9AV5bE4RCb/dV
D5Ps4LNerFBJmyOqt4Jlo5dndBd2vNLstkHlPGcqXd/yO1TgKJHwEEmZYyqz8ZsD
qIRWcP5jPcYG302S4Q7JBe6PEjn0Cwcsif1Ub7tJ/c1uJsP5zvNdOVCRQL9Plr3o
aTtOfhD5JbdakWk6vg46p7zTifaiufzuqqLiUV8n2oLpo8FGWKxvl6VeONlevKo0
tSzrIrZrzaFy4ZawwA718F8ZHjUH24OllZElsba66I6rXEao1gpx7Da8EedNAyKW
Q1FvtXBfYBZYthbksPi3X4BsEKliXqvSP4V+SmtJGQ9MO/LjfMTDItokDj+3RXto
9wEdnwJope8/xwtm97fAV6+gTaaWkPf0/bf93ZpHycxwWpngbct4INaZsb+JFOZu
mltieDjgPp2BbjugjzFETTTjmRKvK4NGncNRxvmI2Yk4SdSvHOhaZjzyNoT/a6qx
P/mF0tGaBG3IKwBqGL7FZ1k+8oyyzFBIIq5tF0e9Z5Qk5hVZMgL7/JhY94DmsQWk
Y8TQmRmEI9t5v/GAjEfsvxZ6HYdqdrNWuG4nXP6E7W25l+mPUuZXNs12Wy9WUGje
XssIL2VM6K3SJo6dfhXSs8yfdRpnO3Gkl/r4CYw6JetcUkIHxc0PumiG3k+sOMpp
vUyte9N2XaSgGyLMUJ0SSvw+KSQ17rAXNbNqj/2mUAzLcfVMXbtaf/2i0OXSNDCu
/8oElILYqZknhbudfa3dWPgCHxHcegneTHJ9qsXvft0YB2Uus6SuZglkb+Cqb4MQ
y+GYgmap7iJ1Tqsd4CtexnUdlYRoLqrC/Z5kGubEMEx8opdNcNJhRScozFGixhxq
ogsf1tXfqi7KgR4rg/LAQ07e43O/gO1kMAdjV/DTui8aPB/Ab57/8nsG2XVWUUgc
sVhqG4tug2RE6XxurcogJm4SFFqy+l2FVTsgA4fnmAIxDWbdPVkFYPUDttAVBs4E
6KejTtQrGe7umoFODabXSarndDxdkOtd9kalyqo1UzvOumsDHHlOU313aZ34oqqR
qSSiTcJJdYT98XP+nijLYTdCCQSuKznzJVWYTaXKveeHcA9VEfoppkGpjDaZEu/m
j7Fad9geZRKnCWxgiyA0ZBjS6dv0jPtuK+KAuf4exGUtEI6iEbLcPynG7p/qixZF
PPkYmjaDagN++kVpsGZVbpmx61HG+o0m/Ek6Tr33WbyywVj5/s2tPNwBPkMPQEre
Z0Rv7xkR1EKC6teZ6ghlzHm/SeyZsIADescBa00sp+AFGRZS7yoSPsab0Uw+kGjd
UFxGPHkgT7lwt+Df4xNVcv+5L673bpZBgmEHrhfTEVmC7OI8bAUZgbQjJTpQHzoQ
9T7Z4RJL6mWfKruH0zT06EVI5Xt6ZTJs4HGopFafq1zIqqrkfNTdVgBBhHLk/0Jp
kPgO92CWkhn7c2qqOwjIK80MPrIv7jx/Yr8LtkzG2F9B+Y9vA9t1oNj9nezqMgrM
4FnBjHo5BxA8qrpwDoltW/RI6e7byTz/50ipszsTjnL1UZO3Yh8HSB8GpWVjwa15
moX379TWk2q3R5wrQ1N4pyP27ptntP0FE4IAkYhoiRN37WLzjCTXKsJjSirMt1QM
Uass/uzIyMpxu0/KcPf/Mgo4n5IazckC1eyJjL6fj82vXT30RnNLSVyY1jGZL0wR
pObsk+PjeocP9WBMRkGSzypnRQsAkftF6S15adM7QSHNGFi+BUeNlCtwFVQBYz7F
mT1AkiTyEi26FHrGUtTjsozCkuTonIxaBXbkLdNo01afXnwvYpPhDWcKZoJtyXtj
WTCqyJKWc9Zywi/Vj9JcaFOUfWMGQM5U8bVUKS1HuYQsxo3oXJKIo+1+RjRmIvRx
weLBMgFS4gBIjU0wjKiQxwi8v08WpG81k3Db9hqmBJZZzb3X35aQbkk0H8pup6+T
QA3EWc2cNFs8kOWuKKFu6hsrZI2cS46dCpHZIHXz08oHKys+Z2Vn8OGmS/MN39ED
il6PCZJyN+Q6wxDLZhD+y1aCe4ax8drJl0VsbkiKK4HRF36yVsP4qS37vcBPCEQN
JQgFqEcw3ZVfFvWwS418d7FEPkfWt0MfNc6oMFG0xAj8dukHU5yiafr7jkARSLHV
4MmR8aq3ygFJQj+JvfY9Ki66PUoxwEG/n/XeXmQRlubOI6AYMCL92b45yi/cqEb1
11AyA+IaSBzmW63dqv5LSAYXYk3eDlNZNFOaZKdCAxB3BRoxDHDMzTpq4QmGHoUU
HXlPT3X5dN885Sey32D6FNAEDRCMK7ZJGuUBkkLSFiGl2134x0Zw74vsnj35rzmq
TayLQS5RZFFrfEfvBcumQlllkb51ubXvD88UwbOLaVDwPpgaEzDtaSokpYMADl6l
AFh3flCbhzCqKmjRKOtB0t19LBb7ISkbqnn5lUAMANZsF/aSguVjofrgZ94XW3W+
pbsMud6ITAH5TVtqqxeDXMQk8/3PNHl1pn4lrL2iPzwey8jh0TBRaZdaxOeV0aq8
0RHPbmoPgDma1AyPeGeDR0UFU6J8t58jdWhKtQ9XWc3Lo3AOgW/oWxTDJb7xxAGO
DWgM81tF3VcPSWFTW43KncfWV15ddBd8WA41d0CHNahlUZvjz/0xUzamon5vCmpi
c38Yoa8nKZRfBXjWB5DK9s7y6Lemtx5ReY3I4HW15LlIAY27lD4uYm06etFluySA
SoGlJPUoy3jXKvIUHFYN1NpBG9mpJjZOJc/uH2G9ARWk7wPItX7eDRX+AUYRUGLS
uM4MSyrA76hPdNWrrskeU25NS1pkxlE51Mbcj+ADA+/TfoAXMHHE5MFuPTNlcWM7
1Rk0IgCzAUcjvdoiH6UqqabCsO82LZJUbQs3KyRfBWPamYhsrO4cJ+JF7/axId9J
/Oe3FnG4C2ebbTt7OHXQwS6cR22bgV2Sj5qM+++9u/7gUZSMgKwD89yMtpmwm++v
usPrw1FN0P2zzosQCBTYMEbDWxxkU5UmojFjnM8D0wW8C6vOwXWDAHc0kEfzJLaW
f6qNs2cgzE06jG7KIc5RJdEfkHVh3q6/sCgVWj6mH5pUqYJG2WlrwiX6dOW8kR5m
8r13HRuiH4/R/Yt7DYuBARKX0Kbm+c85BWRxfufVmzkV32CUe538ZUI20bXxDTRX
GNs+2+oNlGg9tHnnKGi0P8i+zqPUeijaUabG6fx2PFO7Q/Xe9RTvbcH/kE6eyp/0
30BV6C79a9NN3vb9ExMpEy9Lyg96ZKaPliRv+5uPSv+5zZPQTBCoT/wf9uOXtZzQ
nfm7yKGGYdLZOZVhVVPwNwOaRa05YUOqUJwZXlYLlblWoj2us3luHBEmVTspnWHY
UKOGZe7A2U0idvs1e/69qL/knpqe3qL5j2yfzF9t8JGD26LC0kQNzYqpP5O4bnHW
0tsCrlXfyNtsaRAGpiN8xLp7LC5zWbEofN8m33AKX0Q3iVjl/tbTJkpQm7Jcc68K
wlA3u5c72X77Zd80L0pUj21WVyGUTNSHdgh790vsU3OGhDL+h5YJ88aUso87j4Kx
QsrKp0aEVx2+hbzLanPHGz4gCqihxrROFHRIPVKjnJEphqqofq+UEQMYD5xcK6X2
5LQ4gtjO0yWiP4+I2woJz0jvRFGhXFHeB0XMLwkyNwopRFGi6dKKyU9H2mVbE2V2
tf/+ErA/7rbLVN2mSaIbPH9pTub6GHqmWMYLuwXnlXdIM0YqJU77JfTa2rToCCnU
RHrpHl1rX0zcM2jzo28epCVrXb0p2rlFFQdgcCoylRg2yIJSbTHq2C1xfBVEdPfS
bAHe9x4vnwap9UkMkyVt+QNLXhuTYCmEwQ2OEWKKUWF8x1YRciXhcRArqecyVNxG
IE8qqd7YX6zVin758yQX682wBYBlC5XoLUgsyTo5kPePmrVv7mYPxRyrfkwd3uA0
UnTo3nWO4otNrAOW95n9fhJONdw+6pPB0WXD5VODjz7mt4fsswz0XmzpQYiRWHEh
4OP+NpDl64veIY25yXtr2KwiQqdZX5cosX2eXseQzhCXwcK6KekluFttWeig7eRX
VYlRynTXyXkaAgKe1JB3UvZS2kDJBsZfCwNwHPs004QsVFRs0x39BcButD0Dd+1o
fZr57V+kWO1c3TzzTFqobGRna1L/W3dABvdV0FqrUdvgUDknPx7mijYBvuEq8lLA
R3YMrbCjufTVLHb2Dw8dJOsJ3JG6bFpH4W5m25FKGFdGaxebzpZvmJSFUatqMrbC
T6uWa97nxq55hFgkm/x9RS8JXG856ieYThtPY3etKUCO2uDDMZb2fp6WLv/ZPS8F
LPZUl4VdO2dmVNbl/u8gqCiy+vstkj9vlX5KmfOzBr8lizA0h5ezjZxHkTNPpB9M
WAg2oohG9a1BshauMGRgs/kVAjKV6wcNb833U2Qzm7dJTzW59V7n12fLcSPgSU2U
BzgTkXag1LRkN+4V/Ar2Aq8ccdR6Ja5OpAFNCbRcCk+ZR2jgoqqqz9tuiP1KhBye
qNXfQARZ1MkN6LdaJTbX3+jYLMxk1AL38sSJblUkHnudDRt9ChPLRSay8jxhNRmH
hqTQ9OVGFZPe7Ss1CCv/92hjc5zEg5VQa4eMoxKGQya3Bp8XMbsJSVo/p1rZ4SZK
Y7TVrlgqCRRHk7v3eQFT4DYcZCAq2De/bD/UMy/QRI0hoUGtqBPNKYWP1CtThy6b
TOzOOItegPXCKNhWWCnI1fUHG1YNuaea3ZPjY2520XMzNeRfii3nIF7C4neTwK8f
0KZkkX7kNBemBT4Ao/xAkapF0auQ9xQQEts+HWGmUuhTGtoEH88vMXF+H4aWIfxJ
D6iZ9YaYOrh2b0KMUioEKRQeFHntPZLPAthGMvHZQAvL1B5QI5nerygokjWlILYm
2kEaRnwL5J8/d0odF9P3QIbeEpUmIMaswRvEwpbxsd9dPJApFGLRo30GunCdbcg4
f8pvYARJvv8JpG1LNA6nlg==
`protect END_PROTECTED
