`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/iPiPHGVZCo4nhl6RRIwf/pA4PvM13X8a18Cz2RngipcHR7m0TVk0X2SKNVRF3Sf
eFjPxqwFI1r1v7BTfWnKIwpnV2AjpT5y5+0C744LIawPzQ2+DvDL3cspRx2FlYAX
gYLzUrY6D37/iwGyiI7mhwvc+kRhzSR5wmJ6vPGbrpJrYNF95/O96fziQ2r2XOIM
rT3o4Iad2oHNAiVJtBfumJbdXzdEr7yUNSXMaCrA+D87rV42IufXfTCpsm44i5VY
F6ZBOw1hgRtkadCM8zAvt0+EOZ0FQ20r5GTKq0fyGSXBNBRfT4sTlMoMaNTya31u
UnpDTrc1HPkBsvFGcl0w+DL7phOZVLnADw2ZHYxx2XU6/R3YGqwkbeDX4T9oTQjW
AqAt2vGHLKAkML8OkdFWJajJFQGSzX/R6MX0I/UQB+UmRFH7kZaChrqld52jsB1F
ir1RyCWrMifUwgY8xNLUq80YDfCh/q2baA6NBMDSZ9EBTazm9iZ2CIc1idCUIA07
v49R2uTKLnVISz8K+YNvI4Yk2oQkct1wzOOJRD1dzxooS7qwMYwNtNAXx2iS34Q6
wx914fyOUdRm4lcFaaD68K1j1rGdMWRUgO5ZbReDQum9PndKLdWl/jgbWU2RgEJ0
sJOTH0aBQMiXo3qvjBOtwSGSPv3LOdutVJyW6zAhPvrKkyJ++4Lq8BUBPj3S7c/P
nxycWr801YtA6uAJbrJotmiB+ZFfG9LDuHCRqwCdKOZ6G766R1se0+vwxcW34Io9
wpkaEsTBNC1xyN6c05cPEKU/5AzxL9iwRC0qMa1NWKxYJAdOHY1XVO0Gf/xRaw0x
VervgBakJodqqSd4ofuKhh4QKkGI/2kq7Yi6lhfRIJGy+urZBozP2GNsoezdiw05
3UkaS8PYynJqdEmqoUxOH+ERmQuVsf7Fa0KPAsErCHqmh57x6hsENpy92jBWFGy4
tv4D4ykJUpOq2qTEOYwVe7EU7+pTLcqgXwSa9fNUEioR0z/4SaGXlHNvg6sUYMlt
aAiO63Ymiq8iYyzs4WAvtkPApobsQb6z6LlystQUjsRjQSOrwxE7EVpdsIfHL4EM
6aVQ6gfKSwfvPkRfXz1jT+fzSX6gtoxlY5pqzMN/9EiPvPEPGbV/ddGUIJwsKfIR
PFnMVa5Lma80qIFM+4XwhFQXB+oPIQ67MCmHGTPi9loVnekS3WTpdybNSs0Zaqmw
X0wPzRs51dsOBLoolMFS2SSHc5BK0Ai2gXQ9RxvdI/7TO6PtVHb8OzMErVnkEsTq
xz8u8t0x8j9iZeViGOEYBmwT21acLVphQw+pJBqlNgukKfpeqJrtcue92rs9x23C
P+4FD5Nt1m2uEkTOu2e4jBDG8L6e9qmUgNsCQnR73Z+TiecmawsE9+tHhnWdXOWT
3N1cHqkJdkMmjzhK+YdfCVJRvNWj1ATlt406GB5FCFVSeyZviS4g8aNcFBLV7TNP
QLT+OCCBcKuqo0rz1OkFEQj7b1COeUyhGdn9yqVBZKPSkLKFCSk8WuNdssoi5w9D
qoLU2Xn2UnN5vG56aZN64qvA6hfaKm3eCZJpyN0jJPdDP70QRgX3Metaob12E9xi
tTXjKa/V7530pAVfTd3UpntNRVhzVbw4RAVHTn+XWQKmaRmMfXyPg4QNN0E+2wQG
UajGcvx5bVjcG5VjKMU6xo6/FjsZWFw+0FI8uTj50WASq7e6NjB80yNsy/cDewD3
fce0uqEV0hD53ENP+wh9KQgS5PMV1LDFUoz/cMdf6wYnN/ZlAiqr1XVT58CvUwTE
QfIBYT9f9dDm1Chp5UqZJPIdV5vnpM2pMpgiDSbts1mpO5uGifMJlfRfxpSSr+Xp
1AgdVVBdS2y+ZkvaGzG8YLwwytd+Eq41WJ1MiwI93ecNIkVEabU6PxLK4S+rkBGn
9VQhcgq5LVkPcILg0qJTWelLvDgsLgu1YI+QPVVeb29Wo2xXFcrwc2Jr3O99Y/WG
NnVbm2IQUX/92DS0SvCGEk+/yzhO3FcPnT2CPbGZWmWum1K3QOV7KtqCcks9+xQH
0kxoaSFl/bj/fnb0KKplIs2k+kmwoppFkoMKD7JiUPc5Z/66TM3WpOl7GSqgJyjl
jwE3L2wwct5oQe6y775soFk5+vOJRtUDWRFoCNXXa3I=
`protect END_PROTECTED
