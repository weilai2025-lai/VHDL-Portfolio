`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ee+2JNeoUICT6n7DLH612XTyLBWWKtcFNLtYT/kh+4AGZ3vB50rISQEeh0v072R
EVx0Z7zdc2KQOfFT/cE+riGSl5+Ue5k87ijf0Odgwg+uVQawHnV5FyOvMS2T6uil
sLmq/hMLHbKjgKKbsUXuFBWNfwUhWrNvNBv4q5ot/e5mnZFqLNTbEg74BK0Jsxft
Acrl/FTv+CLooswA2A3mfB/6o7ROYmV2eRCZHL0CGd5nugdoKAmyDGj77BwGw8PT
RSztOaYday26+FloHVomPpNhUjAWgw9ULmom8WhtgLOJ6GTMGCIHo7g56LzMSuqB
6cOgGGpK+hEzPZ2cuENYpRKP2nvlkCJt2u44dlgn0Ei9Ynqe5l5bpw5y+qwp/qwB
FjVq/tekZA6ce+yaWSMruFXo/XoaAW+YzMhC/pt+B8f3dCWvHK/c5zfEj1UY31za
mkFiP/ky5YdKMjuZuQvLRj5wFDgIETmMy78TKUnrBx+nJmDhiSmqYpL5vFZpjo/0
ruR0jMFjixOsm+S0q304oAcNbXYB+YJLMSwsvCvSAyvTxiNcTbBcgx6/iUHFUetP
xSDrlY0Ww28azqCXlOIH71gH3zP+VIFk37jIAGjozkdy8Pn6HSk8/IXjZxRZt1qq
zCZaa6AT8kD/j7WZPTn6FLHxB44PqE+0ceRILNsgTsbIjkMdQx+wyA2WD5v5kRzE
Gad6RJ0Sy5+QAfpQ6vS3DOAzB+Os8x8FfkeAV+FoUvU7fbvullmRgnv26vEkMJwI
HCh2v1HBPjBCEWP+/sNFBcJ/9p6qBGB3E9oZO9Spmk7OH2mkh6udWGZ0q1mPaVEw
6EC89fSLTLVfhNcNEIKynqqrrJz2DyrNLRvRZJh4j5CPqdqPwSmh2hPBCv0Et1kx
c4P9jRNLF/sCduPgK5FbDh6upWk4+7rpUsFg/csPF/nF8T+o2MdBzK0mcJ9whyrV
FK8FcFitZnL6PVGA3blelnaanPxw++ZN/PK/KqTA8Z6mdJvO/MipiVmP41q4VBri
vL7oOADKVBGpmjtM7a3+nVAyPpQq9UBIPWwJoS84c49LGXJO86wO72sd+39gasyy
r5NOrdVtJTyTU5r0Uedb+ws8S4HJNIZGlCzmuetW5ekncc2T+MtwsjQim5OaBFq2
ioPnDUNWrdLkZzjg/+CSU/BTl01nEH1dFUu0P5XmLXSbmaKe6TXsW+Cxq34vZfX2
102JKELgJvMhN5MD/Hfs92bpfYH6No7SqeI7Gnenbyv2KkUq93Jsef75tckEyikI
DU9qyhoK740/NlzscoyTqRaMCtJmtr4TrNxKaZt00sPLKWmnvNYS32B/m4pSSnJ/
tHoyLpOtq7hGoCOTzNIZoXOol7ul3LOVJNtua7DC1RMpk7N+u0mXvruX3la0EhIN
xUWBTDjltQrxtSYLLHo0xiWQAPpzhD+idt0Wd33gF+T09CKENjh1EoXe3+HZqN7K
rQi9N3gIgJZjc8YV5zinYylzznLLwXFVm/cFW1NNOEnRsxd/LwLOsKdROih1Fg0U
6EwdTnbGl2TDa3uh+LZbJ/AwsegNdFOTO1I3LDbdMierxhH7FReZZaSkFGwkTqJ6
ymaLSAzJIjtkRBsVuQkMH50yioQfHoi4TwcEKaSO6jEoNeoyaSY/q3SFX5mM2WgQ
kl9akkb0merUP2fUgY0Ut69E+2cSL9M/bWuAmclrpZFHUJ0QVxx8ed/zW+/QyX4W
nqI+bXl9s5TqcFtWtE02iniEd4klEJ0Lk6NV+t3zkWZVmZbNP2jdrEgqFBnfFHcQ
l+AeUo8ZJnOG4/UFPom3gru/77w+CiWszeR4IJ0mneNhC2bh/fOE6YUdL5SXT5j8
ZMtFkifbyTtmDYO+EdqFpBaS1XoNXfQizGYftvLb2zqBnvMnWu/sv5GEsGOgi7Cg
2z0i8Bs/4JbsiWJ9Cpw3zbv81VJs7l29vy+7hRNvb/eWmBkx8YokmjmK9LBnW2pp
BlnmLcB65D3+CjK/r65qIQewmcsj+MpD+2gn4afYzWKtZ2pnvpQgxEu5dWoiFjCh
q0nL88YCn3aPm/pCb/qcyfsgLftRB6C4Ydbh40ktP7kETGev7nfVaybny26nQR0h
0YO2n9+x6lvKzRvc+fYiFbiU9GpP5bPi7dShwqfWvXaYbEuR40ku6lQq/RhwEVj4
s6U/T2dkZgefzQNwr8TIEwrvO4fsap4iqlwX8iXvXSd+Kfpf6YoYTpWTob/fKVhh
Av4hiLkjfrdH9KMbdWeDzHySRxH6kXfSTmjmQV2ScgyisvC5/XXXZ96MdLNq2P6P
ubQ5xCcurK9/XGXbcycQUSz65gLAbSXGDY69EWy4bjHFFHdimFOXPoo4BFAq1LVN
yr2y99bQEXHJA6/kslJ1eudyA6inOJbJRtHDhmoS7ZelT8YQYMqsFG2EQx14Zygn
0pzDw1QFOIBoESvW/lvdlLhDUsA/V4GyjkTRFKe49m+bclr/a1J3jHOfniOh2XsD
X1dftfzNVql7WhcFv/goKRnSIz/dQCD1gNDR20VYHa2h1pXY3kDBf2apQxgV5AM5
Vb6fSr56y+aH99pm9vsm+roOGK+VEfp9TjlIAbA3KprVMuCvTGcuoYbFjJkfoC47
1dxGpR8DJT5gvTzDH4XVSasmWX4+5pAorKEg9PNt46wFv8eF11lzrQo+lu5k8M8U
bmLqWTOPwIlRhQyk2MrNOEI5tHfRvJBdr4Yxc5XiCrFSBLKV2EGjpHs8Yw0gCLpJ
TmGD3HAsd4lpQXQgGInspEcKqMduppKSMWETQJUu67JWj2ZNdgtfq+5T1Lnhijp+
AGJWiHv278OdqEl7hvYsCVQ9FhTK0Zeu4xEIoGwEjt+aP6J8lGnkujcZrTT1SKVx
4FilXhuKEM7wpbUwxsx7LdJElFvYwus9WbBM7JPB7KFupdkbLVyC/p62m0ozPOiK
sqYYad3NV8RK86oDEelR0QxTg4up6RoN4bytkQuTHUYxgA0se1NcFiIk7nMCSt+n
Z/oSxHUdUxOoxpCvJcsYQF+2DYWLYXbuzIGPyu05L6ptFBzuUoUpKqVvMtbT0o++
Uk0bGju62MJtJVTfIBt6OwBZDitSdIKZJuyLelCUcks9VBLQtAmXCWaEf6Wx/h3y
HUFZc16u7jMXSYGdjd0BphFP6eaf/n/+cdCPxDoQZ/qp+R8PpUeGEXcqI8kBgTkW
A1Q/5p2h5qOUAMXDl3+m6F1eU4o8lIxNzhAcCQb0azyw1OD+p3qhAKH+JCKYZR5H
fASI+3dByDx61s+reQTeIwT7L3EP3diVpgjKWUnCkLSOJZolwgl0Znow+FxtpREs
bmBdEy+8QssgHXD1cRCYOqiH19bkU8NgRniT2OlozsEKtGXhoJsTScTFYdiS/dRt
HmUUF3WBx69L/Zm9FoWNBDZq3JDXd44zX9kF90a7mrh1gIuVYQzKb7eN/syVrk0Y
QXVIGY9Svu5MHH//1oQ8h0gk9ysi1lY1IixB6Lc3XiNdjzP4czYhwOCmzypczQd2
cIAwNksx9/8ZdtNRg/un40PDJtsI3sQApqWSgQwdYVBKVq2inAzp8wZhloSInj7J
SURvKtPltrDGYxn0fdjb7P2QaFw7kMRA9q86GKnfs9ez+aDNwlqfZY7bJgYt+TlU
CCNrdQwf40ykITo4+xtsBbsBnZkuASrODB9z1bR+4GoebOfVEEnMvntaOATgOi9t
YfoEjPqikb+V4VeJYriW2gJgmBJ76n8KxgODR9ywdJ09xD/ulFCifwe6/yr7HRnO
FJgjoweFcN69f6jQnaPv4LH/VdHe3vu7NHG3GMmnsDXneG3eNHArHvHQwNkU0fGp
bDeqpvqIb3meWhvR7rkwncLBz0bO3CbD6R2CTqXosvM9iHlHwreGBNrW8ZRtLCsw
rBBPa5fUA5NYYewb8l7bPti5sKqcs9IZIAfeHc0nvitYkNAIO0M+SbZf0lC40E4S
VEsyVVYAJFVd2JOY04BD8Ae9PPinOLOIZIFOyeZ3FerPHBC1uGThD/62a2weGqNd
3JM13D9I4jOGk5S8Dm86dZpfoq76Kk61Rl+8TPeSeC1rBoJvpvcjYKCFAg3ceOaW
tvS5f1wW7swM0SaWZnYe4QXUBSh7vCpcJjdFecvYNqilgB2OYl2p2XH2+u4ihIIP
8x0MNtU9CM8NB+FNJzawzilrt+e3Cx8TAa7lcSVIgAPB9pqWR72LgYtjdf+bIFkk
SAURP9MapEVpOKlVRH5zVKl9YPcG/UHrBCh2xsM5EhRQIR0/Ep8g/M4/SpR1vmpc
N8GM7JhxVBe61MPg3V7XegCymTFrPY7FQTilfVv2Jkk9NHMRYIGPBgnFNDVUUyZb
eJYf8+LRzEjQI285XF9Z6cA/WhYXBjlQR29MN/Jb2UE5+TST6XZhDndkPmxqBTA2
Z0H5peeuXPUzZZRlIjGTrKYJrsOtaAgH4BIUbsHPB3tbRDBiYXj5gZBTqxoc0jBG
rKXb20CFYmD9xfZeBQ2DJqlFbxjPAqIRbiDVdrMKVPPq0w099Si3jpo3QNru871U
98s/jWxxNfL9qk6G926fcRIOsllKRIbSHGb3RFIyvvv/JhOa0xaAwGUDT8GSD7fq
Damt7Iaci5rvNMPB9anEuUqDAMs2Bs6MvIPARG8NalGiI27o1wW7VFQ4yKNBB0t0
4PENimgvXbsUPKQ6BosR7Gf/D/UK+HCiy2vOddCKsVavyWOFrcm3deXf6st6VkfM
IdWmXRyyZL8tUI0CBE9tkQh1BKy/5vpqX9tggF8FVsKXon9XgOuifGCGtqQ2XPik
2z6l9D4BI8MRGl1maCq3wVGmbltjZXYsMgJlnxhR5Cl969kj4/MLyyTVAVdo2kQn
awCWYdSUe4k43LfSQvshuHAjZR7AgjbtogeZKdXtxGVD0tbsYJTbnQlrQ4EgNuT4
bIsh6YeyHQ3htp5MZOUffQe3i7+3zH48QLTxuzWtMX21ZdLQgGI321SdVLeHqMah
5PCrmn5072hbgZedrn6OUqUttwx9wF1qcr6tahCp+2+FDtp5h4Hx2csZlGrqHmVG
gW3u0KMQWjWhkiexhtccy9GGFK45g2P3W13l3iO5SQCh1/9vcK8euDiHshyvnXwP
t3EXRa5mKLJ7KMuvCW/NYLr8XH+1pim0G1EuML0WjBRXKkiX8IUiJ8KRt5ciBoac
6rzy90Xu9JPmUEqsMmaqyeqOFz4pc8dLJ2lG0ZgvbQwMdmAUXFUrUkeYVGLdi64/
ZEjZku1mwR8t/f+wP/rUUj2UpLsSaY87KYd0rLIBdKLmYfx7utscOlaMnN/1TQ1W
mGsThQ/sPfR9/fauU3q95nSAOEtBJi9QQJzApAM5cvbqPUwR2NP1MWrSfvWeh/4T
1VGGV2/r3xxn6Jkl29Gg0nMIOviOPEYVKvd1D9lRAUgQi8gU/O0K/yPedNm4MTXV
cEOdQCEYnHyGWQQ/Fp4/9ocq9NNvMiZwjlT7Ybmj1K+5WdQdLSSpFxkSuBfRhKDk
kZBq331YWxf4fx+C+mcQlf8ERB3y74K6Y7NIWlicgi7WAp1I9M2cBbkEKFIfeU+3
VlmD1hW52TRWwUDnSnZdWz5TybJNh4GviSvlUjXDXb4hG1xSRw04kKJiLb97rukG
XVUwAPhJdXIoWR6ERUy7Rhx3LSyT810fZnyfI3d5w4KnCcCnW7m0l2bU1AbMthwc
Bt+3dvu6Pr8/QucRtUXkgrsvjVD7k7ZBLy1J3p8I1tY3zHkZ4bsTHfSBDMdN+3G2
xRQJ9cvrIlFzkCg/LwDr626YJyBWE0hHci9z8/nGhDDhRTlHMy1A0KZx2RUy2phv
l0Gb/8+mix+7jeyFSp4m0u9l+ZMkNaeBVr1vSKTEGLNAYNIiq22QV8HaQ5R8GX6p
8KYbcA75DVCqDmZgqolt0crUcOiDT34sa9t84SpndAiQyHhamtUfWYB8Ey69YGnx
f+z3SyqBGkgs8Tn6Q1GTuQMOgPL+K/dpGgotCIF7YdlfmYizbiXWcIGLlVE16uOv
HqqLV3f60sdDTMmlqdC0QGY1YHwd8KCDeSkqZujhs5ZYoaGu2W39Rpsjcxo9PQoo
Qr+Pte82LHDQ1KywgVamLMYdBwz/atX38g9YdBa9dTdRDYw/KjRip/SS8HFXfoP3
O/s2XAkEyzsSydmJ9yL1+88IeZYUhApKDGT9yop8hxmCSjzaZPlgisd7tr1QBqOj
cUwMsKP4V7/mYjwdLoEzyv2Y05MESKqQwNL2dKBjz8ajJIJiJjAaaEK1sD9gtkFQ
9mtahK10Z/Zg9PVJ+W63bGXWKtyUTH59WDwPpF71dS2Fi4B5HzYCxAgpXHd0/p0O
PVpJAIhJXl/1bwGXQpK/sewxkZTp0B+iMTyVuQQ1Pu6LkUPAlBAyDmMKchl2UF+d
I5N5yzluJ1ZlhxtAGfd+MLGMhhpbh/YA4K7aNygtcfzUzilpTEMoF8TNNdRzgKLd
WVK3egRm9Fbg2f4JqNWymd0yZauV/v4TTQd1L8i9KhTkwBEMlyQg0r+/nhFzHv2F
GkyQ0a/0lFbnx+lGgVo1Bq1bCTu7jQlfXjcrFrEdINNYEpC60dMSTdb8gMyzGyO9
U+L4CDTORwOgkiLQP2QsolwtMiRmo4xgX65iKhA/vieebXKxRgOMs/qWXpXMgwnm
LZgMiaE0nqtgZ+x0+T79yfYbWgFGcNzj5dPO2LukZZJ/HW9jAk0knLsOUgJmxPDr
oa3+isEe+9wNo/oOrM+Len6lypf3ZFOw99K0rJEa4LkmUwyXI8T012u5OcJcQyqp
VfpvZ3mlf1YlQBaaoe/Mg/J1RSEPJepxojFx1g9L2ydyRj2UToiW4idejJy66dRf
Q3I+JoKvKr5i0JrOICYog/7nRmk6yIrQ+2Z8AiOodjCYtJspQGRl0UqAMBPp0RXf
FezYkGOFAMeBFbNxDIE4t/pxJi6GVpMkDL8NUs+alhjPrjknMYFh0YFR3slV5wbZ
5YcbCYEctBWP3gE2u8r7LMQAWIXWRPS4K8HDryxkH44Mqfh0GIkNIV95J2cyZVX1
JTM+TVyzGL7CtIxmEaDQ1qC7uxaaQugT2mut7ujXu9EQCthpIAMdIcMYCmTpogEy
rLNTkcxTPvg1cxhKv/zuWOGKW9CZUq8EbKTrRlRzOD3HRNJFD+JmKeIjz1esD29Q
K/GkNxJJ6koGFMrJRpNWfFEDgGaPxaTTv/mwt5Uc5+BEUZkcpdHiPY9HJZmFASH0
o17HBoCzisa+MELlp0TKvrum8szOalW3K0sFONBFiwTUBalvAlyCIITXycz6AK+P
2ECdOi0EP8Av0ZyoyJBU2DfBEhBALCt9ZyfmSk2Ft5f6l/1i31G2zYZMCcKjDZxQ
9Fgu1wxCiXN85MUd1fAv4tAtsMa/MDMJHrRl59+/ZMlsfj4u136qoGjkfK8Fc4Sp
+q8bNoEzunMK3Jyez3KF9Loz+41TR4COQeyKeTNgCvpetcRw6DRt+/pIOlROTfEu
bAitdNBRKpUtg/6RW/GSSZ9FA8RnYg/RS96XR6MDEmvXrTp5mbIZS7OMs8sl1jyD
tLSxF2iW5ELvOYv5qjIJawZyn/++0yif6/LFgnOTLj/fd3L5YPqDlosm/+X/udLQ
cOthWDN8lXMIZ97BtMIyx/05ArPEYSkFSAZJwXXScnVakYc/VO+gcVN4a9b79iAX
qKmiUoQ15wycxRxollpHVJLjvRPlVYg1yQwAYO92L2czmOh18//XIvCl3IP4KaRU
NobgNDKdxEHx3jYX5Q5wF4JWNlBMXwKp1olYhljGmv7dmNTNVuZNIJ88OPpVqUXH
BsIoPW5JwSoh5bqkok08RluXmVBCu4r5jbDuDHpIz3cwh8UefTc89Mh0e2cEwL7D
UfBdHggS+YotbB80zqsd6hv69Cl6slVB5fuYlxY9/I3YvvXXqZ0olqKYpRgW81i9
fpse5979AzVhCb1toibmHxvV0sG3pPhkfqxqwWkNK8MzKcDrNhAdEv7+i5UJ0YML
ul+mGzwlgAjqs9+mFNOfr1vSJn+2cnoLRDViIASHAIzz7uHgzgrPgrEl1slBLrQD
SOwiPI0LwVxdtffA7It7hbq/HgHlK8EghN++sHhdUWydYoON9/AoriZXfOFwEBBf
EzldbmJoUTAcAQH0zy3eFRmZTWVQ4cNNrSSt3aiCEIGMF3mfEqEvL8HoQ9P823xH
DI/7Zf5ZrpjV0qgGzACkTU8aeWY7rggExATB4XUA0WgexGE+KhSOW+EsArMAn2Mf
Eq9B0AnIDtGH3GArpe9DcL6b5DmCTt8/v7JL6T8TPuO6fTFThoPi2SaVI9ZbiTcY
rq7GTeW78wfRSHbxIvXZ4pkTwh1k4wdexruxR6fDkvSYrlvoCtYUoLelol8UMrUs
Hy/+18bocXsufqLTi+7pCq43x0JDd5RLx61ZWuvXA5PlIEWYr5jb7fLWuwDN1NRd
k6AoNV6D+T3QcRlNENyn3LW7PehqnSIvnkPjkLoF9Lrd35xlQB+bfOhW173Xrhqv
wQuDCU7qy20JydK5W1M9cbUcag3SuRn28H58akBGGRlKnTd36yli7fGnAaRAgV+b
8A7pLmwMRaLE5TZpcfiIjxYaYAKd6uwPt4oQccK68ajtHw7xp7lvkAVBZ2IvFYKM
bAqv8uA1V2G03pah+zSRsUiuw1qSSgagS+jh+rFKjX2ftTN1G3XuwlHfHNwE4aBA
Pv0CZlAQQkz2F2vdHjVjNq3UdkkN0eNTtiibCOV4fUc4XAe//1g+w9KjVP2ZQX64
UT2ZkOIooR7OcHDo6vd6kpuvcnI2+oaNyt2HlDRXYqcmG7BnAbJEahVpdG1gCqeC
K0NoQY/Yb0Wdco/EmHxd+fer8tzkvcQK6CboHuxHPIshSE6PnG0E6WYP62Ryz7mF
RRiO6IZN6GzApesQZ/XU0xhiuRu8CZo1XZbsoztrf5tcnV5wLPP0kG7YgK8KIVLm
xdqX9MNQoTibJnIHaMRwLkiuCaq1c/W40/g4gDPTwDgpZWzO/mZmotMRdRlvx4lD
3pu0hDIiPaUndYKT/7bamCob68gTwVqBl4XOIJmr8wpfTh3mJWRE4ZN0zgB0fyfO
s+t509FcnyTCn74LilFxaSZzoJpA8qq/aXA1oJyAZKwPCUakbf9UN3cO4WHXEpV6
p5Qy+RJ4AEj2AYqmtmrM49l9AE10zmpanJCDjGK/fyqhL7VL97WSczhr3v8joB9+
KGAhBBRQ6F5Za+FoMX0N4nmsI6EREE2reazZbnuzZUCqa3cVmGGrcnmlcCpA2cT7
ULUGp8SeLZ/rVAcjdQtrhwmbiUQTnENC5ecYhU2l6RPd6R5N40aFT9GXdLUmQ7tY
DhdELniag2TGWvJTmwaplra6Qf953o+yRlyjVZJAVf35NJH0Ou+31J15WtGoXi+m
kvxQq5xfTk+ApQFgsbZgyzDW/Pumyp/ptsDBT5rMKCUjt83m6f2wTf3KvKI+d4ak
frBNvnBY3Ya8fSceI2D7mENuh/H1gae4TSdyPCb44CMBzctb4I1PTYbWCxksj4rr
tVFwC0JanFU+Jly2l3n8Y74HJT1+pbXYHSnLi7oYNbs00yHSb3jh/LzcQa9v+7In
cPyULRpfm1fbcvXDQPftmYIP5vtewL5MiNC9u3/Gro0nn8/lO15sf/XFHY6lt86m
sBKcPZkqLemXhbCrC9YDqOtjK2/KO56XxqQ05GmvJXfmqH3bGXFT2pKDqKh3GYyF
CfU9Ue4T38PvjU6BsciZG8Ghl4ie4n9K53e0fFR/ZwkYG8TQWRxoq17Yk1kK7DXI
mhqwV76zcf47kvwqRKi8bdyB+Hyp+LkC8XVf7ffQ2ldb+qSMOcMoC1lHEa4oGl75
CW2kHXa2Lyyeq4CeLm6InCTM9r/8FspnTs4npqfAoHeqsa7ncB4+yKjuI9PPrhBq
U6v4IM4t8MyUuvLTGRpt+rs/5DA36cOpBD79CXmGN2oqPdLipU6c1nRYSnHsNpNl
K+FMK5ZuugJSl4JfOypFHPnW+Ym1NvXv5oZGc8iuxm7z328Hu7xG0OSsK/w1ahZv
J0WVXv+6xLL0jzOA1EcmjpcCgj6MzjXvbdabaN6EdevSZZeaJENUQS3QUetV2dFR
SlrBqpqYg2WmOccU+JqkMLp1XG0lQUhxXjkfdiwgDLblxyGHZrNxOuHZAVBQ6o/U
G4dJdD5NO8FKVY3ZsGl2fRyIUqgYC1Dr9+MyoYxAAlI84eHYAgUCBWiSvG5ebAht
mhFqvnHD+JEVDK/LvGRzhDlfCQYvHAHWWyMEFHxsY/VceIuymboiAyc0f/KZ/RUe
pUP5jSjUtjf5ei6ynVCeke3t++jagrEQfTGLS1rmx0gmrG8a8xV4HtDbhuJNxQKi
0ZX02pY6etyrRSmf13HEnYR/MXgKVagFuOYWMUYANn+kkXRaOsdEpW/raZZ9+uAH
XZmo2aSF9CVs6BkvBkVBUptWbwPrOWwPN3R+W0X0HmMyVew/JKEO7ey+hQ91qgz/
7n4c7XQK/+UfrGgJaGuSHKb1QjX2pBfmzpsgN2Hb2M46vrzOfrfVzspAq/WUnCR/
bmqYbT+i1k/N29XkiEkCb4vkj1ZVgb/yH7KGwj4pPoErxHDdv1Q7thpHJtt7/2PW
oVG+cDdFOuIuwVgWRnNb28avNP7+OrE5d385H1WZgAYmH+OWWSBsWtJDOYAzzKOJ
ejRYAUBkGcl/1PaP7w2HaJBlM+FoVdlVO7q1Dr22O/9pvBGAATeAR5aVQDqIGiu/
HIRxKqUxYn/l2UIPrQhRUYKGFIpdpk1J5P+QQ74nvaKfiDLpZ+07naad/vargRuf
CpaR1dtfyZjP5ktpCHP93ID1FV3S9p02W9TypfkVa8oEVdrM3JJOKScUleBXcEkV
Bj3QjueNSBGJ3CD0IzoS16/nP2cmq/V76Na39xQml0Bwkom4EH3CWHegjBwdtbu8
/0tSXeCEGX4S8jCikex/GNy0kPxU/WdQNsS/vHDlmtyAXnmwRUwZwuzpFZN5BSg1
pD20VlfivENTUOutmG7cERkleO3N4pXfVBdlr6YBlJoSjMUZEd7+/4VL1gQxLRy3
d1qrCnBpo0MQ/auORWcn+pe5XXMwSkIUZUaJeWyFnjs7M/h0F0+4r5IgBWqwYn+U
sNLYa0MJ/WhwANkeetf+qr319pSXurkr8ncQbAzYqZtldPy5qGXbfFoHHc8widxB
NoC1wTgnhYKjzgiZHffcJSO1Dw/Yrr1tvwq2FVX5RwBN0ZLbbLxNYKCvf2Lph563
jpZYDK9xO9QJuZ5A1iqQwgsthewR4cq8trl0Gq2izH06GHMStN2lRI28Z1T0U07J
ZXCM3RO/KqUrtDqsu/F2ycT8kq4MVdSNxTtnS3h/rdVQZs/sChp6almTA8ByTblz
kXrYGHnBVNOq07ds8nnFzhCDxmnqNqsITnVpXypOHV9f9t1LJHK/6RcdsPLtkxe3
95bICR/FXMyD/zB1NZxPMtc9h9TPvZ4UYjGFklO3C4pPPDEZNYgXrYfGuhiEiE+j
EIPS5x+7IXPJ07Sqh1ZXxcuk2TMT1875WTKu4nJVzFiawONZVTsq2PcSJGnZ+Uf3
gE7bXFOzQFfYo3ai8MHxXcih7Mq8VUCJsThdFc5x0dtaJJ0cPtLnEcqbmWId2FZk
7dXdsL0u22vQi9QnL97OpdVywuJ0AZV/N4uNwbmt1ZDjRmllm0mHPXZly1zVJIdl
932/hyVcLTo6p/tL8Dv+HoX4+MbEvW/9pQZnn4n9fUuX63cuGmiouJOy0TSde6/Z
ZtGHDAemIvsQwMX+ToTilQ6brP2dh+ptzTWSbgPGgtQAIUeUMZ4sDXSTesmtqmHz
alYA9jKHGlW1GeAvu48T5ioESKEe01yiIjRGalRZmnfzB4zOBS5KjxDqdhLW+ZEG
LLdm/rFkVjdCuG69zzzRMQKDb2z9KoMO2jOfxegVj9T6IMt8H6KvKNEXuEr8BZAg
DfdsoNaBTHJ3WHDXoATy3j+nnMoHigETHFL835triNzDsBqliSeFXHM9ya5kxumC
jClj8GU7UJlkhWpYitHHzf+ZWuw9JdRSlA07Sgi7E5bb2fqyLJvLEPVEWAPrI05P
wXJyJP3jKYpu+ddaEZLFoEQ/65MJLqXFsCOa+l1t5uoXvGiR3yB9Z0G0KGrqyRqv
cmydeetSqRGtC/r+nDp8j+cjIPGfJWpysX5q/kXW5k3COA+WEpG082LrKBTbfmye
SQY+cxJlEOgWMzlbtfS1xxt3Ca1nUp5Pg+fuprRZO4DdZg2RKqJ1ovTOLcCQekJ0
j225cTt6/Vt2zsiNRaDpoEpxd0st2PDgnpsgkrqGIZggQF1XJAjRtRBR/wR0Xt1n
GsLXS7dBELLu35bIsFWQPRaFu3NXm/X0lUWBzCU6RldYicL9aEnBVdIKg/efw4n0
Xw02MtyvDcmDZSal3AnN7QDFQLqDRcP06dUJIlP+HRdCFQBpUUHqfhaBFXgwRTjn
W2ew+WXw3fnOZCx3syZNLxw+7jMRv9DTcccw0eIgwibNOa0Nue0VUHrBSoCnWCPn
+s+hHfGbGR16bHqQnoArtWBnh4viHlSPkruZsY3SrFEdwxezFeKn7LQqe5Lb0Y8E
QT850MQjU9nWpjbY9n05ZRGuujY7c4bpzJpgBR88i08pfUFJyvWtOoTGDvZjfJ3Y
I97kmAGb8zlhQzO3joWV6r12V5kGuW4qmoNhRZG8qqUCgD16hyvMC2a5whRgsjeJ
KwvE+L5QYFtXkPwxTfjCJl1rPwF5WLn2e7rFU6C34E03Af4hJ3vqhb7uIMYMSiyM
6ZWE/Zbf7pD5ppKXCtrmfEtoBUXeyy7pinN3fxOKlJFxIU9eKt/uSKMJ5MH+0Em0
8YJ3NsPOnBFZhIKILJFjNcHoGvQxpAMo38ytdyhtmr4387LAWqwTv+jQj7AQlwTk
4L/TGkUWFjH0lwyJhTrERTDfhTwpRUY1QJg+lHGBlm4tkPz2FBKYP55/JX7gocaA
7PKTlq7Ucy94Wb1tmzEMFrLYzMCJzQXkN7A4IOiRrst/FAnUvpfKYUO6fA9vel+G
zgcB5Qtmc4OJ2YerjX+ZdGyeIRhRZdTcbnkVU5g2UPXPUyrIX0AxEhmp36p1Ollx
l+uykVKQU579cdGpQzQx1c8r+stg5Mku+VOC/b4OdnWJBQvINHI7ddogCtzyQ5Ar
CU+Ru/LCNPIfJdD/RPmkF07U6aHwYBz/YtC+TPRGMLNR4oLrC1v3yF9N03mksrur
jZYe14CWXXzZHYtDIiZYIVPYoaIJC3XJobkoflRVckutBWsqdgcY40+jwT5MLNpZ
auc4PPE7RXvzZOhW+V44y4a6MsOa06d9ivUJAnmBHj55tzycyTsxCsHXNT9XB+Jm
EVrJj5m6JH+n+6gatOJ9+/nQzcDpfyXzW/y2eNyiiLtVfqc6nISaZLfvS09zpVfm
5PEd0azXpDTyAFc4H5GEE/wOhQkyxExa8zGJEH2Qdd+E7Obqd5Ly90whfde3cJAs
G3cHV95sTrqe1+EF0MCzpBGcd0BG+CqHtNjq7bIapqOOx916XCAkdcAaDqQrzsiE
Ir4SruAl0M3nR2kdz9uR0CyuTKouQdfFj2PPFJJm9Q15XwESkgwqP1hvU5VDcemb
I7dviTZpZ5HgL07dpZtqCxdRSrmf3KSi1YvsnprfMIluUExPmYMryBgBt1sSeIfp
siUqk1PCF2zH+sN6g9rQKl7I/Bb11gm3ZVHXiFPIEfUnwXIWdLbbGiC1gomh4HrC
/nOESd8fthC7Al4Dd4DMTCmrQJ7ge8/0178vWG/f8TqW7/DKiZpCDqwZHR6kwJD7
kpdwxRn68jRnE+7IWAEVqOGLUwqnpbP26n5kj7rDchOxiS6FKSoCy8r4cGt+CxWu
85rnUrwxh0gbi/bN0a/aV4eWVdBsJRMnnlb0yWnuMcO6zvYqSSouHeeIPDsz+ibm
F/HD3c6yN+85TujyWqtLiiDUGp3TRNISmGJITG2hheRXnbbSM6okdM2EyYxOiEZo
xUcTba6mg1UDd3AU23ft3y+VkqF6A2HJnaOFTqIg1eOhdA0xWA5Qrs3ePLL2jDIS
XPVYFUSSXo1oAjsbkjGA2SVy3HXuSDHmLRlj5JbktGSL44rEEK1RDJnhGCpK6AIG
0cM464dsEDrJCBWjFZv0b9qLJ44/z8OnFqkTwgTMBjRy/B0On+cdmbVazTZus0EP
8fcpYpM9xp/Ps0Clcd2fY4gMdNMl3oAfAWnqSNOzzxpcMRzka5U032jvxEb86cpA
7eLa6i4Ek+933NGU0E96CRZpk3Js24wI+U7dOmn1CnNMeKonJzDUfo3TgFCqUUMf
HgHyt44SDT/BQhYBbspFVWb+Ghr1IqoQUr+DNwaV5/ntEORUhob0DDM5XXshTP4P
P9bWQfe5DrECSYq8EcnbaCYRIxrJrWDM5d9n+KJIB6BrJARkf7EyFsy1uELiyuBV
opElT+qRSysidCDPcCNPVv7kKE7ctitCufAIjtftQXqPLy1eymMlnPeohbG86PR6
I+gOOI/FgEoH34gquqrP/vyA/x+Z9goKaxoIPDFo5AguFuk9gFg2k6NQtdzLzEB4
qYGjsodac+sC1jAQsiQn9x1YIDm2MT6r+ZiFHDuaqbnCwYvbVPU4SNJxnwecZfoG
+XJ3LoqBQ/kcc9zd5UTf6rRblg/oKA9RoxtIdGIMpn3ThAjUdX5Miw70y98U2lS/
68kge9Hvujqlq2+D5oQzH38r1BA1miCDMpOZc3V24+cnGwYmUhvCRi0rhcUGTNSV
NuFE1lf/elObsO2fFro3jZCoWwrD734XsDfUcLLmVU+f/1MQmJGFsmk5zDtULQy/
mH2jnqmVH2PH2evTtKuuEpAXwaxnXq9jVbF9bWz9uzyneG6z9hOvqiC7F/BbRt65
H7KjEKtEekuehxVhLW+3wSIRVhj6FJFtTtmM1sodBIzDy16ua2s/SBTa++zB92bU
2htq7f0SlpnSHmAdRra7v2UmeEdZ5v5Lfqmuz5fyCmUpPp7Wcr7IiD0dnsJ5fnYD
XVvXyZ6pOE2SrL4fOI5VXKqkQ/M865PM0BCTks/DnOzBxheONS2WZ0LljbXp0lDY
krH7HolGdM5USu0ohBsrcfYcPOp5+IE3GnPx+Xr/B572OkhJa8ic3lTnHZfV+sit
34dUWg264X2JuUjLgTZlys+9GoJtT3ZDOhKlPBi2KdL8bUIeribCMPAYYtd0bP4b
2QK463Y4dLcHGU9JqrYWZcM6w72PD86+pZA9YIfZCYAxmehYXJe1m5AvV6Nkc0Nj
6Wbb+x7JOofu1NWQkApFxOIKaq9d+IfmVTdCE2d45mSFmvLozRE/dccU6G/4JHxZ
aa3JfA9xapTDojx04Xbkl71RqUAThCxolvsqPKuoLXFWd+c/qFKtBWu9X1aeRfPa
CidJLC97RyVJlDtZwR5wY6s1sx/wZm3EYu3Yn5GmruLtGxqGnxKQxacZimOAaHmi
x8+E3gLY3p/CHFyL9tua88/FzKwuE/ypjByqmW9+Kco=
`protect END_PROTECTED
