`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
deyO99Iba0KtVacX/Pq/PUSqZJA6D8kKCwZK+jFUfx+g6mFVw8fYgKFjBkqLMNpx
HnbTOcr4ShJbZhgwDZYjHH7Wf9GBdm+hooJum9bBMOzoism6E1LGgUWP8AWZUNtU
NIil3yOpJcpjgQA1J/RRUNgedu+zWl6sO4qYQ170C8wc1C9DjN1k0lcuTOlUU2gp
WBkQGtJghz/oG4dJZ50ytcm7ZZK2QZWuFFVfZCWpEKgKUypO8WUUhBXsc9vD6shs
VKQnLW+8FILTwTiCa4DHEEETroxl0gisSASKdjmTqa9lNJuzZqQ8psyzvfWav1Bo
Qav8MgrANgoP4pDy9FEajNKwDTtlRaN+THwcGAb6NGHZvWPtNDTSiqVsdt1QReJ8
eiJfp6TPzQeqhRUGEdNVpw5f2XsboNPYsxgHti/kF0hk6ezy+Y3/XNRbexHtXuhD
m426uHnlm9MEfoWknoYJAbwvFyKjmdN8cs5Ti9IM+Eo=
`protect END_PROTECTED
