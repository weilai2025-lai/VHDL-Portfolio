`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1suCrijaTy5JdEuHdo+a+o9H3xkJbciZ3j6DbMWH06Blt/PEgkQcA44y+2ehYTw
oUAXpU2O0FvvPS7jGXUXTndBZCnRvxV8vW/TPhd7d+Jy1r+cEvScXJmf40LodRRr
FdlhT0wrkXF8NHHD85USxCd5k4phR85cfvRAyuZH3BGmuVLllkqKDPU0wLhbvbKo
sBHjt0PzNDlbDJnqVTuj59dxeQ5VPcNmDu+C2WsTsjG9dd8rW/b2gY4jD5u/H3Rr
SSZ00TJ/bWzfNnJOWQ+8nPvNrFFnNsow/sZIW5iL/uBUWvmv0vA6dMA84JGLPXEo
2ni6x9j4NMrr+TJqohouOIDEPJjdEeaG/XE1afzF/QeTKu3GMcCJxuzkaRXLMQxx
qWlHfE8Y8pWZVk7Jd8dT+/FRkwI5HDV76fOKYH/WyO4dXSmY3RAnf+S4jTGP5TGk
dWymlVRcCEiHpb+asTqPSWWuDTrC9mvqHKT5hMtntnS0rC0/EfmykxI5kJ5T+5r9
kPiAsE7D0ynr63f7B2+y1TKnhrfyNTj2HaK7dJmE9/mt1YvVrVS/yys4+qx6m4A4
sSA+y9yjXIlEVvCusJ86Z/t/Xu4qtQuTzZ0YrA3B+hauMu/wshBnOf2W3hlMs0dH
8ph5PxlL6knQs8Caw2dtN1lLf305JPA47JbnJmQjRXCXYZuFe5K6HBZoGKE3P8Dv
hBH1ORZNnIyAIEsQeTPgfmAh5LdJPPBFrBT1J/E0F50J4TTXVlJBwcBGIdQmqsyk
+sGMd4NLUdjWDqBnku6f7SrWiuZ2XDGVzCQ4BxMR9zLmmL3ZCdWoAcsQDQ8gC4iS
g/dvuZwh6eyVdX60sKNLsQIubF0wqNppQEBZIhaoiFvho2vzUHf36PHhRsPXl/S2
kNs7jTokNatJ02c+ZN9yghfVLXZtAKwpDHAZ6gbKSnH6P/HYkHKdG8XHVyOOZEzZ
t7vDt8a7FLjafMFsZFZvG5EoPKCRS4tOjhfvJ8tEKQlDqAEWrMcmlrQu7YSK1LPl
jt6XuQvtoSjvQjEUM4pvZMtFHqFe3qKG4PnWWA/HzXl6kziPWaUgzMY3e8QpcpBX
Y4UmtAMz+fCdAzNb63AGKPrybP4UMO5QI9nx5rhfEn9pjTvQm3yP1bkMXNy1i4gO
NfYvFAGUDj5k4E+Zt1cv2vfD+z+zj9xA8SzOzmrvGFGcs7BaEv/JaXNVK4Sj2Eex
VHWWPssUSTOOdSyOr4ND3jF6vBp31xiksTG9zMdMLNx1CljiwTdesJeqdMrD/xzw
C5qc9ezJp3VLW1xd3IAdXvj8mntqYNfeZWfSwzx2fcpigFyF9KkMpKQMD1MjA8zT
DZtWziEPS+frRB9qpzjoFsqVFpvJNkaVbcGPkS6cV+P8070zHpRaMuC6uaUyYavg
QZr0GIKeWfnR8/xYY0cB28kk5LinVOeTsmomLq+sLevoVTMZJHfqSN19hLhbrDqA
szXbkhL+Cm0lJHPNOK7L5xlNUN1UBKC2i/2WGSEvjPbePCHRv6jw7nR/dYmAduT3
zESg4qMUICdwe5AxSjZSpV8A09ZyeN0n0tIAsWGHPqGIAc4I7+DLt79VshZUaU2u
0Kv5fdDpwk0EAWVuG1AVUvZ/ivWW1yFMHVcgaCbIwSlzOtk49tuFeAi9yupy+lOE
b4Q8eFqN+rvx1804sG5elCa6HsAAEUYqnMeYd95wxwQGL9JZnEyUC2fE3Hj93jKE
JEwD22vwUubCAoRGEW/U5Q//VRPO4RE3UAi4m6tBKJFVPKX1FxMJzqaIFe7vWbGS
5Od2XGEzSpdSMDr81AEL48WE1kMow76DGz0XInvjv2/raXd7VTWExFp3q0S1jT+q
Bkfmx5zF2AIGpj/+R5x5eGCyWamKslzInzQTb1XA7LMqo/Znqf/uwcfvHG5i2a9E
4Bj5GlVVH4DpzvgIqwMJrCn/Uk/Csn4RE6jkGJoRXNIrQa9qqD8F77hPTVcvCBz5
vsrGqTQH7XSzQzOMp9KVEdGmCRot+cuB1E79/sv0lRyXQzqZMD/h3uHtdmNRJzt7
UjrYuGurOBaUJ7pkDAn7B/V+NxZWcKwUbaqxUJNeHu8MPCO1mv6MMtnuoWnATQa6
FVJcFkiMICG6Q+9Bro3Q1ojY0gUt1jARhDTN/UynRKWjpgwOwNl/yJ7eRvLsNXdd
JMgh/AzqxcbEuaDqCpRbcQtT6KX9UxUGFZTFB+MCJasIrVh6rtDpZbqcr6Z8w4vI
OjazVxUHE+V8SQaaqQlVNQmBHw5WpKrax9Nxx7Vn/3QEhQuZXKloYdZ03Q53u852
Mjn3l13aLVFh15n79Sdth+ZcEfRlqRbyUNPZliUekG3WSRuo2ROh5hHLHidCZDdS
QQ4JTVGS07iTF3mmcS5m4lAMC6PHhPYl5OKABfo3tRFioxCTOSwHQk0iuPaxGFDn
msTKV9M6Bm7YAiae6Dp8Ms0vVtg+XyPxRa7/xdDHov4IHlDaPkcIe0PgQmfJEioW
01bYuRyvI9F4mV9GGoJ0UCOQQ4rbxyX4JKClOlty9SkOP6qhSfax+VFGRzQBkCrY
zg6lDyq9/LG3A2flb6FAtzcUrlisQPA1B33rjfwcsAQ+MPhNacNA3MdeZXAax9aV
hGhd2xdYNfJUoHWKZucU/8KqfPl+R2RzKTvvjhP9ev6SyRsZQuD04c5m1jxA0ftF
GD7Njn3r03Kj+mLV0yxjhh5+vVYGzdPADkaEGowg2TuTtiNVSdkwIaL1eSxBGFu4
fihIaUSTiuEEJiVM79lxXDO38QzlIuYnElgsQ7AJVRu1EaKh+PctoIVIhob7bdSU
pzkoxjohYX8vadnc1idWYG03iHFLZxmhg3j4ezjQ04UCUum6NYMkUuoEn4Mj3Tmx
p7mqROuGiFE690L1on0ZEwSqN6qal8JBSc7Dgd+yNm2YZpB0KEffFUEGtj58wPgB
wZE6itXRdf4YibTvSR72Fa9vnn5wMnyGAavx3DHaFFONa4BCS+BcUJchI47pevev
js1Zfqjpz6vYy6DpstBcVUnN6byGqGAXx+Qp1Uv9XcMWcEodLdtYVvE9mIhYZML0
RU1U+qF/NG/0+XxfCLIJUHebfBMZZkmDyKcBB443EPcYtN6Pb79fGEtcVJb6SVsl
iRsLFsbPKRXx2WL3NmTQbpG7NU3Vj82tLGh5SJBgD9032Jv80xunrJXzEJQSYiLK
0z9hCNlMs44sPR01Mq+R8M8rHJKt4PzNpKk3OhOI9HIEu2BiQsBFkzzMX3/t2aPb
67512g+wJuIqQZeWXWZ+/Q==
`protect END_PROTECTED
