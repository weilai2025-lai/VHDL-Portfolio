`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZB688mtzBgevcFHIu51Ll6N5MPJFaVXZY480BeCRa0TNnuXxHaXBzjafNRWFQgKw
Vk5b3lQ1S+zRafDBhRGzNUQxuQZrSszq3V16pKL0TV1QFHo2LEShDN/jLZuj3V2V
Y4R4xoD+FNl/0niMEwSYkEEg2Uzf+xUGZATYBw9TJ68iTatIzNzIzxeviVISz/6T
/OM3CV4qqPYERKHj32BPXSueYJpBLO02giobB2JszrCDHfIipxXnLM7OD9lZ/6X8
gMTt+DmHM3EcPWkvd/vj4dq3HvERmY6VsfDGM8Lg64AVCW/GCQwKg1pdXgUypU+G
NWcZS83NcbkKB14S9y4xP1VsyCmekE68zNxdYMgKN62yOvTIC4Nak/DqEhFrJTe/
wB0EloSTVDoaq9meFESVG5Ht/EBygJeOVayU2PzSXfy21ULR622FGYb4IRRcTcE/
VngtE+4pYK1iMlnw0iITgDFqszEQXN66qX0y5y0jDXaa6En/ZRXK/hUmTkeoxAaK
uKsUFFPl2kRgBte9kFvMUZEAKHCBTsJ8ax9c8cYPtyU70sWgQwXfcND6qcMnX+2g
wwWkWyesnOA9dCg9QAYvLqNcCIFjdTnDBUFBGBOq9thzbXFWyOdzmyOnYMkTS9Ep
sCQtBKsu7Ztm98To5Y8rEvLOVcHDgFyrXwipxd8bYWTJlqr+T9P2O+HjrSK31dSI
HrAQCMeciUAtTzcvxWm9GPxkQC4WE26xjTQGc2Xxvuu6asY/SEFt/09YSNATHwh1
XOTeHbED9yPgH0CLpmpif02WNeEW/zfY9G4X+/uoh67P57CauYpK+bVZz3D4i0oV
IDoK+gkBHNnqChFHpb3eUMMVyWTQ5XNxtMIhox16Jnt76rGAiBYhwwZL3h61/ehs
xW4NFo6zXiS1QSjhezZ/eE27QRdOlCFD/VN9p/4HwR9aLtFfciQtjwyWF1uy0b5F
eFI4cgCYXhZM1mc5FIcXXnx0TmymkN6/OpsW5UZykEm4Ikf2eXz7T033YVILhu7I
IOR5xd8N/1woNsWZCoyVw95tpZmn34qOrO3aK9WxLXScCLQufNqDQVixaoZVi8iE
owbxnMEicXU27jQS25Y2Z3cH3d9QItypc6JpH6jh6G3wGCNEjrX+mo9EBw/VK1kB
R9AYMDRumU6amfZcOpQtBePGgoNN++WDSeT6jZU5nzuut4+itQeBrER/h2k+kXH2
rCcEjIgIlRDji0e5PYXWnWbO99UpQ1BqPDQU9FfJJ/7C5966XfMueHDLfAvX6QA/
`protect END_PROTECTED
