`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G50HThTNIUXcnYdvFGf18bmW2c4qh6ZXyz7sfPrJff1hKpjTtUFTzARwG9gcKvGd
kEIp8EK3lL0UOiqrOiABacfBFtyokXfyS7W1ypqzVNE/2Zt6O2up6op024CbAe1R
ij06OCCyflucMsVn4VodcHW4LBsiD0aQPBeApq03l3tA/pRURJBwZPd5zsKqEYjc
Mbre0rXFyVSRTfYYvxVTPcZm8faygthvtQFC8Caa1SVkU6CsWFPb7YovusweyLDn
n7iQ4l4Boa9pPOo7JLHOPlCw8sxpHdXBBMN1M8VsC9FeNJAOhcP+DmFumJ7B9nuY
y1434WRl9CfmLo2Eo7sP7v5Rj85WlWZwZlXF9ER82xFbyKbqyDGPo2l08WmQjdB5
gdEFnGg+3vVcvYDCuEDrJJKJpA9agMCJ21W7G5YN2qdN5yLXuzeNQbv87/GrFSvN
vty5XorKlpiXKFBnahZTegeBey4LcYsWUecDePeN1put6l+AH/P4MUcj46kk/Pp5
fqiK/X2ZgPl6MgQG5fmuNP9qka9OFNveqqzduTBZTYI+iW4tZsYduIzQALIPKwMv
nneo0g5vuVLoUOrl7oj1bSmJPPDsUXtosX/hw8wyYng9HUqNMpopWZW6L4Mba98Y
l+HojVLGm4xCfZ7DOv+SNcG/RCWvjLIA2LG9VO4EGfR3e/IgfWIl6Blap+czf/OD
13o3tO/YE+05iulVZ+VIseaIwUEFeSzH34DkKVCMIHaxKl2FgYcizePK0NY7jMFQ
z2oGyg1ozAkn9/MEy+pZcvxXatM2rLJxmgZg17m619Zv+Ah7r9/52xwaGv7HpEcB
r/Nvp6lwOriuXvwOicn0VoaktsVbEm87C36NC7Eo/c8ZbGalqp3JWWr72iz3ErtL
+Lx0ccwBGFA/3SYbxcSa3icXd29RjU+Lk19UMNti58TzzIB+Wzs9sx6FC+1WgWU/
szgJSQi/nNmz1hDGJ4GwFTzc6s0O94aEU5adQOl7jDuRzFN3B/B+5lXFkXm1I1Fg
GYWJkw/3qrZPN4RVvpzqwkQhAA1tiD2p+aglx1GghNPfdjJv94CL1DlSvtAzdoyw
FDdVq8y4Jv/wDpyNr0JFVx1DEuC4p6cb+uxi7c0u8ol0b1upYdRZv507ns0Is1XQ
lxEIm6T3hHGKBgESaNI3ubZV/inelsnT4hdzUWE49XbYEkRfTMYymcgag9kIMvuP
P5ku6iXrUeSBIQ8oLUYEJNhsw6adSxLOc/1+OaA1U6MGvDHXA+gzmQoSf6ICzcwt
gZdOfJMsX4qEFakdAol8abIhBQikeoHbV/FpSQTKc/ZtM5mWJ3llPZcTuXb6QcKB
VCWp4oH3FoUMrJ/NHg+Z2QNKMh0xqVcvy1VxZ6Pgi1ll+/D2KdxVaFMj+pua0v4E
MTY0NbGZ3hiZl5mhwkyROfAbFvvXR1odsGXCGliafxDc98mg7So9AFX99w5pcQ1P
c1uu9WkAGaFRWilVn0873NH600ZoFNSs7ZpZzFnp3/yDoems2jzRLTYwSOAFaKvd
d69JdEYZH7cYsqfLhmX1kE1Z+5DHr+ZjVnRjpWz93kpvaLir3/Ddt9jhLf71bkXg
kFwHKf8drIky6mHXf8gOrInmfhaFAVk72a/G/nR0lkbK7MoAtiVeL9FQrVyDR/Y+
oJv4w1wZs/emvdKTgEekU0NHkkUm+kvbX96K8Yf0/6fBXFEpnEZCgUt4iOZlWM6d
9y1VXwejNBub8mSudMN0nTyhn+73cih/bvy/XOZQwPw6mm8qVrABQGKeJmyOQLoE
fnoP++3lgDQVWLQTG5/N4b2L7zEC/ZmPly9LIJ9DFFO6PiE4YhsI3XD9G97yDVwj
E1MbhYSFceXJMwBOHYcKjDNQakrwmeOmI16o5/clKIH5+1EmaibSD9k3ENyVFAqw
ya2gl9NMJLny8x2peA6z757lNkb3Rwc+A4VSMr/EXs8t0d0fqfML7vlcZqN0mRNP
KAtEWAZ+eEpxDjISRpBVOcuKvYEPvfOO6+H+/1ciMOU4Gz5TLYInxnk4obN8igAC
iZ3/XWfIRCTYg+VzHsG4MDXSgmzW0uIjq+vMKFNM+cB2Jb/t0lIc3RObhIg21iJg
8IxIoqArKc15QDPt/sFS3Ut1r7vsp3z7D47KVnAtQTar/cPQfu5Tv51kcQ/HJHK6
JobnfDdNWGzr5lkR2P/grtdhUs6NHd+wfcmBt0paCl5Lrus/7+pZc6zvHk88oEiT
xLpZDIpeybOK0Y0dB8Mr8aXd8fXQl+3SbBC0/vNLfMQyIbes6pLic9RKAsouOG6X
kKY3NV1TUefB04F4p9DvCz5egEwFEn0iW2wX/GgNfSF8Qv/fI7mpvS2RQ9rruiBU
jdAX7iV2aLzuQH9n0wjTwh7/RzgbEpQdaTO799NJyWnOhUyYNt45/ycmRfSJnY3x
u9PRNKj2/+7BmLJH6wUWn4zbbwjUhHE9Vhz5DVmv+6Cb5zCYL/niWrQDqyC9b4dn
Uk6m3PJm7LgM/+qzdC+RIr6Cm1GDPQ+LTQEVV0v8FNAHpdM1BeC0diq7GzNkKvM+
GldIWRBOowxJe0mnV3+vhz8tFmcJadjzN+VRDAQKs434iaS4LMTwUgFpTK3U3pIJ
8KfllvD1GcrX8ELa6nxcClWMNVii10CKUFmlTPrV3bO0hWjKcRpDZIJnLdDt4K+J
3ieyovWEMuSoaS74uZVEtEhKdelC16OEHzRYtPHwV2Q93m+4IMUHr0sCK37iqA+8
gbVYPgSXSWyS9XflBR0RwKrGvqDv0BaT3RbYR4PXA6urMJJY0sPy3yE60XlUcWST
7NXKH7OE5dyW+odvkYVN/QIuaKiGpwpsTtdEJwu4swWwcBKj1m+/9fNbJlKfnT4U
nnzPpCtFa6tOz8WKAwCjfDYrhEvOM694ybDbZJJNEhNm4NsF1eDUxSvHVjf7zsUP
re4xY5jjsCKx79puLbRpOPzqCAM7Nikm8vMomYceB9EjY9nk1fVT/TA4zDe5AOTL
45AEy7ORZjI2SvkzZtj/SIXRpVrxKJ6aavrrwaVOUF6flAYUX9mPQrEoxkCa/1ep
dHTGc4wRbqUi/IVXXbbnBfaDDULn21cA62hcCeWQNoiWygQDuSuXopJEhCsJsmaP
DdJDkSSZ9E0a9sLbR/7p2H3ijHsnD2SobqKrxpYJcRl9qS5Sp/OnQBUhB12YXWel
Ro8qS2ySAFL35kKMY+ZVNXtMjwiOCqBpA+BEYtU7cPNvTyjIiLnNNV8Qy5dV+rbV
aVin8exPAZiu7nU5zHTWVok3wceNVdjued/RKoEhvYrraQ8pn1SY//39jmdFTKh9
UL2ZnkkRgkMI8Gir92UJ9Z2o77bQ7gmgkvgrMDOcoybuh51xBUNYYhprxQikc+SL
4D4sUw1zQ5l3SiUZz/aJvJtRB7bKFzGGtzCiQjfElBoWasoJ2M4hypgMBQSeq718
v/OdgYHpFqhlVmXOn6Qb5nK+OVVmmQ62WvjF+7raYRJ39pflZSAiaBvFT3YVukGb
3L6VYntxjiANXt1/OQLkpV/5NVkdq8WuWqKh6mHYjb6XVZ8mmA++SAmFyYeXzyCE
d7m8SPHwsc8a1IBlazak5tHRQYL/vYs7HUMXLpFLwL1nu6g1UtGrZZds5kAClSCE
BnztyFc25OZ4wr0M1wZOk6Xh9Q9CdeHh1A3iX0yrYvmv47sNA66aKSNuH6cC4uP5
/Jv9Wqt9ybXgw65JpDUN0A==
`protect END_PROTECTED
