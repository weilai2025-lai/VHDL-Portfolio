`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6mSaIJvVX9RsUgP/PjlSaEUVzI1Gw/H/fYKvr2iXlENnOEtzSdUg7eSUTXCNMupx
PNeLg+ENgEdJLLwvAAlayGSu/BJ4SyZkYhLSfDdF6i/IPm0k5B2M6gOWs+2dnUEr
qNurVSkvXBnDEFHTyR+xWxhIe9QxlK88fIkhXLq/VFMi4fkrLprt7+p1dCZ3T1zf
OXRdhVcRBVqsZo9MOadd1+6S2nSDBsbL5mBSj7YtZyyZTuIM550N6f19oLcM5Jai
coGOKpy6J3Yq9J0yiyZsWaMjovuTwaJEFl1VNztOJqMLOp9bqmVTMx6RimJWTnEF
8odtXD5mbwQLA2QeTPHPV/c/6I0lpchzkiG64AlpkVaHkB3wDIGYEzgdcfNlDDN8
UouQ+Orlu+3u1oNhFMCfUp6bQPVlrRCRxN3h7PnIdGeyaTVROWUp2R6+z6hyGJdP
12yWpRtKIy8AduqYTtaAHGQO6zgjnZt4/wHXLVal2zd/4/r1hw/ApmVZJRHKV67p
ZDlnI92mF9tnvh9SyAHMOv0au/x0etRzby8pwf25HYUgUC+dPPeRFD2TUjKqlmVb
RFgvD4CW45ZJzlgi8+dKxV0eWGwK+AlKaD9XKtdZmLBO24EChmDiNblnyiVFUL9c
JhNZAQJ7t4e+lOSlTSOqI3kRPiKeZpJXQ6hBZv9+zBXcvY9VxSIk0cI2HAngODeH
1EAICX3cI6JjdxLtF3PbKzGwjhwCy2DS+gQj8zL5I8YA+JK9Sj85S67X5FVeKkhu
2nOnAA+EhbCKK4oCkwXmmMX1mmW/BzzSy7sstZ/GUAQN/G3TNYDHItwO7R1IP1wM
Nsqe5JSWL0cNVxUpJINieMBjnGq7Bl8eOCD6z66xGgzGSJw97a4bNIrJShErIfE8
oWwvG0EkUJvi48THxOMg+sT3tdUe7uJaKN2Y3VcNsoU=
`protect END_PROTECTED
