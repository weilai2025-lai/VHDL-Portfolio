`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVh5CEme8JnRQLEwOZvnR01kdXkaLLznNRDoVTjmbNT28qs/35I4gIgh4tQ+Jmw6
3GQplG/C64R/2fBBaET8a9va2oWY39n4Vhx0uxOLpbdx6hfic7baqo4XpbArXxwI
MCjYZW4E/oJoe09mRfGCFrrPrnauMZKLM5tM4d6c1cKgCRqSQ5Trga4dM19/AtR8
Gag6O+A9Ts/7znecxVDLwGd33SbSYUEKQGfPCLDA7DsmUBUb3wXuMpmWVlGvGsx1
e/5HxG5WWSIJUfbgM8kONCvocLIqsovInzCTapgzFu9uyFSni4fUwg3VFl6LLUW3
L1zRgx9ela8uffxjpTBdEamzux4/DIZ6XL8dc8T2gdIYTkQM6vbJElgtmyELLOEh
IZzvYdNuFd58YT/u3wSW/gZEX8o2Xr+iXRKCHeGzL0H0g+OKxFl46y/ffST5t1nb
BREFMxxNQmIrcepeqKV3ek8kYLw7JRMD62aZlSoZ9tNqNJ3hMfPUUdlqV1n6DjFc
Y4Kxl9D6M3B+TCzbaQPS4UvSR8G1naXTiFUPSrEQhyKt13Wdc1m1zm9C22tp4p1M
cSR4az0AlzpZnhyeiqpuUpWADLAWduI6bbmtYbeG2dzgFvTI3tOa04pKCmRkjX8m
Z7hDscvsvnzXJwA40MYXRiG65l+Fc64Hc5rZ8vTAlMmDr4On8L3A29X5QVWPK5W7
QD1WZEY+a6TLsZAj/DAIoiALW91Uxzpe1yxE2CNoikzZc8poZ29nhyk9n72uzARn
Ybxhru+q/RTruAvFgnGfeVrO/izI7NVMuNjKqv7UrPknQBBv+6TeXUUlyCHoJXT7
0D7yzoHH+MaTClwUcmylD++zPflweWZUmbo9EkKVWNuTDR9xP5rpeeWwC9dYOvq2
t0z8512MwFAPi/7OrIdzjJmVO8Es9378SGXcvpcPiXhhYtwvyEhRlVLNk2u8BZ6O
XpJ9f9ucm5DEjjM+hYjAcou95vhEYDrLLezNR/C+NGfx8dwDIRRx9Bu3rg/3IV75
7MXSwXC+W6Dyh1lzKozI1uY7xiiiNwOM23dwmL5V0DwC+VPQxr4Moghcdl26czj8
QKJJDGKFHknI/TbPACkrwDEIgZMC7afi48B+pRyl3ipYngVsIvfQzCUWNQI9t+vm
NQsgOsjAM77Z9nw6J27Cpp0QagxHki/NDFyb3Dqpgvoq31BIJWFffdVblz7+267c
HREshPHdaPXFBFRjjCIzrTvM4BxsZbYsDBDR8NGVknt7mWXDED0jggzpVz5I4+/Q
lkmVD1bpLPB0KncowzOeitQGdsjuJ7L9c48j1/VS9S3NjEY6ZNHFrWM3s28iQHJR
e3AInePvXnSB5Dg7s94BiAqjRE9hpSpGPDTfK91geXGw3CmpxVFZCRxQYIMQpthj
s3BU63YIPqxfYh3P/aZRrC2edR8SroaqWZtJcAmYQckU3psMnx+Rg9HbQJW8TRkg
vqzYNUYhYE9z91k56MnEXG2bLFFkrGm+M5s2U+6iPgAhICHiUCOGyFjKevpt4MAy
KzdNmdZumejjUg33ADGfyv9knAeFPM+MBjWt++0oWdqH4JvKGLifzjPjHIbi9/S0
iMTmgLMYlr/0lmJkOK5iILizaFy3jeTfjXUlvqoCEuTGMTvdbdrmzIJGnE2SCKHq
`protect END_PROTECTED
