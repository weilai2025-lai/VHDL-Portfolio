`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLm2jFLkZXeZUSVC6wIceFIPnz2M1gc+qZQd8LsViI8xmaOjELiNxEZE+rtP4AOZ
bAYoVTjTmvimGFM7DL0RIWowPjYfogADlI9efhxeyPqJQoc4XIx8ThNXx71iUoqd
cO+k9xETTCPflHd/dVTpR9bld1Mo3+Ho79sA/YFlBL1kJBfXZMQr+4gZh9YUQVYe
0c5N6O0TzZB07Ai0ETArjVK2cfZT06p64lXk1GcUN6h5Omkkz9wcYRlAxoKVLfFX
HlBq30CgJTnrrQJ+AexEXx1LKH4E+LagtShWITQe+j1c8j30j8zv9uY4T6fTZw3W
cvCieNJ5ewddeyIsRnScu3MOnvbMsp1JEZLRT8Pt5ynuACTz0q/B/vBcNVaX8u3y
2wQ9gvFEmZ2hfWX3MZDyC7rvMMBxmgMz4rEt9GN6XOqXOrj7dwMPdeWrFvhqdyZS
MsaQNYTbmQlpxplKQb061uE9omAzsDP3Oj+6rSz7V8WT+trnCtwxEaEbGX6lUGZe
vNIe7LDC0+DUlYCOfBXti+3cKBhC4qzVIe3wC3r4QHf1Rb2VN6/9XBSVDQkuCvQJ
F1YDw0sRBXr74IsSCeCbi6e64LqN0AYI4n9gKLfGtG12nj3OmARkxqKfrwBoayXY
mL2Drpq73zT4F043zE3P9M4vnTlFlJPmTs9n3OJgklE/nSuhVTw+VlduT7aHvybS
aBSMKn4kUHIp4VBuXKo/sZMmrazQV0hoCdkbnlil9LC/mCsew22NG0DNzxiRKc8l
aeLxrDG35UvlzJ85WhbnXEiBbNpjuX7/IReUXaBmUWFtfi/AMSId6Vt432EDA5bL
42cVSnHIC+y864crErY48KvCKeEHpSg9egwAbmM4G5lOipimzkXxLJhIVbdbit8w
wTLEmwShe2U79O+nsuNFQzCWyHuQH5CaZtRI3xOW6kzWbTrbjP1BfKw66ZAMeppd
FFuNwYOPYx8kvA9DYJfnJTNWzmBYzCRF4ANl/xf9fMszSZxjpuYB1W9QtaPHtnhM
V23EEytu/CwJk87xXvVIwFcETMXqXFGjpOVTKzGApLj3XTPpQQ/b/FJobUiLcBf2
zt5botyy77N/3KijaEhG8mj7r63TV848ct+YreQFFnFDpMmW0OKsayEKWdjOm8n/
7ld9uvFHT7lRAYhcSiab/josIcIF4+3+zkb8bMQfSaTOJnsT5nRWPcKHRVRIpfsy
I2yqQ9inoYvsdoCOSg8WclGC5mNff56//65w4m9cv9QAwjoOJiHWouyHLHn5gCIe
`protect END_PROTECTED
