`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mju+lduYHLk74cCA1KAC++EqmmH+uAt2tXz0Rfvt6Pg7B2lusCo4LH9ZT2YTlhof
d9F+VH6XQ+WJMFDMeP28jBp1y9dD/fzAfeZOlXUglRTDYNGV0oeMdo5Okh8ULxIK
dzxCTzFVFL/Lyh1VIb6LmwvSslV9q5Tk96ktwS3JgBL+QgTG1n6rRqdMPCxS8WjO
Y6x7eHOiaSTX5RWFlLr8LpXQ07XiOMe7XibEnXW6sopxsmL3VUpuRkJuckD1fk2m
MVaW3byiEheuxrYCWfbNaOCF7QrT2uAI887wDwTnoAngV4DApvAVlF7gkdxcpYIs
dPEwIIbkCcVk7lMMfl3mQnkHlMc0Pxg8KuLkJVyL8dFhZOZoB65jhrwT9U2p940P
HVAYLo7B+XVcyZi46vfooUpHOiWS4E6aygmjSJqa2HWjGzhPYYs52L38l81hGGot
t4wgTKiPPsnJGVR64lJZf96zP+2E/83Sl2lY+7q5TR8sFNN6u7nq+7NmsLzu3M9q
yemAZm4wg7+XyMV+tIFcY992u2hDdhtkdQsUDUN5tJk7zNgW3JH7E6m45G3eC9L9
FD+ogEY+sNKg7NgyC/8OATXpLmQSoK/It0bCnhF9ABjvDCbWeH5F/BZgceEfNDSl
gPZXscZCkhDPBs5CvPSChbpJWLoq65Wkq/yX/ZTXodcvZ2BfhyaHM3+XSjr7AZLh
J+mCWSKARZGsAYFdV4gTh0IQLgGZnG5ZFqMXd/xCujXxrEaLjGKlf2iyUZimXLDe
2iDv9Dg2ZdhMRyMkYaY4R83LHShJuJ/m+rKNcg9+W4rHMCohGNyLWpibckOXgCyb
L9sblkzcT4IbP9Z8M4uK9WTArBv7yNITzaFNianMmN5KGUydQCwlGO7XD/6//A1P
sweK9Pg2Vki5yjqujwj6moeE+R63bgJe+xljGUch3HGTl+pKB74JtMwda8RAu+ju
V2cPxTgxYGZ20QAK/T9mt69H/u0XWISefVIzVHA9XY2agpRO8L5qCSdwdvegx25X
XDGjmDTfmmGJbiRRu4DBLGoImnSrW4FdvwSBFYoaYvBtwYW5XPtAINwkdtrn/St5
Lc5cZr0nma/VkNdgJQk6+7V8sK+cZpdtLU7fh8lN3KG6SPw/rZpmupZ5nbBTq9cy
8wqrMs0xxVPWHVSr2BOBjyMFSBZarWynrDQSBb9SWNNPdIJppHtTuZUunLDEw0+n
yeonoOVXtFernISNSeJgfYbMxs01t5FKFwqtNGWUm9Sm1Poo2nSGQbg619KvNAVF
8E42CPruU2J6KxZNpEs9XACC08ItPkFS8yRz6ygNC4JXj8NnQSKwDcuX/uSVsjGT
PqdfrAs2Ly1+iCejFM8m/HNJWX2XTM2CfNvMWcZPJdWJGs1c/vUfx/YaeRh4dspk
AkD1bg08oTFtG6XNvYXaatKpL2cfKR2f7sSW2+SF1bk5ZS8+iZYYJx86qPC76aFm
eijzt95uefrlieDC61KMWD3iK+1IbpYPa6asXDEXmVhrDttsFgxVSBTO0WbzLy6p
8RnVuMn9mL5ccgiwvecXvkQ9R4nMRxg2fcihdhsxFw+79NyFRmWlBm34sBLCqWqt
YzyLU+xjPhiJEdGFA3tImh+XZSVGwxi5cXu4mPXY6vk9R9Eq4IDp2Y/qFeNeVG65
26hQ3yFjJuxxAQrESRJqR9TyDk2Y1hj3kixwp7HpQDPZ09RMNOUsjO9AF3caTgGz
28ADv0TGL9lDc4eUa6neW+A3DXpBtGpfEF0aUHsWH3E/2/SNtcHjNTM1R6icUOGE
J+2hDgUDLkCokYsq+Kev+Gwwq/2A0X92r0BRg25otoqdtROLDKwl7cl4FXVQhj2E
1prWyZb/1EKU+tf2cM9KMbiCvhK/XW/xn8kNxOTxZLaRx49LyXj1+no3ejVHZLtB
seu3YHpK6kREVT2AyqeRfA==
`protect END_PROTECTED
