`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Qx89mvoA9qs3epks33LdqLxGSNOjBIBgLG9gI3MwlNOZHrQ5U6bN+q0WxPK1Toh
14DM1pvDWEUrljf7hzzWC7RhAPyKMkEYx+0ebMsbggUQKkpj/rv0ZTvodP6iyr+H
1GepRBywDVbn4tJFfBfCr8sOZa5AlgW7imqRjumeoOBpw3lCYPKoyvfnqdvNi0D+
f51TlsX4Sa8IYGef216ePRAUnnKnWlNhz7GFsxW4ehXY7EQzKpt68N+RRgsHkbj/
/u35M8aMrsTmKAQN9Aul5V2ZM1LNl4mnn8hZYW9lcoahVo1CmxDBnuw8+KtbZ55e
2Z30KFZ4Vky0e52b7LosyHs5MdUHd68pTQoKArK4GBulKLX5+quCpr1xhd9tdqkw
3xI8DkKhcnfwxzqsYpiAhoVrP3q69AEvlgzPwljeAjYcV/MHX5AUQJIwjctOVv85
7uVyUQogqozMP8/zzFZimZIhxs0UYhNiDjVUqIW9Dd4BzHN2nGazp+btzRv8gvka
2giEqGZidL42409b0CuMpYT4aeRFbt+Ph23fw2A5g5dgpNZPiGiaK2myNC+NTQN6
disbzm76fjggPfZk4h4MH5zRkr5qfXQzeIf0LsVoQymSLNHyU9LFAnMvd1icW0Iy
fN5fIRsAci7qUyRmI8ln8PRr7Cp+eusDXa8ONdGFYcQ2ZWqV5auA7goecNruTJXw
mMAaYrYOsa2bAyhk48J1goElg0AmL1Kh5xLqo15LR20j3VZ6ZDUBFU+mY1NzsQnD
cI+qgoJjjSXhFj1GyAaJErgIuYDkqlXupfAlM2Hc1JSccAzHSH0nDzX+WheylGKA
3olAB9lAJmles/YzaoQDOJdLg4VKiNjad6uxk7LkqqQlwSAUjD5iuvbij3jEOsDr
yPKShpuY4+d2bZ/W7C2uLvTRq7UgiFwpr6JY24y2KUNYesJZcJrqQ9RuA4O4JIaW
pKnImBSU4Sl4l/ISTMwHOVvDpP7gZoGRYL1UNcVh7tQzqsC1Flqzcl4koRY9eLcs
GE4FEZ12ZXTO2h7v18mWdop/eXDNPpJcrawC4/8/cunAB49zKKHEQm2EfaJEkEl1
AdABQAin05+6GB4y+xdMvszG2CXMnQ+sC0qDZLtQaT+8cjVlIevBEFgZ+Q9EQBna
BFtvun+WccoH+YVTRK50bisIySlDOJ/gq0cNQ1DMptrSNdrz0k/8xOweej0aCibD
em/6N+0BMXqvMS3F5E4S5UGvlf9AhTkkU6XjQxM9Tg4JqazKldeizSC9vWnyIovi
i7YZ74x5CCObHtuD6yOysUNFTOJe/4aohi9ZKnPPaMJtDxB6Qo3MKkaEElvhkq16
rDmarZMXDwNRkF3PUZI2sK3rx9tsYOLkN8WrGTF8d8j+ECchjCiHuKB313CJznMh
vRtrtYknLmUbhMUGC8S/H5gV+zzSN/gO5sJ1bs2JzqPXPDOf8mnje2Td79aYyv/C
S28IwtDqscMmjI4h4J4JGLk9qZVbr8jX+n8F3du9Nyc=
`protect END_PROTECTED
