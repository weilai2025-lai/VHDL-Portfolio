`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3HeuX5KvoWfWYa7k85HpJdW83IH40XlHFGpbvsEPYN7MMfN5ka65dl+r4E4x9IjM
yf+VYLi3ADYs1nQCJQjfIZRIPzA0A2tiGJUyQ1oyv/wYy8oviOs1Z5LBxjZon7Uh
UomtHS4shegktF/jWWzwRYs8aHua+xgyxhnAiEln3OyiKfJK1NIEC6xaxUkSO4BQ
tkph2jzaf8Ii7BY6oC6fQ5+MoGA4o+XfmN0SdfMWLWrxytXlNKHY9K4ZKgxWAHGC
q53gIR/1yLzQPKVwu2w1K47ep7Pr4V8OMbgsKTbJbFxecuJxdbyUfzwm/AlI48iU
K8GieU9wNw3GoU+Fkymo5cpse+lamHZCL2BG6U+RAT5jml5X2Z8TL8DIgRtzwfO7
0sJnW5YY8MBPykBHF+sJd+3HFYg8XZOtzgvpRhSOFO5X1fXx3FDpY2lCYNdLdX/0
XDV1JU61JMZGIZ1CGGdOt8m+tuNv9ZMCtcOXU+hjMHwspmns3CCBUKZ+gGOeijm7
WNnI9fEMU0howXn7whpLrgk8M6YPmlyzf7WhFde1YzvXLjZJqJetIiOZ0WSGeq8r
Z8V0lF/iH31Sy0i+JGl8xZYq23OYIg4cR6NEIVdkay+7S78Un+UH4DkZrW6dtNp+
bjw6RrZd9NwIXSDQkY6rzJ425zMnfeuK20o+J57V6Hk=
`protect END_PROTECTED
