`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0bmV57yX1p6tasiimBl55KJkjvH7b3HXZKO+lWLgitjRA8VQcDd9DOzwWfj8rga
uSvxW2+NH+EVZdxkZzm1TTlyEaLQdlvE8i1pHgTj1UIC9ntBNcwUDjMsyGs8RBWl
wni2caUHTVsXZ/gluBIschoiK0J4kdQVinwuaqRgNvouD8h+WNQwiHsJ8S2hE9VS
qH4mnCUT3H6fk/DxXrF7AX/1TJ6Xk8nuX2+M5PHGAnB9Zo2hmt1QNkD8E07oGgFl
GabiSlC2vO7WlVOMzOnnVXgOOTbHWLwr6VYUx///UR9wNXY0p007ZCm81Lx+9u7a
fmDdVH808nPExRjlPEf8UXrY3UjWO9Fp297C9xFgRH0kicKBAK/BVF1uz9aCAeCR
nZywBIT7T89VfoRNE2XRK+RbJEproFR/riVis687daU=
`protect END_PROTECTED
