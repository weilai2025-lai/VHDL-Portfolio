`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RWT7aWelGxAHfyrqnyP0Q6/TL2lpYoZ56Jx8lWVYsRgiCFoUDuUZ+HUNN7CsCJO
TNKyecediKvQDJ+nJJlb6LUUCl37CZZykATetqU8CH0VIgBuQDENLaawTyY7u2Y3
RD9WwdZiT0d8eUDVF5I8mli9cYgevyuH8akcIkxurv+9tNVX3U2/MkoZWfo1WY8X
Zz9+4Ij9HODaj77mqkIpvi/oTbCwB552cwz7R9SmVkqw0gr3FYBPlZ8DQ8dlTXtg
E+361skuElr5K791le5WdTsxMda8VRPXQkW5za8F1ibUK+kOwqx4EqYb74kM8mon
xZSRKTcBH3gTDToLUAlHo7LpzJlLCi7ATOGZLUm8Ym9v2eYBW6WTXDKmQLEG2P+S
1Wv84qh6XHR5GW4oO3BHgM4LjKC6NiBRWuaPDFJXLHxuj3PFeRT3m6PIaVNGfLvB
M4FtBITLRdLhpu6DwTOBjrfiyqv1olTgt9hYGaDfI9WE5bFJ3gUuM501T71eZC6J
6Z8qwjDAtYsjMlCgFVlgbbgVwMXxUXycRD7nW5hkUsMVzZVpQnHMfPXmrDChREPP
76cIQxO7YciL/kMk24RBIwn5L81Qo+RDomfqphlRcXcU4yt1a/mA7fn3m1mbtWpb
c7he+PhUkxjv3LbhvmYKSokcMAHzLy5bnj2X5m8w4ggGAk67q2CWtJYT9+5kBxSY
0gtxznDaJnYa9XMUMWSYavxOykBKsu10K+YbhOYg2VADDtW0P4Bx04ie2tutRroO
GjxjmDgHRFdT2u6aaF3Tk1KmzwJm9x4XVbdlFSLW4kmNl/adY1potfbcPUUfaV6J
/aCWhWWi022Oi8+FNY+GReYQTv/o3pLqNCpBUVquQCsfmkAZaNDh/6js1Z5ez3Jl
rAG96Z1nvUnmX+StRDKPNsfWggSqcxxgJ3ysmTEuxEVF8Mf282FSjiIL53QGZ2b/
k1gY/v8F1J7dxsC7vDhXfgDmW2hmZTybnN7Lly+m8/lMjV/W/bkHw0ArDiac6llq
Mm3PaSS1XA+s26BqRUHXpUj3m2IIAsZ0wQTXMMAm0EYE7GFVo/LIpeSlIDyNnHlW
Vgwx1Qvj4zoX/m1RglMo8DGeKmNgUkiqKpP0/DGqe2TdeBttKamFSPZF2tlPTmZH
VLWNpJe5WK/o/an/rHAiJsNnh4WfPBOI46XHM0cUh7+R14np3lw5YKU5EM6fk++3
SwfY8q3YCczSjROv4S4qn85WIOe69s9/bfR2TJ/JZ5yNm0Y1jqHgs/wdabk3UwEY
lplIlE9rKqb2Ol+dhZ2u4zIIUxOGpUyW291hH1DqAMAGD7VUu0iR9Tt1lw/kVqvM
rjnmoVFcE5Auw+SnyjeTpv+bvTGSrIHfZFD5w3rab2xcoeLbYhept9Mz7DEHA9LC
P6NlqI6facELsw4j/S9k4pr/Qh7X2LwWVNq3/QZ7gfI4zYdRJ2q5fEjvdjDJEh8v
uWvl81rJ8W5UV0JFzp2+RwJ0LsekhLuxbm5bHzU5x65Iuo24vvMX9c+pqs93e8U1
AZeWwgEHEKW/ZHEkhTcz8uVb4iPzXZLWIaM+zd1YU2v55/ilRmJ02ldgx9bzG19q
ICMY6qmC3KMb3SSpobarVSI/82TScOb68fr26wHm1768cHffnMa8N703fYkguWR0
BcTZ0H6xxRYaIxTosZvqmEaPbM26zeFb3dqVY0HQBBUDUE1FGgyZfLNk0Vww7xUY
2c1gvGvdIZKLK0KpFRaPZahJMJvQjR94VIg/D8sNtUvGhg/FH5kkQwK4fHQvFrsR
S6ECCd4uRuymvYXgoGJflsMBp+7liyV0GtLmt0R4ufD2OeNDPIj2W47PNgWw56wc
yCodWvhg77pkOxhlQYlKeTemp6OgvhKMCoWMrPJZi4FgKVE+wOMsE0+U4Nv6yxTL
pbAyhfwCxQU9nXFuhvW9X+fESXl5BxjAI2xV0TudcUxF1EA/mjc2wrboFBSmEhkQ
90arLeA+5JHRB3ozm4Vz1/7GwAw8NZoJpyJodg/KC7YNEXA/0CMxkAPxweREPNDv
7tDTplVs4tZfBnW0/RZw/s+n6SVQmqwPLxZ0D+wMKmbxpsjSxJtnIaXm7E51dd/7
+MIoY4fPv3oP4ZeM4WGYSIYL1cweuwyp1SVWZzMw9zqy1tkhCWEc7UdZeTDN93C1
cGmC+TEmWWeXLTcT1MM2eatw3N26DugEoQrPwLXHpHohhEj2YRmOb/0aBBTnW/Dn
nWXlwS4Ys/7nuyQyUQFt4KVqhRigumWW3kYOzj9uxvCVoqQzuKGJwFDe//0c4kCU
Ifa+oO7Q8e72WLyf+dJI+5+X/AFRGJxp9lxk5LH1BJ05ZddTugjb3y7ejxJmjuhq
rJAO2C2FbiD1pxylqTK/wcwDahCGLZ+ABGOXM0BDtB4btyG2m7EmjF/uLyyIHisW
iELp3BpnNcozUPmCkXW07+RveoS8i2PnvaC4SekOrsARj0L8UG8h4GVg19jEkm4w
B4QbpMdlghqn5hFtkgI7cNw/PLlcE79ORGFjZWuQD4cf1wVq3ZlWxwwl+mcFj9UP
Ee0JZNdSmuURZCGP3snNSifviJC/b4GlTusvcyxekFc3TogpfM3nuDanBmhZiEBI
/4CIuL6eqtp+lL5n7YPucc7VMUFvQ1hzrfncFyKRtYWtraRND7W53kyRRuaiUIC3
hA3yVeu1YsBp9I0wgbtXblT2yIabLqDawpmQLfgyQJodl95tqAqtKEc2GoYhARM3
p+8HQmHcnleRjcUtnyPsvXJOFEz/WEVDVMOckSbP9JO6n6nRM99eLyptXDuyatKJ
3TOog2zAxbNR0O2qtM/LzueVLTuSQkIFoVKPqWq9T1Vo6f1zcJREbKJefVdrO64Q
LYUaW3KxAItnx/TQfQy+tVDhr/TWW9xNAcc3qOxeEEgIS3W3mo/k4OagM79ObElx
KUEn/SUyy8GvdA//F2VXMSGsVxNnfn/xCOvuIeapS8ArGiADTJQv3towRSXFUMsV
G2MoTZA1AcpdeaFndf6HxixXgI+4dGeFCan5qKGHFZ083jTKYUaL/mar1pwokqra
VHLfCgh5duSNTiKaTPQ2zwAJ+R5sEGHcYzj4QXvENwbtYK3pQZAk0DckIUqm5C7x
1CNlXZpc0MJ2db+kBesbSyc3F7nBGDmUX0Scxl3s/exr9mQDLwgHg0PtZqacPfy2
KOFiIp/AtI8DqA+KEqorULV9ZyXr6QkOviEfH8ZMz08lpgjlpzCzSVI+cS83ySC2
Y6D+AW89XmNxiXpsghIL8pGM3SSNtR8v5n5mcR5qIQ48XNpD3xupmHtWuUfP89J2
K1m8/iddtZtnB4O0BmjR6t9qfZ1fbeXRPXmG4liIdStlBxkvKIHwjDIvx5oB5y9F
2aUfkBnuLwUdnuB9/tBibS+u5cvLwJ+kYp3UHaqT9J1nT2P9NRJhv/uwtg/XF5i2
fVlmcRZuFmA4z4/P9/y/XHSQBjf05Ux3eM0THucpNBbG+NuRZW//bn5pK8GUPYVA
IMupAZxM2EnpLHd1kg6mwrP13peSiqewiaPqCFIHTOdFYcJ6hjxwYNaRWRkqAYLN
Ih0dybdvkX2dopdzlokylaPc6mT/70ytsWBh46YN4mDwdCo/NBosF+PjEp0sfzdQ
UQeBmJWwUlhA5eN4NmLBzJ1KxrYCZdE4vJst4P79aHG+O/3yAyR4nfGV8eXHRZiP
SC7Js+Titvw3oZlwvD6gkw291/PnacVAZIFGz7R2REKVbGZCgPGlBGnnrbiYSc66
uXNY4CVhulD5iV3i37XiGdMGYxNXW4EUUxV/XCC8Y5GenfdfLknONI4blyLdhWKV
yv2MKgh9XqXIuyfWiZ2Y6SnuhfNgQHKLV7kpyl1pq8O7GTLzpjVCjw/lCpUkED50
lcEkG75YBDkWIEDeazf6PnqlkTmfigyLHqHFiQd5PUpveB08SVuVfjODG6W2WkwQ
IW8FwDaooKzr13J9j0r8lnbnwe1aEjpcf7T7oSjPR45XSvkxfC8IuMslVif9FaKs
cBVvw5s9BMEHo41SDCxi7xGz2SKAnraXRBtu9C1M3brTt55GijCyD6bqY1xi82Ex
2Ee92LNzs/vwIklqGV58Kd4mKgqCEHRHrQrCEjv8AiNl+s7edjWZueLro8ZKmWX3
0MKwHg8TbFjnis3WgKxUDzoUEwFGhepJFKFHr6mUFNPFptXKiRrWk6wTsVomQi8W
6ipcCjda534yznmNvX4x/2Ubp8MThQcUmaAolce/QE/5tCmjWFs9ePiWrJu75OPa
QcvsUo2tdtaI+oKY937k1EkOZIlVKZniG4i9G80FgJe3nMsnqgBnCbOQWQfV76zU
yDVMoDofINZZVqjUsSRhnYr6kd/Lelk12mrr05VwefLVzG6oEtVTHAg+5GwyVcM+
0F+83ZNbVHHQY6/AHhDnMcZASrA7nzdEcyJ7Nu+fXJk3YeF9G/Vqd+Jgnq9HChWn
VVSbvXcWafxEiE4gK2DXQsuun8DdtLKjlqweLAEAp9MBuKYyJ2JwB46oJ/jExkpg
XS9LfEFuAHj+8exq1P9ZiJr3pwW/ZYTuxxVUFhYu1nfEN5qB1ut/+fjTW0qu8VDG
W37/UP05OBNfKrHEoZ6JFZr06/Y0dTuQt1AmZgFDIa96Hst12AQOwkUXXh8VeXni
G1n93Es4EscQO40K8s2pqRCwOxHADZ94tMecZjWamjAEQ0QWGKR9yKiu++7AB9fH
FwqGTMg6yza1Mt7QU0vhAtB5+1sBGy9bv4RLTzdMb7F27Ea71+i9hqLMY2wNIIri
J3sdl+jBk2pll2nidsqFdOFq8bxU0M6Px9m48EUpnIz9k5MYDhh9sYMfYH/I7J5K
vXC0xIMdQSiR5oQGFbPdS9XJrT13W8ThjXp8DF4mt/+2PmDVF5p1F0+PMXuoJBgM
yWHQXakjWgB4tp1kpVl3OU4igdCkRnTojfELroVM1jAwlgenIpRuPkp6n2xdAhSN
cXBXV6RRpbl7oNV6E/CD4hiQx0zA2XWCSkOpD9cyKqHvuJoysiBhXHDMySbPvI6m
ADSOvYCU9+liG9DaBRGnJLRxDucj2yg631ZHE5Ha4DkNLcs1uuveBNjddvowRjpQ
lBIdJJKF8owB/D1ZMgrzU1L0/cTyh3Vr9KAoVqXMeWXyOCej54XXE7A5unyiyRse
D4rF0WRGGstiomiECIFj4u7GptzDs/splt80/T88LNYVGMEfRw1F8+Bsr4tDxCsh
rk5d/RDZ9W5DZyNxV/5xhUYXQz871OsYg5EGUnPuNt/5osolv92mQBSZ3lqLvWUu
PIL0UkH3rmXvwiX5PSb43fqwAtJ+ObFwdnJ9A5C1ur4hWAxige6mmNtOyAETSzqq
1WJlMLxFGuLJyfbHnlLw+JRkMnWIvCvJK1m/cwQIoRRkCt01CSHA6anSYIuqSE/+
kyPiBbJRyk4inDBD3RkYWK3jEJ8ne61fe7/VuzIsKa3GSGHhgHZmeEz2CEZ5T0Uc
CqYnISpkUUXlmmPFsb33aDjpe/CdGF1Un5xdmDXTIp5H9C6FepyFupdfBnw6XM4w
iUOPJYHBkp26g8fIxXjOKfAlBV73QzGoJFLColh0yv8JBaerkn6iiW62T2e5JHXN
1m63qUtbAe1ji9C4R2exnRn2M4Lj2aqo3P3LNWyMNo6V4djlbdiwLS+kjEbL38Io
4LA41hAc9j08KvpUvSv+NPrvRUbTLPiLtuzsOBLZlnWlrsN9YPjRAPseyFK6C2rq
34dJWi/KR9Vdo7Bn47g0Z2yUphHr7Uba6DCP9PbT2yfB6D13YizeJkpPwQubdbk6
m5G8sSyARw0WbR41dYOw8QPVhBkyvca0wjyoWroNWwpKVxmETkJz2UihDsjVlag3
d4g1cnz9Cjz62iH1lWm2e1jY4leklpPzQsepJHjiKoI4YmunBDHW8K7bPks1VNjf
8plY4CWZUMmNyKGB94BxlgsAdsUfxqMucOmqn9kWDSdHQatpfrwbglpKY+jXQNSi
yh/G1pHiGtUgFKvXyj905qEgtS0gsW0+rgahgPSCsXaUQoTAAhrqco2gGTbMIG5R
n/eLm5cJosbi4M7NVvHhLifHVpx/t1zXc0YIYEjdZzwy8DaK3hNnz0HiksxxuS4C
KxWFIEPRukevuanjcFRrD/SEX8J30nRceynknFXuuLI5nHXMa3oh4RFMa2Ucbf83
wxUj2DCWsyxiQJ5YkjdvuEAIxof2a3Cc9gi+aSuvjT3Z/l4MsjfnO1s9plAMRnyK
kCLtltaPIOuTrG6PUUHXzFPdw/i27IDYibMdsaLYNR5Bv8UzGOSCNNa3GfEVJiml
9FqnZ6FL05zvmesxGVHB42vjYB1/nNJZySC7jap8Q9TlgaaMiqIvvd8Svxy5JbN6
UCDl34gxlFvZHpgLQgqoOn0PkU6GKkkYp1qB1lx4frC/QMVCkNbblrHtRvPwEJ9d
1DXNGxwkbGIWfGmmy0QwXYEeJCPXePzZcRIechdhcDoPYCs5NDZOTrqgNZP+Ng4d
XlZO0GrNPT9GgoIf1x7RWJBa9nTYPz+Ucb4uEP3z8wsn6MX9E1QeBfpdw1StNICm
7hDNdWKAo55BRYt114wehTsTKcrem9tMrZv9FQrW05KA3tcBOkjsUrYZ/bqycU3W
KScKjMEtB9SFSIdNfP4su2q/O0IuLMDqQkFg584Q92GMykCT72JlQjzkNDAOt/td
2EvZIj4hajGNjXPoCHGnQ8u75GIU+0Zl4skFKITSnR6J9Ts9q9jOlaYMutYqH6QQ
bIqjiRlwppZWB1asQ5lXXJDcyCnjNB4HvJY9hPbFZ9N7PimhBRhZn8gtlkP6e88c
bLdyn1Vf2aAzLiAmBD89Gu6h7Lx+/Nl2e/ZXbKaTtuj2u/GkAyreUxl6QXH53kkw
7hfki/c6N9QTk0MvgmEE+0WpVAWxOurJ1xeTxLwlSbnXhwfgYjpb2kJ66sslhHf0
LT4SNsWSqhajYVCYls1yhY2E+9z4nvjGVos7tW7Kua3I7z8DZmsba9Pk3CsLXwcC
kR64Wwy1TxvCuHLr0GjYcn9rzqKeGRR+axo7ILxpFapBetjS3rjupF+QmqnkQuO5
cyfBSE3lgYe/HB27viulvpYQhSr/HlhOCRaj5ZlM3a9dk3ywjq2dOS9iJeeewcfu
ReI7wio1gNu65E6Q7UPzir8/NCriea76ivHAflgWJjYkF8FgkOVG2IXp/8/aK/fv
CTMkR2wTmuKzsZHCg7NW++Eegagw9bLCocK3uSYqc+MMUpM/u107lLo2kruDaB1Z
cyuNZjDmRj06GnpF9/8/1RdHoV6FcsdqSqUsR7hFhcUBu24/7UO/FrSWkjheYdFc
RIoLS7h3Xt9OJfBX7YaO9ABJgsgF/W07RqIBKWoIADH9oArZlGGH2nPt2PNuOuDb
Ntr9nUzHk83M9uCkXH8IHSuvLAQw636LMg46E8PHxM2jQlj21gQafW2X9MoagaT8
nhvc5T6AsvqGUVrn/P4/oyaSpu7h2Cu8CE6tN4SJ2EJl19OyKHQsF9kuIKBLxmwT
BluXQdMNvVhCrXSkhO8FZ9BLclDhfCnHiCOOjlI/2LlELebLMyk/hM7BXcXhZUrT
+eDNpFu6WGnEGnffWJE3ThISpoquJFijKEVuHnt5XiM0jChdRrlwqjyG+RL4jsir
KOwTd1E9FSl+dAZpv20iBJhSAq0izziqU07/1u4tYE9WmS5qYWnBJUJN7pj8wVxS
p5+l2NTdULADFDLNk3iwD2bXqXEknHXKO8FMp7/n4LB4vv6c8jVFYEPPmblqv1vY
14NL8vXYqkHZflHKFl/g9ccCW2QmZG9OjkAJ2WMhdhdquu5Gcmi0d/g+BjwfbnyO
iwZBfE6Jh669Hyx5mMOc28q7JcxZgBAEG6NoGdpuIaVOTBZLZiUm3J/sbC9nwN1h
UIcFSoGG5alfF8Sv5zn9jpDtGTQ1l7C3J5m5a7c5l16/NA5U221COrPzNoh3Qw/Y
OmZm4DqNTlgvl/bJ9IyjngOU6a3x8H2ImahjttiizTronr02ueHjemUL0Tbwcdwi
kE2aS+WfMPoe/opm7hYNLJjwMOlCDDhLCCoEHQpNO8mj+pCauy1fMiO8j4229Wf5
rpGMXKRWhcZQtw/FhEN/UCSHVkQfR6WSL+snMIc6KgfR6M+rydm2IXgmT0+4/6JO
wWHAbYOtr+/rfDzmWPiYiPFQGZI0ylsejjGquUqrVbPBuekko50UZRFjUmSRGq1h
yM6S52JFpogRapDn7lGdZZIOUyfMGSSrcjJ7OuCTCkBSYplS7B446dwJMb2YHE3F
jSj/Hg2W7gPSeK2ATpMyfbiyfMsneZkkMgNr7xkRRdkHlQfYFnnHuWTC3/CsrzOX
Zz75G8ar6Vv9kCr6SC9mhn0dcisIiWeaTYQl5L8mk86NZgSc/7f6TfWpAtkMAgCd
/BH2FWlZlfTPqZsyYDD2KhaaNC9k3EqR7qMPwKbGzhF1M7H0qZVjJlt5Wu4OLs/j
DJQGqeCUNId+WUAKB9DgWsPhPu8tqtxfC5B5m1LTyOjset2SY0F49xIFMIIgFrEt
cWA8Q39qclbSvgvipZdHSxIQFMpvT3v8M3y3iAuxSRQ4E9NBkTpJt+KDtKA0NjH1
juj6T+tau0kopLZVA2FgSKIlHHcTqN+IJ1wR9EGcYahvIl3vkWcwRCI37jK5DFNH
hv3Ivdh7/F3ghCuCVUpy61X55cSeye/5le5X8yw7TAngerQKb3z/jhcT3J4oOTcD
fAmQBLLZYvp9S5bjoz+E2Z04Mkr0VgXDtveGpA5Q39RXRV9IYtKCetshWlM2e67G
B9lXL2FRBsL24ftyVUjYRssaSp0u8J7J2JOT0QDVr4F8y2f966KAOYBOz/DUgXrP
pILfhGZVOOnrrFUYbZD6hFwLMoOD3XoSRK3TpABgGLlOtEX9temitOzpvAGQkKVr
tOq+CKyRRFbIhJoFCnRidb1g0TcaDvTbGFnFPHADImq2nXv/vUQaprxCYtrCIcWd
nnQG87KWco4hAKTy/UBKAUy7SMFFG3b0RVEdc6NV+rBvS+wU/Acmbx/BsHfYTw8c
epWOWdIm+0GDYC+OPvxXt7SRULqaGzEmCrsIRNwsEnwo84H5XUYecuY/tNC70ZPJ
HIJNfrWZxGByR6zh64NDAVcaasngFCOFOECB/0XoEAOMfY6LwUu+L8lthi/yyFc3
mmjRl1cf1sR5ZDMosx4YfK0LQ+AmvUGjan4Ep1rjTCwJmCceYOkd0p4M0Wec0uei
fb+zwrbMziXk9oZOelzebpalBeZdSPiodX9f5RdBbNU+43Qu80GYBBK7n/ZqByyJ
7Lmrp5HhOGe5+dIZDeVs3d37M2FkRNjGXt6XCAo9MaCEfIKk8W9pUt+XLs3XOTGE
ThmTAB5BvSZ0bphZJmJSfLlfyzwFrPKcV/xKw53BG4wthvYBDNaXcLhNxGiEwdpX
mrhiLE6krHQibT524tt6S/l+kjQt6mgOBo57Jhd7sH+Rp64jNGziXeILL1oqmMM0
fncvf+X6Lg1o4e/M2lOke7hyPjdj6oz4/NTFSd6Ly7YWMYpr2L1YQ0eGsQYBV15P
LImmj7JK/yiZ4bAhJxJ/uM/b4h+tCa1Idrv7z5tJjjcQV9WYHPuQ4VRVeMvlSir8
Rei2WAENmtBarE52kIfhdVjMUQuxEQ1hd8JMAUf4c39hVu+bXr+vxSehKN5DwCsN
A3Y0xpBqSLPQmwTxkLf3cQKiYoUi7eEKjqfPY3VvIVU1IUWQ89vhJe7wdRI9edIS
tCH0lZXKOauhJYLj9gnJPR6ALiK0n2pthgb4FihBhlpACH9y131B474Vw1u3kzpE
u+9BKCPfAdXECdfH7bbVW7k4K3JvTXBIxxx6T+ajB1atshfsZI0bIjpI2uw5v1mX
np+6dFXmf0qwelKjVhwlLD+nsWzMvrzG4i+yij7aTNoFIVwSPCd+2PW8Ie5iRuR0
StFwXO5KNQjiz5/3K+BRANgXly5Ir+ND8+VTo1e67BO8U5RaLo5mlYcbN0Ls4Dmz
hxAAeNZeZlTElh1r4CyrtZRMd23X8GCaZ1WvhFdyGOihV+hA74zr1psYcHrNjUIw
KRDQ96+zCep0cB5gnxq2zYGHQgEUPtCb56BLPQLYfqYaQST8DFXK5w+duE/VrYsU
4Ni5JgmkOWACbryL/3azVou7LFIGvlDUrktra1w+xt0dfCbkcFQKbORQfMz0YTjz
HFf3l+W0Z8TfA+9TV6lHaVQAPFY6cTKqA68lzZm3CfdzTrxsjfON5T4YcGFtNDDN
tI26Mp5VTBPvLDQPeNJ7b7DOlcYIWoxIW0/yKJMm8+eEjKDwxWKdFfI2RIDfTAV1
R4KxqFWaVlPe1oBGNbsYMDREn/hdfe8IC6W5LR+DUvSdMmr8kaBUN9S6oC2Elgcw
0rz3np+wLpn2zoDEm8cQ7B3g1MUm+Nwu7gyZKCDUXvzdpKfy28b0Ly98gbSyGbmu
1e8ge7OheHuoyfTf4AOGQ1b+qeuZlwuaghzUIwp/p/9iEQphrXbtHfn7QTJdD7DB
/rsUyyC0DbEIWKYX2aYViW0/cHK+yWFJOICTzY8gUCnFgolkb1JTHt7wyQr8JKsl
8j3PdUcBXldKozAx3JXrqa1+m6qV6k0mxTy/ynJXGWbQ5orkdIlqJlZxLOPb8GnD
VkK8L1z+fROFI2FqD425WEzWuzEcEkK+qkruKc9J1tIz+eZJvntDOJ3PvMJMEOaQ
CsTbEznrTCONiEyirKmcmsgQ2PlnyMGwHHpD7+NNP+9PR0WyB68fw7Gp9JyWxnFt
16EVfo8Lva2Ca52IJveIvlay5CPfIuf1htUO65qDhAd11ZDRpZoOMubiW1FDcor/
c2sY8ef7kdKOAvDUuGlZ2qztnx6hQ7w60chaqS4fW9Rs5rYNIwkNkjUGsTaBerbz
gJ/2dC4cVLWeDfPhyvJtJ/8z0i9963/9hJPjPlP1ApQgmJsq8KhEgq/ID/WvObU1
x3LlsLejfc6iCofn2CRWID9pJrAA5iwmobRVdQSRm30/KgUdAQun2+8cQ7RbPvId
OwqhK8J90VESdrl6e3v9dsNY279mWdynlAlLyPXJrGzQBm2h5MGoaYWL7o2/I71G
A25Pfs6fsx87+qPxiIF0M9Mk0siTJ1afgfKqlaAGPlqNO8VaZQvFhnaYOQ7GfohI
vrn4zuYDJfXBfSZ0kUdeBKBpnZmjbu9okF9+ugX1bEZGr1sIT7gq140yz8p39vfm
NgH5wKcGtIXdDZn5WIq9DhmZLv4rdgBQiGpQDuTz/jYMG+9LUFmReTrKvGJlpU6T
5mREOxYVDatKKEPdfdPYU4rnpFBcOPixOjIc+pR2yNXARZn1x/KLDZc14dZQz+PX
Vb15/IT436dNckvzFRuAoeBKkw4EC/Q2ojDVX3s0i+cGU8YFmfww8u9kIPzX30nA
h4++qVyD/uZ3vHF1zBbck7wW/PWxtDtMw0ddqbcsqr3XZRVg7lEMtG3wj4OqNmgT
v6c8p9GOMIROaW7EEld53tELQstvJfFp96wAuXZLFd0SErgAF7muZ/ObKcmXkDgk
MC74QjIL0aZ5Ld0uCsF9QzymikqlQuHyQ+hM4VXW/fwTmu4gu082z/VAy4XGMCFC
6dmG7vlZV+lFLWI1MCjXKJKViv7dzD4AzXAfWPluY0LwurSisNerp8HDk0qSqESm
X63K3TEPR5Z8wkdMuMF88TiGK1nfUBoFtJ60MhJuewNf5f+xT9bWhlYXHzGw2XVf
634Fh2VogensxhO9eO+yZwb6AyPzwcpAWXg5E45ZWo+pK3twL5Z2iPw7KrtfxMkW
gNslHVI4FQ7O5OfkgXWWdXfrhUce/oKtW4Q+fIQ/VaKwqCPTaMais7qKuSXQdeCg
bHR5deuVL1jW5eVpQiXtXhRQnItLINUcXFUDaEjrUZhKxgeJe7QsYbJ/QCirCKMq
gvxmDhy0AyWnKxqsnLMlG9agu3x/+6oRF0LVF/SIzyRIsEwOeZlgjCbmTjCjljCN
cPDimbFn2qKT3YTbs9CHAhivA9nbua/DeFKi6+HmVr749089nF1PlC7tmDwsove+
rLU4MfBeWK8jOGcDY2YZOBVHDt1iKl6pwncgaULnp96JKPred2GnoXyW0CKfLKwn
XgReW2p3yNfeEF9OFX7WPxTeG/dmopYABUGVB8qElLB61wmu8hID2us8v4yLS6Qe
1/USd3tt8yUeSKcDiQURufyqfJlzjrlvpYDtU22kYWo19De40gzdkdJhIFg+qHAD
aMAVin9/Tg5mtZ3BQKf/2ZGX5crwhUk2hRHieV+wXSe96LYdXbOgOS3Aj0aPcleb
JPst3Q7FGRK/fnOcWQgXw4qR0IqBhA5XpHn6yUCDzavSkhPPa4hRvCKfcIbyoFiY
VwXPYz2DTw3c09ag+7O4K+w6U7odE0f2XRpnzbPYzSGuV1Pdze9xIHKGvSSULVtr
2pw/87sf2cWLENg2h3he0xYezpm3HQ/MYqFuvHB7II3EMjWEJFM7DrZD6j8aMKJJ
Y73yI/BGABzt7zWDP7TLGLS9YptSy+Q6eWiktWcrcSWu1t6si00myZq8/MDQHwaV
0cY3hEu9ugiWDyt6S8gAFVUkIGVzg0quGI6rRfwW9vItXl0GNpLwtQyR6wqLN744
cIAR7hFhnhdAveEMzuYGYij030XJWzzXLl/wlnh8XdBv5fS7yvshEIlO/N9jT9Ul
lmDAu2UhEKmQcuoa7Yk6fDo7BEls1JrJd+QWJTEYNZrUMONyVeoh9Y65l1/dVp30
jsnVP6IWlaXfOl4UZL1YD+hjmgDFM5t9YwqbMTqiYWYbJgMIjCufXeiAdncC+8MR
TbmzUCwYFmf0fe5PlgZfgnoJbOOX3GrliaYAp8GJSXe1VtPbbG6ZWTFdfm77Vf98
RXbP3K+jeKJTmHbhx+CohYFZgwUofWPlO6HVwdkALAD/Kns4/0xFPNHWjxp0vPR+
70uZIXXyRM82e3VWGQ2xZQWNHJA6a800Sa4VVcMBEl6fz4qZtnHBytJ2P8rtA//M
DkLDyRmYzmmRAvAHreBl1UGRac/qJMJvvw311IABHGJI50JD9kIHBm42FcvDGBlb
5sl2Usv4vHZ1dpkFdHtZMTC3h50y/wYN3hryHFwVpAlWoW/MK9JFSPRXDOzvvilK
lGY5d61XjBzpjR1ss8pNeMoAAgWwO9ndeC1KbDatx0GyUuqjuADkriO+Ye8b+fs1
kKrHtUG/ThuLxyMjNWPITTQHYpvIzWA1z+l0E1BhCU6lm77PbcQtPq2AeR8Gx31g
sFooWxcJXNNxKdyLLoh/iP4nYpDCHkirAD3vo9xKp70lEj/jCIL/7AkAacN64JpN
D28SI8QpZj+fXkEuOSphJh6+mhUKbhUkQHCZaetn7zgPonVMU0uWJ9TbWGheVCNi
t0oWWZk/SZrj9ZdQ8/cLkqlPNGTCDhIDeJGb5IC2NfqzeRsiugCFmUTOit3PZxJn
WldXw9qCC9ih3YD0qd94SUeI5JEM5eLCIxN/VLwhK5TW0qaq7qF8LR0qHPQ1DVcr
lMFQOUhXgciBTXbpvy7vB2rXHgso4JbvJSW20jF1EcS5BW2BoCjTQ4Ic1xe1cSnx
pYPDVD/kvlNeEnmpStRuTMgpQepuqddDTj4nwLj60aG7L83SVwX3S7xfo/RZb3F5
QbB1RojDV4d9ou87nbZ9s6XtineFWYfqCm6FXdqQOUOkhys8O2pFkfWVUOrp5hm9
ApDPmiZ1Y8RQUy0DOv8JP9INMbCtmOEcadxVNLYSnnOxTJnGXb59DSBMpL2c9mF1
LHiJc/LpIV0+4AK3n63Z4WKzOTVgVHLfcSjN4pdOjUjFLnU5W4gfKzY1MrEa9C6p
mX9AQQ2hi17NRCfQrtl6UkuiKu8iJ2IZE6rXGaGpT9ZhIJJ0AxXkMO43Nb9pjx++
/s/65g/r/OOeljRPbjBoNFw6ziePqfF0j6Yi1Lploq2BI3uI/6xIG5YPvXwBlEpM
/+i8KiOCXJ2Mu0EGO46Rn8T8cHvCK/nsO8IvO7URd9Sapw36WsdakQ8LSJnNY5sD
KlRoOqmaq/eMxxRKn9PUnVA2Ms5stUlAVgtiXwaLoJD+kAu6pzggc+QD+PZPQuEf
uFAsYZj2/+Rbq0HxzqrhgRotPorfyemuz2SbC77D/HUwb7QM5qbtBB/NvZQnvrve
wq8B0UW8RSURctcQ24Bmd08yQLkSzwxFhFK+MW2GD6cyaLu7+ojdHawAeda2Mobz
DG+8OxQl19332oR2ZVTWoR9x9+FuU2JhfnY6PCIvmyN7bB+D3P6tBqSyTsSjnXda
FwtabLnPBSM4C9UY5opPBYqikBbSLlaubULQmGsUk8Uz4JVyigwWgIM/H75glct7
110fKz0IiTU1l4kDfEEHjUD+z5pQspOoBV4SjsPBFSDak1hTGkJHK23pRr51/SV9
HE8sQVeOC3Lir448TOsCuBJ9LlQduItlAZdUoLl/SmBzQGnWP7bUDS0E9DMGaHW/
X0rg1vhLvOXtU/czYeVs7u623yKwk6mIURioOOcCo5ZnalwbTc6qLd+faJuEwM+4
uNEvk7qkWBkSciwQS1vOVedy1jmp3Pnmx4iO/TeyofdD13rwR7uakIWRTzu58P38
l2OnRTyXpugyQdsdBxcJF1lmEWHN+UCz/CC6oJenvwwSv8w7qL5RIwDktZeAWoX9
AZs+TPGE874LhJfska3wQXaQzBPsxo9knPKGUaKqbABt4ldRqikTeqn/e2mBsnAN
QZANJ6927evlJgYBpwhEPTxWt/XMJuuNAKbJKgnjCiuICdhZBLQyKtl4sJpa0q/t
Rp6wuhtHET+4mpgNk3IUbmjnyjCz0QLFZTwRWV+Y3dzpjumRJe4O+CayrFm6p0P6
0jcuyPAWxPRnQB5JCl+wz/WGlgDfdSh6BGvU+NIXp1AqkxlyMq6v/RbozSXQQJQH
HRSGJ1RrOh9CAyJYJxszGq3VZKMQo9Yp1fMpfE3WyMWDT0HkuG5eOMO9KgQP7cnP
LqukmMGARbopi/D8GXOOn0vf7HCNeiWbFryLBbRtM4vYqcQLZpRIQKcBxVV7L5n5
ICjORZvGrpG8FkGWUNpukjLi6V61eJDlvwyflCYeMsiRe5ixJqBmU85VKQe8Tcpo
LPgeBZ0MIA3up3TnRMhuNsIkv/T4MO6F1EPvy3uI26XePQdtdTAvT50WlBgyRjDB
vQch2nBTliBDZfdj0Yf9Uc/1Vu0djPQvlv0uhCPB3FNHxh1cuTQX4zuYaq5TLtYe
R1FTUQhLYVARUpaofxpFFx2pO2y72pM1dU4UkvtjA1GEQeLqMRJ/Dpg0VxRkBz9I
4yof6eOyUbzlvIFOQEASl9yPdBCVa5/qqVXhgvcFgO3ZH62EEpRYociUPeY4Q4HV
cFMgN9Y7dSI3xzX+5R+BW57w3pm4ngLOzNgD4/s4QLdZqMAnm7DFxqzlUVQ82QJc
F9KWeajHE8naLFuYTlwf066rVQzSjV3gI/kSlmP7x03rJO89yxwbEeHGTnjj9Rwl
Zj1xiJEu60MWlHHybflHk2SwEq0Y8eXKGBngUxJMaUrRBzIKacmhsuEXahad5FGd
SEDx9TfDS8qxr1AwWz3eVCq5vuKi/kmA7NTA+UNk9j8paVf+lcpJE537Lk3i9Np1
SkKeiuHVMYi9ybONGbhqj0CR6h7QkjQWL6CWX0x1UkksZaWRm8es2/rpDOyRqgZV
Lb67Ztt9+kuMWL4b5S/GQuQplYP/dzDgU7IU5gqH52eLmAZ3yQUNbAjuyPiuFteh
wE+U5qtO8tELY+nsYXMoJaA/bDZii4b0yK0MKdWtbooKjC/faNQZJuLeImIrACZQ
nvlTIZxQLcTIjFxspCYM8N6nN7yBzlbJ1V5drDgYvRDJvpIiATh/EomMYMXmXsUk
qrUrFNM562OUmjt4F78qqJ6U6q5cMCDGx6FsgmfWW9FERwaDBWCGHKLqO08opUmq
jA3wG0v2kq2euYDDFV7CEROObD3dDKM7cPM8wkLTGCV0FumbtOZete+aD/qQT06R
YzpOg1svfY43CYiZtrGp74P9J1QcF9Yho1ej8iGM2i7GVEchGYA5N7H67sc+tAaD
KP4uKsidUOTVT1g4Zi+RAD+f95cXE+JRIAuQAnPeSzYhBPvE4sR4mrhTwsUE8HHT
lLzv26et1H81ZihbQpROOlSTf9thPTUg/HhHaaBYIQP/bpZmOu/wvkNd5Qm8Vu0j
AH+DLkGfnIOw5oerHm+ZZf1Shcdam73CelKRXPeQZE3AUXH/PkXtAna1y5inmh0K
4BiUAR/EbTGyAsxabOvn3oNpSPoobqBjZAqm9tUKHQOwR8yEYI74nh4CMLoJT+Ww
zGbkuGZIV9ssUsYwMzoB51VWq2xFIHBGpbXeptJoLDbWbFwEXe5FE5o4/geR5PbB
XfGt9b+jPaQRZBkEeiGvEtzYXwn8/acxrDXa3vaRjvk61yz2XFu1/PpqHuDws5EI
JFLPr6ZjKtuFKMIl3LSLqU5HRL0G/JLG9HYxyuycNnSdVUwNB4LUTyoBB/NdYhQS
/tw4JbSuUWFExkPs+WT5zwk5ZmFrl5Af76LUnictj3L/PZeKHfbFBv6B3td32VHg
8hLAVz5MNadpcun67Ebpg3UDUawfL3joYBvqQ82Ru6rP0OB3Na8luWCONm56+g1P
rPeywpD+U/Jxxbygux+zcvRyuezMnL1dCPhTnAD8fs2BBOC6vOdl9XkwSoRCXYHo
ZrLxe98XffgwBb0PIe88n5uHGUv8jbBQS0Q6blQ/9iBWJdTKG8z+canu7jnOUkk4
HtBUsTZKI9N5S6LlPGQ1UgTAtAso4IP7FmjR0dIh/iG/LhzqqtYvotzYWBjbvy/7
MquoKO+C0Z+XD/HZQlyyupeJyxCe+R6+G3rbZQ1ItK9l2QvSrf1ZOxOpdmrrzDOC
5HltA/P9FXnGYfzIuk8xC/ExKMg28J14b2pilB/YaLq/fedMOe22e2MYk/WMfHqp
iPiMZBx+2czoIBhKOTY6ek+RCR2+I6k30uyVfdmdGsUJmBVNIg3fCIKooXfFWLuZ
WxMlyciZpTmgR4+LgPZq2UCYLTh9V5Jhdp2e8VAUWIWs2l0lQkocFgZRZNyPYxVd
TodZ5yqC8R8zLt3IRywoma01tfHcd5O4FqI4te6VM9Owph1tWiaYEwiC4ZBNMoFR
VvqKiUf2YFVRm5WMvitOMT+TIc1mLGCPLIzlXBStLnbS+IylOLFPjKpqv//lj0Wj
jhJa/lvpiUy8GG5GlfMR7Jy432B1mjJC3UlXebWuSJ0csVKB36yu3mePQcrFAUIZ
U31pi4FbpP//+Z3xXlhZnTvjAyM/tt35tr2Mr8U6X/YecdcW+UwYTnZXlCzqdx7d
/Q1zbjwK2XXVfrobdLxP12vIyW8sAiW3TI4gKQ+dGgchKXR4VCYljDrQDeOEYBO2
5LRr7jOPolUXsM4YY0RIm5O4FUxBCtL6ItFKUnH4vZsx7E4imIXSUTH+UbIi6PLY
vSn1nqqmWLfYVvuMf5whgrD5A+U3HP/t9W9Y7KbzVuJaQ0pyfDzcETQlGH3QCT53
aJddCXatq7GA8Q6o6Vhl4Segcv9zB7nMqnvb9VtstLR05XUPdyNjJ1OnaAaxnPUj
Fz2GBKgmJEib1xZdCA905XkerXze3fdljquH9fIdt1UaireoDELz5aheMCQZez1l
ijHaFQJYuloHn9v0xaqGP8FoDUnSB4hA8/d6zGIUfMfY7Nkv/lbjIvGxnIyEEDUB
Nb3u7n+mj94SNn68+Nn3v4eIH83TFU6dLrnKy0Tqs4djXwUwkPrRtrdziAXf1YfZ
Up+L+UgvIBG0A91TSjrJNuqZZTBAaW6gUGUxyW33P66OTfQBVSqbk9/ep37k45mf
I9yNU/Vb7ykjjCI2sDpz6pKa3HmlsCoJBpYAhnYhJSeeM9xwzywxjBwVWXnTOwYN
zB6IoucdjePNSuxi+emfSzMZvDxxE8+d+B4z8LT80tOZkOFAb5Ai4XlToSqfDg3a
eZJ7IkFUow8hIr3DzYngiliO3Ty0ZPTeybUhZRIJ0nElGfZORaBzp0/SzCHrHsoP
GN/ITc+lHsgqEH08SKD+rslFlXcRF6CAklO77yoTo+j2VQWq3sAXgVT0hAWJYaz2
l8xx2ZpMppGGIGaSzR87xq3rScndCWlAfcHkk0m+jDgamxZbAmF0IJnfr0GsF2Hh
lzgOjV2cdH70xBtotyatwdh3CMBaZoIVp01vhJc9IwFpaEIFlvfEHW5dAf3EPK7N
Al7dsAwoMKmvhxDLYFpr5JcVQBuVxNz8hZVbb69vax3IRN4T59uzQN0xMRLdSG0o
yQvGtN45vwjkpnwrR20o8Mlrck/XIIPE3CgAXkA1t+9Peif5rHRfiqEIWu63xj++
fY68Voo34HNg1tf+IsOfGc+ZmtWnvnOC8E2jbTzZCGd8UwUZU5ESX1y51X9meqzX
m1yf4DTwlSsoM+qhM3vX+9Fhp9a8/84Lnzou0nLWqkjoTsTTJ0mcbRPYohKFyjnX
Y2bnqjZwKi9I5NurCg29M9rPSknGH/nukyDkgIAhvOL079cx3qVQ0W55rn/27rDo
Mf7XqjrFSvJeHyhROAOquL/fajMdALIUpahk5xCvW3emitsNNgmzjaq1ooJnTEKc
Mm9b6Q3jMJZwq/OAUXnsPdVFLwZd5bJHvRfr0OUOQtuaQ9DPdwAOAldZxiQVajZT
Ea4eCm8cJm/EVvZVmMzuSzyPdURLMOOZucpzQ5oWL/dNl8JgnmUY1re+F2f4E1mf
oqtJ0b9mQgRZcYuFWHOZv6UghSoHH5/Wdt44wNXsokYhrBhcao04iTInPGELmdQO
brwdcu0tuPnvK9CYX2Uia88wSuQRFFrXLEdEYGgLZfCxjfUvXdsioo8z50YF8ihh
FfVv8PhuGPM76XkofzNf6Uc3+6vPG/LdVumYp8iVDT1bsxQKuKUR4/nc4v1PvTbe
gmDf3YMYHzG6J4EuNdfQgPLDXqpwjI5zBgrMIEB+9Y71DmyMZyM8sp25lJaWSP0B
221W9dcrdlDdOmEAU4T5/WvAUaP0zNJOm+og/XIwbF/N18L0y7h8nt4hZawlAIsT
iaz/iv3El/iHYsXnnAmDnEbxr5xZ+NgZ8wipEgQ0caBcwghSkca2WeFP71nRGgji
LbnZ4p0/5JiviRMkdtZJbAzAZYdS5ra4EbddLZsBqbV+NIeAmhYHwMYFlbr3BPJc
S5A/aFk2xGSldmjzYXz+ZfGScQAPbk51r6JApyM0DrH6rjn4FLVYSTl3MBcFWw1e
A/aM/ReCSHy+Ji7R2U26ZNLbowHemq2Mb6oFVtzi/uQIX39BvamseDSa5efXG9nf
Da/p29NQMbiv9xGsMtniJT3BcHqnypakDgy+VYzCaHGwIbFPrX3gvZhYpchz43ji
5dd5x9wmEyqYX8YAs+9rm13rU7lr9r8hbpMlQivRBJOqN7KqmhfU3U9HiGuzc8Pd
gmvTupkp+cMlGGQzM9+D/MC2BZZp34aIO2GdZc7fjG55Dr3tOFINsFpdbLIH8GCG
1p8N6uxwVWmov6iAZ0bK5Hx+sEgOk9WsMY8/cRFihSaxDJ9tSGQ3W6x/xTpQNB09
6b1GNly3rxm+UD389SXgPxstlC2INrxWi6cC/ALGmBa8LOpHPEGSQBg4AbBkFSMp
4Tf99BckbVhE88MXYq5LKaqQynguF3Ax9knWSYZVQowi1hO/bOamzcHEWcs6tWtX
BJJVsHeUlA+xwitRom02dwRnV+T+mZYtInTA5wmQcM2fJpXRxuJ5i8wEHYL33nAI
svWKz3g0gTgLjiRHcxxqqf13Phtpe3u7TvA3+FhUbJNPU14xzWKoipG77e0UpYup
XwzBN05PuUhHCWxNV0pi2fNAijwRO7wVOr9x4H1KBuDTEASVukip+Jx2sVDEGoEK
XsfQCBfgYvTXYYmaq8kmdzZnhdeG/s7Bm2jTpZPlywNUseHzC1/ctWgnuPmqBymJ
es3iKa3OuBjp4YnkmVgp30eubUmuKj8nqChun/LpOkMQujMIHhzTGkMfKEUE8R6d
Z+QCqzW3QexIUqrSqs3D4gfxq+cc9t2rs+8+H6c6GV4mqRUCT0LBS+VJ5g46H5iW
mnb/jELSDaV17MSDMDNjnrYOmG3kA3bzafk0IGfcm6yCbye2yWHwksRqH2ucXKGX
JhszvkPwfdrUEenLfkYkgzMhLKlD5VkhC047/gO/ESJgPmQCoLoVoGGJG747IYCF
Dx9XMVMaHPjBjdSZu/X7rEDLaLJMcojbB4oBbhvqC/Qr7FO4bsgu1wLn7c1ZB01X
+4/nRHOaGt8b1/ByoeFGKeipNykn/92Ulkg0OprDyX60vUnCvREr5W/weh5sVfi4
zLUCxWkP1Wt3/vi6D4OfFbMIbuLbFyHu7G3IqHYCEvZOQrDqtXfjQAlLKZ5bwT4N
Qynwr//TKkxv8L1nsklkncb05nI6YDXEgvADgjfR140B2hBlDzkIUoWsdZHhpKD9
rupYcxpJqi1nHW6qXYveDYEaq7E+/wk2xqK/4Syil/aWyV0tFG0Sp6o2J2sAJ/Wx
yAw+BOpgw/eszLzWK91sFmFQc11ACvjG0dKwboMMOg4k+Lf7Yi9lf62OfW5fFS7y
NYSNEgOy2kdpnp9JpC0mPtrxNAIj0iSU45WGxyLX11hJ7w9SzpFihfAoydgxV7Wz
kPOuF1sEcY4wcL0I4dkBEysxtkO2MxaIK+D/auklnuM9Wh13z0Gh3mMb/xm4Ljag
0Sq/jelHOMfJ+FyTsTquWQ9vdB6ZHc6ACVgA9PQn85ouPzrWQHkvC1wLfQSgG3Ov
bvdzl7iP3e63ikyiejUeGPkW4WrgZmcSFP//ZGBApW9TaVKFaanp91KOQkcDtUuU
B5gCfNyeae6bN4jAcw43UYCQ2YKmDAlYxlXvqaNsDN0L5w+ZzLHsvn9NHgAeJOkh
Iu4Hvgqez8q+gzXbgGSkrJDdsuW+yjsyrSxHdVh1Lx3b1af6rxVjIAH1bQ4MZPoT
d+dFZG0yVi8bycd5UOevV6o19iertIsl6vOwftL6tfjdkAzsU+OR+GU7gMuPRJqD
FPooZIpZpA3EYpo5c30+xj9xCrw3YyhEA6lNZ47cTYH4dotuEIXQ1XquJKRzf7ox
c7UM/V+la290ivGB96VMihbOkE9pFy5mLcahIg358P+fyLXRl6Mux0XABm9+pa7J
lhTNgBrwXMpMP0GixcW23GHKTpOP5lr4JQG9lKNQ0V1Npcj3+nlfcLO3VET0wrZ1
fPbCVCxumXD5fk+hGTUOaR0d+ww4Ml9DoE8r+YwOvzKm79FQzAqrt2BV1QzFG4jc
OE7x9CmuIZk8pl8iQQiNniDKg6LTfy5ygjGKZnORebaAzmFxJC6ac4Nj4hYJo1t2
R1WjGH5E6JgJ6QStED5gI1z91Gt0kQM/nj1coLIUevdS+ZrlXPETMkD0VOx5XC62
YfSM1BP9xaLpV1F6O6vEPhbEDdur5z56dnwR6rG2rIzH3hesGqgwqP/F5GnJ5QBe
mIluAWpfE/9x7b1JmKM4MVDG+t5ioJe9jE9ORvrpz8twiNJaSUKwDykgezeV67C5
0WFi/038EPcbdaInFtyI4E9DUhNrdy8EF9m5p6s/O3oxgpMUDYfiqQqUP3YUAwQS
VBreQlMMj/tch0OL4C0JgqwOE9CXuwPmVA4xQGubteBucwxi3v1psjOCEEJDYPyp
NHOhnquXDsLbrtGaOJ/H8dKAjl94lkgaT3oeRpqbBKQ2PaTJfVG95H9wKw41W120
UjvzFF1TslzzYq3cm8v85diia/FCS3anuP2Pg7fNRNTjzJLmXNuBgBN3h+W9CmCj
aty9UpDAZ5yLzEaCz0y81DrP9WrWvY0swWp5fQryNxN4rnAFk/cAZA+OpL2bZV9z
GAjsSVZXhsosI09u9/tx/6YXTQxZg6SzY9EiIB0/pU85QlrcXkhHtbUh22M5TlN0
Ch6i0Dyp5iA7erHv7VR9tYDL6Bwv4GFgBoH5dYxuUBobvklyKuddm0WEcdHjGcBN
kqzuAKM7Q/okn4CpF6UesoUAhe6VB8m4Vhw1oNoABv1uZVUZEXSRC7bx7VgFMnck
7OtSIYyGksOJBLl2VUR5l04e/8I3nKMDeMVNO0Slc5q8+mxarQ4crzmMydirZkW5
8ZKJsA7nC1rsvdjPo4pdbmxWES7S952PHbwCRAHdwj0w68PB6JvvkoCapvl2dLZ2
ReZ2EUiF6mD2h3FR+6inGaMNhhonL0Q6OUewxSWUqt/SQJMH2hRdwRg6W8xqYca9
RYLEZYrVCUd7MHkyLxCEl9yhRGlXLUzqEgxyVzeLjbTYscKDQZB8foPZ1IWJhB0P
OiWmpi3Z9++w729nvbK0PUqpFWLxM3cg1dx6Mrgpp8koTd61Ef4KAVuamSLdEKZR
unVUboQh7DLq2gt7sae4AW+HRymYFQfZqmA7wtrCI/6qwQ0Kr2nzx3E1OzZ3I6HL
8BAqera0Bip27B4mU2P6tUAVneVYlblzeHveGCIARpzP2BkgcYeWaXV1OHjYS6DH
i1ZOIf1OieM8Un/JD/jDF+ol2lhjX/J31U2hO5d6fQM/H0W51wdeUgZyglwMwi2U
2uBjSG50tSoe73y0z73sz0FZODKIWPaAkHUvM77yqoxJJdnrCDt4Ou+qCuMiG+re
h7Dm8+rBawjiyZVWqenRUO8LBoa8j1a1SSm6402mTuVIIuiMDmSxG/qWCRHlEXm3
BEKUmFd+/KXFTk2nntIzhlUZT75I6tnO9VfWVLFaNBo2sMy6Zq6fb3XHrbUr+hKA
/UDDC38yhwzGzaIPd2US3lzLV2bt3Oxk+nDV5Hxzicl4+wqcm6xlphEL4OegfNpa
bLoZhH4PFR16quKS1uAqx//wYmokJaDme0FkGOaEmzfLZ/pHdI5MLY9Oz3GuOeh8
YMJ+1HMv9ZJJ7yjovmDQLrIISYGCqWAl5XMwip+69zgyeC1/9u51AS96rKQHdqQX
BDALaedj8CievKywBSCP9cT6BtBHLuDPvsQsnHDQBMd5N3e9MnVBnUEmNJSli8lb
Gu3q0cC5dxMtDiJFbbvdHyPteOjKVPfhlyEmLYAwDn1az+JvcALh+c3r9m+sACn8
1tsYKsmVQjZVXStQt7DFAsfhTIV7mi4GfyiTwwZPlcXXiA7UAcW5lxtfbXDx/R0p
QcQ5uSgNfcD9pN+LgyqnA0vah6a3JJ1Zwm/q5SCPEIBedsYm6w5bEb7Th6hYtsuc
2fuvMchmN7sQsQ/Z7ekSYA0i459xLUAreQqF9yAZD+Wqm5kcobn/8YjlRkTfLlWC
fydxP6kFdboaD717I7MHVsTXT1cd/qMVVLoegRkQ3uHR2V39yLJjJtALSFw1hsA9
MoJaP4+FGy8BNWL+eyR/P+Kso/h3Q5jcUUVVFECQ4fj+wjqOQtZxx9E4cR6VQLJb
q4HyWAdI/8bR+czIAk3UasX9comx378s89k3TiQpQ8DjxeRZpKmovd/5LYX8tWI+
rabYCEjBuJnvCA5lQiXnlaZ5rjY5Sy+HYBaW0v3GlIAm0euczVfoway5ZerC+7E+
q061ibHChseMu5Q7SHrTUpSrwws8Vbhu555PzKAwN4UJcbAmFY9u8/QNoFWuubos
ewGi76nyeOfxbzwQqdNIHiKlO+671lJmbOtFvGLEVpe0Wd1ngq1XjAOM9DdLYgQf
MHJxVL7hYOw+5mlGlTLEvC21PYfNcsmo8Gtn0mF3uv76Gh7QurfZ8blJEWYjkRcT
Bwohyvi+jaLPgm0Wuj6KOYvS5JXP8zUZVcpzvTxmZGn0qWnq0sdElUQceiSt50hF
Rb9YczsL0+EgLUlrfndvv7R2JjFRPxFD4CDDbmm36HLAkurDmxCGmO6ffgEmdsKf
EUmwqZ91pv7g3TIbG/32N0dd+gwNfOwUQTK/enDMKPZaNYgJBTsY3sW1lr9sr+91
+em5U1s4hcySi5p/gRO2232DgkR+D2bSsFOHzwuXo6epGop77WKSQF7ADh8V+gmF
rm7n3uhHwz3XiS4XQsVkvP2n+McBKjeVVNHrTQ2pqRPKzMdtN6+bzB8e4qpJblRD
coAuu19KG34Kur3HQBdCUi+eVs/We9ovpThjJLVagq4yuod1fq0BNoGC77vQAQFc
HQ0koQe5alVEUQon3O4gbElw9m7ef8zagGVh2Lqiiu+hhgPoqJVvrgP+sEMLWXl6
dhoI9f6te5VNe9Md29KxsK+MbKfheB+0iM+kDRucj4a0dkJ3+j4KzeJAkeZBCRc1
I8dX2y1jI/pOEcRu6i+wfXBfG/HGf5Zdi8DKfFO8ojwf/Igg/QstP1IXa1JKDFWX
VUNckOzKblagEOg1UAH8SLiqrCzvYm7gNRW8X6eSwPRYQrzOBJ/Gy2TuEJeec/0n
8d1TsTpoMYoXHugGvOvu3GyX9Ea3iNCrwRtjnf/AJynclGLD/MJACZahZGQhfalp
0ECt9ql6hdWdn5+Q/ky2dM8WNdzTGNP/QeM7HCml7ITMq8U2VGRC3g7/uu3x4k4R
T2PMRkdICY7VKzpyN+Y+wJwfhSVch28ei7XLB7BMd/6xpQhqPx7KCNQrhDKJCfdC
3qHQ62shuM53hJ6NXPrR+4zR+ni+ZVL5qQlGSNTKe4r2GJn2g4IPioaiaHhExlnZ
AfEkUqy8rfjUGWjgd6orgeOPQbMjW/VvpWcmVZ36RlNDp8JLlvZ0+K9OD6e2OVJp
8uorZpPwioTzoftYUnvUL7ZfQMl8bZhUnKkOg5OVRML4zWF/d4eQGBC5E/DXGj8T
PtIX+SySLM0kGHk40gXoRc22TmoybW3N+84dtjtXCqI2enauS/vTQFoPwBv15Pma
iUNmpvGmdq1MP0e4lgxAJQlFTcHQy4t1/33eS3TOFhYnQuDOs2FipFn+goDX5q5U
9k4ruNt5ZAi78SqJpZWQwQkxaFW0iAZeQR82j5z3PeWbr7fKNnV6TQT7Ac0f+1f7
39I//KHfLAXohmVLPywzI8IRPC9Wh/tGtZZg55bDAKd+vCXmdyQhiUEPedC1p3F3
jnpPHRT0Psr8iB5VrhxgjKOqEP3FkRrExS9FemSoaIccNs/CbYqglVtb2HAqO4Qo
Mwp21ZJCSdoGlc5QDKsBo5fPjxZQZOzyjSeqTaJscHLONC2uJ0Zg2Gh0HHoqFmPD
ZqHFx2n7jD14Mjr8smfmyb37U7MqpY/I7drEjPVy8qvPSeN8TRuSdto8PAMwse1V
UWEqp2ZZIHbbERtwsG375VMC5qPOXovZTN/lyOk5nsqvd1v8ZnNtUSwN8ru2Um9u
oFaCjnUhzu1I2PmI3IIJPQCT/yE90ls5tqQawK6zy9hNP+jTMCPJlO0juWx2HaAb
Tv+VZStBBM53J0xKG4oT4naVtl6dRGL3PEcEuOHpQnjR+9VBDaxBGwz/+sltCtXR
dGL18YKRbRCK1ZIvfQYKpxrEO7Yd3BRjegIcje3HnXpO4sVFzJMQWXMsqea2lJzN
k/+VGZXibFZ8mOfOmcn3pGK2Rk8y0xZSi4YuVd6ME6sMd8MOdxFAdqDrC6Npy53u
r9Z72D/KjyyabVqzkeOS6hAYZkh2IoivlnD4S8IUbDzqUhrg7YH7Kx6/tdyoAoMr
fUXlHN9UM+SefrXMpoEqFR5V7UD8f8fCucpKMJ37/0MTnPufh5PU9bcWiyFIluPJ
MsjZ56/KUuVhVsMxRXqtb0jfrs5P2cGTPj0/3HesN2gAm3KntEPrRXYVwmtdN41X
H2nsWeF8e7/oXmupP5bjxp+1XYNfVHGcn1lY3Svi0OsfLGHLE9M98x7U4IQUYccZ
w5A0m9nFuCm+k8F7U4UDQu+AyHzvKFAzoykBHPs0v3IoaHZ/geECQsbbPMA6bQcQ
iNIWspyojj319+30SphvaxkqM4E4ir+ZqkG7qAktPVLP5WGhrjC3Z2Gzj8y5dJgD
EQM17j2wWXWKc3jQyIvKQzgs4o+sagxr4j1UAwAWiqPaJpw7/Ak9FSgZ4+Mz4tAy
+9AAuazItNgbYcT533MIwpbg3+gQie8rLMtjnWSoYU06Merguvch7UpujBH7zcN3
HlCsxQb+5r5suUAySpimzdNWRa4wmuIK4YXloIexC8uWiKw/keitqEXGcA4Heu44
9378T5kroRyfunsN5drmcDXTQVJGuXEvHzZHZcDxdlK6f52fl/bOMiv+5gF929wl
KFOpGCJ0YAY3GzPFFRWY6qCYRd/T27JJnI/V/haBxbQzY2Sbd2X9koSal10ayX/4
hXoVeDNMlcPNvj9XXaXErUCPZgHxL4V4x3EZxlAKp1ZeAcxF+CDZWlJh4r8sXjgj
+o3NwvwYkJeg4/c1K2W/LAcGQwJqb2eilqD7QYVM8NeZ6vXTsouVBJVhtWaLlNQB
gJqrP9dN+MS6rutRCTWc3wXyK9ksleqUJ+Hc4/ldlZJ/dffimgYdlRdPskSVonnT
UyGtVOx/79JrxlPNCkq7IoJ1s/Z41mGntYqj9R5yDfOUQzSy6oTV19vXd7yXV2CU
NIQ6vZjQeKuQ7ZfQma5BZWQnYmJ2m4JKg8JfJtezNgP02kmfVTbQHMYBXvhG5/oI
gdAMn6t+r33073fdrwiFz5sDUDzd7KbprMCuV9NGjiYy7K13Vu5ZCdHdDJKqyjmj
wQtGtOfr2zoCEEeMz+nOrw9p8Wlh56QlFTkdA5wjfeLSrBh1astaQvd3DhvC+R6x
wBZMPmXdQVGhJkT/CG/aB7+7AFpNptz3SHZxLGQRw/eqiT6+nL6sBie3Wfr/aWmL
icqtkNaZjYCCgXgIBPIvVS8tey6D3WDYwdMLDmvOAsvVue0gq5fKzPbAmlnLQ6pq
bsIOOdI0saSqrF2ShjVqcF8zqdrYyOcOv5cPir4pLjicBlTRS/mK4zIHjUDpPqBu
nmMrVq5AFWZSsTAkVBoQ4rl0JW4XuTRjrcXiX+tMC+k0sFH599xYk8MltiecWFMu
Bvjr5Txzk9CfG9CbCaSAvORdSyA0+qVoxW79k9LdumVxv4tz6Wip6sunlOrGeCVm
Hirrb2OtkGmD0PwkBW/B8h9Yc8vtkO3wgahsFXjQw8Jh4Q8hFQJhfFD+8VTuoB95
uomzfgQ42xdG8qqiv8gNmGFW5C/CJTDc+qHTuCwwcfyyHQl7eV9Kx45oaQ0sI4Ho
pFYO+MtRb6jFVbVmGhFOTpniA3l2D1PGtIEEDGJUQXClwG17ok9Io/g0e7+s89dJ
mBAAVQGBpMQxVRXBuQ5OaTV8xEoBoUAQlVqv0jitzRVY0BJ6NUiDKAcPIZ/Tobtp
137P3IT8uiLlL/kGobRStOj3f4t+VK641XguBgI5j4a2Q/yMglYMtB7qHOjHQOv2
CkgUBvQWB7mYRWkYHquB5JxLEFRfuPtqfRJ16WyG29gloVkhzlnt2hV8V+VWIE9Q
V+galGsMbz4WZFJJDg4Y6qNh+Pw7/YhE/AEi5c4oi61gr9fZsH6sERwhWSZOWa2Z
QriYo23W12cvkv2mGdvZcDJVXt9dePLciBK5hgiHnbCDCqgIMSh2Wj8ckP2Lp8cC
klH/ksx0VQ/CfcquEH+sZt+ScNBqFwrVAu95eKfViF/GivAX7qmObiwA7S/o+MY/
ljod3baGFl0qprz5VxZG5YntVqRgDlBiKRkcD03sZzYoR6jhPyy5yc7qa5Y0BNRL
r+Ob9EBqJlJikTF/T2M7zmFOdVgG5LswebaZO3/FLWQJb6NQ85pjaB+21phHaviV
eUeD9gTwH6DwwVD3vOXAuivL8RBl3IIPh8MYIHgwPgAIrBFgT+5QJlvDjwlZof9q
CDx121WSxUgnXBSm8TnRzM4ceKLtxUj6Dn0lYr7PUl/0MMCvF4BoGHQvvadzs+Kl
PumXm7Z6r7Hy2izb0bRxKZo3k34C5zCFvrSeldY+zSVMVCBSiG7/8X0j0NEpa+g6
U6cod02prpAgQwibZi4+uP15Y0stOUcC35zVqxyC8+g5iQvB1b7Fk1sWhUEvLO4x
siK+wnrKUOCtpSzeaZn0u++kUzdNNWPJwByYQKNascX4/A8Shix9HvKk+QXnZ9RN
0jLOX4Hzwx5uBf4qfBeQ1P7R0GQatQ4+b1eJIvQLzQZTCYwQEdZav+6GuugWIJ/D
/+QZXKLbRRmbrQko62hBM+COZEaf++xmOQFOe5SZ76dHlA/Z0jst1ENc6sFr5sHI
jMyj2RnLueMH6tQfRSzZNV9s1svAZsCHy+nPsmxkInFO+Ppj6sdzm+fvWc7jSxtC
Zi/ogk32KZxD2VoTZCcPSzi/JPM6y9paYg2HSAh0wUrKL5/Fa+jR/bYIGjCRgfxq
cxxGR2dGq3sGsOUClrc3hOwClAlR0+cp0oJ1C6EYWu4zbql5cgKFNbBAIg5Ej85R
6cHQEVyY9RMnFsZr2B2DHDxAHtaWqQwXLCmI2i+3SNIZpGp82HUvxJSIpxLkmc2F
30N5VYS7MZxJD75+LQenjtAF9ltPxrz0GGy03KwUjzwJaWQ7/av451wWC2bYU/jj
YgKuljpnY2ByYKJ2YLHkmEeAarEDJW4kHMlct6otnjP+nQ9yRfzpuUPxLrEK/+ah
86oMVRDJZ6/RGGdZeeJGxzqPhV/SYIKqAMUiDy7IUWGnWETAVf8+AQYapv1A2Clx
O+ZYkmLbF3HFDXZ5lU7yQuv+DSYw97oQoNe+zbo62MiVfiSONG8e72PJwb2xxxQJ
GLkUm70LbIdWz0WJkpq3zXOUTmaoVzjBLARB6y9J42GnL8ZCbI3Y5eUWCf2w+lXL
QRUTBLXps+1hqUcZ6V+INmpYy5W0CdA7BYDtd8lARKpNYh4sQK95H5E6PawxbdCc
+kWoVIwaS8vnA8Yjl9R96msJX972OXlVfS4bPenATXslLDlvt3bG6CxTCU/e9bCt
GRYkxtG5zD2e0vGjuv0GfUX8sAE1rKxy8D5kiithFffJFGv0t4AojITWPL4M8CTa
rqpPRPud2uAQICyPUtLK4nuGcg/PApElNJOCefZ0kVfI1S47rei0gZUpq43a6Vnt
DjwDAYWnqzUJRrHUYIPj7C5h3IavoO+NBhZYOJqGHuKGG38GimcasK/jGP4CR0sD
glu2N9p6ofq47Po+yK/PqSJYGK0he9McOeUCNZUfRSgaGd05H+hAFG0QoZxWPF2F
SiQJRpLmnahIoo7Tu4cLj9KpMyDz9VeIvlnBuYXZniQSKYzx8fklNQeeBOHVMgKs
DrhLo/7/qo5ATAM/KR0eog2/aBaVGFkakNb1/R2P8UUvdKl2fmt8gVuI1eF7Q/hg
Z6WAJqM79qy0HC4nG3wDBr3z2Ir43O1RFlAyDP69LXdDCZwmC3Wq7GSq8Noxo1qh
MENMk3haHbfp7orBFPzfCU7qmC9z/NiTmFvk4IalMj3TzksnP58FgWwXhBxv9DPg
K5YFsWQnIaLlbjGC+fHNtoDbhRnhg7BWiHpAOAN6VVl/7pjRroDHVeSSYSlqxf2H
e+RBlNAYPuxa1fUg2QFGO5xVxjYKkUajxgRic36DXpXzbaMVMGy3/VXMe5v5FA4T
xZxTfSuY2HScK9GNlCljfQ7buDK6lOXwhwieCjiL/6PmZ897CS0w6Vgo5+UK+oOx
0MN0YXQqXMXLpItLFOhrw0ytTfe/IMquT7Gwv0SG0JHYlYuhYDBtaRfqdjk9cdAG
eFAq0aDYAixc5hgVSUJGx+BoJZKcqoX8K6GS3KYIypfS8Z+0n2f0KfT714AMBnUY
JpNtOSIV1K+Nti5WGyiP8uze0INHEdN67hKZJrJlGpyO18QK+e6IKDbMIso0R494
UGA4xlCd589aAVWqFabgSPa8Q4L7XDTEbVSnQpfTydxiRfyL9LkVS414hqUFx14D
AlhKfgEogtJaxdKhBTnFnHfLyCQtng+iuQ/tKlt/tkO67a6M6su3L9y0Myi1/7tJ
vFYMhI68hujzxwEUOINkAbBHOMlT7G49AMvOrNviL0uvaIJg3MHAVb9ATZFNIv2+
4E3S4+0AtVHTx0Fmrytj7cA+R72QR0cqJai/pIYGdR3+I+nTsD1L3EQGbpNuLePx
IsJZ8EOn7d0VvFmqdEBgn2eDpf+vH5itSVqhGs10xh1AFr2t9msCdR4ETp4x3M9S
RgANzbTdBO3VbRCNa6cghI4k14erRVCfjHfUTBW2w3nlqVIvZL6DnBcGr7gjvCzI
JRb/ovBPt9v3HwfK2geEb1UOO9nTiB7JXFHWhxFUtV8AP4opN7A8oo0UB28ssgzx
yHM4snbgKoXp9+0h+9oWiONBWYNQbeXwnrcu2ArEE/ZvLO8o91OmlG1w6C7EdiVM
1/N5PW5yRECc5c468jjWr0UhOskkM2GThIE7oqdGQbLT0G2eKNoHGciuDNqKmJYU
296Xm1MWmCF7w86+XhFesxhb+kNKEtvwQpkWdulx5bfEK63SVnZKjwn4PH3bOfyC
Wl6ziH0tLI4Wt5OPentPJY+jxKGK/4gv8uE2A5v7FmuVevBSrx51oCJQoCTM9LTP
qo/JXRyV/ID81skYpIq2aGeIN3eKLM1ry9y6Z5HKaGarHp0dfhY3VWK51Kpn2HZo
jzlzVCZgou3RFQsptOLIn1/o/pfNkIshBweM1/cxg/Thm81oHcwPV4caWazKQSJw
jOivw0hNUDs+BI+bW8F70d8odMzyFnHHyjwuF34C2qAP9pjCinxRBDbpw+2Pwd60
zNN0oksuZ6nUdX70ob/ZXvrMgoipB5oowsk8KRs5oHeMFsVZUvMu6jt2PRMBWFts
WH2sGhKis5IGJ+rV1R8u33Zf/NtIt4CQDMsXAdI3e+C6/UR/EUxkTaDp0rVtoIlT
zZ/Q24M8Sk9bGXmdJTQ1ktxMsi0o6mEXwRuHJ2zEJKwCBRvkWhigA3Zg8AR36vvn
2C5a8gtd7oFNmiy16y/bXhkHc5cizwmL1LGf5fhNnnttKnfht/CcSZM9cNd8dG3N
/c80zPsXbaL9WoV2tysfgZEE9NCct+8ItYPJYaWGV6r0DAeX9LBzKiXzkAiMtkYm
mmr2y15KkIZ+yMWMsSy0N58QlQLM9P3gEjU/wMlhnqIEQ2+dmY1UeX4ky9ZqHDsk
YkIni9Fa0xhTNqwU//LHP70GGVGv2j/7xtcpfkaR4K++wJqEmwPMzMBbQ4Bn2e6L
yUH1Qzv//4lVeK3QHa5A5C9BfvAE+3Cap1NjlXAq5GVTvIym1sn995t524qAus1+
PkCE1MEekdB+Vccox7kig4UwaJYR44tGwCZYLXYDXd0N4h3Hvnux88VRP9PsEYPD
J/2D0IYBYNpf+IHN3OsYWMxkS81Ztzo6lRJoQHFum1Uo811fEf+bMwsPT61RJ78N
Pn7uVlIIIUDB/sUQHmAVIaUSSxVlDZaQkN87fe/eqtEbgLzymm4M2KLiPVlL75M/
SXIpXBB86CCIMJrPIzKeKARToFoSAFbYe9/r6ckzfemPPCFOAXVHT3CniOHFLcIm
Juo0oV83wBhmrCNOlKWM/6L2uTuSH4DCJr2hNX1sZpP5Z5YkiEKfxW7vJ1A1wk9a
jGij4X4v5CyYeZuPG937sPkTlDpNC1iqekBMgwwczVsNe0JeOMzA1H4pS0NN72By
BVzdPqsssntTO4H8YjzQlWqdSdxPjERwKVA3Rx1zG0wyeiEU28BE9WyzyAqitxc7
VTvH7ScwWZwF91KgGWZduG5rYX5aneBcHSFSXlcP5VhZC/TeD3acr/Yl698TzSZO
5g/VXW9C/GcdIhqxT+Xz/Ajc4u7He/s5kizAYP4PkycpcvQYSKoBZsXMj88qRIAS
WXxtfiT54rUPsMSjeXL2wq7xf6HX3OYOmYt8TKk+2mKvOQRyhLaWRZmWHThJqH1U
g8IecGkUb+WFBCeeLsRuY9wwzyyuxH5S1ec96KQOQuKTIJX6MieHXYqJr62JdpLd
accNvCKCdCuf0R7jbF8dUMxoxBqCV9kDCUUq/Dkqq8v7Czw291UqWHsLeUNgQAEn
3beTqQRMkqb3BWqtYPlc1wLEd1MZL0wCy/5K+0s4V4sZWmf5xaKOwYP1jnwNzGux
beH5vGc6+3gc5dua92bAIqdAOSLavMxU8cwN2090Q+a1xLBa9f90k5oX915qC8F2
yXsT891fEOylL0D8IpRI17kfwbKJrwSSKELPoxf1LSpVdwM92+P2UD5oJKq6h4hB
GeU4gqr2sCZ/MkqKkEA7WDNIAvzOFi0jvNNFBZFybKvUMZ09rhzrbczMg5t9lOV8
b0eTQrGJWI/cUmE0NPuixkWMkydtVTh+TiFeXOOotLu0sjovecHDYFEnv0FEWQfJ
+yEpl9nfN84g0cBHUygMUmXamrQGnm9/Xq7wgohRpPj0HHq+OgEsm5+ljrmoe6BC
WHQBfnk8ux7MYDNuMuhbTiB6z4CZTpatkrj2eUG3NW0XWNUCYc1OuvjD6kf6qtPy
KLbBPInjJL7MAYfUHUqUxT8hhSl/VHgR6cxxG28KNJ5szDzOfAwgTYubMuPWfnCP
4e/3ZTZ5Mc/iCXp1V9uwt8eBgeoydXslC23luAltzNMW9oM0t+1W8nHOu3nUNW/R
a3Sd+rcTrksQ2yFzH+wW97c0b3deiHwmvvLARaHYTKRMOnezhV3DpdLIEwLcmTf7
/0vHfvmxJ4LwEwNoHa/QGHQXE9YLWp2hRcm26m/49ITV3aU3pTltNo93141lV61j
KKLLKhiVYJdnoOMDBopxpK3NEQt4c3GO5XX1KbENv01G/0oJ7NMFXr13udFgOuw2
ysEWJzGeO1XCsktqULwOeCIveg5md8bvGekwdAcF0Ba2Mlj9vt70+sS9TpCTHjPw
cNvtxqs4xmXSHKNgXIN3A7FhTbjndnmPq51XqTvxTd2Wx1QkUAGlQh/FV7eUPH9G
O5mmPldtOBsOhRfxr18dY1VmZsHWMTaCrQapT/3gPOn4KE+TFTRSRcZBcUMSO8bG
N8h43msB2qIDuTkXB/BKfpBD1nahWE3ZSar+Zv1qRWoA/0dW+wOUeIK9a37Yawa6
rvF6xEbEk2GgKoaLjZS6qYCCa4Suoosal0v4DsNMmCq9gGqVaBh3ENpgJNY1+H/K
AsLpATtuxXsv5uSVdtcIJf8fZboggRHG7Zd/KiBS11uIv3Xp2C6xZUxssJCLqknH
yJ8VStLTFfH1niRPrL9JWHS23m1jC8JXe8CKozkGCPF1o8/5JyhwMfaUN9vdtvwS
RnyOx1Ot00QXIgvTYz8M5m5PPPRJpR54+VZkCX1uO5gMksq9BxD3PrVdPglt5Yh+
5yiIRwbdzKqKJnayQQMdlfw191oL+drGGsW/clKBe1yFBtYiZSLXX6IzRAgn5YSs
72cUTkofJtGBsvHJkvhhU+fLGtXq+x40m6kdAOyjf9q/uW4V6QEipks3ltpXXIbW
+vkQTsdm9l4xsqmMArfLp5X9OWw05MooGsucs/PcGm5Bakv4s6YZxxnwzZicDhiL
/ClscdEraR/+LX4PDAnwGRSzHoe413blzR/v1d2f5x4YEN0cqLqmWB6CqKJTdJCT
3Q7mpI1gczro0bda5SkHqMPv+Gbq5tqcQH9sTVBuAMKE1djpv/GplLLOPyW7TUvc
DPsoyl2lGw3qO3lGLunD2YeaSnkWgBlMH0zLE+4OC4n7cIg1Ti54+tuHYqK1Pg47
TuaSVqHBrlYJst5tcqgUrIWJJLAhE6LSjks21JFtwmhCrCHLTYtxBKobpHw9mDTG
TiLKxCkRIdrSDTJid7l1LdjZsDkENuKcKzkb0pY/Yf3kcTrpJj/s661zrOxagoWK
mjPDQG46cJg3pe1s1jbxA+Mbe+PFzsIizw4JuPBcMCjWgm+EKv3OqdPgmS8LbbDg
XSop4LDQlbhMmEs4Zr7QAr0xfZ0iwENO/iC5dMoTXQIDhE4RuQP6TbRNqrVrIfUt
DLx8ECptR/wZrJMPbpcVjRhpZ3owgEnmBZzrcfefwV6meQotBGnTj3YdnPhiI3Ln
AGGAlDch8M1SepPJStvy2/g/KstNoyVL+Vp+m2Lu0Fu+dIasTHFFrshpZosqyZVL
WqKWK4kEAOE1jLKrZSJ+g26L8nISbw5krussoPUA9QcgFtKmdDSDqYYbdZqly5LK
MC8o1uG+pkj4auL5essSv9rU8UoDTjwM70CklS2RqqKyVZ9XTJwWkSAvqHflnbWW
efMFzBymdYmGG+R7WV49Whrbpt9mpw9Bt/47CmZrX9s5hrh01+Z5Nd8Uf6tr1EaZ
RxNyZZf9KyW4TcZaLxqc3ebw3t6e886tSzl/va1zdLJYDkcP1MWWUnvKBfMLS2lj
qKmjR6lUrAlyFvPSRcKLA2CkanjY5+2NI65IMgExHgmRAUuTA4yaatrQe4PM+wcQ
uQQty+I2rkRRX/T0LsUtNeyrmIDa+VJlsOd+1dkleSksZMDAIUkmRZkcJgU+GDn3
u+bBS2aectxNyg9Vg5m9bcsE6FbzmVAGspQmIFm5PHYB5NK00Xae/A5KALnnKEC1
C/9U8cDUaClkHRZNOOKK2Mtyq/aluiYbii2LuHla3R0nPXEMWiCDja1UcnTr7MXX
Jbi5vgurQ69C+XTzIveJl6LiTkxNC4zRwCKBUSI+y5EGxZPlCB9Ef8AYFc8fYsjo
ePb2ZPXoN0egEdxzN0EP8DMl82VspDnBWHxRGKr46q36EMQdyzepr5fbNHkwOOLu
bAzjgrSksTCppUYrNHx2xr8ea4kIdcZxv400HAMQIGgKKBRvC1AOusv5I6re+THB
x49inmEG4KAuSkfMTuHG+TiAGq70xk/AWJ7hp4diEvkauQ0sbPNkTPT+g89mB83Y
Mqu2SJrAcbEwQaNK9GgavcnmKBzJeNFAOaaecTGu+tA3Ft1d5oZLSY6qy5STrxxH
rY942wKsrmNgejrNueTH0yOQ2jl4kTokbdxJHW7ReEnUyLZprAwM0YZlFYT43vR4
j/piWpoAirJnZ97E1PKe27MUGaRJmZP0hsBEatzPjXjQIdvsbX1xuK5Vhfdd7gQb
bMcWVj0A9D3QisLPO0PyahGbmpY41ar8luTfbShaaVokytBj8qkU9D+dSTJZsEww
qTiRAs1KZ5LLunC6GFz/DvDigxSm94RcybA9x/STSouJXBPz2ybHAHUrJw7cNhPJ
4/wCuvLgOvJYff70rTIET/Ws1oIXaB2l0x3mZZsWnXbwVGHrNtPnBzDOXHmLENKR
ObA++x/Ki2KfUvxANAEiPqav89FHYvvxUTnYBglN7iGWxTkJZ/fVaEz3zV65FsLB
yK28FgmdKJGZxQrhWs04ApdyVcTCnGr236a1eGiZgFKZkrYW8verOYZJ3hDbrZCC
rPa0ZlcTs6Q3baHrPkqSiAs3PgGbflwePIIg51CzhvJ3Gz486OdtpUfMJpW8Nu8o
gxCw0E6WQ++Mwd7ViE4xFoTE0gyzQZpuaurHTnWCo3fhf5sjp/wX1lSlXVqtaZIj
mMFA/dxMwRJzZ+LCdRc5znPGzJcBvTST5wBp1yI86LBCA4bT0h/w+UqtNph4Pyx1
5cX9Jl7GERJiopgovPJ6QrXyiBPLQJrEBB6/ixPnNke5nypw1+xxoVJuTAN01/Rj
jgP0+/96jszHjxJ3ycYbVJvY88DsN5Sqc5tKDCDE1Dm8tyyMvKrR5oqhvqr4tUNW
3ymtZlLevviMBOttncU3gClNjCvGxKN+1HARfVsTQXasJAliyN2y5bb7DpYl14yr
iiXWDnB6x4dzfZrSnCXKYTLWL0vLgaiOVvSleQX8VtvLwGunrJgn/MSgAvtaYEDL
BitODl2/o3DzyKTi5gQmhHn7ObcyMcpzzD+CvmxNrBui1EX/cxGrGcKBIjeSdfQ0
zC4DsU3Y7B+W7hdIHTgtHWDu1uGmPjCjyeK/WtKwrhmb7ojvIfRuau7B8/DqB7O2
J6iNiLnET3Qs72PM6Z0O3XrC2yjjQh2fAtnWoSO0mq4o16RPhwtPeYG9sj4Q1KbA
92PBBlNQGltrR/1irmhat4SwUhUU6ixJ121QngZActHtaaSHYbqzmgUaz6SfWuXm
uMfRsYFrdVynE51Mn1cWPQIWM8itkGJVl4IffyDzR++cIVF/jtL5viSsH5MhR7a+
ts1k2AMhhkcYUN1+ebEYgW1QGei46jePuDK8mtXYPPjMlu9f284I8eAk1TXOXB3c
Wa7Bo4ILRm/SjdFb5bFfSVo5lBJPp/guYPU+GwpeBvThEoz8lzSUsefL+SEpTjFq
Q1abhznY+Ekg2tTnNtnI3bIyRGepH8zuXORplMluDu9vK9Wh274jiktIl4E14VU7
YifUii6HnJB7Yqit0TcmdrSIrQR1S175W08LN/5kJkwcvdM84R59LRsZLw9oGql8
HK2LD+u+OmyPgZ7tKeep1UhGZpRjXkcOh4NnN1yaHCZ9VT4KBrvk9VEWXgnT8JHi
5wFZiOI04fLoA/OxmzjRd2SmD0V1+62Df0qSFe0KMXzibX2rLB/oHY4QzFrF/NTk
tkypq/CE8bG29xc9Srz0IPXIKyGFmvFyEa4yZu6GM76n/juYKfm9cjoAVFt8tOZS
iOHeHiKDG0wpMBGv0EmEKF64eRyYTJ+GnLTY8hZmko0BkIaVtcxSOQ/9Dj8COStm
4sF6WgXHKC6xFmT4hxBk4YdGRHbMNG8haZ4q/TumpJMKX0tIH+v7mo4TQeqi7npx
+HU+yEkswvb4mNykpTSpNzAkSRr2WHdaVjNRfMUiKhOe+sPsXBCWsJ7Z5apI6KUk
x5ecqxZu37Ik2vH36ROecnCVK9NBj/7/U+oBw9U0FM+IXt6dB7CqikIwY0uZ/0gR
Cm4mtceeZ40gcex97/Ea5+gqj9bf6jokQUebiQzv1kFOi99f4sbw96cIZKK0WrbE
P6kF+g7lT+++qAy16OcZnIQ2rcDS9skI3JWxjrFxkZQvVwy/lIVc+aqRdjMJ1yJX
J+DPt8arFc6kGWwiUS7WP1otmdMRiUhyOrMwt89/o4pIj8E8X73Aba5B2ChrtQFW
DTJJusJLbs2OStbv40CkI6Ass6YW1tnbtECssq2mmQrmGiP4fam16N7zO5wDnyIB
SfnrznqQqEX3dzna4fxFES+5SvSV4g4coUX5cKiX03Q2/CyEqhaTZYOwcaHq3kVd
10xTG5GXaeOE47xzRh/PL+6RPOMuNemDHzcmrnYxP0Hi0Sn1SRc9gB3o/qZa/a8A
mlSN1s+kyFIL4FIZBEYIsaeFus4DkkbYP9J43WDqKk4PIj5vL3VaXKTTP9eXF70w
8mFMM+bflzSRN505ugCUjgL9gTPomDoyHdqaHWHNGiXhlPVEBQywpH0lNPyCkDDi
DSt7HFOglTtLeFJmSb0OitgKuxThQGvzRPfcG9fDK0af7Efgks+YfXh32tcWJUZ7
qiHfb+HWVIxhgkVZu69R6F1nm90rirBkHbmVhgBBfNs3iPyhNb+GW8yDeNTJnaFL
57f/1DVFBDApQd3C7HFBJv5/3xM7ubuAqSD4SqlHO5pLdGc6i9S/aLDOxPTphXWb
IMP4QRUb6ykjwJ6Bne8xzuhfiCz5LTOHIa9exz+e9Eiet46M0iSugjpApI7cOsPC
DxQTRI1nCMEFPDiXnVFHKB+h5vPC3l5P2p3zwduOZuaya2ouOXOJsuBxhyQXLl+x
1SruwbCfLUTdiyVNfPG2uNKlA8aX0FtyJyFphBePJh8l+mZsmkL3H3AeXhLDU846
K8E1Tfwh4ov0c7unJlkE+wQE8jPaugBcUhjkLMj+wkIzTO5VDChtaBNQMZ0bIlSt
4paV4O6GfCf+Wd75/v8AVGfZkoc4Jki+W09EL3a6mAwEUNH3WaQcqEMDG/2YrgRO
Intc+21GU1ZUD4YfidAPqailaGGSo+tADTWPf3XEghxYO2aXMZNQj45/ejmrsBn1
9+lQHyzXJgmTDEH1L4HdBrkqB79SyfLqLOeBhwA58cSEzFM2Rgq8TBuyAgOueAzr
M+pcUBOTIqW0aP4HWqG0uYiDi5EF/YImwGOPg4W36dc1yOMjsdWZcJ9Nfc6aqReh
GinrWPqMPEDxCYPi5JEi+AtDB/IkiOzkbrfNPltL1vVtP/mnTDlYbNBOGT1iFv5W
Ugc7v3uB2ThyMCxS5RlvOAwE0beYve/1TI0tou191agir91YjyABZs+JoO667Uhb
gPaCSCX5e1FQuVrgAgtxr29w6RZy9yZtN7EuwiJ2Pb4E269IGzoJ5kjbHuiF2noQ
xaXq6AHGq4aBwXUeS1VSEermSRKAJuEA5vCLcvlIETMa9Vazd68ABFnvjPBFzjds
r4V6ofsTajTDTpfUMJKV4cX5yOddfrSAyl7IJZTGKrxJOOG4DIVE4VJfoiPzIGrX
6cMGC+IkzyE25hc0Y8WBZY4B/cJYqsUlAy0xookTBQdG2qvZesgty4Bo/aBvYqV1
d6uWlQY1rLbjIamK/xyl6ag8CyLAr7m98wTFdsCWxgQ1iQZry7GsPRnShAiafNQk
tt4MfkQJmwMFMcJw1oKb9+HQwmhlX4LpXW5eIRox8F5YG/pQpGWWB4clxOIZoMF+
L8WnH+k/caw+eoWUDo0DubF7efulAqfY5O957piMLL+0aK4XSrXpOT2YeEezZH/X
BXNxLR/U+Sbpw6CiVkGknwOLacAJkeMe9o/P1OVD7dycIpYmLFoAtyjR+zLYe83d
05UFRgWkbEC0hB52SdNcSlfn0qWpc1g5d9RtrtOvaqSxtbrC1UjucfIlhOYYRRBa
Bw4Izfi8bKDZnSB3hChhFf4AXJg5QUQh4ChvPZW7Z9eMC+wdmSXs6ls6LoIPa/CM
XhnQanFnsZn9Z+k1xoz3ZVTM6yR/ffpPBpJ8+0nZbmmILzkDi7O58cvL5h9wb11l
LJjCbXnErExzkcdT/KbeMFlUm3Si/E75gZMi60d8Ozdo37/Txck08V7MB32gTm+9
3o/9g+miAitL/4W7nuQCn3my/qPJCynKiDuv4HWB5UKgacvBIMvyyKNfMpzYhugi
LQClAssKWC88FnSJfymu5oErIEUBgnupg8ZfaYBsTOlUxboh9KHQzH/mJZEjfjS2
gflcPQEAxkWle6o97zGbjw+noNhOGcmDZGpafZCT5gZ29Ui1dFSedRuvbxrQQev1
MKtXbhLP+Zjp8PjaHbgEZQYNWQ455Lue4wI4C39mhSzn8sYB0/N7a6fWdlJGHrL7
EoKYDRWe1JwZMnmwcy+x9iTkgs+ov4nyMfVwRCCOElE7fbaWlrYGXDLrY7QlIun0
F1bomuQkW4M3wxVq6eEf612DdObDihhJ/Jn4LF68+Wo+zrKYUsU4xQuTU0hwfZrZ
sTb+8No4allaPiELzs282OyRNivyavBGF/5j1U9KEGFjCvAs2iChXoxHKM6xKD/9
fbmRqKgaxU8oW3oMkiTwAEkkjoVlCr4MxuGmryH/MPjJZEfkevpC+E4WRH2QHE0c
DFtrlrQMlm+srpeMtfOTINktXMwExdzD9dPStYA2G/MWC2NmBedwFCg7kSHB4cGx
AW3m6zxeFd3f9ggAlF3SGsE9f3n1B2uVMkkDjQn/s1vMthMTRNPTEWCYLNo64Rbg
DQR2KSMpY+d1W0blwcO+VDVUGIJ8/qoi79KMA8LPbOX6IuX0nnDcs4VvcQp20c9j
OZY6CcZx8rRKZnBX8n8Y0O1y7UV/BRThZxptyXwquDPm5PIMoQ5DiYlRvot4RSVu
ZIi5xz1gd1atL/3jod3739B5nzFS9u57Qpr6aKsIqqLVWNW8WTLFQLdhezsglcWY
agxe6nTcrfP4/xsQot7V9EBIDpd+nBGxN6ug/JpzGcnXeJhMVf1E/DlaUgBt7StZ
5Bwk5sIBy9d4SmtlilunSeTF978G/5NHJT9Z32qLo7ou3vFTAVi0Nn+ncTxSJ96A
0hu01WuJ0WVAG4fOgn3/Fa4BUNpCd7G04JdJMlH4WUwPwnX9KkjLZyL4jUowPmz6
XumjEiiQdy98OAKqf4UKElnAVCChsx4sDSuJBG6kvOy2O59HXPOj59th5i6jM7qh
/5A0m2Ye6uURIkVRll+f95p73F7w1mgilpAUrpXoGz7F2zWC/usrzfGDONoOPHbh
fX4V9A95HgfiBPnogclbs5qatv/4ot7a+YQ4AjDHgyPrD0MhSsDZTae0W1bRBYe4
clioJqOSo1DjfCYeO7zyH3QQRpOw0yDuNxe4Lomg/L7/hIH/cdZfXHszqGOjTwPC
gOwJlUBwgsDZ4XTWiFn1SeE0kGzFpllrOtfQTYjx1b5cRsAROxhb9hdERuz5AG6R
ZPnb0Mt8tjwP98i2pmtlECGaBChQP7FN/u/PZnx4BsIkfWYp+O/PTgFLiw5yliHd
8wuLwNt9EiONkW6R0gVDvmCcNJ+zoetCUKrQYXJaiIcfddK/cO07NSmx6OwxXRQ+
sUtlhQDU20hpZnWzPPtn1c6xM/hqOwekvrKKZM0DRiWFDI1CSemKlqHJ6MXI0wOw
R6hZSZmdAATtkhD+qcyBEsDz7/xG8nQbj8He+jGqsQc9z/vNZR3Hun1Z7GEjDWq5
f1jWp86R/2PxIAM+lDZy3nL4S6J//UAWaiq0IQ5xzfyng2/MCbSVO540z9PC8GfX
scEWkC09027n69BhI6PoyKwAzWSfeGyczzkrQ2FqaVO5JR2BVVA31oyTIsSWJWNR
74YvE6RZIdgCT5PJm+zpYThfvkio0fB6NIcVt8xs3XW7GVN9/RM/5I2ZjRYCGabz
+7efYmYHvVV4oowmxluQv594c+AX7L5WYk5Q7KjvrrnuJQbse6F3uI5X+vJkGV8R
hIBrw28gA77MWe/iSZc2R7yjq1cAdtk8xYL2ozMC1/+2hre7QDUpPFY2MIKWA8EU
nw9/zequekxMJuTmUSn1yjMWBRMv+0iXZaKKZxZAV3iJt2K+naqXnuNld+yLX2ge
g/q0V4yUHD5wlKfC/qITkt/+x8wAevHMvlmhNyP5FGo3k0/B4VIpGa4eoDvmPebQ
JL15R4mr5tGQhbRRFXJJwuDPbeF9Rj7AXjnm6EJofRfD7EgSKeIw/L/kpTut+2cU
90Xu1+9GRrVTA81J6614ChHZUSqjHRNhPaLUOnNpnBjcNGWaE4Rw5Nmn9J2ey2ok
ebYxM0+i0WDpObjyAzwzSpRTkdLshfgAa8ZjxSZPAhC/TquGe68VhepkR44yJzR6
Q0g6ZJzu3C/ekEvjlg03a2weTsH2HuYYsVZQDEPq0jW4W5NYT0A8u6EUqhFA1nrJ
3R1pNhCxdY4SbIthiSToDBT0bgHFCW6nal6Asjv0fHbVjjKzZ9JWgDjIyaBaK7Tj
TjFA4wuqCLvK3dje38X1dkzLxIyCswxK0avSwbbQNojQGN6Wnh0s+cxSP8bTIOLq
HvTALQnmyHVjU3/5q+T2r6zGHV/vkOhZNcFM4FBM/v6qEjJf7wd3O4w3eFfb1kPh
xSj35zUfJT9MwIFhy4tyWusEXDT9G7QHWbPu5HstDxoHKMnduhuPFyNP34DS+tkH
aA377eQ1fBRpeSd066/dW2iYA0nzpur+FFhmnVDUU7tHBgc/fb89sXQN13cvBF5T
nOOMWPooGOP0RoJSPdyC3pqv+tbTPFB24tJz5slk3tEb/7kI9e66YdRL+TYusV+Q
3jhaWtIT4I+evXI+LdWZVGnnbKBsat9JvSpNwlfC6893Ug0bT8bbQQRoEtzjrZiU
7J/FiS0FRqEoouITr+dt+/friWhVZ/tWIOPSqIIjmgSesUJNV7SUW9QLSFD8l1Mw
12mJzBTDYvSOTnLEZc8QRFEFvM2mMopdKIzdjdGmDMw3fgLszCLn6h0h6r6w11cX
mnXzfR/sbpYjRrIFJig/dWl68glQarQD2JbVfwRfwIzsJPxLP3wKycFYCngyLtQy
+/ywUcnhz0mtyV/GUW5SZgTHejkQxfmDz4xchPKnHmYb50fhZcrB+puwE6h97AAt
CiultmIOPg+Gad3wU5IsuA/0zR91Nx1FHNpevIod1N4ABRyLGEp4zMBN/7fFwmfO
qey+pJQRkopQRdgCKNHoiobx+QCIxYQbZNyikPJBynGJxQWOEEV2KFRkJiHhVS/O
JPpokvWoqv+JFBBDA5sFEhOLSxuynhtF8AyTeTJZ4QZlWjIQDjDUWh9MYwdwl6Zb
pIDjSybYBPdxtqnTljPEK5wKb7Kg4O8zcEOJK4Y/E9oDmaXFbYmS/Dhk24R+gkmx
fPQFkJ46IaV51UE3Hr4gc1dDc27DcHHxXscoEWuKeq4kBLfptu9njTmwFxaKYyGE
eeESuoo5xxenAc58eVWaq9euNK2mowmmy58CDGtbNt2d2WoudN1HSPyB9cytXYEF
9kTBxc8KyAc3t4uyQBS9izaoB7fbxL/oR6RfuWqp3QWuyRzbfn18buxP0IIG8Q5N
ubut/osRh8s4hSsPWwBKi1Iuy3xpeexHxTkkb3+UmCvKzLrLTA8FBVt5pLoVCi2B
/eFv3W4WQ6itYfHofNu++TKXPRGkrcmL4ecXlS+18wvtELrZoHT1/FTGjh8SxoKV
0bC9EGv0h1NSqls1kXjmt0LmAhVyMDRUNtU3I8+7xhOZmArizSqYUnjjwGWr6EKh
RHaUcCHR5rlq/CJvBFBzrpXY1dNqPaMUqty3eSaCLFcOjWrn236bBIstlUSZw547
OzsSuG+zSlo/Q1LbxKsNuggM42tCtOpmUrAuZk3bKf59bYZYB0sx7f0tEMu3mSTG
l6PPnC1oM2Qx5Zv//Y/QulPTamvBes7RXsYwZ1NbF6HpSHv6DIJawlaP5Qz4qIdV
HOQfMQ5v0tnSf/VgL2PW1UunfFjIYuooMnPbtf5r8Z22V5SQ1JC3NrzM1VangzSc
FKAJ+UuEcK4eJfWGzixN4Fe+WVSJbbYBiHkiH0wKTaTU41qeui4U6FiAcQiOy1lA
EdAdY3efcwIjbcQ+RzEKunY7iAfFgS5KwcbbqzmrWeVYwPKVYH5iYJrdYxSH3l25
1tQWwL8g+ANjHY0PqOLgOUjOkqFOvoAT9m3v95awhaCCj3rtAknRyMZr/kko7yRs
nxvJyxbpy7p6jBETwjeHiMSq5vnrOkVu6dqLDRRyJO3n9Ml6tKk+7E/q4kZVghJ2
ASSRz6nhBGmxFx/LyHUa9aBLEohYhKn54zzBSwZlxdW0C0qAoFPj2ItAo0DIsQ11
8m60I32EbQxa7qENpC8oT+ZrzAxFdUdxCev7pjR4g6XVp3hq9ijVrTK9YxWm5+gq
Tc9kGoZBiSLRU4mNlUnn+HJGveuR303vMFcRUSV7OAa1yVQsoS9INzwVWV3Nh56G
rUe+WBhO8S0Wkx3uU6t9N73F3h8ePQMCHIBhCDxpvLHGpRJ1PJSOHeiXJC+B41jj
DW+ea/Mg7Kx+8LHEcsoBHKWRF7hkPAIqNst5gM7IqHc9lv0uOZKfmDSmb6leCiP8
OIw87/LHuGIPT5fJfoZn/4e9ObJTJPMDv4YZIGMpRC9l6/L8+2VhEqMbKwDQQ57V
w+4kZKhIva8czvtP1bljapMVN4cb0ICK/+BSfkhFVzBobG8AXjEmtw5vplz1qrde
O5UOA229i2TVpm5aVR5AyYU5+C0FOnZ6w8GuWWF49FltnCPWcglgHZ0SccQP1T4z
vbV0/QlgRQF/BqevRew7LVB/mmOq1k7aWrfHaYED7DyTrkCOkadtCi2bsffkYkZV
UuBlQH1NlHgpXmOU4pNUIMn4llsh2L5SUNfM9q/zk2JHf7VZ3kIKcSz+/6G5XKm+
h5a9DI6zr0MJKqGDgNSMMzM81uOQsCrI3X6jw375neCqZOELBN5uPzFUTaddqwY9
AQDK+FGDBf2OYPejzs/hx+r7cBXV5FnyjYa2+yk+Hf2n81kqWvZUESIuJ8f+uoFS
vesxHku9L2TZcc9G51xEzqREG1SfTtCz8iAK4zk/QWo1hPsY0MfU32+L8r4o70gw
1nvXL6E/E2zqhGrbaEbIsB2mMXM9ybv8NcHbEo9b+iKI5FXmnux2leHJmfurGPBN
BPQaAgOxWE9OtXqHhfcQvDUaY0Gf/bKyA03J/qEqAFMaf5JANWY//IGtYtlakksk
UuJTSaHL0uG6s0TwHefP9iZbd1arno/UmMHkZLj5ZSkChe+NYDaXe5eak/oiUYSs
kdJdHCOnezwb5ZmVDSZVuvDKCTTGWzr6VhtGaRpNCGF50oMfRreW03EuaDr03u9g
72FDyCX1U3vVFOIX57SzkIsP1v/EtSX4+Exu3Aucpg9saHeo5J795eyYUtzCNiko
8ZQCIFBBLNEThUJ2J0UBkvui8IUWSMkNAUCfpiXmFm2ujv2P3DeI44QEqmuKOgTw
ivP4OZUP1Xmk+JSWZv90tt+VA4wnCKGyjXMLOuDq3ht5AigfPRdKXTFRq+ettFOn
7AVhSEaSp/+nLSYqUA5LWkZvaH1ojo/7qDT7QBb68Kt9UFuSTpUZZyhozhDXDfUH
LnQJmOjUFXak/1xdD0YJfQDFYQZTsh4GOLIVFcdgnbq5c08GAJbXKA4I4AhMPxDM
hJI2o7EOqIN1MSGxsGIleAgZdZpcP9QTCOl0kZ5hp2aLy1usUz8Zj66yDYlbwK6Q
cIB3sbVW/79Ak97Qogc58RapiXv8bzH1Hj812PXLVD6eDC4DxMIE0c9um6d8+elS
N/04kLrLidR78X7dR51FVAOtE0UtDlVz133PjwKA7muRMZw1aVphbeVKkRAyiYmi
QiF+2oGQtDEhfgE0IIeAmjLgkAIUHgowcsFpeT//QcNn3G0CJDKdUFQn8WsOuCPo
VPOI1FayVPIuB8AhdsJbLksqWhOXIYbwptU8W3Wr+2FBWt4hsjrpv4YPei6n4nH3
hUVhg91lDq1hhMX9JEn/PzxgPAVGSbK/LxsjsA+6PYmtq1scGece8Z7cpKP935mL
zUq0q/kIsHFlmnDnBiruh3frxsTyPAwoX+SoYtWTHzy7Wo2bPYu16hEMaya+x1dx
fsN5vIXvAf7XhUbK6C3lAOEOFBR5OkSh4B1R1vpc28W6gtlMpyRH5msCD4jnftDu
9B3qV2i68SwPRW3+gQ8B3dpKbztSfwy3V0DBo4dWlz8QOjFOSgIn0wcuRT/Ki6BF
S+Q6upQQKrf3eogTYSdSdBmLhPnrBkYKxres+ouHHjcPj3Ei6/rfll3dExOE++UR
wTWCHM6q85sd437X8wsrhJ5ZHX+YNQvUBY1Y13diV3IB60fkTfnRszz1aCfXvxpc
AnvBT/WG/jOzaJdpEzPU5yf/IRcPucg+NLIL2UX5jZOsizh6efwTVrTNlMF4bmPL
mNE3LMZKHwROJUNHihVbnUCvAxlOVaxUzfGTCVIS+CPdkyaXzCncO2s25m7pAgeI
zMkOjfifBVb6kPJrvVR9YyYc1NLzP++tpmiReTfHaFqe2Cx5zlZIplRLbYo5Fyr5
9ZHJjWMigz1oUpgoPzwwoshMugXZ45vDAZW5JaFnRs/Ko1u3n2hFXCqCFtuIoMji
IH0vHUOpLjGq41WUvSbU8GC9SdRzInFXanyk0buRvGJUCne/r9IA+5WjcsZxsVgN
ecIEhAx56k78vY3PyaWqX8tBucLW0AF1fzKX13FxNsvaKiAkC2ZoSF5oohq6Bpv8
ZS9LOlvberbMRxAmi9yOm5HHTs4ng8zgJR8mQC2p+mvlYvz9Zw13QgiTNzra28eH
SShnchPBPY2OJkhuQMjab/V+FBUCHz2gHNv1BR8pwmbTL1pGPJBi7TUDUJ/h5hfv
+KXFienWsZTs/w4tXoigJitBmY63KDLV4UTLPNJxBVNkBX/W52XhGdhMEh5TmYGd
sJyXb+7ubo2C5XFPsvZbJ+qnw9bK9zE+VCabPSQQm7Oj+ZQSaNdT0/dvgeKxx7bC
H093xw7lWMCK16CSE5W0DNrbOAaazhedLCOlRC68K1HhC61G/i30xsGISm7M1h/K
7WbqXlwm8GF2dO3J8BVnz8Jko21SEMM+fREMPLMs6URnNvRBLPSyCSgw6obnVBTr
SBiohhb8JasOLCnGx3NEPe4P26/7G9gl4ujLIBntM0sVUaRUOwbIM0pws91oSxG8
neirNQMSDj/aeiM3UHNr+HdGuEGA3uCvD1TPHpiEq6Ko2CYXvB4Sso6KAzP7rJld
+gK9Qf0RWgmIzYOsJnaoGgws+EiWkpNnrA0SCRdyFhyK8GsERZf3gtVKUG7hUnt0
4+MD23DNqmZjJejk1xuCIL0fUttWjd9dRxXfu40DwzdV6N6ycgmv2+eBhKGjyFAK
tKLZEjxZ/X6e/e91+lDEWFCP2YkoJWf+7XtahE47NxxAV5H/2cAc4uYjtT3IkZDi
nBFJwwtcd+6AdWnr1f1JRQq01tar60dLhhPBiXZOhoUcYD+gmwYksiQ+semurgSd
zl9BnPhAKQNB7clWx/JMsPGkYMOntJWNxQk4t8UJWK4IXE+DVK2Fzi1m+CMXV3na
yAWD1JAMacLzVCqbNLfnevaMtnDw7rtqm3FV5FfEzjIlTUoQHyYz+BQ0gaedDnKm
3dJ72d9xNowCrC54I9WK/qlrY3lu3Ez4pv4Z4oM/RPe5QJGlBx1PECtXoNrsScst
efj5H80J2Fc2+eRds28uSiAlA3bgyo0rSCxxGPaZfwOrV4laJn0x8yoqL/DgkJD+
HkbNx22nUBmV2+1/SXBib4dnXZSoHLiM4QCNK/F1CalUl/Hjd6JZyvmv05vjrkBX
JL4LM/9weoWEcj2cNbDyi9zI03L5i8EGo0J8PshlPbgm17EKjuqZYU24FV3ErURv
TLY4X2uJSqHQuuAaYLHEZF1e5wq0TyxgbrZSyl6Ndiq1mdq6jdDky5RH2YoMqPF0
YUEBBJu76Ifxhi1MbjSE92O/0VRdd39t0QPxJDt+/YSPnpaUD4C6Nm2/uhQpsGJl
b38MUomS6RG1eabGPvMTnYDa9uLyS8dOwF1QODgRP+X7oZaRMCwt3GTtrHRQ+6qA
Yaye7lOQH14V/87hwAETbR/6DlH3f7BO3pWP+ShrCOfyTCGm9dPGbfeKfB/OW1tp
CliPjTL/tDrrpUy+97JKyPF9gl/DQud/4GWuupGzh2IihtUu9zFZEk4V9DDM6fP/
vQxaCIEi2akuZsSOI/OrP/hyORmdagk3+ocv9ol/yJ7mUr5SOpU4EQAP6/8Gzn/w
wyV+50s8j5+CMx2ao58h2Cq8DeEe4LvTGDg6BUdCCN2pae3YDHr/N59WbwZPg3Lt
/zqZjkpAwTJH1QbXZVGYF+KW4woG0RjRmd9Eicgsc7fIpdwu4u/TttyJ8GLHI9Q7
knaCOllf9DWDlXqLFLBdQJ7pELPRR2rXupeNsYRd9AtzTkx0FQokHReeQz104tB/
WfK0XGhVpcl6fU6duUIXSAyv2JoOLwISaA/ay6Jt1C2X46Maf5cV/RZ9kicP1wek
YC5X/sCuXtQ8pKPzSyZdr5JXQkNurMnoMfKFiUi+iHRcCXDjBvXKibg2605+fUMp
b0wsxAsEWL71Fz5JGUDMPmbpYyVenUxMXbMS83ppxssrGi/maIJ+D+NXwnh1Fyas
miv0FcLlS7DA5ObBTBEW+S+6g2VRq3pA/UaQ4lW5n4B65rHtDCJvNdXgklvE99dJ
q8EkjGWyTORWF3lC3aWtg/FcM2g/WV7DJzf+k3u2LKYUHSLgGz+KDKzeCkYaz1U9
OJBQEPPklw2MCO6jamzm5Pr889MmITUCoEEE/eizdWCVntAK/zAefSt9SUc2mHAU
1CV+Pk2mcuEkq65FnISWE0XuOS51iH/jiNJ9jcKnl+JF0rzBeg6I6qfeKfFrcVOe
h5HAM5A3Crzb82PDE8ZTFLHkStLpw0lMODwSuVAIaG9OawtzmhWnJq2ucp2FiLLb
EBEakmCFhzrBTONIitx11emtsWpmkSwbnI8WbQu7LhdjOs+iDF8AkMR1ty14bj7x
ZnSnVF8thXHnWKRnIRAb04qjE3SKnm3U8V57L6aFXxBxYI5USgPp6K1NMBF0dBrb
cdOYGKW9AGUFB75ZuE1e6JFd/hJ/0ZBxUW6yS2scSnWK+nGXJu8zBeScKUpx14iM
bhGco8zlP/5gPO9TKhgkUcaoh2LdZUxkXWXkQwAalSAfCm4rZz+1f6KQ9CEEY4F3
1dSSG/YKe21InpubWdTcCeu1ni1FCcR24APj5PvsRbwdlZNenz251f5p3kjnMkTQ
ik3vl02LOCDRa6isBm47nwy+++tdJtQ+eQWITs6EZDnZQ3gRCK+HcTfksav2Yg+P
282EG3jDm0JNW4Ys+4d88fhSH4lCM+3+gAh9JcT+IYnnVcWEPXllZmF6m+/xvJBs
uR/f8q44tLUErjDUoBj+z/HJ0szFstJqyyvGG78x7NATVRbrER8j1hg7MXU/LCbS
FNh9zH1PAP8N8K5p9QvLHSEvN1A/hMJG5jLy2F43jI83KKJyOIaRueK1HH4n4iXk
xcE+Q5iZUhITxsRUthv70I69Rq7kiZp1mTtKsfoKe1OIZwiHK4UsIt7P9tf0nED+
4vLX8EejJjum3mV+mk8voLaEBpUN2CInsCZttYARrt2tbmqtvuSqvBvt0Zqb7IKk
c0cG964Gt2s0cUf6B6A96TtWNLbqr3vsvE0+pfFSrg7tL50VcbXWMG2QEfd+Ehme
HFg5n7E7pj5RTRNSchc7ZVepHvdiU4WSvv8PMAcCKZZDKW2MSCHfwZPZy1b4/BSD
e1r/2lMHRziA377jVt3N2EjS/u37wcFaeMBkPVsQWEKrCdOQMsFFTn+3wp0ViJW3
SFCMsLqJltPCM1ZroVJ9oKdrJnF1k33YGhXGCe+yLCrV0QAhF+juCisNchxu4J33
PLNhlm68ycCcfs9sQfklpdah7JmnOe2P1scG3WhRXfsVkHp43gkmFSle4dmiqcqK
U4Xg3fFX3/XVsdV6BNzCWxaaiMnCzSGMQFIH7Rwg7MhCPOsyp38nCtHl8gKaAE/G
urbg4o9MoHu81FPn6TE1le3ZtBsAkWfoZr6L4P9IocPWyAKAA390iHmqhRKM4wry
ptNs2m42a/MGWvijS+6FvTqEU+4FbI0tQSAaPibgKm1Na7JQYx7ryCvaYKsD4jIz
3k//XCXRMe4YddTaVwPvDvQfyQr8EoQ6HgcQd0VpEAL8qHYC1Vlxkfk4a3KLTjk2
Zerjc9uMASURMxpVBbB7ZvIBtHL6vtz2pypPAADzzDyFrSxCqnUViIAlBv69Am5V
15nONj5Q0Rnp4dm6wPkAzPPAfPR8ybICaYrBbDndH2N0YD6N+APfiOOiKun+EvvT
oER8usRe4P4zEqqEpsKS0C5/PY1F/HxNnH+oLvQbPi5bRu/Pbyz/59h0reS0dT4I
He1UMPKY2u52XkokC+vQYdY+X/TOdvTpmTMXwtShGVxsvBn0NmaTGJ4KI0HcAobU
cU++AouU62iNdTIwl+obpCw9zf7+yxPGDBQYRgVFqKaTkvrbwacFmhhtwsX8U1Ov
gnN3U19zGZaQussKP3zRn3G3MysxtswwJRpYToxFO8YOU0eA+NJNUueV/LGWAnnp
JYjWmaxwygX4LcHK2SEYC7sapKLckG2B7U7oSu45o72gvu8V2Rs5HivlnvtoVXmI
/jN8RAgHVbBLK1QVmZv3ulfmQt37e2ZavQgTpzHo1XP9cgZEwFbVYD8DZkSWfkqQ
+DsPu9yLwOS/fA8ogmP4rB/pkzeVQE+eY8482yATpk6VtuPGmihTfHgUmbkSrnMI
oyFtz7Dc55S1qyWCXPMtUF531U8UFSj+vZ+9pUx5ltjKoPkPaOYKJQGvX7/+tbkC
WHRrYEO4zkLVBbSpTZ6mVNVLQuDIwkRlAmTvsnj8rZMvOZu/frH2SWzaCf+YNwss
VDguy8iJdycSwvfol04j+WJt7LKCUmXrPP00enmxTetoZvWG65+ELOq74E4rX1sF
6EmIe4ICd9jcoEsqT0fXg/1c68dFBOi7zS/ZBVDUT8P7UbeSHM2ekF+HcyVW58Yl
AqgWIi1lc46BUakV0KshadKjM2aLnEVvgDHXYU4ulp0ascsy+N2liBqQ+4RoMxMz
Rzs1J4gKvDc3bQ6hZyeZ9/Hfo6mDOVKFmpIZB/U0E2/Gb4vJpeB3mcsdaa09g0nf
yPD0jz5Xln38P8+d0gtQDjsHxJX5bIyqPRIScXrnn715vdV5Ttt//30Tx0Af+A/I
Mvp59ldoonYSd2t9Sn4XZSXB3X4c28WWOcD6JypeSt1XdRqGeWG/q3QGavoAm++v
FWBpFSOsD+5yjonah3Dht0LbAZrNu+K2ktaLst+TR5b+77iAQwScK31Z+3DVLxYZ
TqnbyMITDg/5OeZOWu09umO4C8B0WjK7xewdh/RzXOGbfUeb5nH+ObeHlTXEGlrz
a4jOs2CFV8gYEEzio+X7fmVEyn0Le4cA5Awz5Xmmi5ReMcSxW/s/vcTqNLUvUich
VCMKzdE89rcyldv/fTX7yb5UPhBvn1K8zIptHcbZQgQtjvGKwWsWsTonICP9mIBf
vW/G+lQ8Oe3IYpjomL+mz2U/a2fUzXMzM6TzNAGh1mSImHXpjhDSqtKinSXqcXdf
AWENbSQzkgmUSnwYGx9uqEULqz5kmukeq+C1G905x8wIsiGxpdERQzIOLWpJnqQN
wMUKULVybybCMXos1WyfdAsecVWoMbYDz2w7RNRSp5G9PUgKnKRL8HVXKKho3S3U
uMUkzfB8vQw45LcDPoyDq6MSy0M9vObvagkVao0ZwhxFyflBNY2dJLYdh/D/h8RR
7X3HaMKpay3lWhwQNSRrDM/3JyYh7J8yqj0bEX1y0l+rr36AqrP64acdUrQ1gw4E
nFDtya/3CQxQG+RvjC7kaeRl+YPo45fNAqbSUc0Hnykwe2yxJOWrbdNkEeHouhHb
lJqYIZto7YuUW0F1BeuBJIxmBB9j3U2NSE5qXTmh0nxipWMCj3S7Wx1f0MfYq2bx
xrehBiSoJbvmAoi+KFQHXxwy7Bk7u69TYMCEzKw/l+9KqsWFaurpl8idcaU98Vw3
jRoQRUbHQ+O/ivsDUzT9Ta9kFt6g3s82Fdi+I8MHgTZeLhdLgrOxym9scTL5gmOP
KhVtAH7VWK8Jyey8Cnc77XHnic25qg7okTVZrBh+tZ+KtbCFjNyuY1TTHWt480AT
QV26v/mo/gydx7i7ElQTMEcj+Znk+f9vO2bfIacT7GFvBTDJu1e7fTbuvCi9cpUo
soOldpQeh1qM40YWR4P4zDvDcTL+SpkJT/H+h2R2KaabBJ5BfAG/IDc17n+k+4oK
Vj7GpJQhuUefP8nn9Kv3mejcFOBZfBIWoLTifooiBCDwGUO0a1k8HF2oDBj7pw5K
NAElxXpYnwJEedKXIXc/VplYK+CJ7fPl3Np7hBPzI9+aAAYHwJchjBBucjF+d4o8
pf85W/Lgk/XfcV1xLeLlUxUB93UDnd3C8iQop3aKjG7OYhVI0B8YSJaz1sLRKM2x
+f2tZHby81ANGvyumyiWVJrdIhFGWPcTDvxeK10Jb/lBqcoyYeRtFRPToTsx6Ebr
DIjNH5EiiAyYr00BNi0zjNMYuIC3xegHvEsEgeiY859sTb06aMfg9b2IURL3MInO
nitA86zDSTHdZCCivq8LKoxsOL53wQMP+LxHVskktIFMn97yJU240TqxdZiTaDhK
5+n10cxtyjUDX2Tdr6wf0+mx6GM5gM0qq6bA2WQw9S9N4H9UAR6qAYGZ0AOv8t5Y
rFrSrpR0mttSFZDU7crz6su9PKTvmgo3v/oXvvusomB2KlisaoRRf2IOGeNS/pPy
iGGgVcC4M1xOjMfZijjaybp4YyEINtnFW8n1Y8RM40RbSy2wc0dvoFCIgAeekCWQ
48v83m3eKKciK3s1j4Z1DNzq/UFVa/Gd1LYZLSTbRAtdSbpldlWY4uru8lORZZ5M
LUdEWYF97uIaus7WE8K+tHkwVPsTJqrhweBtglmERAL8q1UWEG0jzNxg9AgBo1K2
pgLbNSkK1NqfOlJI8IlHXb64vK7NrMtx0vBV8IQKNf2AeAiGMQTPmNdZueQPeVxB
2h5vJPRbqxCYtWVnseng5lvUMJxP5GmuPc2EkIITNi7EI+s8lUM+xdjwi+LpnRMz
du8xhPEar+mCP0gQH5hmFW+DkHcrKLOuSmCHCPYYEsW+EoSNgTetu1nagJAH4hv6
dGVzrlJWEmFJVk8hU/szGTt35tzW4jQRMKskN5zW5WD8yMIjZSs4mhf37IFax+Xd
4nf+dBWW+V8jJ+pfIU31mbQNBIcEXNZkA2FWiv0DgQ6/5u79ZWy9HfrLsdWgxZQz
dohIKXuKElWpNevNb2AwFENw2xdZ7Lg8KoXcjluxCLbMAaAO1aS6OibzbdPudici
XE/dJF6tTUDPHVnUSA8SFVKnElQFrnKCM3gOUnStsChwq8UjVVBFGaff1PowdNCR
V3jrZAV9Qq6FkZ4vh20aD0n2NmbRLG/22chpdkg9jF6PwTgZbWazuPzBPPz1pgzY
XYOJ3UNRNkV77SP01g4GW7qug/5p/SNVaIc2+bVIVIUgRavTy4DH9EKDQAZnjMv9
iGMGwc6yUEfRFNSmjR62AwU6cd4H6uu4msu+OhJwMSUOymVaGzsqERkBpmLKPIRL
Nqb6NUJGRWSkf2u5bsCjIcRv7C24onc1WxSgG0G4/q1aoOJj+Z9N4YwrgcOx6JiP
nou6DPAhBaRV46DSxofLI4hrclZAs+a8CtjKmSgomWEhB6s/zh6W1KL4MvmjpI7V
+YIzTNbkNuVxwhEGimqDF9FPrpcfdxbA1qLH/iIlHpOPm1ahu9buI1aU2/fIotbr
e/hUbS3ZybY5UbCzc6KysCbhNFPa+uy6OxAzwS4eiRPC4BBRxstTAp6Q4Eb0fVYG
MOBfcC4P7VEtNep2jTPWjGGY9rhdoq/r/zPRhMe6NDfArbWUsy3CkfV+wrX3e3f5
/xRSKUG1C4yxOLLeOBZzGbIJxrnuS1bjYvavtjwYP2c4e7VU7Hsoan+dHn/P00xG
JVRpmYMERvN54ju7c1/r4i1MI7xb8bxCPWBzrud2K1552LTZsOHH6sPdg0sXtezA
DFlTouFsOIMolKVXrqJJvM7zL4YXGM7ffTeCrQ67decasl1UlgUZRvYGbPMUTDnz
4QYQhcj/rEPNRD7Thu++HnM8sJlH9lLscQ8CY7yFKya2kNm/LhAWkOBGA8vJUkFo
6q1PKrBBTLRWRmPysN7BnsYPABIAEFzjML5Jga+WL5IFttASFQCV6er5E9/75xxY
nZmhXyk5b0SjIJK+hKg/BAcEY3EL7dhB6jyzHAr/0/gYTedAxIFUwH/mCgHdPoxL
8mjYbr3pd5PRfBU/nZzYM3GP0ykhB9dF4usDkzohWbvHsm+SnUfIbDPw7FRFsr4M
9E2Vba6L25AN2xDYJH9+PB53etv9t1SLQ2Rbj9XDcf2XNhH751wMuWeB93b6oCO4
rpfUSTmfdcxMQymJ/TKkiXJ8BBymMZVQqCHLFarUJJPX3ZvubwjgWHUWWqWERcjM
UnqpRq10Q9vPxtwpZ7jY6tzuwMT5KGmAmoqWJr67aaPwLkXV51tucmQN6LOh2drw
gSf9WG1kiJHGgegZB0UpAFAg22bgSRG4b1ayWQQzlXFVlhZTGI6L0GP79Wl7JN9h
lvLftRK3MJ9VSeAPEXKkS9xJ/LGnOaNOr7uyBkWabAflxb9+lkvyXlCyHWuRadab
AWUcn/71GRpz7jE8DuWWocaJILi6seJyZSF7xa6JFFRG4AWeNALZM7y8eXbSejF/
GQ+HxaS+dbFZooBMS66SLYxSgijPDDVHGRs0QmdlCNLHAhUdztgHwd81NpnnJsMF
ZMmCyt04fFAaUSIulVeOzfOGLANaiF3BtfaLAa0A7CZz8kJrBEp2P4e0Kgk36q+0
Qdh45Nxlfl8gwvuvotlLyjY8wHPBPBeZYekuYQnbChBEY42oGoPv+fascBmKymrB
XAd2BMIhcvf6XT6vZBdN3aRao1W8XXIeoOvbPnaFWmY4JHRQ1QV28RofBSSDS6MG
IVU84yHdpQgXkpC7YbRoTuzKyo3eacH+YHSHGruEdL9OP38Z4lHTxCr/oB07UJvM
ZQUaLcwi65kUi/osLDyVqG9uImhH8odFHmQ4HeA6c/dB9c/uIySz6XJVED8oi458
Sx2vY8ZlaFsen9hPuh9ISFh2IZXrEGqOpzgX1iIDZZh9l50IKw+ANEFpAk83pCln
tJatiFqfYPsQbWJIJCtAHrUbPKPU2o4HulCQu9WIzhUjFpubn+VKhIj4KYxgmTek
yOSCFIsCS2sDHW1IWRxEepmgdi8/iEEDwqIX72GTOmTk+ODN7GPZ0sywGvGXBUZf
ICAU6I80JmaS5AlP40JJ5cOMnR30jqpw/vQipA9IMZAVRBX5gWquJR3W8u51P7pX
EJkY3iO5xfG/MUy1VWcA+qHEmyCOFp88MzTa8VS2TLdIaZ3AB1zvHqmxvc3LrMli
8wtYY+ZRkwKj4TSKXoEfka4ozuTbZ4xeHngfSFSyTR04W/N1bzZMu9O0lm+mDYd3
EwpJq0V+aaEPQ4OkX/nNt7stroWuqG6bAr9PBOzklES7veCXXhwBw+w//sIxDv13
c62ghI0o/RY1RwMSsrF08YP7X1HvNEAJ0gWMYOjbSK8WNn2HLUEujqPtPxGHXEFv
+3HiAQ13ltm0n2oS2RmNTKnrcnd7Ljp4EQff0ZTxBpFsogBYB/7U0GHsVwDB6x6z
R4LPO5xIGRbHMPEs2EGoz0+oGRIZJx7lyeaX1V6HNoQTw2RLMUgA9KsGPyQZILYV
lF2292VvxGry4JHt2o+G5IB3xKryH8p3FU8w/JR8/FGMi0Twi1xPU6Uf0CtyKMmi
lID/VSv97diVTn3Iptc1fcloGEuBRSSSpmC65ateO21rpp8GGrwftCt6XJDLQeN5
3yqwWCpMYIEJKzMpBrYhzIRzEronyVEVchFWqy4dBaylVZxQmYdjIcol19KBm4sD
IUcAhBdl+3pd8B+YWpmRDZgaaBEhcoBtM1XJMnjkg5vF+IXvkZzD8f/Vkj0RNZ7U
s1ahvVosBBS7NZ97QT5UlWW2e48QIdLD3Kwni7k8qGHZVOGqw8f+PKDz7Kl1awVL
iydU0LfpN3JsO2bktP9AaXwwweA5gEC99w55/mB1/9IpvtsWgZoxw2BCZ7MYdAtZ
kGUHgbxp2Akkb0wGyJyZxyd/CwcqxaQ8wrQ/ynSkEhVfSXhGSogrSh8gMem3WTWz
6bQtML1k80l1zPoU6+nl9JwLU8t2BJL9hTh2MPwTL6APZGNQLZ2LveCbSdPPUOmn
LYYVczl2Gk7A2ZOP5UHlwQOr4v86xLU66LWNQLHtYnGvkC/ed609qSV3M+kQTZmy
uzdt9wbero/smElDIwSj+KWH/FDo5GBvAalArSNHxazlygNK9es2ZkRhXyLqqORS
qWn5coMvgOFm8ZF41EtsEaZs5uGGJOAVwL8tSx4wstuwwIZDFP0orlcRDEitF4YG
8DZIhgyF36EjQq+Rc1givNGdYoeuHbLFX63Jgg3hBE8L6DynguN467hmdhoHYJdP
3qe6t02gxN1wJHgruu5gMnNj3IXzJeb/t91javlJ2nzLOxnCeccArE14n+5dBeRP
X9BMkelmtjiw+ezlBxbH8zPxd+uraoEw1onrXFrvEgi6Sxe1Aq5HMS3+eMoQY7j8
WGSBmxI2ieVQSjgbrtecDvub+0Y2ttNPp1kHKxv/ayUcf41uTbkXK4UO6T5ieRc/
ecxrD/Rf+jrdVOKupWLDXmJ/ft7GErRyMreLYDG4GQMv7p4TY70RGvmIC1MM0Fak
CQvk9uiMszFUVKmFGY+33ycdIBy9muHZNg5QHWkcOA7zUxi5uAskbNF0f+eIoV3N
cHVQNcNP2ZYQ6j5z/0Dh/TS218age4Rw0Jcno5wvnoBEY1Gb+WiT8PMjtiWbIWKc
Wd0EgoaNde5q8ro8J7oUMnS+JLUWcBa5FF/06egAWRgvORE9aXsMOktWdjlxROf7
JohoURqJN3LW20i52CGE9OXab7lU4CzVILP+xW9zt4LOytN5lnPKwJLsyLWTiLbk
eW8kmWCFPxGysUkdfrEXP3zU1IDLDzB92u3vPaxOJjxS1DB/10sulL29df2qutpJ
8e3Axaavq4/OVhN5H1XipMt3XnrZ7ziG8MW657+E0rpFEUNQbd0Dhx5c9LjOjzf7
kCrmrVeLasATDdnxaSn3QeTRSJnwL94agna9zfEhzcHjLsMH6SbpcfvvXRT8lHeH
xX85p4g8q2FT8ojqTqX61D1keFiWGgWAqLSYkqukv1R+BypylSnRE99EUIJw5quP
lQRJlPdc2fzPCCSQIPinQt8KFq3gbvvmfrKh0U5fzMAOQST64bw9clacsKKU1tKt
av0v+aKhucDhX8RAwhGCLvgGeozEvg2AUlnHUq/nfAeIG7KPU+vw88bzkIWGyNle
TyFvpXhE80TBC83tzFnAwnKMTUHiOyK+VP4rta25FZGzpum3nQ44XuF51Ol5dPpb
1invHDqH5CeF+WUNoFoOPYk8aU9+/F7IFHHebDbV+x2KDQynrh7haQ+HHmaBfKbd
mBs0BHrLHZ0FEu8sDEp6L0EezsGXBy3NBZmQF+3Tt7bhLkBRyOlZgT7WgDa/+x2J
B2GYX1TJo3HcdeAJ8iq5DKEL0z4aMt0YD3WZ9LV6OtJuBNoX02YVuj9op1vBKNdN
PLbD23E+cQe1+eE4ytN2uWozrIwmlS+BM/pIkpzcYCLRFwOoIypOLc61ISIGhClT
ckl2THzZrXdq2dRejGkU9sB+3qrN7F45Kg5Zenysg3Rn3VDjM/L7UHDPsz2C56u4
fdbR4mbVQ9M9CVUfw7bUx7vcR3GFPJ+TatNk1qe2gbqRgQSqwRYiWeS55klXYlGB
WWQAjID7jQ5GQgQ/QzQuQ02FA66VE+Wa5ZGZcKFqYVIAoM0ojTLzRNsRsp4UHB1X
6d2j7ErsFF71t3bDfs8ibZCnaSte9BO7iK8MGgCEP+nGNWlOvHc7+nHqIXEK+FXz
vq+S8ZNZNnLxvtr+z113TPZKkW1rV6cEtCIh4SBTykNUapdzvEYK4+pSxMYc9f4A
eImlZ6X6I8ZMFgNzLT8bsWdkulXIvfhLDQ3R8xQQbnsBS4fPyg4mKAweSLDDJN7R
cZWXebgX+0Bw+y7+p2dcy6mi9wyyE5hSfZS8cB9YnnQkpepBrxtpuUnUX+xV1o0c
9iuzk8RULwRDAPbYdbtpjSYFdLLW4R/15Cr2rGFPed4juhH8/Pw0Ua78fbDBYevN
CkNq2RQ2hY9JT0Vi0uAYmJnVpIk34jEmqKmHJKwV86KIDYLoiOTXU0HfZFEinCcd
RmqLm+IfyjvxPwEGyEi5zOMulcn9RNFKuaXHxzcRlyGA7KJiTMVSlqL+ce9VXNbx
0lfTWSyxQWTEyIv95I2r4TBANst05WWr1CUUg3NTIzMEGsyM0MBuhNZiYWG9Mbze
lmZQlnqIot4SFd7dJrrHH70z67Y94AI3SL63Wjbkyd6aLOV3Qlz42vXn8YXy5ufv
AoBFe5AUucxWgzH+aKRWBMdb5IzguWjZ0MkmzrWAbq9Xk+nEj6ZopiRGCD2d69m4
IVOESodlqbM8pKJJkpCKjKSE6Fy+1kr5XUiAEXiQPoK0nvS34F/tBNkguv5mZX8q
pnNnitFCZDTYIbkw43LyOMwbl37hGlo3YBms/NBYEtaNmsNQbonM4ZlWo9m83qzn
Myyr+4tq791i1c2ew1sYWF+50mEH9b1a5rGPSkAk9Z+pdyuFEfnuv6klUh7S513g
noXpsBA5jPIrOn5IvVmY9gi63UCwKJCI2GkxsqC8AZFe8tnh+zW+6P1HsIquxQh+
F24LEFMD3ruL7vCivifpCKaXYbZ3krLu1lgP2Dm5wN4D3tYgpnR7JhGT6UYAOxZK
rvRexiEnr9r+cbSNnrU1xx7Y6q1UwsWSrLr1DMco37MDe4Yge3BVQvZ9VSkodlXg
X2PYRA4lfpfayebvWxPjGX7DE6MakOCLybWA3r4aJaRMzjGt3wSlmJ8iSy7H79CP
XikyRqeR9lPfPn58hT5g7mJKujPIHicYXzZPoqT91rDkoizbkWAH2iSp4Q4MmHyv
Lpotc43DH4yB8eOb36OQcRY2Bpl4C8QZgl9Y/ii0tfOr2af3vo17/YGh5v//Fbp8
sjUnJSsE+MCxrO+gDm0hDYYKb42YGyrUonSiWrdaqRnrqw2kPgY+ZUSIspghsam0
+r4RCuKFP4l0w87sLOqGdx9BKf6/ARxwz64IH9OKvbUH9Cd63jIF3lYnxCs4Tf2E
YiPqFzVK6JwAmW15qjXRe4ifRizhqBVvcWVgJ/06+kzw2TSbZSGofwGpI2xgOj9U
cErYn6FsE2KjxGCAEfPK6YYCHg7eo9sJZ/psNcPMC1lMrG3LHcU3EkeV21n060Hj
p1YE7k/pZXkPsVMK4C9uO8Cgopwtv1njLReSh8FDeYlKjm2WNhI30mlLnOuw3QEQ
Vlaw4SSb8ZQec7njZZMTut7C7+RRJ1PP3CoovIIQN/ykSYYDZmwWa23nSTtr6Z5R
RBEOffMcpFUqogd39GIxiHW+QZqrnxWcsNMnrdxqcNGLh9bvPQ3taWYzBIlW1RHV
26lgxv+PEtEv9n7By5KHF7JY0ax+KjKcPSwE6rjdSpy1Csza2uadjl/mpqTV/VL3
PEhKbFPZHD1v3UNs/Rka0toXHnbNEWJkTwSlyQg37DFv7mzE+LvDm7rBk/uloNo5
gjGC6fyLublzsj3WQOXKpOk5cccHSp0dQxhVXT8rCOfXnxJVcAtPk4JFB/3dQ9vq
dh8v73xQT1a4LEd2kb7BNritJkgvCvuhWlupQg+YE4dyGJPj/ntTj4C3XOlnr5eJ
N+SwhIRhKw7+r/JBFKE1kHII3RFUDf1bl0xemMjGb4kKZ0H4MWsprITvEITBMhxV
RrAvEJ/qqFMW3WKWS2VO9fOsvVWQJFYsuVEFYs0dmv7zE4Ms7XjVhpGHhj4g1YQz
NBnHsXZMVHIejzfI/gNZlnl9n5f5Jkv6IMQvSLfytVIhemW3SDfKWI9BJzoEWK1l
UfmoPRdS76H9+AryzEglEFuW7Ei4fC1c4rvK3O6pB+NBgieuVOKXw48TwheH85xp
EwNEsgTCxBDG1eA4qjroUwK0wlW/X9Sz32lCmRKwVS2VmxDSynrX/sb4H62vSAIG
8/JuJGGbOqUat5/La3g6ZRM1IlliqL046HgG15peulZRWoerLAMhfxHsACQztfJg
O+YRkExMQx2JQwLpnky5cD3jAiYTcHAD2wSJBP0JRakhXSpj7rvnGjdleu9beSsk
lg5+EsqE1Sq65pR8BtrbLU/JwQ38yCxb2LGjGTtc5iIZ5K02AXlaVuIGeVBUm08c
t/KT4oln864OwOrSvO7jsiRJKimRnTqFCl1wadmZX8GAs2bgfWOw8g1E/14cXAt3
EMzrwDXgebO09mZIkVVDH1J48pm3krNLHQHx2VhihU5ARVX8tpqg4rKtiQ0jNLfl
sSZDWXYoeSLEOBfy4VVRpWKyBTWz7QTQWcbF6AA+UezBahB/p/5DYQ8TmfBhP6k9
545PXjdtUcm6IhuYfMSKoLe/TfdrnmjOvjwL8cLoHUf6AmOqFp8I4BfJ+KV3HVH1
H5+Y/cPZX1IoZ3I8coyWoUkIfYBJLzcihQZCq7+vWAB37V7n1nYZ+CUYGu58qwgc
C02dYrUIA9IX7F8PnKmVNYqY3flRmpgVs4v3+MIERG7OMUgIl4DJHK0nL4e/pYbS
f5kyglIbroGtpxGGyev1QPCN3QOb1QKKo5S+7IQRbWcniYSMQCYy5PlDfk2bTsKO
G//iPgiphrHqhz1areOWUwDY0/ahKQ87oYipKfXlSk0PekomCuC2GrLDZumO3PXJ
BCdQuSBpMwJEpy0iLK88Mpeq+y4nJAYKv6UT6EH4pJ0/7CMAGo53ksF8VZuSNDwf
wYQXgW9EREMFWi34YIdX+D7CDkDjP1Zajjg4HZeVOc0AYzPaxLQOQlh/NdjLBL5C
Gtp1KZa5Z1vWGbxRxsOEyt0BPLzg5oWix28G4P5wHTJ1CUGSrOtXgbb7p1G2CuRD
ttfz3zviI0e8HotUuYI/nQAOM4lPnKL0MsxIrnDxIg8IX8q84EEty9mHQ9TKBBLj
od9+MTt+yYTcQnBLvR+nr5kZBKao7unPehgqA0jEzqOGiREjqsufIoWAdOgaluKp
N+RI4eA8ilVaYMJPPcdDJ2BiVp7oQbrKqSKlptxZ/H/unfJjC7wiHJX+Nidr/P7B
kzI5JLU5bR/SUyJdNBQhVBbTjqcHHs1mqR5mMhrfLQ6EhXucdo1gntnhiQ929vsn
96EiiDncgpQOxHM7GGEmdRww019ydlq95EmCv/Rau9Bb/X7JnfALq9m4wATReyLF
iutjNxYAFBmQFHjcGPz7y5Pk/EnlmajuWyqcgJNOTtAncwGgFpMyfJROB7H50y6l
Kp3Tnlaxa8+BVu5nk+EdOGTS80zCq+GhW7r/wx52wIqkIjiL41G39MwYLKY/NEAD
W+vzi9Kgk5ZqIfgmr44p6Nt+5XhoHPaHkmX81oYKnIlsPHH9A14vfhCXdmsGRYiB
aTta7Cqoinm5qfZCAUXDU7A94roeYw/lTkjbHrlh/ZdKdggwS1ky5HZd5BBzQPRa
BWVXmd1xQxTvLfilhpVHO0WSXKsLtIXmOtEevPt9oYGYHXiZMXm7S13ViwdZdoye
Ji2JKVHA5Drr3wKq/rjpmjkOxb6nAO5xL9hlZTvlwr3ysvypT43edaYFHRXrMvtL
bqEDwDL0jvkHGpBGXIwxufQ9dYAT3q3t/C9DAWIgyrDim2n+Kj27pTdBF4darP8K
htQSOVW+LGmz7UNMRUjCidlpPV7e/wpiV7jQZQhM4ZqTd9h3I5hnTc0FO2I7SpyX
IJbBaaZK+zZXC2Qv+pdi3Ha8UgnNwLSoB4tF012saiP/Sa7PfKbYfdIjZM2nE0qm
WcbiOH2u2/focdMnqTRLIEwQZht5m7W76fqlnaGojfY8N9X/lB5VmUjmFzJic/NE
jTA2kF+Wkm5eU7Q3tadYBCciD3sXsVe1EVZBHsVB5aKCYZqm5AmOTBwf9MySXlfk
/deEEJmupI2/GmTyjn+zwhgrgGC2NIWxTCYjXVfzt8cX+9C3F4BD8kbbF+b7+Chp
UURR/mZ9HiZcpYtcmwMhp3FTLJ202UipGOA/VPeCVZBw3cOyBt2P9pua6pJ63Tdy
V9zRZGlEjSB8PZTj0H6N4ppFD7jWiGOa7O5TTK3yA/0KEHI74Gg25xSJ8/e+jOFy
/QXTv2Va/Lbq6g7cOH4ILNec0MhQQZs3C2YreMqj2IDyzgd7q6W65tL+VrFa6Utl
4Vu0QcLI7xD9Nqdw/5FR95tHnkUKyjc2LCNSr4MuHpPz6wyXsUATw97gl1KWQRr8
ltuPiPGO8HbjEKS13BbScxWYWBUjS3W9kotEokaJ4XjHX/q3Z2krKVzx4g+s0N21
CjExeAoxviQ2KIHupMgnYW9T5m/9RW8AW96T71vN+AoJ7RWH//3zq5IkRnSBGLC1
EtyRKL+7Z9T9RXwb3uKIhFA3T9s9+jAd3QPs+RgXyoWUnUTAWtB2R40Yzx3+QwCm
+nMOSQi2OxenJKEpewYrY+usKLTyFYEcFYgsSV5hyVJ80IEpDhc3LDGnsK6OwA6C
KT6utWDxgtH4TNok4sLiUJbAql96Zj/V6FCnDzASr9z0PSeih8hqpMEPFsAX0CAv
NoiLhjODeNNSg2SXElA/Fe5BKs6rnZt7/zeK7UYJ+aIHEVYdwQNdNJB2enl+a+ES
mg8d3fZ7NeYCn9NS9DuPqTYqu1LpZloa0jkePrvouESoRbCYw5eOmMtbnWrdEtyw
XsZ8fRu6AMqcI/apmRefgQlljsPekLKHt0B+v+y1KpC01R69KbMuYTDl3OgBASJi
VjXayK6zBPyPuqrhy0OTuB7QOhEPc6bCi4R1eJEDUyozm5tzi9ditBUt5KbBJYx0
GDQxdMYUTu+J10zIF0VOwt2rEKAEIW9kSJRzt80vXMFREN5GGOYTY//4gcOI02lA
t+so6vf+euSRYWPLcl3Q6Er9ezwT1TaOueivNbwV/L+2+RzbTDDYaVtcLlKwr9hU
/ewtoM4OmIiuKhjzEI/PQKlrC9dDPrnTx/lvbNzTTm4nmiyEU6047A5edUw7Enw1
wQQp8VbHA68bHzCu32YilA+KCjQHy7kqcDzSUAeAuoPTZcV/seehpEga9rQhkLUx
go9WJudBEOzlPSEnLPzYUGLGv5OgE1YQztx66CdVanCutL1ujjEbeh4DAAdRcXzR
SmSOkQCRUlYIh3Zd3c+I9UiyQRzsHZ72qw4+eV/phtQQ8475V7OSIm17YmWKveMW
a60oTQMWHwCxab6OfEKFpEkoJei9TYBZPhLMjF5igvzivmONJoF+7Cn1nOGeV+CJ
FMW9iOqTFO4NKQcFgDytIdc+d2PsIpmLVXi16yonGMn+QGb8TLui+ZK/fCj3W6Tg
qqATYA+1s7LTp6y7xypoDfTSe6ifnuwkW4s5qHc9giRGQFGFY6n8+KhusICyiXao
L2wTPYt5067rz6U+2nrvXHKjRLj36Ebu9vW2Fli13VbFk3Jm1gYgY5d2C/7G4X8l
iFRhNvZGk+lxESv905aGsB3u/yNETLnyIaIgIAbPhTM+Mbl5lU1qIktPvFCcK3t2
54xaCE5Km26oAslDKACxpCIV3Vfg5p0m4zjdPEu9jiOAlsw5yGmSfiPtUE6JkvQD
fpGyBnLg/vy8FuHL39dw1swL9Q9CtIHe/TScN3uNp2basDhmgPusepdLilrmXDqw
VX3QPzI4Yb5o82mm0me2O6HO2YwSjEK77uVe3TT7DiG6v+C4MFgV+eD/856TgiiS
qDks7HykF6khegVfEm/V7HunVO2ZmRdiMpi5nUa64lSmNvN8dvlbPKn+ExMUnnrN
LTCGRVb5vpnCWpVieKbxXuJdNmD+hKMFMpKxrVhEKAtmLkFDpnQTVONri/3fm2U6
+wWjavsmf2cAlDhHs2odAiJMgWFc9kA4h8wgP0jJuAPhscft4ajTGHc7D5nEVJX8
y/ddEXtpUOCDD0oLOHvTyxbFFPbrrMOoC3PwZ5gXOWAV8X08ZZsqr64mzE3gVYJM
nXrgMA7gpw+ktX3DDKTnYHIFWHWzhSnbgoQcVFvrzMJjx8sEnwfGcnpYC6bXwBA0
zR74sY7CjaoRBgdGu2dkUYSs3f7vxC6y5fP1yUgxpswAD3+/mcPxIEA0X1TIRasL
WtNBC76WQW+pHyTVuPpwc3DfxduuaV0/hc2mMkmp73P92njM7wRcndyZwgmeONJu
fLfsITqkJUFtLIRd/oHvC+6ApuWeBHmNiM6/7pgZSH6uyW/9gq9PHxRmuzTb5BzH
Q2/jC5P9U+kkHrvE9wTAYwFAM1P2rxl+cbLov9POh3Ut0P+BNPvLEWxGYNZM8NKP
AvROM4ITlNnig4DVLiHB3DUYyszj2wiRJUneUDn7aKWEyL/hEgyqaDp65nq23QOU
U8VT2Mp30JIIvNGdc+iv89UzhKXsdFiC42KaT+qo0PMxpvFS3ocC9Wio24TBpa+R
FftsT7J+uRirHq6A+XqQ8+e0TJOh8Q6yE3TjI+rOmRrcRVebAWDeyMoi+JaM01cI
tj0ubo2xghmtD6OdtiObhWPrtP5WhC0R+YfxPE5cPGtGNIg8XbNWR7VypwhicjYC
wM7fIuzyMqlXFTGIPfT1IMokGa6vBYdQddP8HZovUPntKcTUcoNs2XaCXPNfpU4i
DVZ+FNeHex8SGl1hQDEsjkLqhL+KXnH/aioZuFLLMXahao3Jl0UvxzIp5lRRp9vv
mhnBO3LJg0/tw2yp1WuE+eS9IgPp4YVkU1p2cvl1um8c58D9Uy9yODP1NHwZDLeJ
XyFgzHb9QFT4IJ6ceC45hmVQe/iTgFJTpZsnSGxDb9iMFd4ZA97PQONSdi02hPSW
CCv6TY+/a7vAwdpYUWalQNogteP0loTWBx0QlWmJ1Byl+Pn8WFqY1iZ9WzW+YUPB
gtYfhtnWVzoPlpWpesZo+lvFi2O7jKiYQ3gdNCSEnOPLSRnkTA0hPG6rH4eX0Gmj
L2EI3Pvz89FWbd156z2eFUcHsM1MOQTA2HS0tYMPgdJ4SnUCRsMHKnfDE8hXwMl3
1BLOV/WXbMNf7jU1B1oiaqTYpV7MiQSE2Ch2BK3j2sYhLLxXhOucvDoBHfyJ8oTQ
jbbGV+tntPWsP45HJ7jLQ5EQPYLy6xxbm8Kqkur/7rqu3A/gGol58RL1j38Ru4GF
Ppg1rGoJXfda7mVip/t3eQzWs5C9sK4tvSgSs8eUBZiBNqH6vf68DYUmfL6cCj0+
gNQV7YH4cJRbIv36DpzfZK3yP68cwPOHrJtg1fV4hBdfIMkk8VPSI/vISK93P+uh
r7C0fIh/MYcWeE8U8t7uiMpuYQiWEaF5pUOPfu+YaerHxv+Ab4KrBOmn9l7a+zvp
vGGl5we2eAmjkWq6SeoJZFBMQa/a9YD8Ke3R20+tiqD/gcUgK+XwTx6We/85Gi2G
/duKgZyurswz9QebbJ4dcG1StV2tJ/eKW1mbULVc/SHGXBx2PgH47xcS309KxNUR
Glf/ybseNxIRgk7vBmfyGODHbweBXGQU/lH9MB5gIAGyuJjjOuhh7DCegx+HaDLP
OgK7vfVuFpDPm0DYSjNzGYjrDtwDl007IzixcOLkoO9ech4UZ7EK/e1IwYdP4ftz
Hn8h/eVpmaUwlYeqwQ4jpCw9jESE1nBzcJ60eCNxCfzSHp7FohZR0YKuRyqiVA4T
X0gM6PI0qd3stXrthTKChaiHBQHhrDekltl5JpPcnhN4iA1uVqfwrcDqZ+l6JCIt
GGkuV0IVoz6IcS1UPlX1i+BW+e7k227TVJH1L6itBDj1Dr+XgcQeo6Uegu5vI8eG
mLFAaJIyBCt2si6tYMl+rkEAqOWu4pQs/Fm39jcsuZtxzVe/xoEn7MIhxkti3dXn
Cwu9WA3s8eUgq6TMXjfX4w/7bQf+WZFvbjANp2QvSNRm5vWY2dcM+KfchnAuRgr2
H6vdswey5bzDiJiUE6+gPR3m7DNADAfoOrqd331GDVBK3cDcqk/Wg8Pc9n6dh0Qg
IHhiL2wbDBWZiqj0SM4LBtnUy9Fojub1JaLYqIRNslnltEVewkl1Z8sxaBUL+fLp
nIqpIopQfty3/KbNOrpXVE8BW+HVslgyfCLrv3d40YZzDKkKnaI/8NteqJuc0nI8
XkCjbKsgDRz5MMcmAkJr5dJZ0MSzM7VMke1vVWxQ3r9Uok+pk83kHBngHIoRQWtY
jRTrHtIzTYylVj8hJ9EgLHqIz8oPfYZTaH/XUcQbozyydBrIAn0gjeyvgOqSpY3m
2/OfC3rZ82c5eC1TgmGNMlkFUy1og4nVU5zmalx7NiwSjhWbWN/zmxVVxokcOVQo
X7K85MKXZ7bR/XlDADNwb6kFG2w0DoKm+AF5qPrR/1s+LfkwIuo/D3lLhhfMqhsv
vexiv/rXOlnxiH+1BKhbQCVYb4dmp+IWFiB8Uuf8s9KhpH1Szz+W5Iq49RP/Wi06
smYpI0lj85Qu+Qgr548/dqHjzC1vVdmdv37mxApHoxdzaxvTFRBnk/gEaPnttI7V
RcpyoWZE62s6e5qL0LrvSAml1m9pZ9ejSqiRPDtupf2FZzw9Spmk2vhg8u/JeIHi
sTa5CVkN4ve1xVtbeHaGUmJhSjDTnIsQ8XugeLFtzTW27a9OIeBkh3cjR/18KNS/
QtOnRoERRgkgfLVzTKaksh/2mltNSLN6QRuZ71tM5ix5t80vYIxx58RE2s9PH6Nz
4IibPizUuLL8Ho61Xigxiy/o1TVlQBQm7HlPyvW6tD/dffMZ91N/Rba5qOeYgka4
Pca+bfWu0q/v/oHF9i5U3ufQhE2moEMgfEXbI/y8MamFENMDp9bGt2srFcXeRzEB
6Ue4nZcFVeRjcSY8omD4pDZeyzRQl9hxDReCkXojfGq0oqQerJetp2A2uHSCap+N
HMmbyhqsDiWzmFQ6IZz9OqUiu76SqkVTo7W9Ag0lfKRNa3zKHrNl8RVOL85OA0yy
CgYzwAg4hSLvnEHsIYhAVMlZulFmnsrpGc8q8boZmRBUzb128nAYDLQBNS38Stac
ZGRm/hXybLDUIz+/b+0vHvz7oQRlBqqXU1/S5NZ1GWWVbyRqiZtZPdeCnpdtBBww
TSNLx/L/eZVBczfC8avT4OKpEUzYQ6MCb6/05VXVlfU2N6p1X+dOSzLx+qpCgfMW
SPXzCv3wWSv+PWudVziKXCoMC9RkQHFzk2WTk7WL9dSH7vAvujF8MUcJFiCW6Uyl
J51Q08Uu8PjVAroN/bzZR6Kmrc7tEoXXq1Icqf11qAD0uXFEl9D/ZZA6fq/aw2gp
Vb1TA18xDDDIdtZClbpg0eOAPNe6sssDwWjUotntxHYochOvQSozFCLt3kLIA34C
vwPARiI0ma3dkhw1SWMuta91ImX3IHTNtSDTKdyi+OY6uaZKLp/h+9Pkh8VernHt
WKbRXgRQLfPYvmdAxAmZs3so/CcnWUCaNRa5/f/KiVgcgdf1CQw7tBHIHUMVA314
yLxYM7PRTdB/P2fx+MmA8D74GynClYrdE0HSfp54sekp3ZbVElj4Aq58XEn2iZsB
ZskxuKqo9yM5tEow5Aob5HbTq5oX987XtVZlm1FKPeiZ2fbTLKEg25hU3GpjyYFd
9zWMxKj6Z2xRqO8Wr73HVQon5hs6JAHl2RbgPHaIkK6ZtaHeUd1sa/jhduaasin/
ZJUCaQWYOxoh4cbr4bfTMVxFNKxWXoWHL/iZW2H17GfTshyWKUOcAIcaGMZOmoEH
QXroNZkAeCBOIe8TamofH0o4IY2hhaXGshlS2obNZdPBAkEN6D9Q5hEhsuQT17NO
UriIbR1+1Mav/UbH9wpZhIZWG7xPAKd2yaj660upRUeBQEVsN3folbCRv1WZtQPR
KLA6MNorZm2zWauM5fmXALG2XV8d1f+/xABnIdBgM68PQIDArFE6VVtL4XSp8nBf
/sAyR/R0ErPPmoRMpq5PKLw0OiW1FLkt1I1QEp1UWgGjW9x7LkvqPNZpGFtOKvMC
I6ZxGgFGHTzW3gXF5FwYlPWJy5genm26z+NSCtS9+dEichaaQlXVJ6hbW+MMxHwB
pNY4I4bOWqexX2hiGowQPdrlyX0/LG6fDhr6RouSGNpmOpsnOFAyy9Evyl7vZwAm
86jA2RwyrdggAeMbPKZDV7UOsv0M9DWMyXzD0Qoka/IruvOmKlm22l3UG9CsOT/q
ujkehJYnSEn9hrhu5Pk/XD/g0f3Q8aq2AG9u3lMoOdfcPcioLbuxEtgQvU/kCB0j
oAJtDbrBzlceHbpQGS66pVq108Wa26tQFQk5YefWpYF4CTz7TuI+PJ1tfJtMWhFO
dmughzSOqfqCrSkTVR6UcLJO3/GbDj7SGVpCjvdoUo+KMPZBbrB8WHLHV914IWMT
Hhuw3Dh2jCqAkQlnj2ImwT8YHOuB4THLQfNE+UqbGQoidA7rdV24vJCJs+UhV+1S
b845sMJ1opVTw7utFc8z1BzFTp6m9rTDEyUYnL9abu6XhxrLftb7bZT/QZ1UiKtV
WeOMO+v2NDTRa52U0MIBcx8ObaV/JXeoQLd7Otf9xBLHvjiP4y76WjLLnCacWoK4
Oiqb4bIS9yZDnXma5hRZXZ+c1FGX45imEDT6B/imyae6IpzxdbPml2yU7cFYvKEO
U3FViYZy9gnh7L3sq6mNn679FEwc1BWHo5IGLznSrAjNtJa+8OhZC7b+Okg/Oopf
ixJ533lqQt/MhGFtI6VZD31AAatiNLKW0NQ2xRl/FQbZ06W4Iy+k9e/8+hnfSi6n
OXEWQSQafo2Y8+mb9/N2SH6dZbdb06JfJIU9D7Ok+am1IKue9vuJSDIhH+CjYO4E
4TkoLYDErPEwdkpZ67km+c7XiBpYs5p5CTNdB6Ch7nzG9/CSyPmCjXR1bpFrOi/o
M+GggWHin0mxllncPUUwh9/Jl7ko6hCgAAM7H9+NUN30WVm/ejaJAecPsvkws3Fp
sB81c+sRNoHGbwmbr5xB29nGOYX5S1Swofq+F5UNILohCoTdj/hv63h4lpq8vVJf
+8aUt+e8+63JdSYDSGOu5Q1201saqErGBQ57yJQ2+OeBzMx199iV3VDPgdbchWUK
VGNZRhPxSh2UVAwkv4jMJYRJ12XLNwkZ1Q1h1UREFjGesJT0ppDYQnqVapqpG9L8
FzdsJale87W9h1xGsxIt6t0DeVduPnSKfKR/Qt4/WmGdkUqwl1I2K9Zfs4UaO/tK
BBi06PX77KV8aFszBWVicbZOXDu4rXL0At2na5py64DW0K2phfVnb2HwraRvZnqT
HsmdeRobduzF/O2fT4xs9C7pRKORpzXg+zfLIaHxsKUoxUIH+tZ1GgXyG/9mUTTY
j02gjaTW5v+cwu5v/vVG1VszUCPGeqtEfjQFzGvIrMjgixMQSn1zN3GdgVHLaExj
QdUA8eBXdYjIdiXznIW48zleOCDdkhVPTiEexi5fW8DHp+l67ShUY4CtmPtYTE3i
154VdqFeEX9abaeG4vDqmGAmZTv1T5EfVcNtREy4fBkBRB9HmtXaJRyC/nAWhhj8
PTo3N2bCYb1kJcE0NplWSFwX96ijf/uUdI13fergTpKZUSz4+q5zC8h+UPpZXhvd
MH8mR1dnRw9Iabb9rlLwjvPRKvwyx5JbcU9rlpAxLAs5uzn67tNYq8sdbV1AMC3H
QNzAVkiQ2NAXA8uKp8G+2S481yVXie/S9kwLDlSdl4uru4xItMNFXgaGWVUlRhyZ
wYlpjOrHGSKBI7rM/pRLWIh+lYJ7bTwmSTqhci8opYJraBukja0GZVS6d5NPzJbh
PNlvwhem4Gu2zbYkuT6Pdv9W/OIdZLMYeCKEhgr9ap6ubuw5a6kWHTIYJnivfWFI
j9NBYQU8NgT954E73oDc5YzkVKVCduLsvyMe/qYMTpO0p6eQO/jedEQ1sUGn7Ffv
0/7ECq2IDVv0drs7xV49PLPJmsL+HAzU41Q40qZt0KEIIeV8Ejj5oU+5Jxmx7EE4
ZFL+O0YvMC1RbrqsuqDrMN1cu1JtYui2wrU7tjIrFaf/XZKSqMxJqRyfpZ5dM9Sh
71dj2ev8nZLmpsnUXFNI1DAE7JbBd/K2btIdPtfp9E4uPcfWPiHb46wzGNS25TTM
axWtmD57AgshRVAhIuNXtM0iFIenk86t4Alx+We4DnkX9GbjS/LOG0NUnedAKjwQ
IeQvZfs133U7azfwU/kMVm+ibELizNep9erPPg3Ht3/oblzghomH3z7++7CvzQQd
FKyHo/5uHkgYY/xkjQiaP6us6zpXBqHikdA5eKjBbO22Uca//PX+RVjH8YTEBHXg
DNnRPg1jagKrhxeq3HIkMQ0efCf6KUxHjvamVOxnwHdcB6bhXqS4UQczJ2GkFv8X
sWjg5lpGzfZhd4XygnG66BNw9pDabcQsfP0Usd9WKUfD36QEQ8OAdJDAWj4V/3u0
JNdFkXtYPmiu1XtDDa8j08SQZyOAQWFktCLRYKU78d780QYQJEgt1ai7cbPUBKve
E6hDTmKy0/M73g9fD3riecCT//DN1AU9vKW8CCJf11vCdr4z7bx06JmEfsoEGUcy
G97zW+8NtqsA42Uvwzrhk9VhtqAoZP9jxd9lEdB+Gde1UEhOoxdjsP5bT8mDUgG2
tyWblpiKmvNo6BNBgK1KFz5ItHMAd0ErP8+uXFpWc9/ZQ/LULXwsqznr8Nz1VCFE
6PJ5jTSKqbTwnkN/DvpUZDQLn9S31Qvc/2F7FQIqmQptbcZ21q9rag0VapBWT2uF
LadpZ5mTtS6WgO5xkKOYdYKXt46qZ7fcGvoGpTqIog5DV8KAAz4bYAgp28JZ4KKB
ZYVuZEdlP+VneYKOOfMX3LpBWPmSpciNqBHZ1Ys7bCb7QKdZ71KQEIe86M2W6q3o
SJnpRtOyaIhWqu8j88tY7fJxGpvCOrB66n+fz6qMg/WWCm9SqaZ01qqGfzP8c+PO
+LtWtlKD7Wgk1k5BAtb+wAQwlRF6cWVqb/wsGAx1HylEdoA49yDUYpist2pcrtiN
9sSLdtXNjiAEZJCwZIMdasuHE4F35mDx6VU7Pv1MfONdYfNyftky52xSMhsG4hEd
4sCWzAHw5F4nvuQYSGKhWm6msQNfJQ44DkjJ4906n5tqxUgXWyiYhBl7huux5UVz
HgAFx3WWAbA8SS51DU+aoKVHnlc3YSSY4brdH0sm9siDegERa7YksPPRmahA9j6y
6gPIsFbderZba7X9ooUsEFYbKmgSz56IAeQCVrim4WLfqOflyR2vAcHjI5A79yFi
KTLBdvbzQEByYUae02xTuixvnmYv3OkhG4rejKPNFX76oSuhVTJtcikN62fbeIaI
WkzLd3dH/dVm8XB8P24XxiN9FFz2B4AsCC6HqT3OARyIoSdKDmd/cg3C22ZMQOHv
e6r+X/M465TcVWwF9KXabZV/nic4QvYHkXMYL0z1FePxFrXmPHnqWYt1pvkXAKiW
E0WU+Z9+hRycoqL19gt4jt/gBimuUvrIbxeoNbbxihkWFCXdaIkMdVpgQ78/L6Fq
6niebU5jB+45nfnEqNoBZ4zLVn+PN6e2/EBg6jfBzR7S6zoWOYNXTAkLdx4yDZNe
KnVqC+pseVC+ac8PaKEY29QbXrpGPa2GfmGVmQiV1ylrAHNQVK6YfIx/KwjnU5SG
JFep14RNCjMDfx18GiG8gX07rM/+qilSxgojhIDKpFs6Gy2eyfOp5OlMLGECPXC+
HrsaUcuxHFRvvDzBu2+Ut/q1QOZgUv1dbAto94g5AKDdbAamSy1SetOG6MqNR+Fh
niGVJxr6FNtGgY4FRpudkxmth0/mG8NIycSZktckq1zkoBwWNK8l2PhhB95nphS9
NpTOtl8q2DIQHE8q+idY9MQVrqgeYO6/iz4s3L9DnA5wq/uU/QJsRztqiF6+QzWH
K4azsVv/nvUUNkcU7YiJJ8iPyU7qqFmAznTa/EpgfUVLbEg9rSz9HQbn72TtRr2V
3BTC9TwSZEpZ+dTxx6geuHROM88DLQevfR0Bx9LjzDqUBeX0LIqAY80MOFtVwN3t
GDVz5M15e6RtnSgEUKqCBRZCnACcH3A5oT8yv1OMDg4xM44IuK3qCCv6e8RKkj4R
ahN0/1Zr7w8iI2/J1lVggsJ6N/EF3KU7eNSo/YbBZAN3YmiPPjbBos4DFXMHWap9
7KIXXfVcaYSZbaBf1drv496uXpu4yqtgkxiNOEM/MX1cXH0rBYSpkf1lGKwkl7ZH
uUP/kvwuYuNX4GVDH91yeuOF71t1C8YI8RNuIcsGU/8TTK0UyBCCoW1+nQahAxts
Eh8JFpqULVCkDIvosIMTgqzEu5ZWeZMpC+GQinN7QoiJW6fvz5Imco+gqj/8ElGH
paruB/Vp13fqjSF6T3nJTRFWWK7FgkZMOIcQKf8495Qv6XSYkq+MpiCjZgsrvAFD
uiI8VY08hDLPwsIIszOsEVs4ekHS9cXaniw/gqb4ggdnd3kVt+9eSEdvT9mWfnF3
F02VJgrWcZNc/SqwcWHhq7Lun40Dg4Sq3B952x+s0L4aS/63dBYlI7C2eY9CLWmv
I8e3gzDhQSQmH3vs7xWpj25dMmIPQCWQEUxSoEGVjWby4WqS5G976b7jiaB+SYeD
24K4abDBCK3ZBtkQCF7SjiFKOxl8SNFghrO8L7oDwr2nfu8tVobLVF546kYUGsdY
di8lmrWZ3MWK0mpJX7XAL80bW8yEr+PvEP0CYAzno3ggwZF6/AyzJj/lk/xAgT1v
c+iNaXLo8MQQ3sJFLGQoXw5MzxAyVAw03fWAB1mmXelDOpjzqa01/zU3CCEXWMcv
683+Ia6LdR/k2S5DfMOVGVoMNSdlr4kdWqBjEGilhfwNsaEi5ToeZyWxTZDR++Hl
YzfbVygHwAYC6gjJiv4tTtbFnzYTn+jkw+X2yr3PhFrfLivzs8r1juIZGJgFV/dm
0/nUyPM/BaO50InXz1VX5KAPqG6WcAEZ3VoOvlKa2VpxbOXIsmnsewttw47T/arl
kBp9WKoiL71kJoeIZbaZiHbqrCAV8gGKvd7Zw+Z2yO2ynPtB3VKgkOWGPu7B0MGm
QJa0wi0P/BRGzmKtrc8agGYSmFt+sDxXRJw66vHlqvQLBUQEAmdwTAYS9Zl+LD4N
9zllx1KczCrAPAN6RysDl+yxc0CMw9CLKkH6MBeIiF0qMitf3uAZ+lc4Bmv0gmvc
99BNGBj5tGXqkwE+r1rIaDYwwq+1VOE4vcbXBNEkOij90oJN7BUOO6bBWA16q0et
yMgQeJ04neb3QaCYgtFguVlfnR9riETlr0HpcuAnqEyfLKnY1mvW2WKDoT84lnq0
pMEcxB5u22hcQqoPg7bkJ9fJRA3JtOFvlJSs2GRl3e2Q8xR0a3F+Lw3nPJsrHVza
+WJzGeNi2hkrBqDUny7D2n0AOgt5oO1Zvhp5uxwIErmx8s+g5yQsxeVbIM8775MM
O/DhP56/EVHjd/KteDc47XS0FLI2X1/ow9YWXddVWE8lQg8y55s5m47i6/hImRda
yx2ZWsE7Rw4DeNwL6rbw/S4vGrsXBANSD9UOI8Zp+aTAZhVFPcYiJHDhW3gGZ1Ko
lWz/Yxv6BrJEJ/2lzkQkxgfzooWd13bJGJx5he5co9hbIgVY3WlBeu9N/cSwjtYr
QwC7TwdnotHrOO8oB36SdMRPvU1zrm04HvWkEw3k2VsneaHVSeq7VHAo0klNC2Ye
oAaRj1S4m+Hwr1HLKNh+m4dOiVXwNYXgsnjCB9McuqmEF1FAWGkhnKIDBgExKKYo
C3MZXsbMo4kzBC7n0zornhm1JCDBfNkL9Etppw/+f20rmRxy94SqqYKROBi0j9K8
EtwJ/jskrfVINr7ex9gY9uk0KYePNp3/mT6kylx1nFk3yqk3nqQbthVrSDI1qtRM
Xl/WeBp4XfP6NA0gnqrHryhCImKxppeM/a08nhkHrYGUtzkXcMMcb6dZ9qn+wrql
FBmBocYdjA6+vp95LKMIt9Fx0mjKxD4M/6rQ+dtlYkPJ2tt1cTvtOLS8uc4nlzzs
OipLeV16Y8S4xfFu6fkqzpwqpK2BZatKyEvQzcwHzLM0mUPh/OCOcBm8vlIedPzC
9ceBbIw1dK0ZgfCjyMQkpr+e3QHdEUaTui+cv1FrDU6y6sEpV7f8XUyhr1OD+OzC
7B/5A26PbW8gEld1ob27icji9AylfQ79+peKWGofqnv2WKAPNWMKnRWkasMvPssP
E8hMvuLTPIn0Cah2a5rEO3OiQ9+PNSi5suXW/kBNlTtX9o0l+Z1aJlIQNGLmW1oy
m0K9oxT4Ptk0XbK8vpmqs85ZOGXcfDfq2D6fZtXPxRhVkTHKYyt3bCzMEMvYy0PQ
hlHeIyJGpRFZ4KySZU9ZJgCv0olsRHfHext0RNLHWWwaNwcTB03ugDq9bY/8NFSu
sts3ijWTdDS9ZbJrorm6B+AKCvvMFNlJV5gjgal8mZJ9/aO3eBNO27HgpJ5AHLL2
YG/oUzUlsYjXho3mW/H6QhGJSf2tzlzaAeVsro70SZrj6itLE44g3YZIzX45O10P
YnQjU+JZdhTg/jydTetC9KClUYVx+KkdYJOzKN51FprhAj2ih1Vd0rNioCbn0r4q
oyhLWAj+zXLksYq/34UG1RstWe5tH6O94SCAql8pz+t++vXYFpfiaaUWnmQs0ruB
NNX1MZ1C4Vt51HGU3StShnzPUa8BV1ynira56JHhB1L7rZwJ73bU9kS55Hke+IQ+
sN7BmnLY39JNjXkRrj59lHIfpyePAKfsRew/3W3x9k8PiQuXkHX4+xLmrJZDlsgl
g3AVDUO9u8eoKAGlzFE8YsaCw8XregCNz5NKLqn7sn/02OITtNbRu3W2dtWd9qUP
vXZHBOqurwbpq0d6IloSl0uxrMR5cn4Pv+JtT12RodE9a8V4oHDsWQuuvuezDBQd
0xBv4yocnK6kjDtT9Y09aWKLuhnL6UQXviCu+8xKTkIX2Dy8qBU8tOQM/FR46NCr
YfiD2DWYV836irTzoe0bMHviGfNB5IJjncN2jLKL/j+3bWooN5LIaUGkTqTqzHCf
WA0dnmqb2czdzI81wP3oFhJv2CovFcjywyAMjQmd702+uqY9qh/9n41Ma/ObU/Dy
k8kFjyID73383B5QWYoRJ5DNYw8jbpbo8jXw4brELXf+vnzwLmm07VrX1cQDPhBj
93V0CPbZVoZMNZNBpFofp926BBXWdQAeDaHg17HmMy03K+6i+yNM2o20Lsb0y5fV
oB9J0efRc0xAFNyNHTIbgQ61QYm2/EHOrskYl9S7R3wocqxYaV5Anmj5GexyEqUw
hWKrRoITRVd2G16Zkavwn/zT+2LR6BV+kFLobWR4zajDtScOn+9SGQTdVAevWiVq
2YZ1W+QG6MhjF9zFOzhX7Gaef7M88biF6PAuQXiOKuFkyK7em4thjOh5qv/ONjs3
EpeKRPs7oOk6NZwDmtNaDCtU/iYWktGKDFb1URKiULGCRQFx83Wa6It/za9qccu4
MKeTgBszg4CtFkT6cGZStx/9IknJgsrMMcAs3ebNBsMfxTchzzWkVT1+YCXDmvAY
q5yyEQuapcjv1y9BfRhyNxlCx3oLO4MCAucGx90SsZehewGWAvtNre4MYzr17iL8
jMrKEQglK9CJkVW5e1s75if/+HTcA9mb3ZkiDX4O6TiRE4tnMxjF3wr2zmQbft+i
5nUsDb8bbJ4iSMIZMkxlYQ9CKYj+XVIN7AwQVHaK1aF5UWgXlQlhLCuzMinBAYma
RP+cbIm4erM1XPXquNlVO3dNt0BXdbpVgXHJ9BLvPRTt3Hr7VQ0PY6QyJKRZcLMW
JHEY3SLoDvburbODAWQ7b3dkmWo9aD/nusEui4UYgQIzy4zrNygYfjf4GsdsIrtu
J9xcOhMwyvg4TF2WxvFlkL1TGS3Zm6/f7Huv7Xdrk7zpIjsibGtz92s3GZ/UgnHz
wWNCsGDwhaF6aNwtc+V3aifYGVEXG3/SxX4+s+wz+WoKvy3W6K3SN9CS74DMRQBG
BQohRiElDDTMXl2ZD872DOEOujwFJbLOeS13/C6HgeDAY1CkzvDcV84+k6sgDVF/
zsLJOZTXShYDt9WiB8lBvh7kfnVf6XYqQZcWREr00Jhoq4jMNBmSaydfcxwuh4HD
xPlu0K4ggBr9e+l1/8Wsu6NVVMON6epeJtv0blntBoK76T3Gs9hvLeJvHAMWb+fn
1hT8mX7uzaaTVx7Ho8souM4q3Xtw67s1CzjYe+MphM5TdlDYG5dJN0mWJXsN+HJ7
blEnninUoqaoDY+Bt+iNHjRaPNkoSVwLbVNZDaJbQUNvG5Q6fVU0ZbLLQ/esHGAF
AMFxFBA5/0ljLExFgbSyG54s8VKiTjjklOFcHgr4QlFeEn2iTmB1PfFGDU3kIQ0t
uKcReJvi6biOoBHujTw8RsjEpUZ/KX4dZfPir/dm1KsYBzKbA299MCDxnK4oTvEX
W25ULCh2n/M1DkvrFWAx9g+r12xGaTf1DkYApX9lv75xHRJ1QE8HJBd6UWMV4LY9
/oEOoQ4sptTSVpd+eLHkxtsu89H/mRi091G3tsLWourgeCfBBfb6cRsYzHAQ2bA1
SF0apyE9g7eDy667ka+yq2QIUBZHOdufpfpJP8ydUO8WGhTXsbjvxbfooz66WvCR
IT1cXfOHrTmtJE+KhbyLQyplw/91iPyvdlYWV86MFU9yzV69/q0/0jN0Ze/mkwPX
Dlq+kb+LO8aWmJbJxXweW5qCYnVZp+bOHpw8pT3G/kRUaxgA208r5T8Euyz1NLZK
A1IzaNCSOEZG2jhZw+/lx5uy1i6sWEpLdnVi0rp0f+tc5iyrMM660i1ZSeFkGrh8
15Z8v9EZqd+5fjMfIh44Lvsw0XTZmMJJuIUYzxsjG13hPlrPQrRmJZEymmK7A65U
vSjQKcEaqL43Nc942snLiV0c9n1jI5nCw0gg6UWPAA5ivQq8X8Jv+Z9OieixDp54
H37BzZDSMFFrY0V8hc15hsMVa9M8+kxnbqL7nLCCYBrryASbDgi+qKdIxkVSVPCa
YN84GnY2i94ymjKBQ3+OWAmAWhZDU2iQ9tNlcHmASvwDLg83Gqi4Ws97Y+47iXuX
bkDzh8QdTZD+KJNtggGqNm04J224SUE0qIWYcVEtgI8GVtNMKATw9+tf+b0an1Yj
O2LngWpzvCipTkH10RKc3trhOsdBK4YuDuR2hfU1PdmwdldRDE1//0sjCLr/LNDn
jvC/Tr6YJs5yrDoAZ5gZALhCkc+vhDyLo7kWf7cZfxYFNEBIxz8t37zD5p4w7mo9
IXJzMyAO1TMPGuSwHAcu771mpQa4DySzjBcH/CBVKxET8xEndPrPp1olh919FWZ9
/kK5esE6BDR9ZFJv586BtUA/OI+Hs9BGBuqKE/FUVoyw0Qd6OpZvTbZb55hM5aZY
/XR8MK+d3K87x9oUSA3AVangOGSlGi6lOX3O/i2JECI/rt7gCtjBj37NN5seQDXg
6kmRmAEcjSRO2vXnYqIv/hD0cJS/Dp4kmV0nDFle7luyxiuPN1EK6v9jfLAc4nDc
NQL17EXQ+PtG9AN+2Hjo+Nu3hXDgkVgJkLgeqLTw4Ixh5UzOlAM9ims2D2Z1cNzU
8LR7gzlCD2nid1frVhzw8MSTzhIYLeGFD0e7ni2Y98W/aPAk6YOiRT73dLpr8B4O
hxojaScd1PXsZ/xYRJFQyi6zHcjn+u7tjlMHDRZSsUmoHDPkB5pwvQUcrWbzqGhZ
lTpYZBt08prD4YfH76hy5WwmZ9lNWR1KoyEA11IIz3NRVIj3oqgWDtiJUiIT1Pg+
eGlBGt0kO97LRQHYj9ZXUQ7dawI5kU7zU8hqgJaw/DDIBlzB3ZPnZHyioX28yqOL
SGSsse0QxHV9vtzPlugR2BL3Vz4CTIKPEwgThjZtlgdKtroppPQLzQXvgDaUX3VI
9LPSbsz8wkzeBuHWv2k/tcokBXdTJ0GWx2aqkE1li3dz3plT9JlR6B4+umEM44SI
8CL24xbevPsfoRDUF13RAIxknqEpk6c3tiJhMS3AM2HpHB8EXe+dgpiQRlCYG4+o
jkjqXyc0e/O+Ju4jiRwrnTIdOHKam1X9WawT36e++dDJwF6F/etISUiLy4tzTVeu
0EA3l/8BYzwsgBxcI6nj6aUzeu4P3LfxH6xlmUwgFmilelFtUvJig041aMBm8aNv
6Jbs8ZKdTNvjnljClk7p3zEg1tIqhwCrgLV0nLBkVy7GBHMOrpv2KBeRN8XbGrVK
ihkUvYzwI5Jq3IdQJTWiYMR8wyTSbBnk9WKVx1fMu2MPLpW//J47DI1x6k1sExZV
pYmXgfyziq3gJiPg77HIyST/cOlV0jTpOXBVbUc4nCgwvGGy1APvb0FispLCmIja
O1myMR89LIUyUHJmFphONZHFKwv/bof8ReMQE0Y2k5CZ+hs872xDJo+nqezRgPFL
q6VFExp0N17jgRVNw0+oAlofy4s8Q6IlfJ/AL+bAQljgCLz+9YoeFcV7dB8kLuSY
h/LLB+aBvlYvBYJs34xUiKierIiN4c/USDjVGG5AQT+fBs8l3+QH/UMyU0U5UkIF
j3jBY0rAB2meeXdWR1W/4nUO4c2lLcV+TiQrEAiufunu0b8rIppk4WMkUXvs6RBn
ndnyX8ZuDHbCF5/BDNOknct2gb9seLU/ellehBlLCOrGW5nYhNO60nre/YQHoWA/
n+2vrcdLVLBdBBUhAlkVAzQpieO0LzdWe1x5E0gEa1srFXubFhFzQusgTlKbdDPZ
d5svuUbGhiXWUSZ9FMj5S26GoZoUFEvx86yKOEiBvA/dBYgvyV0VZguEypvrVE8u
mOg3NIlBYe8cQu2uCiaAOIr078ggic3OhYKsportXW5fFCrvaUixY/IcapPwfAXx
UIgb20QGYy1kToqMpjzVf1Oz51+4TPjFfT3PH7qXnjV1b5onstlwRsMTfzwz47Su
zHG1Kv9MS2K2QFT9J27fLcurWhZshFy0erOAwpf/YDYk8PQy7ZdpLfTok5GRbdaP
30Yn5Q/p6Hov9SDAy96744moEN0MykhMPbEShluSqOHycxVVXFBeeHCIIuTzNl83
jj/mJVwfMbZ3d+av+l3qxlkCG/oy3mktjgYmsNoHwrP+XbxsvfMAMLa9Pgo5vZWe
bFSQNMoh4+76A3HL+kEhSduvz6Dv/Ld0QHKDmZdKNYXydoOq60fHjG5QZn+Q1Zsh
YBvYbPD/X0Yps/wZnXtpi2uxW+oB/jJ3uhSM9iLQuFP0HeJRsxILohVihlWgrtvU
5RpZhJLg+tKQjBO7RE1COyevTKpmxGT7IGLlW3wYMAUZfG+W5s/9G3g+gTx/PdMK
BxlPPoJ2jtcPbDb1meK/Y4IaxA2Dj79OMYDViZX9PSkYvm59UIIzw9gN8gJeFzKK
EBKebAzjS0mievXb6QrqOrzw8F/OrNuwY1IMvFmGTSyHEL/uMESergbvbDViiH87
hNMjP0ttssw9JVKeMaO3ciiNchKly85xZppgto+PHsinBU1oQwzLmVajYndUGlQn
RVUj5OI7XQhbhIkGL9OG+M5YlDDNUMHhyZbJ9CXN+u1AlER4kGiu2+aZWrm6A7dD
Vi7bzz91iHVkr4DB0UomROyZENWhRFwnjhJ8RDceelGZ9EqFFzQCh/epMgTh3y7e
d5BIJ7qKo98RrlxEvFrFZUMYgkPiV3mLlY5+K/tuq67kJAP5NFQ7zvgysSdgmgUK
+6Ujvt00E5V3kysnqYXBv0HuBP4UgrVMls9Mvo/0xmwyke4PIRr/uJe+D+hUpRRt
uc2TywcDcyqhosxZyOBfI4FHZPCK1RkyKXGGM5G/SwUhVTKIzeLtg86rvpxFRBgW
R8xPo5ADgRuw1kgob9hRIqvZLSDwUqDH0rJypTtB6WDTCreaCGChk5Pa9jBn6POH
EMsV6dPiYZc79uqv7SG/j0s0Jpq8f0/8WhI1WcVd90Klqw+dfl78cmQ8HItHMTUY
fvAfZxUerVjpo7upbRO9hbluvb+kkUUsKr2SVbjntcuvqsFo4mrtgCBKZn8wq9qd
DlLfdJ2wl+D3Ul9Y+I0EFpwYZ0ooKSbt3AkLgfGYsqei9b0bHQsCDkdw7zFLEjCP
4YhsdxcwdcpP08z51y+cUNMGB5uj8c0nzWq3z/n+L5V0gb43/XwAJMfkvNGJy9ns
BICIFUi7feUa3+w6h/BP7Z/nNs1hwh5xPNSY+T+h+Cei7dSSJXl/1fZvKgIguz/a
i7SJ/rLvSlqH3K1lMxbyQEbnnk34W/NiV+Z4Fg9Fs20jid6E2ZjfvfS3pRvL0Iqr
DeW9BJkKLaJh3x4Y/cUpu6FaJyCWGUQqU8gWA+rfl7OoPPZc4EmEJECF6/8e3jm6
yqfhrZIcV80ZpoKTTDWoUsXJ/F3aYacmnIuCC9l7b+9zFzNcrexDjKHZqjFnBj8Y
wMZBzL0T5YZnZXNS7FH7dRpoW+RdfNHFyv0bjcq+lKsbfxPdP3yl02MLJGHNOTd1
EoopXzTGVEfLF/CRxBGnj9oR4nsTDIaeR6WzrINCp/YUVrsfowkREvtWHmzkpxzo
Ylq1rRb0qNPLFI5+XVH3Hle3IltUrqEzvlQD4JgqNiiXA57zZoCr1HC16qMYq9SQ
K1C57GcVplb7Qrqni+bUJTLHaF/UOnzbu/alwDQVI0q3cTtfgUtif7xjhMT/hdlp
XqUTBAiNQ9I/FFnpHeI1JVCdGak1VClMOCZ0tsZJ2j1HxZA7YhzkNX0S5d0sqict
4Zw9EiKnI3t0HCg8HkJL8vVdHv4r5Nf6rE9FONZxxkTK1gKjTBtvyNqQrBMhn1m2
Od2EEuS/YSnGupLBwcHBSCrrVQlER+QAJJeJnc/9LhhA9LjAm/EqpRGSgTSRHY+g
C2vgcuoX+IvZ2W8SUk9H130O8sD71poCm2CrCu8qB6m6Y/DpOue65R2ao4BYnWIn
sK6s4lR6FlF9bTkDzytKzSgUiUxYJIg1Acp01WO3w39ayMXEQgvSXpt2+aHd21A8
5ErCK8ZU9Kag9HcwU6ID42Hb+IszuT8hxsUsoQ+trm3ZST3hCTUnLycbDh+pzKn0
LvhGOdOfYqIzFxeRS68pAEl+9hLrPTid/EbBCiDef2Ja1PPpUTdYLws3Mhx7S5sW
PZXcVlVgFTzIKS2l4b/4ZjMvixKE0b7uA8DclZfWTMCviUylKYPFYGi45X2N8Mz4
mTmuAS0sGn9YjspWd29J/hJ+XU9hp2SCkC9B6hEFM8txX7C93e/52C7zxXgJN82+
B+ARBrrXb0PljMocFVdWwNlGwtqbLMDV5T+m8EsJfKbKZBJNfQQ1uRtDb0ub7dGY
RNGj4IKnDpwiZN0bneO76y53XfmJBWEDNti1586EC0kXGeg52TQ/sWYl/boUpuEy
z162wIjW+kGzr4eja7ojrn6Xf8FcbNjiRJabnKCFLv5iQOdAeMlgW4BJAS4wt04A
m1yQsarPtqsoc5yIrQgjNac5YsRICa0EFLG3LkQhlMbDPChJXyIOth0b64k8udda
4tAJp3sREIqNq7U7S/04SA4bwVMLaT+kLZ4xBSi+DL8+fnqzjdwnekDZHMsshlZR
DJ5ORlAttDVwVIz3ZzVWCuRVrMWRbmsuzeWB3P7HPFDk42U9XXr6PDrHkaUvs1cl
tUwfbQpgPnEtnDXryrgQ69yj54XXiCqAy8cVyokm6eq+c2N6LdRRqDeog5slgdtk
fcGbGg7gXOzb3suJNOk9u7GaThogUOeOgySW7GptQ/5+LxOVKnzbU8R67WS3Ubm/
wBTXEiN6yZlnVvlTNC/iUAL+qUqJpdGmOV52QpehMNCZhrsOqaEisJAHoC3h6iRa
fAxNXbcC7NotZ4znGupOCiRe8u85hx8Xorh4IJBnsAH/LBISJGsiZJT4jkybL0ID
d4piWFQgw0S3Q56hzE/lz2cef5SF4UZvJNvpZ8az5DbA0GMByoF1jlAYk9UyGW5t
hBPKPVkrpJm74qp8sG8PWK0wFZf+SdYaqGybt8OKt/XQ9MgfHqjxrdZYrKN+nbAw
+QbVlevDEn/0ybEpfuVHRQljcWMwDRC6cw9zkDuZ469eSZIKnIi/5pGdi1YAgogp
xUslr3wNBN2peMd4euCknwCi3fDq2PSJd4gNF868khxjA6Yoau6Z35nFCtFC1Qn2
jX/VsiOkgrwqGqUELl+jQLugcryec2AZ/dY6KYuuEAdnIXsbcA6Owd9bRem3gm1A
IoDuxWRcBPeLWdgczl+Ssk3hzz4u4FXtf02mrGf8jPor8GLfbnhZ2GfhPoU37YkO
VXmBwnrU+QXzSg1XwDdC1mNNtK1+1xPeMsoKUZ6z2dOp0Ih19k4XW7wDf1AJ7KWZ
pHRzbEzX5ns2ZY/DiPzEmOp9837+7z6qMocVs7ARXW4w5SzXcsAMySaNWO9jE++t
1WYBcS78qkRREqSk2uq3KMPrtS2Y6RipsEyHVYH6MlngyTgMtk/RAc1QVcmOCy3Q
h69C5hiup+MAj21t7KYdFhIcD746prJS+Cko8AcXoE+4kYWnnJOreSsL86zoNDJs
bV9rxHQaI5gyMH31qvDx+7AmFCjpChVG2/q+FAtPE7EFxyYDZiUKYX0XcAPK5OJ2
KtuUoTvoc3AikCfmCKLAcwYFFCofsWLCzs8JcHy05tD4Hp538Yhq4b/SDSwan8IL
0LVy1r+4a13I4LFsPNb1cyy/AMny30BzEeX+CHdNnr1GCCdkQA53sAoBM6dZ3rOr
tR2sAE7WpY+L8qznSTnMzarvzPcgOl85ApHH6HIBew3I7uvQTvOibnElNma0XhGo
hVsTD+3A5PMtKFHzCBLQqThVOESNIiHQ6pve7jqrjp5us6J6rWnPP35YCGhTAofk
3H5gFmmTOn41S7qd4HdUBIYSnJdswQcOTVbxEH43JXx/qTNvXgDmBQbVJjZnyKUJ
TLfqTV5gwQGYx9r3wwDdyJukR+tt5Ni4kDcnVWEw7568+l8QCdIsdHOQmHRMIY+m
WSi+XRfReMFjVvlJTkmUdKPOw5atUJA5mtShHUlNOOu0Vu1DJC5oKGLXXZhN0ncL
o1FmAFHGdhutFSKNOrJ4NxFh6kXsJrVV+BgM/CgSyu1ejLfxCqlShXbxBS0/xPpf
dM+WIIR2jfVoNwZqv4+2eYiDAmgYe1+ZqR4ZYcfILcAmElKEVp+sn32fV8NYZMY9
6fWUz2XiVQWaE30WtApdq07fUY7X8OsHMOGaxcH2H+HK5+1r+gDZ9s56WEm4jg+8
8HWP9MvFM2/4uT99Wf9RKn6A61EXJweYb5XpsEnY28xqbx0VtmrWe1MKHEwj7CEp
sb785L7YdqczGj+w+pxlJ3jX2EHmI2PlZNgsilH9BsOV57a+ut1g2ZiBOzpVCSOs
8+0Jxx2RFDbXbma8kZp1aw6ZdYzJxPFOww3TGjWMWKOogHe2u0OPyORUZl1P7uFZ
da/gAqJhmEAZABaKYY3ve/VUVV33dFs+c92y2VNZJMhV0fUA04xZ8lLcqQKChZyW
aqxYxKoZjTKAjjti8bFle+yCzeDxmnBHDWeFa2UYSZfUf0viJYbFbn1IH9teb+dC
uehpKV4tZGiymkRkOhajPgDcQo15fgMHH5AdHONbA4XEgV3HYDceyo8x7YSD08dz
r5EZSiLoZLqOxbrhlKoKpW9hgkvGAMVCtU7Le7T60lZ57Aqm1EEel//SCv01HxxP
WqZ//4rEmCKR879NVUltwtjOASqJGKdfFAFVnP4pnDMK8AKkO+3H+nD0+uIlWhIm
3G+TbKHIiIqz6nEvH6mdepP7Wmou3AxJFGcLxyXbdnwSGSZL45f0EnKSC1jPI223
441wUesX80gZqhhu5Onb5m8ZkuaBWPVig6RBnOzyHlbBmr+r9cxnzzTmonJJySkg
4JFyavvSRlwvxyrFgrGApEjQV8xKBHTFU3MKuxR0udSKpHBBzl2tq+jIk/dF3iZG
2btMr+xyS1Hw23uqJStUUSZbcKhqrtKyiRmUokj8swgxNcx3BdO+S9Q1zQCgk02G
ZFgT7l4O9rM4E9jHW0p4WxrupR9cJudFZQBwgOqc4VbrUvgmZGHNLkZ31xZAtc87
ryS256YQY833p9wie0BV6OoDrmd/JK7CB3LBhn4wq/xgzCxMLSpXNEyUV3wKlTly
nUn4czk1hDexoR2DQaoNpeUwmaIcK+yg2Hqbxj8AhZBp2r6ksbMZOU8esyPtTtOR
HWlc20t9NZv7wGilkgaSD5IC2V87encPyFw4bIzGWI4x0r5nebJ2kTY6VKb3S2AH
69S8O0RM23eHtvJM+DypltZC6TPjhTPG8KH34bVGR4XTzvw+uDBWack/dPEaVFfE
m1hQgItypMCX4b2PiwXhsDGv1lO3FImEndUzNFqhwqZBjAUlKtJyV/CINzt6Z7Ls
SEQ5CXUzxCIOIdZNB+1N2D6dwYDejM/bLFqo9prqFHpnpJybW6enwx3dStc114v2
zJefdgN8ArgmJ3t0eat7PhLIyPs2757ippamUxBgMN3j6GA9pdnQAnlzpTKuyOX8
2m4fU/yIDX2OIWY+pJUwQau6V7p8bYLKETRM2dU8T//23stydqcbdp4qxIicdYEn
VFCHG2sZ9nY0v81v23hKDJ59xjFLE3Fpz7KiVfp/REqYRoJOlv4H38PqJKCtfvag
ruciUz+vF1d/aaPkBPO+nWN3T8niOR/4iOVa1BzNOgeY2DTl+n08Md7Tu0vDAe/L
rjk0ApBl1XJyixcSrdR3tXkrDnWIstGKJ97JIjEiIeHSsTTbpoD3hrOKu90RLCV/
j1oDFmWHZJbA+Agnl/WBgPP+RYsJaI/3mEdqgW9ARQU1XouT6T5pldSsjEaE/NMl
xkUXpt25vvt6LxQkFKP9Vf/PG491nR25Ad+PqM5t8rH0Vq07Zfxk+f1WjxHTTl/y
pBX8WbAmbwHF+4Dwkn0c/NLNmmCL467VdZ5OBa7zQyk3y3yMWyCLF6Payufl+oXa
mqhLbmwm0SeBhDDEmjbbXSHYoZbuG/m6lvIFFV+T+4uyDzMeqL8PmKd073zS2nvi
9/brffnYnAEytqV+bWufY1nsaUmTH7w0t+/HjJ8cfFJlMwvXNhz6xfRLSK5OuqBt
8KbDyTOgprFBI3slteNkIGQuZCznUuetT/rXZSeH9gF+J3aXUJ7gq/HsqzwpyTWv
RztueREzrVbVXytRL1z348sf0O0eg7MSEREkaF55S5EDgGzwPKSEURUqkys3D4FZ
Hw0HzPUDLXzDaG/Coa0zDsfd82NVsUFHT8GpWXr90AU3MfWE9RxfuThgs7dYzC3k
uwiZgogO5/X3Tb7HAweswFvWU+JO9j0zeSDd6sPyjqZwbW9pSMzZofDtunvdL9i7
SaO/crGJbFLTOjesUh2adBomuE01z+C5buE6hXnxaEkmtYHxVUb7Bz/lSmGssiSm
61MZ1qmA6jCQ+mEVzL4lmdbK/IX0iUpxLdPjtCNwUgt57vnXT8RqPILSuZWjUibO
d8iNEc459ttZuecrdZJ1Ap6iEJtOxDpi1R4pEUVORN3bS00SVRATpr12ZVZnsouy
bNMUjJtBMItK2PZst0FmfMlFV6VJFvOMeZA0qCIH+S7uu/uwEFCfqEPzyNRYdod/
yoIj3DSR3X1e5MxonuX4b3BC2QNBAubyU04/0/Q48x5BBZsp6M0uk1tj9bzNsYEr
8VlldEZ21nsDSGJtlHCovxvBTA/+nClqsuHoeLh/3TNDpoq57MQ1rdBrX8VJHFXE
RlPU9HOIp1RKK320jNGTbtGzyt7GnFVlHLKnnzZ2z0Pc/2Lal0kuCVX6fbuEC7o1
iisTd6WauhpIhy1nxU/cJeTuCoNHtI6xNseKG1g5OG9CZ13VK1TECI7DUPdeqZb1
kfFedn6tlxGM5JBQaYaJ9Mvn+4rTKkFmiuWSwfIRg6HU1XIZEG8O3b2S5kTetunF
NpRkToFmngYadPf/U5dXSkQckjmS6hSTPJGAOGRk9n0EUiFq5l8xYyTD4VCqLovY
1b6iQmBwu6JrOdhqt/oUQiivWzlC80Yns6ldqeS3jGGTJS4bH5WT9fvo7hizg/Xf
GxPIl7PGLShpzMCy1qct1/MFSqfpI/aYiLQfWQWancxUW3YSzUxpZ8E2XJigdTbC
H14sc/HgIHtgHEwDWLJW0upUJMi25QuUFToOzJrCf+cJ4wObiqi+PzOu3JpmAHRg
tJb0rWLyij+ayIRaURL4ZgpsqXsgB/60k6YVrsa19lnj9+VjW2NU53YRYXJVUBST
Fw1ZtWwyuaCOMDRplC2CrXh+NMTxh5WY5ysn0vkEzLiZ2KOdDD+/O0B5W3bfunJl
wXZvPOKtKvz/6IPGbrJmbIFMuEPXekH3+wrWKknOhHQ3pu5eABS4dtzn/2yqf6DK
S4NV/tLjYVgZupMb8eAWYkgAnXFccZkKzdcQilrPlWIakQo/B4Fs+b/FIPEbd2XI
ydmXZC9t+Rx4fQUW0kjQjQqiGIDWW538onqjpBlZ4w/Br3m8wiNsxN1PwUqibFqa
19i/KcwukvQAADYiUXPu3yX+13t+ulpNnalgKfqkg1AW0sDjMAQlr1saI7xnNKDY
jJLi0VyNwbXqqBsQVa+9fLlBu5bTFOlVbkNqkeSGTBW+xS8FhmxXO+Qt7ucpHVBu
eCywsSbakpAs3ig6BPrSoPkDqOYeWPVhfo98UqcwYdtgqxiVB2RXu9TIZo4kaDAN
47sH+TYVnRjO77lIG6mNgQFikyNRi8cu6N4HDV28tkd0lAC7efBwjYUHPIP2+DWH
ms8GQLhIgmf/B5L+/LU7EqNalOiwjKLLBYSr2ttgLog2RFIMq7Td0NXBrEPBNdZC
krd/rPB7L+X+OISBVljet8T6Xb+HLmOnruNYNlqgHfN56biTn/4+nL+Q03ac2Ylo
6b4WkbA2igZRJrMeXX08eTodBjgeNWoaRQ6lEhSAb0FXdOw044u9mY9FzQ3cH0jH
sinwlRthXLu/pUrvKjiNtns4O1ZYSFAfWPylSFur/yoBoZt8QTREv5D+FArOqxcC
I4MqQgLRDCvAalB83wwL/HOpc2szPE2x90g+9d+q5/Rn0gE4XIeBU1CQTT+OpIc/
gYZGTfD4D+nkJQB6bDqtPAcVKknS0+Kzs0Zj0jBIPa7FHkMSZ1r79jVl+zPSQ3iM
bIljSrv1RPG7o6eZ9W4O/U+ikAhaT/wpZrBNLpPM+/hd+z5I/LdtxWbgsFLoeMJ2
J9mt9qCydwgLViLTboUIFZa+4UmvFXiiY3I7eZOgNEIqjvayBPqR+yG+PpQBVlie
1McpB+9R07cgbnfd9YHJZ470bh+kpELsBZMr6F0QDD++WPOW3tw1ylzuGBYBVBz0
RDtFuzxBrYKMptFM58dnzbfWnJqCWJlJCax6MqQDms76xs3U5yO+0+VaIBS+V6Qk
6pdmxf2Qo1itutMHsDb5eQFyhsEsX04Si3XPfHPeIk6Nl8JNjWZKwpOwCgaqgij3
D/F1l6a9ZJWGpdSxZiMrFLe9RnmUAaAadMr4i38aeUT+6QHvyLua0N0y9kiG91Iq
gyxLvH2DNIbhTO9AxjPFLxwL5OWzWlVJ8Ek2ZIkMfmUfQkrjmMtx4X8K6XA5jblr
otxoU3J/uLJ5HQZ34zCgQtukHX03X5ZhjFzWlfB7fBtpCOPGVo/10mvRTXJF7UG5
ccLN6RhYQF2LC7CcQPMikYD5lSsRa+D/0327XpxMT0CVdgXV9p6GNBNnlNkOV810
VDTdf3LOxmkP2u5cpTkogpGNcC/b2TvU0Q9DLuGZhmspVoOa/aiPgKUBNs+wiZXd
6/DKyc0Qs/iLAN4pI8qERPuKLoGWhjwtZpw5KzhPyE5EaC/SIiiDnJjXhvrUfgLB
Y+teKxceP3GHulb5/3rVUtXrBbzgJGantj8sHVA+2RDWjTjVgmm/htppN7RmjE1a
J/4tpJvHC3TIzwFrpE2a203jKBdJEZaM9zRzH+2c3FtRMF/2eAalH7G1glZ+KdqM
5aZJcaaSCiUe3cXKjKN5C1mdZybrHVpgNEx6l99TI/d86VWNCD0iOQ2W29hIzUs1
HhRuCKdLBYnBhVf3THd3zEDWr6OcgTVpDF53oJsbV/3f3AUlVu9nPJY+NS85hhus
aI9+naXLnTSs0nY5m2UAriDvCiSUsDGQU5CveFnZxMZxUaujoirL3xhf704yqKma
0zVvH8gxsQfzmfffwx+xd9LTx3ogbLoE9o8F1EEs2+82edFdwEI6GW6rLf0//IVn
CkHqEZkuPC4/NP08/pd9FFNrI+HSe7q1ofHmGVNft4JzVZhn9Tvk3EI9LG0iucPN
Aoom1+0F9gLLUUS/EQNDaWrvBzr5VzQdF7wGojOHp0EJirpWFTLpr9KuvQFos8NQ
JCAJntTBmoWBuUQt53Geo6FkxVH5se/haaS5vt4oYGKSiDYTHBO+ZmMs3kFN5xx5
6MFXEdsiBDnUPP0wZN6X7SmWnD+GdPJywKBSrZLX4eC1cQBqdweRycVPBjGtUpBb
huDq2KqW13dCucHNaRgOTV0w43NUh9gD5ltM1cL3jEI7WNQh648/yK3EkAClUN6r
foFgEFB0gbFuhI945Llen0ES+nofQevOIJPIIg8UxXKXnILPbpR4mC3hANW8imxJ
8MvnURQjLAdEQVohuRQl5ogs0WlLNC9br9W+GfhrwxgAy7Znl/nnZaHRIVVg24Va
2iJACALr5G9WA+noEO2nH3s0G4BZogA4Gas3VZM5GfNAlQYS7gcNdydbGFr6lK0s
yqntIM2kxmLix7wivdA7+qrE2yhaTUN/GQPTyRzszxumM9JnSZ7Trfg+BAlcToHx
UShNeuMjNZNJhaOfHK+cqj6Tkogx5MyvyQYT4XQTt+LeSMVxTsN5s7Xf+59nzS3c
ZbakD9nd9wX2k5ujFQ2ICCnC1qTdmWRdYz8gXzeYf7ufjjdbeBNzyEsfE+8Z1PIw
T5DS6sKJoiKNjWFq6CiwyHjAHfR+k1KnkGjO3Z6YB9+StmpX0gBZ3r+w2FNlNzEF
+UJNGyceDxYq9OBiFl6YCOis1/Hbvhu+og0xnvY9E0pd5hjPTdk8EB4GD+o5LzCP
sqQTeYuf+vnXcwbcwwd3C1RZ6XUYo9S/UvbuZVmGSKtnNZUdNthM367n3L9LZcKJ
bJJNu6CHVlwWSSMnIMs3cNzWOon2yHGZpUGZzth9O8x+2L+2ylIu0yv+SLeUuy4z
dRZLheKK9jYZFuHNxJDBHdpceuN+yFN9krapoe/8WmZHAtrzZEn+FyPgBfEMZvyo
SkUl7112Wm3BHe2hSm83r+Xq9ZqhaKYzgX41ZkPaQO5XnJ4lTFLNyDdq/eJOVi6e
oG12TWfPWLpbxjntzsYTTnKdQlCmt9YAnpbayKyfJsdLAEnZNg+xsVuyaOJuibFO
Fz61vhrgYooLA+DRNDt5leeVPm39zmUHLZ8W+4eaSmlv8+Z6JdL9/Bh/ugSiSN/E
7edSodJUA//nYQoaUjTz64ZkVYEeZEPX5EXEcj+eziYSnTnlPFZ05XXAP2uDtHgm
XCMRfHFve5ObfTKoL4I/RlN7scEMQ9MOifFUIpDBCP59THqcJ2VL+tiK3C2k9EhK
A6W2d7nU1JoVPKs0AsiRoBD+sQ3w9uqJy7BFsynFTHJ/nT1dHsZTnrguJBcMEaqP
VLZnsGZwdpj5m6KzQSTInbKL9F+Jdivk9CpG8ge8GwmTkZmiJzFLSyx3sxLC12B9
SUrAa/MTGZiYoMM6QtqDCrw+1kNPbXXAYpZLdMdJ6l5TzT9uUyJWKoH7ePMlbgSM
JIdAUiAehwHcxthh1r8jzY8B4Wbqk6sQDYMwglPG2scL6AP3++DEMssBYxmYFPRK
cY6AbxyQmDDLiocRJYSWrkFX+Q0mbm07PsfAc81yUABvcglonE849TToncjF3Wa6
KOyJwZPY1dqqdMnPDLt3KRnt3sPkxcKF9eYITLfZjlOCMBRaHIq4lMLJ7OfhMS6q
TRTZ61uETP2KayYQQTg/DgsFMeJL41PFYvdFzCWrl4Q+N7TCrvMnej1UwPdxk7b7
vAsHMQawGu/NNuoPnDX8E+I5+X0j8KADzBXwoYo/Cyv/dk3oOr/p4Nwyzie/y0Ki
ITDrin2GfdBywTZE+9Z7RBwCiRYA8n3JesRtsafZWEzUe7QXPiYpgAmpGymK9Cya
vipRvUU1nB1msz/XctjBjYkfbD6IjJJhJ+6+/OxN6qJq+KAWy1L2eStX53SLCVyH
0A7h0cns1Qiuickrd6YDGd47Vudj8IVaiCIWazn6YCbUDeEcN2CTqHUBuNxC80AS
KE8VO6sFIqHwbS9iExs19dZFYTBZdmCcOWaDu4Y5vSl0jEpPd3eUxF2kVP6D6vcv
9jbGSIo777Z1hgM2DlrxgaBuwwXdc9gtB4ESuCEScVMcNJnLrSwXQ+mPFIJuQOEl
Ueud0W4O1qECKw5MmuD88YJidM2qZc64tXl27n4JZddlzloJWsXc6kf2IeS5vhQV
+9/7QRLW1AoeGryxQFpOzgEasKVnyX+4DajYiPXdvugUdx3M5tBO332fsfJPtiaC
/Yq1BS9auI6rBWbanZ5LqXF5Bk5ICOkv77KAMv2+2SrmEXIbCCG5N5zsb6De7NNS
mC3WAXEN3r2CBwnyFJwGlLXvrnlNLr8FsC3O621udUYll7ySe/XGjJ/OgYboi/IX
oHeN0UMoAHPWSwVzrJ/ftW8XACid4U6kZJkZ5r+WdkGjX71OgKg5CmAX3saLO63B
d8EPBJI4W5J1HJwLUkZnTDRZD4xB0x4tP32g1de6n5dc4pVqyNYzPOWZ2Y8KIjZa
XbrKYVbj2hvgXsGuXEbR+C/Ft8j4b43EWeqG4gr+yebANCaVdicAm3vsdbIlCVqV
DllFsW51NFYvLT6ltUhOShBw7S0pYQyc13LuXZNXtAb1igu+xdqHqJROU3LSxI6k
sRB93PT+NVX6e8zvH/t95CNgb8QVPTy2aCZfvx1TBBnc5LqhEblydsIGpYMyGJZu
ufapY7/zyvNHD0MIU3hT673VmspFu/u+MPTfX9O1y1MIPLoMMRxVwICo+2fjk2GG
2R5h4vmVkhS+7Yum6N1RTHewZ22/gXpoDHveRQNWJQgzs1BqieTZHW14VX4QQzx8
iM5EuroyacznO3Z1MT56kA05oO1yZckxwsdlewWegTsX6r0cDh8A/LZdXu5JEpWU
ViX65tWukwJEL/U4gC4bV/umn91QeMrlmsH/ig+JfUy4dvlZL0/BJRaCwm3tXay+
sOnLCqhBPHGb8QS39klyrXjlzTa20g/bvgvxeggMjZp8iz3mXnQmUim4AGcZpCGw
1K9Dql7zPX9wgw96+eBFXFchvdbBOHUaC8gbEU7UlldM5/be8dlKX3PdGzUpZWpx
Q+i8V9HZwcDVwTL0JXGufVgh5a+u7lvG5muiLxm+zur5baQ/3qIjcxGduCV0+pgD
MeJ2XwHZejuogbUfoniECDmf9A0zpUMpexw9zq622LOI3798GWoDMFS4CEJIPiFU
YwwZZg736mcjYZgvItpiShnbTo6nmJ8yEsyaY8wf343WMRpZMbvzB72laZqcRM+e
VI7q+nxk11Kcd3LKWbMw1SKa9T7lZKuDpx6bXYOnrC4l1F8e61opyyaFauh1cWvf
HkYk51Iuvkn4nhnS3uRJDBdqyMKn6tjTeIHQbFYcEwcIOPidcfXcE6ZvIrxTWE3D
4Qg8g7w/8+VipFs2JiSLeM4T45X+m5zNmMKB6fu3enWkXiDuBvFfL5hb/WIozS1t
RvKRJb9xpYKgYFht0ch1qHRIQTVb258BJKwhiPgIS/dVjsT70z0KT+UYvogES/sb
4vE3Pzqz2Atmq35Ja+g8hb7dVSzhj5vcDrJmCO2gK3irzNhEn808iobTtfWY1+1P
OtuFRy1lN345rFGH67HXE+GauaK5hGDOg+Pt+nLHVZ/JhJHcDoqzMWwSi80mkDy4
PKkojG2utgtNfHUHrBOWBBU+2jBHAvgqCp2BkzRq4rACEi1Mx2NUTPGsiakUyZuq
TgufhFfjUsjgZ6ofdAgFmasdy2uUFcl3qRCyUJ+gDoEs8O6WOLC+LPpVqvHoP3UC
HWB3HyH9ZXARbtsARqO5rAiFFQFNMci4B9/Q6zxIbu9uPI6ce5Fq/8QH9E5J8Czn
swb38bBbAmZRdtLatdlJLC1XPntL9+Tamhuv08nyOmGSMBpU670j4a3wLnzvWLkN
t91/+Uz5LJggpAE5L/VCnDppJfllW330HB12kP1r5gQgJMTC30osVZvrL0q2rQOj
vIFsDfADSLvq+r77+9mSrel/avoLskcvoCRlHCHkPDUyk32jV7Dd7maoCS+JL3bi
yWC6rAX/xNZuJF53Km1wlVxwPqOiL4zkKXtRnhnVEUTNkP/LvFgYGiegFcfltRX4
QB53DjJW0jpZgIbC+6I3VSneR5jtB8ONTw5dxR9hF2krRt+zwby/gs+72BOZng/f
lixI8lpcN7Xd8zW7eYkFEi4II8AiGMGJ/nsKhHEDLhhzfbMQJFGBuZHpxYgyk0wD
eCgtQ1CKUnP4tIkF7D8BYEqZ3LEM7hzqu8YmrF0e4dLt9L1Y5s7Xu8RuD3ysvCar
spjpcrmsrGeXmiuK3ng5t8PywoCc8o7ZVvc0R2P3zUvXqRsz9GUvo7ViJXIAKZhs
a3MCFieCs1qNVdG+xFZT2JIGpH++2C7m2WTjk5PtdQ3EQXA6mtlg4hnQ8azosJg7
t03aFaUVgVrkCKaWwxqNLZHPujLTP533zjW9UNx1qH7DJtzOqdOqTlV/I1JbIoRp
WwApGwqoycjJ5Q0AUhotzSF/wcgx1VqDywKMRNyW0cBG49tEoPudXvC5e4ynCGED
8Ldl0/XLc5cr42aDdiyGgkBVShThCFh8pXXjg5lKDpox/kwXKunFrDUsPCpvMEJ2
o5GegTilnpRzIlu/sRCdDBBpzZN7V+Cf3JhBJvs0OeJNRrLTvXyW4n0XN4jiWJ9P
01heWFl2a/3+p+EMT7Fg//M53wz8F7FpLghjYmNPxGE0PrmhtF5Py7fAc+Sc6YtQ
3YFwVMK7wJI8Ad3dD749i8CF6TaS/jl/jYGbmb72wloHClPCtwM0G8gH2y0gVa+b
1nR+psv8k/vGgXuW3rqyL3/QXiQI+ZqfNbZYb6Y0AhY1BF+D/Q7/YA8v8sXys4Ac
mfn8jpUbL7T3HPuBluyW/kjt/IqM8KL2evtTkfPTudz9PkxtM7VvHWbHdVhDi/YX
5c0T3MCgc1Yr8ZvgH0n9ogM6EZpMPT+Pw2mnRjcy1jBDIwmDw/zieo2M7tLwy+zn
WxVAL7lw8TkY2b4TxtBvsoUBOMweg0LpqVPdIqC9uI6rw2/ocncCLTEd3JR/h6zM
YUR/P2ZqBi5i7a8iq51xpWx4dgvEaPKmrbebUq313lOTGKiaSz7e/AI/wlrYosKs
TjQj0GHNkwYEzO5mVPTlnND3mPH94L1LDfKUBWDkYu5O8XjV2Fj3OornFuBaewW9
+TluG1XvHyGyT8gPzuf406SeU5GK87Lb/4P6moUXisKXNR2M5VNIKvetFIQi62fV
jfVGk+vU6ErmpVvF4qEFv2D/0v1OF/Es1X3D4DVnWhHEXmFMqP1K3BkcRL4HTbzO
+B1B7sFZtT0awc91eAeLESSob7dYQZspRK+jAxxS8UGDHAvdN6uAUJ4m8iSvdUFl
rn8aj+DyUtC2GFZ/nUfYBW199U/xCk5sKyq7XsA0RN2jlG9iIq5GJ9s1QsVpRjXy
a5zR9LTu1pkRfH9HZfhZJAl3OAv6pv+XFrub2O7ZGwsz5k4aWxdshXLPD5GHy3nY
w2lFSvMtPM3iv5kJ5ZiQR1YwXzSjXVhu+h/vEurVUwBWOpDTwiqsLCHKHAvLTYQK
fE7FTzADkFEoNGwd1eaL4NMUq1Rndaa3lKXC15A1TLH5YduF9gfkZe+BVINtmWJb
EullMb48jNyg47RkHhZXs88Bn42NhTdWuu5/oRm0c2UsQtv/fWptI+FoHYuHaQq6
ioNO1RwJLfpJageRKPe+v/QerANcroq2k2wGJOzC3Uq20LtG17e3bqgidLLLGqQ3
wfXnnkT3qzYvo2tSY++Vt/QWCzYU7PYGuNLtYRgeb77LivkweUIgpuaBMPx1W1PZ
Tjy8+JQDuEIPrs5MhJcwJb7d5VCz+9rmydU2N+CVjUOJeydBa3JWIHO+o0pD6NBx
bV+ZQdo1ApKk/bn/2FwtZhhTlS6QdUCRL94F/Gzf2E/cC0zj49Z13tfptrbf1GDF
ixrqov2Z3syNKblFWPazHDKuzEvIXI7QHrlxcMjOGN6I/9pd3wk300q6fVK1OeXi
DYcZj1/1I93cHiqZ/UH/HN+3uTwRLnrv+VRe7AY66Z2LoxkZ3c5fHwiVMw5PW8mr
NhuHG8Zvk/kXlNGM50hgAxu59PS73t/8OCs/0A+nsTaP6otzULfz+jUqnZC8MmBd
fjgo87XBxIgv5f/5UrInlMebcFpwI4DS0soIUQ3FRD3saC3JALkyLTD7WVNEBTYz
BhoyqKqGe/GTHrGjkfMpnPPVYdv1oZ/d6nKzUth+raDkU7O2gVn/bpk76J2Xx3Xj
i7dqBmky61IX6RjFERSp2u8o0U63DQCZby8PfiImRORAI7HWDWmNrfunruL6wmDC
3UWQkwI6BcBwnNJXWbDvtIGjDSNmMfeoVIag+x1vLPgypTUcVP3UTQFpJnFSEpUe
`protect END_PROTECTED
