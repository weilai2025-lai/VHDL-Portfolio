`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jigccYe6YcWr9rO8nYT3ojt2NxnoGQuriKjuB/GFe4xpegK15x67RKP8ZH0e2Smb
hIIUwvVQ9HwPzBYn68+lE1fSNts1foYx+crcsukrOCaEYZvZD5BwtWzJfX5UwyrE
O8ths7ecimXg05JeKxiV8ENbk4ECViunSey6QZ0z6OM99ZFRp72Guwg60KZgD1eb
MCwXr/0b/aef99Xt/l0I6tFy/J80jaZ++WlRo5Um7cwGcczJtv5Ts6kAvelRfgSM
y/Abt3LNqgsxe0eMl99A0aLIiDLtHt/pZ+E/4Zy+IL+XQVT6FxzN6xsJwGUC05VT
qiFYvucy8Gz8Ff9hi/o96/d/1/KnamwdUP7iHKj0gAK7dqqga6HaPBYu5g/h447w
XrdbMYMYZwHiktU+QMyR9qVZ+Mxw6DZYmIcCLNOwOdsqwrL1hEOXbeDcFkm6xHrP
P3Zy5ex/b2y/1TwtL25IkG6ZVtFPpry02Dl4vcraat+J6CE9Opjssr8Wl2hPoVV1
aqjsPqrY2IdmWbxce1YsvGEraoy9AowJ2M1yBeJ0BVQHDdhO1SWZLgX3N+Fj1YOd
SyZgne6iWtHCDCkGk5vYXrnTWWAGGWSO4TPjzE/3gJslXTCqI8nodpMtSQHQIKln
K97Px1PB7eKZ5u4BICr67c6zh9QorxQA1k3kjK7N6ioGoU5szEKabGhBCa/qagJ1
RmBNPpUtPQkg1doDqTF4Z//1qZn6EY50N/b7fVFvTnwLoUnJx95NNYXrtJ3a0cdI
BCRVMyOmUTppyp0UoHqaf4GZawRjQ0wq55VDXUzD/wXAUV6+D8CWnOWKZ6xD3w1c
UK1kFgvoYrO8fXI4TUjJi38WjqlcSNpu/9KSHy+nnVfcH5KvIKiznDpdwzlhySsP
KOkg+F/z3qusihNOPrMVO+SlY5f1dQn5ANgvzG+VOWOgZ28OHYvSLTLS/KZlA5M7
2F5QuJiNVgnxcZoqE0XbwS6WXUKkiyjwSyAvctIUl7kgRomci/I77IfpzMp85Ix3
3+54PpH8PQn31u736daTK2m8y08Zo7zNq32QJhWExQGp4zkI1jP3YXCQQXYY9Nar
6g708jTSbmxC09WvSV2QIDQ4lnUSYwjbYfGtblV2Ib33mimVbeIyuEabq78sqUo6
llTX0TIsui8oT0y24zVZ2KGoKCJyqZSCo97u69K35A/fSv2AMpKIbG3sKVqEnwu1
yvV9Y9MNF/ZDSlhvLcxAslAYLl5XT5OMS9X2pcNSjf6rcRvBcDtkzJngMlaym6N5
7OKXlVD+a3rjWo97PFmQJ+HBvMysDLyR7dhSEHqK5QTYQHJMLHsyHUZDf9P2jxaz
2owz5q4hVJM+jBCliLPrWCRvgJmRHbNTbm2m6eM/acct2j+vzOP9pD9mJBY8A1V9
V47b1LfeTCGYXjrJN+70lMgBgs8l533n9ufcW/ZOY5KlIqpRsrwDnW4/ROdd4bzn
xnP7trCylqYp9HR6yKaifOuexUao2srzAWLvrampygE3ngwGyFz5BPYbNk2K5NZB
69kGXzpe2pnunPlAuXprDNv3lNOKyt5wtJTHM7gr/U631VQN0YPVmFF7sDF8yGjy
FwrIRWCClSebGjPmB6wZSGpmb17UkFce1mCJGDMJ7wduRGqv0gGokUj4jcucYZOh
pU7LchV1DsBik5NynDWI72hr/9t9LsRdolbJot+UlJmuIykvrPhvQUnsG1YTKqa/
yu9EttrkEcB9HBPshVi5DKYSwJZ3eH2ctgIqHsnbVRECw4KI/tuAZA9v9FF0g3e2
x93R67k7bWmcNW5Mr/MzGPpFxZVblKM0rWDD75oLwY29VJH1HsvC0C/NIei3mgHm
F4hrjBLVnsJ6/tg83TUn1i5t2rxQXtbNT3CgrznhL8aFi3t5FgQXrh4bGiT9ICVg
LKmQvagLLwVhTJsjzOrJ/oyyRvPsEyGh7XIKCeEsBMmADOOCQQhQuX/xv+OpyFQv
f193MiWUxjbfB1Tm0+aTeNCpNMXgz9XFmzNB6cUcaf/qdrpuCLWs9oCCqldN73ww
yiw/jXWOAi8961UTy+lner+WL2479SL935MkMPWap7xEoAMMQLD4Ih7RcaJD1JzI
5uXTqejd/eI2mlK6zen268BY68y/NrvdlVmC/5AIxBdRmHdbXPslPkC7qDHoC8tc
NqQ4ra+/eVpo+czhfmhAp8/NDWVJGtCGFOzP7YCm494=
`protect END_PROTECTED
