`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vURVbIHftKrKerKTAL754R0aEjViX988fGx1tyQ1CmymMQbCw9IALOxTZfM0lTwN
PbAjwCv/fpxWh2SEKd8b7fl6zU5sISUWd+EYKFwKDC/JrwF2Ig5QBvNWWYwBy3+k
8Sye8uzKyj63/7eqz0AEJrIkbfSKWNrxv2Sf5slxRcFfdNIQCNC+mTgKvgA2tn2h
kG5Z5fbaK0jet301K4eE8If6GPcmN1Nc69wN+Hj8o/1zWzvzGj0/5gtQg0q5WxvZ
mv+uwMBfQVA6pP9nRPPhJwnan1LVJ2FolSrk+bboOjVQahD6+Xu5sRPtB4TmDeX1
MdO0Q6NCiirYhAUlsAePxNL5fffEJwerkT+0mmz4ogP8ZkaCVaP/PxNqC/59Vy0A
jNjZFL33gl91AdGFbaze4/uA9JxMIDxIkiBmWDEapBMHlzY1wpX2pE8XFhwe6U/e
UfW5tBmX8J+Z7P2OrZZsNSKsz1ENkUGmxpNaCD4nz/LjQiHyBhNOoHjAHDekwjMK
YAnvEUgJU7zWhKhqmG3RMIf8lMUjbqP2KWEJQV/RF3QTB7hg9AC9XLhAG6wb9zGy
M5BkvT4tUz1D9KNuUVqWWqqGMKPHMIYFjsYxUeuHivOnrYUrWG6llhn0nzdFlSmF
PqJV4s3VL0e3e1QbfSbEjdP0J/gJL1EULSdZP5Uwd17YBnk2sK5oRBJ+4zfMLWzz
Fkm5aL+my4TQqJfQfM9tXLYWJnevQ4rXLnk2l/I56sl8iXO7gPHtaF0M/gFHarlv
07mPtqwi1fEeqeyg1KTCWuTdBL7KuyQqe06aSGglEP4brSQL2BqTCCwwKcJgvN3a
xGDEN3kFDoujzVmOCAF3wEgtGANDAJqDaDpEb1JJd4BWF+e0KnGJol8Y4gRbJh98
UJC9r/xD3rJj0ZDp4swyGX0ln7OgT8kS87CK1sgIF1rJLE9QAlC9GSoBDZRXjb/S
8kxvWvhLSTojd+hsIIzFp9srI63oFcSbDoh6yInIkTXq06ILPunR6ZCQ3y4XwKDf
N0EGmkklZVYM4ugME5NHte147PR9ge8ITWwUb9sKE9w1xDF5a92hVntzit//Y5Th
GvpQ361nlCLffuyPLV1lovEnj4hSZkXaJ4a2UOY1M5q6COGMLVXY7eVsojEev+hQ
w58rDP+CQaYeztkyZaGT94dgdLqaIjAx8xdssdwqB4Wz/rxU4knDkTz3q4LDjRow
Ys1o789+nXwGPZ2/AZKSyyBHWd9cuhWQJP8h5/ITTyZgIMKzbiYwVvE8JaztLVUs
`protect END_PROTECTED
