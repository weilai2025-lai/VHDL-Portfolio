`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PNhEqyw6PAvKgvuFMnGcSgM82n/vWHpVpvJkAG6iM+IiG1UYudcu7pYa6VvEzUmT
3C6tfmTcRM8LDdBei20TkHtMWk+C4+WwgowDhqOQgyvmSgitEulifse3d/8YiqL6
net/JuISnOpmf0k7LKyK25o67FzwnScmQ9jVySz7LiA0PMWCte6bEHzyvNjKUH9W
fgNSG28lgvi4ZHc6Gxr3Y6oZaMyY0aPPexJkwY6KGghy2Zwt+kS/UQQ6PU7OdYGT
OKzFMXMDqK0iWJxFZVOZ7OcWbnpykN4bgc+VuzLUsLWvH2cQL/vWs2RlMsxt1md0
egSflMZ1l52lPgksa7j56FNGYDDqzWKYqqXuBKDrZQp4qkiZVTSCVOzFcfx8vZXB
PbwM07/1YRvcstyaEgD76qU5ailWG2KyTRZX1Ik1SQwrpRbwk0rouXj4kRAQU5N/
WkL+sQGdL21S73gM7SmHbfOEDe0WsPDQn6yd+05AVBVPBX68iq0FDf8KOc6vez/t
34/jWVPxvEODMbopSaBmew==
`protect END_PROTECTED
