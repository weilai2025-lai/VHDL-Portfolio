`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEELM3HPkIAFPRJF6pp4MHZ35K0E05Z+YanDXRMh1y+xc6J0gfZy6CgHANQiZEuJ
1MdtAvK43V/+x//D3/56N1BjM9JiuDEVZ+QyKfbyz9s+bKVdyGRS5iQ2Asu8ydR9
hzJWKl6A3pqhrgcnO/xosJxv9xnjCiiQQUDPHt2wiItYNt99DMD9/UG6OCUIblC2
BjkYErajOX90ygK0P+q6niS8cReLqqMzkcUZDQVxfKV7IYYKXXuCBxAuIbNW17Kj
GtI7KgWHpiglkE7/t3+ofbaKaFxFkdqLdh/ta2GcecdfALmQ1jvUO1Yaqq+r8ohD
UtriIX3NeNzsXSiLnfrEI8OvcznGOUyysaQUaF0oHF9rxeGivX07s7hb9wOVZZGu
wK8uk5xqx+CCo8yeqdpxF6pHTHpuc+LDSBqPG0G+tcCznk6/G/D+2M2QD+OHsIGi
hkRkqabJbzrT68v7E2o5tSLScR7MS8LC+6UI+kCEmyHfM0nr1NGomHedbCXGxCGO
3LeCe1SjsbyrdwhQPrzNV7YSdGJ4vnyCQfYwZ0+jfw31g2FiNZHHR4dYaJ08cU26
bXQRvD+cMm30FRYO1jBOSWM2xvhDXyX4gAVfURVQxpxDqhH5KNyGxyegovcNZw93
qZIMR19kF+L2rcLOWwNQA6k4lRRUTbFED4HN/fJFJU/RGypzJj1l55TyTrfmWZ4L
tUxhWgO4GaWL0YgFKo05aZ2aLiUwP1FFTIQ4w5Yk7OfRx6rhNXWqjMEAybUtxHqS
C4ubHP87jK+vrcunL5r0s7qo3lDLjK2x/vTO4xwazv8ssDLVfYC1HmXfD0pwJnwY
6+/Feltj/5YteJDxj6UY4HC8aYlhYFplE/WrvRXAn29N8PKomSGQJnXvg8xRzajF
pOf2IeZlmlW2SmEAxF+zwjtruTzkcYbWTwusRn1tX2s9JEwt/Rn5VmWTmrgFif9b
ZqbA8mkclNSEY+xxGbMij1DjHDqT+ZborspyT6sD9P9mN7hM36UXxYAa0I/o23Su
uG0Xprtvl2GCcaD8/ULWnn1w0WopS8SgBezBhlJSjyv0FY6biYKsVPwLAAGu05mv
u9gC9G2AYdZg1Gp6Ur/e5QNgC782Ancd4p9luCH5iOc7GmlGT6NCJG6YhWlh4Uhb
gJ0831hepKsoOOzXeip6afoeaLdZxosAAPsAvRI/qf9FV/O0ib1IQClR19HhkFwz
Gcc1JZRWWQv8BICfcutfgBtO3PDvQkXRFg11e/GSQrc=
`protect END_PROTECTED
