`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ndkaT42RQQLUSmZsIdDqQEU/agBa83cfR20imZaBheAUdQ9yka2AxmOocnzmK/3
j3JE55O603wc+RkSPSWLDBWqgekfyNgEZTtHT1/hRwxTdLz5BaEvMEOEGw7LNJ/Q
BzUW13tiCW3AuEVAp0NPEgJWBIuLaFROutERyVU0klBjmBACr6Wd208qtVUrhGFt
x703U7nRGZvV66/FprmQrPbe+0dzL02mpPc6Bx3wFw8hEDrqLEWTPSsc2cSQUHuV
uplBL7T1RP6kz8LhE1ulgP+tQ9Fg2xV1hyBl2CeILFFH3BZXRw7Mo3ORRSTV59NJ
XEaxCEPTxuqo16HFHnehWJj9yxsNbLkALBOH1e27PfI/GHqD+J5vT5Ddk3XzJs36
lXkWAuuCB/7DbxuqLLUFa3flKsb3nc6PARem4vRPmhh6ibH3snvupuxmQ+bwq44/
`protect END_PROTECTED
