`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rtgMuxtKlukhw3ONgHnAYDLB6CaV9fhZCmi/SzCrj3opsKzCJHGpn+Czc/Xa5BKs
89pusXrCr63yLJ/DxGv9U+bMXd8PgaNZ+h252IMU+pxQS1DmtKC9MVbkhWMs2wcc
QueWIjmOQBOM6NUpsiY4pnSEoMvBMxlj1Zf2INrH0MDI9lJ7w8hKRui9iEzP2KRt
UcZN0s/Z4iOqOU099XV7tPtTyueJLdeT8Iqc/3bC6yzVY6u72YAtU0Hi6h1I13QL
YMc8S08RJF0Ytw6yyo0hoj/QdQYF/nWPn3hYCMtjb6y40ueSlSkuGkWnVAVwtTV+
RN3lioenV/fggvTc4AuPHh2dP7aKTbA+pJZ21YkVqB+TWWmbJNVZW6Yha2r2Wcg8
Mq4uVWVMYF/tDxONe7+Sp21v1byz/f+PT4OPRUakP9Hd32emqgL4XJukPc7j7gK8
D/vtv0jlrlKcp0rblGjqHsxwqySJfvRwNBQKdHJEYunzAwlFPwnr4SD6Du6BH+QB
cqRDDMCZPkgAoUXET38QzG2BZRQHxJ+9CRflGYUOz3DyQshsOz9rQGTX5rD5e4Y0
O+3UArp/3J9YhPBQetQZDZFdzxgXc+mQXzL88erBaXNGmMSbqSJT3ygRjPV/9urS
1cIiPCQszJMCdpJyoDCwN21TpZbEt0S/diDaFjCYIO3KiYo/J1t0nFhPO3LgS5yd
+7uYsNp4U1B+E04RobqEmGTPsqK4nqAw9+/EpR6Qu/UR5LG5w7coeYzvSViR/QP5
VHd0n3+1Av6qqcd/c6y6rq+qRJW8Gx3bfC1qkSF/IrepU9DjBUSi3jfMMrPaDVQV
l0wBRxBl7HtRy9e6XXRBCAeSkUfHGXMpFXMo8Nvu2a/mWGyfLkXCy2UTEc+unngM
7UaytXntbqkpjvh2W/RsaoBijbxqgdrjEzFO7Ome7m1oASeRUnDFV1Wl+bE4bkTB
BWWhaqCfXuMdOKTb1YgKmMMO1caBd0tg1n2hZt6UdcLs8BcxJAQ0KoJdf73R0HYS
y5y+v5anGOGruOfq+75iFk5i5skCUCmeGD7HuWwVil3DFe+XBwp+FGCHZbd3ovbj
M9n4rY+6uY6KZlo9zeaZH9hAYiqd5v1UxSVhExCguWZ25fPB845iwRHdemooxmnb
ypNHe2c6HeQjUDl+eGdffKA7zOyOE+0bvwoHVHDui3XCE6IT1pbiB84VrsR3Y5TA
om1IuSpJQJfx+ioy+gSxq5/l9KH4JXFo2QnyK/TkU8g=
`protect END_PROTECTED
