`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQeCpFnupr6IuElgFlUDlNll/HiQMCofq+KzAb228V99W+gIn0nVJDrRTdB9aorL
FL6m5CQFzE04uAJvhLBzHsB77K/Aai7oykeShdjMrKG+avtInxawVaAldiO45mMr
90wmOjsNsR5aTWmOjI9uDqZcmc5VBXJ2IBo5R2+2NTIzurcVEcgvcY2PzaJrsQhT
gKwI926/Ga4sz+n8OLJsH1gvZq8fXl0HgFI5enR2MmIneAx0ehdYcDSrdGSZKgmO
WIkvx0u+Dtwxa1IgAJx2qnHutC2hZLYLdJVfgo0uHalELiL9pUiyY2KUjV7tvvLo
deDjrPxLou6RoKO85QGmnrC9S9bJDgg/Vy7vScZnDGaD6u16fVDXt/xbcWspGdTj
xkZUfrP5k6++jYKUsm5R/JQRqNvH5noH9avz04vIZrb+e/4RMw7YNfSmp6CneO3F
lN03JFMunk4mi8nV/6IDeTept5ldBpRVE34vgF5ixHKHHULfbke8UTeRmjmlT2Fb
36+LT4zktMU1LwbX4kZxCspXmgOyPhA+JJ2pFSxzBFpl2wxezwnB+bM9WdnGBfwy
5YU8BU1y90XYXAp/kf1ScIiltEehlS7Vs5TBW06B9KN0drQHg+D2ru6O/bwtvHiz
V8e4EcJygrJsgB52fDTaNMu67ApYvZo89DxUv+WTgmWqGvflFQCAKEV6/Qv91Ge8
xEVHy1PynipQg1Jm3M4KMle2i60nu0Eg/OahbRE2L8JqJjqOp2ueUtTPaMObv4Cg
j2E1pOkEW9JBsJdcef9c1k9T4cLfYNG2FTmJ4E6Ys2HtzgWGXoVZTx6bf7BJJ6SN
wzRkYkwrtGIsZkFHDjJqdHQuKEkurLzIaZYAeQUPqKDQzFV/xYq6yTYBTg6r2+kj
a5LL3iI9raAm9VE+6IzwA9PWxt649Iaxh+EMqqTeoZbPx6kR9HfAC9WrGA9G4vth
QJNnlYHnEY75uBfWOPm1VuDwcGV8IvPn4jHt7YpZmemkeMfM+W1h+ucAr095SqvK
IwibPnw4a0urkgmrHR4u0ijbPLogjZ8AyaMfqK2sBhKMfCgx/bwwbOvPh0xGaUyc
CHrrIfADXOL7VetoAjosWD+df8GXtCOjLMmJAKRf759+aB0trniaueGOzoND9Noy
H/FWU+9kFwnaK5RYLuVnQ1Yud+hFB+OqGIsXr6iUI0vvbx4vFieFzSNyasAmCchf
Pm4D0RbQ8ObPD0euslbXc/evtxoQk/m0cfWmm6ITF4jj2Ip5S7srUXYUpr1ibTUn
ZheUJZiR7yKsY15xeZbLs60RxpwkG3x4ykiklybXbo2HmhVDOq+DzcSIFdHU8Mw6
oiOPn9WZz26fIMPkEQYeJtrB2DcsMoYOA7boeH55bwWcLsP/51O+uZv838Gvl4RL
P+BN26MxCzc3MHMjhhGL23Q+VDMlHxaY0xr569X6R24k9iyMnD1+dOUzrFuTJxA4
BDPNIt1jZs4YTC4tIdH+8seS2Rr+5dbYfQ1SQBuJSEVF7RzerOt1GuVp7VIWLJxJ
mZ8+Gn4O+m3aRsescMpKOu2o9vXgwom0w8FsIFPj/lIEWrMSviiA0rbYT1Y/3gX3
SE1Y9K/sC4vlYog694cMz+CxR+NnPssw5Jhm7QT2bbyjdivnYGCXF/oTrAYY6vNm
cBQbfvCmLOOufv+wIhGy+Y+XslEcJKCuIsrBZc5bDe1hwodM4oWyZ7JJirDpqWyZ
s4PL4zAwm4+hwqQUs1BbtSbQougyjCwPVYJrZ+pprVvQaa5O2VrzS4A0WVpvu/1z
IoYs2hn0YOFegjQ/YF0V0gATZQL36nGN+oPD2N6SFAHVpP370nilAbJ8snQbJDfN
Rm2Lj68zBnSuFCMU40eIzFC9wL4YVRUWLaerhxlnSruCZWW3YqSq/pPY+YLoGKxa
jWx3nsQTIY6lU9VV92o9qxBrRlA7rTHTJFYIumz0L1k=
`protect END_PROTECTED
