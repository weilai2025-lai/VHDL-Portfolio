`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BCxe8KduMmPoR6KDo955oifwRVUYQ7tNCRXx+MWPDWbQB+yd4kSoy1lAjyo7c7Os
Q54JtX7x88VeeR3Ob1s8uHRKfjV/CKB9zA13XkntvyWZaS4P1zYUk70xUiOWNIl9
5N+eEgcdVgbddtL2TeZwZ8haDhrQ0ENCbczrOTVuNJ/IjXBUhq6ziLoDiTtKrlKM
13MtwtqZQhTIROYjfMGYD9ZNcfhUyl2iPbPoN/NwNVo/eyAuVgF0VSRD+ivFgdV9
r7r1WquejFOud9YIElu6poqa75LUaUVDvqzY7JH0JQGqasmij6ccmDukuKoskMHm
fHUGQmzS4J3zq8Vry8HnewE+XcCih6+cLJmIRlOIdu0KVpByzzqgZLGRDY7F8g/h
jCndgN3sVpTZ20dWOGgD9KRxptvXVrOATSXR4CxmVVdnr46nJJ9Jf2HZuRUY9nXO
nJ1RPhfedX73Qbkw1swElQ==
`protect END_PROTECTED
