`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/z5LZHLJr2s+RbitW8NRzJNI9QubTiuFkDPjhrP6/kQeVl8Xi8b/F8ZTe2cQQslI
FWSZ/01hvr5UAXFtl9/BjCkkLLxfUNaeoLkg3/L5MplKYjbHS0awCSzzJjiEbrRA
lnoAsP94i9nvjXnFbXRmMvVThQ6XPq+CLQ5OTG3ekTDkspPf6kRjb7gSH/XIRmLj
`protect END_PROTECTED
