`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WYVb/99wScodEAQ8AmaoHYHmAAIST4lZ1gDTjfQ+QteixmmcvM2WzdmORgGzqS9D
/fD7bzmaBY6P4xXKVFjNCXJd2VmBOd099r+inZTW6Q/uyIlOh8diOcRvPr579iIl
A8+nWi9gJSD+hdowRQ2KHyvg/BLpBn8PR1YzKPjlv6xREs3NriUyhnqLeTD9WpAf
xHP6yjAi7HqlepGTnPo1LkqvcAihdORp1PeQzvW2ZEdxgeRUNmX/CXHRlQqI2me2
XM2K8NWWx7vzcmZfGqq6iNDZMYwfhxAlGuaBRmfb/ite59DNroiprsioAkJDrENf
je0poFmeTAfNpFvVkvLlU95Mf05NJnhjaRCMxK30V+RX9XKJDpFRZpFzmnPNTh0H
V36wgW+sJz3MuQgzhNQuFyG5OnPpY5qmK5O4b1/Nxi2YFIXIzXk5zonqMON6qp5m
UzpUYDPPwoaatzejvpYdDI0sZ4w5++fC7K/KiYPglmsqaLrH9pKRcLVAA/nGa/SG
4bV7KWfwPLmVpE1+NFRbynioZwRQqcSjCZMQgOJE1qCTve66lkchL68HLjT1vTg5
O74iY63VwJHa+1LHaAUbjc3b6S8o+JGwdmnamCvVNKJ8zp7t232o143vRZjEsRHq
ERjRIm1kbKiGspSAwXpO7i82fY6vcWrjgY/4tdNJYPXHGPMeqIUYOtAu08P9TSaU
RRMHVPrXORes0xVpGmqYv+lylSkadFEMX/UEUhx7WEUg29ccgYr9+w46azdQIzLM
RrFl0H6cASvBS8d5H5lbC+a8lGbFDijHj+zCZnKhXAQxvNtKYjR5TFvKGn+xDdsB
HAqTaPJHRS5sS1Jat4N17JrYCgsEaPcm60eAslhho35n5AanOmQd+dCrc+xweLv7
DFx8sPnULVl/Tgq1lPvTr1r0rA04xq7yxVda5Z7eN14KjYhBR5SraJbHnCBNwJoE
Jw6Bi1J8KQRvZXKk23EK/KLTRbvt2TLjGFFi9nujOxlkUa9Zg9JPOnIHPSilhj7s
aJSmAx80L8DNh5sj0K5qHAmHZsUM4qGMhTiGG2Y30U4yjWj0Q0BfreJbb73CkgOC
/OXckfBWcYzcgKwbj440i3hkEHzPZLFOfrfKk/j6AJdNcXOvhrZFob8SMEpfttPA
pfXiazbfdZQvK+NkYAwkmpDFgvIc5lxoZ8F6aBN/u4LV3p035drnGC68cnyGUXFi
jHhjAk4OfeuhnTXo6Ipec5esYpsU9ktytC+8BRUdS4Ivd72dAjjdptZ2NlnVG1MV
SMAPXocXhu5xzMMyYhGOyXRar9jG+mcAJhhLqia/cik3P5WMMUwZ4oV/muatq8a2
eeLGND5W+uXsXvc1oqm4pJwfBq9nN3shSwgzkTk0KpLVpT0odvOFzvFYmqACfeis
xpzxIAWSZjuFzml+OCH9y69trP01J2VZ6JGNPHF3PAE4nHFVMEf2mULTfwYr0X3j
xpffXNOk0ln/n328/WtM0p0+rm4Mc/Yxk/JQr3/DOn2YY5fC1X/NgFsWErtl7M26
MNsO5C/kMPKSo73ZdCOlPfuWIr3RuvxSP86bUzCzuUBgNmKfq61Qk2TQIX1iOLNQ
QncvSx2/GacpHK42qWzRMP7NYrqxY1KFZj0EDSxHOytQ6LISpX2/ZNJivM1GC9FR
d+Y+1artlzdaayQpvplo5o+6xgzeqQUCabUhFWSOETFOSPiK4LZxKPZG9VS23nIn
1/uK6AYf7aMGVsskhMe1YsEJxZJj/khY8Xm/NverpJmwAwaGx0lUCTok/nfSiZJ5
bJiDpr1nTtYZmrvTK6ohGpiSLNkBBk2GKfFQeCwmZw7HamRPuU2tQlep/Hs8d54u
SHi4dfxI352m1GtzUi4LuB6EHVtleqqVXL+gk79tNpjniWn9MlfJ1By2uzPG662u
3kY/nMa9I57W2c+Lvnwx1Gl0LClm6d+whhofFCwgVld8pJb0nVFUf+p7C+QnBBXA
y0hSf8xSDjZbC81yNtm7M6qk+6J19P5Zs9cDupX/XfDc4vrTealZBJ13lnLYwFAr
9zCQPw/8Dhm3la7SJdwEJHEII0vXwH+24MTjYCv788R/gR0SbdmE7TrLhxdgS0au
ksvWaAgzPav0iKk5Jj7puAd9f/U85Hc2YE/tFj7NhGAhgFBjmJN9xpVwvvkdau+f
VMS4rD/2dFUSPo8x7FpgjtfpxlSfcCsF1YonD71uAOPifLKv4jWqUZXSZYqCatKX
o3WcBM5q1FHMbGU0eC87lHXM8YamZcb5GJKK7VBEP/NrzQ+Cnio/85OVosPhJUg5
pTqufbidcaDpNfvkHp0h3VS/KNzMNSOWUAubXiIaA4qoBHANioK1e3Csreu6NSQ8
UN21D7iGwoXJtR1u96LlEiNWnnm/huLO0sJ0E/82hxvhhqz+HmF1rEWv1toiHBkF
wkepQGbm+QRhq5jhkmZmPIm/A/mrFIPU6nDTEvYFSx8Oqets0R/Lf2Gp+r8WOEO3
nZqion4hWGCsuUMvI76iZ+8fIx7ldYtbXkJkWJZ54ca76RTRgOewzFwrEZYseUI8
HCgf3Q58+0Cxb1pmYR4yPqpugIR24Pb6nFFniFw248e9xhMimKFfkBLVEmP9tZI9
E+IrL4dxww8syyHyyeMKfKrx7YoNBkOa0HAhzkHQ1mi2jNEJrMTj+MNK6Dv2uDdn
MfKigPUnYK6P+dO6Z5teQhps+g4IZX1cEDc9XGvhUd6Gg7QpW6bFKFW+6rzjkHOU
ekPPDu5dsDdaTL4+Ot2ftQ0zxgclpdK6y4OrD4TTnsMTF6WB4AqHMS9EBUQoGT/6
FNpUO4dqY5aCpJseKs67XgMXGyXU2OOoXqA1mEdLsAIuIjufcucXGjzfJ0I5YIfR
Ot/VqwKGps/MuFBE4TcKfuBv4jOB7HTEBD616YBdhEwM/b+F0bgp3UnMImse0H5g
bequa683VfrMKaxqkzBJjQS7aqQSGqwPMpBopkXuC3A8XymnDfF2Oz2uAw2Cu8TA
FUhsbo3JuYJKfQ17pslW0GVhgiVE4BE0I5PIa/eu88wLbGgt0jwZSpWibiPH1U9x
QmcwQAwsPCiYeyllBNxcxXgTR9VGYmaUdvXGPl3e34xUkm/2/7wLv6OsprYW7tXb
330dAhNjOgd7L1iyqGwlQTip9jp70tgXUGpswrEXBroy67/8farVgaEcbkGY9RSQ
GUQE3nuDY7uB+zq5U2d7S5rFwMTTMVIhCjFdAHyLELC5pOUnq6UajUFVdF4UXSe4
DdqTd+AyNaZ/BSXaXhQst/VCYSXzDMfPoMaJFH5fqD11kzxPc/alskZVx1H7cAm9
med2QLbCMj6B+Y+57YqTSlnjw8HZXruft/XrHvOikoBVK+EM6BFyw2c7w178y1WP
k138xFSvPyEGNcxlFmHfWIfz9iy3LiBBR4y54xPmPFTSQylgypicDI9mtLlN2BsQ
w1Elt+KHL7fBb0jdty+3rLyzCmPO9cesE797VPtozRxJwwCeIoQqOfXdxhewUOBb
jxJ7gzJNJPoyRJWWikyWR7bLn0vlAULN52+LC2rqxovfTebdsMqp8iTTktLFfsI4
Y0MOGwOnZj1Y2iDv1JY/IBitD9RaJm2NODl/zJUADJC5itU3nQJ6yaFLZJhUVSqj
XncypP+fZrkHuvKA/nYFZtJaSGryNGv9owWeQ38Rqsg=
`protect END_PROTECTED
