`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pERzXkrhOefWYJbxEw0nwnePKeqrPDamIkScqpa27mVqeRm0eYx37OIu7cyy5XFg
tdcahO+U+RpZcUji+adieFdXjSLM84iYveDyRndLkRajdoeYP5wpUjQzJ8ErgYYi
m/B4FVacbxgQK+C2VgisIpKaE6U17JA59tP1UFee6ID4PIyat5oIhJRuFchA9qkb
XlJ8PJ7O/yR0/diyH/uXIyXiFF2bkmvh2leOxrEWA8WWgGphmlbS7dl4a4b9uaT0
uMYoWqKzbFJdJZ8yTVUrAkW+q7ToWFDlntXuFpQSjBS5xMtjOYuv6ygV6WnJaU2r
52GllZmrbgjmVwb/RlisWXb0Te3xIVXaDGq7twKfUFIdRHFzdNEUthuEg5EbAADw
OIjhAMcNwGwk5vMWLQxDWk5aoM2Vvu1cYutWJZWOjJStcqu3bRoPQdsmGSOSmvx+
HzqYdiPhl3ZBp4ANlD+mLSe9tvVyyuKPqmAS4oxWbIBGplc1fI6KfXXA/bgWe4R0
d+OK2bCykgouKFmdx69Cc+e54MnxL26KuBGYcgmDnWif897giltgQAR690yK7/XT
mhAMEp7IGaW2xoEBljn6gekFmWsMcXYQ8UD39pQ6CYkHpHXGHl1IeX6tBQkPne8e
J7qjyzrj9Xusugp1yTo2XAiknxmNyKaURVutqnx8lXx5i55hiiemPHT9uS0eiM20
E5UOZT0xN9Tu+m3lUwVNVAdPRiYMpfleL3bVge/O1icoVmXuso/ST1OdKjSHITI4
rFkwiYpzB7gaOhxvJPtCCC/ODf9obIMjLfgovPAIHAJ8X73DCCrXhULX/wntwNBI
IXEuBdgiwwCw8gblIIcmT557Hz0rZCMf11s7CYXYVgdDyRSXs9dt66yoeXgIbzmu
OsVkSk0t3gYDXneZ3X8uujQMhS1wj9iHlfzVvcOz5fx44LIFRiDsgKq3XgAz3nG+
cH2xPnektLYpmZkfw2qSt/XXtqFpFOTEFCgCYwpX31n4fQxLCl2s1za53/S9oWN5
glpE57A/YenpqZNOz9i3iQoUZHnn9yaF+k6fHoxzeTExyoNEz2hxjBf6Ti8Apao1
3lp88AsmYnpb9KRUk+qmldJqBubzFjefdIs6tYAbYemo6Tltv6B1dGZ0M/S7fGVX
Me5OWXdsQD4WK8XOWXn4m5jAn3OA83nT4B76M/EVlih4FE1yEIGiIwLQGOZo047X
JPfz3O4cxNaZESgbEz9/hq/lyiG7yinK3dsYbHCkbKPzAXlw+SHElq12SVugCuXi
oPnsEsP4xkJB9Z6zHQKNmZ9Q+XiP42UPW/BrPvhuBdp8HxEATia3glAQrQ5pPpAJ
kvnrInEp/tb+T4yJgvlDbhAz3pTGAgxfUBsL/YoQfu5MoG3hH6jCZdo9I/lQOJqi
vRwwVpGZJwD/zsfFr3/kDV8GIelMUUlrlg96tvKs1tAU4VJl21Mph1m9lajnD/bw
oZYGPivDCPwhW2uZgFGMnNYnd6ICkNspG1DkMHk3sW5xCVy1VbBzUJHTymSm46Bl
SoD20wgUGhux5W6DqFHCcc5yyt8RzB62AYNFUr9kYOfE4cJl462nFcHrXkJyN3qp
mSVNKcC1P9le/QrcbUFEHAMQX16dtN6w7+NRkJfb/YQ3kXbWt4uWwwXOFhi+kTM2
k/RtyHuDrFDmdSok/ZHEe2TbuY5Ojj7eSVmr6yvUCa2EGNqDdjgou9Gvw0QhQ4nW
/4lpdtp7FLJ2zii6oFVLyUFwZczB1wG0teivmTmSmAg/itlJvkIpm+bgwg82GJoy
CwAEzAJw+uvdJu6nYYASO9+jlZhBlqwuEHqBt2+Jo7D895a6+gYgbvZ/+wTlCBWw
ocebxqkJpaNQxEKOx54y5/KhzD8OqvH+9Ve5PIwu1aIBKNnb9qBwlER8zeGW+LFf
W9DnHz0iJZ5cDuLxgJzTtGo7JGzCEIsLfxcfNQcL+iXShYN6zVnVLjzD6zq81Q0R
+Ybpz2kVhu3nSjxXWkRSApAuXjr59TTupP0ZdibRar23gcvPmfW8+s97C9nZCz6F
crUhM5SDh8bxTQ1Z7vTt+qfDNThVNE1jbb5FnxVHwQKevgYaVnZLoTQV8IWXzZ/J
zk7fhCmVjnlKDgERm4vv7xSidieJWumPjq8YUKhqXP5ebE2oAeI8aTYxToUjT0wh
xWpYzmAbDOTT3OtZD6cM+HXMdXbUq7Fgc57r2a7bRvaIZrJS6PYMDLCe4NAUMja4
VRKXAt2Xf2hpc5do13/s6J8Bc2LHGbSvjdwxGkkTIXVH4nKvFXfUZ92DBgQ/T/AU
LuhhpwNl+fYb+BgH1ixItiuU7BlVBYrGEMEmRYCwri+qw3fI7ejyXk8WX8Kx01sf
SO4JbTGP+6Vahh0/9GLqFqBWGjfrtWF8kmiVGFJ+d52w3ZO6srYSH5hzfBDD+i3Q
b24KUeqfyC05xjX9w8gXTX94yljtJTDytNUxjRkW32md006ESnWMEvQAgO6qQl/7
2LIhRi7MHG2VLKrkzdw76TFbAQxm2THKRGx8gKmdnXmPK3gTdHI99oPmBWfgNRm/
FUrcysRV7bAKYj3FSqPpOhU2z7aKWpATglO561jfzMreNU0FX3oDmWak8gUnO+Kr
JOnfoKD6/7QGNr88arDcuFo5jFheKINiMLHWgcHau5y7xM94Emltrb4mQGiCquDH
UPPiousYYD073J3+v3l5r24CZKCXJFt8DUDcUMlDqtGJZzonrFsjYL3VSWOypTqq
Oc4/0YgqBr6uifHIxyw6VWpiTiPkFgCNm5ww5Pip4b+P+ImwcdghUH2tRxlWEZV9
GJTH2BXFjthnmHWDkxQZv2WvprKKPphuMJEnfnTgaweXNS2utFO8qy7di6/n0ndv
QXuBGQAtyexR+AbekaL94YhA4/FqGUcWRzSQe5HM6R3WxGq9dXjYp68sErSmQV6s
kQxoUjFwj36gQ9OObLJa2vEypsKH/ZbfGajHzIDdMvr18F1zvWxkAbSOgpSAsT9F
H4z/JbkEZX0ofZVzQaPKdoUpPaXOYpnVky/7/Dt8TAJlQakV9P3sP8i3vHkKOLL/
TNwYUcY6OYjd82gBzSQLkPgoOtfIPpAUAe7ZCuwWnCv1Vl812bOiA6li6OrEj101
YhpUWo2wG7sOhYOanuFHQWl7OwBcRvmK65HBbDJ8Q1MqbpPfdBUdXKzv8PwQekeX
lSER2GYwlTrNYYI28sWDDVic71lxUONQMhlHJqKIvfgYOvGG5jiGN4F17dAkaqqU
fhZts7TH1zdKQOGB3XFqqOPXxxyaOmLLCHOFBivFDgjaf31osWHVb7q9kvaJTB1z
lyUa3VWxEmdAya/yDSFRNwIUi4eoHa9NgRP/dlzm+NKi7hUfpFQXcdM2cooz7O42
N0gNGotLJzHEk/HwjVA4GAEAZIMucjmMzUWRA/nqtMIMAb1cJBn7RxeoEmfmSWDO
RHL8ow3T1+qJ8CMTSTFMu3P0xNqhmFFjPmPuFbcK84Xo/4JCMiuPsgeZhk1G9CBx
uE41c7Jk7IjoOmKNhPbWBt51EPXRAzQaj07sBT+/lLoAqh9T8myUs6OUau7kQjnx
hAQGqIoaxEkL0wKlZE59r6cHsHVmt3fozMAWWx+RVc3IJK9dxIfJACp7aPgK2m9b
Tk7ITNP35HsN4FxSSWhIW4fzmQOavKvbmsoFlCUvDJAWZQ9NFoh4lMUcI1uuzo8/
3t4g7tenDA/alXNgZ8UsnX0p6Bbutexyej+8ImuUFm5px+8J/zI1465ZJZZL1MnB
p4IKezAadbgeCuXFos7gCTpXulBBTIBlAqNf8p5WC/R8/UTFlCUrYnOVne/hNhPy
DQxpc1CuAJh0XPAvyRc2wdIctT9fukJjYm4jiE5x53CrQYp3b3K6+GhbzZSVqXC6
YP7JoKPyjKLOhkb8ynvKPvQm0FmUzdFaWNhFpS0mq9PJLbKYDJqSoElCgHtydSU5
bu3wNWR7JqT78tswunqCJA3omaY3DS+c2UoMUgKT9p/+ynU18VuIHk5L5rd6y56Q
V46VnJqZESTPW7s7CqoJqcsMQZuoBeSWmXgRAqmtvaY3dF6icanaWpnkwOeocUEH
6ymLuHezwqP0saAm+pCpaYX6vYFcYATcrZ5WncBADuh+fBj7aHhmlDjqV6X44YuW
84H/WRGwZLJsnT2vaNXV+ipWI+8tfmTwu4mQwOObfmyVQJ+asiky9pShD1SiGsai
ORPBgnRgDDqNG+abRRe476JV+XMVFjGhRjwzxMxERUYdD+pCBMBiHDwXEgZVEkeQ
XvRRI6eisATp1dTk6NqcMYqvUHvuRR70Asc3+vSIbIp+HTUSKW9X5pPmoyqhaykz
eZxSgYy+p2W8uPjaCX4ICSKefNn1Pm2AWvFGDybQ6CUaTYMP0MqY48GFlchgkWTZ
gYl9Um23rBOj54aypw8D+4QNZnpqq+rs13iTqBaU/3evy0HzlZyvQ3M9EnxXp+9E
80CLvhD2oEHmwlTY9OitELu26LZJnhlLu1M1Er7iElwXxiOogUvVzHIp/XLeHbal
iLrUNnG3/FfyHNP3fhEGJSKweOqTAwoZhoE5pFckFqF1EiNIn6xYDlZ0HH6GTs/7
jQOIDQ8SR343JPPU0zgT3fdXsRH07CqepjLSVp1Yf5lk2VAz5n3ZXEOuHapxDkEj
c59+WHtqzoKoUUZfvm4p3/MiMZC4p2/GUz9U8B5L49k9am3TEmRl0oDvYhxWEtjA
Thefa+82eIy1Fa3fcSvTX5cEKYi8v/QiAX0zIKMq9XpEj5VgwX2DSW3rgSD5C/vB
`protect END_PROTECTED
