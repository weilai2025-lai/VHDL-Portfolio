`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNYZ6Q0oiy8K+Y3Y3PSQAkrHjeQ4cy3+eY9paa6p88uLNnsCLbGEcE9oTD9vKtvu
8YLnQXtM7ZYUgQbJI3ab1EvSQs+ihU5QiRnPTEMFS6OhPqqcKh/lC40du1RO6Xdh
TXq3RmFy9Zler7PeKCiGxJKRB+EqagHZhWE/eMWezzYH2/qtZOOyfeykeM5nSIVF
a0aOxXH8YjgwfnHApOoZo1ah+SWywnEwCH5yvSczju9GFttmgqbZXHDwnlVswdQE
DnSE7itxEPMrgKVJ/JyzT+He7JD69e/SaqUMFuLqYvddCIwIBRrtf41FMpoDwWq1
wY8QaUf9dHGnSA9C9GbsNQbPluvSxg3VxlgC6KTvLWvtb+CjzrcVkh4eLVxzrZOi
ywS5JiJfIVvDBuRPIi371IUbT/60+oLYkIZDTvY9FxekZLPAPvHJyCYNGOqIwdi0
3JRDBv5uA/+6YGE/a9NosHo+3efkpO347A0N15q9GGUOCLeMVyMuIY2G3GS6m5gd
N5NtTsoh2Snw4IMT9TIrCINeNri+5vjN6F/g+6eBW8kmCBja/ZNt2pw7w9BETxvs
t+aecAiDqpFsHL9Gn4yil7y6MMNS7z5LGIEIJ/wwkspnRslqGl+WexIUmJvjSGGk
Qjn6og/oVmQpZmeVd17hw1nShUCkZsBO0gaso2joMju/FD2CLrKrFE0Eha5LLasJ
btBj7MOdAqBehhUp4Lf44M+31gtAWeQxQZmtPJ766WM=
`protect END_PROTECTED
