`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmNhArdfV26kqagln1lLBcq/Id8gaI8ZDOKxFIbSPHhTx4psb9dbQ3DZVYZ6JkQy
Z5H11YjcjIPlF367Rbdfhtw6EdKQFPu1QsrOR5HE91Of5JHEcWYlec6iI2tZyTxR
aHPFYkcZyQ2LUqnt/uvYvGXvMwXofJ7u29mR6/7d4dbcsctNrrpO2brWyeizK8W4
cgnTvFoiX7uVpQ3uf+8/0570bdQQqxQX9FsqklbA/SrYeHgskHRsriPUgtxJ+jqU
WUvUooOrlcV+cse6oz4UdSEUa6yBkPwf2H/0xFTmYbN98l0ztyqMA1z+QHkdM8n/
D0B65fJEeyZd060CRbe4AWQAmCxesaIDN3vKyxmxqg/Jyu/C4JOaF70tJAjYSY8Y
8uu4ECfvApbuKYYqR2kQ2whVOmGo1to8Krf3y22qxp1vAOE2kvY3xOlE8WhiQYsL
`protect END_PROTECTED
