`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFtB88wzdSx1sClJS5P5iSGujiYGeAds4w7TYCsstZpDRLUlDssG7igAKwp6xvkm
zf51QEORYrfhf+BZwFmCbDmhvGbgmCGeaQ2Pi4qbN77dvvyOFiVjkG60lGXRk9vr
DroU2R8Ofi6oS5XN3ZAMjbB1sHfdqwTIrmHDW2lfLBjnpBIklb9uaJD8C1P2tEB+
CtZp5d+mAFAMarPDY484W1QarZyQjoZYT0cHLwC6xnh0QzSF4hnh3bFKCMpdVi1A
A3GW1ItD9T8UA2VbLJ8MGjyS6kEySRqVREVcOarDNKkWEHzHvnMQth983IEn2r/E
OYGkJvr7azWSVbbADK9BtM0ApU9Vl4BHNDSGyI4FhlolMlaLxRKI6b3gVj4h2FCb
ZA/fghiQlzXCls+9HGRVdsfUa0bP3evZI7e2v883o5pJEfQb2QPnkkMTEDM3fK0r
xLKOduPMBG/xz4UuM8iYyfEAaUinRUgd8+bz6aC29i1HdUfCKArzRd/WED0T25eI
EEFb9erz1a3GeQ1F7l4p433GFUJUrgHfcimWY3JgyAVfWEpDKUFa3wb63hhtE6P5
r5U+fiCUxBs9n8toNlJdDhkrwP6rqBBxa5ZDF4Y7MrNWYyutX9NopV9UjG0U036s
R0n1iZytttd15q/zGmvHWlYEDl7YncV5Z/a8xkkhRLCQtApsB0tWzd1eQ3LyFlDH
VpSLM5xcfhU+/uTsFCLa7k46jGqZf8jLISZ+7WIHPqON3pfKBU4v+iaQj+mkeBJh
CZ/bCB1ZGqkmoGX82vuasQ==
`protect END_PROTECTED
