`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iid1abh4mCSAhpBp4iNVfBCEj1DsAScbPD/UA1ITNiuRY8iLtqsAhF4wichVHmul
Mdl9lCk4NuVtccMvCBozPZPrjRfuvYUMwe1FctMq9/w4c0QeEZLLbk+jaNBo0BI3
JqhPhyRTdlotupxfihzd6RJtBxuR9MHALfpHWloxyaIVSuarzo8rhZQlTLAwv8zo
jcrc8Ovy4kE3I9IIAduxmDWrVbljDbGLIaL4KVRwE3nbjgEKwR0JlArtGUO0FkpX
Rqk8sGQ3CEyWleM51sguDKG3YigFB3qDwhiqk+/cBifbeNJqH5ChMrrjrczoVtzg
X7SmCQqpNA4Ii+Wnu00/qVY2EhzLUNXfYKd6xJIroQDZrX5hFeB17OeRiXBTqp8P
1YALfEZzvKIIe15CsVjp4VRtFtBiMr5+8mjYxL++SwarB/PF9Y5eZsAXYfnlqdVX
8bSt+b6kGMTtxPAXKwPmecjKyetcVTeqst975hoNaVchpla+kCrG8vQYQFbgfMjJ
5ANEnh6M2bFDMLyqh0PSsi5rMlh3mBdPPUvLNoo06yM5AE/apdAqwjU63uIKeuW2
ctoYljSUeVgyYUmOJdi3iJ8GpDbLjpt9KV8rJNo/ayvFeFTxEIdi1C6c7ywz3vbD
jDb+jp2j6nPoaLtc5ju3eiu+/sIJC4a6if7XhM2GCT2b/P+/si44gMu+NnfQ369T
Vef0TX23bwySSpMne4qEOKgmIEyudFc5eAi7fJAYpgTgfCZUHiYCola7NzA0+qbf
x5VbWBnpqcc7bHuEdxLyLZAXEI0ggms1ieqMRNM8erBOvQgzxCLYaU5gQu6wHAG2
iHeK6O5mHkHtcijTN1nJ5Zkd/m+v3dZSx5K6MoH4Hca0i8PPgLa1cBoMGjcfJ5kN
NnGMmkQkkMsaCmAkNskWiYI2BRBGNB3veb4/vC7N7cLiGQ0ufYaOPqwVUJTRPofW
JYn8grBKiP1Wx8WR4qx7ugpCRYqcUigJ+PSMNiPr0Uv5Prcd7zd9BbsThYjAfzSF
0aazBV/O25llDY2gqidhNp4YRUt1JBab+3v0D2SHndqHmRngLAhtCVpvyFduBl0z
SqSZgvya3YAP4JP3aQlNy3sGuWmISvC+uUv8gdsPtEtfEbrVOcCBDlN4XD3Mwc0R
leGY78SYsIPcb1NL5Yfe0NdvpHZDaFAY/ukqEUK0TqzeIQfMjAW6RdG3VmQyg6ey
IwhAFNQLmCWeV/SmciL1a/MvPbMO9Ab4rwTqnSgtcZAF+qAvVvAggqgJ1Z/nb3Hc
XIS7DhpcJWY6WsfYLiw1NPMwpiMVj9KPjkjGwdcvXVLBNMYBdOMZ2ONiHuKAxzru
xeHXfPdYgBfFMf3hjEilvH997VPhWK4ejcasvnCwYrCgz0soQuVKB5598E+sfjLD
mG1RQRJQy1MwJvf+y+RoAAhdYRVf73KU7u5A/3cRqqHKJQ5ugdfxZm2xAbyW6ctH
w/VD3XnyLd1Ig8wl9NhqjrwVxmDy/Egd+B2jPH58NlQlMChPDwZcfj0zwiJnJIvC
Qqe/Ade9Vhis+eVLtkG3ARhRx09/MGhsvh+TZU254vlWfDyofJZfH+g6+JYmfNgt
zzcv83iws7QuvGir5MrpSjFefiSacnGyfgFaKOOHUgk=
`protect END_PROTECTED
