`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzb/o1to0ww7ljsL/t18f3T2268QmSagf0WB646MBncz7aWCQpceA43Bqacy9b0Q
IbvYNNkPUiRgshC5yN6DB+Ie0qXZJAwMiiwZGGVv9ZKHLevf8MHh6gvAz2MuX83L
xl8XdHilN7hM86pG7vKltZa05aZ1tDXa/QxZS4UYBNdWx4mPqMovHCDYkrsQKgjm
tKQyKFxcmDEnPvtSZZboQkh3b9huDbQnyqRqmYdmCIFeKLnaXv1WyQd1FrTQAb1E
lUKi8dOK0y9lf99Bgze4LLYWrdQqvyaTPKB9ueunXGaH78K73xhxV2kk8wSv7hRr
ECqOjw5YplLsGriKnM8VT3j6hhZmlfdl2BJBszvdXFkxuCljgpkZm5C9WWvCUkML
Xz962ANZ3JHh9ALMtfD7GhhIhTY14uAE+nDJsuVYs/H8Jfb9Su+nPAKL2cHUNnGS
GbLdp7AKtBNtwaJA4R5pjvljxnICQYCHG2jr0PKDHTfh4AE2XpjYvL7XyU2RIThF
ra2DbOZJkqksFH6zPG6G6NH1FIppkZm9DVMGrrckD7u6VcSQjAnzUTIARTtr3fDF
jRDxad002mBQjH55yDhjtWRpA71xkNjjkZOj4dMPHceOWcGCzU1xCJwJXC5pxayW
efFjpZpLdQ0gFhtJnfZH7vaXOXcUbzXWCl8hlEAn6oUY0BD40OOYvhHQkW2zaA7P
xg7e1YddOR7QGwA4w9I0xjbAUrrMEyBjMjMd6ApQVN18mVEgGNxjt2Msm9j4NuZZ
bsKESstLFWIiOMF8SBYr72IH05K1JXzykNA4/2CSaAdaNWEpZQNeaEO79N31lADx
Re9z39TDJzxrUKBM4MceNTqAStqs8V6cTOZIiZoUxgiujF70GDa/4OfTCTObkBdS
vwPxrTH6FCd/zJzcbQ8Kttc3DTT3DKQYu0gsZq1E29p2yI8kMSSzsC/xlftcUQV9
j3+QqpBWXmlO5sjU1AJRQuSTZgH0ktjIryM0Gd4NTRprYzGfDkmnGTln7uq7wJn1
YwA7jEdD9AR7K3fSQZsgQKemZZLugQErxmyiAQt9kT3x+utfdmRqmQWY4bDHgPm5
ZQ6Rd3HwX/A2AE2UmjUQTQbAyfVLw1o2e5VOBdr3hG82s24VzZaPLlnooPlzpeAf
DmChaW3eXypZ5aKHoQe+/TKXturZ2sM7VPu9HcCQECxEXwL8n1bPHouBFb5V/1GH
mKdV7mSc2tNJozKdRG7ReHdqbJko1dpOCOSbm1kotNYSoDe01GfRsvHT9x40hSOi
NV3RBz9abLgyWYqnmvlejXe3v65hZVT+Jd98s5rXEE0Z/HsRgGz4UbqA6AEI//26
uC++thXayzvO8nJNZYn0EDF6ibspTfLu+F4bJytupskhD6+Va6Z65cLzu58UEZ0c
USIfz86KhvLWfvh8H3qzyiYvMvfhivNSPNt+r+pgg087GmdPYnmfrzb2mJEpEAFg
zmktlz57nismkPV7mqkczEg4zowwIbkrePfQIAOkk45YsrCefDX6WzTQ7SohEhrf
Lluz6CZjdIpHz5aKnWzwm0h3hAB7KMmTm8xnmPHLMEaUujMldgFwZEL4DYoygxBg
SW95BmyW6ZiRqGAuzgqmZ+wSdw4eZjPMxF8k8oEbzbXVfrAQm4Pkt20rQUGqsiHR
nb3F0v5gElS1kywJqDxiKqwBhHeCD7MTFuzmmseZ52znSKAVyp94SzWL1nXSgr3+
b3KIC5aqkr0G/nH/Dc9nJNEp5ydArnnbvY7yxSth0knf4VXeHEU1752Cu9NzD54T
XWrxm104zB5+XSfENvCyjCBWBx8hG9BLotYNay7FlewCI2uUBF+0OlCc4qohei5R
VfYk9AfQW40kGlYIiz3EGi5j7/CG9+k0eDfWgZOc7IHF3RDz5SeLtIJJ7eqGuP5n
GY4rPl2hprFXObUr0rRWqTLHkQ9rkKeR+4yWNJW5Buu7WM8gnb4FNTI/fuLyTpBe
1YXHOkbRfueVCQng4mbl3UGjZd5CgUFSGCbox0x4DXSkP8vskV9xaAY+RJX4IwQb
R9tR5im+Qr9ZI6Va+hO8OM3K8NfHWmiSeigaduVTEbV/j8WF75BFtTATWgcX6qXQ
uLDZuWiKQa0Te6erflQT/3R8Nq32lAllp+X+DaqFBLE5WIvETxI/3cB2G1DmRl1/
qJRWkmpxWqQX170KUAsho9QMGFXiuwNJWdFHProFWts4lbA8tfq38zBgAK6JV4+/
I3S6p/8D4Kq+6ABOObVQdQVeLa6E+nQwUtpAXsC6BjdqmmmxmiW3pPIGsby7iTWA
HgY4uz7zKK0pDwD1IzE5GRnGafKtg3I6CpSRVcOYX3bPDY2ouCTGYlrvwGuVCa1K
jaTcTampmVWiY/pdqPLW6Dsw1fTy6/C2ONd8/0lgcR0zbIOptvPlo2m48w8oUV0l
90hpi6jqT8LUD9RBzhlazFfNpiqMXtHcRqLoU53V3lW8S5xsUSf6HDslZQYgDhei
Y5cmgvpFBiM00ZA4+sgjNseRywiwn9Pd2VEyD+fH999w5NWa7UQZPpMXkLrKMnoj
WNhyAKQdbcgVUQethw1tnKBx2JHF5tc8cGKjaMi4Dkboqnxpusanv6vE1tb7xNoA
kpUVXdDKEWubkUSYrJjSsv9deQ2A/P1rzxBItTrRJmtXIcVuVsU2HOBguN4Xzgjx
F4D0Xos7HGGRQqRU3zVe7vqFxZxyC2hX+7rnBheKQ5l9L+n0TLbRS9XW7W5WF7jW
4cAcdYUWZP6hVl3jaAQHBil5UrYyyzTPTjW+A3L/v49AdOqzsPmyyq2AWbos4SwF
P7eaIiUEsu5AxCgFhl3MX5hHDt8B9VQ3BzXvupNfXG1VUwRVDn9WsRoOBNNj9saW
ysNz+N+SKdBsBVLHdPv29APks9sidWCptnaDVX1x7xR2TeiMJAyagtOtc8kCrFkJ
RW4k7BDFcbznptk+jkZpnppvTaQudD9hYct1n8dCsKGqgHIQCz2S/MZQpJTDXZuW
RTtO+2nVkmzlsvYShgsfEBjivp/xWXLEJZi0nqhUico0X4MzNCAWiY0bKdpDIq8j
RxdpFU+Nf5ZiN7rvzaq22qpxdZLIv4nfNsjj4ZOlLPaCQ2jm3yH8RvgVW5NxEYyV
l8q5Yj079LjUR1KCfuGPll5i122vI5Rr0bHCXwo7mczwmOFIfLp96jrDwGJYNO/j
tZGmd2yHckRkgtTi16sf7uLivEdZIwkv3Kx9nn0zHbTuGLw3offumf+cJopcNRaK
6oqBW26Ay4ROAzL6eXbZUdJgl04oXDejLMmtUR2F4V5AkP2zB5J+jFhZY5qZlhlx
hvKmg8gzLLxJlZaLYA8hcy2Y6Gy626pMx5TcCG3xDERrH/ZFyuwvKHrjRA8U80NO
YZZL3Q5sgr0l0lTK8jFfaTT5pGeriEdYnL8j3xwkirrXJmsjfG83ZHj7NdpkY39S
6BZO1GDXI66GoUPrVfnhnmimfkqQvtHBI5xl/tFRuFVwjGOb2KZ96mpwEIU4z5Vd
WZhobV+51eWBVmKCStiNAROeZGAW2LKCfdba05rVtXE+jb1RsDYJd5ne1ofbH5EV
ilmUYk1fj5zJwnOFOb+AN/qoYCDF8cCZ6yTRXOhOAaUrxlFzn9Ba0zoTUjGEjSXc
RZTpl9gPGTnzrnhkpX2hFrgP4uQgjkDooFKked7jvJSwbVonFXPVCqe4n5E85ctF
usufIRLJJB/QQ43Uprkfhg==
`protect END_PROTECTED
