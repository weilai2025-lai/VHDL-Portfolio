`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcMCrjku3qyYxygLlctzQjXT1hex5pUbWoD02raRnq1VXS6KUV/HBrB0lNYWvzry
uBQD9N/TCjI0tDhBVLsmofNfJiPF/YBITFW+f5dkz3uz7ukF+IAucCBQiMhxA2vn
OBDtr3S44AZxbaa9viV1JVkpAb4rfYXA2NLinuTMLtqFLdIYVxjCJASveZKPrcnR
Ez/ksjvuuMfmT2W+E2dbO+t+8OcIPKSMKEpRtxJjC8i3UsH1xzQJJZZepa+61gvI
4ew6vpupf1zGKwVXsy4O2E4BluwDDP6e7ZnyIvPd/P85Pg1VNJ642XVYD8VQr5cK
HqPraa+gTbW2CygGDMDw3FHu1sVK32JUlSymEw42o0Og5GVaD8Lxxfy28awOrVn1
3OyeHTbou7UasCryO9bgEJ++dT4rXIIFShPTvoT6hx0wBAh4jUdTOH8namPpMMH4
g/iEa2gh/Ji4PnoHzmJfHWbqWP5pmWQ/ma4F4ptS523b9P7PHcRaawzSfaUGVeeL
L87CcObKBUeyoluD3nyPiU7Gf1xd1GojoUm7QEwrskH8RbINiHs6bMopjO36+ujt
Fz5XjLVXfHLAXXJZT9e96XQ8+5eJ6HBauqSWjf6YnuApLU/QKAlEeIFvIAikePki
5mpFom/xkPyf1lKDE7qckmVJWbNUwDbVUIYkf8+763EitIcOyZX2BX6FoLvFaV+z
hgh59TAt4ILwxeqrAhYm79H1+L/HjmcAbLCOFb2iUMOTiJTWeNvN2Gf+GEiW6/Xd
prlQ+zdBg2NJJ+3Wy7hLtzmaAEjtgyqno+2UU/U2GTDqmp22AAjmNt+PDJ/GRFpR
l0WUeMKXbg5mvvpQoKfdY2tiDEf5QakpcezrZsAaJ2K+jQkjaVduQV1nhFIBf6TM
VDPEKdsxr51UVlqUnZhRi+fWJX817YSchb67ns4l0UYj8EeDQYhqWuDiQfn/1GmU
fxU6Kg9WyK7VGZnMyLAp0+JDe2YTZOyvb6jOM+SR02hqYgRT37IyccobiuPyKpPa
xH4vKDATAiZPJAaX4cDLVO1jOTNxxQeEDSK6K3xSi2RqXlqDk0tPEBGZpJQ9YzAv
LxC1RMcIByH2qLV+lnjl16pix5+ojnpn2iYyIk6WXTvPkYwcSyWm/RvdnwjOV4MH
k2cpuyZnLr3JyBZr3YarHsSkg/sN/966uLSbj1Aj3hHx91PdzpPtxQJZ+0LPRjQB
GTF9aHAbA6V1XwQIfi0UbiDZ+8rjtq+S/YI8qDgQ1u4btvPV/9MbDpttNRkwzVW7
ToQkGHr24qmUJPFYKFPpWdvYjMxB+yC/pQG7SfuBtt3f0VRDHmNYp3FQAqG0kTMW
9WczMFlHAS5lNzROCNUY5im3aMSi735geKAMnzoRSPnJ0uHYBYsCPIUaLUpSHU+n
0n+ybHrlUmBS4J29limoexQ3BbYNJiZ5YxMUE9uiLT38ZsJYga23C/zri34cHsAR
piC/X0ZWsIg3ke+5FIOK7MR3XZip+SOWLJQVLEIxtdDQOdP37cB1dqDC332lgBGV
tngxlQd4FimHVue54h9rSK3oD6NgmTXk4Qmi9jUNPw4BgRevuS//IM0MbRP7B0do
4U7ijMTMikTEglanNnFvdp7RBLEDeSsp+4ctUSneEXPIfMHi50cykK/nPQdGKasI
Sj8fndoFGzUOm/RlIX8B3TMVr/rzzT++PbBcIfW60ig/Sq7QfHNvCdqyJBa0TZdX
/gmO9925bF09nxSjgPPIpVcQ6iOpZDxm9RyEGFjHEjBL1bUlZ6y3kau6zRDT2HuD
Og6ranPB8++L0AM3XUxWDMZwkzy5UJLhbeWxeNdYx8bsKLR/lYge+v36OF/fn43I
XvjpUgBhwetn8veTNs8saEmIpy066znoIgw65S84NcN5/orDMMbPelNN9wS+S/Ku
Gr0MeU4WCEhCXgW6H/AdEpgBwlfXUX6x8JZbri2TMjxNc0mqOKU3yrLiPWUddqCb
7fT/XeMjctJsJiYMXHYXWn9jlTfw5TdMQuew0fvLuWsaaMu0VdO0LIfMzPq9Ezjv
3bAE8zwgeiYquL+MMX/IqTkR+Lvuu3RLke95UcZA8M4lxgO4n7DbT2E8db8YxaPw
j0NApCS7S8Bcsy8fWmU3ROnA7Y/MoKhau+S1NyQ3kPW9jigq788/o2fndrER0HuM
uOigt64Mr8wna/ybslYkXkEk8Uk2tpBQ0LRqGZUEDGhfVmDEAa24Rc/Jomp8oWbe
rYXYCepCSGzbcPKvyL1Jb4BfDoAPwwZwcLAG7yNr2RjUPc0W1WsqTBaIA+mSkeTO
A9YQmWm09+EKNObCahpGKKkZ4zkseASZhmwq4MQNDUsJOTMjN7KyQAV0Vg7lMdHJ
CVQtPGAqE3VVHR3y2G4mQK8a013V85rIM0o/SPCm66Y0N1xmA451XLXFsdPiv+dC
JfwoUzL/6VHnOWD1omS0pjVFjNcozp1zf1ePlDIkPS48pOjEd2ZhU6ZHT03DwLD8
XToozkBZhRg+0m+s7BsZsPYrSbNj2R+GYrbL0T39HHfyhipmydol2rzklxo69kD5
+3JJsORzZJJuKq0N/gS1KNMq9e1GWj/32qczuxEWh+0t52N4KMDZyvxauYEFuyVu
NcBoS5rgPKgeWthddmYFzl7AR51bI+zW8Lhqj9gdUbq8JAD4zzDve59I++rEJ6CL
6cnxdsIKwfvAVcC5LoESafAOSZsKd2izdd7ZF/lpjuIOHkYI8vsq4u3nZh+fBAwH
U+OvSuDz8ksXuejztdHzVUDAyqTZ2q0Nda3msT+8BI0f16cwrRQ/7zbxUlI3A6I0
/EhlyjXL3xBIfKo1T5R1TP+0kF1O2anQk6F08EOP4YJMdqUF28JMrZ/sbB3+UQuZ
gFu18k1zGjEjboyAYaE8LZoICWhFTT9fFT6O/b2uyVr4kudScQrmbvXFPscazmnR
W2UhUWS5lggPg3rKScWccksWKmTcR2B0wxZ7VUi8EE3GMgNhbVYdJk55XYof7zZ1
cgucQZn1OHs1iO5MaaDr25eADuDXxnmep1++aZcxqJJxKiK5600mXF2P2ba8rV3+
HspddRmncOg6UuLoPK2bv3C1F7M/Sdzwn0YMHzNYTk+6Qd2x9Hf8gMCsbKqq6Ka6
DzhdzdD1/4NP4E5P2+/1qJmC20otN4FKQWEap1YMQ9fxioJ985JxTCGWYRf/JHKQ
YYDHRp7PsLv7mg7bCWHRO0FhRnRK/v/YZ0VUd846MemB7Eifj/FHi/iL5RankdgY
snxM65ByNY43c6mUo57j/r3Ml/D2azQC5/iAlXEYCK60s6xTPpBEbWu+OQNwlyQF
luBulC0RGwh004Ov0f0FaauJLB9kWmjjO6rd0hxSFGx7hkfEujD570okDyhGd1MG
+VWR7Nb4RH+q0onkudyT4Y6LbNveo36E0nqXkm1ppGjNzaCakJxUHCov/0DCWhj3
/4NtfFDklip+Z3gMZ5emFDXhbbA4gFGz5O+OUtk/bWA1d83qdsxPz4iOlQdaS1Ap
NEumNyBun0/4DE32PB4oNqv0SQw2pa13msaTmbRjsD6bl3t5w31WrC6LZvVw1cVc
gc16IYg6zjHCHdCAGm2tmOBLklEpGCvxhMGNz9CcSfQJHfves1l+EigwpHQgBjb1
BL/i9i9kQwOkiwYIt96qE/zLlHsw/rSnYnFjMNjQpDLLhLUQdlcZyiTP6bqdmisF
537RhD4iQK0Gaa3RQJCHDl0P6PyJivQh8IUo9BpbWXfd7Ap9TJ/J7wgQ5cmKfe2t
mjEzMmIIu9onLxLDHXauv43G2Gcsystqv/Vn2kzcZv3jm5BVrMjMddZoqeVbKlBM
lIyY0Hrm0wpetFXMnLC4cdiRkRf71EBaJmqK4kBdpM46gb/gdlo5qkuYiysSOuLw
lgwYYNLDaIuC0Q60087552mf0CnuTvpLCChwv6psJB1yhEd2Sgtu7rUb3nex1I53
VB+uAd+nedw0m5wFi60J1/NFgB1QRTJMyFPtXNbxCFeY9qrtx4udD9M4+xtrxnb/
qN33NfBy7Z/Y4R+XT7eb1qpa5EV0UGTVzwvlu68a95XRE96fMxde78ezws1vTYDQ
YbY4GDAKj0MhlJtosb2Mab3rRhY1y7p6eGkWgYfI4Jfe9Z0lemOMGHQWt0ILmcdl
eGZ58pqlbCfJJocejccahSaFrsDlZCrtfT6ALO9Ke40wYrc2wXkx7PaycP+ta57Z
6NMK/nm1Wdxshu4XsgKf/VJl37AdXevO9qVH4kiDmOnfspI5d4ACEEtZf0woFCYd
xFlnV/oxreMiTUxt2KIvK3S/SA4FxFhJRH/SZ9HGeMDQ84UBIq1+wBevYMGeOfPU
TV8ODPkvlTWyanQn4NaMlBa4JgoZXUQdabnHl90R0WK2FqltQOxDTLDZs7BQEyjR
NUoeeTvaUFped675uFxwrElO8Wu8704nKXVJszODIrbrEgF7hfcVKNq6ytKjF6ka
UrIhfufpz+RbKnuuIndTw1feWTMoVW1UllbXQnde26fzaXeSyNFohAtv/39xoaWe
o9mirNgIVvgw7aSTb5GS1d+ObZEV/J815XoSBAlIIOizoTmTloF7Q7gxctuuqSmY
8KRmfvPMfDKng70sg1C/pgwe9BFuwCrjdHV9lZBMAru/OxBV3fQQbGpm08mVrtmc
4aB3An2L3RLsJhJbwGI07konkMiLl8DejB8C4Qmct0Gd9CpGuqr1rf8okR5TkX6Q
S/zu+jqsA8HEsX4P1IV7X2Xr1SNVc+2nQJ/lvrkFRo2lnHp2SKq+Dm/cTGA0+ILA
rfadQK1Dh0E2/wI6Izs6zAZzuyuvNhtTAyURyisroqZugT9HI3DRPcf0Ere94bNX
NkGqX/+oC2jWXYEu40Lc7X6FzSPM0xw2ZEMW9spIejMj4O5qzA5fMHktEi9PH0mA
flXIqogQCpbfhv2QF09NkNpa5jI3dspW0sfoCqzjEJ8dJufuG7GO8XJjgrGpSryv
2xCx62Mg9dA9PBuMVnf/FWYtFk/6xaUFmmdXJ+JJap4alSFaZ+VsSvBG99EYXOZB
y5yhNIkHkGMgGH2cCGxuqajMbQ6/QogSu5yIKMtdufN/1ClZx2H7D2t3ArVTq2yB
xixwA81FBt/Gi4rKSBRGjOR9Nkq2A5q68If5KtbYfR+b4/NGuDnj2gb9KpN9GD5x
VzPaRu5t2vsBbZuZ1fZYWAZ0ZfS29U4wjsK9jO/ecw+KR/n2fgh+AsrRv9pjFnlI
5GjgGOabAd3nhZH1+PBiPT0tRh42+eXkAT0X+brYFD8A60lO7D+kFfnqpw5Uc/Tm
f60v5tIWTygN5jl4PjcU3P+rabceapqbDvaB38B8fi9rnH4Egm1XgEm7no8MI0kF
g151Otfnc1Tb2mOoZx9DbnDb6w14VvchuWYldZIUcyK8ihNmGJChLczqK5yH6TIL
fgsTMf+TFW03MiADeLpEAIiOzPmQt0hPbmPr3SV18SL0+OxFQlQpDodE6qlfgC0a
Njuy460W3Ua2MCs00L2xmSHs4RB9iwNCTWF7kfJDhVEOUCFnvYoVxPA+aVErnQc+
hvEPdZytMDCN5mRv+9UXnIFGlzT+yDyUhcxVf5xiW3TV2cHLCTmQNHg4gS5jrfVI
kXGSYO467Wy9R7um3FP2Qr2Tv8+CE3NX36EOlcDIy43Qoc+LwDb+iRMYqfhQAKVR
IIHBGpIcLVN98bHTo2zJmOFsQkl7LKmbPtc1LdEax954Zu2JtFXc3IroEJHqaz3X
uGwa4iU23riaEO/QGS9SG6S2GAuI9XK2PsbsDJyYKZP0BOhdaUqnqZJCP0YUqMbB
eRqi9xDh5S6p+4r4S27Qbrthqv2x4h8UGI6LXZzkxy5IlKRzwnSwz7qxyeFBVnrv
LhTjB5wUbLUi0jqND+SjZFvIisDF0N6zFida8ltjjVs06ehsh1jC8/BhlyeZOw1c
AQPnRZ5u3LJRZvGB5da62V2KDL1yMDxoLtHwt8A9oEEnvhtfCwgokTS+h8bQ4xif
Eqb/EjZHbLx4QDE2pgLp7wMs+7lVka7RsnDsWGTjmT1LEeiFiD5ll8/+TaSyqipV
SX+G7IEwNLL7dCOy2gzOdRBBEPgUSXT4Ipxv/tNuL6E3+UaV8TQmDf2RSKXCUc7c
AZI7H/iMHjV/tz+5NCiWrQz330TjjhFU0oSif4FNYuha6h6XmB/S5dW5nDhYzL15
VRWFxWHop9zTtIYAKYHSW3r31ZODutZVQ8PC9oXDaOakZbisGZIePgSX03j2LSyr
RdEeLfIWlHKW+4iwkpHr7UyZL1Uk8F01WSi1pvuhJRhnMTtPjoZ5hs1aOQ9HU8DX
Y6WZQawdDy4l/OMtcwweriLEN9l/aQNXPbN9OWdfCbztDkWpVxh38o9DD1L++7yK
L8BBJpH/dv+xrDKbppz7WnX+q2h8ASt6O8TJJOKaSVma7EnwWK+WbpIyUgZQlZ8+
86+O48I6Ct4OZjLdwGv1KgVheJBx5vly/clsapusfpIy6NpFTVEIX2MUaLNg3Dwq
RR2yVVOL7002tbvAVLKyAXD4xtV6wr0GE6ZoFG98bRWisM+4IufCq9B+EP3ei/7K
vWYuEEWU9gT3kJ2hqlCnxOP2gNI3bK4FFY3tZsCiq2Ynz5rjiJEq80xuMd4di049
GlOL3XQL5dcbn6/NgAgJvffx9ufIyq/g5x5skzaanEnwepFrDzjfevadCQCHIm55
NAJqilnEi67V5tehWjTL+FKrDK40DdUBKSSrQxkMmzlkGmwUH5/6UIfx00pxYXm6
Vl3uR/5Tu4jxbg0wMEqr24+zM26hiOThLlGBT0c3sD+PEXUQLN/Dr0bcMuKATztD
3qQj9sEFlBU92y1Y6uGtTefKW8c57sZEockBmeHoQ8ACVmx6xoCLCs7j4ojrTRz1
NW9LVvehIwt18QiXobdZNgc4xhIuy0qMJacHZQglKh+sNd1/fo3KoG/0A4lx7Iqf
UlDGEHtjTo8lnjgvBZygV0ksUvixbIBl42Yx7kbsb765dXsMgddVj8ReNb3u/GSJ
JWoDY9MMM1CBJdxgzDz5S1kpxG/FIXWyRKO6novvpj7LrQoOeXigvOpsbMJnfZ88
oNDKVS5Jcwl70qTNNFJ/hqaFpGMovyYTa+Y/I/+5R/MCxOOUtMGp2aKhzUHBWxnE
CV5hh/d2GnCk1uTxhHDceFLCi8vVJaLd75MVIcnjycFbs+uC24Nydidz6EoPpage
f+8TzEs0yVgn4gbFJSqrqmEmZoy6+F8qu34sPw3CkyeTRN73VHLi+GnYjUy16GFr
kYHPql8aYkeijHhE9zxBuLTNUkLbWDQgBUap96MlIyzSfMJksxEj4E6fjX/ON5pu
ditPdzbKADJBE8TrtQRLPuO9NFQBjpkvp4s3UBOmmCRmi+uQ9m+MEXCfvpQCc87G
kQFdyzQpyvBIrR4+Yfw3gOqdqNNzuROa/h4TxzBo2ePlRtT55ayBiRttJre/vwCy
E1hIotAk/krCHumtkQIL3GwKK5OYAqDG5x5BzxOJ1LaSmPV81fAKMQZ9NAwg/LtL
7u66aBQ6tWvMNIUW3yKjO0V8Oq7S1Bzcjf81SDZWo1WS+Po7dee+FmWIxoEBJhK1
B+pEj4yV/AQjDHUvU5Kja2jGAGlZi5hjqwrvNkiWijZK1ZkU3/bpklVV/lwWbPMZ
34OkHgY9NrXRrU2uljpvJRR0sv5lzmJASizo6G3kZYJFLNIHs90WqydrXvKMowbG
AQqiSEYAelOpDGtcoTYQ8v77HJLIqvBFoWUV9H2vMFTOi+LJLP96IXK03oQkpnlh
nKwVigN7A+Jr3A6+/my/7WjbhiW/+zmwCAC31YxOiugT1gX39fCGtpUTSmlCXsm4
deaYdUmQ26EjCt8mqwGDaBHUhdhPIkSQq+5LfDemU+gacyksilbGjZv5PuH3WK6N
Cia0ax/GaclSbw4FvDDmIogqo1SrK0f85wJ8R0ucQut9Er7RROlCWaiZZDy4rG4G
SMlHV6hfreL+2ZnY6g7lTmCPngRZeEiB3rTfkotMgniEPZhFD2tfQmAkCm7hsjyq
EsG/RHVHH0/rEevQkqENHsTy+VgqRSI8p4WPP+7Y4LY/gcugO2Nqv92OF+CUOpD/
xr+d5ry6TwETPBBEmR/oaPNv4gDX1MQ71e2g8HX7ccnGO/q9KFJh+8IKOsQm/1sr
Zv4ijE+B88plh3o18MQ41Izi723vB32dUM9yoNnvMg2o1+F+106OH8NUVOCJq6E5
FFZw7ltlBxqGhogXAZ/sttN7ZFNFniwSze1cxIvBaO/ToUFcQXnohdgdmLhW58JP
QXTKiI39KhYeL7zdL5FUKcAXKqy5v+KWuvMllPwKy/6dx/cxppeDy3vnH+XxsJvq
gdpNvy/9/n8y+Ve3GQgsjsN++UNfO1QvNGPX00ps7vWZF5g5qq81Y6brpjjkNJHc
fXDSmQAs+NAqpMKigZgIhw49vvHo1GzW15l2sU1ukGfbN3h4W9pGFI9ctCI9R1hy
68014HU/jBAqKPeoThszOOl98tUkZnL+MhJKtgtmK6eVd6ArloaJg2VEJPAyudxA
PbUqc0+AiQVLJA9sD8yhBkqvtmMHG1AotsWYpRZVAFkRu9Ww+TWwKbyJWuxvK+S8
SLfI/bnEM5UKlC+7ypFH4jjeAyw2iWwF3xC+BPHTCPrAQ6tQNJFoEfsCqQjmatqz
jNXezfxYRcM4F+AVW4/MYE2UmMD8a8pR6MG+1OMrAcLOu2+OED6cC40Xw2LhpA4E
UqL3i+vNv3GIY+c6Zhf+cOeiwSkbe80DfC2lDChxBNl9tWqiwnQZ0xO0Q/cgZubE
1y8gy2sh/wNMm279MIepdDPnCIzKbgYg2K1P8XUIrlRQMwMciXqaH5i7QUpnhtRb
Jce5mPEpuGDglCI/tCsS13dPqlw3EyY87ibrr8s3TqmUw/dLq3oZI4wJernDPQjG
KW2ioJJHzPM9BLWbXdy0Z3D2OKC8eBVqsz9PL1VEbzsKMFnj7p5kLADD7IGbWEEX
RnI8oY1ZXFbj/mPp4Stb1SqLgt54ztJ0k6WbN3mA3e8bY1zTX5Az1U0ahkgWzp1X
V6RKnhLrHqeas1K+un3HIj0pD3t79ohah06cjsNsBW+R2MP8tsAs+gJactY+Yz3r
uTsx0LXcP7hlzfK/GgVL39S06bOOfC4nPJE6z3CTThqVwCW+Ch7veG1K3ivtatrY
37q3EaMWse16g7VZwNlCcI5PRrA+CJQIDPQyQ8qzeiYaven+ZHHz/mgYX/UbJTch
9BIe1L2VQT8Yxzjo1KoIGIHyS/7CNqFtBsIzsUB8VKS7QvsBagree8agMnunuDb/
A19Sy5tkSb5Ll7o+7UcLU4fnfPrGApiIc/ogO0+ebwp2MR+nGhm4aElnz+pJjWVz
Tamd0BPg61aqvVVhTCxyPE0HAPkOBYb7mToo+/bcuV/vX6QCAMvfFOYZSOYXGkq2
6UFKStxgnBpjGfIOcj8XX1pbksPU1IElBNBwMG7WBxWKEt19tgYzqSIIGyXIw38q
qsHp3ERFjBzoIT9llKFghPdJ02unDsWPdlRfPbEsice3UWHTaXbXJF95PJ+kzDAR
nlao9UAQsUSn2Uw0vHRU2gBO7LC3BRf6ao6A/WorfT861RN4SWz6jiLZyEdhBJh4
5BvX8fYOoSuttsEn+Q2ixbowWWjbYSUz+ZtdRo/lkyfsIJLmzOJK3CYvNw5kUqgo
lWcY3xVG64k/YUgV8t6Y0z4DQiRIl/frSpAqo3quHpGlsWjvTdfolm5GN8ACA9Jn
2ipOEP2VEUtAC9d0hRDRY2/lCwabPKKHOzGYj2kW09wtDVbUp137jeQ1iqJqLaWI
L4UkDeltth7ZFNvHNiNDhEhMopb+zWoN3GP/WHEUITppD9/L486GpNejqBn8jfcj
R/FtiwIajJwJiSHRtGJFcEuvI3ZdaasSCl0+2fjbVN6sZq27OFqxYTO4zm7ynm/x
AxcBRtkebr6C/WQY5SFzCR8zxM6Ov4MmHdxgS0vquMPtCImRXOnItuwrZMK9SGyL
nwwAB4s5XSV2py8/MXQbMAMbC3AQFFZajIofdfbdfoaEDVc9+3Zf0FxCoya83X8/
n2euosYHTqvAsRDdbkQ+bsMz+uIYmpYXTXkdZ5cem6bscg7NyEbkTuvaqstDxf6X
r4YhyXawEC4KOSL49gYUVskK/unhvhsM1aFDdTePRlf5+6/vvFQzJyBHLNcv/PXi
i45mOElQNlPLYOQCHeLEcz+9uJ0POX1RWlXvmp1KLrHXFEsuhfMEHup6Q5yp5D+0
HjH06y6DBPBIpvS/7ljUMyStx1gGdW1ohdA7potOpRC/RWU4UO7yRtEwv4g7wXcB
wV69mfglAQ7XM0LiNQGlKFxwZnhNnBQmRCgqEyOi82R8d/hMwJBi4fsX9nzh6FDx
yQ2RNXQTr3LRY+X7TrjOAHzQgWpe+mJJCzvvKa9aj9uUimZ2zClUQ/RUsND1ldHP
EKsYjdyqK8TpfngMcwj3oNrEdBNG6eJZNqsupo3TUPFAM3ILMyrliCVFzAPjd69j
K3GfM5F7XwaDrmGGIjMclTc0Wm6bWKTyPAl344z3QjV+jpubrzLHe3zVn6juNsku
GMksxHZh3eipkHNuqyiReloSC9bzjs8sd6MnutZGeB+5znUb3awBQSpWQOBy5fRS
mM+VXaNSBeVYB3BEjbOGy0WxqtGhJaNayjrYI0egr0nXfv5EivZdgOAN3U5oxFTb
B/i4bHdTshG4uwVOqAZLxpTSwVpWhLY9tNrDKbiiOb63O0UxxfGnKa8wkWKkBnJf
juaVCB3Ppj2R3JPP8AruNmpjpAJrftqZ3iod4OAYxe4HyR6gVIZ+uwuPBvaRAYvD
Vit+Yjh/dwa991e5tru44t2txLa5bUWms1dg6M3gY0rMEEJdtykJ6j6hA+xnK18+
oKTu00RkEhUrAhovlp96OunLVRR9FSfGOd1HMffoYZrSX6zIpPNVxcghpIWvM8V0
N6xOxxOm7DP0QP3Xx1ZRftOLgiodDWheiVHAIbBmWN7MUMQ9O9PyuRWD2G3UvSEP
XA9CiVX9g83VgeATvmTr7YQr+DRdw9qjzww7ZmAlwHBe7x46aL3bdAz85lfvKMjJ
BQx80ftiPxfdG9FyXTTWH9FbLdk1/W5UaejIEqB9syj+5zQKe//YOY6Vzz+uH2x2
3vAcpUFcqjvJUZYrm7VSiBpq+nIg+SAXpxjeqHlmyKBEnvu7umNWRAxRXf5b40AD
L8fXbLUyVnhN5/cksW24nyuQZ2GGDRItFV0hbbvfx4c648E1jw4upcqV9NvDXJuU
93NAyxLUgm4dRtJRu6OCfAjtjAvp6CPlRglGZ3MrXcN/q6pj583v7y002PYkcdgY
JFwopWoBR3Xx4j9rfBIng5YMiCmP9p9j8rAmwG4XYD41k8yQdOxgeg7ibGxXZW1R
w49u76jXsSw9Qicq2n1A0Pq1lP09IpYDkWddI10hEVA831qikOlcGSnNDP1h49ov
pvhbOEisOUuQY4k6Shh/hgL6VHjblf6u25cGNs6CJXbTgBFQenDwLxkJ7xnw03lX
TWIaqhWle5O/MN7d8eOkOFH4DqVAi1BcvtGNjImpVlEoBmKs0TV7UnaL/x6IXlYt
hsWtmOFibaD0BITVjQBxAhLPwlml6mDbw/pMikb3q+WnP6k+TRMnZMj3wnAYsWr2
G1SkgULyZkC8/QizyKQncph3To3AUT65P3iVFqBAlWaIqKTVUGI5he/XvGvLXp/W
fXmthg0AUjnpmuA+ksei41l8Ya7ycAPCDUm0b21h1yLltykikPfEXWTRh9UQDcmJ
6g604hhTzIZ+59REgW37jFi6OnJYylqbFSQ4yJ3I6loE2U2bHQs6jXQtEmxJQf4Q
rGkInl1eDJY7fAgI4O2J5vgF8IDLu6nq4QQBVMzmCiY6ip4hOOMUec+cymG3bVps
FsVy+Q+IgrSObpCsgs/NHdpAoJBqIU4hC4yrAvaSle0emC2dzb8hYT6qgbkKSL4/
Gr1ILV1h5VK89jG3gPxuZTfmXU7Y7I79qKSyFnEIwEEOn7ts5V4FTc5OFgqO2SQD
z/MKYn38W2wF0RoYKQWvwxLQdSdoyD9ajrJPrGTfYw9U5cp4TU31HZTjesen4ntv
42Wjd/Se66ebecqzccYjxGyDrO6MBSsiJkHrPd4p7pXCG9+FTCcN6pO7a0vHOdH9
5YTHLyecSWh2H8LiQtIWD6XWURH5fOuRuvMbh4/ajhDCm82gd3waTWUFs7+DBoi2
UszEBLFC2GqDCmRF0KLzdyszVkBI2FS8dtTdyPsaxj7Uqu9MKc5RSQ82v5AgTn3J
sxP+rN2yMpBdSx97P3CoKuFcZI8yDiskX9nAkQuVErqKtf2D/3zsfPeCgDyiTne3
1ExIZqxQLDzR2+R2PAv+ial2AUsvTvGHYKafcG6bYt563KvinFlxoNMrJMy2f/tK
C01tk06iOnfDU8Mi4fJVdIiAu4N6BNHyBMWML8YbSxEwSXwxvnDLgG1XzDiBi/nm
CTo2Ohs97JjDXKHV7FDZLhZUWa6x1vdV/2Lx10qr94Je5ShIsXxLRhTIYTAsE9pA
dudajmFMTH0g5uQtdAbFQnH0o9H/eCdCSjfg6ijx6j68NnQ7USBzvcP3rNlgzdMr
ci+VltgZ2saoBwsCAS2w4QSJ+8RhBZ4Q+2QNida6r4JR8Vqm+yH1bMdrzg+cmYwX
+M+eW3gWWU9yF00knvCmIg/wCz4F6mrDhJkoh1Nh+Xk1V9xcaNjdrb9V+H2p9Gzz
oQK78E3vJG3tC4ruIBlPpPI71ty8Q7kxo/2pGToKGD+2BHFlForO9O4CFqf5VxVu
x1N/hrx77F9yBawjqHA2jS3VsRpQdBjix8t0swqodMXeAa91VwcDZoQ24El0AUSo
FRa8uFK39maLNBJ42g3TW1tSrEOKzgn3wP5x6Urf25jjwL102GpY1VtaXfbELjCg
h9A0zssCFMz/KKtiiFPriv27KMhGNQLt9fTy/bkR5tH7wDIq5ot2E3rotn5fx1it
aiTsBjM6kwTc1WkqFSWLs5g7yhtMCOzMXiBlJd/y4A+Ai3yOQ02r1AiXbalSL43Z
huxmvs4Rx0Nyb1UqzP1w4tt+Zk9ZmC7HCi0PHfrxYUqKcghj4rb3SaVU9sZqHndy
ZwLX30beWt++cqkGT7yrlSMFOtC8Kj63CU+AfbFEd3og7fUy+xiJrHPPnnj2NzvU
9BLpjs0ubJ1mti/WHBoCvF7VjDOTrxJXWIXhh0/FjmL8KEOnlDji8eZTFyc0DqGN
nkrhapyfXrOvGbS9922l6KwJ4ED+I+go8fAtXAdmptbCRJ6aaurUxS0wX2/zQQrD
41N8PcFbfyKH8oa0r59lF3xA2DBDQOR4S3ZhvaNz8OPH1N6M+al2rDRLC0dZS77u
Ljc83WvZ6pslHM4d16Mt3BkMvA4+xoqO6dDP5LOc/r13OSTOsK74Oni3yS/go5ah
aid5+z3BaOnCw5k1/Rz4QUd/+yfK8/j1uO0aZs1nZcYBOeQUCFew/0Vn0woBS3ke
UIMMofLQwuuJ8w/g/kt+TMoIMwXL7OceW6K7UgVasy/FE9XPtKA+EhzfTDWmazIn
qqldeIUGch+zWbiFEZ0DEsFJvJc03RXU38Q+egXylmgszZFLtpj2jQtKIofM/z9u
Ezf8oNTZum9GZWTTzJdiH2VmD0AMhveGatd0cKQf1mFHu7KwSC9SvppIcP/gMFuB
zfd0jBIaLc0zlqMGEUKAeS2jpUrauq1TZZEkmG2Y3Q0xU0lPULCfKPPrTygc7BMw
GXn39tjfBHmR+njh3XnDfOfQI79h90jzD6/4S+c3A4iuQHWZA/ADu5WspCEfDraP
tK14ZEgD99gmlJOB+6XNUYIVlIO3G4fhxIsKGov/pwRaXke9UAZjaBqA4rVxiz6U
EHpb6pDszP+nYayhA1DY43Pcn13+BQaKAK4T74nOdSApKXEUrjnebFBfD6UnyNHA
SPzZJE9807tBV0aMpfKzhlX+kPu9uy416beKNxLrUajmn4UMc4y6o8uhqCGiUBzz
IGfXH4FPK+cSJ1jf/RFNi6Ue9RNWHyv36KAL2Ng5FUFoxIW4H84LlocRrwCsKyQ9
Ru7jwc2oY8CpKhCQBovJmLI5bzpEB8wZITJV9MMgmNTqLjABUxynCe90xbuofwdk
oL+UkZAxIJKuZh0XLDdXEbD8Ow7coEWzpz33QRbI3Jdw8EM4HXz/WA62rgO89cwS
zEaNgZCmBvh4OAiRtf7u/lYLP8LfV56LS6PoRuDLaYiKvJJXOhOARwaqVDPvmsc9
Ub+pNDURM1vH/jfooqdMd3Gv20VswLmHFz3pS10Ox07fot8bhOVZEWbZ8TbO81Xm
IUR9KePdue+OovTl/w4fF80ovtwQ9aQ+3gK6syXDPLVWe1O55IMZbYUFq/hu3MHR
yK/D4NgpHKVDjLoLDfI37BTRNMJKmK1TnfQ+fzXOdntwglnXJ/L16tQl0X8wpBjb
jeIsMFYOK4dTFwvaPn3fG6FFdRl5t3cyCEjeqfoegdtdvtpyesW9wLiDPv3a4sMl
4hg7c0OYjNuZFQbqlkja2iZsW9dtro3yjP6ab67zZRC+1XBF5cxPIb43LTTb4DL2
uwJOigyPqqk9vZLscv915NtuRoBm/B+Gwtg9O/hWuqQd0ykf/MQV22xLIeDkjjR9
35k7lGjV03EvNmTw5ndOVR7GEEGU75H3E3oFDLjVxHdnERdFzgVWNot2WTTu7N5l
esfGB4ayZfoXzGc/2qElnonMzxWxuuzUHySvOL2jTYp9V6Gn3P+45W2vOWsxAEAo
Pcs41BVDFVlIs5aja5qQnE1/txzMxAkphnAgoqstR82JlkPClzb5JVBrJaF5h80X
BN08GLQInK1FNDk4AlyhR4ukuHUHlDeXa9gKe8qLB2szxoMqWxn6zE7T4SZOKj7g
Kwvldpwa/tE7wvtWr9A0eoGYUzMwc7LAUXsR2CTdjNNeKh/RA54aiSDZuOfiKAV9
tgOH88exXj9R149xyqWRC4F13D4/LDHb2+Dot5p3FHUjExFM9uFRBbtNLXqupYV4
6/A0iFkRn2jsFIyjR+dTomLmg1AuECybpgAC48lGo9axjW32wvT4crczZyPpm5Uv
cvRhvmyoZsvk19JskvZKKePzI1BplBY5EEIkM8jCRJWTl3n7oJkIW1vi1yRz6keb
/SdUIaLiH+SsvpaUaKnTR5WzmHgfHsDL/2060SRGIdhhH5U4oQgV8vodepR9wTES
MnXb1kqULRVyGqlMSW9d9alUFGw8xE8BZlMr+Kt11xJYjc19wM0wCE3/Nep/zRiV
BJMJaWULs4awHCkmyDWge0ulk/2a9jx3kqHCrppriduEFmzxxz68FlT51vJOLv/q
UEDnOEA8o8xgwBPCkKYPbI5tlz4YJcFvmz+9Vqc6Ly9yxJ8MYBs37XCQI3CO9e0e
iPTKh+crUd4Zy631afp/F1LeeImfN4Ze3PH6vI9pmDG/w0iLOKQSsh3aFl2+RgBO
ZaOiM2h+rQuQBDw9ZC/6ZeQ17C3cxhQRpnHMNQkVgsXR56/dyYLzc6GL1fK8zk+S
7I1djmUny81JfMZcoBtukFtSvWySRpQblU2g67xtPUzdKt9W4bptiK/ydpOWUlDK
il5CvigfgUerhgDuDAIZP+6c5CzHylMOgJxuP9dwy4JYGZU2ntHBX5afp0Xps1PI
LTufec0jg9SAjBjQOX6DWg0/t3aHiZowL2ViRYs+0k4olDRV6mdGJ6cnu7kTXZa3
PUlVeWqFdqlRWBuKSxZpTY1K6gVztbmTgIRegb+EgxRis/4sm2/JDmNtPiDzqcJP
lvQFBr2TZTYehTQFY8H+Z0QjMWA1k8zjn7mttdZyCoJ2vWn2RebhVAwkvkLkTIwI
irYOoDgtogxqX6Vmn/s/KLpoygVUz0PhsPV+gMLMf+Jnn8wuJ08NSV6wy/kTEmMY
g4GuDZKax/YRdo43Bz1HDTmjOHSJN27MabykBii+sUUR7pP7TY3Od+CrI2lX+OUw
kaprvB0WfvSFpfyEbPHRIOP4tGKICVRefrCsqL+/F7yZmsWRuPL/hz6ajcCzryC/
SHXM2HaXlLfNJg2+4AEFr25zaRJ1tgbpUOlHR3MX1F3fyruQNcM+rlQRFBZyv5RK
9oAL2IfmbtsuY1gurqbdEbcmdTcu3zodv9IqF1x4XAIHqKLKrP1OoDVEiwlklnKe
dM2R4P/9Vyi4+VZkb/M+2IUCsvobKU5/zenaPcsp2/wpiNsd0cCIy/8pEyMFKYCK
nvHkDe/xaNKb48Rp5ldFX8GAbKbBWUmNyhSK1+EIJbmSjjg1i2LRTrEgwBgwZTAA
cWAySyHHh39QmywR97FKqFGc9tT8IMU0hz399vXiAoe+/Ked4WIbQuHMUk9EXh2w
uqmJtVz6B5jhEjsy5NhkviG0B2mOfvNmSIn46IACK/NMWgmuWwTvQN+W72g8D34g
LXDObhecKZXk77Uq3MXCnk9IH2DWmiwLr1FkL4anOb1bBxF73dcLqepZryYUX6wx
Slz6RuN5gQn5p/oOjqbHythjRYRe2YbNQLQz3vcqX8WYUwew392g9dRMsBR69jL6
lGZSynH/Noaj8dJd6ckw83+kekVDNIZID91hers5Z7ye+FtqdIpsl2Z470zJMCGR
aPw9qIRBdNKDP2oBpvgsvnU3pxltfH1DB3eQeeRT92qIdbUSRvSurVJDKIdw0Da/
XygvHPxpnXEjcEGslULCCns+7uZwVyrstL8aZ8x9MViFBvXIdE7CaVIRbn5qwHh0
1JmoSGvxsN5pZKUOvm1epazsgxijZeulL8TwlB1oJCFmH3bdJmOSboEDsjW84bGG
oUX6zN/lYP0+De5RcZVZ5smKBNSq3sAOFbLft0b71UBOZEUsUCKLglcl8fd2boJv
gf6+WOngbr4IMIaaHt9pV9AnNqgdP8yfAOQhllCbv5K+MmF9EwFUhYbixMRUhClP
rDkPbm9wl11F5H++KgyNy9if/PzlsV/SxvEmAhF6lGVu7eEw6BaijNyF3Yg/0R5+
3WGWunZ5SwBG/8VDcmnsskfw+S9ebpRcdXMEaIWDa1xZUQhDP3YNgaprIkYPip0o
1Vda+h5uDW2o6btZpd0JVNS+TFn4PzngD7Nnp4aJtXaVzR/MUZ7m+4pkxRfViBA+
pe4AJzEUluAHMAit6TY90O1oCmhlGHf9tlG8DlxTpUwScGHpeovzE20x7tyxh8QA
XQmKz5DIrwd/WEaYYWy2mmsdc3/tzLmClbW4ng98KmJ5AlOE/x3Cm0NzIbURMywd
UX7n0LufZo5OEWyGd3e3axIsFym91ZKnD5aaMoQQAgt7JYbwCz60tli0PCfkDG6E
EosFI3ATJw7lJwdv8wIqDx/RXO07iV4VVofif+q67Z7RfmfEAisx6+xtaA1waWBB
L4w16HPUF3GlxaR9ELnPGTcSV+Q06ZoF1krBtaJIrFwxCuA94xux95m4VyL/UaDc
1fO6iE9sPzgaCefm5kM0lbf4fYh6hYL4S5pIsRWwbdTPckh3J4lT5cPqZs+AXbhu
cDv9RfZAz6Z6dlnVn6qOw3/aYcdWGmQGzIg/XbJXVi9ADSNEk/LiuWStCd0QSYLN
4YxVFzRaUO/G4RdGwTjvE11uX0IOPobRljFNOcJ9yJwxOSCyDJV88RxAOVezH7j8
3GURRluWn+Z61G5cn0ni46JxayDSDnJqu+v2aaoVmI7VQHbXOsUp1UaAITAfEqsn
txK0u01qACN4NbIzgrooHaFHATV4+1rm2ckvW7jlZQNwlPGuy2vAmA6LXsGMigiJ
1jQWfhVOOaSH3HfEisH82B+EwcEEHb3MvwjwfipGIFvi+J89tXmVcZHOk9PWWQUr
pVA3B5In7oMHMA6F6PsH8QIRrZphARXKEfqBhxn3Jtxn5xyocA8CB/I0BFHis4nh
/fL8nFbxmgViJtJw0zQAlxYIbVNop+1GsW774InRyfrkgDUSC4eBuITIQKDF6ShO
Tqp4Wyr5TlLmaXG/SRGoyrqX055+Q9ddTISuqFfYA9cjws+Z+l+piXEtTnIQI9mX
Vk4XGtp0UJqfMspss449MFUpyiHOP87zaAYdpn0Aw2QM8IsconwjCo2kqeliPj0A
2uCAiftvIhfEQ7X+Y/JUguE809272r8dI3cvoj+Q7cIpQwltoCET0vOW7dv5MGoM
8Fh+vqpqhFrSrNYifJMv1b+cGyJlBov+422uzM6JCL3orRgJfnYzFMN1lwgU9GMt
fca4ZGjHsNQRAIx2WFmGR2rkP4qhTz6rif45cmRUczAOaV0v9MTdgT/l1iocJkOz
DYiq8ZmSFE7JXpm22T7yiBmToDfeYjgPBv/NBG7+7qQxs0sdbA2cFTp7+muwGq22
JIRDiMOxYZChCSYYjmkR2CF5NQuhwNKbbaKMy9+ydQuu0VXohncst3NqEn4XqXy8
ZJI/oCwPpuIfT/Q9yGu74IK+qcUj3YTYtlUkKaF1TYFwjze2sjWUy+Qf06V3pO2f
w+XraOXCx0FRFgGPp115HZh+KMAeeOe3om1AJ7b72+bS8itIGXc455CJZsJtEPxu
E8Z7dVF4YbsdTpPzrjdBlHpEIl6UAvFeZhcmTQK74UokC0p34NA11byiFXCs+Fvl
boLAwukM3gkjQdUQ6Ktul86hhi18v4clNHpRRuREPbaiWrhawr3Ubwuujj4Zdu0f
hCfWSNMXPdG67svdd9Bn1krekMwea6YAcf/jAyIDJkRChjV0trZICL1XobfLC469
FZNNQiYR1LfvHIOZrQz7HSLlHXxuluNsRSUWyzcCy41r4sYS7SfkXHnRkRw1vAF+
/PrwCpK+IbmooXxQcLzQmuCK9L3LoifNdx2ieA5q/u0rmgoanUP1TbQn4ii4xsRm
L8FuDlC8utZbJago6ZWOKdLayXZJnWaytzifXEskHlm7k/+BoFY168eeJO/JowtU
QpPjozHA9jTMn3rkj83WoYrMENwAHRcHRI+9okvJE8w6MDfQrvlJ8yz6pBBSzWIS
cY8GbYqM24Ym3HKJcQQxd7eGLxvkxOu0BWRLUFgXlYRCzbGzx6DmVZdZmg0RvlLP
r9qF4FWQSHVOHMmM3KGqp/FGIHcqbWn0zhwurBUjbXNQh54XHGlrLpOi/J96aQCM
tc0THVdT2mhukkuyJ3Ivhe285bq+JB9QrOwycnjStg57bj6crNU3327PyyhmJ3oS
kKPUfut7zwTGPE30Km37o7tezn1uhij1X57SWNWp9CfGvz22PtEikvoCxSLxeQBm
Rk2bJhMpbstQKKEJ1Yr1ge7Rqic6rOMjzeUx7XiiLwIxkJFrLpVBeiOsr8ZUUN9/
Kbmdffr2Taprt5H1va+CiztWb/TORzBE+eEwEYkje818TNCmmdMu7zZ7Fq2TwNi5
7j2IgHc0flEpNe7WDCnvIMwY6XcvON2livApvu1vrGlzMDvNZ0vz0ENVVr3A5bRZ
Xuv1e4/imzCliPn98flZZv3e+DNo4/NlOyYwSCilr3gN/7+kw/Y3okGZKDIwrUCF
IDuLBlIaNjRv5ncJK+xeDxewBGUqMPniPaHo4gKhcj4D/JR03PU71xLm454KbGnq
rcrq4vPaEYARcfktaZSv3NrunsLKeG4JZ/QoIuCaq9vVqe2o6imoU6peP1OxAN1A
/WJpmg1Z+gLL/IrfJ8FWVbJ9RNcYYJBk3xAgJB+UAVFnyPRRC0WXB6Fdp0+qgRar
pWaOoVrNyIO9Wdg3S0Wu5n53ZkpVZ1pCN2Of6Vn0HfRNmqcBPJe9LI9taguVQ31Q
Xek2jsOC6V6mLODsUSFAjoOj9k6AeEik11lhHI7AgK4iPOkmILECZV8hSwIrJDon
2HvL6+LyPTBuDQzbQOifFBNKiKnKe21ZSJYPZSVbArxRBBpele9bzo/M61twwagr
08u/Dh+MB+ceWVZBrtWRD6Qt7EujGgBcg2w/k8lteySOzrMs3S64aA9B7gZ8lloD
uzM7/MS772TvsTx5Mi4cnWzcfEXX2IOd1C4Nem1OSH0+E0ir74KfxKL4/0o7syPi
GbbEicFqj5CKy/UiR8KY3wB3CZFdxU2WqJkIugWio9z4I9Vnl9uEmyri2IH2CCVO
JHzDTr9EvkNw2aGUcQA5kqyIdvR0uAu9LnGj2y2n6Cyhqr/SmSa46EtUpQJ269Bb
zRNVVL4NvJ1Apd/edccFHMlmI+N+5nKIWr7PNZCNV4hyKGwU9fPc4zR0acnNEBrf
s1/inAPVNulad6Mtq2UF2usXB46LgzhdKk+ryB0suuXxXFggllPl3HXU2pr6q3XE
D9EOn7DNEFNEixLkhYh85KEo8LRjKDheJhtRXRNexT/VLxJJruWAenpnAcG9Hoan
kPMqOTyXi+AtrSpnOSGwfTc9Pksn+IWePNyXuxTELLFHHXUu04L1h6DgcVKVR+fG
06ghgTxIY0C0N+JRg3EcC6dn8/DZ5+78EKd6YIR5Uts4nnWdDAk7wPT5l+THbyum
fTV0A6TnimqHQsryBZlDBJckn/eht+dt7Pm8EQ5PqDqC6Wz4fatcjaQbyFHdyEnU
zWX/24AwgMyfrrGK7FNAOfSj7UAFlIQwuI+4O9k79IxTVOsk/ObtN6ZlP8Pfh5P0
By6L8aFQMDtR/86EwzoWdY2Mp3zNMPASA+u2r9rFj6n/SfedThaWX0Usd0f84deS
xgukFLbfHxcBBXJIkfipm61WDY3m79CtHp8wRQbz4xKKknX7JsFyiDuR+rzTIQUC
hy4anj8BM8q0RpItoHClNRg+u0AI8ELunn1Q/WKG6FI0d0NfesdfqFPSXX/wjVgd
CEGHL91uxPLdNS2s1DV9lJADDSWmPSJp889WCn1lX37Svn6oHkSJVfafULZ2rp1t
boKE1d/mWMGz7u2pRQaPrSuk6ADkpABLl0EXa/oiZjjH2wpltQa5PkrxVnhtMCX0
ZjBS1fsdg3nSi0r0/8EFj5gYel0TuOX1nUWoTyElZdd/TDBdt1/8TTg9zJy6Mgw4
YYSIOMR1JFtzvhePo24ZCR7FB+wX3/UtqdPMXkLmqKOUeknVBk8z/XKNCKsbQxWk
3NdLFnPV7FFDIg2331JFkLmyOz3Ut+7GFRKRIHmAA9rhNbpV++XYm8uVK2TcvtFy
adzWMVj0Qgd3vg9wdpKBPzLEKUXO+j+S8W2Z1OaLU4m4z//4G8O52nJRroOGUDjq
APt/fpXHB9eZYB/DEaqsShus/yhdGZsC+yIqfGw8yMOaQSxqCUdK6PjR762ECnSO
wH6ZKdotWlNS4h1bFs4n3FWKnB8rWWICVn6kgOk53tegCvxkokVQ9kidITAp4Sdo
qHtoR4f7xqgwlvnmdFUYXI9plivo6qVRRjuLMBGg4DFMZaY5FY9IuRTBR3SFb4MY
Pu/3a8eyoFyZutHvnOMhA4VaVSuraBY23cc86Xa+8tgpnHTc6ueb/wHbXFFXk0t+
dr5okUaLjC6xQd7hkE5y67YmoOQuPg0dxMZxS4HGziExw8O2etiqm1JQccQQN42x
6vqjp6iZCxnTnB7dV9JBpKobHdfuZ2t6osKxqcm9QLDT+E+gasF/5WJOWwcdYUdg
dLCQDbeVPh7r/hIWNihLtqdEX9TQ1I50q2jkQVsHXsWEJ16xojzM2cwWYwGSvkJO
nAIec6V3LtitgCpfa/JwgVEMQOr//8q8fYrUywd0a1eubtsR5u/9ZFVWXzcqOmIi
MU0/9NxIwgZuLzwm+evMgkz/jIfYp8tLljK0XKmZ3Rpo6kTnnIaPBJBdW7o+/r21
FzOTggglWOlPer9QhWPah1sd2jsspzExNEsUevsBa5dCCSCmISIJg1AGdqTX4tqp
wmWvGohye4lwceTNwNH5lWvmgKbz5XZLWhUnF2ZYG0oF8h2w6eYxqBHcBdlvQTMg
Qrf7qwwvmVorOg7Yq2dS8+Z5AU3v5oa1zzi1VCz4zdIMHgJEjsr0qSzFzzI+PRny
GwyOD7ZKcyJiePgIMNJoMm3RmbnFv3bCZRsXCt9hb8QXCEAV0plGgd3JHtBRmBIj
xgLG0T00jSHQY8EwyRmG4JT8vGaO+t9aeFiutpooUz86fhlkxi0cusUifi5ZvP99
24/MooB5V/qFsJ5sgkXuJdvZ2YHbxSU8h8Gd0BTDLYo8fQTh7ZtBg7Gss2cleRAT
D2KOuxWDugKs40RS7+aerofpiNeK0Z7drxtc21aEe3g61V3340O8ptOThfzEfU5U
rfXq++rnLzIHsq+sSJHl+NC2YZGywkqyATwAxKHSpnjrpIRnmCj1VDMMc6R+2szt
BBxd3VQjO7yjzNEioCEoW33gsBobHERn95EfHcYgEOPSprkb2hO8WooCX5QiWzIJ
hF3lO1l+gqqMvybq4a8PD9/5FvWGAkgL8EcAliW5Ze/bTGMNt4eHlFr1Hl9+2ZhD
J17tSps9B4MHqbwfgwGGLms9MYZ/5Sx1tykdvZyfIlIUFf2tqGIqOfLOiEOC4joI
rVLraCQkS+a37MIhPBHr93O8P7dcjUN9+HLZicqQmcargxnXmnSfT07tTQyln2To
c6JtyskucEigBx2Zv/P6YXx4OMFz5v5IF5rAvQf7MCsy/wnThYb+bxnnIpLHgCMk
REv4YWpEXGvpMBpln3ek8jEZcVL50I4xxnvI7jJ8Wn/tRlPm29JFMa6+3i3HQLAp
QW+vgzmkQ5JIPL4vwA2w7Y3Go3kh/VbDD5GpyD7ccYhOWLG3jm9LAocqgee3GlJr
UBYLX2Pr6rkyju2UrtoIkFDzRiYc/awW9yWnjAJiep9jaaX6GUXYwQaRl1H5uMUi
CUjXV7GkLgrfUj+RbFW3y82jbCYirb9J3KHkoXDgFWXPbFm1dDjcmdNIhbws318I
kvcFRa+TvNJvsckgZs9f6AAh1BSSPsUDFIAh2Ulg9Uta90RYhjLOrd3zBbH6RK0w
IO+Yj4M2b+7ZCWk2ajA2qCjCL1U7RUVEUOV/W4qlJ5iUEHY2pw37Fd+mpZEp0nei
7X7SdSAd1aRfVNOyioyFqJtL31kTosIrY7odbJgL4S3OoKm8qMbyfXqr8AmjwiyI
VaFu01F5HeTztO9nKqGwGJ+exZQ4lzRK8rfgYGphAZnmiLyu74haGMz0K/LLY46H
dchc1mLlmDFQyw6xaw/5vQ2e9Nod/dkYhR06k0XGXrt1yQbXJvsaE/e/kBw/Jg5E
obJe5BS42ZamZF7Ufaqi5kEsx4/OlrrdLf9GWqQNEa4ZRyonTxj2cRP+7ATlGeYo
mVgAVOYCF4r+dy/RaD3Fnj0i6a7sVO5/I8hESA60uVKBW8TdynmkYmeyaU2yjpHp
m2hgNcOGPBQnPQJ0RB2dnQIiaglaHGg747nL+xYhRmroCzgw2pmDCyn1Y8Gs8LSl
lKA1XR7EIZQg3OR4GVsKVPcSXBdjYkV6IdcKf0rpKHd6RwEzSdt64KF7wDJb63DE
MPEy9wUcQT7LkbAvOl/YGIZW2VAj9jKdRvmoiGSu5Tg6XUQED/DZaQlAj0r55UYr
E+iR0KscOr5zFiax9+U7A20/NfwWaL197tZz76AMt+BpiXm7A+rIG2O6Y16k4r/L
P3Ek8IGK3vMoOPhSTr2v5oxbxlgAo11U5N9Kq7xH1SEGZ3AoA6ruPYWQoueshKen
LR8GZ1B2w5g3KxHfyyFFiwHzyv+V8pzzD+OnbrrlyE1qj0jkh31pgTUeAPb4UdTA
ayQRrnt4MwvyRotCBuaYYhURIapvMVVE7/vg4bjtcykC+uFms1DZyepp6WQ3GGV6
djQXF2ZAxE9Arw9HJQSdxCupA0ujlXhs8xwuxQgXkrCgths3TbguuffoQrvp7aIv
Mp/lfa+zOb45UsmE5MUtZdgOrc/LQAZAkF78WbKP83Thu3Us+LVhyeXmZKqC+ZOe
EEhMn4BuxCLkKkFL6e5wRF5nKsIo+ZXqoCKGNOXH1HqBA78/KyTBx9tqAndfnlU/
QC51mI5ssjTQ5RwtGa2LdkWdKxCkBKVz9OU9s2RQyEt3320lRmZTvdR0oI8hNBnO
CjcQy20+rKQ61ZwElJk4nYnAcXzxRKQxIn/Sd+M2rBuKa+8USWWMwWIRXNeulMaO
s1g5zA8HJofJ7acZ1naogEMbleojVaSw0MYvhs/saaJ94EaS8xytTNNYM0Q5KAJ+
LUTWnm+z8I4v4z/XsVWELk5gyUhCWztV6+hdP6uI8UjghpwmH5xqoSLhGUdVoeZF
ubl5IWXehs/aIh/kbLDld3kj7h0QOPusGxxiS+1nhxvqAbnSNv+sFY7Cpg/lwurg
wTCmB9LMFKirmh5vpQ6/dbA835Ua3JSWV6M/LiD7tRdKYlUHalEUG2w9KvtUofk5
2roxPYGflA/9dm89uLDDsR+PQ35iH0o3LKyicSBhPXSdL+Z6N7T++HsVFr49a3Eh
bmfhnR+T8qWIeLX+vzbseoh9jclGTiNOaAB3HRIEE5eMZgAfHkIENnM3q6RTIja6
lPSbgT1WY0PHq9sfL8O+/dlvIwGSbNHmxMW223Vx7x0fTrXQ5ltL8Ap+JRCF3Jzk
XIs5Tw58owbvXtavUp8kOd1EmzYTgfLloCMeaebY2tNqMooLD+fkUY9rWKE5n3RZ
YGk00+m4rbwRWAY3EdtHT6sHdNnxtUKI81L5EtKUAxYiecxKg68AJNRsUxPKpGgA
gQTk164JN/bfCQRzMJ/jvjnlnjID1z9i5V35AQ/ZdHCMaXGbbMuDvt70SuvzvS+q
sA1xII7sPp9cx3brAqRLBGMzpHaZaa9IAIrHziVoMAV3d4G35Q1jxRGD2ePT4C3E
vmptabeTcQ+gpnGJJZgAdBrO5Vz7oljE0Gueuh76UjgufHT7RVjNLIbp4NDp/jCB
HgOwXmVwyjCothIOuNe3NuGmtkAU2WGmnmiusisrXA61rBDPm5yIPuF1BCWussXG
ZWCXfwJG5HJUonCXTnJ7T+d6J/aDPnEnEdTiPGK1i2MRbA5P9OK4t53mn8pWc4dn
KGjbBKj4uRyloMsTMLpCTh2txN/Dr4aNe5hEcCrEbjPBZg3YKSv0geg1aRNP5Mzz
Oj9/DfgOVakjmSmVJU+IZO4rmZvh+R4BuKn38KOK1+6YQgnxIOs+uZz/1ty9bIK5
WLlpLIsQR1PImy8GqPl95ZzO1fQoTWQDhFGwr5YUBBCcRgrNdqGXZ09N/jd/KAWA
pD7AhZavOGCTwKj2qVir5AY9T7m505B8q423atAhKkU1ZdpxqjE3rL65DqL3wRiw
o6Ykrk7e/Hpwvb6PcrKPLvQxNGlCpSefNKxUKiBRvAPCIdWBM98qTdnEYOAT0n1I
IGNPTL5ZFD9tjKXPgIloGHAzVMF3L9II1pwPs2FAHtS3d58BWdOXTI0oknGw+Y5l
EBrCmQCtPb3CcZnYBxlegSKTi3EaW0BN35oNFqkjAX9WPwvJ9E7j/+k3gaOLHT/k
kdJv5ReOQbbToSdOINl6GKuvihB3lhKD6q+/H1s1jDNQLW3afX1CpHBNFi6AoPd9
Ake/iEdgHSh8uK9ZHUprpaOPBIjKeLM6zLAzB4q1/2vJXhvaAJKb3RhL0kBRtTSv
UzTJ+T7Uliz77Xmgf/gUToeYAZeO22HlMNPAjZ4gAWuMLqXiJNdYBpR+Q/oMgSvc
JRJKNWBRycIjxaIxSHtEWGj/Xb/KFFfjBjcGhaNxd9vNvOv6Q0NJlRRRU6TNWHTH
Rz3SDw+f5zhLsIyLL+Nzfe1K7Ix//0dvPVe8EABTGQuJn85HXKR+zEValkD8uwQ7
xjPide4yvi6PkBMXSpvjLCpO7FcI8LixNOtCGG7RSIQ6IEXNcNYD40dhs6ugGDr1
Y8XgVTUhozGc06K8nX0Ni8t66L8ywPH94EPihb+DGEIJLCNpGj+/+gyQPwBVriGl
6njvm5i+Xc2KcOYckEw31ro/VOquxQ2ZlnyDu/JuPBwxyfg4qKhvjIlcn7/yQzDB
xrEc+OTGSt2gU0V/c0nEzYausFWr/qBzvgxoWEzwM0rhbgVirR9awhv8VFim1M1H
ADzRjAwBQHdQSbiwlw60D4P8Pv3nUYRuBeAr7UkrdNbQ760j7TkrZssA22d2QWGW
8J9zMgSW8x7rbnwqXC1qMxOzD1Jm9q0Y3Aj55Rx9kp4j26/IPiLpYz5cKlzHklLw
5gaBdg1t7gDDtxQrtwXAoXTlmfs5nEfGOlf7Ri+x85Qv+8KXiyJmLui/9GYsm39U
ZYt4qjs+bBlnBvmMtkaytF92FidbSbvXPzq6o2uFHiTBtRVGjzzviSc6iA6fM/YS
IoRh8Nb++/NUAkvJbRTe6jS/fdh3h/ukt65pSqJaygFtmIyaEz5iZ2PVwI/PUhRG
0xF2GbeWJsq8+0FsU7/IP8qUuDDueLDogQnSt3304BYocrREfkokkmDT7BdVRNjY
UGXDHSDrOUUoRTFmeB/rIB570cYyd78mBbPv8XkbKVcW2QjRapP2vAUaKlUSE+/Z
Ij3Cip4GX1yd2JkUcSY1y6/FJTprBn+QfZ3xVdKUHALc/D1/c3McKmabWzmaXHdJ
5srsPLzUVUl99bJ1VYBJ+SEU0avIBnlWPY+gLsbWxG+64wcmhdCYpl90ydFo8dMW
PtEHPLiRgKZiDi06CUh2dup0wq6kgInMmIpiUPM/4PVR51XqhGjSFbhSBQzBWkHz
AXVj2jlRzQEeNkndhtQM9FfQJDdDBiyErBCWbiGQN6pzxXYxJTgGnUKaqnykI6Kg
cqrCnhqfV3WXYmCy8EZubXvQRHrggM87E/AJ7V/ykziM+F6MOWrDYAAWMCpLq+v7
RIxtC/OKEwS/MM9m+y1Z/eqF75/1Xrv/vJNlenI8MoP2qbHbqgXyXj0EYK2Qvpzb
SLGGU3hl2KnpvwdjrWPF1Pinaj8g23q2epTBL8YAJNf+P4iQYU8bNOZFddwhC/OQ
feY87L83QoBC0sSGN2U4yW4OZfaNAXkMR9/ICFUBR0lu3Z//Nq855pHLUlRYiNOp
mNiPIdChZcAigFiOKgbmgdAeqg3qTQdQhSN3t+tLJZOPOhHj+MNEujdMDhBC1n5n
bn8ForFBaJQu59EsBF/CY8UfGn15TJ7V2aP1Uzz5JBZydfnff9ipyyjmfr2I13ur
WolmyYfVT2KLpKjCYdgPYoRCXyWpQ5DOP+aZ50Nu1HcDDk7e+0u+CgKKXyDkjob+
O3T9TV6F80e7fSdh4EjAXcDD4kepQcQhK0pGxAFZz5FP3UrHupk3wafIDWFLi7pU
YsOYOflX4A/US/NLLET8ETXnuwsc2o+3Si/QX8hjKgbIC3XW6xOx8yMOqhgZ/eHn
H3YkiQrGtWoNeTHFnczLt+ElKOuhq4V58eX+JW/PtDefr4/U7X2qBBMSeJ3EdLz2
zAelD4JB6nB61aeQCb7it3jHS5Bx/GfUO7Uy427MQJH46SGVFoIVoGEtXmS0C/9J
zvkDE4aJfZRaUGqtliPRq6kSaWyfhq7kC5sonopHxxWABnzwQYOcicb5CDL/sRdR
L2zqPn3LxSUlp0HUmokAlnw6Ya1vJD5mrkxZ9txpufiecmBSdtO2qqpcyNxlDjmF
aSYEh9FEXMLcsGI0dkGCpbimFxvr6JobdNYT8HpI87H5vemdcZ1zf6bgPS3hJ/pa
IP7mLPtEOWvGBpSBd2e08oeIQt3oUZ20mUal2JpfmZYRcvuj34gau1UWHFTZrn6f
VnpuAnrGuh8M7PfK/YZmmQYDhvuZlGn/8RVgjYu/bb99KN8VLGLyRZAbUw+HT6kb
1NrE0sKO7PVhZlguNPUWdOETXOUGEFd7UkO1bEkiHXIdRhAGAo9IDCOXKK4AKGBw
23BeD2fOweV/TVyNhkezpptER6RhORog5sIJS9HPUdu4P3wpOtJftQOo3oqXtDHh
pSEZn/S4sffZ8bx7oj20HTFvJ+OzC+2O/n7s7N3sJWeOCRhYLJWcl2/pVRtL221e
l/yrn1SpduJNouxTl0ycr9WTfzd0F9pIl8j7v3biIGJh70ei+lZ+8rc/CCQEuNls
51+IqZD58OrmJ6E3rCkDWl0fK4gMSl1w3ARIvr/ygs7iZfEC5GFFjpxHRYKp2GQC
hkbFq4PH0pxjxwv6561ycNs/0OzFSdzTkdz2csC6uSRFqa7nnnr+PLhZjfEaI8pV
R8jwWJObq1DwEd7QmkLKz4AXWuCgESAtiUutbE+ehyWsftXg9msw3DcRUPdzhRS+
8bvJ5UXJq2TDxmgul45D1ENjiCDhgN+eZ/uD9Qdu2APrg2+wEPlL6DanWQl8yTBH
BXTZvfnLXqZlNzt887MeLiLKYwz6/TzFHFmuud2K9bKiPBRTL4DNU9H6tmqDWGsA
D08mX5oNbwUCu433t+PkMRA8bWPG7Zio7JkvbumQSeEjvzVjkL7uXEyExtymMf/B
tNSRrSZo4wTd7UgpMmSi2u5YqKEIFjPs7Kc3pwUKpP4N55G4qIdCTSMx7OR4eGvD
JymI3IUcGCH1lXMMJV/bMAHEQD25DOAvFujXaSYzXMW4WzUtUIZnGkVQhCLmut1R
yDfh9QoePQk1BOR1lMcXFnEu1AC6yY9iYS9uRkK6S3hSyWbMu3IR4XzsRQ9kLRRM
R6Wv01CgYCcebHqk/S6Sb/YRyDdNXgMBJJTLicdVsQXG162baztcWLuRv4sFRaBH
KYKcNajPY6yVf3rSlBzLTEdasoVliUK6vcXmvGNP1iti4D9I72BvvLop2gEte3jt
0R9f+YDV8wmIG2vGYOyxq8ynYKEh/FnNJff7Qx2c6k4GjU7bPKn+/z1qvR9fz+iR
u4+0JWjEem4SZwCzT//Hr2CwoqbLqoj8mEmINY6sR2AjKgdJFf2Yj2CuZltDFiXU
+99SvTv/9B5F1BG5PCXD2ooWEmGLG3TlsYPGSjiR25Xr9wJ+ENArlxfeHlwLrysP
f263CPW8JdSy+exiCJs92PO/8Z8kts15dqst7qUDe22XHGgYu+BUC1ak4bPrulHl
mjPBwVelvYWDcItDjjpkWqt6J6Mt997/U3H5gSoEEwBnOpiMKT1ZDCCe9uIXqrXM
568+PSkTz4Tos3HvgpjmMyDFg7awYYUcOOWo53ERkrgZYUdlNV2H/SXmkSu5nQj7
0n7jZkbm5KVXkaKL46cD9BO6DTshl5zPY2+kzzc556iZVFjun5JsW2iwE5W5UWWR
A+iqeZhvuMudowAYmh/Yu9FVm0l+2ahw+jpkClu2CosZ3PLZ9ib87gLoF4mqdCfD
pr/GBfWRr/fGVBx3TAuo8xodfO84MtkCx0LNCtOn8eTnZEYgFV0rJMSFHMaEuy5f
yHGkCXG3ttuwJltJbVs4fUidoDx01tHv0CiGGn/9D0yVbiJCz0Y3GFNNfS99AXIW
OfwScgs4qXMnpdDtNJ49HkaNxTyTfT7YvC2QtyDu/6V8xrTEbNaywuFuX/0xZ25H
tFSl/jHCvE7A8/mUVTBBGImS3iNdKtLiQ5n6VdRW3TR6CXKIs4n/r/c5su7JNqXr
QEBPEuh47q5qRkVAsH7O/bz0j5SMPfIsJ/KUFKBD9KtuwXUWDikKUYDtjhaFK+H+
BJG9Zr2EgseMHitaSdlUfPUzuKdwNQi2582UU/NsJ2cJ3ePoqVW0cTT0Xf5Dl6ul
nwmRSHDwW3egl4nvJIPaoePdEAfDqBgu5BOlbxYLlOiN5RuGsst+cCtq9TqlKdCO
NVdbeMBP3qVmP70GLtAJnKThuxqr9DMcSw/YcXMg07OTa/evcZKmO7it/VyciuFM
3bhd6/gxlWwRM9Bz824BgcaB7LFyuh45ILGkLyvVBgreb9n33rJRd5L7aOcyBSKK
MwMSP8AUDJi4Q7/Xe8iJzImll+iCevBeQjEapygRwCCzJowfhLgZ/qfuT5I/Ia6P
t+jTav6WvdAZKnI3QwPdM+zQrp9KkzpJjhQEgXluB+HTNZm2v/nuIvFBvotYD6Q+
7MNu9+Y5udYpJtN6Mc3T7OmPS+D3K8lJSpf1leJWGHMo5FMgUJ6PdotuXw941Ykz
L5aCcNf/Sznv9oeysfc2zm7HaTGPACAS9J+zBc7/gH0MqM/26mUG0mSFqk85mQ+p
/BUQUs6wXiLSAS56D7zqZCL4nFbpnyAjVqwjGaPLdVu4leY0HryxTa0I4xndQXh1
XcqAUi1tj5pHcfxr6yO3L+k06q9//LgI1U2Y0p9ku434KtHgSqa4jolSNOo5RFIO
eBbOUsTvpakocEv/WpfaNjwvY+UOVY860BbnynaAQkLieMotdjkRoKPUT67nL/aI
CSpLeD21bk8OhGrNcmhspgtpFlXgm90DvgChEh1lj8zM+lfSAZ7jJgX8R3NvHnxa
ET0+Fj34BGkx9D/C9QWDVwn6MgK1We6y9DX2XohfjDxa3BJZI0MXXQDa0XS3dkrf
qFDI2Tpj/OaR0zCu57jctbqbyQ4FgPFwVXnVZtGbA+R+E0RJFbpXPes/k1yHreZx
favwGEWb8NvUnEXWrJ98dp9/gA11XecQ31qJaUUWML/6XlluoaKhXMzc6GpLavO4
1Ok86olHXuNr+2VMNCEabGtziRWT746ceCKdlPwWoXqvTVXPIywHqaFrxpwmH09X
c4HdPmq6uOuDMaz7dxZliYJ3WTKZborpE4WbDT11x0jNKEWW2scDZwwTj7SBaRPI
+Sy/mGTeYrFfY5AtyZCd8hTYCG8Gx6rvAvIs2F7Gwij1fBDb8mDj6oOYTdtvapc5
8oVQ4k+9feLvh+AkcSWI36a1o0Zup6VV0rSNJaUwq5Jv7bUFRWZZG7sIVohZH/FW
bqfdd82lId+Nf7eH54namrs5LFABF30dfAExnA9Ijh1Jn5KOg05cRkHwhEjkOBLV
/mQvTciKCzTVp7y5MrygUpVNiNveaSutemdz9MamOKZYt2RsDurYd1ZUWx+z25Hj
esEq8l8E4I+sFxkIqa4IEcP52Yl3KcTqXUSOlaNjNEgqYb/kAtQoksH57MZgBno/
38y69joSLdnvdqrxDkN2efryrwPWVbsi0LRevYS4Zpov1UWNHonJC67f5zLHfMbR
YdMMfhqbSBE/l5RExkb3iIg8RN9X56r8Wg+lp4iq3GSUo3fTHby1cdk5Bc8wi7Hj
GMLepxqi4TdKy6Us3mk72eexbQHrIllsYhZafzNxO1ilimRBTiIv2W7ZUTNAfAit
J3yKyEasnOWmM7wgjcs0c5hpr45WqqrTiTptAiAU/VqIhDn5AUGiTi/u/tzrK1iX
xo2iGE4lVzviP7ADJOvIVJd7MP99NLCwDK5lFaztuU9DBdI1cL/p5aV5f6BR1fZr
XjRx0WgwkNHF6GTOT0mkWt9LnfJ11jjHp+hdWD7XrsiNqGYgOhlXcbFhjgQOfkpn
4eqOy7l6uv3N1KuqMigsQcZeaKS5OWzFXgzh8QIgmxq/iKNkavCTY9MqbzAuD5CX
1vsc6cAsIy1zO07kgRcDh7gmN+d+0yt65lDis2llGC5Uj5c/b17tGf13qC7nZNLF
GDNY0qb3Dzk1j/adSQn2wk/o/HZLqZUfxp9G5AXYPbsHsldRWv1ep4Ru6c3XlCiR
fBPHWCJNiXAUXY5pDWuuEIvDyxEO+PKMHIHgfBK4UvLOud2DkD8aVaj6h1y3yk74
DnuP3Uq0+jrxrurBST93q90eeOLai9S01Subegv12+qqpohRxADbZpdbvGvo5fxO
up5awpGa0t8b3DxkF0LMxEUvyjQhTVcZBMKUt5DyA7LgZUnh2tacr6T/3+Ii4ySL
k8atWzlRNkrCpIyrJy9+0dxE7Yceh7JJb44IR9qf8KlUtVEBW2Xm/3hUep7rBhIz
jgtYMsuIZhuEwTvieuSUOVxZIJwUID5+J860aXMB/ucM7bMgssZojBLQ+D+bqccE
YrFd3VzVDO+i4keRRdPnpEcJJLVwwRFStFUmwT3JAfJTa2TAjMj3LeAg9H73efxh
2Cu6Fl076sARVH4QUlq5fLuriWmTId16D6yhiZcV85/26TkbDc3xaidoHV8JwkkW
21FTh8z11BWKlvLUbyKwqsCbRRcBjXtLBPfiHpOl0wJbD6IHnLd16dPbmY2D1b0E
p9GRejXkaL94fWFdQoyRavv9N4ULURjKWs2pC6Clkpk89wjxDihjKdxXAvQ0znEp
kHGpSmP6NwM/QwcOGN3pxdivKct7QVI7aTs7z/8zHQSKvTqpQae5ELLK7CeNreU5
KqFpmbOGvO3A1TPcAUZyKgbeOY4RzGGSwk0gg8tWayqdDTL+CcusnjTjy88YGv+c
Hwq3rEmPklfSse9o2IiJ5tEMxpE4dGhQTU6tBGjrMUkzAxdn0I0V/YAsqq1gPGEH
9Cdf51JQfBiT8loyl4QaGTcFe6WCXQwPW/lUHkmDhcqD7+oP02LNzYXe4iU8Srd9
6AVcPnNJ6NYq3ng2pFP4ZkPfqjttiuOvPNK17vVPulczgnEUWBrXXd3OPdrLLF+v
We/8nHOwQrUe9QYIE9IswBLY4RKMn+RoCFDjLQFpxMfmO2HhfM47wlT5138Kq+rL
dmmuOjepR7teHEBNVdP93jN2AqUW2Bdy8bUEayKvdzfDoID2JjcJLSgJWu+snrPy
HFVPICguqhKhMHbxcZzSWh+3ugE8cwEgDSijRT0cqzO8wljiqVb2D/1RMzaXQ1Vj
JzlAXOEhYqdieHhvYI3p7d7NIctQ0DAQUB4HB3M08k0p3sMiKqpge7LgZCHoBc1V
pnPV4/d/rx9NzAZxiR90fhlBA4uvofbzpnpyrWox+CggDK/WAgfZrd2EpR34tunN
sqGr3s69AJ34c4kfg3KE4rLVV961jvBtkveyoUIkx7eXsVHCYd8moCOaDS5VgX8L
QxffQJRVOrPy/mTGRuraBV7TgAHLxQIMt7i0BSC+94oEuRgYb0Yggcrl/OP4955P
YEvAYBHVVFFPQmjQVp7HHwF0Bhcio+uqohioKogFAQqlP6/wg1xUxg48L1YNblyn
RBJDbH8UooZ3nXfnHkoGdce83yGa8wQCzCMmqpAfK3VTDs7XBi1XmJYTU7FY9W0u
kZn2J0uHfPJlkGDLmuvpsT9mZfAzXLF/fRd9LJeZ2noGfc7zMS5BKnlhTFspaFeu
53C86O294DatVPCI3EotKM0O7RyrZw4rAedJedv8uhTz+7ypeYkP5QWZ8vDR8Bwi
owdWJvL5tayJKtU4ZDvow3TSMg6uP+Fogo8QKhmz0wrgsSrsd0UPISQtfaSqtHAg
Srzz1oM1fwgzPAWrZ4Q+mx9KT/11cNjEZwL5UoVX2XJZUCTYFQSb9o9vWEw4Ltr4
jBiNeyIAC001+4SV1hFhUKJURoHUz7mD7Ia5qA2/BgWYffRAoOo6KQD8VQiTld7q
as4LHWEOMRYN0HyfeHBZBz5Ka/wsjP6Bke2Vh1xk2x++L2qKPAUoOmLF22cW47O5
Mqi/ppNnDCGw9yL9pk3P0/y9pyMSjFuoHv/NE9Ywme8/z/pXhmCzRWNyhhpDJ5Nt
/gyshV/EKqocEhQv0roUMqpdh+tLMgq2ZK7epUdDJ/qBWwpC8+Oq5Sfba0WGR9DZ
VIcepKdxKfsmDGeiIRgvZzpNP5v86y+Mg+dXn/jtxhTOphsxFMI/n8MKNLRe9dja
01Ioak1XgFTTFm+iRttCMzylvusdYHk+CI989KhUnBOEqXdBCslOf6IyUvsMkiyV
/Iiuelpa684hgE99V2e7KOf9nBpObAk5DJQwUeI3a3JT9HMz/EajVkqbAtlMj/77
dbAmlrQiLgFu8izX3I5FPj6kXKdk+mDQ0bnmr5ZqEWfytca1Dcei52tNr2678bod
oGKuRRs0qgaY4QJJHL4FtbR54easb6PbLwfWHWa8ZBNYH2Wb117JBlMshe/h4nU+
gVg0aGYh+wF9oR5r3ynLrKGojZLEQzhf4yiDTxE2oWzOTPZ8OtrpUrLfCqnWTaO/
qJJc39lYOyxsIxJ5U5aTxpdjrgdvRSpes/7Ab4LjF0CUb3Ke0ZsGDrcoX299M9ND
p5dGMVQ8xIyEO65cNHINUdCgmvOC5MSoZyxEGVU4cuoKJqB9ui/jG7veAylwneyj
Ag8nnAnyvRLWwwnXY3ZSfTiUaZ4OplRACWAra5KSzl+XBY/z3SiTXxN2MdYme9Z4
d9SsVmys2UrO3JKOzeME7uNLdiQlu6S1UxXh2Zf+csnkqbXzCn1vJ3zKt1SrqGiM
5DPtlmrhaxdrMdnVt5u/IcV1aaSXu/hTh7q/a5AixmoIIA3/N0rEWDHxw4SZzu6z
osSLksZ14kAsEqviokcDBNs0pNKfD867jDUA11O9Luq+EVZLISZ554kYABtEz5qR
B7g2R5BQR6t3Fmra+C2PTeTMfFBe2vWcpUtZJCh98TFHLtS7wKU1nh6JnC0olsh7
sye8b8XhfTL6djCBZANZ1XZUBQ+m6wHUg9EZ7TxlKPozYsxUHbiOoZqlW1EZjCpJ
7G5X6td/FJdAdsq5hiHXl555GSJyDiKV01745Ky2PSpUGsp0A2wVZ2col3IPmfWk
03XhBTyLdaiNmm0FxpzH7FzHBvtBx1wi+/icnXNh4jpjJi8C7cBHPRwvUWxaSoPb
prMWcEJc5wjHEEGijd2fVea+RGjM0ZKfFx7QKzx1H7bYqPCvVJkyJlTH+u9mA+ah
MXaVEv+1Kc6wqemlTBi8nszae6rD/56Tp72/wdlD3MU1xbDWwuMFpmqk0Usk8qI2
EXUWSVSs0b+yfTFvO2Ux4o+JRConrqiYPSONX8UgDrg4P3x39TdqhlKo6K+3J6JG
rBI0ru96/2acX+6VURhN+W4bBqeqS+V5SkVZQxfZAR7cyCQUMESMzHC+2c18kWcq
0y6m5AvalaEFZn/WcybkA3UcVPkS0OsKCGqanyHlZM35vuARq8zYIBI5t4tlQA14
HefK+Icp1jpbqNqL/DZNyKfIg7xP0d/c0ZYyI44yicijxhA74Hn5AnE5P9wp7znn
a6PoMz85BqXbqsv5vVD4cbwnM3AyyF35KFg1kV4UsNsYws9ve5KmNpbPNtyeBSaB
6fIG94aMXe3EQWluTlH/t5DvgDI5uDqP7q2B3MQutsG3HgdKYbvHQsmrx1zfPM80
7Oj6hm1OgDRP7MnlchbCvWlDssyRyAWjhtqBaKxVltnFRvea0dveC99FsQH/h7aX
uBEKOgIfh/gWN+JsgYwuO/sXKNf3o9uE0wCJ9tX2iNqRiIQMgNeGBlqooVDdIk9C
B5XmY+v6BIITsjXBm456JDXLpbWZcQtllxFdlrvDArVH1F0CBlQH4bk7HGA/U3sI
0znlIHG9TpQdnUNJVvV4BoMPCIDH5t4UcMcKoZgOE9IYJUUV5Shd3waqCZ2ZkT/2
U4bizt+UZGqNPpWTMFSLalaYzNIJkliy19OTZZZ4IDVCNOPY3x3sC/kUy9SGBFvd
pDM8anQiGLSPJgMmMmpdQlM9l8OeHLBgfW8x2IKXgGU3y2dXvmGt59enfCzdfG17
xNv5xxFq3Ggz1pd71uWFVJeABcd/Ro+67WjYc5eNiRh6gviHGz2Ysf7UiZ1D8Y1B
X8LE0HiSRm+oW4EpP+M85nwLLhjCYXZQbW1HfG68Qg3NzfCxuLfoLIVnmD96nwk3
yZJUEiI+UnGnlPDMikMZ2Ve2LXeD4riaaxDdDbyAA3kK1EYKWHTXKLBVJ9IVRcxH
JL3G0qflMU7TEoIAHp+/LdCNeAf3vUt6oZfcd6A+IiYO1/InFTon+k9qOosGfw+R
YgmUmnriIBHOBjF22NCmLhpabdtbVDT8hS0pESuanHyJaiR4s08nTZGmNPv+qdYy
mEYKrkmyHiFhhOurY9ZjYunU2q/YMx373liBETxmDm1m2OxQSEBMeH3uOBFbp+Mm
lmubXUdZqiQP7vGfmJmZy7KjhHK6HYeqlWFxzvMXIDSNwpitF4JSBTY/JHUxvHKA
gs6pV2WFRe2C798fE4X4/WaA34JM4XPsHAHS4btVcV0mAVPlM7dafN8+6jgKJsbo
yfA5fg8kV6iFIrA1PFebjLNoyZxBPBJRqM521Jzui164mvvc6p3ktG1PtMjiOijW
sjFTUFnGL1Ltm9Fj5GOaaygJeq+3gqLeVLRFFfQFqMjxTni1oBqlz2YleK3Lsd0t
7F/3PsEJg8KN4STFRjVqRw188Puq+xnXNp/VwU5uXjVoPBuC9gJ8f3nH5d1Twgha
NF5VPdwU6Q81Lada5+O6CzLGAKV6m02tgt1QbBqGgktZ6mFhTcw++901EGfgPgZd
JklN8mkDE8thNlobQ/yVQn9aAKjb+meEjDateNLeq1Hj74wKfc1c1A39pB2h728o
acIufGbzXPr1Q2lxzOKQMB4ACTyPvKjC2/VhQNzNIqDxoogouu1/uV/IGigx99L4
6Y5WlPYgFfbl9wbH/I3fDbhOizKzUuVJf2pq9j/BiQ4xJCctxWWpMr+wKEmswswf
ZP6ocdi6QYNbY/XJ52o75admYLTIdzjTTppQY9yaefuix/saKG7lxJXYZyG4kpho
SoxwpieCtc424wBIS/ogqZn0ctP54Mab0v51VbF1/F/cgYSLEzy/oF7fzJoOEnOo
/xe6OkscAEHMIKgPfcDTzF1RNSqROyiyRRl2sJXJ7GikMoP7oPjQ9+feomfzAy3t
7OurfhgrnCDbLyHsgIRQBSKOlOAn8yEvIliROdQKkQV1MJ1NM1RNkU4pwpUeNLCm
ydXaaSXKNrzIh1R2DjfztUt6gLbtvzAsWh7nuG1zQaj1Flvy9inlPBgA2AAMz9ym
I9lj8+/pv0JIa8XM7Z35SasoVZpk/TDc28XdiubaN35Z1FDR0uU5O6/ki/Ma5WTh
jAejCC+3CmGh6AKEuA51qkDaoPkvQiV3G4kcGKVKML/f/GhMIhDpbBTBoI0tK4C4
IbJALBkiOCYRbc0QirHnDA5g6SIO+EbSP5XRQoMyC6SS9FNjDOowcf0byQTgVLuF
lBFxdzcjdxHRVxJYQsGnGIBn6Ptj2ba3RS5XX8Bw1OMhfpRsxDat7s+9eMwNadqv
vCUDmjY/Jj6KMp0Jj00jtKDzyRftty0/bE8IhPXVzpfz250DCyqS8blo/YgHQxMK
ZVCbdWMz4lZwl/2HwpgX69ck6uvPpRNjNzWrA5ixWvUebOL9cT4mRKKC3AppXiEC
fuVEklbhMDseKeeiApgdT4/hT2bbEWyektzUZXxjZW3DopP36qqfSLN50qk0Esy8
Ssr0UfIYS9nRoN/VVZNavJlC4iV+74G7ZJdqjPr0v8vv//1mWFHFLQDs87F9B/7p
+BtBSpxy2ztZv/9VpzBSXB2Aen2+7KYr3zPIxl2THQevRDI0CG0uOy3AQ9pMTuqH
lI/fJEfg5QNFZShnTnfdlMsSnrHVajP+6Gr/zeNnSTGex4o8jKbdM1SbMu6Qo5QQ
Ew15meOdIIKht4Ju2uWIGu7jqAhcNsb3NxhTlvsNYMECcFpGw69zMa7bHHEvrmLU
2pU984RGoFRrAsq43RAVvs/8EzWOJraaIQcLJP1WT4EYkCnaLqF2b7OYNRp31nF6
8/N4tXRGXvzgw/vJ+KSvmj/T7z05v021n5yXQ4fZ9MgknqZ0OhXV3zrSimElEA12
zYBudbaRyizj2xpuurQalWlcUVrHuKlcaxgIEZLGXrOFdw4h0qX2vx/7LQJ7g3lq
Lmaux56iCY1KnGfiw5MPp/wVm76/u3Uam4Zm3zbyd+ehKR2oHRjFWzb8r4aOei61
h/tOG6tmfWf4P9WqHBWCSmYATnrcSw0AvIOcf6k3byuOwgvYHXKPqQfT03d3o0Ir
9NOf9hP8lA5I6TtOqES9V3WY9Ge8f4v0ppPuoHrHZpsiS/0el9dvjy4vzZQl5Q3S
LXyvbU9Egb5Vaotll8pAZWc7zPJvGNP7qoiEakZSeSsWfh37GohIUFkfX2ov98Lq
7TzuxGBCR2JvU/tgjrgiXimHKoMfTf47O20GXpLPM5aMEai3Z9zjdG8NYq9wEDLk
gwNkGSF2VyxHQr+80ivPPFdR+CURNFLPLd4Y4yFEUiMIvcl/AY9nNeFYJF3tdBdd
TpPF2jlhIMXBspT64hBTtT6xsg4stQ/wau2gXovO559cAxN9j8UUJWkDVvaKaAR9
o+VynWcqZ54akZnTJpteYz2Jsjxpn52X+mL857Iyguy5rZhryYBs1yAUGziLzVah
inaUqr6tlz4TdhpX9aPHjasnx6BBUhNFYh4UNHjQorCF5JMW3KsI9PHkF9jeJCFH
1RPTPr0oT7jy/Yshw9twojy5kwRxVO6vezq07gSs1MrQ7jiPk6rwDrevwmmNXdMR
R/bm4mVuig18JH3UY/ynurZ9FN31NFnLKWpbHtL5aTb55jmdQtZhJ31EWJWdJAh6
vYw0OLZPZRECSbxtucyeyYHjp2J4wRPY6NoO8mPhKsoTZ9fmam64aH0FycVfOhEv
/Qek7nQZJ/viq4GT2ijzygsEEc5c1qufvkjN9L3oB7nIy0lA/RpyKpnxxH9y0Thn
bCy5MB2aALwntWd9ZDhSjA5GCdVDpml7N/eHjothUNJBJywDFaXJXwPwDqdbEZws
ACE3OqC/kDBS61DqoE9LKYoZUkLeE3g148BTERnbzcsocqwJEhRchHV3Ar4sJEHs
niyxhD4eCa5wtLCnq8NTAakN8CdSWcZ+2j7TQaRzKVIA34GljMTkkJT6Oe4AlD4M
EWKb5ZZinGgk3SafGuxZqAfPa40AHkY8tOFuiSAXnNvd9DF6NOmT7vYwNahdU22u
5Nv/ZjpxeqjYs4rnObP5Jktzsu+2/mrH4OMKKPh9Y/8nmNU3pD7Lbcsn/ziWY6XS
CuvlxqfKSTQO9ZtW1CbWEGOU+kOsxd8K59f1Y2VmB9aBPCrkueHCkB3XPwFacoT7
vCeSu/HfXrqz6RvR5CZ3YbUa4O2GK09j4gpQd/0zMeaCHm9TvE9wqx9vpKFhl901
OY60abzDmBCJ6TJOurUNcHvzHVZsx6effdY/hE3XLIfU/H+MXM1pjVI3IaaHfGYK
yVG6bmaEkmMonHeDhYHHQAQzEaj2fs+xH60/55ZDn20Ss37g0XTOvlF/AxiI8WRw
Q44V5MvJu4TyNaZ2bE/0ElzFSZUxguNDsRG9vYa4XUnJFNC3vCEKQhEmqMK7XYon
C8kFKxHnzAYJ0Rh/TwvaHMrCOqeRVZfD9NSSaFU1ggbQys+teHlVdzr0xptEySsV
Zep0Ptg40EBaiDP9P4WLJqQu8KKAb53/aAWLqg+o2W9eCkmih84We6LU3Lorufj0
UdnNwSOOwVw1pChB+5WGi7Gxoa54fFhZO11dsrbBdrAe4hMpwG7vTkVgz8r2KIU0
qd68+P08yz6UC+qB0jJnjFTbLlzpYF/twy+372NgaS79X2yj4osRaaLpnKbOUDke
3e1INo6DAaucsVlbNmPH9nKnklh3LdxXe3qSb0xqOqCRuEXev4t8gtaFSnVWHj5k
X0FCZUiE1dV0X6beu4RPck2qJzF3s87OnR5Ht/cgTyOmNRu5Zr8UIU8+q7wTVGrE
lyAiRx4dniasVR9c5TbWr4oRUW8imOs0cifCh0Ey9HPxWvxdbUzKp5SbRh0FtrEe
XBfscqFxYwGWEtFeLsuQA5BS/m+4ZKg2uZG+vGv3NzR6tK67NmJnD/PAOdhRhZYj
8YWgop69msoBXY3GZ1KFpzYnUAkXBDpxAvTfgSUMx7irNm4w8pCa7LxNcZn3yqJ7
1hJhpNiu8BokmfjpOd5xr8w21kOvGMJxHD0Dyd2Zv8eZMBX1aqjgcglc2Y9Li2lm
1mfYIDJeB8s93hUkSDj9ZMI/wQUguPs/rprOyG8xxZqCoKXP0RAvg29FtSoMeLim
yUHRCnA6n0Q9+ucGioWHt95PYlV/oaJju0SrS3xurBrxN2OKeMAipXyuD+Tb6JZW
SxGiJGlT889P/OQ4qdTlY0Td7DUgSculQ1D2Jwon0cJn9fIEBDOBoDYCjKMNu0Ig
TiHgAhrB49G41N7QXhYY1mc0JVANpHpr5jV5rUSjfKKo+/38xdvITUq51xmeV+J/
LV2IYs7w+U0ljcI+o41JDnqqOaL/5Dpmys2+ruVwzu8HlO8iqmjgBjK162kK/zJp
nCKNj9iymKRS5AlGFipKzJ5Y5HKZKckwPaRanF1bUsEhdooymiewDLFHGP1QVN8H
GV8/87PrLpSD6G8HkHBEBp3H9mujBPf8vv00ocRbRuGOwdSdmiwpCS7+dWM1ltiI
eS/h/T78YXeXd3gJeXeaje7Rvss0dAY3T03GwYqwK+XZDBt6IEa9iYBQB/Ibwq8j
5XwIhfmBLZjmB0WFrW/b4giMstwqDeK+TmV/DsGqebsnuzBWA6fYBGwqLy2YRV1p
HvrjgGy4rfxBqWwTt+qQhU3exNjFdr6mF+7NA9c6qG7KJgW4TR/MxB13T+f7AYm5
FWljySriu6NJ7rt2ULNhabc4dvygowwdNUX8+7udGsSAJmGSD0FMNx3sI7mQTplz
fF2Iq6ixZ+2LuahN7pYd88GrRyO/bVDGbcxqlLX6rE7wydl0IKWGCfdde8uQ4jlV
BYjRK/NoI+/uCL/b1pAudd1g7Ldy57/CjgIymKaLYkh4WlBEVNqYecGHZnRveLaW
ABmD4khpinLTizkjS0BFPlxwOKHTwrI/VF/rzfMqH4KIHpneii1MgjN4aTF9vVni
iuXUOwxxbbQ8PeyROb/3vHrkPgShMms1Sfrp4uliRwRu818cdMbUHSuGJo6hV//j
G4xJR12WeUVVRus45wb+2NwMucr5/t4XCLiqy4x8lE3tjqhacGpxG9agNlOmfuNm
+kAupEZc6S/6/XwhP6KKlshsk/Ntn8htiT/5etPN5hZeCncP3DgGHrzYatvdtBZc
1Q5Ma9iUT9usB2uI+VDtqrLpZRSeQzVpzoJXy8E/WuPoTIOe93Jvtp0NmkjVyuRP
+LABHo215CIYayOHhTg1curZWY6L1LHbsHrcl8iEnC2+Kg3gU7ey6QiNbQxbpLoW
ozXK+lRkpDlcykKFVa6OIHGMVKvdn9A7cddzgK4MK5aj9O1/F3vln+RL1dHgNCXh
/bSpIrSagx/OzMcjgtpG3/D0q+VHdWZYlh/t7Iwc40Klwx4hHK2sDKbtNhD2vY7U
CjnpfAa0fpPScALlCox/gQLK/ltEzt4uZICaKT9jp/m93i+xQGJxOtjhUWGQLnJM
3xW4Qle9YsfkBzANlFT1ohJUeSvrxUkV620WlVih2e3+UpY3Ar2w9uE7eA0OF4qr
nOQ/7sB9rzOPLdSKz5sBRQ6CRBwJIvbhToM6OqZ7crSPP1CY0sljxcOHdc5HeZ/z
b+Ko0Vnp2d6G16C52FhysU1ZbcRhVNr4tZa/kHmKS15GKZXjYSVTGeH3zUY1hvtp
2Ui0IfWsAly4WWfgrEXJX10FH46jOgQH+GNu8RBKmXWDvptKkwJ/u8cfeJyoVjuz
tc/28qeX85caqbN/95fH6W5A/TXoiMcKFTBL5sD+KUEQyq3ov87YLxKOIhY2YNpJ
X+ULFMgFKh2aL/1tubJy5Dc0FK5VS6l2rXc0/S9wJMEVtKi2zT3TmI4UW2Rm1P8i
PAp3M1tUltG/O4lf834hV219qf3rY8DV68psbES8If4wtAC1n7ysnv9ZGbpTfrnQ
+nzLFJJeBG0bYMBUT5zAVr+hZD1vfSVeTLF4LuU2wk8sn2Q9hxutHM2OwOUSkAM5
gzIZM5lAa6b0lYxXZmrI9KZUbSYj0RFAv2OUhUSIBFGWUCyYFS6fqxEamfblDNyq
rXUYzecsIpqvgOe1OB47FXvaRtMPpMFuKBlV2S3QvUFcLkII6a0QDEyEuIjlOTwf
6j3H5uotBaWsYZIEEGDPxAXp41Wr3hDsP+rHx0Tu9nMraaTjuqC/gj4lzO151dlg
y1dhs0rsWmhOvPyw8LJZ8TfrX+PTgUAMVCHxzTu17TeFxwnUkYirXvtIgZDi5Hgj
UE4IPadjioEt88GyMOVokf3zthb68rNI5vhAoo2xmkLcKzcLQCKU0s/UZgtNfiM0
+UlkWKYNvf/kJFkGhwEuDsCWQevWVBhypyH/wdeeZHk/yIJexo1SsFes+JiXeC7d
aqtUREQRU1JWBzfvG9FjgW8H4z/yFMClrySW2BHWYbcpCSWXgbjhYtiMYHtRJq18
WJC5QNLxGwvjeA/DlK1idwSmFMKnnmL7UCeMssIEmdOt0KJg4posnVPtO29UD5si
H0vyE5dTJA4OOeorvXbn0mLYsdYMTrTk+J5mmB4dhGwC7G7SwFe/6CXscYs8yge6
MetvTxZVcDjirUMk7D+039uzS/4M+iM+KvHAhQ3y5hXsgs+wx+F2N7lfM2+Nb53E
XidY+VxvlyL42x45xu3tkl7xpMD+iA2ny7ecHFkaEq+zpi7svj1OKg8X6n9fqUGq
cmUd6kXejjlGRu+CbSqDZr0JGvCogtMLc4Ztm6Pdk4J/UHmTXVU63tNXYUtfQODl
9pW7YqbbbnFbSlPimg4PcDqDX+Uc4OwLwqXuWcdbGcT1RwMsqsVL5rgAgpblsN0O
EPAT/mcjD8e0LjNKYZ2aNDTjKJXg7t2xmT7hSyDpWgL6G9iD8zy2Ww5sE1IdhtDc
64gxzIrm80vEAvvwMDvHu1MV6aM7j6m+Lj+AXwI/+PhhfkAPibwfibCYO3YdkJpG
YkbpXJN01Ck3ti14E2a+11PVdK8CgsMgtihRS1qLzD+niB+oeU3t0o9IDxcCjPg9
5/6vHzuii2GtqnvE1JN29zX88t/n4JhxpDtIhtdg4qul9/TOf+Wx3Gu4MpdJxaoE
+3Vjcj163TyWhgjjyzP7+jPSh/QqGHM9wJzHLGiwB5CUZy0or25W3HeeDAoh1YZ5
VAF8R+rXWCGU6nWZXoD1I12igg0UeDYgt+CkgqENTx27gIqINS2djENHLC37NDpT
proIhSVPJ6ksjoMecnk1sQekLlnOK5docVFkQin19iRv0udrVZtvSgLger9tjB+E
8znyqG/mzD8JAb75LkbUzGKcCt2rwMLCWGn6UJVhsiGq/55JoHZ/ymeymor4NlgT
jX9I1B+izq78rWSZeRkVpFH/nIuiolOA5tGlCtfHyUOEu825+kPGXpzfdsNmHnZO
TZq+kllMXnilmafDil/xu9MSf6LZ/EkfrSvBCz/Ad6v6L1fKUzVd+r/AwOvg5GFg
nn4USqFMoY/EGz8sCi3+jApt6+qfQqKhAn16yFADa8TLTo6xGGhJZ2E/+ld1qlA9
B197cX7Ve8PTrAE1uflWMFhSgzo7YR7D8N1yvlI/AyLqsijZ9bDqdX5d9wfD2Uoe
nE9k4gmvHUJgMtWBDc03mbAX6PacR2PAH4JrQphBN9UWL4tBXk0NjUd8JNy3zfoC
PnMUP4v5tNWnDtZhh57aM5jU3EcTCGRKdKdAH6G3RTRInsij5lk/qEEyqlRnlxsu
ojqfwAzT9QgkHDREUv4jmq/VZ70DVM2XNHYg2Y3UCQnaIlXgQoFNOIhvnWlwTgfr
ZZTCQA9dM7OpFqU+vYHylxV7PlPZRbU/+94dlFC7hxLqAmVHwGue1IMefiDouS4D
PTsnxRxg9HdTmlDDSp6clNVagUo224XBcaQic2PBlRxPg9IFmlQBk3y3g2L+d4+F
MpAKCgEgWCUhPOGcw8Rny9reJRvBMQcYwFdlVj6N3R3WNbq1vBNPsillCk4TdLJD
80TuDxFVVQZMxxG8tTLW0Wst49GVSacReHFHdL77PvYxL7exohy6pR7ND/VAMoyH
oLnzpIUBdx47CX2CCokvw9LiZjpFgvuBKClyq9LR4+rDSjavrShGyfo9+7ZnRj+4
yhvKIQCOfaimyQJyjRTUF9MHkDAv0+7dj5lp9hXELBqwIirMH5Hkq3o1EqHI1AkX
Bt6cX3W1LLjlQU8618FpjuT2fQ/33aH1LrLSAWa9LI9vyOLBtkaMae+c58TQ5av4
XCILhcxtEKCDDD5Poj/vEiDX4I5g4JhV5eVnoUYxavXq1/cvTF1uKg3fZjti150Z
8W+SF1HbCI9Knyxe5H1tr3wHHxWfYDvGtBSRDLR6COY+mIMy74eqZt5Z++4erRWN
x+zHpVLUshIdwyC9xRsAwPyA2kVPajeG5AvFEqlaaBMzjeQ1/1eoKVzgNYKBmiC1
LaVbV2AhwCBBmV6WG6rm45XNnMXS40uPD8bqXJDnzz1P/hsaZ+5hz0k1zVVyD8yq
fterK78gX7ijNujVt5jHOsnKLBYkVhEjipeqFn4aZhnX9cD++SMDQBkyxs8/4LAE
eEN7hGTQv05+vc8dq3w0UxTOCT6wCJ58gVAe5wHfIR4/HsyeLf9CdWN5Nj5WE3J6
g2c1qZ9AhArEL8zfdJhitytoniYZJ9sqdeMvEfUwblc8Vc62PAcDI58Y9J0NJTkj
YH2MjqqEKhDUviafFO7xAC3posiAzHXK8hncBZTEcDrD05JwD2BeIvDjSFd8VMKW
r8oXvUyLcffqxvKeHjwfzB7k/Ga+jdwgSLdj5wOe42+xCvi9eUizJI48KUOZqQk7
GskBoMISjF984fdCz/MJFDe9kUvNgJMAOmTLzOiD2NEM09eH7AW1T4/fLNONg6cl
9DobhfXs3cCfzSQSSBbDU+lJwGVN5CtylE79LpEqNtKTtaulNzxAts73U0G0NuTR
f6HYUid4wnz62jKu+8ii5WuQzwnmNSnbcW+IZQ/R35JlPpjOcj/u52+nW5MUlHK2
vjYRNVKkJ4HJshJTEVet/lU4m/Po0clBMFJAoN491yGr5IkH4oWA3rBhA8d6NB1k
YtnZAv6/20qOt8yeV2KCE3KyNZ5MYqSq8dvjMmmhlX9bCaP1QJMom3o4ycRuKKmv
/pS20hrDWWRHZ7mrwt/rzK+SicLfSiLgAZigpuIhs6gx8Va1pdY4+EvaIXSo0b2s
BeGaCTIB1bxFofCYPxemIrNWC7PeODjm7c00S/FLE+VFXQOFnjjWoOgnqaQIqf7u
e+K7GF2pUlsY5xe91zVC42iP8LsQl8M/CpKKthWECfEy3zDsLfh7zUlgLF7ct1Fp
noy8XgryycWvvJ/oEpVP190MHKhP69MRJvC/7vnDugGxp9rCsN4697H1mSmAyTdP
pbE/5lqQhdo1iHfZshnDpsCSP68bf4Eh/2+2yl61RhxAApybpEzQHO0DX7HUA6fM
j3RnKuMjo4jxuXElcx/lGJRyWyoxoaZDCnbsYcezsmHsaBBiStBaBgNgQzxEWTAj
6emA/61gxd2SeE3gynNNEAx+FF31K1W9Z/1orZNtU6XJ5jGaugllL6u0Tn2wGWMr
QFL007rUy65XvY9zT1mqJJ72tbT5IuBC8QpvolLRWNSZwgqQ1Zunbwdq1RhGc4Tz
TJd6MKes1cD363dIt5CrwoWX7bbk+dUcnpjcecrI3U1tpoBCxVQWU1yZZjQlKs+V
lNnUe+dKR0xnV2T7e0aBTACRoZ+m+egoNh9numpKaUDbSb1fpFbfqvqqBFhejFtQ
vACt1H5bDH1xvxKHYSemWe/3ed4attKQHWqn3V/fDJOBVMcfb1pcZceIZCuiF/JT
BDCcX2kYPrQs20Msa0NvT81chQr2BN/D+oz6bNsSHDYPA8g+twRnQSKf0s+DcrxB
5n4fXST/lRhLrqeoMyGuh2zBYYhm2oS+TLCDDNwVi+yK96LqEhHMgfqjSWEN7Paq
qyrv2JzlSyIymcvvAPrisn8222iXDlFagYU7wP+onKfIhWZiEWO1h3V+angPHrUd
R8C1d8yhexy/7thTf7SHSpx2izeFWghiv5gAXTzUfaV+viJJ9ps7DZEqmP9tdjhm
QuHWBXL5C1pAjmo9cR4iccseehoI8BT/3CQllg+QZTD76NOhO70Kc9UpLtr/P7jI
LPc6qWd6srS6wr58CmPvyi+r1qEItY4KKIH385b+65F+CalMPzcpk2VXqIcLfsAW
fPl8ulyHNXXbY6CmQy8K2MEIdEe5sOPQuPNruJ0LSKhqoY5ijNxdlrzD3G9WCFmc
FOxl00IJDRXr1zFiuCg4OxmvsWNilNERAHeJbZs+rDYcqEVGl9BqSGnh6+dkhUiI
bub/tREGmBjp6Z4V0C4PL+zgJt1nbXVRjUUEslM3jAXLNQuhtJIwLFXfG8jVxCMv
EMxcRV++dB9BD1E4fAi8YuUT0jdEOypd4tt2uLGZPriy3wZDs/bdvRc5YGd6Q/QD
y0y2hxMgJDXPnAqW54ndm46BSfF/RW2DZb5Bna2Ht29UTWXUMqqLK5xMy6qMMaEl
t9irHlA18sLlxlMqH79VuvEVJf/MbuqJ4KQmo4VioImDcYOPTaPMW4IFZAgtV+nL
YKSh0HFVK1V1lqF0sJrRAIgeotlBuf8I8c+fWLrNA3ZmQCjX2V4atzosZjn/KuTt
q0oNihbKGOFrlvS6JV/E7p6t+xrhVi5W32RDQl8tqJpSqFG4ibc+NC6DVnsWf0R0
0NcnX4SohRV0Ne7DtmHav14HOV04iNVhfyvnwz09e58FIyqp9xu8YaAV0M6fboXx
5SU+m109yZe/T/RV76Ixo3sRAQ2ZQOCWU5qN/rOyrCQpHUO5AKXT9LtS1WyfFX6r
OC6V55tnNZgLNzH0+GtVNCWM9Enev69TSZMG9ivaiF04DmWJdfEFYfb8XctBBrOh
e9l8yB0pb+KllpUPtiTz0p3VULQbNsZRNrBKvbuZsLzf8CbZiHr5TASQ8leUtTze
givK/N64YL7OgcOiCglOj7U76k8O/6UFaUMbR1X4aFtRMpLy0ggjRom3r+2kD10b
RxISlbcRlk7Kzj+MAS1Nw5BpM0xez4Lwh8+F6gt/Hjf0NBTvaUP/ff1l6cF8LmHE
I4011bveeFub9fQG9qq7Q7hcmtx4cO1js5qyziudY/RJErLqwqVPNRwMltV/EGYC
oYYBfofcsalitffxDsuauxfCs/yvtIVm+495lorogIDmdPm51QdsaTY3ARoA2P37
3Ln94zc0SrcDIA0RDTB0TI5jnxKas/zrRMIFKBXVnj3NkNcPq1q4/7Yss7gqhE5b
GYdRvSqFbLdUW5Q3odiflBNvuDpsJrDi2izVCafQcEI+ON3Ij59y2548MOU7Os3z
KngMZH8D6jIonEhgI7dRgyPJyRYAL8k70qcsVSCyf15miKOZ/cPRhGImVMtzEK2h
rRuIKKosaxo1gKSbfncZAyn8ZSUAg2vqb44WXlMze/Eqhg+CyLjrtfpJUe549/pl
cb07Sev+8kQjmaf0aZIE6kKlj0WmONAFOcCblgjXZD4iTGmgeyloVImibJw/m2OT
mjZNPTWeDwpxvPX+WWN/QsDmgI5zmeO/digef2pVM6dvYx6aovRzkW6Mgpg97kHe
nmkMky8iUaupUG/8r+g+QzW810dnRr4/FQhOjTBcYY60ffsCXrIB2Jy25au3v2DV
pCjB/UWwPQde5x4SZqxRE4YpE+I2ikkW5BcJ8dYiFZuyPniC5LqG2CR4uxgRPuLb
D877OljulhymJLjkNgsOZrGoNbmoeMPL/jnSuAY9XhXd5LZWB7WZy0sIqmXn58k1
hxR6vLvlcmFtPJz9I5lRF8OZBxpJSL1oDfCpC+IbucAafQXgIGNmnUl5cUkhDv6d
q169xvUENgr1IL80s3Ql7stcwzbXl9109V7tQwSM/gmaooZvWF+mABXaaEuwLZFd
VK2gkgvzLcNcVCKRHSOfjnsTCEzTSMiU4GujsWDpaam7vJWJ4kyBXyyS55c0BS3l
uL2U0QDcQrSimNEmnBNs21JVphe3QNGgGew/MF1WVDbHiiA6ntRo10xPkclzE+0+
3wocsAc8zXJ6zbLEYXpbcoB8zjllu8BAdHhTyaZd/IOE1nqeCbFpeSi9vSo70+6c
iuKPa/OWGdmuQLk7RLhj97f3Re0zw/CUQTuoqZ1yaFzL0eh2o1IxGVcpwGsIzWdl
e26L1xHzoBkgTtVduDDoDaTwDm8VoJOW2RAfBnFkMnzy3vAouafQf3OQhhk8Hozn
sopy9x4oxeogE4pMo98wHAKk+/E/YeZJQ/ZQy0Siko+77jAU3DKA6pw22w9D78Pv
kDuC8Lx+E1eXvR4M2kIPuuPqbohMwPfMaY77wIG+pTqgv9UnGLifX+7wzT9bh0Ct
TaqqaHchBxu/5mBt9kv1yiQCQGRnLG11YzyHWOi0n29DhBnM5klOEvY2Tc4A/F/O
PYTq1S5eesv8aFI3SbrwlarojbKK2mCKHGxFIfMPiu58uTifHYIop/WfrRFMVZyF
bvbyYkwa2DW2xixh5qLqbSSv3S839gifFoPdVx0xrTSKhlD4QbvewFlCE/nBZY4h
gDHyHGUXZgatZH0+WNJH1qvz/4TkQq1MknG8fIhDLb7wYN2xBwqn63x8+O6vmu6O
gyo9BX1E2ojhABIMMDPB0WrVls5cOgFgFiOJt++FydlqncG9pZrqgMfzAr5rHHxf
UAsfnPLCc7NTU3Q7q8kNk4uipN3rBZ2+IA4diCyonp+LFbi2TG2AMgqUNnaCVXFy
QoVRQd0xnAxROKmwjK7O7ApUzF5kd9Z64uro6VEzQpT7SDYDMKGq7ar9i2FornHQ
thzA8M0SxOp6i9tcUkOohWu8iyN0hfkTbekvbAvQ0qbVNM7GvCsov8XhGcxvwbIL
caXBKYaw1GUbEUlAhBwB/YdD3+FF/7Wze8JwUL4vpGm1S0GAwNQR2u6VeodkNss/
T/r1BepUyrfLwNS9GXinPLf/4S+C0K9cTT6RjRAA/avim/Q9/I3sD9EB51LuWQ01
CqWU8/UCESp4aVuDbodMV1C5Qky5A2nFBmwJNfcawwUt3eHe+ZARcfJLwaeoS3IC
Et21TiFObZbObUQztoTNN6aiBmnb/znlnzhjWHNczERfIvzzdF5gOFYqElFAkQkG
QVOwARpkxP/8DQ0tOMEDljmL7VIrktz67lAuMC5TRqUWT9Y3a4jn0f2z5lyCwlvI
sGg8Yc8k39ROT0YLwPd2euDu+DR42LdFRWCGB01tF9jhrNG5n7hDuP2AXjCl8/fK
+Ei1167PM/leskvqqsaqgeB8wEQT5B6LyVEJNFGK2U50KozhmGqwGQGlsy9UgyeN
8Qh0GEHj1AjF76RSPVPcFIkwAgANq7R49V4QQt8Suu3rM1H//hPfOIJbt0zzOQ62
hxglG0MAgRInc8gAJ0fVU5wxEMYmfm13NpL62Ili8dClAkUW9Fcz6T62MnK1v/ab
2vW31DHKZES0gM1+8DpMKOQGz0m8duV1/aP2EgfEAFijnkMvmUDD6S9bCVCSsMXF
GrinQU+gkp5xBPmSPeeJC0uuikD+OkHzgs9ACOnsdhWi5n/m3OLa9h/GPZAbAGDN
8P5RJZE2rRayO7J53692tIc9wiRFp0jO5k7+PestHNBudVK0Z7UNe+YvzAZLkGY5
UsCjsm0hkQOgXzbmP/K7RKkTkAwtRBkUM54j2HzyKgutkCKoWjWtxNYudDnoX4LE
zUfb0OFglW26mwG4t59yO0FfoXIw8ny1kdOIZ1TC2sXkTaOHMxchil6Us0BADwwj
+gMgd6nWTStU3DBRI5Nbrtc5Lb2euiSkjOjUUBkzNYIaUrDC4hwEPXbE9aQOPWOD
C59jdzjeG3c0jojQLTsCFRwfaNAGDdFVf6irwW9k6iZp0CyIMjCogCmQO2W8HRWY
XHW6K/mf0BMUJ2Vq52spgwg1DeRFhvI2gF01BCpHe4tJIv2GROikNubMczA/xlYT
LqL1ApP7wFNwsW867G6Xl8lvz/GctTsRgJ55mthv3OZccHrbOiYxUBZTfP1ACdi3
WF82zJVgYFtZyeyMZ0RLcLinvJk3MyPBsXMx6Ew59NOBq7RHu02YGho6oK+mtu/R
weu4v9aiyMj7/6ludwqbSk4i3NYsuSrVL7NYNRH4gSKD8FLqI0YTOtMu3GfM2EiO
LHAtpHkSY6nKapyJXzW2b1McodkK1gb8VdfdMTlRgOmdh8bQqVkmc+7DuiKcnjkV
pFL0M183M+Yi2cWQ0fq44dZ869x86Yb24i2YfZsABZgkMy343L0BKEKAkqmhrSD+
FS9UQWgF7mqJodbLuOEgZXofb8styacNdq2gwhO5QRBL5glesq+l2dDpTeDU0vIj
Oaw+6o9vOJfh9hy+2+sBPB/inQ0y3re6KzfnLifwRj0+KjQodCnCgQezZkGxbQis
pBzUGc0EkuF6jxK07uZweibdDMA0MDJvGWu4Ph2gCkixTUx9kfetCqbuHvZOJy0h
5rJNgVI829/tSx1D4luOJft/YJv13g3dKqo17HrgG4qxFIkew1pBULNONOskhiCQ
Eqanm6UjjKWWPoLuzdm1mHDq1+RwkYtf7jaUycBuY4X6Q8ZZpqUlw+0Gl2F1XwNb
sxeuOIPxWWDrfQe0Ohnmlfxen7cA5HHdHnKCqHGinKQsTuJaZZhQyh77+Y6g/wuy
Av5DAF3CIjFV0LZk/8/H9bZYOhNJptVAIN02DSrzfc4zsF9TDjgih0VHQP6Yv1qJ
4DKcDkb00UIexeXLgH+vuu1p1mVFOInDy0OtFpHjJNiCIHWfniq7azBBycGl9p/n
ilsvRJ9vEvl2SOtlypKGYGYm3gHHKKXzviLF/7AhsDBKt3Cx+Rp+xm9yAGv/sQBd
LW5pMVIZaDi0yRLrFMDjaTj+XBr4Kw1RcOgT7v23Hl3bWpM1BCYy/2jULCMEXanA
y9qnr4Jzq/KYyTdzdikRJ2DriT9gVHEOkTNY0QxLLObkNA3jpBGMdjkCeWrfcKle
JcNJtbPxpQ6UKX63bZbli40G6mAAS2ltJ6qlqBQa+RQkl20XkFJDq90KUJL09DGK
tOOPojgzirTZe7LxWLVD/DdHCvRgKhqTvBCeJyXkLxjLZAZyviaFnMuNuHgT5Jqz
nDsRZJO/hdE/TF4atDhX9xCcFix2/g3sJPylp8y71L6/jMN1XqDyhOy0HEskSJuQ
2Yl43h+ynWgt4A3A/mtaEyRgxDRV3owkJCuvwibMqaEDKw838pDnlmVP8aQmcUBQ
kI4M0XrvIgj9EMIEzZiVYyBx0qEv+V/9KM83AruWklvCLJaSYwgdybOq6M3HsUQt
cIF8/KaY2Hr1Xwum1bpjkrnqVSYpEgwQS1jxEStkTFBAtH6U2Jd/iV+eeayfX+Sz
u+BtO4j26qwhxlcnVgWqvkMDUiZazmprmv8f3qbmb+6BmxpjCn/RqBRLJT8jw3mq
k8sUjIiJOFzUj3ImWJ0g2pLGx0XyeCIA+WWUCTxpAt8O4N7M9Dk3lQyAWEzrn6E9
OJ9KP2stbOK879y6q8dt6WsRxPUvawoecwRdTzlqFD1MOQ3tlnDe26rVDkOiZ7gm
gRTRkCBtY6KQt3HQpbI1mkSREX5Qd09Jp6rUtc90vhSpCS6xChqFRzwBsxqUbXnu
mHkVasS0wlReTegydJAlzy5dfHMeYU3lpaMNdZzzBUU5dNBo7VMld50UGDcreB+u
XpsakX82wPFMJY1+RW9jHVNKiDo7JROQJ9c0Li81Vww3ZaxXxCKHXNGMGPiuaZ2D
VfSlKexOaRKXFOOxxYuwo/Y8FTgM6PJ/Pr9Gejfg3ZBiMKOrofZoUqw4wmNWhsJB
5iK7fsORadhLOKDwgp+ovcJtUS74pgWnrMxKRxL0X4TgXkFz5ab7Gb0ORA6r/k0Y
r8Hl04L8gj1PZJuPdhLaF70AStKWxm8GbLbfpnHtzjE8I7eoD9IJZpzu/tJyqibP
EYN8+2q694FfxmGGR2B0CIojMd7LGdkLgpKYgdP46bqHy+9thk35L7gu0shHXrC4
J5ZtV3FQGixbPuYLTK7GW/mGQ9i3ug0pZCmQgGiO+4KNKE5Ex+WYLYP0GkOutRmI
AZAe2k5xRewqQr1sJE5wGoYcpgSQrMwDNeWxSjyNgHGo4ykkIp7ChJ0S2tKWbUyp
OgOOBqjLNvp+NZDc8GD7ar5aJkFwofX903m501s+5LLm9aRBg1HGpqBPhRZw8j7B
feQbPSh/4IRUi6pweCVTorCVYf2NSAjg6T9PbJYEor3qO8QuJeGLHp5nBPlHbHsW
6XyaKyXmGsn5rWvb2zghEZqxX1BxYWawUxJrk5Mvnx2Sjq2KSnuJeU2HXOpoehxC
KxjcISXRAOWxyn48mmFJy2UgYikkun706msSIRpqF9J0CzOIgWhRqjQLD3tEMFby
050KfGlSzeiMeV+6Zkwa3PWS7Uo2fpB+dr9TwPJPthd+1fDdG7sTaSQwvOFV9x1E
vD6ELuqZ0TXApYJIi37HJBjAqWKoQI5kvsUjt1KLDzC3XJKX8kdmYmkqaLC58+fE
WS7XMDYNbfX5N1Xa9yAKc/kFIq0fPilZEISbwhO5APArezjrOj6qnnQjRs2EDWMq
ec9WvQZXiAp/C8dRTW0lAR8hpEBCe+PgJqQ6y6+xJ1Kqw9OSF6rrkWSyFMSPdw6/
1lypenoGv08AmAa8ZQjrz2IMDCh3Q3bjLI7DhZDk5LynQDTZ6NevMjQgKdqqp8Bx
vMFWvv6Y2V001bevpduF/6Rn6C2kDo7CwG2xsAbp8TCJYzj+dJqu4AwX4XF5TBPg
q1tUoDL5qXHalOrGcIvlo/VtVizhl+fmprbr97hHc4clqoRVRYhC/52T9cWIr/09
mvV4aaEVXfeBVR89Xvyyz1UAuaFgxnvtRHNrdwAuorPBhbdt9wj0qxBIQwNt3bZ8
UoxvTDvUMVAxxYDBuQ4IBC/6AX0C7sQs5FAbE///jGXNm8EiDlrZbCVEQNtxiRYu
whbNquAkWr8ncu4wLUcVuLw6adsU3Fbl/Y29V6uwTLqdQK1yS5Y1+nzkfS9n9gF+
y+osth0W89NYSyPU7aGQt9doLeHNmU6Im5naDeLhyRH6CmAhIpK2arh958z1KPO9
zEO61OeHojOdQtmwEkIi1wOGIdjLGJDuqJEEzKqWNVBa5WE3YwZ9WANtYZllzkZX
iiodX1u5ulSplwVteWZHx541RpGB88iw6uPkbkfGS2JnKC5DwT5e4DMmS+1zappy
9T1xty5aQo+gSFrCSlBbRAKa/LI9CTwMYJPc5JsiPrUG0ShvLjmWgcSvcuzI9EGE
Nv/A8t/7LrLJTG4zyGbhYcDfMYZ9vZ9s8Zh+AF2EedB/Su79W8SIfJBvgEYkRWxZ
EnsiS08MGxEb90SmP8/kxNiTOgr16pVgHJWDj97Sj20R0r0mko3p8A7fFR838A+7
kRWa7zROx/yoiN19krUtT4Fep/YnkZHbfzOd6p2hu5iI22v9wdeiKiJpMLx/d0rQ
x8McAK43Va9c4/1JCuFS8ODs2ZHFVZxfsjpvUVqkjV+zPakw+22RAaXC36mCAfZN
++xNfUX5wHK09WJfO24rbTQrF4W7/TFb/Gnk3RIUMKO5yAifdV6LSrrEAWqL5mr+
0LhPnXHA/Sz8E9ZCPwGyv5AkXQDNtnwY0MM2Z8+MQK31nmzHBbFwbmiXHwWL3lwg
jpFEjwlMNlY/V0oF/ynvLCYjQOY25VrG6/XhWRG9Q2XJwUe9x6wnT35sTjBuw4CD
OnbA+VTElsO0IUVRgle6dcSvSyqW41KUwDxWEB9nT9u3ueE08gXPNk0tsYN/Rj4D
yxP7L4yLXsAZNttRxiO7i8Ok5xQ0CFjfwu278FvHwjZ98Wi5qO11K6cUy3mzuMID
2PurDQY8m+tgatR0aCDPf8j+ZwVH3fLaV34u8AQq/0PS8JCyd1XKnJsR5lEX8zIB
i6V6zKDQVP+haWr6O3MYJrkSlWtSM/tG/7/ZMDiqtg3ZVN9qr36Sxu/rOnTgYTG5
GfnAZX17KN7U4beG4WJXjYcjpFqcwrWezu5qfJ/lXOFvqj5agsu+m9aGP90Dd614
+bR4aTJHpqbI8+1/h1uy1e2nTrhrq2WSHsAGU3eG8RHAXwGjfg2Z0G0f6199fU0s
MTWW3he3lj9FKTdqpPLj5V8KRDrnARMJOoFg20pVKAC0IKOTdsKLuiueVto09/Pw
MtRgtouD06VpQBtpsR5FHyou+bI2ADr9MzXG17v7CfVwcvpdfT11emeTq3FRDoSM
toJaHVpyRrwhEB5FI3Mg1T/MmLycdFsIv+Xz/TxkLITVOx3HNZH+VqDFtZNRI1tV
zbZpbsmCeI2sJ9pP0YDNW/3WQbN7sZ+ydgHDXrqXVNM6+rUHAAMnV6wSlyvX0yUw
e4pz+znfy3SSpXPIfx8TEBIdpRLARasQEUj8z64SK5p0/PAxpXpyS49fkbfF5kkE
pH3HtfKWe0gdPgbMX9lHnhgIWs3Cwd3MWcv1JALONvv2A0kxmO4pV9qHEw5oROhb
IySZsGSVJ4SzaKC2DrFQjw7jOqLSw8ckTcvZWegouzO9xfQH2n5H1oz+XzGB9GLZ
3XNuJ6UjYNgfCQkaioZdzb/Y4lUiv015IKOy+7px42acKC4C1xkF/V6H9vi9KCVP
g77FZbTDtBBtcksQIMyCzDJnDqZirNeOFoWHvwZLoeWfDNMKtRU9EoP13H3J2wvY
hs71y6d/fVKyr7relHZ10+YY8A4co8w9carkUQO43GcP995J6DbseQJ1TSYzh2um
owQnOLJgTbhgHni0ccEKhpeROqr3IJKPgHuWvRenLNGm5Fk9KeCmHxLp/ZpooST6
rOdeexK1qHggfsSgUHyb152JfyQwzOXMYRZ1h07cKg7cxC3nSyD76ElqJk8NZOBN
9FXPy5HCZQOd8CTPgt8k5/mAFWNJdxpCjFTUAd1tTfpaey8jNzf4MiskYBWF9NfF
tN/jmA04hpK9s2cIWU8uDjfhVHqkmOOCPGWP9+4zvp+tBSoFS7ij0bxH5k7XPu3N
2mUXybWOkg64Nv0SdgkAArxYc75Nf6nDEwObTZ8LbPpXxVqbPxoI0ygkRwkuL/k7
PSnb0mlyaLC52u9XQggRVwAxJ6UDMStL1mq18qX9tmpGgJmIyT6umq4YsMHMRhmH
ytWtZuzw1GOYeI1BBDXwq13SHSjqexdm9h48iQ1WIgJsLCppWJOzI4NL7wKz5SCI
YLfa+McXK1T+bzhdbdpAFPYVj6sjZbjifHV5dCVqte5Z041p4gnmDqaw7bGPGQo4
IfNc8TAVyUT7j0D6807ybpiJ/8TwjIc27bPucO9fpKosknII9UsGMFRFZMPhvhqH
ZeZFBOFSoh2G5dQ0O4kzT+6eu/nZDbNudnlEHn8sxD/m4CmHOefTf1WFydLixdFm
XTO1xXs+Wb9HjGly8SP7kL8A1CQKt/WUR1ZO6XYIBtqpc5iqT3ZE5L5JUZJhqnec
oX60dulINyMnHeo8FQU5lMrYH793CCCmXoNj8k1wSGQlO1kxEYNDWV1YB8p0yugW
/1GVucXOV3fQlvXyQik2bKxQYcuZqsckjvLQZKNGQwLagSKg+ilxODxbUB0X4nrh
UhTuxSy+94XnemwP4voL5lWbPgrle2av4BbQ/9CMSG4XMaidu9ZJu/Ybl2TIFWQg
0Qb5/pPWJt73uxjShag4NS63OioW1DJffnhPCjiKAPRYgUcuFsjCEryCrj3ttXrL
K+xwgIrXZyVvJ0VU5VHpKg9hLMuI7dtL/39JGiBpPb05x8a9LWRXBLHFDHcSbC1a
lCNpyqWE/mQsW/bI9uv64aPsJ8n+SFAxHw/KPbyHb/zPXr58LLEjHkictEC19w+u
xiRiYVe3EiFxzZff/sG6rgmClIHVGKhgSL+GvfqS8g+Lmy/8SyBCARSHo4mSRrHT
s3XD8uAiGUz7dD0Z8+A/RE5cT6uEcdDD4k15TVEfaljGehkt4XHgkvtlW1lkNAaH
3OGxeV61fkHjlSbzdjIGdKYCrkP7JmdTuHWL/EeBknD+NM3QSqhkAoHXG/EAKTsp
8rA3pBhPoCBvrYtaodBhra4CzYIFReF1lpjt4IpN92RgiQHtVGaNEoNmL+m05UAe
87wOvDEDfpvYrzjAwa5vek8Umvo89o9hdgorN7ZoyfvU2JplriWNCIbHf3gOg2mV
/7Bm19zF7trgUM2he/Sna5RUGKXeFgpi3MCbZPUfsxGcG5kJqmWIfCTCkH1KqnUs
qrjisfX0BqIJVspNcuveFRg2uXwova67crYjraMbO1DnAhHfGNCRn63o0T3/wkuK
yVWDiox4l6L4kcyNmBlu5z48iDXxc4bsOFC8KxHxTGESFvhtTREGTRlgr9Bq5UXE
ZXpkyIcBkhtMJzTKqwS7kN91oqSHGzf4BY+Q/ZNhfeY1uLeeNrkLTF389YBQWbFj
mXBW1NPxKsGA9zRRXlTRUBzyH0vxngqFwKbb/Ak1E/m5YoS84lGz65nHjftuh7R7
ubw4znU5Y+D3bbGPqWaTXjmR+GK4KRn8fRoWwgvgiTXBRq6KOKE02ftTlmTnjIWN
m297Ct/mu0+uElJc0WUtmZIZ16kUVmRSh2zpokMNE2nniKlYopsV2/na15zNoSek
nGgnAEyd/wNgj+/+7wXCTVlRJqCptacQn3ExBFmD3hLfB0CNPMljJvzy5ahWrhfE
giRQOHpyTQ5tcBnK8AtTLEeEedAu7KicFbAOH8rZTLkXa6jX+/OAn2njFI03qLYX
aUUw/rZ0T+u1hjbdkC0zg9lWyv3Do+2+xRsClFY3v/S3G84OCZQfG0h53EK+Noz8
wrxNS0qQ/6mYhSOly7awod8PIb3YzexqvI7UgDbHC/R0u+z0FtzGgV5XLZ7H82mF
wTNx4OEjLpYz0irhxvViR6+tmGbhmoOiBtcoqRYcq/lkrDdzYcbzTaXhIdyO2pgB
WF5WdsgNoLfW1XoL37DiFJCRdJGyuHLjTXX/aJzYuProgL9q0t9lS1gPL+PJ04MS
cTV6616IPrv3FGaiwGY8G5lnLZX0w2Wi1X/9OJCDWKMB03wwUil/vfPNw3prLcQi
+U3QQtkPDsauOaL8C4v5lZidqEZrdRrzEZrkjs6H/92Sf5ODZuj8+Xp8neHj2189
U8mlJOXOqilD04IAHxD5KVzYySk3UgKPOm/mML2SZ5MOJhEufwhS1vTRYnvGwyZH
ECqUxLl/aFFAQvjeEGkuDBkILlGtenSAt2mIApzOfvfpwzw83US+bDAeYlqULoNX
sF7Dhs/rBMmZi+05lzXTRuFfQ2xSAhJpOON3iNUP6bTYc8vRYit5q8jsGzRcPrZa
UF2S8fpuzIkQMsSxVwyc9FLyIgEQSMiIILZNhk108K3LUlVmsWW1SSLn9ETFyNhx
Sls39PctJp9iwi/dK7DfyFuNiLMePCJEa5WIAEXscHw2UcDB99yfti72+JvvxQVa
lnYkCMG7jQSTdbwM2ilhwoKCGkKT5NJK8/D44OroOdU/UK+LLoFXgfVJ0zWnqRtR
TZszJLgU/Ub8mIc5vkF5IenFJpEhTf/XRwbn+oDWrvu9gCSTwA2ce814Be2n31PY
DDepw6fW5Zm12OVR4JJGec5FNjcBOcN83RZnvd2QxVSxExJ7aYUNNCYbwiP6Qvc5
Clcg6smUogEil2RBY0rgtbBPgnZS+dE3yEsVxCgrFjmMo+mZWeJau0oVfRTTD3D2
ZSkKoFGgZndJDtSivfEVd8Ogf9fduSFlTlEnD684dsCo4Ngoj/NIEUzUsHO3KDoO
gsJEBOlhg6aAuZ07oXqm+92f1sTZF5jJnTABS+qsFGtJWmCGswfyHBn+RT+ruP3j
pNR7wCOGmY1i+Yw1hopznpNIgOo8iz70o96f3/vSFDSydgBcvn/WWE1SX5zmAAId
BFcDkNuHG8dRSATM62uUhPbwLe52YgO0UZvmHPW82WKG015E78ta76Muwxd2S3Ee
nKgxQoszEUPLIXzguYi4W0gCIOCBn0vmcENgomsK8W+waCxLzothz1D5asi2PTcB
ZEXaQICdeM/v220OStKRP3G8/hIgm5Hc3dCfB9P2Fs/YrbQKiZgrr9/ad4i5osa/
/DM8hENhQbFY23X7LKibX+RpS4X7ww1aFEydnlZTBlV95LEQgN15c70GnfH17HkI
htIQJwNpqpnZ8PNDrRQo+I+cd/HcR7CxpLoGXP6f2Fzb+5H3hv042ItdCKlLNDHO
2Lw3sdSMqVF/uq4+mX66nGwXzw74CKAiqKJESWl6NSJGSydB7vazUncQJUeFgrLX
xkmn3n4EFTGPyLVrUgUTKm6V7LRS8nW4wDaRRjLgtMq9xn99a5c5xfAtMg7sYXH+
xDXMonh092zyF+vriNBE8XvWAeuHvewV5bfSXIodtj3o76rxj8HcRtF1df9X4e1A
XFwobByS+PpccbSyYLLcnc+IIJRNt1iVhfMHqOzTJ3v9kuFdjJ87R0G/C63qqWZ9
2LFSQtAu5b+L5/SsLq50QSBYCWINxOTCZYTXUnePwFH9vGT4v1lbzdUCklpltrrG
b689+ZTT7oCAnYZ16QB5WbWQ2As/zqOsfalXbkozopu7gEdMRMIbURbC9IGM/jUX
K1aJknm003Duc0VxpUZC0KSrCkm8u7mTmpqReBgFcLS9k7JNnbi4LCFgnW/j7Da/
kudNHrxJneB0A17YSxdpOaaq5JG7tb6jUoAXu9ksXQvkNYDDkLPSmaivpuyZHRsU
5MEPyNxlwaeUFt+8VypKqUhfBQWAVChYs7tiODKfJCF6lBTEDdvMf4DHA1T4Z7BN
dmVzCiuwBSqzpREhic0NRQj+SF5d163QtS0dT8fwz5XU4x9If0FKoyWe6ZRZkhqf
dn6/7nbjhOgeq3RG2ce/etpAP+V78civV2Go7RxP/rnZF/4jCByTzk+QITj5Nu/2
QF5CdvPHnGRXMmKkqPgB8Xaq9jDemOUnrRuaIX4B9i4dfk70LMj8Huc87gQBDAln
eUDcUza4k2U+3YogBjYVmakVmCdtXtrYmE6L1r9WiqFgC6a35BcGU22whaXV6sTy
/n4waZCp2jFJYHQnKYKaTjoYAHMbGCaxmXhIxRPfOEafeOaa5JCcqtKYBDZCs62L
kzJMzugV59xNOYJtpyZjR6I6+ZqSrpu6DhWPllisMWXl9kX92xI3GpQHsJPrm3G8
VTgWW+cQzx7QFn4uHBO1cVyWcO5llXJEN9gdm+EIC9sE/7XP523/h3fhT+8p70UT
E3bfYVsiTA5SqhRHhC27RForsXk/R6WFl/90ewg47DbIpOvb2K2DJdmoeTyr7o1Q
bJWDVQ9yN9IrVZUNTyp0wJIpL+qo2OXbfxmbzPfXiEM4wIQ/szM9vzHJd79AURDM
rOut45fQVG3giBSY8yvmDV5ap75j9dUlibHajtif2k/MmrJfpWfIk7wGYpeSgc2Q
Yfxfd5PVsyVGRQyaCNO+pKUuOyvbNnmWTrwkQsnwMCRIzjc5mdlARfOjT+gYtR7r
tP20YSy54+bysC7AAeG7aG2ok/hjRMtOoBWhVcHoNX4q60N/unLmle/rMxgvnS3s
n3skOaw8djzmpi/r42i/PkpsXHL7GFPsqJCQODwF7I/+hH6gC5N4iSgoQQuXdlTG
gLxBwrTlbHBTwYHz1y/KQyucF88CScglNCXgaHpZuv8mkraypQXdQLcKohtl4qnP
ASxE4VGq8hN7TqUIBYoitxaunzRkEwAGemt1XwVnrgLh1DLF1qQRv7RehKhqxYif
cJNbF+SpiPqL9U7+4jfLpMpGcMEqUkERi+A/2ABJWMnIbv0CcJRf3OSVBKpo5MdS
P0UfI7AfRzFKwq1kqXfCjZo5NlID/bjw0d4rgG31x1GjWqCmgsDMye1CFmeRzxad
grrWGNgkBWvTPgu6p7Ik1/QFYuY2ftFh3NXg4pJQ275dYpwGgPg/Kpqa8fjtnDAT
lIq/SdSWgWjZyLp6CgaZrxcGxmXE4xFI6Z/m4QSktPbtMqM5rzV/lwYJP3JyaR7y
yBoBJcmvwP8CprOxpMWX7UBDcjta7B+VIcSCG3dOo4z3zcHX5MvT12LjxlYSgdt3
Ru70OEy9IiNFbO2gwdLTFFw9Wzqwc7zh4rG4u9U5ShVRDH9g4TpLfy4GedXeORRu
HuhANTZD63Ka2Paq418SVzstSpj8IIanSE6m7gQMAESeFber9zZx2DEGBa+yl+DM
yRkreA0abW97n7d8LO2CrlKWixvU2Fwag5y0/wPRu0ZNVyZJFfUcGTIOGJDshG4Y
KHBBcMuWRZHwVG0Wr2tj6SlCyXQDbITFDZJmJcbqOaQRTjEqBRZjI3PenJC9+SPk
Y8kBxTjS/23qERFEhNnI6/lzegDc66n8PPyv1AzNG4ItBN3UXQ1W0N8ihIWcmsLI
mEhEGtZjSuP4A32eIYfO1zV1KGeLzwJClwmTYhwp/ycZ6p3jtrEvJAoh7Ke+tei/
ctyjCeuqgJ6SKgcDOjvuFiNGCR2LnvCX8G0dSmh8v9otxg+3DTCTi2gTw8hPGFCk
H4WqpPSY+ZOGhjz8j/+BkH/fGktfEyoAkvPRuLRqC3DYDvZWRItPcBj+LYoOBCEy
fL9UqJxTmpARYNzFBuIGKgXWAXziLh5VpLpOYWtJTvmR2wEEZlebn82qC7PACG70
OiSegn0y/VXqV6c02xrWb/sbpbwXZQUrGo5HSgu7tH6sZy3ubqKGZT544366WPnJ
xD4WgUEGfQ/NT+5uPCq8ZPQECZJezSwG/5u6z4aAcPG6iXcKd31T7RgeQqNcQ3QM
eGBQfLmQRr4qrTpEgnhZF7d9776qiBEzXSF6LtW8d9KsK2AZjW6K0gEpx0A0BVsf
HIpk0rAOzIAmPxInvZA0QVhEY6ZJsG+K6rAnsaR5eqg+AJ+5o2Njm8eojLSRNDfO
V+xi7HnWOpHY2449jM4Ro2PcaRFkADFzZLKPxqNHGhGfZO4nWosvPv45cMSBWKlG
dVBdTJr/Mu/eXV1U3Ph3PRBvw9EQlhqi+dzgGSBHzF/cvduc8ltvattmlFyDn+FE
0qiUWh+GjF/rcMomHRDxv8/IutUMvQbnyuj6Y+PnXtQQVTAXazSbbsOeGrCgN0x2
rQIMb5ITbocbSoqaSqmyDGMsKagfy7QNPQJTwqG0L+J8Kf3MfwBbml0lYycWMr91
lER+IJvyLnwO4YA5XclcPH58WEnHGD4cmA97Zl+ygwIzKtYk1elikm1UgO0UL3/2
HlPTlmtVgoyGXaf4wp+dVfMY0sKFp48HO/NAfhzmRQFjYE7vO00JkS38X1gPZ3fm
XPrlvWo9/YzvcWy0y0wYRrZebxbEOF1Wi7mM8Vd2mHtMCIBsrnioO0t1w9a+y1XP
WkgIExhfqzbIy/pFw31Hjx73G4ja+N8MwFlNjHBLL2eK72fQPRAGv3JNNufy+K9r
ED3v7+nMMSlllLMzalKmPWevLjnDi434RGQhoZj1Sj29WtjLJyjnZn8Jrs4oOfoW
wQH4uvln4D9eeYwCOL9UOcqKSVXaskoMNJLgLVzbizIQLkwY4XCmWYwLxTEOFcWp
wjbMSn1xoFqvVy4pHnqwPqt5cMp8AI9bl0wbqqX2d5PmD+P53DFMEuIynTziVKk/
6TZPRytf6bxidajSxlWCR7cH1tLjRm4qdaEAAfrcJCD2LNPzK/KnJ0GojDbnJQmN
i/XeVI09B8r+dXD75hTDhffH8t4BhUiPHa2qY0lMIalq5O4lc3JCdAyVt4cUxhYt
ovrWB/guP54vBBL2clJBiK9p8vMeQkgGWUv/xitJLDpgNm5ECJnk0R9882P0Zz2e
h2dc7PfTWoLPYnY7+2yDamxCby/26uW7UHgg5nVZF8Qvmoy6eo0+mqOgksz6NV49
Y7mGEe7THIONZ15gHs4hQs7ukPZmDXA5t+4XwysPpM4z144LFidKdvlWxCLjqPKZ
+V1p532j6zl928g4wLePCXedS4qKVVcDwaLGfIWolo5M7ZcR/O4zykFYY0JO73pc
n3BhAls6n79LUL1xDnBp1neUrKa+TGkpBtFrIuTbx/L046h8Wj12jVTekH5EVzFw
mrf+BkGIg8VDPsEeoucNfhK1nscZd5WXy9YRXB47MZCK2eepsfV27uKfj8hlDW2I
EuujnE6OEeuj01/djBOnyQGaM3aEhg5U0NSCSDWhMSaIHRX2W54yH+56eNEQvyC2
VuCvXtGZQgT5IJuZtE+KD+btAZ2d4n3enAX0Mj4MlifpJ2tdFpQzevVrF928wAI6
dyL/UjDcP6n9maC1pnd0DKlEA/gJQl3N4FaCtj6XN/D+5IhLvzREwdL8X2ioOZWj
KuzjBmlcNhk6Dr+4XcGTC74KgL0IvulX5S4Nch7VB604IWaiBhkxWKRdVa5LCrKG
XZEQ6pUohL6mK0kTQcw0/Kbb4PmucHcZ00EJv+ZWYQXiFzpPbZ/LtTznEIfvjvZv
vMwFyXE/sNY3J07ENBn6zh9+bulKH5Einy5mksd+01wvGlP0r/oD0HPSJbWJRhn4
6agAqOcbHAHZ49v4z+5s1X727SOhSBFm1ZSHdYk8Bswe2PpX17zbBr7mR6UmX/kb
Tz+eIlMZlbWn77GgPZV7VGeqXB6xZpKf6BIh/hwd41rW+CRoeuwx/NFYMtcbDuLa
TeiT8M7oeJfpCJYkPaw/Teh5cxWXvSIXU1nluVm10ZgwPuDNWWZZa5YD3Rbcaji0
YA0ckppMfGcoBjolK5VPI0S5y8BKgIVUrrdeSEHsLDxMrA/ZcL86hQ/Jtt3/fCuF
P3Y5CD/nynsFw4bIx5MQrm6YD3VYGj7XlLgKLQSBVZ9MKNCuDmgzUewzXHXwsf6A
a+PkCvU8jfU2nisJJ6bv2vapUCgKOIZoTsU8FN5s5kux2GxsMrqShSaQpqUR7Vjs
wqZHGjE+Wt99SfBwTrzKCtiD9c7FdyFjb/Bf2torAHtXRdOdtBUtq+W/+qmyhPom
AS0xzN6SQi275EWK7oPKaAm35fyINJK7D2du9qgLcPWxilYMRr2+WHn/zMVE//WD
EfFkyiY9zqQkeofdt1UfA4pou56pzMY48PHYX7MBP7pWYmoeOcuAQVbz/sBAXoic
cgt9EmCOAM1n0BtlgQCXg3SNoWm3W3K/k24C57EJw6PR1GUfaGTtSq83RDCMD43E
kZbOFFtyCjkooz1+JeUgLd4xo0E6JRa/sbzpHOUH4WEOWvZHY11BUF3SRQrtnbPq
mhJaU/RjYvIH+1u9AyERBaHrHFM2G1Epb/ls1HiUYAA69lZqvoZ6jfbj1Soci0Dr
KdI3rlLtd5c7pcpka8KDNnMWzMWSOZ+xeE9RyP+JR4LlUsTyPf/a4tf+5Gf9mPEN
KszILiKSS2qdQSgReCiMQR+Ud6ief9/kKAofM9/Z4aGxVw2iJH7mAOalWKGZFQd1
GbkZ6BChDmaUkkKaq7LL5Z41np0NrYaIztJFtduxT3LnFP1tJ+fwOp1C9JIsvpTn
PLf02WGrZCX6toeRecNSDZ8HoPcAwq6feEU9s8wjdUxP6ep6yBE4/hxFoTj+n3Ra
q+RaQvYLrehoCgLtsK8meVeCqEz8dmAnwqPVMdhxtctlhJTq9Blg9w1F7fbwPGT7
2gqTIdr6/DoxudvVeEfNgDNTNw2PFkZG7u23YP84pyGeub2TRauILRozkQXcepkp
uXxqPANjh3vi5Jduaaiys0CmKulpdksAiL2f98OtZ5FY19XbCwGKjBiRjf54HX3d
9jmMtKaN/gxaU7Zh+j6XoYo8ANM3pxgJbp55fHXGVBPC2RHS38yHoiv5PPpX57NI
4om6ZaDgpS59Ec+mEFwibFuB6NW9u1vfHuFN1K1vVxQ3Xs99I5AHhrVTaWzU+ZSr
Lw/p9XN+oKP9YGXp4FH98QqhyUhH8MrabP1oI2/nGyCCTUmrQNyiwraRRsONTc43
fY5DYz83F2FDK72rU9JsXh7rwSjeT0p2zRb8eiZMkvQqaYsJIcbMdiWKxHr0oN5q
sZfjhGqOE1ZOO+gn+BgTLqSR1tonJH3kSxfpnngl/tQHKiyZ0Q6nNhhO7e4EbcBv
6/CG7Ue6pf3EUbewOU1OO7AHqbnhLleuVbRZqeLrpt9btcgRqQdISXdRtT00ZX8W
seEUhBd4zBuaSYu6JRU5cHr6u8Zb8j0b9grGMz97kAawI1KBNOBUbvHDe3EF55k2
WQlqVACsLw1CxNjxOZk+o04jFMHQ2Jl4qY1rEgNrapBP2cwO4e74ZT6SRosL26pA
96WXup8hhRsLB5pNnh9b9z6iFdez7j6tCMXZRj3H3x/z2d3OJm+her5cBNOehv04
osRQgolGPWoVFuJaDadpxeBst+J3sC9YLF253qri8x62a7LZP7Wr5zuWXc8kHBeW
furhYvg9VZKXU72hcAq9n1auxEbUQazJRLDVyZtnShno/pEcu2Mk/dUz1ZrwlkcW
WNylI1M9RDGKIdjz8VxOGReh2GeulewtPRa+6+xy8euqvOPvrIKgzeKevdMQiQds
nUiz/YqJzkvkuJ3LJGdSaQR7YsqMzHuAOkqsD9JujVuDd3z0an1b1sbDFGPsPmdk
4thipU0NRYuTFdy3AiQaHB6uEuAkhkcTyyjhsY0te6rchInQH+sMXZi1BPYVf0g7
+q7jM9bettWEH7zLokirpY+v7qrazJYuQIpLdWTAB9sK8Nn52pdRc+ZsuwQfcnvo
noF6aWg8k9oYQqBZEFzFwAH9b6rdLnORxmYMBtAt3AF/ZA+Fuq+5YoIoGUEDL/NQ
zpFInDVWx/jPaWtkTr2xUedaY85qi0+4/gHx7Q+S/dvQCKyYRUbUlkBAGiL5ccw3
KL7sl/eTDjTa6uz5YZtmGlapRDkJexl+u0PxFcXi2enYAM4MDEeBtwRa1cP/9oJO
hMGVgB8kBIJnMFEKM3djFgfZtMHFaqOXEatYRV+Rat/AiuamunnkYyKET6G+yxgV
+SV5ErsFv5FhYKLdN9JGksAHpH43qtrKxAAJ3MYd08K//Y8/0IxhNJurYtw+TQHe
qtKuAto0hCEuYxiz1h0UVxkRMwEMWFxn4wvt+JUQ9Mm5oenGJuQ1qqmrt8nCA/2Z
OHok3ZC3fCtgkTsRnOTiHXrK2JnLKVwkEcyEvPvrTVzcvCheP8IcPs2zQjd5LiXb
1omcOwsKPOg32WxdpmNUPryU5o+VxDZndv17eA3S6RilTYYFO4wzp+H8wJ53pXQT
7tE7aDixaPpFkG6mtCZ+vwWH9nvkrKuwg7B97D217FBrZM1pkDCV9sFonTXY7jUL
ui8A/luIAG8MYjQf4ubZ+/JdZ6c+fbdAxVy47hN4JC+6a78iQ002vxi31FNdCgT2
RrubKSpUrOh0fhmYt+JYopVcWjOgF6bIvRWDYOhb33E663QbOjpOwBkIGzuCCOYi
0hzlUf9HRuFTMy5I+YjHeaEJsNCtIJobtqBYZRHnswCMht2kSh6/ly1GiG2wSouq
6TeUJnio4sI6B8jjJwPnznVx+UBKZYTM44ZbUPn4HeqMS52+WCMJ7tZfSBC1b3SX
fNsFJnlyE7iivq7KQhgxzpPZKnxaTRrKYBvybA6kp1GR7GJN2q5qYFA2L24xIisi
DGWkrv4De99smPwJBX+qqKncNX4Ez/mF8TecgR3H15Rx5d7UrLltydUjRaGktN/9
X5elmpGKecq7rMKtex1VXISGknFUkMjW0g7r65JtXeBVmjKTdYA2nC9hZDATG/VL
JnK/ahqnRV7aMKgPdXCQxqRo7ldVPXS4aNYB51GQK3QPDBYJ/tkYzyVroqnHCmmt
EleYNG6Km3Eno8EWZMcpF1/rhHqACHsjoxaaTsaOm74IIg2blBpMLYKrIPMhXcOr
zp3W+D3rph51sdT7yPCtFCNIhLnlrhh0RGTFu+CaTkn+IiSTtSdhAipZo5Cv2Q+j
WSIlLrYiIBLxuBwswA8C2sTncBNPNbQIT7TdbJwkCvFg2doM3zLsJ3j0PE3La5Uz
IyCrHvunbwdOxvFyqTJZW2EKMQvfX/DozFnpcr3pimu2RdyuZSFO9oXyzBJ+ZBIM
WY4JHF1QR5cIdDWXqqXnAaax4jLfjv8yVbSw/ryUDUCveyl61fHXm7hUsTL5jUPQ
SdMdx86xRysM0vC52uUBrHkJv3ZE1qGs73OVq9BeGkPziliLUZzmmgWFEsg4rO9b
j8BlLR80d1kCWj0Q+MqUsqvZWRXqLBJ70YjiEhHLM56q/sEZ67VrRr0Yz2ZPQHV+
FpBYhM4d2loX93Bn/CrzRirdpSBz6I4sqfwBkgMap6opbPl8s6IBkLIeWPGjHg/B
uBzU92DrJe0/MQ3XSu8r4bRRnVZ4HnEJV0g1rVewYVXTLkjXaMpVnjQER/bhFfJB
4kSQRa3XiHrNXb2oLsM1L+ax2F+UaMRlOl6ugWm++66u396mGMsvhyz4eIESg5hY
jUK3OWNmhGuYnYW/0JXJADBjLOOVyleSlZ64jfx8UaIwEno18PeoWzm5Ny05No/N
5zHADnwnJ6zazGtRGF5iVg2adLTeDtM2yNVCNex9T3LjdFaWermLyD6fhJRlY/Wo
y71iPuf6c2yGFvNydbmivfbktbwq6Wb86dLQ8rJj/CbF7MQsNTBle1UE1T4m4s1o
fHqSLA5K5gAJw4711dZVNr6fM/OkQwJEGA4fAYUEanFxqwtEabDTL/7AUE7axdDf
SrO2Ua5kvhucMaXOfz4gTD6hETmDKWq7uS6Twqfa6wH5oWKm66J89QbE1w4lW4u5
7JGaBOoE5cHzWM7bahDHi3qangzwwJNfsj1uTsyUPoRdFGOHQYChmv6srL+MfuBZ
DCbfY6tb6YgP30cvG6FywYptuEhu5hwJe3VHAeKeUzf22zF5faM1wYvxEzmDlf3M
g02fdlQWvR5xfuNCIB4VoS8jBzBK/UJTHtQAkpNprT3/z8LWdXv4xxNWF41gFQ7a
nvWq/1a9F+fAIKB/+kAhRZv8AXjHMJN3vBAfKfkxsc+MHB801B+syYWPjGoeARvx
HQ5zYOXYXYE/ADimU7NPctAN+Opz3Q0iSar3er2mYi500Z2QJ036t+eemHS5JlJa
6cZMxfWAtg8yk2DUqDZ9njL+G/Sv2OPt3A34qVONmS+2jXeqli8mvyXAYQSqpCq2
2Vxb6WrPe3TU22dcDVrP0q51dKshqtMLUmucggUxFsuruiONWvnI2C2MiwR1xcgq
lIMPCY5lLoZJOr85+Brt5GgOjVLAHD5+BKLNL8SjKsaEzSj3ZkxQgdB25hs/VFoZ
4IYr7w3gewUgYxog5jBNQigsyvwIazqAWSmXQxn9+rdjPP4oRvCUEsZRkY/RmcSg
4HQiNXkRYF9v8ZcUMwqFAeGFZiNIfrVppagUNF8sMvXQ/WW1hL8iIC+JD3lQWRWe
atO0RzKLqQsMRKwZhJoSAmTAbtHrktY2XXfplFUymzBPB+Bqh21/TRVNOFyODzAF
yKm7PlKTWsFKswNgRLm2A3MVwbVXPA3EhDy4XAzNtvTefd53gneT1rfZwwa/e18f
LMhXSRxc2IO5FzBLTp3TOElUxB+/XEP4BTHUGD+NbYmaLB3HWpiL+zsiVlz/wRp3
Lp3JbudsUXfNgRcmPvs0rECRniT1URXw6L1rlYCROXrNlk21Fr5oNE1TTa+TchGU
K346TIw6DhUexPnuEtn5I5o1QBFLWEhXXWFK4dR5wPO0v37wlEtUyIBStgRZC0dB
5JvzaMd9ndKgBMvRs/arF7AAsZ608zHtQh9fWyJIKEETs0y6iwy9etBS/ISrLwAe
W9z5/G0Nk5wbVNTLA9mHKwAmuw+lAFn1vUwzpsx1NuV+nFnGnNaifFzfxUUP5fga
Ubm32N1bMlii+mx21fiKoNmLIeNhfchPNEck5mc3i6jDJRTVe0TcaewLekPTOAae
eDDjID2XF9KZ+GSPhaKING+VqFPHWIn1z+3i81+VLBuoLDhryIK24Mt7C18DmfKd
cgiGQv84X1Y47vSnKFtQ5+xnEZQ2/CXH3yv5omVax099sbMSEl3zmV/Fu3YUwfnc
+351T5iM/HYgVHAFClogpa6eBIB/0og3+K7hQPBjMChSyx+vAoko8wQU2S2igsB7
ctvd6gESiTXa1QH9f2byQuV1qSnxQQZU+VQqB/6Wtgj+JwtSC8q9vp4EAjMq/tKk
Uf1xaiBWNTsg40BRpTmWLICgPWpXIUhLvfCt2Ub8gLH64FaFLsZqIBjneFVhHpQZ
0/kBChDLlCQb9wpAkLx/NcVGZrKpc+75Pj57ghv8kiPiacPSqIhgO5MnoqO93C6c
urm0lAyswJdM5Zq992a8VRM0rqyYk0zb1IOdNCqQMMFnsEghYJfctSLUyCY81mV7
qk5YxC+07GNPWhxgZam31BbT0BRewxPljjSsN5Cqvn6iV2krnQLc+Wd+F2/UKj/b
/Q/lYRYwVbdPXWBkHz2j1v0qtOKM7i2FlkK+Pa50kTVoneH/hWgGVgaMRxA7BYr7
WCPOgjX2/hR/3ANfdJqo+wIIY7zFOKRC5r/I4XDWl7i+79VcTIBZ8RB+nPbEdkZB
UAjuiti8Sd6djnbAkWeJLvE49vkQfA8A6wNrGChezNw0BViD+dKng3xM3qyGIxKs
477aqEU6qdV8sOWoa+g4c0hdH3m4f/N0rNPABgfnZ8PVVrETnI+VKHADwDWA3WMO
ceeFtTMeGhNINawwu03Z8XiW1UrhfteeM/N99f1aTSyTuie75DXt5i9DLUl41wNN
8mA/Xp5HruSrr807nCvKg+Ibd82eyvsXFaDNyLLPWRs+tdp87cIlfM0m0/eqKiIZ
/DiiOzZFfg6qY5rRCHVmVOLRXVnW+Y1w7+Ptg4UARtRP9xlSROCqkIgja/uS/Xoc
hPkyL5iP2NxM2Lf9c+l8qbu2a9MddwiyF/nQMBMBoN3I4yybbswXg3ffR3fAcK5F
qhXJZxz+VdZWUKBptP0h9AynPYj3UurygUgxyuDdsni3z2XNJG0+BgyrW1gTGjm1
QeCDjFiLSaGzgcKlLvQcVc2jza1Dsl+r24wPDHAbi8A/WHCdaD/MTJ4RadVcsHAp
NldjEEZJ2Y5uJVfpDLBIoruMf7S8Mz1fgcfLnfsSGejqjo02bt1Lm5PIzbXiBni2
eAxqd4dLFIH5aqoeXjpqI7VwOCisH+ojcoeTLdHTDLZyogPw0oKWJm8vtUmVlHDC
HsP2aBXIy+bjFse0hy3PwhH5LD+ZsO/wbLzGsP7nTc7SHCJ5K3M2jd2fVpzZKaVh
s6U9Ak2Imcn2HT4Y3hrifpAxdKoPCX47ag98KB/sxeuYFXCLO8/+NvqWuRaJ5UnG
3nx0QnOVsYOue2pC5iN+qgC6wWv0Jyik2Y0vAymYoZqNOtziMx0Sw6b3+fa77UAL
AXdh4cBEWCxAoc9TD/PKY6PNOm5TwDE9ZLwtZz3hfTWFVZ8eoVVvOdqmywIwnYC+
oquYd9HM3WCXqz5qRk8rbMPgKoXm+8MqxI9O3qtxD1dDHRzs6agoobNs3w8AC7b6
tWETFOYWgl+E+fm+028DFUpig+1sjkGw1REYew6gJVL4UJDwgx27iJZqbv1/QAR4
ckYEiqJY4KaIH9tTfsWw4yjdKDLqpnM2AufxftPepbSLuq/eE9vdg8s6imAXAB0Y
77DGmVXerDIYg15ZcEuRHGQQY9zUMufwy4RuiBSTHgeOzxFFiejCSv5cbwt7Y6Aw
r1/9RQpsGB9s7ijv5TTgAYJbesBweWGSJFDFomlbJRjkCew270JicxzoIxQ9bXyH
9KQv2ORxeckjpy2MtTX7b8LXMw5Vv6DNfOg76uq4U4FsgYEFtg7m4azVCrPrdL2Y
SeBRjChTePO7lqh2LbAgn7N6LliiVQjoasA+Sn/Z3AsyxNq3u3/hC05N2QFODQJT
GMEswzJWCiXz7eHvj3W1PzRdFVryswgOBBctfrauVt8s7NklGemb7ynVv/C5DuHI
dAYWbcfheXM5JJommp8E8eSKlCX+WkRt/Vmj9ft1JBFkzOXxmhRQJKuxnTlmbUQv
ydkQEIgCGs4eQKNjL6n7W3kCzqQ6/FlQwWiSunp9cITCC2nFCrFVLPfjwqE/Rfjg
PVsSz1B6pn31d7Og6PWt39QX/fBn9Fttgm7bNhZe8AnsmabRe8XO5EsckQk3oayh
4wtzMfcQC4y7tF+25TGQkmrit3LYo8z3M10tauHyQpJYkMnVwsrum7F8HglKXAEc
pp3Xdepp9qh6QCE3gs4QvePUn4yHppMe6CUnkUN2TzDxujkEYvdzYRFHuSsf69gh
tglbXmqD7JKHMpWILzjAp9c8g6ON7Xz0IfutUjbQgmTWfvHSk+T2FwhkGs3Z2Cij
6kpGyXyUgSRf3D+6stAfcxIXfSp26ymjNhVpCU7vh7uU6+v4FnvrFFZJ/Ai8F7L/
1n0GSEGxz2tKmXTuw1h7njD9qyHg9+DAjBr4tlmbgzsSsLlHJmYU3FlqcvrAcqIN
3K2wtiBW8hQVA2zNubqWWOh1uO8d+qvEnG1szu03dvalohMeo1DiB3rk5rxlIqR+
rKF9rgSRpOeps6ynAFkV6ysAiordBfiyVvQwtSFBgilhXhI2WVKHiSVYnknYv4GK
9iZG2MKOyat6y2pTeGptzAdP6MFqi2PM5HDj6qPIfaTLbdnwSi9j3qQ+j3mtq4gF
D+vq52NKvUYzWwrybT40y56fxR+tORQpyVd4242dGw+NpRwACb2CwtIBonC39OXD
+WHYZdmQyOGb3ubOCfA8uzvVEuu5SEkKgVMcweP3XybeiDrMcHKygNKVVVfrC3aX
sTuRxTRt7CWYQGchI7cUBtEj0bvSAVWV0CE/4r2CNppke6k9YdlEg3MlSlzla05K
9hloS9gL/4oMF3215QReXMaie3t9EwCjpm0a5NepTy7BVrt1Upr4hPd/qMW+zsdQ
Q2VfjTtfbtZD8RAAjFcBQrEnFfjRc7o/BBrOrxddM8JgZZh7Cf5e//dGNYyyFKIE
zPh3T51nTa63/kbhMBiYDGg9b5YvePKbGhB9yEQ4nCl3NxQjEBtXJYkP4cOptxYf
z7frkhBWFwAl5wkbsn8VJPwLsnnGPMmmWQKFLCo4o8oXZL2rMKuXH6nCPSSBSetC
++Ri42h7GBJR/TSoTi8IIMZK4/8EkBykjZs8PzDsozDCm2KE8LL5ETxw48//yrDP
fPPBiwgiAGuWi0qT8uyHNHv2MWN0uo83PPJMuC1IzO5BroFRU3PnkGOodZKBaZC6
JoWUQOh6q2olgiSE0MpRSoeuNGsUzoKMOa6adyBe1ktEeuLBLcz98dmimfAy2E1Z
aQ4GMHaok6CzzaQDTwTtxzUULmqsXgSVFDXjcycn8348CYXnDYOLjB2wHXzJgw5q
ar2L0v3jHasCrqDuIUN6YRHYQ14SBT9OouusQEN415sotYZJTLWHReQxGVwcrpum
ETj5tyoCpjn6hRS8qlxyxoGkTs0N/EPcYQX7Bva5+HXZ4dqR99X+6yAFxgza47hG
QbuvJ3urW/KxaHjU3tRgoGOzK8ur69kYYyrAiG4CufTXOxWTcMaV99QdmaICHprH
aGjDu1Fed4wFmsXyKE97iKFiwLMucembcwl0lvDAIroQFD+h4gWC6JIaqoQUMz9o
Xr5OU9gSnVwt649SkesAxE3pu+GfBbd+R+F5BQbN5Gl5XnxL3vczzb9coZnzMrOs
Ni43vNYD/dYIAvZg6GIrDKLgIy30EoGZnVdIhTWhE5sDGyFr6SjEtOug1uHTa6W/
/WRy6xgqXu1/LsUHD+XSlfsEIUq1gpB1RVyx3s6PmcPl1QH5LVy0z/N4o9s1MQlx
zMj+Z3opmnsgf7EqKKYXuEkYPKxfhJbnbDEQm0ir5mnt6W9lNcjuVzZKGJ4C4B2X
tT/77LngYNs4ySKyYyZMoWiQwS0thZalVv6xlTp6C/qQNu1JqmHcO2YhWIreJ8Cb
ccbVi/ZsJW++ccyzQwzmCxBkeSkp730jG+oa9djjrg2TjlMne2A7sde5SZ0/hPG0
w6DycilWN+SGcm6NnIEH49N0BBnz8Y0Omy4r5pixytNGDRNQ2dsKhQbNk4Pw7Mi4
vdr1o29RBH3Hmch2D2JnzI7oO1ZyFg7dIxKOgEk+SottIef7rDx5DzZt6GK8au4/
XsuKADWBrFHs/VbMLkQDsjNZbFsJ5Gk7N7NILDiXJikO7+M1FpzLa0NlDtM9CyDx
5ftC3Py3Xa73SC8AozzGpnRDqSeRdSTa31P5jRsSScdvfBzUxuHt2ScFCXW19ZX5
f/JKwbNRXVHPmkfB42Ok+hkiDZl6x3GZfl17iCAdmdWsVcLk/mFVny8LI3tJg6hu
eV5WR4RdRcRTMTHkHD0CFS/KPspPZuKLMR9VbAYfzrc91Pdk6OczMbCPQ0YUv6XA
S1840TEQDWnx4wFxJTi7W7GzGeD5uzRPe/IgQfCUi0g5tEcwjWykpkJlPItnX/39
g7e3qxpGl88NH2+JLRTV0PAP2fUgygGdrXZYzkqiq3O3rE7PEYW62fmRFtuYdLG5
hTFUHjM/U2/7OtTULKH7eFVcSKuUhKoCHVugRFj1de7rIJScEjpczF1xMGyjQ4+z
+5mr2TN4W6sNufcgj9c1zBxMivfD4ks6EoRWDM3VvDerTTVdjb49VwvP2PmUclnb
Ch0dZW5c8baWI4sTKdpBSpFlg1p7H1168dJNJXKxMhwIXKC5gbmEyMj3vuAHna1J
sZ+PZfVzd2sHxBjI6geO2S9LVnOn2xBoCP1PAd/DU5bKinbkUru2yIIS4Co/ezlI
YPhlANFJIqg/1pLph+i2Bc0sjLBM/6BdlsEbCJeZVdKi8w9Gxx0TwcEqT5UnFvze
d/fgsH+Sv2OEoDWZwAZf2oyKzTKfDwrhZVxzAoY96sZPbH/TVxN0pquKBY1bM4P6
PZmflf06eWpSiLImXdKiTTum97Jkbl45nLAyzfUM2Kzphfl6cis09OAhOYNYifKA
I5u6OLsraXgttNp6VO2t1y18IgYwfI+e8egbG/j/9jdfUAbzKhjItSW0A7Hq0qQu
fuhbaxbXgaaWcyvK7p0uKQFzuJ9nrotQqzCO5MPmi+x93wpngWIf+9uylDRI7p8w
y3B1FeAk/nTYR/r6Kr0bdqXLPlpZT3K+6TJTN0JiAuUl6UeecSbRvJQTX5QoLO3h
XqcSj/kS4PyKb3lVIe9HbNo4xPprCSFZ1hLKAXyXKTzIzJt+Uur/zGO1v35q4yuN
tkcqKkbKX4tDw3KRpCAs6O+LeczScfp+W3rfuOeUw5nm1qFt/1nvOtyy6Q8IVYBx
WaG5Etcg8eB/Z9sFgVFR2Jf4tHHRrCZLN6qx1dYHvISnmR12ZrMXl2IjCN2EH6OD
slSPAhgsb9HElPsqRzJqbAC98pHg8WSRZwFssnUw1LPvOTH/v1GtSOqMXg+TL6uR
p8pElefJZXaIySaoz5/LMMJWV0UX3WROFOF0wGvsVyXFKSXZlcDfXIqnWscBqPEp
JiAooqRLyEDgN6xz13X6jYUXA9EF0rCjmaYHyA+OpQC+JKy91EqbDroOlL3vhYLm
DuaKmH8ZsapkxJgNRSDnFjupmUAdiR+M7upNM3TRcxzp5c723N0e09JQ58oV0kPa
+9XgS6mBr8jiuYQtzZhdzQ8DBaVKeHvambg4gAQ+7YLJrBEbTCZkiNmtr6b5Bwj2
6lVrCigWTycqBqYqcMtzibQ057FiIvXo9/SVxPeMVwt/RroYZX1HnFEuxChVOZgg
aWBRvz0g8G0MDBKirUQk2MsufIHjaSNAeX9CWXYCqQa8dfJK8sEYBVT4V8n/3eH7
1bEMxRk1k69HfDy7vX5tz8M6jGEt26ITVJgi94RQ3b5fxj9NPcxmtXPaNjTyvWN/
EF7poZJURtTEVvRi993s/BNUbaJ/5WlexWlM5mKM27VmaabtYhRsvb3vetWnMUGe
XoIGBvB+FiD7c69uwr3c/8+zCH0eenIbutHb/Pnkz8b7WQyp1Q7shYz8e4QdfDUV
jO3EvLDv7+qsugQMlEGAKWG/qj/BI190iMfXUnTvfCNwBumnVVWL/rJvhI5V6GRv
BT7H2NXWIyMbqC60ylszeRaZRSzKjSoeGp+l/KHn+azhh4fNxkZI3uSDjyT/JJV5
6mOrm9JgTHW+ywbqHCT7WxBv7u8DNOzriz6wuq8mo/ePWflOEX0Y/nPiyeHRS5FI
TtYMbSQnodraxUBQac7WIi4ODbWnXooy2yL2qB693Mk8BwSPvabzQ06OcB/TJk1n
/W0oaqKprFXrYeVusSqR0ktb2HIZqtMbJGUs5f0dvHPoArVHuwFh/cy9dAsiU5Cj
tr8vltoK0xKAKVwrzkbOrh+Cjv/JjUJcG0LZdGzTQkbDWcNlN4CLCBdE3nhLvkJ6
E1EFuehAgk6ADaKfEb6YW/z8zbMF1irbdPHLIPM/iT5HvMHOLW9UFO8Xwrg6UpxX
LGGkglsnUa1fuaYZrF8X4vq7C8WmsBLFwSxVk3XBk5nuTqLEBZVhQBEsTxHDuNUd
G/vjTr05F+RnNC65Kx8GoTm1/UOBf4VWpJb7VD+Esso5qhblsG9obOcU77P9Bkar
5iIlK5OJGiEP83o9mQ230WGuVT0N4z17npNUJl9WrG0fo3HxJo86MAbCeLOcvxfd
U6XgKJLxSlKxkG2JKiMywkQy6mwYrTgu7CaSVxTHb2ePXsjsm4inOQBZN+PewEfl
lGIAmzshOYwVHeotGYtgSjWryAx0dQtmvKRunGTsuli/+Pm2JLWYvj375ZmXkNYT
3y5V5Yp//fK6rU3hISO0VvRDfShNlK7/qnPXc+T5SnITC1jT/q38eH5G3Ql5Rtsw
/azYEOJCZpkAeVQcwTIXe5sHEQqfSD+WTXdalORd/6two+HKn6x+S8LybbHl1u2F
PQ+wEGMZqJyLId/liVGOBDUtQSOgT5V3klLaYkaGkDhE2gERRb+y9R88Z71l7r/+
mw2PYF8LDh9qtIT4J5A29ob1z8a7wbdfCPe7UHVr30GUcvYKeS9f1yePgTNuowcu
RMte7dmJoprXUbqfebPdtvMtAn7Krh35jHhAYSWVxSOQh1S75eljLWzbuoWxzsyn
c38timc0Ib9uCQgj0V7jgGyljy8tQrkwkzcTKO3sjGADXZT6zC+L6eM2Zi/DItzz
sOaatkM9aaqvCKaFEqb2v7CoVadBaOwY0dmER3PFPrkSa9GZ1Fo8yvaE2wpKi/f1
2d6M2hcrAK04kbV39WmtLMSywiLQFejOMY3Vo/xNY2jBnC+dg7xmWJ3gSMsJFDra
u2UsXX+Soc2LLeUNMi6LmWYpupyU1+cmrPdOnFSkbki/S5kf6FwQKCAzzIE/XkLQ
ZHnk3GNCLpCTgvrCkZNax4cl1a+zU/4hHKpgRBmzS8ua2tVgy9X5Cim8Q7zfHUwf
/eGaEZhkDifzdvITdSZ/8Yg2JdTig0Psh8fAOXVi04/zWJEKOH+oezs7oZ87KSVW
gU3Z1VxMtyNy0x8QSajksrbmFhvBNFu46VHsE/uwXDxLNPCB2tYDXw4nl+wI/C46
h57utyjTtVJicCRljBJRWENndDJ7C8pB6JDqRsvcf0xc3AhBvyrG4Jjoup4kk08d
pAcT0A9s2qWL2ngndJuvhyuGkKn4w7A6MwaNX+M23Zen0AbcgDQOZiUVYZfXEaef
M6pNJoUlGb1Nmi/C0e9zP0eptfa+7taAJLqmVSbNuuh0nAWqZIH0Ipk1iDlyCFLN
pYHhXDu0SUlLUA1R8uM0ZDJ4f1v7+PIsOD4Gzvc50eXwoOFX35p3wI2EHv1RERKe
4mrc4S38+w6hNpwfza/f38yFfsAwquIFKZl4bLbj8saINPzfg3q9uSl3QoK+5lan
sRiu77uEFJL1Fn+vd1ZV9i2k5Xxf3YTnm7uGc2GJW9XwHyUQ23MkruNmx6CrbX4v
btKu2FQOW/7H0W17RonyJY7VIkPbcyo/RwIPua817a7KcBmzW2uNH+Rbti2UutEB
hSR6Y06Y/4/AG7BlvY6ioZ55IGSGeXl0v4Wo/3y0AptBQZlRnG/sW+CXwkf7dTN8
8DBx08mSLYnr3/T32CiXQHOXG3CNBdjTa4BUijUkgo/w17c4VPx/DU2cScpWApE3
rIV+LmFzV4lZjeEBPs/G8TWQ9bgXw7FnvrXNpet+zIm4gGeFYz29a09VqHcRp7gU
fgZdEhDOEmL85juO/EtoHaI20XAKyeD+b5eGbqyV5LCVnmM525WXwUcaZ8B4H56o
50IfGYfPREZfjs5SfAGvN8abaSyH4dI3y2DXSRlH6WSVRJoPETktG9yyaS/j/UCt
4fBimCe158YU2VERTm3hglNLT8vnTrmsc/3ybp/nDYZBEMcmipJofY7QiwqG8+Bp
NjE7qD5chfBoIbIa4ROnGTNFB+PxYZ8Zg/vu18g8BbJi97TVE0daTZFKD/RTC8yU
U+nzG1lIPNOLUUFQgSYb20QACydA27coDQqmDICq52fvJAf8QBJNNJh7tD8sSryi
QYIbFmo6pzqtDhro+OgC6gRL3juMXaxex9166zSkzDYLi8nte+fz9b9Tb10uxIZT
J1klej98IFGyctDiFY681HYKLs6xe+h+bQnUW8OpzVRPhotc5qCBhFFMYw1L42NP
aqTT6mW4m5cdJcYVvwORe7GiCOOUdaqeiI6C39RDYvk+PHa6WdqbpFNzcnrrw4Qg
OJWQKYANijTbgtcXoueWRSkZKmuMbauxftlEMYGxgGF0MT7KQBuepeGQeChzLZjr
wV4C57o/08qGEunpEwuCTFKqxXuQHk8dAhEFp+9/kC9++3wGenogKACTzDOE8b+G
ukbZFaAJ+EILnmpOw2+tCU1yRdA4v5JG73fySkBuEKU2wbOIgV9lOXRCymWFUnNU
/ZzF/H+ZdGNcLd23smICeDdjzaDJ07SOqDst14Xawkuko2EW7zY5qgxlo2REansA
3AUb3EhlS223Nbw1GvMjSO5MjN0X+6a7jJddZdWpnTk4rk7lTSvqFWl0mARBx1Sm
E5tTVfxRvifCcYj2FXJa3QBk+WLufRmlFEOsDcHHxuMfPl6YZ9PreoGktVnweQo3
e91qPsF7VaUGkU5bTm8B7qiJC71JrgCDHneVkQPfE1A8FKC7TZGEVXbu8t6scld0
/geIgkQc4f1J/Z0xB7rj+jvdErEpp05UVdg5nJSVI/uDUW6ScRu5cu2WxhbQIOF7
m9oDyuXBd8HdAXHiiAfi9+kr6laDlWWLU9abHT7gimuFULJvU/RYfd8umN3UooFz
1L1lfQQ9XQjTlqYkM3MYExRKWtau9Dj9EjmuwtyOZ2ahTEC03bkJYegAJljqTIXa
pJEusZhe5aA9Q3yeM4+E/ynq/oVxVK6i4NVZ0kYQn6dc8DehrJMHbiBvzIR4mnz/
apN3blOOHg2EWre6aL2nOUPjuGCjJnego7VkvzhMxef49IOs3D/DZ9b/EY024akR
qSe7fE7CYsjp2pQcSqI2IF5HaH49eEwjhYsJA5KGB5/8ujO9+DuSNqHZpMtsfITR
srSZAilm2NIqHsQklb+pOFJgnEqS+Amzyqo+31vt6n5R2EQMBoKOUhw10Q/UtTXc
gWsbrkHPYvFVkbTwQzPNPQ+O+H2hPO/mGbsgBJXSfevggt5WjZ/RVAAEAuHaFtfJ
/hLyBSYoKg6Hx794rL7qmGHm+rl22jjX3OI1SidAjVTo2sAzFeMF/tI+t7WPKQez
6EH97Q7w7hktBnrOrXTpiTkgZWQRWkSZJZAJSu3VIgAe7vl0r4ipbS1uvW2Dsn2z
6jSFusgJ1o9te4eJp49C0SVLT+XVsUOzFxwvbmtKPd9vfGhv/puFi5Iu1y9272nv
jI0LlX51qzd/Far7HX3On7OoCz+wH4OsFizU7zzFJAiop4KT8zXImDrUNILmL40E
bvvnCli8hriIbMbZAUxb7W0yS0xARmpfeH4eVvDTSF8SQxnthak9HmKCFQp5jvIl
0sh6EfsoWNgsieNd6aubdqPHcmfb4/mIqPHlBZPNfe9dTLi+QkjzOMwbRamu+prl
B1BxjVzvsji0pqThNvq3q8Z2IYtYkza2yxPNQ/u7Uee7cTXP0T7r3WuXsOHCMKzs
qwwgWCigvSE+usYFM0uiu2NUqHFcNgvbJGn67mQh7SPupNe3nuHNOeaM3wwF26MV
RKnmt3LWR4KFhxSbl8TpZeu+JeX+rSs0ybveUSUyZh8k68n1vngetOxMfxrXu1L2
mzgt9KhDjRQvpLiDP63uFCL7o0s2KtDRRZHjyr1a8uDxJn5ytRwoKvkqghbfl59X
vP8E48eINBBFpFqjZcZLyaKPhIkZejb/KTLrKiFqKAJ6mpOq9VKm+ggcL202VzpI
Q9n4WY9SxPS43fmHppMI4yRUi99A2DgfCdlNImfgH3XdbDiVJclLxwsPxWYYH6nr
Gr4oGl/RMx/tzI3irRRGbc78VYSDEURjGLual1MXq7saxfg3KixnFLwaVfvBCibh
xMyKElIJEOdPif4rMfGHclCWhgrzRNd7Dj4jUFT97aNqsUDrHAI9iwmEjEw+ZUDG
JmhPRNvcfIpDrpqjjuT5dn5AgEj6i+jq7LSg9qylvbLOm2G1N8VjYPW82dZBnyEV
uB5wbe9pjRZQRXobAqRA92Ipu4XRdL/MR9E3bSrW100p46bgYpmTcM6191VZsXXo
VvXLYcVQcJKsMgAGTPT7NcOj7lTpCc8eGEnY3d7MN8tAQZpqtjqS7Z75Tg5Tt5hx
PIhgab55ttcEWFqXPZDJiHbLrO5g3Jnbdcfn5pPrJhU+EMDDoFUe2cSs4RQfgqN9
ieZs1q7PrS0dmDCc+gr3oY5p0P2VUM+I9m6kxuMn2Y+q9EjGvmF7i6tyAxLv+weP
5VdKGGlO3dvMfhI89M5KhDZUeDtm3q2ivKQr30swMF46omKGZArQgJln70BB1RaC
9UNK1aejBUb3P+AgRw86yFCwAXy1uc9pI6Z4pdf0XhdSGi7+cno/YCaKqYpszemH
i/h4x9VwfchVBtqRRSzO18OUa8ALX1nW6n3zxnHP9NjiKFEGxmN0pPBLM6Fp6jZ2
6u7j1QkNxjRszixp1Y+71zn82qlYGiCmSz42yU65oKXCC50L3Qj87OEu/CANQfn+
5wMyrfIQ/Y+G8cXBzmsYaQrIuKhmP2JuGZJ6PI7ObgqmmWNfMQ1LPyHG42tdT7Dh
Vw4nLV13eKSnN4yFFERrp22HhwP1LlasZrMw3l4rNgEsRHPjvZwH/9ePoi3ewHJl
bW4Jsb3npyOnu6tr0ml3GuwuCDhFyw40Bixu7UdcAyiWA9r8CLmJpyu7rmTR0K0l
JidNblxEYZc0JB6/FeI7xVxqUGNGXJBjAP+C29KHdNBVUiR6c1wRt43U18Qktj21
NWX80Y3EkH8K9Wr8jSvfVMWQyFg8Ztgn8lX6OWkOS1nqkCdz+kAqiv8uiEFIsL1X
cnWb7XqqGn2z542YXYUzyGe4rjNs3a9/jsd/1jdhtt7HubfhP5+Cs6hY8oeHKBE0
9zG4GPvfrxlJA0IqwrCcTAzueu+FUMV52O58EqSP8132a7sVTsIrdNVsfrmdQOV1
BlljYdeCKbUlFe+JfrznhfwGhVT2VQMSeHLvG6raLzzWnpxhTNXDf0vLqLPtoo0j
8v+qv1u4yloPc5pXsyw9muXK7wHei7CQ8NQKYIl1Thab5B511MJijDd+kvzwyJDL
S7lL7iGoLSVXdmmoQIBfsQu29QjNUGsw38ytxtvgBNkSB9w75kyK2Qy7jkSsKiNy
Uo3xbvtDj4kzEYtw+IZ0A7B5XTfuO5ArNbB/OEWtJfhYGbyfYlJekbjXecA92c2Q
sR6x9YV1QuhLKN32lqrlXQq1uS1xNu35X2fs1JpONrQTW3Z5+svNV9LnmbT8bj1r
rJ0LOKeQZC7tE+fh09MkIIagtAXC6bqBq3WE9kWYi/sBth1aWVOdkicLCqQqhI7T
ndz6YsEUY0M6tGGvXPb7C2bUQp45kieiEd4UjKIp+38aPlvjAGOIRHf2bXK1KOyM
HPSlm4xKH3/LjzHC+xhJuHxx3RFFgAA/Kdkn6fSvO25KDmtxEed1AtBMN/++QcgW
+sV7l7Dl5bzq9K5AgubA8o9P4A+eOMKF5t4OqecSbxJa24dVExORI64w4Au4aOU7
yyaiNyZcRTD/WcL+F5bov3998A4QsbphmMbkNLrCF2xIr26Nil9URzzVs6EUmfMf
Hp7xpYh1qO+6+pSrwvb1OQr51SxSl7PlJA/ZQMvvAgDMQeLUJX54VbK1CbRhQAB4
TZuVEXrYr9ZNxAL7g+TSJ7MDCq+K9puttijTDHkCraSLjmALEXor8UTk0ald5nFU
BPS3y9MBLIBypGbfTgSzn2yYy0kgimQe4naYu/WutwUpj2+qVVaEXdbKFdwoIDo2
UEm01wA9JQ3UHa9l0WwTHFeJRyjCbGckNkqocimBg8TqkIdqgqkOKERJjMjeslJQ
RIXC+fHqFfY7FfFa+GUOCByZB6DoYN9z+xxQ0nYok4oxF45zu1Fk8acyGQjIM26I
9p2pAOslevpqqWokIPwRzByWFkundfp8HTqitGp+oXivGZPQkSdnv4eCRxvSY4sp
RywOfVuE6Rs9rWo0kOJ1CiBmIXURTf/hNMpQilIQhgO5JxUsGbDoXxOUR4XgAnQu
v1XloMkyIMctRWNguuc+RYTK249GPy+Z83Oxiu5FWjWaThhdeUkIzb+3pSSkpUxn
iMyeZx78Pt2/tzx2uiBiCvt3y0lFwHJ1CXZTZIqKpfMZdij6nwT2/xuRid/JE8Vq
4vt+6MHCUBeSSiNBy+jzx3Z58/oA9132c99pqgt9Zt6QnmHYJD1YB/D56bfuClWv
kmtI+dshPZJODcI21z0r1EV/lejeAiXrh2xAqLN8CqJbeeCyJ5/Wrx0VQoU4TxH5
5v73doB8kRss16u1+pC78byYPOFNJCYR4uhEbn1VkXykd4KGODi/aMJ/69ZDsKJ5
5yU/8A380btfstsip5JMGh00vR/ENFcqwvBb449sn2tAPdhNZwfJFSASPamRQLDu
y1YizG7ufpZXvFzZ56OT1/CBB4E1pUQWfS2TxzbQtD1BZrxbvQ5ap428GEA0ZfTj
4nceDIFviUyswpIJftkDr9D+FINVgnpPb8k1Us9orgZi9SFjr3wgdfeRaYNXSKUD
+RRuDWTUSnK134jq+SRcaoX24Fnp930xXsb5l0++2XsYDufZAfZI7jWPh0Iv9yjW
lw1PU4MezxL6CqmViNaxyCBG2Jt+4mJ3cjlQphGU90DuQmNzW4jXOdUjMH8HOIzp
A2NbnTESaacGwh8bmi6ctzFwPvEkn4yZAetAURENzgvE/u4xn6vG9/HG/Ll9WlJ8
t/DaI0FWi782hnp5IBVejkyTQP9FGwezoA5pUN6y3biZsRHxnbbUUQ3ks67aDB7N
7XwmBt6YxG1wC4J29XH4EgR1B+hD+Tdvb2iKrJ+q5VAehJCtpYjgHSHNEsUyyX+B
aRdYJAjbd2R0eSuUDwdN3/NsnV3iPE5y7hUQLNJp5xjxgbwWjRWFqg9qTj54Z3E+
hCZbnze9TjXaelHnmr2oyrvl6XhK+uKWUoql1mviA0A5BRfqBHQV9BYaCZB2XIZg
RWI+WqGjL1jMKVXV/HLDCkRt0vkQ+9mZZ3TAQSBEGZ/75PGQRAQSbttMWUbh2+CF
zfA1JStxY3jv3vWRiSJQDyiW5x8J/XYHxllRkFuZqcQrGjEq4VV1MLMF2ioLo8oM
nQ7GhvXbGTlGrWzQsMOELXjqR2oMyI/hPK4/ijuOygJXquzCp9ay8mjVI9gdRdgl
Yz+8iMQI41U/dBXCMe1WosqKVL964Uo1TYc6yKn+NsMNaSEy93uy343I4Cytr1Uv
iYr/VSXYrXaX2o2gzMOJASATKUqSbrEnphlKiVAokczPZm2j8u5+LymbZxZnl3k/
c9H8OKAVjzyEVrFnV3Q3b/2bzxlI4a1sAsvgA+lKldS8tr/V+9NMLUyEs9Klayzg
6wbmXSXFaCyahLXxHYG4nWVp2xwb0JwE2NJB2ZC8Fz1tr0r+HtNUgCDJJn+rsf97
6fWsnxhVO1YGcuJflUpW43TD4VoYYquoXrTOwR1NrTPRmPb1GtO0179jnrqEOQM6
jjK05LGMmo+J0nyaVO77QQA8WCqbrMMwIHJPeHYXe90SpVIbJ4VpNSUptchIl2Wy
EjwYYRovEuKejIVKrMSc5HRmHCWMUL+838efuAw2VkTDPI6mu5efYpvPzqy9trhS
9BYOg6U0umwqr/7v0t7NX8bRzHRQvD8XLWMCG9T4SWdcURA6HMqfX4Hwy56D81+z
5Sx/Wx6Gix5Wag2NC1ocyjpE+htWR+xsA8o9hIvlJZ+E5VGUSdMtMwIfZhQtmnR+
0FRZKPjStz2Z4SLch90HqjC9/72PaVg5N35qqnjCbDD0oxmNyds25J/ibIUHtxPg
8CY3bg49ISBpxTeLfX4+/kgAqyl4GL1bawne6jhxC9pGXHE+HFOAy7v+KsnYmD/V
OuRtFe57yn6bClKwVcD8FHsLWcAUkak2XqwOOCjhOX2//aCjWJRoCAOEw3axxE/n
1pwKnioY9xjh6hw/2IONmwFRXdydKyNTS9IE5eS9fj6U22Azh/Jmhsrthz/s+en8
4ecnoGSyiSBl07YfVF32MZ7O4dF6G0ltdXMKCokZXQnOlEg03ZxGTpaBDdukdqvF
q+bnRZEPDEQAXP1Br4Z0/NV7eAFPLStChsgq1Wbb9Pbr4xn0qSp6ysEWeRF9+yHa
TG+0RUeWnJpI1+noex+CL6xMq6P9B//GI3gUKLMoxZEB3IiniGN1vWdPiRA97BWH
6Z2GGTOPZPVUyXarJdlhqXTwc7zLHEyc9113n8A6jB2btN5Sq+lLyObJdUfbGhiw
2VCveBbQyXWj2u7sW2c5Wqvk0WVAzgW0gScpKb2o5N1zvMZQZTcrcVd+mESGTZpE
fjfZbbgH8tfv8BQ/7v6HufRv00+RkiP0frikv1AvN0SWF1DZ04lDoOa7QYxAH9Yz
F+/CHXP5j9ZEK9Nua7DdJ1pcYqb5xIKBAZPy2ihs8BTvkDr6OY74SGNbh7I4ksFG
PLzb1D4eCgGCrPV4SMuwG9IfRfORxo0XvlfojLQPjxStmJsUMQ2k0InUHFc+Q1At
u5pEqLiwOqbNaxAbqTdIphGWubWVnEH0rU78hCGLvFqGA21p17Jhq2lOQhWOXDai
cZkv+H81mdOQ0ITpvP+SYWREPIMebf/U4ArcKF1WhA0ZB0Yj/2Ss5Hqhl122gYOy
S1M0PVoocqqW23wuu1cp1sPCEzItf05J1bRhzfSVrixMQ5fVdyyQ05Gh8YrvXV5M
gQIT0dWAYup1NHfNvGygzgnNu5okiK27cKdS3HaasWEN4nPbBmC9F3fXL5MJAVbt
fXUxpt3uKz7IX/WheiiS3RcX6L+0NgK0QzuHZYRh2R6Btb5UsQqfKwQYRGD0//bz
96lpqlJyojyQiuzsjd8FZ09EUlMxbnVXQFxtTwQb1JcrZBnAB7MkxjIseNRpYIxy
pfaz0561Xx32IX3cqaZom3vkVftTuFlsotQJ9tTdy589VBxqN1nFwFbLSQZVj4XG
z/2DYZbHj8cbBHzyGyBzaSgllcJEnkMLd8+YzGqpySGKqsuaVRMHjka7po+7I4Xg
jf50TQ60Lu+ylayLRAP7Qw1YExHNynx6JH6HGKW9rYPGqqSAnS5hcQKMxgJNy8Iv
0LYGBgpI7Vv2kt7ls9RI0iO15AmfWsTTMN1RO3PVyvELmk3swHFmQqcOLr7sVP0E
IeO5l1C1u7aDUsxzOz0h8OYs3fxRa85jE4IO4NHPBHQLSiRe5La04gmmNFc8NrBZ
oCs1SYLc/IzQcjPFhBqqROxkqPDLm7byRqxdcQlY7A9Py3Z44yhcv22cFCKTYxBH
1nz2K9g2fMqGPTcut1Ro4vsgp9BUa+zdQNvs1j1asW6moyWe40C3T5qz1DxtkTxZ
XvkQCztlPEBPedOzxFkOICQqxTtWg7SJIK7z4eMuX8VZuZkMEvEQEdQ4g6qVLciG
xTKNS1isWpV2QEAj3BV4aUbT9X3MvI/7xVHYvV/COBweK6II1ZUIiNyCCSbHg9xX
/DfTv0IyEdkLGCXrd1eTTXZMhHgtLUL8v0gazp2UWXPXIsrdv1OEizvm9rv3zWt5
1LK/xOBAit3oIZm3a75bTvPXxz0i0hcvKOHZ7G47BObwjyNUT9Dgo5SH35zZOP98
6Jxycl4Babx44CPoUWUfBJysyLGyYRgzfy3tZNcwwMo63NTngejeJlbkUb1r55+N
AcA1C4IPnC8zFxvIYy9nDzJm9z10wjID9pmfFJPW2xxQqFDfnSW1Lv4AVblJymSU
C1CToKPPQ8qWrtJAnfsV0aWd0yCHuRbshhqRvBloeHCP7pGKBlvAbDLNwb8NOG+S
NRxn2YYUpsnxA19RgJmIgFrOGyIy7HJz//LNp0Bj62njRTTqo/kaXdhxIG2UueFu
vcAd7L298lWw6cHUFZyQoELVwPvZMisUX+dsEBulr1XDZz9gLWpr9xD6CsidGpeh
uFcsJgu9oteOgjyqzcFbioYTTpJppOiW4GsafM1O65WNOM9divZoVvH5zWi4+7Zz
GhjH6OT3iK9xG4jxxKZ9jzWNB3WHb+h3ms5pU3I7XOJXaVRWX/2hAu3EPx8FUJ1e
55OGi0U5BUJlPVI/KArM0yLORs88CxTvoWW5HlIau7NdVO4kdtkT/popqWxfkfaQ
s8aJXclK6raY9RwGO1JrLHLKfzv86M/0dQh+1mtmJ3E+ZGLSGU0bSRWhnWg+DBAl
li1RBCGbhfCT8NSuiKvfIfa5DIZPHLEsIF5rUMqRceztG8qZ15HhhUrTL8Rf/L1F
E7dPUxUVL6IIs3LUwX08XW3Iv/C7WsLbAzKduPncdBIkWQD5pT+f8AstKb4foY94
oBtaD8Fck7J6O0iSNDgu8f6PLQYApgzPRAf9gcuhEaV3jDf+xeeuiqKOc0S2PoWt
SPamiKU7slKSXWId4rQmJsbiR7dbQAkv6yJCbhIkPJaMYTyGh8s6qnXI53Da9OGb
FTbZoNhdVzG/vxp9MMwd85bgHA5yszweMj9NpM2Euiph/13Mb3STAv9+oAqtEaDo
BiWtm+y7RnX1QcZrNFOFCwfTMpk+rtJDRDcoVUVSZEak3wpWaz0sMVwtiE5tgdoc
j9609rBHXb5fhwZlXVRjvedZ9dgo1/vdhtVNPJ0J/L6P8W5+UtwXjtk64RFgV/ku
jK9m6uS6JfPrNjDCEkVHs5GFZbdA/HM4YtuvlU+4W5fhaUWqpoJXzgBvgquCp5Ap
Qh3xGaKZA1rb5P9gurP1pB189roQaA1rzmYHs1kvfC+ahRzVX51KqYvaa0mOEST0
t1VKGjkY49pt/zZm52EG3b9lvYAZC/MTrxwVCPVVe4DffMfEY/9hrPmcTxyzmHAe
zKpva23LJM1wsnv3cfC4cgZkspVSAfNSBDKcAoKILD9DuC0vw8pYYDp8If9coqBK
o4x7eefIY+yYJYaTUvPZG1e7it/+DKCfCdyC2y1TAw8pAsxZ1T0cUdxBcRDEhqZ3
05h7+IsWmhB6EKVFvJ2iP1lUNNhBhE9U8ciQ8TXRfFn3TIU/4Ch8JIDOFKCBcXWU
CQ/79763LohAz6DVgaXVAtjWAqD76U07H7KpSqwiULaE4eCQ2CaSumu4Vbdhbqfb
PKNqwHaW6EBFWnyO+pqex1dIVMwPU2yhYkzaNPe0BvYxcG/5Fhvlx2+0lc+9KyUN
VTIWUKpTMpaFOzCFgMjQT3axGf1nysfdTaKPiR7CdEYRRhJtc4JYAKcKmSgC1GCX
IHFN0jaVwN8hGPwdd3xAhkL6qiURnCr7mwHa3t00YzRKLf+bKenMxBjAGB0vkHZk
YlRuVn8BD9kBInvdrEg1VytUnoTjws4WdKaLl3Lnz/Vf0Sqqf9heLi0GGBd4WHun
uYCxre3N8pAKnUvGkrObWIFWtqsoVcEfUbb+/ZTDiA6JZtU9LE8RIf37VkTd0SRU
aPZt4FwRXI9KJuqOXoYhvmd5bgo51gDwyrPm4x3Ooj3IdprI0MpsQLr8gG1O3oI0
J4Th4swkkKP3EYkeXyQdObYyZ4XEeXHJQMw1weQED2Q6q6LEpQ4I/yeydb5FS2AF
PN8EMIBfIzezyFK2ui3/4zw6uUxYwh+TAh3pcKnuTZqMFDPyYHE3N2fH3UPQEBoi
hiHZaOTFkMXswxFwvxLSXzpKB1PKzTab/2EsaAZTpIowS8ixE8dTXMIlRvTnugrE
enLt+HmrTXyqAEfzfVILW2MzB20uIdp5+xyojxnaXBzjz+lE8o95f3X7wOBYaLDo
EzqhBA8953FSdhavVQUPOfBEiSH/yH7Dx0EqCDGjkQsU7BuEyrhNgM8MJOTbqVQe
BqHzMpmc2Jztq39Lu3BmrLZwhdH5fKq87bgmHBypkAgJC7rbqKPcRWDtnjB5doSf
rrDVwr2B5VNlxH0CfcRqdt+FTbpgRcl/yXOhV261FXMtrqL+EaSaOd3jxHvIal59
PYEyBH64sWEyFy5YdvxaGIEbdPQWqVwi/3uKbKlEpPdK1v1GRH7XDFCBzsLX1Dzb
sumPIGDfrswmS8G8RVlR32Q/n7pDb2aj+z/hcdUfFUCt0udVrCFUaLtOsIbT3Dxx
qwLiTvj5l0mEu8lzQNhNSVhrdm41II7UGyyDblg6/d6/TDqL6b4dNkNZ/BLRIC0m
CQw3rVttsQcIEz9bX56P7YbsJokB0KEg8gzjKJ4nk15AzwlsqXGkZ39jQeVHtYX2
+2OQd8N5Snv3wbIRywVd0sPtSCS62veX8GTjFgdihn0bQWmDVj6Ukg6EjLLrl/Ad
6hYbQd/dbD7HHY3f4eCJZRXtXgG8dSle0VTyu6NhmISGt/T++fEYQ1kXox1RWB9a
bSXB8RhZ1F/4cYyTMuvpNtITl1gg+m8PkeJvWhaChacE+PM+0qgndKoY+EHmV8Ae
m/auaBwOGMwb8F4n2DJm76DLr0ICV5OrRc0UuT6cMQskoE2m9YicliMRlkJTuMuU
IVQ8pvVPF4mRlZFqEoYEQTfQJ34iJNKTv58MFFtWWJh37ripbeHpAyO9crpr8HIX
BcPbH9AQGgGflsbjB9+Rc63wBnuy005c124jvIZQkjfw5PrJTbmLaSquvEYMg8S9
gLCJ++vK0dClQeRZRzfrEG7cePzdGQgOaEJLXyTrwb5fL5lkvNVxFOJ+j5gCTmFQ
sCHVwquBRfN/pTUu/AD6IhdMnPXZ52iPc4ttaMYgHpKnvnbZ5wmzlPaC6cqMNBEX
ECw4SbomBWm/tQrAF85resfIuL86kOMw8VSn3G64LUtoBy2d60h6HaNwzzVstNYb
SvaV29RyFrfC86O9QwpH3HckrmTfDBEOgzMB4PQfPSP+pEIH0unB4GgBsZ/I1RKh
NO+7GKtLt4dD0REKmHebpHzsX1ttcFZUwPZ5cJq1iwE7zsTpmawohiT390AjyG5i
/Gfma1kfPEGYm2DFrv82AfpbcGceEuyeAf3ls3s3Z/fbhh7YhOwJqt1NcHp7cZ8f
XWJtwQGXolSs5XiroATXQS1xqDzvDioiWfI4zsBuKHGC41KtU0sOJZklE6gCKgu3
B/imKKwlbRpkd0UQbyfoqmoENqcuslj8f51pDGDPzAuMUzvROCEiAO8JQW41a4Vb
vKhbk/9PtSbhjYuI/+JpJ3zxy9naRW4NXwQCD/SiX/v7P1qsO9LwWwB82Z3qVcdW
60iFlOFRgmNvd+IP+Hr5JX2ZssBmAA+qyZ7Z9MBcem+C0YfsfS3Jx+lDfhNbdBPh
eBe8CfFc1r/YahVKnElf/4pFb9ha3IUt5RuJeHToB2CdKr1k37UUe9JbV+jG1GsX
xdv3J0jA8LAKVfUten3tSLCty+aG8sgukISUT55yY3oEGIrGrfHsz3/WURmkC0Wu
734YELTXtBSs1t2xSsPzsMJI2jTPF7WDKTFvkiSG9gkiYDTBxU0O61kEFocVoRiv
A5q+ol9G+5G54/LGia1GbPJ19wv6quEVY3gBuexNJ+tN0w7CsANEvo8x3RQihYv1
DWyCYiROSalGm8oblA52bDiYimBih+d3+o5ITsiEmzhLHZ1BHz8AF5YreUnKwA/Z
WrdZk0OKycLHD16oJrkvF2p03zvCbuizirJj3aUVsFVSViSa1Umxz85dMzIkIbwC
yqGSM8Rqf6WbKCwcHADVwaUpm4kVFD9jjPFDtwCzWlI6MnyxlND8ex3dMzPZqV6E
aqDNa0Vz4uNaOYoa91JSV9/d7fkR5nzn/bROCEoinxZUlZJ/yxxDIKB3YZk8UcI4
K1OdMDR1kt4owJHuSYIyP9Lm1NTqLg8nhcqeOJHpOFBp6f+zphytIRveb7pT5g7T
XabuUcvKlEmGZndOeJZ5ArnQG6Lhk7WqNEFR+MSV/nQ4yPSZwrYzuRdMp/W8ZWQ4
1TouEcO5sy/2kJhA7E8MrkN4u8Simu2lXRUcLwps3TxlMSfE3+kfbq07lBinT/2+
jVtgLyLtrBNJ6V11+PB4QWux6I7uvZigKukOKEY182fc4yS52P9x2Lj8K3iOZSph
mJ0Y4gJQdzfiVr24w1L2l4xZXtZxm0q2yvMk7/bC8w5NZw6m7xSh8tJw5ZYhvMhh
8CthrZo+rxZVC5G8D0diqmFlGbQjmZnST++/uaMFjadq16csa+gZsulkYfE6SekZ
jWLq0ITIQjwWmFvRZmOVMJZA7k7wqT5hSlSc7pGJR0/lJaTUdC6CXb0zU6b6toad
eTq9uy0/JFBlF6II8X+iBPexmtK/S+Wn1W4m0HUUcthVWhASxmpZZQ9q5pmEt9jI
MgFejiYexVahkQcDTezcgef/edWNuBxtWXZC+hHy24GAJVFNowJZzI7jIP+a5cFd
Y+nuEpJEGWzhUPohhYnOWuFto5OWXra6kZ6BQWtudIVQXH2+ZjJE2QwpfjZDwBj1
AbIfTq/9KOMLD3Zz/HvX3E82X2eTuG7UTRV3RFGKIJvYgenHS3/5o1YlIk414MGX
CE132MZCTuaJV2bfC/5oalNOaHHIN8zZPSsBWeUClj3D0x6bUInh+ixi1Yn0nsI0
mqvU4oSpO9+y4CErrvhmoaSiz9AnWgzOs1YcOMjG0NvDR5HNMYMkAAecYY5G7J1r
CZbtmOrUXNqmxPc1f57z3Uzj9naE4NomulacwkYzpu2tWc4X7y5gjKtjnWFgiO8r
cCOMo/7glBKyMywqa1JnNnZlCR4Kq1aFab1rbc7UInoAynbCGOMiowrnSJXUNz9d
YwHHGyIxRWYvcoTcs7ZEnAKYYECY2gvMcOP54AXeafU19AsLfvDgFeL2cCkw8dqi
qOZxu5bpOyff/6aoA+s75V4xP8hoCGZESPdKj7MGUA7u6N6ArjP5ifTdXBcgZYzL
E4l7kNN/E0nUmOmVw15VrxohCvL5wG7PME32AmAldVs9/DrvQKVJvNWr4nNp5l18
yPfsQ/v39lqKHN9mVkOe96hGWTM/4t2l5fvWjaBEjwoRIUxyXz8Fe4H+Xl0h8/xr
IBGppnqWt34uwaCVVSCxuN9WkaBRV2gLkuH/0RMNdx6h6K8kKyQkqyP/WtTY+WUn
NOYfqzJQcLeHIgti62Ou+VxqIuB99Q7SW6Xt5txtMDwjraYaqwS6DaBFCnMNth6o
Z9uXmE5ZRecUijx6jjmxj0WWxVePRcuTpOgcyN2+jEaugwJEjPhwTacINADtSu96
ZxBcjNBHQybG1gBOdlr6gejFpRi3nK0ZGMs9hkREEjqWfZAWY2YMmCEHaplTk1BI
Bt2svra3yFSzJVO0puBHmDyn9U4048rCZ6/YRkpGElllDK5H4o1GQwYlnZB+b+Ha
gwIXwsasO/zkFz6aKd7trjauQqlNFyaZdrs9pvR/OK7YXyPeMgno/sMuALYxY4BR
5DcK72iMDWTw7HuVdX/Sjk+T+GhPYOlLRyuw6iSB6+pXuzUFQrhZoKhBzQ8IFxSe
dfG4updhKbyjDcN6VFyW61IbrFmZyi/p1gY3JYWJqSneHFCPe2PkyFj2wdb26/nf
4VKamho5c2yR9r/GswBktSB1cMhIVw0h5DA7fNBLzdLTeve4jbopTnKb+/MIDFfd
jUT9zaMdk6WE9o8pEu8j2OuWporEqd/5GCpq6oM+bsqOAcrNs3LK4bdHqHmgOFuR
03o2Row/AhUjusBi4jJ9Rx8IQcsq3cAIgkZP6FOanGck4tsXgT8AT7KfVAqT4IMl
Y333ohGyQXMaFx3+zROGUXdgKfkc+zJt8DdwHDzlUSZVQRhiNvKmrxFVehQpQNPy
yc8fZwj0UmP9CVzggF0hc58F5oEsL/aPXOEfWRgsrGWqtyuwnj3rE8GzYdTKKeQ1
ZzhPBNrIQYgBpqc3gqzXb0nxdsfHIUOShxbmrfW/RpBblvTINBYsM65TO+K8VwmB
UxhCw0THblY9aFjUP4n/+eidZUuzd+7xBVz1ablM7ihH5+hEq3RnkR9dKlcBqQdk
v8SGCRZARcdf8AIoz3ZqQyDBrrthFZO4H83mne3P6Kw/ix07EkrQ/chwL5VNkXXd
qaBduHD4ixETYnAv25cl4azTWYu+ooLu293RQ/v9XTpqZy2AOoTxDgw1V+kxSG+v
UddCEuorNKzB+HAMC01BbRbXQEAydiAS8HdNFYkwLK9Q9tFRmLJjYr96jtJgkU0M
tXzalSCsQksTpVmDSNtXC1R8PKzukGWHJzSKuEgN4CMBKRa4W+TXMq138blIiBz6
+l1RsIbAsbpNSgwZXbP1NbLO9hNYc28sgAA8lkOvYbyRfA/RO3woHESFwDr8dD/L
iSqTJ+evm0gl+ApVEtf28/1m7mMBrk5ybnTwsMtvOm9wxK+NFlyS41fkm7Evlu03
vxdnBq0fHLyvp5u4EliqZOCVnUcFghaESU9IkKLso9GxOj/Tj56nCN3PhhXg0bzV
hg38wTGjeVjhRMWmemW5jthUyLhuR4hYbeeFmNAOjjUDa3g2s6iO4SekKzcG+4LB
WG6w1ceZEwI4TUIpSqHkNzNh/qNAF5aidGW5Atou25W+TiemvngLIoA09m5JOWZM
rLCAi6iI6D/nkyMS+Qo2T6dCe06Ajn0bojg+koGcR5HNHhx14wmQ9dtGL+O8YkWh
U3TMaTOmCyEk5CbEIjU0leOguq7NbPhZeiOwPuXEf/iPADKxrnl6U4kRFDPTCi8K
8qf1LVJV6sCuwqTtS5mfdpZW35CiP2wcK7EkG2oQNtOZQrXlttBy0PAGlgVXKcye
HAlLZZ3QsIJAIFBFqpArzHTEBSpKXiHBxs1aPFsFc2QL5IITpy44XXPdKNvC0eGT
es+bikQJrikTGCdUubbVXW1/FzTcWHQtk0/qw3Hu/Ce+M4Kn4nXrdEeuPNQrHiOp
ci1IfENSf92w1C/lynWia/mokcihxfQPnchx0WbzsVPR8VxvnTM64mHuTCVM8Oso
55hBpLTOb+P+8SozPCPbwM4XhYd/iLhj57VocrGPDs7JvXcHlp1y/cLZu8Y9vyRI
fJZRliOgZJWzj4wYd8ASjmjEx5JUEcgWmH9hbQvCNod8bFIX9NyqR1Mmco0EDkgZ
lLz2O6m6IBE1PNDiWsWbn4GuXWTqQyPHGumKULZq9pwPdnj82vg2pILJdmkgvyL8
LSAI/P9PIkmdEOG/zjmcH8i11g3p6aXWS152oMKlpllejbhfDVpouBlpVmGZVXPh
RvNyvFP41A6/iWxCjSEXQq2RTGxrIOnLYr2TaY+IyU03z8RN1mEoFFl3woChoHZU
SbYmWJG1ohS0vS7qIAzewpME9Xk5IBZZSZHUtbv2j1RBBael9veydw1AE0Kf9Fk7
bE9fDU1yskeGO67rKYCrTMKML8opCv38eNzfUIyszoVO6dC2JJCSG9r4OmxKu3p4
Zgiv3uhBM6URpqt6c0Nsq1l7CqxznRS9TtlwHxfW81wcwYC9Dw3BpVTFaItGyh6m
lchnFMFC9JpB0wIVh2hVHMGvhmTJ1wKz1+tTl/Wd1j21/v4oZLwBRpOg/PH9RSP9
A+6T0AXQc/RwQt+NRvkZqhNuXNr5HPi+PKVX8OzfsLKAIWrUuK5Twb7eRaUeJm6B
mnyXj86Nb/zky6GaifWN7VjYk84cpen6kbDrzVRkIqFu8+eQ60ZzZ+Xbvsn7s5qR
A0jswhTl+rCXTKFHCfyOKUrFctScKNXTA05gZv0Bk2Klq16jJvRq9VxFQiw3mwR7
9zJTWyalhhpxBV1O8A6fde6kEJuyZL2lNguaRGvicPdP2L9c7B+7BSj4ukDgleTy
jYhbjnO4ofoMoWw0w3NFq1rUtDK7GvFiladIo7/DuAF/j9NDyd6TJ5rQ2rszhk7O
JeNq0aVrj+uU5vQYykWNUe2A+hpq0FvsUh2x4//8XJm2nDlJt4hO6R5vmFtOORcj
CtRaXhtNiwysj3fUx4E1WowaUWMqSNMcn3ucLFhPTT+A3bL89yrNMPOpmzyCpHZw
/GT1v+Prn8Y0ocz1lm4rCwOsc7Bm7exaAT7bwMJ7mMvVkvGL96Mq2S8snNyTux3y
woa5c3+sH0dLlX+gMwWTlDBB2/ynbEJl0GuK2IvrJAYZ/MSmsvKdtPMcva6XtCfQ
gYIsHoKzby/BcRstgGbuKKz3+eVBGhEImY/RG9mDY01P7TPv4OG0doISa5dvTnbl
Ve1otg/mQ9707y688bzs6yZMLlIiCTKaduPuriBsTNlHSWhywUWnP9OCQu9bw3cW
x48HEZVjj1b1JHiBWtG09qKbOp1gGG8TClt1NraPVne8okSm03p5e9TsIcDuWkbR
nYdmRbQwWTpkzZjNaf1S46aMxZJFj8GFzYiQSZmO0T8pwLQ+74s4cMcVEzH1f8if
gS7+YKcjDPpPMv8B9YZqX18AfX6EMYUYRYCPmI4MTSR59wySAuu2KOPDlzbLAZRZ
+DmQIhA+s49G1mqtfzNwbB3+EuCAycFB2I8FS/Y+0S9tqDRyIYRwmC4sfSDdD8pn
ycPRxSUuZC5thLHfid7ZeKLDrXEeQBdlLQJLR54G25Oduf70nYt7HlDNWOIde+0b
SZ5Qrj75kFXZ84Rl1wzvw+W9BasSXE6zVT1s3fzcTO3D1M9H2oHxGTILA/KiVybu
mMXcfV3Al/TmYcdu/zzDXn/XN4dPUn1ZaR0vdminrroJ1C30b65KjlXKNm62MRYe
fM9Ut0h3w9+gMRAZ1JcOxOKKlLtGivILPRBqGggJHIPuL8kR3bwTZ9ORsFiQwZhs
opGRO9dcgeclMwpMBd9+aP+ihbf4txkQ7z+hM4ntKfDpFC3HL9G6F3wuSiXpY48H
1aDSC4170RUGFgUzXUEjQufYQWTuZvd4zzIbt5geXfwLDi0VcugIBggbuAg/F7yN
hI/dW8MS9R1fp8Rq9w4TSQy2ewoW30as9qzWv9Blcw2XNJr87KWPHCW2rYBTIMiY
huKJIjhftqUDtnnAPH1T36UFZok+Q2ZEJ3ALd2vxl0EnMyR6ybFZ1qXicT7grGJz
FYDe2FKLC3OPTK+XJYPDlf1AJdLJ9ahI6XnQBQt0vEFKlS9dPy/2J35uCn0lnmCI
EsbZqfb8ZvO2w3O4TWb1VqpjfIFlftIJ6jdHWGdUJIN0Bwjt8d5GluDTY9vp0DTs
4/VzRfYa+okY6ok9kYWLZh8aM+xSIY6Yop+eqJsSj+bM7/nW1nTVg2z34WnzbX+k
q34dXJQQFyn7NX3uyufaClx2oDuCUq3OCf3yDAlY/KhszXJvmjHPWR3+E3MgTw0b
T6V8BU/5h2Y6DjcwexMephYTsfUuvRMmTmOg609LsJbeejhCj3h+09cqew0Wj08q
d1tq2VvIvjv5CgxZxBKoXarFdUewx2WNJ6bcjePPEPM1SZgW7QpuF1GtaO5dWn+P
e7tGVBCpm7hQ2ItpUSCedyPgHRDyc/qcbH2c+0qdCdEBe0Wz/Hps42AfKYIaasGT
jsgTUVqEbvbxNm4NLhE6hV3NU5jl67YdY5ywFnez7Ss0Ks/qga+voK09JBzhHGda
Z2lCoLadeYO1mEj0qaIKvQh/nJb9BfcfHkTVINFznRVeZHmtWLMFjRKQIIuvyNg3
`protect END_PROTECTED
