`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGWhvcjn/yyo8tKVz6BNRTpWTa1B1fmQJ1Uydsb9rzqt1Ha8dCTtyxqHzcmYZuE6
K6qW6cmPnlKex8bcoS+0WOtrocR1ZQgweB+CximZ7PbBe2xac/8ehloleBfZJV50
zPRaIvzPumEWUGiTxUYr2T5qJI2bA6rFIMogfZfhFfSuhgJP31jEdCC36Y7xYivw
oWHHCBOja2DhEaarI+CXXoQGqHgVgi9Oda00YTwaHNzck21I4q5sKQvIzHvClwFG
Q+pFNc66ECVq1h3yBzGYpDhbuZtTe//NiC4M861DmgoLVqEc1glRpyzPRAddtC7K
8MTpg4jP8PumLAXxj2KuP4391vQvsRbyNU4QsdfZnVvw2ScDp73NMUa5pGL344yU
xxeDDhD81CciRQPw3hutnhoNCYXv+mPUXnUKmjT9R3okBzAl9SmhBACwqD8W1QKN
7h10wUh+G5bdgI+LIOLH5qM5sNr18Z6ouyqdoCGHGTnlaEsPbshyHdQSVSP78FTz
mucDW5QYVdgSInzybcMHGCzGlIeF2Mkb1FfUIFsiaQVHjvNtDO4u3fR/l6s6/3ro
PcWLQURacLk6nAwkj2do/arUD4Qbzn/qJwrd6aOBFKYgdNf8Na5seCt57hbLwkdM
dxBLRJNHYDNXqUeIVOS5hyTfPpZgStw2XKMjXfanBGuIbE9+v4k+Njhaq3UTXYOO
`protect END_PROTECTED
