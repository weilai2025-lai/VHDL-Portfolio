`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LEg33tFiUbzGkBizDMFpx2uv+CnN/A2nQT3eV/7oq+mRQKRtSstUUIuIhJQ9Fmnd
EazTTKN6feRSSbvTq06EDOpKqLo4ULwT7tmeLy4CQRsVwmFYcRAMG3KjLuW6TYen
KpTi6hlnDfrUfmYnv3HsOEmKDxjo5+E+Zoq0lSqovsPrY/4xoYw1AW2VWlrbDlgH
BL3mIfbjdEpRYJfIzP3s5skP7SmmVqGcxD2sMmx/OPp+7sIZ+mUWf3jNkIg2WN0K
CxqPHGFNJxeU3loax481RGElI1apJXgNyA0fNFA7wPjkYKyFGMqYoE1o+RmXhj9e
Sptb2fYZ8Bla9SXxjLQJJFpvwGZ0f5tLTvrWKY6bLain03LZMRMFqi/PqRgx05HD
KMu2tl6k1sTCma6o/vCvx5RNKwhIuQio5nIZnslhhNfQoM6hUhUOc2JRq1rwrfCC
yJZdDzNTIC6BR5QDv5BLQ+LZBKzt+8p1hx4dKhoLD8WGuKeb1UvYo0PqFa4s9s1n
+7cCorIL76bYve/QB79/WImDWCfHm+zPP1YW9SJ5he5p6OflpRjEegIyRHWrb4Tq
mjVhbsPjzNToyi+R41mrS/WV+A6nNEx/PoNrwTAJq7SUfIUuSAfEy7edWsc+TMHy
+BPpMZ2rjhsBouscWgcpx6RyUvgvz9ytyrta8+q/IwtoV44x5rkd3yg7nl3Nq3r/
Wr+j1njEKXsodiVLJEBZXbrv6GB46NWpxkfGP/OgbL7lO5BngksvIgNa+1iFxi7C
zCdkKBAP2ZmgQchA2My5Oasaa+1CDAwTxprWhD3rglut5Gby5BiWSNNoyY0Ij0YQ
5JKtG19WxnoWG2zRx8klUldP8dv11TVFXcDBEZ3GJDTnHgY8dxKLgVUnI1SClCr1
uHiAI1Pv4PIeDMTkiScKnlwG2dkcFV8M2kljFTmClRMDHvSrwNqTVrCiI07w8BZ4
MoE7A3wzkZIlgP3IIqMrcxy5tab6VnDGZK1aonakWl9r4GJxpCHGXWqPOtK7irup
8D75Yg58y250jZkz3rhRHJzN+wdxroJDXjMZkgmQhSMRj/TuyQSyJa4ihEL5aNIR
WFIrx45uFqsSTmspNgVxdWwcuK9PT3DkvgOxdG36C2hM5mVwS8+HjjCFnQTzdW3t
0OwS4i/Pl6Dm8xXPVIWYii1kPdqn9VY8wDZcGqHBmFPPo+98JBH8D/5Wi7uL2017
Qu4y4YUZj2v9Ej9w+hBeeFvcvl6Lgb4fDFLrWstzsPr+ym3hKqbAO3vxSlYFbHM3
Jw1rzsx7SnO71hyI16WWsTmzTbk3c/J4VY/EneZd67X8AR98nVEQeYUV4VmOA+wB
80czPknBlKNG4iuRU9InaXsuZQr53xjpkiFZpjmwo4UNhvmN88IMcWNXO+QkVSMY
M+dG++/TYWlXHqSsuRmBLGgrVHI+dgod6JRBU520zsr/4UOqRXP59WDn7nUUzcxZ
nKwOxrxLKNmxvlNjLtzmro8IRhdLzADj4n5ZtotceFUqVaBpfnhhHsofOmTkP7ox
+ybvfJbG/1J+DC3gt7npHgKxHw+icLT8a5YpbLUj53Kj4+hPZOHsOE/H5wADEb6K
4lms8CthpizsKwj2kTsnVr//BRinbH2W2M6BsTpRRLJqtv8ohxyTkbUbBh8i34c0
gWqAO9FKoK5yLepImvwPKlyhZmbLW78r/uKpg0W8VVtJwMCy/EqNpGGzWX8EBjLE
AxDAEsBZuYKWY8pnlHJ4zbSoNLF8e0TWDrGRbsJzhLHkTAnoJueC5GC4HPNvzEp3
ZVsETicBE3FlmmrOK83FK/bThMoST0duyOofGB6C0UEKDPeX8h2WTtF2nqyMmibq
Z6SS/Z/dY4D9OIiOz2C2jlc48T6vHfBmC3NVfUYPW7kNPPLF046+RS4VnSksvvfE
fsVIzFKwmRGaxfJ/dYDxf5sRv2SsdQFU7rqf4mYxTJX3pGMaUxG0AcFy7rCouAYJ
Xg3dPJjE6fPiYs6Oge95i2Wq9F7Hw1Zi4JrASzbqL5or+YiUgqL7alVCp6dJLDrO
J6zqWGr0sUtirfL4VBeXzvq0jRiNV4xzt1qqedF3CFox+nskQBY6hEhvZCaU8Vi7
eIQ0h2vDtCGgDNSwX74wmDYCueW1f/rcoIU8A/8CIFS2QQZeLMaJ/qkB9Rd2x+Gx
SU5meS1osVnYuNWJ4q8vY37syzbjulGY2iUlN+RYQF/B+TMuTsjxuAM/3q8r5cpD
0dMvAjdxWL3lCONgUkjdWqb9fbcFqd4tMvtnUV28wfoC6nXWNaoxOIBv3hskK8QM
nbCkgcUygwQnhqE3puRi6QsaYmFo4+OnUEgxeMkRviVHu71oeX9mk1hT4iUVXg3k
a7v6vf2aL5sCoAjWE9CLJYNgE2xuD1GNXyStkSbmtYHhIu8VzTdoFllW8upmlsSN
4N5uOwpfc1EzDs5t44I97p+juQHSSG3mJN2jWGx507bIe0U2U416klXUSsER1duT
MWCFi5BAG+B4DtowITfW6+2E6/tkK/wjsytl8hKYyZzL9iOFdGOe4b0BFv6rCVLp
azgCF5JhzQ7wXApfxZde47Gokj5EIe+69HjDF0qP2a2aGWqUrOX/dJ+t2GSOkOwK
+aLj19yHjiDmViMq321yEjuIdXKIRyN/yssilMFIAPS5n6+o3bP6N+nVFVoWBp2P
kT4U4BoriDmWg2DEo/xxUHMtHWt5deydplbe70mqlb2W3UN3YKKHhldYGcbbuSqH
Uu/m8bHOCN16qugGpytMjdoZarQuySD4idY7lWe8LxXQWB3+EsFFzv1UjMiJJki3
2z0nt4e2VKiSfH0nSf2fp7LrExaeOaXPV2hoGlgT5rkZLRNG5pJORBHPLFBeYfMk
y3Nd4nx/HRVbHIfA4EMesrqVW+pTX6mv07Dtydx+13GZfiETMzQ2scH4eszL4IML
Wy1E584O/CGOIjtToeqhO3TMrInTqHwIorOoaHSDibkKDxMvatn+l2NV9Cka8VZB
OefenfGL+qc4GjfurEkbbuIPNGlKYB1QEE86Ufx2LFG/EO5BYSMMrSvA4SRyH7eU
Cj56lJX8EJ4ROGpW+SeQ/44E5y+ldl7ZhO9ESBrnkSvWxQp8MIkd/W2CMCujXg5E
ghFI13wnlSDtq4zZr/4NPusdUhmRyAOViW+Z3WUGExWzAgN1HUTl4TlZoiNgYyfu
56Mt7g7VKu+uoKL3hu8UTPQxfX0aj332fxD7ME3JpvtxgKIkpNcGNnJSWaaJm33G
1psCRsjMoAFaHPowkloLQDH/rA2WkoEOO0P4CcRDuZ+4bviY/eqCsSrCKTj5MdLy
DSB+qDMAn9cy4bHyvIFnSmvaDo7SEboLnDKr2XBKFjtgilEZrru8/EKt/B++PnTI
qQ0Fk7RRsUw412UC/iG5b8T9TiPEQPdLLKWlGGlJWkrEFxIKVo8NtZZrRXD2KnwV
avuSknCMoT/gGQNgquwfUCekk34LbfIkWYhhnyKwr2tVVtp3Pzb3CYkm/QnYMR2J
bMPLiW0bjtIAr7PPMe2WnwpqH/G4JgOxt3YzSkn3p3bxYhi5mN//0mNKr6I1qOOm
JIKMOuFkPwSlqgPsEvAUcx1n8zLn4DiVshmi8FBQHafa42HaLxlpemsGeBPunm6r
aTseD+eQgCrUsyFJjbvesiKva/G9a07BU/pyKDgYcgrcOP3VqgUKpSmFWWwVXRQ7
Ktiaedkjl6ip8F2aE/OT94RgSWUd8Em9iEyFGif0vim87CcnqePtK+DP76xHCxVB
ftHpcCoV/peXqkK+Q8o99kelw0VqKeUN09aOd7L5vuYspbrVRYyFq02oYOTvu6IC
Es27S/2LQrX6XwwKZRTt7b9gOTUItK9dQb6ufIa1Xz+Jyqg+5UDeUmo+DLNxwU2H
AQuVyq04yKp6CXBU08wqbcC1Sra+j71vBKhTl5W5ESOSsjf2xYRFRV7Dni9nltIA
jUzoDswU2iq3WsPFeNhXtpe8OktLmGq66v892jySTOxkd3kV0WGJEFKPAiOSsbI1
zW+hLvMeKeg5CG+Tz5PZS4QxX+j4dMFEx/TTMeRQW1TTdTEkk7JBxyYC2Src9HCb
U4NoV8QOdIdWvGa2+i7ULYxRxFczfrs2BfkDI2Bur37dpVbb43f9cbeAHxPl/qnB
T1BALQqfd3uXvZ9lg0Ufcp8TpFIMItPb1oDFvIVv1ByRbgZZi12eBNCg0aYwJCtN
DDmgH6cwNaJfWyZ0jfHCC3jvzhAaBv6aWQQ4KzwgHI0J9YXo46/EddIYjWzXHgAk
lcTKbqP/OW1jus41wT40EdJsUQVeFjbC7d9nNx5EKqjs3DMQDGcfLDOMewm0+wNk
1Bs6J9Sh/9r9M94QaI+jbQKq4e/4fRBhgLPhrx8R8j/JcixlXXTWawHctRju/pyk
6oRG0wLTT4os41MwikjURYTDvltVe5OZkJHCtwoLNxr4P3bJ7sfkUhaZUbvwDY6d
033PZtjEi5clnKH1kOkPnIkTHe/NNWqlvVwmc/0qLc/484iurHRsFwaZi/5vGkrM
I5l/zvCq5rNNVtob3fVrWqpJg1G3RBj+j8UzdAg7cYuBAZclz2UaU0ekvZriSm4m
5evArGf4ovNbByYymYTjlFzCIa5AyawaoHqHggWX7wd+xC/E3E1FydjbqZLW06Yx
59cTf38TA9CPfVWKnZCOrgUvSucbnbCaur9y0lF3BVSFrXsgwt7Rhgni01MUaUHw
oTLm+5XIpr+EooegrQB1hDhiVBI8Ik94T48XKthJwHepTOGHV5iDlmSCAo3ZO91u
kRH0IsLKqfNRuACd4y+DITWcEvHd6O5ang+GBNbCw+NokR9IBvgH8hsxZgcwYp6G
0EVYRbof37DM7gpfKr9DDtkEuCAgQFcu7kmwfFfZN/oUcEWYR9hEc35gwvoM1Mcv
2dyK07lz8yggKhNwJjcT/EZKZ9HoIfgSrdkqz0scRs675ZMddGOqTEyAzq/wLyHb
roEFUZOSnZu34Xs0/pcCAiPeyRD4zOaNwcTqB35yeOaZmeDGOlwj71ZUMTXbXK4A
wKzJWuYoeqJo8QSB/eyndV2i+JkxKqyoiu7RN9CkGRVlNCIc5YSDdFz4EZ4laBIu
0YHCjJMpehH6wqjztdgJsyA8IAW8Axu8kE6mjq8WKDzcWGo1etZZms+SxMUq6bLL
CQyFl3s8DGSoYmxigOiJtpAHJdrBJooQPR6uo9Fhjta9yLHDFHoA83nruH7ITtFc
gi41cLpUXdeZqpOIjj9y5FDX+Q9fvyjxpd4aADvzAIe7Ax0mPlCR++muX8aN9521
QrQtbwPR6iInmW9mrQ0T8eWcxO9afAN1GueEMnKBiOQhRhItXIawgyhpwFLeP38Y
pHrVhUMTheRq0Jn/1COWYcC5VNQ4CKOYB1niSi02+1OoPH9gcAYCxqszmzxGiELq
daDdBMQDR6yv7VS9UO+vXJQtzV5VpnpPRdPbWGYd2dgpCFODR0hq0mKvL6368IAf
Ozyi8QwAhWwSXZKrsxLebwNE8cLfGNPlIlUcr/V/hP/p6/3uSVxOltn79LR2G/vo
q+h4Hg3hCsqx2IXauuoeZX4fynAzWZtF1cgkX54FSGfppFuNXS0X3qFmbMZda92b
8Cz36cwEMcD7yBGNY3X3jQ==
`protect END_PROTECTED
