`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXxuec9EW6uJTGFtO+rSdWGaN5QJc+4lnkQ5oawi62wNgbE7gY8+klPfQn3vXjZC
ldSC5E3TLAtRQy07SdVzUFIiDtZVYBeGW5kMXzRWys/RH5a3olVRFOuf6yIPh0vI
UtGorVRjA4qIzTjRUpDkuEQtA5XTj/VLmg13EUGKcYHPFaIQ0nD135Nc+46LAmH5
fZDJE8djjHruIzn4QnMtVKrThjgnP435EZGhpyvtPeue/ntzTMcVaWEaxJsD/2OL
I1yYyL44k7A1/7xBLt2ocB2uX0uLgxzrFZE5iyUxyp1Yd0PtmFQnmtzDtXiXVZAS
CpdnJo0EUzcWnO6PgHfestumOGcCwoMNxPn8HL9ljDXEruiWGkfvAkNNRY2kRfAj
iDV3f/oTIkbUnZ2PADOW3/1T1zXT6QlHjb1TCY+nxedZswSsQEQ7pcH9ztjZ8JOT
LrAB/NZ+Pyj5X3SY6x+CeYf3KrMQzk3Hctk0G53NrFjUaQzBLSu1q3lv+5CJP9dG
DuwjCZ8uvRkk2Fbg07rahYflPZx8DODH3im13BpDhGjQ7oXw6Vq2Y7Mu+yz5D8Z7
eS+5aLFYjlBuxJ3m99wxrQ2ntsr5HicCZo6XcltmlLxcBycTq/r6SZXMtUrxb1AW
8Z/w+k14AdQNnwqnDo41WcEoJ9NZJsuJqzKeL3ZOhIrh29/CcB1T5AsyhlLS0lon
942/66MXKo+lAzs+beFRsgs9NL1GBXfDbWI9fQUNS3kvEEI3JZabhhBNV2sIOudG
OM+MW/G8PQZwe7UNlrtkTSw00W5lGopBCfAURHot5yQBNQd/HTaByVUxgqBaXnPK
efdoRcgpUunbDF3UUYn5XSbCA/sHJFyxudSr80CSDe+56zRyOV34+FhUe2fFTKaL
IVlvet76g20siECevYfUxeCKGoSQBj6l1GGCN/TWziuhrq54gbKH5BkQoQj3TzRn
BVcIb0UYmV8r/DhkUdRS+zCDpY8gMT/P6C62G/P07cErW2dPEo7Micb+5U/ZTQLK
2Lx7AqEF9uxvJMwWVgm5IsMMFQXUAJ8xmhZInAiVJv6bDJ064f0f3ruuRMs9h8rX
edxoI9kvx5rKFJz05k35uZiawbS97dIkTgFGiECI2ZSmcY3DRLJz9+pA85QIqHKc
PmuCOpH0V6pAUj8snCBEYcpJd/0/77XUG5Co2SpikhMJgf0MWDQpzfj9hkEP31ud
NLV36dmbukH+cUsO9Y92YBUpbualOYh4ADiJNZv1AnzpBULUUBgdXUT1dSVqEg97
WTVClAx81fyJ7gnNfEIgGBBtYdFvJeNiDKJ1tqVvzWtVxiJycWdIYnSOCPb3IumT
qkTSyjaoElA35vMkBfNrHI3nfbKGqdPoItB0yl3fcIIQ4aJ7K4X8LpywFEuNfT6E
HIX2tcZKrwTRN+YZp56isb8KmrLMfLfN6QstX7hBsd9tTLoeOpjOfyOoH/kqf0gl
dT5QqxUT2G61h+MEI6jtxbpowbsoJkvIgNRW3glFcU2CI1ottFaeSk/e46/9BfXr
HteS5+U4VSBeHbAefsuWR8J6BusuqsIG3lRg7RgdKHASaNxcE+Tc1oL/aVQ6ocfD
oV3MI/hPqPyZb5kDmSe2equF24/Q+AqZ89/S44nwTp0o9RfyjyWxw4sH0JF/mFm2
8IUi59pMKFG2TXigtWZJO4NUPFFZ1SeHTFDSlW4m+dewmXhjnfLuYA/zCLQugHFe
u449XVIsS47kMGsT4+/SsiKr5Nd4C2L9BjM2P7ORT27y1+q5PSwG90jIyQUapqDm
mnmts19crlv4mAGj68/JSw3/Gj4npXSoPvNB/KJJ8T6biAqkWoAP0xnAtOCJ0I3q
DeRWvfFMbYUQgXkS0GbsyzmHiDZIdknPRWmB/MXzgXGeryALtI8J7mtCYo7sEyJZ
sMjbaQs8Xd84Voakbd2x/LX/Kzs6m/JM60Rr6IlFT4yTgzRyOd16Bi5xRDL5ddQG
NKCd39sAgJiu3LgO/OyuYtawGyQOxXWdYKR11ARxewfJ8+QONfKmc0R3kJRLvkRD
jyndK2OmoaF30fF8NCRtz82+8R7800j1Ow15ziaiUWWK5OGSw9Hu7WJwblMdN8sZ
tBpHW2+UqMOYiSXFn30O1kJ6ZQofI3S+wqrKrzf47ptCvh4QD26bSQ4Ki+gxJ2vC
f3QiD8jaeMu7wgpVuUFc+oL80n5oOhm804b5z8PivgsG/OBHI/qrCi1C78e3FYZL
HoOIYW13gpM31WoEpRIKLuxznJoP0+Y79ngLalDp1zRXGnimmNbX5rLuP8HqiXMp
XNjFYLRiFUNwGUyQTCrAMQCmmU4G2KAAkXozCzzE/9t1pO4F5cVyla2AB8jHNnCm
2UnqQW4eLQnAte6ZrVSrPz6Sv+eNcrboDYyJ2xKrtUuxiBUArnRH9/E2SdjXpBsv
m8pnvxfes3D5ShnKf2o3hZFnq0gUGke6gZhDnG7TCUBoXyHrlC9BFV7g8OCpsUZ8
WNFM/LE1BOb2AIGHzxIlaRqqSTrx45B1V7RZZoTwhP/aZcasMDjwTtJl54GJtb5m
nNlE2e9F6JG7Cv6ZviZ2IJw4cjpPbdIu9wmsPgXnjUpZCET72JKHIejyoZZvJ6mz
F5lUVVAdUP5rV51hCC1OWj0Pn+x7sT9snFPODp0uRVMoZjfsn3mjEpWolA8Hlq40
ZXhzTsYEUR1V+XXRs17py69HxogGeh5jipiWzzVgr5qEEhbUDepOMqCMZsp04Fjo
HmH6B5/Ai7zIldmrN79JoGgd0j66IMKnZv9o/ZtkiGWV+g00OSXbwll5GEmAyeth
lWiPhxcADwmfxvXMGlBdnqsAXQXbCbgbY8NLIkzaIhpzi+jaFtkWx7D/UaUfC4+n
G1cRRYKSgZkCsn10ZDl97/lbTbgDIuRjM5y05Tzl2lZlGPpwaBrG3SFN1kp4/nR+
A73GWCfH/2WcjidZKtwk177k5L2s2D8yiB664RQMdLFd6aSd2Zlez+HGIA7mSPpA
QtQrenvdFDkbQJAPV8ZXeQ2Lm5uIRO4/RYlhJLry5m1cQtmwEZ/c6T83Ndqbhb4u
dtgKuDWw9F3jwxdM6fUyFSExvBQ4Qz07c9H/jsCtwmTyO9z+0aGdAoeaHzWERTqn
qhC/vYOdIUq/MzBdZHfPLjkStvL8GYU7cMjUmNyzd51C3DtyLOtQi9CsoJdZPKBp
SdEr9jbu6LbbBup/DfWouUjkkD1GOuJ9KmWYLsSg32OUtJwdIDFM/vZ3cjJmOtKe
nF29wknvAm4uuGGC9aAZKMiNDwoPiwiI7B6kzsKhoB6Kn7lIjpv56khJ3EFX1FO8
Z0ia5XINf0GUgvl0ioaalpnRGphGy3AKbq5AI6lsr1NpvqY97vh6Z3NECg0r8IJL
4Ak95XMyQI9LDvn5B1pQqyQcgcnRfKF2VOQ99pKrf+GNRTYVHPSrOGU9mMTFz/xj
4+g8lzUoDk8cQNDcCkC21MDp8TU1U4n+xAvZj6tZVv7qwJ1b6hZj9PWGszvZy/te
OTc5JJzO5QoyIdDQGkUJFXNlYQwkZIYbOmuqX2FsB1vAUJw2NfgfZDcwSkmI+Z4B
NmcU+fqV6nRync57s6Gw5Zb2scVaB47YZ3KDDQ5U2UeEIm2O3y7SHj73sw9Wu8TQ
YQu8/XvDVL9ko86+1/ZZ8sTPJbvYJ5NQEukoDr/vFEXn5JZ64iulM0YUz1ePq39r
pz4sS18UxVfdgD/XZ+2ptqMoHpduTC0oZY9bSQlS0cjNJ+8HRI4QVu5RuQMwxryy
ZMnAzwYL8kdriyl7AT9oyMyJbrApis2GiLs/LCD20Sf41DcOBr6bQfG6E0mtEzpz
9HMIS8xFqbvnaoRaNmRuajcHa0ayTKk2azoYyIQzTgphnDfNHykfZgVzLK/oTUfo
BkNOBWy8NUnHpuq8yIZ6rOTC3gqIOtuyEMdLSHdjfCgqIE2o1zQZYZbc5ETUuFLB
W8dZqQIN0Bq2Ob1bG50AXrMeqcnJ5eeO76ke9iaXCicMHnmDGDwo6YPvwogZfvMp
Et2ouo3kYwEsPljHQl7hikNRtlYMo+nz/vA6TwnnShLoU260rTXfENMY255TuXHX
PLfiwaV81Ms13UU93EEicmWuxAaCkeVdtnTrd8tjOHQsKvCNzhUZPbV/xkDHxBiE
Iblc5H/dYVO5D0ha3dAJwQMUdnELQ8Aturh1vIVmx0Xi8HrHguME0JLFDpPAJctC
12EXE0VT4DB9eDxcEPnt4Bjv31RkZzQL51O912hqAgd1XpyfYpRJf5xDQ49yb2ho
6TAB+/PGwnMmOwLAlhipdk1UmeGhuro1XEWbIKd8yAKRvbru7wM2tsVitgxuOm7Y
uikU7C0yGn9wtXV6SmkgEhvOcTmBxZup09aS7EnAgLEHjfDemb0sxs3BJQiFOtGY
2NNfc1lVnopHrWxm+9PV1rxrUsEgxe+5/SnplpSLGgLijE4ha9fxoLCL15/96/7a
tYroubnDp2+0GhDEWbwc23XSXVJDNigwfyK0ZufzKPKeTjhbeHGsqjrgQe+4aebd
a8NI61x+TYvLpwrAXgQcYg==
`protect END_PROTECTED
