`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1uWUqnO27qfEoGeB5TJvTAQ88Cwhz7aHQt6vV5OEzIse30MCSHoYGD9gEQV2nvQ
vOqUbehN0axGROxFJzp2UEf78PmM4dAi/rx5G2iAddKfXg+erhWAB1Lu0xacpx5q
5DusXuhbTRD1oWZ0GrpfQm9ZcDEju1+WBNWbSM5qUvsAA5IkcI+dIzTmh1oCpkKZ
261+HLVoBaKWk4i4CSzDiYGqG7d+NGrK+TWORXnnjGKfcx5TrJZ+Ju60LvRdqGRS
+rzSNdhb9pwPmLjfbGDvqzFksLf7hPpxvv8VL2N3b+yzKxG9Tq1lGlipI1hhMTQf
gCHJzHt/1TN+d6ZMcq2s7Jk3afcR2xyTRvKUuV9UTEQYOpXz/NedkOKVehYLZqD+
x0vFW6DALQKWDL3wSs06U6PGvdWlUojWCNjUFucek0FATku5Id9zgBCWSzaOIpQC
GZMLY4Vf0UiOBlkVGutJ8ky4JxDx79xDgFsw06PqtmxSNVbPEJdzIYWKb4Y5oJhu
O8cZN7ll1NPbS8Odi8+4zdwC+z6LT8F4r3L5aGHN64sLKKbuFsCB7iNQZxaI0XdI
Q0sPKhXrUuo2eNgncK3Xjj1HnWjaeONMncvifWgRb2sh4p7qQeSS8shwPUu5WMgq
CcV3G6YAQ7vRChA+0bNFVtwDv7NJn6YNHh8hj7bLQM8BbZ9bHFog7KHnEwTImEdi
uD7bBhnsqSRAwfvamAHEMB4xArWawTAoZHuFBNjTFuw=
`protect END_PROTECTED
