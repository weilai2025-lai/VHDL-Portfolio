`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klCt6EWuFZG1UnHJV/VeqevrcWy1TroJbb9krFzCIq7TgWlYZR0YzyrG3mQ6N3jz
b3x1rEWqV8Dc1momgOlnqu1P8xjxmLKIELpPJu91WCsNfomoMIGikO5A5I25iK1W
6aht5/IPShqya01KEf7VguesB3dnWjI2Z79El1zkvPBirXEdd5GBxI8pYIopLkvi
g7Dt3Vj/j1MNB4hKc2OGn3Eyaz8XpCe7PLbuxeS7UKeFsrcwxUgxgkokjWjvG+pd
iI7D7GAd7Ds3rZAwsknQh9sq+ujfG4Xd9uJ/gczxBHX6FrcgYAVW44z38PvUiu+6
ld8TjghTftm0mDhsi7QGS+vUhIzpu44wPfgJ6b/XATKynNn4xK5qxFfjjEhFQ9TJ
MXi9+j9VGRaWvwt2elQ3NlvdxPTzz2jRgHKxz7yCnM9KyMZgYmuXpbQ+ed26CJ7o
l4UWL9NN607KYMMxJvyLiEr4hHWNY5m4x44L20bjMXZqqa+TVY+Q6Q+Fr/WYENeO
0GymxAjMgcf1XsjzxWXZsToLiPc44eYj63Wt394RO158pcNxaeotmJY3eH9D2llV
drqcol8YS50VsPY+zYPJ9tCKXyvtYTJzGZwaWqUXy39YodbF7DSeHQoOWuqAssro
sefMc8FL7scohPAIlyfJhzoOEZn4P3UNQwPltXLNirToMeDjAVds4XDmO5B3n5nw
pK/dRCEaAlahilxz2i1AiPjjODgIAtTBHKRNphbZW9whNP6UTjN7LK8M7keCC96j
awSSbz663ipMSsO99tqFS+4l7UE5NvQEwrujuXsgL4/V6bTlX0KpMVoHcdtNl2RT
fv6HcBfNHP7j56pN7flZttb6NbTAs6bBBIDVvL+658k=
`protect END_PROTECTED
