`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HIg4+FjlKzrc+KroGZ8v5tSywX09bslTfu/kt9203jdKSjV1siv1Jz05vYmmmV8
m6fjkqqw2qLcx+iRlijjwOfN4ykc2OKQwCoFlaEUYGdS/95a+Cd9zbd49HlhtNRZ
GKNfd78bMM2hksRMi0bl5GhoK2AU2IwxNXxfPo08/em+F8UetrAk7qQKedRlFJWn
guOsYdl9ZgGzgOH9Xh8A1d7sCn/26alIES6UigAYCKztyhrjdwu8uSI26M5xBcZ/
+46I7vHMV5y+xoddQxjPCdAWDn5JHhFrCSolTZgh97OMKS6Wvb3L95FEfD8GdCXX
bOcsrHcEhFHVh7VMYM9jlEHtlQTuKvXfd87Dtf6rLdESirIYNIIo2IVepOjyDr7J
pcq1t602ei80WaWM11nA2ZJrbnHGX1qHH15qTZQbw89cz/ScL49Uj/+gxsOGRY9u
NoqkwmR1KepA2tiRosnxVFJQpnNWqJCJnM0dplDSANhpycCVffR4fBM6o80+yqWd
/3d3nHdSfpVa1rQLXomGB67sYCJDjQ6Dqwcq4cZy5lCsn+InBl7/VcX1MwcRVPB4
AWyfODZno0Nu1Py+kcxWcilM7vOjkfk2dWS5UOz7tgdMLvxlh2FDPirqr1jqy5MO
xwAx9HOVwkvuUVbDh9rtIZX52WvymSrrt3s27+rNlaxWHaQwc+VBsHqePkcGvY0D
HkfR2wy1I0hAbFcf+OLuAI7XGhlElRJXu2Yn5N8/yyLkJP2j8TQnbO9IMvScSQP2
rSDuRUBaQFiBsZ2jgLa3xibjBJmHlGizTOzBhHxp+VKUG/3vJrIlGARhNLKRLs8G
mT+gG+dUtJzn1N9/HXmeX3XC+BYwIUqZHedj4ywSAWWWzoK7p/8FDiMetYGO92sx
L8be0ER7RPYEnsRLo39iHHZGKysDoRREfapNXLbwu8SnWl/aMRIRoK/eiAUw7eq7
HpoUEk06w/f7VfNRtthuIDa+2E5LPiG5arV6cLcCajkPhEpIhnbCw9nXJFmg29sx
/fMQMikPo6D0/pmjtxKhSzzgkNNrmojsyPg8m7yMDZVq2zCphWZQd0vJcFAtX8xB
sLsYOIC3qugA7ZlxwxIeoXumrrgMVF7AqrOVw8rSStmcWfDM3kx5DvCzV5r5uY1e
p6LDziiImG9GE4gk9VTuwpdb1VFN0IFjIOU2KHpQdcMN5EeV6PEskg70X6gythBT
GxqUeTS6a20H/YRYaZQks3h+GX4MH1wW7eWH0f/CCvWuaKstuHz2qVrwy3h5XhKX
Pmb+bGjo5ilXIvZH51s0J2MrN0+2F5oXr7MX9JQDLU7fABKFz5NWA8CGX+iD0aS4
A3dvqQim8apYt5iSfNTwULV8FnEqRvGfrKt4IywqA25Ksl0keklpam6g+LfLYR/u
PW3TUhmqP3X43qVWjtJk/DtXC/PBUJP1JEu8UK1nc+cXFXvcmkiu6P2Rsxs5srEE
TTxfAhFmYtZcIwQC1SGfkVaSzGvVoVCUrJdyDpOCRluhgR1EGFP2gDQk6D/WSLVj
Ve462M2vvE6zb/EGPC5Y14IO0/cwxAZdPJ2ln0Idq16P+9M4Refs+CfKWQkZdedK
MhNEJjf9/AFacAp6BCmyOwh/hPHBsY33PzvukzFOCzT6vqTziFqdYizs2HMe2xcr
RY3v0CX7xpJ9znZgTzhRd8XO6L4JigtOr3iUMLuh96u5nSXzpYP7xJyMWScdclMY
BXoV6wV5FBwkDgsiTG0ej7Q4dLTG/F2lsbZBb2HRMwbv8xujmpjSRCZHYb6QySNy
RA/6yZ7+Rznw7lOVmFWGQvZJqzUaMd5DCrP1LwFP+T6pl9IEtH3fMWVyobR3lsCy
MfA+z60nkcNAq0OsltP0D51yQG724DftrnjHcsfBYy9blADe1vdikeLOWS8bNgaZ
jS2nv/1g9kjRNxWpEpA7wBcxzS6Ft1pS5hqhjbE+aF4VqaLMyC3tIpdXzXOcSff4
rOsHpzcPpsdV53NQ7WFkxhohwda73G5mr7F/RZ+2rJRBzptalzrmuQ8Uyxka2shw
HFKEW+iN+ytyF0o0l0W32yRq4ZPjARBo9JXkyYCiHkPcZBQSZHaT/2Gs0MNBL0M3
s70BUEvUeXIaI55/0Nfh8oXz/K/1JF7cdHHwf3PaP8CfzE1cYULtcSey7lc32zpQ
P6txsZOQRNtHGtepdOmLuX/AnTm0CV3Xl6lYUB7CpocXlrvQcgCuO+FcxC+0fyer
3nnhogBRM62sTHXFnaY0EdXBTmSIQMi9QyuCdGxdj8Ct0O1/KoqoDIDL6b2r35FD
cfebVa89oaG8vfLp9YZS8JORSmdaMa/Li2NBggnDw77TwXWqSfX2niSHaIanXHnr
YNO3CzS23z9ZuwQ/meUhluYallYiF2WW1WfpQKgX1W+qMoQf4EPCshN18sQjC1Zn
jdftT02OEHsUSsbWJPmjH5y05zC/moRqk84YTzwRsWzr83emLmpFp3cWYOIUhw0i
tB54LLO+3xap2DvTwlJTZPVj7LD1WWtpsIvieXhC0UUZs5xvRiV/P1u7YGpRnr1V
Yk93UfkAkRmRYt9R8UcGG1ijc7UDwhxJ5QtFn/Ydzm9e/pRxtk0SEGdd7Wb2gMmD
Eco5E2AWkWbEGRvznHheSXr0aA/Mmq8XesEZQZM/PM1pFg5qpbRDF2kVEih5X3gk
QhrvlLxKdrS6ECpcga1b5t17MK/LCLJXpd0AEW/baO2Fm7lXg23eMtvoeyStWuLW
VQb3+N+QLR0L3l2gJswpnBS/c4eUmLfn6hfz43nofPvuQsb0eRouKaq4TvoEle6w
fznZdUfAwt0/HDPuIPOXcsyN8SjQ12o9FL1lyo+0Ia7J/Mp3hCtzWthVpseMtepY
EOriNnamrMpqhDgLsztbcsPU7klwJrqJdcSiLF0Ds5jeJ/I4FwXQFtXplsWleHGX
0ia2DteBvG/dfx7+pjqGMeu7lPKw9f4nLb3dmKHU2P0JVX0j4S7RpCXHCgotylWK
bXbeIWaYJ9MEhC3RF7zkhbgDqN/LLIhrkjpclVSYvocrmdFU0pGpM1aHoh6R1cLo
2xIIm9kgcbVVnuPci7tTINr/qOdhiQn2S2Nqg67OChwkzPHoYBFJaTrrVk7ozXel
h+h9Sj9nO0loxbvIP76L5Oa5GkuDEoq7JhSpWAcO7646slK0Y1JU2GyNz5HL9Lzi
wZRNC1l1VwwslTZmszuU4QzmNwwAQBBUZIegJlk7UqEdumX4vWOR+L6Yb84dziM9
slUvRtIQNie9ieA0DpeqVDkvxMvb6TLjDJ6s1+KNHt8FO5BiHyZHEQQBL2dKQdAC
mpk71AGLm4PCZyTlYUpb+UJNNFm5dqdtLPxTfkq7Jbiw6XaItlntzsACIrM5i78y
hajA8g1t7pk3nFl9lRYnv7r5Lpf/atIyh4LvNszg0cXukgw8NBV6409Zqa4ABDc2
cJ1llIvcM398YXZHvfuCSfZtBQ8+MFkv4r21w1hWTeiMp1iOdi/lHfMtvZHbhyzd
C25gQm+rt+M0RCYYa1mk2NtbHYZ5dj8M7TME89FiwEuz7KQWkAAoK0z0yeevd0q7
v2lvnFCSa86L46n5iu0Om7C9CN88rTFKwEEYLha6xv2qrznmijkblwjvy6k0pA7J
tJ/Hgqk3LkbpR+7TBLytvjik2ckrAOVwI1kntyC8SoHxpFt+KwbecGOYDizlesyp
qe2cBvSgnK7F6ANXwBp9Ohd7t+37p6/hrFUM1BQve7F61wynAYmYj/P+hj20LKcc
ojFhOjh+QkmNbjhqMV3aC4rGkKytox/lldxX0CgWELO+2iAQo97KgN0JXkqtkZg3
To7bTUPQZeKLOTyUkNfyzN05+EQC1d8KiacewRs0RmRbojLjVjmbXLk+6NBoJxrj
XIbn/RFEHBJkZhOaZfcGtgqtW7hfVLHbIMGClIe+AdlG+YzcxrpsdEYZRsopQ3Js
+gkfTY9sO6ZvOmoMRZmQjT+Pu6mv5XWlezdgJIkXRZ065ymBbmDfKQFao6f7F3ou
1nLXNgmf9nd1x2auZtT2RNCnOhRUXSJOoMkM9J3p4o+QjZPGJuQoJiUOQZuJGmyV
WSBlvt5ZzBCH36vDo1EfUcR1CS/JKJUv/KCG+3bH6AyrHO5VJkr3y5nFzwOYv7yK
1obCccmiNGgxDMQJC+bbKEIgRzUL7C6plk+oM2EaTRFpbWG7BDlTMMBlxBdGKhUy
hKI7sXT5T0NwbtOrtMPah9vlOKLoPpQDpb2HZur99g733hg5h0TrXRV100HwqUGv
kl4CsdmpakK3webUxpliRUWSF9xqJePdm7SMFK924nY3ur1mFMPqQk9uNR2/gkrI
ujcTi++2hqLdo4VN7/mA8CS4tngN7NlqJEJZXY/ngSq43Wv1DYrrq8zB9HcLlu6u
gZ0dbUkyA/6PcpzqWUhBb+0hOC5PJQkd+Nrw03fh2cH69LQY9BQ4BgzZrEZneaEb
8Y/HKuTAwuRASXGluZ5qBtCQNrDW9ZpIX/aiqHgkT0q0dmUffxUuWtd4tivepKSI
97+YhfmMA/l2+vNB1YyFDx6kjw/Ulro1XBNzB561orAXkvlqo8NDH7+Ti+FMxhCt
BgJyvdJL/KKFZfleUsjJnr1Siqd74FMCp+LO0VakmJbc+kgBl9+Smn4p8h/HCeIv
F1sbu6HhO2k+hlZELthJQYFU+amib90D5wvT/ZO/rxOz/pP0CSg3CPAt4dMwMDR/
EDymN03FuaNZbiiFDgILSTTWrwI1eMQAeb7/Hgu/UyIsnrEA4DM7qqjUNa4H2ZVm
nxbsJ6LlojKrNGZ42U49j7TZ8wYBkBVBm6K6WukOEVM+OPz3TW9xYhOZQeVNGlu0
gxBpfQLzxCzt7NbClKhmDH5uCot/wVQy8aVcqwxBYhd9MJm4pxsZR4UxCIDppbr4
v9QJh2oT1o+lRnnEwg3sfEtx4qeX0TKP0rdj21FyBctlzMyd2aC+GMiLJBHf3pZL
/mYXxlyE9A5YfVkSxIJrI8CJTPGoN2VHapE+00V2oWZQbHWNy3Pjbu7d0zyJY5bq
YhadUpkJrtU4NR1GtMpXco1k1p7+i4q3LiT2XkKr4DcqYizIdDUeSt33SK/f+ZuW
WLvVXuVHvM0d/aDal5hjo3d7qhWjRCRVjYRVpObCrXYns4e2yZC/EwpMM0WirDp+
5iTIajUpp5skeJeozaiLr9LPvfHye8aK1gpvH/VY3aXazkz8kHF6/wKcrr3doC5l
kiWIEBvkqV9PfY5b/BjnASXbPrLOxMxIi4t6krUgvhthqLEfgvuGPTqGQ4XysITe
/pB/QGTMuMFjZzFt5OWfzz6cspnktOMoXxKAMUIHNgFZLMNT2tAzXJitWpnR+VKB
d8naik+E6BZD8GbyK6vxahVH2845FWhSrCSHiYySOEGg9mC/YLmj2ZJ7WJGgyGHP
O6Dx2eZa7hgzyUM9o5a1dVUUiwtPptrCQTzXeBqw7dlqFSGMBtfjbP5tABH1NJJt
xiFNH1zbQ+pE5dQuIosCq9ooPosJ9q9nbBWIXhZ2SUg/hJRwCwU8zT1bIPj7EEf9
wcmYchmkWnbwsRuA5tXnyeoR1uMFEv9ZFjV5U5csm6GcMln2ZoD8FxiOV0rW+I5P
LMu0MTrEQJ7jX4pmbKXHuyXEdijLHS9gQTIzWmM/1yGlMAvDSYT5x+BZMUPkIiTR
Su+iRy5nnxioPRxaA7RRNPoIyB7t/hDCSR6QUzWU6ltxyyjTYy2sS4a0rw9AOJR1
CTdDFynqHn7JHunpmGodJwHl2EK7cFy0UsAHkDSRb++5/QtaXWZOmZaMkp1gFj5F
QAzCjIxAIA1WAGVbp7sGGS+XN8GelBxHbzkkdQWpwWPb9t70lJLIPAKfUzgKaMjo
6soUeBFc3FqVapzkWNt3XtPwanqn0gydWG6OyHfK7dz2+uQ0cyhOAEZ3EV2Op0c7
rBmRiwDhWKtJTDesKld1SQOVk4jEUvQRszXP0A68adkWBfMkdzyLpgaKXVquomk4
Y155CX6ZrHI+PzJSaOLwZPnWR4uxwqZi8NZWfyzg5uXbcrZGkOV7l2ThCKs1r9X8
UB0exmMJjpDUmmerXvSWgsD2Uo2KJmY+TLC7Zzr8NmtHjj1ca1h/ien5EomTEnbI
ahe0MwCbQ3zrpBSkTFMddZg6k3JCE20MUy1CWY0DGqTNHue6wVUiguUTrRCh+b2S
CmsdYj9CnRgH7vx0J0JPXea+KqzblO442N9oJc1pLc+GN1WMTKUt076Yp3p7hu/F
bkUrbIPOjqfNBkNrIB9ZHu8rHD+2sRpNlkHA7OIH6d4ZNc7DBsOCzVHdUNRXBIzj
HlLJuc66z7XadMh6Ej1pXCDRX1xMyisTZ98eYIOgQ54o+ECFtyZVMx+TWsjfDOop
VJhs6mkn/5ewOA9S2208DyUOAtxzoX23V8TDqoeNv2O8d/S+WHvuYsL1bzm72trL
Ey7qHQo3r1FZSEYjWKj6lIhkB7pC9X2Fw4zayP1YSYqT2+1Z7X3R/JfTVYDZQjuf
rKs+hYQYHn3sBCMLKOYzY5om1z4/IFUpmBFDEUp11S7EIFSRixsW/dpcKwgGzfnt
AFZ812l9DieKhsDF+vhsIr0QDC8aGoaDh0dqF2oD7HIf5LuX2R7va7bNLVNVV1A7
3qEcrv92Dys87MOzgDYmwY/vCe3THZ4DruKrkrNzLQSIqE3/DbQ/prLfCLwoFpSa
lyfo3trH0srBFNYoe+f3reXvvjd1OWPWL/nwMVrDzKpdVgtSolo8YEcCUTGE+NAd
hFDQJH6X8TZpRQYWLg2FtEdPHdU39awQQvD2AkhDzBp8RNbiG/MP6N9Huq6BIGef
chUN7HXcQm7jFPoYvK/+kKnoK8UXA08oWcEOkLNvlNkU0uBeMv9hR3BlV0Oz2TXA
J0B8uJ2O1KjOahecbFBL785Yk6WhZwJZY5dcNT5IMTo2lljBzAm2zun1nZQzv8ye
+b40504jDJBhcPGSqHic+di95q/+KHg8tciLZRNTgDB/e8xYsP/KtCX9dP7VcSyo
1EW7X+Y9ps7wRtoQGlKvtymAdYIXZZhKrLITPPb2E34JZjjorKHiSUVrA3d6ujUR
WIhWdgisiDtILkg+R7rXKSu/kiyZJZxTrswb6/QhRygKXJrIlgXo36A6YUQ1RJI+
EckyYPwz94KkPLd3iWzd88OlAsbE04SM/PHpRhtSlhuGg0+RGNEPmUmmEu8Qsoit
9Mh+iUMitER9u9kit/TrtqXeMRJ+6aPS23mIwA5+Pi8wQ42Z7kptNRtwSlhlyLN7
eAXsVSTpb8E8mgRO+lJJkiHt3QWSv7PbjYjeSbZwTcZFIxkDljWUDhybo3F+RmF9
amiAQKrc0WvdsxpzbqKyNUixmNs21PgoXfW+nz/oP4EHcym9AIEzvNvY+7Opxp5X
ZGhyRKPOd/OSNUAci8X2uUkZfcwkczBhalRfPyKw5BV5aAnXOmI09ioXFL+2rPo2
G998sozhF9x0eYPkDjRJf0H4SWMB0RGgUXmZ+jUrQpP+zBckkqFul1sl6P4O+YOR
nTTYperCI9gSd41xmuL45y++mYCh9GdSc9cfNrE1iH+cqtojk18CgKkB/SKiiqJL
bU5lqrbzSZmXrmHv3n1VKRa1LR2DLqAwPEV6SWnspYqaZ2Cfmfmy/twNqQ8Y3i0d
gvVAlPS146X7QWLz1pbBj28pYDY/TCp26WPYKiIyygbjEGrbU3074K/klkA29o1H
AhQj80KUWwkEoeEmANy9Zq4d5JONQPeZi4CyizFFT4Wmx1wzPIVPepBRUzooml8S
LV2s5sxceNPpeQe1UGCf3mpZy6v63DIQRzyinsp9gLG0pXgnT9opHUBAETcfmerY
eWPhmp9F2lI5Ki/J6Wlcc42uh7fznQEPjOsZSnYg6lBlillZeO36DxUF5M7NKMyJ
iLCcxIGcWdJSNEFA9b0Q/hKnDl80SeGIM2bKlV56AyMJCj+S4D2yTcQ2+nJiktSo
bx8NUHQhf+0OcqL7SXb8RFHxituzhm89mXw2p/j7XReA8V94zlhCLl4I6g/gt2Oo
N9TGGdnMT+1thNPyg9R89c1qMSFo0nPBe2mEv4HxXhqGfko4URPEo4qZBL5nLjwF
O0XhRrOUOQko+0zIdehJGBjtGoIgYU1hhysAmvjYj49T+1jF28daVvAdV5C8yaKi
a6dj2wyY+MSg6TN2OIAnXf8ntFXDVcuDXORRCCP9Y4mzvAR8yEeLyquVm2XH3f3b
RUg3iV1BG1yeCEt5E78kBrBgSfFypCU/GmUcaQNRrIzgyibnVWeVo2HzI+U+WxVz
PVOdwDIchmZ9a0wFAp1EnsFjDlIDnaV8Hf7iarXi0LWWiz2m9iuFTeW//gpnE/01
8dh4dF7OJQm6j1ZGyVE///g26joKhhZk31NeFoktuIlWkM7SrF4d5TM1ELplfp/q
6adxMAiHyv2vPTt/IUs7JS91eF3dCOmZlf9dEps5sjcdOPXYy9IPgkWV+t6APG0v
jKHdciLilJmbpsTHFYqVYTteUrHYUqwEhp8ImbGcxh2NDm+BPmVKanL8I8y72tkk
VoeT6A+8f068WweLak6H7urKbYk7tmKzpS6+Nu0N7MxpxGbEAwXiG4OCBSjwVdXp
xHNkWRgOaGw8jIGWSr+S46UY1kGx4HgMrN4/GtcvbKAts+Rrp+huhLcuFwFhZ6XG
gQDsNXaQQ8Lpey1+C3bOy6XH1mM2V4pJR6vNFZn0GHsThgBSyHEYHOicX72F86C6
5qEypNVH76MwHSN0TgQoifFkqWaTxji4947IwdZb+Oj6K/iAKui+XSsgsp4E6LCD
r7OJEdgDjVq/rUloc4wNLXbx1lv994aJBwow6U2p9TlNnb5tC/padydWZO+JQmMt
/YQ8yZUaIzz0MQ7nJzvMYJYyjFFfY9A0RISL+h3BbtJG0qxFmHchHgJbuQ3Ab369
lz1qQqL2CKvTkeclWODf+fTZYf6C6Rn5rlXpKpX2bBYvn7kX4E0eARHrMPm5wbYO
1uHDVphi75o1rBJfTtLMEjbDxPpicGP46mTPBfZ81OF9wjF1Osq/RR7AySu9EloU
g66r8xZtmm4wgu7iwQKZs31/uWYJVWP6DwHnX41VZgJ65aun45pUk/K4UN8AWEfc
sH4Bve9rN5jG1ezGJqk8dZaTBfdTelA0FLY1t/qv3ynGSzU3YeyAuZtfzfI5JG9Y
tfv46+pHBmCWQkPIt0bSj7PBMPI/m3bL44DJ//9d2r/TIdbH8WVQtLorVbK6yFy0
6aJU2jf61Xmaylk7rpuy0x58unPotEg/+XZZFI3LKGqU6b7brdFpEszKwbOrZU3t
gLinRYfdhmO+WNxa+4MdGjJxyTwRfKbwZhIXrwtUR1yAJS1Lsfcv390O5/p6YR5+
iFiFFl3xb3TXnBmEW3Fh3KitrODu+7YDZjxIVmUWCg67raFVFGT0gmKeWqyNW3XC
n3I3t7qAYYOqjZc/Qzj+JmmOUZr1YI4Qml2E3OSbSubX55NFkqqlw6Zk6uKlJLXP
XWbYsdVjofcIX5HLnsOQvNvIW923kuZ2V+S33jPldhChQ9iTkM8n5tDOJ4Ct8wtM
x+wcHF46OjSX7/wJNMKkNjrduN0gvyxXm1uoR+epL3fvvU4UCQNAWNvH/TyrOIGe
AdOTsi8vPG1Y+bx1hSj/fQ8JlU/FTNGG8qZpWsVQLUOQIxOgK479fDGDQ8fp/Qmg
XQqHzMEEAOgIp3KWp4gM8tcsLzoX5ab/8o4VOudsHvKVCOmM9CGsMC87sOiHSFCU
RvdBZVwIBBUm9EG+6pnijGZo8TpBXPy93jhobeN+yQok10q0j88kNTSQYsrnyoUn
lFKZhzIndTvxTdmVXhuXDuEx9PmEYLqmk4s9ESYiXUgkwHIFKTw5V/Lm8yi+GE/x
cnOdKwsO1wu1vdAPp6eqqcnoc+tqCRsVuC5snyHM3aLzPab+jiB3Sgc+tDBlUIk+
Nq3uzdcwIO6sBBi1dmQOx+Q0H5IhmYiEi7FiL8CAT9raXQ+ikBzlYNDtnseSQe5o
q8vSjk2Rle6udy+GZpQk8xc1zjHBDya32V2t5GXH8d1Un5mZQxxyg1mwGeMEYilm
VtbYyEaQ6psGV6+gbLSWKMCHbny/C6fwxzrpAOEl3ncFp1NkQd06l0bXHalZhC+e
ZTx+S0Ekr8Pw6gA+sRlqEtSGv9X6ty3b/vMg/JHsvgYfWicB4cs2aC5w+mV9SAkj
8qeizbj49KbOlfGSHUHbXrbRTUFZtFNP6BwhrPW1zHNHJ9K55dIMsRHlfSFCgY50
ITUEaZ4fegleQesQ9viUl/3mP7O0wG7YHt2tjCeiF4FIHs6zP8gcpgomI8EJlIBw
yESzwzNDQsY5d1YR/+RDA31O3dLdyGNzAaggoIx23JtOTPTE6HMMn+X5GGqLcG8q
aI3ll6RSM8lhUcMa4+DhNtVmwoJpSPuBKiNiQ1ydNxwi51yRwCmS7t/QwmiJeSUT
sA+6CIJqP81kQRU4dqdYqhI5vfoww7487K0/T9y5U6WJYTFcrIM+FAH16qaJ5Kcp
nRxfBtT9vH+9uzKiyMlpmNGegZxMRvhgOvIX/8bL5ULL6QoUwUkMkTpeZWBCNBlh
BHJaIwx9Ao5Ex7mNPwUUwc/PTChtUhVINvf1iBDW2BsYYoo0FG5iF2nf+OHpIOuC
X6ChLGBKb1JsKoOEioWNMwpeY+lf4sQp8T0fXfE5rR4SzP4hHEYyCkojcTbHAiVZ
vndbMu0pIJ9p07/tSN+yiEKdNALX1nCFBN1pqXOepVJVDncXypxDjPH6DxYo96t1
NY4DCFSg4GTFsnQrRSdQBJ92jQNEqFT4pH+4e67H5S1v3ziLGtW/VUSh5pZzXIu5
9OHaxEHGcbJ/OzB7PH7JSgymAGIpkvc+5dN8QJ69YS8xszWuOvpWYgV5WF+jbILn
G3ykQHud38QaWnpAtOqx0ZTjnBLeQbMfyC33tzDkxSuFMqUnAxQ2pTlsszieIw1p
cLxj6P8zdt6FMmwAmysHfqu4KzdGJ9ym8y+3Q0QbAWXI4PMiuPDvFxyTSbc5gzF2
aTM06wZ9PBob1dB4kffK5vwRhEuK9R5eLQKG8pzIqNJAnKcrxXKH59EzDJrIUtuO
q5gO3opq0LyINv+yIsImvDWW7hPQq9KqMUMATFlbCO5HmfvGy9vfwm9MEADWIMnC
PvK9FWc59vvYuR/1IJZUS2Ma4IbIy8DN18mAqEKNi5FcqiT9UfBLAI96hWJiRf6X
dJfZkbpcwIHmbgH06+30BNOlapA1N9S+LXS/b23qxxJwFj8oVsTmtL84Kiqg8lnI
qfympARYPcNabRH8NS9u7IC/2Xrs4PRvI54flbmEym1TjPFjBgXLcEEQp7VXToXe
h/ks6HgI/ucO2OM1wnYErmLd3GCcq/+46e+/eY1x6LRQRddNH+nCm7Ruu2Mo89oo
UnzwLhAZ8VoJ8kyj5IKoRheYeJQbq9XX+YqLeC9VTGbru8C/S13x7JQNr1da3T6x
wTERx42YE9BtiUvZ780erkJgnnu85a4HDZrfKX5tnWNVNeOBr9VoLt9dbXnNin1F
1EixCFvoTauGSB1JDBWi0apcFQ/coFNjV55WcQp5tclWeVILyuTXOKD2ABOQUcvg
EYWUf0Vm1/44F1ZdnGBQ8pktHgE8Fv1Sp1xug7i0FbnkeGeKh5DAGAaEUtsQE1jr
QqOQvfcV7v/CVKv6RocgvIJ8YJPZCOUKW9y+c7Ayb7u5gEz7ZX6dSN7NbFF95JBq
WQth3FHRcFj7o6As/8Enr7CtDZgRZ/PIM9o+D/WEbKnqP/GbftwBZhNigTv8+nKA
9nDxInngLl6C/wLoaQW3GewKVq3LE/ve7eCPr1sfwxvoeWyZdWYyxfPR8YraHpbp
Suczbj8YfA1bgBMuMjT9kfwvCHSBGW8+aGplB0O/4jBF5gyDQYJJGTogG2RlM5UQ
BeMoLAUgnhY4QeY55rJkuPCFrZYuSJ9gxAtw2pscyCd6a6iuR4QjE4SzRhnw8QKA
EIWbNUeA2jyVt9fXjk5peoEPRqrMBPcNqUkfy4Nlbjkpf8YPfYRq9EFrQtqgPwSO
BdWLH7dJp/hqaC8p2LTpIE0biUjl5R92wgeMiY9cPBw4Lflm81ss5fo1Ix2hR1b9
cqzDzfdfVB3drO80HFIVpHa5n1qoOuJo2xo7LCliG9Xe4tqHo+xErngvvbHn5xlV
QuVnDEE7TTu8BtiueUDkslwq3qSDsB0xykCSXrGbX9ZsdYRSKw+iUb2wheCyySYk
uVJ/rEqPk7eqSzWC6kzEmFO9cst9n320122Xnpxgu/JOIonlZomyx6aIG0sg4AUI
r+3RPJMS6RQN8H5Ev4+HpGGxt7dy0MC8hqZI/AJL+rxCzliMR1UZEt7iroz3QND0
V2SOS7pKhEWF0jjZZIsgQpYlPspBPdPKpZsENbnBHgUWn2oPZefNodb2MEt25cL4
90o7iMZAaBaPDwJbL2xUSgAH+EeOQQeKFJTbDtd6dqsxCCagwt2Sy4QUBi2vpgGu
4oSGO1xPLHXYsPlZsXHw44KsJH3M9lMNTtwbIo20VRlTIA+KU7ZSLU3ZS0QJD33w
7rF5BaKHcBm0VQqd2KxtRxp9rq1MHdeMKxkxkxtkXSIcZdS0R6cGgUVE7V0f6coA
PyAaDbSEaPhrLzaYL7VllHH+Ojua+UMNQJQhjlI8dwLg0tYae9DEhZY3LJ0Xaoak
z3FKup1xJpxXmfKzgtLNiLn+ECpnv8mnNL8VuHbJYvllA7sE6b9nmrlzgmBYsGIu
rJ47wNQ5qLBa1kaZwHeZE9a/SRzl1leJTRQoMX3XZoSx1iyFZ0UsrsUZ+P3PaI4B
z2cRhEiFhK6aZQdeM//Aj+JyvHW0ePyRMBzXX59V8qVgT0CMZ1T/kklVSiBBaTuw
DNZSjOxXl9raMm8jk/mRyGeFaOVWTtGZHPfTWa3XoASWz+m224DSvzZ4OhOG3K0m
YGAU02FZcY7s2apx8LCGDvt0P+ifpZG16faYfP1HkofKJp2h1Bcy14UnFcfB94fy
s0I5Fp6p3s5dZgb0tdPbjuPYwD8GLHX+vgodrq+/s5XEGtg2tOOgmagrZQm/Gdwf
kgN3Qx5B7t9ADhO8iGjXT8v0h32JqjOMxul3HuF7eY2QYsq0g1y8UM+s1fw1baQc
1x4NkZt4xT66xmy8CE4p2yjI3NjiyoEviOhEIqiwh9G92ei8XCGl5DKDBLZrMMe3
mhxSsRRQoTHhsHxmZL1gB9zsJYdRJ1tR1VmgGsH/9bU2NhQTYercETy/GgZwCjS9
sndyHHudrI1t29R0Ry3lUJWHAFehiN6KhTbx3TG3vW2VZW0GesDEDtRwLQtlqrxY
cJiHt7TP1d/vjxH7i3EwOgYM3yW1IXu5suNCb0iuC4XFFyeBKCIQoAm3b6Pmoj1f
fZueJQmNJAqiRbp1fMRtqTgrk3Sfniu91AOFqJfwkNJGkAikqlhmha0mEMyL5fXt
wtmZwccVabR8Rjc9un3B6MQVD/JPVtwuUxrrIIQ/PT9J5KlFBKgHxSiyG8R58iQE
8M6maDqpTRfdlA0pez/rJjVjemZI6uaPQHHcIMXpvNd6Wwi8rpsyKw8Dc2es+5CN
rAzUzsxhV+CInpixHl2IgC3azTKm6WwGddJjKC1Ad5+JdbijN0wuLOUBRJCtGrlg
LFuDbWWWjX7H+0zk0ERrKggfAQeBIHwyf3h1XFVheJNJx9CfhZo2b3fr+qy5tXOY
Mfnp54/V6EyI+yVv+ncJRxuSsPyT2TovrDCWzk1geIlchPfuc/2KEDUJl2VnAaHL
33rAubZQIaCLa3c72DBe/5sobGqwgc09rSQiCnFSXfJ33ht6Y1ct3+YOn9DI2rxl
r6PM2riwNuEvit0M1s9zsWOjcCBZeMHVQvXhYMmoudOFHLMvnesOxey1yU7JvUmQ
+QzvZ+Okb1txqgmdvwT96xyW0IohaMkzGicXek1drL3fXCSMCjsV8Jtn4pMxAa4b
xV0AwKXCAbEQDfxGpzPzYbv2cH/NAaJdt0Yg8SPGJaJr/tAW264a64L63dJwQkN9
ECWe30nTOv/LhLDkjtonQyrS55OtowLDDImeOgRNZ7tWf/2vClZoMilzMQeIpQUG
mW8YwEo0N3MDzf+/qoaxwSsHYZllGZtW2SMyN1hqbXa+yTUiKXy8CS9AZ7Zn0tDj
FZ1Ga8PSJqR0J3o4xjk6cK/ho+GJIb/KPsDJs6CUML2QfzBFAgpS+BitmjxLXjFa
SWwglJb9P54WZsEBE/2UoTcOgHq3sd5BPlnYUi674k4TXFBwEecFrogzBuf/JTZW
IniVGOiusRro8omd4Mf5424phVnhpTxeIQnUPluVLZST4Cl+WFgQhtkCBMg4Jfzp
5cvYGorX6wJT99TMXtEaISCxOPPtxQnOokLlzgsfxatXhXC9OYUbuFCCLHFB3K3o
+DGodO0M/LrRcJ0brkYiy1HxIhiCDi+w/S3plTPGmzTC6Lj9e+ZciXwf1oZY7BL7
nwHfYkeyuhbapYD4OFWp38BwnNjpg1j9ZN9YEf/DH/jg9l5ka2sGObr7uqiEaHMz
E/CBr539/J0cfZPIXNMXuF7n/uTsIgiMGYpiq35atQYdVBsqjWXW6NaAUZmRjwi7
u3riRoO700Y9X1aIXuUu/Vaih6Au2EaU6sb0GHHhYOZEytxolaSXVfDf9+k792qX
BmUL98cwBc46jzuR9I2Qwc70fAK26uJVIhLpYSQe+Nw9zPKTThefe3X19bfodCN0
9GlM6IPrFStsQ+uMuFx30K3dmxUATMXOtD7W5bvUlrcYQMO1IQ8/MtRidt6fwkdr
XBsWH2Gt7kUAb/atFF/NgCRBk13o70bDA1HSY5kZLsDDrO0i548TJopFZuV31ixr
GBwTgBX+CTmy+2RyWNXj7BqFKscKJrlvZKUDlIb5I45J/loS1g59MSDiq4DBI6x8
`protect END_PROTECTED
