`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
svu9dabr+VmF2W8l4fk0Bx/psofAbgES+xM2qaItgujjUuWyyr2dIKIonCg1bWvq
jjJ+4bc54dV5IX29GTkNxTUczypVbtbCubZYOXXHkpjiLLRylRJRnTltMX4z3IoX
FLle5u8wDRJBR4NabWYcaaOAmT7Gbh9njr+8hsm03VNQd4CwEY9xb7SipLgIS4Jq
+1/0k55dAueR/oZnxMU5GUO5nicXVzvsR2ivz2n06Oewegb7otQh7rYzGvYLSbLj
qXm1XtWOjcxN4HPXnWLhP/QaweN+VXnKTHOg7RDDIQHEvkOpnlmlgvuc2U4Bm+15
17Ia8CzLgTgbZwmA9o+ubd1YjGJ2xBW4TlDXFlweCCFDtTgBGh6WQTu9UD00vCC3
UFSF/z/wanehEyi1AbnKaqrypJ/1nXCQ/T7Q4fxjc6PBAgVmLxcBGjlMDksmdikE
gpU2YgqJqnFluVCBuVTsgXqVkBvUtZ0eOZQ5OvAmJQm2eJmLgwnis8z0GpVckRRa
oymLvRTtj/BCr9Dvkyz0yIvg7TTpPXiOlOeYrcjdEQVWYwY4VqH1tCZkADS/3d43
h9XRxqpkbXToTMrpI8Mxr02hoyOUvTn/f8sjGR8lCxXG7ky96GQiKgEia0Bgd70u
6Odl1fW1HBXKYf9Dznf0o0gaMo5bpEpDlGGLQsHQ2VffMH8fGkgrNp4Q7+eODB0f
WyaQjj9uJiO26caAhj8/h6YNK+lTrar3jvBGHIbv+fgVWwf0aU7gagNpKI83JDiy
thdj0/oqheHocORdsmbNq4J4rROPJF3HgVyOm+vA3owfLU7dE3tyWPjssf//YbDc
EUdDpXnV7WhtJBOy8GVTWYw0SrehHx52EWAMiR65ONFS9HDhQv9TTh7AarZgPZbO
`protect END_PROTECTED
