`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hoNMgn5LsZ/e9VE3owJIYsgP+1FcSQu4o0ss07m6JDrA0PyYSruAUsVzlAqKGM8L
9lNwMKSYqoFU/wy79tBbZrudLgGGzWs7N9wJ5v2i3AakWx2DtnlT/HELpk4Q/tOZ
6RT5sQHRssCumfQgWaeYmyZCHHw7/XeZtpvyo6GRTCLurEXNYipFpkYVm/rdpR/o
7THS/nook7Sz2eIecdcbIMj2q1fVdEmTj0GUeYhKvq4UwDkHWoCNl2VMFYs0OC6n
vv5TGakofZMWTV5Amds1pqcgAYYHVTwXQbinFRpyZiWof0z6uLZzz7opsb//7b/c
p7celwtCpy3iipZ19GzF1K25oPTCevLS2Mvbzp6wXruzEPTYuFE8lbaLSEAa0cSv
dey0nvG7tnBuGJo+izfD5o0sy2FT8Sb/+Ycm+W+TEjIRISf6Pq6VW5uMG3dbI7Nt
tn66VXvVqMTpBZpGScY8Rtp1tkdv589plWaFcZW7weW2GHYEXzqiwXDCHNWYoTy1
ns0/ZcSJq+nkUKaJFYxcRocpgP2V1B9rzl7Jce4RnQwYwyORebvFsTRuZm0wAhuY
XS6+h5xGTPT9Pr7mSkUEXTx+3vFBtujCqCN14l1GHSTR4q4LEPiw+Esmz77QuvfE
pVT74qcRi0BGgB6tL2TrUDfxFLRN+zsyjBuoAAnJdE9cklXu/Ad/osHtkyfGkM1a
9/f44X4snQ2LEEHmoZOwO/UWPeKf4Q7MqYPZmP0T/XluE9JL12NI2RpNpIrgsXXQ
OWKbE3OD6AxKYGUkQ3ik9QS3qboY736yLdS1qj/nMWLQVw3J7GydJ02kVsBFl5N+
7qZ2AzvTL46EUWBDseikSUkX/FQ1lHQgk6FEdhkxMvg5QCZJ5d80n9fNP10BurZn
s59yvs+JApQqFoQ9VOBss3BYJ7t8f/Z6yD4afl9H2OO8iv6GrxRz5GPVei6F2A2T
Mds8peGP4xcq0p0962dUjydR+Xwiyt0XkoidQUZQb+5LOSKsFaD6g7R8KWWQbFNi
ekJCr52aVxBMoHI+811c0qf1ITJaWdIcBlbRIwJYp0V3k/Ifuvuyqlt/KsYaWGj6
QHAu1k0OzLz9rM9xhQ091fiqTBojuwANxPtQz3Jtb/WgyqbCfxXwxruaa6GO6RW2
1u0qANcNZr0glG4e+rWBIBWPScr0vevsUwYUIKaUgm8E/f6PFR3hP9YQFczoX7hp
oPihjp4VOAFVU85KKf7bRWDog1AiUzf8Z+tSQ06gFcMHoHAiOm9gpEQgTchoUK63
yGPuRkGa45eQPTWk1NDv/gCmW5GXSCvDchGE0dSAi59k2oW9y32R0LoyE+JD4ohJ
eftwZkbruBSCGBJQoQG352k/KdXXIh1WPHRbYNsfVt+SDOLx74QRYYba0iAMpYTG
hg2ARgxJUvCl+nYjQm2MkqrcMHPEyKt+KFYBhNw6bZcNYDz0a+nJnb/ADBjm+BDH
XCXvZfFx0p3TVRRs5MD6kDGKP91tS7Gn7SZDglHAviYmDxkGPgtjK/IdVrKU5jq2
UTndiOPlXsycTD3Y+VWODP90rmrqrhoFnuVNy3DsiiXEwk8tQk+y+1zcJmvu7ci4
bW/YAdWo7y8BZYu7fGiBpKYc9Y82tD9ntOt4pne2sptnrGDmR2LCEYOdsjNhnCku
cd/MBwffbwNoJFFC/8swcjE1XQqTFLfxB5eSKmeDVvXSY022TzoKuYQ0jVQrjHDa
M3MlAZBAqIaSjEWN+pjmfHy12oH34lIbBBnuYHz38fMSj2XbujDBhklL/0eBdeKE
/d04C0brK4/o5R6BPcmEael02AwB532iLaPnhh1GVHK8UPJT+Cn7CV/1d1Abhf+J
NUHNqiel35KmEdvMGWfMWphRgQT7g4APgvo2uZjmS/KxYsgUGI9yJcmwaHYKYApH
5+QtKUYXUIn1JQeFPi1BaFa1BTcWsUyAp+PbyARfbZLjSplfpU8MaAoT7u1uJT9/
JFqtfjfcOBxLeZemXtqv7jn5ukbE+AraIxBkm7XurVRn0rYZL+46Sh2kbbMce6Fm
DafmOWrjM5BvHiq8FZwBwUdXNdTrwwiYNkW/dXPkEzEdssoqoi8I5Ii5PoAmESQ/
Vgicwfs1WDcWHQR20G8xxCUnLZhpjz+U/rRtOEle5aywI5Iafj9z5xpSxx4feToU
CY/aL/mGFdsiBdaoRQoXQUH0bCfhjMyS6cJQHRhbRx+ILvvnhdL2oF9O7AjWIC2i
3wji0G3GN+N6sTFH9EekC9/vXZLx7P/Pe88MTmZMShz23A8HXvgVtEHEFAiCaoPR
W2q0zaN9HseazywHIC4xOk6WZH+CmVtTIiRLaOF47bTtQ1ew8kqXUJA6P24m1lFO
gk2LuezQeUm/Cz1IViymgkSHhNnzpYeiEF/DYxNpObOvqL4ucGw2MBeXEgbKon47
v9V8guZAIk66iguYVgv1/u0Lp75ySbn/bHD/L7BaNKaHdH0vQd5y4uPMBam+HBJe
IVXtJNzqUAbnkftV/T5r9q7Zm9k6hYUcZAN4OojFgvngQAed1GjKxpq7n0pZBRrC
uBM5hRykjtaybS+5KKPcFzL2cppQQqaZ8G9kFivGQmcb6l5e61ty74DkN3OaA/i0
L1McuEJFQQjIpz0hgaqQhkW8ecSIw9SZdAxhImZL76l7KivruU/zK7PUIDrz55x0
Zv/AIgJwtc5RLi3r4eZhVKjzhJhz3YedSssVOVnCdmMXA3mUGyFQkvnsURhG4IEl
d0YS+fsvEZUClYkxv4+Jo2uz0TS8xmQ8oMAvwOj5N28HuMIddhFtizI7BRDBq8OW
g+U3QTRqGJwcZye3lS62KAXGhyTDFqnGerGDN1GRYCV3TsZRpdDhC6UHwL4yeAFb
go6Yvzrnd91pFCRAx4aQkWukj2krt+aQbItQ3r7CvluM9NdspQeHSU7XpRYhE9cE
CYWVbaiMI5d1nE6X4+rEzvbCPSbcJIKquhJ5HRo+77MSnTi75CdUVtUfRfH+GtDv
E1/RvSQmoWoycvBxAlYLUzAE2/ScPyHPXSj8L98saz9ehKCM1y+ooMLyKoE+r4Oh
ZKjZLeYqWGzP1ICoh2FhPP7ioXM2Rc4T/dcjlNckmDt9cH5qAcOT+gydBWIiA+xC
yYqu8WX7ivrcrg3kULIQ/B7a/Omx50c9/ORUoMfEBtavmwgz12GoRPCoxVsCcRT2
xEKBaZ+msWrBScYhLZljYVNc5w6r5l/cSrJ7MQZWtdkWg8Kjpll0RoA/LGEoo+2f
lBtRCR9fv2u+Z52A0zI5Q/rryGvTrN46RQkjcdsu6wyW6I66jRgpGmqKASY78x9V
Ek/2lf2/g2LoV15XaHvXWVEmQEdenyuhutoMPXBTyL+/8HSww6NEy7JycTiR5aX4
P2vgFUqo/88+EVS+o0UMr6uy7Zoz2uvCFt1g+93ONk0i3MSzyCppUvoGIg8gHFvc
RbDppCtfQ3gnM3s/kTePrmP/K6e8CLRxvrjeFMNAOUCtl6hEHlEHnf4zGLN+Mpr5
NXrCX/jJIZeScigkCqy0C43xZlsdBEJ9mOtwGVYMdQ0ZtESMog6PZB6ymBLcHxM4
lZxI5OMFVByRaMx85l798HnOwOnU+Bf90BKFf3ZBTpKGGmKkwawD5WkXe9YA3yju
`protect END_PROTECTED
