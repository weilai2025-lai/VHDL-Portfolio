`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4I3f3SGKCmqft/2r256U4oFdNx7Shy6LX/2LoWDdLzE7H0KQbmXbrUD2GpFalh/u
n1YAMlvnbXJH+GYXn82PwHSBiPuAcsP7ewWXmMdqNTkNtOAwyvCG638IYowQObZO
tG7QHt+IcqZkFz0N2BsGJCzpbsKtfs33VHfpTjzsFRfuHEd4jwJJCaOf0aXxyeAl
DjZOg+puOjhb+ombFU2snFt0MKXzk3apT7pYObG3sgG2QaCCWfg4V1eb1wWGOFqw
vvIG7CmlKdgqEYLF/5YkQ8kWlafb8tABgYwKZrMPjoiEMP7/dbgMMbKNoO+bWpMn
DxGyjW7EfiAzyKJdUfvhoto98GbGO5LmGE6kxu+R2nzzqevlNaMdvFjhq2a6p8iK
QgQkPzpJqRn1QUbErsWZJZRxqpqh9l6XQgrAEqAE6L7AIyBSTBPD9BzW87KYV4+b
WDY+vifHCJ+oWNXt7INAcYEa9kt2G9O8/5SNGK7mEYt5e3JzsO4ofDFOa1jTkG9u
Lf3kBYgJ7QikW4q1ZGJvuBlDQyOgZeC6Pv6nVloVSpFQruOIldVgDKi14wN8VTAw
Vya/a1ZDlrX1dN1GodrxBMb+O4kxElWPnoEI6TZCqrmvimVe/sIwjqgFuExmMYvD
9WDJPhZJc2g6+q7NyLA+b82/vxnFzLhyS+cHtpb5aYzzbYPfX5ExVv/NflFToGcc
r3v+2iNiJA99d0aY9EiphhrJfgjcFUp/+artSP1VYumaeZ+2VP+RA9yEKDlV20h8
5IlvdX7zF+RUx/X3slewh/tUkLwPPxtCEq740xDbSfMjfOR8aQP77OxD/HgAnneX
1Yb0zC55OOvmgTIWPfuOrplWA7pdvt5exXZ+IrbAM1vdzYUC2HsZu3ZmpgJa0b+R
Vd20AfO3VHsKx9aL4Ca9o8X4Z8Htemii/TyVgSj80Sce1YM13rOYR5pOtk9R09Iz
JHaP9UFiqfqi/A0iFPncVp38u3i8wplzR3dcMGpd3wtpGw7rGnUNfPUJD7AGQ6t/
SB2cEY6OPiY9ip8/1OuP9bdYf9Hd2aIkEGIYOIPhIlQZWVnt8e9c1yTL5NozmDph
XEC8n0ZPsYHV+YkxGB/PQHRG5drT/3jgHE8jpWW6oAiHMoOW/Lb0fXnrErTy7wAB
gDZsrk+dRMk0U3BjCb/gPzon+XSWyvLheQJ/gOlGsGxS8bKlbwtQJSAfav1gE8SE
5ERF2ljL12ZWMpXx/3cuis0rj/8lfr+x6JTz4TQZg1PbH1nn4TJs/ftmtlpbJC8e
kH9TSky8NkdP7A2Ba2fXhL4aGtjAc3X/+D8vIi2OhB1RFN+yoQAnuFf4e48Yxa6e
+909arDAIgCNuMKvxbN0zSBG2BWxqCy8nhYQ8SapSJ22oQpeDrxE2guTxW38GsG6
X23DYhsoGooNjn9oqzX7cjudRI4qg6s+qJdyRzDmF3IYU6mXpIfZk65cTQ03SCD5
RMEwNNgI3CQ7KUE4FToGMf+JpnOswRFnukGrdgPwisYciJXkW3AfXN7+64yQFjh7
rNDqu8s1kkwrpzXADSPTA7eQLhXXUI5UoWl1ZnLuVRUSdBvf/a9ZHsOehZHOXX1I
VdVPc4pxizs09MS3XznbD617edBz8QMcXMBouFsMfDras8oTYgWgo4aDPR/dAxLL
koNNS3dtZLufR/6HZG8yOO/8jKpFEQmbJF7w5N6VOpBHo6H17BKyDW/+92MRtce7
07hEItjt3nWFCOfmLKVAwbOD2kiQ6/edy2DwpImStYfYq6pSVrhKmLAvenc0qR7n
8hMd+vDDr+I3jfONVW/BiGXFepzO1fXrrSCzIcY+c1HcFmFCXw7pAMoU2gnh/6UW
wMXO/1lyEtctZecB/vX1dEWfpzxfBeAHc/qLmCJ+3hI841IszR2ZK3+6BwjddRSp
yt8C+1cVcyDiBsXiaTjk0s3u8CxctkUDXO4fheyebh+Iff7bMbeIjkKtajkRIxK5
alPs9pQVnt9O7S8bR3JHw27gFAv4cwFlCxB96DxrIsJgCaIGADtwyZ2HPj/I0aVv
9p9JxzEU9DzE658o+x4/4oQZOv8r0rDkB3/ee0SX/jfpi/1KpJoImYS4HkUr9HK7
Wc0P8qSQCSB3N0d5/X0KLPdJ1zyLaYRQid2hig50uDq1u2MnTyZTQ2NZwhBc2c+5
IGOjLQ0pq8xtXr33rpwJnIc2MCJdmZ+8yns34FXsJunp5gUxO6/Te0IIgSsXp6tv
WO8Hq8vqMyRZbHSBcMGKl5SVrFqptMwA7ULNQxvCtnuTCmYWaSIpAyGTPUr/Zoqw
SalXpxEX4RolnzuvNHn5JA97j6K8COT1jbu3NDwtLQpJkZO1pVuObTxhNOIPXIPU
5ry/LPWzqsAiegH4tCl5Nl/mHEMM3uhgMMVtS/kkYUpJSV2SpHlGISKoKFB2uUHz
oCLFm9U3A3ItCulymXoBh6aptsH34BTmtWI3rUaDRs9cuKyfPvaWVSJvv/hZp8/p
wnYj7zlsnIslhH+fVUmrhl+yqYfDm30DRvjsciZ3z3tthvdjILcFBn3Tmu3EiVHx
nzxHuJL1DmszwSiF4Mning==
`protect END_PROTECTED
