`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ucv4ny6qM+fsKJ1QgXAYWi9iuLLd3EJSGVoAxzJI8L3NKElEPtASYfvBC6EWqXu
9TsB/SR1+RKkgafdPNqFiaHV24A1aETZ6y1keiYt9C2MSv5RsoyC2HADTEu+gGjN
d4kr19NnrJWlN3wUJG6NdkNC6HfPHJZjpqIJnF3Zn7JjUjrNJBkFjcME/EO326Cr
QRBwRPFGnLXP7ukDwqanAPA5mvJSzOlM2mnBIfwYiALMh0+aidTmk1IFV2xxB6xt
bLtvEQ732+yYnBPworXFz5esCG0OmnY3rj/LAQMAXfYcytiAixp+IHzMu+e2LVwZ
AeUkuu1dhbx6+EFMn+Zj56CxCE0z06qCPht4M9FxiYmyO7zvRKR81jDcUwHTj9wQ
ieDa2jndi4pHs5kh3R0581rSJH3sUnRdVyAWgWzpNTg7jlPybjLknApeseSMMERK
rszZBYWzgRGbTHCuziA2clKNOwGG6O/ZLpltwhFN4BUAfUMXifM+cfEWPcE+v2i7
Q/a/mcMyodEbk0R4US/dMIiu84IZ6vdIukae5+XzHDefRxOrW1QFgsKLSENcQIlu
I4cXxDAFrDFYOSH4EVScJ154rTsX9+rH/k2jArGM+LvXq2lyOVMhXLh0U9lmwsrR
K8dOOHEisUarXeIqCDkEe569dqO181XagDEGhXb3m6fchrP3bT0hraSKwfGWYciT
xWh6CyDgFw2lj+9P8LZCUQ3Rt6mTSZTTgsGg4+XyreboZIQd70UHokSu931RqlFZ
WZmC6/TjCt9onoAKrO+W1Q1eXU22pRDUyImfH5wiKP7sunI87642XQePO2ocGKCy
ChY3EP28GAB0KEnrbEu+pvGRryeR7XCoWzk3RtfkJNxBe4+Rsu/ETgMziut1GOXH
Jkz5xyzNKhyCuaANc8K1zBRNAXupmv8PP6XZatYdPb6/27sXv9NEpLnmlez8VBJD
FskEQARnFIPuiWmFFsphoDeysnKQVDcrgfE2RgBftH0/pZmQkZcxhFsEfxv61T9V
u694fYV8MVUPde0d3z9mD+1+k6krD2JOFnWtZn20T7bqBqRSvcfN9PtDzjXqaIJq
s9SwSyr0SQ6QlBdufnomAZ/fZ/PpsDqNfLrSCRonttzfnwiA2G3JiXpmZNnntUbh
EucKPnUG+5jqS/JPY7N5heY99coqOEuqVgAXaGkCq9vZRa+aSjFNeS8rXLuT65Pv
2lJ0PqRxczST/ETkab1ocRom2bjmppkrM+judgGbCBmoCFLSR5DgKCIEYsLT5fyM
oLiWS1h3HrmfWm1iuZD2PyWxjHRWWc2q/braDF/0Nk1Hf6s51VInL4TaIN9alWLg
rSlEYUwkmncK81rT49Tmi2+LcUju3b5m5FSALRWAZwIoh1RXREyFbMNnrsbExTbr
7QhkEjJKAwkZ8q1gU6qNjWsgBxxp/DKP5A+nkLRYynbOBnDLfwwzq2n857JMqYF8
0E8jZPgl7Fpchy/JGnIHWAFtZBlQnCABUnI4QUC1NlCF4kPro8kAEE7OY8ALLTGV
Wd2FNSH/Gp6uz3tE2Ek6raKaTWRjcWMMxLmmhKUaGXcNYOw4KlU808LN90iMXJjS
XpWr6QrsjEEJvSEu5i3gtFa404k5U6pf55Ic4jIBY9LheWREOq/FwP6DenC3cU6/
CS7p+JOayDwNCy/zklmTPnoy5nxypI82OCBIV1mPCIcwZ8kJxP9z4H5w7zrXkqbo
xPkp2p2/Z+WqxOtWXp3CF55BLjdukCvNEezr+bm/pxVrPFHOzY/n+Y1h64rP8Xbu
akS0e/3ydSz2MLIAY/ABBSOf1Nqezbbi0beF94ET+YPHYMet9yxa+97rsGYnZ4yP
38UHXi1Q3gfDRy8WEgt7U+9y6E+RwgJ4JsZPDgvhLexPnXbCX1ZnnVp9K35fK90d
6Jj1Y8v7c7ReTfsj3eKqvYN8p/G1cOqWsks+XMLMJm7ybLpQOzMCOFn2a6auJv4p
SEhB9622R1jOt//PSGWlhrn0zUEIdohEA8OuJK1YgamQOpt4N+QTxct9VCf3punD
13Q2VvKUcBIoT1hvdlPscPGiTqXzaIznbNZ49qs2lqFyhDY/kE8tIHHYv0j201jp
7jfiafmG363+GlavZpbU3+yDWFYBg02VbJsNqmeuXLO1HPecR/ecvUsuH70hsjPF
RHrHj8tqButnKAV0FavxHxyl45ZNqyLhMKXQMVasQLjwqChxiNvOkleTMZjyh7I6
wkU/y50Kd3UbARR2N+LRI7bGe29yf7iVk1hBeSCXxBXgDreE+ySMUCdMsKR5BaPu
lHrAo6Qhhf6QT+J/3tSM4MK5hQn7l2HOACZko129ZI6OaAPZ1bjEzgEn3XQnayQj
s2EuexEEV8gLylnFNGW5EmDzc/AYIoAXKkWomFiGfrw9xi7Zaa7HU8B4usDIsGix
agZBCoLhye5AAdwOg/nihsJTnCaGeJfAM3sXsSp6yYyIuu143/TEiGUKNWFy3VeM
0m1r+t/2mKn9TR8KwTlzijkbge2AZZe8a2cLc5j5NtaKiGgCvWegHr1zcRCycLak
S2OWuq7Pd7TfOYL3MDmjlrsU52cN4qABXQzdhEsMAwlP87qhasYbTvDF9tRNtV7u
W+RlAXhJMn9IAE9Z/ARDq0PyAg0psQqW50/neJZmVQ1CjMh4Wp5kZKBf5zRAQfAk
RSsZZkPPWSPZRkhRpLDariNa/2QiB5qrfhH1K1RdclMUhCylWxsoUYNFOdFz+/Hv
w3PqseIDKwgCyb9peX9uwUOdabgMeD8MIity/a+fwcUYjBLgx7qtEVgOabS2jRX7
zmcraxI2Cy4XjEaIBavy/pZB9nCT8cBTNUhY2+hhabM2BK+Ic7Gea3dHP3+npKaz
bp7RAIm37y7rOMYtPBNFXfMkrbBgDBG4leF4NY4W+xFEwo1hMJPaJOMCH/s7/htX
dzRWkf6ztNjWBtENXGw6V/cgwrnQvB91ythafbGwhqdS/CzqPP1dIa8s+uPHxbq9
Dwgq639zewCiG9zv7RnRTaZP/pvGs7esWClZ4zyHcwZttf0Rmc9q9I17MbcjHS6E
SkPYZLIfVni4/fsHLUo2VDnbLmISdCQgHz+GyKREv0wHyrPhOzwtGl1jI+0igloK
VuwqAdyYvIg9htrFBWGJChvXZKfJHmzZrn8+TaiB5kEbGvUnmA6axXKFOdX2/kuH
L2d5W5RDdjGjOaeqONW0C5jyfai+FCtVObadUiMuSbobHJ+pZsn+5egCCdfPqIoW
1cgmRpb/yAWadd1FDT+zfbIBulC0qglNTa7UzKUatfco5ouV3ZFcWpirGWUJ2Lg2
0mmE0V6WfUn24594kUdkjR3Fu8PKR47h7fdlFTfaDQCixxbQQcvUfWdyCULJdpZo
rLQaeAJgdaDnQiUk/mz0/wsXxzeRMFww/CdQpqfBy3Tq/etn82itOw86anqCWDq7
7L7jokLq3rMZyTs/SqeH+7SyjTRDdpfe/8MdTelzGBz4SPYefu1CnKCjLIkGRr/H
Pstoljxzl2kx0+Z3ArR+qCwonbh+qAbVZXFeaLbizMSRKFfvMOsv+z7wM6WBURJp
t8WwAjdDxwOJPZtpErt6InBrT2Xs6uBiuzEtgFmbLsCO7IanyHieWjY3mRVcl3Vo
kJw8TmZaEZX5xHow0NCat8vQ7Fn1T0WNFxoMAnkrze9LMvrkW849lukN0bMvS4Xk
ru7Doatyuf+ntzN5EdA0Yrnu2qONFxyOx9cssICQVia4rjN43fqK8P4iPT7bGwuA
M7BYXVs6dsRTpRCJIWolJKW+DxZ/FbO6Xqv8wFQQaz0HPfYUsUa/FJjWRIw/HsMC
UKw9+X4K0YQi7ZkHIXA1PIuP3V3nPA/CipEOFecv83GPv5IM0PoRjZsMId469SMd
TW5ksoOdOQ4YjQfhsI5RgNGoXjLzr9LvMcnKa16bxgaTs6Kw3gQToOXe9kTOqNHS
p/hF7bjWIZh736oydlP/Zd84XzyB8WpIIsQ7EyGvrUDm4Zkz+OnN/sqXFHFyNb10
K6+WDvERUVDvPhQ51EUFUblu4yk4jFRvxMbUojjSoZ1gGuGpYOuNNFo/X9QtZSLQ
+mIiJSFp+Z5xdarYGzBgdYPzrByw4u6ObXCv0X1dHmkti3wBXdpKI03C5jBYYLX9
6fOsueIWkLt1Z2iUNxWQMByPeanuISQSVzme85G5wuoTx5nQIx9I4UBTLqeA9MVD
jdspMgnjZahBTUNGvHtyql40/CNgz4s2uG7tB/aXeW/qh3jgC7g2dZuJXOj43eeA
t9BvN3FyIb7eq8ziXxuFN6znmcDVS8pMxsKN3KRa8Zl7tnqXsYUwRIBjz+tLykes
/i0ywwGGIFPhYouCGGJrQBCpKAdc6IeioVHnVwqYDdNljN5IDmwARehBAUDxc0nr
6mH/OateTFsb1r8imjdkKgbJ3zkVw/bHnECpFj036vmWCcs/Jl5rieM2GmVH0MZF
qgdDtg6M1CMcaupofUYEc7NsrmMyabrMUI1/LAb49g6eqJcNIt6MPzRccUgGKemR
HdYDnTbUukkZp5pJH/oBvj+3aSVcIWn1TFIixwAwDv4SYEL0XzNvVpaK41icBpLL
GxK7mozE68/46uIeqI/i/i+Z7/8V58/u5Q3RbJi9SGkqChPohKIyt6SAldrlepaz
XaoLgSn9OCtqMKJ54UdjLOanOhPTkoO7/jNq/sKBQFY4/WzmHmX7GggZOW3VOa/B
HdXDsYMVNGaquawmNGqc6y3SSIeo6RkmWLpGNJAuby9jFCprxnSBQwWGeN+wYne1
eSBOob4GEgXV1W4Rd68uUaOQdvzhFs1G7kFR7JU6UwFpZgpWFjFSrLo3Y3Qt4BuK
DTlnZbfKireCaZqKBJKFqTA2cANTcawICYKrF8jNpKJnGQmOAiEsJUsVmtFQW+3x
yJH7Bj58gmY3I5Mx0i3iInKuVViTGNLd3uTeIvG5p8U4Xq6S5HEGHqNlyI6ka9nB
zmr4lDVC7edPu+o4j/fbvdF54vlXXEGNJTgy43GhurqilNX8ZVpanfkD4XXJ0UpI
AfNB060jdYzsJjx0yGL5YJ/laZ9zCcd96kDRp3j4LC87L79TwW+l2TDScL5evsVR
YyJkFBIa9ZI6/rDbuOS6khQSnxw06LgE5lZnVINut9K3Pne6Do6CQDWcGwd5QTqN
XVJZlSiJzOlAKHeyHkO9PIlOjqieWZT9EjNIg7NffTAhYRTdGpVEmm9zGkWPjzRc
cPTe3kc3SeyRHdkU3EPlWSAKvAAYSgVuMtq59Al1aRvQWoJa+Nb6SiU3VTxf7eQQ
97cABaMmP6TkCk3fRuQo0diky6aiwzSBsFJ0ro+u8DG+/rbXZIUAOd66dlDbrcAS
UYAEsrVfgS1pKBFmTO7nA9ylVYJuIe6EU5r8m192PgIsmlT+aaifpfBflImnxUvL
IY3bp2j94aaWpH+cDTIHg8+mNTaUW0UC9u0UjgCArHms/Dz1s7gxds2j1ZYXcqWI
jB33AAQVGCvEyKFUTu5Eb7sL9MabWJnFN/GNnho0ehyJEIbJikRaC0UMZrkJt5EG
sTbBOWRNecrrD+kZT57kwRg355CeyOXiCrgmKTB20vDEDLZEb39r86Ww/pmEpHp/
DLwWp51um/W0jrZPpI6L6oN8SygdhHXLSfrsLSQZ0eC2RZHQP2CVmHCf7gMOLJ9P
F7qrM/RcQwze4qenyroS9BvwQ5EAe/yikMKNx1PoLQWkRBhycMBP52sPmekMCOnO
XED9SqZn6nnsvBTEhlZRyizzosvyrq8jNYQNLVDZvVJlwLs0z7asNBYOHkGW0jw7
ruL47M6cERb/WoXjEXTcb+wPw+cltOH16QZQ3i7M3kmi5jENAtgH6uWNzM0LuH8j
/jnZw9UQJKvu5Ja5piH+ecof3dqLe2yadoIa1dxC8Cc0dTgpZYXFeFCkykOj7B+U
BBQvqvxynd/GYG5XdcMC9sm47CDB46NbANEwzxqS5Pdxql7beEgHElQG5d00Sdvf
M2LwAmY7ytVEHJjX/lk/SyMCCeXDcvf6uRY5/ShZBq4fDzf1+SbnlsRfcDpybwkd
6ibieGxifv46eYs1BS1ly2z8tOWzSYTSnRJ3NuXZ0p/lhTINXDEQwVuANs733zjb
Cov6V3ZveApD4FwFVDGRopuZP+ehjQxyPR6PVpJjkYzcqy6d2gJxWIlXxjVXHAx/
HU6FRZ0rESriFKJELxX0I+x4rnBc9gYYL2e0VVBu8olvK0be4Lr/EGEocXCvbd3B
0r/YXVznlfjOGXyCoAnO9Si4bD+V8pJz//OcMyV6H320SZD7FnqxHZYeOcLYuQPH
1U+l1gyWCBgR/Hrxp/xEkaYUafuDTx7hP0norOO6Zzl4Pvb/4oFDTI5YWB5mELFV
ed2g0gVyWYUVpK2ELUpxFzQXTYcq8y4D48L8JW3iq4cP9MMXHUWnf7wX94RqbJQy
nl4qSCGO248VU6LGyaOIUE6U2GkBufpK0xmpl9NisllVH7OQdmxksCoOhKFnvwga
g8eGbnALBoRjLrPO2bHuRI0IKctZee7CtGRzg8Wo+p0X3dyHMifypzE8s2Cpu9zf
JQaepGAdQcC2hodgWy2XN/L2E1Ey3pY0ljtxK0DxpMbtG832uSNLNxG0VXixBvoz
1k53dtRuuOtI1IZ/wkMRvLjXlnijVikTN/DAkPzrzKAZcD4tcIiwozY9P4hCSvy1
aN+145Wd2TsDEM56UcLKo0kGkQ53sBGDrEhIckLahPT2lOhyuJ0l0PiVlhWPqaZ1
stxf3ROqqfn+kTbuw2X2eLzCg47S2LL1xeDN+rnO+bMJC9xT9xgLqCG2WXVItoHE
nJCDqPDgFRh5tiETaQLPZKAsvct9H0JpzXoZQH63FaERLS5Dnlj3WY2VhOBSE+HN
xEdNG0/Ut7CBlQMuRIdWpov5vSkGm6zol+n6+xucxfvUbq7YqfT6ysc07xURxqea
lhEFVUVr2kgPb0mmSX97Sib9xP3I9Yw5A/vugoXL//Rh3Q3gmH9zQuVPLk2UCIm5
t9aX/hLL6eRXKoT4psuInOeXWw1OCB/IUgUqR1DQOY3kVNGlcmE5WLqjANIo7kdj
qyxSzimp21h1fazyPNdHYtxxjkyFhw2jZ7oas8eI8icTYafxSSepueXTQckr9na9
A+wNiJFPhRa4hn+1ZOc5igkIA4akgPNe1v9ZRFz9J8MczEqstkHmKKhaUWbKBFY4
XzJ5Y0MFQt2ZpDPzg7Ktwz6V2gNXS6sv12ucgP7dKQ5oxiIxIWxEqLn+UO+VjZir
stwSiGOwr+WcXgF677AJz6njXBKgmtaNnGhz1DuenQnCuM31XkfBh8umqGk3VLHC
HmUjKSmc8d+26H1IrZnrmiRSZuQ4MHOZX8AnNq65GnLwDk+G17W7Gkf4udaKLZhg
f7OC7JuUmkZY/yHuvqlZ+xS4ks/Q+Wl5UMVaZcBF/4EAjbO4gl9fnLbgifp9uj6v
ap69QpP9WBPjNeSxWiDSyi701pDjZd7F0xrew0IaWshtsXTdsKAwB1HDqnyDH2kX
9SUg+F/gPI1cDEuDKc+TuXf2EiIB5HCw4Rqw59NjYA4hL5Dz8N1K7rPVNkbTL0z5
3ncISRIoLtk8syJ5UAx35zo2l1g+kSCwr7CNj/ARw5HutLPpL0prUNJ68X4CQkWZ
8xWp13pVNfNF5ObqxB7f21llDKQGji/I/Pud6cBX42vBMFHa5vTHZQcdFgr7ByBO
KM+L66fwplR/wk/IXXhhi0KItevhcW68OE3hfo6X9vLhP9uTYQ0iAPWSFfAd3pLy
P+qRsbyYoLI5n8Rbp7QECZdNz5SzRggThP3NJAYlx+aJw6vtUqjcoQsoyLjWbRrU
iKsyasrym4IwGPDsyxr2EjuVSarOADv70xoLJrzGvUBAhPmaV3rlooEBsAx2DsH2
Rze2JfegZRbgQm2K60wZxwBnJ/jgoeaMOEVtt6M4V52pzj8zpX5NGeuSBwF0ZJC5
kByrTAdo6R5UFxZ/AuVcYLI9/3kysKjqhbe9/ujaNEDzlC0khqWNVy9kP3GdDbNP
sZrbvijdbOGggJ7jG0FERrGimEWbG5GRqY9z/wg4tOcCTl0uZNLv3clOmxg6DMsD
VS7J6PWvBZSutjyrF89lHBoWrFG9VdUX2Ec08IFbyfrk6Yfrig77BkH2/LHhcovA
YRJrfBb34MZzUm6vmnWuSrMv+MN6Tz4btwFyuMKF4XsGe5V+6fcHqTDDEssO2ZbK
Ux2SGr6Btwt0Te9o5/ACC/AUIdaUs84X+SsowX/iwUgtT2ryoCqN2UxU7+Tt2aZ+
LVR9B3In6n1ZbTU4yZXV1fBbm5vcLkEbyZcGySBPZ0JvqOMap5DxnRtWOv2uk/Y7
vzxpft81W+HuSmwZJZNznALgrYYipR+eucHE6MMi0lwNFXWtPyKbh5VbVthkY7/K
JyuTVZS22T3qOTvhYsztvekWKx03yRYbryoTqgCXXv2kiC0+VFNorDr+NQ2Tim70
xSyozsZ3K7GpR5UGIgTo+TAIDOWOecR8KpbJtXO85JgkghTuBYxGMMp152BSrQ7r
L+KNWNa9EvalLf1fzOKQnswSgYn47faZRMGtmCDR6LBDoh5YKGms90N4PhfJmpL1
dC19SqEaDnU5WfKqKZI9q/4ax3z2UsJu1wISns720TnxFVHvj6dfWkXlciKUw9oj
y1tyVhnLdoLccfh/sSy/66xlPTGsJAKt+7LsQfmsaelvgDaoN56VFCK/vnTXGV2U
Bt2yq+Sci/DDGm5vzPMxKs9QxpExqkfOBqR6fa2PwHwbZEd4gSkgMlwYVkpRR9kv
8DXxWjdqlhj23mSNRds0CnU18vFuXlV8YmKvExFHsGMCx3doxiMyqeiEFNO2f35P
0yR7NM+JLtnsSswJm25pz75n7/mkRkZjTP9Xu3ozjQtFiXtS82qib8dhqbxxXK9t
shn1unERZiZIxU17BMZ7+8PLSMvUrFk1yeLU8czskU29u/Pyk7RBhoJEHw4ZLCAt
wv9PrY9bh72YmSW3cVrCd2JBniFYJyv2/G19WASMwTwTnImeefUmG/r6N0fSh6XX
fqpgpb+MXfZUCgqv+HYHQ4O2r/IJJZJGaxjSnt4MTVhwhpmtqnlFu5SpE2Y4sIBk
vPYvXDsyeGMjIMZja8xyHOK/JoqsBtcayMkm1C9tVbgvO/fyng8sgCk5Y8qg7Br+
ab3S28QFeyzd6McuizIvzDbwDfrQeOwQU3SaNXK5l7Z+b5Mql9aAWDnOoyCa6oR0
xkn7ga77ntXosQ5FndDy+aDKkjCCq0544KvrMZngoymLtqsqrP9IRVZFhLVYWqK2
AyXIRHoL6G9Mq3U6gUuy0CRU++qE9mH1H4YzwyqfkdwopERwZQ5wOCSlYjiMHbMA
erQjnxENUzKX7aLeDX+yE9mSwSiT6vGea22rNATbKosN2n0JT3fu1bM6BpaeqhTP
Pi7N4oyHNDrhO+vnjINxqyAB/90+pf2CWdGX+Nd6gJhKdTyJCpvuq1uI8QD5OAFW
7UKFyiUDdMdy8BE1EYK1VzSg2Ceq1ppHcG2smfMEPTsDGDTCNBhnUKWCvkxY4Iob
miPY2Srd/u+QaVTUULuwV3ZtWBxy444ouOvVz9d4zExLnwem5nAYE777mFOa5Mq9
7CPNo+O4HrVskwEJCWF6hgp9TtZv+CmvFrChY4thGcDqdaBXABKP5IglHIl1EbvH
krgL7Ye5VjyCjR8LcnGPs5MwLNVp9LHzgBWvvsSlNHoFY3Z8XDj5AfFQqfEHN9AI
LVeNkxDgadL1/5w8QFyN0VWv8B4JlXm/qtZuPMsqflBYjK4i7V2cXVK1m8EOyKqu
KQNHb7MU9AIkWftyCdDs71EBbNfDn+OkCU4NUUinrSXOTJ39FGrZGJ293jLArf0B
xrNWZeUhLPhUyVBNjTZlfOdKgioiLxyFXDgaGv6bb8ujw7GBmEsdm60HgZ95g6fb
702xOBk/HTm1fKrpQDO3UaxFCIadoC9D6nDhqwujzumTQoUhUDTSV1ywXL8MpPZA
O+Kql3il4neTycEUwg1nay5RCgMaENVVTrWSfEAXazGksCfJJrn9W7qJDXKQ5EgM
1ximnpsIELMdHiLxAl5KMAL7Be6Or137/drpCTNi5exmvPJxQ8jmc8DQk45FtWXn
gYgVa4LiqgnwnkG7zE+hGeeDrq6t5h+VeQN4C/ftQGZy6SxDRqrTf+A20I2YmRvt
azv2gA5D1qu1//f/2r8oC5RA9GzQr5gP1lxaB4OgQBWNBVJ6+6gc1x6Kl4+Kt0I4
1WSP65VLe8QnuAez9QKA/qlrc5yS8++nOv/p4xoIpxFUzPWoZ23njGS+yVi2eb4L
5tYyeRXDllHR59dPPMPDQnmGcrePLXL08hchRTo3vT+Vfsa0Klm5iK4WFdPOXrwH
G4s/QVRYrpRZ8qZl23hgxVqUCl+X+FxKIvRY4luZxPK28eGLe1+rAZ3X/TnbUTXe
gb9Bgf8rD3lkFGQDIzSVwtH43rrIfTjPbKah+//4yfIev10jtdCVa8tC7Xqc/BD7
DorLNrGZ15c8bPoDosN/RhOwg5VbsNRwV4AFItY71oBT+k/K8NKyLWXL9rlFUpsd
BmskwU9FyqaTdXjDJbWy6aUuP0ltis+vXgoezbvUtA9pJyjmPYDyW9CVSKxaoh/r
+wXncIqcldUN6RsNKoM8sIUDeKfDLFePF2AmV0rdSnYdFrJ1bA9UIrrKOw685WkW
t75ElGDf1uklNmt5Zfb41fmPMTbA6husAxTY7nV+sGndNGg5eC53bVFw8UY92/JG
5WUGmgQ0aWG7hqw7yBHAoUXhzqWA+WNE/IxBcaWd5Tg7SqhbK8zAMkIGxKQ0ZEsQ
ONUlLcm2i/M2X/IYqM0I7+JfUKF64JFfONPj+QRoSpa3WWVRXkXiTtjg2/ogXiI5
V1/yJxTffo1xSOSN3szR5BrSckYhG54Qaoxq9Ys/LYuVU8qSC6zuNRWKqOZtxoED
eVl0skAVzNruMgFKHkSLHXWqhFXVtfRUfNEi0q86fkTTkPZV1dcD8SZeV/DYn19h
MAHIVLzm2x0cz6N7lOhVExiLf9Mr46eTNWuXdTU97Z2RLyynLHuF4MVALxYJt3ZE
m+oaiJ6edzZxioO9ZKvLGI+mOCQmB7W4G9lZ65TESLmfqR3k6PCOltv3HvgS/b+4
kd6NZuF5R/guG6MokBb9Gi/pJGk20oeCJsdMBh3DC+eMawzhbann+tq+6xOs0pj4
toJ6g2QBwVV8sa3f4PdxNDHdu3zyfnXbYqQZ0WNuIWQCIQ91OxY4/YwROAG7gxSw
f0kGcd2ftYWWF2SoJ5ngdAz93MzksvJWgm9iGXgQRNMyBX2hlXbFlZqKPEMnVvNy
TJALqc9wgCxu8W7kalYToY3RKkZPsDzfoBgSWjl7WaYCBAIjeBpyz1mnnJR4ntPo
ea/wcq92PjIyFKqqIU53ypRGy7+/rJRic7mM/GnypNi8NtOUZoVky59j4GbOMnTB
HaACb9+7m5bGDrnVAfqc47/iMPf1gA26y7IyLKXw/NgtEe2/gUutYs1VtT6+LyXn
zTy8LCqPqnnCu/MUjdOLRJfJU6ln5FMABRde6YNTLjTSMT4LCTy7w0Md6YhkSL5v
HmuDCEWOOOk63larvk7i8XOyX6EhU5cUcLyzY5d3LAfVISnivHEiJxQF5zLHtuEi
O4drZuDVsFsrFVOXGLVo69nPNT5Iod9LsuxmyPzECfJWLQKDXU9wbmBHdQ+Tljl6
ZzaHMdvg2bRYy6/YG3bwqQgmhXNtB+swe4s4sr8jeR3DXP/wU0UszIrDXA3mGreV
M0vrQeXasAuSF/bd4oZvhsy2xp8kig3R0UH2B8g9jS7CQYRiwc34gpTJP35XgvPU
oxgJqQMF8amVIwKkBUsfXl0K28xrAblDCOmbnfMHJGms+Iyj10eMdETYwrfoj+Gj
0/vCs4JCI9KDiYKh9HDPqAyVlOhANi+Bn87lgk53NuaiLv5H5KXXVTieNjUs/zdg
UH9KhqT6rMdRe9OBCePgO6bXLsplKoY3QMCG89S/Bx3OeIZfJrnLAnuKs6j6K/AT
3VVb9m9E9odk4bsJBzPhbAErF5uEGeT8EMwpYUPrDClJ1dCnEhvPRuWldtuLEOdQ
Jy8iXszprt/0GvM+vmfdTldTm3ROkQb8eVIhDp/pcB+wwbRQqOWMmDkPJmxHSyXB
dzjlAjj1D9pli69UnCnTikwW+5I2WA7kNbIUX0Aqm1flJU98mMTeoxyRXW1KRrl2
xhb4MX7mN0i4YG7ztVfJNZWiYgk26rVUwULX6dLe40JE68bl4Qiztu9IPxumxJLP
9A7gQogbK3BXT2P/R3OVCJmxZzCHHiRZgPg6z8MOAptsYfbqCdsMsoLrnEbUbXvM
elGqqVKlpg94DLnTSJFb6XGZVtRKIIPaWCWXdL9VJpZ5CdpGx/bUZunCbPBKKT30
8QbwYSRuguzprfISso2SlBxxtG6+Diu9tZb2Ua2W2Sva7vj/PoAMD8ZWPxlYzsyA
XTzWTC5komkiA9ld3wUbL2ksxfRYt22Xpz90PvUWpQ3Cy+FacBi+jMLZUs1wKjnw
LrGoWfJLKbd+YWjOFtk2wkNEeUs4GwoeWgvOBDKPXmYkqjiJw2DMMlLcQ9xwiwAv
//C7H8ua2qaUpFAvuY4RMcb6yJRjlywWi8fqlhaEUWgLgMjXbtU1mngJ41SCAhlP
FyvhM6fq/wsD8zgVCrk3z0QBP8fiH9cq5IpWU+6iGGRHGvk2BXGrFBkWdW1GMVGW
igQ+nezfZzpGN2ZgwyhIJTjw0Tfm8wDVncTt5MQ0Ucap2dVlNtf0vcAsYez4R88X
EHXJUsqfw4HZ0Eux0jjBtIziqkML2fFQEFS+Ph8U+5a5LgMMMz1BsOoBjhshWuqw
a/5N3P4eFcnutNE9UMHx6qCjIOf2PDG/jhQBbv/K22LiniVQxgfkbDcku9cRGWRs
Fkikg1gLXCtA5AY8WermIYn9VOiM3rgV7JGeFqfaiLQlR+A/wU7reQImgpO3/wNg
rP6PbGowbNyCkkvPW9+aZG8v4HE98LOOeUsYhCy8TQKU3RnlzSp5J1iCvwoI2z26
LmzERR4P42cAVJ1WUIhm5gUyPEESLjflkAqJYpCdjvA0zUyOUgME4j8ZBjDlV5kR
E28Jixm9lOl/LF9SSLuqOeEMmARPhyePC9x5o/rH5Hb6WpG1py6OVr9iIQ860oXE
FbjaY8Oyx0SvmKXfuAEbOxO02vUN0Z+xxR+yjuA8WKfF0PpwLLGjlfLTEXeOPhRj
tPt+f3GfuFMbqN64G72ZyMbWxe+5Nj2LIWGbmfDEnq0lCvPr3q7x667x6mC2aplz
BpT/+MjaVsvnYk5/V8iOid2MWdzfGk3Yri3uRaursfv/5oHsLhVzF38T9hEWie5Q
W/f4hg3j7J/0/COZB4YieNdvIKxINL8pJPudjL33SO6lYCqwgs/tBaWHFYKyXAYR
OFeQosSOadivM5D7UfErlA0YdgPYP8oL4rtrJlRcgUM3VfOwMQmulEnU0Zb9FSPD
Cd+LKuEGfiVJJByWtqhXQeo4nBM9Y/0oAphf1UsxyvF9wtdK3G/FYJO9tRzQdTrp
v2JSV0vOe96jhuDOcxyH4FRKv8T1TRS+ohdbQfGDq4HTvEpDNzA6nfCGw262XMaO
2/h6mOMTJhjyWjIGX7aHzth8u2MRHjpTSJPPtF/2Ppd1w+c2I5HB7E5ojBi5Yk0d
XtaKaDHbrxvT9vPBdeEydHUrzIWGNh13m9+6P5zcdBxNHlwvjne57gEgGdT8jojq
fptmjvFBThwJW3wr/rv6JRwi3EFxTP8fVAg8KYY8bcjiQvMk9GB0j1Y/m46g9DUL
gUKSWEKEHDIHrhjfRry6U937kulEchHUUyqPWWCVLdpTL8hWOKc3VNSpne4iRj+k
lDjnaN5uSiZOqnz4zswYugEihXv5mU6E5ETdmTGZq+njPzmwIcC0aoMtc3l1HAIr
1hicu5/IrkIYfW7pIMbwNZL/4VfdhDVZt9vR1/kP5zxY+9kIunU8L2oQgFOU/D2g
x0PDZwmiIvzuGML7SwkKWCALq/Le9EeBykcBVVkI1j/QkJDvzrjBRGF6LsurrU1J
UBV+xMXxHxla/0sewSHhK1d6yyJxPqJ9XtjhbbTToJW6pZSQmm+0A+e60PXevNjV
pOiWSgF/SKUx9173iWTXf9lP1suuun/InVVrL6tZ9Uc+1uhUGbppvYS31rinDjC5
PWqmjKFeWy6lmSKoaMkwX827YLhdZTohD9hmnpsX55dERiOUGgWVUbYRPrg0hIup
iXeh4pM9H98VmX58GKJvds7hhnCNZIa2r2mrVljQjH9dwiNL7vXSB5T4lrGev5ha
mXSep89wuPe7WtoB5Y1QBZsXyu33DFzi1I1ZEq1IrQTDuMrGSwSl+jGtfFNO6wwB
xdBxa42tAlN+NjzDmJYwiSQUAFqTr6pLcpP8jyUOcBzTPfDO1A+09krOxpwEsqTn
nnpdRkm9oYqtTxzYDmnQ5ae67yMb1PMG89HXk5T3sqIG6S9rrCMY4IdXugrXb8ur
IelITydjpO7VFNgFOs8c1tKWIdryCxbIjigWENREQVrObN6jzmVQ8Rw5OwWYT6c/
nsDKKqXMjNnypdk23BJedEfayaRexjQvlJrhw9NyMj+3DcBVoWlqZVfYMrY57adX
603rMrEo3+JTf4EIXTVSzx9Kh7JYsjKrm583N+ldrMV3HCRmQREQ0PZS7DX9j5nv
zbvg4lEba2GLhOmF5rtaZGCy6PGiurQ+9vCRUIZtPv1d8D/BnfmgWLqS1X7yMyj9
P4Cpnnc0O7sNEs5SVFZHA/CSUvKL61yaOUKrpVws/TgzjqHeDoQ1eAROYsjzDSFU
zFYZYmI34nrcxN/vWV62t0bOOlNFwuLVHpMXwYItXEJXUHmW0wEsMznIF47lzJpn
ndHlMabAEkN/MHuOVBFiAiADDglKWlFy08Wt8QqrQJFMdg//tpZa73Cr7CjJxh/+
OMgFcg6YdiTkP2gBWC05CCAQCW++xEMsnwi8rCceJGqAzUvyxgXQpdsjOEZ7G/xy
3hlJvcNJbxy0immj6LevHdYjiX+sWQKQuJ/m0S/t2RM6dOD0AURAQP5KfGNs/0kE
64q0WcyJKCgwGdc8/nSHQTbBA2tQmQ6ENV8mG7tjN0oZDiIblN6hzNWR0vtuv62n
hVaGpVqJ6HULjgaE2Ep+Jtz17wr+1Z7AVbUbU9RTkVjMrdGapyDAST/piVVd6R6j
Zyub6HhLUJuoLhEGw36CWKjQjUexoiyrwoAbXazx5AQGZHSKQljnG0z9FImApvOO
vpMkBxXIig4W2REjXQOSh4cHnrLDxb8nZXyuc9cwmrOd+QlQ7SwehfHAVLLDBS4S
YQD0zhR+oDHLkM5qV/XI3b5Xu/qd7/RwRBU+VghGLStvQKEHCXv5zcT4Tnf2HRCt
y7wSjD0L3b7EI5qc14Iqu32+PXdBK6tNCb0LlVYRfbHBr3PEEr58PUtlo9+LTVHw
Q73g56tX85Is8NbFFlgXssshi2q2pgsCH2FtjqsqS1HAkib8BarhigaszSe+qRYS
ce854ca1EdcwJ2T00KhzLpELN9rXquqvnOONsi9lgpjQmP5+tl7pvH947dRE4ZYt
IML8ix7d7to2zKLd+bAXxqXZxZSLm0oglW9tiFmqBy9AljD+XeADnNsvBV3Tua0T
s7Ri7H7PI+lzuJESIteoIFX86DfUrj3O6aXjowQaC3MkyJbOap29PFNOPMwiZTKV
NOg/HzZoR9rvCHE7zfltFJebEfo1bnXE/6UaqEr14lkkmc9rPEjBZc5tTVJB6GvN
J22S77FyL0ZoAkKEpoklfo5kv2P0RwdzZAcdbyk0bA51YeBanPaCWMbSUJXyODkS
cVvqUd+rVCavfjZbtDWrN1rAxdORzWtR7jKYSisQBFaghhbJq6AAdiOclxkDM/y+
fucAvCkhehEK+9GHi3YdQgXv9t58aCK8WtLd3craOnIJ6q7nm/UjFHIvHEt2pOk8
vM8hvHbK70IB+Le9p8RlSHH9lKtfbayYo7dJtD9e4RB7tqZ99U23KJlDDSHHr+7l
fiEQFJQFVYHtooSb+eErEiycFNlT5zdmCdBr8qRvuclfDAlhuLPQe56Qc1K0zSYS
lUXoWlwAp8FwmobSPvOhAwAsGkhP43i0basz5ZDl8Ni9nY0MfUvgxt2MYz8DwPhS
ExlvqFhuFx6vrF0oaQC8IPw8zf0jpbl/skrq0xVDCpKW/NaqtN5UGr7nJLHEH9ks
iymb6KHffSktU8s/5zviWq36NjtclT5C8X1LGEvSpiN3DdBa5+KPtYiRKOTGvzmu
Ci8PZpXN/PHgWzWLrjGCB7km2iDEtkzLNf6O6uC0KAoLPSF+qoyRqDHj8gdd1YwN
vberw5kXEysQB7pINqUIFWIkbCWNLPC+YTPhe4MziH1pGy99HTegwHNP/vpGy/ay
89WKvjRp7xDBkqww+tf8suzzj5yOEldkD7Je1Xb+6cQ8/J2IqrT9y2JVmHcKX2PR
GexldfYvCsz2IHhZl4hQpPyauZxypGk0Tjt0nNW8LPJvmQj5DCwe+iGSiqWnRdXH
tqzqkDU8p1Kayef+Ww7xaLr930UDkYG/6s3DOnRlN1Sf/cvJuPQ2GrbH5BU+wRzs
XGvlKxjX4z+DFkM56+9ej82estDOesUsJh4gqRW1DbX6yM51YplbxclZucJFVWMW
FYvNBIuJ1MbbmczDhTZ/dkJ5ZURfn4CbkFLTquAT/Yzdu/NVhyGoNYm6k4h6ann5
/F2fyeWn1ws/S0NZjeu2nmt8Q8kdVEQeMjX4yAycb+wC9Fa+i0glhPMZURfrzyB2
JrzDFAtRBeEfn/Fca2L3NeE8w/wtJc7U5NdYnHW8yNTP2NND3qS7tRFxTJ+ATZWG
mKaL8iglg82tvvsRmuumKvpZtMaPY8FTBY7NsxMuO9CCwoEjang4z2omqdZI7qmi
X+4utL8H0Jsdy/uNI+10Jhyw9Kmt5GL+fVVQpSmz4QiGn0CkO6ASbBWYhmYZRjqa
9eVD8ntThww0IzcA+XiiOwbzrBGbpgl99jIi8KQCSNsjp4iFgrGArziHU1zCHWRP
NFDliNvmzzclXQ74kFpo0qY1VHm4Jb+p6AH7ap921pMdrStwqBuy1f5btlkWVD1l
esYrl4AK8M5OyJ2UyoGTw/PVC+9ZSG7FwKghoKU3fsOEQ8xmKvW3A3yNoolGzZ0Y
LLsqs8tjKJwgSeZMdBta5fBtbhi2pxvBavNH1xTeoAVAhqnt87qW/em43S9FMCWP
haqNRMznYVnN5yIo4Ue5/9AYI9fO2qo/nRwE7eJq9/OzTBbzOaY7xHqEgWRJfLpq
JzL+fVvzIgFEQmwj3o+lVR3vB7tQuy+K/mRwqSCDaL/tqLIbxURNpAnAEqiVzcbh
hdxkXrMnREWRYE4YYRHRj/UyidE/15WkgqP9yAHKPn+pAhkZNrPRqPb5/gEBq6cj
FrbXFQ3VbpYhA/Bio3VnbylLuZOcrpoMSlpf5O5MMbSMvmaygnZfT82E1VyzbRGC
oOt+0SyR1ZlLSfMJHUJb7jVbfOpvuiBUFAt21S32Lfo4C7hP5dObWdXJDa09BnGc
E+dEszgQGKqwfN0s7q4X21SucdoQkjNJBH/vhnzvona5IeZQTz56jMh5jIkNzPea
SRH05WiLz712OLXEMM8qNSWJ2zNiVJh/YRluzNTddCgqoEWtTxq86b2Z0PlHychB
8iUCB3e7mCUBhoDnt2iSub5aFbMZL9uH+IoOYpztPK0rotLEuakY9qORCbEasl/3
/9FTjQ7cQGeWG8ykkBJwv/6hwT7p8Z/JE3LoOzVJtcghsoQYMuXkjl/lhjgMsEVf
lFXa6XJfBZQCIoYwwGpOfX0iOgNOVtp+mUGp6Vn86mS2PB9Y0hZezFHcCP67TWcs
G01hUQG3vRmmPFh8WKgf3juXxge3m9cEWDF5WL3AsxNC8EkeGoWzMysWBAx9Lfbi
RnG3rnpY0tRKuYjjAUmCvbfEnEUA6amhDOjI9xted3Bu4xqAf2Iu/f5VGNQob6B9
fg73ZatTbFgXSIrwTEpZ+EMh6c/+8HzJB3bDJbhA3RNP10ANhcLtJ0EzF+lgU2LN
UtqzRtz4DzHOLnw87reeo6X+qkvl2exqGtBwKMZm3/5SSiHs+9ULYGZpWGOxi6Wu
EMbqbirbeU8SWL7k/+bX4rsQk57RUGDegRaQXg5tFBe3lCNuTVeZdTvCJWM8X5/N
eHAVuYmOxxU9EbsdZYRjJGf8JaleJujBH+joDxI19DiV6Fm59XGL7S9GbesfWXem
YlkZCoq6oOZ7aE9khvmW+Vd2nGWW0XqoQHTltEXmIqR/YubMKYTY3XuQOj8AFMD4
G+pKOsjvIX7vGbJn8TbhHCyelfVkNNbRj/0y2DcEkT/oQ79DrgZq768pnMuLK6dP
tv+pcoLESnOCYGmr61bmu3DBpCtoy3A9NbEM1ICHdEXkyMHqatfUlc0QIdzua/kX
ECAkiet1GZQiS38YmVrzNDy8jCO3ypyJD6z1LXtRbWOdiQ8ID0JfmrLFkd0VeGrk
XQMYFxC4yWKuJ6kiXbDKubFj25m7bOQRWEbE6bK2Pt5xReUmFrVQrfwmW3cvM3Sg
Sx+lY8ronjY+rqsyowTnLvnt3kna2u7ScrwR6nZEWULVgBuuem7sZCKxBT7NqenP
3WTqicXzoSW6BZRIjY+DMVO9xiGKonVBg205myWklQ95yXgmi6GHzf60TJi7PWjw
z01tuFoJwx1MumXhnHeYp73n3QydxZh6glrL+kMKt+BKOOA9kENihMPDE1A9Uh5n
G2Y4776MS58gvSfPbe9JNSoGdD7DEY873qLAhvsdF4/HXzYLCOm2NE57IdyRKjSG
Wd0+jhS7WRqHrAmcsxxaPnVyorpKCzipd+EhvH5onlUMYvv43LTeX9eqgagBbuRw
EWF6zKagg5zs6RpVhYzxN2762TbTqMhzhT0R0wkhMYGr8liQoxozOafXNthuoDFL
BsRj204/H9sh7m4hMwmzljbCnCptjOJrBn05rGtajCSCo8tx/NHQWEMq87RJJpec
SF+CAHLiRh6onN51Pe1WKWwEJba5nhazy+qPz+AkYnjBn0VE8L+B0kW7PdWenGa0
YraVaD9btv1DLI57NYgo/B6IxD4qKBijDx3hqWVhaHG7nB2HiH49SGRJanB5hktA
jNT86lb6F1uqxAZ2NVjVfKIno5PJhaZv7OficGwk1UuYSfjjhF7YdYIWY+usDVEf
E/7y6jNbrjbjSZuJgUTKQuR0EkTDDmppogbVpLxl5xoy506tO/JvT9viaBrlI7K4
j49/ac76MGhFXE1NtqbeilHt+1ZzgCsWevK3GSBmV9ol5JXg1YbKhsMcpgFHu03n
pjjWxRDAuCwqBmuG7/FCpLggLYXdZMzoKVamLt01apTP2zFzegKrRXdJJ/kCkjLO
zPxxFBeMGoQUMcyH0+fEmjdtPQTeP41OpUCQRwdHdou+FN7TsMf/wC/Krq3GiJzl
kN6htc9kEzfAh8pAsA32jrmLKwouGAxeDtybKsE3dNr0juf/qbnqcioHtggdCGyL
aPLuIQjfE44le3V+polb0Nny4mjhHYBdrk3BYSsxCgeb+sKk4dOjGFAk2P113RCC
I0Ah+xuWouUyPzEpNGY8DSQuXo7ZulZDIG8ngHOyGiCjucN5C6Wxn05ovfwWBav/
LEN6nJxXSHodOB7oC6k8+HZdnogJii92ua87vNlvtpwO/gdLj8H8ooX93vNc2HNc
scl3ZVBGVP76LY5H/5G3wkuh6pnI/7XI037OuKEjsCL6zfzB/s+Jjt1ymTaCfEvY
+8wOwAYtz7OtfjIuxHJhWpy4CWWreYK4qWer+Q/SEhXqwBIuVp2WKGQce9cqZUTd
Q4uRaIAJZ2TygIkfV1GUT/Z8YQyUjEfQNdWJNodKAs09Vx5/ct404mV8hetDYwnB
l25tldbIsaQK3nhdWUr75RxYVy4jwl692TOiTd0kEqTYxEcxACht5gKAMGz91IGz
88wxRhXlIl2ilLwNRgzS0E+6sJ3U2dhwfZ1wwQykZ2RvrkKnVBzDee6NeSVGWuHu
Fmp/50Ewuzn/52e/XMuJJyBXh8Ddvb8Nr7TZIVzsqM8RyIGueXIphpR9Jw7RsP3s
ORpXWYrZgxCVwUDJB7zIPeFcj5brqXJS9R3qOxiLiTeA2ZaeSdIi9hZb4vJR0624
Vkn+h4fDclIrStZaqhRP5PggzhTcLRVrhR+MyLxTrUnuWXmSRsuK5M4UNUfFRuKw
w352Ai8WFAv4PH4ZaR3AxM0BqmNeJjibo82TIu6/8GR0lv67sKCFMvFku6k+ouFN
W3gQd3khTsRrNVdgqmrF4SvJXXUSHeJuwz1F9+qSdiTKHdjXjFmG6PveBkqODO4n
W+YsfxNLVen0xk0RFvhw+JlT7HBvR6hGHI91AYj4i9BjYcOLsQK50zUVaDJq8lkt
InXiAB1oDnRitEW0aW7YxI2MdzYY5485HbkSZC3b4TL8CkRjOb60L+Sce1U+ngOC
Ej9tm3N7Ww2iDaQMtn606aQVcpesTP3mibEY1XTwEs4s1VIovcG30z8198eu3EAW
NaacHy9hiVrNMBd1grGTryEvIQu/Ct5kviLEoFCZrN20w2We0pUGyxeQeqrNaNZl
C3JCn4whpLE117WBJ3I/6Jgu51StDAouF8dDHLK2A01HXN3kuZr13MrMjJ6c777E
5s1Qa4+Z6Rbw8ioVZrugBjztHHPbucGQg/0LXnfiCfpXPB1I+N6QmCvyG0bNTf1U
eCcvIO6fx6qWOM1O8JD5GeJdN9fbdS19tZ2EDej9AbhwXLQst3I/uD9MkypkNhmE
Naa6d9/3ZT6MK9JWYuyUEMI9bHEWvcS9j+/MEzsF/xwJurmKin4ZErmjoJe5lWna
NkxoRhNia6O7bb5XbAFp54QIUQC5M8LDPirxYFAj3YSg0s9CtYh2GMRTgBdyoN7s
kW91hi0dNg47lKaHwU96qhQeQbBITXDM6JLYMSw3uJp45KPFH/mAehKqTCEswzkH
EWGLXFujT16t6BDIa/w86mHCh2hqwZoWIV3I6NUahWaeOs0VXeAXv8YFjpy+bkWP
nf1h4/fIM/CcxINUEOY3yXKxi9Rpx4SGfNYwj8RmEYi8VD7hrewW5RiQ49njiXFA
0G+BTeiI1J7k28NwBq1jj34m8SoCqgorgfcBIdoZPnp0rT3ax94ZZbLhKF0c0FaC
ryXK08wFxgs0d2BB4mXxzQCy+k95LgdwHEJcp2QwJaUY3ENg3N6MVYrWJvvWCwQ9
wKembKeuthJySm0FC+/5iMU0dKn+WBollRm5PLHjvCnih36a+3QTW4ThGAMX6o42
NdwZJ/9Jn/XOUjSPVtaIotfyDe5BAjvhFFxbLBgfc0S89qoYfUUbcwoFc4dc1YaO
Oz5NwAAC9rNkeqm5AKmR6EV1OMZmES0IkJ8V3WwFkUVYOUGX9zEEJ0f+niBrcVwE
STqlGv0fJae3djwqyW1WU3GtFrLj71BOnjbUQMvzQqN3DN5htQwdbw2nU4DBIwWl
lc807lXrGv11HdoAnPI3J50mXl3IYDKPzZjp9gS8gcGFe3QC98lDnSGV1966GKPA
qK1Go5RtsqhdS1vu/JXnPEDwCOtzkqdqLrw4gNOkWDpBjSPu9CQmCnTMlryhHfIY
d5cEThcSokfe3OBU5iHe4D6ayAu+Y2Xy4Z6rakP7RQoOvkQil1+uQ7Hl9Uqe9pbA
jZYPefzw/DtFwMq7aNqrpDSjTUrYsj9V/7HMAbSqoI6ojQcdcPNdg9DNspNo561t
C5nLMBXSWFxFU7ZaO3nbxIWgCJEF7H+4or15NIwiSLS5t0o+cjIUoKTvTITiD9V4
CaZmz+9rbiTTO6hwMJ2We3DWKaltCpoFbajyGttqfQEpYWJOBD6TVXxTtwRSHwO5
J1x8vw6JPWwHOJQ2VoBkly8fzX2ef11gHqy/ndolhIPK+SxXSOhwJ9ja56ef1rA9
Fiy3p8mUC8I24sy9xo4PcPDFUaoHpUd9d3bnc67pSppzl9li0oW0QoZHW0gWOSMR
Nqs91x3lOdOuE4owHzTHzSENIrUk0jNVII1fQYKhp1OCJfUQnnrjWIUZiX0IuP0d
5SVQMcEtTp4t/wsS3PQ0ZyZ4756nM9jdIPNo71PTxa1Ymt9EYHIJY8dgMWA0CjTD
8HUMUOteKP2n0ISHRiGFozSTqYtQOauKcBuYC9/rupi9lcQkclk/NPTTjOXoxh1B
t14sv07BKYblxMoIFlp53xNic+ejyekBGJSq3RgG9xdEsxwFMtvRnV20t2NYWw3m
VeW/sfXV/ZLZ1pUwtdUHMntSEMZHSeF1WzcqhfDMrtXxUgVX6wo+oarl6tntbBAj
irAf64WAT5j3qIuMHl1CPogoqotUePy0mnJTDkeQONElLXSDHPIZiqyp1jJzrQZv
uHnKnCuRnCxUhJA7H0vlxYhEd6d23VEeCpv9cXv+pRnVj95Xk5Qxne+BT1IuiGJx
4Ec7fRGifQ+M/zXNLiabbDAMj3DXmocDbDT/SMyWhnVn7qvLrIj/OYcOW0Cr/BA2
uH5lqfbEtWvKIqtfbAFBLlSdDHjRZcaEtPMa0lTY1x0nDnSGOJUyQzjYGtvYLNoP
h/jwlrmFv67La3rIAezDaMdFsZ7lYYA/KK3sAO1iI7i97YvvB7Qjtv67NqSvwCoS
X5VWPQ5pAiK5HBKXuEYFHmlM4IqI/nUOvn+A8tEf/X7TRGENbRZC7jIyk3xYoTgY
2Af6Yw04n9pKy5yqIF3C+llDys/+eXLEFh6Hz6W6f9WpNXOqktZFcx0DU2bjIyME
msS5kH5V22YygFA0efAfo4KkiCRb+no+ozN7u8unJ5a5PxG7ljQVOkqD0XRJyuAq
HIfHXm9EkdniJ4h4guK1wRpu8FHcXL2ktHrs8dg/utxRnHdHGO8O0Wx1Rhzysbz+
m+CHwuUoEd/PAxpxpUxLBzjRmVMa6CWC7D9rTfrxpMCfViKnsnhnbOkw7VntNU8G
MGJ381QkYdGuEACXJ8DSoTm6Q7LewB0sxTY3gHnAEGq7SfgBehZwd6agSeHHGAoG
1gawH6RYz4zX91OWdtOdyqOF1ChTazYUggdJHR0v7B+ftqRMTZt2MeWBOyPIkAbJ
YgcWHeUqtt3Ru1J+vbvazjoKNgJ7Y5sXw47EC2nRi/h6WjjwR8+T+fbs3nHYSUi3
VucS6Grnya4lTj/aQdxeaQWd8HAXUpispWUeTLEmXHb3WEuXYIVokMi12YOoADM7
HNSVrsJHq+0OSy/bf9zjAlvlb3mbsd2fmblfE7/KyLK5YF3/4rUUIGCY6pOY7y7d
nFWY0xOSLuCp/7gXLg1bx3EXQsGXuhoA/LmXR8efL4gL4KQZaGs0/GAxa5AzD+NC
BmxJs0x2t8d+Dodm9g6Mva3AJ8LU9knB9x4MLC2FhveimQoF41VrTS6Tc0IbSWpY
nly1ZZf0r9cAymrzmdg5niLsLTxQcOqyaj/Ugj2DOAxLKwqH3FKafrcwi4c3ZkDx
MZbp6bJ6u6VQZjXYf28os9q5xc4vCldu5pRBCdZzPJF18iROHB13+YmBk2u51SFR
lRH8A4V5bxczyylr7XNM5jxa1mwKVW7e6q6FHwA9kzcIitrhQ/JaW/OyEQ6Xk9AR
QDn4u+g/1MfkL9Yg2klRKBqYz0LkxhPN7wOdfRxhlS/HhRtGr6B6cKngKivfr35l
9v5wUsQPyRHYewe3SiNF1+Ewt8m93fsATW795VkvaKrWYQLBeeaVR5aoD8wfY+nN
1JxUnMCks+na9YiJnsMss/XD7+J61QPT1mm2JHW+xxbiOdCpDVpUhqt9asnqvRk8
eY6yJ4xPyOI7g73bjpxcOO5E57fmKi3Gpr/M/zAxhyQ9LefiCX0qnjK/Cf8+vuAo
T96DornX0d4RxkXrw2rQDdiuexo5I4Vkk6X1akirPUWaHoDQaLx98gM44iIXz0yt
ml/MnkTekS1jFd2l0YZAWjKg70Ty48BdAXUo9Ny6rf+NfecUtqicFGhQQK19V6OF
T24b+g/SGX+9DO62XXjq5ESSBDHmEbFxqFz1D6sZPHKrEb8Qc37sj+IiJSKIZzPk
Nb2DdgwLNzkDTLq2W6R2ssNev1vpxeLlgWVdG5BG7qIUNDMr4lJ0MOau5eTxXlIP
YfnxHWMhlj0zmABqs+UDNmMQm5OGSwjxoa1Qv7fXE1dMyzG6su5Nh7bYuQPb0jSq
wMg/anDrgF1xMgG1Kkm42CSgONgiNUm0CKqk+Aw+U6MfDhn7tM4aXdxTR5abYTgf
YtrDNJbWFyBs2EgKvmBipcrCvYzed8bdBDLal9hy5IMakxaeMO5yr0EbYTm+HBQm
gbAwrftW91cA6infkS6BdaMUTi8gTwgMuDMlMBWpzic28mbcYPTFLkPn/K1OhaDL
MqkV5fAU1jp5nChuqalJj7GeJeTOfJEvG1Nt3YtK7XdIwNbSW/fQd6j89KuDPsbu
CG6OvPJ+o8aCth2haM/mI5GteyfL5vvLC/Hho50ac7Wp9/5UN31O/pQKq611gm3V
SUwJtXqtSDq4Y5Xz0i6i0WMTZOcnXs8K1OL+JI4XmjQ5DS565OXP1pqVF6M3OhKM
4aLIA6xzGZBDSlWKt9/FCz2HJ6VsoXtiC7Fb2B6m0yk2L5BS7+krRQkq5ybjI+sI
0JFeAdZyHfk4pAtWdJj5Clhku+xqcy1vRYDaB4iXmnbC2oIXtnzcB3kH6avFaovO
MitWAho3/3Q32/RrllGXO1Bfdb3MBqw7hQtCVFbsb1U+yFBfqRayyzqV+Uwp7VKd
S474Jx289HT9VxvsufXmXHe4VMe8JlwjYjPdRx1USlgCUNNFicKLScxhEhD32XOq
I2fyhv2hiHJs4mRnmDazPnlhOLDVqM14+HsscMN6JF0nIEqA1TBBoQ97RsRmooqS
zbCJH4VCAysvAr8Q3Iey6zXy8aV26TG020pLr9ZxvdiPcXQe4QGHlhE41Uh8Lyst
yMyg2GFodmamDbiLS3tQgZlxblJYQ6gfy+AJXgkw0T5hXntTQqYkI+9W4AZWLGZk
grpPfDs8qV6eXlzHz/UJ7bkXBU9ukCyCgrx8YBNxDjS1CIu2yWqp2HEcSNUc8H4U
zkvLQJV6da/2A/4MM8/90fMrzYG0ugnwhpN2BbxexwiBMSBH9PKX54cTZlrUhvtk
OhMJEIt6jOH6TZJgvPwiNq6iVafRO2f2IDMQtP8KWobHe2ly9w/KdOC/LPxerZvM
JIxR6yxJ+8qDGvRoMiYICGyKPu5wDeb3xkyHb/V+Sc3qWCfUiyIyH2CGWA02vy6g
k0zI+BawVQYnYQz9mmf4idYI68zfixDh2BrqfdGxnwFAPjVo95CxcwFxozts0WdT
tb2kCXks28LML6xv1CdHd07+cofCg4llLnPe7xX7g6kpYuD4vFKd9sLf6T8WYkom
Cqm4+HSyxHbwJ1QR/QwMld23CRBIkmvoNQ6IdUqVUE4ByzXNoifU3bHYsU9Fn8h0
KVZYK4hM1SN6xwAECZYoYYhIQL8wbfSVpMOoRdN6NeR5avMnq24nPx+hp4QF1SU7
XRqM2C2x1Ex9vAeHCn72CQQRfZppBs7AkFOGtRkQom0BzSTzWKHUr67FVDW5pD54
QQE/ooDKAuWDhBQSMdgitgpHchQaZWAavJb2UluZesjscMMCzQKgvex+OG61dBUJ
24KqFmDTEHMff6CnwOVQN7CPEJLTMBGjdDhDiqWYw7jY+qYp5iiXLiSxro/6wu5v
BN5VJH5Xfz2TN+OUrxtiuN7prhTpbGxG2cjkr+FLGvHoR4zXN57OwKA9c7aqyIyV
1v4I+5gXizbNWcfzwh7adI4lun/Yb4d9seaCPXmRxSB6LS2hjBNQAdo0+Obaao1f
wcXzbIhMR8JqkLGh00TXLBnc5yzv179Iv7CZFn/mvEKOsnovmuVvipGU+HWZxL5X
1+AvKV3eC18lGQ8KajLXUacUbI5UCDD4qbQ5RR+EJp8c8dDDVqoBt7om2yhtNUMZ
HPXKr1LaK1j7FEUgF5qehEeSU3dvSoo2C3OusC858v1l6EK+qmrh2jL4ubnEKeQh
JbQa9Dv6BPJGiyGEXzTFBj0zrZIDy6qjrLeWNzWS1GGtvEiNO5/DkDmn/pCkt7M4
3cFzSB2v8FaRUH+SPxUo8Y7tPgm8FXl9QwV0iDHZEQ3vh1qLN5DYdNhUd8vOdJO8
lR0VM0a0zlcgY3fuHZBvnlXqExt3XKrI/zIsmoynkSg3VdKMud9kjhPINMEM8kzh
o6S60HiwvYAmwQYmvpaiEORw078IBy3/M65SgpflIdzkSOG4FOfT+xoqEfBk4e0B
kFuV/vyGchKkPvvA5vsGKfCVZe0LjcXc8ONM+Q1zL9EVtZZVQNZ/rSeQsmYQJ5Sr
hcG0dYvo3y50y37LSPmoTMNeZ0HaGoG77KCdr9+mV6wd7NPWu4JI04MtzZ43VTMO
wSLPt0TnhPnTDNBeqqZxSbOvcu4KOw11fRBlc9GxtxbDbmBbxsWdut/3bD3wZfNZ
vDhH+aTzqSi7o22QHmfzDg==
`protect END_PROTECTED
