`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuE7G3YjtZH/imQ/B0LigSq4Codrm2kOCdnBpYUnpBmBsWewDOlJwZVJMp+aAffR
+oJpVWCe5eVwRrWAL7t6tCudlfA5BbIPaFDQ4RtDsDorB5YpPh37afV0NFWIFELI
TMwyo0WI2gkvGCj/JqjtCRXFzhwCQjJJfWweCPdiXHTkj3MpQpdB5ztK/Aa9wCDC
1okZQYjdQGEUWtH/n4c7X5Cc8bZmPA4VF5er1RLOWOQvjtDiOrGrKVozPY+SgJMH
GhQfdtKFtBYLP5K97aA/4ihr1Ko62j6/EgBobLGdCjd57c+rZIXqaxehfEtGq5rD
QAV6lscfI51xtgWvXIDg81+PhZwLvDLPNfFqOhfI63iRHEQSJkfUdMxV9CG68ZHK
b3BWqmM/Jy8xZzXC8g4HUReqGuK6xCc9CQYUm1vyuPpKVNMYZO6k0jJQadH74dAb
wh8lfeL2ieQk7YD7gkmAQaKEs+jWpAXxhW5MlmqxFGyHxBFVc3AZ/QG/i13PvG39
pYpayC9UG+WgsxeFkL3QhhNSB0+FKIlxq8CFi7KUJTOXvQBbbQORsFnAVE4bQFag
r3FERE6lJ7VFwwR8i0KLH9n9FLphic93WkvDUOBion9u6DGQSFzr5iTqw4gy+2r2
Gme2jZRCm8cHwFhFnJovxmFzEM6Le0HQ0x+0aRjXs5Z0bD0zI/I7EvAZMF7qR67f
/fLk3az96cxfC7yiRGXTFOUNcJu21ORqdYFNf4YyDh9KA+ZMMuzkU9tQSsnIc7Nl
gpW5YcZovxh1wTsP3SgvPmJOZrh7mUdfSdRF/psek80q8Aj17G3y+4rIGWnWHYHq
hsrQ0CGoD6qTWWJhnXwC2EkDS/8xSaGMpcif6Qyw1o4hN/IVQMTmgBTKcIwd3HIq
LkrWPGYmbum6Eh5Nkb3aRGgvSTSTR/lCLG4iKjxu36qvX9C/Dv6ppI86L86Mt4iA
xBno1L4gdSg20RUqsnC44ENIWH5SGtGlQED2aR974hrdL3Z41YON4jIolbSPct4w
+E+d00WU8sRnCh9zaKq+Ol0BXx/ssR+5B40NVgL2BzXUmDn/6GYy+GDyP9ZqE5e/
4M/tzWQgGlgk33wDUVSj3hRjMDRH3hyMaE2SVDyXYvUZ9jTv/r2Kd04Rr0TgThUV
x1mAPXaGoJ8RgWRdbFP70tho+ozjLzTbjMX0QGoQ5VnoXLN1OW4oF6K0f7rpdhD6
XRfOwOwRteKMouuqa8q593I7m5oVkpPOxPU0mazDbxHW7SueKRGHpa+IHC606T75
2dpXlbrbrrHXdSJnx1zVA83x471HuVaJnvuWW5VGXzWp1zjL/58mM0IMa9LiW7JV
AJzvQnx6KuyhK18sSs+6AP6Eg6qX0zNfZPwW0mJOCKcpizOXdCEy3mNGe+zT5joC
VJg7+YRIzsL2kwztubUMp+NtiObNgFMPAwJuBusi9CMaD5TPMTjxjJV6lEjgocEs
lXrxb7lzVmbGqvgvI/5p9bRv4BvDquUOLVNKIMc2oWvZQBGTC2sLvOvZUR/eZARi
onc65z/VyshRjAvda81L1uzAdyYRLluLoEgSEp4OVEEL0g8f5USV1ioOuH/+S0XO
7I926/RiUVr2PZywxXOYDIheZpn97mAD/IC5/A3YRH3M+Jec7rUmvDXZnrknWEvz
kSp6UOw/D09PP2k4gSLsLU/GpvD4AvlOniblHSJqpBVUiwDA4CXYeh8LMwe6dLNw
cJrHxOpbyULQQI/hpHi2dUhtyE9yaYtOJMZBFEk+NRg23uZtUtii4sl0zht3N/HZ
VdyHaggiZRuEZ5bnLfnsBq5vLb3J99cLj4OsHpZHgswVJNT27VN2WK7pADRjdrcJ
mpO8DPAUgZ0TKyXuyy/7WS13vHDh+UhlPI2KrwNfMDO9AkRgrOamnYURM/u1lPms
VdcXsoah6zGkzqN8CAdAr8++JqRZGJFw3gE4Nsdwt8Qkfz3cibgDkqlsh88yXiE6
LQTQPNzxRik3CKg9fKFAKSBT2oQ8cLTqnAXZHlTQEphZvLDBDNGRvx2tiwxt9y1u
H42XQssIG0ycNKor3UXK1tJ3hrR3+GTJOBz6AsI9gqHviktL64ul/Fy4YqcxIFxW
enwWXiaeyPIWJanMD/s3bCkkxT8GCnHWhxhbrHPoWYd43wu1Hh2SnlBQFx4WVuSP
jL7oZ6Ht91vOVqnVy5vRaoAVzr5BCwKf2/wnXJThj0wlHjogQHD+U5LmRa1srk7R
QK9u4hn7feOYTZJlrtFmKmd+0emTCn/42oY8zLlVqruwTEYc0QupHoTJnQhaEH3+
R/Bbtv9CeRkbAZ+2PlYLIzeZ5BT7MViFS5UGWfK2d0M7yPGt1LvBQqpMe53mkF3d
CPkx/R9uXk30a4sJPy7vqEqFjm2RfzUigoLS0JQq3UHZR98sjkW4cINjNHLN7xsU
XzFY8683FagwOpU0PlyzyK5Y2eBhD65v654N8JeCGqNWYN5BXH/vfg64JwtlvAIs
AAqQbs0i0NyFOpScfmrYKMLTX+pxRyexZqU83wQXE7SFQ1xplnhLTSR6aX+Be6nB
UjQPEeIKhyvy60Ywa6fLF8wwn2sPX6OT67OcxDMGYEwZG4XrBwdzJykvv1nNVBKB
C7Xmn1ViSCFRuKn+Kc74NxnwpgrZ+y6e9kdHkgi1CocIGRhwFY8jSN0kZbNhpkIQ
WMxDDmmWPTnsO4I1QlFuYZeTiEBi33ZZuNJs35I6ZlumonLAtFjiAhm6oRM5gg+Y
oU4sRtqg4dBi2VTiMIW54jDXX55ygzLWU2yMoaM6OVqpz0umIjWqXioh7NdzSjJM
H36UC5gTBFTfdNJUIPAZLiM2lINL/Gob4KsC/0nPw0kZWeJUUSTKVxUh6QvreGEF
8UdQa+nUcCW1p1UCI3OonrKrdnC13C+Ho4ERdMm89vYl0k3PoEOiurW7ANYGcSY5
cLtuJWunXa+Rig444a6TXkVKJSAMXwuGjyEm2UvAZzGMwpATHUG5gXB8VWyZ1snU
zJwuRWW+Y+txrq7lE/WlaebbUuE5ooh6qq7Kn/8XaAwRY3uoV7urSaaZ7u9aNQ/s
DxarTGUR3un5HabQLLeDx0OqM6SUFxMrySIvJgKTzQR0Yqk4qBCzBgnuS3b2X+c/
Iiu4cTAxqg3HXHyqdCuJZO7Kh1iF5AGDrcdU7LNfRRhtp+YaZfBOUSZhBMhounhb
wpYmDqcXrC8kyI/9bpzCnJuDVm35DR7MdlT+vku2ekFNIRSmNDxJZTpSB6dywj00
KOek2pLOmbYvDkKaZd/i2qWayWJpYIH4XrDYxZjlvRAhQrA2UaZGyg3pLTUnZkZD
3UWNUEpXv58fqtGtZMdPPVDKPEvMvmu8440fTr4z/X20Mli+SlTsAfMJnvNL6eNj
9tb5gsALgx874jXBb5EgcEi33hc1KW133zOSoQoUeeU9mK3kUlk721FXuQuKu1oz
AKkrOZnOL5+vF7SMo9ASTyzEDS0Q7TtGq+sLICmqjJANK/+W8qzJi7FHs9Y/b4Bd
4o0Z4/9ijGy8INWlTQiimSV31rbaZjS8iCW8W6j69mSIyw8dFk8KiGxzHMl+QDvm
blu4dew2LzgK+Brv+jAre8MEwpjnTNu1UTF98OBHb9BYHGJYJjBserrRddVXOX6B
Y4jFmAYG4vVEds1YsyZUY6Lii0W6l46Qt2k21ZYqarVo6FZyoRvyucCliiHL272t
it9idksZHyRxeEO8SsdLf1Sn81OkIpuuTLQtusboed0LhcT2Cq1YtMcGseaZXQyg
y4TfqzClYRjvR2p8jCHa+5MNV7m0D5O+ysJRKeEbSIG8FTc4KeFO0GaWP7fU49WD
Q/fSQKCUdeF+VpYXzVZUYX9xZTxUQ7bzWQ2FXVIhvb4EgA/91LsLF1hlbfoI/LDA
O4xfyKgVKj8793q8rgXvYA1soFXVrUcH/PX0C2344gZ3XdRvSRDz1pSY95hMTxIw
nTFXWhDl1K3F//lVnnYdwZBvTA9Lm0jSh2e5eJAL0BQgyXNwSOuT54R9uaUN5cNy
1wJMBqIhLob84+3XVQ8P+JCTSZf+DAKwMRuQAma81kAxSdjzHSIXpcdAkGPwNV7Q
dP44akLHR5e33i1JvxesnLeqoVyuA5wGoihw2mn4SpVtKv8HsETWHIuq/5e3vi3d
`protect END_PROTECTED
