`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jN/pq9nrerp4qlIVkItWanNrYUt1SlMy4nN3jV9gCfX/ztXAKgWiDlDtRb/uSTzK
TnjF3xazYB8uzu4HMv8+fxWJ1MyMkqGDYkmWXieE9+M4Xo6z8OYrTeAkdHdlVlp5
cTlxsDxkf08/R0MbfQu38n3ND2bbIpqWwYYqZbhUJ02ZLmZNBnAdJsphHUUt7qU+
uEdyn2khrPO3eI0G6O7GcafuA4Q1uq/MflvcG5NqC9iaDR8IU+KOzrSlN31s4hgs
cAHrjyDqyD94HWkRFJjnB8uAKX0ioW0kOdqQBrXqrNqDlow8FZHgs90JMPxVAv63
pS+Umoae1OdtTh4ybg4SScDKW1C4kGD7g00c2zuC4ugntufsOYvHCaJXhJpike50
8m93Er9gvqSUV8DBwkvS/Pubz2gYi0BvokJIu532iwi0LB8DFj6epf82PnSvY/l3
pypZVrQofFLuMdPkRcgDc7Bzu/Qc+Aw/ZyPFHZDFmO4=
`protect END_PROTECTED
