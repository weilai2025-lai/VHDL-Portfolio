`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sey4kEHQTCQoa5rUfpQRs3VBYfig+6JFbd7griTimx7mUJaHXIrIfF6cLRwGDguA
G2xPrV7nhnEVqS4vMtDg8OyGIWPneGMD4fk/FD/2qQmN0dN53+4bp/z6F2B+2EZN
SuvT4mFBLRlIVm3gFkzDXiW8Eje3VFxJwMFoDETeoxlxvIslp3dEE+XoI53H4SgR
lUJvbTYzlCjcqSNtLxkPcSdlC5OVx1pxB/kvZnm5+bcqQVYgOIIxiZ8vMZojYW28
f1H7lGeVmzoxnWu6/8zeQnzTQy3Ydp/v3Q1RO5y+AM3zRBC00U8qSTDnFLPNhSMQ
C0y2ZZ8sdsIpbdYm4n3ZKOjyAm5nKiACC7Bv4K8kzOI=
`protect END_PROTECTED
