`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HoOoMSABEcFx3ySCRecQUb4TLWnbUM96wl15f5RaddXVyxA7LLNZqi6jsaU93G7z
em2j0Bi9L5CuuURbFRNAx8EMBsvw2Ro69pdlRRmIZ2Go01Gs5tYgO3jjCpF0TXdg
TYZjul+36okfiLeeSz5srKKYEZtxEAKqkZNnLE+a2EXqySPzYxn9jfR/IpfgF3sl
0FXhK38jEeKi95i7zeVUAdujhe4vli2F9ZDxXISHF4jirgljIQRKRjBKEw3mAJzF
TAHswp8GJQiijaSJIkRhSOKQ6c6SfjFxuOWVIfy7MiIfwXyyvGUy8ipEoF7LW8TI
+zavxCQAHitPpEnbllDDmvWV7assL92vAHl9vlLRcozF8lxHCIP9JOemn7454r2r
rRZ7jDw7+gZ7NkjkLyHPS3wAPRYGeHOy3Sn4zOTNy0ljyo+kOjoxIUxgMOGlGW6y
kdXgItOfskI5fJnNTwrjO+GG3ETt24AHkk36nai1kbJWq84QtY7KHliEPif+jG+2
x+uZ3nrLHlHcXn8JZ+3GATf7GhJbiKRE5ygxB4vmbRlEGH6j4Vs+eedBicaSEfDI
edbTJx/UJRpEv52Bot8oSUxjZinWuk6W9moy2XlgEmatDbwotXjHwRjJtcVP6T9J
8IY7AoMsoanaqL7ev47aN1+itpOBq/c5v/Cd5H/d/OdtGPrwF1lrl2nmak3gPhNi
QCrkXppYwf7sd4CO4wDwwJLxFvmOCOGVRtU4Q+UfA/QPt0264pVb/x0iZSU1hnn8
vbson5bRWfvEIxAonwsd2DhuCbz0q1jurOvWVxArYLSmg3Os4mqoS15aP7zJm2Rb
qdxvx+cCbPnse1pDFbjmjpC8VUtm/32XrWt1FnAwxmyeucBO2ILKnsY5M78uzRum
Km+08H5v/iovIsSh4kTg9RTDu02eitHO+78XBuKIi4ulcsHcwcAB65J2UWcbUWdN
aKdNNitkItBc5tTX+eWmjE+tc1cMgnJW0s300yy1Xn2918WtJTzM2jwYY8LCmujs
TQ6p/BHI9Uat3eOC7wLjBSIqi8wcbj0OJ/4K7txXQyRZXfiyoQ28AEC1lAIiee+C
T57IU6LTqhERrEG8x0c2m+KN9ptQMXEzc19Jx6vlNcF0ua/a4bLyj6/02c32ukQ+
1svxp9YUtB6+f5CiTdj6Wll1A7Mj8oKtzbak/4YdJsfJhiBTEXyNFBDz9nOQ0+IY
DZbxq79XjC2bHYnPtVxHmL8lsO9l3tZEWq63pSvIPUv4/NSHEF+a7BeiZx04ipAa
iUbuPU4R2+KyM+eUJy0kbxa0e4IJXv0kpssC2DLojaX0M+YDUMnP2JLMmTfUWpur
gsOurqv/fUpC9eVZBb1Gvd+ev+s1npP6iH4ohTA4L14QiZE0efyShMJjLDh97UB/
U6O8GU+GmfTAr052M14dyX56j63Hygl1C0WjpgNOoPc7L0VLmeNlpTes4gxpb6cw
py2JsLKNO/09whyXsX2vMz6RsjcXCkFEFTF8VyhLwrgiIG4zC4f99YZ8z7tRr1yU
YN7AWJ0+t1OEOemN59e7iLBkL9g7P6u/TEZaXc6vViNPfc+acp/lhnemGHLYSJrJ
o1Y520d1hm0WsecS2zFpxn/I1izVGAmfxjd2UZZWnkTRXH5+u3PSWn3oa4EvsBPq
CAy/6EVAU/b4In4QKGURMDT+J2CmndYEmExqzmtX/gyflWHYOhjHkCi4u/aI0d4T
ZVId7TsbvwblM7jXC0hPFR5bZVrdOqIdF4BKRjfpBHwJvktNaAOBAe+NfGZmntVv
q7EQkc2aaibAHUxWZckulGmOVroR5vJ7vc/xDgYwQeGroDD8LLJK51HLIuHuWHs2
S50yUBglE7zuV8iiNLh/lftBUXBZM2Mxge8VYer1yqVsbTrrTRFro4CU/ntHTwny
gs8/dXqVnZ/5Nsikj6BlLNYDyXb3vzxAIuQGmT+Gz2UPJLjehfDowIwwfP11X/jO
mWt3Q3kkkJRyTGvExr1UjH75RD4Eks+neQeLrPKq32zCUVQttxqOpL/eXimvxgEG
tfTyCE+Lw4nSeUhk3WdBK+r1sFkpIOEvS0uUoyD4VKcHre/m+gUMerspiu1+l1NN
AEe9ucgETOayuiWP0YZnTZkUnYbfR2zqcYlIN0gKJrLlygox5Eisk2C0lL9Z5vil
5wCUVF1vtXp/LfGhG1TSy0aaC3Wx56LxMUW1PIN7QiwPHDW7GV3sQSup/jBq8R9M
Zlc2lZ/B4sE0NvpHdhZbEV3crFTSAhKKV0uVxprr1IA+cpCVHxEAhoBXDE1iBcTe
r9+UmhlrJkStFsesYP4IJ544VcxFfhOjIZiBcaFu9jw7TKh2DyA3f879zSAj8p+7
mK0vRau5Z2FXW3geTQB13jqbDYm2wyMoDJTRnibcIg2qPtgyjyA1cl5X9koGIflz
Kd+EK+KlLhFXoyWwda/6wfodWotaz8F/zcZNx7BpLCdyFl4qOT4X9RW4ZtMPQblB
W0gb1RBte8c/LoJ5DoAi/M42AiX/LLKaJH9SKU3dlGrWvZLuaSZ4ATyAR5IK78wR
k19KgNVhR9u1o5K6O6nd69gJYQQVhJt82y7CMSVb13Azjb2OIlbZIyzlDoJ3xYtl
WM26go0VcLW44VA9qu6OVRSbcgD+cUHldiL4n+goTPAqY9vRPhzxfCUPzka5g9Ya
W5aj//17wQiUvcXrvBhuRnSiXmb+djajqBXzlOx1MFcHDXKzx/FNKnn7die67AM4
SG0tteIVaSXiADvbvrSa4FBm8F6j+yYIqsV2qFw0UNFjJZlHMVQW6xeOQdltRGEt
jjSchtPHV6nE3FBzaOTYcsfdUxeTgjqjmzTUTv6wDIMpja6J3CfMnQO9+kUzt03J
CC5szfFeyn4Y2Jsz4GK1pv/+/KO8yszDphkwTozfpdrol7FAUU9Bs0O0tDhfD737
25Aad2ia7Ht5KjPNsI93qZ5n6NrPu3AmarpTUG69bNC5jl2p8qNBmT+78TxCIo9o
hP09BFuM9Zqj/mB4jAEBqIe8lC+gVUrBSDVg11VQ42AvG4FFzM6ii2YKDO6GUX2A
vilm9tHqd42Kmbpp7L4BYqji6gMK1y79EYPmAfC1rH1tNbIG0d8gBB8+AS50YQUR
IlyNK5twCp81m9RM46dQIh71wZFST+9RlPeCuS7VyDUjU0tW5xe6dOhRP5B+snEC
Rwhy8CRVYClMdDAHkm6m9xF85+OuKqxWHtRh1UHGDwDfBCetVBz6uTm0kd9McWU/
BL3oCEPLXDrUmkmPnr0Ia4YQQ7JsAJdkvVDLybuthKI2E4XQH7bjXHFYDlNWVLF0
6cG76F82D8/S7QqpS8/iipzgwgZ6MS0yp/hvn00NSbYCqGh9Rhn4toVMniyn7eMr
UGvVU/UqVJ8o3ccDQ/kWVVrhraVbZo5CSMmGLURC7wK4xEVf7MTe3HUoK9ADR01w
T2Syjae8K4lxK6LmIjRCXhiieRYZPZ8fPQtF6ck64R7KEP4lRKFOjR/fMSlbACaA
NAAKtrx7Q9FsClTbMNUR1iLj3+LQhJ48TdQb+qpj4nPMB0Q+hJPyA50E/W7cvlpY
kD0jvTI4Bx4U5k7vSTQucjyYJB366sXhW66lrI92DHgW2hQo8Fs4MbT6L+7HMh6+
rKHpJyrV0F5+pj0J83GiVkh0TNTS5w/UmBAZ30qj04a68JOEnVuZ/okBKyYTpNIx
Z7eJLetgCHsyRk5Q3Ho7JkDxrm0mRpmuj1x1jkaQJdCK7PCXR+QOUB5c7YEmiimE
nBNF7KOE49TJztRt/Krz6VBFVHMKDMMVdNFQP4npy3KYF7mWYwPsQKRXGAiWYY8F
Q2Myz7If8jrk2k4rsBLkzdkaNZ0OkGIcBK1ieW03jenYOD+NoA7OvMH6JRlBM5i2
NU+Tp0VbDukBmCxH/9gyml4yfYNxJnlKIfkVGia0hhMlvmSt8p3OFATDR32VDQOW
P0VcEXDBhTXzVclecSv5AVbpA/iQGuAhb4Ppl/v8t32hgpmsxKG0/6+BtsHvhnUF
Aqo1ywiKp/1BqRGBaSV8mOzS+CecxCdhTWhG+vUqdWpbjyKryr9RhQK+HA3ahpLZ
oPz40CYJU1ZokmsORcU2kQc3k+8q9H2Hf0AueXf8Cn7GNIYWsAzWd5tksVJ5/BJU
KQ2mLxWEGSQO5UwOZXUKw1RCA4CkLWuPVEbBy26KFGE2e+FXIJgLYo/JZYFaK3cu
NMJFMXgUMmsL1U5ucdbA7t+uWB6WBX3/11V5JH27/He5RgDuAUSzpD8z4i9Iixdj
jrIPhu6Syd7gBuJlFevRIXU3YuwDCayfyvSxK8k/Jr4FXmIMideNrHoww8v2mdm4
moYf9roHy152pi70gH1KyoRQibUFT8nVBQ3VXTmW+39ZkiWrlIDahnKI9Z+i8rbT
hqYQhAnO0+PKKkPjY7ZWukztO4fhdzhd6FFhEPznSS+Sz9UTS06iVSoak298ydmY
7FnVmnoHIxFR6aW8Al1+UScghXeo2lxXiRyX2O07J58ZQ3vfcB6XqLLIANBeK9TE
lOh8dajyIxO16b4yLNonwdSn+xbih5F7C/vElmReupx27MH5KnCQITxiHnBvt3ap
qNe2mcLcwXQRDkLIgMn3JkrZTPjp568eSqQTZqE24by9fAAShDH5/r8FaQACpU7V
eR5cJcuQFFHAKY0K7GsTiHlArywEUUXz8hU6TNOvBvqrizj6n+49+41e3l9nic8c
peqgwDrpX7ruxqThO5IjbwDZ702f7klR5jHITnd9o3B+4ASO3x8C8r+axDrVQMw5
TvOmKg/P9BHINgXtHxzYH9JOdlxxMKDEVqU5036Wv9vRX/tTdHZAPpq9V48qQ5Ka
IU5kDZ36h8zIxk5bqDG95yzE86K7pGKCKoF7G1VBsL8arjVVtxg5VnHYoEiPMixu
bdwGlmdimf6DHMLI8xwGa+E1YEMvixOyXoUQddb7bR/6CroRc7TpZb7aaavjValn
p/DFi+HPU3scZrJ9MXDhPelkCePiJUGbp68iBtNzUiQtmA89ghQsWQLxNn8mSau1
41G24vPQ50PCb2nVak51ioPB4uGZ3T6bDwnqcHKHonzkLbJO8Q77xKty+0lb55qV
a2NtyxQUlOfKDcj0QyjCBZOPaRcDVByIYpq3FHEsCUbh3Ffujzw9iUSsWi4HpRG7
R7IJRG7x/Pdu3QS6Tje7iuf6/RgVXd0Fjz5RYBUt8N1fC1neEz+6EguJOUFZO1Hl
qqzzM0M0fQ3XD3WaUC3A1P/N1OtBGpGDjZGMTDxIDjzMOHEtM77kUQLIuFf7iYac
9OQbzwEJr8lXE5DfvLHC/Z2U5OCvzff9jqq5gYfANAClr3Xa2p/R1XmuVCAKRZn9
4a+120wbkGyLluDmkLxbdsCXOJ8r85c0nUzgXDSDBqNJFIVaXi7KRpDVewpY0P+g
1a+ipO4VKY81FgaV5g+ia0nwOHtssfGNJmu61B47IOAgth+6Bixjk2BQ/CkZ/M7m
FjHrA26Px3TfvEMGm75EIbbCOTvLcV7m1auUY1iKdwb7Q+Vaue5lFbEatmqgS2Ns
sfLxL3ISPBLi1x8Xa5Z2J91iyEJmtf2Fh6t/sz3PHxCx/9mccQV43f78AJy/FXk+
gBTi3nkGAeeITEjSt+SZiYh9g3qYJogYJJfwPXiMvJHfD1YNchGF9/ftBOwkdHV4
Id5XKZUnbSGUzkfu7M9LcM0wQJM/hQVcRqFZi9FS7FaRscP6wjrr4jCPaBQFvEbF
WSI0V6tvZiEi5IPIiz+Y1knBT963NecyKuXyycEp5Vmqevr9LhvgSP/CBbCFUd0V
Tk3QzAU2+z13ltLsL+0VoDdnEcS2KOEDLmAsnEZHD0fvetp1wUKZ/s/YcCAccjhs
8QnLX5DK6B3SGCrzRcBnjK6OPmR+4bm1ovEL/H+YfSy/vgMPavSWpLngfkIwMNqe
z1+sw0Sk6JcTfaO/QzT012XJq0nWwOjBz9P1ZLiL9QgyumZ+mMe0ZOfqTnu+rYKO
ifZ+xXp+hPpb/+XwNaUaGZjUewAlz+0v57shb/ChUmSzRb9BYgl4nDQtg51MENcp
0WsO0vfHVSSG/QqLJbKHghnjq1wGBZomEsJy6msppS//zIcP0L4ws3aDUi2Vrt8T
QrayLeucWjc4Hz1IEhwt8ErKrYKs56DbOiNDhyCMWpYNSuZLUt1nILOgSVPlfgky
HVGJ16I+sRyNPWUmDgUGBFcDrfz2StP2lixCRb/HWgoO2eAY0n2uan+7dDj311ro
vxkAkxfOyhjYOs40J1F0RYUnbne9jIvALNW77p9ifyQmsKpx1vGI9G4zOmj/Rb6L
UH775Z3nR9wfIqEZ4RqWs3KEY3NiQmCpa9PGAGFxWO/pxfbooTYVIyxO/+n8DA5o
K6m71NkjGp6KH1GjdkJd4I+ChkxlTdeSkRA3O2Usb8QIvNY+KHbUpqI8ZR2eLeGk
p40p/C8kgt7ULDwbdmxLmfQMskOUQV+LBJMe4+nTq8C6cXEd9gYYZPWy65ChJJUS
TbKYK6UshCCCXVbxOt9GvuzFZWYnRNpjcHhTYD1rVzNfTIT/X+Pu7yvnIcleumGm
oNfXeBnQayazLS33uydIY9YucRVmbXW8FIkczNuIIHSevfiIeu4pJ3lp9LVtCB0j
0R1VAlik7sGTaZbLqcOysruEke1ROAA2JGKSlcxad8rSZszFRFIw1cRiGfA3geTd
pVXaeJQIZkHhM5xobAs9m+rGraSMn/fiiGQVdVmCrRESASY/k71aCzSFzBaBlTde
gl4xIbWZjPMeDoZCufzKFGp78Uurw8bAXFUblqx68HdVxvBvZUwiQTXdN9GMnSk1
p1ceMlfmo16biaJtzXBtwXAIiiQHjTsRuG2Qc9Op3tqO9OuNtnPH2k0r4Rth4oAN
YOQWD/KcQJQKogiH0zvBZEPvOS692lPqqf+ijNaZaQsMok4YTQ6qcnxVz5BcKBfR
n3Av6QZcKmmgaCIKVF3Ls8Mymw3os2M6xR2otv/WH0xJBXZj8sqnrVMEgt92K8vB
kFfhOEdqudzv0MYgmFUKeoxdjFf5DPh/o2BxLEUx/WeFIm3OOp6QHf9vu18pIDWA
2iuV+OqeCw69qYEFx5pU3+DscsYq1GGO1cyanyA4r3msZj0VhA2fL8UcZvnbm8ks
Ibn8yZGXs+Wg1S0RwJVgLLHxQMexWEk9ghCMhxIrI/fn38QlWE7g5SAHKBAaETui
vPy2pZ32TDzRuVPjVYIIxzgHWHUcZToGzb7ScSylgQTL7luX7KoS7WFXYOuY/LNe
aeNDFEU+sgG54lOHsHEjVtEN+9YSp0pBj63B221OPlXjoZGuy1e+hmEgwrVZFJ2D
2vwFLB+N4duCgvTlRgbuUuIenUFvPDmzShk70f4EJqbHZcsYvGlacW7TGwEJ4IlQ
JrNB3z5i9iShfAsYiEsdv/lnACisLKusKSr5IOmL9uH6JhXMMd3XpDcJ75uQADz4
R6QkDiyiUcygyRyIAwGjBEcLswmDkpCCbv6adjsLkkT3enao1ta5RaqjP9xyYs1j
aWT4xzn8H5ANhfFeFNp3r4ty/RxCZzY4N05qYXLaGKKuEziFzYTUHNP0cz0qFyrR
PWN56AI/NoZtudEvM05LFPmSnRWjTFyusB9xvzIhmcujXQQ/j7BqJKOxe33FVwln
E1sFdwLjlB4/7eM8DMoGLZfF/e3pJrXTvaVY/lWjAS896Wj4NloYafJTG16yBg4y
a4SXnwmhHXZ/uVdkM/C8EhRvbj+iyCohpGFMJqV74+w81aWPTbe30+7kXwjx9VC+
YkKrdCBHJcLeVR0prghLicf23p/eJE/+GqOeesYSPiqIao4WDvL07FQSwY5APJZM
CQRaKDL3SxYIIjkw3AG/TW+pnxSqGlSnY2DT/FqsCNIMxoXFfGu0Zr7jS7NQmisg
jb1Lyc3urrrNFCS8hlglI53s8/+oh7T6rLyuvX1MewCC5OP3Owwm9QN2Vn5tdKP2
Pho9qSofCA4IO4YxR6SKNHhSpzD1fap6pOZ4Yr61FTUhk8fSIKnK3TxGdAHAMkBu
A6TNdNfmWqJDx0yGZT8S+qwOHMKVcrGlumdo3nTF5HRCvYliVrUBQqG6JOFI9YgL
csno6GRw1fpoAcDsO5s1HNJIBG9l0M1OquK8PFOMmmgYJyLzHs+jrtDI6X1Btt15
hOMt/9LQebF3OPBaK1KLZOoils3qnS6xJR8D0dPCcATg4z+pvchwBYXGKX4096uG
zBC/oRLurcDc7MNby+e5xJejIlkntg1fBfctPu9WGFIjf2sf2iZ9GuxOJulmCFzO
d8Qhc6y7cH+Zt/Nx7boq2l61ccyPmp0AD8r76u4LMgoW97yKUr+omt3giUoJXruy
ArG3jgzv3QkTpWE73NamqmGs4NjJOjOspNADACSJAwgztHl5nIjW+yUBta2m9lxX
/i+KlkqKZTxR1HihdhBgBQXE87qWBeiQKn+I5H46eb/5VAmmaRBETIYzF31J9qOW
unRU8UYNDdbaDJptmbf4gnBGWeN+g/4q8zKA7D1y5VUS5/g3Z2eWwZ+IYcF87UKu
ggP1dL0XUF5l/72l6nywVkB4nG8KZZYrjUAQlCZ47griPZVy9e+6r5C10iNkP9kj
jh3an0dYYunVuPQmw4lJT/vY+ceg3WlfEFXCV/JoEhkCAiL7GXmwRSBq9nqeSXzE
QSmZIbz2gTp9Amz15T3uh7u83BJT1SGT4RZNnQJ5cCxUq5gpb/7wxBab0igp587/
4kVDqdA0qY6UCez4POy3AerXvqv2fFlE8DmK1zNEFVUcxTEWURZeSD9uP408jy3C
nIpcqi9FWTCMMx1L9etLvQ4jSkLcWkjq/xVJHL/fRBqH/S8hcN2ak40IFEvaNPtl
A/oniqwtn4N3XFa1NN95MblhITpq2UVylLTuTN1zqZ5OLB3WfEO4m4RxKqJRLVPO
TEnMUb5o3sP2N7oV6lwgmp22FCKg1JwMiEKzpMlwodi48jIIML1rLDeMspaEbk4u
0GiGod5Xs/v4YQ1U3SCjQj+7Suz76IvT2axt50T9nTFpP0+SW2DDw8ZOAqZSv6E4
bBlE0CT9BZoQYzveqwUSwkYINiX78mzfX9g/Dp8Ks40s/kyyOBzsl3tTfW1fVpMd
v44o4dfnkdey2xQO8ll+z6pDFgrhC/aKvWy1o2gyEEYwdVhKzwAKmQRO87irU5RO
wL37wWU0q4oE0K+LmCUSuyNkJrKTfDBfhJaQvhVum16oD4RVDnvEEeBbaWUp2ReZ
ssStvEw1347cPTuf7WQS/AQRGs4c3plfz+nw9U3jyKpcRBgdc9ELeFOeh0meyv+V
XHynVhS9x5cmd4I8l+PxmDdHd1NQy0qG1cZJtsJ62TG3aHS192c4YEZSvDXahXGF
sLcN+Py5YrdfteUt8jRP5Ubbcej4UIcGM1HbFy32BjITdpanoYlQ0dY0aYMgxXeH
W5t5luMAmcOkTRMeT5EUOH7WxxATaY+SIYiR+w8cWodA/H9xOVsQoBb25u6RJjK1
RmVKu7x0f+cxM12kvJehwSQt9Xo7QE8anby1EurMHkTVV1//EHHvycqeuvAZqug6
VdCCdd9pTst+N6dNXJzFMXtPqrjpIH+6AE0WrZhupDRJL4QQAX9uTbYrw4Kx0hYm
4YaD1XpEUuuc4bpgmWXaAL9s8x1xZoql19GDfMP3Ehr3AQYYJL4oj++V8xt6PptX
ke0iTQCqVVQ0rqbM7x7i+ma/5qC0KZgCXJs1kqpZtVF8ftQSsrqHal4JGNQZHtV3
EIUTP4Fq71/B838fOsVV/K74ywyORxBEzfVbO/gVOsZplu7chdSoqylj0gfAFGjy
2/5f3zCA751TQzyZWAkrRni9LcJcyiY7TOhQG3omjXMnEwlGNWNfROQHjDmhopvz
VExR7ci9lt9pivNfCRej5P0bFTbCBzJXIpO4PBAEPb0qzPQnvGh5n0wo6liFmb4V
gCP4fLj1KmZbFfBxpHjkk+YqRIt8KS+RXFzHkr/rRU174jfqZkI1Wec3P7ySaKBZ
9qLMDCIRTs9zBjStMzASLFzDRS+Pn+kR/7kA+AhzXSqtKNROdpd2VNk4owXTqYMp
7uR1dCVLz9tD1nG9quaD8fzA12Gd9d9pgPQxVq/fwmcNFlM567ebOxtWsIKiBOg2
TlOPaXlyMF/9Q5YF0ytLZpgXvsas+tyI3L6f+u4hmL/7wBAkhoWtAbpfuipXh5A0
WFr1JjFxjnzApV/N64BlzogCdk4nF59gveafR+UifT0DgFLIDWmTTpdXUQ6z93x4
lFhgZBtoGzckfLjzOpmgY0icrh0mlAbgC/xKY94YSj4n/wNR4bpOCusyEaKNoa7x
oTC+Bd5CJw2TFlYnrbG9GrZrrDgE1oLtho4/axhWSOY3QgX7Id+wtILT/vcieWB8
+ei9joBqOLNUrO6au3v4Cj2gXDTfBkA5wXfI3Xzt4ZeKnoif8VkK1pZO22XjlIJQ
t9A8ZRmbAQwo5978Z3WKfWxwkdX+DolwQgf2hrS/3HxtdQd+AGVIGq513NWrpUeU
N8AW7NHSvUHEJsW8h8BJCJNW7BN2IXoKUN7MJeTOGS8ubzV1G93Ge7AsRDFU10Ss
pE5pwnPz//mowcVkLfhgun6yx9nwvliwToI4ERWXb5NWUglXJYbA9Bgpl/Z2OYzZ
1M5uneIe970tCbVB6muRXG2LnG8F8kdwowkwARInNRS/HuqZMRDIT1qdjd4sHB9B
78QI0P3o7CPs9OURL7VZttSlRMCfhtOXQJ9xeiGh8+7/RqaW16QnOmDfzVOD8ZWH
TCJy87xyN/c4qoP4AjzoOlK4cAakbK+29TIf6vHdshjHetVDMWbY1KE0BynE44Rl
SFnxe5Ag1Vg2NXDycXHv5X6hRoauqB8U5zQn+kJ4D10=
`protect END_PROTECTED
