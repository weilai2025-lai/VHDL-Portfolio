`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kaUYbslsx2O6m5HKo0hc/RJEXay7yR1Qzu3qvIAVJKUSeuyh31ozxGKnVGH9MNuj
dMnJHJFc26Bq1LCEvAs8ztWJqWBi+bpFaeVZXu0voOrpioAEBsmjAGVcY29RYGIc
DnLbJ07rPoO48/3lSvpUhPFfLXYMfkv09n393+bXTtANB1ddAoli/G/OKaxo0lM3
F0SObk9d18A5cMjJB3P8NvhH0yOeyJ9oNCD7KwNsJgu6apAhuuza9qMtsaURojmr
ho9Cl+mfPvFYB59bbJBU0T+lpCcD2ANh9XbpsjfsTJPTrerPpw/e12bTlNuZqCxH
Ti0JBFEqXxWN/EaliB3xasPv10EJ35dE/Ho1b6iDkO05gdClQqM3U4y4aLbkIrC6
aDDC+eAn8SIafw0mFu/VXeSuBKmBTUCzH9PErwboRgxDGperKKFQBZXdBGwieDMu
cr9uAtck3NXKZ/VbslGRTrIsVApcnz+L5Vr3XNBe7FLxFlUXs466EiNk5y8yQddZ
axKb9Y+ssVPqs5puhDFlJm6Ns/DQwHXwaQ2SgC3B+LxzB92IoGoAn0vhsdc16+1V
`protect END_PROTECTED
