`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GcgjtnMYvEha2YnN03mFKJB7NoVacTwh6tGzeABOAFdjcMhdRL/mISSZ21MDGtqB
VyILDpbzGsNZHYykEKYVVEpvdnIuVHumwbXz2r2GFtlLT2AsH+SVXVNwNzkJtuFG
VB243zJyMRbWaQGRLw89zjMorMD1DP0E/AvKxmMRQZ0bLiuzLSVgsnKSy5wKP717
`protect END_PROTECTED
