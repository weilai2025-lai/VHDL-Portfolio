`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzIHzZIus711C0GIGylnkT3C+L9XF/yCxs+2xwF0mSNKxHddgQ+NBTOjD2fwFQjY
a2SavL9GZQT/W/cQ1EPPo9E9CfuZNsOgFNEhmizjBtS95nWh94mlElqjZG1JmD3q
1HP5jKp5rN8rt9D4x9ttpOvVcqrM2tHLAuWQJwz9OnUprM4FnDZy3qev3Kix8BJr
xe5I2UJvUHQLMQUJS3rbvlLaVXuvdOiLY2+jN2djOYg/SIExzLmQ4vOlz/4T7kcq
hReU+XbWp9K3wmydnRUNBAm2fcJQWT+X4QCRXlNPDQYCZtHrKEG/yS4yKkCVMq6B
Xiazhn7M5cIbQoG+ZE7kHWDrk/IbJgvsoK+F00Uyi39uVSfmPmqpHETPBcBj99o4
+q+p0dnwzxGdcU8z/U53xw==
`protect END_PROTECTED
