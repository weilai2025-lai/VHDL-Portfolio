library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity fulladd_clg_withsubtraction is
	generic(width: integer:=4;
			  width_gp: integer:=4;
			  width_cmiddle :integer:=3);
	port(M :in std_logic;
		  a :in std_logic_vector(width-1 downto 0);
		  b :in std_logic_vector(width-1 downto 0);
        s :out std_logic_vector(width-1 downto 0);
		  cout :out std_logic;
		  v: out std_logic);
end entity fulladd_clg_withsubtraction;

architecture structure of fulladd_clg_withsubtraction is
	component clg is
	port(cin :in std_logic;
	     g :in std_logic_vector(width_gp-1 downto 0);
		  p :in std_logic_vector(width_gp-1 downto 0);
	     c_middle :out std_logic_vector(width_cmiddle-1 downto 0);
	     cout :out std_logic);
	end component;
	component fulladd is
	port(a :in std_logic;
	     b :in std_logic;
	     cin :in std_logic;
	     g :out std_logic;
	     p :out std_logic;
	     s :out std_logic);
	end component;
	signal g: std_logic_vector(width_gp-1 downto 0);
	signal p: std_logic_vector(width_gp-1 downto 0);
	signal c_middle: std_logic_vector(width_cmiddle-1 downto 0);
	signal norB: std_logic_vector(width-1 downto 0);
	signal cout_s: std_logic;
begin
	generate_norB:
	for i in 0 to (width-1) generate
		norB(i) <= M xor b(i);
	end generate;
	v <= c_middle(2) xor cout_s;
	f0: fulladd
	port map(a=>a(0),b=>norB(0),cin=>M,g=>g(0),p=>p(0),s=>s(0));
	f1: fulladd
	port map(a=>a(1),b=>norB(1),cin=>c_middle(0),g=>g(1),p=>p(1),s=>s(1));
	f2: fulladd
	port map(a=>a(2),b=>norB(2),cin=>c_middle(1),g=>g(2),p=>p(2),s=>s(2));
	f3: fulladd
	port map(a=>a(3),b=>norB(3),cin=>c_middle(2),g=>g(3),p=>p(3),s=>s(3));
	c0: clg
	port map(cin=>M,g=>g,p=>p,c_middle=>c_middle,cout=>cout_s);
	cout <= cout_s;
end architecture structure;