`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpKIYS/VgtusNeHZALlUyp10Q0VttNgwJ0NgmFfFVjrHBrpyft47MY2G8v+p8u7m
CtIGmEFY0+xZSl2zfQHB2sgLVtixQi4PdN48mk/cP94gXewfjoRzlu6aPgTqMZFf
WuVzRJgSgxE8BPy2DwZLNnDYmeAoc9gk+23vo8iws6KHOg7bxCa7btZrijC4MB83
FadDC0c0mH4goPHa2wEjxMkrY3UeOVf3o/MdwSJy1run5caR1946aR/C0SByqu4F
YBIq6dhJ2UVNEhnX0/VOWCvHeynjjMAVH6wPb1o+oiXwofS5dzbyYtjvLk3S4wwP
lAm5E0YYvIa9Ctjk5qupvqZg62Oh+v06p+Pzz8BDwCP2odGcRwPN94rllrp293Vb
b8pGvvZaN3938udS5RO3wahqLgUuuhv9NnDoo7WoNpM5jQAzLYqYkOj8Ck4k0WwB
klJxn/9zqkcttVo3UCVndG8sv2kC2Yq1Vq/PpB8haQEPc8tqzvglEMjj8yR8VGSL
KjRn1/BumxEtKKeM3TXGL0XkTA5h8so1RYO5CB8usRDD6jHyYm62nEGT8kA9xpZA
NleTDzh8PIgVNE5O8pvYY6Uq8/QKBqPH/U30P61URu6naLy7KBRAdfH6dwU2Mlcs
igOfY9BTmt60eT3GzFvMJx7nol6VfNfbzMaHTL53Sbn3z6ztqLpd/0Em4VHGSXoi
OzBXf7kljIWi+8sfnlaa/aiM8KIHv8j4kygDymnsDvV4zqt/P+LeJTl2oUdlDoFw
PoU58DyEKwyzC2tTv7BhbdwpqBOl2kjszIVa85zLH2rIV/nrbu6ldkksplt4Jf1W
b3UtwpHtlZcrEsO9uCPZU9o1H1uwsARTwlfShU/5BRIxsiuoEFUb7doO6qERA3yV
V8yu7wf86eKhs1zGlla9RKhIGdBo1K4LMEdXSZ85bu8FefKeYlLv+nY9CnM55SyC
HUJ4rFQ1gthQNWtsarn5cnQhyMQX4jocuo/jdgZ/rOJ3xhQIZ8ZH7XugI4NPey6z
Ov6o5Cyejk0KFgp8rifFZbp0fwyDnfvgNV0uObbxZSZK/auuL293LlXbNti42A7N
sG0X4v1ovtqRfb2/Kh6Hwun3oWVWAV4T6R3JP3TWPhJEYLXuV3UjaE4RZJPZV5k8
38BrgzfgVeU3aRRDrIhCjjZledXJLnYTXHYi4mUx5o504r454UcSnkGyabgeYpK5
TTIRf2rzE6iJ9y+f/A5Rx1H3rB2nN2HnyQv7/pRVn8eOh//uP0MG8wH/VJM3H8HZ
RDBFcQ/zKTO44PtdB1iST8/2R8FjCeapSfKZY6ehWKm2j6zAz+d4vbS5Wgunt/i5
Hr7OjdWG/UZzX94z0A8d1C0tBGyiwzJmUREFKKAJVTGqLpJKalzGWxrw/2mQFQyO
gJlFEoMLlIuVG2tEeNe8NvfpvyC3WcyiedREwSRESTgy24pmV4VNWBjLIhx16NWh
242C4WYoRb61BGJc7KNE8ckhZclr3dm5QLmrMMP1A9s43anOYI1tfMZrEvqU/0Kj
RzrSrrS5kmfY4Jd0RFal7C0P3vuUx0GPkApiJk45OhgtC7X8ugVPwTJaUvhugL/V
apnbfVcTKvRIcRCk6HcBOQhxoPdao4kIz+Q9InBMil3+eXPxC16/26dfYvDn8WQP
1pItJHKYdpXKWx5ZdPfL8WkzIAkphPTJbAc48AIGLJxRIRJUjEAWsCTfuaoS6Rcv
mBa8fy2Va9y8VYMv0AlPbV8PZ/IVC4H9zzrqgSytqqOAWcZSnqtxo8phrelUm25Z
vPxfLzx0+I/Bdia1EMuc0udDBOg1t/wW2PTwK5mPDwg4Q62wXNx2ZwaYt0deCHJ+
IuQceub5cq8AwrX0MpxhgB5UGw8m6uRBN2ZuM93YprLD/BwCkcDu7fzCWk8EtFOO
geigxJhoPEo6PEaWeENESwViE7ezInNfHnYfujApAOC3/ORM7cTHqjuAtp+TRUqn
Fbs2sHwcmj68iszExk3uwdNTdwUGYUo9xNI8GJJv+gxpMRV1keooYlRTkfnzD4gC
LCce4qHhvg6Q4RtxZZxLqonBbvKiSGG/aYDYxeaxjXuU2zODwLPptljdmgK/iD23
D5z8zoDe43xJFvWM5aPSFEOLK1wJNquJDwKvLFX28n00emUPpWMpgJKpqec8Vzdz
RELapS2mNPJg7b5almFu1HKIIxaRUyui+CDfKqOPbbb6AMq+rMvjYUlZ8ua+aF30
kWNIl6CaT3wFuCIwiyIVqzY3sFBc+qG4InfMnHP3Y6Nu6xTRskESO78W2PdBUNXQ
ubjg39l1odb5sx+QZ0FGW//YeH4OcpboxclqQS30QrbQjHqjCxf/jccdRtq+/U3R
LUfRO6/nOXoW5R05xN+8e2IhO2gL3x9t/TpCHusDsaq5h/8QlS2cXyAatNEXXKnE
+dYb4l3kSuWyYzUmQZhKvHO1jzKbuar+E38eF2PC3D+BeEwXezsFxYiUU+hYLW2g
Y7qAE/yT23iZO0/OzF4VypNO2uWRecTVmnAEuD6GFt2nebM4R08Fy/dM85sjWLC8
WX0GpApdXSxDlU2gLRNOLMd8zgJCWT0Ft+lb/kvNBGqiqzcZ3DA7PzwWsqxBy9d0
lTBEftEkrTkzHqvXiL40PWc7h4zIxxg/HgAWLEqPWA5S5+O2w/YgAku5di5tUyqF
zoWtg+td4elfQw6DAjKYpZ5mzJEez8no84wQOySBy92Ots2ai7qBKi1sfmd5ukdd
qZgTTTKDbMYr1qfnBhX23+Yo/860u0ctGGJnH2OPvI9uJps+TLxQmPv/VhbhsY03
PJBG3kZEG4Ny1vUN2KEsL3f1+FnwcEp/T6f4F2YLbqWosuYHz7L4dfruPE8Fpc75
wJtkjh0kyvcQZwXltocf4mxVdeG+j7TiD7z1GkndlhuHwinXGLKnybD8Q0YhOWt3
+6nSMAf7Ebh+0r+jaxfTjEgULs2jmDlREd2u5xrbC0aX4UW7g9MJyAYViJE80xhB
6oZzhu5+iTuKJfRD5oYPvDyLIT6sGcXeofeeTZlNCGXr8zVSTtgDU+y58xKfcAh3
bIVihtMzeHMf1I+DYHTQ6GsTbg9/KhcooHCyUWxvTAPvnEVZmT61SlD1PlyXKo5J
jS5rMupQt8LSX2SExNoCoci4GFtmBgWWecJ/tRXlbSiHJv3OP578/N5hlQRKNmoG
7cOCdcLH63/W3eeFhbMxK32inGjCuapns9XYHcSd5iDtJ1npRjk2BsKVudWc1I3D
lxVFacY6XqIvnyzEcTdePz9cYUNV1WltxM/hOOh4MGyKFM/L1ONSuh7pzq24w6EQ
Ds0ByGr9ME1Hc6AhxZK78t2nFscguw8chW/IxGgu28qLHghWuPyXlIvB4cwA36wE
174zqswx5Pijc4bU3gLt8icQePVqRsSX9sJxdud/MRwQjnqeC10gW9oRLEdnwOXd
lNXF0zRO4pdpU/gfTJo279L3J8lSUFoKdlo9GMEfWy8=
`protect END_PROTECTED
