`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dpr7pPIgMo9bvB3+lmzGG23lrw5PE1Ez04UFphukZt1mJjrYgr9UQQrkjXO+A+oC
4ZNG3X0EjJy0nVhkK+CaZP/IoYY9EHF9SNxboEC6eNo5+LHsbhRAj1MLO0obGZ1e
RebSZjMOwmSQmkd1dNbvqYZsz5VGU3fordnDi+QeJO8sYibwINig+cOFoJUMf1i6
9P+6E2rOk5pnJPzCNpY1zNkM3yDZI78ANINlO8Qyc0qSKjhZ7FGdySqDjAdkS7Jy
Jb6tPUgzuA2PTok6g7SCHVGX35BGA/GhqQYsJrcqZ7d1E1nd03gn4tBJZ2LoApCR
NedyPaW4kXyswEn9tzTzLva7iDEEOUtqh/6VJO2Irp3+iGlfaojnzy4d4ARtg50c
ra6qIr7SNyukM4ZFk5kQE3Vbyll6eV7I6F1m+RKCioQ+TkIHL0T+S0dlC/DsmQsk
qbFgUHjKuJhyLdNGLi5AJXJ7tdxphl4mQ5QdKcHxnYQhp22gmmQZq8s32aiXz4L1
i1e2dAxREkULfeC8h6r1tYrTkCrjeHwtnwbGiOZvnj5b2D38wPJKgOaE+0G7+p4m
0Lo/gz9WJtcWc8tN8jxuytHtLYsxoFyCahSLbCWPuFTpgMLuYf8m8u1gz+Y7ACU3
oCzl2HL4wHSdG5ydLVnJfoOo7W0iKpS9WedxpgC5uoBezgYNE9tHg9dV08m/ocqd
quXCSCJ0KsLSuKUbO6IOoraMGRYOtWwhw5c4PX+BwWF9fLWIw598EnV+mKQPrS4G
iAp82/V6WppWLOovvVp7cZT/4b82ywsxmuXjqnnORsX/T37IOIGWboL4yD+YVWgT
8HoI1XR7BefttCJQ1rxqgw==
`protect END_PROTECTED
