`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EdAmt8ezr8vgz00Q5aSp0X6Y9I5lFqjtGdy9eECBes9Cd+KDqT1crJEyKc/t9Ic6
2oY/Ad7gdrzIZmWksgTLKVNv8ahmgVAaLNij69W9fNG5O9mMtonL4mfZ7UOOmswF
DV+kJaRY8NqLqM+VRHZmENKitU7OKGDINaV/dB3rKnJT7vIbrfLu2TcsbnL2e+qd
OOEdFBbZhDXptgn/iigGxA0l/uIlh/fw/Z6mDbHBDGJ6/hCh72FvlE5SeQhmRcRp
R/Pd7YAXqECPXuo/v+UrAJiLy8BQgbrOi6xzguP1k+DWPraiBenFpS1vZJKoqpip
p/fR48dcVQatlopnz16BUKO5ta9gTBXq3/k7iajfOA8=
`protect END_PROTECTED
