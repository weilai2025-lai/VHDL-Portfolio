`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrEE/YT2TY6sE4B8qJiENWXr1oTVTA8t9nQAp4MJMGvrle4qBWIPvzImeG2t4mjD
Bod3tpidpvuicJoEHvsmfvL/nQHWvMm1HTPnXs5iflGLbS2uzhXh4/WEm7Qg9CbU
lXs4TYeFHDYGeAFIRyUYmiw4VKqJOD77d4MxlyG/00CO4JU5KIqn8ufIDMmGT5X9
bwDo5F+0xQKd5FCge8rMYnNgcxSzP1swqwpPeZ7+S1SJaRaD8F4ohrb59Yi/b5+T
yn0OyWUBKb7xn/+rlBPVdsdvCJKSfQy/2OQ24rTk/1xX7pbuMZwbAND+kvq/f2vs
6HbjUrKmUyuhsHQeA7dCpcc6VprMfGmEK17MmUtkA0O060ggc1rici/jGSHcnrME
ErrdUEer1LNy4PEiUWnAC+LsAc23JPYhHWVniRd0TuEDDEkXsA96WPYzJ2kaqbak
vJHT2r4eYGqYb+BK28w8hvTTs4lITux3UOZbEKm4pqwDBYNPO1KpnTPJtiRYZUqP
UHCjdurT06r0iKTVOMmQfPNBVnZZSw/aYpibezS0FbeU4P2OVL539BL+XZfx/M1n
Bmek/eSo7SNesB2tFXWsJvB+JoH618AGA7rNKktrnnlIxp55Ua6HuwdadQ1+xbQc
NWPlTFplZk8MZSCsvoaJEnXsi9hjgneEGoyY67Zkk7QCTxKVURtVYNAtyjA05GbC
4ouZNWh0WDTUJ8arfq6fF3Qoh2MnxMVK1m12Q3x2ysSifo9tlxOWSPKrR0E7Mv9d
3uiy5n41e37L7dO4X49pXIPFSzT4GNbVc16Fk/yFqwidG0Cd4ZYPj8TTG1FKa+tj
LmMLTg/s+1frH5y9luq/9HpbN7JSpxsmLWo7LmYNsSuQis5ZCkdjYPirx1KjoWAG
cMwMlqsIQ//sWCYxF9hypbrheaMuF/CKVP15uG/t/o7FoZsOiDXo++gSlwtRHmwq
JDIOgN8PAgitAdFrl4ZoIRq1lSqjmSCTOGTWs42LBV9DdD7LhpktLaq/qVInhBU0
ajcAobvuXYOOMgZouBFXukylAz19BxwONvpwEhUdybHi/fuCLBcRbiKUSD2ZSZRh
qkYCmFHVQZ3nrb0Cn5PaRInCUQnE0Ey9DcfQ/w0mNiIq7dvh6mvMiNpQxsIirSy/
DjIGTCH/6xsw/OQvPcKoihRknKt5yJYsyy5mh6FSpoKRJaCcxiWp1AdFXAoWWkwN
`protect END_PROTECTED
