`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LJU2ZShnWQAI4eWwWFo6FeFHK30woagoX9YgRIrnkvYX+E6zPeqAFLacoj7IKfn
Ir396fEGhPYJSBt00P8a1KoQivoAOHlLp+9wgZ1goc4kjJi7rd9qfKmt+0yJRSp2
K9QpzMlOgEfJq3W54hjG4HWZYxP7Lhpk77lYbRpAPwqihug/Mx3IwahQ4G+36i4G
IEF+uF3D+KR3b9rBD7I6tCWpkkcWFrmks7mAztUpV050HGzuHJfrof6QS7Smc6Nl
YJ8nwBw+GRl8E9GP2s48RL6Ud940WZtu7xrtKakuzAtiLYmrkWCu03YDjX+qY6O8
A15nxty1CbxAIOwncAhDNZu2TUk7Z9/5zt8nXwsOq9TNM4zfPc8Hb8VEzlLfZt3r
shFYE+/z+8tHqjYP5E2LkhEdnDpva8sUUXtXyy7XBD9wD8h4CzZp0PIkZG2uix0V
DEFMsryYQStZS9+eHAvTBvPTD/58KhWB5EjPIcXRB2I/JXWbXs9zAEoiM7slrrzj
ES7x2OaIRs9uZmiDwB0GprNOM6b0wvRae85B2ck1B9znmfl2M5J6N6FqQyydI/2l
rV/DpT9ezi37GGuRDwrRB4TLzvS9XrdALEus1gPnS9A3nu5iB+Dk5NWdiiRSl8if
neLuhI05FS6wJE7itLLL3+1AekRC7kGV2FTjNgZkIpgMnrBewghNFk4GZRagQbSP
nRqXVDaWnXzFJ88VkbTtqJZgbW7HRqNj+hE+lkI7XAH9zyDXN8f2tECaLbZM3+ZH
Ec9sdxLhh4d8A0RwH1VAYLHQjHwPAJS08BqsmTOGd3vXAQrqR/3Risda4bGICcTf
2r2YRbCDy8fdHkV5tpJL5Jxo5Gm7KyeHsz9EjCM0Oyr9z/2qhIYTBt6t0+VhItmL
HyGgzHXnenx/SVOX0955P49Oz0oUhhXRszWhCuF4KFg=
`protect END_PROTECTED
