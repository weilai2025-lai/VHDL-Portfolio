library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- 這是頂層實體，名稱必須與專案名稱和頂層設定一致
entity fmax_test_pipe is
    port (
        clk_in : in std_logic;
		  result_out : out std_logic_vector(31 downto 0) 
    );
end entity fmax_test_pipe;

architecture behavior of fmax_test_pipe is
    -- 宣告你的管線版元件
    component mac_int8_pipeline1 is
        generic(acc_width: integer:=32; sat_en: boolean:=true);
        port(clk, rst_n, en, clr :in std_logic;
              a, b :in std_logic_vector(7 downto 0);
              acc_in :in std_logic_vector(acc_width-1 downto 0);
              acc_out :out std_logic_vector(acc_width-1 downto 0));
    end component;

    -- 信號，用來連接到 DUT
    signal dut_acc_out  : std_logic_vector(31 downto 0);

begin
    -- 實例化你的管線版 DUT
    UUT : mac_int8_pipeline1
        generic map (
            acc_width => 32,
            sat_en    => true -- 開啟飽和，讓路徑盡量長
        )
        port map (
            clk     => clk_in,
            -- 把其他輸入接到固定的常數值 (tie to constants)
            rst_n   => '1', -- 正常工作狀態
            en      => '1', -- 永遠啟用，確保內部暫存器會翻轉
            clr     => '0', -- 不清除
            a       => (others => '1'), -- 給一個非零值
            b       => (others => '1'),
            acc_in  => (others => '1'),
            -- 連接輸出
            acc_out => dut_acc_out
        );
		  result_out <= dut_acc_out;

end architecture behavior;