`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXUn1Uz4F8szlBzV4wE11ccLOeb19FTpzFSFFRto9TVh5DJSMP33bTius3K3azyE
WeWkoWCg0sSm11CEX2U6tcrvd0zyKlj1QkETLpu0zFR3nIFAP10RKJPJGHxLATtQ
5Q2vVsc2Epg9/MAxYJo0bu6PWTAYWJlW1pe19nbZmxCXGmUkVw6yAHe4QLolNfXc
oQdd97gY9H/El30yPC5sQaWLka04oq1/LMcs+ew+pJwT1wTt6orHeItGoCn2msWN
8LzafjdBJZGO8zc1cVbxwQi0EXzlbxfl4SsqvAZfGCXg6CP3LlpNQBcETIz8+iyH
xaYhGZKB3za432y9oJY3jCH7Sh3ofNXoloEJb+AQo/KCMcQwQUHaoSjZLf7sBU7c
MICiAIqaCmPXJUck9dN3MncDTRXG9uFr688P/gMuba/aD+D4afqGrunFar8E3j0S
Y94ovvN4pKRBpYn6kZ+/yc8Gk47qv4+v9dpBJRwEgHT+uD7ac1sZt5rhJtcLWRDQ
rK//llrI+W5s/7tGFc7VxFLxzsHDWasB3YXz5gG2nOw0/gCV2YRu5+Eits9M32tr
W3TLoAblnOL2RgQnUYqLmiATfeu0E/Ur9qEixhSsFfkEm9hX0Ikg6ROjQdQAPb+r
xUgSw3uALUgQZlWbJN5vh3Fb9liLvi60KN0Ma7MgDpOt6jay+w1a2ZgJy2IwGAw9
LPPF1nQsDyHeIaMbZlwAOGVqtf0qJEgm4m623igwWEr/IoEO57v1KIFMnyhq1LeE
nO/+OD4D4mN8dBHN+ksDg2gjnBo03zaNV8gzUG1TQ9QhpgJTTemChbJm6upE5YaT
GwhQ0eQnbwGpF5JkF6EW35JC1d0F81dsf5NenDMW97z+MmrMqaHFhBZTxavASZpf
Acr55sNALIcdz6eNT7QbwL+zZ5AkUbp8yZ0/ZC41fVM7WZ1VD1B8B8mWGRrZJFRT
bLAkEAzWirn91sWiPNlZAnRTFKXFc3Tip1fNVkDCJ/O4puUVFJDpNGTTaxtUa08w
xYBbQbd2DwmBPhkkK+DOmVZASXBwkyKl2LKzDnZmf3H5QB82xYT1nxlBBKKK43iM
eTRyPH5zufgYPZZajLzvg8FiUqi0ZBZaeGrpg8tScQbZ95eJetdyPfy/Ba7w2Q4W
JBRreh0u2DuP4lTX/bfvwSZ7cUQ2t9X2rDCaiEJEah6nCV8a0rOdN3nJc3OqM3+T
l7tafyhcJz6YSa4EvAlh8G2gnhWa5i6/+jnK7G4vkTZf74JhzO3MJnCfj/uXLQ6w
p8ZyTjLdU65Xd+WrsfmB80cMfiRHLQojp9x5ZYBAoKlnx2UFclYoc2DEqYjwgdDA
W4nGpPuXLAfxwJHydyxfRumzCRplbvPHSvTi5VmRkwn2iyYJFNIGEXlrIasQV66F
wdfpD1DkQF81vCjfglSaq2+rwGHokhtqvhCOAieW/1iyvL1hQMR8U1tvENaz6Zzc
WREywoDkZzz5HCAPWU8yLO6Vy+zILDIKc6ECWMc8vTv+pZcka0OhzmRbOTtN9Vz8
N7wCsWw4TyMOPr+TU8hDwDMQPLxC/Tqvcia7ugNFkS7BP5++McBFcvOCvUh3Imau
gFBXkIqtTwSfjQYbYADlfIRbcvnbxBTwJcNmTzIUfbQ=
`protect END_PROTECTED
