`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ja8/g22MubfTUVN6bzwEnwsz2IZ0CD02x4Hilor1BEnM+LxhQnkEX4pfL6+MIKrq
l8B4cIdwiV5en0vnkLYcketMDfuboAVFFnlhhKIF3Yl2tP69Ja0t8wVllKIiGDEZ
8vAQz2ZIMml2H8dEOpmmnyiIOKjff7IKxwkh25TqTvRuMXDEfNDZdTJe6DDgYA9M
8Sdm5ASfGgv8hieSg2xez82cnD+szI7IHRi9Can0KQV7dPLuuAwTVwJAPI7HicXe
HvzaJUt4hizH9lajMVSdaVG4D16V9et9cDf/oWScVutfPkoQkZh5JnRB0KXE8Hmd
6badw6GpoEgInmmqIW7uOcUnT73O4zzdmA7ge9ABmYfOvW4VfPMj4vi9Kiqi3rL/
PXJxy85anfIMtV8FKHAbYd8Xil/w+mHeZWNUXS8kX1YqhiQf25SUS3UZgXzYvhg0
/DcYZqWscxL8lCiaP7MtSX2Amz5nO8OaNFkUC9Eu93nXUknnfOjZPaqrAlNH9ytp
qab4CvESbEZyr+miktmCuqIJKb3OafPZbSqBT3sr9DCpm4cMs56I/xdjdPmlLi0h
hmQek3pxvuhOmRMEumUnwky0NvyY+QPnhjVSi5rjwSogjeCFugCwSqx0VcuHsXWF
5ZZp9sIq0liKNp8UhA5Mym51V26wWcz22gqhTBmjjsTPPCZ6HhFj/BcfYR3QyRVJ
GPT9cKVG8zBR3uFw49EHIHWSD3oVY4h3vU+qef5qpV2tVd1Ry4JMTusJQiPwMfkd
8OdNj5t8cBRofFcR6Fu+Mq2yNohkz0Kw8Hu8doavQuvClNCk2kd6UKlOUa1Jjq4J
Cw091LsBHPiM69NvRVoYpjTNEZr1MU3VRCULyhuzYkG/e48cyED5B0dG80WXvnul
Xf2OzaW8b6ttAgtg+noaLwYzYZQx8fhlV4re+5K39pD40w16kRivquK9ZPyU8w/x
RxAO+3OSjHO5thB0erOcU3cglmqC7Tp+9FDHv6f7OM8oeJU3oVwhuYpJ8Pl7bA0s
uCgeN4bx6kKDZnMSxTrAtFEtM9tL3yerJIELdIMQkXMuhWa+FWfuB6Lca01cSmPO
hdTyF6t/dFF19Xq4zY73AVLn+Drr5F/+mn4mBssrsqQ=
`protect END_PROTECTED
