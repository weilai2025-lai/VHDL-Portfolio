`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QUEC/DIEdFUl7YsWAVzpa9hq+OriRbXO7B/ezak6jnJLJBaIbxYZjddLguWz4TQQ
Q5FHSvwfSverSZHsdQTjf+06q+C8eU/ePaC+ZI24vbSQV1Mrm8iKBbYmQ3RJIYrZ
VU1+tACL743JM0WpZR7Ac2+ufKzMqKCVi0ZMAf8fiOjHZVbVRlIk8qfBOB07hQ0/
BpLmcf070i5HUXCsht5zKh5lj/iEbk+MkHYaXr5dTdyQ312GmjsY8WJRYrQGkwtz
eUbextgeLgWyas8fO1fXrBmZmdw0cdorVscloG84UtS6mW8IErlaFI/HhrYS8+HL
zXkVFDH4oFn6DZ3IYyhAmfeDQcRgOLpeQTf8ph7bd9jgZafPeHbr5xastfsCNo0s
3wBmitc7FK2Q+uxlbSTYs9lAZp5r/OFWSjdSHhNoKrLkt9wKpDEny6+72Otr/JoM
R4g9esenjO4okApmoEAOhZbkFGfxVt5cQUo+ucDieegelhMiAAIP5jisg6RYyGEr
lr2xBCECgk+8BTixgp0QiDKIIRdy/b+jiBRCvUikta3VWNNU9U0uu1lFWDLH+0Oe
SEVgqNPwap6yVWXlqNcx4Hr9kFRqXrmKI7oFRivZEqjEYQ3nXDYVKGPXzHfqkpqQ
hCFEgiFSb12HTzjuxphg3iovb5TeSFO8SWe+IPiBWkBF39n49pZJ7HmNMAoQ2Jlk
K4cfJN8GJ7tvu8tzhQPzZ8bcqDymfCN7rrNEI5sU1gkZU8PLd785AL0sjwo5Agvm
Atyt0zrfSCvacj6EIHvzfthF7oVHgiE99t9NJOfz4VI1O18p+8Js9oWn4K2bE97L
OWK1fS9gOXM0phSimcH7SsSavBykz0yGzJyp8AZqLmDTuDdfjAyWg4diZjxOT+mU
TDPLyUXJqQlMqPgKcdqozUGXY7utO+xypQp6AlKv/kOTq5/lGjOXLEdT3HkcWr0N
pDXKxtR+cYpdqEHmiJAMTT+oDx0mGcGDIbPfRMD2fIVKMILUDtjc97l18mhIYUdv
WIsaA5R/G83/iJrQKQkPBQHVnPGhXn+ulFgZhePJo1nUvSWm6KdgKOE2lLrzeU9p
1rNpWlvJXPO8iW3WT5+7BfLixEYvUd1Yufd0s8uA/DwRb0JpE0grtyNwpVT9jaDq
a8u3h9EoTfPEdCxpkRtlNqxDeEWkO/xUiyU0Weqm/0iFbFwjG8mmtzMLP+EgUYgC
fqxidf6gPuku2G7M2ytTiGMErgLXKnj/wBDXiw+89UFQiJPco5We2JqLNWlJuMLc
+DdrNBqgZNqIUhobWauRWPQEjBdCs8scg+HLIxvo78n5HXa6diDQ6On06HorYA+X
8zZXF38YPUcW01Q752/bYgWOaDKMNKiBZ8yk69vwC1dnE9ufv8xMYLfJDNswfJIS
MuNk31crWnqlbO+ytMpAvA==
`protect END_PROTECTED
