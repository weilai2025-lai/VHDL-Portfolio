`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ryIDI+y2v8WvMxMqtVhWtNEZDKFqGEGGcfz9XoXuubGdOIoqX9rFO9tn/YQcnBJ
+eN37neh0jUkcx1FH0HxQiiDnp2NqXZjZwm4tRTcUsEU4n/ZJ64E5IDy9thOkLJy
8NACeUMqGgKC70PbnadN+s8NWgOArjmhY2Eh6WvBiSu/aicuSRd/CcOmVn+YvpUF
eazLe/s9T4kx6cPzPKY5+Diwf08wGPz50FhWqzjoP1CztkJm7/2wTewdH7gvN9gQ
VnsnYhg72SUN26RhADBA+Q/xdlr6So5eo/cXC9xAOgV8CCHJ2cc002NE2PHToOfD
6Mnpb/KnGB+LA+VXNuTf1hnzBuWgHZwr+NFSYv5w7RyaDjx6HbjaR6q3Egs3uVH3
X27RGEG6gA7euCd5NnT7WRlWzXy8SsHaO2uHQ4QeyAeBBl7fEkE3+JWhPbP2l+/d
MiN0RctY2xyf8IvhwHSA7gZm6XDiHicIpw2KueYZiFHWeoxGRLiOdH9dglb3DGPM
INS2q3xvbdnZ4BMDtuQwBHJ+dMgNjFjHIBjBWPc24JlAK9lgIIV4frfwFyYRXRZZ
M2s3kQ55V5zfnwh8aCA8TK+HGhHm9pvuXdu8yPTmB8+lh/xl62F02GAdZvUWJjlQ
F+kkGDbml2M9Ov/LdJDlheBt62q91LQBOMyBpoX3cRZ5ngvJE4mAS4KLxyxUti9e
FPlWIgUFU76ImLedbnpimDYV/uK/7I58/FfsAtILiRR6IInZ7LTWF55I2M/EkQRb
vEueVqcP2IP6+T+dE3B1JT/KtqfkoTjaCkqOxDj0w2t/XdTbiwEkTCyp0b+oMfEs
sh+H33CixyF4Iigri3Jxz8+xwgsMyJUcqKS+7EVHkTe06KQKIE2kTXlCQMbmIIOr
Hr7O8GmssZPgSrKOU5/HtZ0sCrMliLyRmePLg15DlfJ1M7Lt73INEd3xYhIQlIuP
uKqQ1K9qpvEPI8Dn3ZvGAIyl/2jfgoG1EmMkn0Rzf9c8jwSEv/3/2vwBkAepqu1G
ePJx/G8dQrNSAoWSOvQPaPkWUksk38OUu7PZhdGSff9bz1f18++sdzy8VGzZABKw
I1DsOmfIOY57V5fiOAPBjVgxvisF8mDXZpdSGglL3y5aMICB9dB5HnSoMapZphas
WTrd0tJdUtAsEPzzHsQcxG+kzP8T5mllDR2lpyaSvZYahGiHC/7nHjPA5oflHSjs
1eOFSZwPB82IzQzifi8v+vxa1n1X3npajpHNAEq+fUhrmrXS2zuA5RlZBs/7ABhF
tuwvgMxtEjkIRJkx6cM+aMlDl/PPwOankuw1V5+55Nykixxf9pCPEvBy+j79lggt
gR/sTjP3U980n6RK8YWBRHz1rwEUQn8giQVNT4aAz22OwJ087AI1e6YL/8JrUj9V
B8rsbz/afuqENj5mrMd3QmA2R1+bImv8UMfHlInbM3ZkqSdvS5+Tpv4F1NhDcu/e
hj0k/ldrrxME7Lu1zGsgurf6uaeGnvXtfRGmRTpWMZR8T0Yio3ELJmaQbHuQtKJy
uIJ+1BKtCHtCVqQTwbFiFVALtp5FP3ulc0WS6dVQHWrOMi68FGY/Oxuaa4SdDdhW
AB3UTSW/7hSRMw53t5eI1KCdhUX/r2A0uhjE0P8jcXBhHYfZ07+3O+eccRXFsfub
sf6y9eG8Pwi+z8A/OJJhdly2GUV6rfzoRU/TzEatNeUjKhSJo3Y7+ewOvOKhn1bB
YA90qjq40WAlf8DZ54LBAJResiFpSiPO3COqmpczKYbtzOosf1HX/RAFTPyYI7Pb
YB1mo4H6xqH3daXgFba2a4tPMUJcJjOrKYxBgxnUBUPKHw9TG2emTsOc5gZ9PNmY
28anKOpzs2m4UsbKsgf076timm8v3xkJI5KEDgilGMtaabmJyk3s/PrEGustv+fn
0aO938K7lE1zLFbRdCuD5k+91k1dIvh+F96gp64XhT//7x7NTv0cta6i6beYcuNa
CAZIQeVS5cm6LZU9+84efeiAHw4l36jYGZbMtZL5Ezzl60R1knue6pEtrvtblPZw
tArVRvJqfXia3XiG5pSwbxAD6isMexRCT13qgWlTifczHQNb53mOkMsZeJgtV6CW
eaIpPP5WGTucPEvrqitHOxcnDGq1wHG1Q2oRpKERGTcTdHcbsjeuUj1LlMn8cvW6
pcWEW07FozADkj3nE0Rn9fRfEObJ4mm+RcQ+1jOhY8KLCqOaq6i+WvjFoqejcNtv
RhCsg8KYrsA/DAAv/IqkWict1vqj/WGwXCS2U9xu7GMdnNDGhMOGpVVOPX5Hpuio
X+xs5A+t82AZ4wIN9AFQ55InHQovbd5XTPujtMprig20bGqoeJRXb5oSujCp2lcb
AXJPDpXx8njPNZvLMExW9VnyFe2nl7wwAo1q889V8fIKwoWcWrWmj44WvINXp3d3
n9BBXfun73l6ni9VRAUOxyn8iGIPvmH8lR5W7tWoFvHkTK31ED4BNDmtdtlN3rqW
8jHkkx788hTZPKmtH4MFS7TPENE3HzQJG+lcMNx2PgHMiYwxZsb3jV+0NasECiTK
d42WCFzW6xA3gdRCCocOPdyvDcWmrABgwAz6LUzFkqYy5BTjBtmYyFNgS1fZcOw3
FRxXBAyC9DN34jQHPk7vkiAxFMEHEYt/IFo2+py3+WtFOM4s6ECtNmRA3h90vI1V
ziB4MHVYeBIuXh6zLmkyHRP74CRSQWDjYrkHasGbT/Sl4Lzus6n8hNmvVXzl5lrf
KYs9uiuqXLhiTobgvoVl5iEKtQFfqQoGaNbb9qyfI1BgAI7bjAUYuh4tRuUQ8ua1
+0pYtHk40jbFHQ1G6DnMe62duKHmz+4JUVU3hUCGcw9v7/tb+POpGOMF/GsQw/Do
Hv/Prz8tAUF5VGDNoKMIq2Pi43mqMI/gxRB6lbKbaIMeHNW8Vr5Xqx1Rnz1NI6bC
5fnBncLLcGJvsHdXIY04z8NBkxCEH9Ppb4doLcQqAjHx1Qi0jSRQLmDaN+NVFprB
NRedGJnVHOfkOKP1ZtwoNUNQsxvQsrfh9TaKl4HbUFxicbQDxdNyj3KeqzIjBcIc
cHIG9iEDJWcS67Cy9Nplm6T+QwKUJIVWzFnn1SZeQZxbXWy3iRefKEL1e7lqHAYe
oxAtdw8aff59vN3ZDnWFijbvfl56Ya/hmEqJZ2WC0Yra5tWQNrUekGpCdWIfF2Ie
cPisgCcFBPaZy+Xq0ImBmJoI8AnBfywqa/wxKlvPwPNORg5MM5Q7A9e3ygKgswRg
7hNMupIV7qWI2LNtmDflDLrx1iVGK7wYBFOmMaen487dTSGobtQO6+mTBjmjjTki
QZWbYqruu8l4Up5LWiXlPg==
`protect END_PROTECTED
