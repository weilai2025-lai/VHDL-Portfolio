`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TspH0GBNL5n5Htx0UHmBPPd/FMhutsl3ozqPkCZ2cNQgpaXr4eBYDDkjNeEgWaw4
F3lVFRWx0msdMecKfHihvCIzrIN6GNupSbBHoky/jBkJBWDmsZryNhepnbCXQE3s
yDNpsgRIdPVWoTC0fv9iv+BgprigNxOZ36uZSUKbGugsTqFCEQ2igBHbGqVTgsBD
xwdMS6jijdBH8yAFoi3e11lc64DVmDwTDihQNqWRLz6CGS+bAXs8w1IdYWEpnlHG
rDA64FDELatZLaEKkBoc6SGGtm8fntUP0VG237cPmNO/Y4rMy2Wo2ochIkDo8Ygj
5sn8cSlMkddz2BSAkGa11NBevuGJ+ev5pRaoJ2mUxXJOoXRo8ue22hYUXPfypA6A
TQqtD0Q3/WtvgkFaaUkNhfWChOVGS2HOgeQzN5uE9E3x+VOICOh7Zks/81iY76O7
wsUKM01fikhUNbndbt0RYsc6TObq2/j/sxGBKHd9pBH17Jav+JkNhAyMFii7b/a4
1uo0YraP6uV7kHEyLY/IedkiAiFN0WEo9GgF9YTYuipm20cQzxwVnWQHF+QpHwya
hTPbz1GoXuQiiOw63ivM6XBHCwLkLkMWj8c/o1cVzNOGXOH7ukAlr30dRq7GfILl
91IoIIXcFYQO3l0SNd85o0J5RXffWkXf029aFCa0AN1ACMHJsM448/4arHdq3Ocd
dVa1J7mc16w+R0lJnkAUClSkVyzRwIThq1DkTbwMPGdmAPxIaXXwTnIExfbcxoeK
HWDypuO3Hx949AUE3S0yoK+lgFJEduoi0GCP4XMBlvEJ1gC4Aq87v86WMB9g06mJ
ixpNopBmtmNiYGv8bzjNRux4WX6bVZEGpVUZOLdh/nV8U1gVXyhTi1g4LfnMqKqr
BF9eKTnYte8g7ygQBU29r5N93aSi4IpqpjFegoI4Z9xbsMmLAb73BTcTQRWSmyTo
8bVqtQU0zf5o85lAweimhbYrg4E0IoYahDXkF/zmRFM00t2fLvKtr+rWOYlqNZzo
KtjLiY7swGOzXpL4k+hi+hnCD3joIjQWkUWNiWuZZupNkQycvO4jH6W1eGduO9FY
CjYtBNdPzMSxV/Jx/FHzVyqRP3bURU71wNcrAWffknSN5cvVZDjnT9VZUsUquT8U
SaoP7l3HzjRKUNphkkhTeheTHmTE2XCgjjwinr5en5Ufon8x+523fIfgWoa98asK
k/S3iPgpDT2ovMMoLqKyH5Iz+QgPZMh7puLOYItNTu0e9cJhSle7lzwM1aQOIowC
Mv0EMENxmcx6jHtubkmX2w5cXARYEg1C0XY2Na7crmBMll2jnND6C4rNgKpFGnvp
rG4LEHgy0Y46+gK0zLCh0lTX61gJgYlK9k7tqnCo5NUh2pfa88nQ/w1Mxd41sMLQ
FiE1I9OcZ40Ui9If98LspviKOfH6Y1SNkqntKwZNrUorIrMNQjkFivN+eN814ApH
wPMKjwD0hsdX15CtelWd7m6wB2A2zSRgrlyoHZ0WOJSPJsVsgKLovtDl/6bvVLm6
4nC6S6jOxup328aC1XJ2CoPtaofK+tzyGmWjBC3ko10oIle0tAb0fs1vjDQCa6bW
19PA+n3ebV2hhi/ucztkeYpgQ4ZPIPHVVP7m1aySgAbMcttwB7aQp66zqHG46AcD
vnBGxX45Eewu5tbJRrFvhE5Pq8Wejf/nCmTmmCapjyXGJ3fgvwLMgUFMDTVlwyo/
tewMgOU0Bt5OEE8oPQ+dcEeWtH+J3kpJx3+U7X2/GvgS2c6E9vpKKojNh1qS7Vo3
rB9Br/KpmLyzkCNdnDESxy5j2twrNnK/yRttuucs8Wd/IcDFLiVVLUeJNDXcCqus
alJZBC2OAQsd7NzA5/8Ha/BIg+2rDNHxv6/t9v/sAoUt+SYUzsot7x8E03b2GoV1
m2UdiBVJpoZeXZDchaifG/5FCbF47foSevEfWGj9o/aOxXzTn3I8bVmml/aEkfwg
EiCL0i/VJfG4V5SLKQmNQTYn4olIqDEHbfNP86kSSbevRZ9Bu8zVUGbtmxQ/dUFf
HmY+urQne+T3ay7O8e8aMuZNyOxhJSBThRma1u3hS7AxI+5kzunNlpA16kenczBC
IPJkCxvLWdCQBAzd4Lp4fTuUNnKCm3u+M0h2mO1hbx0I4S+1PZ7xj0v2kIVA1CD0
3C2qRgF9FVNWJgNZk5u6sEbvAOHKTQ+1zhNe+QzdD4hFk6iYyKFpWhLIP/zwDAUV
A4G0dHPRIgWEpHD1+xbDHE7DbbNsroxjmnPZwHjYiXgQJAR9enwlgHPpWfejBsor
p0W+YvupweF5tXrtpp12MR5Wr865emQ1/8beJ2L4dbs7eA1grTHOouydng0CL3rL
`protect END_PROTECTED
