`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XulIVD28Z9h3OAKlbeHFmopwezape95BjftXn6ewY2GIFJhMT3WHBYMOoQdg0G9T
eMBkMnqI/vlQXOj8bdtRtbrfFtRD/oodCFsVutLV4n2qr9i38GR7P2K0ia8whnVb
pA8KvqoJHSiKzRh+WbiTUFXH7GX3nyQ+A3dh3CnUNQNKNnNCk8VvcD7S9M3Re8Pn
ey9FMAkwRG6CoUlap/ftsfA7v6xFgfLaMpEAgRbmyiZ14Yl6aPHoIrz+2AuRTrMu
ZUhaIWqJxTLu9aAYzA2lFPn4DKJeYMcQgL/WkPRQt13XHW3pKk3ZhYtUCH8i/hPj
n4Yv2l+qTTWrKdCAUmn2ty8Pim9qlU19fa981fr8T4p8r9NnTP3AaqbOE3NVrULP
7tuhl5fgtSocGFjqyFsnkGE2ogRBQ/U6H87W553dOeNSkU8dQb5DJVQ/8PEFhy5L
+Jbj0HcwhJScrBij2nP/eJDWEJmKzhX0/D98UkY1avUVyOcT+4bAc6YvGwZguqAk
rvCsWoLXUzTPZjlRWHWHBqbQgodKki+r88WozwH+pbggmUWT9f4jesIYYdgKa9Fi
AZ73P+APYbBN+4Pe85KbK2j2Xf/QWMMsYyOkG4Cpa3OISDrhrgs154H5/6b8JXja
K7PhM5Xi9H8ToE+aXIV1r6Qdges0nW/IK7N+Q13usv5VHZdfFce5EjZcaZiCQBD2
k3r75s+bTppXfjhtZtxRPZaQCG6RKP60lLrJXQG73hVG70txUpNgeHdLFjYTekfy
cHwK3h4eILplTDg86YhYe8ucNWWgQbzPQCu0tn5bvXFZl8CPVb6f/TD1I4Qz7TEZ
o1oHiS9UmyRI41tBuLiq+iiRTX2eTSyNpOxGbFpx/h/GIgepzQ4+CjAAOUTnkBgJ
/BuPE1BjQ7H8N3VZoFMPyomHr1JNvMfXKhlaTLswQ02EUhjgVFP6Y7/lH2f+Hw2r
+KWTnrkBPATgzDOr93sJXY191SmW/OTvPa5h0T20fEBfowy3rAqjBbIKJ5fzHbzr
JVRIdE1MO4mDwSojcOM1eg==
`protect END_PROTECTED
