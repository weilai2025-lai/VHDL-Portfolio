`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ozIz4VADAXIFCKuCQr2j13YKS9htnvXFDSwV3XtlJ0nYN+PajYpPLkdvDxMLl4YT
9w7pPYNuTcfz3wO6+zJpnIMLyuvmnM6VF88KFYpctqtkJvEG/4ojo8b75PrJEORT
CPagvarZ+JU/ZRHFQ2z5ZWmNkc+0Wq2msAfI4SnqRq1QkU24FnF1IBMOuTwAChBs
z2xj/wWavDQcJImZiGWCxBox6/Fzh9XPPnf3d57/gb2ewm5lwZ0/GUXVIR596L84
SPscL9rOd/AXv4IvcLGrPICI1AGy4shJQ9WHGxYkDcLm3CHcxETlFFtrelQYuQLU
lNRClzkrpI/vsl8BQVRu9fBOo7C/O/WlhyW58ikX7qtcwKAzHxUTxK9WnXkp6CLD
2Eo53WyhvwGXlnyzwp6nBb7C/7ZMRvMjjQtm1X6sKaBQ0up+0t2Hvok5tmXm2Z++
GsH/Pwd5bFw/eq2XIxKKNReyNdsWA7/OzEsSam/VbTSojmpirer27967XncnMvTF
YewhRlugaURkXb1MhaCGPBLyon9rpU9raJy/DkhSm0rrOipTPlJ6Jy+knEKVuWUN
O3PSvDvB8Twfo4NUNhf84pPK/tsf5YzPo0HQHfaUczwWx1pg8searT4dq+qCc8Th
yGsPmA8yhrrHsdKryd3edTPGqcA1nmj5i1v2cn0/Gh1MnDy6McqPeyvwt1YUHu0y
MMHRakCEah74lZXfwCep2lA1Fw2U6/GFBmkXGdXUD31/AlerftyNRx0MQ3mF8aGw
XH+qUZh7KIPU4esPG49EfC7gNe7AyTSe/bjped7ZCvasxsE3ld4PuKyerXEXMHW6
6yPbz3VJ9uie/3gXYsMOhrNS9J2roemVUiytnhw0t88hb5RFMVpfjGbFp8FkUJHE
f56J/hXjKF/nVmGMZtzImiXJcV0tpwEMfLRk+ZO6vm6Sjoe7ouUyaW7tMhydQz9k
D3cNLT7o5rOc/qXSxcvFjazNk0E/Fhx5jyVZVc/6KI/K4cVQBmwWqQUEoemXdlTO
b7/4HZ0UX0FRLfcBTCt5M7MwhHc2sBT6pHjWIRPRyKUPpIKsnD8/C4OLTBa0O046
eis20ut/isG1LrWQQOChC2YbE61EfrlpfnXOMZpd/XV88/+FZ56vniWe96N2zrj6
0nvSnLR7YwehseddhrRJBdu0rjwEaPCsJAFdipfXGBEh0gHkfa7eVWjACsNGCPoO
/CR1WZqM8ZQNsh/dwNHLsVqVGAm/V6G84XzD+DM6TFe4357lD+1aqt5LIBDnS5OR
`protect END_PROTECTED
