`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXVk4qr8ffsiurgCgjaXxG0X/X1BODZXc9FWru+v0+NGMcAjqrSS1vdFANF7dxBU
IPHpSXlkSGGF5Efvq/9SLms4Ve1PrSkAMfw5rhOlNsOrvsRUIlHF2BRq34BekVZ/
8lJJfnDR7y46V4UKHR7Z+VlldpJaI7L7VfU9S85P1F0/r0877ymFJK89+/eCVLYz
Z9rhfRHuM4lkwzHcFKT4fcM06Gm0OC+zWKNVumMFgsnY5ClGVe2WJGFQB0QivmnH
U9eSsrP5cN07OvJPURdetKm0XEWOBJEaZheerQ+lSCJFsCzPtxPoeQyccJyJdsE5
UXGDbberigqblVISj8wx+3kpQxkaWCXJS0Z/JknDqfuoHclQqXO7MBbqgmBAt56o
Iip5scg/B6WrjcpfEpFFxQ83b/olaMjNYb+sD3BI67wLIqwpAX5tBZTMYpKEvTc5
SVhVJHaSS+kKBPGRAUafXsFXRDo6E1ZUDgRaPUGZSpKe/G74CK9Kw4Tj1j0vQoyH
Pu8nmiwzkePVRoRNxzXb46IvrAd15WUWn6E5mq0kio6rkWKHcEUQqTDaJhn7Eo4k
m922VYgFpakcBMCgIsQSY2c5jvy5KvaarAwhwTdawnE8c8NwSbXFOYlcawT+UWHm
d3xs2291gCBBk3HX72+0nijrIrC4jFgK3ud6gj8AgJAsxiqfDvhvbtg0t/WruC1g
NjnXDvqrB/f8+Vg+RIyr/sbms2YMQaUxTDpp833rIDwrjoaaJIzMTKL+NoFSjg3T
tHvOcsILtO35j1q0q8eA9iHyoxtx5Qp/Kjl+iRJa5hH+rOy/hdcdPrZah1q+Ykkj
MPyrwW5y1BriFWMRWYxl3G8ND8l2tamsfdtLH0uhcYnyxhmUWGgdMwtA+pvdQjiN
MyXrXQjCOF1FNfAYwf4+kOS/YRn4mKi+UuS/NO6LJ7arCjGd4FWsYrURWThJFbGJ
FkOz3KX+puUSZkpQfAxe299QKKtXTsxmLpeinYIeTmOaIlmwTUMYzMmTjvFXE5nq
Q61PLz/TA87DGs0tKHezTJmGu8B3Q0QFB2XQ1mYwS/onk0+6e297pJDO7auyLu+Y
mofFNUNiQlK6VgxvfCRSlnl03OMPfX9LzGAg2foBLtHd4BK17lyj2BdWQI/he46s
vyPMkFmyHxjC/JhfsGHTtOZlYP0ihYX3YWqQz0F006DNC1r+nK6Oqt2qpf+O9m6z
oI7E/xdnvF+sdspiBdH2iKoThfXLTkcCpCiTXZuFIiQx6BZ4tA/k8O05T1qtOBrq
adIxGBzsm2ZvZ/Qc6FspzknbbDzFR9+FiBHH31tYwdjMEjUh0RXFO8mohiWbEzZr
wDNVB8vDFTpOtTdD+lAqxYbkkuY2w7KQF/SKyfJWJz1yHmGT1ynbrDie8PGrA+OL
+3N3PRhKBxznLa4mrmme00pMmUBzRelKW+iS6F7LIpFDU4nbMmEr9qNKipSFfWdJ
7AtQ4rNODDs06KMSeXW3kI25Qt/OWSTwdwFzuQ/3PuKAEZtNewM5OGU60abCjAY5
Ipbh+KZAWUfMhPo16FNLUd9P0IMRgHUVNA6UGrSHoOH0xvL3xl7EsS+RNersIYOK
u7DGVo88KKUgbvsMjQ7VHSQbzJtDOxhh4SlbgP6iXqiUZXBtJFmgVilyd9/HUxEz
IszYj0HzJCGr7BfTgydTeJX/O432UNiCTJ8Z5qwEZofyK0wVtMhoTZDX0eU7VU94
ZDV/Ec4iQUsVMBoDyWEjq9CNCUytLsQ2bqC3alvpifx2wzgUrdJF9/gVdv9z+Wz0
iGyPf1wXnJ1Q7Srngtv/8+6SD3cB9vDclEYNfwCZTHTML28/8RMgRJ84mpITs0GL
4pVu47NRP8czXf2SxAe53qc2AIys4eoUAI2vvz5Hp+h1lWvhO617wBlaK6yfO6j4
5gqCnCakBzn4ar0ZnECBTHXpTyn12cUtEsa3AI0vSuPQAYpMAel1JKdaD9pOEfuj
I8WL/Ge+Z9eH25q2z3lS712WXPYU9Y3Yn0o7cHVLIbidJCE5WfXhKy7hdKnMi82c
O1vvfbvWCM8K+gnpNA6WMGOiLdgZILylU5bF1i1QD28fsXBs9mVWruuWa70aCRdt
8YbZ2oDWIoEcXVujix2R1IfqoBHO2SggFTeMM9b1E3m9qqBns+/hjC33GxVFQKgA
clIiUXr7fHkDCzaWhVGKQEatIC71QOMx8A+D22+Wwegpf87JkgwUPY6DWzWCKfXk
Avj4r4L+SrSsJWhF/rzP5zv5h/un4qw5IAnH/N3DDVl/aUge9WzsZbT/06EtpWxJ
tkSkSWFgaJpeQJoLyZhjIGP9ISoJfLRlLVMPPJTR0bZl36zXDsb2CJS02P0c4JU8
ITvUwlnTnWPWQuJy8veVe7Myr2fRpdsVX1n5rJ00jB58wd6rfdvizEp5Zr0eTib7
DTx+JME0IaSn3fsJVcTSjmbMfCVjY7qcWsI6MTcJLz8jcE3EygP8kAJzbq+tQO9O
h+AKcZeTILdlj1yS9SgzTA==
`protect END_PROTECTED
