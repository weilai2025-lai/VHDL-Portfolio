`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oT1fuzK3rA5QeEWT/XwP/VgPkY65tls9HolCwsZh7PD8huLBz5lFyC7BNdytaWKw
eI+Wv7ofTACFd2xZLBsoFDRO7+hGZpgqMHB6MscIy5Pu9rO8/TIE1OMeM7VU1tjJ
kQIYtU7Sj6TZEGmJcP4VbbMFD7RGcFGKdSZASf4heb92eylTCGyCGMYPY2oUJkh4
FQoe3R2IFTX3Qk/VvB5mH6IMNOVh7BJ2ybyUBWymtkLG/XHgd2e1uLSlVIRH0Cg3
w071PFRKi5Z0n34HMndwDcaNUDNeMKFkzMrMQzEbQtxfIkJZDTGy7vxoABxiOutZ
ahpcPsz6Rkg8vyIOLbH2J5zbpNOupA/g+kmv1NNvb7lZi5vAB3tUjHh3pkNIZPRs
7EN373IHQQXCzNkAAEE5bg2hp+fK65hxmTkVBjoEWk74FQEUaz6pK3qh/iz97Swt
UWy8Zl6xy8vpo9kUgTHjzGUoBSrXfj5rxgs/7K3++KWqFsbbn+OcEoyGJ66V/3EU
+mWgvSG7nYAkBE+CFKs0iy6nDWPgMp0JOx5bUrogIbkrHX8Njx2ZCnj3BprJrB9Z
eD8OaRM3wGQ77A22p1NQ5XkomqLmJc3luCb3QN7T715k2jYp7k/8F6uPUbdgHcED
mbg82v2w7uvkwXxb75Fth+ZlhSNFPQveIBcJb+Eohj2c18jEANcGppRo5SmqgLva
ySaX9AhtydL37bf8Ea/2vMeK8lljm8rcvvin2guf+NGMoOGVAzSoglC7rgQPBr3W
2aZ+meSBGhIcZyv2CR5Y6g+nyEgPJ56qDeNCP9q2zdvfpIrZoXlq1viJVfcISXEa
YMsuSH7jDrcU2zwyocvFlW63QhUQMjuZ4Mh1EuqwqU9h+Qbofs9v6t6dElVZjIQ0
Pkx0bwvKsU97qrk2V7qj2SIRDItYnJwUAVpx45C2Rc/5jQOupXyYVo763mgqAtUf
aFOPujdW+REdu1EeaDAkJygZTXmP6rH8m6b8qSbBT2xJEX59/x5MxSmVr3A7BlDM
LNRHGZB5sG9MWMuNen9gUl0ZtVMea2GHu0lwpOK+m+EcKoY4jIq+rjoHiPuYjryZ
xnooUF8ASvuOhC8C2COHyKaZocuROgrVwSK5r+A/tF1QYPq5BlUyffGaUT3glvDi
zRntyaekbRotLZcfnImF6+szCi9LAfVSWoG1Wnz46tyRWnSa+e9Z3ongLAkPOZIh
PXVcTxycjMkWzSxTUYndNd4ykFsqwByXgIBqqItYK+ZjLwgF+9FtqfBgF8rv5SUr
M21SD8n76afjLRtGM57+3bnjI8ochY5YNztjfnWukMmCoDu6s0Ask2IzyTDQ02fR
KpeNRjUbf5qbiHE7RieDHasHHTbDjRJh7qtn1UfNQO95YAqNCZ54D/darMknNKj+
qj+fv65uotJNnSWj6xO0tByH7nKdYSQM7nBq5TIkqqH5B6APEZN3HBQL1GIwuw2C
eoOsCQ0OUAZQHc8+Gk1W/GM39foiWA3ybJIX2AKGMZ0vlY6aJdoRDiiT+mrz1BtT
VauYnQt/YWbN4kgH+PZk5TrMaI29i/41BthTJ4asPV6J/DXmiWqsbIc+lzVflAZ6
X0GAsLw5B6H6gDQyR09ybiZWZ3YzaYrVo3EFRgpsm+IrQ1wi9XeAIaFxB38BfrdO
CEDedsAP3GsyTYI7GtAdqCb9Upb/H5BDAX9DTDTN9HPiTR7+O5usTWNq5awHj66Q
dSSf4ak5XsGHl2Cl4v9JRbj+xxA0D+LbBxWMNP3BbXuVFQUSFslBlrHmkg/LvDEX
N1q8I8mBueXRssH9zCfiJ+0RI4sYJ/vXiMFO2gdRcowBZocbQ/7LGvn2x+Afi17H
ZrqvE0jjxUJJx10Tk6c4jDT5nY+j9eyWc1Vz/mWzBQEFFFNrte70GEatUWXYyV9I
3fX8dPZ3FW4LPt5cG3aLfHHWLn3vcnoe2ky1uAvvzycHFoLEr1dLMM+LMECKSX0x
IQas8/jzvuIyZQkiNBOAsULJiLRS4wDo7st9j3CTOdCttFV9HbwbZTE/ISPAWt6H
JW7uBHTZSNn0nG3KLtVY451VOk2WGp6i1yfCea4QnuFStPYRm03kEpoptTZSN9jR
98nY/ZYsm9SQvN15RLPaWoXuMHU7OD6UOsccCa2dZdCRa3pCD9mdeJaC2EvU2/cT
a/kKHK8j5Ti5JI/9f4ArcQyS5r6Cz/O0jEhlPrZNj0NxaAxe/Qvb7xmQU9rbIJQ2
gsq1bqzxrgZLV+03mNeJaiaxY4kNIJtGsyaktl1tG+XDT5pikESN0tFz+7t2xMJK
DTBzLE35Aad+FS8wEJTg+2sPsTWnMyY172pgGgem17Fm13AZcypwv0yzfmldMIKi
NvrcT8xE3fQ1jQ9lrz7Jnv1k2Skq7f5T4rPoChTAt4G204Y75OzXWB0Igfk90tVn
+QkslLHu08AxTpJErq4DEqeBnjMoRffx9RFsTozsdkbC/97Zib77fwZq4sSbXbd7
GLYhpyfEikRjbzXmN1wnXSzrq3lduPDpJ2KzibSNTJ4MX19GfqULTeF/TMCWVVwO
m11aA8fQgmoro37Utu0U9g==
`protect END_PROTECTED
