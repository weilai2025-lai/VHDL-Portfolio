`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Tmgyp2lHQvWSYILWA5r4jS23kvWb2l6Z2WJtyAiRZyCqkDmAgxVvefgHU0xJN/T
GTWChwi4+rG5ZYpz8gJ5ydEcVNIOYXEBD8RLVJbAvdxaFQK2uJTqaLsiMp7Y+koB
agzjdwIYPZiqjkb9UM0vN5TixX7v21/dYVPec/FsvTyRkwPqL7bmnsQq2Iqr+RuC
5ZXdA/AQAuIss1oPgBtuB4XhJL0QvyL86rhWDFihsGU1QGEE6pxfTKeNDxN2IcXk
yqbEqBZOiLlsy2ltVxRXZ7Hjy4IwF5WTPPBfpyAtzsYM3PJLbnYLa0aQbJD1J59o
QJ0rfCB5QrWKvK/SgE/oS5OdFUT67ree9BzjXHm4TYhLApU+02oW9K/lweuW467h
TXjF32ARuJ5veB9BXQ+yPneCl4UUtwPoiLzcX0R2gVgNr48D7WulIArUqqPcwdTd
s5pMgkIntFvR9GHH7xegaqk6kbfT6KrvhuOOrk2ebPz6RrT+q4R1297EBctHnb+q
BXTPktoIEXsUV2blw90hGhGVPlbWsoiIkPosq5hW4etK3ZcxNSNtvRejynLWhGFB
p1FSDqBM1Gtggh2zKuXtBg==
`protect END_PROTECTED
