`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAvaAoLlWHGR/SGvlMk77SDhFllb3HyNC7+YHNP83h4yTu4BNl26VNgN/tL0/bc+
lUku/xdNUDIJNn1+rKfJyhH/9x/3Njos6pjYTkme5tlhHDnQWjAHaQdOXTs2mug2
LjCKsMy1+reFXxL2JEUs8TF79qN/yfzhAJC5K5lmMZXU0Z4JcZQU2jePaI195AH1
KtddHplz+izFHMbT5USVGNQJb3UZxaHYkVmi/XUg+sjTMdtAxMHBBjuUNhsdJzih
4MUrJpwVrRqI6D50gript7lREYqQWf8ig0vaP6jGzz2y/5FHj1Nm3rOKkTngzxfl
x8G6XMXAgz+zWePSwcp2XtgmqbaVxe4F+SBZN2apaLeCYMgHRP37U2e00fDjcm7/
0pJZ/TjIMMdt7BKdZnuqw/I1vegZK1Hf0A/nsLJJFQPKdBRvdCRt3kcCkky81Rqw
zBrIZAs1jbYil6HWY2UAeP4HKL1HNRIDiYzLI56bhUuu3PQuEclAK9YyNY24ttnU
vqW4Ob+xYtN7ZcQig5hc60/syXonX829r10iZcFeq8T3OiFTROOxOxAJrwyLVXFE
kQRsxqzn/RLvQaMOZ6+0FNCg1qkhq+DUJjN9H0IZDx0RD+kwar9d4cAYuK7eV7hT
+3FrBZoHySb6Ms6GfcfHaAaFATP8fXSexlVNKU3D1SevwvAOFCiZOTkNDgIUurj/
xM14LWsZvRxaxix85Vqwmab8BpxGV8yDHojaH/zlpx0apGR7h3PtooeXDT1NAk7u
J3oqEFPgXV/EVbSwygLIvSeVHRSb5feJaRqf3XBWnk0NNqMNgY7/3M6I6ZpYpe60
AsOtM021EHNDfx3mkeNnPqeRBH35SoEQG0M8vd8mOChHsjWfFkgpJxwcc0OXG+V7
hBQU1F7RpnoupoyGHYm6FYgpDdGH+oHjY1gMpb7spqPV+LxZnVxbDAmvXiLbZTyr
3FHvnzU30vsIJl2n2pIQwIEj1QflLcMlAwph876BozLSTNA1Sgvr2B67L2hOdTlc
prdYUgt8H+qo4udcpHYneIdtWsk+BTl284if9oFRxJYbM6Obfe1h/CLasJYQ1QoH
tytkzl8F59EN8mAueURpp+LA4b35HRN1IKoHTTrusqAoD8tqNXp0SAz2Mcma2Ckg
OVhVfsEJh1NrOty3XZEN8shvyaCZ0b9ut/TVkKZnqKnoPgpf47uixU1ZtKp57I3W
FjX4xbSFuikyo3a9P+vCUln3FOkmCU9k+BQMM2felFSyNBXF2uP/lnICpfgPhhnt
fDUobnu143BW2noZ4PSmZsJ5a1KeKpogVHZeURnI5e428NiWiZ3cBaRg0fi6cTGj
X6JPId84T+Y69KaSLH9+Eyx/WhwYhd3MfHy935J9562RmS351MGzF+7D1tnOdHLm
KoDOnrvhP3S9s0cmkMQR1/sgRmJFzJIf+RVCyXgwmtGAkRHWuIrH2Nv/sLIyggQl
dQKxttB573asoh82V9pC+B/fBhE2I50iFmbLmG99BgKWLqYyXKFnF1/5zHSiOXsw
zbx+dJgiY7xa45LRTtMnYTxH/PpuARlgiHDwdS7OvmGq/+bFU65gs8LS+ufBJt4u
YH1d2snHCISl9bCH3taK2tgRMscYmGRMUFdojwqK7WYwHsSmuJ++QLdaqhkhJ3fh
Dw3mDjSQsCuw3uB03+u9z4GppTFNcBuW1UvmUTUgl5xw6KlRZOhqOMc0W7HerdLn
nKWWD20kEQA8ZMrjVsXoVARNs4M3VU/Hd3Ai08oRZjLzFzbWPB+0p79CTw120q2K
P/iZ33YhjAksSemQ0g0mKJNgeU2Y/ghJEHbctYtt8ucOcAxsG7WOGidvQJasTqrc
oZufEYzjod6tQlWirjoyI8Kr1owDVs9f/ZcFyiEiQH9WQiyzvRekOcOo/3/xuIqd
TVcO/CfSVcaSvEgML5/g6wbsgYKDg/XLBj7BOHLrDxqHP4fw036WbNT4tm9XmZdo
lbvTvutXRMLWEp+RwrdLvPeM+wFCfUs6wLfys0hr95PIQBb5/Ev4HNm4xLSzf+6W
yUXh/O7VVXyBGFBbH7fV4aS31b90Hn4cNlslCXaiaQtxpesFCxRf4siZxEws0ajU
L5Dp192ixeOg78Vg1v2cjYqHYtCyWq64h6jYgurSeOGgRoLmjDxZcnDP5p00ID24
bE01lrKBOxpxB7JEwpnM3wLuWlP7GFbHWMvsY3DpHIhAtQmS6SVmjfi7wnAkLib7
szyGhcSvB3v6OFOCFJYwBwTvtfyCSZbReUb2YrcB5iZmrcUbiOSokgrAk40Dueex
F62r0GLYEz3OI82DFnwNC06gNlq4TezuPX48pGUegsLNVmoLb2BcOlTuZ+hu+4pK
pMZwxSVXytk1BKPpaLWm+m1KJancOR5bWcufSphJVa/DCXkeKThzLSk7WeZtec4b
ZdQOQqU6/FQQJdIStOCBYr+l5Tg8G/Euf1ZgM/yGqft1s6ZF8zYmN5MpIh3naaUN
HviTF/DFW4u8E3+q5i1LZ1KHKr/3xLM/h96ewoiv0qYqNywYCV9e4dMxAMr9rV2t
NUuQYbXM5G5Zqz5gHo3lSUwpNQZWsqINPI0gWGpDxAVapU2Vi9M7nHmEy5BajKic
zvQ4l17tPMbXg4fqLSrXbeT5ROs9U3ZxhjInuFd4mnTqBZzDjldDy55QXGY643rL
LSN5BwYLkdemkLp+zbwTpB/hZiVSXR91fr9tihDRZAKommzE4SwwY/5qHgA3Uh00
MzncFKLaAJhwcRp+/MDrQRPCYA3B66D8mh2b6f5s+axULF3TnqdZDZ2AFJSMkBMU
aoSKklQsFWaSxX2M5T/bt0Wk3t0eWWFgUsn+Fe4NkjVHBKsYcZqUXW6g8oZdYcNz
yHoPMGl8hL5YE6aUytgQmzLnaZyQOkgflJTs1CzIE/t3Q04G4dz0wwX76nEcoTtN
1EkpxIbECRCb2UaNHUOMeK+obpVpHidJi7Fiav+ELvim0dwvyZgCpMjKQHt2Yj5w
VUhuwOaxEMIszwps0L/O17ltze/0qRngvPjue+MQqYLPmchhIdeGl3CvUgKfUMCB
un5x4h0fRdCpFgmjs49q6VQjcfwSLNC0XHEPh9ArmNnWTLP3GRdvMCv8DTr/XgIC
AF74n0iSpe8rUmOAmsyvhofyRor69fOZ92LQhskKSDq9uzLtWm1Suw3+0K58n7J3
OLOaYmtmD4fa/7N7755TmU9BTNf4/+GoRwuPyCsoRsxGZVAjrwXgMHU24b0g3Smt
W9B+fAZeiDQA5FpRwCwXVVNR6E/jU4uUXAVeJyoqGocNiFuACKkQojqf9D3iWrr1
nxVOztA/q6xE/Xde6yt/1C2eVQeoELUyEUmVgaaZfH1oG05giuBYGKXgM2mG1jgy
cDvGfAkjRA6BZ/jEVC+rC2OFFj3WajdRpwHMQO9rgRgyg9Skir7Ey9UXwa2H/xGE
nO4X4bxNvPk4CovrrI6GlmOfM4ruXBTRiR78ayI9j/WXxVNg/o+zgMk8T/WIs0iZ
Y8P/oh8ase7rYlHKrxmrK3xYfTh8w28mJVoCMyUQAYlmk2vsFPtYrv6fYcnK/ant
59owi2PfRGh5XPzToSWXBVcVl4jfEBVmjfO0AFdWiCTPVh+GC09eOkA9UxLrGJ6M
E9pfP8jM3zxtW9W5G4cHPqXHFlXdeK4oDOurrkFTbSBxcikHN6hFiAHVbPxE2/LL
gya4pbGJoilIPFV0Cb2UzqqLRcz3UgrC+nCak/7223OGV9myUCRiE5Fgw1zDFK3K
jdZjNwEc0wEawj5kOaIGRK45Ved4DGFgwJ0WTu65ubpPmQTnuraRiDyiUgYkbXZE
/smQfJEld03RlbUPwiPLacHcYubmA9khTTR0DSQPOI7LMGWAZTHEyFyyf07Fp5FM
2q7aBGZPc0tXGIq7u2O3weVoZtHV4OAX8gjIbufBZ5a/dq8YRsHSe9RUkrrowBYZ
B3vtsbU3o3IT9TjCreInxeV44kjEjkjS3lpP0DAFwijQMtNQTo0qsRx/J4Ao31Ra
tYNidCLvny3WP22JMKbyO9anIL8xEOTAYJ0pdStyrLW4zXMHLvWFeK8uPwVwC3Tr
uBcXjcw4oNAsqdnl/smnX3VBKmOtDRzhw6h1raG8DaSvcCBoKfOm5J6ou/uiZsBL
1o8i4sfm2ikwx/SMcEVbqTd8DeaKcuf4uh0sLJLvW7OLGEqLB69YMHcp6+7zpJe5
X5Paji+mY34YIW4k/8QGXRhKa/xQb46pzpbBfZ7LNFcaJFnRBqdd5UX72RI81ZtI
R68MG08HjMbS0ddYjWd+LC3cBGVYWFfgayEK/UnmSu81tGbmpsH7D001uJkcPtOj
bb8sc3dfbbDQ/d4YHOSAUyp9D9b2BKJdcgHKxAi3fFmCoYVlzOGsPGYmSAVMv7yw
9nvFrbTG2BHMMwhM+hyADj0UfcuzLD+te6Bs2M9WepVT+QJLp97lB/p8MrtNuZgB
EbZ4Ovqj+11OssoBjOO98cG2CuqZDHvAeagb21VAFymcUPnTcLowbQVtucP0rSxB
qFPYarWiNU86ayYRXouEqv1w7s9Q6kaCzQzTs5UHigZxNNEjFe70JdmjxTvWWbHH
ZfW7qkN6O+waTf013MIone0Fg8AQncYH7WpDGRM6lsXeJ54NlbOh8j4ERaioQAu8
zjhflB/ftm9ZQLNqhC+eW8SiXf0DWCfssUfXta59crMm13pyl7G1U+f8ZotvCmim
BsJ23WyKKWsHsOB/KZRjbBGrwxwVCneQtsw5WO5HFGkQNRLqy8B4u7Klsyiazqh/
xA3teSrmnnRPEcch7x2FGuPODaPZjcn9W/3bsZfGaPQ/K1CXwAxSDogkyP49uBbH
xymNh0ASVBIa5EJvj8a53x9AdxDzllGp2/37XbNna0p6w/PSFvcM0GJ0klb1hk2K
BbnN8PG6WWRmM2il27C1vOcQX+d1Mw+rHmj9+DCftwdXZNbhwJDNBGyX8BkDKPB8
zL3gNXhnvwN7bnQIhcaIw6mwDHiY7twDCjLC5v0fPmVdsZlLB6Y8cR7rmBPLlhS+
14EaU6U5lI3iChklMmvoktFfAdaVpw92ydICTF4nx8LChWWKfiBQc8pBzPCp8wgX
O2Uk+MqImZzUkqhYB8Ar57QmnvmM7rqkdGDpLBIzn2czTB7fMXudpXLo3kcunylw
CqyirgzBtM+pz5GSt5PffNCZdtylfF4GbrWwYxowQNKGBJ981tPYa8QmgEv+UqYm
GNztZST3r6vGblO5uYq8fA2iNrOhfT1fmLRIeRDYhAMQIAqo8MA0evZdP6An2n2S
nFJFiRANPLGfhh7ZpeldbOST7Qc4VB5YDlhJq5tPlGWciLU4ohI5GKvcOa8T/ASL
q2HyS5H254KiiUH3fogUHDZcnUXWntS3vw8PYGWtTnc/p6XLJ5pC8Ww4RRFxEdWi
G2Ha2dcbZXS8N4kumHrZJ3rDlybnhgmkYE3zExKJQucJvLsj0LhZ8INl92aCO02W
maqsgrWBw7CzTpQ+/mI4gDAWT9lkKRMOFd/mo94wX1l4sqPF4VDsy3onenlJGrf0
EbGK9/TW/tJIqopDy3XyiFZUqQXmwrfoWMxj05I56BsNnsyv9VJjmtkytNgbgtr4
F2qeLT/395LfH+rS+3P0Hn9n4rU02koQpTnCj751Sy24M6DSarRWcQkjeTgQP32T
1WeO3cftceYen23ktxBUC/VP5mDN6yhvN1jDf/tZNFygFq+S3dMYNf3xE+NWqbJO
zDJCf3IBiZ3rP71GDhVIbEHV/mHBt7G6+r8AGgixOoCMhROu35zcFZCedsWboQf1
1XvLihegEQzlp9hJCgJt9q2PpwQJgRDRyXDwJ3knsLU70HS/JJHL/aaw9OAnQ70E
7kHZF7r2sROO/AMP9M7Q9BHKdblDQJY83zaFqIsW/eYhmwh80PO/ux2mjGmrzFF6
tLRHmR65cgWFytCQ1LRMjPnRQW2xpUlSEuSAbfeqDTPXvt36NHwqg0pTH01AGKTX
f88oKRZIAHPr34hoOmmVItSfTVszNG3oiZCItIj4hr8EPPkq38/Z5yPdaEm4oDPu
SWQp989bk0Z5WLGVZAc0yD6q2sY0MeSTUjoS3YZft6gf7vud++PyVNqE45aSkBKE
/IiLmal2KPAlCL69rlSOLiUElrCuuSUXEEbzskPZFuJrJ0GcTAD4dNscaZ4F1xZ9
WAwBE6UtEcJOPVgMvOwT9AFPtk4J0BvMzAXxzH3ZMg+3EzZozsbPjja4uwwFA8VZ
PNyJ4rSYKPKomPyOSEnr8LhXb1eZD/f3bPIpDs5+2L1J+KxXNKUJ9TILFucRJ0+z
ZPJejRp2es6R44ShYZ502h9F6nLs+zfjU86GGl52D5NRLqkTFEyjWHMvSVXXakxm
yZ0rcbKcu4pg7nwIfS/VbXlgokOUmWMNTFWfsovjZuO7g/F34tW1nz98cvsvus/q
3O6bcl9g34K0hAOtuSeVbOcbODyn8Ur8kS/z9YLPYnTa0+O57K+EVOc6RnDBT0Dp
q+d0hMVVnxTswhrOaBa7xA/C9YEgTeo0pl3fFQ+D3hhq99w4WbZfC9V/lULnTRk6
VQbA/4tBRab9MQF8BR7jEJte6Wz3+Tz6ntH5/XJu8raaRy7QRoj40hLFavxmw0Aq
HZyUC3ZPU1cIMQLXcS47w3rfg7POF/9bJfUB8FqKCKiZt1xLcAQViUjrePNzZk02
g4DzL1fX4PICpA4QZWpatu7EsQoL6GDO4sa2lwMLgOBO/1otIlhKHQmmxBwag29j
mMnJ0wTVp1Twn8q5USXslcACFRT7bxY5Fh5rDrvmaJU8f/veuO1YPKyvY1Piw/Dr
rDlavmb6OqLbBKG917+d0doFtZ7HowKJxlx+bU3gYy5tHdSn53niWFtSUir439dn
2qCQ7TIIrtlEUixj43iRzjWzepsUN5T0K4ghi9YqK0xsFbipf40PnFxsRgr+LWGH
RZoI2mggUC689NB4wHjpsM21/zy9B9Hy/x3LK9ioheeJyvjNgqEODCY8DRy+wBfz
c/OJrO6h9si9UTbXsDhiwJ1UtP+D+wmYE3xcphMF6VsGz+wey1N6jOukXK0aobQZ
RwS9wz4OJ+Ppybsn+ma6p+EuwdVnDeryfvJvizlVHAN9hoknu+8YVmgc8XAHrwvP
xyqusTzozh1f7dX1SHbNWZ78yLA6GkYGz6yK24/cUHHa+DifNnlpJTKm5fWvfYYe
cfFzEz5Tn5o8FfxdrGwpn5365D06zp4WpDRB9uoRgtocTm3ZDdMVgAxDn0W5KQxH
KNfYCGSDovyKxHGeGSTIZsfCLOiATq3MsqawvM9YkggBFFVDbg5HEaGi+WmFREcV
fdYEUMhqDf2hS8Uxiv5sGen7tSwqooXASTdGVfolIG4zHBDRKdXgu80jAMU5yg0c
UdpK4es9UCyyKPfQXACn3NwOavE2TuF8JilG4skijxBq6oPG/WiOVcWan0drAL8q
pHSXFcXxr0yoog1X3DKhxvH+Kx4JDQ/c+ilMT/RrVJ8KA22g+U55lCfTAtirBg81
SKeFeu+2IPuXrGOl/lUMZaW12AoIM5l5pSj1TJG+dLWQibgS5PWdebbJN6NqSIlS
+KyiW3XmL8q8gOaqZSwjSqNcxqrQ0z6Air4RS62Th6ZotXnpGMAVGz6z1kHe9H1d
YrQ7ZsiKMA6pitTa8JtgQwWC1JBJN8YQTontCs53kie2jvnMmj+jEeSyUjxm6TzH
D9H+tfdjlzwKf/V1cT6oTP57qkyi5uFK3/FTaSONnCnou2Oz4k07+lzENNdfaV/2
Rhn+Hxf9b6DDfUs1SINOTk+08KRuQlmLR31MVdECUX+yZuKxEwf12RDW5Pq0JhpU
SXvrQLK2KOYRZPwdXc+GD2AQV1+KSwEE0XE/jRwef8FYN555iNsxKLLr7TkWJdv/
PtjYxz0D+CEM6YeMU0i8Fq1Kq6SJ9yB5G/tqQnZS+V9CylJ8G546ZLbPR2epBjmH
1aSWMa4Nb47PJeEB5m9gY2gVA4VVTK3H/UaCgoGmzx3NaTOruaz7xNQbWTibX5bT
8fQMn6FHqZuVCUurSqT4S11lOjpn7HujdZIkW9lvSNFXEYL1fvNsU5blxedL4PBN
/Zb4SPsdtKFLW7U8hta1nbJ384ugMzoa5xjwdyKMk8CHM0enddqEvG3SD3ra2uUk
99l+CpCME7ZoOck0ZhWjmcQm6mVqbxkOnLWlcGkV0W9nusGcaGTr423yRfwnxezN
u74KNWFeYRfcMMTUZc+3rAi8L7rTgwQGIJEWYNmFdI9OpufdcHCgNc+cWkHvuIsL
9WXZoeI7BKHR/8VwRrEpZb/MghJaNg1m+I9ShvCdLuhW/+sFJZX0fzPTz3oReQAx
MEY93nmkJCfaj6p6OUBlAqxu11/kY6P7906LkLfBy8Qondu1UcExl/0QNoKsKree
9hctSMrltKBOP92epovBBQlQOYttrKC+5f36d3ofAWfzRnEeWV4KKVTbJLufHhrB
A8E2Sp7dgoypcjNTS6RRnDe/er9QfHxv1V+mr0SPnWg/tivIyuW7hcPLJRiFU9Am
0c6Zgyd+gOhhZWzgg6B82b5raO3WNlUyzR+A3J+Sz3JYSHUTTYk1ugMYoN+Vb1yM
fHNFmI2rHJa+UhHJE/5Ckb7bZwI20VPwQt7e7BbeiehTQgZhYT+UUlUbtpPOkL9A
6cg4I7rbY9RVqkgtoZ0BsPx1Up1I2QhBRtV3fQJHI8kzxVL/84NJmh5s5H+ZjK6w
hE64VRGy8Vek0pw9xU04Mm5STYxq090ekW2qNNyoaWpezkFU4HgcJ0gIqDTOmi14
pM2SJwn4CaBb/L8FtEWQCNnv2hIkaDutxFWNvfUjUhZTRob9+MH8w6jyGr4sYsql
ez2w8o/3SUQqJ6Hnw5NWtJW10WNAb1/Q5XnLKaTlxne1N6If/2+mJise9AyUvDy+
rynHYr2pfUVQjuCmDNBWrkLAKcjvjlgbtgqCHO1CCtkt0u6oYSPCBjCXSLY52izY
1BijqPaADzJQgDnWRVXsznUKLEFFybEgXcGenRJRjvnB23p4fxGdAfHJREUrGk2R
9y1yIYjKcQt1QwO7R+UBPJpWYB2fVbrNnVYSBhxkFXDWKtGCycxPbYs+lLlycNTY
+wvFxzOKkMHWyQkiPmDdimP1Ylp7mGqxizJiT8OR6GWp2rUZGdYEmtQBEcwaKjdM
MPNhuo0OuL6SV7GmHgOZs3LsyPGOij60PVlaly2zL8g9EeqjaiL3ufbkOqVbgGSB
gxhkGCICvNv4ngsDNu1Po8MOuywVL0FP9VW1dxJWKadE8xMZp3p50dlC4SZoUkSP
KPRUEdtKse68LL+NQgQGZGFecfcRS6X3ZdPnLBrsy6cFtqwHAhA4vmP58yx5IDnv
Vg+r9k9P8WCpqY7MmtLimi1Ys1gckm2cQWIuDnMmHa1v0eGRESDXIEA1DJahO23x
NBrVLdMR3lQTMsvWfoP7eHg37Y0aCObBVi31s3Eg7Vdm1tue2GXVha5LJXiM13kP
iGYlPxa7ULKiI4HeiAKuq6l2u1tbHmorIjatBCT8C77dS4prQ7zY2QAzexF7YHYV
KkVhxT007STMEhQBMEmwMGnEHgw2uVdnfb40dYAqHou7weYv34VFb6WKFuwm/OL9
1Jw8UgmWy01bXG14baLEm1Bms7anEyfN/FkjIJVJdB0T/16FaeHc6CxF41JXaHJc
dp5bgD3UatQmEzC9P79im5wVy3juJ2Nksx6mjkAmRgWQY7BsMGRVi66ggziO4Hbp
uyFGInLZDJuT8NBE8jXbxWZKfnCCUkw5MyeKVCpzyVaUIsYf1LOl85fPqP3exhcd
w7Q1nRuNnJxozxZ+4ifZtV8ZrasggSWlar5Hz+GUtgC32CRUhME0y+FW1xW3iioH
LIBal0vOu37NMoxmmOVw5my3nnh8Ng72/bbBKkLpJSb4cMHGscoRWwXmTddAnjVe
rpUEL4Sed7BWU9L8BPe5f6E4W//QeLBuh8A8zLz2UZBJqlGS0zzl0WPhucn8PHr1
2gFNzBRjqF7CboZtK+u2YwNXelAygPrPbVH6pqjtktLseUa0pOWdDWYbkhrIBhmu
0izeAFp7lK7uaamzSCaMub6Tdnrv8FXl4QsWdE+B+AdPuNSlUdfseVetZZ1RtXyx
0Oa5E3OM60ZOrRP6gMixW9HmtvIqj/dKBmsHlv46tKg116GGucyqnZ2ruG5VnqaL
p/s0KrIDrisUO/tdHDQXMKhir7wumC5YQRfTE0BsciurSS5ibRWpRoTP7hpUT6Ab
UJRgZK3nikGDB+mEBOdzwsYFBxuxCmzjZD43KuTy/e+O/0Round+oKzteDlgPfxs
grXL62c4d95vwvwW8rLG5x6NYD0wtofFhpON5Hoe3F0sMCdXcWc/XTETGtEWfjuG
3K44XyyUc3CI0d51QKzMevkAy/23XoivySgM+ecyzmKrAhDF+zZRx/y904EPXp90
6wODOG+FgBofYuktcFYEVj1mR8A6dL8xOGf5AYDPouYLVXdKIV7oM3BTtaFkEVOz
TeLVqXy22zyZcXw5CC8DAek6JqHiDSJBCP5W7zQqKzM0an/cmrvwCRSX4MgnbxXc
YWk9WG/GfOInGmhgIPcL/jlPmqYO3Hb1mXkp2L1+EB6jJcSqCG7YgRKtg+lWuQ7m
UbwxCfI9uMZgrC5uzGnZxEablidY0cIgdmA51BgyUJO30HJvclYfERVK1eBIlrxf
/xSZ3DMibk0LVVcW8ZImaMsVY84xLVne508pB1s3F+09U7Uzp/R0F0/qnp95mEUu
1dfmnB0iL9ac6cGWON8GII1yY20VpN4TdKady8oEpD07l9cCsOBnW4lo6g8VAWIC
UnizwhczMGtl8pHolqOxYhMz0cz2qfp9eO4FEqj7ChZAGmeWZ0LGKwGib6dNo0uD
LdQc5Vvz3p3oemJAttvh1BMupZPY/+sxOv1JTVuufpgSIGKlZ4/8vh+rMAzfEk3C
Hsr/rzsJR+hcNrBRGSw3xxtLOQPE8ylaK5obOaBVH8tei9QDU6+oBtD5JPDHitFu
iIzFr4OxIEB5d5dmrF0TuyVY78bF93bI2q4T7c3507Btnufap3EBgfl7f488i/PW
1JF1u0gcapC5m6yWax1zCl+mEmfCpPrH5OARcl/Yorj/z6Gy7HCDgr0X4AKisN7j
KNpZ9h9LGhMai4g5euZKb2HTR0amIzMAOPvovsaFHJhZ12RZBflzJ97dUArVvEil
E8ZVblFi6OR66VNwH9/Jx2KPXmNqSrBrRuGuYeAuK1z1Ed/IczvDdSc1wcC9ap4C
B1CBgxhVMh+Svr4V8c1Zk79YPqvJ85z8I5zNPhgFKJwXMvAR3YZqGmfBu4LksNI6
YJgrKHP66c05D1ZnrAoEmb/IXlFElv9i5zOmVB57T4l6oT7zCkiPkY/yueAYkrqk
Y4nmBc3SD/f57mAXxMH+SL942oG+V0BrZk9Cd464uJ66ySNrlkXYZM7Qj20PYxd3
wu4Bq3JU4kKS5PS16ehxIOHAhX6UsJzMESkvF1qk6Xfy6ZycLE+i64FEl+cPt0Ki
dhuu188799ZmRxTUXP8615rBkL2emmK9kmoB//aQnKfOv2rug4FWPkA6VOs6d/w6
TeiMxCF4K7i0UrEGGo8hDn1hl4gkEGAzMF+pd0oLx5Q30lz+I+XnNOkpXmCL/uP9
zpN0VHavotBVrZKMKJHN3KlMNYAWCdiYYG5kjdzFJIuOyldqzGpeDdY4G7jOHPGr
DbVjc83uBZUEXYLEzc1KIAcucouognbx+he5xRNv7blkCZCbLY5L1RPpcJMtUJl/
DMaBy2r8gXAIowfhrcQYvK55MZG+KCsq7d56oL+Cn0fboEBhFmJ7QfwOoaHnZ15C
EIWLapAAHTOOVF7xQscsdkcNDhUBzPwnoUluftFEAaoWcI44H2pY7r43Uhqzaz/j
QWoz+6h+tbYqJS2RNF3Xb6XhgSp932iD3dmlfU7ahgwIsAG0NMnbjjYOsVXshge7
N59iE9Q9P62/jl2Td8WGWb52snuqBvkwnElTAEOYLxELe+ty7e9oES6ZNsSeE3MV
KpcnxfPNozokl+NlSxKMu1ij+2l4S6gCtLx0W9gyTVs74BSCK++G2mHsKf6Ms+2n
UNjtMAwNjVy4IDkfh7KbKjSLX51cFC2AV0n+OtD4FN4B27Cq/BuB3X1ObnIQr9Ek
HyBg2PjenJdcT14N74+Fz0yu1bjsWbrZX4/z8BFY5f45xTwQTaT4jsQI5RTMnhgW
3D//jhRo81KNfaOcKkGyURkSPmBimbPFfU2+0Iwn9NWfX8ge138/XTKopyH58tRs
T4XFaq+2v8au5oKWxRu1bqZ7zlePHLhVYAA5ibHnSrdtKSHBJUvgOZTanGx4vkwm
xioiHKUzLdNTEZayH1nRATpZi6YwSBqXh6BrNPFZrEvDw6tYFN+9HO1QnEXQ77YC
ORvtkaXsqxWIdKpBLI/92H4vZggRoBN2GVtcNNlvBeKLLx8aC809bBeRJjPq0mzH
25kwKj8fX4kdFyZDD1FpqD8SHLqIQfbq6gIjBqaiP4SETKZIRMhaDq3anZj6J02/
MAwOusqhqETSdcSkWOG+IOj6Ix5D4hVVQ8e1oAZVovBKbczqFpfiVMUz3rQSFC11
nJXeTJRdKT5l88vCQNPRPAoXlf720GAL9rsqoOkqMcv35mlqewYaFgsl/weWou9N
JrqhS8wgdYpFpaOjgqOgS0mVFr4I+spSHFyTtqfrc3kodqdBJmyWsd7wApErWgq6
1FK6UMd+IgrpDUazj63jYiYcO+yGMkAl6sImFWk+ySHWK8TgnvM6+C8Xf9WGjWXU
nCBS8TkhhqpvAY/hjnMl2NtpKSYQv18NsUGosCBi6TYzi+/j8sJ5blGT65S1GLNd
IdzIRk+3B6bZenBBbky94J+MF5ZfQETO0C/sIS/8crX2ozlyNqdC6XotoYtY6Nc4
3KUF7yDzi3dmNjfXJEDcFwy8oDwxly7UunLHixZznWHBxFbwlW+qTIJiNGZjmJyC
Z7OSDDw7EUuAEQ0A+Y5T9YHdkPDZYJutoHphDX2X6SWUS/AXSkejNBHK7XPK4w5u
EEpX48gB/VrmrJjvaap4zifaDq6oEgW/GaMxJZMw4UXHgPVq/u8kweqaG6n7+aan
RlELexUC1QgfCMb0jwNbf9nq/15gzdnE+pk5hGmIf1ECiNjrj4qQjbrtuhtnPH8p
1cog/JObYvrwqmqKMfQ7tM0Dz4htfh9NUQAjUTlRRaVHh6FFxKoPQpstuQDF5VSb
4X1P+bTRne8YaOKc4BaH1g==
`protect END_PROTECTED
