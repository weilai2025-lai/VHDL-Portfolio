`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agOHGv+hm3xDhzqjzUekwJ1zM9Co1Cthh/tUwIV+PvGqCjrwlwxWDLwAIcOtnZFY
tR/eJ3wJRgMR7R8EDxcrc7EXZtAB4bjQ2BJgrFBzi9kNG2zApO7J/NaOE8xJCiTv
FaENj76Se5qxNF7x7KW8PRwHowHsE1Oy7kVRBMpjJjvvb3qADZZfQAwhQ37UJGv+
xvgXeQn8pGE0osrNi6ys5hzdcWbc890jP9I5k6Jc7eZ7xbPR4fPRjn4VLjsjTlGt
ld6odVIkYeBSDyON8wYX5dbJPszRDwZjABndYUuwCT2uTpP5bSG6Nk5Vo7zW68c8
9R323zBUUcelOnn7Y63TO7jXZuRp+pw1Ns8us5g4uTn7Vg1aoPIHcahbO6GPjOIO
3bb4GOxS2qoakrbrc3Ri4uKLHRwhXklN4Zh+9GS9yPYj2uCQOSnHMSCts8b64hJ1
`protect END_PROTECTED
