`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/rToEYfgNpgKV16CbkXz2zWst/kJKg8F1a2DPDd+vYWq74oKJbMeqBXQQdioJ4I
gmve2TQAlW5lwybhLzYYwQ4YM9/txizcg3MBEuLaCVFeoSzeV6kD8BOyuvkLBNXD
hqO30fDV7iGQf2qNGj/9iedJakW/54ZBqK0fWITpG2HVbXt/8Fi0W3qN7cZi8Grk
20N75b5wU80PXtBZxwZOJvKuqh7pQxvYN9pHXFYADUAJOIUZQhkbd4d+v3XvAy/+
eE9N0DAfm2XSikwxLtyAXIeZfxBclW97bWOM52U/NmYHeqSi8/f7x7cnCRDkOAZm
OXl77B4PbhclhTuDZPxGRRCTWaRZMrLS0J30RxbY35i2VACOaQKaVIwKgXLsQRJK
tNrYpS4CmwsnePcZ7nK0ADEfTeIUhEp9AA8/j+n2ixmOjW4K5jh2/A9+Oe+qPcfL
VALzVL4Z9Fz4eCmD42aQr5YMszYwKot84+PZo29DPaHKdXjbA+pEplLqB5Succap
OZBPy40lUV/4IHCNVTHehtxO1WRop6HELaX0lrfOiYptCqWKmHwBL5ZuqKdeUNmG
DQJph/7JZdPPsABIXqpj+Vg/jZPJdOxbXW/Jr/gVnSFssW4Z8rUOrEDjtT2rSlpK
GIgCxU4EcSnrG00QEr7rRgiYQNtiJK/g1SCcQT/ONJx6nsHyPLu43Snl0qZNm1vh
+QII+AGshuEskWSrBNBEBzpYbtJqMW4DKa3hQP2rCT2j64Z7uQtE8UKhTDiZkXqN
Ge6hyI0Y21Vb74EA8xvX0LDycdvLiknb5MlK1n/Y5JoBtrApGVOpQXnLm7ZfjpsA
Q8yc8w8im07EsJ27Gy+SwZR6YfFPYk/+yQljjmLnQYFYK7L3FvPC+cnYfPSELO6l
9a0OFEp0uIPOyhB4yN2/9pH0gY0AUo31nDhHC6Gsl4wbjJavqhFR0CfuugwVRRLG
En0EbLhYBxqG689aOQVnCTU2cnAq5Sb9e13R5ociwhKV7TFzSwlk/GRHZWcazTZG
leBBbdBwycr4JUv2eFDBFhLkMRoe04LpOeBmgpoe1r7EgSuUF7sVAtC70j06MWcl
HrCsoCYJijofmFmEfzoANaRbjLZiFrpBC5AiQNtkR7lP2BbMaPzr4mCr1vHeBENK
LjzramrnUJyUB5dtvG2Yt1Ixs7fvnksAHEHmV0s6n9z5tviWW7bcC1jtgcCgiFky
0Lu0lqc6B4B175cBu9B0rvzZCPPqpRMd94vmnMyLBHUhw7CwShvTrykf6u0LcDaA
42xmMgsTPvPhCFGa9acrOZVMPBP1poNytH4+vRs1+nxJTQXg+7efGYw/Ut/DL6UD
OfBTgIr1yx8kgQp4BDIxuY1qfEcWUm9bGOK7dpQHeNwR1m53vuaWZj1c081JiXSS
P9j0ASZT7ymbbmjjDVl6pjXc8GOznboEEEGn6AR4bhDGx2KNi7HlL8slx9BfSK2X
2XT1PdTwMb4/NRgT9OwUNRJPGwB9lVxUiFmf2WSUlltpo6TmW28NIShrsfnVGwx/
BwS24iDT3XwKKQWvwfEoFjjPf2Kq/Q2HLkzULkswKlgoXgATet57/aPU6TP6p3yW
Deshu2UTR9ETCPTqEqhFNvdIXl5MZzJf55ODT4zGlrzRZllG36aYV8PGOPdmxkbm
ARSaOQK4J10CbRlS3+PBkhXX4ArtdX+jS8zFDg7bF4NjVNczulB332u/vipKGnaF
rJaPUgie2PrGHGb2CfM0wM03vXfGhJpqef3+hOwlZ22zSVtFq0QTDWQevjaFgOXw
NW0l48L5KOz0rhMIRhQbH0Da4K5zPtypVKRfR42GwpoZg6NhyJJ0mc6uQFzpDiAP
2DvZkdZbmvuRDSJvZKFXgsP8x41FPag8wIqCQZPUtxRvC/nUzgBXx9rew5sQeOBd
HNbh+OT1cAe5PjeHrovoxQ==
`protect END_PROTECTED
