`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fwPON+fgBfcGVj9/+AyAUcF5c9T4Jzhui8uTrjJutImr5JbvZw9y92ARLCQ3vCT
si0HENmAN6r+Hdxl13G2C4cKZxKgc7sIdyXFk89pisO9in67a+rPLf47DBAsFToq
yHTkNgNV0/SHGBfhfps7M5IwlsQBZuN02kgUTBNBGhLUbTRFyfZpg2HjKCjWOrgH
ncP2JU34pxRcTTLtns2s7DvPbV0Wh07zqgsuqDxdR/3XTP0dSoNmaiLNAsQD9mRl
sNokOwEaW9Ao4Su0WBvNKnCD018mMsIjFJjoqJBnfTalhv8Kq6OX3WqsXK0ELIOv
RTDglg276KxQUI8sMp1uHNzX+YGCHYHYNcXWY6l7Hb68MeHzatCDqZdAT7kxwDaB
Azs0helwdM1Fmy+LB0hYgWN0e/Cp76joCcAWA1tUkCqo0AkNoPcs9CW5yQBc2yQC
LLpMaqeD78iuw9/kYnWhCrvC+xjE+5iAKhQGzBuRMWOHahdOErgtuf+WVIXPwTgA
tE38MS9/a1QV2AtHKcCx2dawo6wi8QG5DxEpuRKkFaJE9GcdtZP2mMAsQsLCpgfF
gcIf+IDVtvcPdN7pX0YxEJyaW2U9bAQC69W3PrEwDWWT0Gx7nVkWvk5u7amw5w06
Aa/zrGAthwnnSTZdCAJetbuJgKBz/olMJYurU898O7tWZw5K+m64KdqIDC6Tq7tO
+xQy+A8GyYB3eXJmLxelrYk0aGBfi0jOvz3a2J48K3i/KjAHROsFZe5ZI+JS6RNR
am4tOLDK2qhOJRPIhokdnaPcFOUz6VT2d1qg/MSMCoIiV6QQ+T5MSeLAkaEB5f1J
Oso6Sb8aJ4R5jRtGdcq3EZc7LUO0tH8x9fmWb7+qEiL26sIqjGKFBg/dECNxLNRn
UxNrPtQALxFWqChv8gHvCz6lQDb1SuK2JfTx9m5y5/I=
`protect END_PROTECTED
