`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/MUTHU4F65SiE3Dy8zsN9qeM5Wos6u/nPwhiQMj8ERvdQNC1HUgp2xmrWz8ewcR
R1OEbNoErijz6Hr65XFukPG+Io4hYpldKg4+qXNaSgRrAm4YE86DCMBLVsDkSo6P
7VrjlgG2xEB1/ob/qJFzOixgEMgy6ncBnfztxAn5JABO9xjPKfdiK0PVugIN09dI
kmwQujitceBLWlEtkTCNFQVhbTmUWQr3Ka2M3g2Mt/41iBnwzhcj4kpKJPqitd8m
hA4YjAkh4Kq13sGctbEMvJ3xb0gQ2CLLQ624+XW24paBNd1hhq1ny84CvoNzwNwI
Haq6BNmNQuoWDdB3ycwad7wzyIAcaeBoc6XUpjz0xyDk4U5N9P0xQ6ZsJ8rWfMYg
GMFEjOHkJyvsNaS2BslWs62mP9UvHPmBN6vqKWSqFBCqDNPtOBxZk9KG74SgXd3h
0f6BAGereajK/d4u7l/FcU4mSifGhf5CAh0ugRVr491vP7IeuS5m3kzivVXO2SS1
uMEDBvu9XVRKHD1oKttBEH5u3qYTCJ+MiXVU8+aa6ivc8wfQ8hh9z4Mo2Bp9h17M
MyzISBDlGG04+9aXJhvyPF3vXwI1twba9XpAklhirRVJMzNA/q9zeAdsYd5QURJr
`protect END_PROTECTED
