`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8yzIKilsWEPYqt0dN60HogXwuFO23wj8iiqSyT7W9623PGCkZ7DTz1E8D310xAbU
Ua76ChiM3DM8LuKynTpKaIUqaDySkuZYTp+px/x2XgOTscZKvGli7N1L/zzNcQil
ShkXb8Ozsh/sAGsD0YkjyqKd6UT3xt0y8WpPuN8Qlc7bOELWXyaEiSrjL72x6RJb
XSyoZkZy6MXLBGfdreCLDjSN6wcwsJIfliRZ/FcUmEHcAgFL36tXrvMLZl8V82T8
hMTPtmLF0fnstjtLk90v0lFR3rEdkrPCRooWeH0QHkpF0/esin3/h/hJeU07t85g
65UTP4XAQtloMfWTnLftiSI6cdEm6zVRIClzo5di7M5HBqVuHvaj0rqXq8agZ/tb
REU/fEU3vuDbdM0osTHcKlgBiRy7UDpW/evACIcT8vCnb108tuRgIcW2uC3vIqaf
4Yl//oYKLYptJe3kpjjS21TdLdk+RRNvMAyKhqv7MwBOpdWBPFaIohzn8z8F0r1I
eP9asI2zYW8jDO+KiYQxagbEc9grQxYlh3FlXiw+OXwiRXr3cTWAhAwGG3FXMj+r
8sIl1jAvlr2z/PxUqzy1eWvPI5vgzFYCxzwDwg5jhULne/B0upp06DTBIRlLx5nU
Tpn979+PW/IfdYlmOa2HEfsmLat5LddueyuJggIsT7FBB4nHr0zGKpVZh7O16k0F
eh/P6uPS+jev9MGFpdZmIEZCsRiYmHlStLNtRPuixdeD+Aac15cReLfm+JRI0y1Z
rCZEkyS1pjZQtHxCJuiw1uahKoe1Y3IzCwSlbgnYb2nJhvGuVFyBjY55AZ/5deb1
4J50SzUIIzpNK5LMAWhbOL3tXjXImFPHqzaqCkSs7cqwXOMG3MhBpNwXHVrGpvC3
ObxSDvkxUMc6cdD8XQExFNDDS8jlquPKMk9Q2w0nDDBRC+YdvWN9lUNyRgRXdFyT
aF6UwXYHXYH4Ow8Zqi4vo1Ulxti6Hp9BeW6Y20MXAvKIGgKQ/p5iWivUaduXsuWb
aTXfBUnFrPbVxxGu2cXlwSYn6qpAEfkGOqwtbQxmBP9BZ46veoLF4fpuHf4YB5Nc
brUXWcah3sqMtuIM5xCvYZoPaRVdN682FDUp5rW54iJBx1DYxTDh5Uy1yNeIsyk6
ayitI/Eg4T1a2QaJM27ZqLl1q//sYVTbbS03z1rokDge3pb7yb24mqD4DCXaHV+e
P65Hlp+oboFNXfSe03pBKunR6H+RB4Um1tdX8wSzQv9URzQeLPJMDdfhSnzIUeMa
7soXZBv6ktn3QP9s72ncBt+Oh+4upufHpXxhen7AeuPPtM7YCHeTE+xpSB/Pvqto
50mlvpNFg465Lh3PMzCaRRVrzhYfmr2I43JfzqUgTFlNAdWMuRTRqE82cd+MGUDx
E4qLonqjXRLuUMIFEudoZmhjo6BHd8WF2DyKPHxKKtLm0Mq8P4H50x89XfaOfOJs
siUVMWNQTtqmb1vw05Nf8ZWCTkMt0gwZGZQ6CDbbUMGoH46+NdmppWeNKVSKFJF4
6dEDn5QBT9nFSLfmwjcaYH2leXB90UQd/FpNlz7tYxkAc1U2lU0pHmpWTpP4Y/1g
AHsQCyeWQoH4FgFCH7WxRK70DnjDh1wWoTJ7trO0ofposYax9pdMI89cQJJCVD6t
uVUBpCrEcyyZHkmJqRG+XYVp27spov98YbyoqIEhVqmVUZZezYWtY4I9KphdiinK
g0AJXFfYCxCe0WgKeCOXOHW0FM6Pd1MHkxCmW1wcU63Dk3Y2h1g1VVjcUijHycvU
wxYTmAFjBE64rhAbz/CUeCMAu4Ai3xz51nMyYlhH/+LJBTdmvcBDgfiW0UwEF26E
ha6Ufw6N7uqc4MJUPjBsSvaCXumVPzPWs4wSUVLU2rUZcCT/N6yQaFHd0b4Y28WE
ndbvBq1lgihl2+83yY1d2XJDsU8k/sf5aODaxaxlBNT2me3+Faw0AGD3Lh4Pfx3k
cQlr/+bL0B/Lapdi6pOmSDx+vLw7EI2gEaFdZuviVXQjyyMGz2bkyXKewT3qXFBa
QwcJ2z30s7IVSc9U2VyfyBoUttP6N7TYVlFzUQ7xG/CWixs5LZXD02SNes6C1jjz
ZhJY5mQ1jiIs0t5Evg+rI5kiW6UJ4le+VeJn27/SCBLzsQ6KX6H/eICuHJDE9oVV
t3pOS2yJ2asH+ou4yS6VfxFLPq9WOSLuootgD+eBEahvBbHA58OhQVhpeYoUqKhA
ENs6zh1RDsY/jbr+5oX90Li/M3Iu/DieCInbYzs2PUjKTL8iGXPDBLd/sjjbS02A
bHVOwCTaf0rqs1kF2Ynhxmxbi/vsgUA1NQ6dp+aKpNiYPmJtAvX7eSVTa+mB1BGb
5hXHMn68Pi4i6pmAaJHcxmTCtZdlrBW1jB/xXNXTGXirH3/G2QXxfKjwowAV+4Sl
c8TMdGsYNdYMWenV5CypmKeHBov6nbUxd0MON9j6oXgVJ7vLREShDiqlzkUu8ZSY
ZAN92pSsdXgTh33ZNXbCW2FO8r7XrgCQU9LPJwe4tu4ZF0s7V3/UM/rEnJU7o+e7
EUJAX6aULf0vXEFPyDyHztkVlQRs/UBJIvc02gjT3yoCqU6oAPHg3eseBvuLy2G0
LQOSTpgv3eYynanCO3GTYQhw/NoSa2ubDC0lqjN0tsdhGp8k7owV35KKWgOPvB0O
7bGKGR8byTf+qlQHW5OZY5lIxSKO/i2vGFuRRaOmZ0GyW0mAuy+rpuHc0twLTpWR
2Ezjhq6qY4sDZaoe45AvN4qVi/Cu6p5H411lMtDw3pGdVjpEz0KN+1j92fy2/2uN
11JDz/nImw4FVvFCe+5l00y0qaepzywD74OICowgAcdfTxFl702chp9DXqQQsNcE
DFpnudekPPPpC9x7X3gv/xnqF/+LowMqiYzToZ4KmpcExn0vD0MjqwDAs1axOcL0
fYdKOoGKvlmotYjgnG3J8Gvrtcfj2EF5bVch2RCzbe+ZDVlAWIMg1IoYQHFiT7/+
m4qri4mVt265p1kRoCDsylGkbT+CTvmYNExmyFuFPLf5jyFNM9f4GNUCHJkSFG9I
tTC7ia5Kp/Cs0CS+8tKIy5l4INZc5w+OixBILWmx/RUC+CirS3OmKL02WLnwJKOW
BnPskQaZx7tl4ynWeZSuEG4/Wwc4C32SjbkNfU1sam9I0xF3RdpUBiNO85MnEZoN
22r9jtAbJILXhO15OB8BDvIs/i2MZWdo54ugZAkIGmzclKcErZ54OgdKwfrqheyc
VMWaldXABLNsCwjpQcz3NNxYwJ6Dltj30p57bBVToVl83jNEUlk8knJFefd53CTm
mOC2Cgme+cw6uA73o+wFDNNcskl0nhLpzThXhjp6TbLOncDoMHE2NgyLeAwIJ9F2
8ubVbW4/y//B+B9ioNvQhOcgvQheyD1SDSQNbe7/Io+l14hEZnxyOjIFU4p0Ps2f
7aHAiPNwTk5JqGoXX6pP2hFfBturO9Q/EPrO2Ycj8lOwemgRH/Nz7dOFK5drpvH0
wL33x3ttB4G/VCgmFzMMPuT2B2l6yDYN6W3KsePy0eklx2bM3R9jAq2phGxBIbPi
G8YqAAGUpBITfviPghquZrycFPTuPR52d5oCUKDaXmpReuQTQDTvE3h/hbt1vYJW
z1JVgrrHgJoQHBC32ppiBjRdbJnHgfdzN+YkBLv+2gft/+xBShHsVgNo3+hOzNUL
5P6V+BJwHevwNJ8F1C0eQnNcHnfYxRdr4X3sjt2YEZbQ3mU5qdWE0RvykAI4iy52
M2y/M42Rs9RoZlx3ljVmSS9aK4QbeXm7agY7TVlayaQZLfz5ZTME4FvlkaTZYaka
DnPGvcFvRV39BlL5QtkF4C7sk3SZ9mi/sAmmeKUdz3Ozwgd/7G/XwCgCVJlwVcn/
KcYd6DZGm7haLQes0+lZgQ9PYm4p61ICFQXJQaKlSgtY2biEcnTgx5XNbDpr8Hfo
Q0ONJwFIEHpQRdMQTPqcyw30T9rk9ZmCipxPPHchYyxPD3rdq5ZqNhluDgU0vmHA
ZdSALQcbfkqu1F5c2vl5fD/SgoCQ1/ZUOXEwV//YoUKOVvfojDvHl1KRX/L2hyO6
Ni1maSf97SBOmMYYWZYV9t/ESPyZJWSZYuG3lQvk7kCe2pnuOKbHd/RbiGQzDYRE
lkb02gqgqbWhZDbrJ/NhcqjwTAcBIaIc+5/MHy+IO3yEY3w9GqskA62jppMNUl3o
2lZkQdCgxyFI7a2CXHrBsnld1z6NgxwdYQ6/hQ6gCIpqFJXAdWJwAOB9myzBr1oS
D1BcwtZvZpkjixFgxMJ7EYD5QPVUeqtHj98kdjN1h/mnbPb8w5YLsK8o+58IZRBi
rozmnamNSnoJLDjnk54iKWs5vM3GHsNf3kQThkYOulQwVX0SToyut+Ks9Clq0HvH
f3BVTZY5JeWdMXq6KlbBltqR4Ilqxnsm/xDJEBMYoRPuDX9Ej7FEKh6Ab5AdTQS2
1FnXdMnn7XuAPYpqYLKEpA8XYACJ6RnM2lCPYXxHRK1vTRj7S6VyYz90DjODzeV1
fHHHVeJ2vRZWqSuvzgcluH6bBSQ88Bqu7TXKW7IN4fh1rkeDbEZbBrTClHSVICzt
3xwifVBU5Xc8aCXJ75tvwIFzQZCCJBPA81knUqwOEdXnV4HK1dbPQFD9je/c54MM
Ax3yCeQC7pDMR2Hg3j3hjthyoPX4t13GdM03Xo3VhAzl3q7cjFC8mdGqCepVvqEU
N7I8ja9j8VS8aT2qjEZseoQAIK+o6W9DoWzmPn2WSIMQAH2qCdI6mwBVTHEWywcY
/EH3yGnCwh1QVUOB+5KbTnmgU2wfmb9qmPkIT4We249iRETM1rtBccQHGkf4MXSY
djNLoIFNzIB6uo00LuDW31VzbnFdYfEfH1b9snp3GtCiQqNY6f+98MLY//1cf7Kx
ldazaU3GJ1qlYMkmpSLBeNiHwzG/aHXB9uJ2h7ymyJ+P4s51mUoFQku7BMv+WdGd
HTwh6B50+Dhk/MI/C6gveIsfvQy5G2PZ/prBtNI0hyUN+KhcIWqH3bxIPU8jitM6
9rzRXXPKA8mC913kaeoYSY2wa1U+86dNidCyGkPvVMdOfggGSZJoqxgXaOgJTejk
VSMWNrqDsg1NvopN4zTMBvkK/riQl+IEo+rxTzRNbua9AcKd4ilI23ToiThdQRSU
+RlbtKAnFaF0t37MkKnXRWLmj0XNxqeU3pDkZbjfoPOOm7ff4fCQDdwjKnQ55gel
tEK02+DKmYyE/bBPrqoCDVHQTQMJGW1zm2EqB9q4YP1uVjgJNgAX3fbLsNWJvrW1
OqjLoalgzc1O5kXehKseLXOwb4S2jrrf3Hm/LDYlt9IuWrDIu1+S4YqOspZRxUjw
LeC1e3ugP3BWpxs6SySNslHQlOsTAfbnkhiQK3stnOqJwkgyiydyCpeCnID1Gj+x
s9VKMo0Gmk4NFqOgjfiDsfBJios00ItIOm6FGCY8/h4CD8Vh+F9UcAFdjcS2RjO7
V80aIxoZtOErTWTlz31esB/K3jX8G3NEA8ktz5vCufQJ6MmzUrJmccva1NJjVJBH
O5YDxPJ2NdeyYlfAeYweEEeF7cpcoUu7WdBrcGML4yjC2gGS8aWrWEZkIVTTtEQx
R6g99nbLDEM9jRYemlmIIcw6NSan+SdCeskjOuTmaCP4884lIz3AdsvdHXx4Dm4K
HiPk8XKQE/yHV01QsFMpi2wn3Ha3Y2vJ9V0cYxWjGbgJHIORIXnGT1/xXLb3u6VF
Cu9gBwle6nKRxyRofhRHAb8eMV5k6EdkYW0CAXuiP/49yEQMcLmfqmBEpNSYyhEg
bhFtmDUfs2LV3Pjze0KtEmYhptjCa2Hv3JXH1pu633LoHvxYjgSR1LsD+ZZRirSi
kJyszbN8FvLfWXu2EpcrNVi1IBHNOpSFNveeu45KuwRGb94zXQ5OtUS0HA/vw8oT
rNMXcPP/7G/ys2eWU5Eim6ffCXbGHxvbL8hCdMSlCHI3dC5GutR7ajfgddhkMCzy
BelTgHDUu8eqHfTQV8pwgi8yYuYHSbAg+HD+46/oIzkMFyW3BudoSORcfyRtXUb6
hwr6PUDsqY8AMFTWNz/HPfsolKg2uv9p/24u4VzHCvK1qEuhCBk0ACKhPWM/6/Zu
99x53OLv6WuPj3Pj6b20Dk9TSuv1DHGnLgtKiYo15qYdCAgEHPoXL52lLLaj8T+4
45dK08DgdCdOAwke3zokOOuiw/kEK/wqPCjQmzoc2p1rk+6YFWGPvEu+2U7qcwdj
Cbi5ehAtNq6WlrPFDy7WRwnnS4sW0nT0HrJG0VRizlrj4oAq1/5SGAOv/LnfxWnG
tbLibVZbVxKSD+M9cRpDpbx+wwsICw2v+KvVK21dElM2y2ubF4vE9LvzET8BXFf8
g42EOoiEfC7tAwSsk75SzKkHYzXac88CRc+2huufwCL3UqRTnFfSH3wINTvGEAjs
EW8bLhWYmtzSbZztOWfRVOOc/5R8XWpqIgM56Wpe+I58q1F1mykzASLuVBQiLdJp
lc5VFP/BxEjv58AGFkcMBpM/cU3RAFtd0CmIgdwdTo/ZXWPmuMiNh6bxYKYmIpNk
UD9uok2YJC7hiMggfhkUznO5tpN9ILNiEhkimCZVqtOcC4CgE3FmBxdF5FL7fLUx
sLcLJp+QSGs2dhB7LnRfrPNZiO8BqvrnaqHAAmlrWFI9aWeXTcLIJPE+MfwbWVO1
aNATkeylH1+QtbmFbGR8yEPN5fhM5Q5NB8KZoXm9gZ+BhrBRhf1zts3kmn0X1Iss
c2HEAxekxZA28L39Na8ssqUIMLLJtvIu8HbEwVs+It9JQw3acurBc5lMmynkm/Rt
zO2KddQ8eg3j2V0Pxgd98/2emOoT6IZmkaObuKjMtFdNXpC/Ug+GD4gKOEARbyu5
QQdTQlvpdcDtTqU3cX4Cc3vkW94Z67mXYVRPf14t/rV0J47QBcyC6bOzR/tolClt
lOlvzwmUaoXBY9QSb7krSzbaQx78mWswEqrachEF1Utvs3/UponQCTUtuJQMKdha
TH+EHf18PFq1E7+TH1no8RCaxrRrS6TMBCq7rjPSYZSp+u1lSUjXsL5R3hVGlB7O
IAHu+Jj0zLQci6wpCQIAXEokaUZiCq8lG1UXO40qSG4dE1a9b222G3cM3RUYBj44
N/s5n5GRJim3cE0MlHPDIpWaGcP9PI/UJ6/4LHXEp1mAhZ/jXrHfor/d8C6nW/Gv
IhRgOFZCSUJn7y+370mfNHqZa3tl8scOiB1SWy5+3UG6dLd4MDQ1ImeMUfpu1jjt
P1tNFySmuc/2fMOpGfe/ALUXObFwFGY7O4LbWVmCIz82z4K5LSN9i+FGcDXUJ3jp
UR9IgAC0wTDEttvXhdQehzCNgKftyLtVV3qlkypahenKQd1zhJS0Qij/wQ1x5fsA
k8x1sFV3k94A0gnwjtGFNASbFwFaE40dHjly9wtOvzBDJ+wrCEJtU6B2MIOM7xk+
UcRQTMdCnN19wExnyr1ipKzC7IjWEgvWPQol/KEE0FjX3ysquYctaAc4Ik5dJ4fa
y9PyjHG8hhm8bII7RoLGSL5g4T2j4TazeR8+c9XAZ/itjupRHBi2Kx3sPwHivnQc
uz5Bl1tvRSHB0aGSqAQeLiEQXp/ucJV1eWTEhS+Hknv5JVfa+Hjgn9p/Y5ytIxwQ
5HI2q06P/+8Xeb055YiKQQYyLIgjKlhTevZQk3bzSSzBCgtVCKMutNfIMd1XrnnE
CQ6VPzhjUPhAKLpoeD9sRo8h9Cfmoeja2j+0XaGcK4Ges4n4dVS3zcYaboe91QF8
rZB8aRg4oYzSaxI4Ug4XT9H11vkz6sO1AZJaGwxETkE+iLSmCxExGMx/TEbAozJL
zY86cFkebeCK6dSfoAGpfXlN+Qbek8alClL2bxpbOpS9NkrkkMllqSDDOW843ZAe
o6CZFkM8QsJW/2xOw1wlCaA8DvWMcf1Ce9g0Xv3MLvEIrl2dXTcik2bbULIdWJ0d
YY+aa3GAIjIDn1BRwLMTscqe0ECfwIJgW/hcWhrHHGzFLnTkNG9Rm9X5ritkq/EZ
WavY/aWzjYadg0h2FQn26V3xO24ObqdmcqO4hjRcaT4VzXYEzUg152UbWQ7dJFUB
QZgtqnPszJvZj8ESaAehSjRoiF22FiBi/BfwygNnfPa+nYSvejCcWbKhY1ZaBKjO
rrCNCEIK6BEw458nNyT4cegdeiDxBmFEpKpoSq2pzSN170Qoi9mu3Phv6B/nDdpj
xS9o63hzRywX0fmsrw+CgwtHaEMsfmJx997GTo/WTJ6MCJntYKBNJeOmQwEuhvG1
qKIfYgri583JLZ45b0ALlV2UuvA/RIDSN/+BzffXcKwxrnpjgA7KOx2MkG9qS+Cp
1RrScjoa3PFN+4hTVDYi8s3mUvkOTncPCDQXVPJErRvkT0aRpbB6aLf/mf/d42Y+
+BSU3Rft0JoOuw8HWWtJYQlcDryYwAqrbs/y8oV+xD77ZofHVf7KdSoWF5mFtS25
Kn7p2KOasP3iZsr+kShaLfSrT7lr28F5C8fs5i0aTgxvIhJik/Y+TRRGbwB4qodN
6gIxZZNB/40di1G7M8/H+8OAkQwVdpUGoPZJQt3HvwEBEB2tNKvrqTTXxtlemeOE
CIqyRFnIrMGHocRQnomNvTZxC6mf8WCrNG1cfoIwyFxxHqIKTRIq/WTGd2Ph5u94
ZqZuHT9Do5ejYoQTAHyydKgmKO51634Zy6z5AEDhn5/TNoSOhcKkYiImyV6a4yGE
3YYKPgRgVOmZrdofPVlGZDSr+LPPNPkMN5OrU4fHEnuAy5EKblfQckRFbZTqOKvc
YT5Lcf4CrxjkKANiBF04MEwLxJy1oBbFYs9YCFxdnsfLnlfMuEJJQ3qkQDNyXdSz
aFsCpG8Px8wxjtHuIlg5yAeQW3KupJvRDZehF+J9kO1iw/eKH+ngSw05pz0atEJm
XuubBJWs/K+uTtBYP5KthYitivGzopxFf8v0/RxNMI+bfjlHglgFs2oYeiFxSjSJ
6/ZQLoOQBPorsMYj51OmtJ5ktG6ivfaGfD6yw/XGAmB+W2cTfvQRfr9XAPqYDtek
IqcNVBZFuB3a+RYmD7S4u8mQOmQh1yTr9NPMQ5TUFHnapV30diynKRVPxInOkQDs
7JyW5FRw8Ukm2axmuKMwJP25+q3AJvmwtnbyT9txAKF+d1IjA80dpe3DAMCqHAHv
We8S9d6rhxIN8VPD0aWRauStkUDBDJw0Va6pw0KmfB3bEB/fDz/Gn9pFV9ujz/as
kshrYer1ROsqICxxW74eKQiB3XwBXFwQ9bV8jAoxG85v6Rvpk2i/DFNTqhZnkIdl
eUdi/uGg3ID6w+aB0+F06cwOcEmBZiuLFWxQR7BTPI6vu6X2L1S+coBoceU4p5dO
DATwxanF/SXgS/NWpPRDW3o0z51nSXCnrFBGcSon1nUo1MZIdM60at9R4aHPzc5S
6cb8GQC7gbIE1lBLnuJHVHs6s9atbEPWy3UaW4Duz96IpFR8xT7IHfFiVODO+mvR
D/Y14pUfU6ccL/DT8ODO4b18Dp6MPvdzCtfImFkbdpNllWNlErDDbzFhEf4VbS8h
YT7a1WcdR4RuMhcWLk4uLvz/VvSM4ZjMnPg9kmWzymUrQOTrjwdHaN8PfkDgUbAE
7M/06wxP2OkkISoB8Mx5uUBbq11DY7FrX4LTyYIfZg0n5Z312QmnumwHwmiCFotY
/iGn2LT0/ZQRjtEzaos8uRBXXzbYs0WocGb1J/Dm7IY3i8eeKsciw1RTCV/xMPg5
geK/K1mhDrl6UQJKd9AwaDgxsU3xkotKTNsUu+2tkMWS9FzOV0xpNGlBv5usjPYx
WTrxrhcjjyjBRXlncVIhxyUQ0xj+qX1c/LRyKEV2ZdYcC48YsDiyHFRGpB5BDW17
9k5it88Zvp9CObSTIxlemmSE0gfNUVKnrUSL9v3MfazjJM5qocBGy/ii80zMBg7P
kgTROHqNwTuaxBtF5o9Y1Ltz2xo071tKxN/x934xUOitaVlake0pzxwbmE9TQu1Y
0ZuDksbg4jm39Q0tF9y0jMZ/jpcK4BlQWFyOBVyI0l77qIYztfs9tX2wrBRKhiK3
fLUrBXCuTlSqTDp/v6Kr+y+66Qp8WrVPI8yBsDw7eSso8rnHeSxP32mkdH+dcmuO
sLEe3vQ5+JqRcYe/rH+4aG3iXzTgZxuQ37WQr6Z/cDwlWG2vIWExT8DrQaHEsXwd
+BYC5sw5B9/8S/T74f+VOzMH/m6HhrQBDOm6R+hIeNJ+3l0yfRDjp9RFojUm4gQf
SWMsoHf9MnKBPeqPMz4Ow9A4VkjGCtiKIAoUrNzXN3FCVT+cV5HoQzTJ0mOHT2En
3ySYoZhCbgHaPsHSSepWl7EY3eoXOzTeenUZg47zF+eI1hcfa1BLWg6tlXQrziYH
lxeiSr7+r5vNoNg3mSGIGGsSMCioXEAlW6jY78DngSvCT0vAvcAuGhgUewkqsEu1
6nlCuWL4nIed4fVO+7MplTwBV4sJZTdD4QxsYkHLD9sU0dsAb/jH9dpq19OwKIJy
iO6u7VpWNYspcAs07yYYzMTM8qcrYjTEM/GKcVBhQsnmsyW3Gc0uKUI5lvKmxFVx
f5jUsMurlzguXL36JEJWYBZbD0INhLWO7yCf17pD1aepCs6Rv+PqQZwuJltJlLg5
bOQvBJjpQeL7S8B+aYpE4g1KYk5SwNaRW/nbFFpT+C+ZOPgruHr9RDL7RfN2TsFy
JIbf+W6+0CwvwLCBZ8kudq+mHNYEhjE4i4bEdaCz1fwjvQCmtD8Jxx6qkXLeiqPW
QgN6iJz09QJBC6ds1eNYFeRW0w7eofxIMziiKQ1SLK6XnuU9APRL3nfqEtvCuXU4
togVpO2h5xSNqGIy5GhwIqFWCHV8fKsyBBNurS0wc2Ls+VoAljc9rXwXxpr38G1S
JNZqH50yXzw6WmTLyaZAtaGahR9EvQIgorrN3SMH0AksOIHY6B2HsmEWTfBufxOE
C5HjGGAYCaPI1xuIRl9Ei5DXvElchcD0GDqU+1/K9az+qyuLeGuIjzM8KgX/8bAB
nRiT3b5yCAS0GEJYdDVoW3R7L77u53uqXjtCnqOZiGuTrHJACC6bsXxzpqpdsaCU
pRNgzqjwptOjttJIQfzPqh2OOOlKJgD2Y1Sm524M/Aam0xVO8fRt1A7cHtWXlfp+
zvnnUwk4Bqr0MUFFk4n3iUUmqtRNzJwoj8ckOmJo/cvb9/YciU///v4sZoOeh524
bucV+k8GQDIxJ98cBK6TVJh+A5imDDURO9P91VlvC7xxSMXey8hAGcCS/BO7MtNX
TG2iMx+BLimsoPleLgmYeK6DBx/gUkoc52EEOm2B8pc3edr/4n8OkwdIdzsFZBRp
9y7AxzCVYhiYmar9cp8J9M27JFCygoqipd7kAGsfoaF7LaYwUProCZIJRs7I0t0G
bjlv7nFLdeu4zk/cNagJEpm0cGhplNVBrwcltVF8ZcjCQDbXQgicNt4KHLl5+ntc
nYc82w7NljF0K7Qwy7GpsluLqxuGAgzjqeKtCTbLBEVOy5XUPFReU5/ghbnARQS1
pgBPL1GkiiTw6VH85s72S+n+1R8CCtilnLr6HvR5ZPFtnOft7QvQJw2neoQNJglq
nQ5PEegDsEvJyGALqYd08+b6Mw1Ub+w08Hpm1hvw7e0DUwn2N6ah4xaye35w0G+x
sWbRAIK13bmDM6wH82xYUGRTAvL4xWlyTQfZNQr/UM7wphv0BlBQsUF1JWiU5h/5
IkJuK+mcqO804qX5sVtZeXhFvTzHIzw23X/QAYJCw5lY/cS9NGZTvyX9XDqh/5JM
m8NDsDj6gZOLGxNjif7NbOEcK3XeoMWAeRksw/azD43VkZH+bKi7jO1UpDi72N++
DqK7X28RXpUa4Jajyxz3fgDY9liJNBk190RwjdyIfkH7C2/IvUVFP7UvW4yT9EUV
TgxbAZ8PHHnH+o3vRnptnJr1vEx3NveikfSGR9ZN+vHKFm3o7WhXRTl6gvRcIVoD
EWXTcDEoB0tOI9K07ngGJC50KK67QYKKiCEl47ZU2cUg/YzZYwi3GJYpIYiaQjR8
/YsU4M1x786YzAt8LY9QSl/p6Nm6Z1NvV0d+33K/aT5Fkvav4ZKvzH9jcazUwtdX
THZYBEycwrExYfqVUXPy4oR1qHJEHcKTH/H6/2S3e0LIwxOJgDwfUwsV8oBLki1d
hKUcGBL3ln/MbL5YZR9paBnBkvFw1lIVY4g45f6zh25JuoBawVmqB8m7yvnkvj6X
d0mF2cx4V63og7cjlsJKRislJQ0lqlCyQcY1d6nkad9Z/0GtV/Tj2Eif5xARFBJn
rJUslA+a9Bb4/jWMyguF8SflfL3md4j+zf5S98lsjnTxPI46kdXn0FA7pbF1pv3q
JDW9OjEGbzIcCQf3N+fBzPID4RHDzLj4mP6a0Alma7aTAZ39ZcrYbPUVr0u2Vg4v
KKl2ly+Rb6Rj7vEY1fTLmWnhIm/gcxc0cTdMksZqgJ1dY2cAUbzl/YCbvsYUJFAa
xj/C+wCQ204QTVWmqvCiEr2gi6iByOjHcohFsU/UkHHOyed9nlV+gns3sbeYB2Za
6SU52D6GfXQsM9hRFtlLG7sRXJw2B8XKil4rrJ8oWV/Ish4gtbOP3ugAquelJZmS
fnbZjlIByF8kUzV/xtLaiulngske7T+RhE1BX09SHyHXHuqFZpWsbzEqZY8Dh08A
UMZFkHWaRkfqkG2GKJoFIJsZlKw54E8yDJUpovtodQnTxLYFfS/4s4TwKRgSp2PN
OaLXhkuCggDVqksimV+4LMEP8ef75AtL5LhYiGVeM/VuWqzazMXeJwpO0mvNJ4oz
UHXV0Mc0nMd8UhJlAlGpKXFVPPukn0LzaCkBqOvIfNhvfh9BHVq6Jc9vYuEtpCxf
GdIpRQN4uvg2rkXBAvIAcNuY6TnrS9+TqqlAqI3bv/MyloH+30O0bwyQkIfD6Nki
zdPSGHa9ln0z4zjZtDjRjXBcixzLOv8W8sCs6fEFsNloMPGWwSJcmFcxIt3QKalQ
yTLd2KyqH3BAa9eGDek9gdeXpxpFo6+VIkbssvdwyL3T0SLF9Ho+fWGF+qzk1V5k
VhAUGnxszFbyYVa2Kmm8lNH0aQ6m9jGChzoSVXQWC87bMoSVJSIKyNzEdYLTvX4C
ikotlUIpfV5YbPJoB0pCH8IAKhpg6TbYvhGUtsrC7L8hVrg4Nw58OiE8ddAXDiKO
/HrX0/G0H9NA47Z6BgXKKzIQNawNUe9SZZK4VOiOoBMMjyxEnQo3sbD2JeLvdNlb
opi7ULPH4D9ZtHDNnoJVBHMoWZx8mdtELZ8jOFzdy5NcxfAJsDRf8XWRHlGBHWrh
wJ1Mo/kCiTpjEBH7DC2fuhlFCJ75cgxc9ZYtYn0OrF0GC9rXsCiF8fi+08Bly+J4
5RY2zeQxXAIK9cCO5+A+gRxBzg9VfQtSzIYl5ex0VLHmrKCl4z7mLUC2A6BRqi7A
2PMPpML8gtviaiqd4h/baxW/H3+r3g/TxnD22DygAYa6qaBSxQF5cpB3S+/1fp4r
bAeSFW23/UAAHzwDuPygOuMtVMhOASsRpRT14rDsELncWHcMO8XLC0yZPvCcHk0c
v93zhF+AWHNfB3zjdU9PJa5GfXZvggxt4tTOceWw+Olu6OKfnKD2sW0sRRqcXBdK
D9fc4iDRs8JTtr2GkFkq5jZfIAG3+l97mta4Hu7DtwtTR9DIvgvwS3TLkipMwMhj
dNuwPtyVldvOYf1jHY7oRvp1q7RqCFWVXjS8uVFU8S71QNw9a2JJyBCk8mVoXbTL
8NbSD3okKJeNgZ/5CSKgmye3T3WbcoVPsilmxGRnlsOeSJH4zCIYXYjVeXKc7o/u
ZIDZ8XNnIxIQXkZnZr1c0CV4z1nzoEW5Q0AWtxz4f5OTt0pnxLW1r/fMaiECGPw+
kVXsCizGqla9nLJ1mjsx+QYSZtsTUfFXjlw+N9LjH5fLIH7FqtL5Bb/4UmNWUmYT
OvpVxlsa2+uZ1gpRlIRuuTBiGQNt3x9VyPfcOVbPKXrJ9aH2lsUEAxOlP+4i6hOx
v/RYOJAasYfDWG6336FTjLV+u02Z/oJ69TynXIgbuGDzVrdy28EiTqEe6yZUjd5D
EGtlTq848Yz6RFWXiRg4AIaTArSp32fO304mmcDooQBXAfcsElAKwivFN4KTjrrD
VIbw0SboEkktJKY2BfAZHSnw+6gPit8RAHYWAp9coy5GtJH0zv2XA6rpOdEawDd4
usE1E5eH/N9dduKUxDVYiYffIg8iIXcQ/gUZJF1nLccW2kEOw7rPHYnoMh/OwAmg
+ZU0W5pwTtV9U4AhORrXrzfunsXEFN0wk94bl9kFfcyS6Vto1sZKbjJoWoPI0HxA
Hz248cMJ19ls4Fd44rH3+PuNGLiYPQy0HVVuGpDSZBEM0prTr+ZYzOKprtAi1gp0
+RnbBVtCDyORmP5260q8+ex0YCn/thHQe/aZ2m8mmLJJRLO8N5+zpozhb8mPoEgZ
sCWJS7z1TDb/AeJeVzgd+gJxFU4gu5+f8zc25PHY7iA8X5m9V1P+er0/89t8/oXN
D6BvlQSuCjEebYWeBpzZ/tI2zGV3ibeh+5zI/uxLX2n/zp6iGn50MzwpMQRumLop
0pSnYcb6C8Hfgy7bibQhX7VDTCfkEbRHULAM3uRGHO87z3s53q0nv+wm6jSkWTnV
BYE6S/XlOK+5eDS5IFgGt0YwI/8d03JTN7qLHGx9xZxLhPfmvdMT3Cqxj0dgKbZw
10viAFVRh3Xcssi17Hp8BX4vaWgLDo1MY2ulHGFsknSozS6SJ4xI4eE0zjxZbNht
1HzaByYpE+KqpD5PMnQkzChGHeJ4nb79uDh4co2kwSQPsd4/Xpp7Qh6LK7Er/O8K
efkGIPujGZk2of1UKh1qS6vLEcsjE9bp7W+IPy6EHFY7/83j4C/nm9X5gooPnHZ5
VIza7HFZgPI8JVydmMBIZvx63WqHRkjoeaWJbDzyjYhDs/OYRIs6byYwH77mfeWv
9lnXhxczPab1k6ynmdfQwfrsnXJNoJ4UVuMbESJRhAquKJ6z3us4zOLsrFegB/xQ
uio+3ihJnUzGzu6P9dGV+UacVmxPERvQIsRQsR2jLa9wj8KeHNtjJe7fhUhWKYYB
8DCGDB2OzrM1TCHAl45fZWiaJ8hYQSF032GSUNuV47pc7aWTrkVQX/XQUHmI/FZ3
fHd/q98/CjWhY/Sh6Nha3fOt67GzszEr8DusvdK3xE7IytJDCSv0XwwmTw/LK7r2
t+gMenE2Pq+F0PedahtUfYarKtNF1HXJbI96Wjke8evGURXgAwVpx447TmgCdYQ3
GXQZ1ameX2F2K8G0wrdUgJK4mO247UA46OtBJbPOg5mYdNc7q4FokdQYgKnfzAVu
KxdRN3JH3GRvZpgxA7hLYzhY//lpqoLJbDn+PM81nhA=
`protect END_PROTECTED
