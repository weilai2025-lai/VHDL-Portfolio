`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRn2bHHNEgk3mJHWdu4p8jVtI6u38xg0CEoqgZlXJoN2sufzpEzGtF46o81RdbAj
gkT6qRcAd6Mpcsg6N+XC/bq0o9l0yzz5wFUn53saaa63dI85vme301tGDO4ofaKl
dskzbYxHCTrR3h72kFpqCopex7kVjbQ/hIaLLU3MINUzp7aP7uk7kNjl06kfm/H6
b7m5QyMo61m5JyolGiaHUc4SUSyEH81kKbnDTk9QotsnLxdGMBClqYJ34Nr/sJhd
Mw5RGZN5xPcj8oKe4/HyNFAoImiXT84dthJl0UNyOxL4R88m/Br1sr1wiSdQDzWg
BhX4Lokflt5a/tmfrDmYjCEIK/vCekjzqyHVqwAGflECNGkqdY8xqLTlJcpkgrKh
c/Di6JK5N1+snBQYS/F+HuxS1Ue4UBDb2hnofysyBxxtUNFzZvak+sDy7ULmBW80
J/qEwaZkTj7+5O9KEJBCxyyRpU+PHzS2jRT4vSHzcLGdLlwZm584eUMT94s/qX6C
dl6dvll/gBgYpF+nPOObELRO7nUxXTAbhAVgk44Vjf2HSq+jazBygXjpuoSYcRp0
wBCF5dgpslIrkZYUlMr7zHNrsPRArs+0qWVYLm3RfTb4xkj9B9ucZpLmLrl1weN2
fTcMd6OAruoICkl0k0sNj7b7Km088P7lKiQk+2erMr3e352zpBg+aq2rCkcQkdZ1
g64SHSYAEhjP9KVfQv+2bLjH5IiUkgYmQWn0Pe1q/gmx8D1BOIja/xngp4yoUEcO
jkeYDFA7dVN/seLkF2tZKOyV1Id4LyPP476cUMSIJPyIh4+eH1HCQ9+pZWlCabez
UR8T8Ubt9ylEhtT8BsWRG0BHSOpG6wbVfQ68BAyR2OoJpR7+973JaEWr9Ldzyoea
R1pqFvmwQ9DCcMovMDfnA/ViGdwzdfhlfAptUcrBseecKw6DJ1M4lB+svoWI6JBS
FVdqPNjFPUGyBxXLuJZm6mtmPJz9EGZBpHIOTdinSqxyma1+kL3XDx7r7HH5XN2a
a2cx12kdJke7ikWBekhN5KoH3GLBFzRP+1Isu4eaZLO3EWzGy795EjFVIkv+g8Mr
op0MDpoCWgds2k7XzDd3ooK4Ps6wEUoLHjxaYRM+5N3ywf2eYRbDKZzVd7vote/d
m/5qAYmcpb85njtMx2PskZic+bel1VX6HvRYudjOcQKBTaB2h1rw+/TdMwlPkTGc
pQHZX+gALluoX9ltxSVZPHEjX3DeNY3b5HpRH/1My6rMadHEuMfgssZH+oCEERmF
cY4q8iyii9HgCfqZ6NGpxbSRdhIxfqypPUfTsbVVVKX5b82hq24WHbYHQaREQz3M
UPK+KBS28xymG6s6PUyPWtn4cOJdcR4uljiJ3THtwPlcHvBNH/CfjHBAquhiJxvM
/aBe0NSVsz4JXErah3WmEh69LcEGE6/PcTBDtQdIYPaeHyna0vhJPh/8W25kAvzv
yiBQlzrxfBE8WeXpCmZlQahtmwJMqnpztG1zgxH9ArVPeK+rjFOHKfJv0tBLu8vK
SliQfQISwXN0Wwyy4lqJQcDSSgDf2apIqh1duUQOfbHaNQoctRnUt83+f4+RuDCG
Q4ud1FHk8ADF3QJpVdQS5yrarFcHMW0o2snHlftBg0aEU4o3vCMOyyjs0mTtWqVd
BWeP7P5QluG92pBDESeO9exQ2yP7R8rZYfBJJ09asSaWYXpf5OoSHJMol8iPnnr7
+9NDI8UBQ0Zt/63R2J2sT0yyPkO7Q9si1zNufv3zhNIGt+OUy0Oil1FaKdTPKQhe
CUC1lke9+qlrZqV27MZw+ECq9WukHAiKJHqZiSaOXGF2DhEfCKRoxRq0FCy9nZwY
j/Xg2UM0J6mvEtALEis1KWZrrUegka2Oc6y51B5bT5/sj0fiDytzBjpYltAax9Yr
H0G/8MFkP8znIEcozBjt5laVZ37to6XVKVUz7DGmSsMBs5R9QDAL0AqiyC9UmZ15
Ifv2CTzAEWsqJ8yzi9f8P0wFRMs+jfsoQ/npUBy6izwC2b5eBjqaiwYmrHp5q2bY
ASrn++6L8Ap1g5RksdWI47+f74s7nWljPNTvB5jsSJl38FcwvQLR5logvv9YbYvI
5Fv4+2z85X7fjhurcQb8KzLZXSxU33XCJzzPTml8axYH6naYzcc3FyN83/gzjzMR
9jKEp//Ed0Yun8PhBSsZnUolNDdCBiDO0nI6z2Qk4N/PlqMZBLF45bkWsfC6mJ45
FCM8ZWVb/RQqhaLaaPO80SJJXfe4lvwld7/vaeDecpr8vFW3a4JT9n9hejYQTbjG
h2m0JWbm+YtEBFxExIq6JTVYago4TCjpEw0zO/3049vQvdASDufH5FNWZUQnW8RX
IAjDNHWvWKdm4PTqNGgU8RkoP5sGKtaxUcPBDBupppHAEz6WlInnTaEbyO+SxybW
UDw0L3a+PPvdNz6maBnKvYx+DwGYJcKOCnpWd1JOqp9TJg+8LhOk49hCOY2KO5E5
8hPyqeNLwtp6Xg4w+5tjOlw/bRz7rCXjlJc+xJs2+rnpCQDXUGpErm/RXPtZUr9a
XUA6CssAQNxAdPXh2gbqs1Vm+NuwFkYZPWBKXGW8p3oKAxI7Euufl8Mv3w+1I2RD
n+FN0ASRLtTqt10GEbIibeo3GxfeHA6x6vyx5+vuSKXw1zzN+13sy0HRjwUVu5kl
/IXErG9NBcgS9qhskagTCGtSyfo3k43LenbL9WYQVA+vA+iUgHC1Jv1aKtEsKONH
mwatexBwAIZ3q1HsNLFIta/8keJ7oMWQQBXx0SzS+PEdpff8gcpCzsiYsaVFLcZQ
wgWLMRL1e7f42Ghi+XE4FwMdqZZAgdPyJ8s1OfwS53vWa2dTLe6fFAZ/e1oXnvcU
7w9DZ61nIRF1u3gy3W3QbId5mKljwhpwr3vTnFqV/80Hn/NK6lTTHqmHALG5vo0d
xAYKphPnzywkSza42wSSoddWfMA/wXyKYPxhuINpEKl0MMoAVsFyE9Hjs/67Mki8
8gDs9h5kEzKSyG2gwdz/jLMS+PKMCD10hfji07WTUAnFMBrpQaybUP5JPGJG8rLv
J/GiYQYr14xxykKomyRcZkly3dBGEiyKkcgNV3g+tnyFUrCFkrYqYudqJIEPszdR
yOaop3aR0JNVHUDa4zYIUBUbkowt9VkIUPWm2prbUrY4NZmGL6OETUAGGSi6LsYv
FYIgcSRgk6SFm9daTxg6r7bFMxswiZYnZ0hsjIOglrdbsDZbYAtxyK+HSPbbPIax
md/3gPLWGquGzgTt7yYvj4m97CEiX24iQiS33EZj5VTY8mcWrgVFsicf/+MdO5NF
89pvMjjehnbnIwHwv5ctV3ul2kA7jBvkfchUFxCm/4L1wjgk93jg+raNZuLsX2sr
Aoj30CVdvKUdDbvZTP5yuGjjKV4AwZ4utGP+b+GrvfS7QqiI0tVJxMKvsyJV6+nT
Lf5cKBFDxbxjzUEVwIsVGjK/Q3XpLGRDlEkrsUjCSL26MgCrp1Iaz/X3ev1R0fgv
S10ZCsOC4bo6qnLV0GLwk7KYqpIGdLvv6rQgQdnMLa+u9hmApoI/wTTSi4orGluW
M1W6u5f6cW/QwCCB4DeBaFfF1+rDmhJzRAQRhc5/ES6Qt3oBqW0kzwDwgAWNIBeg
1q5DgKclfOxoNttL+hR7SzQxJTSUVDz2HH4J3IYN6jqrFvoTsMqBD1upmtPGAkOj
wDIsYx694CRzrXxS+6GOKobKxLMLVgDRJatnedE+kGkcxQG6h7htr2OEA7lABnyY
/pNwE62y4/3RmJF14eNXVGu7AeJKV+aW2HoNr/xpglX3IqTub2mbTnuLvvYE67iA
BdTpeOSaS70qoXe58Eqww9Pqe/VnhfGn9cwi3bEXHmlim63wnkkgjkrnGAMc4LPb
/wrPJgzFTLxPYIfkcZfhCuhEyIoeM5WS7c7IRXb3W2r4hIWrJ4Br5K/KUgm/z/Lw
jLgPUteYFqRVxV/xNhsnKqSF/SUdf8p5rPW9SrkItIhazB7J7wk01AAovLl2vKkT
usXJeEwor1nQjDnBPh1eAlOKUckZkIdxlR3Dt/sRvU6i1m0PFMmel/osUVgPbSDc
SqClsXTrLbtNqlIVHJO98AIlj4oOe3QZAbCX0cV43+qoJSG15RAde3Flvieua33g
YoqXEQXTt/8LoKaOP6HpxCw8QXvBaZPbGQIJbJeTBPKNdDzzC1Maagk2oC5q4rCD
D0ZciQSIT8Abz7FSkOVnGgmlhSutFjAFZM7NqZU9uiX7OaD55ESu85LItS5c6jSW
N7zxn+5ZXXnRAgh8yxM+JiS9+/9Z9tEmSn8Coz7xAVr7eH+mCRffIZ67jqnX+v7N
WNH6YhOlX0Mx16wZeEZakqw91IrLeDn56zhA+LHhloIYKccBv8e1wLTBDtVGSgNQ
75QXzub2jItpxvyX3TqhhbgkxyA8anjcLIrU0xaID0wMBKVFgGmXyZ8qRJZe65UO
C73zEy1JuNcn78PsfComWks00umc/fIEaIkEhY068v2J/Niw/nOEGDN423OPHEXV
6z5I3NuZGSbIC/UfLeG/MIs2aF+vWM3QSvCzx+ZVjXd+kkLwn6XCYFooskGcLN1p
0AEVjuXKhS9GkRyGjXvQhHLx6WhXm6/fp1lpCiuZD/VI926bpEvEXYhm6VmApfAn
HGXsgcKEI82MXVYrL2VUM8QlHgtSWykxpOGFgk2oUU3+20bnoWQAePU7dxWERaEY
vnrKJIg1sAg/Wu2abCvdZlCncvTvLdpF2xG7KhjFH4+F5PKMJFx7+N5hVZaqn+An
qXBY+KiaS1Pa2660mPuOe3Vl1tMnF2n6IjPs34X62mIUX3JS1BQLhj+Au+KvjceJ
ONkslXtYZjLFWI8Nw0o35CF+IyW9sBRVx+fTbC8+VJqkHbRvmnJBqx9eXUMrw3iS
3kBqHb2ple3V4dlbfQ6cvjVuj0PnlG15qKPzd0YejL9dh2fSvjB091vrpiOadtxj
a4piibXkxitdFagWXk+l6wWqvCI7tDyrEo6YuRoxsjtdNXnIrt0ahJ8eReWLzNlh
AQ7pL88yjz+IrpCImuSyg4usDgtYe/z3l5hAYBwbeLQ9Lrxon9x/EmrlSi9LZjJT
TcX+TbXFprJCcpcQYGqAsTwCh/EoSB9u15GylHlwy0yJ6SkvzkBpkSVxZCrKexv1
okljFkH3N8ploxW75Qk3ruK8+Txu6kP5O/ilvokqjcvVuPo2bmbbqpApQ9eLXPW6
gKPHbuqBIRQImvHaVtkfy8zxFITupPLAlT9KmoWrzDzgLucYBcbSMMX23hozmo+q
ahwdYFv93VkthfpajfVity0WcFhAhYcrAc8xtpfbVJ6F/9IFZSJqwRNaGUXLS4Mf
EA9GgRLAj7ZUyU/mrUCILPV8VlP6SARh+V4u5vKbafOwk8JRvGDNUYTCZaIjMnXz
w2h1KfEGBF8h7ip1PaSwgA2T+hNpYUauj9dmvi4CmazeJKqwUTjagYwkyLOlXxiq
I4DJNhaO2EndWMmugHth0WZLN31P0BkRO4t5oh8mFQwdiM9+Z/8ANcDMxOgL/LK7
tf2ClikvsEVQ3ssvA8wkr6GpB1u0EfhGNdvVOp2F5Ir8ysQ9/2okzAeysCZp4VXR
pXbSsAUGqocBBPoiuzlEikLpoYAUzFKizs0O5FxoDw7IqK303Z8bZgTMtiHBgjHw
caoLbk/1xxOCKxjtqIeYZA/DwMiV2B/VTvnNzLklT/AqoSCDD360EPBmz3LPlWFm
9DSs7JGpYXJ+VGhPBqLQaLQ3gZh8OASIREZG7uGRyBUw05RQviTPLXgG3rRPbZms
lXyKTX2rNQE9kT7Ou4TY5admJZjTsVPG9uoIm/+7f+QElcA/LTjNLPifyrfK0r3X
yIrG6z7yDpcmTK7eEfYAXyaMifMI9Y7ZJ5vmMz6+ChTYvEE63l0zhDyvZ5OunW+m
mRN831UAeC+B/ESKuViQN+c1i2Q8N+3m8wM8j2kbDl0QNxj9TSbqgOKxnUQwyqse
mR8rZZYohjMpogtJ5QLfj4H1NGl6XGo0BmmdyC3L5KUdvK/TQ7wJjXhs2MfSizW3
if3w0xUB8QwfWGh/mBSAiKPZPU8ZByLGeIetmPWm5PxeLp/Hj+A7glKadfZCrGNM
rR1gdMy7NwxOkRiCvYBxA+qsOuveMoVWXo0vECKNJt2NIxnWIRcG5UvEYzokVfxL
+KtNRq9VD/H4Mj7thGujhbyHpaNbKKakQiRh2TyGI5GXIc18lALtrup3XjLevMc+
16TM/GjchDmv0QAsc3r64j6n2lDXpHYY/hHg78TE3I8vqijZkqcDNEoiQ7hu6ZGN
bzKnM6/0KfcUMfJyEzMcVxi+9lf3DEdwhu+RlOPn5GZojU7NqXuzLLhGgp0y3WAb
85BoLvY2sFIHdnwplOxAZmLPVWv2Osm4lUmD2LjpIe9jHqemB5MyAeC90ZFfbn87
sf5r89dZiZs7B8hzMkJv082PBprOMfeZP61qGVYxzZcycoHc0fsp4T1bNWuJ894p
GFBlLrF77znNY7cdirNTRGpgUJrr3bU1GwGqYsrwsF4yR+Eoy3yBUO7MvOhAy7CA
FeH4PuGRud8SITbqL7SZALVLEBwKcWakAvDZvP9Y/GTyW1W7qJlryByfOzU3Vwi4
G4IoPFGn5lOfmadw7LeskPHWWLiaSWmcS/torg+qkNN40osneBra5TRKxEN1sQ0y
aaTRp9Nw4rrlBtapzJEXjtsuWfkoUhybu90N4uuoAeoMwqzAfWrqKAEplZ9GCP15
QAEdx7GYpaL+pzmYmFwmggXQNRXJxa1QJx0vMfkhWjYaqSF3LZFDifHgHldGcjSz
IHq+uG7L0XxjAkAOfamQ8tk7K3FhzsQrwaugiqNqH2d4WTaQEOcyJllksd2lHahW
HL1/EmyRr0wBWwtWVd/TRBPlPJnjWdjiOpZnZxR7ZTYbRUEiVZPsv+Un+0FF4UhL
8aj0f+K6xMqFPWdjW+Z8PB+eP4+wUFkuCTmZs3lDKIH9XK5cc7+NVR2JOh0YIwTy
/l8u+C5tVc1w05wr2cAHiMABR6bV113FYL7j7ZRjCrRsc96JFJ5GUBVqQ8PXbl+H
seyloDyobYxXNNDtLqXgEAaPa4LhCNCfS0NTnwONWBfQCYAP45aSgf8WWpphfLEm
lYJqNq2x3wtICrxRBvrQ9HAZbC0FxgvvR2J/2wdmpjAFb2X53F4Ym5sKUw3MXPeG
q22teKkJxco321MCAbZrPOG7OvgcjDqspkw0dlvI+p0q2F92X85o62wukmBtooTw
mfIj4MQppBUVQ73EXEthnT1VujZ2FHEEq0PmbDHQo0+Viq62Gwyw/59u3fjcbngZ
+60+8JTcXIpcMqF7J281ScP73/hYJp47LhEXzJWz48a3AxVr0tF1uLAKYQt7eSBA
/TQRJmDiCaP7ABMuVZbnzDd10qhDGKaHO9nJKRxWauE+RcHtiWWDUxpmq2AMNNGa
2fWn5+asyy5X0kRr5BmDaJQM80gbnJ8ureM33wUSNAv3Hneo+DEP1aYwvHvgY6YI
bAZ/q3wedQLsUz65qqVyTKBBjrFMQN30fEVcdG0OPdNENsomhv7smp7LXbkkciwd
rjqx7GUlSN9rHX1aZUZpOmL5lII1gD8vgNG1Bm52ONjTWuCPZ/PwtEDPStMNC105
t4fuHqDXWYytt6qjmijnWXF4YboaiIOc7me3dObRK9V8XZSNcNz/jkcdWcB4s4eA
m3mLxmLFJ/1iEw+QghjoivDuBh4tVqu8kQA8+Ci0zV0vtZr1olDLiQoVFdIohj57
HJu6oDnuuLw2kmv89dJQJD1WgI+8BB1hacfinqHkMMjeEqdM6yyEj5z+nqcFjdvM
LXGLSV0hU3+HCnt37qmzd3zo89sI3PsE5+gTb/df2fx/5jYOI3A/KSUg/jlcsWiK
73UW/BuHfEpoMKbPUDKd+A8QbTv93hchhvJpmX3Wdw7UzoHNfIhAdiyGwNxerYZH
TSM62CMpJ483snNP2/tzB9rmL0fr6h2y4DeZcXyBz0PT2aqXUGIlWzS3S5TmQc84
XgMSLLu+RWZ1P6BixsW9j9J1TrCdNDLP0onTrVBkfUBFp0LfRYtJsE1xCTx0kP4Z
jXK6Zvf2rO/6ijHs3EvDErCbOFgjQt5FusMJAfAjQimh9u52CzLhhUVF17sKivHx
gBBl91bbVddf6kdG0Dfr6uqoO8u6bgS3kGL5YOODNF87RBrURqCz5AyVb3GR6NpW
UIsRdg1s3eXLhh+8WW/COjOlox901vnZy7RRWhNoxHGknYpgGIwXQFgYn6M1jKIb
ngKJxuJTsaV/c4RCvgl4nl2uKrYDxQqWtgzL3oQCxHhv08NiXcQwBLzSe6EVxrV2
80h35+S98d41NrvSFjnnLLizLnmukjmyNDDHDYUKUutlsIMb/NTuW3MSCHeZUx8h
/6cxVAQeoTnQhp07YdDP6TNqjkAo/zdJo1zSEpgl/AiSzw2aE4GkNMb3sNMa2Hpe
AeQHNItUb8avJuxv6WDIjmzywtsas/dPHH28Y2i9ntxdgW+Pm/2BL/YKBbI8X2dH
qUb0hAwlqIrh8xURQnfhDCJ230tBUCZN8A+03Sy136p68kBGiYHxJvtP+cSwRjdU
me0+RQCIGcSUkSk7xyC2KgDhXwoi7c/br8BOqOfDIcnAfKHYkwrTIzr+Fvy+EhCa
TiN1d/EaSO8rE2P87tk2cWNkRJLX3xQB7XkVJMcsTh+gONU2Nr9ioSZo22bDicgZ
4DGx7cbK7F4b/pBamFqPdkI73VeMfvsyNOWE8QieWgKV81U6QiYZsNUhgTl68ZPE
qSmBSQWpdpzZOij8e4EWQJAu1XXGarCyCKnDcoKcVe3Yu9saPE76O+mrTIvNEPaZ
fOpRF9eoxrn8Z/W0JiJKGcE37BaUEWbH9C7setO5fpkvKf+oATyT78XCC/srfFy7
PO22uHgMa+qTl/34JRH0p4TJyFUhIb1ykU8ZRmbffe2hq74v4CwQ1TRUiHD0wx9U
x9pq8cx+ZUV8ziX3cbtGk89hFZHAIX3d/4teBbXOTX9M+BKdjXkhg+KsdHlj6t+y
G4YIZ4WeulqyWfgnpJscw7Z0tm4KcHgkcpBcer0F8aeI/2F+0Xtl2VwYprzo1Vws
E7RmpaMxaJmbB6U/lzHF/W8O/+z6cwoalrBn4oymPDoCJZm18dCNTN0kYVbixy+j
OZrFi2DizlDptbVpdRxLtqRykMgQDrClZ04bQfkZRyiD6+5Tz2yHNSiMe8UNXgHZ
5C26B8HJ++1AzsnnTViuisSojL6DBtmrKhN74ICM88rHvS+spZ7hPY6/Oqu5lymb
X/ZtMidDMlu6Or6GeKnIHatfJlx0qpiz/XgtL18N+jdaJ38esQNEhXmjH5sOYAAb
S7wECBm332RHveuNrXsRjIE/MyFWLt/qQklQLHQJjSLRvZA4vzfMdLjpeBHc2v8Z
WCx8GmQUG2Hq2CiwqICYZjK+o5GMVgu+rLoFud6/susR1dqZ9eu5YVhQ8/j2k13R
WFh0ByIZIHemLGsucdx3jIS9FoGSmnQWoyI0ITbtQu1Rpm138qHL6ARTAZt3REDu
ssHX8W1z1mK9wn4zPFPKg+DOqYWaWNTJ74QXcT3AMgkY4fSK68n0Ciyh8FjTPtk4
uVDJUhmSK7xys1n852V/+bxpQWmNnVMJNWg9AZG8iTUZFIlpI1JTwThAtIPnL6GL
DK1gPIG4dgRj6UVJfd9YfqDdK1gUAnMVyc1NpRVkcSvML9klePD4/jGCRwYyccB0
f9AraeaEITJupQyG0RvitEL4araAMOfxxEy1/i0gJ6q8tWsfuxIYWRDINfG0fPj3
dmbOlDi0ExB0HutevFuSNHVTSYsFHKZRDD+A3aOBKLPa8oucyoZ0NuxBJrWUoyHA
DCvbM4AbtDR4VHQJHeXbO01Lh0fRkbyRRWDQpc/vO7pfPji/c3vrf9z7hcHVeAZ7
2dagjMJ1ME7Dy9+bxh/USkFSbjGhrkmeELlXpYCipRBl8ZvdpPISTA6DRqTwGuHw
aKKRgGttuWGu4hTglGCMkFOELP0giMMJ7rs39nGjcvPMUpeJmfKtYSs/DXve0O/r
VxKGwJuD3XSyfVC7+JJTMP0ddboid5IvrOd0x98XQytlFeVcSqTu4TF0S7RKIRcs
wh+HvOj54VLrsmP8a/0u47OHMl6JFMPZeFam7KM1QTXKpwgnV4DD0dtiEQRlBaQu
oOYJey2Mre6piGU8CARB31yZbNfiXe9Xp0zR1f4PLpKS0zI/hcw2fpHQ8iEEDwHI
i5TDxiFcHhKmSVtOr0gW7N84PdH3hBNB5bTcOi+CCwsU9HNZJoOTNmU144ofRqQr
ig/46NWzxZDcvOV7gqXnaLAFVn6lOx/Xbzt5ex/Rm+/Dnofae1ur5WLsHlHZ1YTu
WaeYvZ1awUUwpMHpEAXv7TldZ4yXBu5DLzbEgXynHDUdTZPK6jsHcWQ1CkJflYOr
YFFdDeyfNk0/nxio3VvYHTJD0rIIf7uPTCABL2RtCubg6AQGqIKEFEZgMdeF38vU
Zb/8kqJuW+LR2GYxPds3yEEsQAk9995tNDCtIvehNK7oromKxfw4mO5YXUE9Cp0J
BSeB34ITO9aC1FYZ8A9EOK+vu9BlivIdHlS6pvmoh6EZm7XjC1jav6ad2sGDVm43
kq3Uh9+SepPHCvpNG9BnLTxalmx2xLaV+WxIDuDijnqPMX6pyr8lpD/+EiYLDhzi
Qz4WHjaouGKEHYUBOyylhBqQDmLwI4kCh17uA47esyvNJAAEG2BQepoapBfWLzTY
NfOZ7HVxVuY0+nArcQBfgiZImjwXNSx3eLIctWSFcGC85bXb2gFZ6WJOnEsWAdQM
gXvqTGOtpBLs+YAQBpDCT41qawMtz2hY9f6EUh4HLpAtVJq6O2sR1ouBPfljd9vl
SIDRUog0awCyoqeNOPWMN8lFad4yzU3k+jZhdgR8Qkm6DH/aaX2C/+2SHqYgJ2+g
G0K2Z9MYoSGscwmYev41BjQVUPxsB9Yn0m074OSuE03AlRt2RZ2nHx0LJxMP5oId
NOBfsTfY6zlCeBLlAON6fJpGRNQOjO47vVzPRdRVtKWaZVFQKrX1+VSEqedx8tmB
fFEZPdX5/X+c4XiBPpQ3ntKp189K/iPccXUdwKOHloJ11tHVzswU5vhvQovOVZAp
kdmkbXm4u3A21JpVa3PlbpwyL7V4PXmIWejsOgStZYb9w3shthT+6IjQF5fvqy5V
vz7uslg86K2bRqmNgFFabyLgIlepL8s1Jfw8DFNlQMul0EXSFetdrVlI8wQTNNti
7jIBL8CyDghAd5iSnKOWUfZQhKccUjQyj498DJaiI+i7e/jRVP36wCKtM5D1rv6d
jwIGcXorEO9Ex5IQ1R1Vjkgg1v/wiCWvAPdLwdVq+wwSckdC58Fn6kKg6dAuvGCH
jTwxy5UiWhx5OYDVJkxdTDmmqVNqnogBwJ3gXo14QpqWsHpY2wNr3K/rZ0k/Rg+s
sStXKnkwCAypwKTO++YIr/bZF8eYZqdhXP17VTIgKtXJRefKUXlnM5wH2TT/jGpX
h12WE5s/Qt0GlLEoRPpZxmlmDie1XS+Q9src5VF9Wm3zLV+f90yKtfvXc2WcNhEb
QmD8qlnrUwZXpYtkJg+iG5vfI0m2tvv2sWxifO/5w2U3leLque5vjoDQdmvHM/Az
BZoomZVHpa0/BgJLtIbMbeIqKoQoU9ZXNKG+p53y6vGuHTLzLgQaYgfF4c03beD9
9Bo7zA8j0NUikP/HTlws2LL7DDFtiOTvn2VsUH265P5QQFtxaXuoYknYNbPnXLei
1q0ofA5HM4/9jxPR03rTHI7N/MvZBn9T7sst4tP7HvMS/wXaJISluXnIpPWBOuH/
SmCh6uKy5AEdDoPPgTetK1VPDhTfXiuqxKZhvCk2AodPjezOr2ztHu7iZUEv8fby
lws1RfdhcOVydmE6PVZABflFXbynrLtVhmj/IlQPKCrsB0sfIE/wpI70wYS//RLx
PtKppvBp+KW0vMCzKxyDY2IAS4rr3y3l9A8wFqozIoXWo9VZuC1VZRjVZOS+sdjL
VlZhSJRB0wIwTtPmzDnlZ+FhGnLNrBaiK3teGD+JkaPMeIOayfrBMFwhIlEGEhau
Gauo0faFfvIQYWaSMNnR+Ld2uCm/B4AOD+BMrdhj2V5/8MaIM7hhxX176Yr4ZLiW
qQ1ARD/avHHt/RfQLnJvB+CCJuHqsbg0Lc6cAin8W9sZolL9bvvUcs1rZW0xj7SH
73d0xr6/9doh14nfaDEOaP/cvpfeO8K+atHtNu4o9yghVsk+mMJ3FJ8SSnd4MaN4
0qwWAuWojBmkV4fA+kKSOG1XZSZIlaqHSvpUmF8a/X8eZMeMEVuPz6PO8mZZ1qgT
1+IogGsnEoe/6NPXTWiaJBIqy3Xs+eYnXEEqJoOvfEsQaxbNcIewv6GIwFvCQYYS
/rUXkkqWGZrTo6pE+wmtAwAwPmyGPuoNl2bKsFZf8c1NNOa3lep569igO69XUQv7
gNadQs7ADZjBJI5CwiDQLYU0gtcJjvL8J9FsLAca6mKEVSiyM1XuNbHLfrTtRq4U
nBmZclP4aCtX5sMSwVd7dzFfKVqE0Dse5Q+f3vHx+PzqFYDBIBdKvb+v2DdSU9lW
WMFtmak0MHAkPTcwdZC17huK06CPpN9Z7za9AXw7ZzISaxxQZExEmxcYZoPXDS/3
7dtdMkzuWgFo3xsx5cDl3+oD9t9FB+GahoUqgHGeP7ybosM72J2sodCT21+kOVnK
3/PvZWEu7EjPK6AU18CR1Be0ovCjy8J1hG5jlXE9P1W5moUCBAK5qarnZ1CaPg8/
A+P0h94toWxU9S20ALGwJqH6gImv5Csedd7FDd2/cxkRMMVR9YKkAyYynF+rb2pR
7uA3wJhrNm6m7OFmYajxASinmbN9/aTaxXNftwzt9MRETTwgJJdZXsbnh69w1Eyl
INcqpCsQApluhSkaith+7f3zSRjz6Vbp0qTcT8sZLYMgS1CVGGbJ2A7jEqXVACAr
XgZGZ/rDra++esLLoBa7nZhX4ZJeTCayRTlE0psu5shkF3fvfg+4SrMmwtjNwWJb
MPW+Wjj7I/dkvxjSiGK+iPcanNDuvRJLCir1NA67Cv6/gOH1qUmdja7TSxvUmfAq
qZshibU66DDXoNHKY2JZXLvjbOV/GMcc24hHNJDhcsAd1oTE7KFPOKqOCvWDNN6S
RV0hKyFovqyF3u+bK6FhljMhaxEA0ZuY83sg3AjB1yO/y+FYGerLceW7JJtc/2Sq
U5KVghtQLXBOJqPS4CORjXRQhjbkWtBz83V8Uo4oA0Ti9q/OOXY/qT1E2dJckTec
dujCkHBkP12zeF1RYp/SaalvGdQVOQxiS3j8jMpbsSlsitABRgnEta0KwmKb6gGo
uUVZ3sBhIac/9asQRxMyg2R9UFvrIZUTIuNQ6wo6JBVD+eGjPqfMglkqbqhj4nOK
k21vL9GjqbMwJJiHfbKx1Cww+5DxumyTLhyHN/bjBMNKBL/BuXq42de9uBb7GJD7
GaXUBndFssKPrfCyu/OXqw7ey3SSgPC/PCTekfDda9heUMiJ1tE+3x2vOe76CpRc
+1WX+gniPiDdMdBUy9G2g60Wc8BOiTFo5uwQ3i0ZtQzMHmRLZCtnZxKNKRlBRyVR
0PtdryINMTT02s7XV/3XBnsTZKM3GTXhNrpe+NNA3FWCHkJlwhXYtAQDlr7ZbQpp
pAKvxQcgvDm8S5SbqcjL5ShCcb+j3DuuMvV5nESDvV5yKiL4lVnNXmC8xx+pB4nz
1bl85AneAVpAvTlltT9syrJLkHPPgX7PQuAMDTU1qOlirgFQ8Nt9bHSqHl1FfW/O
3SRYRWUgiuoibTFcpmy/TWxp5umAow4T0hbA5ZMIDNZyN9FfLof7JuR4JZOUxrUs
Kbi+fEOKRYAG6NCcm0Om5GTZzR4ZUzpkw+errVeeWw+VmLxYljL0ZAM4cLykVnGi
R94tHJ5fztnefV8jYj9pEIE8KYJnog6RFTfbb+Q+vEA4YQL6GMQznlHSPNUQoF8z
yKVIEdTmwhac9MJBKyBxEFrJxxfRELNo92zzY6QDx2ZyjXIj8zQy1rivYDRzL0JX
kMDntbvULN2DNHsqz8WU9dBoVLmZfTe3xvEy3XNtnzC8MyrGt4u85uBRQQuMeaP0
8EIruaTTNT23OFyxmFeGhUg8YdgHKlRpAzFZUiX6mdt9xj5RtFWVrebQifQ9FY67
3qhMRPKe1WsfAcV9WHV+GmnxEIKc2lC2vdzRrlJPC80YRM5Txdob1iaD8RCAjOJt
feolQr44yocteR7Csrp504OMDQbaJ3NwNp3B+ci2Nd2C96m4ViOjTDiuM0q8YjIZ
Ki/U8R2OtX3z9fA4nq34BP0RLQ3gb0qqZUI6Ix6ueiCZayd7YXImwBdA9fPScjhD
qxmHwhgdM3bpSIJme4fSaKBUrMPfw9B+nj9/K6Bt0o8/ZDj1WBuGHjiIGyuk2oEB
UBVHpfzExr6HdfFvCjbDHje7rZZGcdaFy92uy0XSOBbywl5Hdvjo8fpUY2eL8XTO
/8ZMYHC/1DRJbWhKYOFORWD79a3TAx2JlLqQxZZqDdGOwcwlMFt8k+SimGIzRaGZ
Hq1sJc4ecO849If1SxW4fRZ+QtCWjGg+NR9HlPEfnE1FoTvffty3QxUYDgaoES02
p/UzrKFtLpuCIPTK7U8A41Vxk1UZLZMGy8jAAR5eV83lW3Rsvm1nrLDF8qkSFn4/
vlrksLfETHX2zYnwrXh9v2xEuqEbKf0+9SX3OPbR3YPkxWIXyxoNbtyil4CiHvoa
M45veitAPrhHToG28u2eIjEM91Xk6HdDNZ6gCVZdX9eHb7c1kxsNMXtWfAWcqacA
nPQgdJNI4WCKW0aHSh1dotVQ7DvE4GR0ejUG3zM2Ubm+PdwgR+1yEhPumUVZTDuG
tJJihKqiw6iXBKcKTvv7NRjlGT9QA+VQnWBiC1Ny6Ng31sjsLd7rLmveT4DUCzC+
8EMHIto9k7p9S60tZWJsML2kbqo+TgZHSeRxhRz6rKQTOyQtE/KGM9HhGm5VkuGd
TI6KPS9bxaz43deLpTCRpZUjB4ael6PvRaSI+/5V9mMzZ2Ad6pIYbZ47V86wRmmN
MPFYMy/bLGgJmYp6y82B4uNLhtcb9Mc1ChzkhGogsMh+48duv/d60jXI7xq3jcIY
UpTtLGxooDJEscugtewK5A+FAcvxBlOjk/SNIhzQuwuffpUNcx3DU0Bbdo+fA4iZ
ATP6vU/SGcfqslcpuhuyMHfH9RswIgFG/Oydx2TPyOmNYs3abX3XEPDd2ZhlcGvL
RaMaDUEFKiBc3eS/kMJWe+h4oi2sfmDqkm5ir1TEH8l6ddRr3fEDv+grOvpBqbZe
qrd5hnggQ0sN+kq2F93Qqrhi+c5zxF0nrBi+BL46JIq9FIwQvdMOgmQIbHzIPnPF
zYzw2YOJbE/tiqQsY6PooMNPT0QgeG1WOQ1zvg4LmkxM/LguS9xPX21923fdhwaG
16xfHnAYmx+Duh7gQc/EWggQxqeFg7TeFG6CwIRgn9DI77Ijw6qcO9VoT+KpYTYV
wnYnRyzfnGyBBnEYShVZxexe5RTPbsS3eGlsWJ5RGnUT03TnqAuK7zlH8Jt/fE6m
dx6EljPSIEtTfvbrIFUABnGSs0L7rcvNNv0oTIxOUjbu4Si/hhBaqbRZGuaZrNMm
wSv1Zzrhev3XGPhO6xthRKU2n265FypcmOL5qOqcdksHsLZwOE9Jd61aTldYw4mt
3qXCrfb7yf6rY+FkO6C11emQtBs77kmm8NFsx0ao8duBwWJcY/+T1QRVf+p7H6SL
EEQEebfO3Za+uZXCsKSqXBBN0Wq1d0WpfZpEiF6zsJwmXool5Hq37qFioZKQTs1d
8TSuSNRTjz1jOowcNx7znatS8nedKGKfePumRYEHSXsDGzsGqse+skjYQMvq0l0S
9pclQzStuyT3nJj6IfFkPuFuGnj8cNbHrD+s7Utbt9MCV6z/L7V/FnvoqfnsWnIR
lGhXui2YDw/FqtECzl5JUQY2p/W0glquYIQDUbFjpp7OJGI5mndl8mISManB5GEl
m3HSAmVnnKHBpd4Egqkkx12YJdv0GuB+wwL4aurnuYOZzHhlBc4nmfYn1217lWQ5
+lK3BWbZ7AWJQU2foU+60kvKvwvd71BIYaiQklJd03Fk25ieidysxa8lVK6R6Kt/
07xfFO7at1BJSE3VYKEXUb1cLWiRepps5Y8J/Du0sigt+GorVlXKy+FPG0IH9HYv
Y8SeAQj4DtlN+KqKMmH00G2JSQIgtfnIfnb3C2ooRho7yt7mY4jXEzU+FjmGZ8Wt
d9eCAqnf5yWqS1b6dNM7KkXvSBbY0G0hkpa3ncmg+yUEGhTvyCz9eJ2hicYr3y+O
3m0oWfssuBuEwJxYi/1cpD/epI3WXsph/fCe2Ecm0stsEpjZfD2OBKfAJ0btK6Gk
7XCx1l0hp7MHUqEUF0ScZXiE+ypeA+N+eomnci0LnMwro1qTWLWkTNUrASLHrL92
FZUALmIOlE7BUlLp4/Scv2RWA1huHQYTnDyUuAk1Ou8rcKIR+0hWl0K6gQKQpRSe
3F0/nIwiVny+einxZo2bjHIJCGK6ZqFfo+pKfMHxVSelE5kHgEzYHv+JM8MAzqiC
J3OBLP51oEGeqpXvrfOpiF2hicRWv8P4XCPn7NkDrwTmg1q4U+buFzglPqud5sYx
nLikEINpdnEyVQOHkMqMhwN7THo5kseo59MWyU26geZmSgU4onuZHm/2v1NLYSXg
w8HHZcIdcgS6nhjKZV9V7wWuTBqtAc5REdRmSHbCdQaZMzPh0I3cHE31jzWHGnuf
BhISaPHysBA4xsjxP4kdzwBd3LpnwK4qh/8DlhM/cYT7ujzzb5wTNA4dGzGWpZoX
O//HULavZUap+m2hDtL41KYO5k1tRhSZCKTWEuAbGs8scXWa6xD+nUBs6/6wDxie
eJ4vy0iYOdgiOf+0wlpPssyFTicLmyvq5OR3zMgXUPK+VN4lQgd6GKd4/0G6Xe7d
C/MttID23G5m5ZM/UO6ydKnnSqwi77jeK6lmjqjQPw04K3X9oUF4kmwTZSbYMsFl
+WfvqImVFXCZOcHqN6szBDYqScaG41l/YqNo354obNFPMz1NBsDW7CUZ5bRwT4yd
2YbJcjkJrnvFtyU8kqIxnPlg8MLhQuquk2uMaayLqGBrzAv/PedgX5HOUtJXfEmn
jKT19VXgvK+uof1vfBqmFxt7WjdxE5j1dyVKMoNAk7cTdgktdmBchDrj5WA650YV
e9dxCcfQfl/6CkSmHhPHnqi6D86p0jk1HdGqiNFaiR/Q1EMNqulzwvl6M9O4hzsG
0wO6ndR0TJ68So96zHknTJmD5alBvMq6qe30kV4izWreT92hb27Xyr0fn/GSIiqE
MUYcIg4OHUSvvWZ8xrkfLWqgk3ktgO6uvON4pDcOPvJT6boVDZ1Hso4TccXRWi/+
Oj9RkYm8ey3B08NWTlNIaHryTUTj29LkjiRu7mjl0iICQr+kBsdqAECdDJwcISfW
kibi100XLT5ET5tMmtXLAEpWvWZTE9V4eAwz5DtMgiviCT+JJ2iV+T132LcHv1t4
vVEy2+5iYBPiL9hZfi8djNOEDcuZx3pgHQ5oTq/COvO+MVwts1n92HTAERAYckzt
5QrXHZvx6i/t+ByVc6wxnTQCalIjwpmo3DcReOMbn2d/wXp5uy5OF9pNK+zTt/GD
iYLYtSLrbrW0sV46P1Q8cQnBimaDWjkmoJhlhhL9G4pKGxKsZ2VOF+2LV+oyXKRq
qPNKL9AHehBX+bzRu39beSlQP7lLid5VPqZMyO7af2QJxSo1JjiGpCOwMTznO9ui
FUytCBmLkj/QyYVm0pCV3rpbYlqiU7+mT6JBrSJ732PdE3F+1tRwQjGRxW2nXMZG
2KydyzK9fpcQIpC+uMbSZ9O4vN2AgG6UkwwjxbWZ4F44uo84AEzyw1x1fPLqL/4c
2DpqHOe3atAmGxN8rPFQCVH7Js3j6YFMtxG40W70xWnzYjC5wDVv9EjDFZ8870/0
gYtMHbWi2HMjmEV873EU35DMCcqcEcTRcl9BHpGv/i17YOmgsoreG2J9wihZTet4
Q2vjjJjVldBz3Owr2TXVN/XK4KPkVorlB1W6kb9f4E82ISsURLoBi83A1niVL7E1
IqNzomgnhssBoq3G5wCOuKZthSGASH0iRMdQiKzYDLF54H7Hm17mJFRZ0wdo7OqU
b4eejLvTDh8VT4p+InwnDWlCh/DsL+zGUNicvlPOk+Ib6BOk2DXxPakPrNHE8hyp
9XAE1s97nxUsAafQLp7gT9Q8hFBexY18hKCGIrf//iqPwSGwtqK1wp8PCBvo4vY4
PvDhBWoYPJRMzqJ30AYzux5XcSi3zLPNTRtuvJEtzr83TOkLEfgz56fxe4GJU02y
vgPdKcgGtupauowmsP+9fbQijZ8VYtmAt5zkE1EE9iJBF5mjfL8WUNMtMgKESUg2
mHlyNWdOElWncH/4893AmfiEKoJwbrSiYJjD019LH1uthAOZYK8MYD1rYrIJDDRF
EsHnswGZDrBpwMnWQoIOL2YeXasuE5nXtTvRmkIP1c02kTs2uAajb4x0f+MAq1vw
RZo2z7YMeXWyv97RpteoRq77EnCbk0N1EdpvgUrJRHEa7k9qyD5TJLaO2tb3UsZb
erVSVWkLZS7pBe3qh0wma3LxuQV9ceJuPs+N9T6vB49u0jitAm7+ImJtaMUUVK6Q
Pkl94gkGXBeaLfjyX3Wa+V+tnP5nVOEQADt2i3YXaObgpHEk1Ph++x4u/Dd1TK3H
3K8CHKU90PPBxOaDZammVwNz1uEp1s6HUPfvNB9lGQPvDJuuMehnGeTZpcAhnedD
XD1ZXWIbdLm2aF4HBxc3VSvv7SrX6E7S0WGTitgoR9Dr7zeJZERjQhB2O43MmrEe
YZpBbauNHHvK80pFgu4URYCsPnUBbPC3EBbt3tdqN7LTBxocUCalFM8B01zx6aQH
AxYBYnm0Osp6lf5YloHEz53D9nTIBkLxSuhgljXG5uznsirRB485HC7askrsXuP4
LL52dHlduoYC8HqzLO3Ijl4FHheNzqa4OxX/4E8a08pWW8P54iliBdQZuB+HDYED
EJ2aDjklhCp3YJ37FSVw3DWRBiSRkVez99IuTNDrcwdD8KEzAV1zR/NGqvRnWTDI
WpT7s8ctmY+Snu12lHJvpasuUjgQxoeH9mbksbVSfPY1rxji2A06bsFSAX1BRaUT
4g/PTekLOSDPD1Zs73NPekA6jvEAWxHxjUo7f8CxvTbKAMkVq7uBgfUMGo+fVWKd
c1GxVbGuH+y7zbw/GcCRV18cr6sBO7naiDewROjeW3Pg9wqpOIG1Zb2VL0gI377H
MTnwhayUbsOEUdPAR+H1Z2SO+6doKCaP8Sfd9PYoE1ILkCXtfp9GgUc6bvCyQU3L
XQJFepC5r6E8ncZRhYoNIAi7KDYaTkOWT5t1PRqD6URAVyy73FqfJ1DXNsdyKHzm
v2MKXYwgD7o0+swktTgifmTwWuLGmw77K+ObBiiknX7Nu/aunMbZTovgtJk7etMk
B2DLE77PePLl/NgUZoBQCkwlloQJ+fZfZVOjtMKc8DwrlCxPa9mkHIKLsoSdyDqF
y/2SOA/uExd1MHJvXdhuSLqeKr9dion61khswMyXwRGgMpSD7huHsB6YVHF7nd89
Oz2OgfzD26qmb5sYICo3awcTndIhQSPJNg95EKawyMhyVeRZGnWmvPl1L08FIJtH
z+Y/y5sD9JR+LRZEdS5E25h9oaz4e/L1zj0MvEeQ8KBAVafe6/Kl4Th97muPx68e
dm3hXPcT23tX0B5DhpAqqk/jUKtLBoOfokNX8hZ50zGS1Y8dZwwPJjbOgjuExG94
G3y/APu2NOcBBg6E0M0JKmus7pbnnX/n/3gn0WgP4kR4AntLdclsKQ3zFR66Fzij
F3XFhMfCg0yaWNoyFIHbXlnM69VATEqd6Kw4cAS01ONrmAMK9/RijEsB+fE0YgXe
W0qjqgvf6a+L/PZffWH8QyaeEoAqgpwHbND93Zj7xT1Qkm8wTCW0aFk2gBRxY48c
SHH69lRrGL3sqMPMtj/knTc17ES6gd064BGa0iOyxamVlV1DgTe/8je842AwX5Gf
IFSytgd/xiST9W4o4+kDp5xTvjebz697E9Sm9DEDRSu3C3bZDA6Bo2S+X7/ha1yH
3UHGYSMXuGwjX7tQwUxmndXmrOOUD7mbO963bPaMYODtDSz818glH6qnHO/gVmBf
S3ifZRGEPLFW/8jArSlSA8ixcdX8UBsOrjJ6AuVD5b9e4KYwQPpL2CUJgV3FZsR0
rQU3uVe9lZJpl7pvjoQ3oqRh2XJ4qffXf/yE4QEcvOKoDquil7SxIwNEK3ifXNJf
Ljtiq4Y8Nc4/HOE/lE1lgyn7J+LwBC2R+Q2nWtoF9nSbRfbzAJu9SmHIbOGwYfkQ
BEonh7YXgObRMdDsGzCEosrNw/VaZRvD/xtZ2P6goQeRy/C3q4GKgnZs8plbCE3W
4hxRNTDubYn4iQV5mCJ5dlXFUdlXQFyjb3K7foy+EwFZQD6rcOHs1ypJISuCoVWs
JEcYo56HIO88a2kLldGEuHSaMrLpsSnzvNCoUi4HYB7ILmRePilYVL90V3pBO76n
yxArYXi+twbFcG6wrzHxgjxz7GrKflOZYn/57ohncP4qWShGOZpM1Yh/rBm+IJhj
X9eD8ZjohmryadhtcPKD6K20XW8VDZguXB7TWoGP2eAIoZmHWH15gEQhsxAZmvts
D4Lnc3h3stlbcy8i2ZrYbOVsNJTRv+u3w6oNLG5s6YPXxJm6ie52BDMXNGrr3Jdp
Z9qpZ8lBNpdjyPPAI8NZ4g1z2VTcgGtovraTxirX4g8LnH6qm7+ZdZcOl4OslDGx
s8FVqybpON3FcNRxa24xeyb8bAaK55y0Kru/djrKbfusz/MlFNbGPAPhbriuw3te
1JE8vL5wLYozYtyt3PzjMJ2i1K8w6b6gBiD5PUG/poNkNtw9y9kbXGZdvQqhmvic
Yg47CPnHL2CbsKe6qTGLOZMQagllVnn4cD0LCxQXqjiFDgYddcfuKHpGvhORvBDV
pGSEJPwuR87t9YjQMSqxayd9MLsEgg+vCP/U9L9u3i8F8ogjgZAWJg9C0BBr/4iF
dngIVXNDDzd0DmslJaTBrhg3Jna11N0w/pU0lZUXTJ3kXdXMbGYoferxbuqZ2u7w
5dYkYxkmGgOAIDBFVUozJECYlIrKdqjfY0i2Sj3lbaYLAmJiZ5+8LrNccMwC2LIA
EdlMufQB8OLPy3N3hfE6JcJ7a7JFwrc0tonln+lQ0ywRfQm+56YJ/5PA+rtL2cPj
vfKo/ulmToqb6nrdx+xzc/EHJJqexHK6F8BwoR4HY4Xxou5OSDsf7lU55pOuUQKh
Ht0+hPGbJjsP05O8BgX2LcFtOAhm+jFPZVuxcRIlZ/fZFKmRSSS0UADrc5BFn2IY
/5HENUgtVoXqcTe4kzp6CJDMRDLc6yDLovOIDL6PcZPzVTgTfAw5mXbaRladqzlt
SYvVB3wYynC0PeFrgudfgArnyHVnsgovcqr5kTVw7E+SBSRWCpTslANhOwG0mAy6
+z+G9+thwK1R1MBQY8+9TXal1iWv1kVNjIk+rNSyIK1Idzabq2FxUSRj3sZn5Bx1
Rh8T3+OaKbZR/bUPpsQZ1f/IOnZqWfFfpGGASLq7mL4tKdVC7vBtDoeEu72qWgis
taJOwDsIh76yIUGa0CAnuWTAf5D4c/Z7VPN+bHHTq8qvZie+zwq1jFDF7CbKC+RT
+qqIDIVmJczlPejjJ40QucffsT7iE8g7VLIl/oYWTlsdHg/XxgusqECHFAVu5Xtu
Ua7Lv9tGdNHE0SLs/7xCkSHIopBlwGhtIRuf+GEwoOHdzd4p4ilzC3LzeIXNmKZf
YykLhKxYkW4pS2NH2vNF2dSQ1bLU7DjC1b1W8K3w9lWm0c2f2XbR+zoVUL74+epk
tHsEqREx60cCcvWXzEWkW66nWoYUrSQunp6PGAhyYg/0NA0wFE4vyDj1uhJpCjLO
1HtUvLE4dD0M8TbnL/RcsQyo91sDjhCiuLB0mbEIKAvy60q8OSZq98BgNh1Edij3
E77zs0+Y4VIrt5I/+I08HjLsWRt26rLD5t8LF47L734CEuYC2anncA9u4aevPopN
o/Y1ldic849MQ+eNHWCFGAHnSCs+EKw/XGJqgHLRbBVgQjlsC09im9xWAk/645bg
til5ojtEyIpNWfwrjsKJNpFcG1Lxevh/tbgKChwEJxLqitsygndoaKNZMCnddz0K
xqkUeLXqv5CBEllXeY8k0ofzGnfngGF32gqDYdklQ7vFge0MfCEuvrafoaG49X5j
S5dydDhBP7fUGiF5xW41wwvKqYqCfN2P3NpLq09oKTtYtC1Yjm35OJ9yQWLigyNz
iwv1CzH0WHr4UqvaN8V+Jv+L4bu0bn9trpIEPMkFAl5EAotc74DR9X+hs07DjxJz
Mx3YHcTaH037rL5tCCRGssxQ1+hZFv9rT/kHcM35cCJvoHoAKrkKHc+09lQ5Pe81
LQJ9mLF4yPhCHlRROAOppMJrTlrG7xIJy7BH/IW23kIG9jWwrw1ix8s5eflghS44
3UUsx5H4zym6YDPDJrD8KT9BkEBCIww0f0bDBvVRWQAQMy/7arnBkxmqxHk4XTuU
SD+XjPtw6pNqabVuWd6xkuaQGVJLOzTLuqzCgbouC3vnEkbFJxJCXr+UCjPNwTJf
RdLVCK5LCb+3lqPbs7427WKRp6iT/nbypzM4Vl3gJ+vzV6K2avfmdR62HjOD2zti
OjAwfOzrl1Up3/KNbKKYIpEpALv0nWAiC9SJEp/COSuu8r/0kQLkh4tjGFZ2zmUT
2V+LJ1wOA9VdeNyIRSych6VmSloXyXS+G1+wZ5ZNxyQb4jBqHPpEtKn3B1ggZq9n
UEyxOg2G+YFFamMqZwKEt7NgD7lqDVKqaHXSmBvTrwwFgReDZannLfZJm35PYLen
zmgdEWQdryqEFR5LaXqS69XL6wnmwwFUjN9BVwfxtlnuyYUC12nwP35l1Jp6V7KW
ZrqApYGlgu4/Fjy+wBVfjfc6JBrO+W6N0inJMZ43TKRuS0LWvJasoTArPqNzt6dH
ZlhgBf+/5v/H7RWCkLaNWu204HDTWN1XsCgYrUQgaLUHnKgxQ4gc6ujbyOrL0SCt
ytfaZjNWZe4E9QJmwHpTYs+eImhYuJW9bBPAuaI3wQ8XdMq5SOAzBhaZ5XM7SxPU
/zyEYIY3FYFj1JkpIXmFtibq/7/+bm8SsMJSa3hgeNqeNgmFzt/LKB7SyDPnfQui
gNpYKqu8Dd1YCGC8qXsZOAs/ndXZw1MOVCySQkAbRCdM9s8mwhsUELGeoVa3Vo67
JC7gcbXv0thyn35ICcLCTqoQiQU6xb9b8HdaMfRbZwnqu7mDflGt+/SY4hA8phxQ
4lxxf6q55bD2g0C4zrULScD1LUqB0in9uVAyBF+jmf/DGOR0PKJuJBTRMIZjyBBh
tmmPVJt+srY95iVcUuHKLyI8SZLw8F6h27EuEEQ+8ZY6Nb73lU/ujwZNhiWYERTV
gFF6oAlG1KIGqA42mmaD6UPdWUi+H1FYR+hvJq/oN7Gz8Aqx4dYKiE+LjdOos3gc
vLoAGj5JB/yJ78Lv8dKd7BDnlgWNxrLhm1pAUARFXpTv2YF6lDgEcGAllim/HKS4
znryGjVsvdpILrRqEk1i6JR0YO/U6INHRJV0i8TMfirhOlFKIwcOBrl8nblQhdHT
lspALtMhyt4pbONIANcrhdvwBqZURRQGK+KAjeFYjb0I8ZXUQ5W1hDX1qss+tKUI
r8q6Io75RGx3pXwJXBhKM2Hlvoe9L9AhmTNX1SCIvi56yDsEss4zxiY3yhAaliFW
eZ1x2IGGR6Q99pw7FM3N5COEr15xQKPQsps7JBOzZ4oAubRlzQq7FcwmlI9eqY4B
l7hLnVPG0ronMOt94BIO10EeL+vGoe7SPbv/Ef0q5v/aQMnET00pHC7OzsD4FZYR
EmxFyMv0mqHKC7VEh1HWYMi3FiUiYX1p5sJuV+c3Q0DFklvt1OU6N4Zyi2XCvIu4
vf47EaNqT/pWKeF3BzucG8fbiOsHIZ8b+g5gzqthjhkBXgodmOUtCSkIMN4hvOEw
rblT922y1YIr5RLi/RcmB+uzuV9t8pzlYoVScoMZZ2wR/YsI0Cgmr/UwouRlk0ZV
GHRKNrzSF9UpnAqJkbFsZ0HcIYyKPP/HKRrZnwyUSRL01hb3hdRwbku9BbCutEg9
Qd0fxV32CWWKljGeGzrn7oEJn7/xulYcSli/XMGU52JE8oQQatMR0ejyDLnBblha
nrmeDcUMPq5PryHjrSRjjK4NMzl04cBaCMbKRaAyDCT6+aWBPVeXi2MMkVQICutC
jzF7BWrjKOKl9VxqIhxSOIF7xzobnAWUfHRzwh0WKmudc8uZgzS5fUvJ5gBQhh1R
jPKJELDMFBtKSFbBJ3BV/sYLi+pCJ+EY+dhJPT81Ko+GS2ugR8d9gY0mVYpzmyl0
im2hvemY4cZy6DjegvicWoHwc08R6QOa5ta6pWbbQr8VLXyeUxJGQP5dCbvDqWIG
MmKD9YTpvlI23+1TsCWLJvDnKkM1L0iiMYHzLiMAaITsaF6Nx0oKroIfg6cdZ/G1
TDekMBsMk22THKysRGXimsraEJtx08jruCGBn1yRb1IvF+aR5y+9RHKWGh+3Aez7
qV5OXUjTHd19nr4pRdY57s2Wb3eaO9LoeaVXaCqI0AaHKa+53V/b4kTY9HNB58uM
UTvpHxp61F9GJ9cWzjmMYdYJDxH1wJVf3L1+XD9NHLxovSayU1+Zavb+ZklhlWTW
UuUgxwXcwwcZk3fen/qSyI5oEfrfeamLlCZ87zYp3fM5+0HwMD+K/1IYj5lpezW+
QHiVlmKQOQ+LZBNh3jItx2SyblIzhnf7/TKb/1H2w2BiudplwOURMrMRtV7bNty9
vL5EP0iGcQ1jUldmVOPlVswne72IUnjiPqLhFIl1Y90fHZQgqQnPpmCyCrmGrsdj
fUgEV6VNkzR5ycM+hfRYBg8R1ml82xJeCxaIuGxz/EpYeJxo0KWrZH8ZIlnOqrWf
/y07/LeAHKm4dtnzhE1BBAQCmc9t+PMc+W7a3pt6PTV699Pu2Skxkfj2tZWvzmTl
eN69PZTShps8LxpRrCZMyFTJtWU5wghSqk5g0hq4iyLv/3jtFlH2dEiaQY+oYNLN
/4nYjwldb4U9KIYVcdrKhP6IONgKfW5FR650P+YyQ23ACsCHNAse2D1DY7Obm97O
9FXdc68NnzLCMsbAXW+FjQtpquqcucLGV52N9UGAGNGNHpgDb68q3ZeTRaGm8kcc
Y+2nVn+0dNxxKHeDJwVOXtW2RUs6rVKxbpJHUQVVq88teayPmMOk3VmtZ5iDxzRW
w3n2gBMF3+K8bWTOaZqgaPfRLx6gxwOcK+jGAjxrvF6JWAivniCai2NDnXIhAzL1
baLf4xDkhV6VdcwiLGoxqb8pwhRjCIYWvCoTwTUB0QKAMALP4JBgObbVZW6Gr2pa
Y9Dr5jpCrdAbLy86mbytVuSkeEYIC7sueOJPT++KtbTlEcxv88sj0kEQbnByFi8d
IOg1rDWGvTPyp8bA+hQg5nZypxUITflXAB7cuUd2tUrxLKJcCRfUN3UIvZAmHvxN
gPQd6pdJNE1AcuX84r802gbU0hLrYE1yVFNJ5TUIkYMJjD3jgZ9miukRm+mOQJnc
/mMChN1UiKT5VnjC23KlX8BzpZ+EQLO98rLYu2IoXwF0D08geGdRYZoJkIQk9wDZ
OSw+iJ+jEEMLwvsJ3q7AOOpAjS+lqsBHQw4fq59+NvTmmsFxCkKvXuXR7bf0b2S9
g6n5XRLj8Eb+zub399iDtv2jJHqif7TytK1miHEAKTnGrzTvsD9rAiGiFdo/R75u
fUhC1lDwOTzOghFCHZAxiS18TDc1qDBYUJoXmGvN+KJ5xnM+bH9UFnR/wK5/1lBe
IidamVYINg1nAXcQgl5lXBOx7ix08ptzocDtLyxpq+hFqjrP4z/JmU9x5TSf7SV3
C/FSznnDno2skEP+yYs5MtTFU+3OnIN2Cpj49uAdZ/cxwNeOaBtogLXo+gMUYtvx
CrGeHobAQy1ZFeNoQfKtxYO8yDfO1jELPv0he3j2pcSMgIeFlmtJuezq0l6JxoEZ
Un9VM3ok6wLgooxYw1Z7GxRKQsTdaqB0SNwrf3So+WD9ux9tDTzSI0eHV48AIP1N
XErK3xZD+hFYjhj+p6Zx4t25iYkDo6pFQre3JT7rimfWQNkyRmApUa+paJNUUQ78
jN7Z68eP/HGk4I5dGH42u6c4U8UrVKOldevlX1jqxmZzjD1q9FxhZJ8UlDstKnsP
JNZ10nZwaSwl4jcn1ze9tKa/NJM8BR29Yrw7i1kJUbRsqVVrmNlRuMJdnR8F6P3w
1s8SGwGR3XxYDogGD0J2QKo4gln/r+6A8n7LV6uFcs7O69vbUqgmes8PPof2+qb+
0a5At/D5bXSFB538Sgl1rFX6WMHLmWrNeB64OXfF/61fymb6XbRohU/a15IoNnld
6GPcw6OvfE0SeDytDz256uDrFQGWybO4V2qCrmkZi7TTtKcnC3AUsoQ0CFUEbLKs
PiC0PsxhNx4Nh4zKAjYMV0w15+L6zPeJZIQeE2L0fIZ6L2PNOTXcTfD+oqbjKAQ7
P2GTiQ63Xb01rDJJowC3KdGVR/XCL92jDP4T1a3DH5AvI9yn/fZWBYXbRm9IP+li
IZyHivh5xXoXK+yDEPFf8wm2iIs1JWiX2/kr+WpA2PlcnnSDWXqRrwHtRk+x7y5t
jdzrWSsDIgtIOlaCS9Kv1/u3CpLWic1H8uJUXnRLMjb89uIbXN0hpoixgRfk6Z2+
A2/dfshjqaheYilAYULhcjAzSUwRp6pXcv25Vv6aHuwBdPfyzTTPmc+Mj52+AYVc
CMFlzXq1VjLbk7TCHMh103DwUB1rS29KfP0O1kSY60aVTJpA0o2/7B+4Qqp+2dSu
2dxyQCqqBO5wmmyWiGufHCH2snOBWjQKwB8vJBI46BRlZby1qdprZHpVo2cCkomK
yUBNBb5/11J3N51+5qMJE1l9g21DKfFpkYPL2zxIMWE47tnjPuV8d+IfJBppuAVL
Gj5W6N5iN383LZ+vHm1vnXc0PT3yFcw6+YKDmrbG2m6RMX0Vwis3/EpxElT1PyST
+xX3hPE0lVCOxp0YhUUkvXl5Boquh087SrBP9IR9yDYRFJXmG3R0rvKor7QA98LJ
eHlySkbQoOqmKM+79pcH6dndEZNkd5bN+VkuQOBXM84CJBVfahabNFuVtvVSruFA
kgT8VCGRbCNYXNHRK8OkqPXgbmlaGuhjeunqpPJWnlXRLw29HDZbELDuGXmbljaR
qRSlh7Xb5j+UP9P7MS24ZDW0KFhQGA/BUvY05D+05EBQucdZN5tf1lq1BucstKom
BaxwS8s5gWHCIOy2BNM7SPr56NZwoxPAHviYXCMTIeUa03l/xZ8q94BxfpWr59E2
lJQnwu2/uqrdSoL1fnKqIj3FRPURrsESrTPjLWeAYklDeNdne+bMZgSscTySXITh
jycDA1pQeE09mR3pEgRxWyOCqM8DSonEqXHWMR8ZPlLWXpU/vp7KPNuz7M1ljxci
4b3GDu2akTeNqWEtn02N/okJplmzYFQAnnLQJedboWAuwqN+eVkJokJnBgiwGCat
cGMngm3TrcyIBaQQ1Gdyq794tYVGkJZy6GGKZcBziC+yRd6Jiz54/1P73CZz9vwM
wXY+yLe1+qbzVfK8s2xmjlsGdevVJecjOULzfvHZpGVUfVBStLgKKOBNlT4afUrT
FRKiEubBNPUrombYqGVhlbMy501eJazd+mViyKY87ZbaXbAf+pm4geqhnOgBFl2w
w1odFciowpIgP5j4BE7iViVgButpUqTkt9bz4E0sXLWwi9bBobkPd1wScxsHuyHk
ETuW6DdksCFVMs4EfkW5YGp4wtM51qCVVXRzSj07EnWHQowLZjk6RpbgQFr1MzSR
vig2qC3PUti2ExY7pB6MWG2RJTDjkgOVOiSeFIPDz9cFiAsgB6JZL6yN/fJza5PA
sUhJ8PmUrEANBPAqL4yUm80aRRxGucEqEQzj5hF3Agoko2URNquwik7nifr27cPN
7yP7XURVJCTVtIWBn6LzIEYaNNGXainhiJqob3jhyCrCw9hiC2wOAyNeUfE2zq4j
2qxqTZHBet4cOG/9RFhU3BhR7gOJmjGwlr7mJNMruRCXBTzDw9wLB/FO7TehhOdQ
MvsbN+tZAdckWdNg51biZM7RoQMhwcsop8CSaCyz36AGSH8a29MJI07Imr3mR1gs
c+I6L4aJy40FHLswRBI0RU7YUM18z10tFTroBB4e/Gufek6QBfCHQMUe/jL96o1U
8QC/eBPlWaqdg9ACm/LsVAytAbWlRFJTHGyogVNJfpaY81bxElgo57vAR5PselvK
Vml/HTnhy8pIyrrS8olJp4YouCVHKCxTN0IBM7vSdv2qN+gylFiqIc+mfDLzfckn
1xJn/sQjHA0rXzgHRURSXE85qKs73SD56kiBvvxc5IJLxye3KBfFBBl1Kc0PUgSK
Vb15a41fygitgPEYwlpJXI2PxI3+o1ILy0Hf0SzYU9UIFwoRszKj+YtBxIriBiFL
MR+k37V1NN1bxL6KJxdmdof8e7pF3uYsipNENvilz8SpNywVc4ARz6CrFfvGmGXA
C1G0YDsmXC7sT9APbDeTk9G/W3ZTZUv/RjPNjbx2EtUXRhlSrIOgiCkSg7RmgQPx
+qYoiyGVhU+3mvfhwEGvpbIy8ngx5Xxsu9Z9NhiUdNFhT+f5RzIqaKI7MJ2rsq6V
uN7guL0vwWwuEEmaguJF2nXHEGwWnLn6YZnQQr8CbPhu7Sb8TQCvyU2k5I4tj5uA
Nb5CcAzj6QYzniQgLnAd8XJy50qFiBz7MRpOrinwZ3bhLRnyPpW2pwgqyTszQ1eh
SOs2AaibpBJKGQ4r/s30Lpvhq1OgoBqCQzYQ2ml5Bfl8tgDQOyMjiOHAwCpTCbg0
3C/Q2U5Na0PD4xxC8brrna6IlSLpheF048balDGMbyFqYWPGA0vqRDPYDMRceS4x
XqqkuN1H1bL8QRUbQNlzp9y67Hp/JMwEXpjPRsZYTXk1friRTvFUkchKOzSsWD1r
EBIJzZOQZ9GGUQJ1I8ISgosLmRvmkIlgCwgC85XJ3+e+zMEck3cES06CT04dCpKp
3Cp1560t87u37PtTk7WCsBOalTh3B46JV8ezSR2Hohl00bKryT9zrvXbdAkTcADJ
O28xN/l54Zc/kGk4TbvfDAQ+CeS3oPaD4LVTgv8MpxpBo5qurJ4NNeOdabTR0dWt
3QFhiuBZy64zV6va/5SOrd3RXZT3fSNKIgOUn30hYXVb5IFY/HNfG/76XRaZyKyt
F2NEVqx9A+rRXWhfV1Rgnq8QGHQz3L5zywaVBXC7x24F4jrc74be0749uhAGG5te
V3Z4fUSzvrKvUxGW9VsHImMIhkDVR6hosoTCdVBbqh2fM8S5BqaQqRWNo+olm6al
oClvoZZcdXP1e+b09kwCLr17LAzZlGCSLPokn5J6uBZW4qHEScshsSTB7SN/0cWL
IeiglJMgF3OwkG9hTYAwvvvUxtAQw/YpToJKCqEUO1EzJM+XUzoQmFa3syGFBqh9
DN6BfnMssAtPZIuEjbvKLEB6x5NdaaACrBriIuDkfh7m9gWeGV0vacG5A+x2T2pg
mikRJk0/ASuwAtMhZAZ3YCVOj/j57EXvY1uxYGJ3Gaznr2NavTfrIu2GbXVR6N/A
/ZVCvqzZvZ9shw4o9OzBPQOzJRzwZaYeES1dLJiFuvPB0qsCSIQtRVN0rf7ZTMrz
Uh7eUb8Rk6byEbKJwkKsQnrGTu1PfjJvAziReHjS0/N0RmrmMh/sH6X1v2QV53wm
2ojUBwhZ2Ljo7FM86BECmuK2yhhUjjxe0i36wk6vnnVPyZUcLSlM2Tjr+zlpUZsI
W6uIQBtBAnQz0EUCkgMxtm9luQcntksNSLFAz+WD4KX00l1e/Uigl+yYd04ZLTOZ
yM9M83NOQXsKOzYqY7ZZftt7lX1QGazre8Zoj5fPI5Xpnv9z0Q9CnscFVT63mRzt
lDvO0VzrRPaxNrAGhf96tI/OEy2Ff35UsH317BWxtoZNj1SWSN9qvsyXQdhAZLXj
wdqOxk4+WLn0DDUyumVLf5yq2M7Oj+cCC+tWDX7Oqb4UmfGSX4vt+JqUVn2YkiHh
84m+/uJ3kS+kIQi+f2jKBtwP0Nu2AJ9Qo4LLH995QJ9KyQ1TQnTNEE05fWug5B6C
xcQIrNEswjj1mot0KkhvQ9KCr6/FgDx9yuO7pkKkqhLDCEIfu1l9UCJZHABGKsa+
IqpURltQx4gMvqzxHJy2YbAymXulWJwt74xaV5TombCmhely6QgfrCGfl4W2Y4NM
XZJYAn5TyOJfDcLO4L57CzYSFkHesdrRAQ4Tscg+o8Fj6GLvKwC747jayCRRcNtL
d97Prd9BBUyNmAfQkijN/ALLG6Ie2rvajP64xVDah7M9ZRvNsjQW0Ou4rzzBMgDS
0hvxQAe8KAsCRtEqfg8/8qDAUXujB9PJ7PgeB0opu1tPLHrL/1kCBIV+7PkWmqgN
wEzGTvHekzqS7YztwUaFHHpwM6QTUbqbKpfPvHIPGGH8mii1DOJ+y8OjehpBEl5J
bW3QYaeWp35gwp7b7ivVA5VGP2EAah3DMAMxzDULiNFIqd0H8NHH0xZ2D5BWrGqg
yh1DkNalXRfEluN8wv0DpZnSnNlbsYMeDTlqLeR7OuvLsfTEu+cl/eQbWa+d8Xze
cfxI/b1cqEOvxWHdN27sLDha1aicxB4rJXqPk8g8GyiFnN+DzTF5iGGwCBmEOsYU
Swl5p2afnsZyDvB0BXuPk60CNKGesc4j5udRBcDEtzEtq6c3A31MdS0o5EZr8i6I
/lioLrovONHeRAlOeXeYdo02f3b40nfD6biQVIgqvofppgF/idvs6bCZAgV15URs
kkZYlLC0Y1X/NzkLviyGkfZzr+RYHWo8ZHhxrZHJo1A9mGZGwVppahkv/IKh12gn
K5LT0cQIn4cPO8MEiGWFwJPp0xyyHLwfm/3L6ExKtpZkJ97LpLpjfr2LIggVFxT1
oIJtM8BK5JxZulPrbwmUxp243BDPY+nC8y/v+/YIwr7x7NWVE1OZau1sLcawGNYh
GX1pjNek+NgM8At89BXuJECqpvpVlfFAEBf4ManogZpqi5Y0z1GrFKFlvDJpijTM
QziaLbfr6ftDuZYFCF49Yt0qiMfG2o1caWnzSt1yv5q6nYd3cm/KpPNz8eftw5GX
S0j4sExPqaHXD3dxW0z5M4uR0jzxzn1cWHRTZ8kltAoQe+dONNpKm4Vf4TZ7Gwje
d43iEv6zoM7HP06XZ3vrQBZ9lcpOkOGwKswTIRmWOP7PamILJYqEVi4LLVVGIqHt
CiPw2/bszxiMTSRWS5FNcLvr1o3GO+Rf9CCoLqgVcn/YNVdAyUsSwh6OFlGyVp+v
orDO/P/5p+yJqEQh7UrdId4yIbQ3dXqcJUKwwLylhr14Lo1geO9H/J3ZwzD9U6OB
EqlUcjyRZ2bfQd60ZHIkL5V8VXqimMPqOLQpLZboW3dyA1WQk8x7flKXvfWv9x4y
qwlicMa8sK26osy4sjY9vYoJOJAitMvI/Xk3GUF3V9rGzQKahKl7Pzlk4mohq+bD
tCcMmYulLLrCMHKm5YVr70v7bY3o98uZzXwrpe6ZDf0=
`protect END_PROTECTED
