`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVgBUNYRvgiJJZNhJHFWfHa6kuESYRN/19DZdi6VnojODzZ2B1ZZD4OVOOc8qKvo
yeyYsUl5IRpAkyLzkubJVc/5MZAfPERVfRMZea9oa9b3Ppx/yAbDR3c8BSjVxXwq
xixiye4W/zZqQ+fQ/+W1w9kR1COVNmrkLgzlwjAMwYOIG+wMsabyqDCeZet5zVSg
vuhhi8M+zkMfJyL2hfQc9o6CDmQhc4AHHpubUcCag7dG5pOEC8qFS/NhQLH/55QC
toW9Xd02XKXhZyBs80RIBihlo7lm3aW3SWoR2Qqo0IzdDJbxVCkNAyjyp2E6z1Ew
qbNw9IQTH7BY/QT91ap3eMBfxwSyovHgWamxlKWFsNaxfb9klPqz5pqsabRl0jh1
2Wzk0iHiTAEhi2BRAAKwo+RvGsIBloG7Hvyj2Z9baQ21Y5tOG6xX30aPQc2eWCRt
BIJoYSG+BfWKmFCQWhoeBapNBt8s+Nb5vR+q8gfw5KMbEElCHWm8VGWipY0TJW7B
OGFW1EM16Y5WzEU63ta6xMYV7cknhKUREbf6xTAqCGkFA5GCLEaiM2l/QWkXdVXv
wh8iOw8jrb/5MJAgiDa3f/v+zbtYv7hZQFlJg13MEwefItU8OHnTQhV3nze3f1Ui
J+ZMkmwe1C+X9fXUHEw7F9GFo/scXOFgYPnSgBG4UWrUF8kAV5FoXC5qMu2uTXxu
PQEsIysGpp213ip+TWE2x8LROC+8QbN2qwE066ocCHmYQGvr07PO90guRQfJTw4X
8YHTsR98zN6Bu51TakKBWEV3OzXWmq0oZAjXIjFjpDdognomtPlO7GQ5FZzlztni
gmS1qoHQKn1N0WFoJoGnEaaddBZb6fyEWt8KWDMq4bbvNV/pgMpxgsQo4KzRUxJL
F1c271gi9jmg+Jz7Vlnb7wdvQCyv0HohWjxkYpn45Wnxm6+mQlAH0gHtD/xJmAFf
KFP9/zCtzyr86azl6nZ9DA3iEKXctBc8DQS+BQDbF0cM4pwr6ZZuRX5TNuHdkbnw
brb2SrV1eeHz3jocWluGfnN9iYNu/X5NCYlg80TROgi9uDhljF5cQRStSZGrFQqh
jssxwITEmAoVkWN5I/6dX/8lxC4pEAR60M0UNX7rwKXf+Zk3yly9NVS1SiuPlw8Q
BDKhBsUMeLUv+vmA4E+WWXaE5OyzT70aV8QLmrOUjhy/K/iO2Gw+WS0g4ovPeaU6
Nm1i1TUKbrhQbFE2sydnALg/KIUdZguCpB6uoO6TMvK61rGJ1V0qEk78HPI6X8+M
BoRux6cD9eO6eWpmwBy83asv898LwgSc/RXYxYVdjeerExS0obab0A5hNZ/x+PcG
oYKyrMRBZJTFje0Z01qzPaqT2031ONR2RAWT5wDE5fYjAaw/ti1F89Le1ojL6tEZ
vz7t30utyp4ADarldwgwIqhFY6kqOSLOToYqYudV1efm0wt7Tqznmz8Sqdub1vP8
h+EgETQ0eb1k7AFCmy7hVE8Nmvqc1u9DBFhSdVKpnOSa0qSuQPJAyvyQOQEgM5EP
C60hXX2kho9kuMRxBRYrrXNLDG8+pkuXxih5s780nfzo/wwZhZR/UBCDYT9rcFRq
lwIjTfF465+J3e4pdcpkeUFl7L3t/mIJwScZZNPrxFfOZX1AZMnTGIDPKtQsG+aO
sIbdgNagLBZDaAXE2FbfrfjmBqB4eydAMfEbTB2yBUfk4C26jPZxMOYBsyr8MXO1
uvrw7YntpPoT1uOgSS+osgRXmSUitNTbtJpONtwIFGEuE74B6ndXoJ7RASMaInrd
zGYTajuA/217EomxDQ2oFlM01NymHl/NcLjdvLAxkjCyIb5gfzq8EvHmVImyAqvg
X5/K3ASTh02KKCraPHw/PM4P9mH9zRv114iqJ01v8WEhz4yFEu+xQpFUoKjN2BDs
T1GxZzYzvNTYeY6ndFhKpHakxYC95HTGocRohlBssVECR2/tisdMXV6hId6FkslD
l0CS1qr4T8Neaf9urf/Yy81/lL34EJo5+cWxz+VMmul3zgzeIUhn4nGaSRfNQOkD
/IBzh2D1Rq/IpFqKld9+PJQ54OTGz+vkT3GrJGLgwEIwkY12ecxX+SY+7dStUQ0B
F7rTMy1K7QKTBlO5HQKX61k1Ir56ZgSm6fkiDV+7YV2HtA/jCHHeUx4kRKiQvBs/
o2+lA3EOiBGN7STyDrIpLqraVrEpyemNaebfP/Y9hgEFeq6fQpUTo+GRnXQ0xDQa
phhyqFR3H3coEbghKZqUyy10hFZAVNGOKTORTlKoSbiccXhAA+zz0DQZkOsufA4P
Jj0SwpFI2y7M2K//tqX+C2z1TNg4f2ghGCUz74IRa7S9AD13mG7U5RVUQCwyHGdv
QB2HKaTF7wNrxK51RTacfn4pt88yRE1Rn7hSioE8H5oufTn72EAbIYXePzI+3W+U
lwDe76QR6D2aJf+2k7ysQTT6aRKYUjKidRPvWsRH5hewcXV/E2+A1NpZI/j3rXH5
qWrFz8elSFEg2nZmeutUwNNjbY8U8ShAWkbIqx8zVTqxDYfi4tLNGL1+81Myyltt
/4vvJAmo7eurYaYOdg6tzTaP0TfbDA3iweI2REYB7l7ZL4v9cUj5cYQBd0mcXdGP
XZX4/ujvrKAzwOw0huaP4ANhmgIIHcHAompNgiWQvxvpPUt+WjfwMSJi5HJLR5bx
LutNBv8ZnFBVwJb0kaakTs5+h2+YIjywIimunAA3MdGPiRzK1d4DPCYcQ4pluIr0
TrUjm1FVh6TTzwyKR3AOPM8rYU+Ufo6SCYVyjio77AEgWAd0f10V0b9bYuwEtKQC
0g36kxXMzidNdBgL56XLvEBJk4DcfFILYdNKfnVQAqDnj+xfa7RDAOFN68v4lOGk
pTOdx9QC2Yy49UI0it3thi2zTBja5Fj8rP8hrRqufLJ5lvY6hgThfA6mNk+q1CFA
IRP5Z8OuhlF4sRdhsV3GI/6QSXjVxTtVQIU7P2FzL4cwJf+4vgHovyXV0S2ep8/t
RkUvk1ITejqJqp32LZDavTtuR1K3K2jXbnaSbOo7NaNFVvj3H+RbZO1pu/boBRgd
SASoFl8ODdrKhfzt41+5qhoSJ8goVSry7mBwlKVDGTO2UZqqF0/6RQlsODC3aA46
wHM0iWqVvBiKzt1QhCApT98reHJF14lbInB5nm72rlM4l9NSJ4XPR7+Y4ddsb1Mw
mbym3S0YNMvF6lU5dSvQFlgFzAPEtpWJt/87Ia1UmjRyyiOBtfRSaPRhuEeQZbpB
PSZZDUUUy203CFb6qXLh5y/ioERnWYI7iQLyvC6+4y7RVRT73Wq17V6afBsOySdo
TIbaUUf1fOeGDlcAHUthf35m2aoFc+GM1eTYGirwc8sQYP7QKjvx7lh3ldMvsgIC
6xab0xKnxdrBwmO6LF5npsoBV9VWHGKnk0+Ifykj7VLya5VmhPQpMjXpVAeXY8rT
vNU0Q6wRfavMwCD8WvMIiTZ+6tOrbIO7FfjTMMrOG56e7cIONrId/gv9oNTvAlML
k/KQlehbvLna6KHqftLMVR+Jz4KZxIL5jsUWUVuBJzUNpxkquzdTepHxudCL/bng
G/YmFUA25iIp9iHhcn0LYFo6h1gLNZwhLxvJ1PMX8XB179sYauAmd4YZ9IGPuA4A
zG6Yqd915BD/yCjPtPvCbzPbVoSD0iFx71XF9qknMQJfM/5+cf7RWOSe4T/cZ6Gz
0pSm1uLPvVj5zL7hdiczHIkfrQGRHhwYwdPrXY9V3AKRH0015tDd0G1+ZXmMqP3g
XsoonlwQgoZX4CM1214Vf0KZlkwrFOwrt+CCpn60RK3s23nGbhsz4AxiDkSKxKba
J2glQ26EMC1lYswc3RTHtg==
`protect END_PROTECTED
