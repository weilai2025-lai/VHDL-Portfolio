`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTeVfOHVn2LfyBV3q1wksql2nHERVyteEGyGZ6bM9SZ8dX40yFu/8BDJKLjtzbVS
E+9EkMRZAU/CrfZjc/2BLuGadwC1nrI5LrPyZ2XqsMf0hAgF8o3dFOcw8pckLBVH
vK9t9nFlq6RC9Z23tmPYwQPZ0ab/HDndNvIi8ta6mw1ZdVx1A0SNhSfPEnuCZaln
OThBp6NCDhA4jwR1gR240MJuTvAcjNh4CgyCTDxgfWwJ9dfuZ7pnKOWUYHE8CIAc
oNBeGHfaFOrsiXa5pPDeV6nuD2OAgTgjBZLlf+p2bTWX3crgR6IoZsHoJckEFxLZ
YJSiuaX71CKzDky1wxHUoZT5psMsrWm0MYmEFG7uE798uXoZVoGBQaWd2PSjO/LS
cuPKCoth3G90svks0QX9IVyAIkULcPaRIHioQmQKcaIJZPim76V7tjgQIGu7gyQz
gGdQbml5PWzFKGm03ksoO25YIM0exdUAsnfVcy3XKN7IRW56iZvNE4PuU2bqfF7R
bA/i1EST7x9FHogkjAu2/F89PU5uEzLn1Z3XbquI4JGGUxAa13HRvDIx+zYDI/hM
M65s1f7Vn4zKE841+9M8c0JLgoHNytpNALahLOoMQsDUNNZGd90hN0XdPmcCRYYn
3yYOGNmOl3AKkxIZPFN2Tmql8Y/EXpVKI0yhAD4iH8Fg2wExqiaOz4dxluC9lYAU
sgEhC53zs7advZ/gVgicTLx7YV+bJci3rkI6UiylEss3fB2nxVPfMO/6ci2aDqdJ
1Up23EhC3sMkzAgtN9T6cjCMr5kvAwO4guYniDvGhFHRMt0jy030jhPhQ46mMy9+
Um+LzsyeQfbFZeBjk2NDpIKWcUqoQBUCtlS/4FtOy8694HMoudauJ7PD5zK4iKmU
3Nu7Tjj2kCE1iTF96U+GjvPD6NvIyGP6opQdXzH4LL85ERdrM4QqC2xzMUY1IOxB
t5IkP8FGaqTNYhp6IDRhUdnm9dEZYdNhCJuMOxKScYo8satSRDE316RnmMnPU6KN
xdLseb4oUm/rJros3Lc3HCVdk81o7RhM2UomVq4kGy+EevJUe5yzAH99lw+HzjXl
9NY4Jl4aWquKON7GXBMsNJdPqIZYF5R1opWjuJRfjNob/g2ZnJHwhe8VHf/yWaX5
3oo9c71CpeI/WOyl5r1uK0Loob4he5AIScwXjBesc3tQBDbC8mDwQOwvNrfbKHgT
YjvHxQTccpzQzFdTYkLMZpHNMPDG0Woubys2AdY85IaCPvmh/m6BLEMC+as69RiU
vYfy1ICDVLO8yWabZ+uFrBE2bRcWL4O4ARPmVlc12Sfgvi9nM9rpU92hjHLXCfwt
cs4LlJFkFb/ubhc4yO59DpUyyWmDCBcwpNUxh8MKCDhYjBO7NjZ7dbYODTjtOCSP
u+0iR+MVxIdNVyWfFk8AQvQd6TBdmAhFdfIgWni6NHJ7AdY/UAVi0k4oCLjRtYTE
RtzBqxVTZIvAesdd41RMDWDZJMpEUO8ihSUpiLjlsiEP2wPRl8yu0EhxV36h/8pn
OSRPklVnAf7rP2HxOOl9+OLCo2OOh9P9BfgSBf669nf4h//0Wecb/BW8tRhNNPMG
wkOZ/DQdol2KyKz6dNRiny6XG/8hZrNwJHn2qko7ECfqbA8RjmDbFmOj2VQBoQPu
MchwE8AomDJQPv7kWIeAk6sJDjqoXQp5Xwc57o88TsFf2jXTHnIcrzPbJo7i9Qpv
rCiz91BFZIdAIe12GMEZn39Oer6mS9QnwM6aEMxE9EO5+yRPSFfO4z0T4pCHIn9t
6ZSdLG1qeXZCHsoJ2tQa48lAz7o9O9fASLyuZtMpxULBoIt1zKOPd3Fy8umgklri
XDM72AKMkAi7r8F2fahC4jtmeLVRUYzhaxG3rg1WIlIrKdvnIQwx8vV7FAtFWa9E
XnaGsi55B5xUTmiOG/T/plP3rMCpCekLVSV6Br4muXKSE9uEmVXGyINRgFnKeQsm
JwdE7hyMnxAOZLC3oOQImEzg0OihzzGhod2AGZsc+Aqb9fMnfpH5Ysoe4AowwB7K
51hGKU2mSJ8a1Y2Yz+ibVBEThU+PWVtfxuMzdJQIMAvbXRfrV2UxbhxH0bL8N7pO
CNDyqahDz4w5+Z9ltJN5amBn5W+P+QXWjjLfZW6Jv2wg9iwy+3Uq98SNR4CTZ3zz
Q7h/sqjduIcYR7c8iJuwGJP9ZOfk99FNaMsRS85kxqU30DhtFI4F0A/jgc5l9WTY
/ixs0VDzsPAYK+WgXbPr2x/temOBqm/SmJfwNJGq6bAI/n45O1JzWTQ1L+WHgRi3
eIeqwAnEJfHvswOEU17Lmz4iGRaUpCVF07yGNZEmVLkgo0KH7dZM0eaBTJxySSmq
DQsnMVy4iL2v09XbQE76OfynN2LLsiW42VTKCg9suSAE/Tgy2urDEqqHl2ITSE4T
Q69kziGKZgQuF/zjriY8S1HHid61pKpq+s6w4/gGfUW9yqkvLRzp0gjUWXXy+nLh
XdtYezp+bJBahNS98InB92Q6hH23pEixg8kGnd6LzgZ5Mg6hi5A1Iz2G8jyqUl54
EpyiVwkvAtaa0de3fPUtojUy9bnG5KtonuemNJ2hkfdNw1RybNxVhCirY5cGE1Ys
BJUAuQsPf1P9y7msbZimxD37180ZKwNRTwEh71fyNfZJBLqjqxShKultKRweV1Bx
D29S5UwUctJHNT63kk8wSyiN1yTlviSXckG1GKtiQsy4kkk2U6nTin7bJ9+COj9Y
65XURXprb/SYTulSbWwoKlQ9aGKJJHo4GeesAQONYAws5UzZUVTXd9cfB9/N170D
Hj0zuIv1lqH9aUcSMGHSiqso2bYEN0hVmyZubSAl+QUTSkLtG/FsL9UndEc9yoep
V4ykIBT/SbvU02r1j499fo94JKup+7oia0TMEmM14MqS029o3OrSJrr3TjujbbDX
L+saYuOAL+w7eFjtXQ5MGX/AVzd7MAa3uTlYVcxg7k1QCtCEgKu/+2x14pbnsU/H
apLCVjYZXnFWJlpubaux0PfAFvcxLWLs/x1MwpyQyL5puU8jyQYrLma43y3V/rcI
KxnNG71ZZ5FPUGCofhF3xvanhGVLai65Jz0p7MfXy/EKkk6J0Yv7XA/HsPFe6EHL
ZvFjFTKHlK3LkD0djhpGGUepWs2aHay5Nwd813ZjX+SzAk7eIqINqJV85DiduTdM
iwoo+TZNw0MwxvRHxJM+Wg10GsQROeY+j/X377KdJWYVtvX7wPVgZSi6cOcYghgk
OrvLCzQCtLBqRhSiaqgdc0g3zZ/GBc6LBM08iSv3qGcflzV50KuJqlduCJzJwTyb
9mi9XYSXAdSLdNkLtU5GblFLJxhlw8tH6liEIR8tVjePtanU1iR/hueSzc267YcC
Bc8ZNEoxlWbqq6hGlmEO56GSWTNge8YM+g+FU9PQiombAa+TbBmBC7tPoDzE/etU
5OMsonD1bbBeL+tg4nqw6YnRVGEMuRz8L3PIZVMj/i0W/Q1KsSsCD54RaxPW/+CP
FyfzcBB/ByZ0nKOdJcN/eL8HIG0I/oUGxapNuZtMAOtxTonGyq2NFQOY1AHxRuSO
0IfaxoH4IlB0cCGk20BRlg0RxXsTFyswqZVf7v7NwsKlDB5Rl5sYFwzwsWebfBGl
TALWbdM0wEw0WBvxUxjVWSFoDmTKJ8+CReYbCZml1QLUKZo2/SDJbFXcx1W7RUuZ
K3cOSPxUynx+24/Atqmu05mOuPR3+fHHWW1TJaaywiPsoaB2PbPE2kbBPc9eWm0W
qK3JsKT7oSqZgBp7G95idGETZkRUxuKOWAOgX0UL+N9fHUXPBTPs0tU3cQSk3Ooo
oQSo2dhDpQP7KNpdgRZiaOTZ0EyYbxgjySbdN2HqTyBos/qSmMBNnkjAWfKxP3vQ
Y5TYXrB7vqj1ePK2Qda0Zu0Y/UB/VhQN9n+Z668lQYtNEfn74W/iBrTEyq2EFw03
LmucnpW+YzJEniME9Sqhe+ILw/XKHZPhlEx76XLWsng+5uHoippW57fwQLj3Etxy
wf6SXCfbB+DEemxCzWXKHCpM4lTMZFLD1SdEvMTXnZuHlcuEpZpwXmCaLv7uj0t9
N9K276xulDF/W8XpKxX80+AomB6l42wshZ0WhdfiLPqmhFTEOn+tw6xpM4ZjqVLA
w7Ezv0UFR/G3bUpBSHSfflX0hIEHDsi9H2eo7wiUfOAFdR4oXpIDqLP8obq2mu7T
vEU0k92UMLH0RXpvl0JFymd0GXopLoFAJD+4z4Do9+I5AS/V0SqbM6hEqpQdw5Cc
ClKBDHIBnqunIHELY5frKelVcqB+qcTj2hcfApInM5BrFLazFjMUEO76PTH4hbFX
N8ZF2dnV5xKP+k0lcsVjY2AMpQbvEHV0epfQv7Y/4cqU3Ik+Bt4AMFr9yaAzLNT5
bbEQ6hLNs2GM/wMFRTYcLU9MBlfvOVU1jgqcFYLaNEvPSugn7Gj2QQl2gEW5YISr
c5AEJWuER/lO3fDyt9y5T4rQi1b8ywGAE+4m+FgjnUmlGZLZI4iv/G/ZptWneJXi
cHBhY4ThBmrj5dogILWPeE2UZwRaDc3QV2U0wtQL6j/CZaQ+Xgwut76vDGXvDRbF
bREjT7eK9NBVSyBAdtNSbvQTIO8DPQxLEZCyux0iAym1Zf4rH+Te+DtN6eAHetor
l+h4kEyLLKaeIOh+5rIIIr0eiRG4WFQTrQZfFyCGr4IYPdxBlieMCsgizGBAoCdE
JwhZ2bxCfAW0Tijr2BNHpz3zXqrG0FfCt3CITLLxdzZ72KgV/1Hj4sj66O005Cb7
9WC5+RdocDByWz/Y7a+TcRVo7UkJMtMujwI2De+MISkn41YJ88/q6iGMmp+8JnH6
qeVmmZ1HwQKYe1yoLtRic3aQcBRmw1mfC41DROuqpuQb4SLOmHWzzN7/A6tlL9D5
bePaS58pBSeZ39XJ7YSu6xocYFv+oCf5OWNvOhq3q5lNWIHh7+poAPK+3mCovysY
qjrbjGF3g9hIq9L2KuIuL0bNuh6Z37aCw2jSqn1L9Fgc0CWgCvh43Y9Q9zohIT7q
Gtk+NFzbKkTflTh5Vg4vwULR7yZpmPxK+XZPSl9BxrRDDVRNOVBb1+V4lmyndqW7
MhSiJm5KNusb6jRDWUVVA1tsgigB152KKjuJDSIUh4ODUwe02kVTI9yXdoIChHW9
wUUCO6ZCC4gNPkvjto4Zm+AKXIahKQUzxC4uVVx9dcc1gUydRAuc3rMg1AlXusSO
DS8XosgAXq9nzaqLQkCfT1UuNXzbpmdl+zsx0XpybyLHTYlGje2nMOz0YaizZDyO
hp79sWI0TWwoVf83UNxrBu+X6hAtfVynacI1fFjWIPtYeoXKAjuwNZBz5aGU8RsI
XusDhuZnzvLqr9pjp6oisDmj0X+946lHxCGdpuxv7PET2tKZ6ACWnIbVzTT1mo32
Bc5FvfZCKUs4d2kv0oggw2aNmS3yIloShVyY9v4uOSyWJh9StJX8MVpi+N0O4y3k
giNMrrO1BIaRLvhjgWpw88vILFIAZO2AN3hFjYnr3dQK7H1xVqRtSk6MCQ4Ie57W
4DRo1ou5jcBVeuVxdWP/ab3Zt6iXhXJuLhkSqNY8SsDaqgi81PiS9a2RE6PyGzHm
rIGxQjdiB75BjqZSGhkw/L7RWF0i22JVrVdKn7TOvP8BMRQ9nTfcNwuzrPo9kwvC
Z3uBjtzD9GS+omICL9hMoZAFxIpdXrdDgIM4+oiSjmIGmGVhoShYliuA0ZE0RZnh
OySIr/k9pJ/M697FJB5W0N7iUXIAOv316yjJX0XrmobCwSxAqTxFPKBwejUiYz0T
zASuESSCIiwEQOM2k/unKEWAUybpm5WKGzId9x/iUu6ix35mKIgOKwTRBZUXPJem
8qum+2OK1hAT/rmQFTLTPs7Eis65Z5dkl3XUTZtKks1QLjfomBzXegD7iz6Bi/J/
0BEzkbgIm4lfoWNa9DFFigrtjx0TgM7JLMG0zAtkqvP3KvimenxOpLddZ5hWgUHC
zYgV+X1pGq45paO3538Q7shAH3zTdsroFlDDcfA68WcrV/Udbt6qUQEkq3f/zl/0
lxxsWahNeb9nSTzO/pz7U36Gz5gortTdzhzNGwesFuFqlMWyN50R35pvayIqTUax
R+Mxd7NTVcWGMJRuoBdkoKB93QUJmEDzn1P6nBuA4goyZTkiAQRtgk5nAztjY6+J
a7Wx859H6oiGBT4LHh55Y7bGHGJRO9yTpMNH+4uMaBpjIRWOLdZgKkZUsIEwPA98
sfwb7SbhQPixDj+N3oRE18PbkGMfcBqmy1LH5pRGyh2TMwv3joVGMnSVmP3ebcNe
b2SzQIbs1r74Y4Q2zQELQG6OZDTQZs1GInB8VsQHiKiIEtxEiIqbU/t+WvsE0u9J
D1Gz/0UZBPBM48T0Odwhb8IbjROK30odM1L0DCLHamv8LPA12jbuf8eGcgff6IXM
oNBwjHT2T6ga7b1L9Od+3egb8g5wL+fuy1F7bjYaojyBMg8Yx9fYOLQ/Nq0S5JUE
jRFsY14knizKfaTZETU4fwEHVRHwd+bkusSsdMzncHBBbgH9JKp3/Jq+R0656sMg
s93Skp9Z2u0ZGVkgsTk+PtyQc6ZEo5ca0r3K7h6bKR+3CnkUtz7g3tU85jpFVFdg
NIASxXX0sIt5CfL93glppotZaVSuUBhu7UWQM6FSnJi1DZIJ+fHeVdEuCgEUQoox
qu5/9BzEon/VTKvPEQ0LLovjUsa89ti+L7YkZ9+5V9rfOv/g2F4JbxwceO4elG2c
taLg8Nnd3OpmPRvihxkqeNFZq0KxlAoGgqmYo9IF4yRpt7y6lWGbm7eS6/IoXQRx
efgczvrJ9PjCU+AqmpucS8sNFe3YWm4KSPOQwwtkFvSLGnGUpTKXw/p2wJd8zHRe
rBDO/BDJHUEQrzZAN6x5WdIiw3++KZAgpggyPUO97DdvdOXNnzASutf5HNWjx3L8
3Du7Plbr8vgDzfZpo9d+TUzF+TAkIoTJ8bnWE5Z2Lb/u4eLPxTkdnbKyji4almr9
j73a0Nva/xVJvsGxTQA32zdnU9wBH+473Q9IWmAsnEuYUyBpFTzSlfgJHXA2RhsW
z1VK6nevpeEcQuha0TAx4oB5UU9PYCvCcBfuT6TkrALkYCY98D33PKq5Oos2TaoT
qt6TydWyXZV202/F3hDDWYKx1FLLplLUJkOf06kYXofSAdFGincAI0tslVTbVRW+
24Bl3qSs/3n4t09CnnepsZH75TDU48ZnQkoneQrQsx+3kcVmfu4gJFht3i4nXfK3
X/PlXA0D6CVfToM6wJ0PDeJPVYLOsx+jcQ6FvJcJ5xT2D6ZHMe6iPpgToOhzr1k9
jpRMO/1O/D6++YRohx7VF8vkuok1qiBDlqaTmHuoB/Q19F2N0UUhWlOCS6jyrf5r
2r8uU4y6IQ38NmfCAof4NNvRPhlKtTO9p8agSN3HbypvYWoUTqHEWp1ya4AVShpc
z5NMP1I6/8bp4qYiLYXu3fiq5oK2NaKapR7rWOacuFJc+L57m3Cv5DRybHucSfzB
TMibWIu+7ZFlmF249ZRw5XzbG7z6dfwQ7JxBnvxuBG+dqaVKErMb29ihkOWeQg2S
ccbzjrLB1WDD7L5Xt0DSvXXmmZudyYQfdukZjj2lRkJPEKKVnvfvUM+owVKj5cBz
8Qri7jzllHajMkTzUVar4swr9O1fO/TrQL47FwWnQO/ktNY22azLA5XLDC2QMwV8
xWn2XZQXQIWtdRA5SHNY5sGjqf+CzEAz5iCi11Hall4MPhTwLFuQJP1e9ZMd2ARK
wWWd9ap8+2KbOM/zHrdKLtJdnnP8Vuy3mOqdjtClGPcvAK6wV2Kmov1dqz+hEE7P
UhmY+8JHjI0IP8oj7+lCP2YZEBM+Dj6nNOwhoWNNXuTX0wazu1D8aohA8Qzc4Ghn
7GjsHMhPaDTODdXsOJbZFdQtxQpBgwZ29s1EMlLrdP0BbHK3c/KC5h6Rh5yh2wVC
MlUhT6lyKAFs6d/0xSqjS3OIda9cbhQRWt/5Tz/v4uEfagvxJ+3bMNtk1vmpPQ6m
5oiz7zRt/Okj444JrzXbDVH5CnEWYnBfI4MHw8paeyZ9shSVc8vWyz0vPPeqWKmR
vUCJ9paiTAaeLufwTo0OgETjqd2Lvoeuc0mMHbcXWRDzYkVuHYJYsWUTrfGe1AZv
Ih7d7BigtkPOKiTwSNk4Ya5hoQrGRPzjxSVXswINtn76Ka33GAba4vVaP8pUTDmH
VYM6cKl/U+MAATyYY8WwMyk5bscfVY1zjdIuRcWplVO+NedKABsRriBZsmgBSRnP
xFRNBDlTq9cGs1qqc1IqrhCmX4cG3efxlRDmiz4e3vGT/ORRbCe20c7IDOfYsfd/
yzCis9Uj6HyCAesz4kg5cHgciqFHMZkC+aAJLsh0nFKgL4ETIFsA1uGcO5mts1xx
VZ4hzMqLKwR5Lmdm5LcuoLueKBYOonxAUGzxg5swpuFv62JNzf1UbuW/qCPHfsSh
oopdj+7vkrzkkHCvkxBIDPSBD4tAS58EaE5eStdFYuEStOaI+hy/acjiI0knKHrx
HsbOL438Qw+KByHPsS4LaoBBV79WhK+yrqXYx1KX53+zpuVuTBnjDSg6IwyhejuA
bGMXQb5jCkVkcBSfAUYNXeNm+vD9HhFd8UnEDUVBeNax7JfhD1KwRR9yPOyM9Y2o
Z7OOhJs5gK56ag43CBU23W15aAn8lhT5e+w8VFltpRjUJcV2TmJO0GhqqoE4evQt
jR8WSel1TfdB//5oIRdIX6zDldlkw0/SzJSRmi3YnKEq7EBP44RkXjRoBCZ0o2sP
exmeTZ/ulqxufPpS6vtThlyItq3p7Df/lxm+ogfGcq9ZVP/S/i9CceejNnmiUHaQ
cke3KFHAS9tl90xWg0CASsmIUVqUZ+j55jcde4UQAI0AbPlaU6jHfKGAuvZXTt2h
vo/WPl0r0WtUIXkTsoPE3jiLMIyK6SFQgoF/K0W5h6cs/ej9aiUkz5f7U1wf/ga4
z7U+TlA7U+D39APlT8tdRmJxL0khTuHhGuj0DEjlWGylLYaSWubMb6UIFhWaf3py
FwQEAhSSnEB6OpkdnUzCMd3lrO9utbAWBeSEo6q0o5vfm/X6cDSuBDdgC73HTXW0
1Wf+L0Jih7wNfEPV5GrLv/9C3LUDmDJiii5IrDfshp8hesH6lT1umRsQrl2cJk5f
pU9up46Y/r010lKCzckeM45DTW+AhxzP2fV2EK5WSzB2AOci94sPj5R9VhxwIS2l
g/vc6Me2h9E0oEjkhoCSwBmV9BDQM01MWmjNBrUADH5tkckhY5tGnz6zwvp4aZr+
hyVFkwSMZ7CDsLVA2eI6zJ/VwFOwbd6b9gDsKnjUjiJ6MSo3nG6h/Gnos1rZzILt
XULOuds9mVUBp3MBLEKfJYL+G6M95R+r9s3af6oSmuxIXsS5DJk9qNR1ftBz8W7E
SFqGhXsYxVEIfo1XPmsgQkCHXNKSMg4tZYj0MUKNfRPggzZzfNpVFvYXoZhrR7Oh
6hXvb5j/HjJvV04LJkg9Mf9IdPC7aLakEvobcOLiPc9MPxtIkcuoJYtN2hhGAZVo
hN4dbWqsHrPpe87Xp6g9F8dEX1i8nw+rZBuqQQxuwGi1b+ZfdblLYDdi2DC3TM+1
JdSj5FS6ep0PPYo8vmkvoFEUnSRfSrtTV3QXGGt1E1nwuY+V9+arY4c4tyrh8xxI
uRAl/upOf5Yhca3k4bKm+UsDGkGGe53d5/ERuCQrBj0WCA6KD63oMyh3nG76epw6
cWR9DznvS83q2n/qybyRaJ6RjVS3qOoiwkPKKCp1w76GBUtBWBREI9Cq7HELUBX5
GXsIssuUmgrh7ZQmnCDptXrtouOub5pninKsb1Vx8+wlXjvF9+njGxvaKs4JbpWD
74B9X7Y8Oyx+28wBxfOIvB2xmX0hsuXTVr8mCvb6CYZS8nI4Sw5tsxf6iMI+pZ5X
WmQyrkPh5Uu8xfe5Esd+KoPEGGjNcMGm5PRso/vOBlSyRM32HuP+N8duakuUwj0R
Bmx6L5pdKi/SATkGqteNr/V5vm6MARbqf2pxBA7bXuhadoUeI/hs+QBZ/sZg55YS
KD6Xu+2ufMNPseEDy2Q0fwRr4t1UtX1aGgVYyOk1eQPKZO2YtS16K2rT5Rbi6Eoo
M0SQWdh88MsTjQafo3OA+v9cwjOw3xwcykIAEqLCiJSgPWA55kEbAAu0lEjgjzmH
FYqcN8TeTcHIvayeD5O93E1hHb8/WViayBS1vbbUlGKQ9PMtwUcHxl+4pMxXnSPA
oBWc+Yy/36BgQfiL2gjal/HgHivQAB/3lbJbPqtSEFGi9jkF24bc97IqUx2CYBch
jiqZos2H0xRhWUMs1XmLvVyB11Onr289zYXOfuZpF/8mIo/LWxFj7HGqQxDOCyOy
CGBTqm6PMtCEmnRaGpgUh1KYo71s21sphnyULpJQ4NWhdd1N9AaRFoC1z0U6Po2Y
AebQfdM5++nPXz0mk5hlvLUZXRjIhq2JABRHiOohkn+0vPUN1FkFlPWnQga3gBlh
/3P1Mp+TSZeu2nHEk2sVX2UJ8Jze/l4I/DIStvaMPVeQb71vJZKiYrf5Vec7LwuA
pOvLMRQBiYrjKl07IHadFtmkwt3vXmTLj+QSVUtc3xa6yW7OBVnNHHlc8pHifM4U
QzQqUPocJIN4vtEgWxdlFclZXGfo68oFdS8HIbqsYl4Vkv9xAgTlLAZW8YUF8aUE
MyCxQGH0ixxYglk9VR+vJu0fO1NFcNZhOm4WPZ1unpWVmzYuCdpBBZhVhINx4I28
3xJ/UxJoUw8yBJqtBU0ENGW0zfE+0wccnjI/et3nF0SzkAxvxJ9MZ8uthzK3wCPy
TyDAp7hs49qpNCj6WcMNfo8zr1QQWh0U8HxZIUazZHJU+t6rbX3kbrAys+Wd272h
1hpl72/lw9psfBL41+PnBN4srQUPuB9a0yK1atcF3/W24DPMpOtgdol8c5By4OBf
XhkKN7Wmzqx4SuXK2R4iBOSn851/4HzSTw8mhxo7NgQWv6ShVrSEhTtENk9F+hRo
1pnCt3Na+9sjlPi7aWSla5DBbVE2YQGDcM5m4Pr1qGhCV3uz390VIO9Zj78VdIId
AgPODQTR/M10PdUNls9lAsEdmiEe6mlKq9eZXTUweRzir3Zm/PwnbKJJGUyR1YZf
AqFvvlXRYGyu0axljYm2ZEddcGw/LPUsK+VyKhvXe//rr9JEQOL25saaTRDX2VPw
vRYDW6ZUZILTgGvTGI27YTPjv2bI9OpxOT1QDcgjd6PJdRYoijGsK0wEj38eBtOt
3ChXTwz3xO2gG8jkFE8gqW3NqH2DucdL4fjIljdknLed4cN6a4Gh4frnYvW2ZTBg
2UFBqfHAKgLV9HcvctFLwVdOWJ8tpm8OVQIcnmmrBkKyy9hVXZCMqVTPUtwOHYcx
wWMu+dtEli3BhSHBnjECHpWj02FBzicffv9ETOqxXkBp6v+k1lW8ur06roEQ4Oy/
feYHU2xy2R7Y6BKXTW46FMUyln27lHzh9LVRaFLJlKgohMrHclTcrhq4oi2kbk7N
JSWJwLDQmED1ZretvtRnR7G6u2TF+cvFsTtRi+M7HBviB89T5DgmJSwGHIQsATGT
zPQ0LGvPlb3Es3hCrJRQvWH9RzDMl+2C5U+tIiDN9a3zlRaU8bGwjzVQG9cvFYlf
OzRGldyitqDoqA3RXY4DUwl5nFEm+1xbg2l7O1Twb+5xLrv34BAgVykPmDnLt3p0
Rm9a/kD9qlvJ1lOSZqGYbNkDmpXvo3ozQGdmn+0tMcMbUV8zy/98aFp2g8N4ISsQ
wt/hsD7MAxB8+UFDCZvfCkazuWT2kvJdoGANF1o3597c8Ggl8B/dOzXzJWXXCPTJ
vqy3kfHbpGLO4NmSllFlL4mO7Oyca97wM5Co8qyoBkYcECGmsXwaivDVmAn0uf9E
IMyuNxVwMkv1aaCwBvL0sauw5h7XSbLmv/XZXt/KzmDo4nG7iNu+M4HFAomBidqW
cbVJuYSwGYih8WSF5tuhpGqlUZOjK3lyRmSqr/24PT5Kh2GOIsgZhqEScvX9Q3Pl
CkTYPE26wE/yUYWq8WAroIjJBh3sYmsv1WR+uxTv4CuRyUMmSSVO5zeUOAjbR6ET
skKMAob+Ie1YoRBp0ROnghgVkTDLjYaIGpvaUQ1vqlQ/nZYeotjhdHSz9h4MaA7b
aaPosQ+RZ2K8yU5G+pNSffNSl0XJDlNfwPTg9TiJjshSrbpgtWQ9xi0aW/BhPx6j
/x3u7GfweTQrMCxlEI8kna15VQwLXFNxDwLNTRWR8AMaSaE6jFqK0i57vA0Q9Exc
qTCRZAesTn8/2+s3NRezJ2htxa9JrxJz5xim1d4QdrNawbWeQQNw4FMKxEIEPePY
y/3/OSEv/iOLjbN8VQNxczwt1THA+iOoDA/tVMHjwA0nbPW6G7N0iLSBlyrX5i9F
JP9P0Mdvwk4kbrXe+IGi5oJbz3v5S9Up5PMJJ+Mqd6RnIkDJ1OvMBqJtn6vLCOgU
VcqIJCR/H7EJp6gFjNle2sj0eJ7dy1dMVlFmCz+4xfdt8MrIs2AbhUdhyp/o8Nk1
16KJlwD6HUDjSQsjEEMsEOMCJqxyJwgNFsUxnk8EX4XssMujruGDMTov59HZ20ui
hXbH6x8/15kRYQ6YmezgWIu7o2EbPP3PoJ+Ds0rNMOx546XuCy26Dctdj241bFoK
h3pA8YpoV95v1QXocKOaVoZ3K7+rVrjcK9FBI0yzBsBo6blL/6XO2orXGxOsTSnk
m6PuopvrQ/RXZ3fsdcT3qxja0L8s0qXkywviDB+dI+dhGSPl7CXrAFHkT+JcvnQE
ZsQQjg25QcdwrAZI210bRp7507hUcocFa4FiugolD0GJOw23wPw4gvNBcBkAvZGZ
JNtcOJVHlEaagETY3n1jE32IAD5FhPUPW3W8mBdQqsxujC+UmovdlI6O01F9lXpQ
7NXwa7IuiuJykTHOs0lz+K18wazsSUy948NEvtk6lqfceOyo0w8N6TqpYWjN+6PC
8B7BktgjZ7Lutp5qZdU2QyjrP+s4oitF5zrfbZZIxlJLesrdUeMJZRD5taPUudby
cxs+BtUG+zhScAHXGB+v7ysAhGgRvFoWWM4mNmW+MHhpxaiLrgTnxD51jB4/sW1z
LzB87W+x84EyCls7yd7uDHSk5rhJ4hPBtJ4U7smCBDbe1ieLP5p3cN/FYaSapqgR
ZmrOxxRLsUrpggzvD1VglEw3XdVkKFvl1mGe6N/wuefekMX2dgx1JJzKzoIvr5Or
Hj2sBSPLMeDj0USOSrS0I8skXps/+fsLmb1w9qPoRrgh8EtyYQs65DlY7sLKyuKI
/mlQorXyuGJN96US55iVaFP8/V7pYtlIt/XRGKm8eq8pbBiIyaBClOq99LgXv9wU
DQpO7gdYnedbGGJjoxdS5RcwG1ue4zQdVXAf6XUmVViQPSfTDGFF7sULz8frXW/7
FORekHDHqoIiYGxaElR2bz+DntYNlzjkVQVVjPETspLVJRRHPBEJVwvoMcI3JfgG
SpCaR9lCgRISy8dfGBzjsSAhLrPWaSmG/sMPC4SSVDjEZbmzgenMGavQnn0W7Za7
gpUie0dtk9gt1wTy1OMBcNUoTwjm+vChguTC3lW42eOTvdCfENOf2scENRKmfZGW
1ePhTDfwPdvg/hYkYYoDbeSVzhyp5o9EYStTRYlUpim/6QqPlryEl81FT+jFjNhB
pmUPgsNcBQpNJj+9DGysPEjfXiFrGXGz+teYTKZpjpZx6WGkYgpItPmpMA/NySmS
aIyVZ0lJhpcPqcAXdbpnnLUlbMKoLq3CuXxxz0pxr5dN2smG/m2tVMADJ9LvuZC9
WThnvqpLDuRR3MYSAsUSzQrFN1Ygld7Bm0r2K93CoXSizb1rS/ON8paGjC9WlTAI
9f30/wo95WTBDNIizUBdwzVZkHgLPRLSAqXKhm6Xu+/kNXt4ymGmEiOgQpiiosZi
i9EZu7Hkm+Lp9WueLfZi1PEvUooPDpesjc7oM54uBu4pLDKrBm8NYwonXCVruifW
TdpKBZ/K8Ta26EHOQDng5+rDiEYAh2ONk5ZgNR4n4Bn9Vq3ycbfXt0PX3QN8Uyau
n0UFwRPgF561JN3+5gZJGVKrCzX9EBS4OOC2U6GIP7Pp5hioivFlaweqv+hRbVWw
Qok0OVmABx7COvmH4vPwaKDoHfS8/APMN0fLZ6gyD3eJaIM526d0t3PPa1MQRpzp
xMQoTRIBEhCXT3MwHiOogfAe8rRuCStlyzBKCGvwc16uy0twdCV6xR0I5duBL8z2
1hQ0C0z9ScS7Uw+O61gTOIGPG+vXRlXM65WCA0JfdPttHob+UlTq6drleJ6oqRya
jLKHW/UbfHGyLd/YepSd192neMzMw1K/FCSCq/bNxQi+xfovJh7kF6/ALWJx8v/Z
6MX1L65ERvXML6QpRleEhW1cDYs0Ln99Z2GNj4GThcsYOUKac4S68WK2DG4AoXou
FnBOpNl5DZTeaHqAsqY5IuCJu0SvTPJ0wVe5hZoANSKlZiHmXlZOKuxoC7CbaiT/
ccBY6VeEVuZWQidT+tNYIlyPmbQGU6JUnj5TYzSEgJnEaOAWD8GMBh2WPTLp6FX8
9NT9mGDRHGd1UOfdwHtbjlm83aMdT8/nNCgJAhFU+nDK8Bt0JqeMMvvaHV1lA6Q8
EqhNpDsEFquc3dOfV1GNy0TwVom5QZF2hxxn906nt7bnnXg/qrg9RcFxbWsLr12J
AZpi/tKLwaHWI1dq564Gdd/ebXL9OZJ3/h9jsgSp/W8f9qe+3+ky8hDF1qJqV1Gp
RwJFCS7ByRK7Mjg36DP3hexyaPbrfJmV9jwVLyHsLY0SdsXslY/xYipJkLzHdhxT
sS7nHdKjJbU4r1ph7CYJZW82GpHusT3Ssy3JXgSlKFGYI7O96dwF5Wj23WXaL/Hy
h7XoFejTM1RXmLypg2uWkcCEgv8ISzsji4rJ2hXKZrBJEkfJhcbyD4yzyUXVXUcj
GJG3U35cfGbIgx0/9RBv8yDJqKx70Z5kkuVv6FUi6FviZpLbiJKvLYkv52a6006W
LEFmxVwNkq9Atg/lIWFb+ZRDn/SS+YpKlLTRGaD/pNrwEdMK/6EwqPZ/T28gR4wj
Y3PKENo8yz3DITd2mpizjaBLG+J/AAsQrQQNTTqchnOJH/4xZ2t7jqiNmWx+x8Bt
85W0x5Km+ZMl5UbaBHCT3AcXuW51GMLVUSDT9jnqvazP7p3h7HSzCQs1x/CgUoPQ
vQW+mdXF2s5NX37Fm0SodYXNyKSmV9QFyQmcbmIRBFvcW0LLl4cWLLI1mytJQ3Sj
YNLlq1mojAMMlJ2jmRmD97vvuxBMYZN2YZv7r81xZB6dJoYaIbJqlx6iRqLMua3c
qGneoe3E5xtzeQyWdwlrzCgjByvsl5Xtc36nMmo7dr6D84jDRcdFF5TddclSqeJb
vooN+ozytrRFbbLML5YHMzzNPYevChfwAzS7dedOpXMOGaMYTBsg3sU17Kd25rXv
YxRn/Ev/JN/iIZ6IG9qEjkW22QPYgY68QE9F0mtWl7L85V6CHAuA/TshMg2zcU9N
We4GSxOiurDiLTeoQNO1xRkOQJ7EDIjdJZLhS37lwb6tolnFtP2WFUarnfjQuchd
oEE48k8iBd9iQTOzTH8PdSX2KW6SAFaBMGoQRFXjRQuTQ+yhK1Ih3Aryi03dgeTn
PFb1317fa1R0toSGXor+6pQ5F2kQ/YbF/4J6gAC3+7o8eAKiO1oYMxqYQBGG9CYT
e85F7zl6hKcOqpIzv8tcWfN2xXeifhum8RIlp/5JJejiegKR8a6TlpIZSikbb1aF
FVFECb9eaq8zC8CC+vapec9esKAU/f8llyeaEj5loAZiLsnZG22JNwUVuOmwGVMp
MlP39awWOkHkbT8fhqlFRBnmtb+Z76p7lQrT/x3YvpagI9v2g1Y00NwYpP/1fetW
O2gHDmkAQr4BWbMQNb9ciLoFtzTwSjFo7okA6RNDkqrEKmcb5aJac5AS4WGIiB2d
gC6fbcopOrzpu/06jtQ3rkSoIX7qwhRlXtrY1o4EpGSluN4Xhr7sjeidfnpGnHlF
peiNJ7dSEhBtg8pscGowfPrlwf789oZIo+TgEqxpr8DAH7BIc1LCZ68swYv1oCjt
4H4dLCaiDMArANNIngmm09/QvVQLlfk6B+yQiKYoaDFO/nIAyMCU0W4tIPe12Wsd
sBvSE998cunUhfDQrjSMgLLNFUYskYb/VRRP0f7DEOx/Q73RcJVUgtDYsnectUoe
nYzikzVZBE3W68pJ3rcqIlO0RHagBUT9B+IP6Z+Se7qxoKsVhcyawkHyHxyJwkT8
kJ1yPW9bNRzxvc+M/WhNUPS8/2sRyVQzZorPxGR0WGlHRzRNG4G11bdcCLIBsfzi
oVLgkBnVJTfL+HjOx9IUbMXJJ1JoL5RQWtPKGKwm9AINbPAmvrJNgYA6Jp+EzqpQ
3vT582h7qJcO6JnoXn3zFLQWjR3OGR8Deet3vWFkfnxnG/NJ2x+Q7rJTq8GHABOU
whH/CbGJlQfETTTuWAhCN1/5leXCQCMa2U0WOohigu4Lr0xh73rnj0HAM0yIP/AJ
K+UA/pZIVydoMvPJ7J/AhZC+VPCjvtcEHODDNx9vPYyDtKIDMn9Ncm9bNIVXJt2N
H/AuRTUkAO19L2jzIIVtzxdfvKAgKAk6kfpPvoS6psEd7nHVp30q8T1s9an42x9J
Gory2veohrX1YyyjsTkdR6w/+Ljdmwl2v2CC01qODRYxkhoRYSoQ7kbaOa7urpEk
wyFFMgAaDQNDzsWq/c4/1RMHOPECmuAPfjnSeWQGD9yLbwXi1OyEZtWh1xz2iWxj
dFuflJ84xytMTS4v/sjdvMaJIubgCDaTeB3zIaiFbVU14h7x/f7kFMph/gefImPB
pto1oYRcK30b7ExdXJB/zZKjCJFU+9rjxBTf70s69uWtC/SoaK1zoS64HCVNB0D8
3HOUR9N108Hkajbgiudv881IMellUniZzj6Go4KUKLO6NvT9H6iujsH77uMYPTnd
NeXnlO9y01MpsWNJsN0PSjcfPdN4Pchps4YElynxEMV/tX9gyGnsqkPyH1wbv5KG
o7nnzqRDxjqIG126QgMRwaO9fAGJJg0UiWSTZdTHGw8HFFGHvKWazt7vkPk1hp+x
+WXTrib3dVKKqx5Osf657ifhrcPZVvpQrUqjrBt8bXx4o1Xf+QXEoVP6THruCFqv
CFghfFQOsMB9Ib/OOUP9zIxf8AlXg7czpyCu1EZOjoK1o4Pgu/EYP/n+KgHeFBgg
jgOeur5qmi3IHQdZV8acVdPjl9rriGIQwxz2B0wt/Etw7rnGa5fdKJ8zn2neoivF
a4L0p3luy3M+wu/ngpKpOnjVBdVwumdNymy6EdxfEeQYr5HMI3Mfz4AZzmh58fja
lx34UOKvMpTCu09l4PpaMhSTlcrafg2zD5ejrlNaRPku/IZ4X22nm4Se/XmO1iTj
ex2UX21Oxg+zpXozow3wF07Q76pMKh4vfsbViPZDV3Mquld8TkbKpszSUvrgRUQ/
oSme8lb7tJzx7E0OgL3Ox9nO/7BNrYcvY+qb7R5Nz1jVMEzgFz395XFKTDKB4Xd6
zDQZQz8X5t4CcmXrxYgONkc5Tuj1jcWyn5vJimtU/V+lKNnAYRfMHVGkGJYxz0dp
hx5MZsVLTxOm7T+EoO3x7XGKQhpjE13oVBL/fYiKAGJN1Wp90egWDo0M+Fc0Tukt
RdbRxNqCxY6WLl3NL0/EBOONyQS+/CwrMgdm/92Q0UQYsFFP26htXnXWTTl8UCz8
DG9UZGXmCu7/736Aw8H4SiTJQ7NPAzbzqREXXXNUfpZMB3g+USQ9Tth6zdy13Ane
BbICCm7PglnqS6K7/WeVXm3Nm564HT33un5kCGAgPI6Kgh1AKY+Et1BAfM0bQkaF
lIZCrPeuLBkB+jiRi1+hJL+Gu5ohgN71+64/cQJo8n+jKVC6OKxUjxvkEuHqN7JK
U80TJ1Vrw6L3KgRac8wBa7WI+jPKg8yLuqHmseVk3HpgTYhwm05c9aE7a95DHg5F
xCtkYSR5b3ZLygHlG7Xgji0VvFpXv1lGtSfMowTdv72BWBV2qdlwWtfZtufsvuHo
9bNVPNhExXyriIK0BVH+7PPqT4ajoZ3O+7ulZFqr+cd9x9sD9saX12UAdsgwYgH4
qAafM0DC1gDe/xH7VaaTvwyFKVS4UNaYkJbG78RakaLA0U07LgrGkZGdZBuquT+R
RMDkDv/VysgukMUsSLxnQWqk0TBUSPKgqL58fVMLtnTrrdRLBealqmovGxtGPtJ6
G8NgCE01crGKfHEdaw583jIS9iZmVK3KZ8R8tHL/LHyR2CDnRlHYk8uaqzVyLowI
rnX8r8RKAWybcrP0am0muq4cbDMu29XFlnlRsTtyiaazPd7QPjCAYnC1lPQBeF51
lZp2vBaXq1F/OwAfK+nu0RkmkDz3ufK+7tJ7HzXOsKNa8ncKjnKcTjq/t5/8WwgC
7FGSpPbGs4YiM6wEe/MvJtl9e3REx1/C2hcYwN5NUXEUZ+0Ny0jfZKkX4ONHuFxX
wsKzCD97x77Rad65ho2fZPcVgKgExMEVqBg8sKZLksoxIV4gTE+pEv0O0UIic4PB
qumR1quHcDgAM7L81PSdGsXIQQh8DZwAORS59OBT1Pe3V7AHCWnymF2hMdVtg+WJ
Kfds+9vBuX0WCGRtrmZT8Qq5n7wKyHbQNuBPzaWLjl4W74xV/RRVqqfdeKBF67tF
Hs2pwIZtIsRx1fWPlvhUEEhbaTZAyC9Rbgu6fjXOVWz4ORcYCuQeVhB1e2jYRxrJ
50gBbulGPOxPB+oHtKaspypSUz+qGcdeMPeTiZzBQbiP02Xl+5Rqf80VLJYfJTJt
jLJifGUF/Ne95+h1V/adWzT7aSnwcK+ijmf7YjYE+Mm5l2IQmN16WOObdM6Y4b5u
I2j5HxBupo3j73J0xNdeIUMMd4m6pTpJVvC6F4FB+JQzHUhwqdNDsAQ+TTFmDTIZ
KIX+eGLJ5N0JZsl3mWAZbwNPBXn2XvsyBfETUvJQ091ep36qxzkMASADNF1wBYxG
t9G87S3laWpuWLsmpppInrdTFoT+axL97ckPyTiwCKuoNXc5jiBjj48IYBUfpNPa
SLYToIEd44A106xVQ4qDqEhJkr4HWWHBvQEVdkZCk8KQ04ZaoWFNZZjQrUQc/wsM
uPULuULGIal6KBbuvUMHpRFKDocVsaKx0LoT7MDKqOrFW6HuhTnmTWQL5Fm131GW
+ztB25E7D6q8wqC+SLJ/oxkAcjjX5H6spg7kNDuPse90kRAHrcb2XYogOK9OIqjr
YSHE0z8oXAD+Pk9iT5IVJDmgqNtoX8kwl/iAZtUNOUdJsDmvDlGRmiVTvKrAE55A
5Mt+NIAz6VSyvntAnEtGKRBKa0BwsNp6XYTr6/ly1Kv278GpS1Sx4Sr6X5UWFvGy
myISgaWJ4UpuKPLkPU3qDY7XDq15EGB8L3Ayhor8mAa5/7CK+LaT/WKetvKLGMrP
y/UddQHaQZJcePqKUtM2tL3CzxnIS3sbo2tziK6dETxS74lKB1HZkEq1TTGqinQG
1i2+Js3lFYbX/ktv0dZcfr089OADZkZrPn1gSMYznAK9XNoRwnNjBfJbh6zVOLyV
ZEsi2Il8N3/hnE1K2SG7eXbyr/cfRPwiOoNNu3jAIgt8mAnjguUiVHz2r4uGxxJZ
lTAoGpnqG7hbUEVuyB07CnDL4pTGZAm99jkRaTAy5O0b59OjXaeDofhPDhhBO+8y
NdhwlcFWsn5VHeSTHCqtfAtgjlkALw5WMh+NtfddS/0mE4xqlOTz3QmVFz9FHfqm
KRNLEmWj4iPd73r9LyduQY9pZPv6BQ//MyhsPdxMST9mJegJPDcVp6XtJh9+29+7
n9op7WSKE/8mUajsZDT/4AZI8NONGYQ9BSARMOCh5UFB1dKRSeRriwq5FWUHDHEg
PXcakrJ40b2aCTf4LdCuKEOBkSMITckdZw3NJtV3BhMdcSDBuuZNM7yloWUAtZTs
GXW4ohEgegGmJeLQjrtZVrXF1f65p1OxkVYWno6ANJa2jFsfu1Uc4uJwO5RqlOnn
Mqh8b8stTG23exjBL3+9BU5+vKaJAvJCclpIdzwZjA2Ggg0tm+mI5Uac0ZZImW+r
amZzXPQ37304c5jhYt/mdrhrjeIjb2YawyzNTqn2vAdMJBX7DPtTOVAeNPsNhOWd
FjgOCcyTpeqVp19bmRxvy26bF/zqZOim13tayueWCVM7Re//4exXQbRwGODdtp4H
eFBnwn+oEChPz439a9xbRG2W5fQDTdS8/uSC3c3J3V3thG33/EAkx+oeCB9K1lh3
KgEXs4iIyr56b2eoZHmyK7uD/gJYpTBbC1vSiA6t94TD6BXqSpveB6m1YNKOUjzI
TKVj8mY9OZ6vpRqRa0aNBB3qeWODjefoLDaL7l9MUd4RUO5ITRu6jzj/FuxgX4AB
vAn0HcC03g25+7zXyM08DouK3IYaI93IBSkkxoz/86XQL8/l/k2f+aHlXJ8HyV+4
bL7f2zfPQZ4gfzxQlcV6MqP5/Nzk9igHx9WLzco56JwSs+NeUcShu9Qb8HL7x5Q/
6t8PLM/c2xlpgYNqu2csvg1shSmy7BiLwqR+7isDTsRaAb5vn/HzW2NcFCyDd0jD
kOz5gBlCQSPY43O+qHkccabaWFg8vu4h7vHy/xuyl2BsJLi7pSStg5w/J/S6P875
xNq9IJ1C5SHK5guKSEeHbnu8gB/MCOHRFLB7wl0+DdOMKQMNNjefh1oTY1xD33wJ
LzCaQudzx+s4Zs+a7kvOMcWlPXGagRan1B0rZEjphwMhHgbABp5fv3wmmhWMfY0x
lpMieD1tvd6Zx35pU4t1IG5NQhkwwuTXGxXSIkFMoW7VSByNQjpVxRXiRNrcs+bh
Ghalpzlk6cn/XqkuRGcDWe+lQchMZ97DLnx1hPENtbXvhW5Zn24vDeawNNhhPf/t
hnHG9rtI1P13m6R8gEzy0nmgD01E+GkGqeYfenhbhsV/5vPqQz8GqhwxHsfq6qOY
MvHdCC38nOmYeSIa6k+bPmyC43HdxcmHCjBGx93lN6UnDE9Qow1S3RJ/7zoAoZWb
arKJpSSYot5yDhp+OsQorDxqvtU8f7k6gDxDEFmUMe9RNW94WiqR6kwXNDw/dpXi
pCjZzJpCLjxuvXQhHwaWkka4LjYeHZi1tqcXm1ESrV8aPQcLNFg6S1I0xYfwPQfc
G9JKJM8zC8O2uBL4hDOGDUY/y6JrWTNEMAmuWN8E0O2YeRljWyCU1Z9/i70HJuCL
s1gyu4Wc1f8gOQfzA1YcRBCLdwVKCpu7Fz0iF8CaJtdH+o7tbJ5RPUluTDxXqIuP
MF5nWfSRcQN/tj1J3AOKRcJj6R38RGhf94XjG4nmZedrNAamqe5djhtYmNsBWL74
kPzfzCNLUH5bwVizkJrDQ0+3vQwQ8rb6XQqx0LALU4pvfHzYi/VQEbkRfj+6smIN
KCeyrFXb/qMoTryh01l9Ps4nGcDjKDAJHVXF6viVeriqxwLEUMt40XpATdiYZJzg
HWE7n+qpttl7ZZ1WGBC9G/Zp6uRTgWa2dVwTgu7gnTq49KWGarCZY1V05Mt49yNf
+CzSH4r2CqUEK7OxXx28rCzcNLaBLxu5eWAUkP6hq9ZsBgvMPw7jdjs0/bIPZksj
ZaxsTSIVniYTBClpHm0NTkUP6+LMAZNwIRxffn9/nZRoWmepZsg0d8UCD7MoYYz2
TzTxMwInuFRTtmvncqPce0uc4FXsBF9ohzY0Oy4dSqrS0W6uhg143G7/vb21YLL9
eYG2W3AC0j99LKAf6oq51P69cuECG8pZsbY0OFWSc/1mhmRkNcQl7aPGERnbhZ8B
X0mJTCD4LQkunigOLjvmoqGoilC2T0KAt0RFdm6etMhg9Gu6SUtRscZnMsyxm+It
eBx2vqrhNqVI2Zpzm4gZtjWQBRtBJ/2eoSlBtsRE1a22s5Mulfi8e/zmeWArqdkF
CxAWqWV3I0vt94T1u2j2EwWcSiAiEjamcPCPFPmQjJUl9ZUK08K6e8Uk9J+Bi5Ea
rk5W/N9fTsAVDIRg5ck81C7olek+0K1XVjl9mSp8C0vl9nJFMX76OPDqfrBgt3Ya
mABlVErGjL4lCepVbZIh3vZJrgYheIaML3LDl59MFcR+P4MmzVmL8/vjXDXTVrJZ
rMfrxAC1gRTZaYzfP5idIoxdYmVmYz32ZfCkjWG95lkFstn2juy/qlbEvd3QhiUG
8lVc7/MOFdnYzBlCqzvTr1TyaIoyJV6RsS7vTkGEHPUutGLXf+2OLkXyyl+ItfH1
WimajlDmNeBaIA80MsyLDr+aPkJdN1FkYKP6s2mdDFQVJI3hAgnoFtfrWK8w+Kng
My0Gpncwza3r6dZ1z5+kk9sEg63OOIX3/z0Zx2B7G07I6ES7SBH6WhPS1C8o75YP
L7gaB903PZfEh1OyOVBKHga8qzZc5R4oAfV9dotNkDBWJ1Cf/OfOQL/UkK7elUyN
SOPKctchF0/QanXh8u6jp4y2JRtsAO+FejKg/Tw3ePIkS1KGyES7ifh649PVncA2
u3i0bqOWjlxPbKEqpTr42DR7/fQJqkrQIO53g18YwBA2SLCZJ5eYNrGkPLFLYSxF
TTxk9meempwoW4hGdHAUbb4rZA0mShCDrz8JhzxRxeH/+lQtUYq/fFVcSuM3zpeq
glccJjyweOGVOWI52TMrryKyLUd9b7mjzV6m4bXTL2r/FF/MmlO2v/BXDDjqpvIU
IKjwV/ZJOMfZYuamE1khA6QHJZ51aIJHJX4WTfWWiLPo/xin0dzXvvR/TsVby/MY
EsvGf944IExFMC0wo0cn1sP/gQfkuCsn7MaB4X90oIjt0P8DfSKHtBSWxsEVtcJ8
y7eVAchhLkhF37msgEMS5TFOldCavvQKblMVDzc7D61ZyK/4va1hqqo0YRvmdsmq
lrIV+EmSsKZxgcI6IRjKgsjuiu4IZ4mcRt2fCo5btmC4dElg9jm7xM28UHX0HJYt
nUszBY9chjru1r673sgo4oVamrqth/Ckz6B4rp58DNHHqd6cEAPMN3T9PH5robXJ
f4gwQ8AV4ZoCqB4xZMi6Osujil/02rh2ypml0FqEisJXynlAt2Ar6dOPoFFBzr6W
i6YcOLaxm6vTKkuqcFooOCHI2DcvueS3S7whRPsUSzQ5ZAwPDNyGiUZpSQVUUo/q
/EH5dDkWO6qMhBSKjyVoGtpiIjFfee2GDBGXOfj9NNAJWmO+0lHTH1oInujDSagZ
4Hf912wisDtX3ws8gECQHYisgYVhLnIQ0GCZP5z9oF+bTxZHsBBjr34BBofan054
xO7OfuyHikNrg5NmkbB9FUi/2KL3QEJW9C+O/cL/D1UtoQQ3b7exfTbAMJ6f1N1d
fB/qgDreohytl+ozVeyIPxMfZJV2k+eSA2VOULLLi4Hrv650sAI2d59KOVMyutOD
j9SN5bavYhiT26Hz2+5OX9iDnn9HAIwu1PgKrVLQ92dcfxIblUONxTVfFXgOLadq
AyEucXld9uxawjj1pFBnsc7YI2BKw4URVRd0fzeTm5gfakynIarCCGxSyoBR/j2F
kb01NXhApnXxOfuhQKgwjHBfmGe9K9RxGX3RsaopNoFUy7T1OyrGaBcYExdt/NZd
ZOe565ilQ+N1mTeuNxE29VxLyhrE3t/M8cuYpqcLfrdXT5dwL4NumocnXXeegj5S
T46Fw6/YL5EXrL0PGzXkp79phD32P93CnssM2LesNg11FWjaELR/FZyl8dJOMitk
mHtQBrhpzadJ6paQ1F1Qc/e7NjzDTgrbfPFiStiz9ikuMfNfYj4FGynlvIWoDv34
SzDq79B6JYLbgek8LTo5ATGcRxK8QWZlghWi2T9OKD4zJRLUHmCXxuw6clcApNPh
qoQdbjnogwT7YlmPiWPY7eII2Eg3meFe1FyUhHBuENJ40BsYuW+VCALXXLEdy73p
hZFN5Co3l1C/smgulc/MyIFW6d93gYyQUvZT9FAOHRuiuKvItqpEWI5SVX//pF0/
e+kzI6c0U8slt9RmvHmwGfa6iyBdu5CLKQyASaKOSXWbk6ubHf9maAVYrFUGCGCs
Nr0MZ5+vAKorqpQ+C/K2sYzK5496FvGOwoMqEDj6WadDf6DfMwzlJzaTeu28JNff
MClVNVnhSS6sV8yXs2kyqyvDirzfu09PBgN5gsw3Zeq0o4XDSCWkp3Sv92JVUlga
TLGQwpUBmN6EEhz3jfgZGkPQuQ5aNZCKBRrMfMfsbgfslyAl5lghCZ0/mA694NZ6
flF11SGmd3tns2YwOdL4ntUu+0N3y43Z2k2inFwYwzTlnK6qw9z7mDLtK+qrOpeu
7pm+uAQaZsNOSXejQDrWevhuBGmOjSnL15GehP2Wk05+zDtiHHAuZlb9hMZNe3kA
xne0H9VxEzeAjicEanVKfM8nS9VHripwYjb2xZudY14mbot7Z3pQIAUWBEmx1/dn
vVtQGRcv9oK6aiQG7NqELdow4r43ooNOVMh7q0VclRxQFKGbr/foMfLgksSD4y9x
eDISotxEmKkZiH2U0qqX2uFSJZx8ozL0kImZNl75FXW48zwmYREvfrNeYTR0jzhh
zyUvETwtBOmzWqGgn5hP5ItGcYcNw4vHXUjgg5IyMFhDSZCde9erdPlo/oaYlVsZ
nQDrx9+XWhD8+r4hqpCsAu/aeZt4y0uenUeDgVydqLUNC9AEbHmo5Qb4piZjmL3P
RLaYrYocBzGXeo+cbpMu0atlYiQ5KS+7pcN710U2wEZdNUwJ65vRWEZBJagtDf16
6Fj3M+beA2uqmubK3v56+bkNeYyQkKSt1+Xwj7Pr8FTU7U3RKCRtF2DuL8SD8v5g
PDyJGQ/PIcyv9oZeXmreKtB06viif9z0WfGY3hGqjRLqU5Z4C2aMllZffmgnFzLj
uIYbR781Lo1/lRd7/dKCfP3TQLqCnv4xTDypmeNdvwhX75XrkyCtKmUAXX4g0rEZ
LWQHoIKXM+TDiV3VDhlzfYrv1Igr0iIKBspIYXAoGn1SOFj2E8jsk573JJVyiaW+
iF+PK2QnpF7suIj77hZ7w05nd4ElJ+zvzV8fOFPVzuCMJD/Ah3yw5FgHAKhmbzaz
PGBKbtonmWIqFamHF97QuPL8qsyJkHpYowfPJeKJIE+R7GSZ8HPF6pY8B6cqbnQl
M/sYGM1e61YoT597e5CMonavszxizRltrvDnDv/0UI0cM1YypWwnad5ctQ52jrmH
Bn0KguwpINwu8aC3z+CLnEgKHTBOnsc+UYW9rwwwc5Z3tKyHSk2J9FprXMDpx65k
F5B62RL+Qmii+CABaByUWV4msvzvUbpF9S7nHAp2Qx/QNa6ux11khBJuDHqLhz6v
kVF+nBEPEwIfc0ZqrL8eDohPEAyDitZHE9rOF53eCTVliv1lXord94ygEGV3XhcR
3MmFInpR+AJylCOHVWkKs85WTcWGCNCdVyc7jNl1+G5cwr2Cm2BvTJFvHhR7UY3t
CvtDmYGiu9t22eggWszTJTbZCKZcqQADIePbmXp2mCRPh1dgVGyXBdOX576kM0Jx
4FQo5eDFC/hPkdU1vg0o92fNbHHKTEVY/u+YjHV6p4b6eLxmjcI9eolxRhl5choB
CButxB4WJerjcUpwyDEKCwTvGzrGcTPg4o8pBMy9oqMVu/RbSv70Gl5APEJD16Ip
GknNeppIi4SJRZVBOqL8pmLWIWkUImPOUi12GkHHjxswZTQ34i2YZzoSWqgkayg8
RfHVtVRKC6HUjI54DwIc4RDAMJ/0UqyeqEpNtFoYsxgyrH/eMnsXgQWXgURxVpwt
xSYtfLReBW+RF8XDCxQyiBnAzFlYSl3umzlRnaXf4PP/NCImBbwirrH7sfcLhN42
NPqTM4ukMOeFPZYo3IKTa+ymGkZLW1hDuGYlh3ux2yaHSmU55EGKF9wqn11me6oD
iRZU9kvOxd5Y0O45q/5Q5sI/dOddhsgPIU5Bj1X0C4a7eZmV1BcbGPAq9jm7Qo+z
Db7Cpnh9uiufXSSLcCAXXPDzuPa694MYzARlTcCXyfyvHqBc+Kspe+5R3yOHLmAO
H07xAcn3gJJ5UCeo7dGRUS99/+ubsKs9gevzDgdTCfa/16Pfgyr16UyApZ8aPqng
RbSj77Lui/KPPaPpkdoax28mXJcc0fE1VD/a0aXgkdw11iulAwAbTWLVYf+NH7/m
p1IIBQet6TghjxdyK/+qCB3qZY+js4k9WHFXRIbku7WR+BLtrPBgoAVjnnpPfVSX
mx/PADrTOScs1+/yCuZY/xuhZnjWfmHKrl3GOzuWWSy9F4ltP+ErUqAWUx9hZSa5
L6zVcONCZnGh+8OyKDYzg+DktEhcMZnRvfY2HJ+7DbwTf7yztP3kqhY8+U9nim23
rURomr4ltjwr4RzXt+tV9uptokKllm99Wv8MriCw2cJISfomUcfHBMot73Jl6hjs
vlGhvK/bgUB7kmCEmZ7Ui4/xD2oQyhKOHFeTSqktD5ey3fPiWbMswYcoloAtFT+Y
FhgaB4FXxnIKB918foLGj55fAkQmrieiglcDyxCjl2qqxQqdKJ0TSD8ttEHz9jIB
3b9jy9UaLZ9QdAi5HIPj2tnm+UNMzl4OBueWykjLJLDteDQF8MisSv2iuMQIPG9m
oQ6qR0lFWIe3ylfcAseESnhrjDkmUCTv0Wpt5MCj04RqOS+mwahYHBLBuYwBDuag
3QE3aJ4Zitj2zE2MpqqntbnXiqYhMBmHm4EvHAy2Qp3LlWeOakXxs2UvMWE73yry
kLPfA5qJnoTZwG/t78g3ERI25b4/hjNJJ3XPqTGtn9ORSjJ/KsliS96B9hi7fFdy
LBArjTgGhZYvzdyGLsO5c5Z/1fEXkGKgkhuEi8dgsnOc5CNygmj6b6gFbG02lyd0
iQG6/MV/NTjibGrD8B35RDbgYDdEw7/yNQuVoNwl0vzJs3wKQ+1OxypQIMh5avKw
mK9FXrWzwpOORZydqKgFjL5pVtbx43Pd+sq96q+eR19mO+ncSt0brcnwC3m2eC5u
wEDrOfkeZjLHKjn/1CjBoGeaHFmJm3n3Jc/4V9xOl3GbRJpU5R1HGxficj7F2dBf
D1R1xgXvor0Ap7BT4YkQ+ZsuvfkfQaO/PaVcYnGf48WnYnIV5wvzW93U3J7dq+Zk
zKydWvt/64/P1Swe8kfNz5dbmgovzcRO8ArIDFsk383pUhV5xoo+AFNuuP5AU9ZN
375OxO7CkHmG06N1OSDx5TblVJj7Ks7TeOa9WbWiByoNP2gEPcmNEmMv8aiMVfvA
LutWFvPzJJSkn/Dl83AxCPqfOORM0hsE0GyEkB2N9yW+I7e22rmPr4OoA1005a6l
GL7sbcPrmnT+cIcqUio6ch7EUyO4oamB480eHaV2MZykLmuTMtaVu6w+sZEKXZ+p
s0/bWSA4EbsM81eSABNGYvsbKX8AYQpYptb0S1ts0VDw23CrVwNXnAvSD9dDoWvp
6+PsHUgzaiIhzNXJuDgpMr2H22VDQk/u971YJwF+iWQ9wJvdDDfZ8gND7qfk7PJ6
uFvjeQk6i8kRypLOMQb9xVBGlUFcPj/fTkTdJw4Y3j8nUq50YRWbqmPwH6KSBeKH
dHUteosD6YU7dkS/AS+vwaDmlcUgfCghHcxr3LWMlJXwgr9Ax7vEcI/J0w6HdTfn
w9MfZGgtxzZ6YovwUrw4O/3RWbELBWg2wfZX5X4GCkuGahbszc76WMxjfvKPyiTR
7yE7k61fwhLn8UaPEiGnli8nBttUF5OXNo99DmqTN8oOkKAz2it2FDqAOlspA0dM
sOjVuJBlZ+TIBNNtZ/eXX72fEPJELivAJwJRgKyWfKVO1bJxmKQ40Vd5GQL9/GMB
q/9hAmvckC8Uu3KOjyVSafTRrw07JQKALrAx5TAKvSolw72OyIXEpV+Got0/09AK
oau7nnQzHevLlAK5jAOrTBGOG0YediKtbN9k0TSMKTH6ehHppEa4huw9ETYtsWv2
Gn6ub+bo5NgbSZX2RsG033QDuMrKlD/HnoZYUjvWvlKRDNwVThu8dFLuTWkl39Hn
E8dMKfRqOXKq+T33jSeZoq9TAH+cvxL/nYDCaVN4cWFM7NDk5b2Fs6MBF44SdyAn
CxV4kSsJPSWCh298NMowMixYYajdwSzgi3CNYVtIGyuaz/CWnjHSezUkZI+xY0LA
vrxMdQwxQBtE9DSfLhpRKw3G8Kehwj93q9Mf5QTBLG3moJwopibRufbpwXJ74Aa1
LQEq0H/CQamFvgtp+wlT7rIg9J9bMc0APn45CZC0s+Wm7Mzfr4NMzHo43D4tob5W
cwa6Bxekzico5tKcLmCHMecUY6UORywRHi9hFMV0MBYWxULOE60TvSAIyRfHBjVG
mdA1r92YxGnU8lMEIYUilFkKXCKNy+Pw3KDkqZQPUB/K6JdEhsoxD8+q15HFcdFQ
H5vTsNnOZhh32/TFR25PfJtYEbPv33/P8C1jBezTQeS3mHC7r/2duSUH+B9+oxb+
QpAsGpzgHgB00oP5yaCo+Njhkxu7macGcESvZtjfQ3L5t3xh6SMFxR/7wDwP8S2Z
FooDEmPE09069XYhBTH+QuDtk9gXVf/OI0duHMssjx6LkzwzM+A1/Wf6w36gCmy2
Fdwzlw+zZorFfCs01QNEXMRF7RxAuj3y/oPrw4E9uijiJtNX5Vz2khRTLGS/FWmU
yX+eFPTQkRlSdBehlHNHG/rYMXrc75JSJKr9bpEK6iw8pXsRqAhd/PsszrLh2R7O
23ZZFkM1fQ4nK3r+WN4t0m4jN/9wbUWjM5VSfFMunh4KWz4kN4VgTPGl0luMvv1e
hfAYUyT/ninOxF1eLzX+pnCXUTqKfeiOYcNTr2/XJkGvTwXtpsfWAuxNa1Y5D2ts
BcZrFOC6TxtOdQiC/gaaLlG9Xzy0MOdNAmSAbsLeuGw8wKTjOk9r2SdcbCyP5zJq
ENHB3i/34lucQ1nrFksdL+g9sdKo189GuVe3Mjesb2wErvF6CTTVC4NvY1sWwhTu
M0RahzngWrrNbsVO1g3UVZpy1rjJFOTy+7zebXUg4MjjGL0+QkDh3vcNWz93/bNp
dv2YrhzcMjowsmhmJzBcylF6S5uf4fEZ1YhQDfpyRiaUaeA7hgYpGzTp4buAvlVF
BMVyIaP0X7cmaN5t0iuD0LEX+LnpBtRc0vhmrJ+j4kIbSGSAf1wtrxFhqaOIQbTP
jdhQEwlQVQqw6kKiBf81RbkCkT8zmNBdh5Lq8qRxioFr1nFkUNS7ZLkZIOZIL3Wj
aRL+wk2sKkmLklAcu6954/+Wi9GfBIbs9LuTNzcY2n9f8D9d9iVcLr8DWYrce4tU
Ds9S/4Mto1IYKTzWHCdURonEGAZ91wkIO0xqPoMI+kUSkTYy7YdcN5DSDxlF5Ph6
Va10qhf6BK5JqXiYEgaF1oTc780kCXb5NUcbs/YyRxz1Wly0YFMRjsHXNWnfvm/t
RmOVHRyA2jm274dhd8VFp4uQaXeik5xn2/coIt1T6OwlMIbbxP4wubH0frN8zFNz
nhSWDfKHPMUU1o/Kvex7jGMMGTPxuoY8sXG78nfSi0BcvLniWD3OenfoVI9wqfrY
4HvQgLCInQydyU4j0qDsyjJpNBSSKxzhcevU0XiJKTZ/B6eSnigLTY9ZefW64Tte
CBCeDIx7foLq3C9UWRrJp5zKX9rZBEexVcOiQlrQKzupxgVkt6oXIIkzbyJnIOOM
hE6IlZ8lUMQJRuLuxrSdKtvOxGF9GJaVqLVOBKLWs9cQniW5zPswQKyIxdhU6tR7
O0DST9O9tc4fJJy1AdSMN+oznIT5oU46SdIITZEOSch0Wp8X0LWCZ5nDyk6btA7W
RPLKIQJKMeB13wHSQtjGZGfpHRoGK6yvXy0vFMtSiC7hvBlYNeJTnjfjdCiyXNRC
+myJ5meiSmxx2mLttVHp3ChQ+n1Z288gtiQBQE0qzG6b5NrP+LWjYGQlrBQP/bqo
2owdAQOxfJerzLtnx/OsgDnV/qzbXF0UWfCwGlY0qb2EXA1tn1rssekb2xOMK8Wb
yZHTulFvMtvVvsHEO52tAkxYRZQixJmZoAO4LEqdm0fNleN6Kvgb9Z3c0xR+WxGl
iMIT6ZuVWYHwiOA38rUPzLwuni6mjRj4I/UfBvtJREee1vrxLQGLGfhVbVVdk72i
1g70NBig7WLo+NtyBdy03o0U3FKPidaMr68+ENdpHq21nK0cv+JUzEuW65qBYoPP
p1QYzeCjp2xIkCKbC1+yABO2r4ke8b6d07Gh4/uoGVtwcOvzG5LRluL9nwHQLh9H
UrqhIp7OyuRhKdX35xYA86I3kxybMkYsCOk0GMEjS2bmx6xal6nZ2e3k2xpTSn+F
z0s1Dwxh3lNT8zJ/UKHvkhWLYrDVLK6rLi5hLdBO8QU0L/r/v7l9J46KlB5HuYm4
t3uq4TNlWasy1lFTSC8G9dIMKqXnTrzyBGXzyL+wvgisV5p7dawGNy6XyktQav51
Z6ka55IUoN91gl5pGxv++A1Ewh+FHqhlZp4cliDeo7XUchkRn7SE0Rc6EMVWc63Y
1uSjzl4ysQTTAZ+Wbo5j+Q42zzhvfBOsZAcSzEQYeQ7TR1UkGL0LSVHjvevc+U2Z
awS/EZjJYQCUw3jHmcN4SOb8/Y7Qsf3kONVSr4eNBN9sQ8VZn9cGhLSFumEQtjhc
PKlAlW81sg1D+tc2M1kt8G1AfBL9qRnGNXlViRHi1rUmnD/qIaiD63Ub/mmZLB40
FWAm8huUVlrhdVfq5DAK/sPpSaAb8BPXjfuxSCSe1fgELl++S8ULy9K/0fEQZuz7
tMfJL/AdPM39YJkQE/WNWV65BfWB94FmRTUiKXfyJlzZMjFCPOfLspdKRxo3E97s
zlWrFe03Zh7cRZQXjqxK6J08wy4XTmYa0xrR7QohBTesJmLqBkRgGvug18sHwBtt
zXxzt3ZUVZvr4eBtDKTTXojxDX2pvxb8pOJ66S5RNLtEbMG9mDt1HZqBtYCKRlR/
05YGd4noE2w1JghSgS6DVSewKfmLCuPFJ89/yvt6XnGJQ3j5doVmhwXJA4eSwsd+
oITAHH64NPF7yq3soAK4GhQ0jjbLjGLFLVkg4rQXsx0h+/n24M8WnZ+yRi5r9DQj
xhaXDrZ7jubn5m7u/Uhnqucq20l/5j71wwv8pew6q5jIbhGijCKOgoD7HNHX8VDk
Lqrgi3Bp1OevuAFujY86OFOdxczxwkrM2yINqk9Laif+geMms+TfG9Km5fnKWWHZ
e4TcmeQ4iDoIwDF6MBaGh0PChyID8uoWUBPUOnQAt2T/2zIjRSz2+BW1ss0aCBhm
KdibpxWoajmZZX8bStUHWGSXHuDhMz7gb4jI8nBSgy6sDAypJ0JCf1NH4A0XKdGh
U1BU8HUDTtdVYTFduMAK5Zh6QnanqNpnvm00caC0/MFuuYlS+A6Ekt7UU+mflF/r
qU5JDE5QBRsg80fE5x8XLRI6RbUGkDxWnELyTAUYQOLOS8diTVpx7HBlo6kI6rOW
tMr3e5yTn/1O6mA5Lm2RPh90iYC3cC1LJTFHbcLXlRWvCo/ypoDO7ivBywRTleay
yFiN+I0c8MfukTp7OQfxtTVy19QXCBnI5vzK5Qzs2v7MrjpNq+klAMtt7J0f9u67
UcygGwvzTxHRBbJ+7lzaTO5nHJdmHuRsPrNPwGHFcNVf6p85rDJ4GrAM2l1ViSic
T7c7uhNUcKWfX3octGYP5dizyzqRMYvFHM7Nm58zU/EHRf/T3gIRoImdKaUgZgq4
P9MEWQmNa6i1bZ+wjfy9PiK/tj2CKVf/HodPTJfBWrxDDb6d2W7PEJQPK4XVbC9A
uENKFzjnIq+r+xjM6/XZYyLSS+yCgLVV4WOOvXUWyrrFy6pOJcY+9lEIpziBZBNs
1UzvV/2qkgzR7+d5Sxgtw8ov4I4kgeHwEXAGUebK7sGkyuehyeNaXq2dYcFk0yFW
H2GZVf8mC1Dni9eNQHnAgT9X/lowuvM08XtNMapSyJdgJnO9go6hnNHxj7Bx9SPG
qEAdV5lILKfuOtRS+8shdlvO9oC6Yfu4GKbK7uRlfib67QTL6QFrAFEgHU5GWiMT
UnW7G2uuxrP5PTEi+qumIUsI4+fUF6fpnEYmXgbWZ0DMN6QQWNp69QzBtd7lMJLI
ccHyJejtiHYdUiWBCAqn43OTbxmCaPqOP+DK0n8I+6AksA7sZ0mOUU2P5Tn3VlIj
pl1DetUvjkwtkfGZzqgvSDuWyKCjtdAdOSWjcIGtctp8qzjIRO5phpQ828s9c6dK
5/bIS4hDA2pafPMZfJ+7XIYHdGVHc6PNYojByi8Zyv2T0cN4S0LPzUQx3hk13gRQ
B1Zit5bqT8VuRECzYO2QTj5PJ/tbrwWUtWxzLiTeaz5pwD36nO01MZeuMkWAk/+n
4+Jpxa4g8a+IJNHAiVXxEQUhwyXU7w/yjRLQmtcuFXTlK2fekLei2b3I1OL7OtKl
l3tRzvMRU9uWEM4T83TwvvRPep1w3RvhgkzF7CJQ1YRUBEwNBzBWta+fUjXeODRm
G8d32ESUMLwG4sVLH4bH9ujdHg42qce6aOBnkXeMpy6oELc9vakleVL1PeEH3pH5
WV1wKGLMOe5zLSXqanzRLQ3NuLjuJVM0AP+u8l++/MAzEcIj9DgMMnSzK7f6TS5y
3wBYOx3vyCqGgyvk59lcbh+qedn6dpaWs9N1FXBugTDOoc44AnDDWDjH5fTgvRW1
favnhJ74tJYAtG/baJHCJoOrElwL6nJmn9nvQBS9vYglt5OX3X6cLAdxID3+QAxK
RRhhDi0LGg3OM0XhO7YAlHpFwIfeAm+RiqGI/RW07oJocqUg4fRECtI769nG3j4f
sKSMQCO7LjqJjfbHBhmJasJMmFCMyO8wtXPATqrO1mdit/xJuBtyK5g2zXQxUqYx
Zn6lk86dt2vNYt7EEouZJ5iRp2peh2HukHmPn3asxQr+jHybNAMAr+s49IUVDigJ
U+6Xbdp2JdPmS1r54pcVCCXWskT7L405pUwT7+eo7/B8Jwcf1KN6PaQCMshD1pWt
H/frV1PkT9ewK6LSOlmc3KMl/1xDg+XiX7leUT3ozhatzytWK3m0AEdjIMaChSPk
WO71pQJevl/z6oo6lpDjxBbcjEsTlQG6rVGk6kW22PVu3URE06jaeyYRLwvKpcis
oLj2Z9B/VKh1cLfA2mY/ttgWb2aup8Ogu8093jJkAmNrFPJiz96PiVkDs3wPv8dZ
Q9R7ZaiTHCnKcDpvguqnmvo4tLipWBQSJTbM/vylMBbeuM36wBbI2hjaHcKarcZ+
iWlPVN6JCRqVgF9wD6dZEAPw8MbgSYtCPbxUZoWlLnQJ+UthQ/BLqjC/FvgzMpNg
HbBK7ViPB4pdreBJCzN7Z6QbE+4eHGz1xNTCN4N2UH/MRzMTlpYAYlTWYC88OF2a
YOJw60MqDoA9GhdUMY16eeRZJ6OJmoD1l+/mPhGZIN4azv/RSXV5THhjW5Dr299H
U4wB5Tku/Zkp/sxoAEy9d9v8Cy8CJnrw0indRZ0Fq/lCvWK8wzQnHViP1Fz50vfo
MDyZPc5wHwF5kSzV9tRfm/RlWN6mMsjc5MOXQaIGfFdKkMbfbU+2mo/Tmtl/LV7Z
WP+G6kqcMDWk8yEQ9Y66secqUOf9h6PsZ/0ZvZev5eEFA9SVOqUuPwujR5w0KRPv
1z4gedp6S3xUFciMmlbzhSzs1/WvFjAQLo3YtLC/oFVQ+sk1ubB3sxRtSiqA3mvg
Z37ONRRmVS06L/L+QNh2HgUde6nbWWR16ar23yMIPGqgwXpQyu3v18jhSmywmtJu
wMZAanEBK67gaIltAvXXKBFa1Dnd5OnKc//zbmhhn3OpaS54V5JcnV/Y1/cUEOiG
x1tGVnhr8+Sj3dLdG/20f2HBwdGW/EJuIZxGDMJ2+1V043G+Heqnbk9U0blQa24v
yIT85U9jSfC8NS9hdkebD50wz1yQe063Zn+icN6WCPiIsO9by7fc+cMz9eQOHWDC
+m5wo+s9d07RFqMKU/936s6l1OAC7HeccKgLGIhZHz3FoGgPJ4i2RPnyGPQ4r746
Z63FKNLBZpBTJXBiKwJs7zDuIelfEq0Jm8wveDHUySx9SiY9gjxgkSxqpjltn0re
urw8P2adW5JtfqCs7Ad1QCiY7eu56kr1teZoHipKez6HEunCrjDrViJHH6j7/B8M
Q82ttLBi3ill2kkQ8ks0s5N0HPzxskrviM/5dzWVzlOCMFksgxZuCRB9zY01kN2a
3BGGzapUwEq7n7YoLYr4iNrSxI4lOWqHf5OGwLxOOrc9MdvU888q6oqscsOcpWSY
wyHpDVRyVrIjm2ffmlWlT0f1ZtQH/3eWrYv/03icnyYlTdNUWkqzpuuLdCTeuC5P
mLUSIl9HlnPf4fuUNutJCDic5JcrUqafxYXyXi7iF0XQAbDKgOCcTTbK3FoJTmMy
NXmQrD0vSXgCpIgsljOj+WUE4s8/0Lw4xSeYPDgbDyFkQ57PfOG9oXfc+1MKnxuk
5IkBpZ0rtLq0nwmyqrEegMqLFcMZ+O05MnkgD6MGa9FkU292j0dTX+vI75j+fgRu
nLt9eXCifWgA4yKL73wBTNXKlnYQalYtylG2J+cuNqF5fJvwzDPBR7vyupoq9Sz1
JURcpFXGNCoWs0W9bNvn7urmzYGBs/qiXVvvLNot3ybhVDar3t8E8q5HkY/RL0X6
JXTC5tNCZJExFV6N7V2cewV5FcjkfDXb5ic/+0lQc1TSYKERtZoRRYdnI1ooY4Hc
Al5nPxFOf8VhiL6ZfHHSfVKlIuEJr5TJggqGsiY+XeUgXXEPQO0uIGc+SxXr+jid
n6MjslzznFLR9WUYxG3MKXvSVDWB5xob1q9+i9CGZVbOFhAPiSsWbLvoFLULT7x3
qric7EEY6vgde9gZeBMl2fYBrM3Nof7Hb3ZMm2xUddVIZ3TEFZobTkVJcxePbme3
WWIw0PKrW336kfCSUHZKWxylqPo/dwq3EwUO/EeW/8LwwWWwTRzUc2uR1iX+rMzz
2eByuETVu2j0GpgtElrMeDaOVZyMe8A7Gyi0cmH0ILf4LXGN4BMq5ZFrJnMCDlE3
p5lrRAbLy8zexENRUN0f4bsfLE8o8IeQb2Ind5gqUUSFwj0BScAtF7pfLWArArBW
Vp+k1cC5SUWCmDQNEA3qalN9KIuMaDwaIzXZldtlri5qA+DNjkl8cJhNw61HB9RM
fYmI7Oaj2DZ7fldrgOUCei0YzremEPrDImw8oM/Dp/31dDX1Gwi77WC9tQzt+WOu
IrgjZgRMrYXO27bfuxGTAgGXoKXJglRChpgNj2/XTpC3OND4EFlGnnIDW4t298Dd
tQpRjRcOomN+iHuHBcV6FNAb25Z2t+PN9ifSA4J7wcQlcxFo9fBEOKcoi6KwSLSQ
PYgYjhXhK0LV4W1Isr4Wnq+x86LeoOrZBIQ7dsSUF9ARAxsdk9l9qqRyh6rcyqLy
1Cvipb/sDGn0VvZ7FMJISJrGj6s0r4wRxJPya1AnnEiTUtyf4kjuhKBVkk82GAQN
FXIGYOQ041Ap7sNFZFAofcOL26t2V1oGIIBs/+X/Pvu/YhP6cKdZE3yagYXGNGiT
LCCbCgBe8cJnQ3y1Vl7DMo9sF/XsKDVo0WRHwuM8J//3cFNsx/ju5eiBHsmyRqnl
qoUa0zahxFPZSlG2KRc5JgB4ejJvF51EqH5u1PN5E2LlDQAD0dN05vyT0d7dOCTx
LWfWRoik9pchqhnDjyjYslxCTJQ2qku3fhhV7sLqGYwuvAgLTzZB5hDoVSg2pR9Q
Du26FceQCF1IS7W85JtO2EGP8yLRZ9hPPI8Ae1/uk5M+o9jjLU3WhPX1ss0kTMph
H77hkjeVBJNvDmtjYkSjsm5T69LTIt7YLU4K96okIBmsENuqpDGtuWnKPaH2RPGH
7LhwtuRdxibxiyQkEZpZ3ZrnsgbF4/yMAR5MidG3e1aCsakLAbRbwmt5HotP3/xE
RaoMBQMkficAQNSCULGfli4Mw9z3fg1K4oMKGW7Z9hajlp4TOP+Opl6Etlrx3qQB
/LxF93ZCNRekY3TF6EnHxNt4smyUyud7DXlUfW+7NAOlN+p4NA+GYuVx3BNX8vwV
aO8ro6aK5t6TU14BcFlF6QIZNYeVcK3R93u7iixbkpTCMzZmZgr1sdNf5RmRfL89
oi8DlXZUFLdKBVxo0Xl8dwcDNBhr7YETdE3g1rSNKDfaICDim0RJFgmLvGD3iDKy
iM2k+545lcDvNDnxq7+6bojkfFUwuDerrfsQIr3ftpaSkmlae/66WEB+T5xC0J46
X2KfXhEenl7kyL/Ey7da6SG37IfVIXEZBDUmRce/rupJtz1uK20lzMm6RrRz0KM1
1BSr90OvVFzLX5MyNpsVHTuH59VrVvtYPJqC6f6nBqO3VhJRImNvgyB5PFBDHJPR
MflD/bpOOGSJ1fc6aT5OJ9rDJUABJ7JowCJar+a8UDyrcFamoUZkQuoDHY1JrgNq
JHKhahksjXbdcIZwZI+pGfOtMVFKeqEdklm5xnjmi0INb6vYlk1hXeW7bByAdINk
XzeT1z5pIXmY0anqyMVI1aDAQks6o8ZnnPP7MSn497QO4CrsuEv2XWKQiAzctX6A
mL2PC4jTF5dp2K0O+DOxDJ1Gqa6OdpcdvyLaQP0n3yaB3M4iIjVAySbcNe+JDNoy
JtbXuXzoCGzzjlfshh8lbF+N2u6Z0cS0NcO98yBuR/Wa9mW7Ipx5BsIe/JyeTLvG
3FNZJ6P6JIAXYrXG5K998RkyQXFm/j4+GC9H5ngMhROs6/9qqh847egaSNMM2a38
SajeM2W79XEqP1ShVp9Exkw0t6Cw3TAh65zbh71TYULP30WfqwoCIEY2rRm6mwPl
+Hmcz4inpeAeSaMceuUz/GJCpgKhzXX6v/CswPLXxShldaccpT4o3NR0/oiks1mN
TPS7bOzJq2rZp40whuU/VFF+aFam6YB8fvRa3QjwjYMGVfaXM01WuKvBUN91oWAn
40xlvcuthB7+vCq+UEowRzHkqv7PBavlz8n7Z8nal7aMsJ3gYdfc1AjKoyxBEhNT
3fkAect33uOfaqNNXLlNQFmoAdPYdJ4MEs2WaanXJhR/BO/N0ZZMMZit8r4N5JDN
BAxURQ87nVMgrOqq9KXX4ulh4DVFIpG+iOf+SgJW5PmjkZgjNm6UmmvAaNH4vt7D
LoutogTFa8cBa5/x+SwVdS6I+aC5jBeq9t3sLDSQaBBVvUWXsU/gLhGcwRvQMQgs
Ydfh+3KAFj6vK+H/te29t6LHeNO1HhdDO0qSYU/a/XLh7vBaiTUHbdKv6d5d3l/4
oISLzEIveti99jzHyUrCE3vlFhej2aApKvfmJB8TKWAAhA4tigB48UKAfkoUDxRT
WP+LK5RGUKZZDjg+okoKsh+XZQnG6AiodE263dogh2f6bvAyYGcThcUFXZ+MqP+Z
8LUVYYoPVjvJwSct9tqxS+US5yWKOToI5/+UBgswokX9XUKa9xd79khtn8lej7Zp
fb86vPeN+9f2bv5qFXFd8xbL+hGdQ+CeEOvtHQHmNlJdYIklQvGBFEO+pWRhrFvh
xxWUuZ9KjdP+/MbXAQhCM5ckAW1/YCAb1JgrBHdurMU9JppHR2JoXR1symjPwtdq
Dxch5FyWtgVb6x2QIsQM2RPMz2kEqvixARh60cPNTvDb0VoDGuMJVmU8YlYnP2kO
3D6VIfjfMq/KrtEGd4m8Mbj4jpxsEK23Glv5SI+Vnd/UGqUAOH3VyIvpBj4D61j1
3XLpFN33uORhnqGaMoOKI6/Yi6LbaGB9xMbHGTqATQsJgL+O0hNwF9IowiXZ+YCY
WmKsPZoQ9zUpbOtFuRBI6tVmOjnyR33WGHis4gcli+YE2vY2aofsPTvR8xwF6VET
9rSScPlyDXlap/vkUa2a+07g2QmqTR/oFTRzWcecLGXDX/TEep+P0FeDxTm6MjB1
m8E2HBpxcKHdiWMjw7a9IyIeiwArQ2iWoA0/TIuUAP3YqUipWHZCIXfhrcPZESua
9QnAad6F9Ug+CIpzYi4t4B167S1Wy4tcGM/bddQOdZxzzTujzg/pguoIu3jLO9JM
OKo2yqTzq4EcJZdYPvFWsGNct+btETUDdFPLb/Iy+0+j+jLaBOoEzZdyqLl1K5vY
Pis71O5s6zw/fjx3HpnGw6bWRhMKr1Wuqd8k5aVFvlKgl4z9wAHDR3zBOpbLhNCo
NleO1xUFj30VRKl/ZiriZT58LyAeeaLH0KQBd7gLBKI9KY3QuYN9X2v13JEQIm+I
FfEH9GpyE+odm0TEnJ0AMlTlOXIoofvAQrkmSbL+JddYi2zdlnNEE2iV2rgfebCG
L2qBDq9oNdqdygTW8nWL+hzLHc3BC1nLLCaXwH73YS0ByqB1adxCDNvMUtvgU/I4
fPMVTqgGj797yQPhFEwE66iWjBD2oKO8z8iPT4t6YrDH/EzLhVpz5wfxoVtrBItt
V6Mo5XM8gw/dF3S/Eiwra1JZ9eWjSrHxY9xvP0UStdvJ46nxS4oZZIkmveu1eAtn
MoM8RFp0jOEMLCL2PChdjZB4SE61HYdZALOJzi6foRypshpswCuGrEPj6sRhxjwW
UmVSikUybmf42q9LbUjzprbgwjCy0zrIDJPUmAjnFKZqWXg9IkZTSVNli3XjdO32
2ZdDWiOOirtV/DciYQMy8WxondeM2ujqE4EEWjN1bGJq58lKqBl18C5xaHzSBa14
cBvffFdWww4ygdqeOO+xEU4QLvK8Sv3q2+k3J6opwfjfX37BPJWhZs/LVDzviskg
wEqEOiDQAJk22YTQMxPMKh5uCum+3SNBswubeyT/Xy8ME/kk6e0NKSciz2xj4MPv
5mbx2PGlJmslSE/P6mnrI2EsyIADj0i0XNHVb4PJKIbHcMVOCLXqFqRnSrwnbRMC
wHmt8VFpyxlv/P7Cxe1U8aWw0lifsx5fIXhf8ydapGAwSf9YLd2G5osgktuI74dv
EygWYQDdinrUouV5pMWk2qxkepc5fVT26euZr5gMiSlcbrr0C2lj9oygGGXD6SkB
r2LLKrze92OuIOA3UlI45lLu7MDAZZknv7rKz29GZE/R1+g3O6aKmvHWVxIYPXk1
O3zrh1UPG3SneWoItnoXzdgx1D83V1QrvIe243X+VzvyTLsvgsi2yDW9Ot7+u1ae
OJfz6IcuwyzGK/Zr6wmlFrDgGiIebqGdKYHah/QRjf0B1TLoW1+yYosBzC3xYjks
oIv7NanPrT2HxvRzhVKeyT4lOnnGcoBHxCR/KrqnK9Odn7GyLZozJmR9TG/skJ4X
lc15BfC8801QrvtuEUdUBwRl/eL1TzLui/e2/IbvY/e3oXsbROJz1xoF0rfyruCB
TwkrsNBSpQWeX9+BIqXcq2EM1rTbYAPRFh7+kemscjHQE5SrTBCYXHskVYny+HeI
jR6oATxvfalELIqg48qY/PP6SWxTMV6N0rVxBlVwpCl+7EAdnPxhorsEeA+NO9kX
jHX0jfzM8Mrk+LQd/bwTqcFszPjox6yoQnXLUsjaeS2VLe8E1Khh/hwMiRnZwtja
YkQxqKLdLDvQOT+2s0rIxjAvaGuW5z7A/sfVfIWMXtcN6Fc9QQNTHK9rY4QCmP9T
WQFhQj0FgcQUe9dWRG8w4hcaP8aP96ov+ehj16xbFZR6J5AljSfpG9eY4xOuPa4Z
5hJNt5V7uckvpA/imrvvZ6AM9ZuVxPMPTJSPHE9e6ivok3s+63co+7lC7UiGQuwZ
9ZVBFxp93D2Euk8ll6VP1IijsHxP/o0edUF7O4VONODvC3SbFHjhd/zl8Cgn3Cli
qrxKwwj3lzVdDhANlJ64U22P36ZiMy8NGKZvUEiPwda75uM2zs8yI/1wgzsYbJmB
lFyuaJH3fKc3xiMMJQq5yLlxjKxB2H1Gqwfssv0771VENeHzxlso/gGBMAr3H7Bq
ndx59MBjaxixFwtmog0vs2HTgH3gdwJXgQlYK9i5jX0JcItw3U6z2ga0a1b3PQD4
LkH49y71umEftxBMD6eOgiFTye3p4vlgonGcxpyPHAq/JOtyX5Bm9NDhBs2yz12T
3CU7orQuqNahFjKRstrD9sUgRG65skCj6UxgWnjihq7+YOGd+BfQEHPED3vj74HX
+9bwIUdQmpqfOmeixbWSCX+BYhuTIstVUoESh2UzdFgDT8ayO6k0mH0KGddz71dt
6ZZapnvcCkqs6NB3Uxrbwh2lI6Zt1grAKD13Neyv+WccRvvnqIdVgDhcPt5XGuWv
cXIuwHtBrkCg+jUCKDfoSJvEu2a6UG0o3DT2VXf/lcv5rwS0JZcKawI3UKZq7/IG
StrwAAaEEGo1P/xmvR+B6IIHTne3bmmtnmIgKrMh2PJSt/KQ1Zyr60fIqUhWhl7o
/BhoquL3vBpG+L/A2x9wwSlYjxYUcyuciUDU91ASSVv7twwu5em4dscVEu/pZ9ON
XnGd33Z292pjC1UlAealiP3FUS3zz5c4QlvJZAv9hKgc1V/ClZlHiruH+VegP1nS
rq2AGaPDCiU+fR2M8kaQTF3s4giH8/CVLvC/906e2qxHYcatHmFuBdOXxXLyRCfV
x0KEmvyY0kby0XdAwHQ5mjR701DfV59yhqwhXle1PpMYiOBldfBJJFHZsGiJ+rri
cHFrq2uNQxrMsIhZLlxcEKfBZgp5JP/QS7gOZvIEs0ax2+BUm56st4/AbPw+WgXz
XUwn03XrEC+ymoP+e7QfmCKh9PtNAGyt7R/ronYa+mEHFjq9o9cr81Qgww5qTajr
Et1NKdUCXTD0TS3Y+OLYklDLJjigoLdlFv5hjuEto/CesvA2CV2wFw2RygApxhSl
N8U9+l0XqEC9QM9A4FE3dvmZ9ny93ji4d/vfsYNzCONo5PRU0Em4e9egi1NbpRLG
rQzotCRi2j8EFEjLr/3iz1pEYV8GF19oSCNtdovxK4SqEsYObOetrr4Jlch722WC
3r1dGg+WyfvH8BngQC1/gpkXkZzT9n4HSpEneT2OjtrQcT92eKkjUQKRARlUUAzo
XRTkh14O8l2on33LvXI4gSHze4RfdLKnRsGFk8NeGj1xvXNjANj750vtWNYE16/V
XspdDRUnTLaPV8CJwhePl0bucWx9C1FN+RwQXcM3vMNzNs9jiVRGNDGWkIrL4j4N
pqSrhYhlQ81v+SQVjt0ik0/OzZn3cDU5YZvye3opSO12hFeV/3blrGKW3ENBX1uw
LglZVwr3LXiAbQQhGt0fQ3W9EVKTbJMzxC1yVV8zf9VS8TdJuV4xALJ7MEFjwGgQ
zhuNfXLWJDZr5p7C2QoLlGID+1G+xzGA6jewyiIBhYMkjw0pW65yiHycKK4tro+D
4oLUuW0tM/V3qvX2zrXNYIG+WiqHvQ1tP711vipNVUCWkgpKGmT8bbWKpjwx/1Ks
1fam9npcxkPCtc5Gi7amVB/Ii5t0GlAQxAKlUUyzBjsljI51n1d0dDQLiNbQoqNi
8yhRc6RdmZE91bcHJde0rwQ7vrnT0ixbC25DH4sttoAmGZ5I3MJqLWF2fOOlI+lU
2P/vvZi0BFJcNscKo0hHfgI3ymOGAUY1aX09c5qaHp/yFoVjCOcbDjoFPeM5jV5e
uASztYss1Umb5NePKO74gu0ruwaN3PtL6Si6G4Rir4nyvyBUY5+KjuMkzCjDPnMe
F53DMXk6QFW9ZSMGw24KOO4aq3FaVoHengjy4J+VK7GTJD6eaE/YlwzUkm5Drlcl
C2z1uDQxmn7AUrwAezzjcJLC7X5cahnrfHgcBuW5EEOtGW634QoIvhNdDcfjCVHl
XpfnTRxk1oV/NW43v/7Nt8/VUnplGucELUQPVzCz7r+KWbVFUD6Mve0iqX7pdXNm
V/pV4WC9fXcIYyike3end32aEXwfTRn9LVWe5QdH6Iumfr7GM4BpXgehN8fHREz8
zQKwwmNvh5A2e6vSzws+sk0t/nAagCBfZoORR684plFwAZAZa2bguKeJH3VBbbgG
o1/GDRuyc5G5RHaXmOd/7eQ/iGHUVNS7W4+F32N5GGX/Jg0T9Ywnc5mTNIAOgtrN
BsJi9rtFMdhUk3qyuOIhSyeFchZG6JuJpM0Dw0vaQ1P6qrCWclWjOc7MsHJ9MDFh
EXmNFC3nEbps8zqK4XRN7Yu4GRZUdrNroexR76EQ2qhZRc6DQnexYd8dArKNoBdG
wtHvZiSjT7k4z1QusIr6y1nzPQkztljcQnUS0MM/E7/vcGz/PmW0Aj/4HleQBFCu
TuCR7CcpeVlOCh0sDjzYmD1KU0wJ62C82PR84kUZyssX2/E2+6W5iIXuOMMOfIDV
pwXGt+JfL54KyjCd47Xx82h8YSQM3sE7ecuyd+GLqyAvEbkU+adxL+XY/xugMCuc
P9HC2BpOvn/j9xPXmZp7G5g2gxn882sJEVk6aR19rtrTMYMXN/xDJjz3nPMeGVuO
fY1T7cdKALtfKDCWOHufrZG80TKOkFZ4lw7Nwj1ngUkS5xz092UYpa61w6lyqFao
C82Rw+buSd4jHGmSZ1MA2b/f8RLt0ca8UcCaNx046lbUdRyA/H5xko8PM6qDzBPH
1s9TaK91nFFhbuLmGV5WDM1zgUt6iHu+giTsyBgK072dDDgaCs4DVEuNvN95+kX9
piB/Fv5/FvcDWp85zbs+icO0pAHHhLUju+lPITdHeHVvkRfYRH3YSI3dGC14TbOL
E17NjHCggF6PRTk7aHU4ImhTpkTLsqEg/Cc0Bh3hLcW6Pj58JDY6Sqn4rQAOHFJX
xQ3w1xGiHttMudn85tkAvn6eypMBuG4CFH9PxjM9ZmtrFirV64VUe8FBUU2Rdn4x
8oAv2tp1eFUQ0sJTk04+JM+V8UdCqoaM/R7Z2JL1a7dOcDHuZiaZFdqURpwBqeDY
DQVlSNw6Su1moUQ45YyCxHIkFiRv+Nlk2Gg6GcrASm3c+8DtNKihLoMCimbGM8c9
Zcb/q/et4VNSH2vOcRjGU/CctO9vEQTtvUxNoDkZl8g1N0Aeq2H1Y5AKqQOMJuFj
S23rmWzUWWEZzplGuZdVSRpK14MWu8uhcjOps1GKkWVvy/mYUcVeMoe1D3bnh9B2
NPp3G6GL7HO03P/LHvvRBNwtffoY4tqEIyDY4krx8b3pJ5fGYXC8RpkIxZqydmO/
9gGP+pr3i38J+7oAKA6UAY790Lp8iMc6G3thKqiO3bGxzFjp8iSjyqV7hmrybS8x
ZrJdDKFCayxmiVVlXXGU6a/h0i3WOxKkFvqpLxWbJsdCxW2iWrvXfHgRbSPxxc5G
W7oAi7OOZTxTbLYLA7ESVEqya7AF2kfrZ922Ji8YHyucr/OGfAIlS2e64HPivs/x
ukQKwHrQmUv9ADWFrRomqTI3tzlzXzwqhu63hrimE0HTUpiV7WKO8JOU6uzHGCY/
2j/ZVEKLh5atnNi3zkkKUPBQUiJqHFPljUN4t15M8aFjKKqcxSk3GVQE6YOLieDO
693ruS7PfPGxwHRFrtTMiGy7Ke6RNeqBbgjjoy19c1mLVMdqjpCxk6xqUhvSA4Z4
U+1Oqh5jaYRHaqY/AGyl8T+041DSrDR6sVn+xXJkVYiJjzFUqeRjafg3yCw7B4wS
+mc4C/On5VW1X5VeXqXuYzKVNK0Xi/w2GgKvlgNyFQcHEloWDkD92MHFVMhdYXPP
kVoM1/TKeJCYCaIEnhww+Pwv3T57gNEgDKjUN0ysQhGAO2jka2We41o7nTgLzbpj
hwWYaJdugJU9Mk3XQfciyauYMgFhs8tTHC2DeaTZEKE4ICFbKd5JN12PHZ2VA90E
WlCDuVlh6MFuvXs7h/FWF7WTipgnhiKgdKvTFsKVqjaTu8WkvxKypcgZ1ARLSjOQ
ObffmvRDO9x1pZQ6RBVu0+a0BfF/DpkD0ddRaFR3PSjqz4C39uG2OzdPBsa8rjc/
35MLovjQJrYs/cgA5Y0zLkDXcSsBZzYszFr+dOHbR9eqI730kkpZ3fH1VevkFq3+
VqeKkHJC4/fMxcyGsXXkOG9OZf+d972yduTBbJXahiZdvv04Zvtvwp0h0xmdm3bH
n9OQTEFA/h87IuMRa5aU2kVsARCnyueB8F4wRoQNE57azKTMaoCzVnUFYEWzmceW
KKaA/lgmVv3EuXVMwaPUPnJg3p2Mu9I5kqjCkrDLCGQotQ/EWcOcCQDJxPla5s/Q
2P4Yey+ddvlBp1DxO8zwxlOAcAU9OzZ3zaTdsIFZGwmdil/MwogdPwQ9VpaQaPZK
WUQxdiKIrRt+u3dsiG0UwEKJ89b4MIQMls8AoJk6A6ko1jtZN727/TlBPxruqFhn
egrqcBc4o8j8boo494gQGThXqrg+LT/t47U+rMEGkOGiLO2MK2p6KESuILOjVcYr
Ybx9tod6KHmykVWqJ9dgKIwhz86x5KaMI2Thh4vwXQ/30ySwmF7HgUztpQL5PGv/
X0zjOolh2ggivUZ3Z6rpiif7StrDTu9oON1DkVCUSSEPECNANZy0x6ZLKuqG6CAJ
UDTSbhnByYKh3/rUICI1y76yBzmMpMOpWp6l10OO2eMimP+VWKG6Hq3fDrZoJ8Kc
3PesUlIDOcKJlMt30uMQnLhohbDF+qzATZnhY3DbE9QlZ62IKnU/xIpjMrfLJLB1
gra0cZ5Erf4Qzfmla5/G4n6PnMUP7Y0GO3l2Y7+BdEivejaIfjHgg4esCjIPBbly
Yb1HY0GPKlOjitt+fP0TPCJpu0dLUdMDPlYI9HS9sK2yUJaS1bBPe10lgal76kg4
eJJOJD9OpBoFF5JF5L3hKtwBu9L3yLT99sBTCJs5CkmHhSzDDk3QkG0y+dtcPuqR
EG+Ee7mHgrbnCWMwCmbgG5RsXqusAVdOf4e+KB41tO9C00AutemN21zFXEXmv4nO
kQYYAL1zTIWRfiV3/V0NzRppTeJhK6K4V+BE1k/M8p22v8Y8ha+aOX5NyGAaNbM4
oZfqLTCaOCBE7yJ8mtgCIHuFP15XJtX9ylxkCPxS/gWkHXGtpHD1b4IT+JasNVSk
3fHzJyFGXCvaknH3QykJ+28uwilIK945+9pzytI4ETZTqPzF56yiRJV6CzVapDeb
ycB+GLEGHajYrb77YNbVCbD27OXImqAYHzhWVv0EwpwsU3rBhPv0XKfidJ0k+nDw
2GIz8HMIhMU+Ou0HOucX4UMueoLorWvKoaJOY91OCKtyZoKPgXzW/YKDpRLTS+1f
kPGCI+k3cS/4/eWiBaigc5hUU7T/AquoFYJ6jXBd8p9LyJdmmArgwrAYmWUJKN37
QdzaAslQIwKAmBdzOfDY+Y2bj1OSaeLjPdquLZIB4hxPmPcIHO1DrPoNxIKYgARs
SPDFM0hfvWXEP431I9zFc0eRnMilTaePF6Wrb35K7KWs99MZWU5HNtt++w54zb5V
0zqJALbdnlP5B301TLbRkzwsiPpCnoISk80tYVvdACRgsJwEi8xZb0YpLc/Pk6Iy
U0DejzyEUWNr6NR/exiD1NMx2KLi11T5zX8u5aB6NFglCGUcC6YpuP4GPFzjnNkF
IceXcics4lo1DLMLf9elK27xUDwO2FFS2Qs8COQ3Qdq7eNrZeC4IjgWdDHpWzk5k
8d9gYbb821snOpNuU0geGb2q4xuWmJj1x1F33zbfoGuCCkzNCKyXbaaO+8m/llWf
oTejqUStVYFyr+J7ByU0z/lhFFcJ9ZJtGoRGHtNFfASWrgpvmJkeIklQryq3KTiN
cFbYkYRH7JI55G1Qd/SqjdJHJkl4OrM3RNMx/mGnMUZgn7WkZSjXkFFZR+js/iCE
OJq6sKWEbJPOwd2dxsRX8LygJn9IkPb0k/UkdLdhZBLQOK2kbNxkNzn/lElfEwoL
POoO+e64TOlCAdnwDArdaKN0hvgnYQ923UCZX16miiSBgJogSiDVKC/5ZSgRlbdp
o/AsPPFzs1ccOOzfbwA7tFJVVt82Bh61YjOuFqOwwK6GG8OlsOU9p/HvIlviKo7N
j8KtdbdWq5TQub2nBBIEmSS1uOhPxPlmEjmmdWXg+A6K9SMEKK2Qm9McO0lXouWM
gn5Pd5DPlJiE/wIZoCB5jSIKr0E0W2sMoOL0iAFKjznwm6PrgYCmH4/Af3VVc/NH
tvHG4/DYAStGatdW0ca/VimFOw9LcMzM70WUR9aTQgRgFHWSkfqCoTLrAHtsaq3B
PG8+/t6jW6UGSE7JZtj9uhLkQU5f4WtTQrMhMLV6T+GLniRkgDnBwZdoByRQ1a1s
uMTB4BZBy/bN053SjU0R6OCKhMf3JMMvlQlF18oz4JOuWeOA6qV0vopcAcYZ4SsW
7yKMQb35ZW2NBH9W0mlpqcZyHBMkYoJ0dbO/B75Dg+kzb0W/C9UMqxNzA+fS1tBW
AuvBz02ZGOojI3qOIf7JcoPmn5uCp26cFO7GSKLMyiw41E+dLDvX3FW0qEA0nvtJ
v7tptQEVzcMpq2VfaUXcCdqgCjz2pRQS58Wkl2/RctcnbjcOB+RTwBBt/zuuZnhX
NYtg84m9LqJhUTGJey8a7UbWQNk5XMyzYZMBF+n+7p7vtjV8f8ry4jXb0YQou63V
FZj+KDmLTLBXRu/KiWDp2xgHFm1LKa6QnlhcsLK8aLB5ecyufeqnL8VZTYaOR8V2
96PTR/yOVgPqndb3N7/RvI6ietDiKx1S2+A71ql5FmK6gUZm5hviwvH55ujiuuq3
RAuRJtC9wYrMe+wQsY7v2K0SzuS9SEKRdemxcMY+D3WTKMb8MvYJV+7hh6hxESql
cmXS5le0TK8AuHmRAQCAmk4+FkCY5kDn0VyiX2iLicbeCbYG+EJcoqtuFIyM7ZEi
ql/uvnQF/q2C1iAcEm4LPyqikHCyWMzRwQUwkvyCvCjEX0CLSQBnhQN/sOrcQSEX
ma3gnq7xvxtIvG7vmKrW0XH/oQkZoLQiTrAkZ8UkPrOUB1vcOJHZA4Ss0oL8GWFl
x8hPbvANSfV6dtkgju7qJeBag7V5P4gHE3CKJFYfcCH5RHHg8UXlJIT7aXKCDoLw
WuEQvehbXnx4VT0pAwttrHUPrmmLE2rNkqWHGbvlC8vYZBvBVtOKY82+WVerFpbg
bGE8g++ir9k7Vtp7vBIXjKrgc14XBJOv3ygGILZByyd0ktBzE26PkNcDgDoxyGYz
YFSc+iEJMOUS8hITXbm1o+WfeeYXNQFcbMC8htYNVenLA6IDdmBFEZ0Q3YlJQMns
3OcrtzpTkMHeGqtwM8oPglgSmlK3A6LCVSvk1iGvduP1soI0KEBVM/ZZ+ZIxV1K3
CkrzBBtKQjEzI1ywWUaSzwDSy41NBk+DLXwyq5f0a8dSqvnYqYuNdDCqSEraXc33
uwuQ7+U/se9aNZyNiXn/gsHxto/XHDvdmuwTSQVgyHr3p/9h7+Vx9k0xhC7RlQLn
r142qH2lEB2hjtncnSTl/BVUHM9F2ocxlHuOGAEH48+TSGLJykPhmmNl9cXnZDhq
n7QARSKBLgHZd0pm7OlgVppAnWtPQ4fbfbmmLESUxkMLeHK0ph3CRzW6j1YfRXCD
kT7hG3oxi+1k3tdfwYO6G7JeJc9jyRogBQ+KZR/k/yGVThqaidyksPVPpPpfmxzs
Fv7aBP1dS0iduPjpnTtdTrjuYBTtHU3pFyL48BUB/1okRdN/Gb90h5dX9LcfBaZ4
91iuGaaY9xzg4IoaVmdN9W73GVLFHmTLz85ZD+u8yhiBAoR5wBFVbb/hWCelMWvv
Uj0xzyhhTVMCL5nNLe9QnYDtY4hyevW7wHroGEJdIPimLgPODwwfcDlVgdXswcGo
u2pDAI8TfwovvUGKM4pEj40vfS8hJlsH13DiDUUWyx9+6Kx5Syyea1GaXkn1qb1m
EaEdcDdi9L/9MNTZd0pwVlC4sKdpZT3sNX3eHvOsPaW81Q34mKThWzbj8TjqVGoy
68hBLf/aslQoPKRrKD4rhCopHUUJfkPmIgxHLrRK35mej2Kd4CLJE50QgBXpDc49
0ZZNpDJGroGFYO626G8NbCHukg1bpflAesmGgzzl3G7AeCj1laxUNFTMjbD2bHCi
gLXm4FoJNvYJzIvKV6j6rW7N6zcNgh0HGfociVEY3v8TKkSlPxw81YoexQfAGrK9
oKk+GsXMNFRcHwekyqqPOA5Xummg7FMh0aj+cSfjJj1J+MNZYhT0pZ1/EpPE8DOL
/lwHMpZvI2+i9Qila4gX9GTd5W04Ou2zfT82IOZq6pjZHTWlViG7nBz+RnIXHwWA
YCWHpMiFtx16IqdU4wA7XqTJi13y7kxm9GJZWas+LtHdGRbZZovnHpnDGDAfwPnK
pOjvSllkNfoc7+Z1YZOWpB4t0pwllhA2lcaWwXv58zeKs06j3RC7BUNMDfVbr89b
zRjNUJ+barraOV4TwTcwkxDCrMO4KjXcTs/Sb3xzqPI77vGiD7TLJb+JMlVcg1tU
YFuhC0OGl9tjqPZ9FlQqj7KFHijLGvk2ouqhZ7VhyQAAdLnBdVDx4AyfrNtlZhiw
lVW3zyGVtt8NfEp5bBl3jrZXIjqLcrMAa+QfecilXsh0XbEQwYt8smVmt3WR54NB
hP7itjVtpqAPhDWWOM6MmqHmfhTQyoixtRNGzZsaZBPT5yOn5LVCzBhUtyn7XCR5
YZxTJsXBlT39R8cekvks6z5k3mwGS9dD1sJOe4S//qunV/LgF+9zd0Li5uYQxxmM
1RAsWjTyV2LtTUgfHmWd/mt/4DK9At2ClxsGSJ6HMfU92G5Iy3WwgVcavbvzQQTl
CURK0lrBZ13q/gGO/KpOv7K8iG4YE6z6kJ/PvF/U1KXvr4xvQAXv/App5ATd1utH
zBUTuKydLqWDf/22X1MrqjKbAV5Hpm8i4sX11FD8FCobBv4fW4CBEFWVzHZjbnay
PNbD0L45GD4Fe1Q9BytQsIgf6ZWgJOTiJS0noYWpIOTyC1DnitPlTGxPTch7vKUX
A6D3hM6AnY90DlQ2f2oYp5Gkm+k7McnYif3BObMU/c9Nd6QeqArzuQYamXagelcO
8QtdkoZ8KJfriVL1+2e2/G3qKaX6lZg3daOKmSS12nyAKhq0QfmHU8otV6RVYjSO
lhsK1HOhWBghcpl0Jo+745YDI8muA82l3oZwdO9FH9EqBg/enc/VkXuBKHdk/+5f
HLggeyws7g4YaXMYSxvgEAsUoXkzm563M/1OvQywNJgA1KvT9BSXzrS0CacdS9/5
z3Z4lQ6cAIyxdGmNw6qWGhx/RQlymVKJm4hw7gjj6dJPsuVbGLTf+0mBhA4g0449
qDnQRlTiLBTnmspv2l1NEFUriFrkWa2pojb+ZroKaVgNAp2v3KMmYjg8pSVQvNSt
Zyuwx8JERo1xGxNR219Gw4WFfhExdjaUqSPh8nPt6bPEPMg7qaCcshZDrwXRqNWR
Pd0HPn4DFcToXtukO2WdFaJ0r1vPz3O9w5mBGHT/6WtZ+7haeYeJxKeR+VL70hHS
KlmXwrxs10N9cMP4TTFYYtTNuyFIEXFBljtu27yhTyX+PskEPMznF/SpIEwkQ5Ut
KJcKQlOIWlBPrIoPZlRD5tI3YR/jckFSG3I0uC5PAM+nG4xlm9/Zmd4Yop6Oh5r4
QsoplErHjakEAyGkzJJ4noz17vz7v2Z8rbLKzdUCUi9Uh22Xbiysl5ZDbzcI/hNR
c+1/yKn0fFquehZFx7HpjH1m65jLOmhinfeNxJ1AxiWO4KQUpNmqww5A8nMGgiBJ
5PllhJpXEEo7ZByqxmfdikBPSK9Wjq6AEOmsBBll1riII1mIiU9pejDXy413yup3
DU09aU8E8F/nsvKYbgKT8oAS7etkNgdF9xmwYl10Kkc2nZVAVu1wawLT2b06K+Sj
tIAjRvW0dcv0zNOeA2XqIdPemhP2IJ5xAY015AzKsE+mrg7JUFPiyNua3NxbY3GE
lgA8mQJ6Iyn5h1s2/owx72teEQbM2ZgpfpA1eexhECepszn+5eIixpw8xKz8isi9
V+DSjNqjTceZwhjq3+VJyLAAyqstZTs8WkfAHXNH7zD0ArULmWvRhWw8PVPjsbdF
dQs8EBdo4THe1WeIJ/tU/Js5MaC8loKqEPIJW1no4DJRfKmWhcJmHac5JYkO1/wQ
NbYfNBDu1UWkqGGUevprTnUwB2gDgEVGNFjMC+bwQnjlFq+3HLeEz5aG1ilFDM4u
gIJaS4rEBmxZ8olz7kXz4BxWvF0ZGZoGHKX1o6bbC8qxpeuSjBVS5NB7jR7M51F0
`protect END_PROTECTED
