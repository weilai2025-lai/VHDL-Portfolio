`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQNYBq46cYnMeXYxO9y6Abg5d2xfHR00ufkFWs9/4nxx7mk/u5Z8MivLvP/oFJ3a
w3bY/4Hv+vahJImF2ReisBGZfJ4QFkOdzXRRK/OkcYUifmfoAJrwOi+MjZs7sHpp
28AEElcA2oMNV2lEQHr1/t1k3wM++b+BgdWr2HzgCc7q3I5nRnr1FLOCj17fKE8T
I2+FY9SlE5X1TZvgQ2IsloQB9g/j6I60Warh+ogJRILsDudqgItBAx1CAPUnpWK8
jeHmgsBrATRPDQ6Qc870Ip2UCz7k9Vwbdzg3wsV12wDI641bo8EDpc/rD4ZN6cZo
mfCdzaVBuZoUXHC7RmjiVcefWYbaCGt5+h0vZXcxtTPJJSgmWArVmPDexACrMiDM
+Eu5P0RaN4EEe4yZcLYciyGK9jdafzW2sjL07YEhqevBa+bbRD9HBNvZtplaJeD0
WlAvnwrquQCcSoy8gxIU8ltwWgBLVNlXtiia2tZWRcgJDtJ0DMvvzLLdEtWC6AVm
QdhfBacrYHe0/Ba/JKwzcNN8HZ6VxTGG7C/+1yqmlyyEgKZUbzPvAVOX7czUJ3NB
G1Pstw9VCr6Agy7Ye2A9LlUbv/fNvooC2rSa0UTnH6dg01f6WYC5El9fwhZhyZAR
zksZOpEq3gDB8pxRE+g/WxieKXabyWehLC+cP3IiVxbeGLkltnR4bwTQKB4Q/RJn
OSPPcxNREkuWDJX+88MCqzQIUecNOxxQWTrdGv5r+KdoW5cFb2KflLCsWtnwP0Ax
Z+fc2YTKKCNTARsXPdS7hkQmHyzsynTyQTXLQJjvZZT6neQtZZOfuGhDHpB1y9Wq
COjlCAZ9F33H0kwH8ENRtsgrgc6R1iic6XnyTlxld/Ob263Omm+cWX+l3ZOB7x6t
+eynr2Z/G56xkKPDzlTxI+SFqBjsydSmKFSesbXFu71ojp+4dJhsZquXbt5XVqxF
1KlgRXzLddVFWoQDdUgB3N0VkMb+oUX0pnJphn+R2/dcaJGIEvbyaer6R7vYMf+5
7kabEh8ruFnhxuM4xyl9PzgMA4WxP08WgvwebGXtWW+/Hwp6O0urXHPVHBQrebDV
`protect END_PROTECTED
