`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oOKGZGoUKw3ILBUraH2bjbsDv6avX1r189kzNDsrI/YSviZ/zTP9PFrbY7fWNcNN
Aw9rmgnJBH3eDSz0p6hX5vCNWroHa35F8/6IOTupYXthHZfnVuZ+Zjg2jPOJf0e3
XKY5az46IyWGwO+4V/7tvKLfiaeOT04ippkAPRmyfMjiT4KFgdMmL1gmm/Ghg+4A
OPHGtoTxET2E8h3O6CPNejRTa9Sq4L4dtfoY/5YHDfsHRDO7Jtxxt2OCf30RGz1/
E9Lu8HQ+2h6hMOHKJBgo06f+kbj2bBzTzi5hnuzzgWCvdvRR8S5mi4EabolVJFst
3weA2ROE9wFTiimHYRc8HJSXtVYGl3jdjcuq5gaS252OPT+VIMJxM9+DrHKRD2Rv
/aQ6DuoH8usLx7Wm01A7g/Y7+bNThvo6Xs4ARwHm9yIxQGE8buL5SKkfR+D5e7F/
Oqtn5Q5MegmvgIufs6qYJWuRvuhwuuya5rIQogQAHEJXs27bYWYIBUzH8+y1Qnt/
iES2OcSBAkuntEnFQ8BSf/QaknhWhRBEGP8ACKQJIff65lRcLxmZQH4XnHGAEFoW
+SqpQtzdpo6it84ExAldacaSnjDtsnjfj/LGc5LQ7wtZutOrCaGJ0ecVA1LVL+dn
iGJJ2fKRpQgR0ozkxSD58sh/o8TUPniz4f/W7+ewcrbxQsZ2qZlgSCCtXdohHOqT
3NNdOBm2LOqaamYpXjQBNsvgQg83znvRV6raoMjdkwZ4wnbo6G+fYB2l9xxe+uCS
dJi368Kn+fgZLfACalaxGOaBBAxCPVhXBLFRfsJ1Gh2A4d+APWzlajd+rUeKWXzx
KuEaOdkMlZ+LNjYqc/m0proMBAhQIQNkC/zplml2MD9+5DitLt+yWMrC1Z9icXp/
hzMp39WMEzz/u8hWKEcGqxpuFNney5yAN/CKocfm8EiMSEoswA3rur+5992XspOL
8kGSDhSmQaK3VzwGvp0E3UrYNAq6ZZ0kbd8rXSSoMMdhoNuOqqOqSbKPZyGwEJV9
1B2ihFmG13vCro7u45e+tXN4iwvRgRQooJGGd9KWFgoTBPvJw6xxnuQThHkae53D
mwDrPTfobseICc+WTJd/P4sC6rqNCiw1LB4pHXbx/jmOj6NA0lEsxSP5NEQ1PKxl
nJ1XeNHfvJOh31DecOH6IfSP1G4S/a3hAiQcDqjXr2rq/IQibeQdctiQzwT+KAT2
iv3baZwus9AyixedFlYDoMIHJXZGalt6T8cKprKyUmT6vrhTRn2+JSF61o26Q+MW
`protect END_PROTECTED
