`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyFx1KJPMfwEfIsFlB3Vv9QFY0FbRLG5wn+VYEHJ1KovdfKYBmj5ZQvNYTlRM8FB
96wcNARTqmhL0bqVSYZOhGIUS7FRr3CIF2WHzxG4+B0+tB3q7gv44Vqj7mFQXQZh
ItQTAahSz9w7ljhrKYdEX/2Bd1k8hDGSafRiZ+b1gAObbpsqJHTbbV+a1WUtrrQr
7vestF4iB/rQf7Ce4mCc2b6ydYSeydHIElvBqM+PnVRBwT8ZDtUA2WrkShqtgpKN
0igNP9QYuqIMp2mY75ypkXQdGf5hTLBnhXYiQVmyXyon8/f27O41RBuJObnIh9yF
be1fU1qsx1/nPKqGTL68AFu0Bm0U7qhfZ1ZymXdIIt5I4K/zGB+Qumy1+Smn+dqZ
1RBq3x5TSR2YzDlR9YFuaw7bGWwiigQ7guCqSWLKyxouwbvfzEVdu3H1xFXAy5qO
vLW1mf7zIB9i/o1NahPDqmUwcF9nBfD5M45xP9e785+nzdxm2TE1wa87cJfZqpho
AeSs4jHOEg0kHyZw86k3igAbU8C7ZIN4lCWnX0zRlm64xRPQzEE6kp/J7+PM9HJJ
fmik8GA61lsZt/As5Hqx5CCSA0i6BGx9PXabXwbJuYAt39StKu2WX5bOmdSQEpCe
IWSFeiUdJU5vmlrsHJ3zHrxHFh3YQZmEuUzm8t+8YDenZ/olRsRQ0aMcGgHH1/in
YbnMha/bZfKkGAGBarUgxby2JLpmdxv+Efiy9KXoTdtyUq4edyUIJR6t5Z6NSy0Y
p3nsf8Tw/ttR2fG3NN6Sn4e+D4Cj+4DZ/AFvY3TwICUeHt/g/osZ2T8zU0LvRnTJ
yoXGHjGjHUum77xSKmGVWAd3p7cSm4NTFYVinxJ7aiKaysCYOlRdd3aK7bQ6LY0y
mXVpwHU1mMB8CcCArEUq0Khf6wr1THIbe/yvCaiD0XdaMo1VP6x4S3Q67Pz4JUhu
yUlsWy7i3afdTjxcroQJqfi5qlaulIan7wRvoJXPHYV2HtJOx60os1X3uQJOjc6g
M/7TskmIpQXH+ESNLdC/89Z94qyAwymEimHbu5tCk62BmzPZh2jwsqEdwnd2gHLM
n/uGZqo78FGk8gSs9m4gPEuuLEYBLxaSDr4F2RMoxGMZj4ceYFJBB1Mn2ZvWKWDC
NYtTGD6cDc0LzshxP4C/H9FdbT2UNEW8t4jNVEowoXip8FQnB/TseHJ+vz4KyFgB
Y2G+U8QykPk+HSFx9dhJmwvU2EfvHl/7uAhic+6ti5gmWbXFJ7d/crJFqA+4uxTz
4G7G04+iijwiR/3aUqYQ3Of6HTXIa5Gs7D42k66x2BJXQr1/Ced8Nj9iohlTsOxC
DC4MCdGDBjDlqlor+fbuacUhO3TSncurE08t1nvisWQI0+Pkmx5OREHQGAAIPV/s
dfIIahNL4CWYf0tTFtkQrA2JDKnVUmETMtyUMXMeZ9zplVBgh6DSiuYuRWUTY9pz
FgMkQzc7bWXrzoeMfoCRdAOJlRXLag+EXNwal0ewPVmzNe9QhSRF308zObAdx36S
4s+ovHCmBrSiccx9Ts+PUlaSDYu4VqV+gO6T0cmhhMSzYETk5+VQO2gS8+7sG5rJ
PSRmj3AzhUpXegeCLWVyXLcsTXizi6treP/GXBzPto5/nSJju7eivQ5U0RD8LaU2
eGi1fH7Iz5SYbCIOOAEHhkIW1310FB9mNbDNrjsan7CZnqHjza2VdnR6OrHBrB44
66pnl7Qn/39CWDr0ep1KFixSa9nfjHJbLVrSpYyKkRIj5LbNTiPIMZs5Ui6g5GKB
pf48Wtp3FctUpxSOZWmL/6kF5KdPmBoH3eBq6614bdsc9ZvOK79x/BTOMJduJu2Q
+QBhR00odbV7PvkbioMKvK3GETrZWQtNNwJsHSodDXk8G8uH02LOy1dvBvduw/Gr
VaIDtCKtUTnURhfE1b30jYpqlkamJNs2WN7N2uVSeQ4ppOhQKgtUVlH0e0XW082v
nG1JDkG8QgKs7e8nzsKEdaziYtjxR5vNPD8Lzxh2xYlCxFjsTRUXSYX0/jcWERBF
LpR3+WcMmOnOIE62XPsDj8AlhtnLrIZk7D3kaC5sjEah5jah0FgKZ5EM8e0u0O53
5Ypn0SqM5/NAA/z4w4RgecszDxFIjv7oytiMrdQBOTd55eQdMWkT88SRdxJHm+YQ
7bdKI3r191PVNDR+S60oIMnnXd0FsravD6rT9lNWK1mTZ09Af57eNQC1PySAjKQe
qfc0aT8y4A6kNWioFbJtIEC59YvDsHVQEMiMm5ogu5hoUITk5/RTlpX2pqleFs+y
tcGwokdo4lGnIvVCjoOT8pyXiwYITPuynKPsikdKbuQQIdQHbe3P1W+COj0p2YTB
qSQG0VNDL+Z3Qbjs4wELOQgFCfmjZgc8tBbvZxi58gu6o0btLrdWst3TU8nSl/sr
xx+2Pn7xn6HkMzkUGvsgbKuLs3R+Q/NjfpyzVFRv4agM0W6AfoV1rXQ+bhHUDzqi
8D3F7+fTuE6FucbjnVs+d9uIVpw9IS/ahuFqKAS6bL/tiD4qrYPaqP8Bi7ToJpxi
W8nP5HiVvRTYbrO3OLRxrAMAVlZBgGaolNL4X8PbSdS05UjWo8v7fYRHEUfGZHJW
HVUBgXBMAQXtMSagJfOmsBmzGu3/1D6pARdEZ1aglVWeXqYR65AgNuhZLY66rm8t
9aGUzdXhQdqB2H85ZbHePuJuFRArpS+o7rSr6SuCV7SJLJ09RRy04HQRKmvtFUB6
OoscEI/8VxEXihYRN9zNCvrdQVJYPG5GYfpShudBdf6Vt4H12vUyrAxqiwZHYao3
3EM5A4cWNX+V65YrCmLV1WbLDw1uWsBixIHxX+oWFPUmZk20as9jZxLShJfXNQ6O
WUMYnAnl6D0t1Qrt9rl0cgaFpktcTEDqkBGHO9dCxI/XTWx4747xDKXbUw9DaCaD
vsovwfUarkW3xYtK4gxZ+7SjP1PEl7rJlkgTCVmzTexvPwiuseeflIcJG1bl36Jt
836xguRMFgYOG18CvP3I+MsHQbrst6/Wh+at2AIh24gSl57VLjeS57o1j7nvYEYL
21RlGqvdtzGlxeg3Z3M86mKLT8MeahaKNcRcOpR8S793hXybbTjdA3rYS5cafsiI
POnUznvnFY7kgiFmaNEfe+k9Ne9u8C/qRSb3NZ6gBXW031e496aZ1zLuft8SK0Ve
gStj6kClRH+Etqj6oSxXBsH241B2/8fo87WBLKaEGjv6fBCEhoMrcN2I8zF9S3Xq
B8VzceEY2UcsuCXOF7sq73LYf+t/Irj2tB8NAeSL9f6qkgBHhvt9tMhUGvPD0Twl
WE++NCQbny4VqvYk8dIbTZrr/ORJTkSl0bc19vXU0U8qmccgSIbgOS2/c0785ceX
lFcstEPV5tULBGVHX3OeCjQTDvcrLtZ4k0f6QTWcXaCS6p50WkZHT5SWubSze/zU
5nbv0sh66fdbj0zTd/QqInd7e4G8g1DrA+aYonc9/Y4BhSRSxYjp/FkZ/wBDVghT
Wj9bDT4zdrWLpJ8g+lb1n0ICCt0ZgWXUQYquipXKAi8THEsaXgN6WxdvCsaMDmYE
esC4SI0d7vJCnT+BpF89i94biQOzZySKIc7qEcR0tFOjQqpSJ/WZMCv01n2Fl0ov
H8q/XvaRsYywo79ERzySo6IKoQKXBfxeIo36DSKgp+65536vybyD5j3j2gIjuMCG
YO9mt0TyIAmVPOJqD2YvKrjSgByAT67wJpFhCFluQRvVkztpw3qJLOqyRwehSfMu
BKxGDwRx2SgwkkGFyTTi6TKP+6KCaWmekJmfIF01de4joTwlcd18xNUm50bodHzc
zmLnPww77ewmt1+qak02WewPM60wjY/C9xiETL8Jd4P2ZdzoLEeMf9S8CTelBPGD
ESAeDJs/xHuL26QFwql+LwZsQghxIAKc1UKvHdscbX3FwPP3GQtdad2JLlROyEML
uX6jZrSdrG0F0PHVlGiw06Wll8FEwK19HoTQxIHegs/jTD3Q12aFpjS1BKbidBIC
pEgZjmwKfWuGh5oAF+mGe9MW3SmzCwgmjPop5bSVh/VmVYvan2Q2RAaodigJ2d4+
WrdrLEcRws4avgp5YUOgilPAdvv3xpAGeVvt2ZOHq5F8c2yYAcJkjiEGobCODkhD
YbNRygnAOIRVaQtpBQ7P3g6jSxGDsEDzZGv588tUWHFjIMEwJkcST5WkXyvL6W2i
ycfmFjK0W9KlY7aPR9aGC9cBRmYwhy856hhng53jDao=
`protect END_PROTECTED
