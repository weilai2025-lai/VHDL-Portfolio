`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+g/mtWmAkq9ZyFBf1qh0vWqxE7HWn7+YYVXGsw29Lqs+7vra4NaZPnzMYzAAHVm8
lJvbSiGeYPwHezYODzh9CWM8GUWPMdfpzRudnYzjleHbTTcc8aQyF4FF6OQ36KwF
g7jUuJzyiRfXAthURYx1PRg3WVVqDSWD//jcsTkVpWTnrrak7xxHsFrm72YO1nQ3
a7TTdFbUvo87prvUr5CENJa9rbQ0duUei/mvoVtcRkndeMPgEIJrNBu9JDja2/M1
/JhnwokUWNooOauCFAmyuUlP0xB8uvsDqfKDYNCW4leB4gRidBfumnjjMqe4nzF4
OIGU/ZKkXHn9JkcR3CbzrAVTh9MAks4IoxFIxHx6VadHurPBrLBfDmDyTPhHyni+
mHnweYUsCQ1sSkAXbr/ER9I+4+c1g9n1sMlRRWbSR8fg7LuUYnWvEZYB9oevVuKm
7EHJxW7CHnOXnMK8VrLXfFbl6utbPIB7Y/4RYX0NqOLm/9uuRIlpqgkA50zwlemh
pXTzZ0llt/if3bqhrAJx2jvWZsM5Yg9pKGlfNetTXyloaqvbhHEhICpr3ktRBZwo
5+6vnmUzRxsesaBI5fZ5FrdACLdzvD2chq3IdVP6ff8sdEZhzAHqP0xF+mhq3odO
qirGFcv6LsZW9JtA5iUzKDlgN508Z6b1wPPdcsfWR6rHY1LGu/NIfZHvoqvjl8Rx
ggrWT7ThmG5OJcg6347KKIzu0QZsc9HeIxJXx44qbVFPIXfTy90FUEWhbmYzuNAb
g6a1wGRt0HPDM/Z7GzQIaMJ6JPb+L02p7jLVRoheJzZxmmYDnGUqouc57UYHNip8
3ys109GpHYb2KhO5Ls4xKUNg98jFjaEADOhFbDt7BMAMi54QjFCOWk9QxjpLKb6Q
/+TMKH/bzutQPRWdg8WExfUMg2Zg/Thi1pkM4LJOlMg1FroFjNFQMZc1rPuqRZ8k
CFLF6uQcAluU3d2d1sRyN4UVY38+ZE3paRPRT5XjngmoDkbwHLmosW9vaNZMbjd0
P+VEWZOUTlZE7XW4oFIM+XszAo26uxK9Jqz4oQt9LAR+BUNGyN0Z+uZ7lsJWpspi
R5AYTfD3ja/9Mn7WQvF9p132B4Rzq3E+KOr4n4WT/a79FXnPETEiOuLXk+iRZEAQ
4iR9e95KbIQKoaaroJxPy3L/sgfOlkWsqppOkOjA+OVqJOCoqdedAQdlr0dHlni2
X7J/nnhuMoKkUzlJqcC2bqPvJmUJxeeA4DTbD/It9BhML+TpM84SV8VKone1ux2V
XZ7eRsWakXlfEpckvEXz/jEL5gsFfE94iwFyFF2FmBij9xwgE+320VbeuTvZuXBw
i5ZIFylTGqazNoayEXtP90yqMEc80JKW/rr55XH2/8J44likvJ6NY04g89Ug0jTA
LaIRoIolRePeomWo8lrdT6DZ17y0EZepyJ3+sB2IWHgC5H+slbIwb5SMpFDdZtbF
SWaNyNoeQdeyKlk3O9FXcuMQi3i2jvwwHX4Cvdto68IlOUXL8P0Vs8cenZyBRDOz
h6bGFtP54lMU7yu8DiDVorCWAKDRvInE0JWMRhSb+M7PFd50RM8zXkgDDZidhaG0
qRbBYsX221Dwp5QORNGRPkZ1LwCN2Y9dCao9S+2TW/TwYACFu91xeRgYKTZsvTXi
raOF6aCJi1wGFys3w74c4mGlUIaU+HsERaJUFVbFWEIShPzLeZtVAFoAIGdu9fp5
ZLih8hW8sSEHzOD4B92N9AWT1Os97GC/MC7sB9ZK4AtGTv62/TqBskYKN8+gZv5R
Fz72PbxsyVgH8RbHv9PmLO0RVHkq5rKioPIEj/hnycJG/oWJpWRPLi+QLYiByj01
ua9wMzmFxYYB9cnIlm8Zut5IsKm2AtWlbingmuk3AcrdX3EYStOblFi02LNXmdnk
touRuLopurfAHH4TDJPzbeSPYRh1cQIqqoBNdzD/b6zyf1RQlKqzhX0cmNBJECgu
utizG8/mejnWz4/fr4SldOMPO+GimQ/+Wm24ww/Govmth/uJB5B0G5DoU13lIoF+
w45dHF0b9IeWRUBcx+ewJ8yV7pzCGvOwL4S3eBdI14xyb9AsI1ecMX1ffR/vD4cW
7Wev9TY25kRAr1TN8CT+JKJeJ3BhQ920rIqWqeplck6MYwmKcWF8vRyILg4NAXgJ
hkfEkfeOvgALF/dT1qAx90XizgsQ0RVLScx6RcmGd/M=
`protect END_PROTECTED
