`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YsO36PoIkYFfnxgPryVcHMI2g780ch89EBy1RtT/UkKqgsMmriGZ0D7vE3my0s44
2i2bJRraNUMIzV2do3pzel8lp+Qtofs/oKtLZnTd4hGjD6MzlrX7/6N3TL660RZn
aVCXS4BE1Ez51koS5YwzOmHeOW/JIWfusVBfQDBZUyF1OWQCYes3zvvh831018zN
DVe3tSMsfE/KDZBSjnhgqz8Ib9IuKOdUiiRMOSjLzsmvRb2FaKgRbQnofnWHEIDZ
01W2g2yrfj8ERlXcE0Vz1B2/MpFTbiBca+oQ6aiTkG3sa+ernysNxMpFq2WOXWBR
BcTvp2ojwTrJPVfvjllP5mOTcql/pO7zAPlLBB8xA4qLvrefRXsbLz10Qi5AQCdC
gRMn/kLmMJaCwT7tLCKnnuFs9hM4qxecMKtOSCxbRU44jg4qwwjRWIa50/Q9TtHP
nGCbika4wi/HHYC2rI4imcTCAZgzseWSKeyRB0Is3iH0rJeg+Drf/+9TbaDYz4UI
5eAUCJNpnxyVf3Psugtbe2/P37MiDry934H+xjp3i1vqpU+R7QHpp0wjDqeVjloH
QPwrOwmbkjjCY0nNZu43bw==
`protect END_PROTECTED
