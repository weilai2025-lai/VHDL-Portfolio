`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sKGxYg8UZlJZwO59IXSxkSb7r+/VXuj6Qllt4HLWcMqF6VmEL5dYm6igc7yB2u9A
ocuM4FAmLcagsQgTt49cuzkCErcinwHGD8q09+OGIjl3hKnWH2z0aJnXf4Lc3iUZ
aTAl0Kz1tBvy5XHDWsQeMmWfhyxApAdLEzQVGO5AkAYVX0s21Y8ZU/bZF2ImERMN
cqRzO6h0vJSlIGTQiuIJgrs97ozZXitDKxe3MceOFUCZOjRQz42RFTZJBhgXFXoI
cWlso05p4EZafRnCoAGzMXnzfxTgR+NJhaAL19D6eKD950/9p5ifBsGawdziKiKI
p5DSegiMt6qQCVaKOCckhL/nyUEr2wWD/rPi0+2U+nE8cANbPj9ayI/iV6Lk594o
nt4oGH5E/Ac0RwCpFeg+Cy4aP2zGLiVaqe1Bv4Me5jMLSABuUJrmxvZqWk48qgFz
s7NGAhexgNi+tae6E9ewN6SX4AuSvjVLlZtS/8IuVv+R4tls2sV+O03cTcUKXPBN
s64/Bop6hjkCDoldC6Kf5fxE06F7ydS+UUKORzt49b17Ongf8eOrgZSNy7sdEau4
YhS6ytEKjOgC1EOVhdbI5bVzaioQNuZbHJGrukdm2oSpQ3o69vRiuKHaR2vTVgwA
FxbozL8OUslJmaQQZ721c5FeuVWGCJGBcENfkp7uY+JjXwxICmKsapV+YU1e3HpJ
yDRrGiuJEZjQyjVR8UZNbklpY3aMta3/XGx6HpfG7/TFG8u5+quoi0b68FaDwuD+
nKHMe9PykEmgHkDnh/HrmRTSi9F6fonDzVGe2Xxcl2B5w1HixDR0PSRDwByot0zT
Inf+hbOEQEQCkN5ZdNnsbTYL7N8x8YytLtV93wDe6Ebaz9tjwEka8vf4qsEiTl9j
HnXYH6Psj2MI5eAjm+vtHvxFkjsRbNA9Nxv2plO00RNI5jbgcGlPkabkaeG/wc9w
MAYLpD2q4HmtmeBOYbDrfiOQxGH0+ZnpTXFKMhepGc4VPKynfe333ITYM4AUsUdW
nFXalDSO4878WgHWj0NqnzPXBsETf4ZH4AxaDdpt53q6FOocQmMtJqaYX1WLjw6n
cQblkeL5mqoyccyHZ+oL105bA0UR0GKhu7RsqnYMTVjOPcMoJqzB8YMQHVOM2quZ
WZFtVqNYo16QJVmMvpk/WB7/omUm4HHfNV2S08nsoz4CEdG8DtUOUmXB74gLb+Hd
zVkXfRYYrKCcyqfFPJOp4X/t1oIiGVJzeoN2hQJ65tJEmzu9cOLUms8lHNSH6uWA
MQuzXhm2oKvJM9rA29cinKiLNB2RNZAKGpal8uavaWkrBgp+dDoSZFpkGP2oTCqU
RLAymXP0PFmAy4xhkkeFxg0lNv3GQJZpMzfiCOrBhG+mpsnwk4vNycqeRnLaoWB2
R40fGoVz0hqdCctFWHhKRY9zrpVTfg7DSX87U8rxQY93CR0f0Op7VL+IPsN3s8CD
CvcqOyRXcnA/9YpRc99sNd+GLml0Tt3THamqkK2ss6zk0gjSEX1I+XqjkkcrttJB
3Bee4cxybe3unWjItZO8oOAe0gItyp57ER3wgbNYcOtPY89WQsSnaHmnvd46BGyA
9Gv02VhKIyOPlpRU5XBzZn0P0XNPqExQxmxb5f8utu3d3AbYip00MmaK2WvJuBP3
XPXSdSjSoRmCsVCW9H31VcyvDr04en3PXF/yF2IJN8NeQ9ONkrIr/t77pDWOhc11
X32BSezjRHcE08NOYg6+C1e5VUp+xBcpw0I6FUZrgPLQPDw6ARn8x/nF04c+v2pR
fE58opSLcKFuZap5egxAJ8zGr8KPJM0EdoEudYIZ4rV+Mg97/x2e77VxyoMtUA+X
xfgq6Y64nY8ezW5Ge6c7YA==
`protect END_PROTECTED
