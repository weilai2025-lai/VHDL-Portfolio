`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIWY3VYVL3r3liT1Ao9QgPsTjFEadPBEH8dIiRFTdHdFdNwj8kgw7Cd4JpvHNLC1
dIF/n3VAXUBmmZsjCrL3fzqwrtAFckCmE0/WXgZqUvikr+b3WFKA6gqz/qraWvE+
vCTUSUjnHZoml4Ef9g/rJHsx3gP2RRTlH5PLftGQPQllfSrNCPEul6Q73qJGWMrP
dqgFQWfHDW1ridyoZwTum5JwLeKyvtHRsIcdwTwlWG/DVWMh4vZ2soAQxn+SWl86
RXTXVn+ph/k505EO+SOQEnnz3mY1kcewa2qGoblAOKTjWr5gwsTqR7h4wgZCHIC7
UKDoa5SVil319aBKMhd8jdKpwDNBkye26UTM/KeRfd75W9A7oAy1JAFwVWYtuG05
rN9xz6dpllLXYfdcGlkompJUX3uuKSg+ThBfe4CK4QH6+0Ieaz0qnRcZCZV4QDyy
TDpxcdMZw+4UcHov5TL/CF0tMPdD9nRQQwz65FMlPYJOSfRfdjxHa4cFT3un0uln
vljf5m4HGm+eXbDMppwLY15sd9jw9CgdeTpbNxG3QTaU0uVVN2Z2gIabSKTWJsI9
Z46YbawagwM/1vmfUoKAd/gIt8zVmyt7L7uNQvLmfu+03SseWGd5krGj6p28v+8X
yOhvc+fr1OkfjgoGne1EO02swfoT4y2rD6z72jWNZKBpRAuP/K9kAg8rn0nU8xrg
p4N4jPMOp/6yiTJuvqQfiuhyhgsKEVMSV3NllUvD2ZcK1yCr0Zu7Zamyv3JL0ogY
oUxhGa0gjawRjb6L1kARlsdH2UXZN8ZeEi9xsNzymjphXKyT3k/0CEzH9FwmW295
99ZXNQDFGH38FzFxUFBRi9hzqCTPh3VbdFt33XI/njc=
`protect END_PROTECTED
