`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O3kztwinyQ92JSFW5Ep38xv71SDQx39lvXAhznM+PJHpO7+Y2bhJGjOAXQ5IL506
yzQHgk+Yn19nCSGxfUo/W4QE1F6EHfgyJ+7qG/tCgvAwH9PPGQhtUiunY5QYfHZA
QFn9eQ2gR3r2SL1qu+rPBxa7K8YQ/wLSnyQVX1BERb1J2AquajJ6UflPZ42myRmH
sw7o5WmQiPSWkpt58CsGgDedc7McUcZic17hEsHvVExNvLO0EaAzjeKRo9U3zr8z
/ZZfi1SrTmJZ4Z/BXOButMXXOjjIZMUQxlaLqyCqnjfpWvb9qEBWuTo5zpP4t8xg
+R3Bl9trECKz0y4gLdY2HI4oiQo4qVEiZtmNhOaq5R6Is/4qCNXl6SPMXZzmc4Hi
ZFaHT/vYH384tojG5vaGZ04jnMBJ6p9QkqIFJGEDBKYmUGDw0k5gdi+yt7LH7Dvq
mc4X0xtedDs74iYF3t3qakjpZIw0uOzMKdCc0H7bYaJSI3wT9BxGMM2fo69ah3sb
v0ntXw3R/Jp9ZW6uq6Bsn2cAMVeQ/CMr6THa6r/mTfIHT31JI4NQ3xx5THgxigFf
NjH0piCzWQMVrOKAPu4JIO8ykIE9kS0ukSz4ZU7nKyY3rw06vnOMfs/Wdx9jrkZY
KD2D5nUW6j31CuxgfFtQkvKG+uMD3VuQCAC4MYahOJ064XOU5ZRa6ZhLqt/P0Nez
5EA5sg0h9pbDzvz4Y62e7GgxCFpijx9dXxdBBakHRgE6+7AzA0UJPprkKxxTFBJp
qeTlq+iQO82sC2WZFf5uoVtKPdP3D23I61yvDqEj/6/DXRFmtXExRVuW5oAMtWRA
AyepsGo7zpkJvmg2EB1p6e0d2dA1tYYoI3izQceD4Cf6mt357e1vJypOXgYNqFvS
Ph/9Vpv48HoBYkRdg6UX0sesSda3cXRgWOF85xGbco6NBHhjIIuD9RNDDovhyLaQ
JzGPSzTQqw/WW9G36sbedCJ2/JQgJRwN8semHfzD3ZirLTRty1QfxqmViHLRNzie
KmGDW5Jf7aVAjsC2mFd3qrnC8dkWJDM+EjCwwpMSj7NZhtZI4MVoKZEyAEAdLmT3
kjyASrh9/6MA+WCf15kM2hW0OHKkI56KwpK0Pr9BimoMqx69csKd/VIWrpDrku8w
UmWD3EBZv01T7nXOtajpFkeZMYkyPH8BNx5XERNhR/w7SFBs9kgPRgRfStdcZO7V
9wXDV5HtYNkdgEH8/3J7SnYKQm9vzxs2bE4iC2JAdb+Cug+b4Y1lfQ5OAQSHCqjZ
Z1bcHjB/9iaz1SNNSEMRSezyzva/0Brh925qnPEEFcUwo5QsSMmSczAUH7XflMds
TI53ALNX5tFICZql9sBL7z0ts+zo3ffrZo1QjH47iXyRUVJ8uQsU9tSUQwAVtzCc
ydJa0xZvTO8vr82R6RtI3UdQbJ6nImpANsHA2YDk03cs93xTPl+7W8aWQ5jzE4k5
zIbHZjWdy0IY0EQPHGu1BiaOiVVQqVDV/BOVhB9BlCBRkoI0VkOv3dzd3sS+wFRl
qxs95+ES0YN+xpkeU+4QZXVDc6wzdTXXhvgIGx62EeO+5B2cTwnzVSZ6e3nkcnc0
y/49n/deHawTNqSiZq4dy7nqB3zHe0cDhr4tacGzwLzvZzlMORAVJPF5k6aTi5j+
+MxnHfHOsPp3585awbsVcz+kQBzFSRdfQA7aGFUFuYho2ED+DnyTrhUcWrFG1yJK
Cnirc65sQpstqC4yBQ+y4R0miC0lLQkZCpUnwplTB7KRIKT5UjeEWbVrzh5hfpcb
TMU8vdTORTRin/q4/gNB4d52pNPeydb4sECOOmCknV84ExRwvbf5PNUT1BM60vvZ
fLURKCPgXAv41r3k/blc3qC8gok24shiwKZi6GD0DRWAqeSmHrBcZdxCF0rOmVr4
Q33qpVHXqq+BEk+ukAFYMbnrjYJQQ8Y0LGWKtxZ8valuAugAeCMPqZU19+3CSN7r
rz28BcubeL4OgS7BCiM/FkkfTbjkae4ljcYyJvZVzdcJFSfhWHdO+65qHlryF4gN
lh2bWG2znMlLUohoZlC30zScoWSmSHaVY1ARIpgTG+/kzZ830NNG4zSVSn0dmZ7J
Wvirf70bpdgaGYJndN5xHYerFML0ZSZZvwuMlukwS+B0VgApYTR90FX33jOsbiZd
DD8As2ggDB+ZTtQl0z38EvEq2w39Q5BPYG22iCs8zkajjAtTqZO1FSODBlTq02Yf
XAz8XSth1uBNP/7uV3VRjeGHJB4ovGkTYTW0X4HYngYj4V00tge/EjhdUP5f2kVB
zc+Egsg0kG5fJ6f5VTBWgEKn+1GsfOioB09P2NzUIPrVISNxhDlB5RexXGYjoxO/
2ybSMEz7xVisgBOgf09wISAHgh9+vgeMGUUPCT1LROPw7+1pY6DQCQ29UkNDAj8/
k0mGIRMcv5JDoKDKPzPzMMIEAvXw6sYUo+EjkX7st2jrVsrD1h5lfk/23mhNhETt
HfINHGcixVLKatE8OAfUc0p64E0kLVzcGaQdc9v+I+NLNAGTiBPBDf0keLBx2FP7
UE5qBNBro0cjjUpYS2ZF3wYRFTqSsRp4NddjcuPHxp8YKqUTK4SEp9YPdvcrz1BW
iu77yktO9MO9Xk2iyY7TvFb6EgMIEW0t8djPUHvOmyhpkAIs9QC2ZnJ/JGXt9zMw
c1Fo8ESgv8SgOCQZSIMPIGk9lUiOnHVkW5Y40+LilQBCr31gS4UJVJ6bPr8G5sv6
LQbu/BUuYRBqDm5GqCjHxwaLoU3n/mXqvkT/RrolPgwsoY1HFZkyThRJ+vIQ6UUo
pusD1OKsRASQiEqPV7h7l1GdCc3B5eDrQ/HwPXfEC3ADVq5NmDRUhOF1Zvs9Zvw0
/was/OC5xtfVS5gUqHJcQm4ev4tgjHwUvoASezE1ltlvHqdRURh2yS39yfh3IDBc
Cb2sqX4Ouw/aWH5PF4n2I33NgAu+uCHiKOw20WJR5xXkF07U0fFMIDkJKa890I3f
4EUlWDoXf7Gf3cJMuVc2xLfrD7tUdbwrspQ8U5SfHUtVZ7KCsmr9bxQaBEQi8XS5
U/vgUeGNTAE++94zsh3LMpS6jkZZ3hw7OsH04wZkBUiIU/ZXRmFQn7EY8qVMpNqn
8DCbPMe/+KGg3leT5w0yBjFeQ+lnWiWn0hYIeyn9GJE5V8QsAJYNDAON6D080O+v
F3i5NKpgOgNGxLdoyrRff2bZSLuV0ldb6/hkhrdLKwFGAikiZa1nMnjjABQUFOVd
GNUFH7D4V/TyHfeMkvI8YxhkQPph2IYsHGiIBglzt8e4k3OffGmtM4h0lUvofmUr
tTSYcue4qAnDz6O9g4SPJf7zTWneTeaxbyd+4CQkC7LOM4dq8r6uvNjLpyStQ46H
MzsywX30MPhW8b2anRMosQOnh55+Fh7Dv819LxCRKns23TC+2Tijcd2Evx9hMU5E
7dE7r9ynNQ5tmEN+GQdwUZJyHbjc3f0/RWIKAlVr2xFM7AdA91K/r81tEPXIhbN2
/MYbueAE/Qs3VagsRlHNc+QH5DkVbK9fzL4+MXD0GDFEUO4Ni1vTF/ONxnLMxByv
6/yqUhQpgbwM9lXIPpGX53YnErcqI3f/BOus0Ly+haTxYD3pI8GodRTgAkaHVfRH
xZGT8LbngXc5VZGN9jgwsALcYJI5L8MzaXYHjewmEbLAC3AaGOb7o50hqMrHEVh8
D8jcjBDG+0gMgdHCrIi4QEfDJm1sThRmt97BUTRFXO9NVbxOQ7do54PI/ZBY6MXc
YZnPgcaka5/xcZ3tTw8PJ2fPAufbRK7P31edViFej+C7kOOXc884hBb2KQ0UuCb+
T0RowmTzwc4SERS2Tz507LHATVewQxEcfRpxx1KpBBBFnSWx0HUsqP3BW67E2hIN
TdhElP2/fND1PAo3EbYZTs/6TpclYeQ1Vjg9FYfIIhmPx7XXH6eAR2eGjHdvNLvx
+G97JQ1nAzXblpopC1K6/dcM0+kXWCChO7oVKP4WM4XGK/ZIzbElDB/4hKmlKtPK
ZUw6Ci3tp8QrKwdAq2ecKTp7wl39C4XLPyReGvevpmkvagZ/lpRJ6FW16QtRSSfy
vZOqOv49c1VBeqVBZXnFwt+SL/qo0gvfONVDEzFhYX0zrksLO1z8VjkK2vb8trMe
TYQNLRtEGVS/ZbbU/pNNUAg8zQlK4CFkUTNTbs23pyqXgWD6hrF3cutpAKizY3M+
oO1hs5mnDvYAC6FU2zY7u6zkeRCk3gV/8qudJTtM97YRnAFC9KNVg1xjaYcrtgvh
nzMuqZKMI5P3rf+PGPsN9j7q10dDJUoloo38uD9DLFG5WwNSkmuJrJK7umUzf2Fo
DuorvcqWMpx/od9wxd13C+ms0ejJF5i4vyrCs+ohnrL//u/l+gfXRXkzJeSwosrl
35k8Y521OmKwDrNG6dNVyrZdHEW0hIX3sa/rlcoizDp/ZzMqiSwUj2kNcjBj1Tih
XTvV9YtDckT0Thar9QUz0dAjoqmdJZKsLexqEEpQUp/hEL8AfKzal+SXwVe/ufY1
aElNQYqGQHCzy123uG/Upm8PzzN+kK/XHtYAvQTUEUhmxmOOZjJboM8eb2H05DyY
RcugArsGygxx4IRT4dt70XheTySKA0CGfkYiNNPo/G4fUfvPVdOpaF9muN1djQmI
QVXcbb5/SgckFXLI+YCoXeslWfm2+l8z/xn6uZ2u1RPRw1meb9VxbgRuZdGUeVoi
iYwqy1JOpdDQIEKBeuRH33W6OwTMAA07l933wDmRedE76e0x6UVWLEVL1Bts2eB6
H++DUQMozAVwVKwK3+3NgncqaHZVriyqwIZcwDOg64liby8kW4jIvLozl5QLdud4
eUYfK4xO7NESg3nBDQhIsUIf30hi4KQGIcRF67vbwghnsZ8nFTvG409c1VEBjVs2
ThUY4Rq5fCsl43KfNltHQXs6J7OoP54zPPUb5ACYQjBqwAMN2NX4zLSJU666mASF
weU5lijMh9FfDzPCdvjiX06Dw/D3nzr9xFXE5RPWxYD0eFlfb+bu8TyIk3HEbqZu
FpPTg+6CEfDq8CmsZvQQqREUGqLf1VnR6XkxVJdSem1x4jzfajNPowqpcluNLBtz
TMwj3g7P1C1JczAcUVMvyG9QlrDqhqfb8NP2VdkBHrlKozi0qMEBJMEMs5Obqr8r
7rdt6bDkcGwal+RnWFQEtH3Mf+V4K/Hj2fdB0tEbo4Ad8Svy/KcmTj7EkVoLH+wS
LvH1eHMJ7ldsoKnc40q+YpmTPVhItd7jGFm9oC3T2PS+79pCeGNmOQ7pNUJy7XyZ
z9CWHOFxoSzN8Y19IMkc/RMdxNHIprIMsVleqmvvoNyfk/3BznOtSdg3KSyso7CY
xWBpsr116skjeul0PYmE3CkRTLR0GbRPjYprmS/GzNgLeQiccDwFwKgmhtLjBSi4
eWo+33zUIsisnwn1JuEoNVuA0COo4PULL5hiKAC7bnwZMNaZSQTca3mZQIA3DNc1
geRF/sM1zx2/wXWBUqi7CecOJFc4VWuQDWXnqQd1zCFe0JOm7mPWXlgv5PBDNJTC
nt3OXcYdw8BBRPQu9TsDnu/xYsAQaKge/IZDEmG14MIpLGjno4zRKD/yu1BDclCS
OX8w1XMIzro/whFrPyVxd/yX5hccRFBmWvfXU7knL8EM2KmW62hqR4iapmaEKSdQ
jNpubKPH8Riyokw1hn+zYKBtF3OOMxEd++xDVxMNG/6yaFujDVavPtwNJpuIpkQs
x52fRZGEA0kWvJSKvaJnoNmFixBCdBLA1lCtxeeMKhRwacirGO3fy9T+P0oHJIzY
QNNy59CiO4XdxeR+usF0i4tfFgNn/d5ul3VBDSjC2tyntvNFmnq5d/xjFYCaBEfY
IbOT6LrUMHm/h4ZSemXgEcfjLSvt3iQvejQLkmK1s2ifAFxU/cvD7ZHkNJ8R+Qh7
JQtUQb/yyoA/ij4HkntOwEWswfx62uSDEOlME/l6qycQ4TdkD6aUbC7M8JtcIxVP
LSKmE44El3WrTEtcel5MbqGoj3PMo0lVGud/lsquVtPm2Qo2ET2nT4Q6VhvcV6Wn
UpYg9HyULXph8bkVVyws01dphel7SLDgCzhxc1zcsDXr9ablG4lqpfn/xkS/0d2Q
NIPOwiYae7DPAybBJG8A0RqAMfgCLcfN76W69Ajqnh8hAsPPyxkrh2+k9yRqWkl9
xdN0lpRmJ0jlarqGDQ4XWWbu3fjL0JaAa4P7wGzICbV8sol+eW8jpR6ySgG9/1C9
IrCUPtKPxOeBl7RPB/uZ3PAEgPmoRk5JTOUeq7Ihm9TMeuK8eV2NJvomvOmBYyKE
hk77GasXN1Jz4iz7Hbz9U1PnZ+llpQNiLp8+jU3Y47mSjafjQi/umotoNZYZhuH7
fMDNXfMc/P2rGo3WYRfZ2HbnxFu1fDv5QZO/w4G5A1xEvcuANd2wErkfif/AgvZf
DysEuvdzDJNNjihE9tJRP9K2ljknnwx/uAzyACqSXu108Pq+7KNwa8w344mYAnt1
QDbN+ckCVubl24xl61SFJLDA9YrMmlVxtzwupamqKPOvR6ql6/IVUmFXW0R4Y6Vz
+5tMyVN6VvfjXKTgRsRoLig1a+9L85dxpALs7gyIykqEW1cLYtYb1PV3BH8e1aBb
6tlgNN/MlCGkBrUQe7mIRMh/txRsUWb1vSpIV6hIBOQxsenxLwDk15rJ5ki66Uwz
FItNPJDpvkZqaT5WajeBQNT7Wk9jG6hJjQ5eQ8Bk2Fa8X03C5Gx/CKyN3e2yJhoY
Vefnpa5Vj7gR9VNpNysId40iIdPoMq1/F3yt1MnAeg2rPAk9/3DfHnxGlx61KrXr
F9F5UnU861Y4qOfHgvzNqEgPBfZpGHa96th/Sb8wKm80jaicg5t5Ku4DnSG5cEUm
X3V10XslFoUSniJIhXEzWRiYBNoJN8f/HXQwhYya0ey7ZqCrhUHwhOawm5aeli0M
x5KTSUeq7nR1fUVwSJ98vKnJFyAOySQkrw9V2/uFbEr+SUF4JOdrWNWYbalLeQWU
/5iFsNRpbmLb8hzCHMalcilt/O04XupTVAzcTd+WAuF66edbrMJ/cSg+q2Qs3LrV
RrxmOwa1W/4VlM5spnI5X9ZUm+4eqqbHu1YsH+0C3jruPgOLNKQ7lllFyCGKB9xe
skHUGlqAm4ImFRxzuNEaxPHbNhfnA3aPAxw672yiWX0DjEfxus7dCquDSA2lAL6c
NIXcbqdJuj6+/dwbQdNQSPrwPrgKc1kOUMdbsmuA2qD158PFHz/nE8mEFZw4qqYT
4oZlmsS0Y87TQYdvuw0vAp/zVULhmHH1ZfoGZE7tcbGMUNiqPTjFtSCRXr+0oVLG
V7iydCbzY+JiyAj8ORyEZD2m6gEnT97nke2WD7D+W8CMjl2lxRS9KnwPGdcy/xvm
i3bJ5zbXSP6WOtw5YLTmSnq/jhDKXqsp6B5NpzlZLSyugC1+JmcKQwsvTPbA8LGp
TSINaowOUiIQOG3bkWQltBJ6S1wt0M5ebXNBMxT9+jIzhmU3xWmwAGV6lFyjJc3O
aoCPyacici6OyfsGtaymi6I+B9hz7Af7zDTIqE+DJF3lAGqcxMRpgIwKzHDblLeF
u5yLQs4fhM+3jaRJLOxATUZcm20xsAHyCOASmz497W+c7i8hsdF9muuJt4ferKq1
quDZSPh2woYFKuwR7ENhcmjrE7s19fFpIYYci8pOhB0MPK7cVDTOpBxEF1jtiV4G
ps9UcqRB7LfE4NypRHwEUZ6Dnw2GoqFT2rtIdP9F1eI5pz7oxe9FKAL/E/sDTDTK
Lk5WH1r5/WLGNnt+D2CoXIRZy+5JVvNbZLdmeyfpSwY3OQdtgxsgFT+PHIP1bbkf
CsRhcu9SGHNlYXN8YetwFv41oH67rTvQlcTc5Hk9dzz7I3uMl5NQhb683wtwdLAi
yX0viHNbjREJ23jej3kle9kiMLWsFRk1eiZDXEZZsea6qCj+y/dNP0wdOL8cDiaB
hevLKEC8YVJmtyV6HQ5zZqZLvzWoRcCu/lgmtxosNpk=
`protect END_PROTECTED
