`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fTgusHxOosEzwi5wwWVjhdfd/vpxA5DYiVq+jwRdPqYmMBxf2hHAAAtIgEhQcCK
dsVjVDxyDAfFQaNAkuRlK1b0B8h0ITVdfm47eWXmJzQaYdhXVUm4YwZhY7km5HKy
ioOwAN2NmVN0setUehv5MN09fY2XHtjvRAPExhvw3+377vsRxMbkZ8WgY/yfvdZ8
hSCEng2EQfWl8J6MSbsQigMvIB1K//jzYOjLk0IcalGFE53CCikHdtulf6iu5Iiz
6TwHLj4ifXbqQHeL0U1K0+LbSLqUn3Xgfuvv9wp8SL8TaIBFnf6zu/xNABDGJ/bR
7UcwAE5nH07/iNCrvtuftHk30mAsx+fVlP3H5K/j0TSX5oUEPIN6ZoP2kcPF0dZ6
sXS36GGaH4MruvN0RjGcMWhjrFvU5DZk50LhehMuiV6xp55dtHKbhbKr8c44xKcQ
PA1Ap8ZaY8CX/HmT2kBvy/Zz9pwE3s+W1s/UOCHGm4Mz3MnwOc/qteuwXYMSpszL
xlfXA7EAYK42ymyIRrsozyySI001xZDT6nBGnatLqDV1iKlrvZ5ytUSSOZMu6Too
t6xbqgVCkR9a7z8YuJHxzvclXddOaPWqNSlrNzPMKKiW/DC8EPKXeZuzBAMFpNEZ
fZVwcGr7E2mnTWMuJSAWv8zdQJIwyMGP5mdBDpaS1Bfqmzm9SNWTNs5Ikwg21z/l
fFxofSj/QclTwTwv1LmauFJDBxTwe9hLcBgIDipNpH3+br5eVyDmaNfi0e7UGjJR
VcW0OcwxV1QFqYHJ5cmEsEVRQSDYm5nh/8qUKQwiJGb6jpV9O38Zo8g8fsJzHcRa
Hy6SKgSNEysO4k99AmBbGXUB/Bmx/gJPcYblyHi3ENqiKS4RkAg2NypyFi+beyAw
kB1ky2HaHHKgkTm2lavexdyYOxLiq2i8M8IvB+5yaHZn5zBFZnjM332Y7YfOD63g
OiZ5+P/BbmBte3CbMb/ROsHm3MoXCSUT3nPNOATuUVgnhaJJTL+DaVc/kVdTYYo4
tnZ0kIBxEY12d2YcbokueiTkwVPzD8k62MEYpGFOEC6uUgg0GLvUeYYwdVA7YkpT
LX2h4izb2PlF4dSv9q+dH3KpEqZ5oK58YJZ8cimVQR/g9lFDCqMS6WJZt0uU//Oc
DIeyIX55JNQNAHHRxlekiMpf81674xIiwZKL77TukR1gArRP2a/qj8AFbNUmPCmM
+Uu/9IdQ7g7PPtUppfGfawUgKS4KMZz+mhzsP/z+emky8ChzFbi5sqs3jg/9xKO3
EjUv3AhGeraTl5GMBk5YmGSgxhC5n5Zh6boBBSSewMonoIGLcDo8BrFegmCDoijp
rrCcE9wGCiQA5RaYRRK7OTuN0ZoZUG8YAcNUP68tCgvJZwb415BvfQ7MV5V4goSB
ABkTUDcoEMYfomlwDbKJ+PLVihKV0Klvq1OuERWdcqMYBBi6oUTLgYRudrkKUtbQ
bQP/YRgF6O0tW+Ad/73v2qT0BntyLbjNp1J4+YnEcVCzdr3HfijpfQ/NcWLoHo2a
hEUUmE5qvMb3Jf1MhhNadtJE5GcZkK+vEEim9VchXjFfhU7rbPUbGj+KFNo5WUef
KjwrZgTUITYuMGtMjKkBRW/6lSkRMmRNg9FpC8aU7uP+PLlwm7js2P9XxLFHBi6r
xIT00H5aTl+WY8QwTfgDkPKGmAJZFeOv+x3WiHHjdcWiblqVTbBuFP5Ap1lwKFMD
GGXEvNNJlmEApVwS0pGJdtlKjrqzrKu0+nGlPyZ6DT6LcJzj0f5nQFX1BCQx3BBf
yekv/cq+6NsTD0kFbyAY+mddSYT0aO9yVJkcuujTkiyzH5Z/6yptzHLXCVhGLK7q
w/B+gwj7k41g8iS6LfSWTEUrJn5ce1cT4emyHaa8Vq2Goio/XMt8iz8oRM2j7Izl
szfAkxljVToTdlUzWGiv9D4jGlSl2GSuUtaZDaKpReEd7mQUl/KeaImi+YUfRa0v
6o3KAHX5P7eW9lu27i7mM066P8Skz5bUojaS9m908YzbiDf4mYiherljOlwcTTLR
r44r6ZNZy9M7pv4X8hJe42p7tJyoQrDrgrNmADBprFSCCzGA5oebmPnY4DnOmwbS
3mo6X0bOfdJvumRJTrMfXA46RIRMAmRkx8SfZfVLS5MT5gQp4jPZ+orx6cXNKEJF
LWmyENT89rrHT3EX7QiE43DoYxP5a4N9krMgIgJeQjHER9UNp+bqWLqgyufBE5ls
bvGZqqRwCoEZ9rjy5t6mwo7qMihYcwSiMqGWHqWJa3LmV8owsztEcctkDRIssBLb
26SEFIn050zhhIlS9x5DtBgedZPYi2LNY2n9H2FrOs/uNMjCu3WEiNLnZ//3et9l
KwL+tK1VmAX+Sk7kQeV5tORUOr5drCYttrc1Ker/+hF0Zzy6yA0hWGFfzL4moCJ+
B0gb7K2sJM4dzWDEpBGYNA+4T2PB7hsOCyJilK1UL2OnuokNmI52kIPOqmIl6YSK
IEkplNx4FunWjiCpVTm8JYbINFt5u+FIE39qV2+l3uNNoZpe+krSlOB0XYDTHUKQ
jd2GNxtXtYGWnaICMBalISffoefmgawxDn6NwM0sKcpNWs3e0Enjb7KYQvEkDteK
kl7wAyTsgQwtJZz1/YTanHsMkc+qLrxcbrRbLKhjFh1yFwyIP/0rvok+oiUYMwbd
1uabsYoOXcT54VvIvp5INUNYj6qzYPRB6RxBnfeYrtGwCgyBVurwPtuFeKFoPioQ
7H1TV7XajxK6eUXOzjm5vEmIouVTXwvHORKQVxQWhmCv/4elly4IALjjLi+x656t
+5r70o1JCPXpFTdzcM1m+V5tJGQaciwip9kZqqsvN6z9wAnuJCs3PJGyYLVQXJI7
Tr20zA1dIfAj7d2YH1gOGuayTsoI2CnqcIOIrIPcxYGOJCccC6eaUj7XLSJfNOn2
1bB4+cURiKQmDs3Xrzk7kLMaBRFc1eNdx3641HPJ98MqZDbXGgYnqfBQ+Dvt+B9o
tvLkV5GE0dHRgH9BK/81m0g1N/3BTM9Hk3RjxsBRXFNWhLSz+1XWxjXKxMcNuJZe
zbBp154Nmaa1s57fKNg8hN8MXaNPTZ1s0ZGsOoD9X67IQyAqk10aoIhXNme4R6Ab
2GKIWmaZ1BU246p91LVCK9Kp1P1xJk1nkNVGuEqC5275Ynfog09vyV2EOcPJoT2X
yaDHtTbCE6pm4d0shnK8iu1qQPJqXAV0xKlQiMP0eeYcLLSpG8lc9Vt+4ipsFmzP
WbBT/3PmM51mGLVMteTlo1AbpnZUWf2af9Jj90v2zA9viZawZlcJaejlykYSklYC
ir0nQIuZ3LWWo4YqtSEYBVRh+ifnC18+meFS9ZPwteVYIIqIFRNuiAH6HSU1oJdU
XWNFsasX02oxPQr91mzY4Erxp8iNbAN+NyWibbzn6tZk7vB+qbdkLfcgUZnHuV+q
CX1YFjwBGyPiUxJNTSATs/Tk8Ozrysr7K3ZuzWp5xZgW+adQhtO/s1+vONxYuWdn
OevrgzOpoXXa/uyZiOen4BOKUYEE1lQ3cxfMXkwUEmEC16dCDrewBEathwkaJpRS
Z1sZ69/cr5G9piTMhVA9JL33FJi9twaqXxhp1ZMqqX1IotD1hR0CVVfEzhzYYvfR
orp+uN4znFBpb6U3oqjh61xslTh8fEaKmAEfjg3aN4cK7uxxaOHqaRbnhunbrNVj
9TmRDK40lyECdgwp5thpOLSxZ1z8G+BdNmSJOitKosv1asNFGQZpETYoEN41PbWz
hVwTcvTa0Z37hCoxm9PeXUC78BEqM9Nz8GPJcK7QsB6hlo3nkSHSkJ7b0C9higIM
Tr3nzLlM04YG03n+0vU0Pc0oCAEcUgYFp000Ec+d2TIkEe8LhquXeos8y9aVoU0b
/7zYI85V+6zSJuHGOVCqsex2NXvzijxQq581v6PgoASH51Z5LKsmyoyPVty3ZLFc
0g/C14aYe945UV4DmUiTcenp0RPyPti7UxPrUJ9O37sdS09ZPnGfBZllKhvxwq/x
A0BhbnL5Ljp8XEp8iwIKiOEPuezpIc3SKPzk56Yq1Sd9ZKJ9MiMjSWbuUfWZ/n/+
vfdoPJhzlvvNIyJUXAUDmGQCnLU+WiLKsaPVwpEPYNSHBEifnGXcJPJBrVtk10FG
`protect END_PROTECTED
