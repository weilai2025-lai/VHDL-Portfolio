`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
if90monCci2lAk3vSCTjc+p2E6RC+Ze4cXeoee2x9046xeQebluKv9g6zasH7nc6
d1K58GwHAxnj+3juTA5bpI+p0KzKceHpJ7EI5QofyPYnkJJUjTXmmejn1FM2z84Y
X+vrM56SCn6JLuciY4qBEH1vCy3hv/IbeN4/CkiS2iJFxnlL43JZwHnDbu2Yj8Ay
XQOVVv5xW9EaIZqFtJO8tDw96Eq1NcFE60eY7YBI9P1Tc/Nome8VnzeFrYjjLUO8
Wc+6hvOwTaI3cJy51lVhWXYr+Outj/bK4SupMU7UhGsRFcJpUXOobdiBuZMy1Huw
nXXh3N/PqgQUhTibOjkoDhyYVq5/rTRj6vOeedkDmVUtjmv7B3s6PWEhxDQ7xeMJ
RwIRzXRsxzJoKw584qsPQiihbw3Kf59qLhuyV7FuETkGvWLQk3aFcN0djFMGEoN3
m6mq7KZdtyE4EVCkUmjwOGWVYmp3dnNIAF7+5gSuYNtYPbPCRCHLeYiFUNS1b2sz
X2Jwj/aQuS8kkX/g4/m07xS1M4cvdHALMz5gX9Cwlacx+xKy7e3Qt9BwDSqZtMZZ
v4mWDfLuOos5ZZoNhcYvrxCvE2WOzRqaRerQc1DLNdJ89J7+Z07dAJzzx0KLqlAQ
icIyQwF7UPDIaToyCRr3+ReJ5Htn9ZpoGhUqZI7Y2WB4VqILPEN9NKElsdwnSoEM
nvU2kKh14dtazM4+fzFI0BvJiTaxyt7zfR8SIDWpeihX3s7I3NuZUVYDVDffjQlM
tbAan8naNlMS1JP6ky2TZ/2bxrJ6BXitFLDNJsJGzAEXgPyA2Qg1r7q5lgt3P9sQ
rIetnHZ6B/JmaXvaePxNn6WD6pHWBwPk8RqvzM6286PcrqzQiRdmXQbLWb308oNO
+cPUgde06hynEWn6XG1n5wMDex8y4Y3tMgxjskr0ZPcgtua0Xxv4iIaLd7IQwSff
lGLJyL0rwyvD+AqMQgGER94GjFw59drIMrXTqu6E6ndtB3ewK4impWRPoCHT286L
JbgwMadanRS/8WXvvAaSmxt9bcGNnq/bD2GoCAwO7b25dHB/ZULCeWruEjGLfVuO
Nr9uobnE9+2sBfBZMU0OUaeJagW+MFM5oycmmCyf0k6ru4g7Q/erpxcimW/+kEZX
kbvAUa0wxuGoWHaNRDVkmyD7fTORt1HuVrp6r2zo2EbNeLedPDChkdl0ZxXjkdkq
RDa+opGUS5in9nz4pQq6kTDUSr7PAxwsZCpS9OXktIpQCTPeDr83N4tnkyGQRUcu
tXT/+4M78+hJd7CAjUUGWgHKd2spEi84AgUS+e/cSkQ+XrNt8j8MfZjSACOCHLAM
6ujiK/WvOhZn71eOuI4O20HtwUeMFGWSVV31Kup1y74DVwQutwwQR0SiSwIn2lNN
j3Hb+BA34YhyZsb7+2PPaGpm2I4ohie85jNEstIwq23t/lgryzoP8AadCH4wS+wY
YvS8aLR5GUUQ0+Vzm9DPf1Uq4rxjFOVfeA+dad6KmB9lHFQoeokNKy4Oe9HQJt8v
DRdzYxhas8A8ItqlXpUW7CSnX4aeNJt4HoWN1jnSycXAR7xqvVg3sxoQ6r0ZANWf
XhO+vSAz+V2ASnlMmDZqnSEVKdHgedP6t/IE28ns0IrDwdFiS3Gzcwiaohyaq8iR
s3Hiw0kXjnq+PGJjd1yaQhL+S0yzdpudq+ZwwekX2FpfiamsH6akMTGe6JOPBtVd
koYQ0cByL4EqB2RHMmCZD0yxUNEcZp3qa55uT9RTOxpqt9yUa8wssOvsdWWnE8BS
egeeAPgbO9Z8hEvDlWIO1/B7KUspbB40ChZbupcHh3p6g/U2qoh+ialN7LiEadNI
83fcsiwlz+ZQ0cCmUJuP1vQa4tnwkzmr52eMEAdinbIUweD7sRI4p3rLr5QyA+PQ
YrhpJfxE0puLvMecGfzO8sN52tZhP2oZxxO8MrQFY5pI/E9aGD3qmHplVq0gFTct
0X3aN9xCQ5x1q9SaaLkYglubHkmh8n6jW386hKoLNuMVkNbQLTDmXbKdVSHGFils
y4/OYNALqMgI58ROfoY+exoQ3/SdkF1eA4/M3rVVmBH9Hn7NdkXXG1tip4GUGUhc
A2NR2+kiVor6KCs+Q1Etn0hQ0RQguTSuv30xiL20Z9K4uXOTnQhxUxP4CsXL6qUf
jVnBZ/YdSSwHds8tzGFpYqkNxyxrSDnYSvi+cMyHN4gOkWwu7ebwwTSa4J5Y9cR2
TfUemkdVjgxVPu4BYOFOYc0gGknQxbmFdNT1TKhEUl8x0qpneI9JPBC75Gpxn7me
M8T1k3QMA6bcMsGENtO0LsXvQ/IU3/CGYvzi3hb6z+6PO/t7+mp8E/W0HQgctkPa
I9Lff5k1u4i14/jHW/ilGo5kXb8iHUea+wdE37sE/WqAsIlBkQa6RvgK+Pob6Afe
8q1w+mzI3qkaONbWc3rg7Mroj3I8QFvuPmyTudth/PEDwKKFV75tQJ/pqTMoY51P
fJ7iu1WD7YXxmGqQimdaNifb33P9dOnxBKh4u+tOWBOoZhNC3LdfOwC0LIOmYHBF
xspxhdzz2bM2ep73ucolmSRra2byP2tmyHlpJOwUVB7IRfkaXm2EZXP4RvPq18N+
PjgIMUhb3ZG+Sf+7AhCCCVL8hqQPLglMTmx53gsyXalqllqNGKwK9fcroqi5k876
JGEI1PUfnTOj9MoZNnkgmzB7VdgPahjAwFCt0lDgKHCQjs/R9Y6x2dzYZA1yj7sj
mG+4mrkAScqifQhu9WPv+KWQdZXjohnjy6Q4nr+rjU7QLvykqYRMFoueDyk+68bO
NnCRMl+eBGOU9uFQgrBjTKlk4qe/BxXVRElZ5dBPXlTN0i7EGYBVDK9XC1r/GtlQ
vpCNVjmucJEaYfOEW0qGPsbn064BI/RYV8YV7o2ha9kUvWDoMRnLNskQicmAYNpX
2IeuMQewjBy3tuIlbGMV3VfBVOcD8Hr7IOLOb7KICiXQZPLyfprf5L/xA8v6qaS8
79BxuyPWrbkMCieVrGHxIfXzeQxzG5sGOzHFYLC1naicDx8JCPFchvxhq783XMM9
KuCFgHoLp48tLiMoD3E5TiQm5atyvMLebs/nekFx8WdEN21Ho1FspiI39dW7M57z
YdV815EXrCaK8nYMi/aE7QUYYHAIXWp3McwF6uzTrk8I5MchZmws9XiURDLyF3q+
qbtNOibo+P70VyyTrzQpmBThUM4QOfkDFYHzVIjcTjSyu0Bd3S0lWWuZFYdT24Fh
J2qWDwx9Cs9dYC+g9sgLD8EyNSeX9iRwJPu0TfWGzdK/pr1SN1Mf0X90dC0alrYK
OJ1lwfXpMWFkgAY/J+1GzM75+dtVB7mwfpLG1Llr52a164EqpdCgxRBXN0UM8mYI
TyPpFTA0001uqXczNBIgJb2lD7NSBHjoglU0auJMEu1EkT2dOYu5g6JZOAncBv5x
JE4eIDdElh+1JTfDiA8198rTZo9LsoejTgkMie48T1MgBmfAV85Brrzjrc0U1uHn
IoE7xoynTASTlYfWgbi5+cw0+4oPTehBdGVpjc8ovUNBs/HT7t7eDKKY/Cf7KCPU
D8TxEHfG0iCU6xfmQfny5BGZEZHJLI/fVHPogxXDpC/Qmlc0E8SVONKzWv7Yuw9a
1gCCKcGVkH+eROKKsksbucs9hCUej5AQWhANwxLxVGhy8kQBeKv7ZYs4ev9b7Zj7
mCqRXfJ76CIxG7/itXQg0Wdxr6m+rSuaAq0Y48qvaYaS4sVnrRFeFW62jMnvtRaB
Aq2XV0DMuiG8CwidPzz34jSZwjaIdlg4cxJcx4V+hfE3xH/ldQh2TGKtuZgyHiel
NHdli5V4jzVbrs6lZZy/YyTYYycgXguwxtqIi90G+Rfqlf6XKU35Y3mOq6IExUzu
ti3nh/oeevt5bVQizyQf0GxVvi/YzB8GoP03to9s4xgKpejwjrUCMzA+ijxKb/2g
TN+R9+VhbG0k/Y8rVCpJ42yOgsiVZ+9KwVoZ8ikeDspX6HzcQf9V8ZhdANnrw94h
ZT5eJf/AQQGnIjOBg8hxfzrT22cz971JxF6kbPABg6LO4sCuLlUkDKgZFais3cQ3
u5V0emdCsUW0Z773d47mEMrVntpX2nJ5NLY93eVqXShPOh8Fo+Bb6t1M1gmx6Z3w
XwKfLccgH6htWBIe90X+pdp6sS2JMQEz5cZpW5iIDJG/bfPz9aE8mcIZjWDkowE/
34m1Swr8Gn5mULaKFhw02+CWlQBrzUQ9XAAfJ5ccctrR9Oj1Z0NE5Ukr2qU4+b2z
dBzfcXlJaW3d4zSCQLtfcufvPYusgZVKY0aAII36AjvlSoBTvQoVWmbtqcpzvudb
zay7uT+VJZsHWcAfL8VaYtgNIlHpfWNlBZK7O8H7i5iBbEB1M1oEIM34mvvoHDYe
1Ss1cc55p+VH9GVQP8zvNMgK6cXe1A7G1WJEvN1eX5fndaMgIWPuYURT62MV86wk
c/xyIV3KAcWIWTWxqE3SrdLRQO6oEyvYjIhcBkN9wBEuyZQB7KTrXbB5ulB5qlN6
JHPeY3NBhvvZVFrptHWI2MILj7yCEBuKNVz29lXbNYXos/SlZcVSkU/B1X9Wtgz4
I286RLs+G2vTZe1MueOBhblP0UR3Cv8+jNdPT3vtICS8xilH+o1WHidk4T8mfmX3
2lMqY5rkkSKsagad0zX3216XN2J9DDxoEmdbZsMYUVY=
`protect END_PROTECTED
