`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJX7GULYVa8HIvTlDt5zStToQfgLNfoTDcS8soyZsdCqLvcDxeP2fhcqXoIq9WIy
nA0Sw+NMDdSNCO+DQAuKw/WH1TvfQbDFWArusUsVP0MzB7WW+xiRjQgJ5A9ULZ/A
e5TvlUV1g6KZx5IA6mS14Q3qME+kar5jPFaIRY5D7z9NFm7sXZgtDl55FUEyJo8P
9UluKc7yvNUKOmOIOqmUIlHBiQ6MC5zUl56cuZ85Lxe+VON3j/kpZlqnfDxhbZ8D
K8a4VfBkZbiZRrvPX3rAZ4eV9J4Vfw1dtIx0I0CFs25w2oRoJVCkBT65xaxVntKP
uD5vB8IsLpOflt3FsT25ya6CbrXNmzqgg+W48pE3wsL+coW/QD/lIFXrr/8I2R+S
N6epKXLPZoxfnyDEHXiS04Jih/tb16v54wpLPWM+u320zKv3o3oJYcn2OM9ntSav
JMs2Fu0D1NVdbQnROx/4E8yytqSiMVxqoLl4wgX12QaRZCDnkSKodquriH9IJJhS
YSMXUuIpKiUNLVD5g8X3Uw9wisQdGn3y/raZqzeHKsKCHfLZThnvvgVHZKSgXYSk
XMAsRlx0Nzn4QMOCDPedcAgUIK0MCfrKWY8M5dkISQZOE6MQM+yBccPHL5iEobgF
m66+bNyiGJkSSJtkyXmEn0MCgSd7gVPb7RADc9Dg8NR4OLdCe2WFFojUhnHCfFEW
f3KS/fnrC1bZBMXYDY8/od5Idh6SXWVOvF+HKscWudtShdkZyjV7a1Jpy7kzp2p4
f4AeQXrGd2V+AUeLfX4f0/HR3Evwj0M4fkY3tbeybIHEcBMMtLT/e6T6M2ROTkvg
Q122l5XBwCjieihLy4eoFZVkokj5/dMpf9hOkLcuzkdAVwi6bLx5uOeCw/VEGd9Y
8aLH0uYI23j6PNp5y6hynsXxQ2/dITcvbhV7EKGQrNlHERoxripzVQ1zKT3Pykpq
3mbQBBHiee64jGwV9uFYfIVZhp2JJTE27oX/QKu6SZZmvU+nixc2eVRkkR1loeSd
yP1vuHLZByRtFSslREX5NkMhjVLLxq4k8pFoVd1y2JMVVpvCT+bNDJKhDkyESH5P
1jTRecsQh6TJbzRp3D4wWQ==
`protect END_PROTECTED
