`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pb8SNYNVDIb3qIXKbmJ1UtX9kpSwhv5T/yqmSLiQqcGn2qIIIwjGWkwbOAEBrNoT
20D2dha+kH3RNRXnjoe4VeTG8trR1hAgwczUYAI0iP0IPEjhOfhL3gPk3Q7J9q79
N29hHzdhIk5Y/l9FoFrkozckQGSOfKTaguf+7fYwNIHGtmKnacw+U5ZHyJlJq2y8
Qz7sC13gmELPWirY/IECUpkylMp9Uo3gk13b2ZA2CZvorc6zYImFRLw/VRPviX+3
o8/ma53VfXlMmFgSn1fHKwcvJwfTnPEcDt0MgX6HPTADnyP0IV/Ca4sNP4Np1QKu
ALMj9UrEmnOq37PHa2M9zV8qNydbbrdqRCgw1YL6wq8FbZC47rRtaWPne7zH2Kac
00D3px/Kyf/gsm0tJKzWjgB9YCH9kRw6A9n0TAwZn102Io4N6QxVACGK1S/aOg3z
ddVNkrrLH1agtLsWl3DtlobcbvsbhKzyVh/6kMV2KGRHbC3IHP5g2WAOI4hNHubg
QsjDbAmbhJwfXjW5wLs/O3NktKTUAzAeJv4/U8fwfMKcLPTaXJ5iqWg+kMq367tD
GHT++q6p7k5ZNEy3WVbt9vpI41P15F3yTf2NgCVw2X2W3GWR8MsAH4JFi5pWPa25
gpIACEXpoTVg5HsZkyWCYHvFj0P00cKB8lx9T9BkONwXAKgcmdBWRrEPrbrRWW+u
1gf+2zIxw4szju103MgRRIWRpe8b90I0OBCNQCBWHGvE/GsmSiyslpIRVNlc6QFf
a7TGJTcFCXgdWgSuNMyBy7YuFaajse/19yUKvxE8x5oCleMPK7yjYm4ZpTw4aNFx
ODu0Hre8qOJNo+vpftXlwgGRkohacm2K59JvamTLXrXygCLGzINSHb7SrCMui05n
59YiiToaIZ+IzIZIJiXugGfD5I3NEAB2pRsjLurEIcOs7vnWgEQneovzGu6kInTB
WL9ae6HPhh8uXwZzV7iU1Hqh8APwZzjyxzd34/KzjLEUTbxF1Er6rfwmbi8eWyzd
saRAaJvWbcuWaZCcjYgJVg7THXdyfj5eIg7bLsp92ETqPOClfep1rBbwWubxsAa+
xeRWUS/Q/denoflgKRkXpbLWJS8GqaQsWKLsq9DoAdH4F9DICdgKpGXyuCpPyBrK
i79cT0aNTZ28TY4Vo6307uhE5TTptk+wCOQv7mjo3IwqgsZYmLXlFvZ8KOeOlIQW
wlm94vR+XMnxwN1ci5rgFHc9KU4J3qlfkZucBF/sgSXj4j3474IDO769/PX2Czma
wlnrIdujLmIIuG4IuUjNTkYwUygHnFbXT9Mlqn+dwA2FDYnrxOx8oikuV0f9JniN
TvjZHnR4F+YX+yO2SmCG6tpX7x59GX64wmNbSiQwRYkr1QQhmIukWY3IvmeQ7baL
DcZX4qjyRMQ8/35CygweKLW586c0jbnx57d8C+WDi/iAX2endCJhfOSN2gnuBeIZ
yD3jPQXudFdeqwqzsN/iopnk7P74cwPqGX9EtjHxolxfkahAj1eV43gENPIRjTLX
8KaqyzNyyQyaBMOz+9qPgU6Db9GpG4In55n30xszK4eFbgREXmTApfFIKqZbMpI0
Oqu+BStf/+6kPhoq2cMPiVLJs4EO/Z05XNfi8a6x6aUjRFxUMScctQg8tJQoB2Fi
AWq5WJdG+iwMc0wEdt1vbiMbgChRX3001IDWeF+U0F4yixKQtLRBoh3O7NYJahVO
duxeCgj/G5pkhJC8F5ekz6q0PL4G1o1i7HkId/QKNAexBxHtexmCp+eNxKYoPOeD
Xm5W+AhHUcB7czuthb6MWrsaw29Gp6I6TqATF2AH8AGbzBlxdS4Q4gOQOtegC490
M7laaNA3ju4B75Kp9toakn669HF0ROfZcMdx3UyQchdNO3JGRnAGM2w33ZF2Q980
YzI+oGvMg/yf9fHiq71NwSqUf/Vq1lNVoGa0f4p9rv8njbXyokAegUFsvt6CzrZD
dJGPMBDLvgZSgGW/4mxXHPDa/vi8SbX0eXOB0OzySILW85rVSHMNoZ8BikwCb2hw
AB9m+25e7YFsdIu0SJrG8ZseHwkJ8DTRSRsaP3oyDzgvQ/hSfLRaeCSmwJlJbZGy
6DDC+OqaZuCPG3JmkTtLJ8o3TNMpOVjcvrnr40RouKBV+P7dz+9mbP2IDz6+cdb9
EaCHddCK4WaLJl/e8JEXqkQ40fyX10knfm27umtDrUk2YvZmSSp1f3XWUJUL5Qm6
gZSvclDLHNxsfzN3Yf8X5O7BxkDRCfPQa3BG0I888kC4NH+UK8HTr6DtZsT7Y48a
mSXNKBfJed0U/ze1JOaL/pTdIuKDBAV+/gcr72Lf7i2PzlDqrS38qWRpl6/Nm5Ab
Ls+lXKwDP7ASyCO3rGRSy93wHUywykeiTM4yg6YbwrHTAIKFHmKcSWmPh3V1RMD2
8/GK6v+uIO557DfQ7eVaYuqvnewUj81zcSj/3InI0BaFAI13jkuVWKvt+MN0tdme
hyHPNM0UqSSwj2Qp8lD+gUcf1skVyomEZH/W1o5j6tB3/W5dbgJE3ylnOH06BuzJ
CKQcmiv+G3Bgd05WsmRHDpAC1GyNzxOlFsrT3x7Ashfqlbv9ZMVBKsIJPPHO+GfV
Y4GQFgfEjoSKBcCSb/Pq+SNkdGf7a/iovdx+w9G65dCaGYZApYlnRQNHPg69r1bV
n+ySjHYpWIOwVD8JqXwQSpIWdGL6hb7nxSVBb289tjZZF9ujEDtgzAF4qle2BTUV
LNyHpZETj/fWTZTW+CnlmDRh8ksZMqBptE5667OxtyYPBCGD7IdCtdW/3idMNJPY
2MO5gPLqCII+7TJeMfrajF3l+5HFf1sptT9i4A8RCFTXoILD0wCKBynvSaiLXSY0
PTbSD1/Tlcbo/F9Ic2Tm2Nx8+syXBma6mhh2OgjqD8hHGA0U+EgwYFCnbtR5xgEh
BChT6HQv0f7JUieAQ1ToqIofPCeaSmH2pOof7tDEuJCn6wUsIUFIaqd9bfiGkKwW
WBd463LW/CYD2VjDvfiD+JN+k2xbYM1YwTzlNi3KU5Glu6gXDeiddFlJgasTXZce
Q5JSfsK0i0ggUcPxGKQjy4ssjhaqdAt856N6KAdN4jFxEBrYgJNgQefXZ5O5h8Bk
IU3aBWg5/2/9zkoZkIgLHfvTUuRBzVFf31Bl+yEsPsyYm/JGS1GCQIkcI5Ge43Fz
d+UaACpmZBl+OjI9Uv3C0nOD+nytXMBHy+NVIOXi+PvqpnQw0pjCKxpgW1yXmsq3
nVtT0vSJkyaBzOSo3L8fJCM07ywXN/DWMxODoiZW5gW9FlELUjQumar1KYC/u/Tu
YL0sUduExFFhV3vYl2lEAYFKNkACw0hTljFFZ9Cn5HWlDoPnQFyvAzMJmutQuRcm
OZ75cZnDtavM9ViduX/DyDK7/mhp5Xr7pDdFbLHU+g+gqYfNL8UdHIXab1VEBxpp
9tqMPhk6yQjUMEysk3tr5R6m5+m541iHpaorEiJvFYRPoi6+sEmK6XUcP1D1pAJb
eUq9/Ed0Ew+h4zoBXFBKuMsumOYJXhKnuRkiiE2rGYiiy9Ns0bw4kVnslv/dhJUM
f5YY14dn9Iq4DLYgjJBU8LQgCH+QVJc+mAB1PWSnGhO4tD1qS0JchWBCxaCGLihm
xW4ir/KyDQ2cF45zIzlDifx/b9r2jN2y5A4OyOM4Lq8TkzrAFfflUoW31g2/t9JV
9l5BPcASFsz4yA0A97D7+e3s3tqRkhNRlxpEbdVTixFyVmaUjjOnWQejap9QsU9F
RITbT8b2OD5YrhvGkycglERNsEgdWjCf4RekMz97hgYLnosELdZ3Ff9u8349VX6X
Pwri7oEBgc0/w0QiuK0UqA==
`protect END_PROTECTED
