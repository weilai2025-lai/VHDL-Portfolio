`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpeCS7t6xE66cLb6xZTXsqddmsHxqJppuO9o6efeB5uleSLVKhPPpcNYtLdhj1Ql
2N1P1HjpQp/744IpXphx7V1uOKn8FY7fmpvQIcDOnqXyNyWPvrvv3e06Ho5CGnHH
2J/lsnRoLKAt492VWeQAurugjxXWSc16B9aoj+5Ivnp4noiaQZRo2jYsHpxcceoD
bSbv0eVeBDPTOdJSY7qJbxPVtkvT+uvfLQAYAr74WxHzrHj97XL7nLMw1NV1vaWp
yR/RGbLVAfJEulxWccKxT3IBBx2a5ojMq7eBcPQgn/u/Agyd05hD0lVtuXh6s0Vw
b9zn6RBdPEtBCBj6+4GbZZ9ClLuyglefVy7Z/9zjaMNF1sTWLQnbYQp60HQpShWv
+K7/C7HEob2kyBYMyrTZ354zEih//YQNuMsXMsgucTR0PeqEuQh13zo9WYyl8ND9
T1a7EiVdWpsqFX9ts223ZeXUSurp7Y4+eJAF7j3EmKBNDnn1wagtgytE3e35VhBe
vlMEY2Z4DjxY3rRd745hbiJJfmwPxXzYccYk2970pv90VJF80hD2pDChK+8XoCKX
+l2GLkFUxS52/EiaUjSz/McQD6Ye/VIZiAKSQzF3izQZcC+bhW3z2r4bdLPK0N4d
NmPH58e4/kGN8zynsdq9TwUsIjKSDmxEMSk5XYJ35bN+EHOWBC77WDYvmbd0nahI
vryV4cqTRFZ3TETxmUzQMN6+WUsRdfK00BcvxtUpzXH7trNdCarTAvZ+zOdOXe0f
tm1pmwy5PVTdMiRY8apxASqd6A0tWrnrVG1X0J2iShKAuY0LFMMjfFi8gFIx2B7a
yPhwgoAFD6CcWuwstXlQ2/NV00rO44C0c/NEFxP1HZH1FwW0ZTeSmlEqDF2O9ZVl
UsZucbufG+Yqw8rAaC1Q1cIY5fb3xzLWemibF/QBLs4cg++jTXxXEhd2u2ySnwEa
x4JFon+jZjixSmVT2wxM6uUbtDl1vS3g+blu4tkh2lWStuBOXWpYxWKyDhh0duSU
obDvsHWwgOlE+zYdAqusDYf3Kkf/4igaLqxhHxIkGZB//FXI8I7CDh0kJSbC13kk
0VyCFVWvL5rfjbegIdR0zrjtDc4sAp3A/jMycdJyW6gulJJr5rMNXvQ7bJG2FU8p
6ltye4DFBeU9pK0VUMkG3W4BBk7FNpNX7TVZRabJ0/8T9/sTop+1yKFWzYvIfi03
BiOnVVQ1v3GloPKCyyunM88dB2OIYMTTHYGJR7YHVnPLHomBYC2eR43zB4zftJy2
+g/HBOF5e3grxheWdO+5LtNZ6BwNlXSKeugP953YnLrhWpVqh0FPowSglXtRAzji
1f2+OBK1ojOuSTwQ+r7XJpHsh5NwqnXAL8UYZumoDtL7Nnfr01COD7yWNlbzSaK8
GY3Mq6kMQocgzzPM6WMobKOX34B0UDbtyMjkvi5zsanMmhh9ibPRsT9BMAQBaFuZ
09M+tfGqil5tGunPyLaavHx/NCLLi8SpihZLN7Dxq8GnRbwpFRI6Y4YzOac03Hwg
enOQcNUBmQRU1yAOpVMtyH+92BjtFIPaIpluGMaxOLXjcBiw8ByiUgbObODU4Vzq
+QiPjkxXHN8jjEXsBxjwyVrcYC0bnOYWz7Y/ZFKtIb4=
`protect END_PROTECTED
