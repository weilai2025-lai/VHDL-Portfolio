`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hXkACrue0H4O1C6XCpFww9jsC7xUD2opiSFdmRP1OWNb5AQNVwxkMRDAAt0vK+0
P5h0k7eNNt/6JwEvQA6jI6hk/xCbAmTdnMmt75yfhcVQsipmI0uPRcmZ+wibLAaA
FuubOkwgjzi6KIaHAjBq6zLqtFUkbFoIxTZoetI6Mlq00odrNXbcZbTVxrL3nuc0
gt01+ulKU6/bqu0DTNN6llyE3aO+xKqhSPKagxHaBsVuRSHjW5EFdv2o8FGqDRyk
wgyaocyqVnT7JB7CGM3SUFl0XiaOzUfspRVZ3ros2KLMSQawpCAtyhtB2IGXe7GP
Dhz1ZkepusMRAROTmo1VM1e8zTNqmrOT4FPF+JwV35W55K1WOWc8c73URzssy/iA
aE1ACoi9v7IHthrBUoejQvDcbozyr0klzf8VL+wAzKf4HCCyeKa0wWwJQ6Pnjx5l
8PeBDDqVWx8064R3xl/A3SiQZGe27vNVFMCqIcouMqGLMBIRXorTTPnpuHOrOCxh
RlGRtJCbWNlszbhwZenwreVyhUVd2fcd/DkFFQtDDKx3vwAtI7rqG65dRM9n6/yH
6xhf5MxVNQxg51m6p1hJfdsJP0Pm4V8BfiRnAiH6IibO3k++sprHUddoYS3wZQmo
SHw3H3smgTX7DUWMKW0Ob1GoV1af55lKM0F6TGL8rkZzqI4diyXeTXyrBfn+xpTm
o1ka/Jeeimu7Rg7fekD1ou3ew5v+Hytqpqm1TKPuyysGIiuBW6E9rlPTj5zkt+x+
K433txMf1k+Qtf0OhtBlfAYzZkHN6FRUimxqVcnUMUg5mBvaPq3C1PgYSzndJj+V
udD/zLqPdALo5DcZV2cQ+oVUDzbqpChReVDYEed6rNUGk57XlYcrnqnPE0zmm0g8
VjTXBJjxz+ENJ0SfjuLiki70pmaVgiCwR7DF7vuHWi/9JQrYG7vFDPYI8gwLA1+2
FSDOtx6OPyXCRoZ3YxKNpo4nYa6YftGFVHrY5ANREjmXPWErT27rGo0hykff3j/x
T7TujRoFP0StAsfme5oebWQe+/YEvIuhdfHgPRJjWMQGNu7qqTt3s0Xm2QxBW4fT
N72Tg3RanN/nSjH8EoJseYF1XIBfcgyFSqV6B9DhbliXJEtmwhINWwoS1lxfEnvk
ZlmAWKMRRkvPlChOVyS9BUrV7W5J+q3RQ+SvGos6wboPDKv9vMc09DhNXYJx2HTJ
qa3KqLYbfrAD1lTGxLKqvVYy0KvC1bX9tU4CgeFI+k82XtZeUhKlFGHQrkmEYsn5
RhOmZRXQnAGLFprZ0ZlkuOvirGgXEInNAmr51BvEISr2l/Pfy5QLVwkx8SF7O8Yi
Eyh3Ry1Y2T1gE/V//cqNqMys2B54t6Dmiz7865XfbejGcoXQSljhW+Suu28Rpthj
PIWZwFNZVhakqgelQ7KD8VaMn0fZKeW/tIYcyWhdgBLfHdJVlh11Ri+Rwbn5XQ4p
3Wr92gS/4FU9c0zesVdKyxvef6FexsDr8UlZkI4VSfgZdWytrLLQfxEXoVk8mzsS
mDb61yqPMYWB9cYI7mIRULVO7anIdScu7dsQy9b1b06Q8vTQ31szr7Rth5oN4+Zl
V3EqnDrr/hwylCiiIqnmlLrlGyfuQ2HSY5Nk7/dOwrhPyDLlbDhPHZPi46+zncji
IfCkHTwj/tKFfmw5Mav0MhVvD3i55oJBTUl4vUtvjsa0oqJXMU95mFhTbkC0E2jD
D/ntEQPzQcPkcIqcPQ46UEYaA9/eCvu8gtBeqyOuKxk=
`protect END_PROTECTED
