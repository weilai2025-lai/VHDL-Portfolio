`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EubovhhkMLr3DzlHSfMJkxb5rpaItcv3J4LrKPJkLJ0AqEmp+j4MF4ud9veiDw6Y
gX+GEeiUN3syqUWMgVK/ENACBJK1jQf3dYMnRvsfOCVbQKKVd+k+cMeFh5nTEDur
MfRcy6CBKfXWq1Cz1IYNGmcUwhFSNN0/jd9AYPInxeYQ5B6VL8kk6RWv/JjLY02s
fHhRMs0W01lZYE8wVZxQxChqP3ULqH7pupMEQX9zZgxzdxQhHE/iGR6+6NY+N86x
rN17t8GRTMb4Sl8SsWL+AHPd3H4hlFBlog8/mjM9xMRZuhwtc080zQerSg5d8dhh
V97ucl/CKeCkJ7xcvAKLDyaEc1U1eR7jHMS7w0K8O16mb620CZJNxzF/0gHu+MxG
BEL1GLrnNgKSrFm49Z10PjHuOf2f5pClyxhZjy2ekKxt7C6C4t/Ty/DDZvX+6HoH
Th8hebHG1Kxx+RkWUTQ+S3AAKx2byTQ6BANyDPc/ZDLwW8pdNdk5wZr30JcdpNuI
qAKNsY5BhsTo9cWyMKbk6dNPZ7POioJqFxOYYeQ037CKkPrQBbECZFmUUbZ0U70C
6tRxtKmXyhdgJ6DsoSYu+Jh8HCjV611hBZbGBr56aQu/WfAHRcUsd7TqeyrVk1rx
qfiGTB1m2eMbh6G2pJzdCnVPxLzDn/MfmHelAwHR/yQ=
`protect END_PROTECTED
