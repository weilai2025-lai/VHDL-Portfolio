`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abaX8qKRUp2DBlgu+pVmJduWEVXgzjrka8OL+GX4jQ7Zw4EcPTQuiarH/g5M5TU9
pyS43s27uf2yS6ndffDEHL0LWrsRxkVssWuV8eZ85iVHHwZVUbrPeJNb8ACo8uZi
7YmkpSp71bkGFAj/k4QGMaAuGp9gX8T1iYTuDsOthsSLsQPB9rXEGYMl8AYUIbul
urnbimgO1592IkX2ldQVi30wZXwrZ3vykhpQouaw1U7nUe07XWZqgu0MI90y7Ux3
RBuPX7pl+uVRGXQy96yh+EpJLT8HI+E14TOzcluc+ZFLn55hrgcYFjxnFyjH6gmu
WsNCmByV0BmWAyKSCjECA1/G5/NXUWoB78NXnhYaYwpWtcehhGPzym+aGB/mlZbr
UaMlzR8XQcCYLrhkou3+6NFaCdeA8HO4Jnp/RUb+PXnTFrIz/dHpcpJPcHBv71UF
mP7/AiggEeNRChz+kTL7J7uzdtdY+yC4x6mdoE9qd0Wr3VEQuEjSoljAM6sZ5Yla
qU7ESbTzBoXS6xP/XU2HryolUcPtAHJFUw3/3STd7Dgt6UsKzOG0oE0eyIqaJjxH
kCkhgOZyLl6ZFDxvbZUNuvea9A48HF6YMEgggBqfX8CWuC+MYC5x5CKW4s++XhEI
CtkjI8IdWekRI2TkpkKhzFSMRiWpVkOydYrJClDcE7aok2ViD+Rtas64qoe9/7As
XKudztHmqAvWqMh3i6/eGm0utqiYbDATQSrDJ3FLbhK3GH1ssn5d43LDsXDmv+zA
pChhdTTgIZLspU6HtzoiogfKICYdy8EgbjJgYWznO0hFkwQz2sR5PCrrfXVfAcAZ
6ojj4drzsBQmxK0x18jdK23ZVDSEN66+7ViC1JyVyCRlNHTPr0wyQVMXym7R/K1J
be/6CshQxDjRJKc4FgVOaopP+RGKg8EILnxgba94AfmbbRheVJvcYAs7AxiPebBL
0AhZEZbEi5esGXlLSOdKDCi1Iau8MffA1fZD5U8uEgacwVOFOcYkgrWm8ZNj7vzQ
FFh6hInAsPjG8AcRJ/CHrVXI5oHgFgFzmeDg0RIXz4yCpZyn1ppMK6J61Zr/EPEV
BYIL01xbeRgpegFhWPOX+in1odwQiCP5NBSD19onp+PSSms56wZrhvxyMbvOjNgz
/74WZNeqAyWIqmrXgbMgrKyrCuqA6/7s8ZjM1o25PSF76SYao2aJhTveYyfi933K
QkK75Tx5Cth/OmKepLmICO6X07SVvdHKtnnSkARK0qQdOMlijYMbts2ggJzFIIKP
YqXWwwR5mu0b/ba70TTDdwfeV+bY9k9LunCbKVquKDohXZ/eCorIKCiDDQZGaodU
9Galf9xAsOp16y6DkYMiUtx5JILCn/TYWgPw6/ljbthh6wB9cZUPw0qjkATHqq/C
f8XiAQh84SGEbKJFXyxghLZie3hzbrNB/OWPl0Kn+T4wO/7k7xJxzqrFHNiZQGAU
K1Cq2f1RsriTZwqotz9dWuqRZbP+WkRs5Jvq51h8ztQayzeD+dgRy+5pqHW6MT/I
SKZJXRrtCpcqTOlrG9EerEzgB6ctQoSVP6nZSLYPgbpwJHFNrCzbADIG+NYPdaSd
my6G4EkElNB9G9r97vlLPZcbdTrl+nZs+qKT81dZJ1or4NeF0tE7n7V0EBo2fSCB
Sm0zCtoyHFxRje1iLOjUggxlgWVPINZE7ZjhBiSMd2IDmReJwBMg0BbXiWac6KOg
yrnWTRlailiTXytn1hBZxAcoNW2cPoF3s9ekLArCd0DCVwo0Odb0qdVXKBekZ/l8
3NSvFxfqUWlDU5QKK+8FIJNMW9f/kFmd5PIPlGJ31XlQTMs1h/YBZ2h/WJmj5/AD
6dWHjeRxT/4iLaZklIt5wA3Vr9caZeHsCZ3Fpmwr52lrGz+HctkLzKL1omXZzjKo
gk04eXM2RiKV9nBkzF7ahrceh7YYgCCrVnvHs3PWN6mgUi/Dys8jqoaVymVhpjd6
051UddBFO6eeZmowi+Eb2/LQ/D3hduzMWu8BPcbf2nd89u54kqi1zhFsMImynAcu
1EOAtU7zlgZWIlkL8nPWF/gZRyW2z6bu6cf7nshvocT6o4mTZuSN1oulZrTb699b
sFp9bLQpyJHPBD6K7wtccL/UQImfhn0qabFbLUaHTUdAW7f3ju3tGCa8FTarv8R2
CpgzxAy27a0NqxSW1BgV75uRxArJJp1X3MODD6ytaCd7s81p2fBlIXjEN5GmNImr
8OWXPOO93L4/5KzXN+aCRhPSU6MnDai2N6cuEfh1WTx/lBf7s2d/ZG9nY/nUcMLB
02lS7cn4b0RpleUA8srVYHynQJNpHDUp6T92opWrHjbpHJXl2q3e2bUHB+pdrIMk
xO1EnDUD2mDj8P5XoLBfhB5XL4Ws7PgSx6GQvqypnhMhaBmwuvQTtUPvUvrlTaBd
wvpCPtrHeXXooyQC3VH2fosm1H9rdQN3nMz95OI9L002BiudeBsooOwIx/mRC3UB
cDak+WDgVlxONTQhhAhVd3kCRNF4+5ajoM16bXEYIXBHi8RRyW7X4GPoqAvDSuWh
`protect END_PROTECTED
