`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/Gssl7XEWcNt5BxFOhJR+55Sa6fs/+ZCcTIMxDXh+4P1Ne4zl0tkPcxXKC2NkU/
K1+9fVWSkTW3aP9p6vfJ1j/T+g44XKWxc34zAYjga9eDOlQa08M3oo1vpqzBbqZy
xXF0CAeVZcqZR/Ui7RGXMgno8mTmwY2w178vUTN38y2u2z8xwZJVoiuhYATWcySk
Wo0gnjRaBtNe5B5RnnOXVKilrhlUq/p63D73M0TqLGRHLYZNObP2m5vk375k28p5
/SUcRLwVp9wfbMmM97jjQKYcDUIAFpntb13F0gKLtiRKLYs1guC5UiWHn8lhG4A6
quG1ymv9aEwW8MHPcEwJ+WzNsM/RMMIBbqZuuOztw57Bdl8bUVSs7my5rVmk1suI
cQtE2rN6oFAdoMR2VkAtVpsPQJyp+CEOt8HF58uSsCCXrZjjuoWret0hcehNkUGs
pA1QM6ZJzasgRFZELFNAT3xjU5YecdqGY13t4LeQW10=
`protect END_PROTECTED
