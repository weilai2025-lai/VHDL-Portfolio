`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jk6JIAwEXcVJnMoawDeZHhPGskUftSrt6GRdU1seB45y9kmNNLkgJ5bJWzh0J9/n
5SPyBTBzh7XLF5yvNVVqeq1Ba2d7w7eAk5XFpxGjn9pyau3uZqwX4rZeks05z5kX
cDomgpzNAtXejJhuZHxkeqw0Ia9jnjLeKTCxR1A3C4k6vh9XTlgJLhHooi+4R6Em
7xNjgHUEoHVddlz6Yj02w3JghnsDNYcOYMeKoqgOyB39pDDYDXiaMNDRDbJgss4v
zHVk5IpzNIqmGw4OCy5VdOYfHi/1qqJPupUWq64vqvgJZnoDL0oQ61o14mdtuyM6
dNMxY47hjmYodj4flniaONU/ySROoZeUtHnZ/oK0143f0cbWJeIDyc2YDW0hFO1z
mV3v2C13cJexnLFS1VJ6dfE892S6Aw48qcQoj4jZZGkeTbRiKVX6TpninYOoBXdu
IJJoqd5PcaYyygfPVGIbKPaUv8Kq9eG388RfPmA+ZSHzddTuOtKon/WYRkKrBo4A
ddfy9UpY4E4gBHtTi5Z6vuSWqkMGILL0kdb6GZoE9fI/xuG3IoztVNHFsXMyCBqc
JgbMyR15yjdFuc9MTrYy5pcRGLcwGIl/xNEucYQP0TCletxSO/4nsNljchfL/Cqp
99c2/fAlBIntdN2czYCUo9jtI7Tj25MwVhUQJornBaedw07orofQ5+KfjhjNAoVa
mSh0Swvc/CyQx7SXyB2kL+FJYRnYvwqlcH0T0g7PMRuEHGsk3+d0dJD5liOx88p0
Pzr6/OQ1ZFbS9Tih10lofF6h6vjNKRZXhBgXIr7fePwP7zYc8lciMxQWp75uqJGK
Y0K6XOjs6+/GdJBsTbCkLv63LKSwIOXIVXnQYBv3zCwM6laDHTp48t1PerzHHTwj
S5henrHiRavXGXTVLt2rkymTW/nZJikS9G9LaAhPBpNM1SMen4LHTON6yMiWeypJ
`protect END_PROTECTED
