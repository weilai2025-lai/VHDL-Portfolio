`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCz+YkQg4hT01SnhFj0L6EEnX6SKIcXLwC2hgT4Tjw46uebJMyvf9wtwvy2MYHWR
VO9E+70sgnzxEw5Ack9JCwDWke2j7gho0acBwuvOUD2xJHJhOL7YvWMZYQRsEjjE
JhhEXNeRX8b+/qSbR06k4dfve33I1wGEqFN0LtrJAlIQoeE9MAENNcztNoIcgevE
GdkM7mf9H8xlAS3FYcLJlkjHS43pqXCJlMQ2xPKvqJk+UZPWdMIj/lI07Z6jAnRh
anm/UBuo/Slbz5APVEozaya71EsMvh3YX4hUhkHatDXivpLPs0P2wctUfbdG4JZo
Z01rxzkkOrVjKTnZKEAikMpzLC3elaztM2ioF/hRmTZeONY5foM4tSNn25S/GLJj
/E2J1+JDGytFenjUUpZ14vgd4KhhK/MNCv/Jyqen3Zv4p+8enHOeNViWgYtoM5xC
Y2YmYfvgUGBnQSufCEar8uVfJFrfoRWCyoYypfQ9Tn4HKQfekNf2inc3EOvcO7Q5
w+fChRYiNnp7WSjH+9f0IRrVNpTwY3zlwEiZI+W/It+5KWfya8yLYmEnYJ8RcvCK
0vj5TDPDtqsQWAZ3wxPx/RPWd96qDSpRnF0+tkWS9CgrBgxZJbWtlUI4C/W7r3Z4
z0badUTMfcoA1Ol111keKq7PytvlNP2XjHJ1HRekbWpz3QOnJthMbbLIZVfodTln
`protect END_PROTECTED
