`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jy7qGg/F7+iA7qInbMkypGzIgWVqoB+P4sf1xaKUPpB8pJr55mRDDRPmOVrmmCOK
z2W8bf8ex+MSZ96pC+kDq3MHkX8FH90PMC+GxRMwDH+LXTGRrb53VvT2z6lM5CJG
lXEdyk8J6uf7GAQKBx//YW2/dYgqomkvd3OOWAUhVKkcmLllMHyNNlBFpKVCfvS/
7pKy6Ms2BEPhc5gxFRjvU02+4uQ9zeIJ+Jafhd4buogZDy0OFQw+RdaQsIhSm3g/
8JZk3jdh85qvtRA1ZNuXDfbfJ6sKz76hee6trFTbLaJbvFMv22wkc7DkgrOjMlr5
Myja1Hy4wFap+XBccQ6PJlQYvB8NtRcn3mOFeOcFdUVbL5KwtkPoW+Q/VFvhxin2
EzM0PKzlIa7xYeePdEsSAghO41DAGp3wxrS9l9HWjyzNv6EQ8IpPUmbiyT5rlug7
gBVmEORKe/6ivYY7rW3ecNUjoAvDLz9GwZO3QveyYTm93DW0/BBuWLj5t/WE7klI
3P+7YcLkKtv9enrPnH9TZUz1dwmNXEoQwxAhQPuRGIURdcV99fOPAaa8NEG+0BoU
U3wxVdDsdElT/sWqH5ZkzuRLlxWYN5+hlhKB5TijhAPcxW5J0bJqL0XJXG4Wxnpp
m1Rpsz8r/U+wHGuYnHYmJOmTcopQ8hgsZxDwNyQxBZrSXizxNrN5ktU7Zh81/2K8
89o81YYqLCt+JhFxEdsi/PAMopyW9cDkgi0zyteVAHCpfAzacHECD/PynRIFFecl
B09KepkJfmEEm0vBvsoohJpg78+5GbFlsgp0ky6AkVOOWJdcUQFqrk71F4Fi5vCc
KEdNgmu5IRkWJGJJTTMqB7VCzj6OoCaJ3GtJzANqjqb2F1yyeRkFZ0qgYwL90UR2
g8j2C9aWk9G95ew/kjPYgBm3+MKr3jzQRRsCwiqs2kL/spymGT1lVGfKiYxx01Ui
vw7SgX1OaLvKweiIyebdnwbkmIcuDQbKwqWmekbPKw4ZK8Fg372ii/tTuXeVKuZj
+mtvWcT/9t6StXOVsAAdGqQu1tCl8LCXS0pDyJvIHrRVF61KQmYS/RHu2dtRxMSa
mbwiDHbL0FhJJv9d+oI4ZS8Mjnk0We5spi/yKHlB+eiaw9N640ndggUXpzNvMwD5
9+9PMiTTMo5exPGazV/nBqjUiMuK5DMBkKEn9ualFlFv608vFuM9rLZXT0JWAVzp
RA4isoSEiUHutLKnUwip3vqBV6t8j7HTSYXMBCX2hxChrqFWi5Ta6bJlaj/9AuIH
XNATllfxjbn9s3y/baQSNYl8C/1OoENt0IzaDEQDICNTSVFU/EKLoiuThrPrmDxg
afLGdle6eyMhtXi+3ICJWhAKK8bBna045NCkUK9sKQbXhSSYgGvCfEeXepYJPYCB
Ei9cWKTx4IeyEB2ZYgvjWKW+FMfHyrD+7GccpsNaqqP1xhuzF0ob5Dgsl1+MiPhf
Q7GAp45Fp66sd7UW6ObtwJxomcxchYrtX4Dt7enkuc0bBbGknJmVNDnH121CoEJD
XNKRWD1+drZVTR7h9IxSMGFPwCrxBf39kak5j87jNoCItkdjNJiRuTWyqPdqtweT
8MDCOr9LMDbcJervhX8xFHZSGrOBtg0ZZX7m1/gq+64IVe8vrgjkaujL++sK3fSI
uHg2s+N07HVLrCInOR/LBhLyMwES0rhOBhMPseO+t95QbZq7o14qWycLMjmHyW/P
7c8vmEuCq5dJQ4eC/JaSbkgftK4OYyC0AWaRVekWaZB6tuzUjN0eJ6Pfptap9HEh
aOj+dVT5X1SeYvgLv2PPemyj9cNO3REekaNzeBxyGi9q/W3hitVrVgfQm2F1qzVP
zgLrmajmcJuj0dgWrVwC2Ni2yxXsSKX1emJjD+79FE6wSJB3pvABmYv0ElJH526C
aQFm/jhmj93A5O8SFu1ODvVl+5ysihxR6VAgU6OeZrhRWQW/Ll2E/UbCi44ToK1W
YuqoK3yCY74Q0EGyt864s/qFRclkT+NZcoqqJ+JVDRD1WDl6WXbPES/9OeZflf9Y
VjiC7QamDilteZxllYCnLix0RRav5ztGiNEcd5nx0G4/lR5yMWlFbd/CXbaNZXMD
KzLbz32uXSCEkKeLJ5MOH2CIlPh+4G7KXvSbyQq+wr4kr7d6CT+xY/hdxSUGGOqt
3ekFiMOW30can6K9gr+Fbr60eHqPgNODA7jH4fA3C7j0dUdZEEbII3lVVumos48G
7TzaIjFFK5oqwKhlum3HZ2+ooHd0IZZLL5J/vabivAPLnR15CfFXXa+VlC7VwLNd
XjbtcaE6Y8RoWfglPuMV4HF3wwIpERYkdfRwUi6exOxR73TzEBTBhlFG4mcWm/8g
2oAGrOPuGyKvcz6OWefNB81CHTLYH2dn5IT1Ohnx6oxD8nupJaOCCDnxwh+tmg0H
gEX0GcDhwhN859p4eR66wKDIaWH7qlzycxR8OoQeYm5igYgn7uCFLhY1U6rWDptH
Jedplm/vbywwM0eZIFHLA8cERPPSxSwF4RgLo7aoMeMCSb4KVZaJva5wjB2Bhce0
gCS0u7j31siOX/6MkSbL45gLKoaS+NbTQr9ucyQ5TEO1H3hzGbXNjdm6GWPUILTZ
YDCTVm7lMlQnNph9t0tZBzyBaUjL/Ncs8zbhX+LdZ2+45m78lRyf6X6N7+xN0tuZ
t3fJzngkm553xVgakC04ZWlF50AQpzvscAJaG+/2zIRDAQEijf3f1mMv7emfvLcX
iKX1KE0UjfImpXFXWMKQ4sd02vAQRDNfOKLBSIL6ZggG4MczYe5dk2Y2+8YTVHdE
RnP0t7oLs16WKXA+9Di1B84hHjLBRlinD3u0pYZJMhRS06vow499LxbIbi1I6eOd
1wCNInDXQfKrJzWDauhUpclGuvBgx0XGT7tUddmpK40NL7AA/NwNO5Bs8D668TA8
3ThFzdtjpYVd1vhPFkhJ0vbjzkY15fs0/R7Ihz7G3D48ezLilrRlcqgSioZyzYXC
fcCvC+oO6Ptpt+vJZNmNhjrTAr5LFVuxEMi3WADPVLy8wKDr7ssa7cgp5B3W6ha6
4mdnR6Tl7J03WuCfAYizREbXEV3VtlKs4zTVqz3NN/bH08D/vWbOTnEIEeUaN5yg
Uqq8I6/WvvL76HTKbyjpHSuzLkWxVyS+YFr7HJmB/UBhvkeJm/ufyI4ipjQWWkY0
cUnePy8g+7r2rxggi7QPx9UcQuTH9iBDfNOJGTrGpZT0Tpo3p7IRkAUJmiHILg9o
qZMCaYUmtkV6gJQ7uISuUlwSinbyM0MZ4pqppaZmLO96j8tcic0sulbgaoERtvSh
hj7Nf/Ct6QndGE1nFJq7kzQaYkRKW2BQvDkEmRY2JagDe/gP1b7vAceMnSq2Hfxw
j93KPRcSeNdFAHELgOVRbloiAqap5q3BcTHWlDMrgwfGEhRoQvtn1f6x2CRcfaEj
quKRXbLvJ33Xo3HLZnWx82jLdI7QKJcZqGDtkIfCdOnt9przHO6kKU0bSXaK6P/u
74VlFNinUpz3WrGxAh+khy3Y0u9WK3eWOz/fGD1G0/tZAAcrTme8tIXmFOGIId8B
twYku8PS+mTuzTXFqOAvbKrmA+1wMkjdizLj9Js74ynyPjBbiH4duUg6F8wLUl3S
3RIDcCL943osidcysBStO73f2WsHA+++cxlZn5IJY2AXkHybHOk0Y0Xk3L9rfvDt
l71sJdUqleGAHVV/qVgHBaEY6HFR2YW5S7ZZ6yP6qAFfzDwWEDI4FX4fAQv/dHSy
KJKpbOgql+ftQWa+jg+QYP08NTakEAGp5EI7mK9s8pOfLyivPlO/VP427imnfyIc
krFTlHpfL94wnqKihiU1bg/Bg+R6EV8MIt1gccV1mz1EJVfJw5tQfyQKtfI07cnC
pDBMeoiiRi36qxMYFNtuE3aOwK+ll7bHYgDZ937YT/ZYRu8y9u+LhafcMWcsxJnB
YnZ67IkyelJagJ3+iuiD1J7l8LIeUe+AtW7lVK6lBL5lxVtqEfdxaVHhlaGFz0re
lFdf7v0vv4jtIVrss03dZNpyI+dLHbG8h1tfjqeTIO3S9RFECgdQZ9pRiJU1tOn1
BfRsP+lIz2sNk0ncYEEikk8/NTojfIFj8zssEqDWh8q0yiZO/RFpoC0QNMVh5PhT
y7XztZkQJWZTeUs/I7JFPt4euccVkLB6aOGbDNsCCVAkn6vGO91tNPqPL5eWrd+1
FSV4+VYNeFp5/VEhODYBXN8ydzWuM6HxK2up8HZZIIxNda8+rJ6SyguDSvMLsGqe
7VBKTuUJOa196xVMwlMYx8ZAhlotI8J4giahzJjPfKB7ClNFBqxj40znnFTeWxSY
EKQ1nyZnoydjESgV01i9RDoTurmSGKsCk0Wt2eTZ2yUgV76kLo7nFP+CuLqwpq/X
VAfUPHP0kkoB+c7ticLZZZBXt7F4BqRoFT0F2s5g5DDN5J5bFI50Vd2PXLBbjlFs
14uLLZdAaSO7ii5EQHd5hP1N+XkBUt+tr69FbiAqW7tE4I2tOyo3Pu1L7RVIcJum
/bBuO9yR2RTaaEpMvdZDQ+qiTzJ6uHiiK/8PyJnpqWRGozyW+b91TYqViq9HcG4C
0FRieAOqATkiUhgfe6FaMsVeCstlAfMeviePNMHsXpcQYpt/YleKnUglmK2Uy7BK
yF5JdYYw6Ug5G+VYuvWU7XWBc0rmAmpULE4N8fm3pn+ds2bpFA4bK7/8dfWcGsUv
6Mk53iw6tFad7fre8TtOTNzGDhGHdiMZQMqLBy6wzt6KGk3PkuiDvoWeWzlXh3Nz
QRH4Q5VEo3PHWwq1/FQvhAMyNVlbIcmiyEPJ5BKjmEC1cM9++54GL5C5sXv4359g
8n+iV6MzCNz4mqUusTs0mMqMfWJfMPeYRoBivH5ojQhQ2siG6xJYRTn5wZFE7IRF
SxnuPGNDQF49SGYjfBDOAVls9RU78mC71Apy5gzx4cvPI0rf3lIMt4m5d+isY43A
nl2CVjgdgKPsPSgDchbdMTWYQ/a27TgVxK8dT6bNfFIDOvUUlihpWE9NauNPvLeD
j29+vje2xHpNRHCvEvSi3hU6Ebk2XVZ6ccclYLIdDIiseGn8wiQet4fwl7r18Ine
R+kjgE+wzg5bhpVNfqQ9De04cO76fIWUR8wxCGKw2M7U680WyQlMScBdCxvmDoHz
xxOrawVXyTQpPuWbFtIj6sgYfNKkDqol3Co2ZPBbPAdg2M/CDvGA/8engzTZT8+B
FKbmLxRPlbY1M5LyR4WXAATTREmQIlyaJ7iiXlZ6+4PW0PunbhlRVM9Qi1uAqv8w
gct+1Hax31kWDlNq3Fj3RbSuOIp34HqTzaq7IigJnz9B7Sz0qBHsElqHfj+M6xIj
sscmESAd5KZ5i7KI64m4MJ1T+qUZkZOYOuSR3FKdveyFeSEtwWSPaEC3tamOqaIE
RTgGc3M9evPWd1/vkas/0BLQmTagXyYyfx9KUWophs2k1/H66H/hVtmpNdla6VT9
DTq5efnuJZPoqA05xzTW9Dlw2YNG5W7ov0f/an2vaa/u7k6OF8hhLdsbZKhK8E/0
Ryls9IH9cZeCiS1ITFFWFVdj95py4UqL9Q+/QeZtsiZBLIC9Xf/R7QRymoLRZQsX
4+qVm3rJYIlnpRdc4+Jy3WlEX0DDCEEKd2nCTxIc+PxE90i4v1udZVpZgcxlfUJI
aGOJTg/+KEHGuT31G4LknOmaJTwLS3izKVfjSYZu9fpN97tthuCOMtWA0bSlR4Sn
Iz0NFS8LO57bgbnIDVUKYVo4kQH8YlkJmRYPyZfXeG3V0dZEZm94efbXJmD4879S
FSJg/fdf5QqMDsFQ3Gjl1OA4QA85tHZfXXXg2pWOASp0pc29zTFMEjr+L052I5PB
uSSj7gz/YMdjNRkW6yXEoCEf93hAQnWp3AM64/Gdg0104EsnQqtvp9d2bREAdHwc
WYI1m3rYAgck4OLk3ICSKbT3DDZS2JthgTM0DNlpsd6Cu0iYo4m7gtPNyTLNyOkN
n68IhFvLhKpliFcr8BfQxm07Ef2eKf5ZS08gdm9s5uPgzJaqoY+6F2toSVsSy/PJ
lbWTLf7tZDIu9jDPaU3NWeueB0InCKQu0q4Wk3J3rjZ0xa/cWWe5iw+DmMA/EChC
J+x2QTRsHxhl2sr7yipJfXPFIM6HfVPQafZZuSeZWVcdAcj6UBPsdEJKy5s+2i3p
UiiMYT3fxXNq8wtHq417aeTcjhiDznZnBFrBNw6q+4HageqKuHzw5KUkS0P+U2jU
g6S0xuXPcASn9vfLqlOYh79H8GjnY9h4pE5gb5sJgbQCGra/rjE5Kg/MnT+9osVd
ZEmMh85F/xkDnC00jRhWIEBk3nsPZUvpJy67JQcxbofR5LrpVLoglIz7xHJQ19gh
Yv8Ca4juut5QTPHOIlUKuwKrPR4j/T8IpW6lS9jB6R9r83tAaFSnKGTtYwIYzmwj
bYUtb/qkgYWmfl3d1bqZG210V9Ube20LePKQdbF7jqYxrcq1oHK9/EwMPJR3WBE+
v5BLAOraC9QKLWfbs9tm8uT8JrAwxuZLVD4Iog3jAKiyYISmvl5z5ZxyxpRe2uGy
udMV9ZIvi+qnIn3Ee7tuaxz/7Nzap65GlIUafyNMVwJ38JEPzpIdsGFd2YX3loms
hc+CpqPMM+Mr25MG1RipiljlLyN25vvzlWqarBFRO48gYDWcjT8yovo0wVTyEgAa
K7niZ+7UDC6qray9IJJYlRkm0Y7UERRogQ1nIm+au8r03PNff1R3MM3IxLILoTfg
LY/ed4PZiZPSlutrq50RYFMjc9/skos54v0GPH3d7FcTcnxJP6OEBV6eQr6NajqJ
oAigGdwxT0ZVoyA7lsPD0Csm3pYORknzmeneAT92Nfg/ytM9kIK1qHQB/Wt4UgWb
NhjznRnNHSC4y7churKFF9kMySwvNQFKXnw4NA6eWbso2bb5V5VpjouwGRCf93Fu
+KJ74QIrJt/ouxR7VuitZYVhcYzs1/6xT13fF+2UJTgLETDwlKVuCmvw09uI9HQX
hWNXybQwFIm51zeXX67Vl2sg4YvOXAFBRoejAJcYUIYdMpIdP8poHKvtpTfk279Q
Iw1IRIsCanJQaHlBmkBS6OZUTkqt252JIHUVq/66PtUE2PzFo/iD/1i/4YQtmwKL
gb2Ku/TxWMrKXC7aTjoGK+ydK78czQXaTsyfLG7mV0uxyShAIttfkKdQGa2an1nX
DLnXzTQcOzgQ5AtWctgzoKTnv/HUZ6cBZV2Z5QUTBqOUoY/EAEoQhO1jaJ2JE1BL
Nur2u4kmBzzvdsnkOMIXuNzpP+WeOex/Zlrd4/TSLjqTd8m4NvYjk9N/BcUtxjJU
WFWqe+z+LbsT459wgjpJ03rFd+AVLK0nIBAkGMimY/638oGdwLy6293aiiMjOp/r
VuHQws0cerPmEv5xdT3qQGyjKcNaLJcJLbpku93B3dCv3mGQ77MiOF9A4KRvC14S
rN1e1rEybJXEjORoSR33KAcN3+5l6PDmkoJh9Iw0oOMd9HGYLXzmdygAB1bOFYn3
aWSs81ofq3Y+2NtEtbPkE+/eF69cAGs4junpRxN9V6DNGkKrotvME0bW8zChdlR7
MeUzZ7u88vlywZTUOBNn/2G4r5/ZrVx6ODsSCMdVKc3oeOiacTp0lDbEdVqJK9mp
HnUvdiO2bwRXpYPWHIULyEZtwZx80AEo3xPxbE5wYSZ8hIKqzPpYfkQvoNQhxs1/
mXXFOmrIqgwkFOSNh4BKsutW3SyFZrbWv/YlMT0yqWBPJSaKZh3Aeboumy1FHqVi
W6XH6cykkRrUXixASVCcoMNJr/8Wq75OM002ytZuwgEW9OeHplGhIfC9QiKcxGb0
OFoAX7fKGnuLK7S90CFzV9oXaUZJY05EJEMd1XwhNtKGVSw9a9Cq1CsfDg319I83
ErYy6QHEQ9KTGEMeyKJi75M0EpKHTbytZuqTffe/O/xDKkFvhkDyNU0mrwiCpvE7
KzBSOb+BW7O0z+6fqkDtSYzCDxAH4xptyFWPqvDIJg8t95WmYPlFDJx58YCoOZr6
/jpJrLOf9EeKLLaqi4Bmq92WtrLHcNNMe48QDYZA/Pin788+w5YdG6cFhxSaunxB
5KSBcBpa2CFoMZJcXWcKpyQbpslfhzIagxTih7JjOGcrigtMnQbCMeFqG0my0NGc
eu8Q+XsUC/21yvQKdBpwK3Y0qZigg0W5ZhQkvnhvfIBEgE33houEq1XOX7OL5InZ
Rn/r8Nqu/K0S+4sHieLIKots2wfEUjTSUrh+GG/BIjx+QBhpgVSvQbRNJGPDURg1
EkkdAvZcMGBYpkvSZLGwLytueb5BOHq+3GgzaFM3PzS1l1d7h2l8qCGQm1NKBzTe
mCLokLlzZLcesoJxQdEUaMbEeJLjAeScyjg3z3Xn1exmuzvhb+2FdsYuRAYMBATh
Dgh3dQsUXZ/R5G8zrNfV2JkAl4Yc/1Bo/5P7L3kMisioOrHKhPC42zbcZBeIlFC4
ob8zW/yUjApgrxA0SPL/7ElfYq9f3tR8Z7SmXt+oEO/TrGZihtibvwAnneZpv9et
qGGBht2/6QOcuTpXhtXCIJTTiXJ02EwITLvZ1NHS/vxIG/t2ZEOnA8WP3Qu8gJSr
KJfyGnoowmjp/8pTMBz7ftHEpfiy+O+bJRAWpq0xGEgOshR431bIaVx9373TP0Ze
bKFI8V+zqZ5Te1c7bc/mA9E3zbfJj5uBLfXTS+TVVG3tn73QI6PEptyxiy/q6AsB
xgnNZzH1nfsh3/0N93bDPwooL5eJXR+iiNn3FA2hX/FVzDbsIaxmH1ZyWTqzKrSb
kfsnB2cPfp0XYGceWk28gvV1ghA2g4xMJ+L+5hhKfdAmW42BO0kY1mtdsq0Gulrx
4jgbtebnw0Rsk4s4LCWFvyOe+QrGq7W0X2KnjQGYiQstMtfHoX3C6BvsrxD6V5mw
psBQpRGllwGdyBPGJ7iUcMsgaChZqzHwoHl1eLBRdYZx3/z54vvIexJCXPLLpVfx
z1allwfSuRFwEMmo4vCQmFMDcubQ24f0VEuntEPo30JFRoSF54T4HOmIpFNqLCV4
+D5ugu7YdB6u6lKsaeohpXpbV/ZsHBA1NpvaqwMmLEF8gjXG0aDhMjOV2j/wTQxt
AAkam2ADACeW0x0ESNUFi3NGlFTK4DXzPsYKV4romWnmZQCodRFzjqZ3V0QIAinX
uOT88ams8JrsWf85OI0b2cEF3D1qnA4mKtRMAOmjyM/c//r94Xmxgu8q2uTnauRb
VUcPsX2Q1m5VVWZPtI7lYwz8VKqILUOuZ0oVLm5T4PvSDmh/EvtKT0x58s9Te0xE
7T0spien78NQJ72swSCVuDgb6EZ+kCfvWnRlpwRAmEu2qgSskC/ifeiF//8sW8Lq
6z1oGbsrL6EdSl1J3p+g8+zoH1Z5MPCRX0LlK92cTZUDrCOqi846VzuHqypqjOfm
c/+5p9X2Uh5Xzz66jUkF6KXgS8DKyyjaIEWNotRDjKvxeIkdAATjg/5lJudsgsp7
16zV/qEczDw4e3Jvv8buLWPbAopPI5+GCDef+J9YvSj6QnF06TBfr8e3adWgcqHq
0vJlccTMPdGJICTsdKUPILyahCq//mNK4XVWwXVbGCwv7R+YRCsJI2pXQ9SisoHl
FmWins1FIHy9cVNgb4W/05TesiLlt3zprmER5dbV17KevPebWjEo+GS4CVW2DXNO
buNqQk3YBDwsQ1skooMdPSmctjiZpRiXA7fT5ZgfxQLWW7k96bgxJcdhl7ilxnGc
3+YF3PUo7vX7SJFmwvtWWUX98k+r9Llw4z8DDlCnGW1WVPgzxxciC46jzJ5NmzTz
FOmkCcDvUab45PXy51VhXP/ppEIS4yjKUcVFoT7rN5I9Rt48LSFQTxIAVLoxprVs
nmZlzOWH9+xZtkdFi2HDuIREluB7tVBQl4np0kFp/QNRp6SUgjkjoz4AQkG13PcN
JrxO1zU1UfP5bp0PryRzQt1pfypF3in/vvjRqjyV3D92vagXq6EPN9TkYld9kpqu
LHYFjEsKq3cxXOBp/p7AQQQwPK3VLxrX6O/s2s1jieh5GvI8zvjOmiK/E5edi4Jv
8qtduo4d5wuKJdlEuv/x753joa9aT1tptEMN6oLXBavnb6CW6Vq4YcEOB9aPg8a5
rNx9BEwDczba9utKD/OSx6z8VgZq4tmt+Tt2gVdiJFZx3SFpPcTgV6qHgwrvxBaU
VzpnEWUwqWf4B4U6yvB7eYMbJk+l3WVBXH4fYTnNtnjNGa5HoRkQRCU+o3hAj8od
smioMjEuZKFhSgjcZxKF8JjEWudOsig6HN5SEyeP8TGzYNdMWFgDPd4D5XulYoeJ
4mQkhRCYsxeM5tltonoREeyIcznT/9/fKizoFs3BXfe/s/o9fU6XtT9QbmxcX7dE
zQCiTwpbNma5QFnJPKVrVxzzmsH+eyKAEAp8cxbN2J1z3JaWooEEKOMvULKjsJFC
Z9oqmvDPZq+pLMPfZxathxdRu54srqcnvH4Knj7R8ju2QW+Lgfr8eXXdeGgUkFMk
TSUUe3JLxgkAC0cNzWHjDdhJ4ByLwZyx0SHcbq0vD9pqurc/k0QIvQyenSz+XBHa
hEY8hzGgodTjZZ0hoDOZDHjIni5MuiTkW33vdfgyhBWx4sBDoq7w24qvxojKjHsg
p8j2fWnhPP+tiPYbemEZFu4GECTPscs7cWp0luNfQ6rs3VjxKI8Jzj5P2+xupxdr
mkuhUtiFJE61xxght9YspP11Jcok14tWoYn3O3Wc7FRAXV4jPj7kQMYuiAY1q+dV
Y3DBTNaop6IavkVxYiTt75dOZ2MOySU9mv+G/iUQSfv9IDgqczx78IpxTFOBGsJS
JKPz1u94EeoD2Bfcwus2O6iC6+0QvNJ/XCPa8wKxOdWzpkb9r8gjVUSAZSrky0f/
ImIpL/PnkAam2faHgfFAPVKBzeUeiliNs0sZ1eQhWas8AT582vkKcz3Ly4f2+mgA
SCPwTltbYn24uyM1I6S1gXNRPjE4GvOymgPM3cJ4lbQ3sKWy6m57Z1Z8IO10u1AH
06oz2wEgg/dc4shm9PdkvjKTlQ+u/d1IKVMveWcUnwsnxs9hvKb4QZiTNgCCIX/D
0AHGMiiTOj6ZY9Z2AmJao9oRzBVtVgzUOZXEGngNihPD6MWApPHQ0zCRdMeJJcN9
cBOujcm5NoDQ2fGrmKeLI+O3yYIhQJOFdJYUlozoB16ijD939Qsb7GeguGOa+zU0
gRY+7IGRSrwCKYN9UTonctoop0/gmP9sO6WzPF5Dy7sv3HvCiZOPkDUEeQaw8z8L
cFDGuewapyIMqGI9D0RtiVPz9XDNhSTeqgVJ1lhhcvo/amILUaCi0mVrivoJi4Id
H8dCCHQl0TK+QWBmskYxfxccgSB4Exdx/oeEVzKaH+6A9jXUPYdgY6hXjxiNONui
VvmwbBd1SU0/AuDm66Tn4/ryei4qw0x62jiyg1V0JU0zQNtatc5+wKI7KwKXK0Wk
bedtw67maCpKdpODfXOtiwxoJr/tQrwO1x6zXErENxkckXbPd+4YgAADV7Z/m1Lt
rZO+qh3+bDuzDa9iS+/KmsUtZ9rSmxImH7SqzBXxXN/t6upLgNwLFIwgwC5A4U1x
JIcJp4qyLK3JQ8oif0zqG9ztSz4zDafkiwmV+IwLyGq3cPk/8+uDXoR6gxzPP7W0
Jy20Hid6Qy0BRxVGvGGULz3oFT8zQxKNgQIdsAImAd3RBOnZLoQOn064hHnbAabG
E29jGq/ouHEarvQyM9IV75i0PpFOe+wkpHelNnsN6yrR2+HZdgK+F0GabPENLTbU
M/nzJq0UNlA6//5sxN5Cg6l13jjncprVx0mO8yNzUXIolXZC6CmhXhKDvuVum4K8
qcDzYqNnd5HG+rsEVrfWj8V11KkF4E8VPVD26g98X7QCNaYvz+BztvHjKnXiBvyq
teZ6BdEWwtkkpIR2528gsgar9YjBQHbE7FLMs/FrlWBVMNKzDcsQQHY/MxUhplfl
IgDvJOfBnTWY/2p9VY/pvCm+yFs/hnMueTPqb5DhzS5iQAw+uVH3ylVPyGsxN4v9
gATtU0vZ0ZgqafD4XFk86oK7tfrHYk8+65Pqas4JiQp/by+GMq+UA9m2RFS+Ianr
+QhSXLpgOsDvGCUdRXwtrrT26ySZpM5LO7D1siRdo9jr/i0G1yqnc+Qgd6IZMOFo
CLI38uaV6jUnXzP+Ia6Nkh3o2XhMZpECJyFmA8wIOeKjYCMuIs98xOoeM0oOZ5CF
igcMWRxdIaWtX1qJniFtrcJgumG938O+2SOnPnuLASoFHN6tg7bcIZXqL3Bbs5Yp
Sisjw/8+lPWfRriBpFhGGNRHIRSa38CiocSF3P10Ic/rdelXs8noWr4QF+ZcxfEo
u/U53vKMX1Hre6wGiH5Yqnf2Rx9DomKswC7BALAXTzLfk7ihd3gdq424wLRdbezO
1FZNTaKMouDM5PKL644PRRmKdCEtL9u99jeFK7qfBwQroD1+a1HfTc5mAPLmSolK
iLrCjIl2fjf4pXS/GYp64vUjGsGCbk2ZrSvRLPQDE6fznj/fxzurykOdMOSd1Zu0
qPRfM6TI8vBT+W/WxZCVpUZO8ssncGB4l5tGDn4MkPdW+VBU+LqymesqjxlvyUTs
vN0Qa7te3jEF9NpPuy52IwZaspzPM8rRcXtVsVks9/mjEJv/gHkwLlt23hFVulQ4
Rj6yoysQJsPi1uL0sszhfaj5vByg5KTK+hATQfg5/VOP5dAAowpqsKYy1vbECA/w
bKi1MQjY1UR398H1NXuC5cbjYr4x8Ml6fQxZOT86AOMNnabv9Vd0HhVsUbu0q/TI
/Iqrf8Go2KjOOeffPNXY693/24qjIXEvOnvI52xKDXci1Vt9TT4ntUEjtMloGzeI
8jwpepjeglaFfE2d9Z88DfoQIFSsHSnsdqGHrYoM0YvodIWy+7dHnFhxFHLctwgZ
nNk09oCRz8EgSS2j4TZNK/8iTdoH+R1uveVSa2m9yU+o8f0CByiUR7j7DVpwCD4V
9yooKM+R6ONhqPTorbWPYL7ujUZi/t72XPK5Jhw8rmc9kF4Et6AMi7qg77ddOeD4
eRLjtydLWCvqg1a9BXJjik6v356E+UWGevxzamTYAK9UEwL3GWCYilnOUNA2qr79
q4LvNn6dgYJBlrJ3Ux/J8ifg3bhAXDKIYz49o2oFeZ5Q3k0Ta9mOa0gujnMe2xMj
oLTsCst93PWfN4Z4pVBiC4SzZ4MxSx8J+8FbErS9cH9qh4xoBphrvc5SjhSHGDSj
yuBpNGL/NVxWqOKVCZ0wGV+Z3nR3CURqW1z3dHAi7PGYP1emtZc8f+r55441irLW
ueOUatZBRZ4eMWOVwj8yqdDMo1T98b0cTTbhvbWrGH+s/KdRKqQoR7vI4jcl80YV
zQxb5HVTlBH4ByogPGPdJ949m2T7Bhr+kV0TKVXmpkk6OOcIUUTjX2OwKrZ6F5Zw
m/P3+P4/fkuev/bfEk/R9cOjqPRMx9q6rJuXKsOTroGpQM2ccC6V0P4bX6OxpG3V
y9fdvz3UnkpNzi+1HO7zobUma+By2mOrv2nbN6H23hsBnQTO9uZnVymPKcRHkyPP
Tvl7Ulx4rqBeYsJppWnjsER27MHfaWq5Jc9bGydb5I/TpXpRA9mityP5fIyQkf2C
M+suk88UAEubThtK5FdVT9yhTPDB7ff0HdBZQhlJl7UdTv2kA6EiRfAxxQG3eyEu
mj7QoqbUgS+GgP/M4DllceK7SeP+dasfX156NtNcd7X8lP1BWMxcQ+pgh1HT5ElV
4DkeE62samfCji+KT3LUcmig/Q3RFCrCUxG+V6V3mX5wTj52o94mbRu+spfi7zqO
E6HMopjIOUNSw4bivQsvXGTxgIAXqT+9VUx21TmvvgeAPusFj951E+TtHi4408TW
Io/Z8T5q54ZQguevRnIswmNodNNRvnD6onE4vvzIXoNkWikVd3pXbGkejiQcDFSE
JIcpdv9pNhMjGl0MfFr+iEv/M0JMXlmtHwbkE/uIJg1u/YVm7lwhMAv+gHHvHGjZ
EUymP7YN8AIEPgPwLKPEmCfcPjrJnJu0OqwVfQmK10UIzM61/Cbf7I20EfodtJm+
RxO+nN+ZHYdUDW7e2PxEQCzDVOzUTok3I+efwNidvjyWEInZovaBeZ7AMO19babo
Swrh9CZ/k0NJ8nnPRUEwOt+/em9peEPMbuB1yYAF8NMTMKSvDAz+3IxSSfHSjniD
mYnaxl34uGp/O87niqrytJhdx1KXX8On84j3H04Xbgf+B0fvTNnoLr/Ja9tpyhPA
yvGU6rYhuwSL5DZ/ZIJ1BD+FI9BnlFQsgoeO8mrH0h2Lnf4D9lhx9eguzVzqE62v
Okfe9yxxwhdrKvfjdq/Glg8oY3pdSU+sGXYvYgoGz3LJimYYbCqmf1+oBPv8oGT2
ukBwTZOI3ElbDCp41ioXlRwaVY0J6RJt7qtIxqmSgK/hwhGizO9BSljcnF+lLUAH
wjSE9HegI3YRTpX52FynA/r/PnBKzztSF80DpO8doWY6J0BGMDta5fkPSe6NReHN
hj7jw6iP/558sShNSZweYvzhdIXBiP6SHQ3lg6veeHAwELSw8Jft+pe+JM/gUHBJ
fJPLQFFyw/pcOiaW5LRBqcO9Oi8bCijPRxW4XO4QOq02wG2aTHU0cltQ19069dFw
7HUJbBLm/fKYPReuLAOWb48nhAUcOijuiDTmtFfomTxb+WtLVTczVicXWi2OdCHt
PuVro/xofqs696JkhJLTK+1bAHTvm5QpN02xZ3eKhqDXUP656NJCLiZ+SHrIVQiq
3dBYvpz8VeCJgCHs8udN7Pp0P0hb8r9oZIV9QA6v+/MGPAkqJugbEUlKo0oHMtL4
0PcdpTNJlQyB/7rIaYBCs5OqUYEmVh8wTL7HLZfTRMZ5HSv7a+dtBTcwuAjlxZg5
qosDwKAbKIrWwPEm9EaT4blQfjrMbBryLviREVqfZFmvK77kA3me0xa6Pm6L1z7C
yGNV6xgNZsGAgxd4fjAnQNLDnES9S0yOvcJDzcq2oaGFeJ3lpoj3LgW4nscHa2fd
HUtA3ADh4puArA42zFwp+j0hM54qJevFZsVh3WNYXVlB+AGFAbExJIA2OQy+jz7c
odiEHNide1U5nLVdJorxPzW5Av/ITaQE1EU6eTU+YGOYgidt8uiSCCT/MX1D1cLI
ObHrwAwWwmBU9tPkE4uIUSP/RYposJA3ij0BQtFgkofgpMZsQgCnS91sJqpNINy/
uRdV12KyqCfiJQap5QNZYIG8CZ3JkOYNuRKQDk8J343wUlI0NMaaGTfwXGAqJbJ6
yGWoMYT1eIZcq/e+atAWUfphSFHF/JjGfaWUMTWapgnabk/R8xaz1ZsuE8MT31YO
Px9DKVE2ikBJwXMf60bxvupgZIoGWOh8EvVgjNTvWKl+WguaFKS+SuPRvtRqSTe4
03+iJP9UcRvA0uHo1ENXSwjj+ao6iJRjLYmrgMIThG5NWNRR9iG/AkY1kzZKpv2n
xW96xMQPQLWUFGVts0EJhsy+OjpPdIMOlMGSWHIIeJpkm5dKuJHKZMcW91T2rpxz
5Ecn3FocEoOXd3kKQsYhcjIjJQrOh489OG31iQdsD8NDyTh49IIPJtGjtN0HzvHq
UwAZKbTx+yJlCB7hx7nvE1+6PVxOrQZVgwuCRT2ph5Yqy6UFBmK21EWPiP1fwpo8
9qfQEtVP1Xr7DmsotCsn5NmPNSnyTpb+X2KB7Hrudi6bsy8JG79oLnniEeafvug2
Aj0pSCNkP3FoKyAhGz4HYRmpyqJJRHcmLtNresq/w0KZPzBSZvxlsKmImHsILjjI
Plp+01O0QZlq9+8GX2JzewbY/C/2Qjdel0aoq+LdkPUCh/WG04UleOs1NU/wr3bU
yB2+CusTiarMXD15lL8AdDfpvtpcW6Y54VKpYIDI+JAesAHRQhqpKdwTHXuLA2WE
nll4o2JG1J6/SzjNq4S9gphfS9fIaIwXsgg37SXRTyLWU4zedxDlgJKbQOML+sZW
0dsqnHjwk++Lfe8Krk1klt6XLaNpJBWevKq/oGbVPwSX7q0FVI93i4wENtVSG86S
QczTJ2mfI1k27sanbo56s3KJBh6vOwvYCQ3fsgYq4a6iIY80ZQ0qcEWUkuOC2Rhq
E2bCGweN+wN2GPhlEcoQiJmyrlYnaQ2fi6ofKOZQdQsWUFAbQl3/No4sIh4AYEaK
kKdGdth9vLn4Lsm6IxMBIMrw9wNII4Dv65YZeMlHvMDIQCK1AGll43O5rVIO5gTm
Wpng0slATeurh6+K0SEfFHOvrrJIab1FW6kIyJKSPHaiL8k8oKP2ACZPs/eI1VsT
7xAzooV+L6AL6LFxT6nOYNQXdmCOTZkkPjVG4guZJ9ESOy51+16kxefaULKHhw2R
r62TAUWtcEb5gHR9XLVYBQvWg9xX0+97J/3/IPmcw7q+lFaSIX4gwuNGDofbsUQX
wPGtQ8g3JjwXEV04Za1a8z07JMCteP1D54NK0qpAo9AD0nh4cu31eXJv+RxGQqzd
Fg3F+0eBoquAA8qNP9SNyzRjqcHYeJQwQNOjTOMepvNwdomNNDNBQvEIrt2iTJ8X
aC+SYzgm/r+a/YEycc7nSDdMLx1YMlHTeteneTTfZ67298te+K3SUlEiDc3KY1pE
C6oTf8nPubzXgqDUD2cDCj74pcNb7SAi8LhQ2TyEq3/slLLpuPJyRCOVemWFzYwJ
8CLSaI1BErPsNM/zIecOhUW8OSdGYg+fq6Q/UNU7pq6B3NKs4fCv5GzNf42ePrYM
RQWOyHTeTe3s1XjSNN9PLtql/SVVd7RQzWlh3B2htYNw38ygQ8WpFhsyuE+YVvOz
JiSjyeL9WJ6S6tehp8par0ke4S7goiL3wBU2YTAHNgZdyt8dtINbz7cqyqE96Rde
Itul1NKM2B71l/DQtj+ZK2sUumgCF2lnTvwiN3fKrhvz5/jVBdUeRG1JzgNYny3Q
y2oOS97FDLvGL6c05Boe5fYENizFd/IMQqxjAZy5TRRpS9a1r85BJ5jrNHuv2O/u
cdHOCM3nsX7zHFYuUPhmp6xRBpdGbhEWOQUhsPMLGpSMcQu/0FX+Sr9R4/V/+8gJ
0f3S0zabanc0QLO8M+ueO3YiEl1/MwmQGzddylILJHKpEnnGe92G46i8FMoHoFOO
s692zuq366jbJ6vxkHHLywT6leaZgkcB87vzEtuNRx59fm4qpPW2fgKOPpRVKHGr
ZFVFrlRzvyAe8Nk5sruv+zi9zTu7wtIRlbJVsHdEvyboRkSRYwRADw3kL6bV/VKh
UlvzuwbwTMWjJI30Alg4OoxA58Fh0e1crtTJOxoHtSUYKNoyvUBKWKu/z7hWJLjY
LSHubOyfvcIH4uMUmFiwq/UyIhTxf2vlZ6e0DvhEipqwOrG9c2/MyBkF0CZGYptj
NyHuh98w8BHjzFufu6dU8I46SRodYEAtLXk5eitd1mKJkLJIsX+sJ+Qir6c5VDaL
RRbypkDnvd/8Nkx2cyzsrzXja08afE7xzVnbxGcPnp9u4VMPqYswzGIWpq+tRaWW
NzJF7xIutqsBZVF1nqSzXnpdcvCkuVhR+biIEXaMEl0UsB6lFUisFxupOdrml4SO
hvyf724Fw2qsrWvYK9+VkqYritmjtfn2/L9hxQiPKti6E8WNPw/c7ctqwAQ0FF1G
EU4RVM/l6NeCJqWhLw8+C9ECo4a0SuuKSP2+MuITjm5tqdZgR2108ACxl+z1MXrJ
05FtoFXSiFAgX+/EjCtWx6iX7GW5wDDqFOl4mqGzPgXnbRuw0QFwnaZsOJvWhOF2
ejeXCZNeJ9IjusawsukO+gl16iroZVbOdUUf+nq8aUANoKPSoGl7bLGJ2cAEpvNs
iv+769qoxRCkq5h8YYH6gLWWfdr0CpICMSHqBn87SlAlWG1YYdol51PlWcQB0ke6
inQrzS+LOaishjoC3FS+HRj6hjtOWRmzJKSTw1xvDzwHy6ja+92q8USlRiMhKJ+a
PEVrIVcZhV7q/OhCfJ+3+HjCTuS0dEnYjwVAlNcALyP8+y5i9Ba8rT5yNzTVErP0
sCJ62vlLh79DRiXP6rYGt7e94nYfFHcbVBJuF7IJ9Xlw3Mg52cDbsYLbR151OA3P
YSvkEkPCNxMyHWM3+iUriNy2kPCrBZxEGrWrP92abXWUOVgZR94zB6nLmW2ZBJmV
VxtT07dcZGFQ5kmT2TiUEI6pnXYhK6n5JYF17I332AyF297S2qv7zaGYS8v+k7xb
QgUcgE36tb1by37lgONuvYIuJa3SE4Vqz35mrLH1b+vMoRmOLMz1Hi9u2Qg4iQlZ
4LIIX0DoMLnC10LMILyShahlEx0C9WJAg/miOP0oWHE6rggWCXhoKqDgAC1vwpml
f0QCjPqo0myMWPhHZysekYYxQy2RMZgvr2yp3zEoMoDtYqlSx0irEGywdOaS2aLC
HmhQnehtbkQYf7tstBnUamCDmLUEaalNONBXDtKYjJqKR4hMpcuWsKt6pVLBWUJt
aVGLdIce1CZ3VK70J0bZIWoGlfaUFcFJNhq1R1mZDag4oic4xPv/v5DDPHWiWftc
seIEntnVWRzMvoAWUPB8IufUybaQiSpgKI5eZt807ZQD9rqW9OZyurvtOPEx1PrE
NspBjuMl4Rh/l/iK4kAZOMUVAgOlgKDmIbeu4MY0SU4BhpmUd/y+GpXhMsRZRNQM
iOaIiJPm2eaNvZrY/ff9/Yr0DNjPyfixTYKVqraf5S1rFkc8iacSptrouRQSMQYA
yQHbyrEq0u4e7twMiD+cgl0Yt9z0g+xFspiVCG/ovorViL/vwYWvvtbKESgj01/z
kulHEsZFzkGagZYeD5ms8F5K+qKOn95ZtkCyCnY0GTiDBQ15kj1Mf0a4FCBedL4e
IdrKg/U2l0AqbvlcGx26FXOvvNXbgi8RX/79SkO/I5TWBG5HBisgxJQxbbpUCeF9
q26QWPfzWi3xW9Ji1qrnDs4TTQwAYHZj4brKzn2kYMsFkAPTnluIwuOFEU4mV5W5
jPFsMRfRcItLGWrOaFTlVwOGz+g5jN+fRPx3I4qXQGKUene8mNzv2qbZwEUVGyoe
1qzb5JtmTYRdN99NvrIunZNcBsaTv4qxI5fRGvavOIVbGdtlKL7dn15v7doQUTzm
lepPigy/jAjWIxc0VW9hQz7CvzbpFPWF/TaDKEtbfJq8nt7jcuBqaUX/1ihcSRB7
geKjK5ZYADMhfvHjcPuDgjUNu0bO4y14z1S5C54jS27NP1oWxInlDGLJ1ZClzAbY
Ixn7JRoEpKQqU2DdmFElV9AZrkD4W+mHhm2qVdoAQbh9H+E2R7xG34nPJa2j9J1U
yutSRbBnAqBS23jzRUd8voHhEyK/uNLrtMYYCCOOBAJmM4Q6UFiWSzeoBimXW3Rz
hp4iD1Hye/nYM+U4IT4u8vNgIqBbM3Q9Ylu2BbQaxy/l/WO/86oLZC8JxtQBzcZh
mtKr8S5cQCFEMhAT5HTzW96/BtT3HMos2ufpRr9RczqMpnO9KNc8iFGJOnWa13jw
l2zad6efMx1y28uQK6wFSw5ZNXmoa9FfuXU8JvbODxRqAwenalIu1+lsMdIaD8BH
PvW764n4S0lvSu4nt20DRjzLeg54j5ShWDsWZtl6qR31ZD0qc5ir4Mhi1n2RoZfK
2Q96D657RP6ChaKVIvt6cR7M8WjH0nqRytxCkaAdl7syuqNRouY7A6hWxglyQX64
DkOK5mkyQ59rYcIA9S/1cQi0+CTX9yD0GZa43H/6kfIVYvcLHZiOJZLljuLfLWBa
3RmJZ9+2n5Bo9z7R25SHPGrRTml1haBdcB6ppM8qLTkLg6h1yUCfFFgVIQuvE1yP
TfWu8vGiNBl+tjK+0DJQvI08TOzOgzUmB2DGKp87hiG58YeNO8aBDt2Br4yJokW9
m/3AUM0Od1i42EG+Z/0n/T0wRfqDDCTZ5zN4Jxu6Zmo2Fft4UCqaf3V2sKs+wU86
NEHOIRdHaZmwK8abFZToiEs6xIGW6aihmAiMzLg/8SVFLMBOchVhzwdb+gQGF2jE
hYP3N5VGW102Q1VgWRl//sFOg/MZf8Wttd76rKqnfRMnpzl1W144lpfcgEi6ouYn
XUDx+YpuNA+BAA07aqvJQ8OGuGpXmtv83vnJ6PQSPNAJLn8voXz9mTo2dICSn3tq
tXSxk2AFjxvo8okZyPq3s8xBfywFI3+PkXiPd0qIT0HcbrAUbUB1gs6BFpHD21wY
x/UBtqwyUxxD6AApVvo+d0JYWkSo+vp68M3NBAsGUTHSl6kdndTHw5OsKITAhi08
ubZpxFmSMk0C6Py6S9tBOywPjtX1+OFSZ+9UhWcHB57yd8OuZtT12CMYY586SUSt
Cjq/x26qT20yMGoMSqTpdkvwFIMZMtHUuRBhk8NE+PvQx/jGxlzaHFwdfhKuFNhg
jL71Ihapg7GLUec6iwCO/563rxWBpitQcFdu+8fZbQGFwY0oeJuvwiDSSl+xMGnO
viZ8ri7v+Hj/BATAqIvhAgqLiX3OzXit6Kehr3NoVYZdcYDBhA/WVKQH2hEel/DV
+yGY1QuHGcqieCa4iwFu1vclX/vZnnrhDTe2tF6yL+XzrpFUszlr0PODUHWxEfQ4
x7aolfSVmjyJW8BszHOMJm9stTEA3Z33rvE3Eri0D6PFVqc/4yoIYSRndEpkd3DL
vTUYujR7SX/g8DvRQIY/46lTHJYu6j7qLgJIK26oXGbnk5jF6z2ivWEAtG48brKE
KzhuByvlLEEOHIFOElNo9wYJcBD0e0yNSPD7JgsUFgjlhnsC9cycqrG57lvh2MX7
J0FdzLOR00RF7GqjuHfHnr5xskv+6iPqXizSgitTJYxcQcNnu6+G0KEvHvg7X/qk
MhgcSQh6RV3HgUDtR6/s4LzYBCIgkQw500/LUpEEBfa6qfp1x7UstgcT8nSvcjY9
3zx5xMtdEpiDLB1dbzHW8kpFZ1pfIlesa9nGI5utwHXJ+QSn9bg11B1UVLxm7ckV
prlPgh3QKhaclH9lH4Nm2oek0gB4qpggx9OVPx/YMAkMbcR7wIEqKVC0EbKi6qWr
T7xngmvOJkBWLlHhYdQoE80ciIxPwGTsYVHrbklid8Q4P0BJIPaIuPHJB++szSLm
/sB5RA+xG8cWeJxAei8vNqBQFwIxKVOEb14ddm0Kd/+SNGEnSiiachw63Xw05Ulb
sATrccnms3R4bmIR9d9hixSAzFVFYH0fCd9xUFBVbzpyaIXmEbczpa4lxpeB8wka
5hpKiT2FsG0dCZBaeEjzz2yiS173OrQ6TqaO4+P/bG8hJ6yIr0Hyupq13ljQhVtQ
f2Y4oF1We8znzKZKWBF11Z9d0VV3hVWwSxece+99gloCDrYBrzXRXpoDvh5FdjFm
R0ToVRNZkn8W4csCdrdi4MQE+URJrY5s6Hdj9PGI4ekdinjClmM0l29/H52LlB0A
xSN3O5hxMxGF6g5ccO4Fxjs1uc8WFWaUQM9p+GtBzvmS9sxdljFFh0HA+N2PqmoK
/jM2nvnkAeDi3ggf/rYBya0VaiOvowvqjXH00KGQc9JuufVFV4iHazxJHKRq3GkL
gYMkvpWd3SlWl3c+Rw6j0iVYGZz+KfOPocDC7xAT0UbWkY0F19RCo1Q53XBJ612l
fcfiPkuRbPcNN66PrYjOf+VEPkCkwB5dOuWhUmqfD9Nd0/h71lbl9T63ql7jGGIa
HMXAUmk0i1+rLZqhMpsx7XqQ4TgDAbSgdt2sZ8KkQAjiCJpKe4FRs35HmnGzqYKG
CaEu5pyxjEbNyFYXzLZ5eWmQD4xwejGmr+ryW7r3UMv8Q+dRLYBG6TTVM643y9K6
Tt2qGsiGs7IVJAYhx1BvML9AsEqzkOLocHaOrqiinvOLkeNqbERWEJIRBncl6kPt
hWYGHO+Wm0oI2sCCo0rr/eXQZjDf5GXc5yNRKnPighcoMaPDfavOwF4cO3IvbUzK
Oo5i3mz/YNifWyepphcmBTzTC6ZJ9iZs0sYasGnC4n4Ell7Arlplna1ne97/y7ia
tdQZUlI6dHTs7AMw/AeXHPcFl47uTG1ePuoShPfRzPnhSStkNGNMSEUbgX+uROg5
iMEhGR0AkJSGhZ8ua5DjlFI/rHR9gbyU6BogMWXNVDuogm4YDksAiswHmuwCrWJS
6Te1FV+ZBqyjhtB6l7YoWiWTofliXcbj5tM3Rit9rUp9Th+qhG0LGq3yw1NTX6hd
8gdUPQ0gRr6o0aJqZdU3nl/uIQkGM8Z7jP4DeYbgkaHu4Ts0iCownOha4Cp6asAA
LwduQRm6p1QrsIsYXMWSziqYNh37XUvYjJuBzDLQ2OnxgTliJZ7LlV/sRN2DJXAR
9uc0IelIPHieSGHctT+8X5zDtp7iFUHfcMqte/uDBosM3wWCEeifRuq3EQMiTuOo
l2kmAaVCZ+g8vsp586FYMbehZWrjTtNO6QhtE1IQUyUratZGERUYK/0K3mEYlYmQ
pv+ya3pBGW9ofveM85OSpGyle3laL7+Tdo4XRLOM/YAUnRCYxfZH44iRrOGB1o9x
yY//xpA9hGENxKStmC5sAgI6XKtwrVZFLDzvj8qaHHxQdTZUsHbyophyYYauQVIz
9/P8QUbHjLnP+n2A9fnk0JKywW/t94DeDvGxXwflMuEmLs1fFQbLcxuC4v8SiQtA
r8rA4CCRFOKH7c3KF6GF4V38AEWqAbvu4kfqRPC2J6rSiRajgyYQ8Va+VehnbPzS
OkPO+vsqImX+CzO+UAuJMTlcUYjKC3ph9xwBmiXfTEcdCxgKeMbTIPajKbPKHx6I
68f7l+BYFXGm6d4rVnnpwUS+kokostKFpCJDWOZUTyacIuv6nzLARkpZFLSMyEWf
6SYo6IpxFlCQzVbCh+ENs9KAPRBv7mjOgqCrZ6FBf4hjpz7/yo2epa0TBWOpVk0E
0dFslxy/lmO/raLfQkv46PGRS1Bnz7ISLypbiR70DUEZdp6aB4345J3VW0ygqIzg
u+KjgceEh2Nmw7DGOoP88IDOgGipysSWIjynRzmMp8WHudLje1dE+9cCGywaXiRL
EW94y3sfsVkOB/dg4aH8LS1iAL+XGN7FLHQrzhMoMPZ5wzkrt0REOrJOxPkX9Ido
gYp/teBAO6E28/x6QywEKRDYg8ews3zryYVhGOre5Jts/JjU0Wjnx9Z33xiLjRDE
oWL3Ttx8SaLynD3L7re0dIfNSlzBUkCX4qHZvKEgVTvZ1Od/xAFLmoG0EeDRndjV
bUhSPYvHAicc2DdOhwgGBnnROoTqfti6YIqhplu8QiQA27Xmegi7xQIF1jvLgZYP
8uxdRq3YnyfTq1CVZcnztmmABTyqHu9XnfSR2EZp7ZDDDKjha1Ui9uZrTphkWvcs
keVaQtIu+efRar3pF+tPt8LZxTS2tSQc39R45ka1RzdlbZCmO7uZJcbjN9Ez8Rno
fQyp9KQxasxeVRR0asfH8DDSY/0aVUzS7GtMDDm+3SbpY0KII1QDNpj6ywbGtKOI
F4Mv93eq5jnWXSKQyXeSewZKkJ9i0mPsIUPRw4dFH0vrEX1Lt2Ha0IF5D1HXYuEQ
q8Le7R3oWvwcfdDepbQ7V6XEqqo4jpQSBTo/IIx+w2qbM4OWM2uIShVQve0PXL23
BZcnPHiJ1FavdXe8a28wrMZWpqo+wi36cUN+jXoVG3UFhl6ZTcnQgJuCbcVjgPtz
94QROsxL+/C/H9N2f4G/JLTlJi399gjnw5Mz0cGEmQvJHVE3Y9uE/8nVsG20d19d
v3xsdFiD4YTXAvYGI8lLVQSQXq+JbfumCDfSoXUSDAb1K6t/JWYPTzqU27hIYOL6
loPCoF1B8502EN+ryqkuz5KXtM9ZI/vvQSqar6DLISDfXvTxljJcOrMcTRkxVvmK
PoMK9CqpNyItgJjjzdej2OAytsvayrG5/p0RS2RSe5fpeuDGGAq6y3dfSNw5Yw7L
UIiwKU3U2NGIMmz9LU8ijIMiFeYQpj8ra7PAW5+jaOblw80gzPjeZEGvwZfpORsu
zuqlRPtybuZamRC4OYCO3SkIvR3106D+NS0MErPYITtbOcFbdgxyZYYOomSPUykc
rY1la5kcyB7heT1Xd0rlYsG/mJ72621RycAtu3HEPR0IoSQBEmYD78sThlXPRHP5
TO7n19GGqL5z1swqE82om/FvjsROfCbEtl+rqJkdZ3QAmfQj5NguhHUY1a/HotfZ
o+0x8pH+vkU/zFFZXapGrk+ayVM2WFY1oLXQgfrxGIMfFCYX8Qz7ZhjlzD58RFPa
DnXSkbLS9mfGSHM+6o0vDxQRP95kDcKhlesMzJuY95ia+dSO0nu+mBqa8/kYXI18
+Qt0IINxX2dGMFSRmVykhQ8w4jxQ0qDgAbzD+TpksIk2BOOJ3DLDuCQvfZKC1/V4
LwkEi7SaaWrHCOjsyWGqQ+wgYzzoU71SGWffnCu6h5/d/Kuas65a3Wav2z2wn7Xc
sg6BKnbwCH8L3oR6LCQckjFe6e8pXKbNIt75FHRu6lhtlnQxCdIQYxHHTwzL9Cs4
AQURGqJH6pGn4qTKG8L3dLPfJYx/p2+h8wbh5UZdjmXtRGd3pV6dUQ0+NaLrDbbR
Fd7mUlv1wpaLHkbut+u38DSWBc7aMuhYdGaB4d17GyfgiYoIBxbv7yd/MqsV7WVw
YSKkZDhr0ybHb4dChw+N3AvCr3zE/eOUl7pX7VYJZXQfnOWreBWQbUxO6A8oDchU
Us0ndOYWhEB0jy0Ay07K0VRU8+wC2Cy6CS7sqeovJusGPqvhIpmzK4TDdfgbPiR6
Scl2ogcOcGbmZCAvej93N/Mk3Bkwl4HbxJ6rHu6SrEkuHj6p2vROULN3dbQxdmNW
6/t49QEFryut358YoxjccHW76PzzUekomUet8NoV53Ym0h7UjqNnFaEJJuczcf1L
yoZJcDA5eDUffnS7BnYTQTTzA933GkMYiYlw2M1PZmnFjyzegpqTHL55ZA8BlA6X
FLPqavNegoh4I5EqtKbFZUX/8L/PTwcCEkb9dpRubUuLODTbka6DvEBWP15us6Ib
bSJ84WAK29J4oWTlPih10ZPl7YM+M+OoRycig1cI8HAVJkGdpwiQwr8QRF2seVJJ
qWYiCRaW0d2mabps+Tj3nSx4pzgdHvcYwNx56O7z9Kbu7ED1F3ZrKvEiZNLHsP5o
dObB1bSgLHX3Q2hIzcp/Bi8RZ3mpOjkH36yQIwjPm3Mfb8YjNKHOx+dZXgfs9mRi
O5JCtzeuKzQ7+jCxMwrPIm0br97ft+ip8ySO1T7MfUON7xpSBz8C5UDqEOgjeCY7
8Orl/K8/m56vclTzndwm9IUldOnW1rvWRGyAS+QNaS0bcu4p0ld5X4fRrwznatH4
VHk/IcSeTPoIezf5173JvM787FcXIvnWobv5P3Tgr9WHmvnm3p8z3Ow046ZIXccC
nHjU2z4JmojC9iXV9PqRuTo4Ensf+6rjOnT1yPL1njvoVEEZGfwCzWFcP4Zsvk9T
29urKlnNOD7yEo3WqCX0MA/rD2t0LuHdicT/0XAUzlzJGVsdS0GBvgWWnSi3Lpq+
UYg9W5IPHjvP66EOFosRNX0QOl2fUTN1m8Qe30LXSbeZJkw/MC5zMu25+8OfWLPm
GAeCT4+P1Rtvbv3vcX630hpTkJBxwyBo0RWordSMNbV+7/GD3rdYaQafeJvvR57r
Kn9HS5x+7l8eDxOg21jAjnq/vJbbJuxGkHzCXH21anZehPBPcypXWveZukgcJ9JG
Um5pRvfZ6mxwaDwf9NOChfhTXv+3D2sPX6jCpoO2R7hKiZTBHQU60+y6+/T+KwZb
zNTdAqWrviRqnbyZVTqiNTPvOPpjLDlNpe3d4qtOAFVbmwDrZfg/yyM3BkxeUdiA
wA0afCv9o1ecDrvProoZWpOwS7AEWUD6BoFglIV79OGpSAKHeXLwWXyPxbf1UF/6
sS0VBVzLiZoAmw0UtZTvvfXWx2v+C8miEwt0yibQqCIULN8nrOYf28kE+tpqoYi8
PrjKuu0tIDt2n8b66xy4Eb20WQVJSSjYMAKMmMTREAtX4vfsXSVMM2Vwk6cY9UyX
azlr4ZBZEkX5uvMVP9M+Nsz+MwRAs169PMsTkPYmKNs6xElAF/7zAbvBZN3Cj84b
m+uU3PqaSydEsdK8B97NdD/wJyaEpdKJCfZFwJeImlTjfADPtXDxbG0HPghRezXU
MMjrGL3FXQP9juKvmCtnPzsrv0gnpfSMsGsd7wAOO+ZmCozY30G/nQG1ByjrLXuO
anREcvBPGOMWMideNrhl/udfFVbOI8DH7Tn+bwNxz9AwRVzONuHKrIkebZHriPyp
K3PRtaDJVNjQaW87qTEBoiqFT9R3aSba1YrsIkPFBnJ1NbquxqIqL957WG9uRYao
L9SmZpd/EKR7GvyE17E5BJX0A3Dg1ExPFv6sR6ouJmx+zO10jbrE34xJQWoSrMxv
M7onBUCIszVoy9hK6fPfM8cG4P4hBzu+vjQ4rdn8kYY6LJIwdbEUHtwhMuWYv69r
+xEhAtgdDKK52e4i336KBfokiOSRj6l6X1fZlbKrwA7e6urSeEugRJ2+g0tyKqV7
on2GCChWrEcWRKFKZlL/EqMa2n4k0S41KfStBztoiT77AwGetSkVUFMM/iKs6fIe
m2G/CTjaZXJDm3SAr1LZL8ca+ZMH0REOp5o1wiMetmIM438ZKmhG7X4B9SSDuvkY
gX53o5+LELDbkRm8RLFEONkzBnS0H01EO1Sc/beguE/cLXyofvakuBt8BCL4bYBn
jw8AkrQ+btZ+5KAq4bhnS5wnZfx2sZSSV7eVd8oYsItvVF/ilB6pqSQyu+v2NKsi
GJsVeYIvtqPKEwcL8d93mELX4OlDdXYRg7RGIyc0+AFvrOHJFMIQ4RKWy0hR5TVD
eTOThWga4e01bHq/rDyHb70/6O7OMG2STvnXI2+vzfhc20JnT5WVqdus4oDiCnXF
tm+DX7QX++SWzDjMsqDva8viClTMUmz7fIQUJW4OkLW/V9lseTfEsK8UTB3AcjaP
aHAms6XxoBVaSjIq8RgBfWCEDwikIpmxAPPZ/ogDSOcfDCGOQ34J5VMC8LZAWpYH
yPuS+q1l9jrZMJaYUXatxKG88AlP+/YKufuc2w+VhxfVVukOrPb+kaQbrzAZO/Wo
WEE0d9EgIhXgBExm9St51wgh7Mw9iyLNSd7tc9HUrdUdAFBSXFPGG63LTyxWv7mA
9Ir4MgelbiUxnQqxAssGb67bO6kpv+xhyLk/sy7seTGQ+warqH3eOwFC2iRnhrk4
dt2aCvKUTGKpSa79v1ZMP/h1VtxNy9ogggm0BpZ6A0pBMQqjWh9PsqfDqkKf9MiC
7QRCuYJMrZMgqYSCRnI7WRDdoxePxLbfN2ShSvmLcrJ3KJc/du/lK2ZqMzAIXWxy
I8bvLFzOlbR9yd1wk8ZQDc2TPi1YNcbcjsRbHmrL2Js7UrBhhixdyeBe+8yrH1pz
gCpCFSsagHU+KemxtFTmYQTt85VnVoJ5jStuxFpaRnCKZAdbYpd6HkHtCbdBKNKX
uQVz/LJXFMLkqYbxMkM0BKzuGkix3kdQ99G3g0a0iW/SHcB7PAhZMm09xrPV9x77
dyWKAlFc9gnpQC/TrdXh4SJ5oU3vGUmIveIZZiK1EHT7xWrPbdMol7iUB+N/Fvxh
L+ivQ6GdCIWsHALn8XWr/rv7AVdKtC7h+lR9dF4J3LxV8jfxbj7LWUKSysRpiuvO
fBrVPx8qF+rXB0ITzVs0YtCvDgXEBtx/6BUfvwBDUhFApubh11gk4iDq9lUAmslE
c33/7DpuO3kwn/Qr5H5v5JR2ANNwD7CnjrAhGzx1ZtzLwdFwqGXCOprA1HOl6I8J
T/ueVSCYrOfQQN1HnjNcZ7wRFWQuzPxD20RZW7BC74J+lEB81WyPHdvtlibAcZ9k
5gxf28MTfPxbBXYz7q4gwbW0IPjFEUAF2wvbKrKeVFEBzuCJZzQZA/TLf4u1mJlP
iplv/yTs+Qynbm3c8e/eugWFnYT0Cbge5kg9Obmen+E4FcNthcvT7a1YOEeGODyj
CGAnkkKyCagJBdPVuy0NhD1OmI5ah17YyaH/I26s4kIabtippWL5EchDBpcrDDaw
3VW2HpJ1mSG82ec3JwqR7sviR7tZVmpSPn+o7rlnGRNshN5mh5uNv5FkXY7KjkZR
JSj5aCqee+M1o1uQ7djxiHUEybNq7o317JRjl/6zgTNGYf6PzMUr/Y6mBKDvhBqO
Cy+CXwFtmaLxdhaG0Oul/OWMIWXflzK6GonkGUxMkO5x7ceAPwgubmsDWFlQ7W2Q
69FRdSx1OFk9mbwyMBRxTW+ZmH5qQtePv8i1MoakoJj8uirPShQmbSN+FCX3W3uN
PtV3ZGxPhHSrcLqBTPX9lJTmjjPwA0idRIDevnHEq1Uvs8JceIuzruAZEl6kHrTZ
5vDNWZC6kkMDIvH/jGWLNq7RQlmQ1vdpIVgg3URk69qS4M80XS2h/MoAqw5xXd82
afXSu9nwbs+WCnoAsNk8K3HTjnQsTVriETe3W6/lZFS1yVkubuaTRwhjzq1uofm0
bHJK2Uh+3rBPzQ1LdJUASYn2FN//J7H5EKY0W4jm9RYfkuwLz6pBUyHBYp1NB6cn
MLm86M8aZtEMfJINeIa6AiKq4vaiIu13UrMNnGWmz+4OZvBPNl3gLLm1MjzIq2KX
V+veZfQdLlrGylP1FvaUeO+p3HGaQmBTZVzXgeUv+xTQehQRPFoczrvvXoiJdRoo
nf3oFGjwTySReui3QsP0GhBb9GhRi+61dGuruiWZXxaOxQkyptX96KiYVJYdYcay
I91W9QKv4aFRxXSwPr7mfnrYrro59hJK9trCqRqN/XDfikmI22nhmh2zDO2/+3/r
w8EEC00m/GwCmAnwXDz64nxi26ei7bCPnQpg8XkBHIUs/YsYIgw7l7SYrHlFq4EX
7QdhLxbxm+uBBdMQswezN145pAJp4wEoUe2zje5tBbE010lCzzpYST0R5YCSbGEC
WzvPqxS5Tz+spD04+yQlxLrG+TRIKTDzfBBljp1x7HJHynG1Xq5aTrun5GVrgssZ
sycY2UKiHoiKXdVNbVkvacAFColsRx3r0OLOLTuKYMbMJoSnxGzR1feXD/Uvm3X/
AjDxpTJYNR+p/zL6EG7IZFK00xgeYvwwKjqYUusxHJDqhJ0ZSCKb3LGPKquk5qCK
Uo1Ja7fUzQHq/r0rvnr1PMrsu0M2izKpMH8fEDmmyP7nHmxCjGnMqCAKj2x4p7QV
dD000qnySZgDhgNmUjBVVS2+MdkiFZfH9IjBxyDUwZwpoRFpgkjifS22fvBBbXck
iVdmXHyGIfiRhm3VdRcwJQs52LuI3i2embGGA1zkYH0AOlXE4x3P6yFig3cd4vcp
2a9Dkl6kaQ002n6YjVeV01m+NlmPmOgZevpMNjtyKLkmCtMl7TMUkF5rngJ7Zd7y
tYfxoZnV+J/rqZU3TqiwDwcrd+75N0PXGeFuSWFYPRR+biFGwBR+gqVfJFmSb/ui
Jg5Ul4dr7j/uxMRkVWvz0N6L19QuGw5N5lHKX/JdOG9enPABfRLue0sXERnD67iL
hK10RBTD4N+Ljp5dX76KR6gMm0vim/MSaeIXcRg5R4RknFJizMv6BR/nw8pSvmWb
EyBlLqChRUEfakrB0WQCl+VxgyMVlOkgZauxNhBR240/aVI7diEHC87A2v7pwU+/
v0v2TQIB3SuPi2AcbDp1WysdlfWnl/Qj3H1mz4VPTX2c99aQBXpOp620xiWQoICd
91PgtCPhO5jta6C4aKvOLyYaWak/7RihlBTbRibXw5ggdLZEkd7bKpjSxxHty/or
uDABPtciqd3wUd79eaStkXvoDRNbOkv1l+VV6VTFdCKFS4s4Azd4AFImRTmIZBMc
f0Lf8V4jfxj6bA6kdj//VGi78iDFjlxJEhXnzUwB2lnCHITi3/JqucI3KQ1ryQlc
YDOoA+39+tlT9ONq3pUqsM7uAEvR11DhnL/YX6FK9pP65s1zTcf1QoQ0zJLWNfhS
GzUXlIcrOUTEwJuEB213jnJfEER0NVd9Mwqp5jM3WMbRXyOOAFKlEfsJewGqrLMP
DkVnbhQHVso8OeKieZ06cj+plHEPehKquWIzLCXSGuFsjdckeyz2zIYPci6Kp2tI
VAJDEzmenydl0c7VrMPkH400BBppokwXnf+OQZy8dM5xMmzS2814EjkF8TwWlHwP
wtGMLtOkiOvQr3/RvXHn00lg2/fCdc/MSbOCfyEvd0hNbXZnLBI6HOg6u/5zAZ0i
ZaMFUFaja2zqMP9UWY66v5yRRZy3+XliFwaCpTJkQVr48mxYIMQBgeWVqx8eybyH
DG6/Z7vjzDq6raJIfTOEo4mkuClphTNADcY6FvYiFVT/7xKVQao5Mt2QCrUpmfDh
Bhhsme/WnznlWOvyRmAr+ArnMCHsy3BQXfLucQMCgUQ9iG6DP1wSRiSMk7Tk/i29
SA21GnKAmxJFh2SqXk8VsIba5n7xPd7OrxaTZVZoGi3EQbxoVvYza5ax8aRkIb6f
zY/uUJCK7f3gPvw99r1xo0J+I2sjgvLVlhYcINHkdinYsufGl7A2i45UDC1h8jQO
VCbKtpbckM+o2ID2tLsLbvgoYOP5CI9FBClAco9DjhKNfmlEHwWks3H/fpvWr7HH
1Yv9QjBjtJxrU3SICf83GFAS30iBYFGVNHe27V6yCD9t53PIKlyX0Oyczz5GQJD3
j6n4olKzBC35i4RTd3sc5Gw88N2I4iES6uLti3J7t+f/Qlt10yKwGVoKjX6wyX3N
d/8cFC1rVdfB0wABAvkF7jwKMmzcTGlTIIDZq+SQ3wzj1aqrnQNlQ7BuKrFZP4ax
yWfUovxAiNqQnMXHLb9sssjNgGZJxSMFWxswvQm6YMwVTfgJXrIU/8Ee1v0nG3Fa
g36ded7wZCUChknktMw5j8S96YiMaGV2pkW04bRf9nNoE0jccO8sgzFg9P4loia4
v4YTlQyz1PZziFPgm94NidWGL3+VQXYy5LV506vwwJBw7jgYRLUYQHHHvnjHKQm7
bGUhkJG9T1jzgdxAlPKhLAr1EuR7HhPBAf07MFXOMIBcCRjw/buZuK7EjVkHTHuo
HBc9ZirpwpBsKs6KqpOPY5W/OgFNZDvwhaejxLoyzkRZkU/sR2CXEKYLkm5vGGqe
gDGOYr47vco06DPKRoImKm6OlGXU598Embp4DXTG3hNTCvNA/SHEmaAlqArjzgSR
sYgCYN7/r/EcqSHrH1aDJe1tu4d0NPQPkFP3B8jUitKXOrPZLTuhQqj/u3xpt589
oreE9uuCVddHG+vvfYwQUeWsURQQZ0fokBiXWJTNsEIHNsMuI6lddhY7Tdy637yB
dx0ZlneV/DmS+QkLo6/vSrOvFpKFsIazBk/95Vl1VsmlNPpxzdeWUtbLQD0sieHs
BeKVudtQdcGEPmV6WVZSSN9KNGxv5kO2gXnvSOofmHdqV80ffr7lbvckKN7IoY3T
lTt3kyPgO5QXGM9qL3EWwZQ+V6eoa0RO8vP5/LykfjDmlZXGTxCVBRxVH/K5vW+W
jM40cbujElsNc3ULsv8TgcVO61kjPVlnRCFkvLJ1/Cbp6Zra4JWRVAbPiL3WIdQV
joHsaMWHYrzinVefU54VR5ijneK7bZiI7eul6NEaNORvRwFLaZUv+q96z4hC9B/N
Vju4/8uHIWEtv0b/rGpQDA7PWBHBtrath2f4S2gI0uxsuFEhC2shi86sjzEBNjUA
Rcin3+V5SLMlIuK7jk8diHpBYTWTuFEOCf35KeUZl1+3dkw1wE7EOYOAzDwMQqT1
jeWOs7lSDSl4fCZ/DJKt0vDF8YlnybA9TLx3sloCNezB4gWhpbb0n8jQez0OXQy+
qd4HyBiK0249fILxTsC3QH12xmV/XiN3fyxMcitK0LOjLKOYG7dJpZJiwAV6tna3
8a+VHUg26LGOaqpDbpe1FV4weZK1m77sCTczDy7V3FlbPdsbV0DHbrT///hdV4Vr
YXNpSPcyRFMYqyAt32uQ5mk0mC7hrQfcwI/79cTt8JRG11GdBf6BjJcCgxT9QzfJ
UnwozX2zRrrLT0inSEsneZejF2lGDvODCWtc++fPoZOqWlFDm2G5TaB2oCs90XnD
WgROQpBu3nvLqsE9EEeDrrTqjBEhtp4RZUZafQcHZ6KYe6lHMV4+6Lo/kgXTcaS6
tfcaVH6zNG3dJHMQJEyIHoiv9ZwnMYbUGX23yqtk/ZWfTvk3GVay8GLKxcA2zkBf
t4bbySBkXmjaxjz8iH0xmj7iU3pfZJvKwj72H7kawrlUAMlJxVMz6RCYcx9kFtCG
Dv88ZeR0XB7bSaYRU05qu17j06LDWAe8we0sc5Ttihf33S8tYFj5B4oqlz1GdcTC
4tu+d0CAn/Twn15h136baIGFQB47ZTKFBBFxd57dp4hkO48DtxXHYOMgFdH7hLBp
yMzWhXUtFmU9c58Rpr5AHPh8+o8mj4GXZgFnsZ8hsXPU5C18sJ1/XfO8I4tZLBk0
89RfSlvv4HF9/RMhw0jw+95DU4YI1bmHw/xlgmZI706t7+9xO70Heso3+sGsp+Ur
u40mdZ7pIlCfPihpyBdbq++KXnl8W7WUT2Snjo905a/vS99m53Byn4szSBg3bHcx
6OXZ29sQYbI9K9xui/6SixbBNggAZRkD/IecVvlcMxkN9DAFfJ1aNQnSuOOAdOba
zmXOdNEt+W/0M/fZliWqgKJOpHSZTofHtwMwrVRJOpw1O185o6ERvckEhUewQuWm
lRW/xnth1q67F8KHUoF3L8fi/saH+hNwFWg1ZoOGVs2/GlgVEBNAWfRPuUX3vUyb
vJC/BhugeIp67XA0yxB8mIqfOeC976rU9jWFeSG57v8TME+ZK8fEKh3dKI5GJRva
js3a+OBwzIFPMC4E+KSXY/sfmvqqGzjzNE75q56rlkJacH33RRODYuDbH7ocBSU8
ZkbQG7D/4H7avQEBYmYcYnx40eOPYysrAazo/eSv8A+Bz46KN5CEhg26lBA2OoxP
U6B/gWGVRwY77XIMtouhYfykedBRo6+RA9mz+lhfHKVHDtlWRDJU2HstguRCWA7d
zAQWX78lv1oXsnxv8zHsXpB3IFB9a61z0VZP/Z0KcRQFsnPH5CMHF3dzd7S6/2Aa
fQMQ+jdxQDXOOXJ2IPQT8FfAXUqkop4mGFkh8TSU7cSL5yf/fZ/Weva9g5K3s3rO
Ux6R+ie1VDGLLrq/KDOJIJzbZIPssd3Q7phYA8Su5QJNwYqaG2PVfCtitd01Z5Z6
Z9seZxmbpFA1aUBP3UCi6HhPZoRCfb3qCtU1v88P4EUM9yaS8GL88nG4+W9YILRR
UiI+qygRe7dLhR4tsHzoNyR7+o1ZNia3no+iuuK0xD5EwWls+6L/+x90Aky7WZve
kNORMvUpcQkvWnuVp06vQQAxwlz9iZvTj77tEB05EP8PICrfvLKYw7twni5xsvPg
RROAr61dh7K9Q+uWa1GgGP4l2rY+QP9EE62hxxce8F6ZgtVIEBFUf27blbMXzaTq
sRXc1z/2YdxQ8/cux39MtDjI2nGs80AmUINIitR4CvESe75SJ2BQ19rjDR3cGh+z
ls65xLb1gOejShJfEP9X/0uaUfRGYPl/a/dCqitCVkljTS2uKdsOPolC+x5bV6cE
qxQjHBIeY8MxGdW4rxW5EF3FwxXTLOcwC+lUKLRfW5NAU1scmOkQgCssbrQi9xdw
WxLe1SEMGh5qY/D9wo0Om79bmGkxaZ69t5cq5HYxGghOO+Q45Rx3P8v/5UQxSuhx
JSeHLGx0UZpW8dq0WNaIkHjJ2XY/5HaJJ7MNDmC9mJtAhAP6tpaXarI/Ek0wdiUH
eIk9s2vnlXcsCKLQCwoPP1JAKGJucZeud2D+Fvehykhaz1+Ymaei8DFymSj732DU
z6CIWgxViLeAOjMYNFWCszl2/WQjukNmNz1/IdhHU5EUUTn/RPzqH9mub2Ec6I7O
lj5dRHy9C87FoWUCp3HoHqT9iKnTs9GfLrnjZ1eBLTVznJtHD0q23syrYyTU/8tl
rtfDKWYM98DfjiCkc+admJsz95K7lcAWs8FWtOhGW8+CnJG7ckwGe7euFjQPlmq0
tS6VLZkP91ghLnohfTi7+wvH1wCYn6nfQk86+cxKgbQECh0qapvPfavCOKYMkIkX
e/WBXEjsWXEZb7jGUsfmpIL2fxDiVXqbpoYjvrH8FgFzaY+D0aCHDpntW8xiPxk+
s67Yd402znHRZok9/0VZnIYvOolMu/AMDd/HnfRh9cfKvQ2gS8TlYtK++OkCAfXx
Idvm5jNV978an84B1mEognuSWEjz/sfB3/HNi8g0acwvWlQoqUVVjD7/wBy6Q5e4
GNOLJ7BIHhwwvYnMqXGv7NdOD1+S9Kt52iJPtgLKowjk3AonYwVqz0m1Yi2Eh9gm
TMHCYQlXnU8KrFqz0QlMBvlXF1Kc3gysDa0y0y5r/jQQtKskalaaa6v3aJpga1iT
/x7By9Ok2ZHUD6cuQo3Z32syq97cs9mK/5k0ug1KhMRKHc01Q1r+zrgzSobq4lby
oqtKPa7vORPNos/MAL2RWjiWi0/ayiKK4jvf6jTCpurtxt6/S1ythf+O6YSvH8wQ
UnukT/FgOJC1qM4Pqnra4Da8Z3UeaTfJjaQae0ho4QMjEp93E+U81M38UokUQTmg
Ofca+yysE8ngVdUVQNELfG+H6XHv4tZ4D5W+wgDbUxOPSR0ePOaPMIXV95x0JI++
N1qHDSNvpnEJhhOZFFxV5gcLOwsagGZZOfa5Tcvo41BrL+udZdXDY0M/fUie9vUQ
1CJ7ZiQqhI1Ff4/++J2oL5VFd9YwpXf4Fu06RgEI40fmPneS0eJMhSgBCH00VRpV
9yg/VnnvL8JFaBmON8K0CrJl7YV3CCMwE6cJJOZsLnB6poP7suvLzVmhQaOzrM2W
nGJztwaitVmSvLLB5EbPLSJYmZujw/r6JwUdUtapB6T7SHcJ0DWIDC5lqROJlE2+
FNqC7Y01cYStw8T2uAiH/If2XJxLk/wrQOZ0YrYxJiXVWfNnDAue9c9tIluyT3WL
EZZk3Xs/05s57Ri4yxDkYzyG10qcPke/YKBaINDEUIyE8ISD+x8DgVXdcWjMu1et
yuFpv4R8ZxxNGiad8zLGi/obr14/vI44ng12dfLcQisNdze2lMrYW2H4vFFRc4t/
U4jjEdeQOQJJMV6auk301FaVT2IUC0NWx+TkGuDmXhTT7ff22ZpmZjPD0Bw6dAPs
qIFYvs1IowCC62mBj8sgWitUsOp9HPHyhX3clBRtCr8VC8cpJgfHmM+d/MqXEMqE
/9hy03ZDRbiY2KPh77LLDlzrVN3IWZoVdlyODZeZFw1/x+XazGyEV/P0SvPg0SUe
HGiN4iH26Sfl4fQhAJdMmTy+2m/L+KU665P9/rNhpyBA0z4ujSjNXw92Lczo3/jl
lA6U8XK6t18xr6nfrYQQpTIS37nRh0ABK2k2Wf2hGGRpwfqwPd9L9MKuN1qQSz7Y
PQPQpLEDIBgOB9s6nEy7zOzmG2DfimH2AN42Ax9Q34LUIYP7JnChj7zpg6ci/zeN
7VJxa2SL3Fgv6COtII4/NWLmeJkd04m6S/oa9bRGHeSz1+NZtykxjkvLKVqPSRXI
w6KZN2LlrP0IcDOgHchZZBhtCG4MJyLl8zzxely07ho5Mf3VBYVtuQHI44VpDmNe
RRgm8qkbzOfdPbGmfROr2C8DNLL7qM8latSHMP8XA4WgevY+2VS00FuqJjLvQuA8
UH0jTNhsTQ4T3Q0fzJMGSCX6rPYqTvyDohoTNHZaCOXAUpLEqenVUTKJiOQEKh7/
FCvqVaOWKeLFd2TzW1LLj1do58uMeBJ2LOTDbpSvOkPgSwwFxhgf/xK3qHkgBl60
f3mLpenG+6Wg+NO0aeb2k5i41dNCYlLiulgX02/SM7ejhTaCry/lxstB1HAhsPL3
gu/IuvtATywFjpo0bEDoRvTuAMK7miFhd/4PzlQP3OHmxJxQih/QOJYl7eptQM3B
6erbxnGo1UUS3Kl5ivDXMQcw6eYfz/uoQ4I2aFcFIi30Wg0ganbCbzsqdPXg/ljW
v5waDXQmQJ2TVC7sleX487V1+ov1ziBbjebvPqJIbGHfk5ic8D+LUNkOsaEgOOIs
a6ZR/3dtSOHPh75A90fFnZe0o3y+QLQ9uOhVVmJ2hDtvyNtp+N9gSE9z7KdK7+pm
JxAaE0PelC67yb6gP55/g4rNqdpiwmvtAxOCv3krOWKywQwXniY/w+dPvRpdqCI2
BiY+v8dMvZY1c4aHcLQvj4DrtB5SYuj45J/z5SVisrrCy86d0pPvD9RRzVynjyI0
5ff6m70z7HiNWRtIHnIEUpnM167FX2Y93BOVBMaTjSH2rhVC5F5lZFBHvLEiHxTh
CfsDKDhxejfKsrMNeFUugxGY4OQ/IsfRGYBiRwNlwGuEDGOzxP83Vc+EaEF/aAgU
4tCnldz7P0xdadQqx5hOwBW1VpGAR/MMwoUSKCN1ksfPSkNpnCK9MvYBRCkhnCiJ
sHXw2EaRFN7eWyAuDHqOyu6mtmbGembpUyH8VJ/zeOVVwXoSkKh35yg58QBA3IPx
5emDM1ZnP1RyDcQ/yeRcv8fKM22Xw1WXKH8Imc7i8YGnFtuiJ2/5kgw3P2llFykP
qD9wyuwoNRpQL21GgRLz6XV80CdY+nBmmJkjODp5gIzndIPlYSMvTp1JL8fkFMQF
1hrODY4VWIdktc5YczEN3Z1C80s3KU0sIMAYwdu/aQoJVf6TruXW8gbGqbW4d+AG
APXXqumSsijgdDDVgEu2lWvr5ce+ccNAygiD8emqHZwdqIJv2GrOiYUXEBBZn+kg
tl9K0Ac+JpnlFoVERiZrdvm304ovdvymxe9aQpsGxSUOTTuxGvB49l6jzyXKn2nd
s4NLz9lwxG98ZT+22UxlKjm9LbHcZdDjRXLgOkoBy8nd33pbLwsiletURBtoehTi
xZJkh34RIetoBsbC7XZgYQhpifcJA/FvbTLkh5vEN5IilFX3kQ0jlLUTskU2BF51
X4lJKBK1O+sHFW7UZRFXel6is6tFo8kOSvolKaWSjJtHKkeOTZTRHYH3gs1arXA6
oOmSn8jzqv46pfsymmLUQKWE8+dkJEO0UNIUo1pcIeQ60LQrMGHMsGA/tRxQ4Nmp
e4BKYkEzx/5alHt9uZ1hlGdvaLIChm/J9G2VUx6vFKlifnPct3uyWQg1nPVEt40y
608R1apdXVta0SNO75qEaRAUXinz2bIxyh9dF9Fg+4aBnCRj6s9wKeX8O9+Aa3xY
krGr2JTXYEIEet7Lit7ReDCfTd0Kqct3pjCZhC3txbR+4u8FIcxxhPkHliKrT6OZ
dMh5Law8w83thcw2/7Xs5vvmbUfLH/zb6f5lfYGaw9v+wg8nDyESsiXIk/Xcx6a9
KKVOzGP4aA6SE0RxsdVoVicpVjaRP7lkZZtZLrQgP89zRhXPxYn0qUTH41nasauZ
QOddIaUvA1LJ5nxD126Gae/SWUazQbREM3t2vBNEaLXx0E17D1/q7uvjwXqCcD0j
/C3lBat30nxFA87+yc8juO7b/czRoFPsDthlU4/+oA1aV31+LBADjHYicc6tgGRs
npLANXnyB9wobDAl8YjGI0pnaSCdpPvQkyY1bZUyjXZ5hFiJaVbqEmQxmVH2+5Sr
SzJP7xFaDfja2+FQjD7GrON31ETYDwIIjlGqlHq/9TPjRdvS5y0pmNZ0rqSV7nQP
++45m/sOI/qsdPTqGd4YPQcn1ru7j/itKGnVdoh55IOgHXlf8OzEKMdfgQamlHDl
P7yMNK9BdXtq5Ud4IlR+EAhFXNNfWEFMITTohKytC7EJWbZJb7wRsS5B0Jxr3Avp
alt5qJFidBML6OR2UpYTcH0J5oXeuzwkUmC+RxPbEBJXn+Om5tfa8T3NDWXRYoel
WE0rdTevO8hKq/zwb+Zx2wZQX3IueyDEHrlWyM+BKO+/Ema5G9fY3TFsSLwx9XNT
CJIPvKcUseFBpHlYcUtJD0OZAubGEaJMytSMGMUX57+EC8W8iveTiWnTUyzUg3FL
W0hMictyB7/HklGZbap3vp2rDpv8ZP+Vjll04yN7Ufc/gknI91TWkzeBCm6iHMa8
vu9K1Ca5Psv3E/XSu3nN+4ZmRukk+KM4Irm6OTIoSPJMgMTdNmSlF89zWpXg1oAg
k60Maw52cyYiFgLhSJ99Sr4awgwa3OPXhpDYDJXi0L0XEiEw2P/93ve5CwwfIktx
yN9cxafHDBlCGfmc1fVOK1n9w5+d/Dcac60LFXMgssciryIP6bau3231p0eW1nCD
aDLCzzbP0kjA9m6egT6zUKvz5P0KLchFWjAjAS9S6q8Jz6vuNlS/cytHCATaGUWG
h3dSBVRTqhrfvZaAgT/wDS8jdCIIOwjMIX91n6CwGoDgvMtuRgXqllCzrr3Sba9a
8o4SbhC+Nq+2NQrHZjbRLz328OHJcaVx5QmtkQHxOGNqGU+OhUO2Z8qWOyoL0SOe
yrw81bBXoFGALSTDmm3aNzKb/EV0Q5GqjnVBbqCSjecltaDzPQFMz3trDHeZFamO
mzynDKFXQ+7UsGym8qyjbE2p4CSyDWAOcHJfoj+LijmWQJLUDg+J1KQElusBY4aD
4kuNQF4d3JOJzxfWajuzK9uPqcdbveur1yWQTH++Eha1vDKN4LJH7ryHg+KDPeVD
YttOGV7VM0ej2Gfiwy6IQ2ByG4H5MtFVR/2DXHI8NJ1z4qM+WQ5VxjruigIb2BAG
HbSqUyx97mH7xSRIZLXLiExGWIoofmUQ7MSeec+vdZDeSUENPD82ybYZZ7k8BmNT
ZvGPiKEPU50J9MIMVxyqPYU5n1/0Hs/fepsZ1tJERIsSHpdkmvnAv8jqUX1/CPQu
yFZZaAqkTkgUQuMrXxCGYenxN7h2BC590A2Nvt31sG0Ho+PDgybuStGMONR/jrAE
2ziztWqNh+3eZtEw/fbTNAfb24epnmCl3pUonPPs5jqr6KQjKYvuVdSVoB1p0kZQ
kBFtLBnn6GOElaoXpIiK/C1YLFwJHkYTOshlugAK1WODIVAPBcOnbvQEQKWCzPg1
pPp1457Xxdw/1Ba+xOj4FsfIAapBFo9dE3Wfl0kgEBO80EhlAkjqfL8BNQlzdK55
P/WSVKPIlLQUETD5LexfJhx/XedxR15vGXJwP2373aau+YglInDHBl/530GDHkyy
VPR4i+utsush7QMABOwgT1YHubhCA3rVy0/tXkLWh0/o58Wwv52LO5Zv5CijROh+
NE6Z1cWdGyUMBXAyZO+GmFmEFgMMImq5H+NC40rDBdZJAIvnxXNufOyo5KYMn4vD
/F3jpYx3Aaq/HLGslkx35ib9k7+fcyRa05CJItOk9FcTIwTM3s+wNR4wlDbcqR9R
tchuMXJKVOPpZbm/tiwwEUGYNOHYQO2ihaGyIcI+5xE0hLB8AzuX2TDVod982xX6
G57+/WwC2KSb2VOIlnNN+yd3OPDGTjDmPNdN1008k2i0Adltl+Ngaqxd7yJT55Mu
7HJSepilFRDduG/kndpHxSJ5uhiPytKWO6bgu8KH3wyegQbwuzETETEWMmUePeOT
PvTjbQOJE0OtNLSGigcnM8fzb8VlcW3Dac49O3mFVLQK0WFZ9TWdQawNEmwP+nid
v+9rPWpb0P/5uY53E6JLQSN3se54ZDT+TWsgW+NvuCg08d1jyQSDkMQJAQEiz3nb
TKMf267I7QNFJgn+k8R6/GbXUMZxdjHsJyP8z55iNYxeCYSzsZ9JLWSMOHtW0qHn
S8ZcpOJsRL2OeKkg1XpFiqY8cVuiQ1OLlwCnO1UdNjYoay+75aTPEDStt0VgDU6F
htb0OG3F4SsqWZ/0SKmVpdZNrepB7y3CUvPU8WUJ7BehwcLy8ajM7crCcWIKEDI5
zxhd2PPCBwjwMeFMnjW65egn+x0MWoXi437gJB+dNn77N7vbVOtVLNzNPHdkI58u
2+lY11Z9pFywk7/un2De9F5MCXVu2dJAtARXtIMQo5wnxr+WdMta5FO56Je58ktN
xle1xT+ek07IZI1XG1+aGtfQ1Q6Huyu7/sQxjNMXnXbEBRs4mYWcnS4B9sSaPaDH
Gh/SSenZytSmanYQnifETQqYYk3Z2INye8GeNglt+iNT2o79KtDE/3VmA/37GcA8
bd3MfzORJoNC1nGjf8F6PbvMZPaey8Ndg6nRNN467tqELG/vuHWOblraKVt06I8s
JH8BZK5unCJdDHXEM0aGDeHIVmQqc1U5wCniLVxKe3qJmUElqkyaodFRpzwrM0su
aq3wqeZ5ojWL1goxe84+b+TwbJckSSH+pJc7H3B8U9lljOHq/d4HUUdPvRBFpXw6
Wt9Hw8Hrj8OOpIvKGgQARbd5QYdY8BE8xVvAwCrMf/6CVZ7a5U/sO6wY1F2lZP7v
BYVdWw3kDCzCwaToAB2rr2du1ZNqQaE2wMKJ56yTOl/wiVbqbeOyc3pGOo6rqWq5
vWvwnmvb7gItmtKf5IfKh3WOUqr5di/OTcZhxC4xkBi7U36XLQrJNXtPrYpLnbUM
ZNSv2xYS9oY0mAY5CRej4rn2OIQKyXlfP74Z/5i/8rO13UBHPo6ljrdE6eZgjn66
UJmNpF6D47ClnXkdSIuqFKvfHF9nhO5iNObvlPps6G7DNPUsjvTaBRs+Aey6rMGo
DUmxXG5lelIFVZ8qLbN39jYToIcRhg+s8/ekU5K+kzTu0J6209tfbKbpnGhtulDs
RH5uG9iev+0vtadLPq35QL9UZeBlL4PXbX5uuu6u7dJEA5blQU9ps1AD4b+qhymC
5DBf8z92qgc93lDy7cz2p/Bh82wfAHbsRqHXyOpdYeh7buEXHd25zTcVKEDMqoyx
KOHf9JecCcQZhwQISL++7VkPDWeMklIiWMT81e3zs9FbC725yMCU5orPug6xMPl3
1Shh0XAAzrkYMayAe3Go0X4JfKrma5ZLGG5fq3w3qwI0A7pN96PCfxv3sjVTNj8a
r7Cc+qYYDCw3A7cIDBQmYQCxWL8qV+dKG7UuJBq9jpqlM3XCMKyW6xJcW0TEbDZ2
onwKBHtzv/TJobbI89hrQqlnzHeh+KVYG48EdiDL6yfpmnrIU0H31fiH0JxzYPTu
NygJaudZbkDtzVUj8oTyLngilT6J3uipDsinmGMXfOvAdfPiR5ErWUrE+FFqmfr6
hcAN7+WnblieXDMswYZBC1sqbd9UhGI/wg4M02loIr3NPH9SyvtsBLCeUyqnz0xC
8Kfe0udxphOtSS/ml6ejf73K8I0/vv4xB+m7/2zuSHpHdOPELqGmmMBn1HfW7c+3
PCdWKK0lHjbyyS4moMrmi3wxkYIF02BxkXawZbHSLIlNGuUk33ncMcmHFPJIVKQL
T4XwJ5Y6nWyAfBns/pVLpJhxAMJXM03UhnVUGxMs1Bu6+ZEqFKHoMRtpL7X7ciI4
JgrPlhRJBElloEtjvjjI0FzaZeHDXr+AuFM07CN0cCXPX7TLYBZ2LOTLZtiWfY7K
EVtwguYhbkmJ4EVNXuQnszmR+shu1eelQKaxAYUg4dtNdA+fZEH7WfFpY3rLVaBx
A7ePwsNl8IlYgQY7LGG3DANao+vy8BCya2cKdTbApZAuQDa7PD6LJI2n6IwRPFCp
/bgcZBSOKHIT5y2ZQByssP139fa7msf6hPqYm+epRgaNzQez2qC3x+uLCX2mFVRf
GNDEHLOuFMzfwuYevdh9sOjA4EeRs70Cl2D9wR91sirJP/qQ19s8pTIPCH7mUo0d
KfQZAZkxaPOsEZiHTft8BJkrrWze6ArLxkZ+jd6Qi75xFZvAz/03O0AsQxZuVoBt
WJRJVJVQTrrG2qu4MQHYmj5GROpRFMAMtykjUzXGf2AjKpZdJiMnqt251w1hqQqj
Wf6uCz/8QwR6XCXxw5ZiWP5QP5AWgcMZZJ8Gt22EZce7OigeDYOczlr1aEA8Nguw
HQC3E7r0NkAngd1n3dvlf5g1zFoSnkfDTPZ97mNxLBSryYxufGNnskH6gwasJv4r
OEoCKN3CMjqwXP2zVOpqgkIT/iLE78TRteiJ9thTm1WtH05zyDx9kLohjffmKGpx
bjobuNYDGsf2ezXj7ApLcTVHvpc013bVpaOyBNIY7J5gvEmDMbH/DnDbpiOO96Bi
nLQx5B9YLxHfWUnUQ7VYGydYm8A9s/ceK70CORdhwXW/7jyFAJhhnsC7q5Z+TARX
6W7wIO2zxemVaJ79FHr9f6PJvt3vWeY78GJTveVZpnc9NwHRRCnqnBbzaTGj2pAY
DJgXimD2WktO2Z/A32tJVm16dZWWSSyCSrAOEGLb6p5blr7K4Sng82XJv9mfFxMF
5T0rWmAB/5jeMra9HYLzIIicimu8PiGRXP+tPf+MDG+jgtlrrqB5PcN/NmTlmnBZ
hE8Lv9OUj0gYE9ochyklmJkfNmrcy+j+mKymLZ/L9S/j5EwOpszMrM8vUgzaHWub
97Mv58OZLjL8MjdKK0hoX60jXF06WZX8i5LinPuP81p9U3o4F7wEBhbr4Agsa80F
zVNYaNnHZdKsyqgjyHCK/Hf/1pQ2copcW6izQpQ9J2ybcDaOWlWXXTvEnr22Risl
Lk4V8TGwX/0nAy5T1Md1hA2LK7C0vJdfqU5UGHk4og0GxkK5lgg+/XCXq3EdpkJt
Gh1aIzvDZDo0bQ4G5NOlXg9VXRh8m5lIC3acmQm8BHbRBh1mDBK3XoM7mv2+2kTE
rNA8GdlH2w2YDl1d0vGECJ4GRjqLZOAZ3cBxJ9FdpdQokr3Tn1DUfsN6cPv844rh
TQPzvIG0sBbt8D8El0YmWjLqKbcIFAE0vYLQpxFquupYyPy0jtPKn119qK5KBHfU
no6p0bffdp29+7fWpNUhD1AD5R/sN3eDhqlB9Rzcl9BesCyOvelCOR4vHiIg9cgx
IvuS8WZRE3vzMgR3tiBSOdauh0gmQaHsEJUjlcvatuDAg7Zg4YXlpmpFmdWnZ9UT
SM9PbPDdo31/lYyHvYGkHKWfkBhqCBBJbdCnhNych5vdo4nRB/La4+6L/W/cWi58
mqjlr8HO7tCMVbw8PhJFCdsmTchyqVxP4G+r85VeypRNQHyM0Ppx+6bAtsJNjbJ3
C/t4RbEpDGdQ5+IdnQzud0ufBOplrBVxSWKgwA3KKIa1Xw0OAS2T5mcY6d5r9vnI
yYwDOqqzc4uZlAo3D1CDG/299YdaNTZRu+2b1zxB2zTpnrMpRBG2nVr7SPBfrZQP
+y0fG+xuaDPQoXLHlu5O27ifb8uwQTABHSprs72KYMmCQlWq2qHF7tgytjTkC8hV
OpEjIrxyukbvqn69SDBAivQrTZeHHt5H7FMnkBxHI5qyvIYWFAYLVjIGJF6ygSNR
VAKSRehPrscbVELEhWz/6FgBTA8WilYRbPtcKizzr4pClQ+GFljkMLj7EkvOkyvZ
HfAb7PgQj+39Lc5eYadaZyV4ehQqzAKOu1Jtam931cV5HPYxcxGZPKFMunEFuhSC
KQ6tAWeT/HkSR28UFNbcMkUbbwzFFNyMBtP6FYsIUuMCwZUwhf7cHGW/VjVFav05
gpf8iAceA7tmk/mKRAig/KTZQS+qgqcqWYt1Zxh/VOOsDUhwo1ILfRI698TuH3J5
7YzYly4GQ2TRIYwE4gG8tQYFXslMowQb0nCtePLcgX6qpKv57dZB4RwMticZOq1Z
C0qeNMTixYn3QGIJcLG3sxZuUItW4SJJYkmAmArBL3gqmigJzfU0Jd+EG7gqpZhG
SOvgsszEaHpXu2YBMBdDEkBvWuEdfoDmz0UvnSOsATPVOtc8ZKwUxV4mpqluBhNA
VDzLAMQbEjhvFDuppHyqn69oGlbRETc4Fe3wMD6uqzmSMLyOzr/3Ev6CraSJldQV
3hh+6DO0plpl5sc+fmKNIopewgXT6R0ulRs5Bc19v4kdeisDj0DedreXohZrNPf+
Imp7RYjD2yuWtygQpegyepwTHlaLpIKSfe3PRIxKsK1AR2Jq5MVaA83Vx8iHdpdW
QhxnacJeQz+4qkXhP254Y2JLGXwp/j7IrBIyVBSjWaKzY+m6MTVGRz+aiI5vJoWA
lHJ/RJyZbn1UPs/mEuG3mp1kheBa5/psFqoyvzat93fHIQ+K5KcU3HP/SU+7oGEQ
l4Of6rDFVW0NSoepRTehSDdhbgCC/MjijyjuiyZUV4KmcAUB79ZpSbwyBdDIbvbj
Noc/ca2wC+Eop7vPAwnReDZkSjiZXcnz3cp8CANr4RTXpHfa19kUZq/cVxWfCU6z
PL1sDKkFt/OCO3hQlKTzVH9o7DBcabukTT5rC/76IiTuPn01e+uTgfb20cJ/s+dT
kXyferqdoka96UeAi3oPbV8rNlmGiF7eN0cuMll9Lr265H+tAy1K4mbAu3QrSsNK
Qe2SsjGvJZk6pVr7FxzsjJD+X/CMwJF4rsYc7ueNNYNGlN2V9cHRVhNIiJjwfpZ3
8SzQqFjw2ZVuFkgMekDRvUs4Quwa0hoLSSqfGRLfsbhtRO2qaib3iLxkagl3BHrp
3yOGW7V3iqa9vaMyPWO3YCvu3Wt+nEwanch+rnPthhC3y9JGUPivxFLWLfRDaFNm
qj3gPWaajWRQpBa+2hHvxPoTOJHnNpjoJj7az4xqtHvAMax3srjlmHWUohLYdJ6F
5LzQrpzujG7vi4SPHwAbo2u3TBjjjbrppxxofAjSvlxxyS4t0W7eH73uvsP65oem
GZLdl0gugcBHzAIgC/t153Fjnu/LZHjqoW2AyBVVHXRCzp0WevwKpvFehGZ2V8ng
O8D8KLUl5zaSJCRFuhwBkFJdXFdazcW/NN0zkKQG713T/XYUzrVT/LvBipnUGtBe
PDYxYGqgP+I9u2JmAVcNzGvZUP5qiWEZoQAJS2m/lM6V5dP4oCFS3Tj8PEmKCmqj
VXXA4uzRZ0ztt0i/XiGrEHNTyecaFqt2E8YO1C/UKvnvzhWGxsnQnaEoEOKSahtB
upXGbp3EIOqIjccK5NPShNNTUO8R+fxkbHPiMqBv3VryheTGMSd6HnDMPq8IOq+/
dsCP7FNT80hQGnPYTSuiczUjn5rOACkWxbV/aeO4drCL08TSzdWXZ0gJ48hSvPIX
hDF8aekjQgcztOeHUeqc8OLgg0YrfmJniayBpQw4i9MVu/rG3Sn7RK1dkM8XpfVZ
RyQlD1vCR5mgU2ea3AzAlRopzfSajakSaQ2w3+bccQTfek5pabE8j3dL4vboQuVf
wu7f3x0DI2xdLODGGdX/IEDhWNvF57x/R3lUWeqo5+X27tWR/dHPyS7AqJV99eYr
unGqx8AOq9kTNog+HaRs0T+w8Dr08Y2mOLYBZJVLalwvljCkvr9cdnMQ7TWil58U
U+jOlCmx22YstI2k77U39qDkM/QLnuosiNIogsNOl235XgfJTLSCmQ7bewsLsbMo
6ILWZCbyIQOKuPidDJK+1uGaNr+WD/IvL+LhOm85J/WklrPdVk+yGm0r0r04c5r1
zkJeBHAXsV63N4lJx5N39S+4zVyH1DtlBFQTj5L/jr4lhA5fcHa3ml+T4l2TN5Tp
IKBel2Q7RFCd1+upP+eNWZoJQins7MJJo/HI47LBzQ8fx4IEG6NM96PoEmXOcKos
dQW3mPEsMaDh9QRYBgIzo4Z66x+7OQxIf8IFHqCw6r1rP7nwxbMoWWpkq2k+9KQK
mPg5avDHt4XxPvZM7qr7r/GwZmKu2oa7ltcKXpveEtwg6EW/TGeQnlYc04gtKCz5
+nJ9WZpAJYOj1Meo7bzZr7mgFq0a3sSao5ChZq19uGimtBuZSRUX522BJYOSjt9P
euJ7w8CvCYFWfpoQDtv3fqLz5ftqxXa5HjeCZLlo4wB8BNIAiHqdQyqeHUuHi4JG
yOy0OM9nDvccOsY3CEWHuZaxc3a6Q2YEkNT+LCMEQtNlO0xIr/f6s+98gkaykREG
jEJarIfwK4pqEwyFs85Mc9HtkKsXc3+DXZWIYYdEb/evZeNJo+ex6yCqH2wDm9tt
cdCGcQAEJ3odGGCRFy4Zp8cUW4m90ZucRAzI2ybFaiTiEpgxZQW5EfMkMTFRuA94
6selTi2W5IJ3NVKY65p0qwdioaT2WGsFDIK/OKXaXL2DPTbRyk4BXMRl5D6FN2UE
9soV9kFdxpFn2hUqbvvHuYBytShpdDSnjiPYZlYdruIh7Gkn/WNeNTpVbeCyCdVh
STONwaYLXFQqfej4WAKE7jFrIj5vyxOWf8bghavqrTje9ONlNVc+HDHo4us4+mDd
X39oQF6JxHCnq78XHRTXZyn/Uf5qJ2XLEE1kX7trN9p+9GvELQIpyyBCgWKxLit7
Nckhn0OIWRCeYPELrpER9HsTksvW67u60z9S7phljR250BS3lMfavy3eDAOHS3A6
+v5jYUdW08SHUWzIRUP3g4LA0aW4KNCiWXUmgPnIzpnzCD8bepkNDzErUMpYo8YO
+TN/D4TbRftrWsft3xw0ji+GpRsKhNEbXNaMiwfKPVXcFqRR9BSTi6jzfgaQnDqa
LI6dQEb+difOosxqyF0AfT1MDQOLKiLVyxk/7dePcTaD6iym0mlbCqb6UqBn/J7d
1Rc9BiiRzz1EMawkQ1mY7nAJBXdPTMFXl3p7q3jPbHNUm9G3Mx2nKOxPhgC70njy
z30JuVCoOVaywUP8I2PqkDWIoD7dbSixi+h9KjRKeODk72Kv6BoToiKJcC7rXkLJ
quygQ+qyjrILjpPR56tMfw3xSRJotCarx4WfJz2zMxyYhm7AcfIChIBoi35V86cc
zvJZ9WaVJZA5sAPn7UAzqDTNx1+rFXQ1npp67VqFlbOH2hYW7m+cQ5eaOqd0Xmcq
ZKTVKkJtBvLROuJnrpisJqMIUb3YLwU4Y8UxrCw0YlMSYHR/pDtOKlEpWgie+2Wi
jolKVbqhR4CM3AgMUUTBG6wdDYF0A7/pACmc7UJJpkcbCbzvRv9RH7oDY/tZySbZ
otBepEvUQsnKjTcuSaIMa4UtpJJWtXdF3fs76Loj4mnuXIEwIKRxRM1aE7R+NEze
x9iYPU1wK6pdTT0PFFJxQwfhxUDpfZiUouUwDSJriCGCC4ORp1vPVn+a8QALOODw
/7JhWE9bwx0CROHoywwCU4lve+cOseSStDp830YW2Ihe/TH1iprJ5B6J70uSZI4q
BC0me7keWUtFpCheFX1cYxj//Vq/bgO6SQSNpb+ngu/XDiRvqgzUQDj02ThBEE9g
2L0wv6c+Tc4dsa/Gm3vrofLyAgPDOFxBViNJr/Lwl53ElQfRK30fys0Nusp3KQsP
5bR0oznkjQYydA7vzc/dM5Hx9/1wMhLv8mu6k7mDHXrgURyOrpoNI8tWGlDU9nvi
iJ9l3R2fJESsSpOK2I+q0Kz1Q0/S+e36Pb79If+uyGvz1tmBwaaCDlosMDbth9UB
oaBpMyK4Kgy89FGOtIXziM0ETJYqow+w6aQCa1Sp7lSdceZ+Ftb0HZTPC5/BkUeI
PVmuV/TMCzwxpWmrkmjgHD32FESZ27EQx+kwK1ExcKeK/Ghj1UJGhObGtqBtlU55
sXUy82ChW1uf/spxuv65pFsiZOTYaFVazO1V0rJipLMNhDAA8CGGZPrjGKNjiFv2
oj1AGo5fBtCNeRDf6d3DcUwKsvjzxJT6ddnuuY4j2g4PhX+Y/kKk/k8RNe7OyS4V
vwLP53XLgIJrEOCmhLtfIumPkmZpHmjt7MPyAfBg8m3r1imnXwBfwpfPTDwQa9rf
NeT1hkO+fmGYmZuKh5eG4zlyhaunh8QR27jYNP8sy4pnllf30dmKR453ge/UL0ci
NlTU7ZNv+/fN9sMrAYUQNB2ccp9vqguBhy/jML/yo7gixOxkuAc8k+FZVO/pZMUK
x7b02Un1SAarrIDrn39SPuJYBPzVZp70Ze7w9w3Yb5il0R7EbVfiGpITzumtU48V
zKjEZl3KZQQ/uzUyi3+VXq19VoeBWIxi7Nft5cvQrQxbAGam0LQlpanio3/w4Vd2
YP7K6ItBqrVEuQ3FELy3Zbx0h3jFrC/9gPbMIiaGKAXSoVnJVzKVoVl69N9pqumP
nZu2QJ7ENE0+jBNGoC2Eat9xvNTCmopcMixo6l4QVmA1JHLjiKIRPjKM0bHh9MqY
5qDE3zsf7tkjYxW2b1FQERRgjHQZSxU+hMNMU5NR32QvXtTnv7TtYQBPw9o+hfku
R1f6jDkXRaktqTIpoMNip9GE1yJj8SEcNRp4WN4Y6poNqsqz2rTGAIJYB7kZkYVT
ex8wRhb0DuV0wWoTob0Xp96VpFMwVHUD3yRmw7D3Fs1MOwAgXyCxuQU0/Hj9QwS5
PaRlxwpjxgSlDZvfmJETA9SIIkOGNoqao/ZN7dGCmDLm7oCGKsP8dWRDwrFfVVZ2
aylgoL6RFU3d7M39RL45AKfsUf7clP1JQtYaE43G/N1y0vIAHE11rW5fkt18A9Z6
BsVmKhIsgHMsMAlJWraYdtnVfhJY94iPPbxQ68YUO83XcQmvZE6yJvUflJkiT4Xy
mCJ1Omn7JT/jeWKJ9XO/eTQo0iB6sUFrmqEVxG6MCZSkLmcCebnHNWrIWPQJJfvz
mJ7jtacTBn5JwAgeboXvItD2k29t5LyOaa0z66+HFzvvWWLLgtPO5m1w8X6j1cRT
EZDZ+C1dT9QgvjYKmHzE1mD3mqee+91WGBkJ3SuSzLMv6aVIosHQ+1SAAVHGG10z
KnNBK+lb/0B8NFIEtlizaa+5lfj0hQJfFd7BA6wWKnc5OODcn1eJR0ymCUdieiEb
/w4lyGs90bI0H6Oe/W0ipDHRtDp+CYNGlAdF/47tiSBu+lUTgHt4LAKRMkXshU8+
Tygvj7ujCsLNk6cTPOwQbZtOVoQ3vYE4ifQGbdidqQJWTj84DknCfGdeCDVeHih6
Wl8RNhDcbmE1/8szSjvWkfV7r/L/iA3eI/X1NOqt01Mva8M8ftn01wIwKc/zEnz2
heFjpogyfrZkqCYL9XzAn6ZBJcc1Ow/v/prP9NAgniuAORSWw7yXJUEya0/07Xxw
e8skUPUdMmkc77jCLnMhOPTarte8BT/RhDDALauCflWkkDS69QdtWrfg8Ma2U1Mx
fhVYS2M09UYmAzjq1tqhT2G6HQEtaIJ+IQngd1h+Rq1BGUPfI6XviY5MSTnCb4HL
mVbEdaTN/GK1bffEgT14NIaxY3/sR1RSvar4uWYGI4bDyPavNGPz2plgvqZ01NKG
B+Qy22D/mOq0ffWP5slJbRobPoJxgxH8dMyawneNaIow1jsHyBRn/Ckc87U1swDB
ko5QYwqxLhqLRLmmeeKjvfxZ95YvYG4GTUge0VhrUM9+DXLT1IqmewlxUJJ1syyy
oWQQdsQDgsdtt7MNCgCakHF82FXiW/iZvLgotQ2rrVK8Q0Jfgy7F/MqHNbBSpRwV
tXJRf8rvq4uMEt7MAMTA2nHrMMTB5vGOWKv71OQ152lK6QSdwd+OQ01QMiPxwmfa
EddIQaEWpxd0LbeVNyQU17Yq0Z+6Mo2pCbrNFq6WHC5tWr/0EoCu6ml76WY7Ih9g
czVoKP9Zd0rNCw52/wyKNk2QNp16mV7Iru1S9JhlSfW2SIfkqPX46IhOaqFgpr2H
IFY1TC7u/o2ChWWpLP/voay8ZyMzR8WheJ86klODzHAuJpggO0h1ALpzKJX2RKfN
cRfMiYbSESwY2pd71qzb79TperaT3oaP4GU5bCDtZxShl7IVQjKsoLnhz5LIOd5P
7moEZz8YPRMECBCD+sgVQUv9e9s/20OGOFcGy13qGkUA34TnlQsJxykaR18ECZbx
8YE2BIyXF8KH/dvmdewpVkT/r/1GAlUFwPxQNIUKO+p8AOo2u7vP13WuAKFz5qjh
kLoWrs94HxD8BrMILKk6bzbT+YxtbQJJAcWLmeA1wbP5WazmGTrX2YYrpSzYk733
ZjoIAO3nbC/+S4BZwPdOL2BuIRTHQDzFyZOhKQoql0idprU0XLYOPAhnXEPpfS/P
dOun/72+AwYikOZ1AmSQPoFZNn2JE7rfiWnpgEMl9EGqeMu+HlHYknKyx6exyZ/r
AcvsOAcjXmNulhSmHiNCJLmlFS+l+L0HwXH2fYL9fEBLZ7BBuaQ/hj6cGFxOya23
KuckFEAUKhz0GrZzIYd/Ax6CzeZXzmDuzFFoYgo6AlZ36Wc2jlYznJr/Bn5y5Ns0
95O0D4ER3yCuGIlqBdSHHFSMxKhH/PqtzbImpFEEoTBYKlNZiwbQgEqT/6gDa+qQ
6A9nbaZ+PHYvPEidwLKy8r0ADJtV4MtkffWXgxBryVi0ItmKKQBaWOXlnk8mYZMo
vt8JKjzSxyq4MDpmkFg6xfumM6znjorsNG+s3eSq89wJ/DjERsPg400clgpf3/iT
TlSFCl3xq4v3f2CAbh9+om5l9H3EAWdnPcLAZapD9Gc/8Tk7vaw3vExW6SkySZ1j
BvY5DHIuJf4QWHHT+s2gKofbvAL0Qi3dZzr3XIREvbaL/0YouQD8nIJaSyuA758A
7Ffxp6DlyxF8tGOdR8/tQi2dhEC1e8CLrriPvvFUyaq4hfhYbVW7xaloNN+1CUTr
HPSG+sV3UUtgPczJV+KrG8Qgmv6lMvz2kVU9zmmjzPSsHexwan7y1Nz/cy3rImPd
m2Q4KEHvYfqJIbTYLTe3y2aS20Xx966lYHm1eSvA7yMbcQgwzS8F4z9Bj42RlTnO
B0rGN6ZpV4yV5bD1jpt+HXl79GIp5UHFR5YHOYzVNR3L+MEWW2PV2VHGjE3Tjvmw
q0CaslaLn4hOUSyYYUSZ21b/oF4mDFIupRoaS34lqkUsMr3gF+C1bX0MdSgOmGfz
ubK1rihL0qrg8NnCB1axGOjQYgQZsDHazIy9Qey8PGXLKXEcq6dh4Zy9cF5TJ0qF
CpYN/quwcl2PbMnNI6mtg1b58AjCQx67dRtOPY7wCNM3Vo1+c8CxJ6LUNHVHg0eq
4S4wUXPPBQb+prZQGVMle0tMmrwYROUDz/wPZTqH8JCzFoxlauFDx4ojuq19htFi
b4sd6TkqEyAy4PE0VIlUxiG/oQQxnozqbJqjsOkUbU8sez2XpQ9wiEykzJ5PwkYZ
XBuTPmSIBUTq4awIfG3copuaxocKeRmkR/cjOml5hK+p0ukMIjqNw91ez3uxl4x+
qDyg+OPsEZVmBzV4OYpm8HmaBqjalsSqVmWESkjTQrvmYsD/X0i8Jq3fsNff8V/4
RlNsuPiXKjQP6XOHjWqNyYsj3NCYATGEBddMhxq7NrLrOc+nUK5jGT21tZ+Ltb4y
Sg8BZEkrIR/g8ympwXmXpgIkgzdEBjOFqYcq+MSpPA3f1Dvd50l7J95/w59RMq29
TiCFE+PG7OJ+G5YminMY1A0n2Ic4nXDFMpgH+keA7zhl4cPlQkOEKYLMIU1Bk/pI
AvQwjRWukYfLJOTYoW4A1g9HTJVXtC56WgOkYOcIk9j9C9pXMhNuAvK7hE/x6868
PTP2xQZ/5HeB+htusMTN2sULeDT44HBFNNZUlsjGIe96y1GQ2WJFNWRKUeB6h/4C
Yosx8JErcVOt9bSLY1HGj91bDLaZFvKO7mUgp2nWALTBB1rfIyUhLa2xOHc7HW0f
2cArZAN8UvC+rGFcha7JHGG4CLQTBDEhUCBfwM6WYiFF0FvejNMyy9j3ClfYi/8X
IJC7NJMpZm+Y8tUfAW3NScWBDojWC2msfqn+52LJhvL0+s6Ci0N1nR1ajGo5rWss
aut45v9NPoRKKz9xBmQLPtGRxfyUJdVeZstAEe8SeUE2t9LZiz0sbNGv/XQ3Y0yQ
QV0t0xVDzUGhByPsrjU2LhlsN1fVoevX7GWGhxUhV6mcbDZIu9fSR5Vu9dEnI3WX
UjTEaO4rnNs3fBMjejYFQaXIdJF5fHWEh16Lvt2ugOmdSk5+1kr4G4x1PJ7gaem/
MbUf2MaWQtOB1l7KCU4VudThticIt+nXv1pPYQGNZwglqdAUJt56hDuF25IOcfYS
I8YJV7Ql4UvBvEZjI99xBXbIcMXWWmGTV11UTZkjNB5rd7AnV6mHRIiEcyube3Mf
L/81r2/qwhPY+9qH5RDjjJ6a9HwqPBKo2qOcR+yN8E6yczEAdmvWrBCqbWkgOAmP
AJR2cvsE/dsxP65+BtLFo50pyRrUfhHbQMOsohSOz++vPdbH0Fbe8sLLwTggCFM3
8lieXT+LCmsE4SS1jnckOiekF4nWL13GUC3/6Il9xthMVIqBms4idPujOps/CzdO
s7yUb1el19+5hHTzNosUf7NQs58VmmT3msqqMxh/MoRLYh9xkNDqyrgPMiYZcoXG
iHC2P7zZ8zmXk2LiGU42G7gf0xLwhmDHxnbPJ4K5gQV81xdckIbDDUcuAgWaCFsl
79WVE2U/oqyPBKZAjmcO5DyQMpq9lbFVJr4njTxbONLq3JcbkWoPnsXx4OTvzaJi
b4agxoxvd/fQ97nKeT6ZoEoMrtgjnSQ1wQ9ZJr/EmiDxTcO6gPkBkZUcHO6Nc54j
B9/xu17GnTVuHQJA+RKkxkmj7bP1w5pdkzHqDFM1uwPFc3qBIps0M5SjOzDOwRdw
VLKm1Q3qMPhq77R0y7C450pjQoz/NK1dTgXKDXg33OrJ8hvHl1xukiN/Mjsu8sqc
UDIyIq8v9TYRn0lHLfsKs+6ZWv+tURbnSk7wbLDu0SxIfxeyPx6toc5bOgDspZXC
ygCk3ABfgxvxmJ2cfXMEwbtMPrxAi8BHu66Pvv8PvBdDjntXaYSQxmWTbPvyd6H8
c/X66AoYUpjURKNjx+CNfJpr/yoffvfSmK/0NjiecTB73pncYbQm276zAN+YhiEx
aOBiwXVFiH0XCcn0LiQ+rGXe6/e/Ay69Itnx/vHtTMwqy68G7rX6Vj+z9jqOPq7S
qzZfPtsslcnDf2b6viYs+ngbFKsYxyjUIDRLl13PIKeAlOxRFle03ncaFbVfRjxv
nvXLrBZdB76HfrRdVkaint8iqainu7TYLc+iwbi6nfTbH2tLki43BEcuD6TmMoaM
m8r3HJbQOLzPoL6cfCWbEyKp5L6gdkJyRxR/fSswmgHPWfgs4swCtZMUYT6ljQxu
G1myhsFOL+mUuO+DcQND+1R0MSy71YHk7NlHPHS5DCgoGM6q0by9XTdYPlVoP1b6
P1coii0EeP2Ynr8E1KYYxAXOwg6azloZPxsJKMbDL4UxJyLlJngpfZOrDx3U2jv/
cp/c1jSjMks76HLNyBiSUqZL5qfklRyk+Jc2pw3PviLUFE6iLK6OrRocr0yFWPnh
PHFI1hgft20k+hlcx/yel/niqB3eCbos/axd6a9umCBx74AfFD1a2m5jOpgJvxIC
JiBc1uQKVwNn3aq89riBLKwWqSg1WHR3VO+H/4F0qlTazPpy2jQhTY7O0Vjsbrp+
c6IVq4KF+8rieO2/X5+hElVFkNOM6eQQNj/qT3dbqf33MTCkcS9rYJWr41h+JgEs
aL91Yssyyq1hCDb3Z7jThHazGwyVBt3u5xLXnY6ITcFlCIRTdMsqemwLlZ4PCUCa
TQyg6N1HOZgrrNhp2a7ucvRraBSNgMMN89Is/bRSqFg0uvNIN8+ROU8Ih9k3mqGq
x9y1+pBxrfuYuuWOed5Y3zYUf4eJEUazPDj/zCow5K2xDAyXj0CHzpXRNFbS3Wto
N9jNBqRhIQ+VhLNvmnWGqahpSVyMSL0oF/cpBWkPVeWpc+RnY9hu5vLkpZfX+l5i
NTGz6T8H9sbaP896UVF9xeMVVMnw71l7NcRwu91ogRK6fZ6nPIGx/1nrSWcZm5TN
g7tbYbgopjo5mDh7hSbVmv9HQJCEM/wTb3hSYG81wDcxHxBx0p+4J/0+RzM88ah5
HIu4D6s01CSlQ2blKBIRS/aKDAaR7md9RU50RfAaoYIX2BFd+TLKWTWD7JjdSVpZ
SVOv0kKBPidG1yFvW8EClC1T4uQtW8XM+GwVyWIgAy+CwRT+61tpl/nrFea8Vvmt
22jr1EwMEYGWcizQMh6bKy5VQQuDanuv68Y5miSJ1IE8zxq90XCmXNQQH3vvQQtv
AHr5jBqwJ8uxL9gXPad7mW+7400ygvOZVG+FTkrV6ALCtH87fMwrjGOoJQ5Knrni
O/mYNrYA9a+HXmsUjuQIa87tm85u+Z08HxdX8zLLAV2BuLQk+As6T4pC5pFOjWZj
q5oz1OIMb6vdQrDtCiC8HRscAJmLFPPIGgA6TrOrGwTQb2cRnSUQDDcrrvWerCCu
GlaVLIUO4NDEw0E0Gmxz6fX16VmfpTUWWDbh5ThpvQcMB5UMOiF1aIzxKgHFmGge
kyK08g7IvKY98p9w3YNi+VsGZ4rgwOmdVfFeDpWvdOEUtnlkjk8vm5BLPg1s4EJW
4BEIJgUfZOk1SUw8dbFiIm48lcvGtIjo9iJJyIfidMezXXlZr9FZrwuzJeYr51RK
n6X5F1oFdiAzeV6eFD2NXT7VdrO025o1c7YbkKPIEwDtIS3N4FjeA7ehG0T1RUvC
wUmMLp7XemMF6IWqdO6hPbHm9O0dlJojdjXNzsNPucOFqGGrbKyforZ06N9i0DPk
jHdTkxpdYoJEwOhsx+VMyInKyQAIF3w9JppEHKACT9pjkgBBkMppoM2p6tl9RHVe
ysIt/EGg0SpgEC/xhMBJ070LLgd2mlUTt3QPOS7swqqHj19N7Q0HkV0Asrz7sRst
VSc+oClZZEs117Zx+hNS0VQYO5RDI4Rcpv8gejcQfJFSLrafneJNXTQi6b0ItRaa
mNIncw5N3b5LlZJCj4g8BTRyO3CEtU/RV85D0pNhkSdLafUOZZ8xKS0+UiCfGC8T
y1rs+B8qtl9nEkNOWPc8WCNNr4UoY6/JTzGt7jEEGruvUKG9uEk1PnequnyUViqE
3WRQpG9PV9Sct67TSUyAgx1pCQ9R7TnGOZji/jutUmU6en5V8VYrbl8wp5zIoTf3
pNgW8LvENWSqa+MJ/4xaq33gyb5CmHpr5vsjff7Ag+HbcsY05w0v+ORvfD/vASm9
14y5kkZhVZq6HYHQtD24825opJ/+71aY6A9Em45oAKoHxYrZY9iPL78/QQCzBHmG
e5MdMu4IP5D9qBhbVyunxdS2E5I4u2+Pn/YeiiU4yf4YBpjQ05k9xLqZGc/YwhEv
N03nI4AjYyL6h+0qPIPUfhB3hLtzThVIQoA7I9PQ/9ElR9MwqMz3OdntxvT+NRea
MBj6hHYI99JYHOv3F1aV610TugHxdH7bjIUggvlZqZEHP6YBDYW1FB0voZ5T+Frw
2nI+9LahEu7uKZzBK1VAGKGJIs6caxTfJXcdZS8gu8CQ2IyzlN5TdC/N6OsuGmOA
sw4jFeOkCW2jaOJdAPBhd1b8Z+bQdg+bVrNs62WikErtq/jQc1DV9MkY0PYxxEEY
ovVzslkawd2o5kICHQPNXXLcGsvMiXDaSHpzZWcFul/ju3G4lkdXlZFBnf71uZ8H
HWQx4MdoyrW4OIbBTOQPcgaF0XZeJWPXATNIibHdgQi5tXMWHY6ZHoV7WnJV3VW5
WwB1FLpsk51E94J6UyJ7I1gZ7DX9xsU48yg6I6YebCY2Hm0/l5zKhZ1/BiDshtfh
77HX/RoJ15G3/Unn7YNXxkTGTQSiIKtzA57wCZG5qRwxorzwAi9scGl446P1gNRm
6uJmHEj8zRouFKwSNoAr0sfKSO1kG+tycEu5XDVEUblTnvNCON/dyn7PjSxovagD
WlBdUNHNPcL4ENEzDmMTQ01io7bkM3nyRXt2w1B2MLnHGUzQqf3gYMk5X7A5cWlH
vfMXx8NX3XqhFvsl6j3PdPR00FBDBZgd2fiFi32n7IeKLUidKoNc9W7xlIHX9HKL
a9I/x0X4V4Y7koyg6vpOIhHaw2eJdTYCfjaKND1J72e+fJFapwjif3uPnqDWntj+
kk+y7id8m8BMBIXakKMUJID+LZrwjShsHWdYqbvEOjhTdmNnoBm3Aleo1VjUCAJM
u02LyGtiRiFBI34qnVpjfrVS65u1k+j7rnM3bzgRhBX6UwaHeSGLjP7geywqw4bX
1pPLe/icmC/QWuJJXEnCf6xjKLkRvRQJrAgAAhDHz62ZKolwu3e33MS1s9BrDDsj
d5zfLRpuBcgNabj/b5XKH/TYYvcn1esssnzsFHnnz6K9g4aK0Z7Zbt4fOsiQad6t
F7ZBkdANsnIox0njMN1GSus5fNPeX21IY+kfGZVqagmkvdgSW0SHocc5TxywDpNN
JBnyEI7xS5C1LXupKACtAkKSB4Pfrbwt056QF2PBVJSToRlTUiMOIHRKEifcZnow
HTjc8kNhiHTtOY7jtt0SwRezjKDdHpsGgS5H60U6cQAOvMs4cU+2c5aY/TJ7rpgr
qZIPYSZo/beWnWbbWPlpi0S+iEH9E3fJy7VZ7f6czS/tIb21pY+BM7zQqfw5Ax2P
l4Q7oAEf/y21hoahBMjjyuaaSZl17PP8QG4s2kxHrU/HZ2tkuBP4MKFmIJ5KLBJ+
qItMDEJ9AU3oEly6BNGkoFlVn6Gy5xyUawsI99XkByAzboP8SweMYU8Ms+8x5xgR
ZGZUCwJhTG0dbR4UGWPQx+X+DiqG2IeeJ++OiYUErc1yEBxHKQTrJPK4rHuG2659
d69Xpx5b9ajCZtcpo2gMj5h8ZYKhBz/9ZTajKHIC1j0/y9AytWqR8Glbcq85hYxh
NeIVi7AWrKa5z68URUKXCTkjD2wQEamXjso9aTkAUZA6FlWwlcxGU1ISOPz42Yc9
G/6XFAd0Bg7lm5+VpKhY73pZIazGRWX090bAygHZ0QeA9SbrKVr3hzGHLj/Rn990
yr0JQRq0qj6IhwIGd2CqOf6dPpYDXRimYD31lAGEHRvKOZGwiSJ8F9zENNyFqs7D
yT+X3Hfq3ZtWRye/lhCSr5gSlTX6Dzcz3AXwhL69bzdunPQM5aI6FWNQWlwjWE4A
F/I3DJ8ICfsMM7BwVOdqBx1CAGzKHcORsvI1K6JFPO9mlum9Oye9u+plZEmgUqaM
jWMCvGLxm9GqBftEaMCw7Wd4tMjZ0wFJdoSIVJV9fQ597p82lRvtfHeryljdD++d
Unen1IT0pfu1SaPtHnGkdYsyB+K/KHCXgYprgywgpoamxy7HogbludMlpUMFvmFx
zdHhXhwoNDIGwWk7iRUVNEXP0S4NvDH/zFHKAlHR+tvdhoJcVIG+Nu57xZ4l1snM
rhijRVn6/lxSN1UA4CO6lPf4aXVbY/MRfWcB2GfDvWBlX0yLBQSNgYGwCz5N/9tE
9N4Bc9HamPxjxCCVcOqTjYCgHqtAQtozBWJAkSEKBPfb6OzMRLDO34UsywGhynxo
WRYIQ8eI+5fqqFv68iY4eMs2nF9borfU32e6Y2mTJzwQ9s64Rf5mFi/VZq1DtQdT
paLOlsOBh36nIyhM1ShkByAr78OVzPcXO0ICTc0R3tEIXHoGcXYWD3wUmp8V6gQW
odlvMo5W+4gsOLSZu9v9v5NRmKffUYdvjPqEmEy0KGR9J8HZQAZL4AzGXC0A1iq6
fGxWeKqrnOlsYCBdkU3PCTBdAma7729rkZf32q+A4YgK74wbVkEWMyoyQ25xKBqW
koXDNXDT5L5anEy8s1N7Fs7y5S9krT0la9x0mOB7Ql9rF7MS6RxYG2DwH1qFpuH3
6WgCo6fXCprhz8p80K58+mDzCI9EgrbpOtJACwxdKKockrPuZ4yAg17Di1zZH9bq
TDeHYPRqUGDe/SbpShCq8Luxo6RRR8mez8kNF+lnU04EVVzgYtqjGhcor8DEKlIv
Ayt6Xm2oLPLtCvCLOkz5zr8NjIGP6N9S2WXg3ioEkMaAaKYSpxgIso6/R8hAGuZb
SGfkqq6aR9J4mGaaeBk1VnjuTXNGkp7JR7WZNbTRX3swvlQLp+5tnzQSBT+r44L+
OMp6w2V4qVMjsVh458wEw3aabKuvLE3Hi52Ec90fIvcWJ4tkiOPVoU13N5oSPqST
zbY/7UlPswIhXCMVoLs1IwnDBaMr39Iot70almfk2Rsk6QdrKvyF+1mVCaahXANZ
KrSHw4JtGlGM3hLCHWZJjViG4fc3yMAncv/58WyQNFzMCMh01FguoGjPFDvYYT+w
e8B8MgtVinpxNxpU0CQNF9s8QMpnc2wJYVi5ksAUcroDM99loKeSUw2/+akuuZyw
/fcwEknEgUQXQb1Vvh3aFNAq/HZVnxApzCkWM1RNqqofQc3QkKhcZRafxHT4pwpm
sf/Kbmg+zzqhl9tpsaLxQD/EPXJMY/66upE/nYC663bAwFPDWY25P2Fv9MxvmJWs
n2uZjUaGpNqv4MZXqWOtZG0GPSMS5AScMgoW90D4iiS4yRXM+dR3UcV4SFfiyf95
BHfRCodKR9vksUFGTO5OnXRDOs1sXWW4PBPZd8c8+ax/f6yg9AIQ/XjyMVpAUqy6
/mKP66adUdOQa/MAjSykKs8xy5r3ToIFPEwXUqyyMS00L3awYvD5iBF6ZMYOIt7s
mikr6+N2K/nP007NGr2+i8b5esapXsCMsNvC51Kaiv1JkPKjBBbCnP03V5Kl/vh+
wEwNboXTL/0LZ1hPcJACKbtT24ZbZ0/bShUIToIQO1a9I4UmrssSt2y/ItdVbA59
kJk7/IsCHTpSxlfwaNU/nx+SJC5qkrjS5AZT820b0ly+/6xx4ZD+VjVIJC3XoEb5
Mf3chE3CMeZNujyd0TT+SVls0y4kx7dXqcuyY59QDbml9bEiooIlP42rqKmlstyf
tz0UDDSFlPD2YgzgX/L8jOcZT1EbI0Q1D21Yb/0ydiEeyFaokE38ijgWVjDGMAia
H6Wbyk9gXQDaDKn76N7WzlJyzBdEg10+LJYRcoiUAz8Bxo5ScG2zep0oXdjIj1c4
h4YGrnAFXb5ZvbcB+JSmNN2JFYOqV5AbHphx40k5wUxRqrGxJebVvtZ7nr3zFRYH
KsINedZtxml07ugXj03bC9GP45Z0K/Z2pik6jnHSvjr8Ls5s0kDWyQF5MNIiwkad
U5tzdwr9+VuM8OUx6xmFPghigG3FuuHz5ksw1q//7b7lxvGSnaR99JsXX2ou94Q2
5u3wP3hyN05HEbgLAS1y4tV6xTy09u4BGkGhIlD7qULevFrrRRDFyyLs+KHUmWr/
ZOTwTHvECTxlL6TIqz6V0ehI9gL+wTZPVPET9bQd7gXcTTg7YX4zcLU72rxZAIaG
VxRo9PCtwzIErluxk+Q5ri5tLGnJFjwolZNFBTuVeRFOHLVKaOMC/V4tsJZKDvEm
tcAbAMHCuB/BxA1WajBi+0nqD7V2AVR78a1bBD7vWQu8oqLfwDmzgIv8eWvoq5/o
b8YCiYyBab8y1RdO2VtTrmTBXAaTuLS1n1FTaCUMIGrKIEtYI1mAMRPCQprZkffv
WfVHvB4KiBkNWEpDWii5NLTyfsJ5DW/cwr4Q9mPoYQDfdheoafH7TvXaa1vK+A4l
+bn6XghqwE++kDjeqIGarb8o4/IuQWXafKkWWjJe8+lSSOpKwuZdOSNosOZ5vINh
JHmR/JUUo9PTMzVnu0sQNo6GdXW5699Ex6I6d4w8HEoIepwapFb1ddTXr5abJf5b
KJFIyvVy0A+2/wgyFAJUR0nFU6nMQRxNpq30z3omjrbFGpJ+XCEaiYqCDKEZqCUo
N0L/ooPG4njLlY6yn2MdizVGaaJeoNwtUXVH5UxNAwW++KCo2ywAmXD8ol7PkUeo
Uzu1WXIA5tbbIKcrtn9cLHjSNi9cbmkn7Oc3MyKKv/zPxgTxzrj2zTpsazIuI/Bw
42s5XpN7yzJyeoyU8KKfn8RfJ0+6tDSUkkaFsPyZwkHujRxXyTk+/dkZYNh7JYAb
JsGVGslyq5VS/7WaoRtM1zAVau5qAogzknmXvy3oPiWuB8YfzK4PSM08oSgu2urW
6jjYReQ+tMeWpqZ4Y0toqkQru663gNiY0rt+PqkDGltkeuwvQiiBs9wcFxcFPI6O
KwMEvHY8rL+iJ+Rm+WLWHYkxgWw/dXDzqcoMUen2BLQW30XeYs+9OpieuVT8Wv4w
C6hAnvqLQoFSq9VXvp4CKqjuruUGyq0M73JHwHCDQsDn5KrP7ZJbCUwGGeoscAIT
aQGxoua1PvFLbfOhz1V2nJ2Y0oBWq0U+3E/RmpqtAljxXLcxSPK9Ter3rDrthiq9
d3TRux4fHb9AHWVDCwWbN69AakAqHb5HVLCudO+l4zuVXN6t5XDBmD7GAONM50q9
elXM8LvIyEmaiozcGZROz/epDCld1zcl2QiIiArKybNbiIaXV0x0srdCcSCGJ1El
AcB/ZK1Rv7qPD3MS8vj4uuD5E8z0mSx7FKEmnQ10IexQ2clWkLY7Jl8V4OlGjh6K
lFrMb+zM40Bqz6c783vhiRFrW6gAsRoNdoOxmJNgJupGKdTYdkSZkXYbvY6x5Jrb
kg9Ow+7L7YdbguQ8bPbjJekB+mW8ozsQ81kPTKLIkaNk1VmqexC9Ch9Wkrl7Nmkb
yKPVnxDzAQKAJE724CK4WSur4YIjpcsZ6DvAGzmP1xFEUPOnL3g0w5YbTnXdgk8/
zOe6MXYn8fL2SLIsFLpavFIa3egDQLeCfmn2Ol0wnO75OjO42fYM69OcMm3oS1sJ
1L9adE0OUudwq2RZNo6sjBuy4BbqCpb12myFAyrSJ4HKNjvrMIzah/F3VGl0UIeb
SPHKWg36u+ESAHaNb/IQsnkFhH43xJvfSixpp82UAt4i3stYsvjcrIRLdNvYIbC8
RpffUHis+16VuoLYdXLCcZOmiZ6jveZMADnmSI5AcLbznCNdTTZQXK8wNDuDDw+H
uy4LaRqhl/Gf4ftXFvWytcIqxKBiBeU76j6Qm3YSSb0Edzka12K6C7FbZwop0U4V
cQYHbLtfucTujeP1xhHo1UvCms/0YWAkzWeQAkGKisOxamCkELG/CE0sEa5fcCSX
ovaDhIsyVsN5h0z4g8obm6NPf7eXZ//kY/lbJt74WBil/Uz+g1TpTVIgabHycQ5b
vheCygfnUfoJ21KPVSqqfmlgFMIyqFX5Yh3z4I3IL80Rrx2IPVisA6LJBoRJ7PPK
tMQg2HZrAagnsM6+AyPuOwV96nrunKF0ahcZWeOSywYAnTbvnirX5WdJ3M/v4Nao
xGg9JjswUOXEcqXs92D7Uaurt7J2k0Sos2539ZJQ8+JMF2lFHpIfx/aM2m9bh2QL
lZQnxNFMR7Q+FK2koho9rSukzQUGaoSCBPNnMriUCaBzaPboklWzwhgZ1Jtra3g+
dHEon4jsni/xmzPxP5O/ahG5+dArSKTq2nc6l3VZLR0/KPmUOa5S5yYAn57HtAsX
Zn7xBGZxOnD0rAqYTZFsTgNV7ywQTJCyaOl5sp8SnwIWQOfNfQ98Mh1+/oEcZl+r
gXFlEMSxTKV+liFVqbVucn6BIuQSZscOQN1DOqBq6cun8SvbEuvpx9E/rtmn1RFf
oNrMkz+4I/3kROKWUQY7Lw5lMp6zx+SgXRWf+5XdyL/SlYXDRxUED/tQiP7aA2dl
w6XWjdqx5VyyRCh7FeqNQ/3mkE49imYbuqSBBRG0qe5UQ0pfy/JMAtAGuwE6HCeQ
wSJ1I3DXOE4/mKji/cS/ZQWTVfjQuwiy73lBcicgXXkA8mzPLDuK+CBRiy8zxZaC
2J6meCwMtBpRsCF/8peCu57eIn7HLwkS6hHKo2/Fh8eCa4MSOkrXiPGwsS4t/7Cj
TsNGnbNysjzLqJPKcsAIXGjnQUsdM1kybjmjpHoLSorahXppiN0Jg1HYuCeHefci
q4r0MD7ghzP6MWGRBEnrIgvP2rVF7EQuKH/8+FEKRIKSqW0AS8i0pbroLkM6NMii
5nVeFCpDNdm/e0vgUP8tBtW+Q0Ir40CU8kUDaWSWpeooWIWecKnRQLz86prIQWBa
fOJFOKdZjBCUXewmoRM1fndTYl7H7RJTPFBfuYl8cfA0rTnGvMzl9uKl548Pzm+8
ZOlkoOmCj2SZscLGpYU4efH1x4RCAXuzDvec1XDzhhCvcsBIf8wZOKjX/TswZKhQ
YtcoVHfmXnaXChm2p97kOilrN0yTC37z2vnrMYg5B24dZu9rn527SDxvB9xtows/
vQYBDWEv2/nKTnphL4NXj3tMCZLEN8/lTrHYwuMwR4sl3iMvKkCb0qifv1nXoM4E
DNhbml1WjGrEMvl3Z1xI+JkCaqJqmVuKwQFqpxTYx6ogcGynSwVjsfl2Az5B2ZXi
L3dSHKMMi8ryxq37AdHCMu5QNI0d1hKJm0/OmDrrDZJj5KzDui2Csrlv2KRQvhQY
mNHe/y0E7jflrEJ0cKg5hs5LV9N5g7WRJ5IrIDY6Q0F3smJVVmQsgB1X9uk1Fl5N
X7dgQ7VlYclZmoVFMbYwKtQXz4migS+NNI4Afn58uBjsdbQH2z/5oCs2vJPvBG5x
xjdnIwxG6OTN8y5HNo+ytDYR6keRxdiUiLqFD769qhkiiQT2EFzxa1q0x8NPyZxy
a1g6RlJJAnMiHe+Z/T/nLv3QqZ4JarHZgVMAcnwKP98m6yZEb2BgSuTxuZEFahAe
7Vj34aBkHKvjl0f0WVuQ+HdMWIbSwGIvfrPymbQgdw+JdicaMreu56H8r61YsEET
b/dDhS6hvbXuYy6dMRydSUIuZPPTKAY2dG8OL+Rj0RJ8IXiyV1novDpFE/paOUat
fiLS4jdLsAzhrl4c56ktJ9hNlfAOIL5UadKqkHFaeBTSn3NATqdt7elkr574Nzcm
JNksROxC8iOP8JM7eBb8VzroIhEHRJSZq8bSuxNrPfLuMrHbIUcWskDkTUBrI1ck
tv2X+Lt91UAXAyOukGGroysR9fHqsaWbPC6Va4hT/gY5Mrry9s2cxKI4Y8/tkLqx
Gj/0KBggHqSxm5nOS9UkMhEF2CURaLR/Z9MP3MH9CovtM6uCasIOsPjx7GxmPiDn
8ukiKqJLeJ46Jji3aSuuTBTviM93vRvf7+feCA1D0MqmckcEQOcPztigOvLJg+Lo
GHvMrFPSovxUILnlZKnfEPBuEh/GLaVi9w94yaAJTVFe5TBqGkGCm0zKRt9WFUeh
jQlow+HGtqi9sRweXIAXKrGICcgcKJKIxbndXPrYD2z/mCwLdabLBuAdR7OQmjyr
Vr2DfR3Zbj98ecK2WOA5U8KCQEEP66F2JwZPz/jXYqStOW51VU0ES8feWwP0dzid
umX6cJT1wqKJPzwza7kttbiARiTfe2rgixiK66irBVyOcAPZIs7kpr9n8wvup7sB
eb+3OQicOfDSOSXaJc47BhlUjO9uEhx+3TpnDoXnc1IOqnDoIOFJPx8T4IQVSbot
MXZvbYlEV9R0hC7RE7GL59rV41bTUvnBe8HF0e3366RUbKS/eGYksqIAJUQhN/ln
Rts+w+Zcd0vjTCUg4E02oKhqVgenL47ItOEEpd4LhzSZ4nQLvCS77Be2z0OU5Izq
ZPaFMw7s63OF0ljX7jMK+NGOFTRCfIW5cvG/e9veJDkBG8JjLzC36AlQZuU9blNp
qM3fjyp9MgnBUGE/BSJOnKstiYiQ72wMH0y0MTLrPZFCz8S3jA99P/3LYUyOVTiU
nNz9ojNUpXPXVdTvj3hc/gxqV7igTWNoV7evqLbWW5m8T/hn0av8gJ3BSY37ckCS
d5X2brZteVUwVV75yBYGpRc8qFTrIuW5wVCpK1Zz4BRf3HGZp+gPytoVcd+3AMmH
sUTWIVkg05BPBIEuKrzqStsLScuWlp5hkmBz2q11vrzyO1jwqoot8L0Z1SDvv/nX
1wIliH4CbOhWs74EJLlGT/uh7DOEbdNDUCo4hXfpvYCl/hWdlZqD9dgA4kYSMlq0
pzRDY0pLS0HIVJ82VNW2/2VrWssr/IFEAEcGnDkxsz8YFFsUnKVfdvSwVMLm6+6M
rWHb+4qdhKiH2T+sW0KnWL2SCvkqpRxxLTjWphiusGQghRwDt/egM1XJvg2ZFRqw
mVO7c7Pe1EgKvvonK666BDT8Tbd+MyqO0sCTW7oBzAQNguc/wEq0sNUIUeoOyjvi
t6zRvgWtqWp7mYWbAA2uls+a9o+VL2xfSPZssQPLBLM1PCBnH+Hrtuq1xAy9mbBa
UzDh9F/cTm1057/je/AsJPeQkhreH3XJ34AJL2T+yFmb2WUqJXvCr158nm8rpGNs
slvWgahkJ3FrPoUz1AmILFXRnd9WM1Otqwh+njPADQNe+8i2fR+VGz9Q4U8Uqw0B
TpkyGPJQLLIKW4N1h7Ed+MYLOLSy4mDk4gDh5edz+gUvzvy7PTT4v9XZ2Ckd2KO9
Rpah+LCEEGbW63nyQ1uDjFFjc0jvR85KcldPPS54BCIHOpIxWrG9+Lim1AYoTES4
uP9d95XkLNH3H6te0WOGsb9ilwDCpNhwnQ4YI6DtUVPZNQ9Ek+QGOxpJh16h4BVd
qftRez3eSz+tQjliVcYm6XikupXREbCtUwvez9G8bcviSLkFRnpzDqW4ZmrHlow1
qxiYd49l+vR24qFLZWROexext5xJObtKsgQQBnR3sqw6s1vXv6cSw+HxHSRMPo1Q
zENWHttF5aQpyvDbgvnXK6SlsluiOEDZr/FjvoOuJapC9jp7ekm6M/Iv8oU51W2m
Bi4y8v5FClVkbfYjfRU+IHXsDeeFoVlKkVJi/uoyXuvE3avdCww+q8JjA7SLbXmi
pMz2IQxhopdVrqPF7OCr6hH80snpk/+JB5/HTwzefPzJYwkSnzSuhsXmeJrdvmqq
8q9kvyihGB4glZ9TYuEmz5pIFO50f98em+I93CQMx25C8qL9+6hsGKavXPH5OMzK
qAIspZ8B/fZAj1fTb/ErwtKG71LtW2EhDg+/XAUMYSjT4zkiMpY5ymuBmtaKb7EV
KugGufQYhR+Ja0jTi0sBLg6nBdlypnembKzTSDdTsu8RqQ3s+KsE7F3+zcy2Gj9P
X/1qdEhVwDUvNNTQLayDcKiz+FGwn4PKFEDmnvv41RmO/Wloed7xIUZFDYXnHuct
Iv7aMxdXCWoi+r77XvRQvQJ0FTW75myJNaQGPd5Xx1XuzYGc2lbgDCXmHyUEeLmE
6bax+BJVhvUGFrN+QV5+RFIXsWG2wAfGdlnaPBuwJeYwXAuRVHqPWCLNsCz7eexg
kadU8BjkeNaJ49QnIVuMYngprU/a/35g7OnY82foFIFI7PYgXhpNWhI6v9qcbGmC
mLULmNioJcX44sqshw544mK7tiGe/chWTAe8ADErhc1LqGGEwVxhbw00/huan7Nc
7uN1XiSVpT186RJLt3CKsj6EBp6DXEsDMApEfwPqlcac/epXwwCU5XcwwzQGYHaY
GpL+qhHD64XBUzNTIiY2OSU076TWTXjfs/AoL76FeW2z20ogdLWnFUMrTuQn+gGl
pr46ewvfMYDl3zTTx4dlLi+C50O2Yz47YozjjWBeb1JyOU9PAldiyc6VSqPx7xAF
9KJCalTlf19dOP3r+tnsai2ZgBNLc81A/40ISLK3sGI0wdZWuKA1fxhjoZhNI3Q3
HhPl77kG1vXMCuX51h4AQs0ARppUgeFXp8Qb6fgFLsIddoKvPZ4ZqGBo07CXf6ws
Om8zyYqDASwaj6R7VMG7DZaEZ8OedvLSbjUzh8NNU2l3I8hSntp+fNCj7GnC8OzG
dQF75PGxILe7jnCfJfTVgkV1rH6pL9E6cjihHoaws9iR4ckS5xkSbGFgtKjN18Hh
9dSelZm6DtibZkX/ZYlRHOGxCoz8kGhn4NAaOpB9rKLDcH1XhEJkmQxBJzadg7tA
+ApZNjscIS9DC9DcThcPl7vgTEIgMkR4HKROVL2d19NYiqSgdqLW+ExRzVfIYjVS
DH3Ki5zy9RLS9hfYAIdeXohe/r8rnlKoD/v8XS/wmuYLFOzdHjgZ9Vvm2FFkCCtL
qCgzL+BfDYwBCZuVM1PTH78AYMz/mYm3i1Rdko3Ys6S/e4wc4b6s7mBlE9hQ5cbr
YD1JNQeTgxNIMwxve1sssenN8HdHtLYkEB4E9nZ/VmGZtBsZcFUepZoSStya22qM
1EMxhzQhhCQrLQd9upknpSOpSdeQif9qqkKIkxJRe9/9YOgjP8lW7XpD2Tsd9Kt8
9G2IBOB6YpVULpzhYCJdhhcnGxzeW4a31xKVmZpdnh0T84N2sZtj1XRRLPkg1ItM
gSdJ7aTciKuizCOIUwEYkyluIxt9OmwiUm6MOUaqGS3Ch+e97X4eWhIneTdDJfz6
HAGB33Z71xkS8vpm7CDiLv95GI7y68Xav0uKitG6CrculEaNZgoqieK6nQ4vOKlo
YR+h+8U4yZbxoJF4NuXI4njMyKf6M2z31bHsQEbqRUUeHEoevdHYo3dQD7ePvOyy
olbPFdVKSYbhK2F9PpwbE77aLS9sTECdg72SQ+DjkIcjqTCgppZpgAzOQ4dKAH9a
NhfGoRDgFP58caXJvMh+FV/HcUCJwCjiNcWTDRSaM6O45pGiqNQnISafAeMTK1Su
r+aqM9cyohkdVwEGCo7JdFbNciEMQr2oe21Y2vn2UfSXlmD85w6GkhxbPFo5/I30
BSyzjS+0KNKeq7CD0ZbXeBDfHpO/vPOiGbn9KbgiTpb2Zvah12waPdC0PKYMDN1p
r3CmOb4YCiS+SQ7EQBZZdqEHG8FB78DN1oOglin3vAIFT/RCiltdNZPhc201TL7z
yLa/lvwmVpFiRKdDN5fa8bVZNF/VZTMkSK8gsqEszuA+b9eHNd2WZZ3CYufzJprI
eO1oEQIZ+I+8StlUlkC3eETuggYjq6SzQjjTI1dHzwGaa6uo6JfT+8L5vdv3EVl9
wFKqe0kTtovnjNrsZ2uOYUchhaAN73Fo9j47UY8VQlwlqYXtMKqpHB6QsGeEZ/HM
jtGLMtEahropE6v8RLxZ1ycjJhPCGs1iwyZU5Tq43OzysPM3BJAbbplrtvV3/TnU
kEPkVQCeusMWknmBQVWrQvse0x+x0AAYQBSsU10bKVD1I3z3DNp6My5pwebgVr7+
lOwUGLfHIzmWjsSo7pZSnK80sdk7XBPZ+7I7GMDV921mHMnQT0GbmgvTaL5Em7SR
R0HwkNgzfyAp2VuCftBZyfC/7oz0xCfTNl/yuXQP3BJnDpHMj6FONnmqR8+/Ulw6
Ih7zzfS+jZcZsAFCSxRDNREKp4Ud42v4gMsB/tGjlOUzIQA2yovJcbH6xeQOeN4Y
VyiZ0FxZmZiHaH0cTHox572+25x19Bugv7b8/xaOelHOQHNyl05hWhoTKq4edCoh
hwcInLMXFePPPlEwAdxe6Eqzt/cFIfIITfsuvngA0CJoEqMr2r3z8lM+TCutoIQu
MJ84SxwE/lvJT230ztvNpJVqe1tByX9Hmcob9/Pq1jntkaw8KOnqOShFe9kZhD/t
74Oxsipk5M1vO8azU9BTEvH0jXAWPz+FxzVCFfbuseIYUbSrXKs+MgVbR73m0iQJ
egaDGyfCzjt3memDbWEl8WdHppYIupoQx1xnjzgA/HHQPy6zoU/lCnZe8CjwP+gG
rGiv5Mm4CnM+t+lvwE3w5r1mHE3cnTdWD3QLlanJouatSmte9th1ki3sK4iNTu2s
ha2vGtwGUPlys++Qv8jvbhMQhuKR6DqFfA00d2arUpF00U+QkR6MaRXf2x3ePEJu
up6r8UPAtzTO3eSnV+oI2RpizBkHVk8U6ntWNXXo8neb+jwLmTsAJdRMFdvfYUu0
WSxfxKe2bVsmL6/NlFu8SywDsOhQX3nv1CLD7wo/+3QvyCI++i1Gc6SFL2nZ5awr
GBVAqPpsHMBkkQMnlIdZDfBXxl8i/FnIVVO6WSlJLwiiICpuRCJaRklrbx9VjlS4
lmOHUnWGRrBZd2ECe1PKu6BQG6oRc4g6xHZRAXUfX5pXBG2DyD1niWe+oHiQRbo1
lPD7YQFQ3XoJoyxAM4RJNapIpjLJzmAML9Nxu6xuRMWQipT7IGaMXYwCnWOvAgm1
GmBPdjyUquTzSb81Y1suhXR5q60cYAjOu5Gc06RtD3M/q7rKzSAIcdHT55hywd3d
0lsZbqhiQJsyDounSBVUdYIqU6ND59WP7aegiqvpVrAhY7ZOhNOXNXvsraR++5gO
edPAEXyqUcrzAv3EgSOPkHIwuWS0aJNw6LDB5dLCoYTE1C5tizZwDZCOLxKIahLJ
c+93ICqWxkqixTFBCn/dB85mbFooPjXx40JSGzmuXXCEd6vFEg+b4A1lRKG9WwRA
2rW0SPe4uw5TmcsrbTdOQXotnYSh5BZL5P86wEUNlVkgWas5lH727hTrtbZxjvQ5
P1NJu/u8pVXu/OkNT9calS60xdEhEyM3m2lKef5paTRf1rwIyrsmLKwQERAN2+9/
AnHhICaywTFKlpFcrB0TOrJxSXAnZ75aTTYAfCiknSb25xbuad5Uq6jBAv74qhEw
hJqxyc8VSM44cv29vEenF6PmDUjlxQ29LNMJBslcYxIJS34pfmUDe6k/apzzn25y
GKTciX7tTovwr9a6uKoJPB6u9SSLbiImA09xC8sg2UICM7XYSRfBH1Vy+O7RzhCg
djwhsEO32nMAIGGQUMwPDwXRIUpLHUQPtctmOcNWundsRR97+5nRQF/Aw44ZWIPr
W5cHedJ0Qm35YCB++QoPx1e7BOPtPATmN0T5Kw0vLS8g2L/Z/WuuVQawxg9xWRQv
7oZvTrkf/9WWwud6WpIpjic0e0LavBGwZwiTuHWVOjdfMtZpo+c+RzfL8JJ75fXH
/SPJRYNIIEst49jSOCq81sbUqlt4KAVs6yqAxs9xs1rzSfAC/RxCV4SM3SphsZWy
k+xgRz21Qj0jZapE0RfYaYoPK8Hp6UVFoyNXmnZEuIq2/MgZJlAsCWuDGp6cvXvV
0LYBKQKYOotQ1+1XICSMS/j+bm9CuE8An/cb5klLmbPbaETIsWZWsuwDe6iN2I+0
1JIDOB9wUPq32Pcdpng9w+zONRsPjToCPiB5w3u4tPb+7nzFQF9BIE2rdH+wzTbR
HOS+8hw+wp00CkpOG8ZJQIkXJJ/mnyXUHJM60W+/EnW8+rhzYUDtcfXkVuPo2nCq
LqbcmDuZ0JgRe9DnkqDWy8teOojiJbXLVSMy30IY0/mzqun6yt/UqBmxeDq3wepi
grEm8BEOhhNAsZ6LIMKZPqOxyJSezwWl6gKMOVix17Dhf5iqjquAe6taAUWVO4DB
X4oHow89iT/BFkVBtynC/wFbu3OFa8MBIesfr2Mebd1Q3QuaMa0/QaGyzbibJhPR
cbzNCf5FvCe9UzRGPuyCVYClj701PJKO9YwYQjYdlu1JPm7vM+fG5Z2XvNHOc6eO
af1lBtc1ksCk4xpMlQSQ6ggBnu9gqgvfaf0f20IR79IvfNyNctqCjU2ntz/7qUBM
ekA2u9YaZz6AyaKKjluce4dYkK0tZBSVJnVr8hMYKXt5UFQhWa2wbiUNVsGXLJXo
GfOYv4SKhmKnyoRfjhLLfIAvhIRej7gkNWcak41kEG1ILdbHA3HkZeCRZhw3bJ8g
JgoITOYKsr/e4wHnlxO7ugS5LqihMC2feznwYEO/j0mX97IqN2rrl2ijdeb9Q1Mo
9NxqfpQJi4OEndneX1j7jk15qtzqEWkoo32oXzXl5yawGIYhjc8I/h+GK6RJEYv+
MuhPoQzf1Tyv7lttOgd1R6Nkf+8lJLouTvnOdUcJX7TIcN1VUpKIzsagxNVkIGac
cMxYrU3Vk4Oo9wL+FB+imrDMxJc8fj4pnEacpUS7fXnFSB4/Yt817aithE/rgr9R
DSXlQD0Ku0MUhseSuGDNR0fZ6hTgifAGiHVIutjEzMcjH3QZaG0z6mU4ABAVLCzS
qBpFaiBAmw4yymFqR2ralNYRxw+mogag2IJqRlzP7XH8msmZM2DUfY9yWlpoZv5d
m1g6Ki052KNRCiYy87WpZAjJVzfZjgdF1274Fm2ldzVcqIJ3qE2arziB30oLMz7K
tVeqVmqU/38irr/3/dt9VsBwZLhsWTkeEdRfT81KA+qrZ2z3e3Xu8Z1VF+SFyR1/
UyygAt4s6DM48Vj9b58h2S9n86m020GqyDYb2zpqUBzNncdUjyEpGZYd4B5/WK+y
SlIo7zKbQ1gwWtdidaa+Bf12d0eSnMAgkH/NRrDyZJ8lGJYMVh/9Yvm4tgnlQ10J
5r+X/ksuMqHSAdOck2shcmdXxisQ8+sSuqFmfQ2p44TZ/Qnxyx59dr+LPfD/rWEC
JVV2eSlT9LumvJjX3IKZrzDRDMGUPaPMUacja0jk2d/LGKfZKfq2Y2fTbteUYn97
eofaxczE0KUBX3adctWqiKNmHxnWP6X2r7TyN4025SdH/1in3xC2noX419mU6xz/
6Ig7cAJjYmx8kPcIZTUw1t4wr5hVWObmxr5IdmleOZTrBLUaMq4Np2lMizAB2h2+
0CdEQr9560pdfwMii4QFi2NzwVtSkRT7nWxL2ax/LxD83A1/5O6OPIcrDuyFflN7
68PT9AYeaWOnfHyf4LoIEOTwaDiTlVfbjgfX3yquOrGNzO/UUoFBqAhnRklrpkcm
RdUUdXERn4W6QmNmUBYrelEI0L7qLBRiWPibyLN+AQr8zxmtDetqE4L9xtM/Je/8
mrE+e9Vhy1qhYwfbBrdySxICZxB9NiSHNq1rpuf7BpXVnfFYMTyM8IR3tKIHmAwW
yvimp4vkpDGNZiFCPxIWLJc8XPI5wdSyAQR64fh86B0/G8nGpLM5OVo+kgGaCvun
pb04XxJ9OmQ2hqoSlGn2NYq3uMnLlFaP3H0A+htUb3DjfHMiFp9hrRSjFJ1Px/6Y
Y4/a2oawN/Naz23T5DmKjpsd4ncu3fkGMhPI8ABrNbqoWOBxtEPTf+qyky0vjq/y
9t4S05K5m8TszOYd9xtPB+xlVjHfutxbc5H1QxNoJbPHseiYvDyeib3k8iZQVMpQ
FhvTe6LS28WlhWffvyppkiE2IfAxXtVz7dT57CwZcEKxtd17fODU5SG0C5a4QLYw
9STZj38MVFVl4tzVsKPHHguitR/8iHEknNFHaGFsrShnyEqqwRqTsqan/7chGkps
U8vD5Bcz7LYqcJ2XzxFqsV0uultqQWeHk3kFGNpJphkHyp22OC9zehpLWr+K7z9C
63cMJHTimOlaUlsGVXtlVc77Cg6+oy8yPgNks6X1VItD5Vhx2/MUr+6+qvKZlwzy
Fb647zigVbbnFkTSk2MTFVC46AJoi+qBNU9qRTjL3IrxDnTetaF3r0RkufemnMbM
TrDCikOeWi8ELUNxPRRrXJNscHlgYwbQjpIoTYgCN0YnL3KCmv5Z/c1sxk+fOtyA
6gNK4W8BdyQwhBXfCpB4Qs+thd5EuX23N6uDFaKD7oDG9iMUSqYysf1qaB4wz2k6
JOEBU9EqAwcseuwQbL7daJYnlsz/GG4P+Wq5sNQxxX28ye7R57lfaGWAF0EIVjb/
x8SU0Av0onyoTv+nysX9AEEAxG66zH1QzTcqtNGY5NKNX1yTq7fjU3mSXFPMxGxp
aU0w1EPGvzN6ocfbCQuiWSHUafw6T+u4Y0SEQtcRNy7CyAg+83HhwjYxqIRmq9DT
WjtGQ+8yx3mgCkQi2nXZy54UcuemDiBI8ReDimRH1MDyEVj/PYrS1iWrpn+YQZVt
uhmZhkm0GiTTLvxAQQm2QCVuOfUOQZAoh1GDuGYZxKeMAMKluideJRjHO9lelASs
8Zpk6bD7CkW/lPhrJSzLSBXHhV4xq6yvSe7hfXx7MceeTdRnKMAX56AAHjnpvQzt
dXahwfZjJ6FG28V2quSiWzJEvWA1EguLyf1lDBjaWESnJOBKQRFzhHFIjrjDK9hy
LFwO7/qPAyauxepzFD5j83ErQfPg2agc3DA/2cOynbw6j9RPdtcEiaL8+Gb4MLzw
nEqigXrb7jt+7cZ3OxMwGXMGxgtEo8SZ8uldXcCmJHlEtYc5JuwmYU3i5mO5MW03
lujr/dZ08kIpQ16L422eEIJu9ARwso7i92WT4MKw6WGLkGN/AV0mhFBBKNJ8ZgDf
vO7l5MGy2dtz9c5p7GFmLIa+MsZ9AJJmEQG6TSv3lD5OipBSlKUpgmVNiYAbZEeg
tQaPv5fEHNT0SPna6FJcPZ8TjiMxMXflwROD6bT97s903QNr9XNxy5Dpgw4L0XHR
44wjs7Q0PgL1ejZsfm7G1MHGkuzIqtVUsnoeQiMKzU6Xi4QtV4vuK2ccSoYcKiT9
OW1ClDm9OPRhjeQBx2RKBCHIXGYu56nO4ljQXYBcEwb1gIG1+QtNmQNJydXu2atj
Zw33/nxQYFs1qvg2ueXhndKwyPJ/Nt03pINtuEcvXDp8xpGts6zmHRbZ67N5ukGk
bx53nPDxS5dOz2GFMOe4ghDqmRGMRDSZo1HZNi8sAKHMUH1fvf/VFgkoIlni8cdB
ElHmxkpWi1bSb5fxfzGu2l5PhdfGXu8/gxVy18l9FzAQcecQzAUZdWPHUUuDIzkm
P0NU90KlM+B1g1UImkaNWbKUmUPab72SD8gnlkWL+dRFqKXos3ckn8MC5Mwd5rBS
Ps/fXuHmNaP9hGHK8gDiWSG9Sufh+krh/MqccWM9ZSHUL0TKIJLEK/rQV8phUtGu
dWjteCDzQ32yj542jKg59wVY4g5LGXSEyzrZa5VQ5boKkz/ljfgA0gK9f5JWIwgv
wfzTHp3ypdN0x3AQVa7QE3LmBXD82xPq4oBOdL7Ulh5QFuA5Xb6D5vlTSzgniwSE
yrGvLQXfCY2F9YoV8+Pwqzs5Pkp1sXY6ekFZLimLplev8L2wgMAHn3s7J/D+WlFj
HZv8dfbzyBDLmmuNqQo00bwIULHBsVQi96871SnLK9j9GrbjhQnxWpDWgclNIO2B
6wh0+JCX8U3JlkucNxHjMkDBPw/AbtQ3dBDGZ4NGqQKLvtzsHbTw5Vdel2WVgsFx
knptEr4hiwyHZE+4N/N2ogPsNo1K22yQV1IqxMO54KO3EU16rlEi+2KgINaoj3RY
mODNT/0Ez1V0l6D5kevRBeViQI6AUkfZrYdAvpnnPohX61jz6NAs/K8UPrHCacVt
btiD6FtWpj/DQfYGRfckoHJmtHoPlsxrpJmOImGblljKBRIpRFpERobMGSSxYHX0
PyKW+hAJyLjev/spvPv1PBiqG3GkRUeq9GxyCMU/+QbiHy3xPFABTt68h5xlujd5
CWga81I2AxUrn2K2RJkQfI9IpP6lBjDaHY9l84P3HkeHt1vHGyJTYvTe1nXqzlNa
ph7tMbamIH6rCJyGp1WuYaN94Oc2Q1dzQxbcQ44YjY14HajaTesNEmEU/Wfl1tLl
Ec3MnEuWjXyZ9/bXUHsQ5jDqi34EogmeIEBl3Uibv6y7U+P4fAs8z62sLR6iarl8
zKvhHY7GyRrkb/+P4QCeb5cJTv9fZ5PwnnGnYJckpgvvOFenhuOHS9X+HH6Fsssd
8/5tx4pbXtGUYL/GExhas7B/17sd6a+J6uzxZjuTFbB0XM0fyaGGmQztIpvmpBCS
U16HUkM/Ns2OkJWpYQIE+GevE4V1yWs7KUk+HXnNXSCPZl1/3wsX7PZgpFFH1lYF
cxpE75pYCPrODHLp6r2SYaj3xJhSUQLqJOZ9OsiSJq9U6qxakPemo7SPqlEb5nH9
TdQ71LwW0s6BBkEa7ibD0dFNGRL4rQggqNv8bSEuYQClq79Y0/4mUBQ45szBku3l
32G7DZ9P/gKJG46TIH9sNO+t+G1LRk0qLltBwgN1uuRGi7c77nOYSgBrFareibp2
H/UGoPb1qm8VVgEC0irVNSMu9AP/pBazSwg2xmyxfIl8S/GIGr3NIbG3xvwX0YLQ
4FhQyOlc28rvX0m5LPR0G+4ltOwyinpNsR4bshgGL+7vekTswuQYoAjL2UPkleFI
TNvuMmfnhT4RblfGO8uulza6ob6v2hT0aVA2hN5j3HZbtjxVRI3+ZjgpJ08kS8Ru
WQxDwfOWA06N6+5bYAnkM/eivMbtBGJKiBpm2s1tKliDLj8s9jYcxH/byDOTzws1
zxeVUpVaI9vnc14VPTwfpEq8FVLt8O7+7WpA4ZJ6OQ1otS6/s2tTt9qunP8HRWnR
snURoNugKCuK+XJ6DNghhwY1Xq2cJmzRVMb0cYeQn2/X8fRPWhzgVtenBI4M1B3I
oVQiDLe2zKVtSRJncL3F9pEM0uXXOpvKv1lf5cWsVIOoPNiiOsIF8z4m3gGsK78A
53XzPRQ4odEloxHKNRPwTBAefr1Oes6mVExlMg8Hl64sgWaio1nNCszj3jQnB6fR
lRsWwCaeTiwN5QIo7UTIl1svK+8JzewTV+tK0M9txWaUZkv4o4DyObetlQOVKsOo
zB4UJq2aiXQJo9guFG1ZZPfKRTEL6kNuRryrqhF2HXYdIokDDSwKV7XIC4S/9yz/
Kv5vFJc/8kF3O/a7T/zBlS+Y2xQFQT/qYMWBeR7Dc/xZPGaGNH3vwNggw8PYWZo0
iv1+7Atx4VxP6AgDUloHHFslltHTtEHAKEAbrtiLxgdpD14z+xZCv2vD/aOOK2KK
CQeHNczk5XUcnNG4aUHsZXXDzr56LqCOwQ509ZJ4XtEmq5zv+ygeBu5JuzeBXMhr
rOiDw7e3TH9890n03bph+P3BmGxqAReFOM0XN4WLqHeTi3ah+61B+eFMet1IJA67
VnsRSxpCzMYFbZzU00Ky/aAxv0a59/YUqli2rBARygvueqoTJofnoKV/XHDPjh9n
u7Ni6LF5EQBokcFRZffwYQBD4Fb/iVJ6j4GsXbUnk5Ch0IZQwiESyfy6Bs3UADyQ
sn74M+g5eQYnYVZqdYxMYSlan5gLzke3bRUG3RdaStVJv9wtc2A5Ft7TWd3jUXyv
IKfKC/wSaJqIBwU9KLhc4Xz+601r5RXOKFwHpeKyZ04x12yyPjh9RnR2mEniNZJC
xl1/3dbeeUEw5qai3QAjiIDXUeBsPvXKLkAuPGkPVyg+4BB4rt2jB1gAQ9E4SkTU
VAOcI7tCHasPsM4ZOe0dgn7uqhaiK6LrBD9gFN94Qh2+MhSan6bPuA3AQg7onbhO
CWD5UqxKT588QqOXWQJf+CUlS6LrH4w52j1eIPOnAPuiLWqOwo0DfcpPLM5qFzJm
pv1x1L9pMmfFD0oHasY+s0z5dKEgViyplGtSQdPGsR3a1rMSWaBekMPBuumeu/gK
zWFiSDHOpjwZ7yHMMuzA5EeAdHcOc3mk5oQwiJl4kZxactTK7VwB1hJfJ9/CD/OP
KfDauY/p0FlCAzirFhufvua6jfwuQZZfJ7jA0+3pO5i2VKlnKy8s+olLzpEWJS9l
Q20G9n1jGqjsMYET93HhNIpBDgmQ8GrL0fmplH+i/UfHdMQQGL+dqdJ7nACy8wxM
wZoHY1N++GmPLeZhGnx/Xu81QBaJ4Tc1u8aLqWHkrbmd7C6YdTairlA1abenfmq/
Gole8nwIvnacu/pGxFjQpEEWrhvKyaDZlmOMHPmpoWK2eCl8EdH61nUYbp5zteHg
E9gS0VLdIPN6H3ifnwkQGa1lFAdPLadr2/i8AWd1tpK55QfpOQCr7DuS8QtIkULP
G0myBowrGEScPoEH3ACr5tj1rk8FL2//a0mdu7cp447fNq0Y3DiyxlhVHeQkOeWj
84yFN6Eq0kRf2UBgzJHw+93xMfExosYEAveaX1m+mLdYgcwoMl3tz0GEw5kLYApy
S0gKeYpwMGYhy4kFo/nF1sGpnjbEppAfNd6eeNofwTPkS473VIE9Tlc65PS9uE2x
6NC1mBvEBPaM+y1PCka3WipXJYyegvvBkvXu2AHa7ixI6RMlYoZBm773PnvS1nqs
dFYMkHKbD5gPse4jVMxVNIHO1PZxyXpzQMPLOpRKZj7E+xtL5BLAtQIu7hKDaB70
73DZe5WiOLDVrEQpL4goenX0+DEGslxvP2d3QuW+hbw9NJPQ5FaTr9RexhKYzlFi
g0b0BZMdSzBUiLj+E2dIcqgQg7T9hcMJgHEC40YFHfg5QYtmymVrGUabsKCaZ1K2
Qc0F5NHNQCCpf/u7y9SjaYptrZ8dI1Jgax4leihJ9ncr2+VTYPJQVQjia2Hw53vB
d03eyfWslIedzHkghS2+xJolpRVYU5YLDvwj3+5cwVbIdpWV24Xn/5Hp15ZXIBmj
+8HESrinJBqKzRo7GiKbHfsTvme/cCrQk3kn+DM2aMDstVVKSETZCLsh/gLCorUr
c0IXaTFKjf8ZJixIXPi+8MQb8JHGk6pwJDQFJ9tLqpnt/+0OXrj4BsCjRKETfAGf
XOa3fc4qV6mUgsREXJLx7+wCUsED6u+qTuVBCRKG4rhRcWpEOA4A+1wIU+/155uM
zU5+RhiKMpdbW7C3oodkTegmXqZbyDjN6uNVZvMoS84oVZLPAIZouWp5fir4wcQT
hvV57oXtI/MINmClr4/+TLoS9/MuUAHb2SPhKN9gb9Qa1Rgcv1AFZocXTqQfhnT9
f6WB1+hQjuYW5XxzbfNTksnsKNaP5vCHtGrvIrZxuuXhQNO0VQnOKSXhywB9ylq+
UyYfvDTpwu1ILsJokDMJMlrEA6OlBOSgsIMxwTqOZgB6wYS5hqS6NTSJId64790R
KSjbQn+tU74i32euNO0mbA3wiNEE8WzgBFJQDstfqo/FO+dM6ERTIIhjSS+VrRF6
GGc7xMhyqvC5DYFLwBsxACZ17nzkZMdogzGsGGTXeat9eND+r/IQARDdEDM8u8HX
CX3admm6Hr0Ch2VkNXDbHqyYcgoYTbHUPjSZLkpHG6e2JT2pDvcTZAQ92UfTY17G
8wWQkhHqlRbUQSTfQQ2HvelGwUaxXfSQa6liFE7PUZ1OSlFYz/j7iAzAy42YKz9L
dz4EIug7RmexlibTftuQGJRjV1ic9GVtRwfduXfjf4G9o8FlAJrXx1tHsU4ZTMF/
MFbbKyy+BQ9MJHaonv5Lai6AItXusbQWEy36Iwa0EXoHnlfLCz6FUHzaDDKpK1JH
ymkNY2rqND1/o++6F3aKDlqLVRBVTZ1/rAaxd4u6lDUM9AekDk1e33jqhJtGMFP5
cAXkvvq2lm2emgB58u2pGE3cuO16Lw81hOEd7AS5NqQp/AndyZTimecg5yPH41ZT
pTx6fnG9X+AG844PqpHFuhg2rwvfVYRSd/pQL533S9jIqnEk4JuCHqYvEpQD+UUo
k23RWGpxPR6q4jJXKh/COCVc48EnPNV1UZXL5rEeiWDtz7u058jd6Nb57Vlpkn4/
jYDny9HNzsmNfe/HMqPtBU32b4mOap4MurjBrlRH760HCpFMNv6peDMbFy3X2dZz
tfYpiecIR0RoB5AocooncJTqXY+rdcFVrRgkL14mH5LPaNkA+qjF1jUbgZMz2X27
34ZDmLGXvOUU+NWGxFAV48LJJlH6+CgYH6yqlJzdv6RY7oawUjqT7+uniVm8y2u1
1TS7Z9OM4dii/jxKId4IBWZEmITSTwYynqaDbKss9JuoU1VDW0/z8DX+wn2wHvP1
xMIU8BaR46jcHqtsv93REEeXgV1fWPdB3A3FnmXeQQ/Z50cYm8AUGrNIg9EHwx2F
fvFzAFGCY+LB/jXVH/Eo9wI+LvYALYY1f49UuR5KGsDPIh7Ivx93FhmZKhQDjOTa
qkrerqaHa5tRZqIxVYHmSg9jk//07Iamac2nnMAnEi5OMJw4Zl0n6F5vp4euWdoq
tU/PB0hj0sUu/dDuLEkOAIEvuRul6OvVnHbOzF3yE6fQXfl12K6edFWES6mZAA1x
Hjs0e2QJAvNE7mbmSE7K9Aup0XF44GKbyGXf2wNri+rJQI+1ZXypBt72gb6PD9K9
SefrrA62urublT9jMjobDMkEXoec9jeg4OeqGIkYART0UTSQ5OAvtt7p2xciiAr4
ZWzeDJ5fvJlyktxhkpGoT9xW724/xhS9p0gLDJnSe1p9QmZgNsmmKfbD8GLsXbEw
XmbZllR2HJntxqhfOQzZTEPmKtD4RkC5C1PTUTyGzgp/Wiold1CzUtdrtl/V4Qwr
bXYdty2zyrU5K+e2UgqH/m42SIz/OI4SQsIkNg1b+jMymEgDoXEdlT39AZaufJ8N
iuUNYRaO3GtzuiylMLp37sRgLQRil1KP9hjJqYVBK1pUJd6TibtXS9oNxt6ZeneA
BvYsZU/VtdqU1F9glGQn381YJnRS+wftRRFTd0i0nKFWkGgcKd8w+pKAXovHMwS7
tv31i8vgUyXki04r9QOrP+nhr8o0qmUBiHe/9W4MPwUNuUKkKHKhucQO/FpmoqTQ
tzouztvcC9/Xdn0oiytLyLvYY2gvrYh7y77E288U9k+ZEMi6GjVNyjuaxlPS2GYS
p7zrS2fEuQfjU6yy5ikwZeNLvfLob/jLaomC0NslX0ezjXx1vtdTKd7BslBkomDq
Cxr0wprTBxhyr+MSbYjvwwx3A7Ae2wOHGt656SpM2IEa03GzPIXBYMVJxks9Ty6J
R/UHdmSw2yWm2yIDfRoVflxua3WDjt2gewK8MhQzYZpcnGBi+BHPvt7+yNPBWHlI
6pdm2N3qIATeqdNLY0mpeqWAmbFyIMnHQOlkWomOzPWQxIviAEjpp+KAYUqRWowB
77VleGpl7cmWeNB/HtItGlGFD4R7KL+/xWQurywQQIQdWt0P0n7fWoEU+ogMMxAp
egOCCxlvFObBu9uwvH54k53fOcm5qaPkciSL2IagDzt3JGq/gK1bph+0PMqgLuVR
q9oYg1DBz+jUG7StA/zrlmCEXCtj7Gkd1FWn9oVGvxX9OIO6RNiSyHITQIqqSKuY
lj/apgZEa/pXH5Oz/IekvMOa2JxLZx2in/epgmtRl8Mrm9bqrHifpFtMJxx1xPhQ
mZ2z3sDay8jnnDgfIp8Ey3VPJSCwzcWJcrVN8HF6aWVN6WIXfG/xrS/NlBdEgTmc
prNND7NruwFIGMQJiquxVLYrGskFNn0I/kz5IrAIzSDfYqjxQBipcmaTLaDw9Q0h
kBLQEgDQ/wgdmU35/jdiQdLd6Euzk6awd67KA34EhhRKEGvSpguIx26O2k4HZ2F+
YBAtfwJuuBQk9HJjjE1IDwf3pB41//14bSGLtBARqYZ+6KaMUDniNcq1HYkNh1c9
EdEq98CYxK3gCMRIk2O9OF7+iAgHRu2mMzvqGxpbKirwfF2yXpkFuVgVtQ06/Tiv
bRfpWnUz91+FO7ozyMByKb2fETmEnN1N3ej4oALkmrddsT9J9bNrmCODzW7S2rVc
a0KsTunHd1liQcCtsc5nmFQizSXsb1SIKTKIqvAmSPQmAI41fa7WFEpL/Cla/1M7
z+rtuBDn25aAgHNuGPIB+qNl6uryg4fawIGFSSjH6Putasuu5LJNmFSS55hYjnRB
xQjFD3riCvyye5Rqk8YSeUPfEu49+qC4+Ldkh5tqm3qXRIOxiRavUoXqkfvx9Ep6
q6yv92Qh/YhMk/ICcA2oZ9wNtMFcG8t0dZnh5Qoi/FcLDoqsPbQGu5K/X2HoD3yn
bLvzDzLQyMDL4QfiXq6Oa6BL7bB/2KY/3KpShipCGapOu0hpSYBBmJUuWSobFzsd
Ojy2chNIjPFJDAQYR0eTB1c/DUN7Q1J6UnZsN1dcfANk2AulMSn4GmkdtKt83HLF
zeNBH9UmIyeZ0ozIdd0b2QoNPM7kYL+h4l/pELkpWiKpuQfS6JRGJek+HpSjE4I/
kJG9KPs5dbwQ6aQms7RtxwuB5jg2JDaBKNj7nmFBNWtCknE14NtyEgeH5MnvnXH4
bLAliizIeuoF4T7jGiWCd5cd0uPc8MAQd8Gk/Ma85iUGJZXP2wDDaOpZWMZcS1ue
/JTf9GbT4zoyWbpdFO853HZER0jNuHjHeGk5csxaTZDlb3io4laliEkbGE1/srNL
C2uzk5FEVTQ7tci8zJXwndy/qMUK5pRAYO1kO3UKoHY1R3fwK1Gj+Qg9YZt8pTzw
c+FAvEvXOhlsXNTE91aZokVn5ZS8r9pcE17eE4FZt9r23t4dLD/Mb4ErXFEMx2sz
7gOM6KfmwbPZSRpSShKYqgmpJHzvVTNTAhJ6Y+ltw+sTUNHChVGDWafbHGMCd9w2
A88wF/XgJZcHLlMNpYZ/APIEkjkMJqINPfWC7KNa7Jpn7xutPuEds0p4YfOj+rtB
Qq3xMbdh6M3fZ7j3sTa/WLrCNdLXhUasnDWYQLJMuwUsiFXJSLJMFRQ64Hd3Oh1B
aabVHopxXcO41GkF77YTdG6ThLyL+nNCWLOMfinSHXuWksuCdsEyvJHhdrJcUp94
PA9YL623hvvZXD5wo4c+FdEdY3epSsn0XoRArNmvCVbdHHvJhRhiLJX10ICGIRDw
jHKdw8NGi0OJhYN408V+tpagb/Xb6JyxUBQajDo/LbHvPoYmLeUcYdtLukDLvRwS
n1zhN7bUM6NmgG7l7sqL/53SXJ6XptWKmcvr5pTvcXRyCnhm+6W33Is4enlPMd4t
GC31KA4ejOXkk1uAAj4DYhif/rVFnJMCKvSKy0Xoiy3vpmCI8sIKaevNtG5fKNtF
wruYOQZWQubN8yhizMwhum8ScZfZ6KkQV+w2JplRl9poZsER09bpx0nu+7j+Oq1s
ByMKml1cuLB9H0DZ9zVncZl+Fjop6zU5GE/mDrfSAqIkFWbA1GbkCnstZU6eIDJD
oP16ln/FNSxWq+JjGzzSIhy/McRJiif+W9HG8+4YDwHtu2V6mg2nIhTS/LPRXy4Q
13EICxhX8eOLW+cRy56m6k4T3+R8yMHHbH640lEa9L1qiH5pZBvJk1kiryaZ+MN9
2/FXwGntU5hBKtYiUmVCKWZ6EHZPYQP7g1+aVzUg0Nr3VYhCmNZ8dX2hlZOpbyKr
5T0zknMtNSTQqM/VDNT6Ab9GWxgXT+4cTDmBV3N54ByxxBLFUkAX1KnwBWRW9zzf
FsJBMv3PFaQg3YqKMvF9SIkEoINOXmkA7vH+NfhxHVb9ohFh6BxKZLLyZJTwvVCD
jzDdRG71CtccJmtEzLi+H8vW46kUC+P8dMNFGhgcsgKlS5DFRIoFT65q9LCEtb8t
Wqs1UNlWJbjxalyUC5prD4S466tgp15OaZ2YT0fOESif+SyLhvW+fyzkttNBWk+n
U90X8+otIh3eMMi5dwjIUSMKb2YlPb3MErNwU3HaJUEPTLkOVj+AmMGkTyALrmRR
hg4zl18Awh7z3R33D0FA4o5Jpta49NmkkP89bKPh1D5p82mWGMQwiGma8g/nEk8B
UsXasHmUryRw0nn6eD1xcq9xaEmw5Im2M4vGls2kb6VbJ2ON6DljfYRFC8YJvvwC
7k0/bPHMxkYkeiBaIUuba5bIcdi1U6l8c5VEdaZgeoEK9tVKZLwnYI7YjVNHTkQF
Z0HKYulsXUQU3Mwm9D68jeyJaOC8QRdSsRQ1NmM5U0mfUzAY1Q6hNv/M3WVVi+jU
ClcRxDcMZHsCUTj8fSfbYejYVtj8hWmF1/pLQoqPypEj6evLrsmLddZP2lAF37w1
PjI0MLyOcOc39mz7yNPNdKyEZZmacLPBqMYG6gi5U5qXTe6Yedq6l794MP6r5Ecg
o8H3tSKpmDwT30FeJmzKWErm+c5JDXBqX5s41xV8CTkpnG1xKZORSXVwwQEnRHNR
B5Dfc0HyrFofQnYW9Pwmrze0Y2QkcRaOFBHJR+SRnkwJ8Xgu7WS9w9IQ8bHPSmNE
QHz5YxhG01MFMkq5B3lW3xOp5Efc/K1/KVgbilrjIJkDJbKR3iSnBmeZQPJKNTv+
/xlHZ5pc6GKEo1QEosMeYuk3FZvbboN0hbjgJPxTt1bA6ZDwDH+f0Boob0Htkv2r
Zh3Su+wJyBsBXhdGJAZzxnmF5Y04m1erColWYct9xa54+FF15/i3RfGhgXAH2eNc
425CvoE2uySPrawctxS2DdXvwhGJeQd1RHcraL12Lh3mbJxXnedensVXIdPQ2UKm
B9VoILuB05VcB7pGWPPTSUozxdy2l4cepQ5V2eNNaxB2TWMOsPJE7RUcUz9f6QE2
z+4MSvHSS961OI5qpnhtk4bHGM1uHCuOIcS5m9JdkWrYWL4K8YSnIZrGYEKRFbDQ
NoO3lEOd27jAy0xmrsGi8Rpc16FdbV6WZvGoGQUV8l49OxneQ3u8MkdVxRp33x9b
1zT0APv6mDPquNxp3qOgyCdhJrumQiNzxY68T5hDJL7+19sNyzxRMGFva4F2kdVQ
RG2PfnEE3go0V16GfeEFpVhrNNCbxGnd3XPCBRO+NvvQxGB+OzHa8gT3WkS3npQO
s+AG2vxtIOV811D3pkx2nvIU+FgvMZjDhCOmCeW+0oR/z3hbRYxC5OHvH6PUE+wo
rUd/PvJnA0qy8WScDjNs7LWJgiflsfiwFD3ILEB5IiKbgR1Z3P/D4dJeZfvTQKg8
xmpQltZRzKXRG2n/kfe12bOfrxJKuGX6tAI8aTA7Za22ztgFPqhJfWXcFMp7b8XX
wqGufpnXaFsNCxrgdByo0A1AKRWildZIhRyNEArNBQDzuC8RPihXHenSqSlkPb2Y
7Ief+bf2tvPrwb7mlhwEXbbfHMOji4W3Fc8sJy1LRNShV+lOzSwNPpvgxMx7laE5
4hlM3AYLkYJ2XClDhzf4Sf5q62QyidoNC7eWblx4NCaQUvHo/G8u1Zm12nWVjNcq
jSbySOZfAasNPq2W/9w2hiwOH7OnOOtwy5vi9BY4xfA1S/NL6bQOffRaAn8kKvih
j54AMqqzCOMHmzpcWRaV4+3CeVtf14RhGSlBIDmZ9qazbhol0MclXKfB5d8LFBz5
qHWI86bX9zZQy+WtQVnCpjlPkc3uGgdgPbQfP5RW6pTGNDKJf5FXVQfALOkdMLYQ
aZKvNqy347EgdjSDF6f+QdaWSdyfh51opJ+fswhGSy0goKV9m2HNIuyO0+g2VSMq
oWRrIvpR1seFeb93PYZ2tHpV60cP6gJ0+kEBJj3TcKeug5YfU8FAYYNURj+vqqOh
oUjMoeXr470jMl/8ouKaeDS/WBLzOhZ3nIQtgliXWVB54vcCJF4eJTSLrSNWSD6i
b4ybZX90IOmBp4546xiGBItSydY8JhYsnxAwM6PKDJ1Hh/UiTWczMoq1vTm9o99B
P5pFsOKMelNgitUlj7+Pmdz2qPR+SgogW8ooRg1VMA4cnaa7GlomVQdj2luvFVse
LC5ESHAXdwhB/I74sHeCtdLIUg6f1iMptHRI4xFxkjwM39BHTHmzngTsm8xJCmBO
KpESy8WYjdemtTcIR609tiyr9agqTbIE418L3PzS0D+FIsSApxdY5AhHYx3FIRbP
E8Ttwn8qRYgp2zZNublx16LbafYL1Cvxh4w9CNYt3EvJrwKxaKpxepscQ+vQkbiG
RYkuCCRy8Qd7wuW6aHoJ4Yh5156oXjC4YZuA8lp7pipFqiBsftLIe4T7UfbPC2ga
7uXZ5hiIqXW/KAEjlxrz8z2Nd4tA1637PFlNzZbZj7MX+LjCd4gbPCR1+lt8L05t
1xfFRoIjxKrjBMubvLtzxiON7mN8leKMC0oxD2ixMh2b1I8gE5QoY6GsIMXYVHpR
/wLnQuP3OUbMEMoEEU1iYSjKTw11dpdVejU8tEZEfYlV8ZQ3B7u92Znk45nSQcHc
XeoFgPiPn+UwzZvjzEApK2SgN1EypHFmdRDZC+p7FJ3PjwZb3qu+OcLFa1sqhZCh
egs1GqfadLxhU4omyQaQLRlQjVJjviNcR8h+BviqoxXvlAwERrJp5xWbzLmebsMV
MJ8eaCK02vbSFYTztQCj0YQ9iaYg886WLJG5AsWdTFQ3UHZNDp9A6zOOx8zQSD2b
x1BNrWbGZNm21WbeKiHi/UzfEhmFntXjNdaSyUKpxtY/L1B2b4kHFiPkkTfR+HF9
Ht3opcLz8BgUCYaHbvk8fuN/1eum+cTZD5abHR3xmb3LtnOf8JME10IGQlGwn01/
YLw9zIwwMz58J5HkaVNOxYQeUHN6odh7eOgHFPWW7YkqYFKTuCHYReocrkwYW1gW
asGJ/5bLkGwiujv91GnsNhUBajYiJKb+b5Pk3qsmRCSCeznW8CBy0VWePKcJlzZE
VuSLAo7Gnnh/rMCMdyqCjWQFZ4iMMKinIs1fcZkl4c8bf3zwiEnPVdDlGiDvOkL1
gvJpjpdRFL+gIP8f/S8hTQgUoho1Vt1msbcq6XWb2cF9/LnuEgmYUsNXXgdTADNc
wbOL8f7mwwc0+n5KdQE+xM/ibzbU5sGYu8lQ4UoqPT5ecShcJC+SVjLPbQW1g/0w
OzsNh/Ln+pgQoE1pE4Wb/YulRgD3OaucGK3Wp68p5NSGgWI9IPKQ0cVr7Vge/kX4
G34QfXNw5VKa4h9eCZmHI2aB2xbFhSZSxgbp9x/CLOlP2p4qCrDqoDKUGaOeIcGg
laUoC+jtS1peH5udKCYvrr6xtKdQNtx42CdVmXtMJ+AnHnzG6zBXcaKigj6eMgIx
ullvqQS92x38XrVXBBEuUxnt1dCwMFjVvU3G+cTM4sJhzhPPPztLAAH9FCprSJ15
EQv5epLypr5KSdh4BQ1j+qZpUffkmsqhDXVbQfVqOkZXrTbyL/qu2yFZG/g6FWSb
jD7bAoww54pXjCPh343k2s4U9ocfXpV2+PEL6gHAmFhF4+w1v+huC4LectKKbHso
xceNmLtHkc/ZqDBfOpapY5FjyJD6NW8cddvcyayJ8bG5lbau/DkQiYvOPIOX4ejh
Y0xJpQvVCwDiiX1w6KXv8bInFpHzsc41lkEhrT+MZlmVspoqHl53IjxeWqr/m9Am
SCBvsqrqvUajd9FrfYlWs+QT1Ggv6lMyDwH88tcROHJkagRIDKuduppCAlKEuxYk
sQz9tFsVIM/ekDsyD7MrALxQwDsTCGFp1KObnLm+D7AM9LcryH7E5hMPeejYi3NL
dYG+LPkmW2PJyDK0kQc3E0x/nth1Sc+EV//IUrciLxbPSkYLUrV1QhsSB0vc3ABJ
v0JFCcGahmazYl40ORRGZYG8LwRzIKVHS9yMR5qL7HEryXU0hn7HO8VehJ8Dfd9W
ghm9CYmgXuNqamLA8cwcG/1xZJhEZWgNka4cplyy939qAQiAmELuu2aVfj9o4YvG
T5Hnc50juQQbz3K2WMagu1vw7J33FTlJi2eMBqTfn6vRkL61KkBf1W5RZULPzjTL
xr00/pZkOa/XO7CMG4EVmb1veynWhFh0zyjfdzf8J0juqITOb4r1Iy8Ad+vxlzLb
+GaSHrOh6KE9KdnuyZEl1bNLRz14YCreQAaQtq26aXfMDsHPQmeSTBTI2qobHKk8
Mq+6FxWVzqQF6H/bC+kDA+gOrsjQ7WIU6Mt1QiNrkqWn6plD27S30MNWv62rvK5m
AL8bfnX6FEA59m10Xlgj1fGz0UY9nfhd4TRuZgzYdOKMXNrqP2VwuzhJJW+buqJB
iUyQhVhJibEyEthc90Ea6Une5Mcooyw1w0h22dQCJ9IWRvx03VBPFouwFG+mNA3J
tnnXOzlSuc2vexbJ5JTNW6g1XpRGXxalXsGOw5QX15RKVrbTqZJ9Gj4X7OMQ1mjh
s6V2kpXCxpZL5lbng30SF4o3Jkzc7DKQ57gTqmOHE47ZPR4+pa3iW7vRNfD5LCvA
Tuqf8pwjgI1CW/qOUpNVSZh19W1MME5l7f0D2HsG+N9N+21Q3U4Jjokm4789OI+A
SoQXVfWLPQ/v87Fj1fX6fqgtnCH3PJnnWEGU24wQQZF4c5ztroh9GeeSV8ooDT/H
Rta+FH0DgJtQDKguT+F9SUqDp4QB+xuL/2eEdnGDjuIPg0ZzeUC2SGjRttR4CNrY
a5v5S1+2ufdnCeKivwZotOiwPCuJfZeeLkmfoAE159wGVL73xetLVLatvJbSl/Qb
XnV54l1/cMvPZl9e4Ih2aAbyxHY84uJGMvdsuY+qjK3percswPfN306TtmfaNFUT
+EifWxtg7dSVDc2DWrPSDoFP1Qtnri0Q8JgrEi4bLsJ3xAM+dZjNcm17MTyk/SeV
zWc3GmRf/x/L4N+1UXUgcb+t5JwQ7bcR8bDumCU75JYr0HuPH+0Sw6iKZsyTXRdd
oaLtbnZg8fW+qyrGuIr0Ap/qOWTZKOe+nY/FJRmr69yEb+cpXsWeyT8YFHUp4wMr
utBP+2OLmS391uaZi1IErx9oitV/3l32a6w6WYVu7LQMcX6Swkp1IN1uRn0f1rJ0
Xf7i3gs3ZnndquEX5haHN+8/UCaT4hlqeLomR+yLjO0JCRcK5oTLGTcBnsRc4WaB
qtgBAtdcPVsV7Es3g+Q1dGI9Jk88GtgbqC/CG8zqFxktuYpWXmHkcahrlv3ykkI7
6eMJ9vPNA7lGYYkwaBgcW9aPsQ9r5JLEL4l+yQc5EBO/gwyFl+oDdO+Z0pYMtfx5
JDt2qOhnME2CuPSUFwEDXZgM48n2PH3K/w/kDQDDRIkRAGhbC6sRxI9nGyisxV8c
/7inEUGL1DQOg/hZiQ91kX51Gis+VRY9BQnGtUqTJN84x2xgy58r0Xeh0DychLJr
r410CW+XIqOOHlPlHN0jMvgCTUw/QJhoEmsnPF7pC1v0ghXazpXEB0QjGOtcSQnH
fJmYQw/q8qFb/m5p3rKNlYORpGQpHJSNHz2R4s7YNj+4xLmN8ydcF8S88rToeqto
anlsGqim6K69vLoQfb2CZbEbaCw3arzSyNKb+IN6szM1/o8fi80mHoV/qURwVKPL
dIlMJ+Gjk8nvIXLzKiXiMEsvkslNQQktHw2ZfdqKH5tRf7EDxwGWw+BC72RANyuz
EkLRBDALXKIedc7RTV4qOlkTIBdtnX/UrM11xjCQH8RBDia5k9P85BHahOQjUO+x
3k2im8SilyIvASEdIU0iV75D6TQU/38i6X9geYWRwbFrAY3YsiBJRDAOz04xOHWK
ucx+w4Mz+Ph1hnD9f9d5bThPP2qjzEQsU4wjzIwqEREIDoTSA/ediCMxwMzNZahf
Q6tjc36MijCtWsd2IsHs+F3EkKjiEcBq8xhZnqwSHBIUSl83rV9MkE/wq8WJaBmv
JWGqcV1zQBOMKBlQte48kGf1nDPrrDBJR3yn31O+IawQwn1yxiGYISKHPBREX5Tg
QWLYi3m2lC7ElFUeL9Vq7uR8RbA23O+wg/1YnyeFNxnLt8cfsQmyLkUkRXFnRZXT
+qHCPdCaNskE1oXxgyXHNkEAGWvD5qyIeR62qAtkz9z9KF14/NkWbYwJfG2qakFX
Or0g5cnvdJS/hS09h3GwVXekBSaMYzg8WkZBsY5Nn++x6PTol6gMP4rWy4DDfDll
7DjK4KIm6dgIrfojiUPIFHDNdHGYSTDCjgMGOXWK1xwCUPHzYLKZiw6RxiucbCCM
LmMB8KpO8NuWMa/tb23rvgsZnVawLtkY+KCZInDisv8c6kzF9wags0JSQV1YHqY8
xU696YSk9Bg8u/5EAieThRoqKPnCVq6EPZgX0ym+fxHvUsNjmbY5hveA5uobF1kO
oDUvpiVhqofK3wzBSoq3G/67lKIHrPp9hiYAvlwecW9zZvSVFSuDKFVEI/CeIVmg
ABvA8q5sSXYihPLmoSnJElA5MUTKtjdclG+ne9PgChH1YTV0rAoZWFIuLDKhVmtn
jYVrQQD3ChuzPLJybK+hERfxMZD+8paL7JrnNSgUNQ3ZUU1swLcwXhaMOaEx7Xs3
RZK9wq/fysCIw6RAIBpW15Vv1Bj4TGp5RYwsMvwdCw6NrdQeQk8x9L57CyqnPeU0
GTcWbHkPcbrnK3jan5hdT07wBheNx4O36oFIkhxdGuIkDVttXzdldbjBKfPd6oi3
rR5RDXXDTncFwCwRSfmo2XE+nHk7IulNUlIJOgzLBNyg3znL+oq+fKS1iok8r6KT
Nv4ZN4d4an07+C0WEtQR4LwmUvsXWtat8AaSoem2FbiQ/JCq6az1AngBoUX1/B4T
1pUagI1r+qhwJr+uRymhyrTmjhSc0NTQs2n578gOElQoMmukMHj3IHfgLM5JSBZE
JboLsu5QZpMjdMSScOxBwqOJqchs/187JXldlf+Ousc+PIqbwxP9714VrCZiY7JG
fHD4zH9V1o+XPeQIXTT3aPblcdulDhffuk6Z+haG2NdnSQBZKrdCdac/hcSXiNgo
zY5fK6e9nDZPknaytRIuE0A+lfHeKlVhxLWreLAotemp9uO5jyrJuwpuEdK2h+pR
GbmJHLKMVCFj2tiJ2gWZOiz7rcHhWFeIxgS82ceP5g+B6OJopJ6pHUb89BiYmq2V
yKKIfMFMVgv/YW3NiJKexVxnpvKbfHHgiRvCR9kALKBRJdnX3hVdUQjqgBYzgVaP
Zw4vIr2IK1RrbjBbyFWAsPBubFiKI9JyNtANTMkM+WxcarRlSgJSShhusoRzHcLr
EqXs8W1cIVXY8Nepn2Ybu/vePuiTw9uIgWmKHtbNngONx5FMF3QYcGL2dIVOybZH
y0/HZUYLfwytiUi3ZWU06fApiLiJ8uL67Q1A8UY07UjV+SP7v4uPfgZIIoQhXHBI
RbCp1Zyf+Jv991X11LHmsuhR4P0IWi7au9C3biyGx5BaMi+p7gHLmn5ywTZp91dZ
l9hpZwEPLaNcnYa3PpMp20HVLe9mLcDuSGGKd7QWdnbn+DKt8TcrsEE8JiCf3t60
gddoH/gu8478ikrcZwtTrxfEwyFpnUhORASxi0SZO/zuAJgGFbFRZ44GgeIGzocp
cFn7GEaQ90zPm2pKxB3UJ5HYPLj89Yczcr9eedG33t0ORLGTZXBHZawFYWcSADt/
4FjP2PRhCFaMckqmYevgb5fdfpze9zB655g3RTvXtuxFbalnMxVDQ2ieAO082ZSH
t6PE3+W8LgFdnCfnJyIuBmWy4XKJh7W5WfC6+ZQDEq6QFxuxIK1vc++awehmXFfd
R4SjacCR4PsV/FDZpXm2oKr66NZSXxTm6KWaWmPJCg9+3Wot4MWUC0bT25eWyRgI
qtE5RpKOyPDe655XU6BCbToM66hcBK0Q0rZwlNL5/cMPVHi4cEkZm+wDL7F1ugwb
9m7qdmUpG9A+cmpxco6pcFBxwPS5v4arIKOl83yECzQ9j/trhAJI58LSQctjhrfL
uKH+5vb/XMkuR8TxV7sMeA7h36Pci2KFkUkRsjmUEIZUAJmFS+2wEE0VGRhwghJx
iNgpa3/YWMhAJDZrCq0FF04rGdCQrIFj8AU1+61maK3LNgP/Ty2dhHJ2d1Yetbco
+ji6JzC+1j9AAzL6EnvTKBHeIL0Pr2VA15pFfgVCjnk9RgYOOQnW9Xh/Aak0E+nZ
t+Se9V1+/2vLn5lvbIUJnAdsjW5TXRKKdcTpg6PcD++YsAkXapigmeQEgG3DtG7n
ZQPY1LDDciVzAdhZChxrwWym9Y5z5yv2I9OJNHDAhP6VV2sA8r0rDL8cbPnl86ea
0T01BKwDIDwOb47kUBOJsR2Mmbom5IEr4uke+wBPTVl3EnwNQKQxcQlttWJTtUD4
Y4OLB87kB3+xOjjtqakdmln+IEVm6Pde51v9MI5Q1kG1/Atgs7zDM12rIUb5qDH1
Bl+0mokohT1qxNqnnq19Nrcds7z7X5L2GE0Fev/SOlN+5yVETMZ7urkulBU0fjgU
RLpE+lJ2h9i2/sc1gDfowk6O3S1R+1tct1i6dXIqjfmXdiISxyYhYncuQsIQUUse
5tdicyoOVz1S7GnesuFUWyT9rF1UpXjxIGB6AHVLoBNTii5TOQ1j3u4HGfzut9z3
Ofcq8K4IDFSlrftyqsembI7pciOwFwiqQ7ybZji7QKwIQXomcDw1Vht9rOnV9dDo
UU6xqH3bt46BFF0lj6+L4BwhFVPv5tZBCiN7fdgCVN2y96DTvcWHS6DcW/qVY16z
O6VrKGVxf2UsxKtj8tME5fUuv0zQ3JQUPWXDV4M18/5FbSk6dJTpNsm2aKR9AQd1
OxGJO79mO504ubIaM41br96/wWcYURliBV7twr1glhyPunwap3gFXLyeVHpMsVPe
9UiCnPpfgmJ4s2G7deOaaldcXj2qEzsXvwfXxlKzrF0bOuapAvZNOotbUiei7eyr
Y/yK9DCkTrF7FFOmOpFbjW/UoGVmg5eyitYFRrFyjBIzSGUDB58+SG5A2RfA105W
3HbN/h9F2LzuWDNcqRHijGPdEN1Bv0Eeg2HqziDvn6JaGGHQFzPKRp7+go621v4+
YDChqgXNq+hkE4afK0cfhFAHA/AJcYQNDaJKuQLqQI4ph0nqqQ5FIFd5iJKqxx1k
AWl0AoO1AqL8J0SH2EnGhRBW9pVoQ3myiaPG0f0nCHT6anaHCpLmCZkepXUOQ0h+
4xwXtkbnxfv3SlD5KwTITCmEFpinIzoMHm1q43EwsPDVFJa97OBpyG44AIMFXw6M
xeVzc15w9PdAg33tMov+fw/CgC3CE6G2mzI5Of376a/t0brfxHZnA3bhAtdDs5Ea
iI1tbI1KzXpiosYwWC9FjDQwv34Swgt3QNf31vUZbzGLiz6xCrSTJ6uhUcMVYvfi
MozUOkLMNIM18zTVvEPBsS80Ji1TduBXwkaFseNn0mOF9jo4B6mE53l+xoISYtp4
SWfl8F7dxER2E+jXgGU2ctW7/lnkrp8scyBg2DOVh/lbC4c42UKLapcJkaCjfZN+
l0s8leZyrVl33DQ9Hn0Voyl24uSSPb1tVV8BELJ+UwwOlzkAZjcnXKxkJJWYFr77
AGSBhzltciBG115VxWNs62itJpzDNkAWl8/Q1y+3VgfaTG+g7/W86ZIVtQgKQ2XP
LdYkZ6Q6rPMZF+d4tePWceLfVox9GK9UYelXJjnyk6Zy49QV8BJvYtHOrfvXMtMF
yagZx+1LeIuR5MMioOT+VXACj+YrSURO9b3/F3A5Dqv5AnBi8B6v+EfyKBzSbnMR
Q+lp+0XG/Og6wEtxHfxSjqOk5rrSKNtOJ7DsRCMqjQYy3U1XgmAE/W1NSt+3pZQo
pqAQQ75u5IbgJ94msYXX8HWjpeDq07p+esNDfuT23Ije/1CAihOw/CHTT8zB5as0
f+D/v5Ce2QowzhVEAMH9IDaPM8JOz/Fd7S1ahc1F7tpyJox3IsydO0sJzwBkQ5Wn
CrzTmPlAQR1OAn8YR7YEp6LqoT+fZ/NmWajowPLiDOEKmrBoSIcI2hYzH8NpVCoA
IaUQQqi7h3vreGYDLxNwkkPWjy8YbJG0M40nH5TgfQEmqih1KYdAHJMn+9zn+Lbd
9X86zRysP2WoiPGHT3zF/kFhte9PPJGyRLsRZkY/31ey6yTTougNXmpNyfXGvUGK
pCpfAg2exQM3nadHQSBGGq/PWwfOcAmSHaGPyrR/WxRX5jOAUlWiYMyFATA+b/Oj
763ZYcazXBj3YDOfynPNNv8jB3W3AGoHsfyBNcON7QcBC3i9c4P/oaFE/cKaZOit
L+e7Z+Ux1z4esLVDE3l2ugeP23iniomta40fQqTQpr42tSgW3iiQW5DChomsP2Cp
7GnJ9vsPuaWuz/8upAMlag9sDEV6T2viqbiNGH2PH58lc96K6zQjWPmedgLPJtRa
wJkp+T0LjcqKjEXWLO34ig8Ai4etflfk95C2Il4s6Z/b9s8K1BeVPyi25H8haF7s
lfWHXucHs9hgjXgm3tcUSdtkdixkPdXLVdT5QCafsQ1BLfbineoOxD77MZJWoZpB
2lye7GZyWf+6deBxyQ6eHcyZuXbsmkVB2tZ7z1TP4tZK7dusf9vzK7J0nQ6DeTGv
L2aDFgdO5MkZ/V6Zi+sH/Ot0/SkL93OlM3eZ9yuD7+11thcaIphnCaaODRc9+FB9
c85DlxCXYJBCb6xuFRYsz2ZFYYJg/ib+XXZlGGHdySyIByWH7pnVMw3e/dn6gukp
4cxG+3ysxvlazEQzpP5+Y9QtL/sE3S18ypOhWbUrEmmkLvrKMiEGpfDXdCJwhcLd
1v9SKHHwxNxJWmQP1OCW57VXvPPE0P79J7CPfb/n0iwTBbgHZseNTjUdgG4GerFH
rM6Ky1nV266tr/XwNDnTwkMDPPFZnKYU2rvL238pOUmSfYABUsX1lD/5/VlC0/km
SLnR0N4/F5Gyw2gA2ocXXZ7DdPZtoTldwttQqGoSB9kwyx8sg8yaBA2cjPAnyD3n
th8mb58f+OC9tGDIn7XmsKmqphMmu+3LO71ygxfLEIO3IAF+b7axWMFgU6dM0HDf
F/Qd5CotYim1N5juzYkHkayGiYfD1fAEmt5yZZh/dE+ucicZUDwvHMQkY00vhC0U
7nO5e2zyDDOVbQqzS8RX0dqR4tkjnfvrlBOpleTJFNFJWQj+93cRGZ+PPZE7evDu
gnHsvZgaUVTDL1fV3hP4f7jntfV7Zr0o+AuMHLxrfjCu5dAmtLdvGCU8MlpDJqKE
Sjgjnr3jV0WPzuCh+zv1d+Y7VoBhd7nRyljIWE/jk2DC4aJ6xXEJwyFeUr/x0YpI
TTTmpu1oP248KknduGlrQPH+a91Sct9OYH3X8g7zj89JT/n4+efniQt9CmR8KbmW
x8TbUxrNH6QGobe+C9USXy7QWBxqN+ax1tHCXmJvMCae7ElUvJWJvzxORqAlJ/R3
GuA6qQOdWteKeCQVtXf3jJ2dcV2sqdlliLciCFGCu+4XTmHxnrsxkGlUNFypj73/
0BS5uaJqrnqRbls8mGBcrF0RQLqeq7cmP5BEbTp+UMZvmHSiEVTogWo3BJ1l5YpD
7pqKIahjl2iH14tFRF2Gq2j1XoqAkMJ6LrATv8rUFg7nkJowKVMB/EXSwPvA4G80
GB71xijtDrH2g320s2PY2XOHnDTgTCd8aXwMlkua0Wy/l2tcqDxb6mQIkM2FmyQ4
HABJuPRNz8MMhwoFCsZ9EE7SsTSD1hSG+Xr3ZZdpxWgT5CNphzbQPinzBjP7mm0N
W08AKo9ofWLfNce3FhoFXFXFa5WF6D55PzPkNcFZqqvLCbWo3rd/30VhTWY4nTjP
FCUpXQXDYx5OPgNUT8HEqv/TVT9lDrFg0xGGpi3ZwDV/TQE6q9rCTxi/xJUnidMJ
zmex2UWJf1f06jE+PGpWdLOY9gAhrIixaVEuu70cC5Lqj8RPetzEXoYZD7KJHT1J
X9Ra18EnUjNY47V1jLQBNPy+GdnryjGPPh4HePBMZni6jaF9a2NIFD9aziADiceI
GNV3NZoC9HTJlygGjUXggVi+qSIO1N33UVAzXghoC0wZLfvQNZ/hJz/G3LW+gYkS
4P5blRdfS7a18mhtn3QHVKWihCY/oiBcJjRLTXZ+zjTQte2r9tn031pF34JP13zF
SMJqyV5Z5UTgNH5U431Rgmg1qi24826sVeiub0zacwC9nzQPZMEv7+ulyKDSBV13
mOj0oog26gDULfQ6hqnxtAnHlNIVbaFEovqO/II/pmBsBpdN20GhkMwMPHyJhCeZ
PEBea3sP/anCwaNWF50Qw0o7b5oMUkmLrYM1X40aPwFFtDecDTj6yRLLeC4sPouK
MzGNOij0dHPlFKFKMPaFYs4vaUHimoc+vaO23ocSc2OJlbvYdmrCm0RqzwdI1VDk
DkSXtSRa3Li4IBgjKG+MwlrfVc4VpCXgNQNAMAt1iNTEExSpsUZ4hDcsP3PPEF0B
3MCRqLs8lxiomYcHcOqz7ytb2CRdTZem9aJtemwhdc9yWX/wVUtSscH4GxoP3iUb
co5tt3BbZtg+TonGqUFieYZfczc8/7WhagzI81c6KV3JE5U1I46AOA/9zpZzkuf2
Qg1eUgOSLAB6zknfz0NxjhmQmLswk4XFJ5TfXVP6UBK8QEQcNKnCdVQMS1Hb/KqQ
zkIW7e8b+NQedSYJmOqmCCmx4R+LrfwPYqxK2fTOUw9dohr4picberABellVsm2R
jBkzznmsr8TcDDdyZVQoqc45+Fi+MGI/wXKRt2uT5P0WLwmNk+nDDcZkRZlZjpYW
/7Xn+vFG4lhOaWCyALXZnc0wpave9HqqK+wQJohe25+nzVO/sYGza+CIXMIpofU/
1IrWX2LJ1oOt3OnCnbc1KoVfSD7rF2iT8Lqlh6AXFEPQgNVoXaEN+XGQfkTj6KKx
k8bq5UuwnbJI+3HY+vr6gneAks6cwobK3SCHOe9MKzJ1zopJ3h2qqpBYThqbdpX4
UQcqVteq/RPGVQEBBqR9b+jUrj7Q++3iFvkSgtmSuQGlX9082+Zm1rEhKYcA/SVp
6sJG0IEL+mL9vpCVNJrbfUePpWK0KzapbE8Kng+xYeOTijOuFrxvMwgp6WB02qom
8B+2CgnTjcnHO/wSsQG3KNs8/2irvBuX5S4RejfMbq47SH0ox55J3OMcU80YfKlO
d5rYreufrTtkpHgARZoW5A69zGEvA3EWR3hel6auA3BHZcC5L0PtDxuZGsnpUGrh
lsjoUbJB36QySrpLOZIptFtmrm+mMHc2vXTK360xNJj1stUDODAhUXUb/mOPs5gK
HuxWE9YUmWRNGVKpiTkN5PQexvYGAfE3wddcvY/F8WLPfO80gBBc+ChatL7Nn+x0
wZGGaSUkmYlDvFZw2SU/ny8xGt2/wY9X070r9ZOAphMSh/KYvvgfdyyTWrA60hPe
mGJJhc98sc1ZfsfEDye+X6FFhS1hoTYAIONEwFPdOXZAm/WWme2L1YI6ThxMUcgS
fkdUe4GCFDv3FrXy7DSm2BqP1UQkXzUFvvpyAAQwzp0XbdRqFUDxHcz8e/JjM+NP
JVmo7T+mMGPTM1hN+Ex0hUIBgpmqpa5hIqWjsm1DpI0A1L/+vA4lXVE3kEVw0+Er
wKHGqg1pHAkSObnwXnvKEiZs3s32EUGxvkx6NRikx9XM86fREhAzNsXeCRSTXJ1z
PatS3eCkj9iiCtiw+djv0Yr29I1fC998MOL4uoqxnfNL3QcKUvjwpZ/cZKPq1eA4
UKRsgT7sQf5xm+sH+63NSIvXO+aBiqzu3nWrGYEts3TD/mTMsFbxZ6p69s3oJEQ1
nkdYahpAE2P0XZ8baYBJBU++B51u9tIjo439uFVEHiaq8C1qBnE9oCLIRti1vTBi
aLU+lBvxXbJp/n/JP4jtA9LYbvF8Utelm8MIVnGNhUDSWVfFGxwAh1wAjo38zT7p
EvfCIoYyIWdju3C6346nm+XEfatRkYxkSsv8afSF8r0wbB89c2TpB265+Bcz248k
D2cAIPIWWTD6KHQ6ZkC+FfvzLn56689b6OawCbeEOF5TEpb2NPh/ty5aNJWjzLok
LYceD2bZNpA/56L1d7Yfd2XyN73tRw7kCYQF0HvUtUFXRNR6S37S29wfe0kYGg4+
2IF1okazDPmxCe/zxuee5u67Osg64T1FXmbpB7hsa/F0YfgYM2xMKj2wsFzzgHod
9MhXUaQP1xZrPxNPxAA25TLKA9k370Bn455ZyrXf40uBFHifGYEdpVZEwBF7+9rq
ZSMg5yvPkk65+ii32NFEdgWBuLLGPMMCVasaLymwplNdFeVE06oOlct6QL37CTil
9h1wJoVt56YMrkGYifer7UaKzJg9ACzT+4IYjDSV3381Pr4YQkQMKRgR58iedGz3
MxWIQjhvV6Woy020fPTQhMGlm0Ha1AX6acJrfStd3j+4RVb0RuPXWjgMG0eJP++o
lO4vuNL+gDTTo0p5/8RZ74xXGWOTlSosgyapPinEJaPoCsNCUZVf16Gg+AdJBDpo
SQli80PfAxKr/HePuBYpOqJZbeYGGf2nRDvd5IOCDs8uBiZsjjBKw7WuBaMscP/j
7vimr73tQAxSfv/4dCaz55ieMXq/uLed3Df4FO2aoSG6iemZ1kn7jE3GOUB6Adqm
XyBSEgZKO60dSqYGOYKSy1k0OVEeKWiGlSnMDc2wZ1pwyfVjw298iG2G/3qV8UYO
j8TrZLAKhbFsQrR+R4Kc76QzcVoiAE8rmn1n8PaQRufZB2gji84GskM4S45sxzKL
Ag++xldqkj6G604v4kZ944YH80J4Hbh9BUvojbeAYc87AKSQhlgNPqNLXebDofXX
n6wrSSDxovlTNJG520tzc8d08d2TRjyJAZWccRl/JFxdKoGdinbO9lafJN92NNAV
hMlnGnQDAWVzQTuPollhEcZ6WaiuSCP41kVRTWvvfvx6sP6I8HtJqZi4V0w+Q5P5
JcesZ8zjW5MeZw8iFpRaGljv3K2O/DmRQEHXlRw4NSNJao0b9ialPbk0GgODAuYX
ovX5fHevh7QMoTfdJJAOr9QAvVz5vofoSG0yTU8dbCPk5Zl9oKbmvHWxF9agNWlC
ddcuExpI5NkuAgsMh6iPBmPKSi5m0+eWpc6zIvSnyd2eYbenlhug4YlaIjkoLnDx
IH/CoN12JVbQeoxmk6JINn7xER9EycPXyOL+EkuNnzyN8wAPXmdmaZdyHk49fRqX
wylTFjyW2RynjL0vVXx0O4hQbO7Li8NRBdnxZ7pvQM5zpX9l4xZ3ZtEvklPLN01P
zX+bjOH7/6QsacElmOQ4MuC9c96BoHWF19MF0hHz4ftS75g04TABKlmVwmf4wdS3
kR6tQHzgkRBS0nUHJNqFU/RCnx49Kn0N9UHXraqs8nbzHkrdGtpLNC4IS5gLh9S6
s3KKdrw7cSfUk5FWyc8QsPLE6y2097lPkflcX+GesHUoqr12TUXT3X/KMzJd0mvu
xtX9I6DtoOwbB//fnxma4Ck8b8mrZEPPq6sA1nUUgeI1xVVpHvhis57LsY0FV59X
elPauE56FYWkPGhSB71fv8MDOO7Z/K9bY34qdxtF2M+ykEaE/G2eCE3elIA8uKvb
/hMOBjO0kYcdxX18rlg2Ld6vBcnWOEqX+7bKWBjNUpC+1M/6U6gamrTnqcwiOu3N
A3AHQbiezRn+xCY/j70PPCV2Ki/ucXqHaTINGv5Q43mRWlRi34K4bxHwr9E1BfBR
ZjFLE2HhiV+zhYYPhaio22kRiRcJihlzfyaC3AKnRLaNaBA7EdEKRp1BX2yPpDZu
0x/EHjmzWTCww0LyoJ4to7ObdMX+fYwwkVqGTS19jcXPMSITFrlUb2o1Ezu7EWoG
M4Qj4EpeNm64leLol8JEKSDpyL7R8VZMxO1uSrjHpyZML1BmAfhuXYNKpNTRBF5B
r4cuM2BlLVDx5+kQjo6RU5qPLqn5OhRGXzE11eanaP4dDIMX+liwsWwbfnKDAqEo
uB6+dXs6nn8K5pCh7FWTU9ZAnuJWHirGAfX0Kg+kbxwcVfip6WhbRvv78BHgZE/r
xaCe+oM8UYx9C0s7dsMDl3JeRVOW9gi4zd4IM8ygf12HSoKqbRl3eU1U3xyDi2yz
bHSYNoMF7YKr3xPlUva9EhP2wdAQcaRqtsWqARPW58DWeKSCMJfQ0gSUMben2BLb
scXvKQ0LEpcfrzxns4VDI9EDPItSWk4yHgvt27ub5Q4H6pEdhkYfa6OsdCM6hdnK
IT3J4PgcmgE90vKnXseG6LjS6vj0gcmiad6NNlsLoYgDzZhwOGkKOqNHjP1WIEQx
cJi8fRi6xe9DY5Ay2ZdiGtxdoD+XLIR3EpK5spvUDBz4v1sof5n5dIBCy2O85jmA
UC33TtTBfu0c7O15/+SDfeXfQQGRnrTLojJsjy/WXu6eO5QEH5JPyycZqFJydJPR
YEDIzGCeB7lVryrShANfdKDuMqz1T4i26Zguuj9RjDFJqTOxjB/D6Q1LA7LTYKBr
POJLsKUVMGwB3nfEoHULgy6Lazr72egIvV6mAR1f8lSE2Es7zIafu3Z1yMBpxYIt
XrviUcOOqoLGS3PBxm2kSpB4F1tcHyHSFN/T0V3A1EnFpr0Alf3U3zfc3mfy8a2A
uidjO9vMLrP44zB1Eu5nwazM77NN4PhuBCy08YI2ddHFzag7Zp5W/04+JigZXRSx
dJYq+KQfIeVefyyxdBY8Paf9ZYr6hgI5uEJ3OCmXSmNeOt0WVXI5ZjcbWTMJM4Ny
lAHusgJRholNPvoGAOKm9JkZsJSvX+LYTS3qI3I7/1x5h9nOG7MSbNaqIYwEt0ST
DTvdbv50WFBEaLqHWvw1732+PGQp4nr51aiZNx+wf7HEu07kFNR/kUDhUIGDaDrN
tWTUC8MBC2oYxie4uqkD7X1/r9lz+M1dfeurTEkH0/tz8ZwcTzRSZByUK4zuygJM
HD+uS589kp4aEH+gyIn99OS/NDfrxlO4/pCLsfn0LFqDdeEIQOf7mEiK42Y8tv2l
1JtvKJ68eZxHEmyIVZM58lymfx1djMCGM0JTN94lTrt7gcoImp48Hs9rLK5y+CMs
XclzKI9LywOWNen4LBQYsCPa+vsxgpfQyzjKZssBoaZ3LQSSt5RkI3SIqJSfLs1D
EJaRE29R3sHjsi4gWlPbQvVImpnma1xOWuyp51W9UOtnSzX2b3i+0qW2CdBJ4zje
r3niGj6idQvnJfGN87/mAjI0BXx3j8E4hW+j7z8vUGLBg04Qw1S9/vDGsYoafX+q
EqsNNErr6f0mWo6Unb7lbX4Z68qcn2NMUghgoRRlABTjLFoXmZh/aEcd4kmwCJmd
36HMXvpgjXxTSbw0OHj7nmdqBJ/aCrLkxBcIZfaN8wqlYfPINf6HeLS0rRbkmblJ
hFDtSWSw5yuIQL75fJ2hF+P2A4hziw252QOd/7Fsbw5PZEKiY8JWLgmIgLZclWR4
nqGOQCRiuI8nVnxDMt+E1Htkj/7Bz6yu4A5PWdU60Fo0NaJS34R/JkbJwNB2Bdv7
g7AouHr7Vwy/W1k5fU2zV2UEUGGNNBbCKGfDAX9U+U6nYLU/+F9pA+CYoOxGtJwt
tnHiwOgvbg2Wrwb1Y3NOPcvAC/34U+ak0D1hG5uWcPOmyvI/w6/U6YKpAif/rdd+
Kx3rNAGXbG1V0fJE+c5SK+HXf1xr60yXgtEalj/Aw59YP2n733uUzqhwmBoU6DJe
DbKu56RQSNYO9cNK3tZpkENYLcgRr3As+Hw4Dt313JJD4ntrjsZzitubBK08+Nms
aZNboZyQSyT1IRe9WqOre6MvBzOey4SiDRxg6OMtfvPKr7NOGcI8g72ZmvnehXXV
GR67q/mSDqe0bP2aqAbHdh4rgYmeDcVNdx585960qL6DgDf8i2AovF6soHq5Ga7c
Yd9EmyyXEkUa06zlHw5KEOEkhUhd27Ga2wxCp5C1UQ31ZknA0uZIhZxE6+gg96Bz
e0qkoRQs+A5A2Au3F3pXPxjOwOFM/Gmi7r3vAfGRiqM48jfatS22uLMXuKxnpI5f
r3gV9hHx2dk4gWxpSjZZp7A2W/LC04UP4ZJK69GTHRYl/UIU6tLU7z0SbPbwS23h
y5s2hhjnB9rzosG/WqqG10qB6q7o63jHhVViP255YMsCLoPUkRVv1jPrK9iblMXH
zbP0kDQtKqCGO8GG7f84AXeDY5OvBotkOeSy4CWAGDcRzoc8R1f6pGaRUaOR5uBi
lj7eRgQ4W71YmzEPxSygbiRVun7higQKVTZ65FG7lccLGzwFFYwO7ev4ejdCmGRW
fOzR2siCX6bwqeDeKumUtYRwzUxMfvXBPB+ODYI5qQ3ZUE6dwh+Crn/hDvaHrE9H
c/de9U9WmFpj/tFfxB76w3eBiJGsBwT0FcRGlD77DmCQDKbjsenGhnKOuIza/Ymk
fQN4etnjLYBsUAV2D42C2aN7DPHWoTf/SOI5IJt9OBEkfbVBa2HF9H/9icVyVrku
NcdXQYJR37Eonudft32UA81+sK8VIN6UMi0Knc/gaS7Tov10XzYUbyAfkvnOnKpX
CBy92zefSFIsezIocJSYT9XBb3uqo6wLBops+19tek0Q44DYtpgzxhim86rv3SZL
Y8i65coA1fQYsQJYP38FCiqN14bhqARXErFO1eJDa0FoIyXsWoC4Lk6/dT5PTA+9
yCoLb57xmARKqU6KCT36u7zCNG5BgvwQAS4cCqHBGz+BGqKfimOkya13t+lGE4ou
buhQgUGw8xLd1PFU7WkDntNY+5gsRacQ3j3FPI+xLkUxUAQM7QN2tc9XbZmWio7T
rientzJzMzOF9LVn02EVzNh+AnO48vXxam78Poko4KfsfIaERPvplSsK7owmU7hw
0KFvEF7x8VwUcOqekqmhbWJ9ZVm0wjWNVjMH05DAbcf4gDTHDGd+3eet+BCeAMiZ
E8NGHIB+9T6IH1NPG/hOI357HuqO3JKqoHb/dpanMgKZKXZR3kbeOjIcptdcwlHX
2kQVy1hXZ2EMSABsVR1gNP+tFjD+Zhp4VX35BgKywGMamDViWHSlB5iZTDjySwah
pbJVzFBhKGyT97NKVN5eT2pziy4WE+aSNkMLYDhKnVHG5H4LuAvJID8O/X4lQ+//
u6kc+F+27bBXcacCfGZ/JPSJWMp9qbs58FE/EdAtDlsxOqXiot/aZ436vP/wWxPK
QQtGT6bktL9g7sMAegABAdFsmnufH9aUAiTvStRpPBIECDWIUYf53hjrVSCJ8dWz
fk3kg0bQ8t1YhhaMQswrvAE7cspa5CiPoYcQn+fNZnIQkosOzjmS+aNZM9FU8k0q
+QFW30IMpRcLS6d2D/5uNB1qd0Sx0eJlH/P1J3YO0dTDESi1GzPUXQlgMvKoKDed
KRdMEUlqWSrBmUuqonbBsQt2bmpJWyI4unUbnpQzqjj1ZEqNweBWzV9g2RYz4Hlv
snae2p8P0Q71NBpEjAhpEd5wOLHMlQMuvCPdDhR5bc/Fm8POZ8hvF4nZde2MySxU
RuWWrK6M8vwsk1S/GNDCaLaFZ93upg2PQRywOmYRhisgbktXd3c3a59xErj8Z733
BJoiysAq8+z2qrnbMrjn38guBt+A2QSckA4541MB9LbzhiRaKTw7+o+wEYlzQB7i
9aIMlmCSrgcAYMp1gOBEBbcr4l24HuRoJkQI3jj3uaWOZfQ8n3EFDI9ixoqJqbEL
Lmud1zMPwfm5v6PKOLHQOdxR1cQM+ASB7sqpPpHIN9NcYrrAQuPGn0tLIMI89BhN
nx9rIWRY4/REQU4OgNoO9+b4YiMUZOurCSooke2+89LnFG4ngQ+ccyLRw7x7+9Fr
DIoOu5d6yAJACTr9Mdis79PQXUo5GRpOf3AHJPBnrMlF7neOjaId7KsO3vQ5IxD7
fWQL7iAGk73v+Om2fD+jxz7AOyTzpNpiuMKx/KOGsCp970XUBL5TSwh631oZFncV
7pvwAUo9YKZVlTtVAOEp2XeXDfwAY7mRSuctpShtLD0F8jbam7tJjyo+/NGphg3g
XoHBtc0PCPH7HNdPgl1ExrmldW9RMawYPoDmgjxr9i9AfSyamlcrW7pGSGoZQUBO
EMIpp+cmTD3NPce6Wv/yRcNOL1EBmAQVZ9h0R7zNsOtraghdFTssJ+MTDc3fHK30
tlhkR7rGH8l+HOlGz7BMh+jsnXAFtNr/Qy9rJQRVW7I5PP8xQitI3NQEkr+FXbZR
zxFYrdfPBUjanAaFI/0TJrWnPpqM/Sx4/j73maq27I3EWZEczYK/5LQ//QUgLi0L
pYRDRMlBDf/Yj32ewziYGlFclsosTNBwx9WMJwLzPKnxfdrLV2lLizvzWNXVonoT
1ASbDc6WDDxYSydPYj3nRL9XWNwnYQY8Pspi3UqJ/Lgo5lFxT62d2Y9V2+ZeFS8+
JMLVxeXvg9Hn7amaP5HTsoyAYPv/OUTnppG0VPmr5ZVNi0BbmnG07a5XRbE3zyCA
kFBjnVbDhadPZk0WLbuusWDLxGdA/dqskghGUr34kYwaF2g/YZM1Yiniaq3jCdzU
raSeFsGouUu3Ef8y52x3N6XWMvNNmg0TMy8QqdFZyxwqOXXeUq9t/Xb9S6YUpVuu
83oLIOjZiW3/H6yRrFi2gBfMT48/e2gr9591pNCOpOJnBWUI3Zi4kCP+DLkaqY0p
vnLIrhuV30aFnjHKPpBYW9e/cBInYWtLQiiSMxWXH2QQA6XQjYHz0ZuLO70h0RUI
Sw+1MBGb8qUFCGLgzCvNDcAup0Y0fKRajYmh1MLG7qCcZ9zN1WTdjLWPyYfZrk/6
WdGK0sS+51K0Ccat5J85LjVe/b3wZzGGPIRQiNUy2h0msBC229Ju9jzskD1arzZ8
//1SRqqHVAXAeHfM1s/kWxu6eIKcqqLZFGj5kvDywL9HOuU3IirfKaBm9sR565Wk
RNY4yP2sgbiHPH62ICckknr+00WTNn37p+BGKpsifEpMWGRGULImTtIP5Qm4SQmX
mzPNyWUQdINFAY6srJOTmktjiK/YuIvAVRDX+tZNPNJNjgzFTV4Z6k0ZWczLAaGI
vSEqXC/a6LabmuzqumJzBQ5+9htKQ/oM0kCL+QlU6MW/qhcwN6E2Hx0jjMrw0HE4
8Y719T261s5+HPBVs7fqu93eAFe4ChgyD8Stu6G8Z1Xl03APNsT2Ue1UAvY6Neg0
AdyhvQCB4HgfBz2iv/UyHCm0MMTMRQy+wj+Qrn6ErHYLftBelmpBNA4CJqQETQVL
TM0XfKluWfOofhlGSAoRzx7468rKNdFzAOSf0WFRgqdtGYdwbtC4h1B68Iq1kqhE
JR9A7gg2p+GAfbsVLISFRYzL6beIEfP2n0/7o26rreZu8VbnRGzyTFoToibmi6MG
WiQaZjxoXFg4Clv87ThI8pxhwfY+GbzEFlA/+oIw2Osok1VLSc5RUJRrWgEdYxA5
hn5YkOnMxcR9ZWP74hoyveEylY++5pJSjMn8dpusqDmTsY3hQ/VoewaPJ+tYdjC5
UUeYcEcCCxTWJ6Y75I6dFPmEY3SZ4sU24muAFjIlZCRYUbHb/H83v5axJMFQcZ6b
45fKui1ePRDDpqImSuGM5vJQ8tKbuIYTpBLjqF2r29uFIcW1dj1SjUqS6MxScDxh
1frqGLLTCHUST+I8I8O4tlGJRGCTha362hhkbcs/fnsQdeWmGsSNLZlhvUCfZDlu
Jl7J0ZhgP/vM146TZhscrX6jnGaVfeXIi9fyG/5+vfhbE7BpO77RrbqqHZ69iWOF
xYsUWL7WsJbZURzoK050VrDbVryIWcQcJMfPG7aPOwIaJyqnOef8+P9pTFb/1e3C
HoHZqnre3pULUxl+QvsiloGrRoOft+DzcIALet5WZqvk3TRX+JBAPMS+a42O9S3F
guO/Cna2LZfc/Qy7qYglJur2tDVs9HEuRtdKafV+CrnKvYzXuAqs9ZSqnbRwDbeV
Lv+ZhUQMFe+LV4JAKQl6RTQedqbfsw+tfKWO5ErUviav7lZe8EBETSM/mpiVBE8n
uk9D/x/UMdE6kFyUXlzLOh1Zvh8z0B0Caym6tBOBHIc6+yTIdj9yYnXnszmF5ana
bEWfQXmjRK9ME4ETF9lP9y8sYqaInkTvrijR5Fka5YOVGq28EN5h3/D9uVY79xxe
j5gk94stZSa8t4exYRctL58rykDvS7EFCzYUlIiB+zipYM8Avvc61eovmuN9JtT0
Ick9oip+T2MDfAZtGX6cqD3hIavlP+MiWI8gLmo4H0PuncUCL1A066yzFtMNwcEC
ugfsCAHmKTeVyRLf5OCplxVP3Mx4RTRVCVlQL3Yss/Scz4lWCmpgZeeN1Q3PI2aQ
vDNlgD2Gsl5uuNaNzFzlKw9aaCo1lTnzFH31F463UHAy1S/ftTOMOUZKwtn/Ro4d
AQiQrJORYuo8q34nxaB49hN6QxKzoT4LSUMNvFBkWN0kKbrj3sPOD5Ae/Ndbys7j
4/f17tFNTUX0OV5DUpBOjjaPmcsQUXGS/oTKoVO4uAO3xerLXIuEgZxApg4DdOOP
m/Ew5GwN9xMQtlE3Cu4vWmMOEwCRNALD5QxLtSNWsB2HkOHcZCXkIg3bB995lysu
FMUW6jUDPI1Vohj/3LXi0iSMakCK+GQk+hMseLHbQjmBpJGoPug2U42AobOeIEQ0
iy3l8tCjR9/eV5ovMNLt9QjUKFC2MXq9FXw5Y/n9EDQmNkt7v+QE0yKoT8wrzis7
bp6MT+ioT8kfX9C5Sp+E5WrE8dnovdj6SejBpdd/IYUBaCMw+8H1GsDTbBGNkt6+
r8dwYeA4xmQ51eCfvfwfsiy3dfnspfU4ogp2Ub0gg1ID165dqvStA8fmJWGRRxtt
PeySBjbHYqk9fWVIt0XpDKzm5yJ1Bk7TCSQGbmi0fpz1IeERwUgnqQUmOjqtJzFj
B0cJddJIm2LgPz+6nFAzZ9bJHMJ/tQnmguA6MLxLX+p7iehq6rmj6RppQ1F0jEsC
6PbZlh27jsGudXSqLMK6n93jhZk6+2Mws+zE6W/wyEJGvzlwcNDmZ97JwUJNX8Xz
CUHqo1e5A0b3uM0nbkN2FMpYlDCCv05YlxU0/JNm8/hA+GZAxI24xv2pnv2oK72f
phaJRMQSBcveQWUqj7vvkImPm/Q/uZyyUaPCOpyLCBthV/OG1F/9M8nYB+LwY/ZX
tnC2+oZjoBaUZHkLqJL03RQxImtLMcdjo3aS/C8e1i9qMFGRA/ZNO/NZfnOqUINV
GEsUF4FoQFQP/jerBOiniz43slyY1ENM/yTGTh80er/NUIT7maCXircmoHJyyZEJ
IDssdgaWrf94WxlHUhHNBOw12u7rvdyH3ZYVqPF2gBPPt+5YZeZtTZhOtSPpl/5u
6R/Honly/C6hpwij1eUbaAA5VMfke4nMeW5W8XwMMQ2VpXAnevWexWRy3skwQ2iZ
pvdyzAjbxYloQw3lIIZf5OhA6ulne7s1zEDtZpVcSadVnrvtjg50DDKwjGMcAqIt
SAvbP5A7dcS2HB78EMuUZmJv/YVqNL++7tzsQt4NDy+9sHl8KKqyQp8nIlqSP/83
9sdqImknQF7+N3hEWGlX/RBjWL6GLpeliV08+MbS0KV5kOULuOwvRtyU27hzHLRd
7UPxCAB/WJcBNF92GtVxyoPXn8FAQHfRY2V7U8Lmuc1Mz3gRkZPuJ/5/YUnNFBnC
i8ths4U8l778ORmRHGIrOr0z3mOhRaoJppUf1/J0yddIT+i5Z/L5HxhLLkaC77a8
ZSOAPt4vorf6GzM1CpfF3aU6rY5kiTSD0u8DGKnAzRAKp6NSQNKQ3JItcJ3VH26J
8RsQRtpFw05PqGv8/5kvjMaKA9I5b9sYlzRiMLTX+64nQQ/D5403IQ73cGQekQ4O
x/QdoxBEcIOl7ajpguSBL4DCBQzHzJ7tvEGgyMm7jM/1O0T7eXOLiMW32f6BrtpW
ezFPBL3Sv/wA2cqIqVFUTYcIGFhwAGomQCdnpn7kl6F1KihZ+V+wk2lsuE07TS7A
WX3tl24r47FQ4m2QwNarbv9u22IX+WJZvDXo4wkUokeiF9sqklhyjB6JDimistRN
SktwW/kV4d/MrXVZ/J8Z3N8X6COxLdWkKgNnNO0s2CmGc1T9LiQl0dA3i1FdOQe4
cEu/dgtLqDLijZ7d5yuSALWGFSfUUcxtGDSgMr6K9dlPTvFcW939ohnJ2A/0XlgT
3WJguXbh0pZq0B+Eiaf2ixWKpOWIITJnACj6Hpl2x6WbLfSO7l1I8x5K7yzWDN2n
ECB8R1RSGRRKpLuTybmPOCwxOUMbfMQP6bKQrEXYIl89Aolfk4nD4s1uXyMVk7BZ
AOQSY1WQM98QTepLIX4aed3+d7zCw1wGgkGTLUiEcYsQk1CszfOrteG8I98/uXVt
QWCrJouaVGvVFrqS2CItiCWLHKLc/4XlBq9qhuszfbl+P1JJj83+Dknh0APlI79e
1spyJyFaJkrBpM7dyF6R1GCUS7d0jHFOrv4YMPx1N0xowx7klOtOM2CPHFRHaNh7
CPOl/NkwMnPGdW9wNxnCSWQbST21zy3+0ZOvQ6F5JL57uTgkH0T5xUjX0RtIe3aR
kfnOkF/CC2rSDXoDLEdlyWP/2dlZ8IuyFSGpN/SWVWajLCYvwAus8RM/FCTemqbF
XT33nTfWQ85i9yo70wB03KAW+t6MSDYOa9xbdZkxRsOKivHNKlrg6sRs2aML6gUH
N0BPiPJlslxfAigFrK8vj5KWPgxv92FsrN+M1b0blKcEwaDcJeop1UvOheZ6Q+Az
WkHM1nLgXjGu09MxxSq1SpArv5QlTwCakd+tPtRg8bWHRMGk9jIlqfHEXvhmy/1J
rTDW0vxC/N6yiiACi7x1ALfQGQzRxeQlFMAyaTPlPtJkqqmZTznMkGiiK8DvFTry
7gJBxH3w9PVLm8HlNcb1zEIaJMinxY9O+D8su/ctUz+NG2AAOY0DoXmlsypPGs7l
Id3qYO4cx27Ck6085+X2s7UES+/GS47L6WFbAGRHCwkJnC1NnvJT390r5ZNP2qfb
CdJxEiuJ8SDeLptcsRq+UgzFcDoRbrIz/2rvhxki+IPzClfgXa1PN0te1YMtxx+F
gJQFm5nyCRM+/VAO0KULU5kCx4hb2/6WJCazke2+YvnZnlT1MHNOcSMFhTE/rrs0
TRguRVXFPT359eRvONQ+T6QgM05mpv/7pYwGOUwhueM0ERQ+GaGAQ0J2CQ3MVvm5
aZ3vc2auu8yXgsoah1tgQ7EqxFKYmjnLWuUb+zFApDg63vTx/lpRmNRgPXFO6tUr
g2lquRVzzKAgq1M8bb1Pjp76UM6KKeWz/JRE677rSWwW250Da21sodaT2UisN7Td
QtgVf7/R+R727E76OlFQ+0U3IPzDl7dELc+5hCE36m8YMXFYSj17xQl2b4X3XRmr
NCWlth4QGkAD3Kz5liwMTqqKCiP7Cp38ciBgdC1lfga+uCNnTTlFJn904maqisKs
QhP+vqDQ77cP6kuCCKSK5d3UoQ2UAH+ZsExSix4xAKRLW4AXKMLZapF3mn1DofZ6
dQPOKJ4ZL+IdkblnVBh9PsXSD2/OShUdJfCmD38+kqaLKIx6ul53kk0jwmu43Kyy
k5VFS+GKTNC0+Ms9OBJLn0x7WQy18AO6KmXfFsEGogXLhAZ20pObQ36FhJIzPy+d
QrpVMr72vxMX1/cC4UWrMRt9EO6P5KiPsTOhsBaJrSM+kw9y7yKjgO6bOjw+amRk
lnaPCecyYcE6tCSefrWrfO4d8T47EJiR10pfp+SWG9D1+XDSvk9qzy6nYwcQk1RO
5LsegszzxLkRQNCF7nGuPgwQTdDh5zze6GUznlRhTw6cPzP5xhIAsCz34W86Pco0
/TQ0LGlB9L9LYEF2t6gFElVkgcKu07cF78f/9DhygrPgZYqgL0tXSTXIDHrMahke
zthqjyzya6mtQ32Jyy82bEnrpEHfwjnZH4BHnYwDEGe61lQhzTdgRxgJuaocu32s
eukVYBI5S7abYZh9SfpeH+SbK0oKSXkWO69kLVvLI/uDwIyZ3+MGAQWC/GbhqzGm
3KcFCvqV/LsL+tDNE96BBpZONWLYa+gcnzOlj2aZyyN0/97XLq6oRlw5lg2DrU0S
GuT+G+rTtOdlBczyr1q91gZj0e/M2kwAQ/mOPklt+OuWWifiD0yr6eJnFRneEObo
Omq7YSm08UxI+ENzj5YEKtngo+fW8ci65FxHAyiBgLMMXbXKBhrqQCQHhqcPEsW/
UxxvDOaOXk1lqmzQY91WVoeNRwfEGulOHReNKICb6GRzVtjKU/YCNnA7dPjaAlCA
L1Crz5jOpBzJGVKiFW45NPTnbLs8JQFrU2MiEZucVpdvvbrFAua+HDLBXbtKJ94s
clyZPBRNdq2EknuerRCBGfzSbdRt54DpzrI5IoULyIILt4DLNfAK4bZ5yE73JXHP
KxWRUpHo/64Vi+vfFBIN91fSWfsTHpzeycfMYrsjuL2MshRs001nzgplyRjn0dEG
5rMwLGv6IMTc0By9xs7OogDflT75oP7C3BqiN52ctMQX668O4VIaVB4wgfb9ZMdQ
+xnPCCZL9NTu0tOp/bp9+EOEMW4bE+YHgI052lGEueLR7tfWP2kYPDjczIL3cyGF
jr/eJs76oidJTT1fDTt6tx+RhXyOSXjjatIP69CpLVo2LB8EBYGoTpiKvV8GrqOA
29Al1YXavUrb3yAhDau6MoFDdXal7bCr+trXiNeO0tMQFdiRZuXIigLNNAUBky/x
pMnhINWp8prRYwu70l75vEUzvjMolF3kaWq3u84Hx5BUMjdGT2mvUQ4SQQtsYsKW
UENys+rtGzSlnJCoEWTzR94GVWkU4OU0IhWdnJGoiJzGG73+48q6eaqKVtWE3g8Y
8S6KwsFSUlTyxzGUzJRL6c7EKJdcPOqXPn0lJrhgKTciL9G9A2I8uNfgE6BUgnoQ
JkqAqfdydMt1X4muvbknaz5zdINwjuHjViARUpkszlq2VK8s33b0IF4+GhwYSN7N
bDBDznLEWYQ0H6HkDrjsDORYn7/HJrpwYqytVusjCYBTNjlJGN7uNxW7rtIDikbB
hyfOEi6+T0lHXKwuV41czBvre3ZJt+SwYNvWWfhb+01Fg3UjQ0Y2b2luv8PkVUwm
cks1IW7EOG3QvRM1HZNRzfXCMZVv/wqJMfNPbbWwyZ6fT9xMAKnRfGCcAH7v/Q6P
iR4NVt+pYj5hWyE+fTrEB7VEsbd8H+xmOerrCOTAPFBKPDbxE0H7bkHrtcKS+/3x
NTJXmqtt9sVkX40OqhL6Y1FNhtpWvG7vjjmytajbGwjbGSMwyBoZifI59JSCwT9b
CAZE101qalb5BpKj4iinsXIbpR3lLQypGwmCHGhrZw1cn3stD36swsIuEsT1FDVF
7dvBEmYSwaVH0EBbjiZN47/4aWb29paHzPaW7RTCB8fxy7IjsPTgOr432OE0yKl5
6yP4KHNROCvhLxRtdQRwSmxGOTpkZ3NB4I5n1zauU8be9QHf/LIpYAR+Ox40KLir
VIMFPjYpT6T104TMFBcTWT9H3tUIIqFTO5RFv+VDg5sNVhYsBj9JXmUkvbs1HjjH
Z/nEpZNd3ljJOpn3QCgvUgts/OuQS/TgWi/Z3cPnV52yew9lY9+s3shWuV09FDVb
3Py8sqkv1fdZI4NgnJLoWoH4UTPY1asXdhNReyKaPdUKLEpjNOyTu5dC016MV9IY
ZF3ykwVLGTOkqn1JowyjOQFu7rQm+rlNCWcTnVUusIY666lDTPhWErcQ0CkZRnsS
jFQiL6BCXzWYV28XsrFxVb4777ridkENIKPA4JgOLXT5KhWr0tQw3pWJpuhVUYtO
nej2zYeh1Pe8Uhyt85M2XMmZxihyT9DOa6ZOBlwPdldRX/hFqaUcfq/5SK4G8Ddw
vLAFGqDc0H4y4F4wRjYrjCIU5lOdGDHFRYdMPOLEu4OlSq7SxjE+aqxfiEzfOGRw
aSXqhleVudpTlvfgMrXpw8/P5H2MTojDvG4L/+p5MV2BGLxIvfi15QMpjaEBxyYt
aqtehJSlQqBALuJw2dRTBtklnu1Q7Lg1xTIIKkVnZC+aWsM4zqC9fxVOK02KuAcF
YUvq7MTIdSP9mmFyuUCgUimIZobcwdNNC21RIcaOd4ZnHYJpk/L3O/I5IHK6pzQ/
lyUbTphaQ8pZiKeEwrTcgai+DR3y6CnaOaPNf3meQW1hvgGXbbwOD0CWpmIGUDAl
aiBixnLCWNPoknFbOuS0S+Y/u4AsdJmMD5veCzmpP7Um+NjaH+5jmQebbxtSaFdt
wkKmtChW44i1Vw4Go6HT0xMYCuzCSiVMdQ7tTa2/X0bdcTZRHNth2C10btLHACTX
RHGxZPmnb200hMhuAsWfjoLGNyeNgGWrMuLt4lTI0kZglYOo6SLbaPs7uhGaFXZa
8FHiaw+3nZDJANLNFzrJQ7gOaXHnwdOk+RDlcRCSi8/3aw7D0Vkaih6tQXQjK1DW
jNoGIYBUjPWvSXuGInZNpkteGwfwCG6i9nVvJ1O3VqNI2cqu9yIYHqeuYHrq6DWT
+8dkOTg4WG0HTrGZ5Xh4qYxOrYxbPvMF5IOSt1cwcH4=
`protect END_PROTECTED
