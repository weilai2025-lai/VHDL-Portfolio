`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8tnuXcFmrpsTmjjaFMTGqnkEnWzsWY5OPa7rkxYsDakdGl+XkJ9+NQDHRpoqgxt
N+FEye36nl6YikkhdZD+GEOrEYt8rCRUGGso9ttvQFzrbPWzqElNWfqhyczsQyZl
V3xVdjr20hM11OjYiUJX308iHr+m1ktGCMDuPJ/PKpc6NoQI8V7TETQyYRpZqlnq
loPSAuNx1vLERk5ztM2dDcj0CZDqzDL9WvFYHWlcycHhlyxbUTFHgrxzoi6WBB2u
CFD6ZQ8g1EaekQL7kEWsDPXluqAIn61qt2b90d0jwXoU1cgVs8DYHbrjtidVqZKT
swAwFb5Ykxeyv8gv6BgUc94U05m8cXdvPCj4Fh7PyAWkcgXEc/fcFH90+3weaXpl
LqSWEUbp03poU8zOYPjQ22qLtGqbzj2GRfiUjKQhdr9fEReK8PAee/xU8QAk9Gwr
6fcDOfRGJsEkwMCpxK36CptSnWgAufKVojx9AKYqTqqABh2Hwsl0/DX6JizHhgO0
pOG6bjbycHeURCSTfJWnXJHdQSp2O2pdNLdko/ZUPfBAXFFfiHZBvqQCNU+G6Xkc
CMe0YwK37ItfuMGXsr0hBcUzHsRfDKc39KseTFCShocsb0janEaJKS6GnoWTF7Wp
uOhX2DVxGhsM5QKUa+pMkNMJs1ZAaJ0ymzdQhztifg3ypmH1MSnK0muhVnhNM3Ct
Gi/81Am2lZCpCDe6Nl6ceZZgDKJF1BokAgExJVPmGSXiTzLwdT3P1X09+ipwFTkE
vM7ncWSGe/MUaGqUe30Gl92doUk9aXw67tpEth6a5eZ+JFSSOYifDoYIdA04DBik
YDOxTTc4/qCtVBlWzJ/TJZtDay5Ft4ZE8VdrG+YF+MVNy3eMocxjmjuF3kFmZtR9
qlLXq/hMsnLI6gGh2lIu2u3kQPXDyGUgIfPBW01f4HC2uudu35jl+73kboez9e2x
hvOaw4VdIMm3nLU7Lplhxmh6pMY7MWuvsYODM6aEaM2Mc0ozzCpGE27eHDO8KFDG
bG4FWxC3q3bjJrD43v7CvnP9ASwg8UkNL5YjacYavy/3q/DLaP8DWNOPLC8IJn/G
+U0oB7gRAYzCVaS1vrrdMvKGW0O9s9VUcuvhVKkeoxDpkYalggaO4IjlYKUeA8ip
yICmw9yfOg+isLowJcd96OFPwP9BpbDOJnBF0ouX2aCGNtF/MEZtT+RcoJpLHJLw
74Tk8O1apGEFS7gG91NW9Ukc6r3lqnkncwUiHkNyTDdo/6J+pAUoz5Zt+ZJmJaTi
dzLhUBsh6vEuaVIFJFP26KzHsfK9p6ihPqVAMHu0Sa8xLxC2nEtG3H2Oy2+barLU
uxWjQxZ6kRJGq+fzA/uKz55qa+c9qcrx40jXd0zuinUPfjc2uut7N1x6LPsHjVna
ve0KH59HVImv/ZjoKV4LnJxdolkIm2EY6VwKwxp7UbmNM6Jou91ynqfe1x0yxwWu
ZWAXycG2gGrAYUCLJiISEF/of1pOA1u3FjfN/z+r+cKYWLw0eXZ3kvW6BoQ93cS7
dVM/tDspmyb2vhv9eaYnqZyH9OUHayr1Ftd5KTDRhVa0X7z9/G4tjj0Ht4pZCcPL
7uSWv/NVRLMj+HZF5yfxXfhLseXcf1/rzV6qEZuKoCF9q8wvRWndEdlB5FytqN0I
tu/XSPlC089O99nfHTVIolHU8jdbyT2PwxkBy3IL9Dp3eosmLfNAyUdH5hD0BI4+
jxljteVY67DcPEp6QhgHoWwg93Af0UQsBUt3+DawWjDt8KdXJaHYwqwqihVQ0zMw
uHG7i88UOjt4pinVFJIPnMDD2J2cP82fCSDb1pQQBXL6ez2MALpTuozfQOEx+ZKt
agAEZ4OBe+cPSQsZb9UCREfd77Io6ZreeknbQ4YCg34OYWbHeaUZBhqwmJshswW3
W8bvNKenh2tGN6Yw0cHUuPkFpkV/l5JwJevSjMdS7qjuu8XwBZSTuCjcRlR2GbMa
SrVmJElz1aPF36+r/5B9pk9Y82zREdXcvqwH1PidEddQWvG9N1eGKRrUUSdBXlmx
WYK45PRa2FOCNwDRJNHXeyd27E0CsPbWlXdAqaj/HIEcnMhmdwMkPYMuQ22zWfYj
kdlPltL+Mh2qsbrgvRuz5NuaD2f2QhfHX18uaVwZBQzeW9hrBDFbspG/ukR9S3PA
umvAyb7yaQrH+nZ4CT2iNTyRYoek3ikP8tUhw2bfv/BR98AhA5zEsACSbkKoSOgP
uN/PoltPl4Q/oD4yJsk5fA7MTxtm8ImT9xKnFsb1laKY/0pGHwwlbW1wHnbQoVxc
CzTPDj1bO5HQnSJgwkyO0Nrtrem3gy6lrh+wpd/BP7dl7BMlSrgmBLp9LmFzt8aq
iSQtxiIZvmIQ/KENzDTPDaVjYWOoQ5EPrGVbcWttBvi0MfD1KeYcLiDtmcQkrfkj
6Zl0HkL7YzBOfAs2w1+WqRj+GkD1pDikq1w6o1lzxcU6v7Ur5uftceDJrVx/B8Nj
QtK1cIn9MMO1rqADCieOnZ37nNtYJM5HTvaVrJehCWoUQWe/mhYvto6eUS69CV60
kAkXrnDc8r6hInK6ANiViVgWbGVz8wFVop5qic3+9FfNPCmx2nRwQha68zlHILXE
70cd65PqaoF4Q8v9DYl/zS36s+DTCQR5Zdg/7vcusVakB55JE+m0QTMjmSPJ7SQt
6dsq9K4QBXSFcoskUntUQ+A2ryBNMGvyGbCsZJNd6TTWca1bayhSVt/3/T2u5S/P
UN6KVde1AcRcD1ntVtLVXEz3HblFz852R8cVtJMTANihD4QdgA3LBDlZ3F+1Tlkk
xSY9R04JmiotRNlg1Os3VQeIikyZaj+vVmysHi5ca6EgO8lLmNFK49rclsOX3qpf
yYFYRiL3vUx1k3ATxQT63P+5Jo0Qqr578/j0nWJgQqO1eGYQjR7gkUqWHf/ihDGX
Mn/L6NBeUxP52BAJSIJoRsKGNunFJSVWC7ejI7frkQkJLJC2uUpN80NgaLingWOc
vBIj5lxIrTCjgjJUEA3ratHo7oA396QJsGbFBy5biG7x/BvzBOqb5FKMdjT85hrV
Cnxu7EWSikH4kxs6UbHuTOamTBHItr/H9F2toWQ9aYjP1LizjI9m8KwojMXz/whE
wibbplRjKJpJoMeH40XLE6zdpvr21Wimu8/Tvfhh95PonF3ItSNK4WyGKOMJHP03
by+G0gKfjWIr4ktq/0jQhmbn8SEJelkqNB8GrrJd23owWkn1lrGWbvemTBvy6+9Y
aD5tsblUkErQ0TkvCj+vbkTuR+fGoa+K2SZpN75tubr01kIm4iogxjBHsHZFf6JO
6nL4JoMHBq/epZvGOotkMWDOYqNgGHNlBBjrbizp/NuWL16LZwKCog+ECDclml28
6cbZlngXwnTdIX78gW4DdznVNbtXuhO8bBXYV/aPysJAvZnmsMwpQ2QQDWh1ae8v
c5qXHfBf2dtV/MCOXdPynsc80IjAxCNAYY/+4eqw0ZXKnqIujHP0lHq2J/rrvWc1
Ti8g6X4gjZeKLKkpP2xBg5yqW8EOZNFzHnAH6PSMYvlDTEz3fTDR6ZrH1ejFaugY
AyiEhRyKlfDRFGATWL1ea1gW6yAEtC+O6YPOnOlcw+bXT4Lx890RCRPJKnP6+6M4
DADyDF95VLinXnLZZv7SvYH8JYKP1ZOwE80/zr9HRIt6M2IyVMRGqP8ww4by/o6k
8X/7aL7Lyj9/NWiHWUD31z9jTQcylTYIkHUG2SBhTAk2eQ9Zkbte+Tn/S790Qn0v
sCHcAUC2XWDQXsgyuWGhtBN459PD3Nfz1P0lOyJp2lIhosTMGAohLVEqzrnczebk
ulP1iX5mzwt7dRjUIi/b0llf/Db9/1swdonbshGQ1iwaeK1fn2j/FFUbVsGmApCS
SfQycL8WFnfTnWfTqLKiiOP3b4UMeKiMEgYYNtTnAyjKxl9xN+HYSWwtelvz7gFE
u5VhAuFHvnMza1zGIcc7ExRF+RhBnsRilMkqlsRnG6TVxFlfRP9LGQXpwXtXKw5Q
yIlEUjgjRmw2XhBvYayvXfKzQnRAhGhL7aT0++5h+iqBbDMTEIqq/DfBO/zI3gIC
Qm7CIaBohY9RjNh+soGUAylD3GOGJYs/iKyAH+GVdb56Vx8LW8L2ZqTpFT8Pq6qL
G/V+absrHt7GSvXeTEwRMc2vM9ei+MmVTMFSL4CGQ7GYw+fCVPzGvjc+y58MR4YK
+QKy7SyF4vmx9vCuzFEjY+kz4kZHPRDBGxXQKyLieW9cnTpK47fDX5a50KfxXw+G
GPm6XUK8Uq3cb1YLhvgL8Eoydwti1T0AppyXdyYuUF2iCShyBNv+Igw93BlPkBb7
m7aCGBZ2UdJXP8rZicyFlRyPIeTXpBl50fsP7VmWgwzi1FUbHLF6QmC826uHsviw
xebhQQDOra4xPPN96c0Sxoy9ZC9LhWsm8hTeTZutN+AL2p/1SfDjQQe14ASQvrOg
yA1/LfA5DFBsN5Br0RACMSscJ31oTsI422ns+bXsVGOELteVEKBLiOwv47Eot6aT
ZTQKeWzBjhdtzVsJJ2la14fbLok6zJL4T69gJx8Grl/BLps842NoxL+2/fSqqYHH
mlv0A++Q9FCeM8DW+Xmt3u+fvdI8NPdQgKDNrUeWaOezCTBPDXZci+egyGtMO2Ew
GBQqPsGHlK4eQRqnfOEiPX/k4bU5+iqe9yEX3T4fcAKAW2DRDSGBhIU4+ktqDfPD
BA9+fxG6wYfdtU3F/Fi+dAP3bxA3V8MItsXzMgE6M6iAvuePRwezPLeCyoyqKKxY
Dd6NDuEUweO6/0WdEAG7YClF4yqwa4MtoLG1b/sq3/E9oRXADJM7udoaHBVJBe1S
fDkRbuHQ+4XkvoKJxI2a0jm4keRyQkTLyK06e9qAGscuQSnnKnKtcZLDaZ9CkhRN
5UC8pPPPkq1iJU3MckyfrBQFFnAvP09Ag1dDDdMFRtbXdve4yypUpNAu1umQT6TB
m3mtUABG+VRAGtc7js7xWf+o7oRWGM3ZHUFhPH2EwduWd8lGayUu9vK8rAU/Ff4p
Oaxz3CYRuD/Y0CpjwnnZLyRcIMkRbT0bABJb0k0ldcy7Zguhj50X9+M0+7eyZTwF
KNI9WwA3M2gPl3aLdjJ5RvfLp06ttNDeaVT2JB5Yq8mQpeK1a79v5VVcvumSuAyB
m381JMJZ2ljWl+xqyJgU6YRdp3rMzmd2qTcBDnryzRQ9nUep2Xu/UosSD3HjbfAb
KQypYeuxvbeEew8qXoJzMSFKKUbCo1iivR9J2MPZdW5b3F/QFswleK/P0QAfZqLq
JoLUVAOkHYL9r6Yx6dRT/FImG+dWC6HGeb9D6EIWt3jtYqG9Xt3FQHbQxOxxA2sc
QPfu4XrmGG0aiV7M3KOwGn6Xdy4NlUElYSQnADumQX+lTKiv0Guv7czRBrCUdojf
IQrPiLOl2sXhqjlgBtHVlNodOfJDVAw+/R4sqTK3HGALY3Ixc1Xnl9Co1FxY0iVx
Dy6Tohxa3ms3wa+owqKUF5S4OuFAzWFCG6K9+cJ2EtHvyxaQFLFHrUCNkmq7p/nV
IE0kzOjs94LUJKPPrTR5PN4k7Wc7vAaW2QC/BXL92Thw8Z0JtyVl7JDCplet2bbo
3tIqRTUNPmT101i6P37g1fiJgeWtKQVFFX1YYGNjBFw43cab/I9sPS2mDUZhqQvY
Mc/iR10QcellNAPaWzbxHkXooBPAXnCfGNJr+k4iW2MEOSEFYRy5PXigkctfH67h
oVzFEXBARMmulvFNVmuAFK40w9Ahw0fWVs/rsc4bvtIwiMQys8IDJ71YQmj9VpOY
yj6QOqNUxJMZ8ZKGuwmUoRTpb9fTwpOOmJtSkhoSMLqTs4Emxw5MM4VZ9Ael79k+
v0f47dgG5ey/PTazP0XfHGXGnl9f5kXQRUnVR6wurIRFg7thrOUJ0NF87TpPa4Sy
sWF6t4mXh9SePzlvqfAso8ZTxn5XEHXbcv88+0fUrql86Frwo9M3pqcltMFlR7Ko
MtsD9oIduFsLn6w/0W5WiwwEl2pePu4LGuywpsTztKZ4uwAZP0GUynoAL+l8WsVL
NziYluFpyHbdlla/eTfEXq+IttUsQNbv7mjPMk3vdNlzGww+fN/FYai/eSTYGnT+
16CqGCmLTHMWPa+Bp25TotjbQT/BeAv4udA74zFLQzXcQy/JSBPfFOk7YnOL37ps
86yt9UgjXmEllXuSKmU+dlRypPBqjInfTamJmkX5V72RQGMj4KWd3J30ULNhumjG
AVAJAjmobC/6ZFZ+YE8oCAW2tViRAD9Fa8/QnQf1dAGuHMQSOa1lP64EWVbn4e36
avEQ78Q8V7QPjwjMGstz5cnVzEFGxGYiC/kbRGY+G2AkakzbetdCxAUzryCWCaLx
UF2YLxNXsSKT1cGJdeueyKZCP1w8Yqrh16jwTXekGWRXguyfvrL0Ysog6gweca94
GnrpokdR5mjoyy2HYCuXaMRVFkUPjFleI0EMbTO69KtDrZmWEwnYp8TS/inoQuFX
oi3uhcDImsFjWV8IMT+f/UYvdgUsBODePoLOjJUxl+/UuX8WqrTKFBCPjq0gwyLo
HIywR0Iz6JExKcqFNa8iqe5ATyC3WkxjaKlBNnMNgTZX+2xnEYJySRSPt5ROdPAD
pAHhfznhlBNzJJ0Gy/8BtNzKK9ogdZlWHQV1vvaMZ4bOf/D2awUqgo/nWocCwB/f
n+agJIzHl4joPLdxs942Oc1Ij0LlGBZE1s0izXxLchVs6Rl0hIkdjE+m5j0wadZL
3geoMbbAIAJjI4hYfCwA0y9O12/eP0zBQxflN/GxS4fVerqhFwri4iVjoewpJrmN
P2TBVpvVw2A/H5KvWuIefiTeHA9pcFwdVsofDLm7/Jt7Vjr2WgjjWfZyUI1T7Bay
yfE/TmyrwNdvKHbPZccBD8DUckVlWBdBnvsWC9/KPM7hz5OIAjLFkSOKcVWAncBO
x52o+0vAKqnkb0pvEnJSbfdv0xtRcWlhh5eWYNvj1i/d3HILJMa/K/iSfB2mJpCY
rbue5scZbyZiX+reRPeu3Lc68mNQrpfn/dwom3wvmEZcVi6Ki+jJxV03H21pQ939
trKO6rf6zu1oGYdB46uOd9kg9wQLAdUogt7ULn4a5WISCJrj7MZwCI6aOVGbwB+y
yadrsL3gkhg5Al9JRDIvyHjixakutulOpNIxmqyjxlvsti/sHWZNp/3wVoy1r74v
TDfRiGLleISJY8pkP50mMaItUWZyvfY1lqP8Ono3QfYOWEUtTxNLv9xA1nZ1LM0e
1aLbGlKaZ0g4aG1RqOnCXtzgdAzkqbm+TRFThb7xGcLZqWS0Ji9F4b2+mqeOI+vz
WEwK1uqQBSdcTJyud/EgldKoixGiABRodO2emb2KvDfORdSFkpnraZJV2uxcOgBc
5Y/SgKViw2dZ13coJ63P7i3YNmXCHUjnGFMC7DaMee9UuZCI4qzVh7+E8Q1DEsO/
juzANryoWxFn3EAKoCTvalG8HUnUPeq2oeUVQoqjpcPliIfwG98C8mP5z953Uz9R
Mf4PFZS8OTKZSLxE4BAuV7mbsxSKlyA9IWZ71OH46fOGTyo7vAAUASxWq9/OGPiv
ZIK9a1vTto3r/oXDuX3yjLK0o3LJW05IjuZCgtaHs0lHNjOv43IOhwpB9ro6Imyh
ejeT0esbTqFPO4FiwX7xUlJKLZtWUuo/fXk45rf1CaiTFpC0Im8qByUNwqnz4O7u
XQH474p4AoUfP6rtMW/5gHCDzkZG7cdsxA/wFm0pplC8hFkZW1uTy0IyqXJtyPVO
9ossesJ+V/lcdzm4WGlNT0lesi+5SK/z/9EYY/xQp+WHnfdhraTdSaAde/DOHzj3
xM7ChLsjgWVtARUfA+qoXHInZOLmR1hVcuovRzUJlwS6jSv2XoPzAKlO1lm4XR5R
ZazrNhp0EP+VjdHjLuXo6SgG6loihdSn2jwF2c1GjWsHRLSrEuoe1zbTMMLannUs
VssaRzGthOHk0QA/sJn/g/tmzCWFbMf0QKQDeTwjUlsmBxKJbeZVFgDeh31557o/
WQFH7wwfKYcgDR257q5dWD6SHZUs3HNplLCMRo8SY8rOgbEP7hqBoklo4dCkYpD/
uppuhOPxuIK945ihTcWF+vM+Xj6T9IJffKBdawI8qRfqs/zFn8rClwzBzIDmOtUU
dEKvygZlCvQ6JbW2IO+uNdUlrhgQSIfNpJp1CY6jfnUp1x+P6ayK/ak7wahd7LR+
E+ZuzJvjIzF6fpWHomweMGtZeAstIomlks7LCRdCwzW74fWWw9XjpebXPL3OT2Fp
N4PKVFlO8r6AjB5kq4tyBRbDl4Rd4Fvd5sOISGcajnn/vG0VS2iyEVhZ40sJJmE9
hcbECslXkHgOQOMK7hPFuAz1Oss9SRyz8uF3MMKGatRL6marQucWAHiIKIfdVe6Y
up7vYZ+vdCWK6CN3Un970ZvfNgh0lnmT+dyaaoFVjTFq1q2z6NFuA1xViEJtTuwM
MVW7F0bDaaHm35etI3pcveUF4Fc309TedKZGMmvGvxDoTMIfT/HI3ayJf0z/iQg/
fvXIjN8d5xWJXsqrBTeEtu0XmbSx2dyl/3XYdTL0wHDkN11JJes1bJBpo8v6XWaz
DUW4Rkn0tp6FPD9UUSpkJDAGRV3dhFKHyQkVnGpmWXAm2zxpRq0ZtvLflKjLnrG+
o1ScfnGLKE7v0LODhGID4GKp/Rfi2lTJ+9M7wqGb0KvOdnmfgZ1nQfrHurtcAVLy
npwPzwvsLMwXPmg60OXUPWVbJrsXHV8jY7iADMufEr7Q7EZ79jTkhpWSLg5VRVK1
bs0FxkXQMhot/Hs3BQodsXiN0jdaCMTMtyRM9+JbCfS88aebee43EypX5TyIGb+N
K16NSBx16kQfn0qNBQ1QJxAFnvXDkQG/clYSIlcf9LY/UFb1vAMn0/MNaJgs4SdZ
7LspQuGhey84l7ev3OxPB7qoz4mDyeTDVayWDVCWkNH8esWX31ei+Qi8YsLB+Uew
yK/JcI6vMBpX2kaX3bHfqY3/utAfOZ7y3niKRckjjjI7wgipeTr7HKxQBsb4Y2+r
8U1b5Rvoa1fXcVFXjzCcOWEiop/xSsJaXoJkOpg3CrMZBtq8xZr2ezIaZiJzi5p1
wtWdkxbr4LiiGfmnFlBUxVg/cSAOy/rhYpubAzoe9WDj/P38GYQJshIOwnm1cg9z
HiojaJMJH+pejoVBCAP0sjTgLYGYhsDruZxq657MCgRHcJxn1MIiogoAS1a1n3bi
/HDkBny5Hu3DTTb6R2s1CGkLmUzfzDD4AcXSGDFOkAf+42ysUi75OuDLtEVM+jhp
Ove2wGZ5jEJTBQPFdoESEKi3sPhax3i+H+Prp7cCwAZrlIQPf/eIP+x7TjUO94du
ncu7iBsa35OImqQKdzM0Q0L3LmnunG9sBUO4OfD4EY8YSKyb1RQ08EaUoiaCciKj
h0N/9ODmi9k07D77O6Fc/sX/R3O9n1FXXPKpBv9l+hHcHiegXLSJL8t/cR5fV/tS
7LQrvV0OdZ4YpFoMJb3iXVHbZvJIMPnudJ2FxuiwyISQ6L29bPe/ZFohc6fcyy9O
Y9Zs5iJlkvbDCCos3U8J6esuZh5e5W3OufuF0uEHtgIDKT2wVdo+veRLyoIg7/e3
MupxmixHrxNSJbfR8O8a6lYudQg67lXCXSK1z3SGTam8yiP96AlAnWKLxfG5mV33
tsrbX5Hf9c1TrXljrJJqreXnOSG1idxx7EC0eZ/x/L8isSMh2hg5ocl+8BRJ0OWT
rA60bEXULPrze/QCsnITcswLVyD1EaQscB9l8sStHODuVOHoiidm2eOARwHiwWka
ebQ7kyQMcE4UCvoBypgfibD0IFW3VP2Q8xRFp/+8X+CTYUE500Z2+i0GVXk51oPS
PwkLvGHpQqaLSJCQtP/HTzomxnFI3+UOmZcaCvUmjRXoraWjANceoqvE8pbo7dY0
dV04u0QP6dKVfxJVu2g7XdNDHVdaUB+P5BDLIabRXSJo2QH/6KWlkTeJx6H2CuRO
BMgsNvxsjIOdlDj0zD8w8kb0idS6iKfjZqL725OO0thT3vBJVSkay1zH5H4diADK
t088cUpay6Bk5goTkoGFdKmFUtBoL+SAjJwujqGL3Ft720gh1SF7HC8foWNlOdLf
N0phWT3DfBgUeJL3bngMC+4NRabrYEtABmQymVrYYNrwrlUfwb69yIeapbBbneYX
SCXHmK6H/wJl06YY0fMnjFudGj7Qh8vdGYlMfeSu/KjUJEPlD7XJXAaZvS/Vo7FD
dPmTgH7NRzRmtNvpkxAaThGr6p/ArHsN5Y7EDkGB5QDs9WW81jA3oV7m9q9c4hwZ
WlYbGJIJmAE0OGEBOgblIbMSOLrwpES6EERPiEV2uSeEVXBErJ+ND2vGhYLrM7+U
Ew5KSLCjLuIlWuIYDW95ue18gfSlNv4DQZBZ+b23lAVF4hEiDd8YWnfYDR73S7XW
eBHityYxDCU8azyWVBW1h9jmk7nZAXkv1hNLqhTdl6sdjYNiksKGC8LPv0kLOPPP
cwd3nePfMSCWqGrFU5Ed6P+6PtUn8piwX/Oqp+Vl4Lue9P6OnWOiqay+DCLzabTu
isLT0AybHa88r0+pQVsaBRKipFZBWlvkTMm/nHpGLgPN6WFS9gzmdeZSufFbbslW
fXXaqubbCPR79E6pTDRmuoccXFN06m56m8zTygayYU/XNdUANA7hcW5L87s+vGwN
Z6SgyXN1nVoWkxWZFaP/o92ak3ScnX5kWryL+gkKZ9tp/OinsxPTQbOSMFWRS88p
KI+DNRftVOHitGSSLr7Uez+7gJyodYInNMaO5fz9k0FO4uEp2CzMaOQuhkQqPwlA
SlfgguCqMCIdABpQYwh+thSfJkoWhtNJrdD3uI8MziwOPg4CjJg+VQO1ur/GRg0W
deKdoBdC4nRzZFJf0lD4Rw9/U0xxFC3xtMNq2jK6wQz161/l7PQbPFywLaDxi3eP
pbT6lWm7SYWTPU2QUHxoi/SgHVP0Ebf9OdNbKc5f3ZI00ZVfm5GIaTGJtItPu83C
VzUdeVZpEje1UnhqSPl0eU5G+zbpoXlKImBH6sOAU3mBvO2wJW4+Yk1/lwIfwhjy
CwnuyQqN+ZrreCJUkIuXtozChZ4juE6BxI/Xu0sjbmZM12OdoFSYJpJusYE7XBMf
c5h8hFW3DxC3zJZPQ0RxqhHN45NzmpvB0Nh2pIQhHRh/bP2aVQbqXhn6TkENXOYL
pLo2zBdCU55aLBYmiVgM10pave+msmKzLeL0YkCjLTlodhiMu2ZpI4YPAvksW2nC
JzM8bz0bvtsTx+LkDwnCQusY9lZM9ZTNrelka2rtORqBbyW+e+hvPxeGxgRL53iT
/QVqdBN/U4H3e4e2w6nIvLOWdR/8oS4HzBXv9cyX8lQPqm/IxlhRKgKeExzJQKX0
YAD8ADXVDjnioE767C1hcIkrgIG1bHzt/Ny9LOrhlvpP2mpLOs9MQ2HSfkekqcyZ
vJzj7lQnhXAmoYQYxTwp4BKdYS/B4hiAo683AW/QzDbvxeh+KiSZetGIUE9CZTDF
dum2DTScWwqDlddSov5T5lfB2U091mFzi/HN9sP3WzSg7MZELrYjNzx3wj4rpvs0
GlMI+XFvia9YfklOqq5pkBkaTe8CK9OBO3/++Ir9TNZxlbyS6HVwO+LRX3GKbf9I
oNxzQmPPnKIpWzT3Mi8pbnED1OJ+oqTzCJDWCLHVD1+qp3C9txlwitLTJbwqTPjy
0QRsshq0z7XbCg0Wl7HS+4Qp+ubfmc+48/W54zUfslPCDRVWKkIoKz00GmMmcefv
G+WnHcbn+EHAc1nJr9iIIGajpEC46S02yyzs2sdQGueDnpeSub/bf/mD/GCzSIv9
zFFWM2jX4pROveXJCieVniuK8ebrMtk1AhBQpuulCkKF6ZJdeJqXOW8jfSthRE2X
bmLBN0lhjUQX6J+j37GxTjjXD7I66qye21RmO/sJ0NJpOi9iVU9Mklo0GgrEwu1I
wgtziOWyHGS3uN3sFNCN7w7z9/mDx5xcmXf6NBiDelSS0KTrZaWbK7uvV680FcvY
5NqdWu0vIAIZIIFRfqtNC/UE/6XvlMrNZ2xZ11SUHqgOYY8g2oVUeBOdNvdKNEmR
VpDVWDnsO8/GxYDzziM8VlHVcoW0bT6twVdmVehSTXeVyaSAkX1YklGI+jW52Hde
WL3FpwBrJEuA5DQv/KWbT3B4so3Sgz3yqQHCd7qZAiVU6folHrbAywn70+9jluQr
kWY9lfV4h6JEpmj5Xiv0OuvETYkGF/htquSunoXy7j/O850FaWsXH4e7x/Hu4tzn
dywS4j0SS0ULLjmlGsLMnUv3jOd+zZsxIJdzqqEIxmpZOqyj39BMWxQTOHN/qOYY
bTqQZYJni9EQjoWSFTBu7uBDvENvORcjlQBDTLg+g9h6X+B3VuremtjQKsBOo48d
bD3bU5pBHwTHgaTFbEL9dPP5tdz6Z90xoxvP2CCm1EKMQagTeuWmxssj0jlBNJ55
r4nAb1HOGYFxgAXq6V3kxxUhTU8l+bFsfBDzCybTz1eJylNtGGaMhE0K9MpzWzcP
ZMfyOcBmRCjpjI+VXHVnoHs1JqNzGJyoS5UOh8TgpDTihVoZJbyQa4S1bUS8cElg
6HSgAzfmXIafcJLsvd3o1HhVg8aBVTKw3wxHcOeQtsyzMLUQEyNyzdVlaWpHWk9w
2k2Kd899K1hi/PjK1pnaCg8ElJitfvkrO1BI3di4XLxoP/pGANd5PJuU2UrBVrxJ
H9x1wx9e7p+TpwD2RrOS6suSVkAIA9unkJ37a48tT/+5X9EPN7mGBURB04qvZRbU
imjA9KqMfzUi2wcA7FquzTY8x6QSH2nSDWOdepvwx+doYDpXxtOoud+EXPKD15u8
P1iiz9uaQB07WRoeoDFNtvtfz5IE0BhnZ7kDqeKUW4RyB7j2IZtG3mRm4QHmZlPs
Gq/2zJg3lXPGzOU4sU7hhgXjjnojsNwCCB1+OaHhtkR9oGoIGx+MoJmGgBMyGZkN
iqBc/WIrFdh85n7Wr8POvcxcYcKeOQwerfqpNWTmhkANxIqA3MhgKjsSMYS3veJS
J3KzD2g5SI+erAdc9DHwJuEqy3qptCTj1/H26mgJjHnNNINOqUOQ+OZaOmnol1Oq
JKx3ovGRRBxQqdce11CjnWlS/Ne4rEMyBnmUa5E594rNfW9K3y4yP8DkZ6mx+zeb
96DGoJaAKY6Kej5ZNJd1zTHK+segueukKKw7VMu38NjbW3x/zQEDeEcRNvFRzUox
PEwj0Ay602JXVUn4w3uOAel4+n0zHLqypgdC0tA2zb/a6uUs/9LyiPSc08FzpQZt
N2k2AsidfLmgffdpF5gfNC0/RqK7Ur72fg4NonAG5msXn0EBmxO+7TTB5umN+B0g
iUrzLvEhD+xQ1epMA2sBZpPvx/FzIAzqffoX1KejeTzkSTGAXvuBEnVp65IkWZYD
GisO/ESZ3Z3L0vfWQs5DO12u6E0V5jwza2ums0sCUiGuZgEyNvm1BAsdW2tv2rYO
L8PZQmOdxyy0dys1D0tHOrkWwJGVjuxe2bdzGzCFLEMYdwDHepkUqGZfcjqfXGyt
VD5YdHMgBKZiH5ygI3Y14I+Lu5YUgWsLfhBAJq6Ii1OrTrRtf3XcrR+7rN3TcAIc
KkZZ+Zbr0w9v4Zswyi5TusomWA5MyG5cfVVFApQjzNAq7n7gteYym3Ewcr9YkDn9
OhIftrz/b5yrYJvjeclEborvD+YpMq/EJfoY0mailHvO/9/A5lkWxA3aHN3MbEGg
tEd7d4irmD/O86k5Mr2EEGWnuKzNhG8V3R6/XUP4Nvl5MxT0WVx93P1POh91X1+U
y8KmXZ5dxhiDWOi+mbBmFNupF8rn63FyaE4rXNJDCSx6PjerIFq/SbJfMjRfvsAD
WYpE/5Of4keUabrpRU4SxQRajU97zGqHyiPZfL52lFI3BILL+I/7AibQWhItZK6m
Veh6S5Hp8mS1/TQ89BqXwq+WqVfBpE/Jy/Mc0dwMBGIsJ3QP8gUfk3/nt9M/IV7C
Sp2N6GSqotaivNLkBPCUEVXj6gn5+Ggo0JqdG+di+f5/RkyvpBFilA9t04xDkcL6
06PyfyvgmQXiK9ZecpRHoMcFlano+OQC6Q75005yhf0mkgITGpOsN0ZMAOaBWZpQ
AP8WZE0UVZ8k41LeiVilsiTLGTPcRfQN0/cXUNMs49kHbzLyxzeAeok6OzGDt/qY
T5A3ILT90XVF/GcNed7N1rFgru6trTMwiVhP6300AOPKCKOlifjCg5ZUmSdIL43F
ONpuwcP6qju8wlg2XEFVegx5M0Lt0F1EDwe4L2miy9PKRe905Ndhwu201xdqC65w
NjhATRLFw3CcEfSlG0MwTrKAHbgpgR66P6pm0mDHJYjSzdfaFfk3GcxTwkT8GAQB
NPRYksZTPS6frVrQoKony55dik8vDtIEo+3iIquTQXGKR8yetzCFrofaCdpYW7x2
CHLJQzGdb7MBF3iS0Rs0uaTZwFOc1/o0m0QhehZSjrqHyoEUY/K9UoLT20CPYLUX
/uoRh8TzIB3JehF6yDV8xQZQvaI4XSu5o8ihHQ/HpPkoiPPLqRwXrk1Vqivz/t7M
EOwnKsXhgkS8o7uU7XmpV/psXJhbLON/hM8L1ql+CLgtl9GfzIUlqkpEAfinw+tg
VwUYIlSkDPHbVfxdw1lTnMPBfoCiBYX/XWAVaNA7pITQMmvOxTz55Cu8YK2cpgwe
47MIrAr9lGpVRE2lXOJBjiEb3oZwCpNqp2OC3u+WwxMhUM9iTu5VPu0p/o21xbbs
IKuzeKQAOfFuRw3i4IEEDPQMUp+1OXnmYoGvmq2hybf42SSIa9xRv6qIcm9+G2Q/
+dr4W1LRNFlXSWr6lEHiCTEVCCDYWU9iuEtjNQRM+Bxj2FzvyE43T9Cumdg9kXjs
ZijoJ0rdvdggzgU19pGyPCyjQ3xAOgamOJq8NHa9DwKDrVVa0in4b7FYrn+XLcWg
gvCdP6Ue0UHUf8b0IuMeia8IXOgR05GLaRrjTZniyZ4YzMOplqQ6uVYnatSkv0Ze
NFvGBqgfj2PkVWL3RHqWAhWicX2tSwYu+0ZZjl9D2nz+v7kVVHCyyTmIFnT2vut1
zo60GVnqkLQkm6HCwEDyK4Bnyg1gnPsl6Xfyyb2UtQQCaL1HFsEy3H1TLoHANX0+
nxMvhEqCLVcI+UrNtH8IPhuVmoBjVO+qTqnRdKefXOSDSCk67+ilYMRH6R+MjxoT
dnJI0a49vha1NfHIkpDacXf4ElS49BxIDoynool4YN4yUK+FLrwSHlxlbV6gH8lC
vawcJ+1a61uopvswgeUWpOVwgZ+Zjo7yn7gU6ABd+7qOLGmMlD8VZDO4Ds3hS4wH
FuGyJUNtd+oerdHjlj/JFGjtT2h+eF0iBsWeu1CwKI2CRI8Q6wYhsgMCrYi0/g/z
uztAaKYBIlSGhv51S6O7UTYMDQjIZSTiPZryfn6cC0EpoFTdEVY4i7cCmvNV+nto
EsWvY/lBJpT8PtYnsnOEm/g163Oz35/QqdNWOnAFISeNvfpOg6uSFY0crGslBxB8
/+AXPlL9IW5O4R7Haeul/HCs6+ewrYN0MMuACkjc4fpL5v4iR5CJq2+38ji/7mCd
pikbQcZWN6CKjc51sPkT0O0Dvd3WrEhT+FqGDNRJoRrzaeJpoyeE/tHOogCdMDyt
OO1lpE1C4PDRa/LH2tUgUfq43wU52gsFv1s+uAuPPogCAnQqJ6phIyi1uWJQBHbZ
QbOpQ3AJ4MEXnpw2sU4/LCTq+v9OWlqd0rwnqjoy+ijt9qqnDvu//KzEL5fmgU3h
mHvvuzlSCl0GXnKUXEK9pPTS+oTJ32gIjK7Xwm7Md74HebyLpaXoMJyZUAUcWiEe
3KwtVEo1m0lsaCC3jX0GSII6ZYPsRaqLTGNXkxOUeNh4XhMo+4NMD8FP7FH11Z2U
qlK/2AE/yJNLjsQoZ/ds7Jma+RctqDOcVB89/Gklow+QJlSyf/UqP48/MNX8nqIe
Om4xWLLvpNG9JT5+9QHzc0DOhpFW9fiy/XwIHgM9ysWZBdvCCm06BDdf1BeLYuph
s8i+rWKe9rtUKzG1WvjQe3YfoOoUQ2GafMC9GTfuzk3DIsv+Gy+uT8NXxoRc0YjH
LO+sq9Bgn+sIQPL9UfPlYxviItQ0DGHtA7KGmwL2zDmWxcVH73O5Rupx9TDfn/ne
dwLt5Qwqm0cFwDumVpuMNJ1iC6YS8SoaPFGUPfTzOxA+7USdv8hRpvRVkvl6Yn00
tt2iUo/+RXJnSUmln8pNaaFEFiwjNUGxpPhlBk2NHM2hNDgAt1k6pb0gQ+yUip6I
KJqavfyTJf4sdbbJs3IbydzcSvFd3exJXc1jbkLszE2QIjPSF1jAYuG9Hzk38TGm
7Ka/XjyAMYWSJy9t8umTepS9DKhb7WCzj88Da0agwDPMnSj6Pao/xeoIayL96jf1
V2e+UzoE/PFP9aUHwHB332c9LD2njaJA0r4s/e8t6fjBCfR3pq7FVF9Nd2KmSfRS
7MxrN5OiiQxVG81eDn9DbrY4FAsJkuOOIo41xceWsn9CyGeAt5Aj75MhjpBOxuvf
uMGHWb0rqXFLhY2S1h+LIotbHQAZpx69ZIiEDyjK5mnM94Bap9j3+YdKUrE08/qw
CQ/Ro9HESok6pq1d+Lf51qUyuue6hYg5Nk1HA7hCSvoBo9KNg1gTYhd+jH+TG/0Y
qXboTTVg/+UNe3eZHP5EyCSCjTTfLMBUAZ32iF5AVtHUgkU08jGXdNCZWgHOpbPc
nYZ063lT5fZmitBBT/cii658pQ4QDPoDMjiaPKV7fEBUzCNnOsf/wlmN+8JhZPI8
rM9LVbFJCHTHvblkQwTLpi5bstj4Vf6gGDrBqw5LYtLMrshPQ/ak8h31OCM01xJp
hBwsTsivtTPz+qy1n7hdOCPqsLq6olLTy6ooMMQpWqvaybLOQM+sMdi+VzHXwwKY
soXKNzpzOwsu/Fg1YIAwwfnqSMBdwWchxs265xIgR1aZROCZ9mGj5HA1+47ufgM8
HagAzqftPJjM3hXxXdabR9uuTug3TThiOmqWTdgUXSvFd8LGkuCwad94m9jc1ucQ
Dam94M2QvRsk5Ndc6EmDIv0Uj0myrER3I31LDipVpVEDyixlXzNABctivKxUZVjM
7FnNYRxDESzdQl/4xrLtxqSIti9sasHt8ESllIuQrLSB6eBWLK01zWxGcTYbqkn/
W63BF7/Dfj/r7ai/fI/SRUtoP9OMWVaN2iesEjRqQ8Ius34gi/8Wr3SDttHfdg7t
qTJVNLsM+/8cPAM1CmRC03YoYCcNfUz8UfKor8it3SMn/CfrwJR0AcLHgBjRN2Te
l9NymplEQm1R8Fpq/O5b3V5wrOG3WDQTGvubQJJkq8xkNtS3sTTKEsn5b4EMroNU
olHrPJ1zWXl8s0voZkdaXHdCv0kKIB9GOVYZqsrFV9i60Fdwnks9robYEVhqkXGW
aZGR+YXNMyfccnQIrsfhC62UzwLtSM373lkNke3e2ow1OAgN3FbqmS/8xp7ViHPi
70uUjtzNSR9Ul1ZBGzjma6oHvGMPX4sunMR1GqgF5nikgmuiJivcZEqimGGa1c8t
Ddqwse4SXb1Va6UXx1YFf6uq1z2V71nGH5rviw25LrcXbwjkgFe3/8E7UdU5q88x
ZRiCuxoUNo89hzUYcXN504bqn8Fm8KIW6ffxPutK7T/wGpEBlY6AesTQIKsXsN0d
DFhALCfHxP5q6gyRUFfGzmO/ayapCwm37gkPT3WwBChEvSHUvELYHBqu+Y1QpKSL
qc8WBXOaNbS3auA0knXfO8hcb9Ret5TIiwoFLnsfXbHtILMHu34zuCHSJRyK4foY
qRFnhGYEmwHQ8X1EYazgg8tS8YBpDTBOzOQYs7E/OcFXZhdEog9uY71TvDUsvGUL
sZ1cagRZPQu6znuJlnqOioFKPgAa9zmD57iyi6AVaDgDVXFAX6XH2D7N7XbPWUC6
8o08VoPEEkwZEA+YGTwZ57vOXndxPinsAcM6Q57AjpsngMtaUGrTECqILa7XzCqw
g6TR/WEWw35I4QnlVqM3Nl5ZZCSlNtCfERjcJAqoBwO8BQ8Ij1Ec0Y40Dev9jjY/
VqNGIb2nXu21k+7icbLP9KT6sj5IvND6qzEnzFCe28J8Ey9CifabeouyfjW006hH
aL+bzQJqIi8xdp0XJmDWHVVY0+/bv24LV9Ti9OFqxCt1an8DV7EoKxVnSIdc0BwD
6yhujYX79rqpaBCwRFrGP52mUvAbhDpVU1iTJTx95p3X5GXkxAOIq6xFp8CeOZhn
hZi/vSa2emAuX4FMyPwpikL3Yr8INNtaiknZ6n6DHJOMPju/02+FilCcuFX49TFh
cQPmIuCngtP7PX30pRyjwj3/9tJvTC0T6Py9gZewJYxhJ+ayGT4gC2+c/pR8deP6
b3jZHUaX1lEORD6eOjaZplJqJN/3/mK7YiHDuhNquiMKE/dNNeQzkIUwoJagGDJ0
IyuTve7F/3h1DxjCOiCfzEU27YLJZmlYCsxv1Pa04G4EhAzpgv/L0/GiPTloDH4c
yqYQcTyEK9i2bt3DzOmcBpCiTMg2+ydCVe3OUeogfVrtcrJby4gbR2K47BQoAf+B
eTmjwExgkqfn3+WNkNJIvNNHa7uvsybGmWTNOXYO2k6KLWLrtZRye/mahcBF0amM
S6zunn/SPOe2iGyoq0Lo20Tva43SFUeFJPJbdKm3ypb3NHEMumFimC7S7noyXT9t
4JyOttY7iWbS7D73hqZUs6SEQdk3S3exvnlI24zs7X0sve8RihyW1adHmTSVIQCR
qzczwXN9yTFXsHGPwcmGLyLTLP1bt2+x3te1S6smpQ4VAg8P2lFNK12WqDKm4RC5
bcliZc1xxXSeeFfnhw2yZXd3x/JQzKIcmn5Deg//wPoXVssv6/gU6U/aEBwxOgdK
tQsSUkcma+QwL47R8cVvUFdSW7vvYkdz1/P0tMcR7iXH/3Bo1Pr5Ii9Alwzg/eIy
EZzrYPa5wB+o3uqFKhwDvF+w3/HUVpkmcXCjLm4E1f+fVOqmx3NKNQ+gyewQ7z8G
/bSJqeMy+VPq6iGHUWp6jgNExCt1MTxo5XnmpBClqjwOWpHL6mq9h7s38jDSfwYT
W+2S9dkvSFbz2FsrM/xwumVuNY3ACjiTqByUvu8Lg2/nvLaEqS/b1EhmJGUbdCMD
FURuIkh4/FTQX3c9sjBm4zem3QrK/KPArGwv0A6AwOUsAJbAxKatlRad4+zOXQvY
HyeAleu/cfbezdCzzdJgsVcmrIeKDFoeMndaEQAahRvPSDLyXG0zw8JlX1k0m6Hq
0KmJFko02HbUkHlecnxZQEcBQFOoRH1kc1s+jucZmXuC/zOpYzUjRLsRwG/b8HUg
HUZq913vQPrYjWcY5YcMixBf7VeWzv4dvAANXJ2Kplos4oSTDEVYGtJxMo9cJSR2
z7V9xgrvPWepNI8ctiZUzp85H+dO4hwHQvkd/tipDBo8+y6u9VraNy31c51yxteT
eW+4yAZ9J0/kkgVrbleIw3r7OystFl8eQKXXGTgMvz7NW5mRt1Ih4EmfszFjSREY
NnfYrTkgDHYSvyE4DCy+/xg3EZx+Vl3EK1aHSugBj8V/DHLqxN6f7ELe8LbLXpGD
p2WZxUFRoPzfdstenVF/nh+hVej5Jq7E0MaHYL/d/Rs1Ep1joFNK5INiBBUzY/L7
qlVFOAVt/RyS93rCDJz+/+2tne0pQsDLam41B/rp7CpaE/BYrrQKi2mlHA4j6MUi
pcXJnhXoK41umgpaU1PyAftqrjsj3AT9f2tJBoFvM15DuxGBEcGbNinzCIPdKBvR
AemNhES1Dp2QGOlTpibNaESIz9euerBOipFkG0UZ9ErKW6ARtNl2V1jou++ZtOO4
bKoegE8z5NkYmSlGKfTGFE89gHlERzuJN3Iv3fNwPVtxWaW0LTx7Wo5/jRL2Lvzk
+kjifi9mkHi1prA4dFrZYE5Y4DEbwaLTl2tsLG8grMO7KfMELi9i23QXRxpnl5GG
6M8kSalqXg13XCz4J1nT41dzPJhxs5TI8FME6bm/aZ78Udda3V5ol4MNXbyWZdks
lLirjyzE0q+3SxB/gDg4CR+7O3v/CVFmxy4mpvKPAyYdzRwfuiTDATPnbSI+Z14b
Sv+OkLginZsjhH5QxO8TQ0JPrxg72K/2U5byai1GWhDIlmEuwyRXzbM9OD2pFlJk
VOCoKfz3ic3yzF/KNDx9A6BRFdKT7COuNqVp79kLiijokid5UHQZu/lKcUHxlbNc
cNaKA6bo37ihfmayuDyGWLandJM2kZj5+qMmyVVSfNijuxbl7Qwa4j75Lt7Gg3BU
fYszDFuNn8AChnBKWfXnqUbIfBAlG8jE7v7NIUD31tjOKICJDDK0rWsP1YtghCxW
ExpWHpv7F/s1iKajkSGPASoBwxtMHuZpz+AiF5xIyookpdEnGql/YVvaBUQsgagH
16BFwBE4VofERtPFacORtaPvF6H9msL2kDaJfzgkD/RU946GUpNkvNHy/YSM1iyU
cOGs26STJoH6q1jzxh+CIkLHInbAATWzYL1XmiF3kUFhJZYVCY7TvcG/53ErLA+y
gs5AH5qcbGBWqS0qrl9JZtBPvQETYFHivdRvBePq3qM8UEdt5VnrBSq2z56nhtBQ
cpMQq+oKpzuVlul59Ab//0Mz6YkUTUxjmZ9YdRu/BqPvcqvLubCwbT4b5SQz+ykF
uV46FcG+HmV2UL8aw4pBZMoR9TEoMlVXT0wMOHaAtG1jLgq2r84OxHCX+WIij4v9
aR/kYVNo5NzyNdoz7fe4XzTJHa0r38sG4A8Gl53CeVC9qpL3bzNkbjrUkipjWtxA
V1LJSaCDStqCTWwunk3GObtna+fBINmcPfmGxy7u9mfrqXmYyrrdHef7aCnxkjHx
jqQ+xSZEu9VNAGTmxgzx1ZT3Ipd+S4xMzrlNg6b9ZElrUhwz1r8kPKhKmflqqtG5
KRdK6msH6thuEaT03J+IFQXhqd+gCgFf7WVS6axn0IDewSYMqQTRG/5E6LvJm1VE
laZhxW0qn9AUk3FWEDzd0vnIQTvsJFPn8dlLJzvIAQSJyFD3NVpyAFojUWAlLX9R
kNHY3nIlH/CgLQBoJ0ZsoHzA0NndEJF6S3m6jPUS6wniocaouFa2algppTdqoNlX
PdHecf10Vj2Whvt7Er7zk1eqYaBfS7zK1WTAdrbB3RdDLiY8gQiFkV2FQVlA0Xdn
0OqxXkOQ1+uQa9JigcUf0ICsNJQt+RpWiKGoZROV/kdF6BNytAr/kGYedKX+OgJ4
92xChZ/qpaiBe27rauQku4mKkXS5cRudAx4njwaE2uTPsw3OsQ3NWWqsrCwC/r4r
/jwnL80C5fc6bJYZcAVH7+WBDLrfUi6PfJG17/i62iQLRMCcU7nTmlnnVAeyS8u2
wcxyyKDaXnuo7+Y8dv+iygM64AtQl48v+gSUhGz+bLIJS3Sy+bGMhu7V4As1j1MU
Y7njfOidDc95gmXg3XwnS6txdwhprRPauhoMVl9t9itE57YeS4rqcZ9BzUlyXH8y
VDlb1DPOzMxGPtMNf8Ngl3ZlE/8aMUcOZmybDniBvOMjp+9g+FgzZalXVXQ38aPb
BSgAZQqtKh2lBkb4fvtNQf43ct8OeEMrcgcUX5Hrfg79zKKFeDaNa7i+LXw7vPGY
HqKZT5Ah2NXDn7XLIx07wyLUD8J3TnH3hU9GRqIJuSxQLML8A9fjfWHJJTZnN0y0
UtEWRfinyEBn8gAZ+2MZULbEBmymn8h7ESPFKs1fbV8CmglLDTU59mKE5y6cROs1
cBuSAwR6GTF4gaaoiVsjijRHuC6NoMKEK6jYWCYMAk0opTSz4wiBmI/HeBzAdmlz
5jPpmx1/zenOtCixgSQFKge4kZLUYOzAgRyVo+LCSuVPvxOLIaRfXoyvRrhLGlA6
dKclOAYWx3StXi8rd9xEClYAYBxyiXPgvXdLbRO3thd7D2YILRxU1zfDzE+0wiAk
9FH4EElNUcZ4BlWDcB1Ry9gRHVnpZv50AoW43watoOXnMcUiuWxWHrK/C0jsdceH
N+WdviipTL4eJXXxYyoCcYLP31U/5bC5QkOVDs1ViSgaJevSs+23kUHbihyNHgSH
ZtJn+hBn7uzyFBvG3fvekil2hBglO4REsErv5/2viDhtANBPjaR4toGwn6yvdeWt
R491X1Dp9fWC/EWzY9Ok3+4N8FxxA/dE51hsxZ1PXzKZO8EhjmH2KUt6hB1BcQK/
g/bimS/N71dvgkQThi7b+7Smr++wcEEH6ryBwbrkn9pKIhLbG/Fs3ytwBX6P2w5Q
5F0H1B5fYtPsv+ERaRdOk3ae6FHyRdXOgBwipbsLWhtFsLROYUoLFWmdgiBA2vbD
TgF77Rm2TnjKRMQEuD/KpU3PODDTON1TK1Hiec7o7drosi7Jw3q7AsmRBwK5jGI/
Zsfnfqe6OhmDmLC2qe7G4+J7dVKc4qQjuE3tJk0EnaOOfD+LFt4aKhV0pH6Ela0p
AAhm8HwEqj3qxi7VpK2wxsbMno+7bFanrOGoiGZ9LhFNutBz05JtJqw063UuqlZ6
3d/eVE83PBjKc7omdyS1JoSN8Lqcris4wex7NszqOqYIE0gPxEAPq7KoVbFwLHCo
7d/x1PnGDagNYf5KB95kvpKyF3gf9Wcjip7yfYXNp+R271J3RHyRYzJMvRFVFUN7
D6zalhpSCtMMrHp7/DzYmLbZLU2go5CSqqNuBKNFeZ9lp09vkQWSMvZMq6TRk9Fi
s8pAcr+313F6qSr2q67+dFfxclRb1CwsQ6uDmFyaV8cMmh58LR2e2jKwQh40NHSf
i0sGT3moGplptYz1nijsO4z/J39XwJTkWevgjQN7oRXlDHJNDYAn8N3u5V2SJ1Gw
iLxgDenju2kc1YLMLfBBfJyFKeMHJyRrSdkppe6d6Ukoht8mJ4fI4ROM7I5z6enz
9hjg9e1fKkW7ORZAbR0EwyvJ78NcXcc7WuzFnofNq1L8uRpA58/xDNWFW7QEj36m
tEmo9JsXfkj9FCMB6WCL2zyagNbVxdHu158S2aSr1jsxwxsqtjJ3H5kwl2wPgrz1
aHIxEF09zDuLRPR8juRrCKaYExP5TBTkue7RAyEUg5ZsX71HsQ1PWpzL8CXwx0mm
jabGTCPnptgzJda3A5A6ds+o8jvlxryAwHV52zVB+8ZA7xnZ6+9NnPU5bW4goZfF
e3U8Fne5HG9TuIOIirpqKwukMkiO9jbccxOrUt3pSC4715AmYVxWz8ClGp+o4QCV
fjRQg+hwAGp0UaUGodtcKB0V8dIqtHjbFQep5d4tZKybNjIGF/g+E3BbtEOoMeZX
Ptlv5F41+9B423kOYiFuDh37afUNihN3HGz3kU5ydOBAoa8dSVOHnkyHtPkRbNGY
fM1zjbGg5BKv6RaY9BXifTGUx8dlCDN3z8z9pOdqE1bkQhadQ2aTWqmHT6WhfMut
sMQ2ZJpvToBcO37T7Z4MoMyPII+Dh6fFaW7m6EiW4JR985qFY2Uwer7OzfreLWQt
Dt1wR/R5eousfwEUFkWpnO1ZJqvItMW/KNzRHMDr76DXuoliMjCh0uLxQ8jLhz4r
OexqF2X9J0ZmUzM30ruLu2yMSuj5m7N81C6HqU1M49HQCdwIiFO9NTz/+fmfKkCd
zg8RXXSqFqkHocgHWZCR717lt05HFXV0Kl7DjjyGq7yLMrlO6dL5QvCQObTzELto
gAXHOP5R4wfHL4azit9NcdIlA9MFPxBx1WJ62YznRFOXeA5Q8UgechxHw9gG4Xe0
KEPemh49gILUKq7uZhNYYadU96Tu8NxSqQ1rKsHE47FZqYxytkfzcUqWnlhxC7AJ
FXTysQms2nY8cA7HHIv6re/zRUi3DBx2QPGoXjgt6GUkvfV3aNelbXQ90dFgCxJe
JTvm/Q1g7dR1fGQAY1xjOX5J75jXUZGPCSIYG1NMEjF77lepAjcAmu0y+57V99so
80kvQEayu4K7aUp1huJMhDRT3veVh2kV/wcqmebhgxMhkOa5cWXUDi6NPxAdbrb6
r5U1Pmm0EfmhA2jBp95RDI/3UUTTCXptAKY7iivcBvbp5r4FmiDp7/it6xtxKe+C
/4Qc+zvdxa6WKqUompCkyh++W/XhTLXC6YVAZJJe+Ckt6c66+9/BTJTWfSRH3tD7
PrsqbnFQiq63cG+X2H1rRttJLc+uVTeaOyQGtqMQZrkwvB5D+eEgeKeqGym2ohfg
gfz55/pNjASNFdQ1jJuGBqv+cF4N8CN1Kh7YFpa0KmYsYSX11mZc08QtJYgVq3Ee
dOgFTwus/F7H2fM/A9WY2Ulf4bErqA2+S45cxYHmQHgzEzuzIgnQbvsYmmjmhCWy
QGKnkoEZeF12K0cFESDWpLQFAjy7B7Osf5OwmYLp9NXvEEn6BugpGALju0XKjNuy
y1AfXceqLa0F4D4sy83U2wtN0XmbSu+01QHQOYWp6FDTQOJ5y9RgqWs5iLO/6alX
EU2E+QbL01NvF1p6I8vPhEVdIPKBCzQ1O8LV7IDF/v0fCNPZENAneK4qqOnFJDTN
Ih4Cjp9f4Cvc3IvNlvcHJxCo6Qv8y/RPDaR/uza2l6QZV/Ytp4Bz5FfwxsVqE+GW
K9qOfosT0kPuTQtsAKpDNn4MKSqea3YM0reNPcMJeRIVf+bCHlQbDPIzqJLGBo6m
W9balmufRhrMg+fy9WK1SEp3D885bh6dt8Yw67OlF6QWBTRY/fYkmu5P2mlBjKaW
MmU6GAD/JtEw3y4MXtBmAmEW88KhmXQ3aukxKjEAkO5oIg2Qtt6LVKkBKMiGoDXG
4wFVmbVZ0b6xY1VLMk9bntznd84FN9/C7fyE6XvCycRBfHYwdrDkrdoXOjxWFgme
TVPCUUpwhHCdKtVfcg6j7XwpXgU8UfQg1dXigc296Lvkbk+UR+sWo4R9xTx8WkD9
VDDLokGJx7WFoskpjS1iWmY44zH63BuwJ3nDaTBZ9brqC5Dd0S/VgzObmF2wbJIf
Wl0DwC1IE3tOzWCRzv54pEHs/PS92vEYLaxMTYWKdXAcVw7nMMWMFky1Sm2gDiET
6Dswa2hzTUtcsDWijqf6anYMSX23IfyUu71yvvGxc8OgZWn4MuX+JM+nzry8b0+V
FBhBTCIQ2L53M+Y8tFs5qz49/kWQ2uJKIuvIf4cYDV2FcvMQ96l0NdKIUYYC7qcv
P1c8NNdmqZoi7iU/nYAATWWl6RpuWfE9qzy+YbXSWAEK97boXCRIA3SB5NzHDsTY
hmaEW3Qr5XnT7opz0xnLNppJMxeLGuno/jc8dxF5eGYTddxYWCmTufHUVD3lCuwF
iYNVFQIKObID4mjdo9TSb1c8hxFLplpoVaLz+DCwqvPAzrnb8PcNP3GPyGeE/N5s
HS1XRYYLU28+Fiy17xQEdjlY0pYxn7ygaFh1VjxFYu8ZbN9qYfOO9CmZ7WvksSha
98uuqUpm9Ou8jzJw0S4TOLULIiOx+2W6pRrYf1hhpA3nSDVdOk9SnMGTrrN8dWVV
Qz8370vvXqZDS9mcymSU88G9fnxSbuCWL2TfD74PBKtTT0pSLDBd9n2F+pjHRbBq
Uzhs19oZ8e3iMRYbhVkerjg1CNPz6JOo8Ecv8nioSa2/FTwURLDEpC5aRzRP+bq2
kAj4cl1ZKLTVr/rnBU1bFJO8TLzjjS9mJyjb3zBC3dKbXpVRSQ+MmZTWMREyhIwL
+c2P0lDP0poumwUqb/HqFqq1VSep63I16HmOMvcXNjIqlmeHwhupOo1tBTievjZo
rayUwb6mgb3DruviBPK5Ox1jx89cRA1UZKxboMlrTZqIOKC5gjVOtst0HE++jQsi
84YJHBVcxVT0I8ze5MnxxvJY1gWQR2hY9lkEf7WEuWceUlMgc7BIoUHDzSGOF7TJ
qGmin7VRJt/710FUPBDYXK2F7coBFwJUjq2TW+qCq71uay4vRPeVz/aSqc+Iun2P
AP/R4xWqMwdyop3NjRh3kbw5MlXDO6LcznpCNF+WAoQJn1rNW3vFNpVUEYXNAvM0
FmWQLgxAHDlNJn8NryKdeDMcKbte38OUy/MerS49rX/UtWsbQS0+O5HZ2TnwXVBB
N/AGM0cpLI6QmjafB/jbM2L1sgkv3ByGlPh6EYWB3CVRzgkTXADurTScJmEOJext
Egy+NRVor5IPei6FKXotl5BpqLkWVZX9Q6uu4WEoWLg/W4c8ZYKsTHwMiQd3cVvN
+kzYQMEMhpTyiyxgy402rEZfDhzlz7aCt+0yMjJ00pgAguVXc8CEfaKvpAY8qb9M
ZIYt6Ag3+a61t7Z+WJ22ICSe72xBtjSX4LKJJOlnRcufNtzfWP46yM50jAMP4hAJ
E591xTCXB0STze/MyZ7oWZTw0OupdduHz0eiB/+EAe8o/iFvYhD2Laozcv6iVrAM
3xvhuLmdKrASqtqGykJDOXR4Rtb3iL/Be5w+u0RBGr/x9Jz6F/qJfm29TNNo3Kd3
BSGyBvccLTqFvW67ackvbJWCilajculb4bdTRO9kQPOE/Bpx7mx2NHtbruzMNZ55
bHwpMybBm4uzaptOj9WtsiKZ1UaQ+ZUrUcLSp0nojBK6METNsX5092GvuZp8YJa1
Rbp+StGnbZxdPpp+ebi0Tk9ao6I4Nc1f88gFMXB/CZSM/ybkAHFlcVwr1awtKSBe
qBO9xF0bfQTC9jMzXO9/iI03MiS/Ry4LDUwedAHF4X0Bk+Hc1QO8ZlB5hJLWj/a6
F0CisLWpOg7lwhLYRv6dQPA4uQ8Pm49kSUuqqSwUsVMST4nmm6noWqlSz0UNjvWi
GPWP9xyTjhyvMAoK3z2Xg2mS8PVyKRHZ+Nsa9MfvO+NklyB9XNfsI8le6fvS/9DH
1OmKtmggJy1LvcCt7rWuNuJhbNwCTAILZhgWZGTKXoy9yb4t0eU0cXmDynbVXTLd
9NtAaFLp/nBFBs0Cu1qY1Mnq3aYfsZgYQX7QLgRCUf8GXbbloEEMwImM6W9cqI8K
uFBX1VLpq3Y8RkdQTvyJaqrwYzAdqIKsTv1JuhIx6f6S2X7+HxWQZ3Vf4q9zUiHK
CwtjR1klgyzEwcf5oulWgvPs8jESLclI56RtHdAebRM3VIrKmC6Gt00JyDivfHat
+4ZGu9xcULjXKNFxHhYVaIsGJqLUhpz1dk6UbRSUgr+cd4MJh/14WbhliQojFVEE
c/Xw71YdepVHZgd8ec9I/3W28F7jfZbD5ooQrHVjQWWyGoB52vPBQ+mcPCHjESVh
xzaIk+SvNr95yjjrjzqjN944NS3kLXuY1RRLrjEoNWfqgKeDhHwxynz5+qAJQqTV
suuL5GDH0+sEswjVZFBYHhculwE2KTw7J5GaSmJqFBHN5OcsSjd6Fr/F1q713Frd
N3VtAzPZCD/TDDpAvih511+lnvxBVElfVttJ/ENPzo47zTni+Gp4HvYsULY5mxuS
1uLpxUg6wpo1jXcnlCYXD7rhF9oNBAjsBO+GwAKBoS8CkeHEGp46Qxe4OJPjEUBZ
0SoswdYn6Zf+IVTNDqOroEGS3IW/EcBAPu4aopQQJQDxMcDhZGCis1iAf0PiTdsp
PoUt343asNmdiGCpwRG2RYlksEFsb2PqPTHOmi/lbEDyNRk61Yj4dDYH4FVnYxMD
jocNd9k1YQL6iUxjf29V0VG3rdAaK4lMkzeqJtZJqPMN/kpsuRPqKGxofLa1RG7Y
8KbSJHUF20pTk5Wt/RDUvjIxNPPqDkvNhtxi+NAQ6fC/UeYxLYz30oHzuiFAJpVy
BrUJiBlnniK+6TGfWxqKzVWzCzMiTpxlLPVojyRVDuX1SxNSE2xFR3UCBSjNFwtQ
WkuwfNnOO39iCy1UQpQoW/UJHVDGS+k1FisMIQPtawW1GgzUiWD1SB0n0qLiSl/R
4t4AGEMODtdZAvwyMfsTZ6AiQzObs+qYMajoyNaeBEcGq9Lic/ev0vK7oLvnGv8Y
FT9HzfvNOqhLsmjkKvY4VgLZkmEbHKciIcpPyatbY9G20E9/dp34GZT3q/5kGY41
X2k2RvA4DahexyDE76WqckyVPhTig9pAKndD9z4ssTQTuwKqVyWsA+LoGKSz8tCd
iKHBxLzG5WlKGukgT/PGUw9CMpxtY/A2b5NY9KtTu57uEy3c4tHPqdQ6RndWgH2P
N5w7P8HYsZKjaqZCj0H5hkU9g3JbIMeuVOu71Bno2F2FdDWjKoy6hfxRKZGXiCZz
ArKMQyJ7gsLppDMgfrvvZHnuFI24mLaTMi1ic3yWOB7qQlamPY9Pv9VzVICHOnn7
Tb44se+YmmNAm6CPNmBXB/vWJPFKyQ3ecQtbsD+PJygGkZFToKu5+Pdyxfy//cHu
b0MJQVC/QJYNAEcI1Q2BEL4nqSnyUfresf8mGPCcNstlKB3FMD9F9ot4IZLNIuMO
bvpEOUvtQ6ICztHaqKUaMhOGeKt2y7qX/iD4Ov4xGZBtHkHAan0AJZTtXwG2n3ox
p4cFFc053aW5RxpJpMMiRdpBez9p21wcczG4eYofxuMgr/2BClGr5wq77kcfWUlu
ExTga0t3o5BBzaxrayGbDV7uWir3mj4uBkp+8CZfnEF7DlbfWxda7BZNquwExsy0
/ggtZmFBUBy7DzWoS9wzPB/KXtLKIN47OFm/El3xMgeTZkm30fIvNTa2mT6MsW9n
4IZH8X+N/M24K6A87cwsnMfvVZtwwrZIVQO7yY2PRAc8XhRIm/lmwTRSHfifP63V
41ziCtiOIOmibaeHSQqIHUFQpa6N7pAxwmol0LWLLNFBCy+bAhwymw9FmsNmyzCP
RiLF4TN5coTKA0kCerAm6G31ozkywS6/Spf/V6qmvv/mxfkGGr0mH1F3/CuwC7vP
Zx6bQniZx7mnEyywMnNhRCVp3zJNsRvFMkjIETSRsRo4NUi8ju7e0LxUuevYDPfp
P7f8I6NAm4EgLw3BdqnB3mjdlXY1nONPMv2sQkt4cX09C5x/55Rx3dQGnp4E/J6w
ucrZLlTnUby1u9EV/Hs9cNI6HFCVra6NabN4EZq/gcTGgsiKYc5pqUvV5QhnfjB2
V1xunCwFNDvKF36ZxnZscVpruyRaM/V+jNNr5GpyMQIT7HEJCB0A90WOfIU2/X0r
DyE1o3GnEs5FknCGqnWNR1WEmFKoGeWujziuZtGGL8xPF4sU9SzuVFNgG7bm1Lsv
+JTCHwyq4MFtU+bZZNOmWecPZftIxKj2KDKD5ydjCiiPod3/InpTfFkM2hMnMbit
FDtYxJwjK7TntcMwEvbi6lodG83B24apUGPyXOxRtQephUuD/hW7dXFsb5DEvCHn
o8eaC271zZvunxQvIDFwUzpKnmJ12qZh+/FhlRByittepDuRNELGDNWMgP9mXIwG
FtKzG7peYwvRDjE+WSMGjO4guq7qz7k5b0jCV3yDuT0T/sMBhSTK2iFJsJTdCkRA
62J37aN3zI3JiGSfCzuqjlpV1cMSeIYfrGX69vr0pE09YzNWROASNf5lz3qgDZvK
ax1TxAPv3FPDDF6YKDl2EEoTtwd4I1zKIRmmT+1QxWbqGliAM6lha33blf7WLgKu
1Pic9G0/WgLX5JFodZrG2jPUK+Q4xIULHMnpQU2+0Jf4X8y2eYVDeAatpQBkAlQE
a34ZJnajGoRZvjRjfCRp1jWjvN1s+THa4ZGuk5tCAG645Un47Mz9YODhvJ0vmueT
APo9kKBXUbna2WFrlmv98gpbTGUahW09lzgRIbqWDOA/dAndTO4O9bEaMDlaBuAr
vIKSBmfDhFscxQ7AHEhmVRX9v7/c2Xq5zzsxuSeUZ6QRW0px5GtRQjjCHSisirYk
ywEhBu4pFYmgmrqjOH8ZOt0NClGJXHf3T5rq4308YgbTN8898uOcPW7cMXnAtvsx
3f8lkXJnLWNGDwEJBqGpPexwm+NS21hjM1OMkK92KUfcsjYCtVhZCdF/Njsv8tsL
+YdcQLmUih7nZLIIeKQIvGFIdE9KSLgka6mo6WxqL00ZryoXwd9x1VOfaTgurLcg
nOr0Qe+Sg+X1TMed6omKeYE8MiqtnO4WZ2rMeJtGN3E1XtNdCCk7Hr+BIIsjtAyf
P3VH/niziKa0rRfyhO1wCDzhHPJIvMUk8ly9MjTTFWAtVEISl7kXruJ4yGtae0lN
jvYlXSMMJ+/oVj1OEq2rwcmlX24u9Iwcv7romKA7GRtxSVpu0sSyAYc9NXrOdec5
rq5Cri98FXZWsiFI/M1Ve2wFNIAKTwSvqgUEOqC762p49ScLV9mIww8CrRvU/sFu
XJxQRMBZ1C3pR0yz84lsd11FQOgsbMjrxEcN3Z2M7E7+vXsSvgfMVff62mDT1+gD
llIi0ShmFqHWGTqiI/W1xC82eK+M74+vPHjAVjn//j3uXP6Q4L6GNHPGcb9iNCoX
hAMCQpijOLXUIdVHR1hUAoaDjq6v5k6nDHvHRcQCcytFcE5IhYLDkteWD510r8oN
D1tnBn/e6HDTUFg7D0sFsy0ZjwntSHCdfzKKhnfsj5Bl2SL6t8cT+SCTL5tS71zg
GBa49l0+Kedwm//YWD/hzLGO55oWpH8+H3ZbEQaIDIV3SvyMffYdyOxck17YxZIl
WIBkuYCY+Dsbdt0mclgjZipDTEhi7Y6lK6emTDT0G36V//uMDy1ylgfZVwDmNH/l
sRwhHmV6g/y9ySpDfXdUn/EA/PF4z+SjSq15wllxz9q3pglily56HTioqdbm8izL
6ExBh3QbD7gZMXIcdImLRsh/psQdzr+3avpodm4ql7Nrv/rsw0cDE/6bNIPOMjwv
1/Nf6YbHr6uvtALHWTMIVbXLpURXcbhDQHPOrNsYv84iMNkmyqsjpNW8XKWNo8pO
7hZ0lbLo3OXiU9t2opHiShR7IV8LpzECJW3k4RMa5rSpaO5UM0T1CqsUbWJm6ThX
E3aiCG5SXQElsgrWBbVogrkdNfHt1pCkOXLocooOcXCwCJ00/Q/G6l+7qgjB0uGM
wivB6NWinxBcfGdee98s3Hur3z74oDqS87qrlRp/+5IPyT/sGAQsQfBIKkZUMyhM
OKJNGCzB8WuWBpc5TGo/DW6dY/VJuBSr9jQ3yELWRxrOqlauoXaYvmlBCzdZBNej
lH83f45p5ukpZq+cNB4gPOmdDCknVydZ+KiAjIosTmTm57NUCdKraPj+SglDfXb+
QBkVv6Li8wZSAuSbNmJ94ZT7OxE7sWGBKxG+pxOpy4qPZ+mkEIoDe9l83nMagtaa
/R3i2lHmJqwBvICCkK1UEk9Hudp86ZfhHvvyCX2J4c/q2WW3oo3sbDxnQyzJTrIT
yDm2/yAu6MQ933BbXb+r2naXNkaa7VKTxieNUUO34sAh6QaeRfzHEGc7UcMLiQlB
0QRuAnTPzKhfJVsSOjWqsxTlFiIdO8ZgqXWkAqQgmEaIWFSeGF//cjM8FHRPQHgW
9cDzR67lmZIk1r/Rs00+ImJbeOxu5aHeEIZllyahVA01/gKgUS9yhMABV7zUDFy2
2Ao0fLfobGEu+qotuTWKIN/lsKNR0jw4Z8nWuDgxcPDuHu/MK1HWkSvCM79Jgzh7
CcIfBnbiUUt0F/zu14W8tng4oQcGc73fnLi5JRu83Cm0rlLNSvbU4/SaKPiFu2K+
6aoXFNRoM+CTfE5Gz/vDfmmSsK5wPVhrO5p0J0fv/0urSc4BtwGJtek69Pd+PCig
ApYFeT98EnNK+EPBAySGGJyTNCCkw9UqWSDYprmJsDHkQlw8uOkJVM0dNnxKmzRu
QDVcdp06FPlKHN2j6gpK+TEzhlew1y3aGZ4r/eJY6E+5AME+8G/h1ypTdDaWkuAY
Wdyy4xSE3QCNdSLbUTu1f/jy0fB1T224J2WTGTkgdiNZ/65jPLg+HJiJs6Ag17J3
GuhJpSuA00StUW8qN8VKpNNxGUUbEB0jvP2zJcvTo5Jf4mNQxUGzNNEQbNXOQ8Lo
YAGD3Foef3stEilbGGdXxsZ9u1xnge//z90TKUO5p3FzidJypFrZ33YuF7yj7I4S
QG+GVtAk39mz2l2klfJSO7Q0lYvR82soAyjy06lDCfla4+cW4qSRb/FdAZaCodWM
g3qoZrSe2ZRfY7ycYEmov3BFFJ7YCvnNcc4oMnFDMxVtCEcZ8LvuZSI4QGIW04Yh
QNgNghKHpD22DETkMKtJdFUGj80ytB9QsbwreQSj4EhLrg7JH5o3j2Qf8ZNvgq5h
kFcJGGeYjkl0GW965dnCHflirTgDuwPUoCaGph6jLLclN4zaYoHLyE6x5cjpm31p
qmGi+IOKA4+2rMekVqY9DrsJfaSwaJ0cNnRvfwf70licKEwtSoUuO0/mBbmpMO/w
iHSR6vxc9AGJ00/R1sh+HgViqPBUjeg06xOZC+FTBa6xZzP1WtojbWsz+HMMM9v8
mLMCnAFGNEiYvCbVjpQrXhAUEJzVxGL3/2wz68rrAkfnbq8v+NqExPpAl9qsXule
b5+OG9vWS1N//K3e4VrV605SV1RRdZn6uQ0Lp0iSWa/gUDmWrtKK634ZoGxYhMcj
W/2A4WEvQ8P5KuYFOefphteYukIOcrDot97Obp33z0YbUh4nqioftf9TYpMiMRr1
oKAvae02Tp9d99Pk+y87yzzah132I4p1Fc0FCnV1YejoL7z4JNfAZey3dPMGj9si
hCOSCpky9q0KdE1mlF/yyxf5d1RZET7VNROUYQB5wBHqSZWeTSoUxMN1mRTggVJe
TcMqQpOvQXa2/UsMKz1dbholXVPYnsH/Dhpb7Hg6fHs8OCIQKqbOGRABqwUkGVPg
AYMDio87rLzI0NnHGybtnBfs1CQAAYwPl4mY8Hshc7e2aB/yEateSWAe/QbgMsih
HLCAGksCjNWlHmdq2/dWFgZaZQMcz3YDFkcj95mJaodWL264SGsbqG3Ry+PPw/Ml
zMi7lS+z/AsG8mF9XgQiHO25gj1anx4wYUCIkgQIlyqgAFgar+yZWCSlGttbRmIi
zSky4Y1sHSbu0qGKQWvGvC0RgWS4OkEBpSefdRazlp/a4Xvx9a6fLNLk1jq19mzT
CcXBvRsMgd5ZOjoQL2+2FJ+JvsT1IRr/ynFleJsYGeM2fDwzVSs217aHT9g0+HIE
SWEui8e7n/kSWNTYC6B+RyHkMvUoGbsjqgniKrXTM420wH9W1I/CsNNTz57vf0ik
hmdrK/rv4NfR4GvwllvkKRqPdF0g8NDaGKAryemzRIbgeIwuPcTneYTHh0vmAazm
ppb/T3Qsxq4UHynYJYTEYPKIrAVEnpVCjG7I+v2DxkdP8CEEKpXzHQV8hPC7WZcJ
JTjDTp/p/fzYV94YaJsJye5345HFUbsYYnrMoVe1vDDA3MElqZCRqFX9jczJK+8/
Z6Jsb7BCQG8x+qo8IzNk6jHVvpFu9rHSjkkvffwLfq1k2kxFlsQtDnuKHLLaV80u
hYxje/YFrjF9UWXvLSVKvzBC7MmjoEUnd08bnuvxDdNehuy9qGxRPFzUnPDU5l4x
8rRAECcgQJ5Y6FS10QTMWyKWkpK8k72VJzTosoIpdV1/60dzDo+/ZNdVrtG3Rlav
XlunL8doV+CcBdxA8Jc13/mAYlrk6SWzxhC7fYBXvEnRPZgvXTvm+9rjM64U1t8L
NVt/YZ+uF9FDIWEkTcUAP3qXRnLdcFjBkWODfatzdkqiZkD7huRW1AYziUQFZMD2
dRoxYRfBlauSO/HCFJe47zzSiSA7c2mUqcHg+sp71JkwLMd7kkcRZOVYuSfJ81v8
aJo/bHu/C6jMr/h9phIbjE9FkB3ypmtAm7S2VGYy4nvNsQIRgpQRTgSw+ElFfw++
bsYBrVv+MMTFxTZiz6ijVbjlNSnaBiwME9e5x/UH0VTjH4sVOlDdcRa3KmCeid6S
/qlJKldWlHG+qX/gyns2JHmLbxDfkpX/xq+JfWaCaxSfM9gQ/3f3tmdyK1+jc9If
9o7xCyfNcGHyDhAWV3/szsBn2KrE1rjxpSgFRi8yWfkEfZU4tTgmw83gNYnhY5lw
OgcWKYBbtwXXWM2mk2xL5eMUBwzjx9X5I7dJ6tUsjk2x7fQ3ThSiTTiv16hpyDjm
4JilmtGG6dg/Bna9pgaVme/7nbZjsQHOK6ngYufn0l9pGb9IgXJmPO5amaSNjOFk
/NCEiQe3HCeoN0UxIRlBZ4gncw2Ki7I157WLdd+Xo0iNzY76F0QJRf9oSC8TpZ55
x5QZVPrL15eNoqqzGP6zoRMpO9Z7HktiQJcp45RfGOQRtC7i++0GCsjw7PLV8v6G
GJg547hPwW7q2OHlao22wbVO9C/NKpZDx4sBA8Fb3M04r0ytXeTOKDXvlR/6HQBl
qYJ47bBUzif3H14Z+5EVnymWq79pRff54V0z/xU0gsfsbdCx/qUE4Hx+1KgRx25l
+ioLX+6Oyi2EQrjmHlqyt8YjpE8s79j6Q5ugCcBt2Lb3DoOtbjh8PRs2m26H0sRb
1heQI6iglc1Icrvx1CHcNf6UqCxUCnk2boiwRuXvLYHnIf3MiZx9JTJSuuVryuKS
cYsJF/2htEXVS8AxOn1i6udkGjLT1jUUovn4xfzjsb104dVpqzK+7SpJi8Rp70aQ
D3fZL13fn9f15tsVpufeqYPRsioRC/uZc3jAh5ab/dqcdkGXAjZLOerWyuyAllnA
R0iKURwWTA6/Jnw2ga6XPS0oJ6xupQSC7mlwXmhIljIcwi9qvfbug3esIHQDv/SD
4eW/Ijze7ceyFvL9WJK4m93j0R4v2kerKVXfeDuUFV7HlhoCzodZyZdxL24ulRBR
zDATy+Fla+eU64lZsCBiwtpDDW093yha90BV3z+e9y8swcL7jU5JaGop/G4o8qR2
Vjt5pHzQ76XL932KmK3JNc0PUur+Q5vG+n4dtGZCipEEFm+pcjsQ81qx3oAkK1/S
riFcwQ/Rva2hRZBno4S39qsc9KiZOeAF+u6LQW+/bNLwqcjcOkeWxNwTGrqWjcaA
7nAJD5lpEI6tEZXhh6U223dMwRPWHOndHa+5UCiduAEAM1Xk2T11UiftqOfpuW/0
hIDaQYtSgDz3UuIhfW3qYZcG3Enf3Ad2T93Ysad7By25cfaCx010UMVSFqMi4Hl3
CoHg1167wOJqOQYL7Hl1VYOF7V8G5pl7cnO5ySVlipfPXqRsjiTyve9wU56qPfWc
fDB6p3FT20egaECcDVBitENJxUTs6VBAN36NnA78Y+9z3DmiD2zFvdUcCMqxPHUk
6Ox2RvXKJw5xKLLqcOkKu0kVD334XKJg7LI7o/1TMwGg2RfEh1y+WQIZ1bqDias+
6zayUqYRG/irHJphdLulCE1IrfzrljrrnEpaFoSW7KOCCkP7vRABqSFzo1xWI4gW
+YlNEk5I7Tl+9eUeL/6nuHeja2razmhOuxP8KSkRKe4YoravCgZ025X0ySdnnei+
pfzkcduTeRuqEfvR9yoeRlOTMZUTJH3+rZ3Y9FosULc1D+ubKqAnnHAqbPhyeJv6
fu533WpnuWxe20Jv9zgbg/tTlgb70sFWfQ6+EW4IaSNaT52KlDm1IK3B2Lq5IYBR
aTyctakQFpiDWS0qMrUvUpeOa9KgBm2StXgFAcJsJTA83MGwoA9ot5mx7hx5/Ygo
WwZZA2ZXn4+ixYrx1pNgGOTmuwTgbiNyyUw/EeQ/1mRhy3ByHuPSMWi/AB1G3MYt
185BVkYR6rF2M+1xaI8Xy2pB9Dqm8ok75qhzIbLGXLyFE5hcpYyjapEJ69Eg1vcH
f4Jt2DqQ6uPFvDQ3VOdIW9Vg6c1C2GWF7+VFqGyEzxWKnpT5oLl7Z8f56S87yFTR
2hut4ko7sMd7WRk6UG8PhHqJ0l8vnnKPja+FsAxFldqD0MCtai2ZRhbtwA66MlJs
Olwd/QEz+8RKXe4sSHZ7RV/gVgMNIaMCmSaKuYtEeSLqriLLdud2tTYzu+S1AXDL
A1N+vZiqHGZGyrrI02anbdAFx5smjvR24Yhqhdc3cadbeK0YZVl6JePWpfzT52C0
c1OFkVTJQaLrhBNyhk4n0oe80ZtGUtuMZ2xY7tOvwmkBLhkal6KZ//AgCd8798Z5
JiqPvryLenW/hlysLNalqIgZNO2GezjtQcRU+KZOiP0nrxlnsro5bCrAOter1R97
SPCrOpiOXkERHOGD+Wg6yMNd4oJiKJM7QhDaD9L3gjgbR3Z5AzW2TnOthay6qqa/
7SPB9RicPhfcBEWZNiCnfYAuW5gum+TjxiWFAHP+Ad8odKxoqYRZENCIIxRZkINX
CCNcH2lHrMv3xFRHgm1KhYC2/I8Fz+nhfr7/7ltpU4RF0jMjm2iKR4ipOJDT7MPg
kiPLtjRGmXnIeNOO81X0sW+zDFZeJYwoAO3hFxvCNGuFTjL2OTvlyCbBVAgjZbuv
DTSJa2i16eS+ez5S2euzWcDoR7a7NRixlb9Leq5YWkSqrEqeIPHHYfCwR35Vwt6k
5ptRei0CYXYTwWRgvtWFasNkJFTIQGmp83imccEmbMFkumb4sLsNpeDWjEMihZ6l
yyYcnBpJmln585YcMw2L7XkzHnS1i0YwF92J65qfOmwqUbTO41RQt/udQP26J1iL
eFNwir+yL9f6mvSUs99FSqZNX7ZZkJrYOgZAMaZ2raqi43Crqj78o9d1l2G/t+XZ
z5VL6vJfCz4XfKcncG79+RW8vId/iMamxYGDXS9uxM9aRJaMF5Zf5oOfwb63YjQL
3ywJZd96rDDGo7cRkPOmV1dsD7dOxfL3fZhE5kehjK5Q9ZZgS6Pu8n8OvSyIwAT6
FB3oNKZ558IA9STk1UXX/xZf7MwlGmK9qVPqEk0JkTP5/7jnfkMe/vzm6dS7/31V
+3nbo5JLxaSa69OGDtRCGrUSMPXxHrpq9Snxg3w1BD5YWHtgMvzu1mVHpxqLrbIu
gaEPWJFmFBfaThN4km8fuO/g5W1zutkN9gaCZ9GYEwlqbtKeSamfLks9NTtnulBi
A0uJCZlJqtNodCi6pfpIHZMgsGHSyHiTbM+N48nYaQIxR95knfXopdcpSWL0Wwa6
y6NkFMQbpdLCrqm3cqRc4ORQI4rO7pF3miuOXTsVO14AJ7ukaweDtduBLn+HJ2sQ
7+OsXqoK6qVt3wvVK60ts/pvWk/u+Ld3Dn2wqnbzneVEqQzCs6TIOoJ2femX7yYR
7bRJXNX26v3ihH5cU11ixmFuL6c5olOd/+on77li9mWX4QTdhNw+sxOUPO+KzV2f
WFh7FBgXK1Dbvc+LeV5G6mq6zYgJ8a3URJz30TSISVcAKKCxRa+zHIKyibO/9D3e
mLfKErhj8G8YbZd3nZW/wQ++cDQPn1ZYXriIJjV5QT9k5YurD3R9iNlBtjl7uXxl
V31DU/713kkKlGfSJ2UVuC5RJBNwLMtF5jHWcDc5y1XwFm49rYjUsAdXVd07EE3y
QXHQzRSv6nqUHaRsiYXxUwTxX34G5tc0FugdD4RUnK7Ddrzq7+u/Ppd4IdbTzdZC
f+xkWD4CWEuSZpibzQOCIHIBPCDLu7lNRbFLOjHjeff9GHyb+UveNmZfaDG+gtmo
Hlot8bzJpb2IojH4J3gtdjeSkyO7vGRrnZRpPtJ/OhA7UXTTkFznA9UGSbGWwpH3
WXlMbowur8pwLyxMEfN6evy41D5rusgq2SwNUrDkpJsK6cL920uS1Ed+r0GdYTRp
ftrcc/GhAd9RL8zkMNXeDHbQzuOaJJk3zZjbuH8pXYt5ifZy/0jUjjXTucSA13zo
+ucnzzX65/y1zxoYnwiunCBPiKwOFlBCVLWTFY8XNyvb6J0cUPj2sxEx60T+j9Iq
2mxkYlzG5kBXNPJFo0TnOE5EB9UHkCnbldf6NOAUH6AMoMv4xT5P63Zco+VDqc/H
q1cDGoClF7iizHZzl3+LXWKIdiz98P+o+ZmxRcLDVvryLspc3X8GVkqL9Jhy7+6U
iSiox6o2+psQ00pjkeG7MibyGstYvVTLcN9m9k+NC+eJwzahEl8xpRzTn9OchTrH
JTCPv/gqntW/hh/bV6fo55PvOZqyv0T4606/HVkV1vWpfs1igY03jsNzfpE+RW+z
90nwlkA1ayT0jjMZPpeFxrxtX6zdcZkAL2Vz3M4pb4Bf8xhFWLaVDi5XGxEqJuTB
GQPjL0VtakoxI/xigm4bZxXL3ALX3NKaG1LIje30EFWjT/qYr5KYmsRVvZ/80twl
5uj038AfcXNWvysTsXrbBLoT7iwYW0FKavxfwuj3R1yo9chexHMAgt4GtGEqQykc
b87GVED+y0QctVLUjOisshlaUesvytAb2Cx/m10VIOPuPLC7Rtx2GAS3h/h2rV+W
QFlnU51+D140eWYH+8eN8+k8On+vHeDtXVpBwaV8AecUkdePr+zjaLwkxu99+PRX
aFbIGyoL9OkL4SRWUp9FaugOVUnmA/eIMuhsQFMJI/LO8HWfrihrJ60rRt4ukcjw
ehzogiFL/Bt+h3wVuk348SfzI1BPKjPQTlb9PM0rf4ySoFPP8pdWQZvd3vFSMPsS
ITPFxJyi2eBxtZnNmOb+CqhiM3juxkJR3mQlYVftJRcgxHXQUFEJYssgaUUoUfhK
cEGq4VV6PjtSrvR7WNVerDaksCpxoUpQZpogPZvkl3uENH/7GZ6pcfapo7GA7Snu
iNlag85zosh1frukEaHN2EktzkQpqMQ4OsJedOWMGUAaCIWztzNYak7gpJ0Hwlc8
AG1GWbDZvRoce2yTKjOKgwe9PYIbMKK96+juNK6OuoOxSAj0FXODQrgksDYODVJe
yqwBtl2q2020IraOJKtB/0TLiuoa9ZWUsa9CvW+WpDdpNBxDhCNO1X5ZxzsYovJZ
nDuadEAUj40nSwtfwdTQL3I7kl3kokTBQ1LBM/+HNoJwlv+L4FKKnyu7+dfnHWMc
SXzqmiEKupR7u1FxqwRJQzUC5ZgVDXD3NV/d3K9mrt/R3/dRGNlGz0sZvify4NPl
0IzyPpmJ2BEwwr+C9VZ3oHFw+oCykfpAYkZkp8C/+AV6mK8Rz0TLVsvEAko/NdpH
zUg7WkkwYvNmG+oQ1OS+5FmmSIoqG8qeiV8I1n5rHp96K5MNFOvwYr2EM4GipaFW
KrTlQELz0PVjZlAcyVhwEGZJtFNUWxwU25/we5vOJLk/VHNJ5zTaLvaZ9I6UrC1j
Uiy5YJeiA7ZJUYzu8k8aokaNDIhAwVHrdbE8TBMsr5vmvPy7feeZaX9Hg91jck9J
AmEQRusssTKrb8gWIZa/xG+9OgkR44aVpdZJ3yULEHpPoMVHF11zXRAUx8HCn/Ln
tsUVtFUhAMdoHeXhy03ZT25Upq/r+krkkHw1ojo/o9z8SkH7R8r0ATMrzzdYM8gw
VR/9VKgiJFFYn513gMo0lkEMV7Bmg037VL8ltaZZLXutIocuaiiehtHKvG04Meii
QGzakbeHCZXT9lp3D+O3I+3JQPCeXu2SngkKSq/uHm4LgkxkF8dBTE9fbWE1cVjN
s7OXDprTDeSZdgrnizX8fyKDYDSkeoRnfgDGIuB1VpRitv7RM9sJFQWEe1BiEW8Q
oM3xK/mt25PO/8Q7v+DiqM4x2yxU/P02Zj6U/0MlDg3vkims/wYwY8RCI5MnmnDj
VxlrIVdqA1Qgx23TYkSEGChfUYFmlTqDkT0BMiQV11D20dmvjczexkfZZyWDPJ/X
FVy2zVmgtNHKaH1B0/GnlAnZ6mZ9Mw41dXpgDZqmfFbjRnCJxkS2Im8fMWm1yfuM
jyXfxxQYBRbMSByIDkdvoTEGOuZuF4uTAuaFO5At29EG9MM88Ie2TxvyfyANfUHd
T5g8mWbpvjSQXqCfs/t5aOK6bIJknFNNpm77pFkqoDbPOEOsVXG3sfmOMc6r1YSA
442PWlKE2H4T75l49RwL29S5nFuP4VsInlfcJI+prf9l1kGm+jTCbrUoCL5rfhe8
xI0ko4ydI2JhSY63XVDTBISc079nsl4ba6NcCcW1Vjsl54TQ8FL7DKSDdn1b8uH0
99tnvzO1Jz1bUehyRujApkPFWZEaB2bKQ6PqHzAZnObOG48oAH//7SQN87FCrONB
bRsuKyaKLRhlMwfVS/97cxo97ReniTMse6+ZQ+QIKVuWJw18JOyHXhsCgNJYbdX0
KvOR7Y3/ujE1j9VHmUHwQcIf1n5s5vIzB+sgh5M0ZIZkFbjP+FA0eOz8anvbEB/p
2sySEM6GgYl2LYX1VRQW+EKKE1WP/sa37IzSMWWvcniSztG482jUl2P028l7UifB
uLHi6QrEjYSCH+Top4L6sNkcZwTCjywr0wBB7IucMgO6atrQQ5hqcnwozsM4YcZ2
b+3gxSRy9ZYb3d6amySATgDZtElwcRLOBKiFHfhueAVEQPGafvvql1qFydYUDgn9
mVFReL8igJt/p0mmXhHWCRHINn5UHGeNSatO1q8e6cOoWmncQszeN1RXZezhe4Lc
wchCXuTH8t/HWgwPKbwBUsYaPk/p9UD9qyVuCa4Uaf6SFZO9SK/au9DmXDcbsYGJ
QN2vDuDYdO+Tly4/yee1rU+aE+6Zb7zH5Cw5F2889uyJUuguiKgsVdxhH+O8pRcs
OyqRDtg717zZ+h4XmuruYOicQDFccleS3PPHeJWFWPE8YPa6jXnrudCSCMQxIQw0
l6qKUCTZMIsdB2IaAvN/x6idsae1TySyNuHKcRNSQ8we+++4uqeYMDrhQD/BGOaR
Fg8YrTq4Ugr/uTpc2W3pvfFLV3gBjW9o6u7VW1t/vZYl+EFcrz14QG/dC3cXTRm3
iQvTNO2b4jPQPFClZX9+AJIvjXszXpSnBmQRuWx0/YPWhuaW29sbzqWdvUpUd3ih
G4Jxa+DHcojaO5XwUlW/YYP2aEv/6NVxhm78EejcpioAZmcFy0t46Oi96VZvpArY
I1/mhWfzlrBOp1792MTHFs1JIfF0CfaxR3CBLtoWfRzKvBy7yc7lPQo70DN3pXJ3
INYgQQf/152sgdvSfF2/fTHxkZfnbjyCZvor/w+gMTn4isPtu9mU++m4/8AvkeG5
HenW4rB8v2kKhvHOnG9bfSi2EfUWOqpWSOTxhZJoI33Ght4dGvJt5PU0zy4mM8Ir
lJr2NXDkS4zGQ9UVSi2J1Kh5p8ykqu/QCpn8w0mCc9jels0LIOxs6UDIeheiHMud
51H/JydXK99ozh7VdwD+QFVFl5GkiX4cKP2TIFgYM/z7Zsd6foEfyhMQNKSIsj0b
lEM4KWV9g4zhcI6Ra89bOpKx/m6SSqSoWRvGVjkBRTIrl5X3E2mq/VTyD52O9Cuy
6JYI0Cg6RwVQteL+/YdbnQSL/dinHjjLM427edORFuKrRhBrzyz4CvXbEsFlsbeT
6vGGpa5kG89uuUcXdbZsjnwmN74GCcXcc/hFpo2dgmGmRwtcXKNya/jRteD5lMNa
AM3Fi87hclYM0tmbT1Kz2IdnK/I36CVgxeYRNS7h4t57ZHllSG5FWstMZgCD8Ttd
H1E6/cQEN/WLXgAEow3LlaBv4rqNu3KjdIjkb13Cov3EaYLz7heIo/Lbqbkxkc3Z
81FLyc8W2YmuWorLeCrb5+UcXuliuTHZN9CuJQO0Gl0ecMlvr5FwXoNDVk3ceBXT
WP3TovbSMe+JEtvxTBqZE0mTDIZ+gICWCuxjpxxh279tpEDU2lmZtiKLizLtW5DD
tH2o444cuUyGsooA/WMojJxw4SNLjOW/TjY4X0EV9CkH9kq//VgZsUZ2DQabWhNz
nXqeHw1HbYIdk5am1VkH+BLSW8W6Axl7q4l5xHAA2deVGnC1Wgll9Zfcm6GKU2UO
Xsnr8/sRdawoitY0mCkkkQGyw66SEdp4hrEmuNXSh4dyI4Wj8GABiyMkQnUh8/XT
QZAFslRHzWudkZwt43t+QolnsSJ/96RY9iSJ19y3TdbYiXzI5mPLwFLs0x/8qLS4
SoNhlWqMNBoaS+yC3WBQ+YUwcnuahzdmQjZfsFWCdJ5uRtQQR9aC1ki2GHGkAIH1
9jwJGe2sqg5FwLBVPyUFZD520aid/0ct4hOGb770akOiN543isuhCso+A0ZZqoTc
LACiPaSngdGi4dExBzsE1W3BjztQu+/QT+YBdpxbGdhnz3VfpRy1Iuq0uw+JTQJK
inCZ+h+eAZjxxrFGiPc+6ftx0u202IThb3NHvgghG/D4nIGv6iyOOk9kqFhrjIxg
LNB9SFrxtpLL1L1GOXfvcB6JYAFgDbv6WoDnZtWXiv6hVEWDC5vbKOD1O70qBYv3
TWFabiErQCbssDOlGZ1OMF+1pn6gt6XZ3kil3ci1z1m3ZBowuCWRoKUZaNaPzOrF
+2/JlPj0gabJgnn20Y33c5um87u8JMxvn0r+9vbhL8ffFj8O6By9ZlU9pchuKnbp
tVj2HWp+RhAT2525vDHiBMj4zjOusO4YaP8TwNckE6Dn7xCJdSJ41cJppppBgRts
5aOk27lgndn4WmpwOtIUbusH786pxRgVE2fiSy8L2WKfiZNFHkqaCqKlfE2QgKL7
rcELLpclvQIUMnB5TS/aCL12c21DV9N8c4ABE8kjac64WOZNH0Ueqpe9zy7vUKAR
034rXlBFqGIHDvbEo581I+Mm5VN8xF1Pw6HwVlsJnLScamoiD6m2NCjQlil786IU
87vOxSyMGjz5yLBVft8WovRgbNBfhj6EgaiF/JSpaCyqjpVd63HzckPyReQ4K/Ce
lZHXQFRoZTn0WgrSpjGFo+UArvE4DfdxEGgDA/f76dUyKR1jq5Id7SV0ccmAF+wl
aapvAKn46uaFxQjDhBExdZQRNLoR+GOVJFWOBeBGwKHKdIS+mHZAsG8Eprk9F6AY
w7RMfe1wUVP4vfNOsxwh5ls9R3BoTZzvkHScAEKCRsjw7Pk03kWmOGHZdGdZsWyQ
XtB29esSJfgFQgZhEJeWukxAxq9DS9XB7pgqEd6gl7oGzpDN6w2UkEFEcS+50FMR
yXyBPtM0LUCOj5riKizPEECMkt/nf5BzGa+F4DTSqxXWQ0knMVnsXaXSDmvPoQb5
KNTRQBdUyJUuI0fk0uz/F48P3XA9rOHOGrLvI4OIHYGfQlI7+DQeo4l4G0rz07Jq
F78f6A26COx39cyrldk5BX7CB9zzcGQihTCh9PKn31vtDJLdFj2dpks9YprEpVj6
js7p7WTNCocftKMyTd3hZxO7htfO86SXlRZjpI7ORJRczC1hEtcvJM7eFng3oGOs
64tcjRYUT9u+gpaEqat5wOBRInMcE1zE1RuXWRlE0LzRU01A7mvq+b3MJWxLyKE7
FIl4VC6/kBudLKqVI3y5xjSkYVoWyeQPHEWjJJrqRxe6Fkfn74iGJ2VN/NDWnf80
Qohoh6RsO0+QIdizoW6LwvMoWXjhrGHTagqJHhC1uXzFCLOos7DYORBr1Ep9hxq5
CASo1fRX6sTRcTPN5SgDwW+f4OewekJ9rh+Tz0Z2j9GB2OA8ueZBMJVpdDqR0sj6
9Zqmt2x7lbkl+FHBma6lvtwIuDF7QV43oKihRPrv6L1zquDwNTHIHfqe5KNOjvUz
9Y1stSYRIxnQH1xDAfd7Ds3cpBJHhlODxOCEnz1tcQuafIOCMFRdiYFqa378wyhX
//mtz/8QsF6Fuuh89K5gGV3aykCkyl0bUXzQTpe9JJq6Z+cnpPrE3ZwwGFWLmjGt
bBw/mFqgc2uzM9YAdk+K5kVEhyjYMv41jGbRrTQOWoiuqypQubKh1QuI2sxzFxWd
tOVxTjgBKQ91wP7pCHdTVY4Ej9wvpf34vWso8kH9Nd28Rcyq8e3Mayc9/VHoIZhH
dSaS7aIeFZeSMphVMEemW+R0zesxFJdDytqQTWzCKHDz7lzCEyoU0ABZtvDrWqok
99/kxPjhwZNOr1nm/Mls7wOUa7+7xVpHoKnaFfVofbRWanDnZxGqu2YXm4+sAh6q
OTxQHXxGtOjMODQepaU1UdUlCbBeUzT627IUxiRnavhtmVRyUZN8sQqj9zN0l5fH
43enJibel7wcZPDhoIPr9nU0aG3LtDxdov3+m8ruDg4AIdggvCBAfxcQUNYdb7Xs
24k1VqpWB09gZsGKUbCeZL0xWta73LP8elaJmKf3UHLO/CNHNlMQKYRkXOKjbbYY
KClzOfP6aH/xc4w7dJdsiLy9n9RcpAwybxxlDT/JUkUiI2ozfqn1CMCuKZtGGX3k
ZqtkxxXKP0y7IvioMyWZz+LlkRy4DYPEOlSiGToPRKlc86xaF+Rye1IpBFZsxS0p
HjKNgJkQDmPwZoTheyrZVYwcp47ZYFpCVk6+OlPDS1BscdHdBKKEwE3eRWSiOD5b
J47RR2CIcjsZed7SP7sr28XVP8p2ooUQREdlVB59V4sPgJEo5Qm9+dKPrao407WO
DOOfye74MkGs9w3qBnEkBWCqhK1IZriWN41TwdBMngDxFT9tVVgM6eFsjv19wAS5
F4/Zp2bjcYQFzHFiFOdAxxsukRK2+29UYZpcsHXk1CTQj8n2cvfprk0UNwl3mD0J
WldLzX0V7L3UltaH/kEL3Z77/+PYHulMDQpTQnE5c4qOkCmzeFMf2PRM4qUzod52
keBbOktotq1uncSCtT+nuGbmnUreKFcPv/CoXSD0eiacb7GqF0qouUDSJwSlJ1Yd
QevvQaocMOgNSBwepJ5URvI73qf213x24vZsXCkYP0UoN2HfXhffjhensWoHQ3+k
gK+i3GsNnISvQ71e/Dve3grruIHh9Os3qlptf+wYbxYOuxY7EE3G1PnbWbQ6ccLn
NEs42BBuaMq7Cm6W1GHXzDAYOiEDi4Tjbkk0lfvKAnrPFmDVcOaLg0PInPYKBIM4
/SDGpF/HEwlZ12b8MGchpER5EmRMBDLWs3dhgLeEACELYvD/TFAw+Ato/TXgQByk
bkYpWttaQbNzh99UyaTouAR4VNMkaT24hEfAtE1MzH7VOSs6itk5Jirl/NilM7tI
riqaS8VBPZwxx0ZqNb6KRGUb/erWCNYTko/ok7dodfJIFzWYndYGKhdCyU540LUZ
6EMwBEWgaaGLqNpwoHNBNgdhDYd0qGVmvdna1qD3v7uvu5xaW41s/lTFlhrX2j2J
AMoZfOqJnLmN29Cl/gzle3nYeF2fvr1RmxcUiJ3uq1jlSVkC3pBjGYJ7hnh9M7oo
yQ5l02/eCG4MSsiINs/e86f1nYC9mutQG0GBeyEdmz47iubK/eVaIr5W/HkTRvhS
+9nBs5plbP/36Gy2V2GkYEmSQlmYyT6KXNU9FtBQeCP3CeaulQTNkeofSsZtGLXs
ZmPjTZrqOmwZqrcv8RhNjBvYJJxziSBoc6xiuDBrLllTmetpft8JvdC+QGEQrE2M
Ucx3yHfZil+jaBjGP9ZK4VwSAGt6UDfQcQb9et1BwMbzzZAn6n1sCZ0hTkDBZAaV
ZtHSYCgiSwYGK+lqRUAjG5g/zWwR5Cbc7CzFAcAdnc0xeudisom4/yggzULXXGAc
IWzYWqxyRAEqjPnB4DEEYD29KAnbwh+dZZ1rsaSpLCpGsgr5Kr4J2xaSPtPJKjBk
3cKhXS8hmU5T0krtOW7XAs20xGTRnHW9I3WtDbQwHDf2XS0JqOAt2pWPyZ1mfRKH
4L0uPHw0Rw2RaD266ULT87tgxt1uv5X1VMXQWZ3owhq8Pt/pEJKxq1I/lNQN+7ze
FqqkrG44B7EpxndtzVQcr186CbwLxm4rExvnwX9FUAA3G//f63ZwW7rUnmjiXltr
U4/TfJ6AU/Mp1AxmM8RZHu77LTJYfKslcEfM69jMnHWObnQXs44N/QVCSQ2dIFsY
SY3DFP4TNgRudhJ2sCQq+qX/bJCOLiulpt9mFuCE/9JTLcGHORsPPi0Gm/m2yA57
VKvtMM/SE8g7GbOlfI0QxVWk26tWXKQDJvzm85FT94Dmzc9HNr6lHxBtKMRQiS5V
fjP2xk1Q44EkevYqj4kaMLLLUsNY+Csq+GFUn15rBoZZ3QaUa0aFt1IFz7/mRJOV
PCeD/2OjjJGkPXza5VN0fTwTfBfjCFk93Y7e3U/ZjKF4hFokNYcN54z/C5FQqOB9
otOAF4ODQRrryre0DlAquE0mTw9VafJFrUioMoWFD5XiFPqgC03KgPotfzqOgrSb
KGlfYm4zwEkMtuZ8aVm8WHdvEZ57OeKyG8B7rEig9Xvx7m6wOn2Pfz4+4rgcH091
HuDJI9KwlefIykchJIwodOdQ/fvHyiLoP7vO6xbVcurTXqhOtwRXPaqrKdQBxN0x
8ZzUz3qm632PGbNqMG+786rmNfsQCoNyE+a5Vel0PS3UYwdp8JdaxubPPc7V78JR
wlFAmFqFWgJqPigontOmYF7wF52zg6WyB9NpxaireSj5bb6VDMG569U77TP0h1hU
Qgi1eolHLhU3kD7r+jVIyqoYucRH06zhfUIansjJALTxa4U29CPI8Lv4ckj1IsLy
DVT8uxqqycm27a4XCgmAmAVEJpbwsG/N8d6Xgkgofvt7FaqsTu1hrpmVSFsycWu6
uTq+n7WGtqNy6T4xYCyEj8VQwEmLD69hXrt7G8SCafRBZL3+jRYdvTNe3+i/6EfY
9uD3IfjNhSnIjYu/pd6w3AU+Xt+TfESDpjuahuwcLD5/CGU+Tul4tnR7JWcleu3h
IhjM1SyOl+I2QIPjTGfm5lVSeZjhFLHqSq1P5f31zOKNpia4ctEbbZ5DuSdVMtKV
EkIStTXnNnyFxRFwYpkTAYGlJc2ZjmhDL1NifFI0y9IADY6MKPmEIh7rR4LLow+v
9km+yCiOoGNf8yODSV/KV6O7WHrrC35Rhjh/p7aHyuqaL5+rJ9pOD1tNqIrN3us+
5fLMnFAs86AL88NO23EoBWUMrpEx9wwEBvCcFuvqKkRDz15dPMcCfVrZItrY4/NH
OJ5xXA+IuzL2fZSbUepMcDCnLTpsG9noNoH4ZMvuXLBLMlNroOylxebMWu9T/+kh
jQH56jYoBD+lQz6PmQY/DYc0d2D2QgdiKD3VR19bLRHEbb+lGo3GnrGaf8CFcZPv
2wGVFNbClBjULvuGvOGhfEJZAOKZWRBriBMs4tS66JdOoYDT1N0VGIUneAki0icF
UHRfjvslwpdo+jQqlfCNQW2erdFtIf5YEXWWgE7pgsEMz7KBRLUXuDZs7mUj4hUp
yoLmK5v3dDacC5V+t3gQFE1CMT7NT25IWpywU8/awGrxpnFdPJGwND6AvDIt8Vq2
O9n8u03dDjc4nnSCCRriu15GMG4DzYfbK3Qr5Zla+Mx85cFWhDUOVgn1DiIm7nv9
sw632lUMYJbcWnddCVdJ2Ppo7S/cSH8X7QzmHCOS72TA+t6J6cOl9rPG2QKS5TWB
BkENK9SyAqqFV0Y/3VfiWEBtaxlP8uGwE84RojyfWftDuaf3W8S6MKFFKM1INPqA
x0+UE8L6PsIsy2FPs+nXXQW4cjA3uZ0lKB+kMBRVFYcmynwbqVIcJF1URlacct7g
MGMr2KePLchcy2tWW2n+jBbJJYenN7QuCFHMIoNHLXa9OC6UReGLttX3BcGQvzTR
E4mHC7oY3sMYlUN1qtSiFFXZApPvqVNhMf4zb0ojS/QPCXsKr9NwDfOo9/73aUT5
3tsDptnjtOaqZnR9IDNNFug2R4rS3gcCPSM/YiEBiPnQlMoNPfp1wJggM/3tFfBG
q2awxsro5CmVfDr+r2wfhauaR6DUEdbbmkueTIQJ14bohuiaZQe9htUyeaq7JyLN
GbzBZ0OlZksEH3hhPwTnhmLkmvAaZdxXto7Jz+Qh0rjw17rcwpgwL/bLbsNzoTZs
QzK6jnKX/bkC1H55aTJnvSJtEquDBFgU5YYg6OaCScEU8W7dFfjjwf/Hz7Tvdnly
6ZxPBkGIT3uEYnTVZkzkl8dE0jkaWCVleQjbt4ywRTEusrHdq4j2ilTXwHVQj/FD
VO01pjHL30RIiYftUyBTCulnYfQ+9GK2Str/c1NhiAR8fa+qrPqqlG9+JpL3qEJr
8Bo7EqFf8T6LnMjnXFKM4mJZcP9XyGoGsUOTwwvE5DDWq/1hxfd2csQGzLLCUxzh
wG48lIcCvnt1LK2Oisi04Ju3jyImJ7CkysKGPA9dVyFK8Su/syvQwGG3PpqxrTQJ
/zn7YjrXvm8P0csw+Ff48XhM3AOVErEg1qDWKKc//S9vaiCXIwhS2dQ3dC0ASAzz
7VYt9BMSKY9AkvnTox3/zRnu2I7iz3miZIev67U/HAGw1weD6zUgTYa5Dw88IWp+
y105pQq0CL/CKIn7Wtmx31ff4Bnvc2G3e5dKw02OLSqCmyKYpdDxrGU/vsTWcBUc
8QAODjk+366ALp22zZ/93sq0uqqeOo3lvppo/fUCyJGRy7fxaxhwHmOC5sS+HPA0
GtyJQh2PHU1pAFOhgnQ4TvZI95CLQki3nut/EZFNOLp4alAf2EjVF/fWAs9y9kIt
2hrrY06WqZEA+tQdJpohwCpQhGSauDrDBSe0j7UMJMuXHgvkYLX//eRS3bsSbGYI
bgh6K1aDG8zSf5kRqWmWav0OEdzesHyUGo8Bxn4o0+1cOioZ7GWTFHLKi7AM3QUX
RnoDtjz6Rdkh9DzNPFeJXN5y4Q5GfYnJpGyl95ijDOy5DZVp6K1rABwpuBggu9ZA
idm42kvqxO7p1fjnsnmo46jN5Fl7mU8o9fpy4KNKEsIAXFBhep4lBQX8GxU3sDNt
wh8Dv/fIOZZk+7U/sEXnmWAYf/g8m8v/KQ6qIxM6X4VZN/KNa6dy6g+mxaqoFrUb
5XfkdTwfNVoq/0wAkp9qg22QJp2ATa4HXBw76PCum59Y+MwBGjmg+yuG1r4HqENL
AG7KckGdeYbha0onXIxYS1nDzP4i0j0lrtuaBgoH/S/neXy7JlRWHC6wyZwGuelx
cqlwgtNPI+kRl+xvQGztaKAHn1FBSYj7JDFEWGWp+ZPSlnQspFncOg2P80GpxwfA
givfbuIErxBlxcjk7uaxBy94+Dkk/Zy3wn0oDxf+PWQQEHxLc3P8zUArfFblGErw
sQ8dTtUTF7+UhyWItbei1Y8mgLBAhK8NxDyoqhfjE15/lIuLpKABW0iWr9hl2q81
daA2R8jrZv3dWqdV2S8LTkdx8075XV0oEnAFf7qtCvbbCkf/ypbe787D75YnNC8K
0vExU9EuicewcQ5fuHWiQ7xlOdosOVjV6ogvz6XqWTLEND/Yn/eaRqnFLexSqI0k
go6NB45S2+4tz/wRvfD+baA/2pN+XWHRvaJeNdD7gw4Kg7mSxM0hvr7cxGwQvWGj
EFG1NbuLVMFVgRop6kihnFwD5ybI7fmsRcwQYpY5G3EHREvVClNfCcT3j2WimxHr
dtqNbTbqEk0vgXFL+PXn/k1RALS8Y6rpzRQcTs9hMJvRHUWmkjOT5tIDNln+wHSO
oGnjlsV7jPYhx5vftJMifv2UHiL5pkZAtOg34Q6F4Qn1G+l/O/g4N14Rc5VrvvCR
4ef3mev9tjk14MmeRtU4BGjJRConczXHnxjSnA8elc78sXy5G4faOE8noE2PTecG
pJwdAB+MhhAY5t/hDYRGGfhvdx82VOxX2V6Hx7Fs9OyKzsAzOUNMCeq69xcmsYVd
72NXTJu6G2a9EonG0VX2++9M55OdJPj7EI9pmNzivCikCWyUykbuEdDhwA5p7I9U
rEqRmaZ9cA94UZqxPXY0dnPRXyzXorI6tFJVpKFXrbfI9foC84ErkEK61aC5rjwG
bthVY36LmcRXYI2nsWVhehvOfck1Dcj9jhtX8PFl1S9c663g3xsjS1rVf2+ScI1U
ylJg+/PWwVTzExTTRxjNgw6muUZdyMMXSgKgGfaREECjzdfzfzmT26gC4zLzfcGn
lDT00JCUfld1LCJa1hP0roTMFb0ptPtqLqHaamK2SDsK0hpHHTFrui2Tg7aOMoix
vrG4F8BbMxIm9y24gUMFVR/QPG14oMne7f5FHKJn15wG6q4MsedpKOL444vpICvI
3QBJieHX/0bD2+fm+KCRDl9XiyBund/GoJwiSCN6hki70+ZNGjXZv6XSXabOhayW
rOjhhcKNeZdARITZ76Ljqy4h9Aj0DpWxqduY9bHg6+DG0YUTFcPNZhRMazYFft1s
TWFdxUhOS5w3N7knMOfsA5pr/dYKP4oIVj2VEuf7ehhxeB0zAfodpihkefu8Yylj
JS3ZdapYSbRhHtxb6vQgAzVDwKMg+pCKvNGLyqGdP3ExHacvpcZp0VrfPriUcKB/
eM7MBq0Uu46AE9uszmDCjVhmUvxmGv8XNZuo52az+zoZiTCMTD0olUOycc9qU/a7
I60bjWa2iwrc+/4Aje36tZmOEz3ZPpkWBxLx4IMN6Afz9vpRCkx/TnKOCMSM15o5
r/dD1Y/nlh9UQ3IQ+qehlZpdOgCEsNpA/+t7lme81K031VsHYvfo2FqxNFhq3+7n
FwHKoPIgtuGI1vklJWzrLeAPd5bGZRHE+bLziKaDA4tpuyNYkahq66kF5XYQxFk3
bRPFYqUtJrBRJt0qbLUOC55u4rOOUvv/2gxzfGJYF+0L+GANuFl1Q/CiuGtTnDBk
h84vd6x4UF6tnylAVj+AFTBso6zi9Wq4ZE3iynOBoNTateuQ7AEv7kO3GXsF6jk3
8apceiASZyEuh0k2JaceE20aG5eTky7JwpYKV4hit04SnHr8Mxy2CgTfuGAedi3z
kCR2Tsyz0qxn1zxTikmWAotvZD7RE84RDcFV02t7r6U1w7WAgzExEmVrzsJH6o21
dpnFw3re7pPz/g+JkHN3gXS3fWKZBL9kJjJwvAKSVt/pkBkYVjl+UqqPnvny49x6
zQpsVTo5Vja+Etu0OjR49Hog9EqM9mzxnHYrQ3PEzoQUh6nRUfC7odZiLfB6enEd
yMMO/VXTSj6oLKh/u1BgrkPt4TuOUqoz3kktuaXWWFV+TujrO/lPXmQzmN4FQdYT
iDmCJoif8HzbAymUSGZUS6klAZr7ZR2n2lbDAUEQMlIsDKdnOwbUEUWKReOWlG5H
wCouV79oFk2SdGwCbOmeOC0WiUIPWJ+rCH4BipLvkcW9+Vx8ummQ4eWlfMRqfCW8
C8i8AGY3zpVT686cbybm/1dn1oG5wTB2hzbjh+9RYdRi6YfziKAkTCbirbBql8nA
TvjiyH5k9pAKkjVFDsNOgSYuMBl/PO1Ymnw8nUzZg84EFEdpJOnDq+7pdYLKIvk7
18HBdOxbRS1qeZCgGoJ0fpCw1herBHU3PEPLmEPm/tJUrxKBT/4L10qPzbnmeeYn
lxN5hY+fS/SeCpdp3zPVohfuUK3PzMl8AzKfWQxuuLEM07WJHtW43Zz2fiwUxTnW
V9xvy0MJTvUEGERsKLkS8d55YZ/ZsITua0sBQ3q+YF3uVu6vJxdZWKo305TetIlM
MvLlmLwtuZwkHm0CNzmjTu/C9kV+tqLK+VoolipQQeu/GwGLaIuGgiWH8naBLJmr
eP5Av/4BhaBdaXizVy1cLhr4TuZLnwPlYZ5cn8k/LaWYBMGG+Cw+B/hPykov13DH
UKLwJz8W0FUIn53kilLIGOAUComREillOH5Ug/aXWgwTR0UrSBlP5J3vacGYFuCz
F9V4LIRpmcSg4nZ97G+MyLBkCxyOihKsQZYarvPCBj4t8HthbpuifBp8mXZ73ZPm
2NOVlLvf/1HOaBlffIjWO2/WF3XiiKVs6Rv1VVmY4JEppb3vTr32uTHAlSOPGqpu
I41+FMiZm7DvUpYB4rnb4TGgP3QwM16a+4QdKO+JCNS9Tpb5S6uLvqQznl1lMVay
emjeWzLs/DYYwEpC5YpaSwvU8ufw3Ikx3mtvD/TDAJrnG4lXca+DMPg1HPM0eV9X
HKE7lYINFdqHl0crhOLk2WyVtw0h0+TUwDYijCvL2/BNN4dG0Zg1isnhQ5IJZ365
H8yM83g4Ua3ynEIRSWJa0jc1CIwnG2/bwqayOXiIAo5cPLRzs2A0m5RSz4t8oCEU
Dh9D4SGA8ccl/DHWBBRM9KdhDUk+27yp9t5djC7PrhMF5yIgdTRz+m4BcvK8RKn0
Rp9Ga0aSiz9rb5w8X+gHX4KwD4IjckU7YoERPEvWg3pPqN60ZSdKBF8kFC0wXOOR
dupQJQQVJ3PARkDCMbARAFWJvlHMQDOrWiVlGHOtN9+pPo0KQDUi98y240Z7fs/1
f7ubfVKJrz9hcjMyn20FMVteiF1uzSSRK9KAtZWzEYt6e53Cq+1scrHqhjEg72Hn
7ayk/4bu2XfstjUGQR4fb0vbdKYRqXCwRvoXrZUbdZpIRbagNbtItui1MiOzHqJf
0/sBVrbJzEGc3QI0W4aCQWDYRZYDQC8AEzt9hZzHsNoJ3TfrS0TzJhHKhBYQVEoo
6aa5+3CE3Cs2dgd5ozbhdpKPrJE9K4p0f1GUngdNrLGQquVrbTF9VO3klmIkoaMJ
y5Y+CjLOLemsq6AOt+C7WU2QWDTqNVCjkJFB4kBXs55zSQDdj6r5i2mjxQOH/6lw
dTZ2IIlJ9grilaBD8rPu4t4/q5FSnsBNA14ZH/f0B6TCn6+iHXJqOzHYu5gR6fqz
MOTk9AgOZ5uOnD7VcDlR3O6GI+Z3O4OvwUlEl5kIeibICExTDqkvBRu6DyuUyF5e
phVib1ma3wA4Imkbq07g5RYyC/82WCuJhpDtNj/LKs4Fdno5yoiaHKZVsg2yb0SY
fqIZJOQzfP5qZJHJQpTiZ5mMbLZ5xjOBoaOxNbW7Jtk6IJDMbUm3KHwtmvESwnB2
Vu8YWjjAbFuS8o8K/WbczMmfVYL9a+JQL/yM0qyic7JlTHpbRI/IibGpAN9ZR8dN
eVTVZFFAvyhcDI+04YE+OOqsI97moiAO5OGeqlcdpTMkHEe8vMsgQmpVOO0smj2c
+wodidQZxVp02HJSUvHhbce8wtiVpHsXXC/sfLZTtfyXBlN+M4HyLOliyo1ymXIw
dKBjusMCb4UiDVw8pkmGOrdTGa4GAuNF/cXXdyK6gWF10X7Si1M5TUxpoG24vjqF
xz/P8Kf6g6xu0g8gJH8k5QMsrWo8xVvx32e0OSQjTZCASkPI5AQVCe5lM15cQXrh
lxvKH3uEKeDcrKu67OtgW6tHP+q0/UEpkve2BdFJok7yiwhgCKgLdceX7G3HAlgr
z7nSsqyZebVib56fR4jv9YTD8OYvhmr1fsyhyic0b9dYN/bw9f9cVFj5bf3Q8W7K
oJGDshVcHLbTGyuUzPoidSYF5wAv8kfuu2e9jAhpGe2XYB2LwnvKFKZPykd/ik3w
IM5F1oZZBDgMnLIDZB4/4QbD5sabfXL5AL/em0pVW/6i7bIDNpYxt77ilREpGn7P
RA/Lz9C3yBpufjfCuOGTct4SXPN51BtRDkTCYDbcj31RROwjetATWkCj3t7WIsOo
SkrllieNyzDJrEXrlM2qZlaiyfR2DTlcB/asTkp594EVcinQmXudog+8SM9njY3H
8RCLf8DUcezBCGGVEdqYdKGakhNZgPxSXABtyyOTlArh1HvF+S9SWSFd4PZKa7tS
vhPT7WeWYLOCt7b6jFy3GGp92nbcKks5RLkD1XbgxuRBQSb1K47Xs/S9U4OPzxC3
XwPIwHYoPa0sxtxfR5UQJ3gJ5gz1RnoA/PCwOnVL4qQveQY7Xu6FkQ10tXlf/4HM
3mqJe3S340SpV1csEfRhG4KUpFT5oABEJHtj4Em4BnFsv0mzRH5TIALcBPsld3Pf
2PJfD5BPHjPiwuApQsJwjGCRD1v7wF90mwacnv9t1KVu21bI4gGuufJSErB0koPm
Gt1GStHP7mhKINEFuVqP0fRyuGap4sSKoa3w0lYFVJY9Ro/cn9OBex7K/Q1rfN+A
69RGiHLgdXg1/0ib3xe74M5dR9JIwKjYIuHENwJw9JdQk3Gqr5pA634gdwb+D65I
/8DG5M3sSPjb+aby1jQjgZExI7ELiJu4iHzW3WoG8LxpHYc80uuGIZByHPREZwoE
nno8BjHgLDnJya24RGete2SmyUYw3+CpFMEVTl58mPnh+u9/xtY/tAmVCOd6jcqz
ZFUXGXg82MupHVEYDP8rrMQBfl/n2bN+GyPDtAvL2eACYi4acNqei/rD/XZHiP3/
jd9I7Lkb2X9MT1y+ZJ5VVV3rq+nfHIa8Pj611HR2pTWheVt4THWTY7ccyF+mzJVU
bAb+YIOkUI0EYbTMgaEOUIFULueK4n+tXijfRMujxULU8V09kZx3+EiFFACIiEO0
FFUXxHPE39Vv6PHzgwJ2kG1mAoEmyrxCur02T5EJkKidGibRBMj++RA6cnvG8D+g
nsuwghv058S4yiRPdZfkC1j+5/9ZaA9LhavvtYYGN7eIL4jTqQ37nzwR3ulyMJQw
D8L2ruqrvJ6siYsAQb+XBGW4eVRx0ZP7MY0cKAodI+iaVkW+HPWw5flSBtQ/IXWA
HYodzSN8VkosAxaIX/lVwuRrEt2A7i7UVfa0wFrWeqCYciC6M72ZworNwOxdoLUI
ok70HsfdKOEPg22vnINo52aHJvogcVyjRt4XtdepklP24Rm67lp0/N6SmVbVHr8E
raLypYG097Wrnc5/a8tTkOtX/qzW09Zm6IPGq9DUSFMl857cCSWx2Gb6XhipvhS8
ESW9y/o6cITAL2ld/KVnX11OLcdrmuFDqY/TySRDPpySPmcVkbz6SPhPBY+9alZ2
OoTjt1chg3YL691Im7qByJ9Cpz0oPQCaBdEB5SOLw9dB0HiYr+ID62nwk9IGGKRI
u8LkAMUWXM9Fic4SKJtJXl0ZX59bODY6dhMgtUjI7jvlsdEQ8sqyzDdzmv9UAYR/
7cV+u0GthXm0OP0PBY0zpvxcuo6sHarx83ODkp/sDJjKr17lCtoDrxe9Po1dHztB
eTQ4CioYUwIglQ3hxSBHHYfNX0ZnHsPRSYf/jGHxqjKHNC7m/S+BDf4utZOBrzAj
TnqXc4pN3ZZ/C9f9hsOuFWb//08g00eR/1jliY8CzVcEMSgCz6kh5uhhE6KHT9Lm
s2OW6okW2llY3DzsWJaCswO5Bd3kvA3w6oUZ2kDdjH8mkd2ABxuCaafoYvmHcM45
mBIIJeyOJm596KwCd3cYClwfxcyanaAP9f0nMWonJLQm4jH5DEDklVCGNWaS8Ee+
yT3ZJBAjx/qipRlYCjHLENdMnmu39wcyE/xMAhWUAn5dZWVSKwyNQLOhAfcAKty9
vLPxSn3eMHe2/sTx24CuwhR0vuaVs5xCLunZZVhmTOFC2gCEjMb7mVh/vPYEJbt+
XwfnHWgOGw7GFKiDOtqNfm40hSfGyHcuF0SBpN3+mobyziF4osik5PlpkjvrmeJR
FKWxrAHOLTks8+Ph0PMYV/CkaPGmfxrgACpENltImnU+6+d8FskV1baoHEv6RoJI
D5yvI1TLyroh+yVibx2EhjpQdJIMua8EjhyLAiWCqEaozd1aUR847g4Cn1SOMCFv
/2qGAy3RNwayXzo9BGdoiOCcP8goSsWyBflVsyDqPvUPfVMZhg7709Az7D9XSb7z
S+I9ZcjaNnicN3po8t6rQbI9Dg8K9EKXDIEodX+MxJU1u+07nHHG6s9eLXCsYBkm
dkDnVDFhVAHJz9ZeRsELb5J/3A+fKGDF/xB+l0HCYx9Qrb3FcM2XTBSnFpfwR4qn
NheBF8bOJlL2230wfahUa7zxG4WwnfCTgpaetadoBmQb4SMWD8oshJNKDLmj1zQd
Ltk5jMrUSaBGhd83ar4NEJLBdk3CYN+Kr8XCFohY0+Oa2EZ4Sx/UlGRAXbbGtKUD
GGFEhgeQt6Xr0UUq4wIALWwbd/E6wW5vgoqq7XvFiNyc8l7FsIJ0rGxtPUvpIi8a
VWUjuRIDsbU9RtrJf/muPX5oH6E5xYaOTsSl5S3KwFB39IR/4Cw6U8AU3bMCQQiU
teuTaAdbsASgm9G9EySAZ1cnpwMzwuoauId4N9YGltt5hWGnbxxBUHRGAkEOhiB2
Mjwy7MoAEz1ICrLufgh09JmvagFGvqYnOnCafhcE4gUsIGtxG300plzR9LyeMQ+Y
shY86DeIXyUonHXZlT5Q7cmmFSbZi4lTJzZJMwhQmErRZYriP0wjtYe23iI8a4Fd
9QQGe2YyiG6rBPxFR3sBoWHSZThnVjbOQrYiKJw+CEZY1bWcy3gVtviuH9jyIaL8
041UFtJCixEAPIP93RaK/3XP4tuCs4t8HVtcaeTsXF93KL3tG3jlB92Kz9FwSIvT
iyQKf/iD/xuG8u2mKCUnPb8F6lxK7sGkKkRJCCv0TDr3mQfPqe/mnfpkXd7TMJGk
rDGf+WlzFP+jtPK665qfOUco1OguKVNT20+CZzgvZSbFcScd5snsKnVM/NcrPzdg
2jlIIX73DHelC12HUJcGnGUfPVJjFHz2UzIqEO580IS+30OsQPllkfLyxWQT1wh2
f//lQnxw4gTiTRRtO7CivPOYK9gjnQnc0ofLvCqH7tF+ZdmpmwrpGG19xQH5XiqK
AdLaFwmZ+IcH1W2pQAx8PqHLDQy8GzjKHS+8urgaALjSXQDPhBiGdUjhFRfW1LiU
DEpXjS/w3ewLG/TZo117MhcMq82RK73yYctPIn9pAkzjfyPmNeXs48Q5WAb1cEfZ
QEzoWWnk9gyV1l7w+Jb3smpLHbecEBRB+s1iFO72VvSy2Vrr7/MbgWooEcaeIiUo
l1j3mtrRJYppNNvf4R8k/0e6WwS2hVTlbNFP2P0qwUbSlrnONYd9KqAnjmomyKaa
tGluoY6roAi3X3kUWNjh8r64J/hpoBI38wzwKEBK/9u36FImrR4PEPNrIvZX3eWt
jxC5hQCK0hUN03GHR03f2gGi9kQADMKpkcMNc6VNzTp1JiCJh/ukZm49g+uOGnh4
DZBzYDYl9doLUi5LIdBES7JFfCpV3La86/vMvPWaIXECO3JYPjI/e7QwaYWC83RF
+DtOQvY5n5Uk8+7UInYnX6H4XUZ0GCCk4HgRFxgOUcEjdpHd9Suf6Lde8MvAiG/n
bISeQPCV9+o+I97dq4zuDhoQXEvXW+6HyjPeO285zEphCrDmcL63zohjsYIkiDje
pAA5SUO6Srd59HmluA1DFq4ohMklo6MotcMED3av0V2S1pYlHwjSL6qwG+y0F6cv
yIFD+eMMpIDezXhpY33RWBUGGD3yOXt5QJt8j+BfAESky+d4qIuQ/RNZoFOoWrjk
Sw0151Q3vqRfeQp2rBcJTB+uzkhuYL/2THDSbYEaGwMKk981vk7ruqPhSU+Qpsti
zUYx8xXcybtPVx9LcQUaBH8a8ttdMc9DOlbyUdwbgLdUqnGNfMGcfDLFLJ14m0CT
ORxlrYE4e760Ztc0uaw0mDq9wOc9thMFZBqKBMrpb6A0yMoQWcgMPq2drh7TXr9W
3rEpZfjbtLRm6AwQRf89+Df7L/KU0QKqYlJ+vvEj3asa/g3qrrKZBiHHRgnaNdOB
kb02tK8+V83tpCACktrnR5RkDaHkxk4/khWd0rIWZCXrXejvB7Wn9Uf1HRJmVjIt
AiywqfRwpVSTTXGoWQVTAdOu8GcQm59oXnAxFWs/8m2UiwG21+SVFJiEdZG2Z7eW
m7IBlKQjK35IcvQEZ2nWOYiuPcseHVaVTGG3SPPzvESreEyyDgRhppoYkQXrgiQq
lvyadgovrZOU3wKJtXEBq8RWSASeRy13UQHkJtG/zm28v0q5M5p71AWtRsLwABIf
VKklUk+qxjP6pshuOYbt1YVt19qdf0yhvEZ9Zq1TvLJLRAOYg1fv0q50eA7L4hUB
Et/83K6TcVfbA/EcU3/B7wFIG8Y0+CvBpXdI2VXeexXnuVQZHelT9MhU8KLCZu17
BOUXkTKwu7kp6S4vN+rO+b8brmthar0stkVywdaO5f7clZE9C0BQfoWKY+b51Kfx
in+8V/O+QEiLo0UFGkDHqMna6sV34qQfSkb8WWx4del/9ZpYwnACx+3sRuRvMcz6
ZF/CzvX9McoIjfVgAgBAXs1SdnZ/BI8cf9Tzv/RDOprzPCMD/pZuJValdZ41Kcbf
ta3ffBigAacNip3GdfQvfearq8RVdvAaKVTOq3BLc2/ZuVHZ5b4v0OHRdxgRYs3V
jzdLSRXrYbkkmiutJwek4P6yLIkeVP7dOjGK5e1LJs1lLNl7T7GU7wWmBvT4tPyG
7WI3Po+qwdJnpUVUWTMSZz0ZLeuHOyyhl2LEQZTGiTQYoYub6LK83fMksPJU1Eoe
8DCnS4Yxbhy+7fD9KUO41sxGwdNqT4shwBQlcnbwLfRQuijqqUx+3dLfKZHY6Yty
XNr455Aqe9jEuAtOSihdQP7FydaP/8X1gje+JRExzXYbklxsTRD1fyLzibqVYXSo
QOysdwBl9sFudQMuSli6YSbsxIp3xm2crtyIScVkBmaD0icoYS5liLY7dbJI8czL
SwIuCuF8q3g5KaWeXO8WXj4baaMR0nbYucGamtMUPcU9uHLm8hIykemhJASDz9Ju
dI4j2fw14FJYcfkbZuBP6qu1/+6eqaXKXwjj3zGPgSDizy1StUDWU+qU4oCo/4YX
2FvNZ9Qd10waOyBCF0r4AVZ11vKYs0PMAt9Isr2tKbJgoJkCNjXTej7tK+5Y0fq6
jts6z6edBaSK5DXesthjJiHQ9o2qLMbduZ7w89LU8zIaOHIV56OoW0zzoRyAyNOA
sRWhQYkcYtDM/39wHyH+6jH0P5XZomtvLvAp3oVBX8mI8p+Dgt6poTBfe8LKOYqk
+96WNh/MB3fVm2lYYIUPsayAfryR7fK8vaL0HWxl3ZWPEjDG/ZUOT1uz17qC2YUi
U89S/YenAChpe5ZAmJiWzJkzVsazISaxTg3d2JZ0cJwiY+uilW+15wKAeeZkGs0A
TTYvAvS8KhQBaVS8/1P9DX02yGOT91tAa3SjtFYgqgcZkjN+yGVzrH4JmQKnPTa3
lp5cpV/djf/3zlbhsmHvr9rxv4EoEFzlswuVV2GvRQr9UZ9sO4jLB/3Bm6yA1ZXc
bG/mGR2PSqxwXaoCJRUFXf6+mdcN0tJw4Aiir3P9T7tkj8qolehIKVqLfi97vCCf
RGH3+cjGfnfyxZyrOuTzyhPFIXCbOuvK/rfSKktlIGfBk01ZQio3x2N6iPDuNohW
61wYDDUFGlQ891+f50GZN/jfwjVZ0BTzx1odUQK4kknhPYupKPdPXLqwhmKjattY
DbwfE2RX+K3mTwPfU+4m1sg/ztdSJtrHE9gf+9sa6x05W6tLjtREvXNBwA3ZLt7z
HNiIol22ZHO3I0eHGxNpQw6qZxMHovxYpaTThptYCo7IinEFA0y5s/oCCzvGJaD0
21zOQ9o4qp/dTG4vtdDxqJWHqs7U43p1POl1oriAJ/eMTo4nPO8XRguTfkgJbNsx
gaFwtGp5NXS7LSx9W/HcwD+moMj4G4pFxhn/zqCnJHZLz0ljHkAOnGbHcS+Fw6ll
o2KmF3UdAVDmW/gLXkWqDn1h/Y5MSxSy0MDa03YGRGPrTFdkTy9MAYMzK3g2Hj7t
o36AW8i7XMMPsI7Elke9N5nMYaU1wy5smwrXZPQzP4noFU1flzdOjQ9Naww5DRQm
HIEQaULpopiJjM6bWNxC+cWojxLFeA+i5RoucfrdPqurElNYkTgjSYrVg3bPwoeb
+EXLi4mx6YtHdZ5s3EGhrJ2v7YtcLLQPTkRlq77zxUR0pa8JkG0ud/AbZprQ/TQu
BREpgt8ejfNdTiWy4suQQp656uotDkvgNIOQbVWZ1Wab/42qIZltMUo7DLhrSEjg
jfElEuqyJWoVURJ44pYZ/Q2CLxMag9UFoCIpNdiQg82YAJPkVYS8FZFwd4sy4owy
pnf39ZubA4DbRABh/oeIWe9sg+j8FBxY/23zmjuD8zp7xCmPFGhUZeMX8zjBmUgP
aTDetZp38U4SVCnb0/ebb6fWgy6Sq3h7OmNQJh/UW+u7Qy7MJwPwpa5VrU0f4dhf
+Cjwm+NzoO111jqJ9Y1xR3YhfE9f+MXIwuoQZ/YolgTgxN3hBoCMhF+TbRx/sCQ6
blxPJjVEnaL6ePGozDbGQNiV3FhBFEvWC5voN947Bm+S2Bs+T1eUY87KX4NFqix/
/kFNVmdTV+YWD/YyX8FtHmTMNJa6naWvJ50m/zOVjR2OYbM9+b0hvWEL3Hh0Kxdj
TA42MPNNJccHOWDHEvwv3bPCJSMBdo7CGVG/JJsCEVJI4lPb9J8Isj0ZYRZLJKkB
3n/rVF06Nwa9NJLOKXOPvtKnFQW9qIrRKw2azoxebOSgFhH9w+mqqm+j0wFirCYU
+4LWvrW2rdJWXEOZc44bYc5RbmYM/J/pfSQXVind8ypmezrfef2dg8azR+X86nJh
M/vBelG3ha7rt1wSzs+E3LOG/NELHJxhZVDoc/5WnSrERv7/LzLJR3B7E3KpclhG
sgXYA2vSapKVG3yn8dyK89xSc5a37A/KMYPy0JKNj+nNka/hhpGScgzoj/63ENw4
IueJwHKRUvHJ+8qRr8zj/jcz64QL0VMVuO3teRtvXualbUax+1Y5upPaUCRJaYaf
64sHvaOr3eYL+gYSE31sgYgiN/t82iWx9q1/JQ18rU3Evh6LGA1VXKMfunEVCO78
6ET/rhF1qCGFn6gIx2B3V6e/qMlvujC34Fi78oqrnTmEIeC13JZdYaa1CXWBKke6
4Zz/Zc+Q9eztkvqciHwrWB4RkbjAGDNFZvRNv1LBUmJwNj/RbYMpCScjaInOZ++0
W9VuuWf5mbD2wb8JC3U9k1lRnIow2s5yfqEO6pCNldORWY6qsky791890/ITLOLC
9emg09/e6ebWI/TOgN6Z8CNZ5yDbaBv/Anli9yx+QAjN03m24tu6+lRmCOOsxdAT
ChfBYXUYjIslkJbw6AipusJuzppkYPBAg+f9cYzfZ9OHsAOrwmchi0q6toly7kl8
ZHxvtjpon8QwJdDVFurmq7JrCwgsqgpplECKmvQLehqoCGB7XK4hiQ6MOWXaYO1C
+yHkanVqr3cHRQnGVyvOxsV/c/FYcL8AgLI9fptj0GVkPr9pS5QQ4FObvWR6YYGD
Dw9VFbKsXtcBmDBjWjgRLnxSh5x1ukB3NFyABhK1and/iyM/JOf+wBwjsJiBaMxd
Zq10nnsP6MoHDhj4b4+tDWZgIyqpGl8MKNHgiKIssDIa8P1S0JvvxyBe5mSVjUxX
kH0i7lAR7rURh9r3BNgzmSj9QQgzUmjCZu2xYMWeZl44si2RsRWhokeewYe69wDN
GiDtT0M4YulGjzeZtf1P9ymg1o9Em1VRBOBbII2mR628c6w/+uR+Yr8K3WMV+m7b
nt0a21+y5HfsSJMixqCxPNg4Q5BMux3UiRefjRnf/dBOSZmMeqTgKtwrW17QrRSa
bPn78GufNXOG21JV9OijNnCJSyg/sibRAofULOkx3RqWjM7iFYlWRAprXAB6+Gra
tjQQnyMP9zJtAxBrJrY/na5vFYvS8ADxb7q/wTF1DJtX4XSszzjgbyY4MPqUNj3H
WFMGQIIrUviKoqN5ZsOPb+9F+qvufZRfkq32IvxmiTfjbG15k0RIq8FO8Bt99lxZ
K2DoGiON/iCzmDaX2k5sgbh1HYvzQfsu7EL8s3khJZGaf79yNhoG+5cVvYg1Oful
85ySnwOoPg9Loc00l+TeyW+4HKB/SWfrtF6Mn5G0Bz48SQpzMYPZZR/t43DunwX3
lWIfAtvtRgJSqz+zoNsxKL6CwmTXOjbB1RHlkfg2LL09CC/Yiyjumd38CQ+mEBuD
0j4ht1b3AaL2JRgbTvW9+kEipM7sNlvmbBhA3r61ehlJ3Q1QX2wPb+5FDgijfOfw
7CVNF17PfpgH4D/O/MhfwU0VUBwzDSM4ItBGj7KQW4Stz2XyASx4EJ31w5Sr6Y3e
VDKqQHUaLqDLJ0XdP/fPmnj7PSNVOS+9+xJT3GEKMj1N7d+YO5kMD9GVi9CMotp4
eVwjtCgxIkfS4dEIaawgYxgUGAIqT+o0cNT2s9lIPh1Xj1jG/oCSeeyMA6wu0wmf
ZqUR5k3v669PUpdn/kCxocPTZUfXmhHG2F1yMQHLT+HpBHc31tph+/1V/9lSGMr5
qUemqMuTy0biVvH0CfsqWjkq5FmUDeuQcyO09S5v8EJwi+sH+niMxmOsOCTeMo/G
aNNE3mE1uxfFlfkOlXCMMMuQH9L6ove5k81mE5nEcEjOM800hGuoHjh1ROWXCfgp
nhok3qgkLRAwkKkfelWnln5kKl+C0327qwmyKNzCcUWMqADsmypYXVrl6w4WfMKH
ofqEDSQgxleDP/3DpyhCpaBRys/sFkL7UPGu1NC5vyB4CbCB1FPaywDBBc4X/b1+
ojoyNrrb5gf2cfjmzbnU8xuLYpSDsUpVPIELva4GSuDYXwxGsXoOb44rYEW0hj1d
NOm4b4Q7YVAFARuKHbTnGt/ts0qBWcytzA6seBTcp23+0jXoolNdDSkjttfQr826
eQzW8xd8k1MkwGDtjI75Q9z+X8452aAiDstLZsadST2zxbg6mwxEdXYDqmPlo59t
TvNVOG6RY+jV9c7uIFWQSWRfw7nxkjs/HnnjP4WUs7AKcAeXSOidZXwWODXKyz9E
O4+WqGNVKkaPACV6FicIUBNuf8lTqkxOWKDDjC8y9xFPo/rVcUy1czwwaoTB51ne
N+t0mpxBRb7ree1Ivpon3NFOb6nhDAXY6Pf04Qy2rZCH4ocn354Rvm39ABxASj1R
uMlJbdieFH12z6/ZiIDCJZlWGrc+yrJX4KV+HK7SxJZTWpikjA9MmrvBLgubcBdk
vzUZJbHTuczMiaHNPA3HajUP7B+pGA10mE4gCk81UVe7XjAYawaYFAE/AyXeszwt
TRimcfYDro2RLG1VlnIrA5qz4L60tAOrbdXXO06P4aoC7b3rTFLnE0EewNmrUsQG
BTG/H9GgZaTHn1nDCLT33c9Txw1GPAPPzPuZ5Ouy8ryUaWje+KLsSTnayFJ7BIXE
UdQLJ1wuFDxdTlQZoPY5olmNCebqev0OTo/xBZayl6R9iz6o28RKbc3s5qjmbGBy
zCTDYX4PsDtI1rIHxacK2m1Ac4pxv8mbvGcOGkGBuOAb0Wc7S8ryGQ4jwssYJLGd
1crsb6LD59/rCOkdc1eChR07t1Wdw16h3NaTmxtz07vd4sEZ93qsBUOUWwgYRDmW
J6Q2ye96AVcWqrbQ3WF6dmZK0EcuavlR3FUojKgyb4MrXMAEFonxfge8TChs74aj
0Ak5DTwYA9nfQVV+KdPIKt1hWQbKEzGhPEKn77IWda9oM1GU1ggEtRfiVogHg4/l
SFZl2E19NPHS8NdCGcV9Fz7vJLaRUoeXB2gYD+InK1qwF6I4RydU5a7kxU/gx/yj
Fn7Y+0ZOA8sjAJHs8gDn11wqK23JpwHA7mMGW8lMtjaouBeHC7wlaYdSIYHVbPCH
ogiaFnoDf4Y+MjsSboxiSq/+gSTUVY8uG9N4EtlkL+QmNcgeAyzxqt6XLGg2Bg6c
WNuC2MOIJ/elnhQ707rNXfWcybz8+w2lxrx80HYk7DTlGPhazr6qV9MKihpFUuoX
9DHvbv+VTF0rseyxKdk/9RYpaWiJ5arZrSQXlBNLRAi21F2FPEMzVtAy4BUkKg7n
nh72vImA/g8DnkaCEfD1r4+Zz4gnoBZjFuzAJnpm2MqBWVqr9Wd1GYM6yHIRbPBa
bP4RTzuUwBagyFl6qNIxUAn9zTg0L0y+1Kq3RcQg8WnyOwYXXU3PYMyKNU+AKC3S
sjguaXlmpoo8NmWaHS7SbN7IZrrb1l9qpTWLxmY/ObELSu5V/FhTcQcqOvlFlDxh
wlLWGHrKR1KZKJMd0k8Ico9deaOKdTk4aXOHfx4rEvUg5/EAo9oi3yZmlOgRdlwB
ZhzKRC6YC8fOPDJZajGwHvYddAGJWvsjYSvF1ThhuV0RGujnXf+vqxrYhZFGhsNp
WwS1BFoDkEvIKzRAvR14Rile3EKN3OUiSYV3dMDxBz4cY1ppTFNyJ5UN8XKPgWQe
xJBq8tglCNNFosIMQw+uUvPo3uIudcjCiwYqjLSpLEZV2A+yLmLq53nyDYPZ3C2C
wkfAnGZQ2fo3lrMBaAbyFFaJbp2NkUeBPI6gU4OdmGN9xg9QXt8RObt/ABJv88fL
2vz99c/2+NaqWvBCPgb29yACBWYe++BCEbccPuXdg9G1xPjhqxd0icThwIgaW1C8
xVtIIS4oJy7XSHUUVmVS+K7Tbzc0V2MRU5V8s0bKm+FsjMO4tvLI7czevPlBsrdT
LSjWwiDl6DmDhWglFSAdl0uyFX2oen6XoY5f0t0C2SOVO6RUODfpgcy3Vi5guhAw
2FywH6jCBBU7jKkaCgs24Phgm/mIOqUC+hL/gcuQ/xZ2O/Rh4c3F4LpaFLhX1LQ2
/qUuuUVsRW6bzdEhbacIVAsdljwmnAqtZobjEyQlbAu+RtcWU9228+2rjDmnCy9C
dzvCbwZFWJ5Onj4kcS8yzU3yaDhpclqfAcpJ9SAypUl5nY+TbpMZdkQ4sW3t0Tk6
6if47IOF0YS7uMHgL7+UEGQgMlNRrPXNHdsfx8QAIbgxVym/hGvFaRmQJULjqbvK
O/rTMwI+NYF4yYrGLWWD6SjVMK/EWPifKWgZCku3mGJvXmMR/Ngls9DUO4vykdIB
dQOvdZsbTnwwJ4oipilLd328ACuQoxum3AkDqc2RAXzkuUAAugw2tHGIozk8Nlpe
LMa/IKZu7e2Jx4qUs3B76X+RYS7iXNhjtHO4wN9G8eZMuZNN3TayekblenIBwrtb
ILtiQ8wgUMiO2Vlp9VQhx3i4ifnZeM/+wxr0SyZvEBkv15VHFGrYXhywndZ2z2pm
X/MP8h5NnZWle2L8oHAQkSMwc5d+UPoOP+hfUfQdW7XdHp77LOyFhF8wLEumtcyw
yBItIBQny/tJfr2SmoWQm69L/kZPkYCIyeBZ05Vg/Yd9Zh71FiS59AG3VDKrjA8q
VeCztncyLi9BP2kEGOV7CBWxfOStzfWQCfDSRLQBqAaspSuMeB8huc2aN1slS1SS
+vLwx/1U1/F97SvVYNR2gbxYS3iYkKV7Z6RtmuIvLfs3UXMoJPB4GbJZp4Ds2eH0
ZitvZb6WKD+grhCsoQrDZBDUg4brwXukOBhqx1AANq2faCxe8PUpkFZ4Ma5MG2xR
YUqEiqkAxzlvg0ILG/sqtpBewWAJdsoNiGvfgaKO8YQLQm5Msld56HflFrlVhrAZ
ppc/59aYr67mL6SPldztieXY7Mdo7pRVyt3bXXSG2DHt94xt+3pUZVRXtJsGyOQ3
8yTDMYy/2VvlwsKxn76OE/qpfu1ccQnKcuCt464wB4Dsi0oanKYQBQp0/33/FdNR
UBaNonGTbTtqIYrQNis1gFyRrEgrAITnYFRgAlxEWVnAA24pg9ynirA+gpcHDK/3
fbLiXivdKs0fO4BWgpmZfc7kQXkp20w9+tOuux8zu6miTgZGZ8Fn0m6ypN6uCTvV
clwMFoL/ffLLzxbt6V/F56eOJSGiNZSBfdv9CIeoc2OPpmaQtYtXQPAQGFK4ZJ4a
kyNSNQAlPH0TCJdzGg7tJFvPF6AF8ThVwHjOuFHQQYK+JsSlfvafyPf4+xN5nmb4
MoB0ndUdV/5FTAlLNwTfSbQiMEtYGawciVMMj2qqwRGzCKxCqNoMYMwFEt0bj2HL
yuxfulElRv3QeP7g+ci4ON0HWc/T0W4IQFGNCP7fwopdRhqYO5ueQDzDP0ZSdXCZ
lNCy5WwfRQs+93qSnzgJLwtcz9oHlvpxc4UoZiBPWCgxGTfhcBt0fZq/el1mJ5FI
OWJi7FzMm5uGjWNUcz7c4vFx8yzucCysKhW8EOe+WJHYdh5gkhizrpLmMDqe27+R
veN6svKzrM5ykAO48HXMyPTzR8GJC01oaA43iEcINhF37ak23sLWU7qRZtCdRCci
Y5QLdMObVqkXS68DzeET4Bk2VmuT0cRLGO+/9p11jkGV2SQcVfFJ/WcyRNK1jiXG
th66vfrztupzJ1HSWvWw9mCQLCnREwIwhGZXo8HC8JuUx/zHaOzHCQ1dmM8Ci1jR
UBF7YuVmvb+msSSJaNpXRPIkzdtutppkhf1GnhGGv9nZ+U67jAFkJXFY7q9jAsrw
C0qEfloS8K1UHNg05tmJy9KLiVM4wb2yhaCgDm07WZ1lUgvWbMt8prc05i3j25qa
p2V0qbrI7jP8cXN2LEa5x0rhjOENhUJUzMo2qguho2cQX9uAWC30bgMLSm0fV+jN
mRhHjHeRXfdy3Pcp0GDBkKXroGe0R2x0wbHmVfHlJ6YDIhrpb7+qT3G39RPMB6H0
Jp3eXXgA1iYmR0FCtEF05HBe7njDscj8XF7m9WhXR+WRd0XG4uxytYCBxBnxW/0s
B3GZkHlMXeZiv7wMX94RkZlD8AxfaXgtifYsM1Ji0RIYy6otbJLH8UVpjJ9zXQhX
2XAAOrcaMh9FUYvACTj+T9uwzD906owFNiYdLkNUs6x0y+Q5Oa0FWjt7QRGu5P9r
CPAO863upCd7GPOdp6j9DQ3BzVPtcHCuMgMo58WE1NabGI7WvTjfQi8PDJlE+kMV
qlmrKPZBQfYfySGXLqxUDAt4z1tL2lod2QdaTYZDdT/s2ozPcCV63ZCghtSQviUr
h8+27+lMaAlG4JwvoYIInw4RgjUt0cE/4A4JdkljX4m4p3R5+ct/Eao1gn6Zt41W
jlDMRKxc5//UE0vn9ly4mVaStLL9RL7Fzio+oklLgonhXBe9rkhR1a+zvBe+s7mC
kwHWFcHJ4X4unVxUIKwZ+CmCGvUH3iaq2fJjDoGeWL8z/rtrd/N5ehazQGTTsI2P
MFz+LG50E/kIh1zLnoHcyOY7B4kq+GYzHeanG2KnmBRsqHLKz8gmjHPhVNb9YsJF
yEiFd9veyz8GOhzfIVh71czSMNPs0YDA2vrLVT4vXtN/j782I16bZ49++L4jJgDS
Aq4Ts8gM47dXv9FSiqjuAN6dlFl1fczJ4nCvqIgdaY3leTmlEAbdoS2Vs96dUknA
zvPbwbHcfLMvwI5s28Rg5KpfNRpmAkJB63EyadePJH3aP4FljoXq8N3HH3sDEeda
dRvDo7xHAM4H8tUHYq5YhQr3MvBgWavWV7+JVBADSIzyckHi6nqVcSmn7KC4UbTX
ANdNvN386YWJ166STmJfBdA00UbwPrVBk5+8jBUT1Z3FMmt8iS9GtZPdXHdmHTFb
gcnTeD299RrBIp34KPz8iFimI0KxHRHF229bmRQaBxjdek9cOYawqD9dhbFDq1RR
9TynlQ9jf8THNXjGUW3csrgO8F5bYlaJjdmT2y61V9aIWaWJHtTzgyW1ITHYH+Dj
mH5Z0FKWZxhAUJ5LzbxWJloK/Q2BA3N0oNVcB+k/2Fha/HhMmjhUVDDMhDCiXwUU
4TWHdHoa6rssn0ROwoGD5I7OupNA2XU6qodELcKoVcYmPD91++GbNI7H07gjI6Rf
c6pSFNRCa+V9JNfjL/Oheee+ettn1b+liwxRNHeUDMX5rDfGFTfyw1Pr7a4A9w/w
1MUxg1Etf9p6ZIQpIuXT9aE7y3BP/hT+QQT2twX3HxdVeUBROLLTVApoA/lnlXLb
XC5eyfjC6un1PMx+slOeAtNbTV9/sy8nxsA0zX/v4X+wb7pZrt/2t7qJTPcpdZWB
14zzVUOHiYmZLlES1dHwxq35YY9DZaAcMrwmkN3brltS0scCYRItNPPQtXKnJ6Uv
hqTIUpvDG2tBnNC+DgzuyatSrCkhScvu3W163mYkNmpCsY4RApAGeWl6MQBcd19o
GnU9L2aqjCSCQg8Aqa2siHb1CcSnudGVh+WHYe5oHk5d70bSAXF42aDkGVNB8QEB
tOyCQrirW4vp6eAi6jJ7EWxZfW8EGx6KIr4tnGrsKmf4BlM1as/3Rq/gsjwczkyl
ij19s+BtVIat7352b1nNFwySesaFbFNWgvnHfujwQBdWLBp2W9+B7JKVa2xjWSr4
CK9msNkeePHYIOhZMYGbzmzqbtmjvKSW/zPhPTkqwLxL4MUQruSvx/8bP1jLpofg
fUjFVqzBdSdySVjOZ/RqwpMj+TjnXepaR9LIURI0YEuIY84SJkw67NCzjoxKI9Wa
hKhNqOIxTSFEroHnsRrn5XKehJk3DZ4AOxxHhU+ooUgJUhOMZU0HIK1u/QiZjzlL
Qsv1rOvb8/LAdXETEk2Fg6wO+lXqWC8YYsbPYz6zqisEuWVGYHt1k76igOmoGmZy
pZaFB8r2se7mtrCrBQkG/EwHAznNLC9Mv0QmvpSgtIvOe3ILeFh64B+1eiN74+en
8mlziTneoUPKEBCYcQjuaqeq3dMbGYbOkfu1724UNDA3YLBY6ctRvMMydDJ59wbT
g8h32dVlpuzlyHEs/6bkM2pVHBPjMbcXnQmfUcQKf5mqCeOCj4tNbVuB9QYvty4L
YU9mfo7zcN64Vf5L8Yk8vY0YtIV4ixdm+Wn7szrG4nBB+6G3nTd9Axr8GPveuQg9
w3F6jRN1TqeZJj/v/0qbkcOOv2Ge6aSpA10bjObSWXQNeb6FXsUZOdaW/5neX/fF
R169P2NzYm4IuHDn/DPrPa8TnOgg5OBY6xnC4SsG8gu0EQfYBbwdoOGhVfnYrTfF
2+3ahAls1F2YYBRAMuQniPQxPoPioM/8PvAhC9lV/VrRwKkDqEu3AE7DzZa0FK7s
bEHxJpZq04lVFmq7bT0ALwFcmj4DYSwD58ux+9nLRfbFyTSGM2suPdWVPMjYtL/G
NFlMBjLzBGH1L7RxlNsViInRZgYM4NonOk4RJ+Q9qPJ+lfd360kCslZxS1TXbI+M
7dkZjNukke6PtWTkJ0SrwTGtTfoRdzjnCMEBcgMipRDFa5wTvH6X75PHYicw6edb
ZDfNevMMkh0LnnVMO3Hcv1SJQ+uz8EzN+Ry8T+pv+PRVt+NcTDnl1aMKoA3cR5MK
FiFFFoqijuq9YbUQzskFC9zIZgtqmCtwn8RW3ImG4Bob4HOB2bBz1viFiU6k/fyT
9mJ0lmyBz/NsxtLVBewY56VrMW25PoNwAIbjfi/oy0eFp++HVtBO3rYAeyHhCZtz
Wt780f4eTBwLtT2Kpiq51mtUBDAXe6aR4oh+wTgaVOpm3Y38IHaD0cp61D09PRu2
mQB3MogttKtBDFdEkx8dnNtAof1oK4G7sbEN/EgnHsq1N7eLPdjItFe0FuRVMCEf
dpG+3VyKBx/v5ZX4YsrEvM5jZyDjjThu6pW+Uj4lVURrIvr0/nOJpfbDx/ty4vUd
SbSYgPzPTE72G23ctOaeZMso3EJYzo1HJlvX36iSS7hSrF1yDzGAdeLAWZUXYt3S
JAtbz+3SDEo21xE/cQ0J1dGnhrGEKuALevoaBhZjJVRBBZM/AKMYTLOJSOPpPDuf
IHXnm52OQX1xyc22C9yry/++e3YTlXZWk7XtEiPS3yxToWtzr07sN/L+48OhG64I
R/+f7ubT6oFxyb42TsYYjrNjys9j1YYAxhOLoui2LvgotmBEwXRWwwEn+bidzMEU
z+oXcwDD9JHyL6/9k2tY50QEiY4DYqcLSreZieNJKZ8pS5HKhIN0j6BfWsroelE4
lMamgn0pxJY6FOD5V5dfFK0uj+6EPMJW4508g8OaLRyXGJviJMoYJYhmJ6HGn4mc
V40Zd0fHdTOirbUi0ui6DNkjc3lToYnev7D3sMLmB2Q64TAdbd2JwN3ZyJwKMVDX
zUG/JUWUTibslTL3biEPJfOp7oDkV2kicoBHbS+grTauv7zRLGi90jXxvjgDYdMK
xbHTJ3pyNv5T+nJDa3uXn47kA2ViObPbZtGjb32MRSOtaAl7jaz2IXqx85D2+jrH
OVyQGDrPdEMrW/AsJZuLoBSkT1pGcCmaQ+zazTzwe5eciJ2Ka4Vzpv7wJR40MsTW
aFk36OteBuYe7skONvXqOYbz9LIoEjLaCyP1HDARr0ewdW3ZU0DaC8mYmgH+zrFf
rtMmW+MEbIIM4r6KV9NyyVyWEOAbAgMpl0/fRwKpF8oW6v3DqxRW7K2Sk6kAD59a
CKD94y6baOzcA3p4hWZhWxsfGA7DQwWg1ceFV392rfTS5VRBlvtb9ee/efft1cy8
dPYAJxa+p9KUit+q6Hh5HOMy2eivVHcroV7dUP9zb8J80DF/VRNfc5G6slbpcRjT
Kv+6Nfuzfw5pI0K9TIr+UfjX2psB2+KasHMytN6mUPbnVsyu/bTYW3Uypf/1LFJe
y7JqmUenRAYqvouxEwI+UkZq1I/Y5YKH4hEvzsodjuih5zWL5aP1veuqmSloSO5J
6eRAAE7cKs5zjZnymKXh+VLogdf+66h5N1VdSM0s3waaGt9mPq7FF4RR8yuHEzVV
Aez2Zhqnh2+rRAXe73J53rgrutLXDA6ZBbUns6Dal9lPxculPVUASVnLO47t2P8t
yuwcaTZmB2UkDfyLw6EN/x7hcb4ccnKPrReWpXlBC9etCrpIBqAZHQRyIEE1km18
C+HbOuOd85597KdTyoi292NFvG6sgRMYrxPIlV+z9YUubcccNDP+DLBBmhSMrwdC
NY8Fl6smkqOF+u55EccRF7eOrHWYRolc7cquM2TvrnQIrQklm17pCGuvZdVP3gMR
uKjM6WYhkBRpAU8hUsjFrpeean+BQpZMi+LP7weQkL0PyD4NmrfcbVx0tV9UemtF
iHEHI5z0TJ59iRdDgDu5wXzqPw1cfl/CoOJ+63nfsFt7L8bJDe/nrfOV4Jed3G2l
/tKeRpwUo8c3h16If33W5MGHQqcYWC+Ed9rCyjhNKcfxeJanbKeG1q8/BdAG1ztY
ESMdzzLWeqeN6rM0eFK/YoFbEm/WGkLLwloTlPchFUiwKJOJ3DnFkLtEddeylJG+
BIyKnycOTfFq1z4di/Mn5UvH0dDGKx7KshgbJ8iiMeFRo0vgpdx55Lkf3wPoqx3O
tSeXpcDZw8kWLqLF7hx2E3qvwwbEIfB+urvuAOqSeXqYkwbKk71pmtkd4acdOFge
7EnLAap+LMstmqF4qDLGcR1y6BvD3HgC3q5ABu4X9sO+GExjUjxpnnM++QM7tRPU
WkOnPO/2IPOIlqL+Jluf5KeE75IZTlf2qG7vt3B3pe48My/3B6mfd1oLemAZVzSH
ZjtR/lhBE88ZSb/GgjthyLaO4lq6bBO9V+sA2tBDMV3l5cJD3AZyLZnHYLmKmQ+L
txqpfgciBj7LOpllq3ocUzePjo/VJnEJ7gmPhAtS/C+zUltsTwtRMYiSxx2YMeEF
2Sw9x+4LL16uZxO8K35HGv+rrpisrk548kwq19yJPyqYoee/wshGB7MtDjQ6ajV1
M3Ph28XWWi4m8AyDLWVmjvfKZpSVDZ4tnSe5pe4xYwn2TjTkGoA5eLF+9/jSYXpz
AYffj5Uuy5JBJ37084+LRoVO4qQpQDXib5KGPRRfmjiLaVPP1+ut/zvcXriIY0cA
clRyNExzg1shC6IxU1TK1k8xAc3XycJnjK3/rIOYu4Qqk1DOD75Mxd9QXOqts3M/
jCUsQzTJAsHkDbJ0Cb9chbrI5TPnXB8UWgCbXXolKVPwEyDvlBcGoSbMhCbY3afw
PO8fpNvjKdxFgByy4DV/+xA+eEudrWL82AnsAZtvzQxTVhaan7buHMRFBdBaMkFJ
UYNy7MgTieUMp7BkmtRuWr6g4y+yxyyJkx30+KLinWAHVtPbJCC4c0ST+n4vops/
tJFPSsYlpVI8CXdI/0AX8pFBCh2JQexyddkk+55GV9nLtYYxwNyoVlDuHoHgvIqB
nY/9Xw1l4YHbXCJpRTmCV+7A0K2WeYVxK9wdGIaMsg0LF+xp600Ii3ELhKdpN5Z+
wD1qspZzuUhsP27alnLuenPL3Vwxx/O8zKBfrodfSyTaorvSNTljh4cLEn35CCWf
gIQa5HbLoRU5jXYvbfT2FJ4g1OPSiK+qZh7e9EQr49zQRmfRKzqE6iNV5+zeuM5g
u0fE3fCvpyI7vO4g9EI08AdPS1AEIGdCGzsDZw9VE6H4DeCWCYz1A3TmYI00LI76
XBllkKlPWq2GrrBWHjJI1D5rFzBnyzkZpOYIXEdX74rdOtw++e7HAvtP/gk7h+BZ
FNtG3QvhGXyKDXVvsAvTIRGhn3Rn4nbFD0jdQU/HD9JdtatfXEjzJ5GOWWh0XZ9+
zaF3v7N8WRRO01JSMJ57wTNEXJhTp9hBTsSFKrIgEF42mU0vV+Vxbl5Eog/FBb9f
kXAEvvYTlOQzYHSq1Tq7AnARuVEeCu6ORvTe4PPsRzKBF7exp37BAVOi1+daRngI
6qJdzRsm0rSrrNfeyVMpRaSmQKpbYfkwBEUnbFNOJ9nmkxwHRoHh1GY0Q0G9BZgm
dy9LpwbwXrnpH1NvMZzOI5/PuLuO4dYm1obn+8cr0S8/xc/mJjfk8gVIPT6OqXdZ
QYkTCV8AKcobRJ7aO7O+9A49veCHOPXCYu0Q0iZ6Tw5LuAKrVrlGVGUqxtNkZWJS
CFc/YAXTovZ9mggJiABdkS6rKZbhtdsGk/SC/IrhAUPB7jJt4SPxcFsgFPhilA4r
LhJinLIRXCibsl98vI73wS67AQMyPiL0XaY6lHReSCMvfpu1eVWcboYwsl6LuSdt
2jGlhbYri+6BnRMPwXiGoHUU63TLPwg1vmJHGQNvdgT/zXXIrkLn5hzSBhsVDH8a
+Hn7ryvPGp0ol4+oVyiDMghZ8AmYOwzqnryUSL+bP6ryeyuW7KXOP4TnDkxi1bJE
ltXh+P6q2Uuox6RbeRHQhsZEuggUM2pMOnmNQGQ6BcPPSYKDityF8jPEfsZMVsjp
PDgeYfFZxUhinUKpbh82GIZ6nECtdA0UBPUDkEIGUWvGdK9sT2zCdQ4SI3yhLk3A
cSa60PLD4+xTP9j4mvmjchsHCt1beNjfkbQOYecD4BCRL6ma8XEfJ2dQkrIrQk1T
drzZTclfSofGAsuxhMi7MCaAhPGKWLgMkp3Vq9d8ZdHGAuohJmYpILQ+GI/r1q+I
rQb4pOd17oDWzaO3AfU6EBazfYH69eWDjOVEk3BNf8SoYQsrnfwZaKzeI1PvF7tn
MUnER/CjK6hEuzkuGDAn2WKXWfPAciUC43XRdv+ypJwFZA/wXCiSrY6kiH5Ep2k+
G7h7ggzCQrfrDL1N2NiUScMXwNb64DXYgMs4z1EJgxIsK1Hs5MTr7vlq4/fUJhaS
ONc2A5Rs+p+cjB0k6lrQBOIgvD0EfdnI8XaSUH/nsgAinK3+FkyS0/F3hymC0FGc
XGaN0RSbtlpfgDDSt7hYhdf058+rqfPZDEK9qwNvFzNvQexQSBBO0NzqxRm8yuj7
5ywHQFX6nH++pYxGTUyjeJ8E64cb9KzflPnZEGSXutFseWUv55w8FOi7SbQpL/7N
R7k4R0jpPg/ApsDGYMuGTvb2PLVCSThaRzK0O1TnP4NWhQMj6lZpWhqKdNjNqW+o
RoGIojSI3eJJKQJ4FW+CtHgIh7yPJ/FbNe0s19jzaw9Wd0la20RwuO22Z5EselY9
2P6KSdy7jUrKorX5Y3GHMwlzfJ0X8atAyKDGEiYkAOkRZ4j2sbnFe7qJ5VozkwwB
6tI3xzil2h9/rTI7Jh+/Gf0Nx/Un6//R01fI5EZVQnJe27lJUr6hNGqu8BetU9tF
sOoFs7rBoYiIU7z9o8/E1KLx+7OV23ejBcvBNAWpEazEQ0B3uYYkxL3EAVi17BHk
h6ZuqDYnvKvUMOPmecjV4fw/gd3o9/8x3KVffeLI2co+WycVw8YVoMVD4HZ26q5e
ICKVINagX9o9Gy/Y3AqPTPpinaCJFqyEAdJ8SQ1JwA1Xil3/JlzLi0WD61/OK3ZH
zQ+TF6/jVz+a/H6BKxTc1tn9EMOy8EA07puH4oBO0gpEiqMVt4R/RI1mlpevBHII
EXwmC7QzijG1ojUSOFXNBPK1K1DdK8feil4S8dqYrlAm4aeK/KAlMKeczniCA9Pz
EdeajYuLO14KSly5iiXRq187mtVGW1go65HSbIAKPMFVUw4SjURh4cqpx0lQNEzq
UUrlKF4PfxIbX3A19vyNV0i+lVoPhO/8x8YBljKs/5jDFYI1Xc8Zxx0ewPGCy9xr
yhJc2G3GWA8qfX6tumL5PNsklM6q75SbbN1klnNe9yBRwTr14zA2i7hFwwiy3RWp
RDyhv/F1UllMclQ0vsUEd6UZeB7loq7/+UHhg3VSiqxWgw37AA+Ztg1sSoa7xgb0
17YH2C0dCu5X2s1hJJuQyqTRqD2/nRj51x3ZJ7Fd/aETU5Mu1xfnki03wkPDVAL+
dzPwHl0qdIeUpthLcpAIbx7VrDoqpG/OSszMF1iQMxxYuBhS/vioaQPjE1X4LBzD
vL6zJZlS8QLNza1ZwlOyoEkuyMdzu+TwxX8p05NSkRvxGrm35hIftLm6s2tBc5vo
zi3M73R8Rq41UN3vOd6SsVajHyecBtRGXdscQ4D/AU5+EGVtAjGkoAGPY/e+05eT
PKOj9Iyfd6fWWKNG322pU9Qxu4BVn5j6QaFmop3VnYPSAYgEpTjmQWigttjzBem0
HkxF3dLtnsU/yK++ZiaSB7D7P/6ArqtQBwgwJzUppEDVg5d/7wEe3wUtBE31NEX/
jDUGq0i7yB30GJbjTxfcAVzjiKx1DNvuxHhnxtJes1iW1jq30FKXKBjyga65f/OY
fzTEFuCh6G2cMrCdEtCsovEcl9I6GqIphVaZfrh04JOXjDO+HirzlUt11gAxTzxU
/pCMjxZQ9A/nt257f834SzqDx2K8EaYuFVnvzqEl/YcKlhNj1FbCZ5sWR2kNYRaI
C4bmDHHTHmmemXtMNd+pxoLvZRkhUQ354EhbXXmPMs+7U4i+HvhASEcenyu4OdlT
DXbA170hYg9fdGeLXjS7Qhy9BuBp8q7AdQ3aUnG65oliIuS1zeUXitgfx/NnXpa6
ZUqfi9xHr2FDV2GLuR1anDw/m6pH4AwT1nuC4cboNzwu3dXq2r9TC/vuFA1DYC/t
1Hjr2npLt5nO/1CsqoDDlkQQe9AfNsICPafhI7D3dgS1LS7OoCkAEZDPTEeHbPhS
YFux9ykkVVzR00Vhic5fa1kyLAMTcf9u/0i+ubMRoFYWtlt26bFqBVcOSDqItATB
Rh/QKIRLnQZjSpWo5og3ih5wunETMSy/f7aI5A44i95B9jkFqeKy26r8lC3ufKT3
J4RtP9A+KAzuB8V4Jme5CMK3BEzxD0FJoEcTD4i61MzuoaX0jVvhXlNB6UK/oTIN
nM4hs2Afee7oRtFj93opQeR2fhG5YhYhaV7OfVk38R2KnkYc/G1sN9pbzeiaFWLs
p02JGUCfI5XtfQb6l32EH4gNXAGu1A4/xnuIsO8mqY+vDG/JAxr1PfBTM1i7BW0H
GB/Cufa0+1cZAe2/7OeM4Aqm0QXPtELErOVXcR3EKA4e+BmJqlU+OiBlmy4pDEIl
KM85MAuKns6Lg7RGxU8vmEHMWiwgXcW71GOHnjhQHdv3xafLkZB85TZXwA+eWVYr
JZaHIEFj3bVrOh59SiX4cb696hqLt7xQDjDv9GXm3i3V1CfblDODKqmBKYXXzMoI
kxqT51GAOyzQ/eNWe5wS6jJDPphnHW6D5tmWUbJvoZmSXrjzpblQ1Xjqp501pjBu
bsCyYTEqs6/6YH/dNtb4Rmm5kNKl/dOuejZFpn79aIr8cQMlR0POsy48SpBmSLuC
6ReRwmPqsjFKeFL1cgQmNfEkTNZZ74/A146ForX6Yh5yf0W48qzsbrX0OYwjVyJh
DKCROoR3rfaFhY9833AZCTSv9CiAuJFWBP00ccjSo1xY+hLi9rzFIpCyB/j71Ly9
D5QkxwLH4GmbNrm/t4AWGE60AshmwzRnB8LCmHbUHbmA3pwhuVD6iO7gRzcu3FsH
E8szlwruaCFp4QTkhBJ4eWVVWVsK7jPxtZ9LrWrrC64qixvKFghcpMudGKTnBX3n
i0RswbqF6RsQud+FgXYDXW2P2Vpuk0EaE6ywgC93KARbO+FUd3FiVhoH0t43+Z/K
hUCn1Z0R919rBRmB3AjZhX2HNZBbf4B/oTWQ4jfJy/0Z8vmDqZ1m0Gk5YB67uHfu
zLkqIDu3Z01YVIK7mjecBCWz5XWZZlp3GC9N3Tnhvk3T0D3SlbRftezARsFWSuTb
HpV4m3h5Xha9kqTVH8GoVCH6taoD7i66U8hjsAHtV1bS29SWXTsDxOPErECH2JH1
AJAGYs/9wnUBe1t3AV3Cnm2ocTHW2hndEXc55bO/XbzhspfIrQnoNbniwxo8Op6k
OmRW0lhL1T/+f5I6uQBw0BaiZYoB6OVWv0fjKXC2sXpE8gnseG7lbxS9lYtPT+7N
wOAiivTigc5kzDBTIpEhFD46x0XkPq1aTxcdaANURX2K9sVBz0/CrwAv1ThYYOAG
Gwk4U+RwfPtMtHGr7zitz7Qx9wp7CvdjV5CVidRAjDIxC6McEsawrKwrUQx2+YIW
QhvxI8O03A8CvssardPsLFJGwiW/0ptSJJDtgBSUviVgPXoNsz6s3O08z+VNfm4m
Fep51GcdxKGnB7lh/LRHUak4IgC5taQabvH5yMvsdeJOvsGRIhVeZGX1Nq1IEXYa
4NQfCLaDTpDLx6cqWh4Dss46Q2WYE15v93cOvd8cZB0t365wCF39e+K+YbAfFk9a
RQ/RQKt8u09Ivkk5g4/g/KBWiH+ewVfI+jWNvUSb+CVlSCweDO8NstHS7L4OiNYw
qrCFTO+zsNv/mNdYFOT616a9DtXtXlaQuTrmMEArf9u1c7rA88ExOFwR+8PK9Kjk
/ElJpvtr10C+So6x8VAon9NVQEnAD8U33BG5JUCaN24dFOm/BXxeOxxzi7urkia1
2He9yAP6RMzj8Km7HbIG1quCOLQGzG9/q/qSqbTniVJXfvh2pkDOSArVPur3sADu
sJFI2BRQp/Mh/tocV9RSHXa8sbWIfGrUiXDTVm+YaO62asYRKuV29eSrxAJWFlhv
x3LgZK+8SUkRK/e3W8K7bc50Azqp1XzFi9FbgYBwBPV6dFiNcDrKpuZ/On/DBHiz
tcKeEAI81IKl30V3SzM/MqWro2vyilgD3nueEU0j6zK7yH9++FK7Kb3tWQnJCLzP
9oDrbsn2sATNqFqxOI8z4mZUNwFeaOJvgU8yLYUJyNHw21hTrI2xc/YEupH4DREJ
Q/dMEX5KRU5CW5Fc+mmuoIHoKdc8JEDFIMh9mfDu6mlQvLfRiixvAAa6xf0tYX5U
lRZNjc2f0jDDSk8To0GasjOYkiT0tH/lztC8AftuDTlvJMkhg5OyGjHW8BQ742yi
l48XFpapqklqy7Gu0lJpaclbryDIt7/foLOSpeTrj4Tuf11DsrWcDIMZuuxvhpls
N/l0FxpFLIiR71+Rt7c1cBWSDcESKWEk9iAmtsuYpl8AGMFpOX2wHCXCXuvf8vxz
rkeGLOvL7A//NCG6SYqRE0LbqI8UDNscRUbHDHVRMlVV92eUHlduE2E9HMxUHeyH
h5jDLylURu52tSORqyu7vKnmm+9h2dFFxZFdKb6Ou42ouJSzHObGPVXqkhRgHJBs
0GO3fVLCpkdDYKxXIGtRFsM2WgNz/V2BYabo3JW+BK0bLQXiyyScgxmceLQWFrHW
Ezpie23cuxJOjT4OW3l9/Z2CviK2bUkH1pCXA1kJvHIi3+mMxQHFJCqIYscT5Lgy
WBCIwuhsKX9oACfWMluBMqDvR767Zab/leaY+r/HfEY28sxyKK2AcLL8szE/yoZU
ut40s7odQMhPzyhJMoOAjqh1tuA82LuYV4zbd4bv3EYffRhSIJpa0Z7CYfOrs2fW
XEsecsj+QzaIKQcw80os9RhNRnTpCtJNDdniHe9FulryfDq4LM1ztpEsrpTks9eD
zBSW9+A+oc+YHFzrKuzy9L453ybq13dXRKPr8rQy/1m9LGWDK5+AhunhO5wS2Ps3
ps2rrPw0wS2CcljdUyT2JbRQZ7hGGz6qFtdLNdp5cSM8lYR7p4+Ij9ZgQ3AeD5YK
dfdV5OPoev0LYgNGUQKfU7txcnp2u8RCl3IYoJZT9WpJQSglv9oB4nYAyJqWg59w
F6I0y9+mYIoL8BeOczwHDpgo6c5U+DKf6LZF6OR77KUScNpRwd/agK8VbrASxkOY
xcIgarQtFOxws2048WFpvvtDmkElM89Vwiu4J2/NTIJd30hqMCCK1whV/ybImAKI
0eJS1+FqWUat2KyLMmZHMrSy7IQTbj1xGIXJ7ZDvxkoLLjjxg2IThx5kMAfKFNxK
3pUPBV8/kweTvkbDLpHer1Yhm/JEkY3z0WVir+JP1h0MxcxubFjlnwNF2L0DPDhG
Ero2258uF+M0TLslthmpqpwT2NDU9kK5p6RyVtdiDiJIPmSzNQWLCAci/o3k968y
Mue/Y6TMKSQLJpP8/CVtRA7V6zR+MceuG1vhoUh6i4/qVEHqDf0JNH67652ohALD
290ktESJLmgWmnugcPsdp4u0igRp6Jbnd2/5kz9w5ZD4+Cm4Z5pBJddpHmdj3j7B
AjPVrBC/iAZsi0l+oH3yps5YJpVGeMx0+Js+m/4+CZR868KdJHaewVJGG3O5EymX
Gdk7jYIKKoYzF9zm1RL2LXwnwOtdGbPBkMmcaIsf9iPoCiN2y2Y9/27ePuxTGMJf
+/XZ8tSq8xF2VRgPfDUGbrxrKIhXESKx9NKUO8kqeYQDreQjv9ZA9kR4sWVwVAtA
AkkiHSvsj+RH7K2imLiMsSXxP+K7KM7hyAZ++k7MOvY9IQX0RgMnhYBmC8a/3bbQ
2YzsNBfcgXzuMVEjofDkGsBVl5a9FyNKHB+8uUIpQoJheXz+hRZB3YsrsoaPs4vm
faIXO0yh+xB1FF8nNsAdyX44zqtO/4AYhIWzJvq890jV4kEMkJUrZbpcE5YJ6Zqy
W1CVZxLpEEsOdS0J0QgA8oZ7h7WFmu6kNzMTE8DEdDSM/o0E9sQn8vUkUJKfT6DJ
miPOffyQt+BveFUMg5m1QMJjVCgmyIcD2NohKbwyDLN0VBvQ3SwQd7WMOCPXRDfT
9tiYbSyx4DOAsvofs73w4bMiFV/Oc7iFMc7wzJyDsuxk1z8OVHFaR/mOKgnW1h+q
AOvOJLdEb1eHz8nEep8NDHpS9sDemo1rmDgNT3SWRCwGPp+sb3olELtc3uBWeAxV
gvpDQbbUB1FQAIABhgUii9O3TjER6t32fg7sdPXjsnBDcnfx1sGrhR4o3UU4cjQQ
x3nUK/xRbhpqecncekqq3pjUBwmYRTM9QfRVS/aXpkAeCqy+lf6Nf5IB5K4jTrDG
7/ibACej9vsIArwuntKpZIQeISYDPVNWUEQAMeD9LaZpYGaFGkIuuPNFTOFY2cLl
qf1QPlj+3/mKisn+jtuRVyOIFJSrNht/FIfIj4LqzHYfMva3Rj/WUQ8JYWH9ICSM
qcTWX612DI4carlQhoOXfwtcd+5BauHOUGu0T4QjxboebfeUcK8ZvTQJgEMOmEkx
QDPQbxdNbBT7b67wsb3rzFu6AaEao67oK7mzO2OOK3iHc5n1b3vV0SkDy+oKimyx
Mb4lwUS4oWGb8TkEkoVrTc8JbbVq4wAozpoi4j/qMCKqdtMbkqwOGrCSoYXRxMDn
8IyU0PVrkfb0POXDqUQZwG3rc/N15XLtwIs1lWqErdiM9jvUUslXIOXwZpFK0I1l
ajHf9EROcdI5feAsgweCPotE2lrtUQJFK/1/1CfBQxKeowHupfZP9TizPmbvtBFG
jzUJv7AV43+GAPJe4D1rWIpP97x8djocxHKU8dC0hg3dRUxnAGFhoCsHoF4IY9+G
fKQ5B5IZ2J6fTtV7lFbum6pbHkkFS9Mk4HQ6rghMojSjrmJ1uRRV0oiG5no0jCmg
vqeLl+u71BBFvPbme7Lf3qe1kKiXOIFY4jrL/a7OXMRMHq6jzRUf4ZqJm5YZrSqX
dH16LcHYLLcB31IBjhy1JZ5hV0ssm8tNUWVLLEA7PQEkldxkA2AbgCdaytU0aJL+
EKcNWr2vt3UaIKb9WY84HrNcw18vP/BLeti0UF0fJ6yDJsMTB0WqBl71yXJaVIvx
oJxR6FZFVST/cJtoDWRuPGSxDreVN52YXORv7cmQh8XFTRWbEuktg6s8pUusiT2w
WASgvNv3BVlzJh6ziBeGjN9daEtcQmVFiv4U1rcdaP1/VMGWXfrf2TBbwwDTrGXB
De4lECgWuDwFSFoRnH4Lf7HMwSNJAA3j+xezCjxGcylN32QQpPsBQHVVi9KfTdwB
MlYNbckguLre1EG2ajj7uHKwKnCs9CEZ+nCFU6y8t5sI08ObBWCsN15cFLIQA8/g
+bjBwKQtdXX3WXTmrAy8Pkl64OJAZfdtGnLjBCjwBCJh/X9IXmgqnfrN5LTa5Q68
m5jTZfCFytGpXf7gE3Sxz1tRVVKFK33XHFaaxXPKqAmcwHZGs1UhekMCmlTVPr1C
6A4tytSoVMDfQKlQh2mGUJauQIzMV/0cO6t1INRTe0hTuz2fW1Knrg/ODNbw1iBD
bTNNGgk5Wz9zIpJxsSY00kYHmJ8hWyrre9e+Rk50ebeTQs1V4gyRuSKLJXLE8q4Q
sm8hylkpeTSZN6DCUpUQHyMYkNaAVIM0stxdoApQf+k3aXdP/HvE1OYsnJY5DZ+N
1iiNplOhW6y6Yq3apep8RdOPLZO7+0CTROVFh0ru5lYsZfR6Tndu+WdsHut9ueQS
dl0rOUzFNcAUOAVtj3CiC3i6H8sZR98mBKjAo9Vh9QR8knFH4UNkTJfJ/ZoaMpbG
8g8/k7IryVXDcrm6f6Xci50kV7aVQ7JYGt5RqV7tR7mhgEjajpC4CYE7TcdXWa1J
CeYfshUmgAoOvdDCoDOoZbxD9XDDKJ76cdHtiQv1UEEyMs18Tfw5a2Xw9WP9vzqr
XaDTu9UfzfIJCLKN+F71X/D4P51P3+pXynR+KZ4cAIVqRyEADlDSmsK3pgEWuC7q
cBdk/G+SXUaqHJKaikyJTwksRiE9wTLyLi6J86bOY41Zjy9fSCZy47pzNBBPha3p
YxgNNcm/5I1qa7WJ43I1n5EF/ZqRs8UjFy61IR/aOCc7jFYh5feBr2WG7nLKafc1
HiMyIgvXEpsDIYczHuwvDpBbp1SXJz/6aYhN14/XqHDw/fGwbxalfUTFDctHdvBo
q4sqOxBnP+7ormFeTXlZIywVYpQyYmKh0frfsDV6lZJ1i+pMtGQo0XoDblVQs5gw
EUw3E8kvmyAZv6wE1J2fbcRH/rROKajPmBA1Zaf7m05ylMDVh8TM9iFqG4FqvWhx
9o7tezFvgT852+eIwbc+/+hof7JKlVd8oqffbbS81gAIJB1s72AVzK/dBOeOiRiO
Hy0gceAQYMPIWw/hxAHJ36qs/WCAu1Q50hH1WYvmDwe/w0LtFFVyWrNfjxGDhE1j
SntWb0bZ5JEAxbNoh3O0m/SKUts8Uuve/0EkbY6EBB5VsupAMlvo1lk9Fqrg06x7
WzRNIzHt+H6at8oHzm8oxQWlJzhy+X0+WVbhBKBDm5FsIcGYw9UkD+YDZuPj/D1W
5SrEqSSuszGO1gTb2VPIfZ7IYcGLsTDpm4k4PvaHzB6cWS4l3bg+5u5RmVkkf5Rh
V3RXGiQ/l3RIDThXL6ECci8Ulqb1L45OvP8n3EMox7HjzoJa0ihaUcaRuzeJuM9N
bLsEgJF56DodK9yjXdH9wM3OdGuVlnK0EX0182Og6GXcu/UVUKP+GTceerXN0QSD
uI49Y4Y/C6ndUQmq1HmQkb7wHwDiJgdmonbCdE2IkgHeAodAII3IroV4TePuP3ql
xChDCj4aIP7ApVufey26WvH+9agcokcNhuQToZw0F/p5mkZtWUTiSEbHWAYdEVyH
hQPDRyqvz+g6JRwp4aQTU4RMduNnO3JtX6xKXjDlEAPy7RteZM2FJFCWFHh5ca6m
oetEv02dMWFE/nECdap1GvNDKvTiv5IjncPlmtjdfF1ikbpaylaX+z4EfkPFdbLF
btmqbXIIfxxkMuKFojznOcnfOBZj6G7wyiqws496lTWD7mt+V+4uAGUW1rU2yZJP
6CO7Mwn1c+uZV53Z1EPFqAHYQIeMHhsVZJAaEVAE7gBcAv9YHVnSpfMHpKZFg9vY
e8AfLfNQfVqc5RONc9CijLlrBHkDOffid4nn0/Cavv42k/7BG26nxSRdgP+NH2YJ
EkldJn5XM+3r5TkL4RKM1FqDw+gxCzI7apSTLm+QAMkjwGKzyqQkIU2nOmP1f9YF
nlaZvNKRvO/5xF8sxe4B+RpjfDY6O308yP6SoZrb4rFgL84+xwELNARuECA60/m+
GiRysB6lCCUV9yMrEHEhTjovu8KNPXphHkAPYeD0oozbkgocQlDe4uPSFkd3gTsu
/JOiOw1nOq0Fy0SuZfZCjvDWTwqRiQ4/Rzx4rojdIzgPhoo5ckvBARISo6Cwx8xa
BlIfX2xYXCste1Z0ygzXCEf6aPfJgp4pvrpseL9woHlt3PRnD7sqWkuenLNYCjo7
VvSR+yh58PHwL6+i3AFdpXvXkRuIGqN4tyjJEUUR2zUU0F/4X8SKL2mzpLnNcpwL
T3/bascG/AXQctR3RjHUaSKYV8dsMda2w+TJZxSzORdnJpduGyAFND5o9gFBH6cx
KDOl2enzytV/NjKQd6AwFXPbZZ1MiRpfCIEpm1CmtIeGkEhq+FWmNQUgAhOVBXmE
PSTsgKHTsypDe369p0EvhKh8arOzCyhCHFUOcikq/Nxz1RcQns+eXkVSqUoAWWOZ
SaK2D2Dt3XKE8GXXcPfuWdvyJJIFokd2Z+PLsMVLGc3Z/mlPu8guUNPtdSELyKIh
eHxB+knT5CwdsLbluN3jIGZQTsl81zAkkF7/dJZUc865OsiVtsksB4sdcs2vf6B7
MFdYzXk5vIhpEroSqCm1dB5z4LvQcngnid7XZFEEXFrFZ8XMKsBod5yMgxgy+UMe
2iN20uScWetwA/EaSwrUFnge7mRfrsdrEyRT6HaSmpAT3AmAyKYutYj+yXjMOEof
pae29R6OfIxCikXHEZDhJbpmJJWAjKYNp5piZDikMB4ScYE91967s4mFVEh6lnEh
Zvbu7rMRKTaQT9ZViMgEtdtTzG+1MhuscFR7gxXwiR/uD3Y2VALDRSyiOtFf7S1r
49WWmbujZKh9hty3ORb1Q+bWWiZptoQ5XCE3JKmRPu3UmFP5ar9XwfT7Uz0HABvZ
5FhOvvLVubaToUZ8zTG5XuyHEbQ4zJRlbSHPGR0xvsU8vFOoMr8CXYneCRxp5Cea
l8qqelXlCbzkHhrypjWiNbtA74QJD+80DB6abzpVpotXRikVdUwGikApf65DitI+
dRyiA3u08Mo2N/syIzYbSGXrF6IbJ6TvXh/gQ7kpbkC6t7W8E+jaE+55BJfCPYf7
coBUiKzpJ10QYa9E4g5T/FXz0UUT5V4cn+3tU+cXcCNgIa7cqZbGmneQxrMUHO3I
cG+sR/1AXDtmnaHR4hNiFSAQ7SJNweskjoAECaR0xzuvXFXnOO/vaSLbT1I473Ns
G20FlSbVDwtwMVHnMf0y5z5/4mfRu8IDIo+efuq1MkU+pRg+2k/Wk+qQzRoJg2ts
znvMoK9tggmCZhN8L4ZrqIIEFJR6hH2t7D8BhNnEyNLnIc8sTpqfl5wRIcdvCdCY
JeBHn474Mpj1CXU1kpStoiuVLaS6STfV+m/GQvUeQwrSmIAdSBveH7XDknoIxXic
nYTdYI2YoF6NgEZiQ3OTvzYKiRnq/NRyMNJMxyfAu9hlBGhGdFo0lwdNBIeOxsYR
0r6QB6CmgkfcDjcFUztusqnhe1wor+dj6n2dZs8qU4DDSPyxApiF7c4q9dSyoi9C
EIGFSH2vaJ7eU70+ySMYTsuFybXA+sdokwMCcFF/Ro82xHvIXqrOusbBw9ce7Oc5
oZd5Y9H3a7LG3hkyOcNrvKK9Iofh6adL5fu9gk7I5Y3bwA0aungYjiMJRfcQk/Q0
DF86WXbIzojHT+EkMB41vt3cq/qpu/yPRXOb7uVLdfB7UaIBNljKSo9FW72MMWOW
HawT9nH9Ec2oMD5tPZFHMbrEMzGQYUHdWSCJlNGkdswaNczOrx4bCowOc8TKq003
ijS0RXGobnD9BIAkuam7AOlAWHiv60mIlxLIUeFTUwlCcr0+/gJB2Q4V0wS9bwxj
ld3SXlV5JhVFIsdcim/tiFOuFo6VDPbIn1xpEdlDtrb2pp5qqS+Hc8P+W4FdMIwm
076v4UcLfC4aSLgovCXmyWhr2FZkOKAdts+M+TTRExe94pqq+TLKcTeimXwLBns7
8m5GjV2klgGCe1U3DZJMfYqZBA7kvCU+0fB1fTQa4F+qtFckvBQ8AKkNZiM2Hu5v
or7oFLxjIzMmajh5o6OfF3dZovydC+mMxJwdyrGFsZVOIBuoTP9Mx9ro2u8vH+kV
cm0nf8HwkZc1mK6bcY2UO0l+tduzKF12Y0VmAMk+9/pK6KR2rrKyB/kZ8HBB3Roq
ieHZRCM4Lvw+V231noCM9E9DLCwpr9SQSYLACOcbnlmgBAD2JobOauheE70I4As/
N3Cc/wS26RvJxIqEQ3KlltEepmJztqD9mibb9U9F1Q60rMcVkDbUtSC01idZAMGX
ZnAIUqhIFpaPji1zwxxOac0kLZzbUENxCdDWvvRIVmYARbuY1ENVbbDYTs4N+bJX
eBZUFYpJLrcqMckr7iiKbdU6LQIGkVZS1XapgBHEdIw9+dJmCOU1NN2H3CG4dTZw
YOC689NVZNqZlfQfatVWFxHyJ8x00nrR/LZE3Uc1hQ+9sv2iBny6igahj17NxEjr
qWyzgDm1ZLj034NnD7m/zYH1jOp/Ft395SpIsAysxPNCvC48ZIwhK5Bl2R8w4He2
CBl017tt6Yhmgwznnp8sbXhRdfwNfPujODgSCXgzY08sqBUn4og3xSxPjMPR/qdA
4IqKReaNkWaXlIrrem2be9CvAN15mfeXCgnj749qr5neOuGMTjl4nkHDe2W81fX4
VuXeuWmHsNTsYmwvgyeljcQMluhquZ+egZeTRDEXZBZQDH1k4idpDJkghO8tTRRB
JrO5T9i7RFWuQ3IiuzzsFrzDM6IFEEHcUJ9jWrRPYzNfq9s1m6S28B9atdPQFWs4
vI7WJsrUIpPtpnQ3r2GCdLStcOoxA7mT+DrqEK7LERTNruxBrQcftHfs7TrFQYoK
Z+to6abnrdhz2oFihSvAFDuafju1KjJ33xl35GAp1jzcVMUrmzSXg3JvZbfvWGIZ
KTRwV297AZjV7VQhUvooVaiQWOHT4HUFE1wp/J3ccwKle+1IAnhrJxDqV+/Sh2NM
lypZoqc0xbV5oK2+aZ6jMv9JBLufrdK0wx1iF01U6xW15frJ718ai773233KWBKX
qChccYIf6vIDVv2pWL4blpF53e5PeGv/kiHedfKt5bhY26MduZ0vW+MCbUtOk/sh
JpbjqqASVtcV0JJmD8ApysHwr+07mjGUPLhx4r7ocbEBgbGP4+GXY+0rtVFmJuU5
s5OLeTwbueocwvkQfmA6a+tqElEA82Q99ZYxLFP0btyYLo7MpQbzyyt2flVhwU11
vZodQXCdQFE7T2uHn8bImro2kW/gGCERwJI4L1Km0h2fV+H8WlwitQS9kwvoNwZA
1j0klBzbtPBUqvc5SUZEnBvITzrH6/mUFlG7HF4owrVHkl1V5akqmW/iSafMJ5Jz
CQvzBMeLqrK/FquWX2XvJY3PwCPUSpAnFWIIo/BBiPfywBSMmh/9n/tUDjK8oE8W
6S/DfUw+qQgDwQDzvSDs1J8c2VuvAQj5O1SvPmXmtsOwqmkq/cAaJtSxwRudGOKX
hKpwjPmP2UxfSqSQGuU79qFkU6eUBr/k1YWi1VljjOeI8WkSZ3e2Dk7fOrwZywEL
6jKx5+r/5D2ig49KFIlDy0fExFF9IZIo5vWEvZXn1TjcL4zvz20Rc9elqAQlBOTc
qi18UntwdriHl+yhz5TlltI61tjoDAnwP/FtGVutkgH9CWOYOeDG18qgb3EQeAmn
o76Q+GKgDTOnTLrRyTpGKlOJOrrNq2Y1iILhFBLiB/Xy3qe6jFYWdk4QVnDeUyE8
+r4Udp3vTE0rNRpu1JhZLr4irSGKwFCwwyj+aMCJjSPfUUUWIHu1KWRoiH1fTxr3
Tj0jI3ebzk2BU5oGKldiYCnlnWyyNzNn2FOVXwm7PFD7iXi7iESPIWNbSKSU4unL
STOTEkWRqskddUVbujAt5ZavqZgYqmfA4n45+pw1+xy4rhywD3JFuhFOyAZ6QAiw
Yl9n2nqGSD2T3bct2FfaRU4xVN3UrYhzuMubBIsB4jJSyBWz2Nm1ZCyZJNhdeh4Z
q/rLKKmS14CYiPiUlGwFjOt+dC/QaKZd5J1HVImZPl7k7BDwYG5jotMwWnDx8f3Y
Q1KhLuauWKL3YFvn4iixzSd9RL4FcOGa68FfPeBNHL3Y5CBNsDMvlJ+P4y2oRaLc
JWu3wlWPgUwlFOceR2XM3EOeqUbaY5tqIKmLv3SCCpDafvY1Bzre1V8RM5GSycNs
kDzBAPsUSxEVgeSkQusnB0hKkTAaZAV+bdQcuBEwKFlBzGKi0Ti5NPqltRCSkim0
76pf17tkh92jiqLVDamfxOf86DH1uEhdb5375xdOn3j2PEUT9cCpVD8ax+vT6TDN
rgBXxHFG6GwVrP8hV6gCjpoZirkEIJxl6vrrIhNk1yCN3y0xE1Smluc5OOmMA8GN
BB/LQGn1ULF4NhTi7SGYcZ/FDQhyBkJpGnNjX4LnfNiW6NBMkSnh54U0ZO6nklNm
7FW64mS7RkvS+q8Wxo3UxBNXCt77tWLB6bRHHcp2XXaaFeWs9qJAKx9saaO3KL5n
HVujtu5ExzdqRqchHAAqhN/xKYQP6O3m8fCmgME5EFsusL8J2zSxv5UDQldzN7hd
aRP72bz0nVqFhcpBmteqz52mCwWD0nlKSqEYOUNpI0w5F/vk61VoZayurhGN7moV
5KVFjPzeph9YSrlOu8JJeD5mghU+Fq8sD1WxpO5I/96RazMhlDIikuacHGGXy8cf
6CTr3FCnPOk5FNdue4+xtadWZ3RDGwieatlWGUwMPieSDma/7W7fAYruO5iZeE6P
Rt77FK3ARZHUZx80TeXYDrXLxb5WM2tID47UYpRxUNPDiuTHtNJNORhxKF2okn8h
Oyxj0+sF1+6smTm9WiNefsimdqUIjdo7TXB8SE7aqmQX68qKiAtnHKVtl9OYU3te
WxSmViI9HdJAnzQ7+LUA4WZpsSqnphn9ud1BbN+1d3IyvU1yI05oCz4rKG0eki5x
wuhq06enZA+ApDaLylwpyaSDthjGniS0nYw/CwbfjV5THU3X+j+MAFr+iWxrRk9d
ZJQVW0Duula198X3R+DssQajrRw9KFjg1BWS6y+EjMcQjE/vFQ56PZDu+9nS9V5j
sOd2MTUjxpbIT4DHfL14RzK1MuHSaqYHz+ej6SoMNJld3H7r78mswfboiVVLjEeH
Ptyg1ErlI9l6zVkg5oNf06xzejpZHiO9UI5lzfCLAxUXe8d7JpyW5oOuK7U4iMrG
1pudHUanrMVRKkEbSLeTatMI925AjExRjolWtnSINabDAXrhv+tRxWk3FvN9moG1
e0rOjX1wjm0ueO+3ARw9OX5VH/RsnPsGaAwM8QMlhLX5Zk/nPtBdLloAcRq+pq6r
kxrgcte2dvhh2zDzdOUFEsQ52vIvc9/ltUrgKEzk6lR6VxztS8o2lHp3lYgoe1wm
09toyT7mIHGFlGqpJkNc3FgyDK5QIH7Cmko2KDMdgf/y5kC9WLdTGaJt3+avr03r
6Y82/Vr1Kf7UOUQhGdxmWFcVpH67LYDDhv9ibgcEZA9HFwCr8EdsW1w4ra85i0WN
LIWf98j730cOUYUqwy0n5WMQ5RTyf5Fx8Nh4iQPS+ClgX+zZ0nenbUP+Ce5Kbv/r
LCTMSeLDrcXGBHfQMpxZFd1KOhKJaxEpdSw6t1qaPlyZLxJ8fxtNq0dusAhu6Mdn
NCioSAAPZ+Wtk3sNG3MTjLzH9cRcOiIqiv461HMGIGq2W1nBcg2IsI4w9MoibdRc
fcMGOvO1MdbsPxeUH9npwYOIKvUE0jOVV7CY9uniyjl4xIha7smz4zGQFxJkDmaJ
m4slHxIpT9sKTPhAgLf3+CbSYb7Ko92TYj9OwisU961i9wHl+QAcbPyrYYRT43eg
E8172p/lcexo7tKILvwVWxbaEk5KerwITVBOLkuH3QvKiLXi2sCG/uI+vW5/NRz3
Ma4XzyRxT/afORC7V5OmrzCGGG/MhhFFKV+H0uyNX7jXa5LMd3VuUrXAb6l7xJdn
9+srF0xh0lC2OdDv6AOhnOIAgauhsqfXbzvBNiCbQQlyINUYgjonvTPXJaXXdMfH
pb680ZhMo71vLs8oAohmOqiTzAEXtC9E7rzVBw/r8JJGau6EdSuGnIJj6/J2aXni
6yV1WTtTerde1FpGp2v7GtTTyUTrwVPj9njo7HJqxZeUnuT0Er/vbe5k3wpTNun6
8qMb6ceRxRswughSJcRYMUhpZaLTRRXYVCPWzSv/kYGBuBqJtYxPkGapQ5L8Gb8s
4xVXbE4dxts+Nc+PxVap4doZPc22q4C65UhibSWE6xhqGaR4nQicWSSUU/BUNsZa
/5oXhvdp8uMd+5hvrpjIQodsvUT9XKnWn08egU7PVQlmywND2LDAvwtF6BzPcV0Z
FqjvGdNSidGrxFENKQOA0WYO0eoUSNudAN/9IK8jGgnMepBq2SsQaz/QtrTgW+iP
9/EaM47Wkt5H7BeWQgzRegRkIIAal9BafyR30XAnAE5jgnOZh5T5fHnQFIJMI1f/
vV894u0lP5Y4y3xTEtbbaedRI3+0VbWnQhd2wG14f2nGUE27/oo9AJ4WjbklJiKL
PLpHTCdjSkhGQ1ycjBrIk9B/7y0P6HzNMpAJRv7IC/0Df1tl/zk5Wtaa997djMcl
l5S+z7hJB7X0TQnByOCZO34huYoQHseNPCT0YVd8/OsInky3/08wnutoOzoNCSjc
2bgApEB/QZs4uJL1zDhNzmXJp0JVJsXjZlVFBCtwMAtdwd3tHBRdJisasSvRVIQL
SI1Xy6baUSJc6q/QUJbECrAyfNhYFMYBoIob66DHlp6Yo5zHnAIcGQduhqMm/cfl
VuD+dariaKfHqXDhVRcpbRhxQzRpoP9KPhTY/yp7FIC9cGjRChvrjvfqrJYqAVP6
B/a62zOGaNM1AEQ3u49uvd9Ze6B8hPmIOQvTppXMwZvubj3BkjYyZ65XwzDLbOcP
Hs1bB4iclhyfuytwv78aRQV/XNxtggiia2B6/d8DjeKDkt+rFhmlbXz+waxubZaC
xfrjQDoeIyw/GqB85O3Szrgys9v9QsyHszZFBK3x6BCRpdO+pBSxKOE5Dlp3Ey0F
1/YtpdZTnH+r+dw7o0k6uYSiUCgHC5aM3a1QL3hsYlQKzuVEZx/P6rqDaIpREuf4
gjdAt0Hu+CE5qscZ2qK8q3+cmPw40ni50JQTUUS96ySBxUE7KhMQSWRMEf/TtcPF
UuH7Ik7k2z4yiEKLP7KtOPT4kHr6DhhySwXw936ncLkV7/Z2pY3aQn4retousw0e
aoBG4siKOpq7//hNqfpVmUpOBPsJ8whKBcdLZJSiO2b+bRJvkw8QGFfc3W1zSBll
hDTJqcbBqWIcNG4fXQ8thmxUxRiM4tUHLrW92+Za1u51S91hDNzIwrg58YKKU2jt
xAnJI+YpPEoe0HdB8NPzGVMFqr07bFKR7N4fMTBK8WL5W8l2jm8CK3TOe7rlegaY
E3088KM3obD2m9Abw6P3745d0zz4hoYSnkntAI9FEKkJOgJkaI5PhC42ItJFs70j
AYekvtFFQLhR+Yb4e6P4g/INWURIZmZJIWM6syOPZSDyrr1hkpXCkxcqjnFr9KLu
2WeUVK+CVbcpcqiGPOdBhdfSsYunyD2GTz+2XNhyowRgR6Kpard8Qnr72EQ1JKg2
+ecneuV285W7xVItqVtX32S9Lzy1IJnuUOkrjEk5qxnOGqYuCdWvNvPn46nSHdK8
QqGzloVOmVZRfQtAksRP5g56rGgi9fxaDzbDSQHkrP+vbCaiwaYwVvbB+kAUpbt/
e65U7WnedIIw8mFub+pcv518KTa16qe76kPlMK+tnb0gIVokcjKFPkH2tv+Y6H5h
SdM8y/Zc0EhF+dB0Q4Z73bd0Ka7TuPTBmCNHMJq3QZzjRmkR1C6t491ZPdcvtzQD
Tn3H+q8N/GWB/R4Rn8qPl0SApMhgSK5d3llLEm26DT50/IN+Hi6ragE9mwSA8wKk
oxwNA4Bzdrs0XpOYyTu2GNIMse8/sttbvyKipgbfEAtzW3OmTDqFqwEXhxcK4Bk2
afF4ymgq2WAEuJChMiJFcmTe0KALkJ3jeTbTdD/eDLvq4T42M5d+G2Y2ly1mvnhr
AfpxI7V1RTWJhATlZP3oErRZCfOJIXXWIWty/VK2zZNGhaxU5ha16N2qsbY9s5FB
qSyVn1k0H4CR2UUJK2zgmgj5kdj5I2BkvoERXlKpt28TMj3y9u1Pvg/MVrX4fw92
2oksIYXjSM3k/SaLVqpUyGYxphy4DUlyOxyhf76DiGzm5ED0IyWfIBClml41ti+J
vxgRSlRqayeN7IL1LwXH5oOzPKTyd1cfuiyuWtv/kZBv61/ShTRe2ynk5Tyco2c1
dCWfZyyihDFKM2eg+NPSO08hgQSnY24N+tLO2D4/aGlvUGkJAFV3KL1X4BqIVjgS
Fg6mhcdbJf8oM46St++ZE/ETabxT9g4RMlgihHQI5iNEFBIDxrsy9JI83NO1+i6X
lHWfpTv0dfONcyelNQz4Qo4MFETX6hUi+fMF69f0SjRUsJmftHi1FgEjky2HgrYQ
GpQe3l423gOMZDhxC6veb930FjikCELN9GnaqKnpSxooE8YoAiUxVAt36cY/Q/Ad
vT3BbHBIOi4EHJUjesiaDaFJIUcwTFoWggqZBPNdwjRF0vGA3MAmrfycMeRqlTqf
j+JWBLYABOU3a8rbSFWhUSI7Sj4EPnbkdVDmpGSpskyg34RM6zwMWJUry2ksmxSs
FD8PI2VmzdNfwQCxizBNH/6Ek5KOyxVOgS8/gLDjfDGI9rpk2iT7nsqrQOvxL+f8
SrmclE+Sd81Z/Ft942f34evJDDWKk8qYUEEDLORogkLBumLeLztB+pgrwjnaTAhZ
pL82ofHbhThaSWcJMisQYApinVSjtoyb2plrUBZn54mXPcm8rgUMrYaJHD9LUCMu
nFImlXZ+OQx5ldpUJoUo+9hETu3xkcKtuqUVSVBMjvMcDRLgqeWZmLp/dDwOtHQ4
93oU22FT5gZmk/9Y2mO0gHxkxNRHxPofvnjaIdD90oFe8SNQjUxI9o61i0ofzPye
hwBM9kx5li+bWF/+ahWm5540gHuPxiRqegGwcmNA2l2r8mM4GHyASUeQ9B4snCgv
/1gYVnzdWx1Lq7iFc9G27choTvN19n/Phf0JT2iP/Hy79dP3pdcWrSyVBOPGgiSU
Bu50Fn1sZ9KfhojrJ/BzlUx3YXtcioJY3R95mqXm1T12TqCABbqGukY/+M1QJi+6
Y2Rf0Gm/iotEuNAyr9qsEp63jlc9SXjSxgoMtUdGhWczhywDDJFKFqbyqMbM4tTk
vMYvtx+qEU86cMViZpbVn+56U7L9b7GpSTtovpbPEgtmQ79Dr15ecjD9fKtBF7PZ
wS2efsyugaVWhaOk5nLE22wZa0PiHS/EXauxIynU1NOzRy9mW/QGMY9FV850m7Ug
WhiWJtt6sjB2SmMt/7Gdujem6/XXX30YldljpFHnEzHGOtFMQzcJslbpUc0X9WNF
e8LpkCpkDbQthQEvS5XM9L8mtEiTs68xsw1sZ+WKruknJh17KOR6FTKXNpagSNfZ
AUA4xzZHo9cs3o9jux60ahTT3G35sZFeJNJzWzvICR2oJVNw53bBmNW/amsBVqLL
eIn7JloEU4NXWAK0+JdLCIBVSR+Ao9GqiE2se7akkgMK3JwupsJcFxPtGzb7OUkq
aNYKCNCPQQsogO9NAP1n81EIFo1KRULRjdi/fWi1On+sqFTVDX8z1BpDR61mYhty
ekOl2iYn4VpIogIp/rqjU0nBm0U39nvZgcddCwMF9IzKP9as6QCwiu3Ya7TbZ/qK
U87IGDYqjvDLC1PTFotWbvoc1PH4HLc3ZbAGyfCcKtkKhUKqdXEzta1UMqHKwsx1
SIzUlO+Z8kf7yraCiAkchmEwrMj2FKSjmyrWzlTG/ubY9KQEq9sSDlOtKQrv3S9g
/Vgje9IrHcXlA0m1UJAKS3+oyAtwUILvbiyoQ/TUFINERDwotthLdiFcZTT6o3Ee
Z49jCwku4kawt/addEMSdNmp35tMhbdPQ6QVwgfeIFjZPDin+7Kk4E/mTlQ2LWKm
uctE3oCRK6Xg85qL3bYcvrPkLKnAERhHhBl/CW2nXnAIU0dco8kbo6juJswOn8eL
li/vlcKN8SzJC8eRGfTLudBBsEzK3IAsjlgw/ZuBL5HbYw/8jGG60C35fzmuLWW7
D1w3I6TuuCl4JtugUH5si1PpgS01rln8ELPQ0OL1WnRU4NVjdEPu9W5OMOEuriO7
NCMsOIhhzJEYj25sawg5dwgBSoscTyj9hL7LU9JEwe/SkozTRTmjoAROupRhOcMN
lXVq3k2KG9KD6/DwqAozylJmBCzg7yGfO/TjODzJZxjpadSaclyR8TCqQprD0uzG
wZtch+vMjMInyOUjKz2/ZBFwsncGG7aGbB4xxLmprB0GMKK7LoWcJHOVRRB8RWxe
R5qOllkjSKCwecwrCwMcMWv8UmlmJ0cC6sOBqpYOIA94ZruWJ2fwVa0S8Rv/Y/Qo
a7+qo//gSUd9OuMkpZ44TR1h4HimdS4KsoUynXgO6q0aYtLEkZWLi2U4sJmXJt9m
3uWFqBUYoldmKw56sszY0xKSjwNW9wc8mlOVg5hFTVDDvGEml5NWnFEHqmGmUK9Z
cGg/64YdgXgDAvqkNOGolKnx8sKE2xJdbnRNs3tmtAy/sgm5AR+KTEPpcrGvk4NO
TSEocKbLi70WHB8/5Jxhgdvp0MGOZqRTdW/Zo9ckE6GlQdQLcLka39NIS6JK7Lko
FHimGR+jMJBfFQY0uv5oB/vx7k7tIgU8Uzl2Gg6wEPzgL+lTfi2AKFtJcdBGNiWp
ttExeqlPU8HEy1ozwN4VR1ohxMuJIZJ79zGZ8bh/SseiUV4oRPORzJHQkbZ5yWzJ
Pam1S5SGmx1Oohnmq9qBrOyzVPldURIhOhX1fm86iuZhkBvVIZXnWaz+Vt1Fg6r1
8PGPakz+lmmE0CrHCFDCQN5J15LsmvINlBL56LnKz52xzTcecxrAX20QyChMfxjt
i2jcls91yy/o2UASZq6DIA0mPtbyiliUR3p6sC1xBqTxbx+rl2qAZ78XFtevKfe+
UpYfAEBvVACF0bI6PmgSQ0erWhKLXvFOvfrJjaT0/B3IXazx6TtbcheVYc8MYkM/
1XnEaD5vJJFdFPVJYxUkvJ53Dmpf6lt9UNv7jVduH1LpvSsaDCuTkhHjbGgaj3vr
a+4oAmce4mbYQ1Jz4LM1q3cgnL3YwF5IYlAORQ+hQkckKJ1q/C30o3tMnHsXEZX3
0q2fQfjoQnPdx2Qesi/b9/AqxwvjiOZU3sW1URvx9PMlrRvKHZ9zzt42+JlFNvan
+vWF5N6c9MiOZVL/03vk77S2e/6wt5q8SiEFOISQlcYPHuL10upsMmBPdf5yRmgh
KVRiwvRpnxRjGQ4qiS8P4lftJcpRpbCxBw5iKUIMhG6bRqpsJxE1r4ce4eyH4vkM
LtNKySpukgVfHEJ0RMekjF/tFZCaeMkrY4WX8HVL/oHbahqbW4A5D9sEd8hswPjF
6my6y+6okvDmmL5exqBwzYkp2SrVhYh8oizVH/TI00eym2ZNH8JlhyzBZ+X2ayHq
`protect END_PROTECTED
