`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zLeBvhDOiv75zFOeHwIgaladEgV+JFG/K/pjGJTgcRS/5/k19AnBiOp39uolN0Uw
79JATpd+M+QFXLdWhanh6jV46uCP9KpFDs+LnHTrxYzMMzuVVYvBNfwGHbqyuEtu
h1XVdHdXriIPQwDG4XMyox7ZvSKTvFcc33PDk6B6W4s8qSkAH7qUWHJucjvusNgh
`protect END_PROTECTED
