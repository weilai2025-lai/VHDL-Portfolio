`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5N+cMXdUZ0hUnCYQrfiafRn/l40sX2UvTdh8Q0WlVyLsjtea1Mp3DPQAbO1WZGh
7WDPgEpjzwaxOrNKAPn0A86L81eTEtMlUtsOdadcjuIeS1M0875Ma/POvejphZDb
XL5YgA5d6L0x1kxNqP3oINhempQVWAOyxLZxnP/FrJ5Y63rIMSgkpYSagRZPVv6k
llf3gBj25xWGL54jtNrzyfCg2mLXxdTEJcF656UGhaoRoC1rPdqIBECIAQN15tF+
GwMmqPPM5/S8xiEkFOpPqGc2c6y3o+pCPuRpPgzrLZVWMGN2s3GZA/pEswi9C2B3
b2MAsakne0xL3bE4VU1EMbBycF7vSCnzZIJPy8CzQXZ1sRG02obLPh8fnl4TMvAi
9+pV5WylvbCwAVcJYxHMaQke71Yfi7H+YwnJmNJ1CKJl1JqCtPr8/R1n0CKjWKWB
I4XDa/am1I/M5P3wi3aZDukxin6xsKei1N1VnOHeLFHzsSd2wQ/fJXlP9P4aBFDo
rtcVn/Mg40HlI2M4hL4FLpB286nWBePmUc1kTdwlFm3U5Z9ALdnX0WYh95I93cjp
X5vWfezv3hWASr/86v+ozHxNVZyG59BNaDq0Qo/6sY+DAWXJ6NCNeGHv+0jbQEY5
qRFnNi5OyfSC6suP2Ged6P59K/XvPLAFpItzkIEn9+BvrC+CRP4Xu23ot4+Tr+Gn
tct2XaIQitbYKPq5Bh/v4X2DBHEteXZ1jb2AQI2GwZhaSWZkVXClWpxe4SYXDq0M
2WtLk6sz8Y0vrECDXPWoNn8wPlHSob2Xw/77yQ/7j5O4oZ33SK1ze/U4AFtHCRbR
RD0ZZn3Fnz1JtIi0qxl7NdRr0vsOnAS82dWmeX1p4gz+zNEeGQJ6hf6+mNvyX807
tANbpwfa7Byak+ut2o/R5LyDClrgElOQBBsZ3xeDfN6qAvsDQDfpaSOz6NQnjBff
`protect END_PROTECTED
