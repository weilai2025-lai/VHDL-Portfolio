`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c2yXJx5dGwwW5J/qbw41xkWtNotl0UdXbqPVVgLDJC1lQo83Mq36mszO2fW48FOO
tugORyTLW+oLo8wu5TELJFAgLeHMMaHjiMq56tCFE/Qr2RJrYeABpj8epv1+GA0Y
Od92OutCl1LsQ4cTWVjBbo0xl3BTMbWxLNlut7xbq45Z8qxs4aRtXcLhVHlbkgl4
M724Rg0rFNQ6uDV3pRzlV3KJ2v10nJwGQHLrpcnO8AqzGZRfwAZEfYXPSeynWUx+
Ci5kSlpukxgcqI0B/YZfoxpCeuLuC3lth12y0TGlb7nuzigPUxdaPA1t5mMGjbrd
DaTLrYFBWTVeJjtJK8up7U0TwmyCEsneMXWWzgtoKSuZykhP625Osr+rSGkax3IX
i1NgjQDmKBNheyXO4GLL+NQfHDoSVJdu5TmWGDpq4RekOW1dxiX4iuMu3Zil96Vj
nRaYlCwEUMATQ6iXElD/dZ1kgBN8jy+MEW9DnaQ1yGHiTXj8Ve3AQ+VFnXjAGL2Y
2n7HBUnIyWk04lqAzOEZv3OlJWqDJGwbLCfQAPiF7Tz2c2KPig5QnqJQystWmD0j
M9dqDLslgiwM0GJZHfl/9XNFMY4buh94Tm51jl6BXC0YYxhAn/6hbeNrtBuO19SE
u1PW+2LjtC2JYU7igpU3rJLVX1ONEDlqV2z34Vk4tbLgShFaeLGZe5hMA6mYkJ3E
1BhAjKCm2XoM3W9ekRaYZflnm0hPV+3nFn0L5qbUZd2HQ3uH7gsW7acDBi1AHSkd
WBSCFyAMhJhueP6g+y7ZOkHIjukqOsd+FfpPVMekrBCdQDJt3/q7rLWge/Agw+gw
1cCm7AMW3X6tPaI4eFGsaY4gUBcDlOdCdORS2g+hUQ6Trs4gmuANrRNoyWL27sw+
fSmKqcyKltLKJDsuv5eV8a4CNhbi6PpeJKguS9yOvYb4BddbcVJ3uLXjnjrKL1Za
atEyLQg6220zZqcbeMVSyVXO2w4WO1s3RlPiXYpQM92eU8uSz57cLNLJjzovXKzt
IzTpC9deOXRiAn89qhqBagTE3flAEoUu693zBcH5EiEto0WHpY5CWa3y5cQBjYzh
bd5zDMCHRjHMvJaCvQzQUEKvC2QOiGY6cBoWb0yhTD/KTApJExmJ0bO/E0G6etS7
3iZh/VCg2nQV1aIHlBIvRJLECK4O/86clbozi2Y74G9+u+jAN9SBWcXONZfV9+s5
cO/hDick9bUgzkpP8ltg29Erz431xtkwR/kbdIimOO8iklfaySm03z+20Yf8I0Ew
4v6JDyqMVh3CPwfqFVdj+upiCRDiHXxDTwUrQG8y/Cvxiaia4aCF5pD3PmkmTmmY
IKyXWNYOfgJy0uso/ob9BurHqhAtaCyYu7DbVHRtX3+Hrz3XF1ZvZ+khxP0TQUO2
cvM9bt7QDzlouMJYl4MmOW0qwBisAujs87oV5qfiP/0uvWgCn55wk6g1GK3YFv8L
iMCxUahAEGHpIuCHK6yJSF4u3RCKVa76t/SM1M+GaJEGRF8MqNiYdkjtmS8DfZ3t
7L7GjmMAj6jmFOAfjK2fCNnI0cw8Je3wjsmvbZpJ4azQkEn62LWIhNc2M0KDnEMF
XoN5H8vK1MXpizwKKbRhqzcPTXvgI3QESPrJPJD+IxMvNEoQgSoXG4JPEIFibf+V
GBzIRJ5t6tPy2IdxibWWKzIREAR3ZH1LKoFXXkeeuKU3J+NZoXu8t9I7XONiiXwY
Oplk/7zVhZ2HKp/bPZt6eBhU842Lh5Zw1+texMIClFGUsKBpE9qu+XEtOm6XZ46f
3O43qp9xI0rxTejwZuVz/xIkBcUWccTbNE+zs0BNhtrp40usR7Mw/de+/ofmgDE4
npjj0cPie9VF4rcg90VHjoMj3KXXhztz4QkZvNCAdozwZejbmWUICZnkYak5r6//
lwEB1srnjnbquHR5NGcaemqTEDJ4Hvn2bmLVptQ5bleWdWmA6Poy1ILMLwFaDeKT
9A4k0B2CSzjqMemR9gCo4ccWMRUVuKWfKf/F1euwYqRmT27Lt8ovVGhkXYXHpd91
IN/G1akCN226DSxYUITnvAzGPJwWAmDso51dPIt4/syNESZf29bumRKWYID/xTsL
va2rz8XuQXRkQnkZX1Kqb/HmpAsSvD/8ii1h14F/Xbk1NhMRHpHROLtRD5KagayS
eI8mTSHPF7Uu9LLXAfVUH5mdycMgp7T9MLvXYfgc4JWO8ATOhznfXKqXH/477CH2
FlhzHgcMsTPpUpRmAoOcIDNAzKMN08FRdtKtvipKyVYE8R2W9Y2fKFsLZqy83av5
wDYWkUZtyjJyV3svAXzOwk0iBdbMwBPBnvY4fzUdiYS85SqRO+JeUBcoQbjhucg2
dRvAdZL2fs3wt3zHLcEOWjH+lfBILZcEEKjLwduJdHKcYp/ld6zdGbkgHinec6Hg
qI0/2xftCcziIqCszFCBbmBgGw+5soyxUMtFS6BU0cLIcCgFmdGxStj6oLHOFysJ
Sy+dI+kYtjh/xNWQF64jNN8xunksKFBbHWxW1XBFXwhObW9SeX3rAGM80uVQl09v
ZuvRFdpoYyx8WAlWBWqK1YHC/MW7IDyqJ6pAF45FeaN0HP067roTZV/eqx3/u/oh
0Nw2jRtgYdI8asGzJk3zZA==
`protect END_PROTECTED
