`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dtm6rsKWb9tkzJsnwxzn3jTByvmFo1Vdw046hG7qkYTXlXBcXNbtu0wVgyoDQQus
R0Jufs0mookmkx2DOtyToB2+5yDVCPVHlZLCD6VKmDC99PVg33BQGfL9t1h5W4GY
H6M0zA5QPaNXQE5LkGOF0Q1RaunYG+CczHsxpQSoGgaOg5EErAsB2OXMuMJD3E0i
LFBXTzyiv10C91yjAkTz3RriQhH/fEIflUyVNrJnQqU4CL0UAb0wfukeOubgBcOY
NtLMvyRRVYHkB0Wy3rPwSNiBrbqUYBYkvv3nLBVSR5prhWU2PDpwvRi+i+HlcEvJ
OjMae8TqdlQxuRGItZGfcupGtvJbc8Rio6oBZxkaI7qVkgnpT6DlZ3esZSZKImkg
IEhm1wkrF08rbrj3M6sNJe82axPh+UOW6A3GCkRhrSrIJAZDASg62iUudiLIYEz1
JbPAB1aPBoDC2dU6wvJN06nj+kHAk0ddclk065rD6gSLgBsi5Wzlk6NaSywjj15B
cCYb0qd0NAoFyiE2xJn+7tzXbK3Fj1P7Xwe73PMazHCUWfImiXTdXpoM+C0yOqoj
BLeX1V3LyhqJJmjoxCvnALH0ww1P6VPtjdEiq3lt68AIxHhq4IwmO3lnSDljMnma
vjF50sdShxdYGmAHeNDT1YzHDtNw1AD5DRwxYcljP7398zaIQkg6Gohwt/AuJGTL
YW0EYYxhxR7xRP3u6KhZDm1lziqsNmFPPbOfucx487K1koVUBJkbbH0RpsmGyHAs
H+btz/Uc96+u6F+9AR+05MgjVuh5HtwNmXPxgf9JOU++r4p8VRGETB2f2u9NluVM
r22ke9ZZtdrh+y+hMHFgj1w1YsB9pRcC1WDBXIv0JWI+JA5uXmTktsW12ZeQwiDt
owkpVaAYlqzzfvbVQ04UdO8Fo+QVU6O+JYN+fvxUJSrWiovFh+s749JvVOus7lWG
684ykGc1ycII1wZjtgpyWrphXeLYAbPPRdKikeywAmfJThgAfrU8C8P3Ymzt+GrC
SJXQayRJR8HI4Vf9orge84VZ95wPc4tM860hcOhnKweL1ekIZ9Lpc+Nk4fG4e1ok
lxlOUftmDpziLyZMMJs9lSybTduk63repJA2hN1nN5uJT8rBb3WLk+VLVTCHkWxa
toPpwDRe9qZ4sEEQX8KajQ==
`protect END_PROTECTED
