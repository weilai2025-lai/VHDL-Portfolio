`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v/90vk96+cqPyRH6iVakRipgwA3U2p883h3aPrLik85X52L1+DS/6Zof1U4vGHPe
hs82XtX6PiVGsRtzYCRR0i3egufREn6IxysqKaORYQAONSBjOAQVSwYwMlG5jIJV
Ag4KYF8PBOK2jBndnBsqq2TPt0re7wFfHOT0F7/DmU3mQn3BxzgzVFWe+0SOuC4X
TW3w7udkn+i5fqc2sOpLahExM5othegfPAQAL+Eq/YCBj/yfjvS1gc2OQQZ5RiUH
Sg6yFhv5DIqZpC/nQ575h5Lp4wNCroNWGxPdouXgbH+OYO4il9m1N4woNfMAiytm
8DtUQMyLvvD3+AS4kCuWbU9zU4pytz9f6ZoEz+DgB1LWjC6JNJXFmSZrPjDNm5EE
PNJcwqYCOPCFuqHfqVsnXyaBWMwNhCWib2DDeTtEmWO7+vDNiMnxqsoYOoG6307a
U6dTmGm8WrHTZ6XPGnC9gB/dqLynct4w2kQQCX8gCOkMxkIqi6xde/wb6lsR4TYt
ehyHfq5CKajwzb/tXipZb+v2UHYHGQk65Vi0OEVfpnjB1URlZUuBxIz6xJSFtn7I
txgN8T+u1b9ZD9H/ad8E4j5ceTynkNPbXXD1GYsmVcx+DNPIl6ujbo/WvZfyZjdU
/RVeWxeE6dIOr4NzHKIWM5jMPEYMq0m/R7bWcMGA+0dN2sAkCfeLZl1ocEh9D6Wk
CpcMDpKdBi5+BZnr1sGmPBLn14y1Vxk2r7OL0OaTqL6pISiyQtLbxjOFPyzxlGJO
Qm7qJsI4nksjH5TZhoj1wAg2qrd+YKr+MyFxT45PlU3am0yg1V5LQLpLJjTkW9JR
JcGLC+WwittmXDv7GWHL1YhEASJlVqenew3q0QzSPY3xiExjdUeJlgNpj7EumMDk
27/4yyPMlE5BkIpPlRWCdSmpeQnelvi6TJvUF8vTarJrTTkk9G2WS5zUmIc6l83F
rICmN+wNK/u7bf8Q3hX5vfJgCSAcB/H35g6nV/HQSga8TuIWLJIjJskZQ+eXD60M
YlLF24RCBI0lFLkYaGq9uwyGJYffYKk2KNx6hjUflsKkhqRdd7qXuzsj+N4gyKDP
mpeEhp5mSnaO/JZPQXGTrZCEg21b+GnHSmhhvaQwhopoZbZuYQTfbjRZtYX+VpjO
vuxRH3mrlaXEISx1Ufm3kJheuhHQ8TW4eyUgPFuA0EOl7Jk9EOKQz/S+H/zqut3B
yu0vMA13540OzvWGBu/AS0aO5/udAzdyOHQAjcD0dBoUdHMlq2L+k5QHoOTHX3bd
1EFEXTj/C6K1V5+YdgoxHHI+7nomum9j9CBGEF9S2wrSytjOZGpCm3XwQo+feiHj
A4jj3kuXN0Hd8ay9aYabQJMQHrLu1Pw1NsD0TBJ24z8+itjrqQ1J6OGcxNPawvRN
kT+ApfFdNfD8S+SohP1UwQ9AlrZtzfKbev1Wc8szCgeE3PuG2z9fFR8Y36BkwZTt
PaL3+udxdVB9vgH1SZFPbBQEjktqu+iL0DJ8zzpElrG+acygEuAcdYL8dx8r0sHh
DLWWQTxDlhLgsM3cNTojT54tAg/wWnZ81lDRipnOCPAjmWOJzzhQY82uDynFlM7K
3IoX1BV+ug8slSloO10vYDwLElrzase7S2pULIfpPs0Cz3MUvzT8nmQ6j964ihBX
IBVdRDRdV67XLvdRDOuGoul4immRzLZ6XTAM4f7UnwBDyu3aUKKkDe2Gsru9WXgD
mkz63LANTC+9SASR0H5NhHMsSynGzlBJpAkw7Af0nZhtXTxVXpn9qEl0tPV6waLg
+uEISMmCFh7E3h0YDry52il4+qIDd1NhwEI0K1GF+YeChtefmdN9QUmTQNefKJPe
dQOqC2O1kVX6OD2aYDjdEfXWx4xxmqSH73pbRkvQjth1qCZAI2h74JXRluts145y
LmivfB/SH9QTSY/NlODIUQ==
`protect END_PROTECTED
