`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Zbad7++8V77u+ad4Uu5WjY8raDrhfvc9loPY+4SozolRgAwMfdRC17+cZogOCb7
VAdgu5Ckq6EuwJCZDPx45WFRuv31I4DYw/4zz2i6TjoZIN4CtBtSvqi+KV4OXgEH
3X5q+iWeeN/NQIBLMeX5YvIsZqheNeoDvuPN5IXGaXRClcuGHFTRzhqqiYHGZ/g4
IXoNcrzk5vfCb0yxcxx0UP3gV/yOxJDie4nqdI76aIvkp0MK3D2VodVB+HIw2J+O
sBbeMWvK2nQG12eKZt2CNeXY91iOKKLeFZZeUdkKzbGWwGQGzTZmbUBmqqbCQfkS
Ydd4BanbKb/yfEWWuVyIhNj8fLmHZGDTjvfmoxHk82I2SefNPPddNe95Na5bnG1p
UsY97c7vvrYMehxrqp4EQv5d+4mXzQq4rBsEouUnf/R8VDzbUr0fP+g9ylLo/Uko
INyI4J1mjVstg9CYYhuuPzfP3/3E1mn4LFVNHiTY03gAeGUsoXzD2qFntXhrd58H
QxEfivaaruXzToqoHeu9PZw2g2g3tOVPbCMdz5pMkLVbfdZrAB4aggwNS4Ci75A7
MMx85fq8uXXqcmUx0FtgF4lU3+NotCwApKqG/EjTkPm6KRfPYj34stlGpCilN8MH
vEH0T/R4ANQ1d3m/tzEX25Ah9RxX69I/0ZMNjz3wIb4Lyj58kFnDFyviyx2KJ7Eh
3PH/Yf1n1VJtjtWjORHNkakJdxb/GgpNNZdPGMbhtMM+z7Ep30KVKfnLKnLSv/gW
8xCrL45TZF39I08fUA6ykg42rMdZcfQyCfLZiyBLSfmBexozi0XVnSg7ExjdE0CB
zAgS7lSNrmRdZ/5chcBmmAg+5iR+g57Xf+GTQC4Zw9CDu391TRI2sDjRzpe/GSFu
l3XEYlXo1w8NtV2UMAZWoVivw94LmyH/1lnkKH+SqKSqp6gAL3wbVf7qlgBA+bq4
RyL86/95QscIfYAYZppl4Tw7cmEdkcSasxzLETWwhgU68GUDa+07ptaaiRhJW5WI
DySXlGTSOuK+a4puDY1ZYxDy8d9BTQ0d7kP9rM4ULLGjKAS7kU6UoP3w19ufrJiV
ssm4wITmSSLshjJZM681MANJu8K5BTRzz21YrIokwXBJ/+M0oXjzHrN6A2h/l/Ff
0hztky0bTgGuw0x1u7Nm2W2b6uymAiYdCkp3PgfNsMlcy0m3Cj4MPfz+n/hv6/Ms
E+LK8SPzCsS4FYV+kBPJAfcupZT046S7UACd4PWta5Xp+3B4uAxD+3DyZhhhf44R
iibWsUlQ7wUoCbByBxqjpk3SjOrpeRGqln8CFSU3UrZSUgkiXtW1dpvhHFhoVnrC
3IjPFak8EMEPr2xw0qAtdY1AzxABEke6l1SjQQUYmn+jEPj0EKqLXGy1QNdsu9pj
MObnEDjZY0XR6TMZZg7SwKZfec93Z0hgMSFwLG7KRBnYNGyqxKmFfHY82GP4L0Y5
qv4iXhHLKCna+gLYL14sA/WdJaer22StnTBRbf1hgEfROOiZHvzuvwqgbwzPlRMw
YgCT7oy8PzWnL6vGLGNw/IKS8a5Whz8CDj6QcxYqC/X24i3zabUIALPGdAcghOrO
NnRN9iZ7d129YJ18+cefo/hwpCT/2laDN7wyMUk3eG9XNWhDlaTSFWdf3u+Oosrv
Ozigdbc4IBDE0RTIeueZdzOpZ7yEvqjQHOHEkq8yJtroyHXzC63uEcilHwAyFn78
4BCdp2fmAVth5mZ5h6+LodM7FcDUT0WOYbvosFIH7HlcLBJS1NZ7gvWZqkEifMFV
Y2S3qh8M4cWZySrM+/vieDwnFYoLCKFuacfm2d9xzvVfHymWYEddwayG9Qh/MDHd
vfnhAsmwCdb8730G2JvccTt/Z4IrPxfs2KesHmRYIaPxxjjPnyfFoBX0PSpOTF9B
yaMR9sWpin8VETc/oPDg7Gigkr5tJYQTPoLU+Vp4GVhLsQqIJ8ZJ3u84qa1qfhhw
ENhD92MVPDjjTCYrvwQYLfpVSImpzK2pmX4qUbuJ23Q2YwIRFdbnRr0FbLlEtMIf
dsFq1UurrY1FC69OcB6pxZS4C62PS4meAuongg2+B194ZcIMCJ7XIusBhTLsBX7b
zMO5pyZ1CRdLx/+lJNqEce3tOBRmnYIMCquNgymkyaRE45Swpj/Gdu/cP7+KKVvo
DXWTOkXBJd0JKY5F0IVeODRe7zT4QyN3BdqkQlUIVROrvxNjTTTds42hEK4rCLqz
YZQpBM5XebkHAZnNPDl+6Wq+3Ey74Quo6Z2ATRDCEuh+dxdWZn32jJzKvoXTD+pQ
h7fezsEM3ytY2KwMDbHeH/QaLfKqIN1Qgv/rHeU2nFugrl13k1NXxk/H0Detxw03
nRToSbt7gQ5ORC7+5Px3NCxEEi9Br2QzDa6+KxyDiAl+KkyUq2OoL4tfehKyAQaw
HuCj75H36o0d+AtmwyAxNQq0Kc8WKrVJctDqm7wwEbxMXosEZ4r+OFMiEsNr7Ig6
1KCiV0f/HlHTTggREiV8kGm/aad+rnK9NSjZRzOV8c1zG1N+pfS0t6k2SkXslYB5
ew5HUft36xYGoei1QKKbbe2uTdT1XMj6/bUDYURCgqKzIviDnEII2/YX3ykgCN2r
/XYodQwT7TR3HjlIF7ZI1SR/elGVEYFXA4DuFtCuhprlcX1XEf9n4bNskcl8OpI2
+w9om0WNS/g6rmqYAwKwTua+9sh7Ov1A+c0D11E78D9DgY9Sr7iF6jBsKufqiLGk
hyXiHaTWAtV5mh4uoS3TG6gADg7ZcG/CA3g05oOzbQJbVgeBMmDePWb+4OkS8b3X
Pxjc0ZrCZEdaIKft5BopbJK4jY23Mjm5XmIfqvjuje/rNQEjB2UCfGumWqf4znm1
SRvJ2yE8DE/oQ5usmmATxEuX/jK81+eXaSCTv3aH5KLKIRKFP++OUdgP36QwEJ3X
DfIgtL/Oh2wPTmjm6f5yllR71vXPGnnnDEqxvRaAVzyajw6bLze7N0cTr6/hTe4S
AcpA780cr/CANuSGIfKIla2J5o+H8O/q/pxK4wtAhv9ItR766PUcZZAWzTBzO45F
9dhVxi3VSM3qYKkxxhArVfse6Wa8140+2P6u41Uvb0hjmgQKmdGabhAUmE7mbr1n
Af8t5//5Fttc6+FJ7nifrAJ/F8BLecfJYyMymOipEKyD8FFzdwyyo9jybLkfT4ec
0qW4itIxTOuJiD/HL/RYfhIAjQprsLJzWDvKNKel6n/mv7ym1gXZTefuv5jQQGnZ
0MCO3HTBxh+NJkv/FngeHQi6B0pe3ZNCNAsd9Rjo7eLykuGAODKlLMPKy7HrJ6ak
xKoHhdCjU7LcHvhdhWsA7z7UTs9xSeHHXnlOdWo2la8o/USCI3BHnYOtLcT8BVkY
fMZh79361ly0tt0VIA+/Z8P1684OeYtrlgCekciUXcZTOYnSm7GagX/+DJsPfY8o
I6u8rIyHBqUWQCWixmVsV+aHa9W6lX566vERYJniTdew/FOOPb5Tfq7+EoT5Ze1y
Bm+6vbg67SuFL2uMBt/5AzYE1ne2GqiFctawBrjg5qeOOMsCq+ePYDNjl2rtisu6
F2AbF9okL0My0w6kiPdivI/Xd7vmVJJ9B+/cy+Ja2D1bx95tL5PAN5bX6DwqjwAc
Z/UYK1/BYDXNqeF4CDBg9wCS3Qsv50O0p0X+iV3NlZ2RKfRGvIn7vd+Atxhn+IMc
PceIUYoiZKz6R1tpOTme9eH5FmTx4qnf+4KoXyTaUtpYgwBkw1HuK7d3e1ePg6Hk
qtGJ9stwL2MQH7v5X6I6x8sbQUkpjjDnaeFa6HfjYJUj+KzripWzJJTNnqd9JqPI
bOsz4z254n2bHWzKzCiMSlhit0zQyEuyjhsd1DEq041ut9d1JTNH5PTAXjsYk9Nq
zROSPJam1pa0rj5xbQO+6nBk/JeReYlzncHgpHpJpFWpyrLGYMOGl+qg9DULTKuN
FRhDT2VB8M65qzVIYriLtvDq4VmcqUmSFfxZXkJEKTr9bHd2nF97OCCh8wOe6tn6
/dBq31TBm7BeCHu+VFT3zzwpfhtYHZSk9S1DbjuSy71j31/rY0Cf6wsIEIPZRDw4
kb7lStz5am3fdY7ct/DuVOYXYLlxRKBmQ+K+6V3rRAcImeD5HijLtXLhA2uXmAX7
pyiWgUJ8lvE84fSXVCNLf5I0QqCxD/MdBd7sR+w2jRwrKt3XETT6gfBG4TnGYBeJ
gD0MPrp74ZKRLw5v16ipECyaFuxUNFh21ke0ucfjHE9uyE/7w1wZWibT3I7YnLJf
RSDkrrTbnksKVYOrUV+69jj8zYX8NEvktudOxmUFUffpcQku/5EijGcqFZ+jn15e
MpzagW3/9wlkZc7fpFVMzJR4dbgq+hS4fOHdrBKrtX4MjIVMB+jUC51BxxQZ7LH8
DXTtrIUSamwsISJtITTYtzgmjkS2tIZ0s3etiKioD8NmXp6WmdociJ/8cpKv0eib
nmPECTT5MOXTDxQXGM7A7oRSHJDnbCJ0r4CNKd3e1dGSHQevvCNIplFRpDURBQya
nja78DJBFPHdmlWmb7YoZd084oIbfODF/IOq/GWscNOuM71JAI8yUQsGf7pjDXgM
KYnPVLdYtj8kMVmLFhCTqnAVsD/bVHwj+/hBSbJZsmiur/5LAcFC/0XP37K394Rz
ZD95aYoUXmhqyFQJZz6At0HtFg66bwrdwPOl7IpF0aHH98qjRvI1gc/VYBNpDG5B
LPSC/Pj18HKgclWfU6d4Uo9omO+JImcfHPYqppM72UibpzCWwPjiKghuKEzkxLsj
6bCry4SpnPPQAU+2D1Of3WfZvTuVp/lxeujuQJGuoZfYrdO9SjdeO94n4hZBCGKj
em7y/7eBoRF15pZdQGry4m53QwbLUIhcfGRv3GsUG5C0PgGHbX0kOSGsYTDdTx24
Fb92JnCtiZLIqGvA8OBMalv8pkZMgMhVgxXDl/v+lLX3ludRZwz0OjqPcTp/h+Dq
7rKUt2MlUqTJMyzTtbXza9KwB2BRfG4d6UX00HGsIsyWb1RCRie14qzUIEUR2LH/
keaQOOdsby+HqcwVa6ILYVGKDLfPlzT83N/O/yzWRRuqn9bhvGvTccW20jObsGKw
Bu1BSpaQOGWhd+92RHiUTlPLEoFGdmZDCrFEi7FbQUIT2IYOb/V00Tr8wd96B34J
dmQocf886hxh627LYBN6ywGPHqzh6DVS9WnxEI1P97u/fm606HjkMeFWgweOReV2
0D4Aqww9wW9XHxq5EWo//A==
`protect END_PROTECTED
