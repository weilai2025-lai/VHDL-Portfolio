`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NMtljTS0t8kMkR5HvOiC+3Ac1BNFWGpQRCm1JvE85ncdzhTOBBhO4s+jtg5rD13I
rX1Jf+rW17obhH4LPCZFrlLpeIqJucA/DqhoONWxiAVBZWaLqNHa/YMkufXGFUuG
izUOIf0yhZ1yjj3LiZOJm4S82VjThQlh2T8wUSF1RzlloM33zoMty/lcfdO63wUN
Jcvfzr1XM0Lu3FYVbhLPzPJrKiK3An13RcQCRhLPFSO+2ncZkg0Juf8ZStkjump7
ocfWl3oSyZCRsq7Bb8eHQjqQ8Mm4SkrOWTQuBuC8aDn6gHZLGNEuYMXsrY6Zml7I
g1W08W0TttNZn6AQNli0JTa4/X6kKknXXnfubL7lreKnlvwSDTs2bk+wOf7PMVhV
5dL1HsimJ9+jPIYXCRVx/jv0A602gWhXtSdAsM6vmaho+LA9DDOfkHJukoXqQsm0
ZYANft2sXKouLtgu8q9tBN+fqi3XEMFWgLgq3qbgOnG/waCTjHRXqfQt1qSb3N0m
xW2DPZppB5QLHdj4y7mejQ==
`protect END_PROTECTED
