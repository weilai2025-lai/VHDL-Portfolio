`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFYdfWWwEO54u42m3h/3nUrqepfCIhkWYUdDqrD29+Lr4DZU9uqnD1RM7N1eQ+kW
I1QXBhJ4usGH/zUrdP0T6gBqgi7d+PPsCEa4uDX15QT1hysykW8/2FiQ6XEHXSUv
n4pao64Y9tM9nTKDq5vLOxfZSvH46qf6IpAJzPcVI6DANr29NszwDHJih+GrfiKF
DHuj9YFdPFAi4hqZD6jmc7e9rPD8SRHX/kd9y9rb2bIMx5NbQ50we2yRAcql2DJp
esm8rKTRYwRYsEOu+jhCGMQKvDTZinTAAnIpwkvo+OQWNgJrMWclIzsHKP5as7CL
nyiDSXW17bPY5RaLWkZhhSsLnLvBv+WdlxC1iXWHan609svr1NT0R43ttQJMGmVE
XZTdDBu4nZKKov0iVVpdM5nRrBUglxydBM4PA3W8neYg0LIWpO/aRvarIf2Kep+X
Ncs9A7o3rDPWBaEjYH3GX+lnvknXR9XKgJZL/1saYcWFWgSyZtFpCEaaqt+iKj+e
zVz7Kd7diHrOFfKsVzc1+q1GoiTU4af8z+dAC+Mo+8S9JK8cT1AN6T7A2QmC6o06
QwZT33t3l+vsF1rQADQf7j7y+2D3metAYqRNADIFB36zV3FSV/gbyc2yjoYEdbFr
rvmPpFCwxbmA+mOh5ENJTzmPZMf2cta/Rep9s4XjVZ24DY4hBJptzTlXTIuW2J63
L/RazsbNcmoh3SyGd5Oi6pR2FPnG1C7f2rLRE6dOzUW1qmXiee/KPB2TOma8Zdcy
/YqntqYlmqCL43d/cP9TTqMbuPY0WW6l4SmnvGbIbxi5H8XRRbKZjt35WAgKrVXY
AidkW02rj3olPAsQWKb6qySwIc1oHThFBoNVSEux1l+3y2GT9sMJOMu3CQFuYXZk
YCT7hM+kBF4Xd6OhXA9hvHssid6G9ZMv0Tgcc+mL9XrAcfzaHOFU5PY5qfp96Ppq
Pq40W1eNOyzOzDRMnHTTFuV04GuXHOL4Hu13tCV/owu+QVIVEYLp8NVx1vVV4G+r
s0A5YWbKz+drICvoiS11mmKEq4xRX7D3thBi9K1xYtlZ+CFCCv+5S4/t5nDVB6yX
8oPBMoV41P2aKsT49jha5cwLAmTmov97f8IZDaADlubRwjhaAtv+8NofYcoUJw1N
uVbVT517ZnX34UTl9C10apACaQOHSDnK7v2pveAQgSa7qJkO7kU9WXjbmaGoAFil
ZWf0UKXDV42j+yU0Zz0WviOfnZN7OCGpWhrjQVOq1UID4djgMlQrXx1AlzJvhNQZ
DlwcegMmjgxyykAXN9i807Aid1/tJt6Jogf83g131HbyimZt2rQtVTZH6vP5Xjht
OV/ZAnAGs3wSrrSvrajNBcswkJwDGMAisFokpaMQkCDx2zXxjEcitxdY5evrMU0d
QlngVzt6BOJYo/1uDZvFFXKr22+alp6h6K+xSvRP199OJMThLj7hqzWel6au9/5Y
ZjpAy6XvcB63N2PH4cz8dovETPmzNv5seQB8+Tpv2m1znZplSbXbgRO6NMic2DcP
Jh1Jk/n7HqOhOeXOw3INmaEC769ZSEoWBKPaImurRvtmtM1WXOHxQkRQrnmFbtRg
HN1eRL+GzSRKmVudzVE2r3tlP8QIbWIjbP5uL8HxSzSQyHhBbBwb7xgtR0hII0Z4
UXuZof6oBXhSRl+UQ0r+T/bBOP84NfugExL5ah3yIIo65ZHKRjXnkxgqxzYOgsZl
upd6DLcr2LROfF6AnYhm3FMqzAdotEU6q/dniO7s0m28yqUdqQqE5sjSuUNe0xFC
LQoisOzJyKWYj2htvvBE1NPZhWYCxJUrr++CY4oMdFGsTjEng3/oI7ZZpXzvHYiG
Dtt9Zv0apkkpjNyUYqAJ6AcG812M4Almj7PSCVPBAIeFP22DzDgbiO6cSfgcZE2n
LU5Flj9747t1P6zjdGyxZZ8vD7q+MuoR1rvevj8S/S11YY6JiwCweUZWn8jmRelh
OtB9yNY7yYQfDGOnNxPAtS5Q0bz7zsnZtgf21SUuMl1I/vQkfGhlWQTBHu5iaXlX
LQJr53Q0mFGoZ5Rre3qITFcCQ1QCyDkdNHVvAuDvR46MUFj2zfnriOGFZeziQdCJ
U8fX3N5s0meZXSV0Vf+8LFX+SO9762p+9mQK9hsxpg+CcvIft6ahxpe26skXa22e
tYQ782mRGlIJCow+4RCk7MG2VAQQpkEJeSCJ3xAvAcE74mSpm++amXthAndiGCA5
Tuch2C76e5zIgKTeYP615hahTbFage4vZlpXMY0vtAev3mmfT6M3QaX4HcdZ6t+m
Q4mrLSOoGnxZk4/KxWIu7YP/8Im77GrqjQbPNPHgPsPYBnbcGeX+dxj+FR05pIoN
5rVKfyGbrvXjMpvtnXUhgfvMKpRUx3rR/oAEK41Y2plrgFAFNDoC///YiTA7UMOn
lrFjprguu7JpRQ4x6Alf0Ukh1xBDumDp2rQWUj6V2it78CrrhgQ0qC/6nkU8yrru
nPMuV5SbHrXXoyeFT+YnR6u0Ax0yXipdVrgVlqoeHgGj6RJLcEGO+ibx9KbOjKvv
OrxpoJqOUHtWvbhv7nUtIRalCkV9gI2l2qUOqC+M7cLlqYB6i/JXUgsyhw3Et95r
/ajebGymclz+HHe6K9ouibCoS7XFN4N1VQbfcUQZ/BNiRsgaSNEAI83N/HMWzeM9
ycTqAHJrYqLwplcjBG07F3TRiML3I2DKmZ6fyt1UIUPVepufuNgc7nB3UWuOHOvP
g7jgbr8LiGpWLnEiPVfgu/+W9UD+zfLilg49EZPJDuLC9XiocV098AMQOLazUZYp
RKvbSXw3pYXlBY94ci4SQEIk4LEPsdUnjzx1Yz1BhIvCJO5ay3A+cLjetYuSCIG6
Hcl9A4AR6Kaft1p/oL0p7T+O501t4WEddc1qViKh932OwCZZspC+eWFKVp5JL09C
I1pUJ/U7GnGYchLPf24dwWfE49wfsPYxz4QoXpfO7hTB7g5jJEFlNOQ6eU8EJ1fl
2J4tTQdIbjwom96oMYaA3irHeuS4NvKr/W/i0eOgVrr2Px7QCn1OhxMiDP4F8NAf
QUphJxGM7rTNST5jXKtNmIidmHEeUEWwA/txGk+uL5GobH+XeAvopBfNVWCWRL53
XGaPIpztn2TD0uEQ3fXw1QlqVjgrCzQrHtmyKF5mKn0W8n+lFE3uCAQSB4pq1QwD
4FNFD97KChKiNWdnJDxYpTSN8fhJ42ps2YaW2pSwbKBN2Ym7yOJNztATO51ZAbpC
s25/+7Ni23JSNR8/9ZYVO96dlyd/+h7ZIy+Osd07zKYR/ZZbbx6HBOf0VJmizi0a
Dgusv/MMWZwfextA3dvLmXQPjOfA/2bfmEhuXibhJ+DwerCJflveA/8JTjAZeeA2
3u39Yj7cIE+hZtG+n01VNbAVin6YS6VULvrSWO1SbNEQWoYiVuDCePvvARoipyTF
q16B0PoiGyMCW5SUO2rqcbtI5g3ZFXtmOBJn1YEalmPrZfO/+A4pVHopaVr+9ZBK
cJPEtyel+itr2PpI9YNlkTZ4vjVsKx7NisOWnQyl1dEkK42rhnHMid72jYwuAEV4
HXVWvw6bUvuYh0+sac76o64zfxtsMzwTpbkoh0BjbUrAZOlPItk2Q5IGfKA8xPT4
kmhLQitGjbc/2JWXgSaYOq/stv7FBnVnLCMFpVbxep7klZV4ID4QwV/YuOxFuPaO
pdxfj1HdudlnL4rBPN5XJ67dNnAuB1L44WcYF267vph8ulMnvCiU/qi7Oo16oo+e
gtLp4XWijbhEhRjFkZOXCNBSO7kKhRcggQbJKW7vD0mac3swN0kuaj7jPR0MZvx+
aP3/gAsvG0RTFN5TVSmeU26yK+6yEBVYcu8ZXfZ0lNN9G7jrwnfneTwBg5L8SxPz
BSR80pXEDBM5Oxcjr+H582548TOBsg7a+nfCC0+jxDboTDXvKO8HU715GPDU2+Qf
BnZIMKezzNh+FqUfcCTTgCbr8op5U0FwVEPRPQB8gWjb6GiifjyqUpCJCDdxXM6o
J08ZYPZHeG5nxqlCHoFZ4JSetmmFoRvB4JSEiRy4YZRnQC9TOYLRkqAu7D1LeXmU
PcL5kH+cenQIjDBuou7mMDOCohdTvqMPaKKgTKvkGj5J9Bw7mv3jVbMIvlduRuoy
xuD4Cy8xtMgkc088exb7/uXP2MgvfXTSIcomvy9Fy+anGFPzGjeTyRxvEgSbkvZf
HyQTCOv07e4kEhIt8YstDEevlPURWbKhZdcSLZ8ond3CCz8AxT9uNGTlC816Oa/Z
DLg2xRZE+lG8WbpyFeIgG4A1BfFOF7gfJ0LQcqD+xhO2lQ2scJOCcfpk5ScKRVlP
beAb5cgNDVEnXYOJcZNfzM3nfUN+1VrN1wswz9/o/A+ZFuaR5YVOtsyQTBXX6pqf
Z6xtX+wKpeBbxTyoH6S/hDl+0GoDcpzhdZk6q2hj54PncZ8sQnuMs4TQNARAfZZA
ehCy5nwD3fI8Nitz9dRm4dYHK6GTK+87RSmYZiFZs4ELRZxwOnKq+okya441vdbA
C4Ba47WS0hu4t0LG7E/OmrD1qpakcbI7frBqY1U5zp3FKjsV8qXuKDDcqAAkTKxa
9xeFzjxwVdLeSnq9HZhawNGBsqLoI6vOdmxHc210JZ6HteroE01vdFs9V6s7C/wA
ssN6lbqxHFkmH836vb8KDi6dnEnIcH8sr6LwIGChaFmOsP3DOYKbqW46rFicYnyn
CPKD7gS+hdYrKNwWlmp+9p88TMTGPSUDbyCtZWjSJoMEdtr8SKXcKYSukfFEiYi4
4+8mtwhUpTrnFb2rirN2vt0Q6LNPwzn8q8cjvkWSuTzDK/gp5YiDmWcFlXtrm8Ml
s7Gce7D1VZivjGfgZCJTyg9gvMAwSlr95CAUpTCv5CiwxC54dr1qP0wDSjLWMZYo
Pq6IjoPQbKI+oqkBoLW+xkRl5UJTz3dQkHXgpgw63H8XLSIniLTQREpcBr8CQd4w
i1qGqtuPzydZi8bXdZySW3UAjqvocukRKk5T/L+w39LgxEZI+6eV05m/bk07yMrG
VfsTx20cOnHbPuUa32wTsTYC5/82tjPuQiOvqWyKgPumXIosRWD2ZsTCHQTBHfeO
IOy1TeGyy9AFObCCPDo5GJCecKd0hBdk+nVeGeDF6J/QLu10uyJ6vsqgzgzI9Rub
H5RONTye06Msaf3GVmCzfpDuwalqgCOWspboIwtLH2LzzEVMUxZ67xopCcc0slxx
g8+BumGE8+1675eDuVBmLdIS1eHw9x/fLQjL5ycez8+c+sNJ6etcTXNRLuusCnoh
kY0gEqkuv0ieaToGxU2YZ9KmPGvPtc9t9NDosjPWAh8nacjeh8GeHEnwB5EgbBgg
lvfYHaqH5TnomndX9k61brl2Pi3BTRyIHtB0/y8F7udQ14b8cJpLvlA4XPqu7KaM
QFTHQvC1uoD1RqbE2Yauu3lOxa4YDyXU6rdeC0y/ih3QSbi0nXo2oyxf3bdwqJkA
VhbbBFzjQRwge5UExm6pxEINWgE17rPE2yqMhNzDamoDEFacQHkwVnhytqaFvTIQ
hUxoWmwwTqO4gjaa4g3BK52CeahfrhmKhhuiJ/LBoYwYH8OD2VvKh7JjIDfmBhhF
hbec8nwPDbVn0bFY/Y/RRxZLy1gdo1zQCiiWtWsZyrPba3exbaTxY+2vAfHoOQO6
8Ef09yJxg1xN94Sym2LnBg2dQFDKUh56ycuYcwLcVA+Jsphw6DSG+eI3XhgWUkIb
QDthMP9eeibrGLBUGETE98E2bcuvoDfShfhWoD5sZKbffwy2LHpEm25j/qEZkGS9
dXLyE/CBEBEQbPFvgw2joHjsVlivbce8/kPeGpaUI1tsKTAljBJqrKs864TOzyJF
b+KrvdL05bnGmTHgTVd16FGxKqZ782vhBCFAUZZ5gY2qNcKiLqBBeADD1ixeHQRO
YxODTpY0Yb22j+DyimzQgTzjuRuym8PZlXdzyYscC89VY0TqjTN0u+SlGOOpt/97
V/6KqnpM8luX/5KsE/L1zjd3SCNbXcQacW4OefZKfnOG7NtqeUTtXrkjgWGC6A5q
lkOJS8yGREVuiGkgLKshlWHsReevTwpU3OF7jB3tyIcXEFo4xDhgBIbGkTY1g8bG
k8Rhm2m8SQhrEFT0xDrNjpiwy+okzIU2+Epsw6H1jeaRMGOuYkPHGPag0lMV01rG
l8W23aTEdfkebFqn8bKoOAnPzbzuKKmqH8AcnCskds7/nMZL/jcae6S8D3sv84b2
Yomap9JYgRWgCsukUdHlhw8ZczhgXvXTxhzryhvfhY20M6wLeSyPnPZgtU2RVBYk
fc6hL8EuNyRk2kbywzkmCLvshx2QkhWYlt9K9kiFZz/6x+Vcfmu4dlb4YoUcRSgm
DACBd+LB0AO+zuBWi2/aAV6e5RXtNsCA5f4VbtUELtEHrlQ0bwIVsVzEw3P1WB22
EbkrSqAnOUM8RrKdiI0BDRYXLqEEzVR0N2H5Y1snQznTOKObRn7eBUMedmg0b+C7
Et8yPn95VmhPQHsqBfaiZFvk2QpawHh80S0Ah/Kkn0IIFZgpP/pxXH1ujzZE8UNi
Kpgc6g/1oBOxdsZ8WBxiNqqFFXkvZMt6E4LgeqxeuMpijNDdFSSHuEeKMAfjIZoh
xkh1x/G427tydNGSpwJtazPXEiPdRJohhsxDGM1TvZ0RbBj1vdHyAQhDXWy/uks8
aUTVzv/wAaQz1elY//HAJ5b6E0Yk9+K6BnDtIoS6jQggwryEautGHwJIXKFv3zdh
AVJRt9Ylsodq2xSJYM0HSoohESp2Cg7JFubVMJTOQOUW8FZXVRDCt9z7FBjygCcA
qt8AUVDmlyucdBIvOgsUPv7okgC4TyfuE2QibP/mNeGF0lgtbl/aSeGt0mw+IkMO
P0J58RweZkJkc97nhRxGasVMwMQyEdDNpc9VgVoW8KlKk9hBadccARJrrFKfbiqZ
9yFJes5C2McleHMYbW+Q9n9RCW8+Xg6Q4ZAJzSeq2+gEpWTjhOl/QZJbG2YDE73N
bkGOd6yB+Xp2Rnd9mGSqx6WaWQlP1gUwgm1/iqG/RkGkyMzu6H5LhrHpi+sDCf+u
iyBeKDoHd441r9En3TToMqQ9DiIioLvnt2lpvxXmbsivYYN0dAiQ4WodUsFAbsv/
qGIPlEAtNAxqJ6whsyifI9JehtKfKLaBb4d/DmjCW2lwUkyuI9iUtik+ZQC5YkJ1
aGWIlqJjYOoDsOuLf9avzQldJCLkJ424Nyx0koi+O3trVLTrlcBYo3k1Wpj7THhn
mkprgw/CbLC2DtWI/Blf343tMPNwScWLdLUp92hj9/8OfGYbPkUOEHjczvDKGQE/
6qM/tU5fUbwwEeblBMLuvPTA6W/XmlFA1u6AVnZUxrY2eOAUdZi8ynv1jb3LHPrd
TaLc0/uP9mxPk5e0PkIh4uWcYwvfIuzcXnKVv1UAWMNWMj5VQtcK2fvvdrtYKTXy
5PDOSBxNCxHkWHQ2y0rOXfvy5P32e6RSUZcirg7z+51YYElYERjpc+E+Ao9KKL1B
9mnTVd3ojlKpdr9B+CSdp9HkFCOzhLzfqtXgPwrmoHf62i980Y6lcOq9GKH6210D
SN9/B/LWO6c+vWas7BLGdn3tFwyHo6FOQzU4UfR7gNijZQvL6qdpId5wEbzcRLmj
UHi6seIOYx00sAY+eFNPVEcLNlQxWP0zNhAULo7mNNbu6J1Y3jqUH2wVn5TF1uYr
BRaSRdb5QyRYQz4zq5mKRH/QVn9sI4earLrVWFarEC996l6TrMllaiCwUYasXY9u
pvYcaetVeYcfLSlcNTsXsJXMyt8p68EdIJtq2H5ZLxIICwKiEDDrc8kyUtZTTEm/
JLiJyjJ0wxIs7uYZo7zrmdrsJmFlP/sPASUnffxKIqJJwIwUi0TTcNYiXC3NvNBY
6lJ4I/qdcC9s/CpROZ+3F7PPKzLiZjCbtDFitV9G/86po7JZJzh395O2/SmCrc9Z
Z1iLwJCH44pNvewKwVpeArocMykVMDVW4IUJOH1f5IozhLnwMzEnah/3oz+vJU6c
b7peFpyLpi43/o+mYcP80VgeSz5CkGwky6HQDwka/dUcyUFqgXUeb562dwVw0bum
6OkPyKXpqPftVn/2XYlUHnIPBZxIQvpQrRc4NJaTv3H2EymH4Q9XN0wTSCrF7d7Y
SpI9BQ97tIi9RJ4TurMF7X8RP0nWaPIIRXEASi8QD52Wc/vs4fa6+6Lpz9jV9OXz
vtGoqYKcbLPeumg8gTeylrUcjabfYGGuCIY77rOBzNg1tlEizAr/8oYgOe5OFMKG
ypjL47hp74jY5BzhhWuX1EQOkqcahVsFPBI0MeFbKrOM8lK/gnHDnvJJfOw+/g7P
Ex9MmebkBBXJ7t5BQ4Js7pk20jmNKd8Xt3nV0+Vbl+UVWBU2Cvba0CEvrIzyz8F8
pTVaWqAEw7cchIhab/XYarq5UvJHzZKqMUsLI/m5YVNPstEIWs1hUpxCg+L9QOme
bpr38A4hzvEVCS9IVNXLQYmwmMHJDvPM0pMOB13YxWHNShpbyY6XGUaVUfvZAX1f
B1A6+DcuDA+2544kfomVs7sFDwfzRkdbPI1REYL+Mco3mWqRNFA6rQyzSwj3RFVm
G0yvvr7KOyK6Ma/6x4/zoCt7ZRmdsoSixAKIhyAwAh7wTuoZw49gFU9ke1iNe+RK
62OyLVbluiD6tTw51xpjPAmBj578TCC52q29Q6NonLZ+a959Q5ydPkFzpzz10GTT
sbHHU1h6kBQtQ80+iqk5bXehrNe2tQtjPJ1bqGN36/PJTVFEhQbFv2v29VLNWuHS
WYrPzW9TOAZzJs/Jkpcl3e+ApDNydGPcZJIzIXbidDufW11OjBdXzoxcljNl/Q2+
YeNE9FYlSPHgel2xz2//XvjHAfyL4LmBydzsBLhJihVaCwmSKv8LEeN5sqEfJRsL
Uwmy9+9zconUj6XP+Oy6X+d41G0xclvr2BXICAk2duNgBMLiytwv9IUlYDtJ3mY0
DEgCHr9/xQMO9av08mp31isZGvEF+hpo59BASNnEEEGSqY5ZumAeKmQNLUAt6h5Z
plgykb809rSiwRiOwF3Oq06wf83knx6KS4FiZnN+67r4INMazgsGM6Zrc/WBde27
1Oze1AVKwf9ynkaiSvNpNp81rnhUpqYt+InY4sc0ggF4nK58kdLRYI60wmyZeb4j
G1L9/gh11lDtw/mmCHWKdtgHRi+bIUK7TNNyLb0IZGIQF0hbayE2d3ssKIywHxEh
ow3OQACyrx9pXWoxfabP6TH2WuNDaryDUiaLM+sbUikuqmlFHaMcyXNgKczxtao2
IEi9EjQllG7M5SNzQgzNyYb5FTThhKSj6/cltoK9g+ZW7IUAPBoeiZ6WMaSDWxe1
kAkE3QPzse+WeCqRXQkzWyPjnZ4Q+egcnKZbXwZK/U7IbXxWnL0St4zkt8gZpgz+
2I9mEVkM1sF1ZTPNneZ3GblaFhq9JOCGuX6Rl0yeWNd9XhI9AzgP+e/TMzsdj/R2
vq6dCTtFt8dhxm3b9LoCpeLnvNKc45u8BZtkt8BYQzo2CmADtTCw/mdgcBSRE9r8
89CzG+emGq6OJIzxxCCiW8cob6MphYHGUrFJEI845wpSZ4qG6ZDiYM66AdcYLy9b
YTBcqcY6sFRP+C/xhmSjn06v+nae4VEi2EeejxqzHvEA8wnL6OI1kX2nPmyGBJEY
+Er+L6bR2SRsBuNbwMAXcaLkDnX7xSWedswQkcNiXuDLXD9YnZP42jU4aSs/fti8
ocwLAmXm0prqXVhVj2fHkZwOLDxyeUNqbOhrf7/yhXKyikqwIb3yWboQqobpLpea
YfE7CPi8akmZS9ZEMo9Jh/xPj7HBETztajL6ps3G7jSpEhLYzR36GfuW7iFdcqzY
Arq3o6bS+VdRhTc6HSJVQJeXZuZP6/WpdlXESi7yJBPCnXGe9hf3+5N51UJswLlN
ilZtIQt7wP5/4eSirNB/NIF0kKDnAWR+UnU1Y7hZMzbuBWQp7+WxrznMUk5NqSRk
TBK2bAxvwS7J55YVdGiCXZYGd0t7eqNkBn3ySjGCG3RmztFCsNesPVbq6fXSQNqD
k0xY9v6qr/Idy7jlrpohbuZYyO9vvPFMSHUK6zToEu6u4w1MRxuuoV6WZBOblqwX
rndWQHLpSLPoVZ93c/yZsHFmzbBxNebkzPE+qZdkmBIA6oXRxx1nyAb77UFh0Gfm
AZySS92zy+bhFCmJ/wH2igcOWETRIPelvjkkUXArRBQP5bW3UMOXAhUXw0j8ogKY
sTc8MUFDoHpVgO0nNU4JVp6kvHRwHqra6bMt7j/HvUwWQKh/zzYYRelId+/MPx1N
7VGugMA/SeAJACHre8o/ZSVavFzPH90/7Ma0H06Ky6y7bdMGj9G07RFgvwQBSlFl
HuQQBNcy/DbtClvfvy9cvFUR7XdYC00Oi92VtC2FqRRLijnAZ27ItJfDNDzCMBwF
o2xxgkGsw9LfvX2iPAKQ1UNLSRQaeVGn3Qctz1wFsTuinLkizpIOs8uduBWivfAV
aP8vcYLMHPWxMyHtjH1CcAhqbdWF4TFolhbuyAyVWQImwGt4G9i9gesY1UiwvM+w
OgK/cpaBI+lLrnZy5YE/H16KNDWSKytwKru6iSCT29FnRLEn0jf1z1jNh6+AiuPs
uaV/eLQGsjQLze0/4wH0OWMBWOGVpJPEmpMCFu6J8cayqMPNG7vBIz2N/0msslXj
jDdy1+97mDtEkfwoMcOFGEvYcj2j/m43Dxb/bus37d4kDtelHL9obfMqfqylmv+P
8CaaMAs2zXZZX6IGvDmZwc+e/RmqEYBntKyAfOQl24BbnZURPwiY6jTouEcVsPFK
`protect END_PROTECTED
