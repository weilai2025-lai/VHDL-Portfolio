`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Il6QMX1fLmTZB6FARepT3Er3Gxs0Fj2sZF2pdQZudlFBR8EFH9JmDJnHX7ayx+o5
UNHcxMlmixev/92Gma88TXbo5DOMp8SMvOIXeGl8Lz/tHMBtM9LcDxVZ/FVplFm2
rN77hhXVFUSQ9mBS2xpXHpaiPUJGe6ZzcEp7ATt4P6gMdnUpiY0ZjbgQ5aSUdaWI
d7+9LkVK3vEGlaefhOeKPtQ41bGG9lQ9U9mcWtqr6dCvUPb67zZei0aiLYH2jXEy
O8rxrl2ElLFeVfslA3Fg3iXMMFWV3DvYv91NXbShsiftQTZ1UmPryhT6lszVUwZ/
n5LCjVTDwQvBs36w9kKALqYGywN72E4Wqs0702SJ1l8OfX61A8/5LkwcPVJAL3uQ
zJb/Sp70JH39fu9OCjuKa9j1S4yRYuPmFEeaPGHD4RNDWSoZn+BMor+DCLWNitOc
nnmRDtyYdrKrY0P84PV4FACwiAJYRy52HYNniZ8mUvAHzi1wvNRLu1alT4qBBwgo
a9+j8bww93V2lkeE0Y8MNanj2NqOnaPwB1zckPKTU5Q0QFuHn81uGWpmKw+GeGmE
tEvVyDhfHehW2tufpSY7QYQGe0YezKwwR4mOygY2kIsIEu7XW34kMkfxuA9BD+js
xPjg/zvgx9bYguqDdQA46GarDFO+hhqTrRbykcQvA1ZEaN+FnehrS5kRHe/9Nnqy
EsX8KiJCHvzm3WEJZDIhoV5LP//rPDU3jZaK0GaS6HbF84/c8CWAGMKXNiCYDEkL
dncdpm5WADdDoI90BKYSpYMTSb3gz6eg+5ye+Ce4UYoYKyjpSvJmsff0NXmdvvpm
F+UiqL8fqWr2YW8qOgm5qxJID55AhacLvnPvYKz6Qp/GdZ26XWBJoj385MERP8tw
pj+4cMfomLXW9uWbSPRcKdSRnjkR1gZDwBDKNgMgteSPY8HwzR7yuQzc53EuhD2n
gooTtCQAygJKWaI9YRjiYVTLVtlq8Zsr0ElGe2TEeGsg++GkEq90Jl31tUeoq7Px
3Myb/iS5bt5k+6br9WtMVDDVyAZxPxOPIjSzYLzjrTO29OMEj0R1unbj3RAsw9kp
WXc8uKyEOGvKsYnRXho6v82SU4az1VEgC0g3Uz7qIqmDPNkgND+IKC/so1ya4R3+
SygEh3LIZPpYfedEAeXcFA==
`protect END_PROTECTED
