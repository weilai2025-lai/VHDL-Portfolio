`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6lAAw5a91Rjc4s7orJwQwLbQ4b6YT8yx0uMwnNCx6DNPtYscKRZTvZRhP1e9JuA
7niDnpwQSarSRV0+Jr4Woui5nUsvv/b1DCKOGiKMg48/slVq+29EFqwF4ov62Adk
SR96QmTvLPO7HAyvNys2a99uG8pmfG0cdDiGvkcUGDT4x8lAYQdBmFkrEdAejcMT
XpofbyNmTevlSsWV8IPaLko5vo2vROZB2QTGxb0bcj7gB2mKu4GXbrXY1KpZ1Hnj
/vzuGE+C6BTN+NWpY5dCmYVxbNgUbZkBMLRahXkxVLp+BT9xagsrddM22ae1iq3c
8HDHPbIKrTqBvuKEmDD/W8peifh9IDTTc1j9x0XWB2aldXlzPe+NmF1ophc6FhO9
jB5jMVkqzsP7jC9teNo3wEUMCXKNUmebqY6A0BUp0ahM9ckqUbSddIGHueHYSlJ5
Ak+iHC9sUA4uK8u1t3wqUw==
`protect END_PROTECTED
