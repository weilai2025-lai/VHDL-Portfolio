`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEVM9fgLgK682AVSxrNm0QWzZTyaFNGk094LCeAefsWoyxcowGgT7r0auvyyS5aw
/xn5+iqdzLe0y7EI+ZYLztddoglPl2Tua3sstUk+0E04gJ463oPKh12IRMozT/WY
Pe0FoCvBcKNPptDrRUOe2D85NHtR/al9ucjQUIREPuVsGLvWjD7hxVBc2c0jHZf1
JWeNid02Zrf9QETkIG1WIkch9uzTR3r6XgnNwpZllE3k7PVf3stRxeEqgW7yUJ0X
kVQMGqZ/2UqyIpwazOsvixWOqoErX6F8o8RE2/ENemrPwtn69hjYh7H0aI32HHRj
RNYfC86iOluuayXOwzDETiVvwFB1qLn+AKF2L1HL/uGEuUGVtLSM3rbxkG11jLLD
XbVMHnHcXfRsa+HBYJKci5Ws3O2GWJtPtrdu/Fo6tH0GDZtJR0+jHAYZMJSIUOfn
vb0BA7tO8DlbhhUi89K/FjteYLe+RSpMTnG1F1R/QAabWuGurb42+79VRxzAdWZ/
ITETb/5cSDd1l7fgc4PKFK4vgHKDgx9j+l5zyoxpYR72F6zx8iMZ8dxrtB+eFXaL
lNdnSMXyyRQnP5R4eHKXUO1/XHlCUyzdg3YXtfEaoqlr31ii5Onvp+OrvXJKfDoR
JEI0/SfVZCxzz0yKbSneS8+ckKyGn6t/plN6FfIEsx4/bVZwbDn6w/g8yX4KNx7a
J9qkpEovc/UUeOD3fGqHboWzWOhVirSdX1W4Pdc4rCk37wlv8OfSoKP5maFn/EFa
JuiN4xQcUbbNnD++l8OPGOMXVrFwSWOdmTtO5igUV1TofU+v84ueDNGDhFPdaA5A
Fv+hdwbMTMaaguYnzQ9NUxAwCpixksJp8n8OwOlpF1t3wN9AbooZFc6g3nTaiEqB
anV2fK6yhmS1Lq4wBHpnoMfkOaDLLnxO7SrtZUqZe58laMLnKDc/L1xq7k4575iy
q0qhgq/236c0j4L19CPKEzExwoGc2ZZAP6NxORmGGbGh3SQ4FZEWwVM0LeExyIlG
DBTJ479sLf3Y5yKIy5ny5oDlFZyF54t81HbMJTVgkWd3wXKUrAUOk+s9Rwsh4+lF
UT+1YuE8HysWzlrtNvFADSOveNF5z5uhTm78uCEX3JdSAhtZzQdY3imJ5NllWVWy
MSZxGeq/QXn8ymCMZ/smqgvo9oEp5w4JDxUdRfHYjvMHBHgyTu72IsCCh16l4zPt
zc5qqYrynwq1NeRZA+lj+j5AI+xVBvadbKCC+cNS45LHgl/wMWZL9knQKIoDF+tG
exxlbl/D0Wa2vJsSeFw6v5XpU3l3+cWIYmLsIG8nmAqHskySsql8tWJEMStHkgNe
AzQFCXIciZ3iy+y7hVbq/3amKqpKXEEgy8LaxDqW9YIHw7dzM6NxnnOAUWGmuya4
4C9mMceF2nfume4FxzQK3NGfOKfSTorqf2+1xNNjn+RztS2u6O847UGFSdIKZC5n
uv5dnJIYtpp7/kRIO92a6Mf+qJPELWuh021nQw+pKCOkLnRQvC/VHYltusdkmX1C
r0mOLRrRIQCD24xl7AvRdLMsbPCd3FKX/qwVle4ctCFS3ZBBMGB0VSAyIRHb9pq1
YPo6ZByB8d4CpYm2pA3H2HlQQUxsshcCNATa/0JkmYkXxKfNi8wwWMnA2uu7A1Cj
sRMSUIGeOTSyEFu+vX2PgTb8n+LHtjgySW46VV6unIYxkHmFiXg/AnKIeQRVcXx3
Q+X7XFkWjp8/wkKwX2a7gmoFIIMM5IfQOl4g/oiFhxaMYc7x73IrVIcLSXDub3RM
`protect END_PROTECTED
