`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mV4sxYCEB3ljVwZ2ERfn0WA8lU354+MdfN5v5fuXMo626oJ5ZozoGn+zaiVvvFiw
aIcqXLOVj2EghAKixqBXCan6UaKeMgUAzGrAxZTSZD05mKbmcow2S3MuHuEkubJ1
wrDT7ALFzrZFp9E1rAMVZn4yh8Dh10Qpkw9RoUdmjZhTwQDmbZZH+L9bj2xnsiVL
6jWMX/55Dx+FDqxQG7Ej6Bo1KwlD8sUZxxWLCvgxvGhZA+uJgCNS28FlGW8tbTsC
akrB8ciXFALP9X9sG1ZUzeTuAI9e9fU0EDReHkzXYDN9PRBjTFF0uR9mj8JYH74k
Bt4rr4Nv8neC+txtRJnqZPOFlSCZKkWrK34UzNB9uAWyLNG/rnAQN8abuc0FRAvU
Wr1PGW5d/CRSab03jAoIqTpFK8akXrDcqUhI6BR+JJG7iBBV4Ai1aX51qENTk4q8
V3SlIQXRjLPDQ0yOACH3MIU+h3YT+l8vkxqd4mIOLZ0DcT38tqpbJokQF7CyoMsX
ZRqqBsqua9Nn2bK52xFTTijR/pOPXgHU7LBRoJiRe/GrLEkIHCDRbcf6evrRXQgl
Rsnfm1WFlsaI5klahR5DJ9CA9oxHEj7kWgHyd36T24JfRRdrsNIScdX0PiyJe0LO
/pqZVA19OySLH+eR0aY12R+PSDKwFWbXSYee534IR9BYkN6n1kxQ5m580i0BBGzU
U6R0+aA46toaQ445Fn7uQppBlnVZK1sVnwit8VLbkWOcjrUVsses3F2P6XKuYTQc
4bl2llUmkZm0x3Q32p6BD5EKxLVdb+EeSGgZqCddieGeEAa4xXXyEkKsR7xlg32S
R2w90bvi12iY6Gw4XyZDjnnc2g/D+3/IM1YGG6ifUJOqEYlnODPxmV24j9BsoQJH
3ZAyriYsm3ksI5Al79saCcI33aQManWQUW2UCZSKu5MB8jeVLNKHAS3MOuPAKndc
rRzU8ege3oeLrZPlPweq6C4mQbIS7TR5fM+jw3BPAphAlA23KCBDi5h5N11KrrXD
854jSLT+sekUh+SjtvovCGkMsrTZnmgdRpYLNX3/tgaOPHMG3/scRY9KzYGvkW8M
h5On1T0RfS2qpe3ZMmetG4hy3/FUMtoDOL5nwia0s+MWFwcmVd34uxyCseE2dcQ7
9wDdDNy8CYETJ7C5QOLIV1Cq0dB77jLa2msmCMx7gOewEer0nIbjtIolNUd5Byrq
FFCfUrfOd1mqtVCrHEcKzt1rPWnVffuse/QhkDXo07eGDcrAaV0niBzUuDF56UOc
pYYDoBD9TOROyBYplPOPaD0L/cvZ37jKzUzTM0XIw+VfqfZ44rWUs5xTqaCIYuDY
XLFoSmObd//8W6L1HC0xSBkAuawzbL2m6ht5QWgDdll2aWQjkBBWWvBmPzcCegDZ
pScNLDpBApmGghtDllNXYcrlUcuS5H/EJWlH83flqyr557HT2hXBtgOPtjhoyGrj
F6KKCvjQN97zwB+4uD3rrufQeQmS0tWteTXSQirHPJon45jW93h+D82ZiNznA9sn
qClSbkkcMeDcPUdUaeSMbBo00bGEOsLkgVH7JdsvgSB4p2EFZQ+/HxFm4/yM3mOj
naCOXvO2s0UrwQpKG2tEfI7Mu6Su5TCYb2/mCbDzTlwKEAqaSLJFn8iD3jBZ7prG
ag5hdZpO4skAZJq1wdPIweTu9vXdZG4ocwJl658I1NH0b3aawxN1Fom+X7ejTllr
yIk39GybNC+gYKgtg5c3F1TvVunH3oCjwudP0uEGSADeKhQvI+u9PzgZUhbKHnvG
AlrheiQq8UfE7G6OzzTCwqvOgmDls7zlqeDxAJ4rJ6rB5d1wTLqaRV2QpspM63Ay
cfu6yFKREFapcjdoKnyy7Suf9dMnP2ten8ULoROYkKtPNSMdjFwXSf9gMmLELj/b
EDLGZAk3OUOToT+c1QMIsX3eXk2p38w0NDrEX1ha2z8iccVgDocsbNq3VSKZ2NGR
+BTO68S1zbdJhvX78PK0pm18jWeQiFPWE6NUINrHyK66+OZrKS1tgYagpMPUduUb
9X15ZGEd0bHSg6uwbKgemPNdbFSL8zNE9/k+GDdN8p53mPJUG6m1Oe6zs2MrioXT
wSlq3wbcrFk179cTi3xIXBSX3rMitIK5kZPAOwY+32c8/mBC0XM06lptEBSyLVJf
Bg1grpfqemAhwLVyBtkE8xj2BwEp8jBqWHfbOEzpWYDCfxgAcz17M1ecJm0V0vUs
OpH3rjj7xm91zAoO0tdkgfa9NpszrIJqzpCL3nSp+Fx17P841r+0g+gxeNzs0CMI
txVFStVhKOvtyOHP5ANaf7eVEIqKy0YjgvLGYvMdSYfN0r4qWv3OX0DBYrbg3aVU
rDGIk1KEGthWnyBhMgf6VOUS3hV0QJS2i/eatC++qm09c0RpKEbVYY2XZ8hdvU9s
W8fDt6PyuLXdb99BTN+VL+T5LQW3mD+h0szfSdpaf/MHZwq3Db0LGxVuXkqLQLZk
0Ijwbz1xM7+XLhzpeIwjtbYhddeqtwL+RjcWpyrvIGXhl5gNG8R8jR3YrzjC8GVO
ibd9+J5FBLmC7TUKdJQHGgGUGG2XQCys6qAg5XFmb/TYbUtnxoHtrcxSG9GocswY
VVq1fqgK4qZaZo8dxVhWuX6ngVLbmAJiZ2PgS1ITELs6bPVnrXGobGKT6H399nyY
xBu+TIdUTa3ZSxVFgFMi8bX8MCwEXXiGsfMs2ale7B6p8yNqpku/+uaghuECooOA
wHjCXGWgWNsscS2LE1P8boIFJMGgYUr8xJo//mOx9vfh7D3MV9oBZDRgGY6o6vCC
CXPHKevcFN1Vb4HCLw9fy+DQEOfx62Sfm/j3EYYzEk752wJYxWa6kwyhjyhJ6Smi
ezGJJb2z97rjHAlXsZItd27Z9Ho0bN6F30ru2mogMRp9FF090f1KmUNNzQZrjVhy
f1sMicJ79kdIG2oIbrwsFGOXm045OW4Kj/wnM9p2Rw/a8ODelo5S9hEg2mkXXF6/
LBpRaiNNwtPcsFcuic3RgMxOd5K/CQWenL2rK/ffCGupYLiWDwe5CDZgEQDvbWOi
J5njWM3Eznn5PhIeIsiypieQVBVorqJ3Fu94doqH6QQoZQ8jjegAWnCr1oRUbZNU
fUtdmEWLvGmGSfFgFkfRDBr7il9O6JZE0j2kMCc99NCzHGiiq1pasUWFruaqQjF5
2QM2jO6aNgWz6TvrX5S5W7y6XdiXTXoH/27f1huzEETIM+TI9h7F01LQpmebZOT3
C6B52P8vj0+tQ2Km4vRUgon1lw97rNSF3RLNvedQU+p2C8CJT0F+qVreh1V4rL0N
BycFM0Skt7YvzvzM41NR5PzXiW8UUpPDRGFAfd115PpdxdQ/O3GijY9m3TUew5ed
o28C4pZf5ika8OEgEGn6YnwVB0v1MRjDiBwvL2aSqqcEQkKaNh2A1bjTUOY4ODee
nzl0gaZnGErSz6qimqWZpqaA//4oQp8lszLkvV6EMQDkdCYghst2qdCWZicox6b7
swqQrdwE2Qra8qNXzWOcG6/z23WDY/5RyCTODiPMvI3upukVYq//tYOld6tcy8D3
stgGUV8U8mpgEmJ/7ERrni69o8oDq9iWKImGNLnMf84VtS6OFyMc1t35tx3zvnFb
US5LlVJja7V9jjyJIUVVY6fxbRQ4x8VxBnfbHjV8iYuOTuQfkF012JMlF68EfHDP
yhPu+Dxc9Uj2xb/vr5cbFw==
`protect END_PROTECTED
