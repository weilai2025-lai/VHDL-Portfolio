`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e18QL7+L5z9Hn81Gsc3DRGKJlqAMoZChpupNJTIcdXILqfZhe4+6JnwZtsrdd7OV
9z9hJREJbYBO3xcAHyeNUXyTx7Gz8mV131tx3FLFrtXyWc2euVHcb2aBYvq4XbAR
ngmV5+jYBDS7tV1/cF2AHmjKAfZNMtM8ueGorCcGdYL9/uB7XXVVjtKTUdhI43mM
K7ae/xqIYYfEbHVBFDhvAI0l2tXlcnp5b01n+P4Pv+iSNtceNrG2Yx4cu3u4NamO
q/vODRwvnYxy9pZBq1RMKFIZmYe8OqiXoBsmvbyWcqbCWXq/0VAP5LY1Ugh/f8qk
YwXme4oLid8NJPP0xH2RLAec5s/Jlwrr9azMzA5ItjsE2voz7rQ7hZDCEwrds+k0
vDHLbbiF2DRIqyxkcMef6NzuxrNWoTKHy5SHCSHF9EAEFJDVckydhQJY11WJBWsU
IRQwQuumLSGsvKn6gq4PkoKe1KKpBFsN0LxUABFynUw=
`protect END_PROTECTED
