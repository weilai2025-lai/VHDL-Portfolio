`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gAw7UoYXJo7e+SS4x+mW3wYXLjdwqTCEZX9gg8FA6YXDQNoC3MvFgsqizOI/QowE
GL0FI+2R7CxpwX7vrgL360P+nclXJ5OmqDysFjpYqBCHv/eO0NcSDrcs4eV2kTvn
MQo4LLPMJG90mQ6Y2U4cyqug8YlAtmMe1hljvsYTl1OWs6l18AFf+Z8BaVCkFsHo
JZhQ09t9NPlDWnJbunGxII2RApv4EwhcR0wfTxtWwgGMvJ8xs5sm44+HsETeecgY
nVgKpIqpxL68JEoaAA1OazYK04Zm8BiT/atImjA0qAhLD4cI6M+/HRDzIYHPK8fx
KrFduT5PbQyhRe3OuZc2G/I2m956PnsGWmgIF2+UatC0Y1hfiKMl9JvLPtfHHsGi
aA2RmIA2v6VW9Qo/kdarIQXFssnnaiC+IDSS3kkL9KMqFI5woafQvULmuCRV+cIu
QyyhuyfwICkJ3/tChghT8NWRgiCTVBf651TQDvhAFHDc29FDMcfavfYRSSur/oVv
uvtqwIrujSkzp236JcRd16B/rd1Sas1+pOWYiL5DUKaQtF6rVzolS4inHCixTiuF
3uaBUBxTmbI8eC20SEUh1sRMoMjmhFS3sx6iPOxwJvztHkxHPjaUB47rtQEuraJr
kWpe3OpGT3BNc8AIS07bIBZNbX2yWap88V8LgUvt4oMYAT+FtS6caeRXpPUPkeVM
q3jCib8sQnMFSI/08byGIA9no42tvcYw5coNW9warmifbC+nI7spmS43JyIKDEA+
zL+6jHiaV5kzPe4ft1oVQz7AQG/LNiuG6jRRoUWUGxAmc5eoAGFyJgBgJkcY0T/7
yJSJz5IMBxIXmtTWwosNh92GcfLfa8sg51q1NSXYE65hgLXjAZSnrJl63tMo72wM
Ysk64kK65nWfu2cEAbnZMI1pfkXBup+YBzqk1oCvXdjegoHJ65TsSWpk04bahCWG
gK8NA/3G1uLQ/N7eeH6IYQYsYsKWpx5PSxisGzGuGJ5bmiMOBCNBdZvstQYCg64e
/6TwaoYXbqde4EQvxn8y2AcLH6FTb1LWwRBwwR0rGa5FOJpJlbaZB2Z0s57exjv2
eI1DCtCSaAYKYf/8VDL3C8m/In2yThUSRletGkNxpAGlbHnudyD8SCQdiukWH/0G
r/nIVmZ6xNNCLuV6iUPfhlwYMdjwW0EGpmqWmscaf0KY0Y+4V+KHaZ2Do5/k37uU
SAdSjviiL8aqW1OYx2CsoJSfl3wm6nyMxUCTGh+6Q/f1C/Iw8SKd4X7hMLHDd3bx
VPwt/vhzpQhMM3TITeHy9xVDYPl04K9tBZJqkVpp2bv34LymRI7vqoSZ0764cF8P
JATkMClYAvNhuHhWO7kOhw2F5m5sDRXNHH+EkzvEKlbmp//BCbEAncxexeEdTSGV
Bc0RBEj8c5RqayNbF78wJnZsuCXROg4KxlJ5nw01BajsbkNWKNoijwTLkkogJ+la
OZX8NW+fGRXO7LlLmjAciCzKT/TCb7ISeU3ZRWhQAVq3wMe2N0/0MCEZ7ecVhdud
bn1a8mfYAQ9/GqVQRprMKD4unmRzQrcb1BKk+WRgW0ie0Bu1jBf2iTAJSRWUuaXt
0+074NQnEYLjvrDFVA3LVL5APoCg4uIUEOW/RGia7IS6r+wr6ov+fq9DTz6Xx8tS
93XyQwxXl2aK+eSUppsvqiTio6WRUfAzzvAcsiViluZBKc9akW7O/Vrr+co8kTkg
xbBZIKT6pueDFUkPDaIlzoKZ3Bv9pWsv9HJwullhctMo6sX3dokXpZFTf5brA8mh
oVnMvAFtBsd/h3GX0hT4WWn1lrbCk0zGygvl72Xn/zhZqeXAQ7QnmUHdEiH2FJy/
0KhlS9PIapR802G+iMIrff6rujIC03GsRrFiufwEEXDbArbApbgdcGIBlCsM6q4G
qLSK57HdDRdiu5Of4GMuTzVuFC1Pj4nx70jPvGo40zs=
`protect END_PROTECTED
