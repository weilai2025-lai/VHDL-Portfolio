`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fJS/1SXgyIJ4gY1IhpuJX2AGEL00zHksuyH+pxP9eyvrGATZ1NEXHSAZf/H7vi7t
akjp+jxZPhyvY4g4nBzNb4jm+cMLlbWvNOo9UU4YZ5SuYJI+/SQBr849JbjVYLZ5
8drzZWEtlH9z/PkFjp9Q5IBI5QGHl8RMfdxfisAZ1NaIGLVSKHvd8LAyfByiFDnc
7GmEKXq3JufOEfoGHb9lPimOe09ag+StWi/PO5tv18iEu9inmL2vvJ3P61c5ZEJP
6tMUIAmKY+V4CoOP5IyFqHAlugnXroz/FfccYwMQtMtxux6bmtzmcbilab9hMB/4
aL4Grz7no4tTZXGSJNKhUmx/Lu90HHCkW2fSxflv3JGs9dGjJgnfBeksETFzhh3K
ELn4wKiAyPdT9HyuYbRCK3ZALVyjYqn6qon72dwnu3BmbZ8cPETKJNocgNXIy2PI
rDhPX6Mc13WJXMDNSQMyY2EoZP4cDm+RaxkfOppavmMFsnQrtpOWnJEzrf2oPtIU
HI5lMo28Q1wtNhb4Z74Wqe/chpgQnJm+e1o9pvv4JQOBrSknZgbMU6pWSxqWlZNt
n8MYaFD0kszngQYwWwkFkaVFiOeDt8PhCVK69UXp6bPx0Sw6FT0U1EDqEqEGSSkb
A+7OrBf3gha12UDuvDWAY99N7IAFXmypropD3cckfVbCSUsmppRbtnb1cUTP8vHV
6SrkTsRYuicjO4mUWEuKU+Z181vArEIHjZicw85r3BeH0AwBqIKxuhO4l/Z3C8Jp
aKyXI1Sa06WndHffHJIXCJrSO5qAYrPxk+C7bKPpEl7dJdFBmQMTtTRhoegAt0qX
1GEQqY3B0hMu+QWeZ5mAYCDk8YwqHIr3NMxDQOSSi9/K35sXMlLYG7p/mvQv7QOh
5UdpHzqmuB9Ni9lFtX93qVWzC00mm5s73+g6ALZCm/FRQRfBDrIWDz0a6rCtR6b3
9VqNbDhxSY8dMCDfxw/lPvyA/Ma/R6VgGYk2M50UYpM03scAkJ8IarAYRYy2d7YY
73hBVWdSBdC+EVPQKf+ll9bzPI0wZ7PuUVJ/16fpCP1y1B/G2k+GL3Dqprztrd5t
Y5GOegN0ZGdaKWEQaMvYm2w1NmpBnUPm2+0qdalkZkiaNYgjb6v4zoO/OvLcP69e
WhEnRIdwuKeueXiizSpnO/+XUgoA/iwyRWBuHu2/iaQJusMaVRtwy0Ks//KvMbfG
k0VuNpKXKbjEKSpe0xeOiArRXcnonAuPkTc6txseQDrXsERL8V0rRn/yyfFfdrzW
We/RKvQhGk0akBa6D1hOUMgwrQOj0Q8bedCuPr9bqcybX8Ma7/fB4cS2Td5oSg7I
cVJt31mgnkJp+3hdLOxw79J879HSPYfb+Mxay2EbvDuSvhKa5eiZAcw7yOjo2BGf
S/lSXToPZrFXPsmYSavhJvLBEmMV7JCbQNEDFFUuuoBVdj5F9ft4AjIKc5GP+Fv9
dIW+Yhpmk/8pRfuQLqe3eBtQp6rOfEYwWg6v/7rfEqXNGTdlDEqCkAfjk5k6aPMZ
8KP/L/S5GiqbCMA2F/oLMBwJW7Pp8VCIxqAtIbwmT/73SjYAVZysIyLIpvVpUJ5g
xSy7WBBWl9F0mxLDbVIvZQlHpkE0IJm9Mi3XpHd7QpwIlr7vcoLIcuPcEsnCQ2H2
Q/qNIJyokAuKIy8fkTNa/rTtwk6sJW2S1T58Kz/NSuQAdx/vOZ9sZuu1x/JiFDy1
qySnATU3xPhA/pKdapm3BGMzdYQDcWm4VONptIjRrbV2eFTfPPL0eMlyyHbJ1nSO
naZJP1GiTzdk82b3b0c99yli0SF2MdiCUfD+GVNQ1dSaZDhS8FovnPNIb35LwQ6B
EKABAeFDjHt124FYvSCqs55uSf+LB4/w4G/iwFll1X8+YxVFnkHLncVf30umHPXR
jStK6yU8xV0IfjxHvtWH/DXwrflmcJtP7BaK95vIq75mHUS43H7h5438gddb18Qc
Sb+LkBY9ZAqI3ztK9vlBz5SnTuLS3iuadZKZnXw/7iZRXnLtToCiXyGRsLunBmGa
jbkfpvdZqrf01h/QYV5FwIAI/9EPVS6llp2Lob4Yb5bV26tHk4lIbLIO3oLK3LiK
2jzUdeMOfsmm4+/9SzFPy+rBuyIvs1l4Xze5tyJJOiXoBerwN8F0pE6UktS1YKUq
DiHO5AXN90cPPN0yGUrxDh3kLjA8Ovf89pxppC539K2seq41EZ000yApxuoo9byl
namuHQlUd/H8A23NvA8aff9uEfL89uX82HNjUnF/D/hsndVESS78o64useUye3QS
cnJGHaeI683GsGg2bZ686/hgurNydHq5Pne9oMzjnc2p2Ncz2+STw9vvHmMUCjBb
uPBZd54YTte7UaiFLxUpf19eTXCCPGRHAjTbL4bAJPjoEkt6s/HM2ws8kHVTNGmm
zTD+Eg/wnwW3pPga62hu34T34CtkAuAF5OcL388hGHPgJYLfQSK0dDEeJ3OXVco7
K82jRvcI1Qo4JM0tGXQ8AGht+vSrA5yJk+5GK1JvL98M5TR77dgvBEvmZOu5W8z0
aY0+DVsbanK5O6Pb2cYzu4HD09dlCxpdbQO/1zSk4h6BDUY3ET39yy3/x045YEdP
Vg/Qgqfc07EJH6tbS7RAZDjVmZMBVQSwp/sjdbPRRYOFvXPZOiHFp9mAEFFZ5fc9
Mr1VcSU7o7G+Gf1DkmhynwMupu5uhwSv0wi0wz2egL9o64au4fTH1DQ+7pc/lKA5
6b3gT/IYqH/1xg3gsJHFwhEMMgRKz+fB8716YBxENdyW6bbpaYTs38Lys5BaqgtJ
kS1S261xdUCdns4AM85ZclpiVp1qPGClfK+cCoQcUwddnekKeC7blMWT60EPXhG7
7elI7icr0XhOuvlFvuC46CU28sbMT/R/6HBE52mIkDOEogyWrdDc2tRQEoHN+S0d
9+CpYvrlMbkZmKP2xdG6PUr4aqgU0ymmKkyDjskIpTLFOUpv7bdo/u6wk0Z0L8gC
YZWKMDphxtarjIEAcH8dkcIKVRFxXKJ1yEXL2bXIyWD7kNEtykl6W5o1IKvQHkWO
6n0qjp6HHSWWwje9poEMVaV2INWjQLgzAY0LNImPitCmJP2AizbIW4FVkolV2ByF
jeB404sXGF3iELdNHHm461CRslgG6Uq17BUpwiWLmDk9skR18Fekn+A0QpEd89Hy
AE+juED9VaajLblGAXCkO207pXSvWnzgNcXtWlRSl8deIDAcufGwBRte3GwyuKkA
e4zP3XwE8zJA3AtDm/cOnNwk6WY/5M6vK8IPZKf0dJQ/V7psrxbYKcCvlPXW7Lpt
uvm5fkVmDT3mhXKrkcpHcX+NfBedrp4J9uzze1FNdD4f8ggv1Gk57Hg81Qlzprfv
SYRR+dYIgC2aYqkG3w+sxobEzCrPnIe4Wfp63DgHFhUEvweE6Dd1NWKGSSfBR6hP
Q4RdxCgojZbw4WTPz6oCXAPNfZIIn4xKUkqMTugabL5L8Yn0AKgpFvEIW1WK53Y1
tjvtYvp2WozW22mTzbCK/VyuUi94yrJPLwabojluypn47yBr5a/jyFxp0mbeivL9
xUYEtfVxuO/+K4lp012HbT4RC34TSQhdimdTBTNVCojOJfhEONjQiTVloIPAkWph
d5XWNPsRv/0rgB0hHvK9zQqnUw+Go3FCQN+Q7N+dMOxmZsqfcqMiDdSaDNavGVmi
LEJvPCeDTJuXVm4eTL1K/2kY+31fWZjvO8g8INAmEZvn4FZTQH80FRYFg+k92SSL
8uhqP++dDbZqsSwazpApT4lM5g6nhCazoiRtIWlIGs2DcOoStJf/Mi+/wM5dlItA
oM/0WwcARooBTfydmtDyntAWFA9Aa5Y4xOWzlC4hy2xFi8WhC0TFM68T3cPvRSWR
wXJIbGLrUy1h3Ez6Rvv5BThSkJk243x1FnJC9j4KYHeaXJs3lLBZLJjGdnYuqSca
nJy9yBnwdH/Ig0w0caTvM4HOVsCe1UhhIMwqBV9rnK8LBNOwRFgfAA2/M86FkW98
CJVHuVvsMQbDSwTlZE/iUT5Gj2ipNCw/GwQOv4T8cD9KE6YpPdow96GQ+d67eWmU
CtggA9XZq603ODme+gEZLLQvEiKpHz6h2jxK+Pa70a5s54d83GRinzGG2oJ1u1l4
vPOlBS57cVOIvKczjFUAP5g2c3F+DhLm0fsAV86yP6eGVgR1LhlZarRbH2S7OZFI
mY9UFDviIlqDMIvnhc97a2tiLcXZosx7wfPQEJvj/mb1gVw0e8srgdUdpar6nV+f
0CiJFNGqWwGjCOMvGG/+zUl2quNPivNrL8MUbFsUzMwt4Z6tzdgwKJXmdteelZi7
/JtBd6X0tuy9NsyIigWy3LsDHBaTGR59dDXlwaStjaQ2wiL3awsxZsCrrOSIul1Z
VIYTAownqadj3RRwr69mTv8p0vZKI2FZuZE4eRq1IvXq2zIcEZLhyvOYFYF1Odcg
RrCtWDGQFOEsyOeu2Vyq3u9AM4oKIoTXf8U62+ajQHSDhHLMZMC+O7osq3idzSHL
Au+vol8GhkdcDXlFtTDvihZcWePE6S6RAlb+2N9N1keWcpFHNY/NgVqtetVzsHQz
tsYvLEznEZhUPg/fvdVcz+f6rJvfew5nRSJuC0hcmfk//o7FGxyE0RS4Djvtsq7S
xfxvviXjs6Ue4WSDJBJ6vufnJDcKmF8pYzfiYF6j28jc3jbNA76CQk5lLf+fKNsU
eOnjZ2tbtI3AdAK8t5NBce6Quck6/EjbWeuYmmXp+UwO6JhK/Zd1cd0Pw4bQWHUM
IsP+Pr9+VXdrVvYj3pa0cBSmha3bYnkQDyac++TnASYJKsoTehQjhCOOXcI9CkTj
gSkbQKVcYRK9cqnX/clh+Spix30LeRUzyzjhJsmwO+8K5BDSt6HD0q3Mtn+4Gf6k
+V8VQwc8TtHtLy8VCBdIoMMtlRgMrrETSa7sJ2D0JguCWLkvUIcCkxoORNGAWqyr
1VkZaJs3LwUrZSR7bUGaAyPzazxh88CLM0HxIVf1xSgy6ABEkUEqA8IXGi8p1bQR
EVV3saCpXvySXydPSys+LKMrw03xTM5qoBnOgW7pc5Y3gQDKkwu8+5Ptod84BI1K
3lGLyRrl43gPv1jOpsdSZOBWrMT+VQiNrZu7prGuxjfv86t8XsiOJgFK4O0qEnUy
dUNxotGMjjIORwo9GpTKMzPu4ToD6RZsdBUg3xpakXmwFA1EyIX1aZLNXKF9ZoN9
VAXqiIUIHft5CSUWa4GvcAxR6ZADStjYmKk+DGtv6aBB7yz6HrBw0x/OSRguNfCm
sx0V/qcIDijLZIXBqsL0QiCH8UO2gIHj+Dm7oV0cQEhsN+3bKb2ujzrDwRFyuIgA
G4789kl+Ic+sZRT3/GaFqAiwXLkS7oooFsjqF8TsIx1/uHK7jsE/VpYiG78e6yFW
/41/d/x/yOeVuHoK7IAxPc30yu24jwFFl+0iAFDaifwJl5cZ0gMv5oiZ6QFa1BJJ
8/c600683Q9ys0By8r0mqgZGgtn+Mx14ki+7gRtKneRpbqK9GZFImM0vj2VY6GnF
+3TSEreUDssKdpzNl86FHfHYO9L7r9JGPA4ka8VykUy5POhs7TF9X0kBKDGACJfI
ZeYBtdqfubGOclOAc/bS55huuzfQrhVrneC0yEjHtHddQlQuBgwi+Me7j2TJCRL3
6JPO+/8CyM4DUk/A5qLGu+kMGip1PxFZA5ewLzoCtMoMHHb30K4gSrc/hBpzweRe
98A6TLz4boy0yDCcjdKi/5vL24zGo7enNUjR8U4PfGTSgm7JBIrG6c2k/FjH2ojJ
+xnNDEAH2CGFJzBn86HeD+lttAfP7+tXxgSTrmJAwUXDllfRrkBTjm3AG19AJwn2
UV+BYz1ufMEyoVotUSosWceu30LnR51mbZMgeglbNSRc+/MtQrghLYAbXb/El9co
DC3U5zZsv1BBoO/zJ9HfO7o3A/tnbbjyqri06HI+jATuJwHsS0CY52LO7pGetoxW
fgGJmRsY2oKnlyWihraqs6gR82nC7RlipmdRPhjDIv1Taf3P3FRem92Qcs0tfLe5
5ee/Fm6BtsPnQkbhZhC1n31t4/Na+E0o8yLk3xQ3LjaxJcRPyk2KLopLkpGMesRC
AO5VNONmbuxk/rUGnEQuGGoTASy509D5hOe9YagVmRZASPK2uHKnKQNBmewA/NZu
bo3WX61eMDOXaWAtF+XF1lqiDuxx621HEvEjyNkSJc3ZuJwes9B3tDP7IGb+/KNm
dqW7vipz//jfwHeaDoqaxOfX/5Q7gLdOzPW4N4TzJUqj3B0G4VWtQPB5IjmXkql6
yccfp1oXc/daEMeEnefb7zIJZOaCFcm5rKas7GJ/8egfakP6o15/qqUE5wAVATbJ
lfXQbBeg/X9RC4uSKZykxCLYC/bkGxT4zWLICeNp+qnxngi+RT4OlzuUsMpwsa4m
bp7yRgWIYlEG7aQBR2R67RCqhxiiPQ5Qm7McubV5aCoiv0yCHCyTZakUhlGgSPAE
YdvINrfoYZyoLmxu+LAuKmjCe6huaditrsmGOfz+t5O6yLJhBd76w2XfUEjCsk0m
z/x/i9IseUjOe5xf3CZ8OEboJAen0299aNe6rEKrG8J34Jwf+bGTKUEyABl4lqsI
XJsWlmHzTC38N6pV+KdvC1X4K3+XWm2YAy9BztNLiMNPkc/mkjkwObjQimTQ1/Fs
5ep6jIdWE1zy7ELxFJ6x1OekD4gPvey8tMRYmLsb/N7ev7xiU4l3qilPpUIOSJ5P
1pFkyDEahIvuXCffhMFmfub8dCtNphIsKscAWKimueATSLIhUY4EkEF5h2CpAj3/
NVHqsJYTIQTDafoTdVHahouOMehA7TwoAy4GA9socdsi9v2DMTdEOU7xL50qA9ki
0ghF9FJSI2fmRTwBnOHZDd4jhcSjc7AtwCXUYTcwq4sk7W3Nzgcu7dB1PgXOgD23
SSNHgw3ORBninynkyGXDuVei/55NtkU+nognjd2TadedFusHyV3X7tlcRHTGmF24
aWIXz1V51pHDURwVeIIgTCIHiovGce2Yw6/u/q5WHAsS2znmymyJ+wzkx9wI2uS9
3m5WemouiiJfICxNfMJ3/TqY9r8vqZrsq347+gpMlmOYfFbTwaoeJ0CsKju3e5ip
9CNJFecrCnQAQL+Bif5HESSheO0dOO91B7oryKlbnekI0mcsCr8+9+KcX8NBA7Pc
n8zs4J5Jy8Qn5qrJtlEkpZPKeakH35aPvC3GtWMheMWVs7jrCVsVaooKvI5VuSZy
iVvJMx8uHopHszuWYhYA/Nhoszc8xgAasn1FToduenJ+A4i52akb9hf9cJpSzILa
dBdJCIFfSyOLLYOsomhDuiyDcvKq18nac3HAGXe4Iha3syXr+wtPcE75gwb7mFVB
2fTjvaMw95lTHgd7UOvMCWsd1X0eZZC5xXuJQyARTWcdgZWd0fbk9P7Y+VdDyWr3
YuOPRD4zjS0brisePuRzWPLY5tkWFd5X4251aavPX+EsorOQSe8JNAb6s8P4Z47K
ufKYtukznB0ozobHjbaCPhwbXzSIsKdUW4QnwNAC25QppFaX9Kess4hgQLZ3/itA
zBSPSjVcV3ZxSYqPCEiNgzbP+nuht7Nxi49VPPZbyN2F5TEx7iBNn1NMZZpstKyD
Lfyk1FG/Qnxfr6DEtUC4RpW5oDK2RuN3jfZGg6p2dScSo2tjnWQDaB65KSJL6Wtl
xT7u2+y6KMZWsUAuUKkp9qaIor6kZYIkUzJ2j7Dmm1t7eWCnV7O4p0Q2CqhPWPBU
CzrlaWLyHDco5WrV5ynVpsWqFylgixckKUlTOsdCDq8r5Scl+hKMs9fuhGCDqO9B
r4CGHgjXCun//otnb6223zLSJ5YVP/E86goGFiLoBJzLNem4OxBWff65R6XBeiM2
4jM83usp/MYZNEY0cBwLzZGbQWAXHcpUMuy2brFGxz5bNhX1EoGm9AbBpOzof+CH
BEwXDB3eKECXjCrwz1HfLRHFg3mymAFnUN2aKErHZ/OFjHHSUvDVnnSH7cjU1FK9
yacRL+n2iMwm/QcUWXGI/3b5ZR2+pykkpbdVcCzvC+PtPeuKuKi7Tw8BbFv05LDV
ATgrpOd4EzGzospcQ+Dh2DTrnqcEL9P8GmVoIM6Gkz+14oQYCLJpyCWxBsBj1rKK
hfnVmlirN5Z3NYriTh9jr7AY1p2OjpKAUukZhRXvjCN+0sJAM/DjSydT+cpJb/6z
Geo3KLUWlMMgHbDEn07vZ/pQsTwS0i5igjxi2CKVmrRo9VVD+FwLOqlGnyrN3uBF
AfmhMOtjOh7ZU+wK4POvV5DMN3hYD6ozcMThaNWbN1DHhZE6zX3FUNpvo2/BssLF
VO1uE+LIXYdpIWu1bZqHWAsRFayG01XWCUqJOszTu/Dmau1AV1QGTN+qiubnAysm
BsCwBYHbeXEAYDop8z0JOlBwbogYUCOXGJb3cwBHv0q3m1ruNm4OtfKDfD/OJrKZ
xLhklP+jX6qaN6AxQuQvBEiIqD0VKTbEQ40JHaKW0YvfnVRehTO/eGtwrYNi4oz6
rTotIfvVRb3rwXB0s9pvUJmBvxaI7c9+L5xjZ9zg626ERLzfsmd8TNuBNm+T68Qe
t4XP2wfA2bYAlFoXUWbV2v6aFInY+k3hlKVLztRxCEIm8KboEz9KwxXxAsNgj0eO
lAxc5+A86NEn30abU3h2T9NnzXbiqmCI7jjkZkxdIpS76UcPBmQRRAiLlF77wCX5
peGX/qnoN2Xx7B0jrYr8oVx6R67G8S1zbGwQBnCnHofiUld19nLRVVopgkKZ7+lV
63jVYzV0wXVwm/iHEmVIMh2ftCERg8nYEIKipDdR8p6Bg9FzRE4svDdxGJoi1udy
3UqTVh04oDb0fu1l2zeEcNxL4g7+dv7fjWxTuqRYgSmiAdZDr1nh0sTCS91rS7MR
UordhFTzAsafiViXWdvGXT+sWKOS3m4B6H/vOdzWYrX3oJSySLYZys1KWqhQ5M9J
emIyy2riuLJ1wEvS43wmj97WiAlZ2m/qmxy3MGXUs9n1ZMKjUlOw6M/oUTjmVyok
h8Wyu+BoHluy5RzAFVZfWaL8ReOqcr+kle6G/Jp5RQHiBKjnDYs2m+HmxvKRznGP
G52jsDTWwFLZA9M+sOR5P7fYYF4oKNpYcIRlg4fVsx5jUEJixHgB6teyuYNHZe0g
hN1RmJmwyQnPuy2H1V75oLdq4TXoqnB50Cuo7oBjl7LddyH7gfTldyAd5heuETJD
Z1Bc6MXoxzt7lIaPRELDRP6ucSyrsYfZU1ZC8zGA06hl5B58BQTJyP7Pa3A2pnll
FtQontDY5Nc/9N4Rk3Pe34enkEX1EhqTLaCpXNOcls3qLh4NgDkxHXtke1qaIYAm
6kSYA42HGo2NPzOdOTyuT1pOo0TVBd5HzdtxhiaVbzIG2nt+TNcvWPM+3LfUX26B
C9obL+74XqkorA8IZA8cOT8jnnYwEIq5tSVF15Z99t3nBrmBqm4D0vskr0UUOWlN
ifnDweOz6IX6TSqK0+4SH3vt4+hozxSxu9mmclGzPOjHtvecXpNVyzOAWwWgAuaE
KbO+0d6cmznPHd0XT5BLCtIRjEf8svhZVERYAee2vASac1F8en4lPfctxryJTcWE
mW66xU9xHKsn9ki3ZyyU+sN4S+K65Vp5KcteArHDBdSQCu/+bsY3Fw6Yu21w9YP1
eUmDwijmu1zcaSyd7DE5pjqJ9AMucRHsUFLqueior6nujXOtBE36kUL/ygEkLzrN
1fF/NMbJJ2unn0psIWzdn0OYPiNg6x8X/oF+AWhMZ8SKNBsvYhWuTnFhD0CyFqiP
xKKzjLRozGfCxJrNLZ+32N+LjYWWAHmMwz2whzeVLyLoZk/BK68E0QpLgo2IXOsM
hMsVr7cw72CUjBhqn6/WZPxMW7cFOjVLtz7VA0j/rUwUvFr0GtcqoCARvwv3KSAF
IHlKdf3jl4wrhx4zRJ75EccyuGbW8O3MqBkDP3MfV6jIMGMmyO72ZxagGYed7D85
5gFfH6YCr37hfN+qpnccgfcWz4VyeqlUt1nj3nam11xe/zu+LqbGbwG4TlH4KuiV
cYkbm0NX+3h7qRXsjN6bG615Zg9W7P6m7dF1+JhwCbIB/tcGfiJUmI6p93jsJcVL
0i3Mid88F7aCnD6pFPXfJtUEBwd5lTRn8XhADAjTcxR3SU4RLX5/8vzn5B1F0fpc
0RvX+b+f59ZOvOD863pwPOSetKSSCAiCLRN3S81rg5W2EZ/ksUPCbc4gzNBPbzTf
jkw5u73e44aLQ+fiXL/VdTuuQG/3b/CE3N9BvWJ3ESaOJRph/1lt3EBaIdH5DTSq
DKqBjw7q+FZj/TCA7y9CuxDn//nZSMXNXfG9oVNI+6cExYaH237lnskmhL3s7LJA
SBI/W227XAi86bYxniKZIr3OzwSlgBJb/tuF4dSYSe0W3lzkldSSUNm8GvIs8tC7
VvXQfq73+D8VhnWAX3PEXvEN0Daa7drXEdcrSoWfwJJ+ruf71MQg+CAssn50D+Bd
K2SQPKI0n43jTe8LdQyVxzuGvXVOxswfpFXpezjAHxXAPgSRC8m6VjaU7Ipf+iu+
M+BHey00GkC87Q7TZS1IT7AdfNTmiAXhiQb9PtbmkMM17xvtvu1icTZGED3/xXO+
oUUE61WVk7CQFtaLog+rBQU9n8GEirGSW6PRz/x0rlbqIe4Ef+Aalag6dYIGxnRG
Y8+hkEay/m7/Ri3SlRXTsAJlStrN2hKRwbRZPGz7hjwowiNm97niT2C47C8VkS/C
/ziHASNUC3XjaFzuohaKcVp8oG9SK9krNMtAb/aUlDKs1MHafsXPDt+qLDO74jKi
iWWeFgOIGTO41bqOJo7i0rp0RFULP6pbOXduZroa6oyKOR6BGiiuvjcrcLWf6ZcP
gFBz/RKbyg3UZaDK2i3lPMDcHZ54TfBVXh3BIJrwngFGlaVxRf/xHcNY6/5wk481
QrZ7fNk87Szam/yrJSTNk9ON6r7n6BJfXFG910N8mQ0vW6n1wmmoXr+3OfZxW/Kw
r3zIOuRF5HJ4q0omlvBjsXVv7uHyU89rXElWnEFSHiQHUxkzlu5Ta7y3XgTE+OvE
5J3y3NtvuZ4TbBg9U9kFffV3y0p0yS40m1ZWpDkfbS5ylm7RN7Ga2znhLeCF0VLI
3omBV60CO5JJCs6KAAfePhK3HxmvOFho9+Nf6q+RAyW3fE4P7B9EHUz+UhtuTKLE
VuXZLEHwB9lpRjEJJN/yDUo1mJiVVXllMUF+I9ZT0M56XMXQ67IWy8zeoPTiUnNX
+wGXbNI4HDxaO2UopKRIAIZ43r8Q2dN9p7d0DQf3d4TPzCVOdudKSxvHG8X0kokN
SLF+P8yqnD3FwKgxl5TQHgfhVsGtcDUJ5kqd4wrJ8Xjukh/2t6lMJqRD2FEyHo8V
PkuF/1SQVGrH1CfI9noVOLa8yabb6859C5DlKZyZETVp7aMIiimTY/Os87PfGud8
rt4dBIqnZDJ9U3iCB2BpE+8qxe/bNDOS9AuTUxHEmh8+EGdYg+nV/W7ZLDy5ovUs
o1tChB65WFwa/7jkD/XGZUGDbi+wDS2HkTqGciHpF8ALViKtNq8H0Jt9gCKM6re6
WFXoU9mnIoreB/oSwF8CHmIgdm8SaRxD9Gok1UCw+4yhP1pSN2itPHCB2WdOr+oy
xAXDrZBmluX2GpMI+ejZXfFrarp3LIQdxYs8Q1R+x8kaOYrCYBWZG6wCSOxBo1ul
Bb6Pbb6quWQ/9T7dYrMNxBy9FpN4Hq6+nrBFA0WNDBjwVk9p5x2HAqkZxFMDGgGc
UJYFXQ8sE4apifHJbpauxE6ozmD+9toMfJCuFXoSxDI+e5YoWGgxcCmYcfEcnrOl
a+nrdjBP5MN//i/5rn8v4zL3evhBfYKGK1ZbPbSadUb8VZ0VmPdpq0WM2BPnlCUM
nsXYPCgvHX/eWID9eb3o+HiCwJIr6ZkQOYYhCvoQdbf8l5MkBLs7DHJVSlCME60B
jH2Ze8KTAI0suqGUgakEil8QThiAytlRpdojj7HrHHvviGFWv0XH43CvHh2dHM8G
i/w9zaLbb/tLQKiSWCTJwh33nxEEuZE0gKEJ0vmzquxBzNqZeWij7MRrQT3u+uw2
oizL1suAm6G6A4Jg+b+K1OBOJPBBWHxnCIEFU/U7z9P0UMynvmDPWOqY4qfNr8Dl
ISV1ejzNN+jGeI3TJTphqcYR+Wf958ctMTm6SSU5Gl9iB7i/qssgDxqNiRUnmezO
ExfF9gEJkfnQJhn8Dmf+cC7F4huFTfavMft0UqDGoWfhvMK7kD4getah3bkALm6m
WcMuixguLBG/+3PYZMw++p5ElMiVzDsABmSPkuIJLsW0xJkxO4QQ+3QBs51Y4ASc
bZQ/hIy7hFHqLqs8AXqr0zHQU2DPf5Re8kxZ8AairzwbS4wnsRM1/QTVWLOB2s/N
S3Mzct6IT/e+S3J9UsB9liyUyNw+kix2KVg0/dwkDCKHk/rtPBPP/Nj/e/Hbf7oE
QUBPcgLMsPeJLuWoID+5AHCloP4Xk8HDrruRUQ7zEx0rbyuQyKHXoBoIaR3oHBLU
FWWgV68f2AOKI+KZESmH4r2h/PeQXFzGONQl/y7C3VAre/O4wjUYk/Zm+E/JPpAC
IxXRmQemvgAZ9VwCgbVswDGvT/k6dlgN+OM46USXskPsyKbNQQxowZouyyWLvC4F
vlc1U0EsDjjOGe9ftI08hRLwTTlZzBtkw+CBWyn91N3Vvu0NcV5rKJZFUfPlcBMM
lF7l5MnpANkxlns6/bDOMqDCJrvuDtvaStP5XNWEkarwGHsPuNx9eJj/9+6vYSfl
DIbGDGsGeaz3Tjulujb+6Wm8EbxtgjxM8lzMIiNlWBZaF7pKPgaWPKEARONYmORw
43C04HNkPmdm+UH5t0VGm1ftwbCdVlxtMPNzTOdj/sucKXfuWPSBDCe+sXHxstnU
KR1eVsp8N54lwvDsEJQZUly7h7aFH/w4BBKqWQU7AfzLseT7DNozHr2zijnr4wQT
0Ry08HOH2a6wGPqDflHgZomn41e3CaJoE6e+7Gcx8iqVt/KuD78DvoaLqBZtJTl7
04oaVEc6oLEOXf7YxVzDEwxKhnPDu72ZYnUI+3RhmNRHhAI55Xwt0NSDlM8RH1/A
Y8BwTDsDu+mwY+U5Dw+1Z/jBK93nG6dtproULuRB0eXcrqqg2hLAv8Mb+I7XU7I6
9xzuFrFKc39kcBuTuswxtNxL606esZslOqdV41AjGFeYMnMkiGgZUpE6yaaYw8W+
oozsoWKiQjaYUBm5zN4MSgOTNs/P8ew+GL3fR+PH+2SY2PFJHeaqhjsreq44WBKk
i5svRDX5UgRVW4n5AXeFv8q93DSK5gziZRiiR+exHX38jIXqCpwcI4yv+JyRtkzc
g4ss3YQGEQdjfgYhFBoH3eywQ5IEhN9NFyZE10J2yl8HZFfTOFzYzKBfh/TG6rP2
Wl2ipTsb9wm0CTmWWEGgexAveqSyUfIRYRO50uBQfobnjqVxFXjXYxMrAzwXbEhK
V85NfvhVYrQGqyfN9YoQ/0UigYizsYUc2vxg4MTYWR1HPq/1jNuHOm4rVpFuX2+J
1L4HAtjWDVrfMIKRXvuFlvwBQHlsck1X20wOwG+UjdbMdrYx1YZvsIWTozRRGq/o
j/gsPbLrPBC7gPrnRtuo04ATEIQVhPA1MWl7o45d1SpMzLKyXFpPNbvX6E+u6pgE
cras/XZMcjP6xSPFg2bndTQTrJEXCJzXOOMO0TTwAUW5sOKlIHeK/eBQmn/AfjoP
05jg3DMWlYEOwonQuzrsRL6ti2OJJidlirC3Gh0+rveRCoTzmEXZzM8lOYfAMyzh
LgoxIXEinu1zd48OygP5UWcAUM+X0wr4avLuK+G42IQRGADe7T0S3lRoZximJ4i4
bnr9IMNQZhSfjyUy2nOFh7ecTHCE7OXjFAbeoa9JfcbL930qn3wjZUdoBCsoXC31
MNn0fcKE7vOrur88evs05IdRRWZoGB9oQks1Y7uHPqqCh5ozfnTz7QpkxELuVyth
Sw0ua/j9cf4WvDlUkv54/COv9QqEqlmSnhTeeIJQCQJK5IH66IeTzksGCL4sAezy
UuKS3QGE2IwO3rWRbSzpDk+CrmtIkusjnBuGktmOR6DukMC8ClW5064gVnPeMfCJ
ivJYRe8N+EFfqfeViEi7DT1ENq3xa6m6iCa7GMxZJL6LNIN135LFhNYUnA774ifS
LSsf2z3xA5Csqy8IswQmKS4gqxT9y+7Vtm0fBAdhl8i/yv4bwyfAHALhwIMsrB3/
gV1GQwQ6wGnRFcU6wjFEktp2GFuNolhF3CQIA3xgA3XHYtxSpFTLrxnlM62F6DLM
tCvwKIhvEPC7UCpBTXU8KcK9Usdc879PM3afVkGCdsRBQ6x3iqlMe1cFjkthDpVA
6h2QUzcBJhZVmXg5IaCF+wlN4FYv+a08/2uqoZDLFeVREo7XAfyXixliT/5s8l8H
8RmUINCeHfpfGRDzUxTijFpQa1bABoPqHqPp8jmkXNL7Wjo+SkOPkszXo7meYegS
MR7/AdPrTPEOaGgj4u/QiKE/1C9Nm124UmXkUbS0nv1a380tRj6GmQJzl0DJ2MF5
qDX1zhAJ3I3A2AeyCXelGrX5GqMw1qaEZ0ShfMbM6taPdSb8iN7/iqffCh+MmyZz
NUdo3WiJrUeNLDivAtxl/G7zN/6ijud2cjoIdh/y9CCgQRKRmLAzXbL1jIpILFAh
fAuydB+bTuKvJurWzbHK0jttYx+YCZSQ1tu4NPwZaNFibFr/qy4RK5rqyHgKcaGt
pd3toH/n/BfxFJh4ywbFdm5jSt037oZ7bUNUv/I2FYRSzx+BTIfqFiku313GFqa9
l3d97mZ/RbFhNaabC/07iv8J+XwhB08wQf2U3ui0ZER1bITlEA7wyxD0i2HUisxK
LUWhkvauloAS/aiclfT1gfwKUtM0WkAurZHKk9+e6WEOY75V9fVti3Cp2b8IvCwR
2/72SZDrjlCx99TBBYhnDE/bsN6XwUkcbYwhea7FhrsEvo5DnLLSSrAhCGabIKbF
s5EJK4iP1BuBtPyB+N1dhqAZABLvkoelHW4V/MUJvRWjr025nIrZRr2ihoJCz3ir
2rbYzETYmrRB4tt6kkxspzl7FNzZlbEE/1wkhz+U6DUDvWH8PbY4c80GYyFesQd9
aOrJRhgNO2MwPy/CsDnMKqNlIHCltAGrAHmXG1PMaMUu2MfWTVRlagbPKOoTiHJ0
8mfg33/ZrRJoHVr62vsSQoWXW47eved3AwosQKaQ534Midzc28+Uh63QxWc2wafz
cFiTTJLmQle2IQhSsogfna/KKsTNBVahi+b74dNBP8Y4tB2cy0lRJq6ybGyH0UFa
KLM0OhF3OEDVos6zoHaVemvcLYPt1fFEYylO3NOdcTQe/MPV3Kdurk+6R/TuLVG/
VF+EbyjOGTeUwKvaJGSH8rnpccAnRWfiydS90CJ6w6HEUpLvxRz7pfCj2D2Pfhyo
KOko1U4KNcncZeZst+EdYBpWGZt0Ko2Lo1ishoOxxYjNSxHxZOHuoTW8yGJSNRVm
ImYCGJqdKs6YssL1gvIypSU1ShksdqNJ5RkzIDCtR7EvnUlZBkfxFpOp+dYdovG5
ifR8zEdUM+rIBV8vzOQBsf0aF0sOJ/mhXvlxarCFnrqpcNJxcPrerMtNVlwf0MVE
lqQwiTLLYtTq8QRE0/s5VXUUDgJv6snjTC8Zd5vunPcSs16YJqbQRWA9fm77tVFP
vmfJyCT7FPYQ0EKZuhedMxwfU2e6LwpPRxP6O5xHSOtcPt6iTI7+Kgvz/rFk79xc
rxSoPIEGES2E4V6wBDLs7rdlBgrXsc/XL6A3yh3FKkP4NjTxCdxwtCvv6kwfgo0P
MjszNPFmIWV/6AXrWE2dcyT5sYsXXD0EF5fFOUO53KU+n/h/IDGxd4I2AMfYxj0W
UXc+g+58vKZQQ8g0Nb2avpGYmGN51LW3536CPtU3n5hiSZVhKf2YF5/Rf+0L38A5
3xzUWzghrhW7THWFcyyCqgMRKz5eEY8326xkZE9459QG47YJleT+YhJOoL0rgoPp
B1rnma+FACRCYPnzKNVlbkKqZZEZiteV4Qr87HZvEHTcvAA+iB6JBwZRBx3Y2Yxo
eXwRPX1OKf30OAlCNrvmij92P1KyXgjHGxd/RZHFCr90aLFb12ldJY64NI74JY3f
zqTWua3M7VQue1MZsg0I+ZH5zq+/SyMZqWTFVPoyQ/QH8LFDcONOidHLRV1Ue5ob
uNRWtgcAeXLOfswj+jlrPi9hzAfDR7QkvDSbmaetGloNoEaSHvgR5VBqBC+grkiG
kq0KVygUobuVTOsmYf64E7fdWt0uXhOTslkzGj0YUNuKKcTlw8XDpl0IdgYs2mnF
+U4p6GL2HmygxHxgKT91bvYIM6XLKHE6B0ovtnN1lay/ndlwA/Qcfp8xH94teMiB
4acqZb3PBJBk5xVtO5iWx8qF8/uRYVsdlZXv9hdTb5sDXShnJIbtDcSHfD++7Uj+
/RLbbBUCZc5qWU/WveKcWoaWNq6JxpYmxH8gMsMJoiw4KsdrsxhTrLRm6gVe6n4v
eKTelfAxBuipbntnhZUBe6ZCyFpxBmeg38w70b1Y2Ii9Op+vIGDPVA0DcUQYH4Ct
HJ5BlGcHybE9BEyIRHWPFP3fTSCUrnWvrFvGMOTkau4zG8fXF8sS6b4Su8GB7883
BoJ+JTZWGwuIeNkqgR1QNCqi8z5tPKazYywymM8N/fYRf1fgHVk5caLItUCYckbD
sCMt8acgC9XNlUxbqJfpRxtlWcseRdMKg073UKhBYjfOwdvRe8gYuaS56iOrbZMU
VUiESH5yKoBlnh3+B7KSKGqzUW3AR5WANrGx8WIY5xxD450JeTD8dl09yXEih8pu
23CdkbcCqdNMaLspIvJuMTalTbkG6gkMLdobPX+WS9cGu9ISbOzf36OvrCk4dMeD
8BeMgQUPhhTOkfFW/PvNU+XxjcDRxO+Cf/nCZ4FpmM/Ll8pQ4Hy6tlMcoWtE8jyA
C6V6cB3qaxGeCtq8IJuFk2536w4oF/zM/pRTpoygW0TH8WQfbpThoz04LS6Be8AZ
Pd9cLCEaRPQ73B7GMMcYBaSFqVi2o3wAYq+yTKeAlULYZv9GcaiFvJBakG0iSm2+
NSYVRS8hOu8O8cJ7FU8KnVGFSmsLJmMo8/2/f06pQnQXykxFX/sRgmhL4/Zkkmoi
0QITlrIcyTosf8s/avk7vMzHKAdrqGh44YhZunHtJ18MJ/cFpsKlm2yRFXi7wIXh
gjTtwLpqJLM9XMlfNluEymH7sL8+/R+KfYJj+tGRxvjCbTnYRQiVfOfXgzYKlHhi
qCyf8izHYgJnZhxX9Ge+TxCY5xX5Vba6kyQmHd8Z9tb6p9Ju5U0W2qffpLrSCCL8
F0IcgdIsVt6qpUJPkSb2rB8TAR1hbxFxNAFG9wTdPwzAludH+bNQYw+HMyZN2Zvd
L3mT6o2E1ewU5wxHhRW0N25wjmQzUuN5+OOM/0GlVFg/QwcSLk25BvgGCpLJBIls
AoZMSDrrq9wDEU5O2l8gipjzPm0OyYUmLhKDDD+Tt9TyekOA/8FAHM9KE8tnQd3i
jswhYAHICRoo7YfQ/2tch/cl8TH5XWX8fAR+2nWt7AzlnFlO8wDN2fSocP2jTXP3
fT1EH88o9jJPcZIzDbQEOqvzurvwxLNMih2vQEZcEXkusjKYZDpkSvvIABojGgn6
CgRMCVlpzEKHm4Sl/hb8VZ3Vf6BJ0qFFMlznKX6j40V7vsrBPr1nF0G1FE4SdJ1W
5A7U1p1S36ZkmoAS47sqhWwjFVlnp4UzOOUpplvZm+O7S3Apie/WXtREnNEnbC/X
0YqMZN7jpPx/Qmrz+7T/aCVMuS8An3uobuCE0QKCGzqkGvSHcdWsczDq3NtF1PxS
QC99b+3dSFRSv0fgOMXDQyARSWIrjXVuPAT57NnwCQISxOE4Sm7QO+3Q1GNdzS/n
fWn3Q3AAdliMbwUleqKJa70u2zFTbTx+CyK5c/hSHwnTvaYfzqEzkY6Ct3KOud6s
ozbkFMmnOxwDVmduol/0PzJ5or0+5ZDw4gtHKFTkjCZQhGrn9N7Kd7K5gBkTQSC0
4ZIHHe5KpWBlldtgozqS0MFm+9LexagFvTUx02RvwrRZOH3fmsqrxrGiQoxn1BCI
BhqpKlstJ4bMY1AmGKqXWKbjAfYAITYghcB35bJF9sZCeaqsmubbJJQxj8Bv58G6
mL8MsZLthPqK0QNSZcjarC/JyPvD7rKtAzfwkQyeWXY+3QHjukshScSTXLR7wS19
A16r5anHpqN/6CVrBoWbYoF2+tqtzOH+xp8IUTZr1iV3RswfLhzJu/1EcmNLpcyX
o2HT7f/B3cEIlCaZ6lJD4NqRhcQoLv4mxBJgw7BlzkFG5eEHAdkgV9yXWh1kAuIQ
qDG0oTl1/9Bu56NxTfPw8VHWhpK1tDN7s3q3PsyO/vHJYg0B7SGQhzPoSdeZmGm7
VItu7Q4361i4kty/b72FbCL7RMJFSgWEF7V4oBkcj0QvuTzXwWeaWe1w/nfDd/Dm
tKYAH9WmeAAAthOJkhqIXwoDR6v2WdcYjPcir1XspNUZtga5dpDpW2yZGpMLcm6+
LJ3wxXd3TrLkv98bkpszswpumVZI9jeUSR9NQWMrv37wlzmqtF0U051HVkAWQnyS
9qjH+AeohhQYK+RAaGb5Z0WFp1CXxKZsYg7Eh1gAEwXUR1bZ42fs6HaAgHoM1Npg
31+MPII2wV79EFRlC57GHsumV7Ar/tkEM89YzHyHqgUVRbXE2N30zd8uiBroRvSL
WEjVTeEQ8oa9AUxJYUt27X3hCqrJEbUMwogQTka+VaAjcWzascw/fNFQciNM49Zy
Hf28MvDGA+roMIhDxRnRxalnQlHLK1Yuc0SGlgS/TtG1VS7RlKpAu0xUWu5noMol
uHkgL0PIlAxMYQs/RdSVtPie7mhpbAZXtCPJX/swWwYUwYoLFEZ0L++LK0QG803d
pMCS9W9nRFsVaTvEQnGO4YdsG/g9+Dbsa67hz+qDps6iByFeuPFo2gia3YzyytmB
oKo3y5naRWAN1QZehVEd8f7Mgg7ya3gF2LARql9fHal9qm6jxSRnLfIsN1OwcOqM
kzm6VSx/EtDoKeRoiPZ/uzSXO0mcdGN3p7QNWV9NkSnIC/LbsKJlsYRuOYkEsNUN
buijmfU0r5wzUblo+dKjGSRz18w5i3Cp2P/PtesLaf31iMBjLWM3AimaKcSiER7L
t7rkGn+5rKp3g5R8kit5iyODIeF4Rf7sxqust1Q+Cods8dvNngc2TeBLEbGIYt3K
I33Brmn3IAHoWd2ClADn1yMv+YbD934+AukupSCx8EHVR8fM6kRuyXwFd85HxHW+
DGmS4Xfew/jtwcjnUZJdbkr8nValQGlbRnZxyZhcW0vAHIZ4kZMUt3sDj7lb8tRm
RpVHBeOdSMVmJ8kufUaW2GUWCB+F1CoaoNmYgsXzxGPEOB9+MVXJ+Y6BGG8FU4dn
ycXcNoKTC55I6YKao7037nNWdWE5FDdOqG5quy3VBb3DZEVPJ0SQr13ZN0uVLPF/
aIgLsWhZkAxE4rf/HiYG5yEfxGbNpHM6jsJsOFxoCBQ59QGOheAlwds+tZ/fOFnZ
bzXsJrpQH4++lgntx2kLcklD12x2ysTr3HLDqYTGRGe2psLuOBeOinSOee7WUWO8
UTNM0qHgYxma8L/hPYRX7q7szg/aqItJa+hEjiRtnhWcb4k5x8tifugQv6RrKsL6
RFN0S2G7GCH6txHG4BGipLgNYCyQRL2DmKnUuBqOz9I20hCCCMnFMarNasjH7VBj
Tz28GO06t6qidw/zvPfJIqRA2vZ7NPmZanH2v/hZu2nlV7pgq8hy0druXd5jLVR8
3QH5jvCVwH4myXMFgfYJwfk/eD1ZLpTxAxa0DZdnVK4zkkb3KhauOyi4lDAyAuRc
O/4UTZqF3bSXttrBG7Rmt0Yd5LIwEYmwK8aO3CqInXxj6lel4OlvRMvU4LubAnnC
Jbv23bBsn65Tz4lLY1TAm8qqCbMl/Au1YnBKhv3+pxgSEKZ7GhxW3dEP5JrkcxoU
Mx/vUTwuf0xBDM5tOooDgb12RS/su0u93t3PYepLwyEL2ADOX/mVD9nwEBEwgf+O
DPlRdREOSiiwaaWQegGv3/GpN+ptBmJvCplLUOGE5XRnn0n8lLkicHxTSZxeotK6
qgISFtvDZSqG8jVUtiVtzTvdVvFsxVO0jlDH4qgaG4a9NRJ/25d7PMnNtgXJm9Pw
UWthrodfEFBs4YrVr79bo7FEWmzyDtWTkorX9TMxh1rQevuqEiCh5SGOtMs1IMa3
MOSgJeogQMzHV33eNPBVCM/z5QIMfVvn8ZtPOMYydx30LfvSU2j9XI8mJYt17d88
R+JQPVNP+74ySuAf4APyDM7/rBnKNp82hNFRFekVUNi5K7LuW52tHMxoSP18gKT3
RwBDu5bDt4Qd2swPWAtKmv7bMCpmtyQHfaYRzRtjvnUxYBUi52P4PR8UB0czDuNy
e4EQSxJwDVK36hnu/BYf8lWcGzR2DGmo8XwVvmcNytaqhuVUbk5VI3hc6PXUm1wj
5YEieWcEWqM5oLaOolkQaQ9cf/B57ONm5OajEVJfcbQy3Z0w62fY07ZPLPMntzqf
oXvFdX8Xadv8kiPyau6QBFcf0eG8bLmXUqaMbnzqVHsITvSfj7wDs1JNOmNXH0MV
WfrtaUBNKCS09IcGdx/CH384JDu0iHA26L2mAXrRpEFrVyTsH4vzeESXjzK+NFzZ
BEjxO/jcB6dGPnyjHtg2W8N7LJCrCtHkviT6CbvRmOT6ZcgXyldXEsD6aHlE4z9B
PxaQH/fIOyaAuPqdQU1nnLQ+DSkYssN95KDg2CPYnaYYPmOfE7C5a7ihUEqSBYfm
VZ740M8nb27IdySgjVTMuokQxgIjkeYCNwhJd4AwAOVGeUxJhwBsdFQS+1bO6Ujv
Bn+X+72SI2SNqMha7PSG7ZHNCUl9uCC0ZmQIJyC4y4cIaEovVoPnVi6w7rETyKCO
Q/ULbbbCCSBTcCHJ7VbBffZARxHOqHoty78llchVC5KKmlRfJciGMRDZ8OWDrTPI
EECzpkLuw0VRI+t4w8v4u+8BRJl7+dkAdlreTY1GdWgphoKOwVwgxdyI/TjvJX2g
jBkGwl5mXDeL+WbFhwQMc1rPM5ifdUCG1pS0UQ9hoD4u3yzmx544uXEhdmu+P7D/
AbiYCapQsGrRd/iLQi4+6krMOwzt1gfPabUeFRMnAA8cgix1MEsilvWZh7W7dW3V
M1Q9cMW3N5debQ6hgq+h+fmaTtGtskTedztAIydTlZ49gvPTUa4IPfALnSP1eFwW
wksfJs8qgT2kTLoodN7QfYO+3pVnsmZ1zdzUrE3WDMIoQKpPPB3Sxy+O+Jmgm43k
QAPaW7aPczQk6QwnM4zIcqMBkxLE1Z2YU76KvuxttC1DbledWvgQTxVlQaM7RQPl
DNaPOTV5TzhFNxHAYU6V9lOQDJ1kxSgg6lzdBfEc9HBhIm/jYfv5FSxxujlUJRcl
pkl1uugdRpEDXR+zG3xgX2pqW/LGFuxKVk2nw9obRkwPWeOthTUyYh4Us4lC2NWK
x/h6AiWPFQfJJvJ1ByKtNwlCe4lt1op3e9tbfsUj7TPdnr6tBG6mb36ANQE/Dv5n
PaRS4HJ5egmLwcbLINyBX3bh/2udYqOJaghkRjxaeI6ntqZVeIBz8VJGAd59AZjM
QdZ1h3CoN6ZomJfI2u66vVqwZ5tdmbXSPeYsPrJ5N9tpOVSikkcoqzaU9N8cfsdr
vP9rtQK+Xtx6PnBKXe6qbMKUGu+1EhMj7vZJLbikLaDXd/C+qv2LICcXNGuAee19
ywSq+KcLnFM/uihUY5MgVF7uncu6gA4/mvO2tvw+UJ4XDhTY6C6JftOtSd/0ZAN9
1ZkNBDgkMwYVn9AD7l4h1cMOO4r1HILkXglF61Nymx8YAU0cXYEtDh4BZuAx1XZk
RI7V7ik3MjaYt6R/FB0UsFroHSYrJrFHEm2cjLDqB4G5FGOuSy1CLoyJR3KDM2Vl
kOt2SKh/C8DmeOWs7jwqbsPY8rCc8ZSPM3y/x4074c4x940JqHntHSRTkd8sX54s
GqjjYBhi5mMya8vQyQbizT4MEVp8W6IZdd9xX/ED0XHxDr4WZWUelhcZK+D48YWa
H64vOzNjRQUgO+Fx3dMgdhaLvgO0mgeV1y5qFX5K4QwDysvYrj8fDx85slehyPI9
9byfwOHp4gExLLsiaCv6VmmoPZV08cL+WkARkzxbwKH9b7nr/xU14fgEmaaxlL98
/HuCk3lHjtrBdLZM8nNbDYkV/Dtay1I1z1yvwhNqz2wgyFRzAASUwfPgRJ+Oam8x
h8+TEWJkh8D0lmiYdG9FsDBxk0hIYcDfmgDGPB9S6L0cImFNm52TgJrNnpYRSZ3j
9Ukd5yi+T5E3FIM1dOUt+IrnFuUmnpvZrS/YA2wWj/FnKWhqyFc/6HfDYW1huHEM
RRmCp5IER2qB5zZhIOJYGXeZkdh/ErWCdXR42fL+Tz+DQX/JYpVSv46RbOkda85p
I+tm7gtrs9wZiyj834M3O/Gaj2BobRPU/IZQbeRJUIEzn6wD+Dotfuwzm+vzGp+t
uDuUQzk8Ps/Txw7ieDx+yJUf7PQMqfc7Bo0cjGWkVrNzK8pSJuxH64ioTtSGlTYi
09nZ0fW2Jc/QyMCSnpkO9BfvbI+QSM8td788x4gwj/RJTkt81q68Mi3TJXKbR4aX
wiRLcUbDluo5EZf1iJRgvQ3IfbNvG1JL1CevCrhzfiWOk6A8yMLShVBlGZMr+H9m
PexcPt6WVQyGgfI6w5TeYIvS79JQe/xTMCKTtNE1A5OUBKBIfyYH2CJF+tqLEBM+
1/QFmkxGqpT5S3DG9TJNK4hmalXnhl7b3UYFJ0b3LsZ5T6OkWoOTbMnfxmh8uZJ7
76l6qIKEtfl4ftb96GJSUd27Z5CtTnLzhow2apPo83iWqxC8+sk2LrWhf5918cLK
OcSjPCZADSiby2H5MlbosfKx9HoRQFies9+dTGWv1oGOtfxX7hLoIj297oGuzmZu
ooBrLwnkHgHVMiB69DeuXqHdbQ1DFd8WH5e6yhi/2+5X5l9k7nHlfvwvEjuCjsqJ
rA9u/Nn1V59g13aUytSQ2uwhKVcJdACCNoTeteD1vC1Jb4giyj09WsIRZHNwpbSq
CJva45ZwUUr5CDuLSjk1VUaqs+nPKMsK8SpiA+DjkpsU5Ppq7NsgrMNIpdg6GPAm
M48c0RXBjub0H1IOVNmsSFg9jZe1u3qAw+I8loTZRXMP14mlTeCOqtPYcqx1yzYo
TAJc7K7xOi2QJLGAxDmvzSWRo8hyAKAsIQfIoV6Mz0aQtvyQANOnhdvVNru1Lpxp
qM+Z3Xrwqlskknehkgpr9TKFpGnSfdt4p4BK1+DZTCVUMgw0KnUzKbblIxFxkaDO
UttsT4Op6Xj4qEnUYn4yDYFpwgFKyf1cIBHCEEPA12MCkTuKaDp8Y47dz5GlXYg/
GS+W+EMzmrlluo5kbC5CoavXDsW2Pa7ZzMWcDJQ1jwkMUhGhlLazSjSPxJIcU0hA
xuuKezd9xMpWDApYHVIi52u8DHgfOYkkekcfT8GhBR5hpqyZ6uTjU9TcaHOtgCM+
0oT4s0GsBTE4i88Yh/bvz4rMpKuiGdrQvhWPZYLWLxcwEtK0yQbTe5d7TJZTyKrF
qAHxZQMWZ5DxqALGSssirnL3rrVJMXPnDoCGOO9gQeKOcd81PBRmIG5milJhcxbS
ExJO7B1fRr06ykMgu11MW5qUWbK+FIMEz+fGN02x0QUFvq+F3XmF4DNBSL6FiY88
tffmwm5K2ZWgR5OT1Moy12/DC0+nk5y4wcYpRmR4CuLJeH3cX3vzkeepQyPFq1g2
0PbxfezN0MASdnGrAo8Zj3Pagx2iLb28k+Xe0pKqBXnpsiztpDOLrq1maOS3I4RR
K9CGSwiGxCO5aqgwyzKoZhiG10FuYOYcMwo4bHNFrW5TyaWqh8sZI5mWMyZxu6TN
HgHLOzpBVgfNiQWUJu5OGYTKnq4v0Yzq//igi/p/fEt/D0DC4juU9sONJari6hnr
47AqpDMzPaGe/GbffwWuBOHRb1aa68mF2tPQ3FFUg9LI99+M/Jil/udl0MOsC03G
fnTv+oSFJlM6yBCUC2N/xbltaOmpjD804fuUSgOgMzHDu9lyzIGBPuO3GFqE1WNp
bnQzXxIaszRbV6OVlaqWVHNe7sSnfNlsHnApBuNPY9C7pUk/l8NFMGdALSzf1Lr1
5VE8cldxQUPjUO8mHKpfNyM1RRO/ayX10yJSWPRsoXIKayoGozJmFCMfrtWGBFJ5
NbBJLIR7RU3rlZnpnaO2WuKxXeSk5gaKlK/KHMaxa0Dk9t2A+nO0k6UhXQekuRSy
+YGP2DcIezYqypiXgQhJKGIPNGoOXcLxNf0feFrxasz9BsVH0bXzwu2eXi3IEs49
DIOOKvvOQWWJQgnsMTc3FECvqtmUzZfaNtmaz4+fdA51L1dMTgItkX+q+uO420J5
aUEGe0evhYDvBOvZRf74ufFzCifQ2AZ8Nf0K1MUXNVpQACRcdKGX8o1lP2hxvK+n
F3Bd9n7XqZ7zSQtyVNacSBGSBQXzcNdizIh/uk3DG8Q1xRGXtUo6iW2Wm5wEqptj
Wgbd7ah7lbgT6TKCcD9TrPpdaercArIeyD8yRjNKOkM2AVMdBpUaW4tQFRFr3lIq
xC+PFYidMNF2NrmyhewDI908mUPlT4C3+unt928gLmVFypT+GVuAINDJGMNBpBk/
ttSuPhbByWwB0KLydxl+uEer7caOLVCKHxsLKkhcxX2vSjPBgLOHcaAxW2/aSQCo
SysLCzaNAk3ea2X76V4KR/fCDINEEtUdWfW08130/l1zGmHIfa9tnXObMBifGUHt
BMV1uqaMprUtSK2LPtz5HPBVZ7lEAem4MUr+K5L88G/GhiqpGqXRqjsVagDD9FNa
CoMvgktydGYPvoNi3P/WIS01YSfMmiu8prT+VUD1DUsm1fswgCKb9Y43+byZudVX
ng33+YDl9nHnaOE80xO5FpAcO1kqVWbomn2PaSet5Z5k7P1JxDAyZpHtmBiDZwkB
3S8ADQYo7jpaCltlVIEjTi1dgy0UJivP9JC+98KpLHHmDcf/26Qmil5YIqxZiOh0
zDWkclDLD3SJrV7dFod9+m2YvkvOIXpJve+B5rL9AqtYNMB8hOUqZ7fk+prAgdCe
ZbzR83o7YxN1ttONEwOeG0cl8E5Mj450NnQSLhobxpOgS5bebUXqvjO4G5xhsSUm
E/M9iaFrfmJrSk69HbZjzaX4gLWJxKWk9WhWPsk+XRWoWU8b4K9klcOjPBPAWCI4
DgjGBkLgWkZnemZaf4tpMmO9mbVMAh+6aGOz+Z/2sF80ZbwxNjDnf/Kh5Hu8qAgs
7ytEhwskoaLVTMOcDLng+mFoFyX2kD20IBVs56pieWZyFvn9jBl+7R2oUIOgUgRJ
EAWVU13q9T3o+DR6Lz/7BzdAtTqnSYbdTtso5dDPuL8PCh5wFajx/2ISxaswhSby
68q0Wr56tEoNQi/WoWj8d29mSHOGF+J3yFiaw0Zn0FcW71dQfaFw6px3D12llYKI
vxZHp+y8JZ3E9zxQmQ/OgCBlvp0BjSTZCC8CPk1qVkS7hsGmK1AkgF5FFN7Y4oWJ
drtgmR05TE2UvIaMRbYz4/JtUlyJzsA1SknYiojxFzChSsboHhF6MtvzsWQsqyBG
Gcd43SDMzMQxI8XC2Ht3BfMd3AZP4pFDNwXNKsaxImxT8HdWjCztL/ePIqGBg7e4
XqZ/1sq5Zzj09gs+atvB33En3XHLNQLgSYjb5yXQxDWGxzilbhPH/7tjLD/JDfZH
AROUezZ6F5PseOZTA8so/+hb+h0E1/2c0ZHK3jgTWDjwCys7KHHevDZPPzkbAPV6
Zz/PKHJYp5xJ/jp0R/EiZqpxnD5pu4LPsNLWcXZ1SRn+nVzQydqY/sfuOsVt2Tjg
0DsnjPlrIkEz1eicl2w4mGrkK3Zv3oPX4FfTerExaGnLkL6+/lrCWqi2t3npGXPk
9SJvgnGHHOAVKpvYifv3tXlh7oVl2zYub12ohm+cILNcHs7BZ5hzRMilQfh7uBPb
Pe8z5Q6ovDb3GhTl5TrbYO4TCDxksZWKTeMYl3Jgk4ZFp7GOLrBIOaMoPRky8yjb
Y12/HoAoI3LqkG9mUWOAFU1UIxaX6nbVMEkSwGCn0wEurIirQuI4n62j9IvyD4w7
pj5W23jhLpz+ChjKc8/er5DGuoin8zhPOh8mq87FDVuymYJEjf5nKT6rjpDh9Q61
viR/I8QFCr/hBUgqFo6GgjEvHEYELDqE7/cHhE6L1ysrqEkGscNX19IowHOelWsF
GbS7NxXlE9rVUoFssLpguw2xFIIvYqHmZGRxXnhh3Ip66v3zbk49IgkB5bk4JS7B
YeSTaI/kX4QDlpxnAY7Dzyiemm8s/dIs5RI9/FyrNjT9FowFxbRdKgiQv4aAmjOC
rv5XyRK6Pr67NJudt3ib8eMyOXG7O6FY8j/Ft2HV1zWrTBwnJPWkDBapN/WI2hoM
6O6OXadu/q9+7AKvSpgevKuKUKjg3xa4ADiysYu11aMalh5zLFUKoqOurp02yXHc
71a9FVVz9b+NbLr1s06M62hc/oW5umxdW1CGploKLJzOjpCl7kB89LDfYyd18Pfi
FfqZVx5GoljZbPV0S5j/vYqcrtcLhbm8osovTb40vdbfVFzspKtq3qvTkHlDdfIq
Bj/mQuvZVFMhKibhQBJKXgut9aTQtONP6grKh7yeCw2dkELecXvXODMIEl0mpReV
2Nk4EAKghtBoadtS3frwRb4FDsjQsBqXyMye+rsZuULtcA9i00vLPuLeVCdSz21w
ELZ/AoYyGX87u4oao/AlhO+Zi35YcDZx5mpjzQBUw2ygsL8PFy5pAF02y7M8FK3y
kuvibKw70gLY48cZ9m0QfoLF1GeuiCfuE/hps+wowL6PM3rrsEIl6vLiJb+1E+D6
hMz4rYUTB7c4gwpF3q8JRjONOUya2M5AKvomPORvLP0v2c3uvniZ0uxgBtRgjZT+
Ap+wYeQpEEG7xzmowPwXy2G7wefooMyWXF/+oojsvlXxKkLsrhZ186Yr0+HxoXbp
SrzBPlY1+dRxqAgIWWHAMQhG/1XhFzrARrgCQHXKqnYoSNZqwREjIF1uSP8nXHeV
sEvmKCt73btJo9h2zSKt5f6d64TB8AfbOQLXN28zVpAhR394xJTA49lNSSBDRISa
kFKHKmrW8lgJOWp9Gz9MtSNMN8jGScufEt1WjkotpGXASY+QHgC7xrkOzSiAAcvt
TCmFN3IYoZDWjAByulOwNr9Orr6nWiXX3CuvF3ofPCQd9M+OtVMYx2HqWi975otO
GS+rVR0i5ly6ZFnQBM+Bay6HgWRNJZnPENgLi++2LEoyNPVdnh0m8H6+3IhWZUqX
6PP1aVhQc7bgSJItPJpvWiA1Mz6D8Eh1zlYaHwH7o+een4KUM/fp3OYaI1XIP17/
ku0sI8yERE1JKDTBv8gz3ToXa5VMbr9NVX4F4MXyflo7z18g02fHzE4EO6Jc17Wi
5bJ2/LoW/5PkMWNvP4d/NKgmTcF45qu/Vur7m0yGPEynO/VGxJyxXqoXVVsaupoD
eA5sI9WkAuY7Oab2SMTAfoKt3Xt/sjt7U1WFuGZ7ga7UzhVWuOXW0jya/ovC8DMT
/LkLlBBZuM7xDQHqIkYfLIw0nLfQj4/dJPPXv7jgKGQ9vtZ3dxkOPi5ML+Bz3JjG
yAYAe3PiziFZlRrs+iE507lmSx7jcKXC5cbpphcV+QIS55kno96NFK3BQFgw+GSH
t6xv8QGem/yVvgJxgyHTyySam82pRoMxT8sky4wr3ZPjZ+Ee4+GqNrGO7R+KwzF0
a7IqQZ7+ZOjbS1zU75iT3mLOTpV1heoMmm46bAcfiVxfiooKz5yc45nzFkSu3g6Z
BMvFk7e3gJIUUXD+ficzXwYeJ6m7iFli4pDM6I4BKxZo9WSKauFYf31jqmsLwEYx
tEwErRgFLSBrGdX3VIscrb7E/GvT8owbG2wDIRUOWReENI0d3tSbdT+rEab7Fr+O
fF/te1YACSjcn7FUPD+uQ+f25MvfZB0wpzrdheJKydFcKD9A2vX91/zJ/6rI85CC
tZDELpSw+H3ZKH5g4HiX838kBSUqK9VMDIcsRw4pz16jkMLUgVp05Qfu4tQZLHpu
uA48rm/sZzY5F5cTD7W2+yO3w8PI+G993q5AHwPWi3lGP+/1nvWh98KQO1eZeOlZ
h3ZbgyU5jyg90u3mfvzbbyBtoIkBuQqj3f6RHD1AhFFpQnRiHK6g0uCZnOacdkLq
fW4JCW0sRFw75Zp7aYY9Ce1ivYF6T30Wz7kK33BVs2keNqVtqntRX92WHO+hhxrg
mGfVuwX3T0yT3fd4hViOIc0PCGORlz5tp0tjIYsl2jreZ+1wJblyKnhYpPe89wiu
rmmtHEsW5ArZPeWgebPDutiizPEjJ+gzR8sGzoOBXI1gzeHOx6r8YIefueqy3q8W
34GObu5Qpmj28a9HeaGkPJkb0yQIbkOWUhJGCoxZjseiUuYnOYf7I/P/mJJQ7yDn
9VJd2CHChXAvnC1aAzm3lUtPX43cBBeeBC/DRzOghEDLdsvv8AGUFflQGEVyyXnE
IG97Uo/FyDR/RCfYRuXaMQU2ClnN7w2wz4Y5Yj8xuREDCAiCPP6TuquBUEGQc9H2
lLwcwpVyvCB5MgQBlkJN64kIUF51tqi0toKU/5ueXY9zFEbpiaEfiSQtrKmninNm
izwYgtC8rMV7BhIw8fD4rJ0FLLT/5DTQLq1lkHo8SPvNiuHdiik/w061KiDpxS0v
ekDk2fiW/bKHEdOO+db7kSlFxYikVukJ5xgNcJVjb8M20Zm0+iqchf09Slc0u+W2
YAwPx8Xu4I79mS4Od6w9X/pXj6rS79xFkZLi6qT9RJ1+8glc1yP8mfT9/REzoEuC
AQenAk/b+cwWpfsSgT2tWHGzzLwr3+Ia9CKd3a/3q8xB8Aw8T23PG6G4bCwj17/r
S3dqbhWbLbo1oHZQzI3dhKR0dM2CiL6cTRD6Kao1ExOwlYyP6HKeCUrzsWilNuqR
zjEDM+FhR6z92hqqGrB43B14EpF8nkT8uFh4JAL22Rfow6xu0FP1wyFB7U8Km/dR
Whs4fmeQUT4rXNGzPrrE2aXBGuWB0/uwlF85yEYv4MHn4G7ltGM0M9qXbkninNJ/
ymjrbdKiAyrmu91E8c4PK5wR1Wv+4KJsOcfjQFNHbqkhFV8CxvX3lDOXyulev06L
uR+rW1xes9NlJXcwX+IdbKLuLhFTqQLSWEh8d10uMBGBMIJClke+irbC8PPKPSHI
bjF2n/6q7ixoHwpwioV0Qyl+bAXHyXF8AB/t2pvATSohyeUkQi22w3/lmTrzV5W9
TNklAKPEjg2EPcqJFYFZlqjWkwiRY6/MsjPuNR4c9hxQpOCESIxnmia4+DTQfR6G
eiPC7HRbfxp0jAnZ7jUkbjPIUGXno13F9o9cQQLSBPLgyYzkR6uTtxdOjLNL4ktw
3ineObEmg2JhC0/v2fdVF8NhcWohm+PHfvE9GHRkB/PY7wOcfzlEKX+OumguDM9s
ijVllCa8MZ09lH0wtd06sFMreH9xF0CbXuZlnwepyGH8jV/A272TM+98tN+JQO79
l5pJyr95Fly9oazmSl9Nsjbb56nZgSkozTh/jCCjBa02teCv/HoLG8tLVijH2H2+
29QuuQ3Gp8aec3i8DM+AVoYt0yePtZNvx0ntbPaQh8Xk0JXI097XiYhnjHh382/4
Jfs2N23b0QxqIXEnfVVBYvOOX9lu4Cazp/ta1i78yGngjYrZG0cTnoCQm/CiC3l7
yas/RFSzs6M4flZFcoifoGpL7RlIDDT9VijzFP3cmhcowIGOq1FLgb/3Btez4uas
ieMsW4+jzpiIchTiwrswQXfF/0TBBifeljiAbwh1HwR1YQgAhbYUQIn0ceEboFXH
K2ncz0TiQVl85uHjEvkW+K9Zym8tQ51n39jvI4MI0nYlwvfMmlWhlqvDvX4NfHEs
6JZX9RHCfsRUGQMtYiFSsMnSYqCKHAPmZB1+EswXo81JxWHKMRSoTAiSMFiwIpbf
YnWwoMDWhp9mgdD/16cqPqnqw8hRvxtPZm4wbZVP3/fnG73QRWr164nwy7txZItu
dcVI7MXwmAhK7XMWja/NU5aT63fl8BbD4WX+CCMvc3fUyvsmaTh2TYnUX/9Xm9d4
sUSyxFVBDPlEBJCRuj0WNx1mARmK13c1xSJ0WjvffYv78hMOeB9j3fGS4l2LxOwq
geyyHyn0PjDxH99b8TzscA+B5gRi6qtk5SWPr6P3bc46c0qMZpx4kXDs4hB5UE6D
6gzJpPoHrYcFcvAq/VlKBgQlA8c5qRG28xYTbM+kM8/U5l/iZsjjaR9UjOwrmd0+
Bwr37kPJMeCpTc+k39eYHXU74+hS70DT5TYA5eL2ghMHiUutHP+6kXU+AEiRWbux
Y2pWx2Z15niYqln3nx9YjxNZtrXm6wONgEFjp/jDc3LFu9KmxHBnABTGq9mlbGp7
OQQqjs/NQ2jsF/FbUqdC3wcZqA6kK3OjzlB9l7CnOD4SOKmpekX2+Mi3ENtLtITW
f1ZvmmkmjelUlWIs4xMQAZbnB/YCk1e0KyVA8w4CnAahz7ag1IIDRqz48cReF/J2
uiFEDy2ROftTmGq+cZxmRK+9rMeULrg1lQC7gXgSs62gQXzP+VcfjGImLCqqVmD5
vpjrujWUO/9zsQp/3Zwa2cT8FTw2w9sx26GXSDM3Nb9iXy9tqPpWrFqBmtlUIWJw
Sx0cBYFsL8W3z8kQNRAT0CXz7l56uhXBkyz1f1USK6E7fFX1+aD3hEa4iV/1GFYd
paTdtD9M26WGLGn76m21RjbveGlj1cGeZ574K4cITGejyr1Hs8Nq2ROq/ZXlrB7t
sIVzi/eSW0+WAU0Gs/sUgyLulDcjA+S/QAYNpUrMH67KlsZa/b1Vc1pqIH1NtpTr
+W697ZAo778vSo/XKgQa5MHDBtOOy6SN1ETH8e5wm30syXkGVE4K4Abu4X60DIAh
UyQZn31HEk1/5wX5fkE3G0JLaO2JaZcyo4Fg5koOKV/dmQaVUYhRZ4Izlo1tv/cb
e45ySOuOE16YCB3O9S3JFhMOFRmqnOPuVOSpycfsA2Hv82vAmiVqqyAW0GzbXiGW
nqNIngJ2N0bVrA1zijU6bGKEWq4lMxR2W2+rhHau0HbLr481g/C4FUOsSIYOlHmJ
7TsDxD7+T+AnSpkK9aI3pmSK8NXwe5ZIAQ+01E7LD9r/CkkEWhFULHbTM92PS8O/
B+TTeS/Ay5s6oU/Bjfa1dJgA9Lp6jrVNkMSQrOBVZ7RO6tPcwUeI7PYTYhkhhHfd
tMU4t5LJlifsqSOAkpYF1gZo/U0miSJoOKWg+QcCzFwCaPvFMgUwVTx1NwIcHPdR
EnWArZV6TjT2/2VnO8BtHDdDFpmExZYjSR9hZ5Yr0g0jsJLikjls5WOlbU17hcFr
9N2QA8iuYgmLkfFZaKmfbzsj8iPuGhJx/ZiGNl8UNBLrRweyJ9QnLDey6HMAtUv9
ZnUdbfKt+11A+0Nx5YuCnMUh+Mqd0wTr1Xzqd8huR2Fez/qV1lqTi5xwSgBti0Fb
e/BhftHRgJTY0f71xMRY/sGpTpZVDnvGGYd2xLWblY8hvDhy5uX/fa3LOlTXRiuz
y6yN4QX0GDEBYY1KR2gokslSlN1pxQLM6wkzkrqHddGVLWxvT7wrtApANyQ0wO/9
XK4u740NkQvYsThWzaQlrINwNfe1Reyov9VtRJQ6IxTMD9rz+DR9/pUzBRxVANOB
sDmrnBtv1GTcNs171plBr8zXzg9/engzr4/S+F+ivFfjUKXWQe5XCk1Je5mCKyQP
j6kbIOIzg8kD9sNsmeLUacfiOHWq/WSFwc6P9vJ48Jm1WUqFhNA7VQkqzn3XiKzn
H17IyKPZKecOexMtMvrUtd9RVsTEn5OWvnH8BF5GBX4PyJUgOT/2JYkvJyAgxMCs
G2Tz2U5MD59b6QuKNkFLd6Nzofe+/fPNSuRZulK5DsXx5pOaMislkr9k3eqkv0Zw
b2MlvQNrfvOuAVF5bpnSe8LzLKAHrAWto8A5Z6s5BS7+swCFnJ9wIiIoFfPSvBC2
8kueuWNfGZGijUipxQunIPkDjFtlXJYLHkWzyLgffOeSoH0QYfInIWA38qDX+6Jw
kOTGvUimeapULEuPKsS2czNrGWvoHtvU/HLLDHPJt9pJK1xDg+U79X300SSMQMyp
GcVhOd+VWXbisemwQLi7y1ZKo0pobn3c6mT4zzXyccK5W+h7FrvbajKuCMGEnhv4
E3QT0t54+SryFZAaoOgYZxu4fLxuqby6ubr69uAzZl27wBxXtKwXMJFv3ZLMDpjK
55UAqVzEdnV3hPsuy0WsU+NixSOJXwgDmLOooRF7hbS1Yie6oINeDptm/75b2zU2
1NRSd5lfPRNNnHt0SXb801rjsJtQceuYVMc2izAq8nOE8ore1HefvpPVyoBNWcmL
SsdrScbsu+JR7HphwWhYjTmO47Q8moZCAJUOYDgR2cgowesjCED3DpoVAy/YX/i+
mueiWAh3wLd1K+VsWshEXj35yujMPSLIuoM5COheB9VDkIsFler3hgImnKVadgja
4FetHW3IniNS0QyISBb9kegw0BA3KgjTRIcex+N6MA3Hz/KETvoKKslvS2MNCfPp
EWTNR3N9mPUTnTutVxSLIJUvqwFChAVmQbP88J6JTl2DvMmNVPkQ3A4Y87GXdfDK
u4wHNEtGAB4qR8N6mGDjGQqJyXHGn3eMbrwrAMlt3s/aeh9GQbJIPnsWCvZxb0dF
TafDAh8PiT05WoNQxo6kPerK8QqElZQ96NDnF+rRfeNdEuTxfjeCmLscMVIOQM6l
d9BEte1Vgh9YpKwFcjTsdgOOyJwso+oFiGdJ+Qxu2jvpD13CDYJ25qqIINnRf0Eq
cvnHHtwhEuZU3PFdfFcLbM749wJw1pesthMUAKBO+GpCGZPl18UkCmu1rDxHrUFx
Eb1BOe+pHPgxc47hTL6++b98XoYyHYhRY3StsEnCmM5ZPgHz1GTGWZ6wKf8HOVyt
BCN48d5Dh+moLlWLwAr4CzJzMZP4cu1tKh7HjNMR/LywXnrB6D+rM41nAWMQKQGl
P5x0p91BnuMmW9URu9QgJRIdKmdUyCn2HHgq1WF5Mb5OefRwlNQzg6lki0Y9RPF1
JHcNIgUvX/+0MnP3hPVLCUQo5t6iDgfeMfXRHjJ0j2STs4uKtXoGhwkGDQUdPkCM
okJgVlkEmsukkXVwkGdqpPVgZce1RSERww1FVZciY8V/dlQQ79wbGIvJW1hsJuNR
mr+6mgiTiwThmZErPsi5Viqn7xe7r8xGkA8jpGwoQxag4jf7klMiYlR2V1WkEqQO
GDRpimc67s4x72RW6f4++NX2eO/vsWsU25a3y3U1dVGmCM7e6XOi+gom19/mYAyk
k+F9131CKm4qG8IypVMEwOs7eIKXUolKuH5pZAgazEoXiLoJSJaKhTlTw3xDMd86
PEhdqbLQVL327IODKtgZa0aQLMc2WtbkscQIfKJLCEBqSCv1+N5YJTQ+uzd2XrTm
BRzf7koPhID9DFYQTu3HJwJGgk1dIALuN2PK7qrjrn+u+pFN5DcScvWPxxGJcEBg
DV+9OM8CO8OmTYT1eZ+w2k65D81zxrF5xtH4jlllHX4L/LkW0NobTiw0adCh4dcN
96g9y1jPIJJFZ9SNU8xjL+DjaHcJuchcFaMSQEMqW08cxSHY8xatNTrOlCSprGR1
hzqlv9pQ4ERK8OvEKfvFAExiNMdrjGd7qxJ0A76Qh1ZtCdYAC+9AHRPyIZSVZEJt
upDJ3+oqaxT2Pkbd5tDEBmx2AH2V8mmVv0U8WQVqScfeNAVCnOxhr3qy2RmkztsO
gFH1/r8Z6FQLzy2guD/AD5zbEeHUP0A8BKQ1YC3DYYGG7RgtkyBIcaw2K56Tnqf5
sXil6beVUGmA1tqXUYr9gS+G+CbxTmtSASveJLUcQ5AN+H4MslbnIpN78cObaumR
kKYxJqmwSNniahfjbKL6oWoBl6xA1/gT1ak+EMwPHGg88e0vH5NBkVqnYqtOtitb
8AZN/5oKgJdfXoJ8UYR2DPovcAR0OcEgtVLDJOkeH6wd0m1Z50RaQOpxn9xDZy8r
ygZam5TfS4JD8y6WZU9zekfPIUEoceaLpiq6D7vAdrFrWMF1bFVp+lO3wVZh20wf
cFEALSElMlKnkZtOYuHuV2LubQW3vxXvWUNpDtQV1u6eWZ/+QI6BBFFzww97Ng22
xRIMTe8QCZ+DqrjLsPpPkS+0LcaVEHhgDL6VMoS2LdJIg6z9wUrh5030tyxuDzvn
r2oawgajZoWNz14EXiHIowkvR8+RU8MzeHxUb3BSqzShCDJGWqklMcplYyc10dW7
/cSrBDl5h7+Kq80USKKnatOTNdomHrXs03/CDx+6ZrdrCY+QxzwCskWw7X0DesgO
n4kSdYCA3Xc+uwI+tlro3MbQ8mHQ2zbfqFHKk2wU876DygZC32Aim9HdPVnEam47
5tLUApkj+uWI4ufETmIBqH6vCA2preSA+Vo6Y0o2UEsg7XNA2vCscEIGScnx0Gz/
8nolT+L9wK5DhdjDugDY2TCFKYu6Cc5Uhg6BVsWxTyP2Opu7tvp8HouogbKlH9VG
RRbuiZnVQxZVsJ0HFw9PfD1aoKvAHJTWf/7YNNusa4vnmEPpo8OQ5zfwbHozh99A
crGBng2t0dgXfBVg4KBYhuQFM8BzcdZPWDxiVUeuQrukpUgRsXzKFN3db2hfT+xB
cd126uHVBl6ZM8DFwmaQvDJXamnV+ONR8NNafEr0k5SdvMROPiC4RFr46fEULLRV
QeM5z4g/quiTHlbxf8C2Z6llHAZLz9yrobFwD8CNTEzbyuyBcO/CtE5fLMJpVSM6
fMXbDsAI9Je4KF3v8TJdK+0Dcz4dPjOm+h0dzUChpSDl6Cov3Ad3GD2DhIXlAjo0
cixt+/y22Qzo20ca3DN4R3Ycw+DP9r0wjjwKRjfCbJtPHGmxzpG8g8I25o30WCza
ocDK7urNjY1geb0Om42sOW7SjtiYjKwCN3jp+JSS+U2tchyEo67XVXmS1+j6ZE0L
Wa93cP2wx8yn99nHc+5vTXVfdNllC41IYvq3gHezL3GUbVFyMok8fySGl3NyaHJV
m46WwdsDU1d1ajS1pRVpFQjwbyJPazZMqqIaDuP/myk2O23wFuKhBGXQgyB0zAqN
uCbHiggmzl/MoFTW1YEFJugIAyJcH1Hyno7D0VP2XqnJ0zi6O/QIyb0I5dFYHDZ2
QlfZWZjM0bn+ORZIIHKp00cgEzVfq30+CpmnLP0bHpNKRxirCG8lKjj4RfptiZtX
rxHevSrR1t4YiqpV1ZXCBQ2mLrVwyU1b9Iw1kUyFNQCWQgsPEhuVnHqewuGvZceX
2ezp1pEP2FHG9e9/2yz8Q0cEBB6FG3GZ8IcVRTBZWGPSxJ6VwBuZxkUSnX0XhxbG
eJWtZGb5DGqL6kCiDHulYW+skwzXMLF4zq1QPPPObei/6YuvQIBIptD9fWvP+mSs
uxYAgepFUJ9INjDotx95oZpZ7hQ+Y3aEIvFFmei7of7xkmeg3Khmkj0RHeXff3WH
ykJvM82k3rNbeqd543vgNCIrtU533oxlOVhzn8XZc/xj5mK/eHQEW4DRbyGptzf8
82595GIZLa+EbD3+GBc1t6jWV+cq4p9YxNn7z2XpFVjjOoD8K+VowJ+6Jwr/v51T
lIRHyng/TzYUGabc1CRtIY+pVU2CRDEsz53JKGDk0jz3X4Yfcv54jg2FRQNLizav
YXOggO5219oBDQ8Dcj/09vlqKXfN6lA6YcXwVLTmcOGzpi+iK6/MpSrELwYdVwnf
R5sNTgpYgrFLU/h5X+J6JMsWKx8Tgva1lhR6gHD1ZNdCpG8ICQ5+wC6qCFYHphdg
OctW7CUtGTS0oO1DEFpArsKgtucEfXaL9b7g8yqPm3rTOJ+tKhZOtqtqr8uBRBHm
/r+UaEKD7XhkCFDRrOTPvEZ1VqabipNgv83uHqgg+pPmJngqyEQ7093mw7YQWUO4
iWvdRn4zAFbQI5RP+pZ+cmq6wGbaMlcqX8WzaF2vzEgYcGk6+Ebm7K6iEE73kyav
19yp9xD4RxesvHz5IzaeqFm9ZaCej2g6LpS9omDokZrWC7ydFdmXXWBKnW1+XBvn
cEJGz9PXEmOJfaLZ9TcZx8VxWJteWfdnDz111s+tn62HNpHiia3DnN+bv/rHj4Q0
Kf5BC8vSv9ce+AnYmNLseEGeGqYM2LXN12aiahycwWX0jW4gtUQKQ0CcyRbYVIip
O9Nyui69C0YcQzMjJzjXSfN1Rr3b6E7eUDvngFPm4ot4eSUUFwUveYEZ4yoO71Ua
eUYsbvhZCoWCFelj/yYfG98fiCi1a3TVNO0UBmortZiNz76eI1snDNWcONhOu4nv
xmRUt83YJfPb3pfi1Hlsuclbl4HmPRI5HVzeBK/uSZojd/9pMtHzikAThRC5Q7m1
gy66Agpl/4vExzeMvRON+4aT32U0a2+IEuqZgonjRtcRUrbdOy56HTCiTpx60lAe
mLaMi2pCTIdykOcNI/SF8lys+sCG8umCDG9xzkxBMOqzib4cVaBIm4SRIXIJDiTD
1U11PZlaIGhhIdzK/ibriLcPI15KpqWGQqiud+lPOY6IGGzjO+j4P6tP0rnLHQ07
wa+xr4JABUioQufRkMQoIbD2NpDE5qgkYnvons5eQWYjleqttIsbQ7FIzdbU9xiB
nFcOCJzPPIk/1nzTbImwd9mMKr6D4lH/92rFyIiWWjGjx9Vi/yJeSfnDGlIognZK
daRbRXI5pf+x2g44kgChxn4hrnL4sGCNQKjcwlGK7josOC7p31zp+17jGisWsA25
cMy/QTADLXJmQP57g2lxiwvPyd/W2irSuc3XiUF8ErG+CXoRMnT+MGklCFZJaNx1
gL6BZeUX5An2JMW+yDm6MBb4YGblxSEEFZbP5ZSRUosDZjHJnmAyxleqLtVNhc/D
HcbDh0sCSQHtyMqxNB21DHmkb7rjS6aUSljaRJ5agnm76RlCS6KDGPhIXVGqNfT4
V1CDkYjOYQs1ILCzxVvyGg+dDvUVl50SEg3558s+oNxlf9UM2Gy874VYin8Kn+8n
n9YWCufiZgTuZgQ4DRAW+M1NZLAVYDnz8DcOQ6QRhi864xwc0mLBTMhBGc3HiitC
uGChpb4rJzUhSwBLanjI9N65baEUq8lTPya3Fwol8ECqYrw9NdulstQbZgrScUDs
AvpaXndWk47FVuVIoBe1QRGZVWe1uh5UpKAkwhK2MhzaMaPuQTh/5P7eosSXjAMT
iYk5mgaTg7WABXr+Dzd7tjW3wZM9AzmIukq4YWuWbh5XoP1HLd5xFyFTyECvOxjp
ETsfNT38Ww/DDSlsHixu3j6u8HeESKggJmXnp56iyLGtMzpKSnBwGpsq6vflOl+Z
dBpG3lCJdTivWGv7sEplsLQsU1pgxyQPW9whk12T6KkxyWjuC7JnrP1qvX+nRzZZ
o5dLaMMz7rVLBewndK/6eM7lS+GS188TEFO/73kDICGVkuR64Ov1gxlvKt6JqQWG
o9bZ22KNFRzA26zFks+kKa7D/FL7H0W52VEnuV4UnKzVYZ5siDyXJfBOsoId3fMX
AcSm/foNQjC0XBaOHs8zFAdI7BSTKNwaM53iuqqq8gJ/ZJxvM2k6IuyGF/7sBH5B
mKeMi/jRs5Y1kqarpjss/m3utrW2I6EyMDSDFh5zxMxiPERbDv3y8g6mL+BKGfMG
9r6jKNJRf1fpFcdG5akltKAbpczGleJyAunSqqWDnFYkhpM/gtDBHoj5+UnLD4QQ
Gv6jPssLuf5d1UgqkhSh1gPairytu8jhUWDWJo9+9x/yc9SY1snMoaq39xl/3fHA
2ENPopw4a9fpHkhH3GfImcRMAiM5LtBYQXKDQLX3hEIU4p2r2wqTY34oLMEZ7mse
TOHF4lsRd7DF2jarVm68+SROmK2CtGrah/jevbDsYWDMT7YFMPVDmXux2kF45VPi
oWOvXRUs7VEJJN8Al5jL3ui560k1/fpM81o7/WYcH+ODNlGsm+Eq/SYWbSl4hHI3
tsr2i/ErWtiKvp4u6iOt61G6BALjlQkC/eV9mBZbOPrNd+IUQ0p+xP+GvWCEBXBT
HLisxoKBfONzLtzXnINLZuPEMbzzgeVtgbzQoWV7cNr6scov5zuaa9LsqcFRhGhH
bcZXW0QwqrBYpCL+us09MrNBmXvvVjNqFj23kgzSr9xVE4wLXhnq77v6XlxMAJrC
u7eZ4Le75Dm0dTQLVZjdA7AeaFkIvQhcREZV7qeH4f2dkYaLIwrMQiLeX3S9KdFO
lJWwqcFNd2jPVNumbOZYhMJP6tCM6B2Iu+vNvbfC10n48bTBjZvd8bweuAejNxqo
cgTpkSnH35WxRCMr6wqJSfUjx2WX6kzKxLQ/+yPa+U6sdF305mzj1+MEYGSXNGvX
HtY82kc1J8M99Z1psWWo6rnDue4arAK+LrfCRPPBfvMbfDry2NH+90OnQBukUuY0
sNlUbNz6fRUtCDSLbvx2gM20k1JLIZZ6lN2WAFtRkg4cAH65yRby3mRPIa8d9mAn
MziJW8C/z2SIFcfaCDDv6HOViKJGQkzRtHLtPiLXtmaMdgfzaSOqS8iSvGw8npkW
HFZh7Hl4OuEduFh8fniwGYxKbVpFv5yWrk3YVD/w0yOY1WVTmhLQKOE3c20voIj6
zjiYvC65gQQFGhPVITOG8Mp0P5ClzX3uC+hfQcuTqCgEDkVJ9htO4Ji6JDX1FYd+
4YuSxNaOORK+/4pGShkF5qwfafb0Z6KxNZJ+n3iaIMOu/By0gWwFqhjFSt8JJnxA
crGa35pOrI9DlwZJB9DO3rA5jyLKX64VumZgPudWZcUxUV7R7fEYXOouZQ+unzC3
03d/NZrp6sWFAkzVWMEOIHHQfaXpxWbP93dYps9dJAw25O0gDLZAg6zJgid0kPc2
rhhCI5fqZ2DSujVtOvK20NY3zx3DO0auHwLZdGWBkc9YJnobJQxEcfaV3p+8FWZZ
HIuzACH5GRG+fxHVmGaJsyV6S1S8htCJ4hViv7gzUUbCEj80uYH+YqqbtZtx/y2x
wCSSa/Sl8JcZsIQLVTsktLbwsivp6IaNn62GKTLf3M4DsS7/jiV3OzpkACaTklj1
NAKsqixOxbuUwm6zANbnEfytN2x8UAO2lEYOb2DqRC7dyc5qFPrzqZWE5I3aUooa
cakaP1qnil/ZAsJoSvKAk2n2qCF1D44dMlEcUlrqJyYID9AzWWmFW57iXQ+tjLZ+
k2tpYP2c3QNUdab4CIQwEVbnIOARRwtkuSV7n+qa79q8Fa4uP9/wbdbJJETXtjBm
pEgyXO++ZMm+a1gGXC1becNFevPB/wXIU7+ImmlXYEaNRgqQ2OSgSqjWyvy14Y8J
QEhHnWBWrIiq0Fth7sCS4QUdmlQ+ksFzqC8Lowvt7jIcv/GsA8MMnsceU346qsi0
dqnfZ1ET3ANDQihgEq1/wTYh1WA6Aokcqx0M1C13XoXs3jWU7PILepNmqK1NPRjA
fDXohEnX+2J7ggoa5MwTRfNpf7a+ga5wpOdMnqdt4pCU8xlcoHUQ5kewBVf05+iW
r8B0WOYeVU3rQ1j0+E6nc/+doWF/69U82nETQbRQpwf3wo5QI+lMShVLadivT1Am
nSf3mUtlQPW91P1mt84kW9IlCMnmgFQchAW8GBetAw/Je68eBdhocy3ZZJ9MLX5w
dPzNB5msQB5Khbzir7ysaC6xSq+3M8VqyOj4oVsF1MV9o2lTD25Nt5QW4KnRRhOl
gQp7IPhfNNyQwQOcz2hpKu2PuoIu2Y4BaehTZbXIgNZ8nmI0aCRRiz+Wpd/X/ZLy
Ty6moRsqdPfQUAJQwEntR2X1okPZ3fBdTM8I1GqyGAvyq7qu5ohcy9XbUGq8ZIn4
ptQfpbpN+EE34KTslU9DsY8CWLM3WRsYtF8Umd62PeOvOklgChv4EhtDMGC3W6Bm
G6pfjtLAoEqCYUga/1rAVWtmg/eyrm9c+HzhsrioAzIssPm2WSJFXPb6kX0LQuu0
uWVSewJ61gPl3W0PMWk71lwUQ0VwuwOeXejaHLI5A1bBCnLu2SwAg0i0GWoDyJ2t
S39sGJEKt1rg9tuJPJxUsoYDNCEaRCkf5cs0D3iY7L/OYMXoRcBraVV8O8BvgxDU
oI2OUnvINnC4mevJfYRYARh6D4Pdt903qaG5+jSAj7+04hsmXbn/vNckf81veChf
/vbaBQXMZIQgBLLeWh4UojwckNQBuhhyYiGgC+Zer9p7OgjSLVM/SqZOPEoHv3g6
AiZbMoFtuQYEAFiuv3n4LHKKoNkNepYv/wlg/ufVsZF3XI9odkW2YkS9xun965nm
1CNphkzzU7jtsKeYFfs8HVdssG/qkOf/Km8qhFwOr/nB/6dtsCc+77jLs5JaK5NZ
XHYjYPR+haQhan+H17gL3andozc1L3vRJpu7sErQ+300uy2DJ1Zn3DTlbSuo+HMX
z8E/SyKEQ2+nJRWYZjBvQBIKCUr5EqjfJls9rdQUgAw2IhNQspCKWOo7TSf3lY9Y
vhOZo16apqESzUYX1NyLAxfDpO/TOlmBGsvNxaHbG+h72q0ABJ1uhUpxHLxhkxtj
U8JnG+1sbxR481JCBZndHQyPpteZoOeLNHj9UUjVUMnkglRYy0wib79ZBy15GcGE
rwmPqCzfHlTbeabMRPFYif9euWDS+mXQRkPYz8Ok9GQYC7wzCJ/8eERyU8eqLXiL
1NJeqLI0Q5uxJ/XkW2RVX9K/S0+907cZgbjA05n6YLuDQ3uO9PrwxXe/vE6aKfqg
1ciiCGoCB/X6YelFPlPFLN7de5fI3sIUgF/KAd0DE7PIP2tM+VFLP69OQHCtmN9e
bAFhVxvTSJGZ6pKwCcuoMewwVi+LvOuLiBQqRt5MVXFJ2nz/duJEC1SS7Zd4JPOl
S/EswoI4d0vO6ts7NdbdW1kG6g3KAelgx1kJun3PzRs37u4GNBpRqXG0Rq4Q/KGo
cIM3gw4SEqefuDQXwJ4J5PV4nMeQYngqMQS0Jt+6DRps0WM8km4WWEZvKUfWl8Wn
VwrUTx7jmztTzGwGxmdysfMAcB9EjgUd4Sw+smMymifOj2nwHOV7PaKMhTgOqjWN
62xWjIb7M55eK7D0wGvjowzXJvPcNgM0L+li5sZVs6+/d/7XpO1zUbUCis+W0AGq
0cJzXWmfnNwZ8vl6UU/vFm93d8lXkG2yDtrpD3r1Aq2Ri4yMBBHdRQNo803MA7Of
9cx274y0ijogoa3E9MlnJsJEkZAdHajRwM/q3ZbU82uBmy85r+sYlfUeOobEIYgs
hxF3IEXzUfwlDTFvrZgx/f79VQvxm0JUDM2TexLDKG/SooxUR58R+8JS+nBAcm0q
+T4yE36F4bCb2vwEvKKhOY8TTm8Ge5wu67qS94Qo3BYxDmHT11xAHEMQ9qqT4xQ1
aFTT4gf/SR8gdoW5lIyT6M3Lym9yRBPwGm7xmtzd7qruI8K7ui5SEAPgnAnNz3B9
/3duKlhYpbk8QpOM5IuluvYU5IqP0T4oAO5X1wNRsLVgFLDZaqaqiiE/qFZwAmjJ
VI5zcUkQ/qFe5BV8Vrb5e3eaZxQm0gc4vdpGG6LYnij/vAX++xaNU8lHBc7jDVVQ
VSwdSLtBgDOec85DmHhxHy5rmWdskj/O3kkqK81nEuTImuM8MbDmUmsgIKwA5D0y
tyoQx7O6/is2bswfEO4yjWanbpmomZc4PkuvrVwwcgJee/D5rxJY8x1Tczz33HgP
Xs7lp+DDZTiZ36FEkVBiwI3nFhWgp7pvwN/IU7oodkHfZlV7I9vEM0pueMuARK0e
m+08gpxnYn1FVNADUvKGp8DCTEsEyVrLMS/oUs1joXWC1dFHwgWdc0mGcHaRk/wL
zNDW9S59tW27wR0DSJg6X5pyd4t38p3ISpREmqunktIN2+UmPS5bOw6pwTmBx0/Q
wWNke/iA0WT1NsEuPXrq6r0jloz0H+pXrz5LrmYfeV6UEcEA26BTcUtV81ytswjC
H11NN1bmC5HFXU7juNJTyvmvWluX85XmJqZJ21zXlIQNi2v/zQ9JCW5QuDzrZUne
vlj4g9z3CoyQNp3oogQa3MIVboFeeyHSsE1Iyo+yaJDc7jJO98If1q9ml3fj6l78
ozwtUSdd9pJ1PA9g1mJ2RfAfmrYazqy8Vkmq/Hut/SsUMjBaFv0bXVXvrmNl4AQ+
zL+Geh6YScukXHO0UyTsNCtQH8TDQ1s5hv38v5nB41FnwQ2pPnldEdrZYjrP5Bre
WFlKkHsyIPGpE+w9ypXEGRPbU8R5p20WI3EGC4iMHgWJq5BKTcWPXgc4dfw1B08C
vBwUCHuQNdU7xKC60F+BQLtERiGGweDOd9Dpqy/+JvHS3r8YQQngnU2L8Tjt+WVr
1oiov/MKqajXqdrIOhe0n/Q/bclX9BaECVE/bbNX/it5E9iopaUo8KNuvFgiFnhB
ip8xW4hbBgF9+yA93/3fIfak7LPS5vkOxy2VN8X25dSBic/ZTkk7y7JSYc0nIybu
h5HajX9Pkwk0cpAuK6solHpX6Oay15DdBqV8VNklmByJ9iiYIWHn5cwNSJgAN/42
tiPLbtmYtkhnNcY8ryX5QYqH6zE0Nb85HgQ5CMlh1VlhMbaCpUm0wbI0ccSoOSJw
hzawbuKsK2kHBPPIr91f3ux8511cJZWzdT3vrmWyIu9IdQtldOoSEDPxnL26pCeP
MWFRgQfhF3K5fg88mJ+6A45hDv/OJ0cuHBsseiHFATxWn3XwWU477FFN4wgCVC2i
JcHKI7QwJ0+DdfmDC8aeCyZOslcIFJCcGnD5G9QOiuUipiSNI3xytNx9U1WRTNe/
L4uUk9wZGwU1zUsyM29yqHPLDhFMtygUfZEt00qeIv6MNpfAWJZt2wBJ0tHX2ceG
YnEZRbo1WJDHPJxg7SietkijYmUOyH2M5ktB50RVEkuZvYPZ7XwkLrYEIYDnJfcl
BAbKRlT8XxT1V6FGGGm3LZaIg62i/OwpwcdWN1HrhDAh4H4+NAx4bdyeSdFdAYvs
gMzBJf2LVvux0iVNPagUcPTI98I9B5vhjR5KCEVUEGaxHYfNztTkj6XsgrlbbcGM
S34bN2WL1hxe2AaWVEYAEf/kvvtHdsrcZOmf7iqQEzpasH0qOXAabbI1hZmHtMzN
mM/c4tSFHv+2QEKmHqoyxxttkGj0DqyMjWJEYJyjwQucK2b2dXS1sEK93KjdNwdS
Dsoo+KaOClwtmVa7ymEn5YTGxG5pagR5kedNIUVL6+GpNKAOxQG9F7nHsB5+D+a5
ptl+0O+JdUwh+6ncLqcB3me7AY2GJD9quKr+Di+CNJRexugyB2630ZLyEZ0oyM9Q
GUB9SAX6S5xhDoxyPP0t7Xr7X+7JuTCB6LCQ4zWWlCygIcvCtnejhLcRziDnSYzo
CaS4wKGyNrPpp6rom9ScjvrxFVO9cFjaDK98auHleVBKkf1uRCTZQGsXzZfXFRBx
i42FwroplxvuIamVHZLalOgCP32ctIdLh3J8TWoqYt9ecEPPO/+QnAG6RUNJAkr/
JE/LBNTIzIpS46Kf0UerUKyOx9MQwnudHRPiQKf5+WQ5qdL/pfi6RNZqFOrVbRtx
qtSKYCJ73YS7gpyDRSlBHhGWaI3voH7SCLcY0nWjmNkpbM5OyvOSiJNjFw78Vv2S
3xBf8q8vc9faMSOe3KQjSMZ/cK8PpDAY0JwUmibrtFHLN+jnc74kNwEI+FuRyFof
8IyoW5Qrpbg6x/2XWGxa9tuj0E7BQdodPH0hM8qPH0/OVH/xcYRnOsUnyXL8PUz8
Mxf6Ni2tXMJ+vapDsNsOQluDCGUTvdyQpngpqY1Is/EZ2wlLBgedS9w/Mry3mtsm
dtJNzWGeHeND3IplcHM3Q/ZD1fCq5c+Jn+YzpS0fh0nYf894gAixNgSbgI2JP0n/
H1YaHrvYbesJPHqkJ/oatY/9MSFFlhHbapDX46vPO6Xs7qWeZkMMEb1IOwQwi3bw
2cb4q8dZG9A45aL3GFy1GEVbd2WLOlJpTWxpgZt0KzZI1uWd4aAc6p7FbTobmUg0
6VdYWyvB03zNkPlTnSF/hlr719njDF7B2suSTeSkDr6XueZ0qlbYyYgkXFiRFWV7
nTrtJ1m7r9Bt0iVcri0JJOgyR5tXJAyVJzTlsJBS+H0+QyyyqfREEtovkNhnVLbS
sYWZ+0YhJxORhBN/P9hfCaH0VX8TkbXaY3LaUzZ9IJntyMxdzuricUrNe576jzLR
hyKI91N88/vibUNzK4mSa+E/AAtvtMLdzSwrD4fnkWBXA6MDjYVM5zfxNHtLNENn
TGo8JEuvlJuunC3ei0A52HopdjcDj0p0FKWKza3HiZvz6pG4HgfyvSDbafG+DFOC
i4+CCCC1h8fLKhP/BQD2Qs4lMDFgmsNrOD+N7NoHKlXk06PiNaR5Mje1r3D1gqgK
ReP7ri2dixdZ9NInDBaUfvKH8h1gpgA/U7XUN2boOCL/a0YMFsJWWlPHSThXs0ML
7z0qxWbT0YJz1+Iq0PyTMFP1OnzD1bKuKXvKzlpqdEGeWdQN+rObPmlz7HCsjn+r
kNgorE6TjuNZ+v2T9msvW3CRMsrdqKFvBMEypjAIPg9paqhyQifLvqwSPJwBERCW
aG1pKwJtnCJz1buwhPWLVH6fPPgfbh/L2qMT2FS+O68t5Gc2MfDlKvhei72ZOE5J
4P37qIcRwpWs5R+Sko/m8mYi/vFmRIOBNX+aaLw8o/pXDpew2y3CfQnNbjZNZC/b
jd/9tkBpEAyTzTat0gJ9YiX9bVAKhs/1AxPeLeEpO0Yt2hj82vJuYqHv4l1K//iF
DWODoz9NCMnpr5bUxMWevD2j7UblRewEVSgNT1PvF1CQNVwj4TqpWQHWYo6RAWva
YySPmPPSjdEVMndWC610EUrEhtHf1D/cp/3bAflQR9+yjc97zlCrRf3g5ZKp194l
930qhu/564tLpfPqo96nt9I96uJl3BtzTzcQFi7heYW5vzDp5vJbkrlrZiXaIsFH
wl/g9X1ynwn5BRTwPkzKG7mi2nBuGn23MrmgE9449TBydNZZ9ax4CGkkwnLYg9po
9AflKxtEg/rbA8ZMWzeI8lygMktZ6hbC9jXoUJtPAhMsXh11U57zzAwLIlL4e0Mf
S3gFZAcsYpFun3JNqlx1M5snZV2JYpXdl8WydQ91QVbmeRullGF5jwDgRh85tyuC
R30dMBsd8Oo4Cp+pTBpCeKUz/VqQ9MBti22o+8hYzc1rbIQcugIMQnMg9yoMvUzG
5zaeKYXMPYvUM2Rs12zS+1UPa4avVXrZCqweW2QqQ9B3vB7VYmZzxSE8y21ZUrjN
X7ngRI9qegDjBG7U56lVTqe2Av8YIxzBOSglnEhbptztPfWRjAycmDE2g1tqFdDf
8fZz8Ijt/RwpUaH++hwr8aFAJMPgnosd4zi4PaJHxHybMUD5KVlMckCPMMz3nwZj
WWQm2IJAkm1HoOVxfIFusvMYzM24TzU9WIZZH5uV1nFGcnzLOdUXtpVIRvtPYCWt
+7UlyoHE+eBDoYEZD2Igv6gvI4xDWZzgXazZYj1ZqUx5s9gzJ3NhmhIomBk0Uctp
KFf4H7fWb6z1ds7Bhjde9n81/XKPSoCUjd/9SVTItYlW8In3FpUVGxhicKsvmenk
DDONrtldrtfv2vOYqTokzEkUOQ5TZTw6HVj3L0ANVOuqVm/XMB2RkzceZGm1XyUz
Auu32ks0X2cMCJZBFogYXsVCBCkZWwSHdWv4hJL5N55QPfZNoEH1ytkOFqbDkefM
HyYXEpPhp2SDWEHb0FWylULUwlZpIjvJ+OQGuv85QY0WPD6/2V1pUGa4jg2hoAXp
7VU730QqW8dHnDqpUs4t6M8DvRIhSORSJmBZqRKDTvWNvEZwkHBpbhcZm6U1O/cN
1HGLqI+Sue364RGdms7vX7Nwm9/BGk2ire+5qI7gXn+NDuzq48WCCzSV71iSQ0Ld
PcelsSSGhYRy1uB9KOEnY+QA3eNVsgIYKGJ9yw1a7+T6D5t+/6vAuYXF4HV+p+gi
5tP1+6uJxYYajmVDSXkOFsn0j4S5/V9Dos+Kc00jp+g5dVm2fVa780+qxED64X/1
KR17vh6JPBJJluBY0jxZdZsum9yPQSqlwmYpC6PAoi2NYqV8V4rHvUfThaGmU+E2
1mdLFVrpaiaurlH/F6cRV2PPwSnybaHpNnzbVkz9I/6dS3GDzaVmwD+sfJn1Qxky
TYw3A50FfDGZf8DCvehTuOdnKFhJqTbMI6WZlqxeYSl94E7zvbMk0uaWzA1UcLhU
rszq69TlLlJ1SznWCZ4Ii2BJVV2b4RpqUVAjjhqc9hbiz0MStOpJtoQKMm9ssjhf
sFjk+qsrPCH1+0qbm5SGnjq/Ow02H0nUSwiO4NtjkE2BxskXOvy6YYitaaS9LC0l
3tJcFLVCNlFM2r5vc0upM1PbmWvjGnrhaIi6kvkgQZ5XtzRVf2AgzbzOKE/3NUKT
aZKF/3UF2y/I+BUSz0wQK1/2jZqLKIbh7Gben9Sv+rQ5zBrkrHhaXjZXVzkVb3JC
pGrxbm3qk+UaaNsNHu+1oQb6Q9eETRHI0WMs0uMcnAAufqwEF1KeksptVCuOcOgW
c/c1+ProOxJZIx70wlmZOwRULWW9F3FS3YV+GHWvP7AldeCp9JTtTtOSsWv5Ousz
Ynrxq93Vhq/W3OEW6OLiPlWchkBF3gfbNH/0oDq8sW+HR3I+ok1IMF5pGZbuy350
+WRDjev4z1wbM4oMeGgbEekeLhVIa5Xwc0QjyW2JXvJ+cYrIonQzwF3it8C97bZo
YEqboznu4nGQRtdaD0S/IXKXVynQPxrK4rvAXlhuKY7XA3o6fl+fjCubKAEIbFa/
cQOU5X3Jt5q0lNE/ousi+1C3PJHMSM8AWXmx+0+iG43wsgBa9UWDNz+CvFQ16QEA
wFjAMpGmUW/m+EnZgVLEsSZlMQr3DXTYYj1Bv8zcD2pmQ+rUYSGbNZ19LJvkPZ4W
c2GIFVvjXeBXlj2c3HiroRAgsYt5dW805NXPfWYmGCWBfKEztPyuTenZneney/4O
mDBo03Mz0XWA8s4omYGUNly13xmY/T3Oj9JIMWbRkCFtDnjV8Wxt2LDvyMq8ejp3
QNUtSS3pSZcMB+yW5ZY2S0p4Xs3t2NXEmgIJdje7sWLW/btn/E9MlhHeWPGDlerA
8Q8ePU3xi8sXpvz7XNBF1gW5XN/05s5OvwwXMwWurH6+VPQMxfFzUOC9Wr/w2znI
L+pJFbbnKKX1WrOvEYKIBGbJ6K8LYgNLfcvyyaf3/Wi+k8hkoqXlklDQ6ajxcLNA
4KVHIYlwK0WXKAHFbieu+8iNxs8csSxErj1sEiiXgLQCl92CECRhZ7y763EIdo/y
x/A0A6iDhUyDTAciHetWzxKRE5/jjAMK02+p/jsGzX0bkupMx/Wmzj72wFajIwty
Hw0NSS9pVe9+wOSPiijiP7eTcO3Lw94ZDCu1v8M2s0wanELv0NIJwpi/7NR9Ty6a
5TfCgW5JDNwrb8VoJbUpUsZjMf8VqZRQR+Z0IZpLl0lgwPnA4K+T0EDVZ0vLbVWV
NkA48bXr1yeIGaFRUSel0KFRs+4CaQXQgRxW/E11uPrvXBYq0T3WdxnHVAY8MSFZ
fHhi4lfrhSlbCHZUXuozG5uInVwS31ed1LvMOZULH9CHJyovS6vY8pmOZGp6lL92
YTfyAzbIftOdkRdJKN1OaUa78w2ZQXWNUkeryuV5uQz/RTOs3OV0Q5eglFUQbawA
FPbod4QvtgGKw+GdEP9shPxsHWLhPL5qgUwSC+QOvLOV26LGNJrkKCWtCyERMJg0
67m26+wG6bhG6gkOaW0J6aCN1kitjIu9dK1atqyf/m7urNwsY2uTJDiC1iiR7sXM
raHUeLtARVcNl/K2Zq6Mmf2QNUt8VzN4KGSjBTmn53z7vJy6BO2KndjdLimlgIqK
AABsmGz47N7069mTki65Hn6bq6BhATk27c7UxTaNCQyIlk821n+NftG+giENHJY1
i1o9MofxfVATE8biJtoCzz/Zw79AlvnbK5Y6cB+jn4KmRwXaVQz7YoxVu7ePB+5A
446YHqe8iEa+J4SmC7fcPEBUX2xrpnqeu96GIPs7l90aLk9UbyGVqnnj42J3HMo3
TUnxPRMImwGzoDFaV7ycBj7JnWgcEVwp7Fa5UCXkMLSb14Fo+GFY6EVkOu1L/RgG
KOTlIpEjNerwylLbIH0sUxEsdc/XpRjvOpDEGDYL46TmyAumzW0hnSu2brUYUcpk
M7FXrbPCRrp02uCsKZiBq5hIyUCp7y3FKJgTU0ydVtY5JL7HZDeDwfZoM9EJ7Dq9
dtkXR+C/GuwqPxB5TNbEl2qvcxPearP4o4bxdkjzx29npOt7BxZ9glVYt9QozIRx
dB5Huq53QjfAYUILRizEtzH59xWe8ZA1Lnn6ZlWc1q30v0q7oGSsnaEERZjpAmL2
Jvw8i67JBClXnB94BJoSxk7jTV/a4tetuEmMTeyVt7iUHHPNd4qU+xK9I+/8B2Cc
MsjoG+w9KrHsZQVixxt6GGCarBot2RDDV2LKcitYCFWc/uG2ryQzmp4bA10/5Z6g
pL/kc7ZGBNHa3lfh31sMyOChQAY5vUzMtorNJPxgL+qdO6tOBO84ToC+LDgj7gZZ
rG1v59/LdKHx/hM3zdUSsr135zMF6Rr3EEiLmshavLi7WbBsrVgRorIDt/clhvnW
4U+DOmu5waUwAt6RKyCJKnWRIjLJGuy6x/wuMfMwHVcGUf/D06JEwnXkzPJRxWFv
6SGr3uNZ9mVbIRT1zWkqKidl1C1VOkFPrZWofACUr1gganBOsVnOcRftVjmXAlvB
1iC5rUzUNdjLSF8hQv6YaCP+p/SqAKn2rP2XFMQsr/ejHhBmsmeONuKevIlGIcgM
y8pNmRdNWKnF5UKeYXnofsiyB6xokRkAuZ6a8tIE4YxteRBVXTCc6Zg/fR6jQbP2
gPmHPf2iNtT4o1WfITX89vNHvKjebjDCTGxLFAmNzqpJ5FEjU+XltFwXifhcmF+v
qTiJ+qypqq39QP3majCJ+7gH5+NtL5lbHaNgbArLQdkMIOMCJZbNIJ1xCh765xBv
Ce0ivT6GCVtqXBOAdjsfGqVcJi41VKRuKIwQYRHiA3JN1vqrz3eTklC9IJh+rXCk
+kODZuAEMxJgJm9k248V2+vvqDLwCYzdCajCtSLc3Yy0R5x+Oc+dBk1YbcGQCpzy
16f+MpcM/5jDv2yj5m84tspf8OJj2bJre4xUVpORhFv9loteJCi3b/N/1n3+0ZWb
sBduTpQ6VCMjZbuPrIG1dPWJnqC7udY+2evvR9MsRSQt4ce7UwconjkMKIM33qe9
n7IXSWJULm+I6Ehe7ya0E6NJP8dhOaDGmDv8+jAJp1CL3Le0MAd2Rc5zR9SrNR/a
0qz37fG7mh6zHJKlCidMjeaqDDepEyYS+Rk5WQUnSbXIwZ/CnektghDi6NpdhKTG
/0MbiX9IDPyBIA0B8iUqT9HJWe9ppjH4yBS0VJvmjjWpKM0cC0pFBIyAz8fFndiy
C9ht/p+fSFLeOH8cP4VWlkFyEQvio3wBVpP0Ea29G7xAXF6gqQC9vjRcP7FpNwko
5v0Kjmor2tGtT6PZhtVwRfC4/BEdQRaJ+Fl3ycS7X2Izh0H1fFRq9mf/aiO2LSAV
2pyuLVFTqQFK+m8e5szYidXRr4VNwExyKxKvBK0b9MGfrHv/58JTyZeU5MJpATQZ
gqzkojFXIHIUkIpXQ1vvoRWDW0qYPgM3lOQfzW0/v7+r0mHaRo2rbKktMS0z7y7l
NosyoMxDRA+OwwptATlvC2jqMWjLTKwE0dvO9X0udnpsAe6kcklFgW0SeymepBcD
rfrd+aLblq8mUsKX/7zfcWMhwVIXfxJLqH325hFdIwb/bEzz/q2roicuS6y7QcDP
a2dOHfANRoU21VTz44UK0H9Y60tSzwASz6Y4dsIjbOM9vEPxOUmFeiaUZ16wlDBK
pkqpbpbDU8LgrpjBNJ/whz0Dp7nWiX7OF7lJEY9cLGNF5KBI/uJyOKe46DyHxWEk
RNioOWxzQTtmhUDAtQKxpAvdKcOj7GbYegZSy4OR1xidUMe2ywtOCal53+lOE2zS
Pw6puwkstyfwWxuoF4I0qL/E3evWF3A+e8vcSJN6bgl8hcGn0kMEtHiKajDIMTO/
mRFQT0LIRrDQLl2dgnkkDYEzvOfI0n2cLRJJp8r+sRhTvVYxNwc9KxXV/fgWfDdg
amj831leAh9zBhbdUe2L/erAxqlJRaEvexKE3vggrns7jkDxotTfmmExbzheOr2o
nY6/UPfy5Klb6WYv40DLacjRQDv2N5x64HhHsxvn2appW2pt3uerzqsY5fxhPSXB
J3kt+4A0PsBzfxLHHqx15clYALBnMPTSqgLzvb9Ki2YqQ2btDA3Y3vISiiXyqgxo
QEi9nL0UED77fYAr8X30JsfXz0R0lFj92gAkwkR+0gcQzFZLesil53CR441udLPC
6maoyP1mhPd8VoHdRendIQjt88vW0D42hdAePNLhEA6DZuzUTfrk7CYlGS2H9wg0
HT25EGvy5cWXDKc3DYzPh2TwsOFjkIhBE+lhoHLAbBS0vPZqpmGko2eMEOdTFyRa
7NS07dhqJl4XNqb9u+bl2uRzxYHvJJ/sxjuhYPnKkO78uY8fyeAZMuglBAHtwk77
jWOi0x8r8FAA8Q9okM2GN6AY/uHzN0LczcwsLycImoGC2xnTAOB3gUhroD6SLttN
P7T/eYF+MJ1fSBMs3J2tflCoU5E+VBPSNj87iyoAmlQxttxJGsYTBSxY1AvmRJC4
tpMS8jKNOWEPqGeJa/v2ZVNZOYffpsj8tDNp/oKP4YhmfVvjpGvsJjl6FYdaqM4M
B1wWQzBWtP9OA8fNRtt4IoifQiDu6Y/xrTvWfVfNZrfweeJVuftl4jc4854X7ZCq
71eSyexFEVMuux7eaElFe01aj7mlJPhEp1r5XmQs4SPiFIlc0qBNDXq2WN90OcBE
OSXJK5eABegvjtI4+EwKEmbtjOkHZ+Mmt+FC90Gq1+fFCdP5q0k2quP6bujri+2n
lUZk6nvXcT7PNX42/YCe/ONgq8wtYeDLfUGIDt49JHQ9ld7cHohLDghZaVg0KcC9
xPLaD+6xqE+i3bAwrQN7tcqUv/IG7eK+rgFbgIGdGNMvpPWhGGyRgMc3l55wVIO2
Xl+EnfnbWZheOuTMo24wtSCVCMXgMkDJ7qvs7o6ayTKpMJZ8YgVEk4VcJoIZ7maf
xKoBgn3LIBo89cNv4RJG8kzUvQJ+7f53A50DL3N1/3E+aUYe11Kw2S1qYKn/JOCf
vmtS2Vi1B4ekWLL5Xaligfho9QnarYAHRtjfF+EKZLUUaEcx6sdLKuRX/knFQR+K
ySlinyXlgfNOBNcPV+hHQGCWOR77pko3TspV1+hJw7pH7fxMAhX53EErk2095OD6
e118XneboZJWLpQpQyRoC0WvgRBMZ53DuzcaJPj+64ErMpJ8DZpYrcyMVXPqUgpL
UrVmR+RdkcFBOYMuRxReksjs3p+l3X74Dwx73kuCOmHxhB03Z+9ug4451whVVpCP
fxNOtgJhszX6jmFtyohtYrT2D5QFkmUV5q2OuT+GiCbsA8tT4vgvDMiV0NXAiDmI
KlOMvv31o20UfZku/1HHELsts9oGu5oexgWgLqOKM1UT7wR8HWf79MWHygiTuXUA
QtpDhEEPkQWq7OO6tl4TK9ih/g4m3Jw9pQK6spqbGo0gbpzR27iFeGkIMODhpin2
tVShSBi2oxKpN/qlIUDOeKgLYPvEEv7MD4jGfP03h3aNh8ZYJWoYKHON73oIgAsz
ZQM8WnbdKPaPtv7rS7kCA5M1173A2K76UbzAssCvafSYINPu3EAiXhW1n/5k9C2M
RYhXwmupHkV+54lU5FVZECrPDNzsbl9rK5ohLaaPfNbiaEwjQ64wzMwA4j06s6zo
1WCH0mTmpRDzF5JhX3pgkpSj8+bPGU2t1eRnYf2S6qP6ENBA9N1o9/dJtls3kRTA
KKqATNf0GTkUb4N8G+JlgLY7kkwT1kIpbQbyA0Yd69bPujiB+2Mh8/fo2BqIlWno
Y7gTfICJ8qPGlDf6av5bPQ7brh9NQFaoaLm8opbFvTmrpjmPch8cOZyxhaeME/SY
zstb9raFPfLUyu/JHVr7Q+HUcvJsXvNmey4BAk09ofldFuPFMt4oR9iF+lFoOxYE
Oo3d58BV4440piBimZ6P0FmT9iC636Uiu7ArJOAx9f/5mluvP/75Doznpd3IdSi5
/jOy5TtjkkWBji8evU0fYPaMUbwBOr6Hu05BnEmKcLspBCzZ2LW7AQUk8ue0zgCF
4BDS0uDwI9VJNqknYZ+2DROyi/G3nEA86x7VwsNaGW6Or+eZa4EzG82lVPF/XGB4
rQbSsNZJr9K+qhHbJFwmX5lP7sIli4NjE+IofDOODzcqBbEMXOIHuOjsJAhpJA7O
2EkWEgx8Cm1nKESnPUepSOdbcG9Ct0D8wGHDNHh30pdb1mV6lgNxGuDs94GZXTex
WT1Dh6czTVyS7GSp7q/8icbTlnxFv/d+yKH3Hx74lCCJAnlcZQr1TbMX7K5bV3L2
9UiRAafbCLr2lgEsU6zuAno9dkQrrEwBQMNXPjqFxn0zziAoLeo7TgjvjLB5VZDM
sO+IeKuRH+nMuzRfvifQbyIUlZ5yF69rvfI0SUB9ApeGt5NvEwnogy1f/KEh96mj
kFQGRZCNuLKH9gbW6LQ0W0HvhNw9UB7ahi4lYS00j9pVT9tJXehwTum7xcTQGHJV
t3j90UVuqgP+d/Co2vGIrBdbnyprVm28bDSqZ0i6XnhTc7lchuO6grZ45nZXxjQ3
x9Am//1u7R9V3t/ZOmu5PrO60P/g/ERdLgdPe6FvIoQzeUr+21loQ7/O19Xqh5iQ
s3gdRiGvNF7EWkoFi27/QuP14QHfBvDJDq15jT4tBUf9HvXPaoysPZ1Ehj769oCf
RnP4CUTZUYxYgpmn8SVYdLSfcGf2P97+LdEA528s8HnbKDUKXjeo6ByiAOnndfK1
ne8sD9px1be3/SgyqblcYPLbsxErlQ1GmYKsY1ocJBtGzWqoItdQg+TVz4RdC0Rv
klnNi9Lm1/VwdbjvbBZGa8vVRU+Ij4QOS86QJe92fYb2INgwJ2K5ZAW/hCmL87cc
AzVV6Z9DmqIoWXQoDGccwrQBTYcCpBXNFwdJOn0TYdsR7NthqUXZiv84i7YBGE63
gWEOw++FL31AHb725ewW43zibcCCN9wMeDry6H1X6AmYhMRScEtERVtYBBd2wLr0
/5uhVFew2A+EEEC4vogbTud1+W8d8may7yV1m6uehfPb2+SNORuksXhtQkdGv16h
R/n68zYKpJHPeFKv9JN6afDOi4x3LYZ9lBJmeO/12YumQj0NONkVGnL0L3HU865c
G8gCM3GDRy8jCneuLXncdlFr3TpVimjK4OdaDJ/OvRCK8u5vgzc91VJhivswv+Nm
nHxapn4p+iwAjCA+Dlty01Vw5kbvEdq4oMxx9H9/JcIHdoTY/7bqAjr7dROUxoIW
3OmXCl54L4pOaldPHWX0+UqngslsSkHfQvfDW4qIhv0jocrn1ISK4MNQMT9zrtnJ
DEI3pl5BLyPv4Zth4j8stG7tPo+ab5W3O0/E+PtoOWHg5dSXuNdSCF/6RIShzycM
AYIJOsn0BSVQAnCaPL2DrF0xgxcng+ZG4FuZ679h9A3P2MovzoC9WdEutiRhoMm0
+QpqQNDLIF0x/VtthvVN+144jCkAbw7dEVSquKNvBnu+5z6mUhyRMaL0pVvHmOuc
4LPwIJPFclD3vsK4ySGLgJAHHbM6l4F9kT/ie4B//wME7pfkZZch92vXQBA2h9ND
ls7hQ3WSvqMjSh/dbUFnkcoT+28ioaglHy1LtWtom5zhLKT+4AqSYhmPVARt4AYJ
DgL2UslSoPxIuf6FJsCxyPuz7FTgSId5J4HFrpeYhKtNI6d1LqfbsRpdC0zkcgef
6yc1NXvygGDYKRSd2MpSi213rcqL/iszvIRDAblGGtMmVH8hDfptKTdGVOlo6TAf
QNxhikhHBTHthgm0EPoSguhu263UCnYgNx4V6wNMvDtMbk+fvFvk/ghsXgpcLrhM
W9wGuNAN/jn1UbzzHoDCFBE7Hy1TeLX/gS7/BQ/pRvZQnocBf0uIxe5UoKNYO5Jg
cRw8ZspYIN29PiJZqLBDQbchEWfMGVvdFuerTDmlUkg4y7dvIel8w8GpNURcZl6d
m2udSnDBLIeEDA2ZRkwmXHT971UCqy+84GAtZqE1VWdBNpdcwCBZ9t9uH7laj/LF
IKbqZ4wfuC+k/fjfdw2Oh4GYsjfXLG1iNFarVTbtWs5tOrzkiQOPpYRwqLWhPBBL
vKbxnWrR+5e8owP/MpI+ldMS+2BGMR73PoB5j6hTJx/jcJcEiRrbPCM/BCpdZ+7r
DbpeTay4d2dyZGC1XmprL3y7eQ+/H+SHf9O3cgXvlnnWfeeO8Ae/r/3LZs4cYdmU
b9Y57n9kLwORILndUTPu+SjgOct5u+VMdWG9egxAXuizZHeHhX+EOqD9FWeqhJ1N
caRUsMPL4P7fX/AfHTqlt0DGcBH7GvnOfnCvIR32YS/gJRyQvBJafQNDgG/We2eP
00S8nm74Cs74bwdW7oY0A24Xk362P7PXnbbh92sXvQMD+Ku7gR1FlEFaarpauB0h
NjTYGH4URK4yFKZ7mJlRdwu7u9xjIDgR4RKuuqq0Zvwq+qXKb4/Na7N4xiTy9DPB
kv7tQ9WnAY1lGy4lVE3eu/R+e5Q3cFNFTx5ARo44prIukv2MjkMjVDBFE/jTcAV6
znednek9vk/WbQkWgm7qeRg7o6vJi6MWwtrwo9rhyYZaloO2m9AO4e7inAiDqNpx
rqiA+J5go+61JVdFxLxn+Hyza7Ly86dtMVmZoOUh9mFcjV58lojlD7NcVlDVHtPn
w6OL5WFaF9qrUltcVJ8QZV2AWjwpDyjbpwkHV5zwZhaJnsEcncxxU0xt4uToON6O
LyNE86yWD/o08oqQT7dLKXQsCPfgl0hRKDdf0NVTjj7kqSwfWjyqvqvy8vLDSs/r
7B4DdGbnthZN5XNG8e2euRx3UfvFUQAoWOTivwBNK/JeeM4OkRSqV8LfDpJW6Qs7
KVXvAmSiIEkC3zCXdwtMGiW5cHcJC4KQWdt+Thfh0EPYY8GP1kxzT490dWgkB6LO
NngE8rrvljtL0PrBqykN09oD4jVLMqoBVPL19sgA2xbBUNF29UTXIzrL0Z3NZBYT
odlN9DYRvibhX6na8sFVbrg0woZb4wRh1zVJNfqovRxuMtIb6/76XPpght7ggwPk
HRBvvhCX/oT2PbzlknxhsWn3dkCtT3E7yKJcLMumuhzrRke4RtpVhfITKyW5CJMs
JeXFT/30ScAtYzyvGkcMwk+6QY5ZP+qlbamvqIixBkhGoNod6Fr0QI2JUDFCfuiT
fuak7AgyAu6Mhn8CpRLW/ZanHj/DWhQ3v+nrMLtuLG1lkGGgGL/qQlD3tTOD/X5J
3M5hGAiY7zJC+fLzLrmRR45ihhuwlRRz0Uhspa9ENlSjj9NOTv3t7ZSzCkIjk5qG
wEhNANtH2M32vGw2RhwPDXjxuINrb2pC9Vdf5j8n3dsGxSivfoaWJ0XFRQZCj95H
t56FY7oSR4EzGCUakXk7O1Yw5vCIl7iZ3tUTjuTUq/vE0zzSP6aKtKvvJ0c0O2bG
yASuNiyGwsLsk2OPYr5Mum2PvOtyxNsS/WDfy6U2J3458ws/oyrIqmpJZ5yWVpVL
VB5IssKGyKqA/mIukhppjkUWRMMU/C+8qO5DqcD5umvZ8redU3poaWtslIU4e99s
a+QDw+RWbFxHsCBfmddPOYk+nYeJp2EnCasSDR5B8TIkWovAQj0eDiG5TDSnKLHb
TTDf8zMtiTqYqaLKCLMzhZngzRN2g96h7UdEYDmgG3qT7wF+PhCLmAMu9f1dqa2V
Dz0cEaJ+LspmkfBF31Wr+kIF6V6DiwFtQ1jmLF6MArU/MyyeaMgNq3zD+rVEHCNQ
65QAY0naFvaF3bp+CV/GCa96jvpl+GV55FSssNHIKCowugdMjDnaX+c9bolemNHG
Du6MhI7tA5QI0tef0xMrv2+KMIyZPYpdZ9OYTlCgmbpayGSwMBVKqodfHsqJrpHm
tJQ/dAqkrr3mhReE5y6JTuAKKfJmVmq4L8+05Lw6Z0p1UBfvElblSS6rPvXPHgeG
uQU1tnnFDcn9rkUtuQWQt43hPocgilRfojTjYa4cHhjDaNo177fBx5d8DPgDyeLQ
q5qfn0gjldQvmfygzRRtClDO7r6uoiZPxCNdnX8dtl89AW6G9Jf433LCfqxx/TqZ
+wTIhDs1QbJeUc5cNF1LSJcuJJ7Ec5LBYqQVGTJzNFQTG1UD1W8yamvnXUeer/Mo
nMSkJSDsJpXsX3Yk4nV/zr2WCMREuk58BSxQoElm9RV0DH6ZOCIfvC4yxroAI7vE
TJT9N64e0a7Tc93tgRpMIHIa/X9omv4py+AmSx/NDCnltn4eTVeqY542Dka/ucV+
geQ8VvLdEcn34YGUUz4yJ288j0S8TiATD3ZlvWH7XOtDkKpjZxR2IdKBP4mbfD/p
ahuCaad9KIE4+Wymm4S8VbjXYMm2BwRvSXupoMUUwHgk/eqeNy3JLK1sj0Q+1zNn
OvNH4ZiXETWqlw4NDyVwg1mstlWMEoIicmeYDXLcXziRVAwsZTq0D29g18BZKULt
vkUilVfNO54LR72l6hA/O1aVIDxbxlzclMryMKCm44OuSRd+0BKIj92YcjlkbGfP
zsYsJigLJlFaovBNFg3v74zTb6x/G1SsXHkhqvg2vezOIALKXg+CTqxV0AlpsNL+
yum/3D1nAhT1BvJgkHl/fb4tYYPsaDVKvbGe6JvFF2Eu8RC8yzBF+LPzXlbflpa/
WC/uir00z8k6KE/TaNQUwJbDtuHXdTxVLhCozi6IHNsUj1m52Cymny2hc2BoAgda
LtSyDvT+1/KAoM4hQRycMS1LQridOrw/DZ+nRblcaglMRwzLwkZdOGQM5t6OW6ad
5gk9FYuiW+eRrQDDO3l4X8NfEF27qkDkYDMZIX4xXJLzDCGLxEK0KWJJChJMB8Z4
mDB+e7gn7Yh9Jhwsz8kKd5UbBh1xPecsC0sr6E/nG/cPXeJvrJq28KXo/s3TBv4Z
RABGFu3o0AbrNemShuUq1cVHTmrRoWMogdmfdOahJtYyW9yVvO4l03ACpzdnwd8I
6ksfCwaoLgjIJOm+6no9GHGFvd1T+ValB388d6d7Fr+h2APWw47FGhZyIknbgCPw
45hSdQwVd7xkx5yxjfZR8kqcPPhNVTMB81SGr8ZBDI/Qg4i3ChnqKy5tMNctNFJe
iaNAKhAsIvrvnGjK9SSUO1QbmlxxhuuB4d4hEboLPOtfD7+IrQMibuGX6HJFsvZM
4lpcmX40RqKKcBMMe7rfhmzJmn9rgdd5BNNSTlcn8rt5k2dmtAKN4rOXMea2q/Yw
dK97ZiUTlnV5eRzk3h73R0ExZiWRArF0+fKageSUTGgyLpxQfsYCFbssBpyWcnIT
bR7HiPQR04kxCVwMRV8SKS4kHtIGRBqeoG0+dR6xEY3Z+SlT4tZholLS9Mb5ngWC
Iuh8sh0qRQxNMZyt3IuFfoh1IO1hxxkLsy1TV5i+jj6/9Ml8XLnqXXtHXnKVjrH3
jjuujzmExLfJjzUvLwzwRqBy2NDNzDzz1moUQ/bAwesj4nRfmuhQlD7/L8cjukff
1Kqwu3aoe0LA6xo1cB9VCQ3sGtTTW+wLSg+3g1caF2JdI3xG8N6CAQcGNvRDUFHS
sLl6P7p0WjPf+rGMui04gSqKxcF2oZ6Dd71IyByoOgVSXySO55itOWnf0PGBuAh3
50mxMHAt+xLzy5oWAJxStc2XenmQybLf3vn8LX3o4csuXHJIGp8alZEbwmL1fph8
8ND3iUE6iliV04xnZIVowjRtc+AM8/HXif9eAPyz/NHtP+slvR2hAQu+C8O2OMUB
WoIynLOAv4S+X5IVJN1kVkPLfs1Op3Q6TghhLbnC5Mdmp66Dz8BU9m8nNKO6Be+2
5jAP5fddzu6j9zyAlaz+9Z7RYosoSITilL8BhvWNVCcww/ZpgEYMOHXi2efVrSnV
PPJHUkGWDcdt8BlT6TYIev+plRCZWdCN8pllxQJ8ZCO09z9u20dRQfbuTYSt/qUa
4HKEsa3Fb017ZeJvb2E8rIsgpr7UnmdIeWYFDt5Ely84OSq7XNH0JOVZZoPFjRfE
Ok0daxe00PrlmWjhFWd6klsp5cqgt3v4n9bKnV3/Io6c1bvl0v+0Bp3th87nEGPO
SJTLoDpHbwaGWxGNizenxp6hvgnQxTENvhUlSPKTxTCEpSxqbhAFGP2eskiGcvlm
u+4/pKmIe4vTXRvWSzZbRkPc67Ar76MFvThE5y0idk5J6iFfoy/5A0hm3P2maxMX
YpnsUmbmYo5GMRwL1klg5dAlMqmNN9cyq4olkk2MDGgd/BZ6dwL878GjMu/IhSQr
TbqywwCf5twS45z4+GPmmKzOlOsovQ10jV703uQVQbiyxKNqVFLdv3n8N2FbJqA/
WCavO4BL2GitUsz7PgLEKgiT+49Wqj2m8JFQqmuHy36kHotBpzQpYa8mtFI289km
Klt7zN8ven0V9EXT4zGYQrAA4Mz+X//kyVcXk+EckLRxxGmoHDc3gpcEkS7uVusf
PT/mUautWQkwg7hZ2gPVjq04P9tktegqF4US5jYyObec9PtHUNw7cB/8dgvdlEqe
c7cYYe8v+LRTD7Bg2fPl6XJUk+f/Bzn8MyFl2LVNSRXecxxhcnTVZt6ZRKjFLwrD
SuHlUoNoDxw8Pu/JkJH6QGAAR4NZGBFyWMq1nN1PZ0AabWOCH+VJUpbCc8UdBFI/
Bb9HO5p431U+ieti/n3nZjcpGh2qhJr4iB8kxNFikanbx7t2niM46DhrqaaHulWI
L4N+WM7X60AE6Of8/c6N2Cmy8R5pP32/vucOklnq9i2MXW7Vu7DpSk7qcAZ9ZzlV
oAuYaBEoPXA65tcLMQmbLcV6pYqgIJxbt5v85oKmCuqMCQSnG0LwMMJJC6oyf7J7
8WXR6H1O1euF5KfTFEjsyCQPPeb4cQoijJKxgotYCX7gGb4guPDmfKhO3WRKQcMU
CVCFuKSoxqImeBlcSTBCEiv+Z8NbTtrIkm3gDrWFvCzKACnJrCD1g622+ZrzmwHx
+qqcZ4yfDvQqD5aI+TmskMajWAebKuBKoLquNU5v1h6G3Ri1wmc5xgCjZWVbjbIX
PS75GuXlTJZTrBgnBjbnlRwoHPa0wYHUNn8NrxgMfgViudcgyewYiMFX12HhXQyb
HcJ5UCx5s9Slpe0AJj8E2xohaR2Fv7v00XHUf1H3v6NpSlJb7TDF5TJW/zRj5rEf
pKf2DWtWHXKmHBCEpLrot8JQ4zEaVq20iF0kP2+KAi4b25llJzjYnj8xa1e5988K
aJMqfMqjAimId3Gefc+eYBtHTioTyEFBcJW3Wb1An3IP71nVXIBgomOWS5fV6hnh
KSIVa/S0axA/6vwtBU+DFVC8hblVwhCzkwok0vpmyohvSKjCEQQ3EkQ7lphL0nVo
rpAk7WARN6e9s1kgeKie7iWbTNsvKWwmvC/eYfv6+jLaTYeb7JhN7GNcrjIbvuuK
RDzyJd5EfG8iWw6eI11T68obvVbFyLBJ+y281hdLGIfI6rBe1eyLlXy177uswQp7
Ll+TpniZSa3jWlCH8RqNOuwQnsXBodGb2wOmf81IaQnEnyC48v1hRTVtfulSe19a
CF6xP3A9b7LY0mV+yV4PXRoDcI31NuYq+DiWJGRMigPidav40w/LTVk9CeHApIh0
u+al5kr285x1FgwgrtlkOp8ejoLO/AqrjmCgQPC3cxnylu3R/AXl4HEykitVyElA
FzIb35eIcDL/+J2MSa18TWxAs/C8tfSmZ/+nkStlcsF6QXU8nwOtSdwfcaNNqXjR
444fwm9L5e6yKsIFMrXdArfp4SGQQQEReJGz6bB0RJqmkCGALO3SkGxxC8yMVbDo
N6nuPEVnnD70paCMtZZldvY2MLU1Dduf+aq0hvBi7u7gj5xLPlgqJom9pc99XGVy
TJAMg/SH2Hws//5DpD7TfMYyNE0+v7UjN4WKKkqt0/fWPlYsJrv3tBAv0bZsmKRY
kOakau6SM6Yr1oMGnqqInRUY2vOdZOCZ9KSOi6uJ57N68SpjXuy+RT+2o4f8g5p8
Od+nznGbNKn8hpo2htxBUjBHKtvA2VseXlsYtqWysDq+AQHN77xdrcIHRCv15tl+
yhtiuMQGteUIx0GTsDs65ka+gyKptTt/kx5qGrNseCCyA/y0WZYp2RY+wVoGsXbi
21if3GBYhQc6JdU1W+WaqvZqq8dt6YfGi3afolRI++Rrj111mSzyYsY64YdYHnGx
7CY7sHPxauhCQBbgzBadi/HQs6d/mRwx3ZnguP1A3Ao8Vr5ltPcCuKwl6nnGEeY9
MVoLL+Oni8Z4uThJJojoSCGWdVnCY0l66k057A4EERMxCj6TIT7Nxrm+z8+T+M3x
T4xLTLF1gu2UZqDiKiWTHi2OtNbaedESCZkP99u7jicT+0sf/lQ5ZJ1m6X0PIzKM
w7QPN+R8Qh0ZuKp/0FIU5SXzig7ALWgAfPve+Ab8x6TsuTfaqVh1htLrMdpehmEa
E3GYWK+nO2LtB0cDIc3Oqack3qL7lVABdw+iMYaHK5LSPgXt9o2DzEj403l0Zb0V
0D+r6p0eBqKl4J0DSGmGTXtIolnId8TtDlLnqsjMhRm/SRi8wL2p/J4sxk4gdXcY
GsziLdaUX5dD/m/Gph4diFA2eKFJivbMG8XGwMH3zHurSk7uenFez6fbUJ90Pndz
Xt7qaKn4rpgt0u+O2Eke0jJTxSoC9pUaqHORKi3HSYx+0MoWg2AQm6RRWnImmPYM
dsIGaAfE0F+SiZuAHKP+1XEchBF+hp8ba+evgnSdWLceyZuJoi0k/ZN/SYKb9rE9
O3S0klho76Le358E+gTfQ/wWkcVyKkl8qRHr4eZwFDJAVeYUdQdYtfs4RT7ithgT
ouO1IAJ0ni3EqrilZF2KhZ5zOoBwCXAHUw5FuBeMKaCI3+VR/qpIx+i3iYxHwSOK
7MyyMUHp2vNGId1FAOGm92G+oKJcstbbGXVz/x3SKLrqDzSJgo9KiGY1zNBpVCzW
c5t1dIOcbGKvoDCpXI14xxK5tE8Q5c+jeFjPacXVeIYCPmyAdiNuUv9Hs4uTW9az
i+I0ZCKFh8gmIOqO0sVan8c6bU3WY2rf7QI+e2pmPw2img7GhzpHbubd5w9yZsfu
68hJXAMGIO7o7/fEkaMqwUx4xBObyQpsF3mhBFwcBnRfpLbLYXUazxccDTz7Uj0X
dE6sEnilnu7DgEB2i4QZFVZ/wPxZeBU/851M0VbCi1NkctG2e69JUBjDqFp1rWLm
SWLhxCNkccZZQe3Ml4LNGuxMvdd2qA2qoApz6UCEC8rNIBJKrn9rIwmOppbVvfFb
fqHzdYanPuCL8QieDKxOjBT6zQclmQzHHzDamCWwYBPmerxoQby5sdx1lWAcx4P7
amFjAGoxYE+Dy98AXu4USOJGTMlb3uu8ZOrju1r3vZ5yncETQeH9ZDau9vVMaFrt
yECdVBIFvVqS5KWpe7b7hGzxul9tUYqD25FSYe9XfaEzQbI7/7ZGxusuVfPr0zHX
gmc9EWI4kM8G0heo2OBMJCV5QJuEm9rJ2ZJ8Mp8mg9rZQPiJAqxR9DEB68+DnSro
XqRHTU5d2qzpig3UpH9rtkzXBAW1SxBFR5yj78bg6lKR5EysPUL8DK/fVB6YYXep
vgY4Vt1k27LRfO4wFtAH5DmZtpXSb5Zy6GpfbPUg6GBqL6ewEHyGjdcuKk4ZjvHX
GEWOpgQR10whM3nQ0a+ek4FYwsahSdMFDgaYGHyYdekZVaDC2fetxNv8muyGhLVa
XsWV4TYNIDgk2F1nG6Z/a+lSTAB9IClqRxhCKP1YsoKBL/wsPAFOYHVpepxCqrKb
x9n5F/xrYQH126B9bma68Ks+e0jCYo+Ton/pVoUxnXei4LIeAUCp7mxDVpHLGKiR
UlgPdSU9Yru8vNEOESU9vIEATTHyxl+DdW8wiHlYo+cRYdfIpfIUglvJeZJuUndJ
aPb2fyI9YPx/VDMmyPwaAxTB5DIB4fwayiwfh5cIcnRKAS3dsDA7Ifrxi1LxBrdk
EiY4VcvzBvx/Ee5S/VBbjCVICXkSTargX8nY6KMK/ODdN41Xa9gf0X8x+IC++Qhi
phDauNOR4cJ1yQSPV3kR2jFW2orCMG0iTkixaX8pc+Tax2+bq9GXUCteB0QnTtAV
IbUd1QnzPJPlF7Q3tuYle4B9WO79C91CoCpOJ802MTvURTMxsg1z38wp+KL1yiIt
nkpaMV4VhF/ae1Z6nRZOfoV/NvmjsvncjG10L2HvoyXWAjigIiG0yFBgm0aA3a6Q
rW+YCtvyU2d++NGPxe0AtrDEsW83eBmPMChOq4+3PZsZ/ugBDo2dUcT7LjFYuDkm
CFm6sdKpt3g4H70CvaXblC4dMwK3tVD3mHpRN0v7rqCoDqZ3oEtCEdpxfJwUAJ2x
F7lLpWtZEzVGQl4c/74Z9s8rQ5m5OrHsW5SpZvM+H8IygMFxQ3qtQwZx0elSZnuS
geAJBfvftSeLkhvFC70gH1srUOM1haePt4toDYMc7D1WLgNRTBjjUgBWGdn9m58p
bLs2eK3QQ9cErrLLq5KHNXUxEJdVyrEPjFerUwhDOte+ctGJXIy7S/HC9ouTAYl6
JAM9YCzdmDLukyFpltVTjm7GGpo7crHsx1PpcXQs2W4jlelZKn4YVLWnLWagWMBG
WBPYT9skfTb1MqxgxMe0nM6ZSR8mYJrQwcX7OYSnU1ratO3hFft9wR7NXsV6HItn
1elUaJrw2VjITfNTOEhQ+iZYZa6EhI/A70JYEhqhXoYXw5BCMFWhD6a+Y5v6K0lv
fE5wTTJzybSkn0gkainCRcI77wfVLvRHXXwoEy50Qq2/EG4364yECzI2ydKujQFn
bicy6tlf1LC5BDmDkmIHhUsSAY8IpStNVG0u336ryHulbyoATx03qCpd1ppxjQsX
5WtdFOH/S7lg+vYJNS8thWPclP/kCgplIHC2cj2ZGFP0x0qKHDg+NXkB+1L7PW/r
vg7kFJI9zEMRuAjgJjnifNK4LJ83epZQ+QLToEkBK+FficmTancDmInM7lrtNuEo
X5Q8apa8gBoElXOFYXeZS2+/JvSeWEPoLTtmu/14TGAvXiltYRguGr+doStpSy4d
yNbbPpsAx/AO+zk1TTo5WtQCbZjAggmY4dMDTPoohktYvH4cNj/WrdQq2+oix/nj
51MNaOYqam0w1YqxVC/MBjkkcG81ZVh+e+HuVaqQNxeQHpl8S3UUzQcfxxsU1hKg
Tsa7oVi3vhUbn9v15oSjhAMFCD5iybiLf8U+lHEmJcC4vY1drJdGTvUsjGxUxjc5
CGQhQ38JN3X7PpvuPcTHQKexblYFXANXu3BkBcC0oprnaUtXfaNIqfZP0nDCCvXd
6/ebqmi+Q13DmBLGvaVq+JyED6sTvy487Yx5AG8aVamM8paJ6You+zvxlDpgLRS9
Zj1T4zuTSCWDEPMlHqAQc2ycZM4KQrJiylfyVtK4BYEaz/CNzsQTyGIACdiRWql2
IsQ4BqUrTicE+NOHlnZpc1mUSe0eP/aPkdyOa3huy0gzIBl3ScUx6645LzZhDx0j
uJgLfLdI9ka3mcWeMYjkz9t8KUW/t75ZjvQI/eRn2Rdgi5njORidhDZyOWVrkrn5
tLWFTFQv/KszEn54EpXTR+hxnorrh+mtp4W4QAAr82BDeXRBiWDFkJO5KK3NvRP9
Ub8w7rXEzjRxE89V9tvL6X/i0R0VlUzue6nbQcSTXG0GWcf3GotesuddyscAqA2x
A1nA013OIJTdkU62ZHp+faBkTK3C4VVhYGBivVR9V6tJ0jkv2BGlgRqNgsYCS9s2
YT9/l3fT4gfFir7DnmFbXLGqMjFA/g6SCo1V27C2tmue/n5eyfypJmkvP7feyJls
Q0cKUFKIV9aOYjvjM8qZ01jZZdUlZX19emn+6Vc7o1NZ1ZsOCaK8JBOh9VTrFcUw
yxTkkylWTmCX19wGTWRezPOclmvkkC6Vru5NNYRsFzNCXahpWyr/QcEmfpJS3Eqy
lr4oxBmhjoGfDCxDYDLAmBE6ObM2kPrevbRTGfTrlB0AqPljfj5rHdREcF6O/8He
QdzdHFcqputyNjWrxRMfKpbJo/VJUIR6tNvBbaL37X5d38YGw69FrUmArJfmxsSk
H348SC39YQGpkT4gIEn1LpuJBloMnw3yqJUhUWldYqnI4BKxrAz7t9lkcPtSeamn
MZLdJFuAgX/oQQSt3xnuAkYcJ1dYzfes+52BPLYALWsPxmeqAtWo1ihZI6ou66tY
24Yuc4JRjSUwr6uVgNsjtmccFSftANJGNhvdD6Rm6zE/f9NEIg4y7CcH+wfdSBTn
Q2hvmroe3j/6QZyJAryWAHndyjnJArfupalNebTNlcC2QABOlxNNuMVgH1yl3atf
aoY558TybCkZlK864soZpgnOnOxFBgGWg10wkItVahcutDbZc3NYoR0KFFCkSENf
c+QUpnKyM4tMj27fxIGDEGTSwU8ZbcUNetmSmvpqS8FuoyXqPm/YmxxQGp5u8z5/
ld0EFWldtsp//jUjAmM6G6aPrt1d77OqMSSKFHx6GuOMuXk5KGX2etlByaWoqgRA
SgE3Ud/Y+GH59r3Uh8ZwgoGZQhhdhoIK3AIEUSFxfglW7qO86mDB/mRckIjVFGMh
C7edRAAN3QCq7ds4BRm2oP14Mtph6Ug0gwG6DFs9BaR6srY9QDR+xRYAtCk7W4MS
b3Zr+AOXY2fnYAgkIYSezfNkOL1jsOGzNXqg65FwWF63k34Yxe2K5bN9/96kbLnq
unG2I8vtJpUKVzaXhMxP5d4Y0U349mhoRzDiMz23kTQ6UKSRvl2ubZ/GM+NHEqsK
B9BBrKPM79yJfaedR8WebMe+pajBeGty3unDK+GecHUJETNUU6KLkh/3Dt9Z6Hnu
WAvLWG5poq0a62ciBQ7pfhOC79ZrT0SHpxGyK78z1fSx7jo0w2CvG8U46UQnGb4Z
2j2IahWlMWSy7xJnx3ya+xmiASKS0bqtXu8c54vQpcN6bNFGqr0GWCmvlh8dFcoE
Lmrt+yqht+FOvHVwEKMweXH8pCr494iOPKLSfWUTEDhj0ivURXmI+7YDNEKbgjpX
CerxLF/ibBDjWVAGvuq6FT/3vE5/OShjv63ekT4WZtPhaM/XBXAGyGR/PY7Q8PPH
SxUzCZWfAKxnxsStpzFr89nJhL9AoKx0/6AapKEERotBEibvSSszqr3jNZ/dAHQg
5DA/uxju5CFF6vIEzyz7W5heDGhTQuDCvorAEJGdNeLTf+xj3gtV9RlsmupnKAOo
3XrJy4cJ2W8sqisld4Q4Snn5Lo9/o7h4tMoRsX/aaihbIxxSrauUlf4MVHLCDVHG
iwBopEntb0D7oPz6aorLYZUpBSMllbtykek0yp0nTx7DyWMz2iAiwlDznF6ZMKUZ
LNSVSrAkHEm/jjDLfMOaWFzWBhV/AQMCV3tyiLiFOqUjk01kpcbFG0kGM63Bei+y
b5HhXkMP9imfT1kRSx+eEPqgaNL00k0je1u8L7GsP26OXnA62yLeXxV6+rsO4wrX
tHw6BiwbICooQCbJrotzbDpy9Jq+iLcX/1jGol3K5Qp/uzs7FR7/la9/LX6gDisN
SReCXcDphuMtkzF4JPE8L3SNcg0RstAXesukbwmAp9eZyhn3c6OUQWHaV3ExMK/W
cP657GwIbxNRxVzzoasalidzBgGUxwE7+U5IGTMsraDf42/YaPQDLOrzcPulskh8
4b0C9voRF+zg8zTdzQQuuG7vFMC4K9qRJNGrdleGPctrxekqPmCBpQmsJZB/H+Bu
Vy5lOrSPFpPzy1rZA+2KXhJjxA34uhMivIrljHAqDyhxHDGUCiK8a3jAlpiT+yJa
SwIrLSyC0vK9A9hnqVsRckHBmqoI6zl535BKp5NkB60eDkno2ajBaa7GhAELClkd
WgrMNQu6cYU9Ng8V54nkGZFPda45wqyErymEc6/6O4Kg3iK6zUNvvYUupwD2Etnx
GDnnyFGJwlD+hjvuGDhipvVGGCNYWxzr7JdE8aJ+wmKkPTIT8DpZl2W0QySh9Ljr
EPF1Dz2mpn3x0ONK4PgRFpJytq1hVwnfyHZGTkob9wO3U6K00cw0hHpRjTDgdGff
p15KaD/Qq1BWRwdsZnqYwOE16B+ZKhMEQbW/L/ibEKPAGKoslskkOcvF9kkM+Dip
IVPNDN0ICgPOWGBeheXgMXZV6r7SWENgNz/9g8yZ0qK1GIw+JC69MQdtPOyMoOTs
LYsZ1EywMcA+jzhRiFjxCY/Ovqhr6vw4F0f9mXlMUfJCk/zSTFpxUczg95aGNDLV
YF3ivNdrTlQ1A6yhgdhDbVyzNjREij6+VSa1GdSM+z/wiD7DazTQt3vKzvScHFlN
uhYo3VJUu5AhQiFAv4l6EozLdvoEB9/QJKfNkiunKTcAqiNUDuSBljY0yk2SzkHl
JT49UcCtR65WNjHDig+oooT2xynUGP/KGv8iVtCidILRq2lz/C8+AmUVyMf5HCkQ
tKg6yynwgohUl6imJrybBWkknDsx82cgtwwaZEtaJh1OxB3CWUMLOqDTufb/6o/I
f7Ca1cu2QOInZ4gNStSDFXx/QuU9fj5QVzbiudDDxPRf4WCVuyve1lUvxCnrEEDL
v928BDK7qGGY97sO1psdZPpJDM3GdSnNDGCaW6Kz9iSJRbGQyaTN8+v8GplLbZvt
2KMs8Q7sL68w+niEvJ1to4nWnNVMWQiaDPLoZFEI0y8wvabXP90mWl+8XdWa8i0D
iCfEHWTB74hA8h/TEjgN+M8dWSPmFhiNGWeNyosMhd+OBIdCkFEW3qSjnN6BIJN+
rDTwTzuV2xO0g4dgnzGL7I0P89/Cay4cHkdr5Qn7Juzn4j1wYypW4/OThp6mMSpv
rga8SXiKTWpA+aeEwQFGR/cBuOE945a6eZgIgUis8ayYTFknblEiMYXN0B9e8mWn
8ky4l7t7SBrSV3nH3jiMjy/s78DrmOlriuC/QOPFxEDlG0Ry9ixHcnHauc/2Taym
9UApNypD+qjb3gt8nd+49H4P5iHC1hARyEyqd3f/9s5Vziu3ITf6NW9dagpaayET
mNDJKck6yck5BX1YNdnTiWyfgV/EQxx3QBRGUjna5WFtWS2/o9UCAJIDycEmrBJi
z3sN9Z5Q2bIWC2Synwa/5qNbLzwmyIiCqJImiaMo0AEHpycxYSsLiKMQj6LdqUX0
cZstndRTxnSMkbe3+SGQCg6EebN8MXjj9bBGxhO/VEeEekDnl4BDWmpTJaVixLL4
M2qtFPOZhbPCIhqDNICAs6GR6+qv2GFdBbP9vHA8w/DM+PcL5Nw7XdWoTKZlR2uE
hBRgQa3sNSmw+8g3k78T2X5nhohuL5fAmfmXwUvkZfLJXt+xLXLEkXKRY87v35GS
hYhC4qe020NjTUwAfiOuu+rqr8nlnm0cUfk/eClsJpU/J8nauSzx6ypbOIaYexg7
tPcfVC+qkUEK6pfOCusEoWxB1kXCe5P1dllUlulMZKhtaNruVurr4oB54GiW0spu
/gs54rh5AX5R20v6mMmz0Ena9XQrrKSpxc/HNKktrKifPHla40+tMBsyYrglKWLh
zpkbMsE7B2UR4aemwvMOLVGn41jAGUvJ+xw9gNSg59hCFFhbv+8a8LC2ez0WBygd
06KTK0PfjpGcDIcwFImUDAm/Ak9iVC1qAT2AsBmqRtqBWMS8kosyRVTsuLt5c7NW
XTBOCj5VpDxaHWG5lJAJ8pJ0ZbFM4e6TTN08pP23dtwmNlcMK361zjHiXn+T3LEZ
vjjy9l66+qq38X/734NbdwFVtEB0H6LoI5vLvfw6iMpcryKsMRSGZbKRo4PyfLV8
kcP+q26VjkvjZbeGwo+bXTj6qLkhCB7kRGZjxoLATbX0V9puT2iLzmcHK+0KWGnz
azyYjNhpr/4/TuOiE20M09eTQCMl6uOk5oL2p54LwBYP7y/XF3qvNYb6vohezAmw
pedxCg/GSM5NRuwK6BB/6rwo4VrP7TtuPOoqGVsuVUVMOI3G+TNOyrMuACQZx27t
hQT4AN7rcr64kN9o8QsZLr9pbXy+NylnECIQAwda/LDiz3hio+OmzIH6j/N33Kzr
45KvNN6vclCE3vArR5Zi8NtRAVZuuB7FbX4JbFJjKCpN+GuNik06hvKL3wQwOtY4
XWg6sOtJyGGFjjVdQMQvcZ3KrmvwkzjhU0lIiLhhL/iTJD9Ap7Vptzs5a5m9VRrh
/kh5U93Ac6RU6bcahc8djlGmvoLi084hbLmJAHgWRWBkqM46WHXKaEFF4Fdx5WMA
l4dcrj03HJ3LJW6iWsTgw+zwSKrU5VjQnuiGMQtdypptWJYYYq7uNb8KfwzNkYmG
AE1ftkkcvL3lB65tvZjO1N9FQ37bIrb/0U5sATx1Olo/ySsyeelPdph/6XKBEbTV
5JXYqfSe7Oh4XsYYj8e2yG2LzZQ2+xYzafva6gMwFBCi3w6TVWZ0A0U3tL+qKPGS
Mz2GizWb9vaHkwqPMvn0+6b5ydxg3egMprnXb+4ON1R4H6ncj8KBCFqej5UMYs7F
AMaoliMwNfRMOxMwoFfub/Bp64mMEWS+0zfJC75gmsP+mbtfDogteLAC1BoWLM1I
0/uGooe9di5v7+DkBP4ZeNGUXR2Z0HSBxU4ViR5DoR8brfOVBEF+5OTmfBDcgDe9
bcsmreOkJN+HuSBUWImolCTM45GwOaS7EcTCWiH9L6/8fVorjmZwxt6JlVaNUFO4
xjv/mfJNtF/vn4s7LwZRigvYxwsLuLRfnUrcEIGYnSTbch2aqnb1IKN06Nao1iRc
Ws0wso3oKAuFpOADtiF6/WTI+FYGLIPw521yJWlN9DpVC+vhC87T51rKHrrNJpxA
0dMMYEKP+EeZyZqAK/Ze8C7/GFQ9H6ZcTZd69PptNhdEqeSsvY3MBixtkSKz54sh
r30J0iaNGRDUDnBxZRGp87yhCwGZRoAVuZ6vNgDF9d5nnNNIJthuQzTPXTLmDmkV
GlhA2nAVkxKLX3Auu/ikbqUztER/D2NUEI9yIxx6aiapqn6y76e32H8DbAYTP6fO
DmS7Cmwe9pQfTyUu6opud+o7O4oumN6Ja0uQ39Kx2/bqMFxbEPCEeWM7x+3UhMeG
7lR8pHsvHtZO7so9mF/c19ENR15aszUmw7CQIUEwZdQT9FTw+THYpdLfZDbTDn7K
ftp7d/5MmdnD3LSQoRUDGRHmebOqjPE5xl4hlLsfHrtely7G4XFnyyPj1kQG+ujw
CbZ2JLgV+ZnJtAe54Lc1vMlWTM9Ufr3LVIdPuAPVwZpwXbGYM12RMcWxwCwVws7q
PvYixN+FuH3We037+sCISn1+coG1dOTMCnVSGHjrLL023PvQvgpu9b21oc8vZs0p
dRf7kIgC+OfDFaQ/5BT8qgYdNl3uEEPojEErMyGNhATee2D1N40k4qfp8EtFGdaF
JCdJ3kwhAblPbBQsio+v7atOS/KnZLCvaOs12q9q8tb2uMZvfr8di0nr9jPV4Grl
kXyhd7rsPWPR6gqF0Nbsql0hsZ9duf5eWnvWH4OTZr4csUXmRfJvT28V08eA8aZz
tqUDVgvM5l0JrsPyBxl5JGH0zTtr8VmlFJx1sFt4iflMU/X4KWxyHaoJvst+0art
W2yRodf+APLQuxgvjcj7XXAYxP75K6kKcO8q5S/3p8LEHO0nLxkj5DWEG+rs0jRE
HJOK+ZNovp8Ga5AtoN+ncc+NkdDIR9v1sM8ozOM8QJI7JzUrJb6ExGJqhpeWzcNq
XaA+Sn31KsUCPMy+jw6MMOfzDU/x6HAvKT8JDiqnC4MNwfY3fIzdrxvfKXGmIKa/
DRU3OCt0g7dSHLWjtADZI+Gj6/jWEEttfhyCYft7ygpw5s4P+SBnCloxatlP0i89
TUakDdMyCgKWSfCwti5wuPdTDmjXUaV2S+JwAQMPS01GKNt9Q6zSFLDFbfUgbEXA
Gsd2tIsU5RvSAO9S9ver+OzKrrxDLUAgTNvkKe0U7nvHsGWeU4L94vGZyxjMAp9E
FaJYa7WJlYZyvmaKYL0ljh+JmpyY7XE8+Lg+2ju8j5dWdgf5E63QucnSd+/AzHr4
+GCZzcDhqaCdX3l1q4BHW/G4YV7Y85ROMsfy6yW+kF1rWArKxhj4aKA7TV/B7hIg
455T98qXUa47pj2EWciV3oBUp0Re1fvH3BxtABCCq8Uu7I7b/uH++Y4pYnzTGwzn
iZy1K4Ioo9lImE1MOYI5eRuTFn+FG0jk7mI7/5soLkLojLCDGddoxEJBGk2NETfH
BPLZulTc1gIvL8vQKEfCZ5eK5D/I5YT5TBaC8l1l42JvH6VleI23S8l2iBMCUwBE
TrMENSVNaFqE4W1OCv0J8WJN7tr+JzdhJvxc/kv88vNb0eQS2iW2LCW6F9DpbmZd
UwPgJbhKlmC7iTT7BhwKRQfSvg0NyMcdC2x7oYKrBzm5lkXu9miH1JZOMwFqYnNH
48yzRfBzF/lXaMWBm8IbcJK4DASuOYv8u4tMBiarRRhnGJ18tpzIhbPtyG3xa71q
WLCvF0jOQmPtr9+GNtx3UFLIwbkDXVPUTQOOfwGtZFSwNzsY1+GvetzrQpoTr2PE
oT7Xqn1l7xfdgo72IpJloxDH+qihCRggAvorkqwh7uwZ9IgN6KSdwQdLFGjbyBqi
mtsK75CF7kTNVd3lKkoTPLqJN1AlKunZueMaANJsFiZXEgCRvgz9d0koshY6NC0D
cE6F9t3B/YaHckTTWI10xtsSgQAYdPpNlS+IeTh6fOavEkyEuwazNHEhS9p8m2oE
lQhlCp3/n55myJ1cV+7pjI8FHEmwkP65l+VrabTCTRFdyrmkKXpRoC0JoGIkcxPn
B6leHPo9wnWf93uXVHlrn8K73h+x3DjtIbESbuW6veF9kKw++h9SlMKpbkGSkCae
Ift/U+ttDu3yqSWgKWx5i1zq2g8dQzDJsejI6+ufLuagIEVz1ByUPatvg+MA+rnN
vu8p/rUfhFtR3yQdW+2UWZabOUVe6R7dQNtQ+ty1CFmFVBWNNLbmdIf2fQHXXlEr
5qVTXwzKJCRVX8OaPEmiYjziCcf15GrBt9y4VfM8JK0ADqbASGfIJ4ELBmjOcIsn
VVGvSKUVynN/kOrlnmSb9tWY+m1ACaVw1fABm9AIs9Ee7HYGpxXWnQthIzc8A9sd
cVbg+QSRq/Rz+JRSd9p+mtCWpnlKP+o6rNTDMz3eICHS3CYzOaYe4qMyfaqMG5We
fAPjXXwkEvBme221XYZko3mtx4zFAlhEzhhKITd73XqKExIaVurfcFCLD/tjUpo7
E29nrS+RpADJAWDnsAbkAXUZeQ0k4mLdlijKCfmZ3yaYy6ztS1T0TO1702L2sB2H
WyimBZgBDASUYNgKir/2aY0bbj+r8bW60P2O6zh7/leEpYyMVHw0iWzXnrQkienr
y+dLkHjdNMLXaNvYyi8Z8w7o3QR00xWZ7rLy7vioQVWMKajkrq5G3YyqiYuL16it
vsKS6SL3JlAGKh4jpverVyRp6BfsHwMEfpxlYo1fJluMLQzg10kXNRk14TybLpWp
3GN0I285BExBJpE8x/HLAV2sd/TEnD+ZlfiIKFf7KyBa1hLjFoAzEd8XRrNi6wUL
Ty9MyHg4yrL/HVAmdmOqRrEvO7PLk3GU4YB0Pgr8Nd6MNuNRGeuBkzamY2c5ohyK
DvY0K9U/5otcLgnkkQjhBE7XGFGutWK1H/HCAVgXMRjlpGjYt+ch2LsrkTrIhlzV
lwXSaIzg9uIFmOsoI+u29ygS8G58rfQmUjx2Mg2wePWa5iO9kVDr01zZswyrno64
P9hJll46WawvnI5kFMszjHs5eTHuKfu0DmBx70oXeyzGKISpKS2XGxPcmnB2cSTn
mwAmy06vxsyt+zXVgyQUAYouniymZ/geGIy34pwoC+80NNrj7FvBPUI3aPK+jaRa
aGvamuhsYNKwF6IWMBf9obMSRam9sCPWrN6xREh9SpLHce6fMdp/LyXh+h+ABqbj
HKAllQBVTOpjF66i6qn+f1kaItN8mamxyF4saq+tKxYYDtZK5AXKQKDKKuG1amWE
41DGu6CfQz/2evRow9pmSFvzjzer9WITArIw7Ea8p2irLdRMRmm+bTm32AD5aRn2
w/6fLLSVFYI4QJUgLPbQqU1CC1MvxsP8D+Lh0p0g1+a1QiTSNP4Ap5Q9RLsQadQ2
ox8fKoPNlWrcYgn2Rr3j8epknEH28amAmgnMXeaJq7HbiRee5jloBRompJ0IZCH8
3kadT64Hgg3RXHBMCSHRghULo1b1mhlolhqW6omI5kEljkp7qzPuAqWR5+JvFpWE
XBpCwJcvdJ+eVA6Vg3sWKAgtARsMpOnCyt8T7c4Uu72EVmeDjL2z0Bb8zk0dYcCr
CiaropqJcS8HR1YE1nscpRuOh2Mxp8dI61WRGjLZ+s1HhMf0emTloSpW7qhO6Mmh
5xemfLo7kMKe/YUUGQKqLFx+7i7O0yXlo7HH+xXQ5jjJUKBhyTvTpE9eFkL0fhYz
IBs3xqZwheTJvCcEFBfXLoAfS9uQGg64X/Uhp/4NGk2AppNAinFYWV3iA3IpbhqM
j4N0gPZ4LTALjfh02Dj8wZ5CctQaNajHKz6N8Nr+yxCXuWHveOmWo5xQRcxNxDb0
h1oFT+IFzNQc6I1y2mXnx2BkzyUQX77bmjpVdkuz6/ZbO6fha3Gzp18AxLsa5Q+y
AmMtes7W+WoVku3V7OSHtO6A4EAtPZq/HL44Kp4mKfCOxUAJqt2rLuYlihJCaiMK
DYcl4uYkaCTOqHglNb3kTzJMvhkG/XLugHB9E0xZbxuHPQlZDONGXjjVMdx+nyHD
F6JiNsJjYvEM61aXuB64yxUZR16AQykm/sH/ZAbXfjIYpnp76wdAhPTAnmVrv0lT
Mp5Pd9Z6Dj1RXyxkNhJLlZj0Xv7pLgzEIALSs7yCPMZnsQ16UXufG1wyARdn0FA9
thhHtWYu8uy9vYGFX8eMit87TuYGWFnMbiurvv6Tmw64977DPVT6yWUMJ4AyHcPg
e1L56/pl6dWHNCbQtvOXwOdm339LcU0QpWHD8SBJDgVCHixCnRk1L4HollEUUPul
d2/pbcQTyKL6dj78Li0KwoZR0B8IbNTQbgi1V7fmOZzDe1KXFHh6CdoxTlJqCPic
URcAVXCUkBeOhzKA911OYzHbHm/2FGLRMWwbPu7w1wXSYSyL4vgqe01RG1oa6+o+
VHZ6lVQfTot/3AJiIDHZ0ba1YFOwjazbonVEGsbEiJFvqyDuSqMLc82SUwhx0T8u
9cjIKymU5UcTHWvRj9M74PLO/aGoUF05sbvTiVk7wpC/QX6GCXpZiz5Md6ja/2SI
OM7acHOp1rSlt1cOMjYuw6H52tRq4kxggsSo6fLDBoueHKBAxs8Z6QX4pEQ0o4EV
ELuuSJV8YI1EsZ7KDs0ZJOh3Y8aX5oPwVv2xQsHrQLI1qyjAN7VUqDOKkyQHlryD
JfUlyWGF9KAXSlU3RtHosJ+RnIaIqxH1CzXxlawfU237uhcC7qbXtFEVd9QdpRG4
o5oml9x6UF29PHbUAgY3GSs6Fv7ZB+qCmAcRHXvO4RTaEXqw0dsRgFKJ0fDuLlPP
HTzYCeSWnOVEuXysHUf+dVeCPs1KLhJPjYbSAT8r5J2X29+U/Ry+x6prfsK8Gd31
uO7y1/o3K4Yd8TUyfcQBa1cXjnsr9mmnfB8IOlDjW+dIQLafcdy96PBCfzrI0xV1
HzKiJIobsTH6bP64oxG+F4g6PIaxIDBFdrLmwBn8YvTs5uRNyFkUxiLiwK6QuS46
HMM9sNtze9xQ6a7JlMSipg6pJevwdtF8R0IhETIlXkFSP+MHvbSKnwiaY8R14gFr
xSFOZ1gmaikySax04JX3g1afNs4+yY7BiLzw9V+l7lo+1nAWOCUaUlidsUI7IDhw
0DLCK6asHMPYAD4MTpZFjR0jKd+S4g0wPDUiMlwYt7s+78lNqVqjjRjS5wD5W1h9
IF341ncvMHnQ0AnaPgigJC/6rYwMMCxSWvQ6XK/QsMYgAEr4O3flO53r4WQ1XBmw
Xwe4ar+JXeLoZh5N+gXcd9qP5wrnWvt7Kzp8WFeSDSz3kXVRnwCsLACL+mrSNQG+
bN2rxfGzx9DVmVQl1YLxU5XAvm6BTmJjl0nIn9uEsuSunt8nJH8A3WQeGVrdEVWl
Zt1sXZyQzyTueRvTy0k1TqiEuylb37kj7zczvkMA5xNg7+6p/w8Kh1Ijlw4uHCo7
E/OXV+YrkM9PuhpwUc76bcB5zQDobUv5BJv7owxY4jcjTq6Kgm2Cl/rzyTmdJFMk
JGtmu97uTJfaeoBPVQCINrKCBgPo+rTBefyFJhnqJW2xwMAKJrcdDeP773frfHBO
591AOtnMLX2NdJdsdfp4tzJ4aYMcuZd1/LhpZ3FTwA/7Mk3EkvVPgMBqmvZsarRw
JuAGGHAE0/dvfDhHFuPrFN61s7+GrEVo3Ght2V8zAUHO+ojCa1v6/4/9EcmWapNy
c970X7kM4sDynJgnWFQb8A1k8wL5LY63+bOkatRgTWzXZhp+8p9XehrCZ2o7PIEm
TxJs4PXgdc6cdb6vu5tNMOu1t7br2YyNLsChzKP6+dBtGhl9J3ZFT/+0qDpR4oL0
c1yYBwGT3K7GOjR5kIiCEmu8scyALNBlvOjRIWEppYwzTqXnviAst+GBBg59xCl/
zwKKckSZS58H4UG4jWnV3FsxaEWO1SYTX4INQWlPg0iMH+TB9IapoL3DKbyVmlWg
L/nbm4f86jtpIgM5qrPUWxz4FgVlouilAd88/6Slbzc+ljWNw3Rv7CPW0tdyqR01
MDPwGYAU/d7uaqWMtDbSd4pkQpK6EecvNpQbIgPQe62VAuQNcVhFqtLRJML20ce6
54IRh2uyAWL74gsnupUuZRX8zfxPfTGyecDef/pfxz0TBOtsnODqGTPkaGubFaFS
e22wonvnJkMpOPB7CyEndIl0rovgwtIV0tGjc+x0pGpWX1dq9QMcDcjPWriktkRM
3uPVRKvWdgcMmkishj2+2FDgMtgYYEwJijcsyom01WAb55Hzel15SWeT6Kf6mfc1
zArAIeRRBESst2bishla4mss7Zo16qp4jqppkBN7tIrtM2M4mebVG6SyKjxgy7ku
4CXoTrOUXIH/p7gH+Or6peCtdI1sYOwZ2IXT5zIXbm7mv2K60ymymjqjU8D/OytR
t7+VwqYEI5BxDDcSQz2XZE0ghsoijDNtrt4qF1WTaJ9c19Jsz6RA1c2fZKszKu5c
xqSkYV/HzKVrrDl0hEL2ZydpmcEM1NYGcvxB7xAtKB3ZZhdIqCDdK3XWbEQHZntz
HJoauGMU+1prtHbozUyjPFugXjtwqZz1NeUvM3bzrZoTLaFXi+GUZShZCsQRA1xS
2BgfTEviHKm5driAKlSee6DUXlmLAlRSGzVMNXgfxTjDXn5wUHoTdw4bsC8arUZN
3prP7R59UW0Tk32TOR8ohp3rMKwQqq3mH1di7uSXp7LZtfBIfN1dSHR0BBzgm12k
8itJSoLqUKt64k0sat4Hi1jr185+5hVj5x7NI2GWfAEs9tA97sT/Lq+0Umf5CB8o
C0aVg4M6CoaCQGSQbvkkz1MSCV68+iIor9ai49N36fX5RAtipTE1yd3WPhudpwFV
u19pbeGm4dRlXx1mg7Kue0rMnzah+4KGkxlOdJ58UFNTWPxALzB2JYM9QxTXen++
WCJIw0kFYEFA83idIzxDz0Iy+nubOErUgGg4U6uD9le08+SGM5bi0R0Af9R83pd5
cmFA5jWGclN8LDmokmy7wozP17UfnPK92Mllow6ct0y68QxJCITwzOBO1F1trEef
qtwl8V9gKuglnBV1OMGrSV8qwHv1JP2fMgHJHi7rR9CXzWDK9lrBPYXz/FSnZNvS
Dt1eUFgWGtAlkO9u1k8RkZsvnx7j34ypkmC7pUZbiR81VlzsOoBdwGBFcJDIH7aQ
R5eq+1TayU6Di4hMMRvIM7nxtiY8dSzTUTJmSdYh709L1eALtjWLM0xr01pcCFaQ
TX//ONMmuZoZxna7rwJYhNlHop2hHiYXcUEo/XrUAdwve4xulidzbuqT9atTrKHu
btYKW7TrPfXBHP9wKBwRFuUw3gh7ehSJlGs8FAXplSNolaLp10vW5+rm4jk+3kPu
w9vHBLre0YdqU8S0ckJu4BKeNFOoX6xDTs22J+EaGEsf+2uih+ZkyfPYfzNV/q3N
ktjV75R/NRTEOVo7Q3xU8Fj3R7fpVaiEf2dlY6br7jGJEvwSfEH17vLGUkSLGlnX
jR5TS1FaaQvHIEwX++LkoIKxVo4OGlpsbyQBmg9nc0+kgMEoUGNurM9vZXB4KseT
ZPK9sYgisDhw7ay1/oKSoW6GRHDVM4ZRQOXXeS9SQcDGtE/ioCG69utrrl8BvE2u
xP6PblNbOj0L6/PbFu2JC3bCs8/PAFKQOHFp/6VtDX/sefW5aGKBOczd+7aApj+3
Na2Qy2pf+x58SttncdAs4xKvEz29mTB9a0pRwt5FJPjVZly3bERzp+eqhvmPZL4Y
DQZ3CzSiCZFe+55TKKp4NQrqR62Jxa7RAtpLqzt/n65BB5b569Miq07bLndwwsDd
jcijlvSK2OSb9X+Cz/rdkogWBBsd9uWAKlCRckthYkUDxhotWwVt1nyIIFVKfHSz
pHBjjY+4jpobD3obBw197VJgKjmB89Ks6Ycqj9kN1VOqkZPNs8CDObsuzFysjxWP
c3DgeuT/2lRgayHFwHPMrG+jj6Kmt3hcRzmWP6i0iCFFDuvxIPXfyVi9oii5msjc
dc+LZhXQQ2oDPD/4Icj+j9hisz4evv7uBzpzSPewQoYOC8Z6hc4oKDEbTAQ1qpZX
rCNsXgJFx+BBZykBV+4DF8P0F1+VIGCYIBCF5TUrA1fVzr5G6K8VZeHkjVy9bR15
rjJuJdNO20VPosKY42MOXyXsHkDXjIwnGeAg1OiymOLHzCP7+hP4FTR3EETAfGN1
Q7Fn3SriujV82V9u6sMT1/J8fMX38E9CXW7SI4Z220L2fcX7dCo76bZpE1pwgmh8
yA2XuDMSDof0kV/kvuS46z08jbVC4fOO7NZ5AcGdCUkSLPPURPF7tYpD5U0z0E3y
+tfDi37jGL4GraALPr6zYopK87WIES76qXwwzaHCgcV1qNPxCAQMJPqk4eD4+0yX
l0CdEgwVRZps5AMCxHHtAazScFo5N1VvvwgFa8jrFyEvjAs2hQSzVKDWb1RNJQxN
sRXSM5h7x0k6pHd9iZLjPx8DupHbsDGe7PO52T1osG1zhiBBO2yC4Wgm/rr6GdEN
dJ/5FlpeNNEsydGEcN7gMQZ2oh6n9iGjd7RrEUjq+mgMStUpu38xZM+ieTYK8wcL
fB7oZhn9pqPHk70PCrKGB3bqOmjFo7j8iMO200aO9sAZIN24N1nfBkDL0fMKVlaK
oUYSax2+BSkwd5Tib+3kyKa0r88GZj57ev2i1ejCaMI+/KO7Ws//NOvsEBtT8xF7
xe9RCERG3D8eJ9jw05P9iEF/XYHIIbZf1MWR0CSKa2BsVqzIrgXGamffYTLXY78g
76eofF8c1oFlDp1HomFf5PMqQvi5btDBUoI+r6VNv9iKu+1NmiVt9fYj0ErqI3Ep
acY+N179hUA2fEu7DFykEwZS8VCWBzV6MHwkYNJe/13TRUUqTFaLpm0ZYJZ72Zlc
ZFuqcq3ovs/+shtjRVr+lcp5I/5sSNOjMbLZa42WEg09tHAx1gEjqkseUN9Y4PEx
SB0NL111q+/9LW+MY/7cYE14lAxK0YCek//c8ETX4Iy2cZR/u2v4vA62HBh/UqnV
Pns78ffcdqWCAFWsXltS+2W5Er46+S4Th01VTGw9GIJ8M+kK48/DT8tu+2ovrAj9
h9WAuSmPCokSAFHy1VXCz4u8Q7hIp11st0ydNDk5YxlTbA5Z/8cLKMB90Ab5lVN/
CPLJg894bj+1YcwyxH/xetRgb0K0L0OfNu93DHNzHalq3POm9Uyhffpq9L3WkABg
WGqKxfwYj+C45LokivVKYH+OpMUl6FkVTCu5rlaMIKFxDcWCVEU1q2QEpQretMld
A+vd5CokqeRCSziv12ymxkgc6wf8rLewk2/S4f7POCuZj6w5pihIHZdSglW8buap
UWdpHWOvyChQPmkwdAjtGbrcEiO/B968YkZIGag0TsclvU/vNrGuselxIAl0kxTD
WKqNTbJDYQ9edJGERxovZrVv4UqoHi7d79jFMk3a24JFZV4uyHAdXNN93Ykb3emV
q/ucnNU/iehcq5WN0m6Sc3SOtwlwS6SV6xqFPgp90CmJNPa94RmdWrkX8M5lI+vl
JMDjEzYsMto0FitowbNQJjMJlK12ApU/a4nCQStYMzkD3gvO2lwZSe5oHcaq7PTF
KijU8WvgV04KrQ4lGFnbMLbgQzFNO2f3xJA152s/Vs64RrT7pzHoboPudtwcAvx1
B6QnJQUDAvdSdjvC+QjNJa7suLCo+jxqhaWku8SOoA3nqYjEVyezZKtFT1dPeB3G
J0ILWEvVeN7+6lJWYFPVdzzJLaAVJdQ1jAa1iuzOHwTGniZxlJUfMZlRzkw/uF9p
qANKexX9/D2hUO+aehvOfb8qqKb6kLGM7C4aXpN9TBJ9lxhOKhHxB/MJb+IKPY20
e1B4ubNlKMrDAHO0+H6s8iOlwRQ+TaquLCMsTo31F5bgzVFNDcWbmC2BLKKuvdrq
uVpQdsTzE/TURaDeYUNqekk/t5fiQpRVtdPT0ZuJezp/ZlP6rGjDTV0+vvfVoTij
yrs2C6oaSZZvrK9tsM/xXCjBF7jPjqt/iPi64YbBTt6D5Dm8R1jStgemhxYLpwj1
FFRN1yTV3Ms6O0DavJdr8WKk6x5LLlLQN0aOpDbd71RPNx0jbInKRHe2d6MhGBYI
WM/SnK6PMYwp5ikwV/XmGFTKVAHxMMrcBpY88qhqoo/TDLibDl6pTynG4WbkA1TE
AbIv0BCoZhk8ul1HprRiuVNnN0hcBZVdvmAoHee7j5s7qbx1Kn6thaSnMiJCdopz
wdYf2OSgF4+W8xS0XWyJ03ztLN980AXq4p+dzol91MF9y4AW02XUO+M1sXFf0ss+
su0FJYqaP8xwwIEt6lrWgIVIp/RG4NHONxweI1IgSsD+LZBzABpcdmujBC4N3sOH
c/r7MxoOzKUEF8Tsc1YMaLNwZH4xSrksMOPhd780XGv7rpwDWZKIP4jSBI7Rgdvg
B6erb1yF2u+qlHAXYO2cPa6/58oyJeiTjPtcpCElCwGyc/NfW78YEEhi9CbYTw41
BvBqcgxkr/iP9C2y962k4eV3UqpiNpnQ3FQF0QjSN4gNar+WPZzRAVyhV9msq4iZ
TNW9ghU3lTOT1Z/8+o2Ocs1yy1EeZ42v5gpDGfjko34ZEniy2/z7JaQHIV878mUw
aj42kQQBHznjlYtdz1ZcWi1AO76+ZWL03qjCFYrAf0RamQBW9dzkCRgzjpUuqvwG
jejj4KocYRVs1K1ZBmh/XccK+kwocQu4mpUM07603FCCL9ajuZfPbyws1CPh7xTZ
MiKXP9h20cQs1Xign8xM+pRaZ6iGaTurnbOIOqpcFU0/RApudE1wFHt/qZoE+nRf
nRScJpoM6fI3dgrue8D2AAjqtYwXlynJ8BtIvtGm85SMmeHg7rx/5CaMDEQlj3hG
hDEscmrXTMITvmeH7c2JLrdDx7RDmXIWCE7HQegnovDrCvUKEmq0AKvq1l4657fq
m4XYuGsIJ8YsK5iMeAFzJBPcBQFhvYJOcKmWk0hWCE3uyB755RhsSuOn5qXTvrz8
6iVrWYrDYF2RcbGBW4TD3CKEZ6FmTeyU4DIIhGKJLWxEoI2MSFWbzYojv0w8q/c6
MSYeknWOJokxo1xlIvWi+pMUZcR0k8woZEFx1GJRaBoQeCYko6CaeyWXAMexgG2G
PmnhE9MzMIGk7m9L3J3+YhHoFYjImhv1BKsQdMzN9ev3ZjI3RkVA42zWKOYOcxGO
wubvmZy21fMemZL3ivjruhr/ZPWapGwjsegwhLdxcSCPRwVbV+GuG1qoYPzk2hur
EfHtLH+Sc6kzPJ2fTVGT5iTjr8t+OQYtu1xv/i8vaB3j+RRBm0u1TV5rt6TaaNbr
fnai6ELhzrs0w1sy8rZPKNdtMHjbOj+q38oOhcrwESU5eATKAmGIrUY3/X55PgWJ
jlPY6P9kSQaI0Hm3c9Io8L70GSbgbnLkCtN9K865fg5peg9Nm5vqirnLF02Xj5ZW
BMs4il8jC9I6DgsiXOg/NIFcLQKPrSQr1C9OxegnK2r86nD+G8dZjCeqY+jd7J6Y
IJxB1CUjYWJz7NggV/Azm/VfRVq/i03klkDwRvvx5Tsr+OGXGe4q0Nb3xc3BhSX2
JBC0UXQDhuAK7ovcJcFCJRaDtxaWmJXLfKeYYvAI7eszz9pnaD6BhrW+jiUZ0eZP
vvPQHcGSVHgJVoxbVSt1eWj0xarbuoDkUf0rM6cb2xq3E6TYAv/OMByhhnUlI7Yi
dW8kEE76oQ2R/NVTlIywJAz2hGaa745OawACgYKC2h2c2merE/heK5RH29egw4ne
GhXPsCF/CJUQh0MaQ3jS4NncenkfCMgH+1+boOL3Op5fm1/IvPAVz92DNKhW1YUl
wp+mWUwxh1YXRyGZ6jmL0SQYm2dCcwpCA8caeARQHoKQqsQfG91K8+Wq6QJXYicr
EqN/vnVQ5J69qDaDUXsX+3OjFnGKAELVkjv/VQYqOBwgpU8aD6EYN21euKHod+Ng
nqjYBJiwmrTjksAWqEFciOKevSd9fI/S+J8kn/w4UFe343P9HGTYBQLW+c7KJP2U
2P/J+01JFD8dw6BfNKGBD/iE/UTBE9PQm4fd2GupImFZaiBhORuUiRosECC9vAKx
4Vs5e+Sv8cNKOZWyaJt2mQ/tJFzipJqKCFS6GhTD5dqFRTzKeT13hM9ttJZ1RGUP
aUbcz5Mq8Flr64sGLbOf5vGpDCMdfHEyrVB1ukM1i7nbdaR8vwX4b0Zl78HQt3q3
eN+p9m4EfGN2EQD5G05vyiUEAC2ELVGOsXDiLr4iB2cHn3Ik1Jpj/HJtQdcpbS/Q
cdDc4djYcKqwxtvXe4X8Bba1ze7Mew2n/fStjlg917tkGG5yS4HNKWfVl4/1Jgg0
4+F47+SCf6iYrZEXszwYCkmINwlif1sgbEp0Lqy5FaxTbCam8qTZT7gpFSXXNq9W
McvXHYRyYYuK5mxqqJuhYEC5Fqpei3yZqiRJAWflcn7A5aWeaV9H9ggImYLxpuB+
2sKCh9DFm8QMRAWGV5C3CMpM1fLdzdc7NTpjlh9ox3hrCas5vcgztr7TJJwblYi2
uiqRl33NiVtQUaADUV5d/47g2r0mT9KDbqKCLdGdqikssJMJOwbqdlpu1+DqIe+0
VT0WzlA5prch7+S2Or+HOS3iBj2xnDQMz5tX645CS9izNNslRq61d1G2DQ7H6sQ0
1Lvc6H7zWzjApqPLGG5t1f5wVOXsQ3aJoHs0rszqNITIkuLSPfK8Y2FQKdH+heej
mfDguA3gbcxDbMaNje00TDAHIFtalj2hpp1gJnAQZ8WTD/mXQGCqbaZ8AROpeA7Y
EzALIHB/DzZmFYNuAXu6Qh4P4ukwUWvowGloy2ynu+8efK7GSFZii/dxOpMLNjFw
NpiMLRJLPFT0/eArSJa3V0hbU3cenDrCJCIV6qQyZRyIt504iKmBM7cGax7/YRW9
wV3FuknSXuPDCYEZIoahdnFnbk2JDtvjDg+WjUPfTkrfpXNJd1GKn21t2JCT1wzv
skxnuTbZonNkdm3Q0Q58l5NKpDtm6SKDoz0sysRfa2eEW2CVdU64L/h+BVB/9BmN
uBCCtf1bxXn8Y9IlHc9xLWhWvA3f8+YENGvoO+SvgDsIK4j+50vIFintJZ2cS9mq
0ltdf4X8Tb7ra/NACNBCUSmHhH/FpMkuPbIaDOupDCBm1VAvpYbeWRWOfG1J8acH
9Y876TnFcZFFFV3ekA3cFqntdg0ZL4cSzisyv4lBCxRzpBKveT1Ue4ZbgzxJiaZc
hJcQnfULjOjrJZK4R0OXprAihcw5IBA9MpNElh7XLuRGf+D1Q1cJgaez0Kia2EPu
UJqRKBqECgp1t/VH3iYXPwQR9ddyb6uRC4mLvxWEAw3sulUKa+OCuRbLFuEbEBqi
P9X7xFiol4oHlvBD1VBCfDH3Mtt6JAgdIhPvHoTm8s5XI0lgvtoMvKi4gqN3cy0M
mxoTNnrum+802Pj+OCHYVJ4HndvAas+rgQQl9UfUpL9tNYWqBhSBoOAxm+aj7tdl
DFV8n6AdExtinU8naGQ/mX5hzKA1J14kRHqF0+m5BWBSOnzy9lKCSi7wUP395yDQ
yL5SxZr+xO4S6sBCDWlYfklQPTBmgSEY6bl18k3NIXa+dOqJUmvQNDueMx/SbYFF
RcXWSO//tshi5Tc9AegQwlDt8iGCs1GdUk3MHMQDwMv6NRFFhhYUhwQ4KT+wkdfB
SJEhnVwBq0HkuZb5hgg/jdG5fs98X52Rvmjg8lJhbWANuV2S+xF3ZkhHc3pzszCt
rbcHR2Y5usgdbG/SOAN4bI8AX7Fq26VQnBsb+vtd0ra5SwejmNquDlntbfs6QY6X
cqPosLwsfz0xcZmbUpavco5Onx45uYN6APIqFysZtycLfUdwyyMQI9BJKyA+7MqI
VY/TyMee9lzkXmkqf5D5l28Zvkqdf7SF1t15LIHzBgxGyy5prY52gxgYP0bpjxZu
hAghNiRq53jYZSjqqZ0rn3ocKPAcSBIQi1uRZ+dGnm9kWmPj6E//XPRzZnqRq/0O
nTdL9VqaLSeV+t6t8fRuIFt8aXa3NcVYvPWrkt5cwToS7SvhzVd8LFWcT3V++eS+
ptF/smgujpJevCsbYc28fMaqP0tlpNFDj/EtHi2Z70EceHKgw78RnEDHjeLyiyX6
DRFW6ADC2hMaYYf6frLxpwLNW9F8QDDF2I2lijadkIPxGG09n4lB1YC+2QoHMIra
kq70Dexxx+OyYU/n87anyRLqQnHxd/BSMh93ED7GI2+B2x2d4lPrfkB5c4Gtha38
UYp0Y5L+n2cfbU4iBpeg2JVOfviH/M+py2tADxURV5GffNj1GaIlT5dAAva7q8If
MMB5yTqr76fF+8jV9zTzdjc3QachTOIlLgnr4Qm1ciH0ZvDwSiiPIyvuofzGwyEr
UTKRtEpMwSf9pM4fLai5OHRQJNWLOOQOexklj/HgWAN7DBLiCxa0vAdn/jtqjGEF
4P4wHTocs0xjjXC+tfCpE962jlpm3jGOWmaGAGUbUs81qvDpVwbXP5cx8vEa8N/T
toFafXwJzo/WLKwiN8DnK7ctb3Kaytah4Lsnezw7NPkirXn/JSmELB3JuL6w0g9y
7ehiGaji2MMX8bndWoM3ZV76HA3C56iBWZkenyHmuEDX20r2tepeqyKefOqUKvcj
QAyv8YEXDsy+DmOtptxKKhtpmCN9VHgklSUeozdI2Zt5MTEHaBFZkb3oOAEVC9Pe
Z9Nns7qe3fWMoQWDEDO8Kg+vhbLkE1xrvo2ouWYy/1PpFyGWVCVzQ7/pMMiICk9P
VTrsaYiPoG5kaVgHUS5UM/BQbQgDTR0xOyw0u1T8xldpnq0BDALNHXqc0V9qtd0v
GX496f8sRzHTzkZ8XW+fyJbzUx3/0ig3qzqqS9htbY/KH9WvLWEXDHSmG1LBngEx
BAkRCRPQMWv8JXgxOMvxdojpGhI1Tfm5sWA63Qmdc2C0VCAWeW/0PQpwqjGyQs3R
PvnbGgT1dcACJA//otqREZNvJIAE9sJWC/DSeGAyI3M26sXGclyja/XS4Xsw5Nbr
mVRDFPC4FIWPuXzamELaVcIrclRKJ3r2XdLbC1JZjL43hvtWj85hSc+oYN/3Vcla
1B2lM/k2O9cItuoiFoZh4Hl2XjqJ4S69etV5ULCe11EFhEVc808FjDsWHnyHvC1M
mRQhFL9NjujfnNCUXDez8K2dIOkE2riFtF6maJjwqcvnKQLqG8IWgzPVRJ9y6BMW
/TKqpck4Mc25R5My5CiNogO86AZjdtgVfqT0+ZE32rofxigG7vAgNgpwZjCH4ugK
+G0iW4fUtcM56Bjk1odTuSo/tbnm2jn8Bev2dqHRTqQTyvn1nZkbrRgl4yVQiKsR
rm9AC6MmOHDxdDYmvX4qwOtcJTkTmU7araKWtNaxAgQSXY65Q4nSvMA5TbCFnLac
Ef9uaU5RsfLIKsAK1fvuh+e4x7sQmnJKUGh1YLGv9pn5cCTCE8/5+xTPOD8/F/vI
i91TDjSOZsvMzUsd+JyzNToKnboI0OSKZi0+7S1h6TMrBLqtAqM8rzynrHWRl3WJ
2PE2ckPJZKf6w4NlbW+vup5KHhS+dOA/x686kR1TmaN/RzO62SI6+CH5AEiKRBwK
53wMSh++eq7If8pMsVrPcsmTm1VGW0tJ4OLJ9dpn0tRk4NujwJqrDAN+pCXHi160
VRJCzlQigkGfpCY3d5p28I5CT+Vz436phxKp3ozafTEPDgiUun6+7AY53Vp1TDSF
M3jyvTA3ysDhDGk68EE1f5ktoDbBHu3anlyxxQMv8BX4WSM3lMMY4kbSyiyyywnb
/8iOc/oK2JdA06c1iMaITL9EMCmmLa1o800raqJnkWnkAi8QByz46dhqRVwwom52
Q0e9ogleaHxVDdsRd+TT3gvaJU/MXKHFzZODmKLD0sW1qpEG4NCReFHXKDmQAG+G
y4M6a/j7/jkPa2cfQXN/tHpna0jUwj+tcETGBgb7jQo24UK7uQj+cUcfMrUK6vka
8GQQGkb1aE4bUPOVTjjfVMQ2SpuQX7g4SNXeV3kCQve5HlFqHsmwmK33zx1sblRV
9Q+mxO+0DJrf3YtYEP5labgN8zniCY77gmkAoIUrcv87qMBhYVk7BUDB3gbOEvV1
V9QNoINOEanuwdYWPec7CcXrEzMk9N1Va6XpFb5oEcPnp3g7ZAvJ1uH8go8/OTgF
OxGMu2Isv0BWfAEKDiXwSR83KYKOOe+WnqbNQujdbxI1vnIQ8e8vsqJ6ldbSj3Ln
1/Fmx1VIheZuroQUCXUQoSNaaXWWQgMIUVDU2UQbNyMilda3TEIGv0rzbagJVHI9
senaz8mT8yHg+hPnSIFP3cWY9ezn4el4Rnma39O+o8ACLAFlVdDt5Z13CfFuKvu1
UeLckM0XzjNrVexsnFy6rWpxRmq7swqoGpQXdaMjr9aMsg/MoF6Lwdt8T/EN4SYi
9oKRDV7IekIMU/+do0t2Gz3A+dnDg4ZBTJg8x3nnlRLuuW6KoCDxlBbh8cmp2dJu
hWDGxt0MbznROWWrIcttFsZrhGL4UVLBZH1GLlJKZF380QOXx3yWfkl5AtR1OJb1
GMGR/rtgQT4Vc5ZpzYcryK/KowUZeNNDP6NBPB4ePgALf86YG14G9Iys5crlsmIg
xPzdlKCV5CDOKBjadxlgUP6KfWPl0JXW3cC4/YdPad6qRHKCJAKBY4aNe5yVi2zZ
6++ygvExLqLy+hpdPKSudko6hvww3bVBTbSEWCWXC+qOEQsbQOMLmtjxKs1Dm5iQ
pIjCbnQ8umaTMNeukgyhY7aWLCBHT+FXoPN5uCP4gxVq3EzpYDTHo8aeSOnVEmbk
N8fHJ0V52POtRX/zHHm2Z/8ta7pm8X76MgVSTU1AlLbcytkuZZVlA0hRGmXP4053
SOuCLwyX0kIYhGUOdLqttP1iSywD0HWOpDaVSP78EiBeKg8AsZNFyD6JQwnHHwL3
DtQ8kmNVpIWdZ5b4IgDlK44tqsPe6N0MO04lZAbsGSuxwihbJ03TOu3tS85A0qbz
tvHwYz1SoMlGc2RQfjXJHB6jGLRHG2xqzR/Jus7L9ZfZrprfxKvUhJp4dWxCQd7o
Q2IKvb9kRR8ewBeormvw79n8bTtWHGDXu6Tn4svhQvMBbJW+G1R5eTTlMBnuDNki
egzrHJNDLXx5c0uiuUeZAGSr/pJ4MZOte2H8vb/pB6ZZytWaAn+4smWd3HeLiSY+
5S9/LXcLvL5jXpcSfSYWbZjrIGdurol9+C0Kakz5KZkz5wke70anD/Ntel8AjYOq
6Q1BNAcEKgmq3YhYFfRBz93cEsVUdqh+j5SNsRBXDaY3jHADuP9/Ppq3X5dCjB6F
AfGDmObsthZOV8VmIs6/kGU1Xi1WqBUtlU4UsjOrHzLQYcW57b5LdD+WyemKzfCn
qNpcDcS91i2erWuXWPELJyPAGsubzbla4mZQZewWGrgmeazzyRHe0X3l/2INEGRr
O6Ibb50ciBt9LbDgz9Oy+UeJJ54AvDPWuN8zOQDZgyaxY85vHZffsQol6Mo6V8BU
GPQFcUGY/T7YDxK+ZPu3bg/OJclHDONZkjIV6YoqmcPeCwizjzdIS+LtenCDQDlZ
8JY1rXLFIfgWTOUnef9Z+EHoicpVHXVhbIZXMuNY9WEkSUKGU2rRJbl+XLGNOy4L
FTZpH5IQsq+HOsYzkivsKOYDNCC86deXVsvVOesJs3PY/KiFe52oGp5XrQvR4eZa
kc7/hs8zfkecLuYUfuib6ayqfNNn7ymv2b/pHmlvqKb+wO1QhDKXc47FJns0iV84
1kLEZDrGK0co77FRCfwY1VDiVyMjuIKAdL+fp6PuH9P+oQsn+LZlkDGcJdXTSM6R
MUyDVtmtEfDh7nEddtVTv3+RLm08uzxrBmn2SLkbn69a+0nJoHD3kbw/gGPfPTxo
TwsjRfsKGVHA4gz732ioh4c4INaWUy5NvwDgXJ6ZdxW1dtmiBVir0M4TzhCUZlYC
GF9lDCdc570DDPgoyhdrgkaKJnvQth5q5dgl1nlEn3eYsUvD+J2Rs+MYhMU0A2Mw
+BsyXKHPJRz8NLLpetEEA9IBQD+ebBqxVskwMOuA/qpN6NDmHi6RNYLcl7SkbYUF
Zxvyipzae/klYpgt+5+r6LaUwvKqjy2sK8EdrPC5bYx2vmiJp09tNd9GvhKl8xP/
0jyOD8gGZc5/2MnKrZ0npDWP1V/b3aa8VNIBgfx0wGcFU1XtT4y4hyf2hFe4e2Ew
KCJIN6WuRfg2b7ufwjg0EEkfx3hFf1lLQ+9+smyetnByQqy/PaM8WxftGKvDXpPX
MYOS0RUxOyXK9iViCQ+rKBDzHmFBaShBo0YggWkOzxuRxPXNmd1ZfsUrRGKkmtBP
pyOyabPMMttm9xTk3cX/U49MN5VvSxFkFTP4+CGZMsEsjHhdKzp8sw9qeJEJ8wFf
pDNR0B1UY/dgMz9NYin8WITM8t9Ugz0u/aGqx7MAm68KKAxZoN2tCXKOqgo6TekB
H77B/7lxOT6P/lVda99DYyZ1Vmf4nX2YqVftITx+lUGO3CG0ToahBtMTs2S5GnYn
dmcRYRx0k3h2Uraz8DBpqE4a+7bZMqP7EX8xnxVM8rB5l7rCsPYvx5+Dc9fu2cxo
sK8HQ1A9uu5MJ0dFNrTVzTzf9sJxyKxI/s71itBTLle5wTtRuILDXc/SltPrcGKa
HqXQ62hRY99d7xrHCDiUi0T6G7CiIBziri3gsMTxHj+wK1AJzZHpUSQKbhxAqtn4
MlPb52F92LAK1XXMkvfVAN91i1IsLF02D0prCF0T2raSKzLussC7PTHqJixXLprW
uBFbHekI7m2KXrfV0hD/dvjBT82DDGm4AEBUBmimsM7fefq+YwAxxmkeRfYkUWaD
7fJkbRTLYuTNZoMyVMqxVzYRUZhmkRudK8ZCtKXutZwKFaL2GHY/o+eCEwiTMqlC
6irYrmpuaNTS+sJSGpHBo5z2upaKbinadm7gkNmjHuqvPN7QkT8ZOvHi0ngkoEW8
0+YM8w3ZiQAwtE03HavVFInsfeYCK8NPEKB8llm8c247nfj4XsdD4Bw3u7kLSMgp
NEcJFGvFOTo2qBqKo7bv6zI0K2/HKqYTKMH0hDhQcH+LmCVWqueRga8UZB36hQ42
vG0W69wlZ0vqMz0lydjY/7IvweXNvm6IqOv7SZ56OnxSfzfPHxKAlOy8jN46o6/b
LlsLlhRcBnRKjlhN3LFVxoMQEEAE6rlkPItfSW3NswqXsedPJM/v+VkzZi1MIPJs
QMKmKiyn1JJwB6AvxMkQp7IfOzYnB8dJJ1nPnWTiRe/HyVydl+Pe73uBPR9B6E06
MiHso3/5jCrLD6cUA6d8ntJGNj802XX9i9qoWO4d8NXhuwBfESAo3Glcj2TTRblr
8PhOs9hmCQ6CrEK+vf4BzdLL/OXogh/tYSovzbq9axLNB/XmPsbZ+er2pzK4tzl4
io7u0kQwnemexCoGn5D3e9MwlXwNZqkjSGI5hCO/bDc1r78AvCTyOyw2+h/eSkSi
0cRsw/pF8sH3+/PQ5y2ZEL/xDwhKNVwHoulHoG0KTtYrOT73uXYZ3bTzHPpK4MWx
OOfBUJZ8PixL1KuPm6ozEBWdczVMZ9CxLZseysOcST24Oz87MH2zk0ifsh5UAT60
mvbGBOHRTRuSVM28GoFInU6LOvOpjumgOIorKtInhpXapYKzUaGrwW0o6jA0GQrG
VKzZGD8sOWZK43LLcLGk4xJ7jRyIX+s8EiskPDHPcQbD5+DnlzkyywPM2VBkn4fI
t+GU7Hru9eo15WeOXJp1SeCTtNOLDrMHdV0xbJbA/kkkRw1qb1qCIsMsFnWuhHwC
hmCUbEx0prbrlinxD9a4vpS9DRgd0pndNAARtRKYWQ6JQWyMOKuf+Em1z2NGodE6
6WO4VZDjXgIQf7Xv+uIdIYn/y1JTIQSAFQsj1B0dCcIOjY6AvXmWYeS+XayMx5lo
7IPjfP/DPFbgrKghHcVC+oYnDC4pYelHEaC4It969XXXhv3rwRTLIz0C9kyqllkN
DGIojH81f7xpF2IPAbg6vvejw54R5lLKE4GP/QKQz7sDocXbDPzWEMhrpSAiqFEY
zaUpJlSZH5tE1tllHPgVAz/ckEfcXL+KV2FWrxPQJKGDS5bW2EewvzkNnZbn0e6Q
HlFvTw99nXF4OmSq7PB1ASja3T4HCc8cTa4dWQsAgdq1U1GsVLJnQn6lsdSECqsk
y8rWtPvbqIrN6yZlSqPxy+spB79sWcQXlEVxLHklxOg1rAYDMKUQ7SlNPYHwzAwx
2kkV3qbH7G0AQt9MSpcS8n4z/nRvAHHe3n66gQqNrnGbwWZOm/CGnfklSGVCsw0/
AIM/JtZy9oDeDsrLicsWlHMCwa3azdw77Q+1XPVc0XWIrEZL9b1gSbjlw4V8meIE
NfWX2GDDDoVLnwmF1A+uFBhyxUYoeudlsV36oL2U2jCSYwU9By66A4Zu6YIX+QkA
D2fUdIXtSbjv3CXSfjbvNbH6rqXE+3NV/9XolVICpCc4tMng99L6/3bfLqdnv6gR
RdcFC7oy75wXGSE42XL86D9/wtDmTZh9KnBRKS+GBfa7fJOhkDrecG6G153QouCK
zkl6eRZyernpo/DGSnxWegPTFoWqToSKw0A7KcYc74uCfHF0QnrYebuM2x1jNAzw
DrvNZIxpUm+TGL2/jfQytzh4CxTyDKNfiy2d0CcyfcjQLsnNkPnd9KRSeRP8JpoB
NI8R1QKaMC2uW/p7F0yKAmGgwEAzKDJ2WHlN5bD3szHeWOGdc0OQo1sOgDF+edmz
2cR0R2UEl5mH2nmM9fuG5hWb9PjyG8rfQz3p77ttpy/0gZ7itPqyMs2XeZQAO3sU
jqzN47ChI6Y07ToKgy59/pfhWkTb2yO8cstvAL4g52gQ8QKUyj9vu4/8kca7+ty5
hZJJw/61N9zCN8b6GLNBzOwqsVsswRTRXwbPlnmBesimA2RZXBrcjCd9ii8K/QJJ
7IwwwHgcaeRGgBCB5CYrqEG//GKcG07Vqk4PiXmqRJXMv4VuwknM9WI03cnSsFxX
JYm4/ZgGKmMAC95ywem78h+ZW/xlcSivShf3DFUXGEyxH3L1+ULwUAH1LQ7+ymvH
lPfv1OOWOSgahpiW69qy2BSFEujzFzB3fm9Pac2yUGw8gu3w9yS0b3ICWt4Hma1i
xK2QS7Lufafj/uxMRNuCzcBagF+/7SCwQGP+GWIzVHc3AoDOmBfMrhc/Gses1Qcd
/WnWfJOc7hifmxktANsUd76l5qD2y9BHsaJVowBzYWYGGrmVCp1QpFC0/No46cVP
5T4IrpbooJSHucZZ+I+FXnAdujIcauEOjoGMAjibO1OoUnnS2gq5ccUKKMk2y2l6
F5GAjcFw66cGZ5CtOj2j4Z5AJNoYmZqsNoaoODU/OFI889+X+PbBrfIBsAMBcl/f
CW1N0PR5+mVm0TLr4CN/UtX4jhPg8PyHoIgb/aqoiNEE9mzbRCx10Pc3/dZFklRX
geBlc5A5ZbO+Thl3rPW94HIjwQIT7aO6KEXI3Na1zlIEhdttlBcNBr9gsp71k3CD
imkOuO48WjydBnLUJnFo7KB8TzQTxy5kO5oMYVIB646gapsH0cpaGsfDBj+Ijgrp
1C1c3/sPAlmBp7g1pMgUA7M66NTD4cwxtGzMDVi0jgbYGt1Lr3d5fBp1Wn2jvJrx
8MOWFzGPDE5QGJmJTo8mKm9sJFHDdBCVOzXc7GNYtzLH+GNlKab4CyCaXq/JA953
ir4XSU6tK8dHPH2DZ3laHoqai3i4Y0oU+hsg3Zm6LCKJ2DZH8wGhyZsgfkmBJUes
N3C6+uDFRVuKbznwnR9AX8zWATdw0ez5XnwPcQvYjJqYo1THxko2DX3k0dUFRmBh
h5vx+o5X+EqaQJ6j4IUl+KQL0dkQ/MPKQwhG7DVrLCeOpXwUhtafwU7tCjyhiQTn
sZnbb1YNEzxfEyNUaT2zcxe86zQVl8EUxJ8STCi9RCEh8cWiuh1i3vfQmnV7cZN7
lf0y62YDXyXh+i0zEkFQvqAVfLanSp2+zovlmtxkzx/oIRCDwtQj0qfd1IkrWMA4
7Y6Jp5Y7UfmNXnKTtEQ4F012jwY/qJ39ty2pJPfbt2MhlY7BNnf+DiJ+hyVEfN5Z
AzTgmLDoeqEGRhrLjU8puz+xxlLRcV2yjSm4q/7+fcaXLg0LJX0Yiz6Xc7By87Wi
/vtUiIX8IIlA42vIxYEd1JWx1dHhtObtIL7p6TaDItDsL+pEosz5nuxEoHwn42KU
M6ApfF68xpB+2RkMMfKaO22N/e8VHbVT4Z2YWDIZTxLF4SDfIrpp14TCgvfJSj0q
5T26r70FrxoGCJZwjOiEl6isIXlbitZ3FljK6j684ydlmLLIzmse4dNO/AvLHGMt
awAlrN3BkrWHlc3N559OJkfqfpduLSm1h35BC5TuT62BfHOQsjA/3IijNu8Aa4sz
XhyUyFhDdBdufytoh7+CB+3fO/+R1q5PQGyX7LoiAbZGuf5fam2pdxgICFmvpoRw
nfvn9Kl+ROtT09vpcCnEOA5MKks+39o8MIjJ3L/BTIk1RUJjz9LkjOHIQMK4A6+E
UrVSJE5Un4qXXNNjhnXwq9RFduHu0L1PcMWKLYufTDCX5Lyotw1Jp8kaF2vEJHbi
0TL3z0fEIl4A7YEW/PQB1vj2+uIE24RsD0KVgVI5lXQGNa3/1abdkJ0AwlfTUcVC
H+DOMPbF9NGuUz/2i76pScU106NdLhzaJiAfoZFzCejGpPC5tBHvbK5uWsWftq04
R/BL/87ToI11tN3nn6FA4zieoJ+ZscEK3Wg07s0v2qheKc6YjXCJ639IS0b44OMw
HgwhmGapAgeQClrvg9XPLIEfTpz38FNfg8eqnujBNoEAqScYtbU0ILiQvQnYBcta
ILdGJOZG7HGIZnPbDnOBRb9TA0jLylp9i7RPXfEV4LE/evk/GsxaTXS40naDyu8R
MYc08WTwBclClUR72+NWP9wUpgqYkm8weBWDkEDLgBQuvIxbrqAeuDgLfcPlZ/+T
QszjLkOLecmPLX/BZpDM2IwXarZH4yDRT4fgZHqcDjLCijX51hR2nCnuUWPh2++W
fo63E9yNJ6dTkKjBadDLQNz/5HrtuMF66d5D1kpaite3lYsqik28mvYj60kf/uG2
xOoLXYrjljZUKcAGMMgNaapXSall91sEyPYU2RWJsl7svc8qmQ6R116fZC561Z3F
UzfJu7GLMuJP/GK3l8RayGg1SUZ3/QAo6GWux6bUOzeabdiJvSXQD/wbSuuVSObB
vhrkqZrXzSLjZEhqU0srRcBYdsg0q6+hG2nVmy2SmQMUBimzOUUZ/94cZxH8cSgi
/f54MeDCCk2ZIyK5eybwzRfwOAR/qQB2eAMtLJcNSDOs+FAhfyMukSKhbHEU4rw2
SiXNbcVgbQqMfauLqG4P+rQjg3nxaTl7qw4qAERrLYdD2ojza/MhLud2E1MNpZI/
kF6Ia2ovUHJAuj/GqOn1S8S5jEKdo6LVKStMTA3jUWRFQpp6w4bY0L/USbsggj45
MXxa5WpJlShvTwvWZrkno9whvtEPEoH29LP8uWDcndrd8WhXz7198rBYXioBohe3
CASayTmKefEhaViswUbUoObXW6ZgpDgN8Am3V8qHHjUjXMobsB9aaKG9WYyjfizP
uHXno8HO5byNFC7ROK2ouf2AVcf9IsrkF8c9k1Xxw0VUbaHMt4aT5GxOYrOKma5n
YtQCnBzZpEWfEU46TwYgz8fdkTrc3c7lRfmRZQF+I8uxs3oSTFVSbg9SYFJUPbaM
bvTewp8+NWhsXInM1a+t9zchigauDWw4lilyDNngQl/qjyvrwvfdKD1FpavC3KlP
2J2IQYM0axtLXShUeLWb8N8WWjmSQY83vlLNFAp6/rJXi3Ng4XyBNzKUD4YnbFrU
fX0AC2AhNixcwFwAvgfsEzDTLRSUC6XAQui1IEbcAL6yNEDzM+Wu4wUd97xLek4Y
B6ze+H0hHHgChI4NVkYsM1zdcgZqiO+du1syCGoNabcUF/evrhXb0RooYafUhGKR
OwIWqjKxskW2CeG1+J5eLziJUuo7zNx3tAAMeQ5cvOO/FwmNfCr0vSm8DWGRJwYB
7+s3yA3kOSFnaaYTVKzb3EtkzZpb0GlUo+mZJ5AMcQoa7S/xCU9SKibT/2dkpkkD
LCJ5YmvaCcQcyLQQv/0vgsrCle2ZjleYMHj2U1GHDACO3mptD62960M3OTR3oA15
MjPDC6cCnTvhXgX5Wptvbs7DHr0jXlbvcWDGSyJZn5ufEJel5VvpM6tOnNcDpKcs
Zlpu3xbiHkIXAyaC4lOXPo97ON5oej2KInFiTEXR6uc2/1nXGCVtIsg2idUWKQFA
xFEvtprmrKs9fRfKjkW0+d11Vd5eqIi+Hk+w2YxlSZ1e0MQAKJuotxZgMI76yX/i
luShSDfiSJ9NtVojhe1eOQkXHn3Sz5Ly25BPzi1eiSKH/0YqIjqLnMNlD3IGp2rY
xG/PwVgU/oJi9PaYBdDygGp1Bt/PXpDGkV8RROaLA/Oqh4kBpuorn9Wge4N3S8q0
PKmeXM3wIbrjhKsJPH5dZr492OZA3aQxQDajZiQv6nBJa2lm9beMxtNkIxnbbTRC
nRdkMxdY9r+3g4/g92aazKwGuS4LQr5NF6Tty/CtD2puXS9rF1GXT+pM3/UIEzPn
5VtXirFaa8KniRzl/JCKT2ulrpuvNU5NBVLAAggxfq6jV7hf7RSDvkZK+NKBwa6u
yMz4TYZk4PiqhkuuqgXFW29oSKEBurZooE2eIDFsfrFWTRPdavaqAILT0jlwErtO
oNA8W0ecR6sf/0zDB/NEfDZ+yvxoYiL1TEQDHddICkr+kSHFyXCAcV78RXQ47ZmD
0HVExozI0VUMFKdGrasLea4JWMgz2+t69DmbR2Bwc9vFU0+bwOmEJVeGCHcnLpA4
JLJjqlylRDTwb6kd4PNh9KMdyCMYwhYZP+eSnCVAcpL+NkRr1XTPc1Zl+G4Z4vXS
ml2DQYvLQI2+v+qyM3PsshTAHGuAwq548i4Kcu7MjSpiomCMHRZnhRfJ2FZLOp56
dFiCwFspmrkbVRiAvXD9s35BzsN+HQ+dj2YgW0g6rXgvG2fflOnt+G3TuahcHTtm
alLsTZE2hpwTvz53Y3eiFhns5GxlsULK69fE+28TnWDkmr9H8haq+t9eCe7KMeXv
bBNVZOlDmOTINNRkCBbTQm5UshJXyt/9pqcfu3lPcm1R0Vpuq0VTabi/pb9N4XNV
M8mzdJlcDOxBFhrE0Ublj3TEacDoDo+H5bS3y19rvLd7AB574m0lbHcGdilv4zMQ
BJ46Dr8xE/4KNoZqeejcdf/h4lI783D34zbjl/01WBO9LvgEBgGJgwZxCYifQbSJ
1zvBsq9SeBLJrNLaJ3dpKcTkMDwGHqWRBHoX8EBuU+0nwZtHK0ySrnAm/dJpltjV
VErMAyPP4c1k7LUaPSo/rhCB4x8NwjJ4XqQG8JMHb7XZ7/9VwZR2IklrJq7pAcg3
kybIl8/M5LOYYqvrK4WDTFYR6ncDgMRzWan98vJLQUkR2d2lWtjNS5qIEc/7R7/k
iu1MqzT8X8D+EGZN4hWNPNJObgX+EJwdjpYX+kh06yU5LoPtzSKwtK8+aIn6nVKm
RbXcy51+WESdcw8ycsPe5kD/bqzYndOBbdEVJe/ROJCFG3Wyg+vVpVEC/Q7Zdp02
bEYDyrz+u073/K7SLwV9cdY/z3BXGtTOXHRRnzuCaHFPByWlD8DsDd7hIzYQ3McT
Z/UHJLF1GDbiZgZ3GA6YJG/8liAraIxLOQj6qE5XsMoPMk+Uu5OpJkL5hoXFS+ee
yW6CHg9780jttSDimm6aG5etZZcYy8EUrtDgcUfC3nZIlSr+NeB7TUSdxj31cHQn
odj/TV7kTuNdTfHVqtl4C/93sy6yoVPmhGOHckUKwwSIXtw5l0yVCxr0bW1sSw4E
K96vEzbejZqbrtgtuxozpDvQNpBTc5nHAY1WEHyerePG1OFvazyftXa5Wlup2Zqj
LP5Ka1hJeocDjVM9GTeqA6prQjoeWrZtHuFXgKtRUQnWYzIMuY5+ZXyYTy1loW9Z
ENLZkYBvgfbSGkY9jeDT9Kq3AedwY7dgKsRz/KTUUc8ZYfzsiRt9bzSc8RdDwiR/
Su8dJ1kIczjz8JplyN3Zkj5zFn1pX5BMG0vxUrvTxgx0lTSGyEUPo3JD3zmg3pqC
tfmT1wvltTObJrzH5aGzwcsYbRa6Ux6Lg1LT4mJqzPdhNw3TuvEqQgDmOo6owmQT
KgPaKwZV9UlEqQ9Ix8RYYIdpvjJUNnImKhJ0fbPggoEDdcNJeWXOZFt9kb+RVpTN
KkcaUwL6lYjL9JiZ/6WX2porfHW5Ww4dIVf5Cc8XW/JbL98w6fv/orzyX45TfzUF
MhANTXCByQTag8mDL6j/7Bi0JhCw2F9d20B/je87aczvziBjTj/WKais4gdVYq2s
kX5ZzqE0RRSQvnD4mS4uEBGKduq9+cjbCiL/iuWaIQcItd08HuW95R311UZ8Q0A4
0dXwCDfw0LqnBjt7BKm0uVp/2cdwfh6ktX1rofq6E9Mgt+O6LUoy5oEza6Tr/OX7
ym0CIf44ZvUxG+ii/6zK8vWSxx+woZMBLyC2xx7fJhG79P+c7g0KdgYe2/u1gLLL
HjEcNJadnxfDGYZuP4leDkZyNodlzgxTSz3i2tnJlRvTgvSYw9hh8C1Tvx+ajxij
OIcWHahwSoBL5VN3CMsXqUzZOLddc72gQU9dowadlx8zeSYwJHWKMTRxIgUtWPQX
x4bopocbt5ojaxkki6qozThKNNcyc1cAxorgMCy95pufkZ0nx+j+2QkiFBjwo+wr
0MYvrC18yjRgDE0nOkUdIP8EJRdoSBwFCJvWUtLAyeSyrsdU98tOl+CftsWgbaAe
4Hbww2mqQnOjwaKPBtUrqKQuCbezBM/5JDJYjZG/RVIwdlarElkkeUXKT/uxgJAK
iZsLw8xzRGwVk9RUoIhyYmQPC2C/QImVkWT3fiHJ2dyvNhRCPked14ik6mati9Lc
GdjoZp7ftXN5c9x8/KL3TXAy8y/JreghJfzwjx95QWqSopZr9QT35kZRne45oUXD
YCMg11QWDbNA0b2hAJ54A0ifqP+HGbUYl/wFnrUK1ErgSmz4kdXuL9+WEvj/vRnS
4NbZMy2lcexHr4We6cWWuo7v4mao8YRGStcrPCDwhQIjKOX852ek1FMhG8dslK4/
BRvTEiz6tC8Fy+m81aW8cbmZISg5wFc3KGncA42g4bvXMg0JMtXSKB0JppcWbE1J
Z1CraSNJZDqASpeILfsTBbT84v9hLT0u6kO+PgkqFIvBowk0IwyC0eZ6e/VeRuoA
kTuHfZjX4HYGwOMwL49oAOL0h06yGt0stvMkqUFDI91YxEY6vKad4I7yFa45Uw8t
NKJEfEXclWB/CrbKsVFAPQrLHke50Aowj6RQ/GmWbtO077ERgQI/5j2/bqsVSKny
5PzUcWqYA2vFYu3QpMWV9gzzeMTD9u6BztLj1j8OQqcKX1hD6A0COCVVjG9IEzlQ
NEdKM6PVglBd3PxrOXhk5SRodNM1ExSuGEAH/pOfRgcZOfZKbfY8XIo1Tn4zBFOJ
d1Yvm90Z337Q9f9T306Nt9YTFOq4H/qablZWnrJiVHqGHXz77ml8VUCzt+g5YrZp
g7WY3xlDtPyqWaq6Zu/Jn1LW74M31VopBCW1XbaHoTHmxBpat1AVQKkb6fKtqPJV
Oghbh+6o1vACCan3pvzJx63gExnvMTYkqrtrRe6vZKN+iBt6rGKiqhP+iOUMISQZ
nqcrf+FufLYV7hdp9XmiiS/CDdyOM+uFeBWnekY/qhk/P30BB2leSo9XH2SyEkNP
CW/sBks81UEUa6gaTHua/lRMB/KBzyk6+WgAiWuoQsA8FbVIrmj4VgckFMxpIwJV
TQOyGOIkiJJUKWyD77h6eezTZE1QdbHBJ6nJF/FQWkQXnnjJcY4bosPDNbGkwFL7
caGjObe1cy3+ZgyunWBZFakjJSJ+p+DPbhYqh7JbQqcliD3VS0Rcm6/XSntDpok7
m9uOIeGYgdT22xy4uqpqsFo91g3ScCCUEhBRraoSJcN3Ad39oIh8yX/5HLwh/ZxZ
0XacySR8sxxMOzGX02u4d9/kLE9LtfTgC39X1DunK9MqCFhJlIIPutujFQL2f9pN
7PKY7ns+JwVEebmRie5b43P2ccoGLiZu+QUBo8vV9/Bj7WoMBXhFJdV78kSsoGkv
l+77wS82+MirThh5UVMyVYF3BgxfKmbiZIMZYjzvR7i4ujVRDoFREIkc0IemB/bq
yC1OA5qNk6wigiIts+zxworehjwRoRoXEDpQ3zQ0QFBFmERL+ibrnbwtSmu9dRp3
XnAJiYN+iNeNoawxJrLEtLkA+Av3ysUiWc0bYXTwNig3JagSltVtP5tdODdUXp3Y
XluO3nuzpGzsQRCHyGBEcDv2W1Vehs7ePoZch37oavxEwYXBoj312yU9e02BQDr7
9AgXSDwGr4uVkyx2mzuRK+/82qnz2zMb6skjWR8HC0JavyRtSMhHGNkdz3a3Kii0
+jWlSFkdgkBUSprPHV1CjGa+RST0pjDro2Q/6MaUb9B3W3ztIw/82INKNOb0h3WM
5MHw+9rsbulKVzrlRKb9cDHVGglfJHPkLmbXo1PbpqVn2K3ExOdWzbP+DEKoa06l
RmWnmRRf1yd50n0SJ3gO9LbO0zqlx7xlbfAK1HYGweKX4Xb/MzxHMj2QeA2Vt55O
vUEOqed1Id8th3ruC8S+lJUPoAwDQ25DmeI/qWxYpobwRxPSac9Z6UlfHxRD/dQh
4XcfeDKklemSebfoOAbxrlJP//YXM3UFUiUffD/y5wbXaotJImuFEXayN2xqMl2w
CRsRhbRTHHKTGaepmvydq6rrzZXNGt5kx2gUqACVTigdMYY2EGYKyNBbk9OfFqrh
Gg8Ez09LxRXr2Dr5urbOxKASwnZyR7QFS/rHLFKSxNEGUrQIetyCs8Mi7uhEbiMT
uVCw5kS4zV+IU+wtxpMd/vV7fo9pmu+iqIKb6v3KsN4P8FD8OBbi7b/ZxQjwTNmb
lnSVANv8T4rjEZGOLszuEmX9WwyQO0Me4FxuuiBI4qlhouPNWyPncA0oTeUJFg1Y
cDxkF8heXH4NAveOBvgD+Q6jxNHrKFF8lUMDODYpQ5asNkAhjT9RbvxkkXFx/vcg
PBtqUbKxqN5aCs5r9hEJlHfCxcUouZlRYQxosgJP9vWkNriksZWX903skhWEAFQ6
aUzPa69AUiHScHaxfH5OaVI7iQd9C0n1pMGwA4BcwoTdeKt4U0o8UKU0f4gvAmHE
E6UhoJEPDXRFsNWU1v20R0dKNto9Wi3HYzkutIol34HUQFWyi/6ya3IJlktIxA/y
jS+Ty2ImMz/pMuVWU2dgETSe6ugaPPRogCyOpbfSdKqffmD3DbLrFz1wTB7K9Q13
UPNyAGTkFEQfM/i6R9W6se3e5Gsq62DhzFdcLiW9czrotaYz8suJp7gyZCXuP8st
edm4zPUDev7dt/btXqRmGC3JWP5+jc9bJwBF50uyMMKGgGsC7Lhcbop35eg280sc
NFbWushh8T2Hd1/Kj+XrWur70CtYb8OPlopUQrcnllAIC+YUzyG/1M+zU6nBtl/Z
oZj8CUZsVcLjabwe535umxC8bJouGBZJ81NF03QQ/FqCsK89Vx7HkbG8Ym3kWgvp
v+foyVJIHAxUc5EGsmOyExHlmxpm1IngOXGFRZebmbkLXVxMez9OSvhcQEYqj1/N
7uHwcPEdHjoOxS0K3L3iVMwfzC4JKd/2csktCXsqqwK3KMOmiOzKgWeWolCikCdV
DwETH4j8IuOF/qtluzgszxxc6+Tzk5R9qpqUgEZ+vCeqVyKs3zdj6PAvdJYarSJG
3W5L6hAYV6Xsj4v00ZE9cTc8IV38M+9iJwy41aYvDTsrP+eOIhp9Uksm4RWUToXI
jryNCzNzGrnue9bu5zHC0t6AT+RZJUF+JYHAeBgfvUs/ZmRSkf+ZLmsfSAf7yDSP
pbzU2V4Rm+XV4xNd6w0HOBemAe9PKciB+YlsCv7MLQviO1U+ecIgnRh0yGr4ENC5
kll+EbioR8MS/GxLuvtIw8uchNsAS99qxVSDm3kDOwPmac9ZfhTPsmJHshgBxpVh
f9LBrFjENB2/pZuGzKLvrdKdsrY6df1MSO2Ltkd4d20ANRtCsAUtRciTt6f7hzeZ
7hO1r4QXuo9NkMQyN4JrxuSGmPe9BqLysAx7CSaM48bqrpntEHbbRu6BykPQESux
SxziGFGvDqGvwfK2T435tgzBwaA5h5BGHjXeyBaE/QiXaOinWqslxdBgSdcluTAq
PlY704c7Qs+1F94AsBcxKxkUcbkVE4nus+GQtASpWVEmoc3lq+iPEdwfHzDs5o0W
+GWgYEpvlOB6hCl75RGuEvqUJTOlNKxQiJN4ayHuPi9eDaxdFmylmY8Zv99u8U0H
BE853kW45evzdGTizLNgkYd6J3bzZ0wIAoSl1a5I/tm4bAu4aZB7pq2I78nX5Et6
LmOe46v+IfSuLbXfXsxpUXIKYKd1zC6MYqw3Y4JdYQQ2zMCh490zwbNcg7Bw0fiH
pBR1Q/99MsMLs9sb7t8t37+KlkR1t8seeI8HT+a+g6y9FwlO5F4c57+jaVwUEsrL
NgRDq+McaGiq0mymwR0b5N0VqDivVEO2xh5wba4gXd5ftazNM0E52ccO+YvsfvQV
MvPVJ8NP+Dotc2mHWrZrlsScVuHX0jO6C2cfGOPsMbXptvYQorLvNwx6MhsA8MlT
5dlFoNySvDylNweMQlJTDyiH8qEDRsCwoUP6W/AK2Br20vyalClHSJyVbVdSVCGj
R8zkgpeZRNSJi3IkJk+ls6tx0RSG4kP7/JdKLwiLgstaIFd7FluG/kQDMnbQgYfx
IIK3kvJIrOYbu31O/XjSP1NkAji5hDCeQUinzoMffOOYT3cLEPPNAkTdBW/o8ZP7
wj1scw9er4TZLkIGfz9KRYmYvpfEWcv8hPjDCG1mxX6Co4CKNL2EyoyaC751v/Gn
058zuHIpr0uCZoHib0dQjFPrAJsfaaX38/dsKTACCzOD4sgaRsAUHRrwJFdXldRo
k37VSC+TYNRnhNY77gNEszI6++2wyv3t541taQQz6ba2QQFdnznmVXV5Lf0d7VMQ
NmUx/klZq0CCCCVWrISUcVsMaO1mENLtNC1RZiMBQo8dfnG09Xkl8JiwJPDtz1lp
BpMKYvfpxrWel/bgGolk3PFg1NNd7mGLCgwGYGT1P/dOwc3yQp2k9xb8L5EIaPUj
GR7da/pbj3QyI1YQCJn1rkM9FdyU1a6XPljz9VBTWMqndNf93IpU7kuSNc0SMV0g
Gq52/aTFe/xp13/Xt7QswcECHZbwKq6X8N6kt9GFPXvBU/Ig8am71WLGUiF7lzmy
3Iwzoz4/QZLqdS+qE4cxeLYiAIlmWAAO8npSOYaZJZVJeO594DlfL9gfRymkce7p
4jdZH+wtmDiwdQcKXFT/WQs/hIybbgbJ1Lw4luO13eUXNccosjQ8NyXCP6/Eg3XS
zdKqCJSi7aU//T21xvf23wiGcUFQRX5nSgtdMZu00eghOUN6eBguRf5zQ/AjJlqB
LuM/WyVligsfybUve8diT0891+XSX8WjJYPD6C+aPh0DGuF2+eXw8eWOgs6TDBO0
jejUy0saAGiolTCW48giVEWxZLZe1gdl1Mz6n7KC2aMG85a93KMt/SpHtjqYfRcE
2Yf3OQryX1HN2RYj9Q6ypgrGp++m3VMzDXDbsgZaghE7d7hu/5LzcXO1geVY/fWS
L0yvRYE0GmBXshqKOv4VmXdrt9+lI4SxlCmttCq5ZKNGyDfzcakBNISuK54aZdNm
PWEwX6/9fUblMHwtEDQrsKUUNzlEbI9yypYz+J6iXSdkSnWeeCdxz6mgVB1ouaS0
YA37E8cRm2qxs+C8qBnFOTpExOptsQtLCyklo3HGeXqJ6UEt+HRWedCC4pWPD2pE
sS/9RCbc29vvbslf3SMEyOOFqNmqChx/DVIP2v/fkXDsuu1M4XYNwtdEQmYVJ/Uq
B3UhrdF1UFxr9dSUhbbX4GJlOnKpvxBlKgEQ14jbSEbNdE6NlePqaSwvGYGV8zYm
H49TB2g+fYRfDVhKRWJihUXeE2aQ10Ha7xGi8dD3udQvezs4FCjGnx/rNSVr2Kma
0QLnb1VmJGhhvXSus/HX/U4KGACToxFDzVJ4Fp2FTZk7189bIdhaDSjMZEqtKbS2
dxGbYG0FH43dfwh6TuxuW8eGsB9fEFdd8f/EkxVs1vlQqiEA3WJV9EECJ2U3M9OU
JydEb0oO3NiPHuvRyCJUmK09cMZ8e9ZaOzFWrK0AoeI4/MOZm/AGnCJxgHN/dcXG
RxlBzKgLqIA4IM4j5864zm8T1LeavJFdQCriS1ZNgAFkCdMBhr6QpsF7GNO2m+EB
K/AfIV4NXmg0p9qx1sYTnR86dCEvCfJJWnWVWQzw4k5sOqOCOLX/gTxlDAI6WNYZ
TiPySxgHGm6C3S7O42tKzWCW8F8mJH12aW2TwiOP1pmctQHZ6nXIaUw+Z76mW1Z8
2VdPt54Q8+iSSeVvW8RG6VbAG1WmBAYz5NaLtp9QkdbAtwxKn4VbetHV/aNNgMxX
awSZR4YaH3hx2qmMqAhIcq7UPlr2/NqGo1oXoU0ZMEMdZWUIWJ9oFpKh2gcjHfLz
scURZQ6M4tRZXyLT/fgsp7hIPGOcU1nqc+zdFnyBls01m31UhG3URNJnJYNIFtcl
iFLlWKrysQAJpbeGJXoZY9/ZbHm4xVwGBUaeFv6LI3OiwHpTSVsl1d4tNw7LP6ud
fBvWcofff4/R7mq0PE6Uo6Bb95ex0qpiD2pJj4evQe/TaU4YdKjhaPt7NMjGls2S
Pkhw5liTuT2Vmqg2WMkq5SUc1bc5Tlt7rRCRZ4ffWApvJQysXKsHnp0Yy8OI1Khs
iUaic0ukI58WsPoJXD4LvXHq/ySC/75fGQWgczThSqRyj1SbdppCiQ0N7fdSkTMJ
6t9OHhkumde0N85d/vItxOvI9t8HX+OauRq2UQTLgOpS3dD1/0S3SaIIm7JhwkXt
9IAiP7cnmAZvrIXCU9yqKJ3hVJRSEay9UFT8S1TFEU5Tt7gqOFaYaPldSuzkw9Vf
Ik2cLh1y6bApLfMPVufWQzKRTY1sKgANmr6ScQSi64SWKRg2Tqd/WR/a128Wk8Sc
SYsQpt21MngfS7Eahrl0sDbmqKidORRDS6XLSjx5e7uD8G1ie8YMLxoGaPZC7kNd
SpgsSEEZWcpmwLILOz3tHCQGqQYlRwGeGBzIEfmaIgwwKkpYxidAdLRoAdDVMrnc
bpPBxUx4CP4z9EnMIC818YLt/t/P4FVYjqnwixGtpIuJy55R4N3qPM/UhHr2Cdpj
4wH4H+4kx+AReuKSc1qhL9l3sWypFFjkxtAZVssiU6d4RMEXVGt2DJj0KnQd9SBm
9T4n+a7N6Vn2hu88C7HR0N14+BEi6HQFKLEtFIkAbM33J3YbVRrH3or07PPAKcdW
/1HqW7c3gYkkHyh1xFfkXoTcNEch3yxyYNfvMd4ut/fmpzI/BUwgc0qIqtoI3Tqs
yW6zqna1Q9zVQgxCsxKCFn3V4Fk895QeGrV3KAzTawO2S4kNFruWxa7d/njBCy0X
ryNR+v21aSOJWd9plPjZu0qhprbIrafiQeQH241zWrBXi1kWBMl0gvu6dDXDjasv
c78jLf8T5Knyyg9GtNmFpXhqEP4TEIx/OjF7RlDZ2conshjFLgvY8ZCe+t5PS2bP
h1nvqe3jssQfZqXc1qnZbVp0OXRQaHdkXCdA72muCdSd8L0AUQDOXnmrVoFJPmkC
+NsjS2OxwTizN99x4wMNcLYuz8ROEu3eVRNp9A2/KC0WHK6dpEQNONg04loNYUxf
eeKEi0hkRyDJ25v9D3h9gHi9TYOV9l5BWnHWmMM28uTd2/+Gzi7wFGe8CL+NLwOk
b+FuO6JmMAa+5lsK7NyqapGQM8Acv9iUPiZu0fs63D/zBseuA3rZGDSShIBnAxZJ
wakzmANfH31EYVSCgKjBwnJ1UrpMZO+VuvrGyKQDi77JXhx/3Rc9J0f9c53M8j1O
2suTVe5uwRo55P4LNs3qJ8zuQKRs+vJpxzSc1tYKnOB5qkbkrr+pT6GPo2j+FOBI
bMuQvFKEI6eVHaP9m8LbLqIDwTND1uyDknMfQBS2NNPOXjLYiqC9AZtaoGWi4u00
FdAUSP2HrmGdd7qST9Y+5XtcYzFcIeQYHo75XhSTHOX7I+sXbrB4WzoEU1Hz56af
3zRKDDbVsxqpuvpfbYwBH6pD6yQrPCSMws3N53N2bekJAXdyM6ZQ4CmeYsvNUwUX
BE5lOZMTmJAO4okYfd3Tx63mm6tDuvKVQahopHR9Eik8RBjQ3AkjOrzFOawAKrrk
8NkdobIeIpktIhvpje5kQ97ZayLdHyxHBCyqBhKim6I+tuNPqu+4YQGaszdiOFm4
qMc44fGml33xAYmTMtPrTTc5IwT26kdB6pZALSZGW9mexcqjFuEeKsbiV5JAjv9x
etnGGR8bMLRkesIrxsQq84YWgMrS6sw4gVi2JvSD+GDAh/eR97wOq9tQNWLfw641
sM7aKhrgWUdChcanzY8slsw3DiLvNpwD1Vl3/tgmhSXVjQLXmKioe6xGxUiqRWJQ
7HC1vENcFFqBIvQxSB0xtV3LjO+TyH4lrUM1fXtB1RJ3d94wbj+plOphGI5UbDmL
HOQE6m6Q62FCT/ltZkPHsBMX1AIHSbGqhdSdtGBzfXUtoRJVmeQRUAUxBHcYbBxz
Mo9z6YYRFU3t7ajz7Oj/NBud4tiKo8cF7cbXxiGArTdcv3ybme6LLE3Ak3j5Jr2V
s8nEueUaFtF1vyyF75j7d/U8nU4WtdI8yV9Kl+2z31fuiQEKrcH02q/oAcR0tc4N
ST8kDReEhA+Mitll/SGzKtdXSI9TU651TTD7ep5PQl6xFEo5IzcDDor+UXeI7VnC
ELZvJRThXeBY2DXsx47NS38pitMt4fGHjL2TH95K7Wdk683ZAhVZ2wdAPNZ9KqwR
U7zzehOEVH7ozIijFK6bv9yCYcDWIbDqF7ci959+kKEMjZp3TZmYKPZvW2j64TdR
PInp0Vwx3UQSZeqydvVOeFGZJ+vWYkwUfq5L5fkOrBpztnn8sGxp+6pv+eBK7ulw
/YSFut48TvwXUll27JWj8390HyXqt8zZhr02TATmGG1yCrLY/dyIY4ezIK5wRoiK
ADPWKymaHtaRmlZqcPYrerHAf0NqCERoUqCYIhkYrxUb99hHQifndaqLZlfDaPVS
uA6oadpg12iheemMAf0JYnQfpkknWbzJxPwhj/5MUfjRpvcI5qI3yMU5nZlAX+CI
z7Abcjz53GCqV6NSEykYLKDzVU5K/PzWwIy8R4TZns1pldPeNfkH03lW5dEPVNur
gFMVmSp+MBcWF+FbIcFQp3juMiSwkoiWndcQhpzsRI8m+o18bEvGegsBsnmsgEBc
ux4Fa1FKitYEHRclugoT5g+oXGtkRfdA//T7h70OTwxTEsTaXgsUF2ua3sKKZ8CK
82zLMD5Rc9+8KeAIZmbRwI+Ox9cBXcFBdMGHqtsMjPh2lfIL4m+jvbQF0cZ/Ybf4
b4StDZgyWU/bdhQ6LAzBnE9808ZrxqlsrdHE3RgAHnCKvWg+9yMFOe8UPiOqkhr0
QXb6U6/bWIPOHirwIsRy22LWNVst30QygaJLiNMkIFoIwXIbjery1qDTDSzQuJ71
2cLq6qzcuGhr1XB/OjJTaSI/OCLGScZGMVUwDH/ABBQxWgW5pJx9lUSnomUEj+Dc
X8oUqAoa7YyTers/Aad5e8bJdACAcutzxIqIaG6EweArTKQ/PwSydn4EQYIB4nwQ
P0Vaq9MSYgxoGkC/fzyAmXoJ0gS2F5E39E8SexsqUwh6kHwOT84F/D4UVf2e7QTn
DNAKTw55BiENoIe+fL71uQpz4EDOwGnRNnnqwSiVDy0jPwgTJgVPPaWIgo4zSskV
hFlxyIFaDd+x7KDbrAzFZ3a6pDjy1j9ivGlyoes4DoBEyQn5R4114TKITEpTCA6i
aG7CnuRXLpphD9eXW0gNQCqQLeYcSdGLt4qtnaJKnKWUaFYFoVbaFdt06jDGZ4ZA
SWJRLxTNsB5Fb/a5V3nrB3X6aoFT4v9hU/vf/fDDM1/Wmik2NqQjshOpJohVsBY+
tUI8jXmZKFENbVnoZFSL7qLPsC6lua25NQJzW4fWdavOpCu8eMnrxgfhZ63Wup9v
1/FRf3jLDktPOaSewsImZW9uhOmgoRmF+GT6wLY4mgid56Xcq7eFLY5cKEEafl0+
bQWuu8+kqMHZ+rSe7wrTroppNFORe8LSi9Emw8YrFRLsEmegL/MUdLUM+ZpOsmu9
gDwZEbj9udcjiwZHk4yPxfbwMLVjnfwUhzW+bukIv3y+Kb9xVXWhcXfbAvDab6HI
G+xa0II1gO2QUFKIk0P1zGeNnLrhIF44IRQk4X5hX9ZBcZNP9BDnYsJHYL0gtcOM
q07GdqfZenyXKX0ngmuHMnbVplRPVnUxpDiyK6bljrP4Ua2fdYj+jPbFNnicYcxy
RbeGtSH7Wend2xSW2m6by4InvSu2FArFP8ySACrXewQIzJNNkmjR2VNb8byd88bB
iG0A7E5Lt/db56KqF3DI7R1PlbQmXjjrzDYDeukqjy6WZChnxBJHUlXUCIxb+sx7
mZaM9ChBuq+zRAy1PUTIYIoNAN0lBjoqE/v2kdkheMJprIx34o4Wcg89tkiclawi
swNuOLp9EVjMOKjxYW0BgQ0alvLiap3vzZYGaKy2ACyNhxBn9cDxJtmC1hgMEO8m
st4mA34HiXZmRnJ9B0sSIxVFwnYOpcpoenvxc4A4wL/8Fd//3KIC8KrnOFu7xsfd
A7uLsLiFX5IXwSgDKmq/k+nfF6q//leZp7El734xOzxRbUCgdrebfHZpIreyXXhu
dhTLuKA9W8MAmMgrZLCCP6y4YnFQveDntinlpkzOAcCmtmRfqKrQQC2oO1BWXW/y
3tVpJYQBMyhQNU2Acr4HArC728qjOLrnX8/pLqW4ebh/hrr+LWo31G8KFd2m04Od
4CIqZuhKYTCTxGuXvGBseXvu/oKY7ZhhVtqi69Z2e5+8beQ+RuANyyuUYBPR3B58
Llr6fugZyHJmc9g/mx35gVcamWiveWKNqi8dt3ks5NfjGy2yqvOYKLY2wCNzu28b
KEh2utpG4SUWatxvtB8Y9YAVA4J//PkpuEO9Dj09lcESZ4APhaAc4CxUP3cXX89f
JqIGooW4oUUjt505i2zqlOdosy3GshTZ/PgK0LW4ZZ6iSi67pNhW91fO/KtDjFLE
LSX2S5Hwn4MsUTfa+ig0VcnXLkSc+ELb4+s1g3V/TI9lI21nUqwhrYLU9BSC+rut
HDp1knD9sUHj5PP65LqUHT2ppEzkCjIpvQhBRm0sktO51ogl4xzkBwkrdv80M9Kw
Z3oNa4KFchbvcldg9P+GvSdECFsNz7bhJz//UEH8FRLjMZG0EVf3wTcy27a3YNqP
Ni9KLbdZnmhqq/gl1oj+5bE3cLTLpzKhAcD6w2Fr5IUMK7JMkJ3ILIRVrDC55Btq
LOJlSxyhaTgy46/1oS0SB0FJ5qPtHpRuuDR5WfS3lLAUV6h13k5BI1D0CC0ldlFm
aqzIvkkeP8r8EkStxU6Y4fMfL9j+J+nevuVWOjAcOQkfEiw7Q296hJNrYI4vzJax
75IWZUJmLcA9peWo7ENMMoOiV7U+C1F2lJcTzR6RT18iBN3bInwgjoM/Trr6Yq0X
oGJAfDn7gQ71dwS+Fu11+UK2xACbLpkuH2maC0sMFBhimOeiXjqFJ3wYZV4Y8lL7
HSHKXTw3QFhG+qdPNjWvRdMNLfsAjK4eiqBH/r739MLzqhGkdwfx9RHqLryGEBA9
4lGFQIRK125yHwBtJkDy7dVlOp7JDuZVz0AezYnPux8kmPkRlSgevFlwfdfWd7f/
nUFXMkWdlNw6ziGYb7g3yl23eI3qMzWZBzRxbNzzyDpzk3RpdnSkPlbNvfs109wc
8AzZu499SWC5p09NHhULYiHHHQD0D1KZfO9eVEvJJFnHmT/jZ6gLh9/oR6s3cbEZ
fEcX4VQA50ZdeVx9jZIyI8QfiZuk3GB59Uta7bWvBReIZ/YkfUNEiRRM3vy0rMUg
gALD+wxpKMTaKl2R9tXiCuce44BEvnr2ILoOKyiUHNcbolj/IzweejFWdac2gPGs
/1VCrxJOMsU0jGZ+sHkazNg/NJq8Ap7DhC7NUk0DWomAhRnFWzsGvV0heRMvIO9h
dEOG1pgmjKrC0Q+CBVrPFfnsh8JoP51mJLcdeAyM0l8L5j6iy23/A9I9oEx0lJ48
tzvChTtw0WVBjgyjjQHLkGsVIJ0J/B0IyPPkJKo0YBXp0uxGH3GS3YyLrTyrjdUT
A9HqAiUE+DFPkf1PL+i6lojeCpCoDpDu6upsIejmrrhB3aPjjY1vrpDf9jD7IDkR
TTB16Ns48ZpqZt6gmJS/QH37+nBhlKC3b684s3DJN7radylJXrkSZbJ+xbmvoMrb
lBz/s4dzYl/kEoTGOdMIGQEbGc9ny+p/qtUyvsRCkg44v1+tqV+e/QU18euf+71u
7xWUYwHLEFPzvXfWg4JNLfhRUIWDwUaG2YqXQvo65e+FzyiJY7V9dKWKXK0Yfv0p
s+EE7Yy6lkE/EzquVJ39zI0CSYsY5ThyPp0Mg+CPwEn4R7vZ4Zak4aROKssOzVUM
L3vrXo/gCcBRUOTsNE0Qy422Akr+S631T1UQovc6aF7HXDHbuSDc4AP32F84MweY
7aoIKlev7vYgEJfEltKqpoeCmsQ4hdUgvt3NlB6uMBoDK2wCI6iXVffEXrnaY3FL
nGcU8e5HeVh8xeUWkwVwrdXKdrvXxBPSQRNfq0nl+RI6zwtPMPtF2jdKR1ggNajW
AD3Gi8KtTvj9eJeCTkPpeoVrVynHyDD2hj3c9ERwWB0sndA8IXLuFII63iUVnqmm
t3QBjoQnEOB45wN+pKmHYXABow3o7fYU6kIct2bWUmwgdSE9h8iJ+YQQH5xPQcfK
bUNgd86aDOMTWobQRqYyL3XTkiz4BXnHka7axe5uaUa6IIO3bn9utPJPpBCVN4Vi
ezGAG5dXXV5QV8V6H6bYd5iK9JnCMsm36UHWUTNPAon788hjrPq+P7+ITgIYXz1d
lCCHgDKJV+dvfzS+qaSx88yJm9WRk0pTCbi67d9PwEpCic5CFEb0Wfpxey+Eqcoz
emfHRs5AotRCvhKvpIaYAlcPAjgiP+qg7n5Zff+CldJ0suTBJdSJBop+DtECQ3QX
hYwwwzmy2/eAsSmineWdu6ngy5tjBygqaqZ6szxfb1aC1dW+x3YGLZBEJXqph81Q
ovxQmzixuwOvqbASr3SU2blCEgryANORNqod5nyusPNUCUyhXn9AEsizAYOC3e27
ujdYNiJwdgkpmfdswQBzls1QktF+MiSr+Dyc1T6Ru/DD9jgeAPk3qn39BTBJuu2h
HfcPuZcdmtgodP+6XgRYgrLmXqsDg2pZP34866ELTM8oywEGJZn39BFjBbjw7dVM
/Rha+igGqP23l7DvZtFCRqHaoUUGv0NCY7CNb+CDhEa93xEZu+Hhh1MhlwFz0nvr
P60QHbxZLflECHYIGxnFL1AaSVXl3rqjY0sGAQ2UrtwLZa+MMZ/ivrDXdtdTGFtY
9ig0DLxDzq6e73i5QfB6ZTvMpdZHofzZmwg/tmZsEqc13OwnwKJLkVowMjvPmxVu
RLcftF/PWuNtfvQ9bX6KKzxwAZM4HImbRz4wGY581zvw7enH6w1kYL6wwVEU1T4W
DkLgjpWOXV2vAdacK6vvtPq6gFDLeEbz3LGcrDZVeKP4VCNQtpet2YyWBId7lSY/
sbWa/TAMLtKLzyEiJi9aWoGxfiwL3TAOblcqRqKxv31QyDZHD+o0ECXYSFP+29Un
JCXoBvwWXQPFK5T4Dcz1fpoj3vNZFVJDl2nqpV2IlcUPKZV4OoIcVrLwzKnlZQ3h
U+MB14ETkdaLh/q1dJyV0mmWcopoFy5JavjpuAu31Vn+CD0+uEvrwWEVDaHEeG7v
l94iapzkNqlACmDxuDno9oSfemTdqxHV58KKCLg39ES2hW47MP0GLuAk84od6mzq
QUnp0dvHw0Pi8Ysxr87t6Xxmp0SQ0dRYuWVaK8sPwZiYREcNZU1Pg9pyqU1xBHEI
/dhMyuiOc8NDA+AaiJV7UllRlfNXMaz3YKlFDGt1nPr4nIIEkgN5mpSKdFsnL2Bu
l4z9hijbbZ/sngl1lj1LMe+mh9Rr25JePL8TLAn/Walr9vre46h7RGumLRCWgBY5
jikOj59VH1Ra74Uxgw76rp13BChvgN6LlHOxk8RqkoKXUykhRRLJQWD7Sv/vcu+9
4Hfu3UwQ6hPRF51H2ay3be0nm+a8fIh1l77FZlByBLZ1lPk1UPg2SUjgrGJCmo6F
elx0kYfcmRknFyaxA9ahsFZGsk1UtipcqhuRVf0BX921xwItp8u3uXx7z69LktcW
7hQqZ0Ffdf1tevY6HVOP5CBR8umX15HQCN1G1LyLhLKxi+532oLpd0UlAXAZP/nf
sZb9NbIT8Nxt99nLxgQlMNKhPoIhh3WYEog5RRncbHVvpu7B5lFmX2ElG0xulH+P
XY+woOm6NM0MCSrnQ82Pi1qOdc+qrUmHFnSU7aDZuxxBUusnIAbgZs9/iAbY1Um4
9U19eGTyUUlefp8p96WPCoP+y9svMXMC1CqxI0XehF0l02VRWLD5i7wV4uIvtM+j
O+0Cgi/5J8NJtny0mmhXnKX3T7cUQrStIBStPkCDeiKu9RdB30au6bjQiqL8IY4I
ddSuYqhf+toem4Bm0s2AnWNssBAUrbqx8EO9vKFLmXhdZ0A2YWOu/HMVD3i7gWAv
mx09p1wTYX5cjl5NynarRS2NrrD13JzRsi0q29SWed7TD9yh8hPITZr6IYUExxd9
Fkcpxsce/q4zfncwJYBo4CWdbACCHp8csrNoZqJ/XLbBFVHA/MxQz7DRtj2DRP6O
reNjT6mSA/VuqvkOFE9AioVamQU7QjPe3POOwcOEntb12VI+kxFuM/85XbD+oUBh
xGgyIHp+iHdjqC3PiNtCdetnim3BuU5VUhPJCsmy+GNBg1NZdzNArJY2rOxF+rsL
Lzl6WY/EPG/s3RN3S1/1OQSDQtMxJehIADI/INjU+F36REZKOpPeXKbP2y1nnpde
wm9ZGvZ+RgFo2gDNQUfyxdIyjcgPVOyvkKyUt5QZDq+1Pj/FCj5+kw1hz96957rV
OkJhc9CIjKb2J1XaFCh2G+VE2yKv9Wn8CM3SjqVIevrnJVySceVkA+gj0ctSzblh
k0ju9o86sxum/s0pgxB+quXwHfQyxNxOtrbU/Y6nlayYyWSis8mUKuT0fjAqHYT3
yaowOtucBwOyESvv4UagZCrtnSTklo06vhKzXX2ysQY2og6N6JTMRCDgpm3bG9cl
vzUJ/nPcODh68SNarRs5cG71iFbl+e9QafBE97EwfStF0YBMLKua3XI8cG5EW2im
2NHBgORS+8hlIO1IKjDnHt7q0D6r7zMvEUYRUV2RN/XbP/YJcRu9s/OByA6cxfIo
LoXYDm42rQZ3YA+UScxkoQtFeU/eMg9VeJJ1KdNTaGFOJ9q8KNV86bOfz5a8JysM
KxvqYy2w1E+qJRxyf+7J1Z7p9+P8iOAz91huFVJO1KFuQSw2GdNrh7aTldZ5cG6Q
9Y2u94f0KqvjltI00zcBDzTNN0SZeiFsXq0VDVkuoimlRL9cMn80rmmqc3n4Wh7/
oZK4xdIq1IBGXo7jcEt6siHUp752lNcyp26u14F0r4Z/x8SAAerkC2MjZWulBB4T
yysldkJfc9/2egLWHtOBfVeLD0vtbLGOgC9bsjOJmFBZRQC2rgpoVQPIkWkH1s3+
/nHrs0S9QFX7rntYlWkZM/pcbcql5+wXcIaYki4DnaMb9sw0z6yxwXmRJ+x3CY0P
RxoTurqNbzXMrlCwljhzsNfd6ZIvbhQQWSnNNAqQWLqHBjUr7I6lFnIfI7sdNPhz
ZdqQ7aLcCpBCSUp2+rm+oq84a1WqRPxbCjVfru6vkMg8E/tHNLiDwIOiYhviYr/s
FkAoyPB1Nqt7sWGr0AqVJ7BTXA3oKi/JhHvrYXaTsJaN5ojAjIHVRRbz0EtOV506
mOzS1XcxWPXPUBAqVpF1Qu3xTKTBYDNq4J7ikSS7QhXW75qAoraaC5BCUjsWTJ6P
o/I7lYnmu9JYM8Fw4ybrBPWOEbqUS06joOPIJDuWYvwITAl/rM/s81qqvQcwowke
29XDxOTyZ+Ys/DweAXFTcZrLRcnlVj7BaAimpDr8y2N5uFVW5cmqOALe1vA4Qd3R
F3bhP7bRzMKzj59/rXVLA0PaAH+6305MmuYJlgb5AaA0RyOQc/83b2whHKNlE/ch
mqcIotJWHcklRuYcGl9zY4jPDAbikDjGpI4N04MZkCu13Igrm7IVvSTVj0Pq6TdI
vdGk855zHyqZaD+iDx5S3l1BvhkiEAkHr73x/eq5hvAD0zfoN+8KR+ptjz/L4xng
h+yMBo/pxGmM1d9oOTGZ2g9emzFBdleiqgr1nTGx1qFpA38XaZe5cKUiCN+AnYDc
jGjGmwFUPDlHPlm7fDvE4ykWo6RNmZP30pG+xqEzSb0WVYVV5hV1E7ljU2dsyM+Y
G3/v4To75dIZxPp9PmxNLSnISyxZqxlEFU8P7uXmO2hmPh2WYuPZC5fl669tyAUf
DUCwZzeM0h5EyWYrio8D8ycYHmS5u4Ludq/+cA2+IT6viiSMW2kMfNuRnPCkaKiL
EdleZzLAilxx5m9mhuh5y8gobBUTPW0/xxuOwCa1wsb2REgp85fyQiCqPDLlDsY0
ZqcpI4ltoq4NdWRqpTe3/3j3CSuUcwXryaov64k1U/w5UUIYdfNb7ca6orKt46i1
MfUdShpga4J5TB3EJzPYlTIsSXTttH1y1VA5s7nwvBi+12zSb0utK3csik/NU+Hf
dKrPAV/xNIY+izWR5t/Z8FTJl3zLHy6gFxqwmRK9cqOaFFyufeMShE5eT4Qk4Q+n
gPsldSx3rfBFUM1zuE6r4BJmQS2fcTvaR6oVXJzEB3l/eMEc2Esq23/WsR3M9jVd
nStBleJLIIweS/xCxB7oDflVTgGHUDtkitwJUuPcBheaoIl2akO29yXksH2U59an
L/WsSRETswFhTb0Mm9b57rnFO7Vp+j2l3kipSZA9FLoexEQiC9cfDYB7iBZsSnrU
60cQNkGHI5cUDrmpyfqzTzTB89cBNI6UuCZimtxvSyhXijoamwMAhn9UYbz/wbzu
0Le1Qj8floF8yIccqZsfH0wybpw9035RYYFo2akHtAenQVSJsFye5M5v+vje9CpO
93+QijMx49LOCv+JTL+ksfxGdRoV610oPe3sU7OZXzRAp7+tYidZyvo1+R9dyHl/
cxEq68Avepd+O2ASe7n/mul1CtkENpvL4euYLlxGZaYSEfcdxtONx3f+8W6fk4CE
Kj/+s5j1iIyEA8x1WT7447lGDd1k+rDgWefhFp/lQY07uGOYGmK/ix8ZLCjdY2oV
z9I3o24vbdTcf+u/hZXKX6sSaminjTHZwUGGEE+neCx9nuOJgRBONRYgOgHl6fEi
L+15qhg+m5DCZBcRr8Y4bGN5b/j7aRsKVQoZ2K7y5rR3YEtkKT4KXnv76mftyIGt
FMYoPiSaPJkZ4nABt4lpc8uDGPoQnbfiz8lCEF7WHzYlyOF9UQudMxwfAtGxZb1G
+4mZrILXf8czmTETIoskvSfPG2QmQgaoxv54JFWhqMfe+zHPQ3IMrFP3q4sSn6F6
r91z28OJiirSI0Y86YnfUrBuHyNGiejurtqNxx0cS/MoeaSIT3rf7OHrIL+6JpJf
vhbCgXit++uUL0FjWNYJtVMFw8JxJQe4xQYzA4IdTf/k+2hqymOg7jql+7dwpCHb
KsfqD4LFlleDbC+TS/rQG/RIqpPK8v2uZ2xRnhJ4Qe6vqEBkF0hX6jPgJVDJY++b
rWBDjeJ20yI+RgyiDH4CgDEA/t/7DpeUArR8p1lY4fy34zY9y3RzQRdznHevSSQL
Xf8z+TRA1iSyLZOilgOAn8W5AgoQXUK/1YzYolbmvqI5AUs+tlmhA54R3X5Ow5xz
6GxbqW6O/QiPswTSL1qd0ryWNOGRkR6pOm5RwTurSOnRTNyUinubW02V37TVdapb
i8y17vwCMsE22jwrDqdXF2YW9Ag9zqpjLrNnzdc27AcoSxcvS9BzlsyWtjKCKrIr
78aOP3rbVD3pbAkSqZDvuxIioJP6roIaUh5dfZ0rrFGyuNuDD9ulgKxD+OBSuw8n
0H7hdNkArhm2A6hXFV90if55gyZ6GpQ3VlXxg7/L+ItXmgXaTdWbWRjq/XQC+MA8
3PU98/X2xWY0VIgP48w6K9sA5XNxGLmtWsrN3O8CAiPGz7dbkMPhGbh0Kbqj4975
2OZCsEAXbfd0JPjnTTP4MJ0xaZArPotfkh72IODt4NzSHLZ6BRItBEdszYQoftiJ
BKQBU13pvtQJ+i5YeyWrVV5lGGe0Im+POv7cTT0W3mHBK6aCHOmmtYPHa/+DM00Z
eIJT0Mm36GMr3UbGrE9WQuycXRlbJVuRhPDRMK9Pf5nTN44pMLGWCPmXf0ZLDCgb
gwJCbY6QY5HnacA4oiKvLxr/OYLxjv+uO4LLlnBHT/NdqiyDWC95NVCIuRkAJ9qp
/fuN4syvauZVSsj+wwvVCFlyEFcEwnFIiDz59onohQGE0DvGRDQvp2uAJToewFuj
MfA6d7vnv7Hsf4pClTDZN9b656b/1ZWnkg6lbPhCOMX93tZ8Nus1ys6wNcRqe4gm
+VICbLx9EwZdwiYU6vJIZVtdbf4c4Nki/4pFQpeBPMKqqJW6nNaBS/MCZbkkW5BE
e3bjD9IFJGMy9lv8bVqmcnadTOFpIDy20VbkJK4uo8iiklLVqoqNFC3J1gv8gGRQ
PCe5svOJYOUAaDumHULUG7vZYeSF0v9eoGtVxqF0QdSyp/e2W7SYF3SNX1tmiyBD
kh9gQt46BO02BXgHv6ppYQKvkGGR2VUkgepWcIvxL6YndBaB8n1n9m41q/r2EEzO
zZ/s3jbKOse2TaOOn5hWseBKbkTrupqYmQKlL9oZh0OyVcJpLMnzOl6Siau81g79
u7/UDoAnwBVckBtPBrw6JydmgSao1TRhndru/3C2U/wgMYFHB8guw5gaesf1ztIB
I+r+p0/tqrQnHRMceOrZ8rOE85cQRsZ6JUbpDWUL3GtYqtYPpUZXvKphCkaflKzx
0t8dfxntOsjCbY1rUFeWat3ir1+hE2p4uaGZFOLF6yzjDJi+Hq9SApDAjSuhrhVA
YjFhyLwHdAOES6VE6yWOgqHbsUq7CX4ndRQSnjefOs5azCFRJgjgDwbRCGiZY5Xz
pmD9+P7lzs+jl1v4f4GsdYWNUfkQ17BNiKB7VYlRCA+MXtNoVxB+PY5UGyno/PHx
vu8ZmjU4LAYWFttdQ4br246L5lL3N+88Fks/UEp43cpgsg8GiTUbYrBS1ueQi192
oUVodIoA8QDqiWLvIP6t18wnMuGXILBIKrKwG0gHj/WfZ39wbKYa0zRW9NzD4QKA
BRO9WQEm3jaiG5Q4Gyaw0JdDbbw99iP1NU9IDQUtE1rhgvi8zAHxOcPt9W3f4kIb
3LlEjTiYyahWPKMm10err+LHWK7qZkFRsFiZBeSlwZcp8LFa5qO0jpTIdQhFm+ni
udv0yfFJ4hTnaEdyr5xiGs+3b5uVepOf8LgRcZ3Fqm8FYsF65Bq/BeUABwLUplDw
zTB3SBLsCFpnUqY4ovJrj2iwBLT7zxoGvxjUGEkpDQ2rhZMgN1UPi8e2YHuMvzyu
RNB6uqxDdwTL79RJ+k57LjiWSa8fW3qx3nho9IY1gVuTJ+MfpLZfmyyPFN2DsLpP
otT6p4EacuU9t48l04QfMnSuJm6JJFmOwAHB2t3jQC/OeyvStsc9UMAHkEowGLCS
RCy4hr1SdUl3hR3Di3f7xsu2kuAOssqFyit49DQcXhkhUn6xYoJBiSw/dkP/qKQj
FI4tjSPkFHxPnCHRcZ8lrWqssUge5/j1W9zQp1iLqtvimJplp26zji5pGPj9hWK4
h/HSjRVSC64hb0Jte4ghLxU++fBRBus++m6O78zEeZvkAn0yQYQxAQ2J94DLmaa7
rdNzWh6rpc4oVioaThZZZaponw8M4CS3rrIw86HPsYkyqqJ8Cz1TNH66pGhvhzbv
UctOqy/pSw9fiUs9bsnRIpMvjPXRWYwwmN2eONJ0+PO81Ck0VIokIJOyK1qoOeGn
aSRARoDakz/Vhmhjv+u7zXldiRvZ0Lg6UkkwRO98NPGzQH8KZUkDYVIVRMYzqmpf
hdjZklASFmjoRFX6ao59D4+YXlMs2vP95ZdwUwOgoaay1lmTnXW0mAQlHkuAJuW0
UHbdHudisbUIGistidYWqlrPkRPWBtBY7hvP6k3WPERrGJ0h8PS0RcWABmnMEXoN
vpK6GLefk7RsyfNsZeHrBShK7LdO/DkMgKzpSnuQzwEw0DQeNEbW3b4Hax6i/nKp
O60nSnj8rv5Z707rnhl20Cu4wB7JCJvZS42iUbP6+xj0xtAJWEOf6mcxO7vKxehL
jEnNBQ4SJ459bP6IvulJ+sxTjK0TX7C+O+hSwvnUieVIF5PRmjZq7c42bu8GM9Pc
f7BnHvbOjI991NAANkzPBnCM/khPAofUOykw3GwyfL4+fuvha4vyu0Ph149PaNkD
J4Ahw4OuiCATVIFImt6ftroxxdja02gFsr+hZPW6CSNVHIgx0AxOB16NjuJPe97j
aJEXF0XX69XWrp0Yl779TPaPJlGEOhB8WxcI3fWomKB6JUrZmIOXqpSQJIuXWoxc
l0RXRW7+woyViwkjvI/CprUiL+dxWXYNwxErv02NAxVHcJz49lJlM3OPdo2F12Jc
m96+6x2eqQYSIGj5w1QiQfsIsqZQTupMM14pOhrS3kOs2Rh//CKlpLS29YxeMIoF
GefuUOtelz0KUhIBuFvqouuZjuueVZz60izUZ6EKjC3+w4terIvrP/9ziiaR3T1N
UOOgfPeyzlUnForD3/76Asj69Z6bCKCMttCCdb1yYmHMgrm4riLMkZ1FcyXStwC7
7kSpLo+AzwcgdpxJBbl/fZ0568xIm3lHlf/2PWsgHJJTAJosQAo5IP7WGpimzsHv
zlO/leh85QTkL3cpOAgqZfojVnXfipdx6SOsyXkfaZyRaIiUm7rONqBgXcNiE2GZ
nyfrK7UwQvuTEQt7oWhmowi2j+GFbBA8Ucn4v4yiUCNBDJ+cGat6GvRcX86ma+sK
GsrDW8XoW4nFXdksx5bTZLHDVIiqm+qeav7SnHWcAX21/NbyqA/5kbSy8PAO7fBE
DDqOEscXNYn0VCKgPjjCeefcM3ZcC6spC0U9+Y4hVo0KAyZYnXWuRykmBmGxVNtq
L+XZteUEn37wD9h+MTazoDVg3QO12mj3lpc/ARawvB4JIQvC0GFvhzXAYy12I11Z
brAAHelB/YLNifqmPRmZBJBmKhMpdPaHPIyRLY8ndMFidhPoRQoBq3e5xiA1JNgN
uQQfC4h2y2TGeyamepJmszVuKD/I/Rd21VbpwoyyJVBtHfO8CUR1zuvneIcCM8nF
uylt4DUVovjFhOiphsz5LMtPKVu6bWPRCiQuFmFqQ06D1x5nmZ4Mr2IEW8LRXF9T
OarxiCzO8o5C3FXvh41Pp9dgXhLxAT1cN5Wi9+8wXbNf7U9YXFmGB+68HHl2X5s2
8lPOGhGKR40bn4kw/SbQKaX6DomLsJcThoKIf5epmkivkY4+SXGUHumqRD6/3AvI
E24uRZs5GNp8/01ptuK+ch+J88HEJXk2BE6g3CA/uS1YE9ZDliv13XNxTZBd/7ZA
qV0DqMhTW+BcdapNWwn2CBZvWhLSDWgZlH65XwSRE5b4Zmxt25QmO72LI/opi1b8
eWGI/PigzIHcIkMa4DwmKSiTB+qgxV4IXICrw6PBYs/iKsnAKprZ+GINjeEeWRvZ
gZOJmsyqT329JpAGllsVgmnEjlDlJIoWUe6vkx9/kowzp6YomgHeAUX/Gt8DkD27
0GC6lX8Z3kyUSQis+dSrmpcVAIwLlmEEnNJviRUrK0J+BcotaQKRXeMpQs6TThgu
xlgxSCIuURiuWNJp6h7NDLHSNwPlC4HsyI4D7AuF7YwZHKW+lnrXVkayHHGyK+qc
hbIqc1JK7wyhC1EDYV5dTyQOUzF9O2gybkX65W+77SC5cgsycsL3w3a1iBWLZag5
erxIdQXP3j2HBKk6dVuSJPq8oEPCbkJ62AOTJP2cn5t6s3UjzK963tK0jwMoGp3y
8RpGoiEA5+MLfWddOsRhnY6Cac7J98fUlXnVw+sedoc9eP09RHbqpQK4puzTr5Jh
2lydvZ2Su0VdYhHnGBqOlbUNykKI3pdDrXLHh457G5Z5iDi/yEMFHUjy3iEF2xYQ
PYSB6QQi5wn2/VO8NEqaNc0jyoHI0ppiBORR9T7HOz2QPG+FIlVSRFLIn8l/kN8x
+0FbTJRPirVhHBmwT1quWJc5bDmfPmsjsN/yhqXSW6zfRHGyWPEKSXk6gee/TrvZ
NW54L3RxHibBTtq5yFzrmAj3lxFCx7rEXE09O9jLyKXlBVxhLaD0kFR7/6ZgVqeU
KPG/P4Xi1eFb+0+WdhKbR+QiVN72lzF6uNRODbgiKjaromRB+J8UutOgg8+MZueb
t5+IeOpn8n9ZUC8YMZiFikOIht49yREhJJ3l30tYNZDrLAlYunAcIRneYIxapIA1
aMPLknuPoCQFk0CGH43he/JoubQIfwYgpzCosVRKAEfzNSe/CACtR+capWcASQl9
Xu125+NzlIs2Xh41zO6dHPr4hkIfPLsPlwrHNo+CDGpHlHUrEHCEyKuyUsDjwqkq
mEWS0dzti5UtJsK028Ipe1khN4/FX75J9daSpWp+n+TPedLXasiNov8+QN0ZKmrF
43fCYa+xUnnkdaSG8CuTFV3GnUo1MxNiesEh2x7usN78FM+GWGNwGJuLVkmscw4X
kBOuQRsoiwjbP1Rnkn7OpWLg8kcei8D69l99Vt3quJxMOtMcGSbGge5KG9jXSeU5
zUNFYnXgWADocDf4RyFJ3I2r8LhqMzAo9d6tPtnal7XoxcXvcm7c0STTQfByPxBK
tXzsm7vPIpJQOLwOgPfrypCuKeQ+2EmO6+js7tPBNYOKdbfytUpw8t/CJDpl0KPy
Z1ni07AFlSC0WM7vUaU0G1VCdm9sbK9JPchiZ2K32n+ltliPCXdGOAcW4MS79WKf
cpMZKoVQQYaxzv0ZFmOI5hqYPiUmTEPqc624zTtoxn6buRT1mphjXhCpn2m70AAN
2eaSLWT3+xWJIRFXCvyuntcaUoxtl5oDnbmZvBJFJ88hthoS03bSOfeMmeR5pb/Q
KqmHKQoTXg0FMRT0SP2V0suKJwTlxAE3lDRpb4gyavfU2gqaiSLBb65LCyBpkUGa
rQA238WovmVbXm4GatmvxTdt8zIsxsEO1WXMt6d2M8L2miw2s9+OJeZTxId+6XqY
eTCyObSh0odRLV0tvKSzqmprc8PBh8X6LRFZmCU8EIythdD9S813yBuTkoC5+4vT
8wvEYHcscvnw5qgRj/Yn9cb3IV/mPJNwBIdXTEFlcfFhHxyawuY0TS8D+8/+PLga
N6cmRzLQHc0+G8IN3kpuvr87unmhroxv0EcvvkocXp3Tm1Mti1s0ZHyavF7Uzfkt
OcVIKEhpw5qV4EqnuStaK74mD8gRPZWhlFX4FB1+y7tno0B/QSyCS4bblcsr1OJh
8BzB3wELqmrhn5665gJg+YWNT06pSUWmHXlVjvW1wP/paxYPpfqFdxkDfWW1jRpA
zAFD7I8M1r9Q1NLpZEHP8OeVJ/jE/YGxZh0aeaB54pbIWmDjZi1cQYzmnUUX6MEQ
MVeL2DZRGbFiXBG9Ulj0r1LM9AoUPwVp3z00ZmkiE2CSxOF/QLmQ26nbJANL9qZw
0b1O3gzDjB6es5BlZhJl5GrS9o8K0RYlTaM6FdVuF9jo+PHSbF3ujus4RM85Ke7/
c/bebbTXYwfkw3yuwYR+q9wzhd1/dalRinVjmrT/GaPnNR1VEtMab/gj17jCh/U5
XELqbBNq0Mj4uDCSj6QF2AtWl/hRQvmiCF2nDTsUGH+kiGl6i61y3PX7GvbS8kGk
lfdK/s5uRvZggNkhTiAiswHQtGTdGOkjsq0mT6KAwVrNeIurXL0Li8vIrG3UmIjJ
vpka3eR3ZyhylCCLLvWAhDiz1ZeiCUVs2e0hxxl0ob7yzleAPjn7tAHRRwl8DZQu
bUZw+olHWzpTFw65W5+IwaERJoC5mHpZ6H8KgxRUPGEOK+lqH9/BdDPEfhEKOKsz
UJwJ+lT9Ol5/ZXurFvGxIeRED5mkcKxVkyZJqgPlN0qPDrELDPJEEaBE1G3+KaEI
KJ5sdABqECpO/tPyKbevkL7gJ7iM5eDFSnpGNiD+r5cbGkyStoZiWORIVb7bPiI3
E0xSkROza38A3EB5M5X89E7E21eC0OmHfOA6LNKlZya7jtkIpq5ijFaG+7rGMn/J
sHRI+6geYHc+TuT3Sk6FAO4gZyNivy4EqdpHXix9af3txVxbLYhqS+txn7e2cDJn
kDn7YWK/PXjqUWmeYMIt88ux+B2f+kFKlwbktruI0qCEK40EBqha+4pJ6sBqk5xB
kXsPd2gF1Wf1r/5YIlivHSKz4fACacoRxAbOjmZm/xUE8Lw72GhATA5lR0FXrTQ2
r228KMJG/zTaXPhvWe1mloMtsaKZKXmbYlHiUvGwuX2PSBlXN7bgxA0Rxtd1HG9z
+G25I6f8bwaQVSsvo9mZBXN2EqG/lQuWbCgQ64QKp/GO7mLrBZHcEoQnZifR3nHP
+zMn5XN1FxVdxOpKsQonSsxTGLPYGez8fsv4XYM8+c5hBRtQo5kBYx6JVx898kf+
O1rvxiCSTp9SV4HtxZjTRBg0NrPo64SXoSAwe3UdOY5eSBA66J9MbJp6E0a8i+TD
zqRj/Zuls1rysBdK1WIqj7gHJos56LhygmI1Up8vmJqmMx7vq7M9UmCwIoY8C7gf
ExS0ViO2bY42U+er2ayEOkzewY6Rwf0lQyF1P15MWkCuXYYYgKnGqDwcKy+hwjQ+
InIy1m1xH7O2wziM/q4BIPC6Ai5HOxlezgDJrXFFc3Fz1Uf+L+qN5c9+u0jpLbbJ
jZIhiSOTbxwbdQahruRhtWq9+sKWul/taFbPjrtdxKJ+MBxA4YC8Aw56Wa4Xrhvd
EFRBDpgBv2jaxaEK6aZ6bIcmWYlHscKoMKFvZZ/MzQ6LB0GeC0lBcbtkwVXo5xJB
9vsgncdo/07U8nhT/2tuciI7+BlXUns9bfO04+OVPbS253ZzIw/ufPFEk4GNRD53
jIxXhWeDeMu4TmrWGm6bINFadSOX5pgWWL/sA6ICmjmq97GorvVNKZDxrVTG9oH9
jOmBZD3wcDFV7kDPIJ3hDjQljC4+OZufZhhxqmoVcBaPN3FNuV4COImfFi2N6lQq
A0AAGzPiNXmECJG6nFsB7FzCJb52DfWV3e+bzwYpv+d8+tDmS1KCUV3+DNq7b3z/
Q8Vhbw5JCclpj2Ti1eq0owHFcwSuTgp9qSOXP5F0M8MGqVZ/YN6Oxkz15wQIn367
0pLHB468O09o/ic/YwkaPs8KZkipt6XROt4SBcDCGBneMTzZz6eLoT/H4XH6z+qA
ac7H+2cMr2nYLIY7bHe6ULFgOmDtttqZg04niwsMSBy/ywLo98OXmPBaWLFNfrYo
F+8h51y9Uq4pllpe50US0ine+APmIt33d1RoHRu+DnDFfQB0T2FIQPMx+EEb1W6y
jVr+xYdMFL24SQ39zgqiD/xXcscdem+M6VJTL24tRz13yX5n0D5/BeL209D+4Ooj
b74s/uZ2xSiNwtlCQBRWVQattj6CqdKp7ICKCuG9RSmqVXPyZGEAsLbeQngtPo4L
64Eb3KZzahDFsi/6gZiQsbY+T1sXCT8Q2PuyO0AqPjX1KShglL+TUpdIdlF/oYjC
ipqxjavOJ1pfo9C3ofGUO06xLdbFGYOUU57PXhRIGYh0ZlJ0HzNi5i29SAXg/zc3
83ifXQ3q+/jUpomWgn3SlpHQKsGzkye7TNmxAMs9lYR9cBs8I97UCjJG2296GABm
IbMktcew7jm/Qt0MQZ46uZIfDqcLS2gUDdQOoUWDe9aZ0Th+ZXCK2mb3rL9SWSPF
3pq2C/l8Dl7GESYmrUMsd1aO3tBgSrYZFPKnDeHzZcyTMkPT3YpGW3bNqccXCvR4
9si1DNb8cby+DE2m/WdhgQdbwic4xUF8txGX0PJ7+F8mccwjBitB0fe2hdGXrisE
s4g8O3pp2bOUJJuE4KZQJ/xARohbTrqxXEuM3/ADaGK2gwKBGXkBBBaG0C5pZLKb
KbWIN1Z6LxTBxbfwyK6z1cdxM3uLYQqXmV9XOaj1znWutruz1laXYWiSnJqBOCuw
Ic883MYhQYttkGYzB6dBMNJMSGDU5WdeWccL7oxZxoheP0cNdfH+nTUZvdX16q3y
g4PEwXfAuVfKDyDKTejwVCooLV5R0xhHCM5iH6Oz+tSdT7XcY8C+RahFa3udiwXr
CzrMhBqg9YomKuhrrgpbGgg0WyjQtvObMz4zkyR8SM+Qa6YIviYEDZ8s83630DCE
nuMKS3oggMI/II0W2rNmzo/WcSsLd3zLK0AfAA8gSq0/Z+/ewJHAqt9J16nDXCCk
8edXyD8WCTeNPHtUeiwXF5Q2Ffp1W3TgqRovrm1RHqmPVO3hjvl6kb8WVcTHQiMS
yoff4Jt+HIPR//dJDLZIXsNEMYoO8Mk0OW8/ioVmRYTBE9KA9jfFbQH9EnkrbiTE
N3o8+Jg2AwLcxVFdoZ/yvdhmWMwa6bZuMbwcCdFz1Spm6VDRyath3qO3brfeWg68
4A2L0LiU01jxrYG+8P2oTTTie27Sbf8tP/Mv6y4gDyWEb5dnKclcl+KCcLsj96zQ
hGWAqC7/GjNFoFmeQWqYuWbDqdXNqpnswPweI9FHX1HMAqUj5zflG8eMD/QhJoqA
IEQt0ym1Mzi7PgwbjNMNx1rA/dwpgEbJMbsDWmRbNVRpHarUAaTmZGolbO+rC4Xc
vPAjXenH4gFXUapXEn8Qz7z4qlnEeVfP+H+LrAOZGyaloCuAvgX00u+uaTTSr5HV
aO9BqOyi7W2HzARUVKKiHZwegS7EJcQ0QJspWQquMEf9U0C8bmIq0Y9qb3qJgcpB
he5AeXk2O+ca1Ik9kIhaY11jDq5RAZAYEi6jHUwUskHJm/OHwKuXfHdck8QRk8rn
wBUjhN7rIAdw5DXjgHs/zr3DK8WylTANkyztzmePNgIFhGDwyc5yvUv0nHw5jsWR
6SNVjEtsm4ZDqCvfH1lqlcYtytaYX0nawUsCf1mKqzyPXJptr0Zw/NYe83azJvyi
hJw+zwOVih/q7mrR+LdBMs/qf6GfN0DBX3/YElq+0OlyPuKED6CH9x3a6XZQvFTd
8XTgBCCWhWWfhT2N53bO/yrdz+/DoEIqY4BHGkwUMmQdF/x7nwFYnk72cNQj3vFK
Pk8hMsKbYsNYebYZQFXZusUlADwQNo+nV/U5oDgwSec2Z3NUpzwySLuNKiWIOJ9q
ZmekL01PmMm2/g3LE/t4w/jSmxO9GSqtyUPDH7vYOOoGX984wqcXJ42PNjWju2xh
zg3T+p3ttqGLbwsHrxRM/zdVCv6+Ruta3kP8fkr8IVXswBv6flsMjcR9WQ0SkaV8
KLHRHVc9/+B6XmmyHT3AV8UCIagJyUrT1CSowkw8MzmaC16dNjvgN3L0dA7xtPcb
cGrFnls+F6eGSbuSvdIFgOpSXLkZgodEzu0zefuo8Uk1LPPWrxuPRxuLQRArxvMj
I6WtAtwoC9yGFCXDrORQZht9XZJu/9kUe/ZaVRRQXf3jYnzcwo3kYh8jTKz9fw8a
oaj0cjiWEc85KnH2dWPIKNgoY7pzI1MjJU2GVYuXWvHNwXeTh4fBMKOGUK2XeNUO
kz8ZG4/SAXTEYXzdFWX/IquBTjrdZnmQ37og+l64JpbQZon1qepwlBmzo1SgR+3I
Po77eD7lZ77QgrO1hetworSIu6fshbrjJB3/SJEfCd3KIV4CGb53bcEektNQjQYV
HvqozpNBQ+O0ygwskd1p+FYvv6uhx+zWKIuQmvasY5/b+7UGekSemepkSD17A0Rj
a6GBvcuf4UA0SJU4xRmJZuzxK7i80e9aVkBOzOOuLIu/wCcpn6bj5tH4L6/3w4lo
gH7rslo0KEdUW48JLlLcMhh8zqXp4J+RbgbzOEiNhww3+XOv1PyvJdu05wDpmO2m
s14XU2IIcU6uYsLTE3K3Uz/QtTP8JaxAkw/8I3SKeWt1ZUhtvxdDnUbBF0hnXyzQ
/NIwmPS3t4uWyKky8B7tpxoPOMtl0XusduZ2Vnho6JOHhT7ydYB/KKterhP+a0lv
6DzLK0zx41Gjul6l7iLY0EMS6vgGKn3NJb2eKRjpIpDC+XehBzWpe49k2VSk2uXa
ppn6tmH8/fphjZd7xOAozbxcM9wtR2xjHL3FRFKMTSL70LPlqVTr/Qtkx10051t5
822blZEeulE1KMWLcWhCVyorvV+YaGWxx11QNuq9vNFcXWz1PKqYUdua9E6EBNSS
b61UCEZDOGVDKPh9Dcw0rWEIQztUniOumUe+USC0PoLao+NnblNIsnz1bqUWsdFn
75ZFHuOK23Bwi0NZsm2/nwMjIz4W/5VahInrxJeJsmkhQsBhUg2AzSwm2FV5KASl
FcjUQKw3tjXuIuriD9bopde7xiQKli9H04bVyEfXBZ/W9OURFf454yaCSjTHQK+z
LwsxoOeqRtRCeUhZn6U/R9UU9vVAEVRrEmJqNCEG+Pv2iU93bBugHgjur6nM0sDb
X/o0Nc2PsNvNTKJrvCBdfgS25CYMeMk+Zi9VqSUkTT29YSPm5R/jtRBWUs0pRoNx
QWCpeTYFecsHAbfeHAXDDCUZQLZSholkvQCJpR12WP3fq+jL4tvCR2wUDu1npJJ9
U12Ps+yySqvrMYfoT6kaed/7WUvj5FDOGH8ozutBU3nR/3BF3PwzPpf1ZhVnl4xo
ikKW1bO8k294R/X00KXeloSYB0e55bh1TZ08iXf+TXeGXreke5y8lxxcrkeuYell
NQ9ATgJD9LmHpksL5zEKwkbWhNq8Ul2+o1ZUrhnaI1JNdCcCUMUnWTFmjsiikfll
VhBfE2uCBnj+jyP14ueaf3MoObKNb1Qge+lNHLLEglrfK+SxOjnl94EyVSra6R9J
f0jo3YLDwr4LNjE0TJ56xkPdBEqJUJCfiOlMpP7oOUpgGs5392EUnCjcbfGVJy1v
tsSF3aak9yFWhrUVRwJlEJFdy+0GZNy+iNmSGt4OCT8HWLTc62aNPYiyPEAd/BH0
VTJGB7yn8+1Jv6liAKnqQEJvSnF3qfu+p40A90JSzyl2Y//g2jXztYftZkJFSIHh
INPNcpEWYTNtR0mtevxxY+9Kr2tyLnwlIzOSC//L/NCgG/x4K7QfpYMV+z85KJ7c
FuadUvjazvStvTr0VZ15BAhvOEcgZwiciEk9LSF9As5ZCZzwkKd8TeLl+caNWR/P
ZAJXXLp8L3cdBN9QnwREzd1FHlssrYlN7EDvl6lIBcgmlFYG/juLuWtDnGY4baVA
Yu/KK0qYzDEwG2PElK3Uc0dfYCvg7eTNP5tFI1b39xulJTZ79SWJdRICo+QNkMUz
xLk/rpAOrAXk0HyAbEotqrcJII+OpImwKa6P4kxrXsneNV5sW+GepOIH+FCZDNfy
Ct8GSDtBDAuXKx1B6Odf2ETtgw1P/21KC2bgPObGJ9Jv8b+vJefoxF+75FyQ+VZs
NNkKWl1ODIjwvBQp7xRxJdAdvtHI+m9eNr0bHaF72p/YskGGYMKV+gHIwAV14aiD
aSwtn6mR3CEYq/uXvIGySbO3iVSDR7R0umJka5wa2SnKV6UvhmpKZTy5Mb2BCbSi
k/S9jRFlTbuWbXfgzeOWkE255EjK3PbFQRVPbluGy5WWNzWrR/VUbMFS69sA5ZpE
rxrEXmCaO60b8WHeDLHcxoLwP8OevFF30U9Y9lzK9GQYF0at0agMNc+F4rRUCujA
5k8TurkQJmyom8tTs1Drlgkce765Wu/et2TmJkE6f0DXezYFwBW8fo6QKEtnyfLJ
6m/SHv0wj9gROv3KJJ5+3i9fXAroOzwNlJRTn6+4VmeH/g0kPxR9WPgsMnUmbUQL
NWTx6nE1n82gbQS3Gbb3LWTkzaIHTqxwy+n2KP2vZUunCCaTB7AEGWGyaBrQjNoI
fQhJtM65fU9V67lgySWLLitzSggIQCof3KS/NbcWhtBIP2exCb4abzb0ePZjzUAO
+Qxk4XXVtDgGTQ2GLsw7ap66mD7308vAYPOdy5aEJiyljtZQ9niXtD/Q2JuSwEp7
QLTS29hkn122QikxBNBrXmbITJFvQNLLSJKJZgErvw+f4pgn3OhYqIdvG6kAN1RR
jZg2uFq9BTnlKDHFCkWt1KMVt6fgSgMpav4oiEu8/SwA3D53HIa+p79gv/1tqdLn
qR7F+WPWI1WHuHQnXXJyHuImxlhrqrkqWHCdSL8T/5tLfP1Sd5c+1ckEqmCZqe28
tgDH0qSTOWl/h2QlNPIhsFTyrkfXNfbf5xsjz+EM/qbOXw3hTxATZxUrkVd3ZbrY
6NAE1S2tuZcfzd64DQBjEStvVni64PhOI9FvftVrHTX/6zQG1D+JisvU09gsbAss
PLq6PXvsw2L2r7PkEi6nplRfJ8BH7iUdlodAKAekhoC/BUOkeOx9HTDb8VGRUbj8
uFQcGndaC3UguYhje6K4kUOzquW5S4ONbHmabVlZ5sFBOnXoeNjYfPCX0uAGe3HB
NJYHzTCh0vmaLX4zT1q3+WmIr++M+BEGL7pSdlalMWJEnqQoDQ8FftuA8HX8+0qi
dYSwNQ0+eV0TFzIHl2M9snsQSOX4FX+i2MxlNoKyhjfXQUgquxvMyty87nfvuPym
XmIJUDAwQpisWU0lpyQcAjATK2Yo3nPJCg7nSY500/wk5gE4HxWM1b0wi7LOFdcF
Vo9NaLQaAJvY990s/c0gdmhchW2KZIrWfLBZQua+Wsg6R6Ur7aMQA24RJPk5IX2o
MDN6r+aZDjQicbQErBaO+2aWrpum3DJObw7+V/0PnRvoq9MmnAfJObWg9plp8lFm
LphNqB1PPaA8S15OjoYUFP2CtP7tE5wWLCYH3m7FuBD2+//HNngsOjTmzGyKAOKC
ThuSc82NnZbtT261uc6bKqcqsXXOynH0z88zMG4xsbSGAV1+5PhR5FKRCFoU7VqO
FdYlwp+OeAYky6w1ldptkJKiN0fwQBE1GttWYVPPmuXEszPa7+YI7BQRr9i4ZQF/
HlKnxfdYcXkh9iPdneFICCqlyIcAdf9U/NPonywNuhbDSY/bkKPjJKlPX7/JKI6r
/2CA+uT8hK/qlAdoswDi4OTb3mGVsJ9sbHaCBpS6qV2lM9en/fAPZigfSwMYm8rX
/t+TwuST+Ou1eJLwuWU4zGAdpRKGIkcov2JWEfTtusx901hnGXFXLqcakTywE169
5I2eR899VwkpiZS/AOzgrwrn+5LcAdLQ5199U5m79+z7B6Ci8q8PXwllLRUZ3j7E
ZwHYALnGqQNvx0jxI7TQI4EUMc0cwnc0N6c2vn05xlHtgEvV21+RAIv+7y74dm3B
FhMC6mjoYWUZTnXLd+KuFg15UOf71a6ToRJL5IM0JaR1OmXNOn0I8a1MyBxdMVWS
BmWsUrA6KBFq0Fen/5yjRyF5qe44kbOSue49ziMGVdwrbnutB1sB84+p32ZXt9SP
d5Pyilh49O9+g4yE6u2I94/atY4Dza2h/x1RjNx96KdL/1KAKp9UFCmGP07l3Z3/
yR/HfeiEfZu4JzfBhAvcEN9/SG6rAORl3mxVPMvO4sPQa2ZjsNDl358TE3hcycWg
uyArIjjT+ScjWUl6Hi2MccZ8VcLkpp3PPhr1HaBdXiLGTigssm88JZrYFAd1o5Nu
EY4StNRRe7i+NKI5jumphFnk+adlcLqu74nBUX44h8KaObig3XrFCgJIDAYOd6PQ
qpcPb5DPAwZ28JqWoziGEimAdmH0ZZfHSSTtHIwkfWBst/XpJdefkeTI26hR8ain
eQXLWiRh3T7SfJYSzFvV/iYtt+piZ5iZaMoPeaWPpIoTlUaf66OQkbcU0IIDZRvZ
AumVqjR3wD173esl9vuqdGUiHw9xZRGQQte8oconExsVX6hbZeJQ+GChXUoMzKl1
wZKfg+AbTgZ5Jp16F+Q97TUtKGWIqjnzJdV/VEF8BEmCjKqFPdQmQGwPeonw+U3Y
iLHMyDNhcf0GtKp0kV0Ho7E0oad2ymMVOIDWhCKH6Ntoey1mJrkgfvRAD6NcBJ+a
IYYkcS1tw4aqR80ERdjfDdupppPS9HqlMQ1g5smXNSwi6U16NgP1OVgbhJdNiFc+
nMnrs08MJl2XGoGcmM4fFkJ6XQRG9M3H5E5SBcZWB5XFfuvyz6GGkilznk0P8FEP
tFYoNBV+migrILR4C0qQvom1jUUCgi6vfkGxjiBcjlwe0bKMrDx3u3sSzChEkDbG
5y6piR2VGSN0+GXlMUpA3bW44FuVNRkykYSI9D+7xCSDR96nom/vOmCtpYUZwREK
d0dSkopm5/7AwW/KKW96w9K7aB/43eDJon0Y30+fcMfNFBtAAH13lyLmDQ3EqH+l
drgLLYQK/HWig75fe1AcwQJ2AScrw73GTqo7bTKP/XW4VHdBVGJIWlxvEPcmTOQ3
tpMxyHui1YCGHyu4hf3WSbBd3S1iDYJUkX/pvEziAnJLJb7ZaOqBrxiQNRlsnkPO
m7xCLZ2055hO0JZvIyN9JjJHZfnKKWhg+NZmsK4YHywLK/1q18wA/gpIIPG1kIL/
qVNz6Qfr4cENmHj9kKc7WLhKhsJTHoeKnASgBz/y8ZpTAvx9FLOiPUTOhJbYiJdi
H+yQvNdav7jGA96Ax/vge1m+cGfrYW+B47F/Z8peYmjnGafS2op6LL1llUl2DwVT
SQakT2wdEk+Wm28do/YObmTZC4aOkj5pvb0BUcecgLbgQynUye4kgYujZyM0i87d
pwGsMKcCyjGYylogS9nXmVsOj6Piwg64Gv2J4uELhbf3jwe29nSBrBu9nBVNZttO
cliW4gLpal05KS6NuALyFDtpt9MA3P2PZ77fsIbzHxlPUkoJkXFqLGKBwgYVAkVv
9FFKzFQRJFKka3p6JEoxHJkD+3wTmV8I2lGqskvMZMOe3NjuH6ELU8RaUZ7hcRD8
TqP/SRvGMmVCHC4Q/z7MNp39+WFFTVqb8XgifW0Hf2aLJHI79XZTiiKyWxOIi/M8
J+dkTvyDz7moNNoM91J1P3i54RXDrHqkxFa9TObDo5E2i1qUZHDhZWmWc7sk1oc8
aNif6P8pGO6WlkM6ylH8eWBRorpnSLsEM/2VzV114NuFRwoYCewQM2JqqCveG64u
ME87q7zxils0L2svlxA4BK1bYJ4y8hxZufB69Mg/ZszC1L5BG4L7pAQysE7jNpeD
sQwWiRp0ja0zuCNcaLywYJtnFTJCndkxlJwMjS1MRbfyCiVsbcSVRnJHPQ11M0tz
kve4063btATtl6Hj3eZWLlHH4f/tKBJoAPa9XmF0hZVnlq3GsIFyaouMxqMW0fCo
uiXwWsu4VuOll7iO6pnH8FPcVM04x9hQdJVLwRVywdI8l/IUQzhMbqiohBlDC+39
Ol8c4ffC+THupmhGfIlixckrx3l295jCVD/yuJUT8cNQICEyIHmzpJJJU1d2o7Fu
DRE/0B4XZ1HsD+Se88l++Xut9VqzUT5jchmgjfGCBAFXdRO5Jk3KI1lDNSs/nMse
ztIgTGmERVMw5MeTZyTYdvEiHrPpgksiNn1golUh8cSoTV5B2xKMwsX66jr6eqSc
FR99JDgjGepPlsYaAJZiAYstXrlBP0hPaFc2dSUhddGFK1Ty8XBcHjn88YBA/jM2
Z6AsCC9Y1IRltPrXl2I9kD2HK8CcJG1C40pVguguiR+TcoYFWenliyqRXos4DLLy
A+ql3+0lBPzro9jGpsPF+/tZtv9yX0IujfX/xXqzv+VFi9tEpopi0BOLm5L9oAUZ
oJjngTu54VscFmDQce5nfj6syGiOXLc0nPGndDQq8jcOey7MmHBs/m5IQ9LYetVI
A8gFQf7/7ZJ5tBew4P3niCImvsfwPsAJKaGM01EIji1S7vyAcBVv3lJ4vTN9eJDr
rQbY95amgnuRHSatCLp2IEOc5onrZtYK44EJIs80QHjqC4Kh3AieHv+vYjc8gN0g
1W5KCOjhoe3UjrqaNH3+FmwoV04R0GEWBPbyzYlDFqj613is57I0UtoKyDwV47ak
mU1bVPhfssjz6qLH6c70HjNLN8rsrzN5g19UxZTFiMed+cZjC9dsZmVLTooAMyzr
7fsoJAIJw2ZS7chuCm+w0cFJwHl0NjG0HHd33mFUB4pWbeyX2Wn9PLgkaNAxZvKq
FUKpSP2WYpLq+Q9U18SJm2i1gM897kedycxWCxMFfZD/417bZFn0x3rwa6Jxs/h/
JWCbwq69svSp/FsmS3PkP911BSos6dvD++kOXxlhnV9m2CxNLynpTLzJQEcmQjIN
1E+LAjEPvmdWVIkPWFIT/f3uSdmiq5mA8l3FtHXjDsuIEohyv7QdJ2ouptLF8wke
R2oQg7CJu6DcljLqxE384IzpAKavkLOAKlaSAFN84QpDRIbeZDEnQNcAEX3reV6L
0u544HYRVHFjYDTvp1ODyZAvLaDayM/tImSc95StwQGkApebfs/pghx5Dr2SaM4x
omR0xPm6fvJB3U3tvhWYVhHKSd61/2O1gDB9KYe8hgxFn05TdOcyQE2ke9dKJZD6
1is2H85m/5AFBU9E2cH8XwVn76Gl64bMl9HzGO7AlKShLU8adcFQOxXP86zPXLTW
Cmz+NuRcZMLAJtvTP2B37pIWREyxvkK0adP13Jtks35eFkb6JqScn3qFKhhiGr7Y
lHWSLZmNa/y7Eu44IXDzF+hkUqcC4dRyTFiOY48rXv5uS5LJrNvgMCxALq73hjuQ
0EnA6ViW9qSDNP4Tuao2NutP7nnUghzZ61vPgP2E8+s0hTbPvCsvU+KA2IEwWhRq
BdrrOvDYkkc1VeSbx0U1OASdyEcbgSuUAHASvLi5u3hjPEVcYaF7ZC+dU00R6azt
9NZxakb2yPp5HKDafUEJKemhaXhOAR9T3OoeqexSHlg8vzMjmC/ehxX38iw5HW6k
lwrMuryvpF/rPdMaYV96x5D1T7fmB57IX8qYAll588gXvl/FIGsIzAwpRAdObnPo
uR8RXgVEv3GUZQd6xqLUTfQIM4ndkqkEcGEAVKCittJZ3pOsYf/fVhiN9Rau6q+u
GXk/WHyNS6s2fcgfuQKZ7bgq6e5TZi1StNcX9XLkj4hwCvBr1/L+Bvs56xip1fJI
r24ZFVp6mYxhlS1IqdSv+kPaxW3jinzah9b0GL8Z3iUQWBZ4LTJMcoBpDlf9yQiT
yGNW0a3jeC85mZYsVKUD12TinKBEachjtM/Ls1YXyp5Z57+gfqHitAnEvvpOeIoC
DNTLigkgq5G89wypDiDJ3Om8NPTYHu90zjxYz9GvvoM9d9S0wEMHk7DZQd5LfA4d
hOa2+vofN1d9YxnUc4eWVF746UVn+uXhIaYrQzLJpQUKTtjiY3dHxgAlBBux1mbL
3dg2xY0kiJYWy5ava19UYKIA4n4YwWWgh5c2nReswF8C8uxEjELmw0xYnAia0/7b
AOwA8wseUM0cVBLk3EhaEDXqundFGOagRGV+BDb0WE1VeIcdJJtIa9eZqtgCkQhr
FHdAiAd1YXpn6NEyXsEguFLvyMa5HBwCQIuDSZCB3tf9DC1HAmkBTUW4vHDWCyhp
s88oglKtbvsSdaIfrQxPTfZwrBdsu0L6KiHwHgx/Hv9yNvqps57dykCOzMPzOKW9
NmT/vYFf5oFdGuI70DAA+fr/wzBIlGZ61ECDvpeB8pxt86RhchaZlqQT9EXCjuOk
8VsX2Pr8eoRtOLljcbXYGer/BaizVJGkM978he8L1ViSRlQT8ZCFppi52VIdh7LO
bASPhh+EqnVo+PPfqwDB4YeHRrplgiolAKrQJ+H5DMMaUPkVHkGC2l41EqJ0LzjB
mmr4WfB33v3d9xu3qtokpJo5Jwmz2UMS0+wGc3Po/02/AfeL/y80Bv4d14VE9lc6
PK9Tdbbe+Pvtu83XXyJgtB78B7D/w2H4kZD0nRWtWGrjb5T6M6qpvxwg474ZAlYN
DtL4Ww2t3zZTlNxzQCwpNmbCsBYNGCYlvBl7h8lTZ/ssI3Jd5rUa84XmdgFp148m
gTQt0I7evSmiHkVEDSsgrFvNlYJK9J0AI4bsnJOXDJonpuLtLUleVUEDMOubLcWK
wj5T6kCmX0VwsGUt9RW3u1lDsRRIvDAGAh6JAozWdbTecottz9nolVqFqAVqj9gG
Md5wwtvo1f/t2/SnNTBXBZsi8kp5SWc9sKgpPAJf5xLU9fvrhmDUuqNET2acEP9U
14wonvT7j7eWrXaYneNOqDa+JesZkReVE5TAMo0MajANuB2+tjOPbh2hINRUrKTM
grkimXYDlrWsV2lNHO0oX7tOx25CAhyS1x1md1gg47Wtf0J+OqCf+n/kur8BnJza
5VtWFAXZmFwiAyY6HY66jTl3KqcqNfM4hS/oMlFrDfMtcUycLXeID3jOGoRZDski
vsdl9dCq4CDCapJI93ToC/cq8P39vZjjiQIGU2EP43zrwhApWxCUawJVXiptAY9Z
9PqSIDrGQJAgoGQZzJ5aPj8c7kBZwVMpPXVhnwfSDkRMFyZ9rD0oHcAGHvo8+Fs4
1O3vi7krG3wQlpOJbr0UHuLZuUCi7XMiBIZMgFqpcn+fEaw/9sNy12sWB45M2OCJ
0ifdkeAejKYcMFvuQPkyUPnmLAP8F2ujnbVqQU/zjyReBAWjvYcrEzxWUuUMnEJN
Xrps6mZRQC05U5vvAwwPOLqmuoRi7I196I7schESJDoXy2q4GHHZ6d7tnTFOlgg5
HBh3uLQjR4O9UQifHmPx7vk3mP09XrZ9D3WxUOhvfMrT2+wGVrl7TN6Rmp9H2Aeg
kMdxzSlp4LikcLRoC/y899W5PlYSXRFN0A0RvsM2QdmjaV2kDUJmL3hEn/kVam5U
EHyM0DocIiKtzANeE7B1d+Tf0p5Up0SsO30Lq7H8fATGYaufl5YureAMdOUijkEi
Z+mGf4pCRCGPGgXIfUHwV9xZtvc7rhbhOujsincvL0DwbPxeE/8+nEJ3NKSndDBQ
jeyk0TcncNodcaLplVVRwaOJGeIxOhy0ry8DxaiUJyRuK4x1t1V3PMA9X4eqgoPm
q7i8F53Tint4+LV2P3G8K684WxiN3GzSbCG2+Ckv3pDfeGJYbbJSjBYqQW4gV5ps
SlxVfJr5Wj1Cp4zl6GpwNXGE3sm2NmHX757nNg9YwH/qEUVT5zg4rqq65kKGIBp5
hUQ2MoymjqeqsWbS4c/7HjSH4YbS+oR2LuiRW4rNsrqOFy3n76PQMetMcu1JhRxW
Onymc4h8qTU5/GjHhFfSAEwEbDgMTJ52T6woNivySvqsIi2kyto+yZs1IbYwy1tS
yXEYC9x1hEp+6Fcwr49jkrK4Yp7/yFUln9KR0x+CBnzLZ+1JIWIEhQtE4zh25fOD
RdjMiVrRaYH4zWvUdPNK9RVTgAf2cr2yp+GapwqMfBpv6yTlq7Eiw89eDsbitNyE
JY71Lyrz/v8NSOIBFjs89eqND2iqZP0ThqsDUqOVC80RhJzYK+CZ0ikF9+1eJ6Mt
jq05Nsj7h6cRayNPzbD+QBDzfbiIv2FkZiFJdfq949ZhcITxjd1w7CG892uxl40R
7E6IN2fJf4A72lTHerLFfiUOZZc4XN7+sYCF5B05zjdpIa1npHGg6pAGNx+bjrEk
CocXcMYfTwfEPWshx6LnZ6+KAAZM+YzIdBqgBIz4hox7kl7Rd8mzEG2NKVKxtkaX
sTYSfAU/8bxJhVLuu9Dok3oGenx6052bj79GAN657xV59mLNGulCAbZUswV/OnAW
0n3TLNkT3NsokFy7pQRGNgxlWKcvIE9ExJzw3h847EDhqnuOFmuY3oQfOoWdCwek
BYI6rYEBE+zTWgk3SmEumsYS6PFBs/22l6+omRrk/2paO6BKwF+Ce97yElLdIsCQ
HlymbIWweo0DPdbp3taJo+MhpYkn4mapmQeLMRAWOBBdsx7wX8+/titdt+v6X4dU
UtWc6Vpt8Ta/mCZmBEdTP645T9BATJNTsWw5skJHWA3kt6jQXWA+a0cfJVxG68WO
5gKJtyIIox/nZo1Y9UhMPhWoug8NOBFpaCE5YAEVYVnSDtOg46aEdW84uwZgPTkH
i5x9iHOQAjxZXBnLv64qQf3diq6qTjDmDTuFnBwgbEOCD37xFEdu67kCjtGjrEnG
K9+bmIusPF4WpJ/S0j/JGNDkFuhz85YYni+GxZNzLJDVNBCmTF9D/J/c6u+SrwN5
eLBAt1Qi8dVhG4JDG8rrkMCps19PrOlQeL6RPI8AJDJ+s6xVx1nBNfWckz8D2r0x
2imtzq/SupfjPKjw/V1IDXjjENVP9LLQdwLPZrWA+UbdtVuK4giLOxjW70yC6XG+
U+aqnDQw6rWlwrrn43oG/TcaO0wtLU6x5C3LYxw/NKjn19pYVxbFKvj87NRLxedb
8yy5pTKDnsfudb9g8UJ8RV4Q9IQEZdOTadt8Jd/K+Onof4KhlCYW2qzvAiDIs6e2
Ra4U9CX/gOVE31j45897b1cwkWgAwp08zyyjbIK1FGtaiC0yKeEmlxjum1rsSJL6
5OuYsfFc6WcUJ0bNDfpYzNug29MlnPD+PrQ+kHp62yubAArXu6mbPwdZZqBnSE3Z
r8UH7KMak/zirebuq0NiEqHj98HCU4TrABw9MXyrnFUCBqwpyL6ifzTZlXWVsawp
qYChGKtOH+sAw/RyHabAC2WrX1GgRAiYWFIuTTCI346c11tryeaYkxouAzJkeqZ8
d1aIPYtEcFGHtVPPxvZ45NvpvrudbATH27FHsoqlmhb6cubjPfBobYO0bz2nyKnS
RG5KiosAdH9ztW+rrkCUpaU+AftU83qMRBsy44cMmujUdMqdoQEJFnRDqPuqIcRF
o25pDx53WYUq2O7gSdfWKLzClJC1VwrqbRl/uF7t3IkSsGw4HsqoWsQR4dwap01c
8upQFvVdAUJDjN3QIjUveBSVK5KqsbZSVQJaN78UEuhtATRcKItsIPn2T5fH4OXf
ocRFKfmWGTMmjZasH1JcJ6YIX89eszOOe4Kv+7/P8yMbJBlLq5we3mY98Bvja5Ac
xJKFn5X17GQlcx0ypmOhR7VrTZ+3zEI4c2ITHBHweDmpmyIDRrjIOR5YSnoXI8Nk
rlNlgMeBCxj0bCV5oHzfdmnWXayvxafDJ7iYf+TqaifgCH4lIh2a9sHN9cXw9rIg
lG1BNY6AiHlV+IkIHcptQPBHeOJ5JwaVaW3i2jbT4CTLpxvZbEbygShm9AR5/tHJ
GK5SCokzPeFPS2E2cEyeJhgwevYpzDVM7/rwtWe0oqKeYnzCB7QeJiVRh3IpzJVl
9CBwHtW7Fy3XjxSKOqkBE+j2Rzvx4mNWyTd4IlplVOCqBFrrcbVa36BSClRcUavR
3gQbcgBIAhTX1n/Ec8XN5W5ASAUW/hYMT3UYf6xNwrR/eBGmu6/rQfQPIaj2GVjM
zd879INVBRdixveRoMuRXEarsdkd7+aIyqQSXErotycn09g2qqZhj4DnY60Euzxx
uiWh4hLIsQ1rSmB0GFwMY+Z2dG4fWKElBx7i0QtCrn/yCRzan0nWMGjMwtCLg63j
TTf6YErnN3Hzurn+KGcP4CRuxjlwq7F+yxHTCX1jAWoQuUUmSyTri28euhlxxuLo
FkuZYn5pNLE9JltEQqp5JSsLQAEa8WXRYJ6jVBJqZ52QvmgwH7lm0f4qliFJ01hk
Z4jrIBnXejuj5XhPmCsmHg73XdY3ZLkekdPywbpxKnkZ0G4avgzENnW0/eF5i2Gi
7suZKQEpjISIrz5oo05R1Lrr47CZPqskBwQssAurLA6O5fu8bJCvdgiNc384k+h0
OwdwsMxY8JMvZxkAKUqysWANSJVctu6uy+iC2Di9OX/KqNQsd8KwNc7RBHkHfkZb
Qv7jKHjSUH+/t6N+7Q93ikzY2aqHoMtrnC7Ovhdc+p7mwT2JBNHJpbELVt/OXtes
dsTTPNukWSjUZOf4t3MLGp9Sj3UAuoqriu7wKd6GGHXiYCZnoE5z9N0Jm2Ip16b4
UeY05Nnm4mCxZ1+YsuBwJsRjjqRh3lquZ5GaekQKN0KBhvyaKNOMY3soKV5zEMKz
+32MeYzdumUa63DjRn5kl3OEqRN/6pEnlLe1d0IP1gVCPyyglJ5Lrt0bO6JHL2UX
w6l0KkuP+cbEwSv48NlFrS4zZn9MDPEjdY0eD9us6IPLFeQFLgjY/9sEPyf9OmXb
fI606lPn3B4BmPMjcCbKHwPauJjejX9ZiBMXQQwW68yY2mTXSyIbx5E3nK3r5iEc
O4PLUqWJYTm90rwKK71WBIZE6OvAWppHtPiMtXIYn8nd3eJZyresDS1HIgu808ad
B5eolRxZcsHh9yiTOTwxVfW86U4lV74GXB+MjgSmQU9tYfonbg//MEPBN87GGJrL
IrPcwi9fi3B6/QT6e+R9ubiktBXkkOXUFoZp/C4DwRnnHCMv+dYT1lvDaBDdpkqg
OMxNkNh3vjAhu/7SUzlvEK0ZfopHbAWUTKG06zA+Fj4I45TTbHp85rOOaL+yKBTD
6/8ePz3r1JrtpU/fjGMs3v6gsRrzQUJlKFwQKUfTIHTJivca7s8D65g3InhcZBuF
XmC6Sa04kUJjGKIcVYpI+046wD6xPQymDP77Pw7BWg2E1Rw3PX6lUbVb8AYNm5C3
HxdDaV2fg81dwbTgpyyBK/+SP6WIqJ1sorPygyAWgbY7czcBWwr6AnKyk2k2FBi0
aErVZl4yayG/ZduSkOhMasMa9zJosiTmIKmhoQbqTP6+BOJfazJPuOCfApgROAa6
yB0l/za9R6xNDPYivRcRuvT8JLkXy+Ds+6UliHENNjjSP3F+uOR8FuJBBb26Wa9d
8Mh0iZDfBxlI0p8akogTjAp9bj/c6VNiq4FPpGI5w2i5jrvPYU+Z0mURmqUZfltV
XUX8kMPgUnxThnx6WVd3FAz9d//m5atLMshM9X1wqkGv1kVPGPaWD9mxhq+Y8ipB
O/5t6F2CwOZaxySbUiud+YRo3irn+pKiSotzWin4KnFcd2NcnvUEsC7Qy9vs8eFK
ZNkci0vzAhnOBnrm+wpgYMOBMjMbqiNVbnY70/C4MtzsUvV809lBIf2L+HHmYSo+
3tmy0hWW8lE9vqN0DyAtzk2RshO8ku9Asv8to/N47GRq/mic7FD1ZMphW0eotOzz
x9mn7i5EyGXEgL3sFdfrMs7C3WodbVg/D4W16MsZ/XC16h068reIomep8sVBtKsL
2awogjn4dtz9xCgvUMx61u6jt1Va9ySkL7gAmPDDuVZXfzb5eoDqxDMme00rCLwt
/Poo467TcC0g89osyJNY9+ajHisQFlt/1QcuM1eE874ls+7KREhlXI+UWbmqsMDz
68GXOnQwOxgKtJFqly+nOTZDDJP09Eg8q+0Ej4tHM3/xL7DyHiNhahmCa/9W9Z+u
oQ9RCu/G31eFqWhUew8MQtF9VZhRiz3XHND47hX2XmMCAeIV3o4P4jbcZt1VsirN
llb0u63bTkyIwhKs/0Zy+fXvXdkp5vHr+oO5+dl6B5NgaveQoJv2PE/KUX2cO7UZ
I++LgLkm8CgeNXaqOcUMPU6fiIMP/13snPmo7z6gqzK2IzS+aRWu7o9LklWPlHS3
siFZlpHONr1l8cMMghOBtVo/IORSK80cYCQW2qYpRLZloHmcFvNZ+I4UPCrxdGum
2v9sBzk1vJBO4hQQYD0nM4vhxw+tn1uuSTA8SJm0TU8zVf4arnugPVTQln8Dq98b
WPtWmzime2jlZ1ZDU1AS6hYJjo4MrNZf0224Br8qgKJZF2T2InhgSjkohB96x3hj
YvkpBsLbrtBLcqEKzXWfsARGLQ3BOPh9uv7rRs5EEeM+mkpmlomz8CN3EQ7J6Sbc
SrDg57Obwqm+hgWjhTzyp69vrwj0Kutc23TdjVZj0srcE/aOpbK04OQ+bbNtW4yI
gCs3MFW2Y1s1ERXp454C7lfCfsZzKHUvjzr9YzzPEzc8Mt5pllhU88BhR0H7kmy7
b0UYIxa0uGeQwoS/sgwdJYiYCFPxmZq6FaNI9nRug9397yMlLxJqoIiGMmHITRZM
rkaRPsisHA7Tjtkmec8EeuYXSrcV79JVCB52RkXNwY1BYMJ4VeRB8v9J18mWepNq
WdThNeoqzv8aPLH4OqzYB4CBYbE5F1X3bOywHDPJM5kkcMDr8jiENlKs8KwJ0y8C
W6jfSYSDR1Sm0IVn5JG8GVjU0p7luSxyI93maan6+14Fc/9fJT6XBkdkY+enuyol
iMc1ZwU3Jq5Uwmjh9gIatXuPyQJ7fCw5oCcGkFo4dXRB2EUg7dDA4j2NdXPQHMmI
/h1ZYIobL7HhaezreMKVPQi9joMB2ybb1M8NnkD/Bk+p7//HsBbn7MB3J6O25uJM
YyIRrpfCR2qtWoEwberzH0OZxpJeJbed9OqlF6T3/97B6pE8vFZPhKcLbSiM5o8i
E1xYKuLAHsHHp2eghyQgJp1RVkUWhRaE08YiWNaAPfA3E0Y3K2FKxbm9TH66zOK5
/7NgrCbxll+knX2yPV2A+s9WeTOqOUioERWfZF6Ahj6Um2QWDv2dAIIuMn006tB2
mMpXtk/QS/gRzCljbsncIfl5V/yp+y6sM9taJ3tZiEE4u1GsGt23TbjL0TmFQolO
e2j/tA/WupsYuLryq5//RfMLARZKSkMtAhpG/QvtD93Ihl7/8jkSEMitB9zCLKdq
5LZBys90hj8GBkYwWgnA8ZB4IVcq7W13ZrJJCSmzLsC1MM95Nwban+PoB7/OhYoC
co0Wt1IoCCuG+sk56pLb0QUxirVQRVgosTPfZm0s6Ba21O0tK/2NgRg5eMT72EU1
huwooaKQ5sW4FNlhISawaANH3+1XgEB61ciJYdb3yYBNenIiVwEleNOBZmyNM3rV
46JHUO4+mcIblrAkQ+mkjQXUn03MlsHbeNaSwqlOnVCX4Ff3xvCIqmJlhe+8uUWd
GmHdoa7jAJ5hcEs3EQ9WSLZUxMuSpYE7hcZERZfArsLNo4wbN4y/Eu7Ly+a3YXLm
nroNFGT22+1whWnmwLArSJYHaNY7Lom/nGC4GpqyZhUCrJEJwoAnY7AiWuP9OGps
25iulBh2IKxbY68z+pUMzC88E8yOPXmR0BVke7AV+gM4Y0Dx9NYhl1VZ9AmfwRQe
bcU0J6dVdE/kJvZqNn7VQ4fEa+VILqbHSurt+mlAY7mR6La7dBcsvzpDfY2W07rh
/Xkz/8n0zmUv4UIJnHapOep1YglUoKCaMsxb6qoeqhDhRcXWyNnbppF+tn2/sKVb
Y+VmwrK3Wj5PZE3HEuM2y46xdFsWYAy7hy4h2yd520HxNJB/m4NsMI4zGqyN+NfO
++ciYkQT17oC+fR8mNVX40kPLhDZH4nLTgsfQ2Zk2hyWrB4ON7k6a5EzA6pwPtsA
pfg8x64PBNCPAjurzzuJakLSexsKaQWjvNTlGNA3+eir7fqk1sx/hXDqE7BCW0lC
EuOXfAo9WgL6D8a3OkiTM5Z0XIbnfEOi5ZLTw0bdErwlcIkHbuj6v7jCyQ+4LvkP
EvmsGKiM8hVYqHcA3SEqsqi9TtGgnIIlE05oyNiQSLY34SRYCP+64usKeHDYaWDB
UaBQjBQOaBpsG8JUEbQJwUrI0QZOhjvAZ4ZobZDS6tzgo265Ssh2FDybt+QyhMpc
/2X51AFUZYZzGaPU0Yn1Qv3p3hFNo+rXqvN3SA0xjTZPA5gDshKpPDX2hVDU1qtV
CCcp/kAu9bXc8ZEBC2y9XcFpdN2kS9PivfEl7/wA7f9JLK3G9Sr5z0zxA/8O7Ati
SCNMYYLnTpj1ae6FywWULIaIjtR0lpT0pVyHmNTJWpkpMG43SUEon5u/0727l0sF
oBDy2m0KD6B2Un+XP42Rgg6fykI6pA6jUTSO2KGdHmH5dYEKXgc9HT2CthBh3TDf
G8jOimDYU1u6xJv7JNmPnpGFRkcy3Td6LyplC/M9FkK2xLQPAFpaelzKFAZkxqCU
UH9DbIqUs7nu87z5rA1g0LzaudmQUbDWWELqm724JBKnV9wB+SCvUZdeE7UC+cMB
Lrue6VcEqE2LEldPNPogdlyFAl1OJ6uw0cb/EcdY69a6HeDLj3aUTqUrxeJKfncR
aAjQK62VOYMfRuXU1YlYbHp3EoXJqlb3QCGkLuHtf60cAABGSKxUow0VL6H0sO6/
/SP17dFzVp2AotywYBG49ghgcvGuaVDunL/gtEHjPFQT6moiBhi3cuSbPv9PbupZ
ot0J+9IJmvE2oRcvMWxEvlpH6DgYhfy4HqymQIC5GUllgESLjrlt2Jj3tFXOuTWo
pf1JHBWf07kXOa2BO4Ayz/gnqp4SAUxF+BxZY/IlJqqU21NB55QW8SnGnliIVwWi
6C8UO7GAek8gmxLhpEYNPsWRYRJS2MIoBgRc3Qd1iLyax7aa7FYMGZRpWdB2wImQ
9Lb8RayD4Uw/+PvjEbbWChC8KhMGLryOauoIOm4/yy4arFT1gKGCzgl2+v6jKHO2
sBME45pUb/+z4shlMvLesnV733ztN5giZ3/gFg1FBvm2nKZUftX4DFZagunmCqEO
JN+Oeh/BTCDPbibmOYwPVaWAYq+T6Vyd2Fngm3D63epxJWtbMQq0wNlLIsctmoI+
l1KWxw0OToaUHuWlOgzYBosyk/Badp2Mj1ily8+mqtzKb/g2DKONfP/2esjuob8k
oNsoLsy1HD7CQDfNyeqcsybQiv7aHdw9KnWvOgPMHjlZz6eiyGUpSws9SmJevh/D
bglk0a+z3+Gdt/Wgk3R7jFwJ1MUxj7WRlhYe+evXzfQAZschKXbnhV4eE4LoxSvU
bmkBjD4x7TsQXJWEBI8NmBSS5vcM2wqcWtxIR9BtBvYMbqUJ4V53qoY64gt/PA+E
wFY+HmLJml1ayW0UFajkdgjKh/BPdqzd3xEGrShF1+JseZL9+6rdw2tbZp/5i6Qh
kxhk7OgtbzB3GAxxaMBPA1L84nAN2EOpIjiIhQlYSFNU7fnT7BPBKw98JmM2tcto
QdhsZvH/zk8zk/CoTm9/2If8tJ0P9NDvUiGnSSXblqrBftuqkq3kuy23mN/riQWR
6wmOinLA0k9b/TxTG/ZqZv8txEf6iGWe5vlfMK/shdkDZxh2QPbXKCa2Q4yaEzRe
EcCd0Fp8OOGxhyoMVwr6VpwUJEOuwkgO6v415SdJXWY5HMWFxnUJAmIT7Zfwaz9S
jxnuwWSOLh0u3tvOuznrFneNytZTg7pJ4K3aZ8jmSwxlAKQ9QSrw/ZcFtgn5XMBK
DhG2ta1YmhCl4cPLtPdeb9vfntXI8ZmFRrwi4JdUJh2mx6fzHTfSt37i32Ftokbc
I+yRoz3Nrm4XyNhNk7fQKE/7VZm1d5PiBpCjadJ5jKml3Vd4Wl5FT1MBRkytAnTf
osEagBXIG3JGUg0RfvhH8DUGqPgzwfUfsGGpM2unuEN8IEPsEhAEDL4Tx2j18kz5
CR44hsbQs0DRV0RKK9T1GfQsfETtYI/hiuOOKr3gfUVvnjdmmwa2j1ITux1PiJ9S
+LNtW6tKoRZYk/IZA9YeNxmRIMEK4LcYiUJxE8I4mESzAIRsn9/3RCDws6SPq1Yn
6g9uOsCf+3EW3i2/14L4m77US+zzO3aDAmwWOen2imz1NREybzIW8nc/5PsgJEpw
48wqH+b919JhVTDxaUGeLO+hl78fVvSXrrxTmkJ6DDtVfE4hv92Mre68Rjdz/hBb
0LKONjJO42BCmujfCu9/HHff124PES1bC73ZpDSyheAyuqqeBqbONUoFW+YEsxEH
Nr8Ak477qxtkFqOd3v9gH7x7hU923pYktvp0LO8O+J7eqD9IXhjVip+84eqsiplt
2dxOfmhr6MgGTKECg5hRoXwqxEqtogiT+hTy0nBxsncG3VJnz66xYzZ/OI4GYdf1
UlUUOqfYt3eBZw1qcHQJMngTRN1lqXq0nJmkMu/q3zKGxNzaWocGF0X12oARNjOa
zWLvhQq+6rggjxoZ54I20Nv22wwcqispx4613MdRRBR6FTiv+pxirJ3vslMF/r6+
nAXKus/WuO2v0GWgVyR+G1yI1HKCXeLUr3EtLg8SPCl6CUjI4aVkNKLv7JAQ+ccr
nZb3WJcWUtLzPXa2s4xvo+zQGLVw2oZC9lgJ+F3nY13H19/zDCR2dsL2dFj8FacL
nSvL6LS2cjJ+HLPFtYw7K+aXmv8vkQDN0o6KeJSF1NJya+/8QrfI0AmnbtqFP6IN
P87HL8luss2NQcFT1R7fSte7OPqZFWp4UHfAqJqq/pb2CDA8LSyWwuf+0T9BP6wV
VncmVzp11At0FKrldJHaXEqP0nV0mP4R069bJIafgp0acMTsXBNsWLjl27RHLmbc
7Qa5rJkCNxOyQp9HY8BUnRT9JOKeahnlosK4ZgLHB+epU+o40u4Zz7Uv7/Nq1LZn
w6PP2EtR+IjYGB6/6cSLgzhB8GGAXNSO+Y9p6Hwp8goGeE9uNS3CQhGOaXHiT2JJ
zBfONk1BmAcMh3fPklqzGpRuWMVy3OhdEB9MZURC/SzEREUNVxHzdoOfr8Z0qmwg
YMdpO7TtWS/nFupP0z/6L2iEM0QlL/dYyHFU9iEw1Z9W8DfJKsIAKWFl4HRHI39Q
RUQ88uqRhD662tH83MohE/qJ3r5z8woyBOyJRn0B5P4hjPdl/A18oJI9WrLx8Tr9
psJuhjVAiFcX0WazpLE7JWLoxyVNmFc6VvpTt6E387wD1MtwN9K6iaIS5xp6PCP9
JyrY2I6F7WavYHo5ICiXpZ7r4mPb3necJpndOVQhUy6u0Z8aujLsSVcab6mJE6su
Em/S1twosB2Fe2belbFwWSERRerijMlNlb/KVZCRqbUWVHwga8cSOelJlDOJ+UJg
UdjnAtRDLTsOOcCfDXYC9mXutYRDl/S1pZEZGvUs2JuZXaFkd3q0d+7OrYfcW2Pi
BuBuuG3+G/+jqlvsCh/NZIozFMd20GQb4RaNT9fhTNZJi8Ya5LnrWagLcOFDgBEy
V0krHCPWNDYip4QXVJv8zb7BPs0hmzOuxpAsz48khX+lqc2x8d+HD4BRjyjRYK1t
mQ1Q0NqpccZ4riO8T2i2BS4H787n13ARpTnLbOS3UouepakWO9tnnY1/H+f3xNNI
V2aTSVkE8c86JaZ7fmk58PEqJYtA+OEnI201Ig2A3Ei9g9QqdrvO775qZA/qCaLS
GUh+TiBglONOtXUqa13o6nz0d2j8jeduaF2A/sZ4g5JwT13PbBFMQKq0ymrdSMfy
5QhtNhYUplPxotpilz6gvEYQK6IBmUtiVPYoqzcIBJHKhlN22N5UTKgjc3Q2ARd5
YngLIW3KSggVKix5mJriApJHW/H4LLcBFT/dxV4HRoCVrFENXiA+WNC7BMMAFHgV
J4LkTzqRLw94X7gZgKK+5hxUWKenuA/6IeOMdE0Szr5IkxnOG9FrEGkXLdhZhx50
PzyHaHfZ9RKIB+9ntryZtJAWjdwRvDv3BjxVvJF1EFip5sDePRWzWSZinbEWrioa
IZ1V4RJi0o9NxrzypTL/Tw7G1KcEIUXAA+an4tLCjYFgTrag6eBc4XEFf2/0++Wp
Tj9knb+MquL4wmeJXmMldI2evFlM5HD17wLePy7ekV9yI8LgM0dzXQw9DNh4QwJp
dV7WADRNi7xZog1mk8/Dejf2CMjfrF0CocWhi/e4EEZejmu0oxH3xWEFmWPEwM4E
yv507HBv4zfaAvSyDFgXaxynplD1jbAp30nEve2o+gjGwbKCJ+sBwPWSoz+ED2MH
S4nBks1n0wvTCuqY6Lne0FFpY3m2rSPL55P513c5bVXyr0PdOtEON19tTis2Za/i
C9bHSITeDjblB2+g1kkqzVCvsSkundpSGaknrtiv1cX4Iy6vpS1Zco8WYt7frZxE
7l2J3xmeQ+rFZ7EBT0MDmbtuHkW6gXw9hut49YysMX5CkWwdSuRl0PHqgRVT2l5O
mSteqM4UQri5aP9R85/dmFeo7LtdoR+43YSIb04qWZ8iVj1cSbQSFxXgNNnLCUD2
Y2KivSOGetquGB0wU8TTkS/xRebQXDUpng6H7DJ8tvqfDAcuKqkOJ1dIMWG6KOXA
3Yz7dGY83qeZAaQy1Vg2YmoQ2wMPmHmYg5lQgLdQvtx4JnwqmEX5kALw6M1b5MiS
2gidezh8JX2dPm9qyWerJzzv4kCkvjwN2ur3GxjOPp1PdQhP06I4WEIU5ETQfE0r
AuARAzV4P+3Dt80gM9Cqkz5oOAhB/k4qPnDsrUsr6alvxYGZuEXUqBS/QUwPxf2H
JhCW06E7U2VlfNQGLQNqxMFTY8QeZ2mb+5+e6iFATl1UqtJNKcI3J/z/6BYCr723
HL37wZA/4LI0mZTVMZQaGipJTLelMaUBfDesERoQWfdZNgrh1I0RYlz44YXwkv6l
pwc+6feFWNM9JSVYikaXcpehtZmmZNj+QiWKAK48uShgjWod+/7TvY/RGZ6fH+lg
iG1eLyYe0PbdZFTrfpzqfhXwUC7plsvuP18v1I/KnvNqBmvzafeZrcr9HxvGq3sJ
Wtu+MLXoxbvpNe4vqMEtelOvd9oJv/wm5wepOOhdj/n3OEv+ATBkGkTa8snWpa9Z
xopd+WNGLPsFAIglNBAYY4kp6lYCK3Sui9kRqnuUKLNAP+IRss3f6SLA4Uxo+6xC
Wh8ZxKldD4wTbq/BRwpoYMlItKPCWKXbCywnbVq7j7W99gdj0fMiie3gZjREVAPw
U2XCq/jzJP6+IK88zLP6DuOdt/e4VfL/By0aoY605apvIp6cBWnlDvqh1AtmUitC
6EjmH0nWFtZ/uG0DQRtdqhe1Ud4qmql+I0RIYyqmbKV2pACt6vmstsb3eMcBOLc+
1cVnD+evbSjqGURFyXpNvc+L6BHVTlI5jpZYw1VfVPhxhStj9UPOrO3pJntVXF8J
FSjVJRG/HBauQIlg/j/mkxJZG4Ax8JBPV0pfrAaMvSHsE/5NBMxzzprz5xHLaQP5
7KT9QXwFV1erijgOK69TeNIMnRZAS1OAG3DLlfJslHpW+rzj4fGWWmBs+sgOifrH
WWVuzbVDmQmRQS0ZuPKltUqozm+OfzGmvyCI3gCeXO3WI7AJ8H6xrF5yDvJ1LvMf
kOmzW7Yazbzs2Nq+/ICG90jLmLOPEFCxAsD0lcg5BacB+ZPK80KKn5TaR0/5bTwJ
pYetSEH4+MpLuEFTGdtILcmgxGAZrhxQUaDLChYZbogZCd+xj0+OHX6CLKCPzvoM
ynk+nYpn7W/t9tSLFLjZs9ssLj99i1qFQyfnYWwk28CiIN4QZwmZDcO5+rG2midc
D//B2lMPO49/0KoLxphTXByKm8V5vTS8Tc466IUQZ6rLjR8aSUe/kEwf8wIRtrpq
7Z1xZBUKB0FMKYyKhauOKy8VwH/7gLdf5FkVMM69VX30xUD7qEmYKZq5zxF0Gk1R
TDK6EjMjW/F4hcz+3XbFANhfKG+wPRkNAatrZ6gzrvGJcLPe5rYtq0//x/TWPzvX
YrI5R+yic8LvUzCGVS6iHar/+yFhEYfNuIWF7xvqkiuzh8B0QUfh2b5mkbUbhWj+
1RTsJekIia7VE3foxm2DfMAqgf3Qh7+1OQ4hQ3TUycbtnnoYdUgkObfPibKACjQA
oSnDOHmHOAhszVnNVbUXbZQnb0bJxVTArLonks66YahaDmwjWFU7VU5g/tw4cizb
DRem9p/KTycsApBz32x/WJ0qzI8K2w36ikO6DSai+/rZacJGis6mrulr58RFOj5g
yX5lBDI3wItRkDjf10R+3+3SKTA2wawPNCPPmyB4vbBtL50P0Ds1HrXUsz7cq4hZ
6eiA5KyP64yqlaOiUWY/P9A9jQPpzmsU6iGe8/ygvPk0BuTmoSNuzUvbZrw2exIR
aRDONH4AfQj7cxxDVmKcEAZ0K3/FZXbubc88V/Bj2utkujUpNsbFJFq/wFD47sy5
TXBlAIoNarQPymNKB4UcDn/GfXkWRpHhMwRXaLkv5PibYWTZ4K+90mVYzLp35mG5
I1s08HHPMgLgNzouL9aw/YM3s9jM+WPyzxcjWLj4BNTRlnwA1LCT5HxFw87n7Vgh
oD5esdQnN36IdwlirdhEq5QYPiKfve3ZNFvxkJAdtYLg8eeh9rG66jqBwzlhISw7
1ha8+yHv58XPd84YoQDxCHb9I4OFZPYaedKfqPXg0dsYmhHXFQ/KxT58WEZ/HmMc
7LeY2S9bej0BzIL5q0HviY6X3FpjQGyfB0HR/v4yPcdsK3ooby+ApO55vJgxyCAo
BZRE0afhsDLR9wKcged6cuInJsoREq8DeFZYducFOQN8bMFXnxku9Zqk0Q6Yphv0
dYMziVH3OSq4XUv3mova3bimuqvp9e99PumJJ/XRq2v2Ye5quUaxyBCMgPWp52sN
/t67qspRFqcecZvSrUrAdnudnq5s0Fd4iTi8w1l8MB6ewAN/MlrBGi24fMKphke8
BbnB6aoefhxR3yzPFZAVJ4OcyIyx0OF4RJNzXmt8Runh8JG4z56FaYmly8XyrnWN
YNRqPDtw/8+3MtgcXd3omShk+Jkodvr5LQwxzeS5wUS/Zeq8kO0nvrqE8JA399Ml
hEFnSsnSCpcptjiIpLmZyHSCDqh5Rk7s8EVYIZ289ueKKO6tguK3vsUJCA+9Ljnk
oHnVoIS5CPf9NR5F4mUPEG2Vs1dPWoC0Xe5hOp1c62Tu7Vg7aFKBSzQrKlWuckmR
XdlkFRGOhJSgPNKKpO7a4kYf3vDtPKLp2TxaZNiV+bOK2uEYdqMmxsqNhd3EYWuB
VbwpdfzYW9jc4l5sxY1VQksVzitCLxE76/SB735ByiqyyZVHlJyOdYEnoJ4toVpa
98TI8G5os1KGVUmngL4eXKmOwZqLTE2kEAZElYC2YmeoFT8D7KGLhz1ivYkyGc6p
3tgpBPrWnymPjgvquzCYkBICU5jIfRfuWMX40tBHI6UmLyrmRwRVRTEK+tIOGGc/
dd5WwcG2HZDAZZncYwVqW+Nz4UrseAWoSd/2b6ZBYo0cZXzdzefHfVhym+R28ZeC
x1KpE5wcIPBynZYcolAi0gd4IzTPOZ2inbxioSWlJ8HNTXqanNEgeNhsbBioaE/5
Y1/o8QKNQ/GxAb8fyclbRcqSyCtQ2J2lqVmoSSGp8+ojw/OesTRku+BqRYEwiq4U
G9Lork5yN2MwBh19g8pYSdtDqStkrbWazfie5r8tW2CKk+3/zfYcFr9Hb8U9l6Eb
6ZBVSCvBCtgKoGwg5Z5afUZQLyaphXHEef8idgxtbfGsL81eSXDU3udoFV5rErUV
X/EYaSmAYBZ1vpE+HUYnx98v4S9LFnuB90lt/vTp3Tr/1jTnD7EiIrQcv+aF1aOA
mbLh3PeyBq0ww8mbSqSxPgM49inu4qcI/vRIFoJdr+nuocShYykyxKTJjmDasy4m
XfviuPNYLAbjoC2Cy2+P+E4Hpsm3XJNDTUyVnEWBJ3ZLmpr7TNkeBFmVUogmUfJr
6LSEbYTNFpsA+w47+QpxGU08Hb/FfA/mlugliPTyo04aRGEsHG/8RKfKnbUqgJgH
guQbd/7tOmIWFymW3n0nrJigZsLlTlpxKV1HItR6Tru8S66Bqs/jjko2GhDbnvAi
0O5RcKOqosIT7iADiTFy2vIRlq0CgJuvnWFwBu7aZ+DiCg0KliOYuHVylt3I1UXa
bd+kc0379diuLVKFpQzLWmxTRBOFW8v5QW5Pe2eIjhR8uk/WsNOFMxVim+MMYu6V
RhPjRUtRhr7LuVbye3mWDr/Xn6nO3C2OSsAuNr2eP8tXs+BxzqD45cSS8YLSEvlP
DB1BrazOv1NH/o5faD7jw12cfoYTgF/pg2U1DO0M3sWPm8JecxfAXCb52x6oevzZ
5sYnvgL2VuxWqfpYJ+wH4BzA6hWhtbPMi5Ce13r1ZP3vUGCMSt6CSRXxAamVCSuL
f9Eq4JtwXH8hndtylXmJ66OwGwgw9qAd+u8E5wtr4ZzhL2cU5gCFMRzX5EAw9x0e
9Wv+jpqXjc8uIAyhVBYg0hP048gTNqmPHikBKYUBzW3Fb6S0zJprra6h8QA03onz
jDirxi90tUImUJbgHC4WPlbN/CthGaMlJEUCKMAqM4E3N/tcrG+Y9W13+cr8VufP
Z2JYCMP3wFm4Z7AFe/QATWI0NmTHQDS3uFzuyj5RyqTn8lHztxRx+oYPlfYKMkWn
VWait/+mUissgGMCN707sbh+FuRxydKxx9jah2OFTqofmd0uR/c+6gq1ZWoXZwa+
J3HkrAl+u+9EmFaXgtjPtQGvRLJNRa5ZjmqjVVq2xUB7D6FMsr4H2ltPOJ4wlLO6
Y9fUZ7UP0ppuaTl6XxqP/H+DS92Q93MhaNqcf0vEoeAobBJmjX0ZVI7EH+Z7RI9g
reZk9upOlR/yOKG5zm3TRpquIUXsn9MCegF327P08uU9u7wFN9N93XuFgKnq94hc
zpIiKKrLm3/WIQVoglsgeXHneNyxh0zoJcUYNS4m8Isz6Ww3v9K5IC5Hieha6tZ0
X82L1zBxYP/EdJL9ufLp9dS2Xn+zHjNDyHvbrWDup7D5WM7OMzOtw3OY6Jwl1g6g
ydZSrSy7Faf7WrgqVyimZHB3M81sioCCN+AvvF4NJdNrasM6cLox3S5b21K0K/oJ
k1vZxpfdUgYL50+HBUwciDewOca2+JomRMOWXSuvq5dXWiiUZMFges8gXXa47OmF
M8oO+GyHmOZlLyz2eZRYXXHp5mY236YqL0QHQoj4IurgCeicjHQoL054L/kOeyxK
gvWITzGZVKyfGo3wMcxT5YIIvdJH5KrurOI/0V7eSSamXb0r8ex7MtUiekXzmNd/
bw0teNWBGA7lv5fFCz/9LQ+phEl1CFTmOKl1qSW/p2sGrkDt8fQSC7+TsdW8PvyE
6JYbyEVkQlEAoNhMnfcMD9OqnO2MZVbMU/Opjd0/zS3T0yz6nXW1wOZr2SK/a0V6
ECvV2qiQrO0M3oUEGOBsDHSizT5R9LpKHcFVGW5w54rq8yAHiMdOc8rNTWISZfev
efpEGdgTd3NVWT1dNUvQQ+xWp93kRC/ilNqbqX8RTAVZTzFeEnhp3sbUrY79XrNu
88CdEth4ysldlRB401jlke03tNTwawh2xKJktlZ/lcU1oR0tE+sXukOYI97goVnI
/uW1tgEh9/aBHwYscRnbtykF5UYimH1U6VlkK9lfEOx+faFE2uwueaHq9r52MBpK
gfuiSk2zJzsREMbXaqR+nk/KJGuVTkVOZMD7JEVy/W8lT6ztcf/zokOo3sVbehP5
e3JwXcD31dujJhF5RRdiqEPVekBrcqdZ1aY7w+PgHXwomG2cxIJLbGUeKRQ2uiJ2
cnZwHo+Vk+pLdj2aISaRQG7ejcaTu3aurLThNk00+YcPaVzdQx9KKwgFSo/z5StQ
P6VmoVkn5ghufMQ+Y4NF9uqNaqGS7xYEvbiYErU8wuHOMd37S9vHk7tHqovKd4W8
FNgFtYR18wzr9Z4HmfevlSmWg8TkiEmB3KwwXbWOD/Q+bJ/pm1KQIYE9kIa+egGk
JBMGShCaAaIeBKCSjwPAGKYLRhrjcSCjfonPTeAauFwG2PrEZMGIrIuAW64dLE5t
bTMBp1R9i7zwrpobDgL43RfwpStto0m7QwtDfL5t/n6c0zGLP4XPr/YUMLbHaO+j
f9EjoV56rawOBYOvl20cE8FhR/WsxSQPcaGGPSHdGqRimb6z7IDT+yM0jap/+QT1
kp7gDtbveRCFQNwPYjoQ1qzCn07oCknKuU+sPL1xzISBM40WMnxHMZqs+zM9EvlD
XKkqBw7fEpih074WRgFjpJ/Ssd+NYq5KBaiBI0I1Di6VOrhy4J8aglahUHfwp5o9
dGeSTae2wvnZR1gW+By4mmrtJ9M8dpiMXutAPY3m6oxoltG4jqMX5BcadoJZCxJJ
RtgcAZjKgFNsQ4uiJeuEmTQppEtHKYSST07XThKJdSSEbPSZIz66LsM3/yBOuS9C
//vIkFl6p/s+YJcbfwhpUVUeYggEEHgpsnnxKwndj8loEp1yUcNTl7cMhF0UeRB0
LK/I0vg57xzubfr59s4oIK2FvtgWt0ZpI5RRqJCSGxpl2XPhhj9l/AvkoQiSsvmv
ThsyiqUxAYkxIvP3KCYH0m2qmdTBWgSTqViH5tk2Tt/BBVLIEnJzJiAG2GvfFb1J
77mwksHd0LbIcoFTKyxRx89vJrHExCl9w/t/NuPDZluyW0civQbuziP7B925dj61
E++SIDkyZd8Rs8ZrBKfQfDVn+RF4r47D5ZODxQpQoSJoVy1f29722BovToGdR1TR
FwXsOur7iwpDl4UKj9xly9rUKBv7BR3ZPNg6ruM/yXpPMJ8xkvpS9NLZt/gtATkA
KdyDf853ZFmxrguLuflQK5xyp/TIPCmQp9NZAHt+Hn0y8cV/jkys5/gk6eU3T2kw
oYwGPeXUJp2qdLPyzBOE3t2UmMTgFzxFS/okR3J8CtlFibk2G95PJqFlOgR8pJtX
mc41El+uQuYLhP6j1fZdnntXGRarcVhaf6rifu3q7Fb7gJHKFKJh12GIF+CV5Pr8
YqrupA6W6kSIPJRt6Df2JL2TDDnz441P7raoZ2KdbRqcTuVWC0EG5PPtcGs+ZtXh
0gpKyvDta1xIquPEMKzMg5O+NxTSNAaPtZC/ZjkvL1IWLzk/kdgUBeZeanafOP9X
7fBlozx9b+irKNgJyEh816pOvouvVITJvWGq4+mImCqT3V6djj3UrDS7dytdv8af
E1AC3MiV+iPMh2gCbAS/g4xf6C9SQhqTnYsCzRRLIorl6teQLA4NgstTxrUy5nKC
kLBtQA0rZDMbx+mLCTKYbKdUHD0jjFzFFEL6LCtUfh6EOAewWgutEZuRgpGhCoN7
rZcWZVlMgq8iSvrQNuDtbJIA3xJfy2CwJhWjPFDkCMelibsJTvBYJ91kYViqvaQI
ytqYgh0yPN37x3FgGS4F/N8cUmGWNbofjpaGh3CkTwp7dEK5T03FoeMqynMn4yWG
HL7+LBF3q7M/Qqnt4zvCIRtxf1q0EVruATpzo7ho5RYxAAEX+BEOVrlC6MwFUVtX
9Xr7YV+tQg5d8VhnaDd3Snu8gknrSF5YbtHkpEcXn8wvff9FOM9EmLB7Kpb0cvo4
49XBMu8L1zkUwEx3PRzIDhn/I3mz+Nah8a2hLFmFQY0Kb6ZnOI/EughNXwGBKkFh
hsYFqQtiWHuKPH/WA7vqQ4ZqrTr2PiFdlFX3TgYPn7CXqw2ZILk1YUHrKXbGH7CD
yUh0bZJzKlGTNO6D/BpEAG00iRBt8tyCDGB2YTuM4u1SEbEs/EiT7f+hMFC9q5D7
xls7DxMONAwyH4VwvV8d5qySfnM+1Ci5HS4ivMHt7dRd13mWuzyoSzCLOQ/xSOig
PRPLfn4BSMu6SQwzeTEolssvhGYZf55YU94NGYLTcVznc0EB+HG+Zzgpig8WoMHm
byge3hfMWXrxxmdsey3UVpQWbkZQ9ThgLXhhMwJ8jnM4Bhy88RXj3LWVT2zLp0p5
NWxp9ph4BsRYKRAUSwfjp42KIgUYMN5SEDJxYLJCM724aslb9uC3Vh+TiFy2S8cD
3sYbfkQvyyviIYlNF8hPeEPf1GZUJraxIJvvylQkF8SpWInSEmOqKrbocyH9fhcm
ojLODj62veoBQIYjwp8WOzk/0TkuVQqnaaAMywPppLAK1H5ZPG431CmuiSdSlY/W
r4UjOXEKmVzjOcOdo07ah+IJdMLvB9Kx7RefN6OtB08ghZaFPXPq0wS1OgZIGVsn
nary6rshne9SylSlCuDZRWDJPzVPKkbRogfk/vtkw8PhiqeoAKm0fP2PckmMDxWi
myXnpEYHYsPeNACuf22A/jCErEqw7D0TxuT/jE2cJgvHjzYSCzdJ4i38sYrU97QZ
HA3APY0FALaYLZ7+lqekAz/5zMyZwJPuflUAzqJ5FBSrlf51GILVRJDrLfP86pgS
n1beqrIZ7r7FdYTAi7FybF2xRMiuGshwsbF5RWoEfvhZFZif+ciGap7oGz50y0Ji
Vs71I8bGy7+8xDNStH4b+tBElpiYT8vvs6tIJzouVqCOfgwlnMcycguRUkHFKUP5
Xq3GSMl6dpL+EqLUTGQn9OblQlhuHcqfrTUBlikm/mAntpUhHYGiUtAmuJDlKbAu
ViFfDU2uc3VVsjOVP24G+09aYEROiCacONcyEC0Pa+B3MRobwdiw//rFs9mura4m
tSf1FvTGviYXN4Ek7mi0Y+1j2Cgqy73wH/pdP4XNUBWfAIO1KyAHEgmWk9EgAVRg
+uZsR7Sz9zo7G8zEZef9TF7LOB65wGnwQZTj3UvzV/aDsUtTgAuni012I1Sj7Fvd
/P0w2RkSS+Tc7sIl/qeY9jxUxZc0W5mViwmi+jLkayLcuYY2DAeyzo9N9xNG9iQ7
iMGWerxdiIW+KBH6Uwywe1eVqEcq0o1MorIjKJYT8HBdDzSZQDfmsrvt3/Hkqr/r
kaWEg6t/TTcIqMUfag8HS+3p2GInks6zoL7IBeSS5U2+dzxHnXio6HmkyDQsR+F4
V9aYByWy86/1MsAWNmVUxIw8NQdaWEZh8jMlUqx5XoxFbHWvcNewMMGu52XDdtM0
sn0BTLHLDXMajlKDvRQ25j49rd/eZtfffRx3RcSf0KelK1EpFdo4Ommre7ycCKZk
JXHNlHR3Y5oR9d/VrEpjLi/Vmdsz+KvOrRtbSh95sILQdmfaqm2H8qdxEO25yO4u
YsL1XBlGmhYxg3qh4ipArwtk870xoVwiHoYudZp6O6BusT5W3tCGUZjTpSxkcd3y
tLOM6U2HBEOXlxzhRpQyxw+w/RFDyHAHLoM+9Pbae9J5t44XSs1LTfO3VJ1RPYxI
qvtf7SHrARyQdADPxVwdzMi2sDEGLJrlT2JGBy6OOBlZy7D13b5w7dOKfziGl1nW
pNm6nSOPiHdpf+aSkq6+o+2j2wB24zR4F3GZ9B45hLbLSgSYfVx+CMgz0wrhp6YS
lx8Enhitx+Feqliy73ARYCivKJXseIzhW5n5/3IQUvT3bTcaOReHUnFPLW4DsG46
xFUh7dfEN1c3En5SXFef6dEZ5zzFmbW63AZ4TAtuJ8JZ2SoLoNDlZ44FFIQTRvv5
H7vWE/0hzjZZwl7W+t1dHLPnL6LtR8txBm7wf5zSkq3ECYwSJrYxssEdoqs27MKw
jl8XI0DIgGf1DFt6uTfSceGZl3E1xwqZkX+FSBfxR4DLdGUapxFg/jRhrptH51al
ew2TC8rZvHbo71vLRHbpuZLNnUkf7CyVmHgcbV07+AFAQvXqpGYwzuh346OvWVoL
ACrW87e62BHrq+L0a6rxnvNwWCs8Ii861hjvEsLhgRCixl9cCfOxhAGJqG25Yaeh
6J4WtA97DNDD2uV9h/jwvjk9lhyhPOV4+xxCqDDDoHOY6+qxfzlNVfJXBwTwqYBi
vEwc7FkoCac8L4GXPQf/mzb9Zw77HtuFUVOwPXJEvHfMYHaaeA6p2FTsCb06I986
NXlfXRHNwNu6bs8QQmkJwsngwl5cAObi3asJWTIxxnS0RIp0cu34fuf5WFqA5JUJ
x3uIOoY8GhBbnmLOYyMWG1ypOolqwtpvQEPmcCH2dJH5ZGx7iiQMCFOeXpRGeSTm
teqg/ja0bF4TFbx+/Nmq8DwmUJGTyE3G74+AQOK+pyX8oIfE1+0Dq9l4uxgK+WyH
5W9ePY0YBkdVRtthP4KN81kkk697NBPZpoMuxv5qIVsBQ/2O+9kfv5p1wFPlKaKX
ZEWl6rn8Us2esUSg3HvZI8o2LC7cjOFBvJH6DZcMNaVonS3ZG9LryOq8+fxCj4Vc
1mu3aE7vyW1sDjNCz9xwNFadiLi3+OWvsH5ROiLHOfM19yPqvVzhSd2BOIY1htcd
5hLeyectLPxDs5FsiYaU/QCCXDzXqfpi8BPmEZg+/I3oV1uiW6hnftfvwAUAtrLQ
8XsC/Kd7+KbTa/7ugPmRQ0xCxF+M20HGMuUoqVd6GglH0csT7ix+2kmFV4pfKFe2
NCPlxeg8qYRtuyYeBbEe1wfgKHaQ6z2ZL8KA3AKCsLs5rlgIew5fdOrP3S0ofdU8
0mRcQszjEmqqtJh/4WLwRLjHRZfQyhrN5VNh6bsfzE4H5XPbavy8+wcbQqLPDJw/
Tt2SufFVJV/ZW89XQgGX0KawcTzUerNlShK+y4ITo5qZcOLgsL4vnzilLy/Huhr7
T/Yt+LZ3oV5p2cNzWV1nVheb0rCNM0c5IYiXTJqNbJTa1IjPw8zUq/zycRhFgDSA
+5h29fHXu6ek0MSWjNcA0HdSONkOiY2aotGi5glQA1anblPAk3v8owt7dtM5gEMs
n9CM7ZX8Kfy7PSu436KSeoea90fE9z/cMfB9oniR4AnHRKmkN/J9od9KZcuR1dNx
jZcX/WqLq+NwJtkERgQ+ewrjyBuN7s3aKpV4GFmGxLoiHA6whc7DCWXVV1tNC3tq
QOVgnaXvIz+m+vfmOMJyyOqYfJr7QLqjnlY4ceteN692dPLnxEajQLN9mxVOf0yg
Pyr7uBruvJb2SllAFazenOZCwqCG5DP5vtXUP9SkeHQf0zbmmKJkOchDAWAoTTya
u+FxYJfshahTo4k415P1vdYjQD2zkZtRqxLzWblIlP79TeqdPeb2kTL2rdD0sm2m
hwdtU42EK0IwneZFRhQM9EmVNNLifRhA8PAE3+ULvq81pSARUbLIUd7UJ9JohcF5
kTEyi4VS//36wQ6YZBc8B6DUNMGq8EbjaK1phtySQ8DB2PPg4W71YQrU2NMa8Q+6
uN+qnpDNSei4GoPFi4mfhdrSuab14D80ZDzwJckyfs+Gw1drM0y5gOP2RzMes+St
W22iHkbJpAWzupHuifEzliUfO3IO9RXv8W86T1DGIkFqObDxFB25kC1O9+Vpov1l
G7vXuq4yDsU7gOKnQcv7djTwxw+OaB6sS9r2mn+2pccLnGv5CLbog9oWO9x0qMMJ
UBJBuGPsHyAF2XJflWd89lgjg3FSTea4bIT5SJbdfU9MXMnU1ASMNsJhCd0P9a8Q
2tYSFwCaMV/6eMHOFOmWiRouu0Pust+PrfZWMVr0CxEDcd40TcZDjE9hMdhvM4yD
uiO3X3jWMmbbJzXpqWFMEHRcDhDuZZcQHnZ1RNyhXGJpvAAX+v9WU87Uhy6cMHaH
qL8Hr2RQhIpEvPSfrs/W0vS9YDXrEOb/xNO+kP+i9LAWBf1eYbbM544/VyHYQGtT
TQwtbHME1A9lB/xSBzLgN+YoVWTdfeBbtcZDsAQAk5J6CZGQ2z80I77D75RmZcQ2
8dy74fxho+jKACec+Awis1SjA7dGjdSX7sJPsLK2ddpfEUa8fvHlLbkudVh/MsQj
ZivPhObsPCaQVZ64oR3BJ/3D9CVle0hjmnE1e3oiaMmSF2uvLo+x5MR11zmsoG+K
LkcdG5v/e1f673vj2xMsvc2j3HQvtqLSbLF0h08GFWBe+PKunayaPW2mIn8aIHNl
m/PtLf9exOTZP1VFEnkaZAyyH5vYalGh9nNJIvSmfka7ruAtJ4yzVdRCPpyHyUkq
glHUHvf71dpgRa69mgJdc13o29ahijHUZKnKOrKLjAq1g2prQbcOwJslZ7KtYKzk
wRSnQjhNbgwFDNiMD9Qt+6gcBuwe/u1KfsObKnsVVp0TzPNz0hzIdLKg9HkvLTcl
eHbmH1uKUkcP9/DDqq6gTXO2ozyMTBIbiMXGvaHM/+fWQZeoeiUIBkyhkii4nnNI
coyi9n5g9q3/tVcIyBT8t42XVjgQQk/XR5bkG5jLjzyzdx0WuB1ADf99vlDhbmyR
dIIiq3ywxNROJSZwjb+yr0cVdD7sFr+7+BFDGG+PuZhcMxOgdscqRsaRb7vRTthW
6k3euZ/lxvrOeAHLOc/aG53aJx5kTJwetMpxuSVlEjmKiMMiSpRvjpZ+SoTyxt00
e1PcyJPIs6WdJA2hRHA/+murqPOcXRploGGlMLlMUkmBmrZI/0ynvIEngeoJl2o3
MUTjr37j8PhttKMWOL2fwsyoYFr5CnYbs+JWroKAx59847WXfLQNLHiZq2gnEaUL
rMHZGPYPJb6rn465VqPlYI5HKG+RPjpf9jlGJ3bVIsUm4scCo5iW4vJBzBLiGjxF
kMF3Tzma4R8NSa/lYvpGz8sLqJMvUBObpuMzwTzUnTcWFnt7iTjgxSqSLDLPmbDz
PmkD+7vNN0w9Q0UR1hlChK72BSA3rm22WXWb+1y8twdgxMNuQZxFPuqB6e4GMzHN
lTMBPY776uu8/8FQo453neehnJNymHrTnuCKmFsqwJ8qoj8KyDJL/NrLTUVEayWZ
faZOI4Y3Dm2yj+t8+m3aoGPKxnGVou1njbPSH+d3Ux8YkElkzRT/nmRpCv7Yq0Zc
7LcZoK90EdF45E3UW17HL4zHJ35dhrd/hmGHqe04ZGGD0KfY/NznePI0uNKxQOlN
qcEHNJmUUJQgSqr93od7ebGiPyHv0WeTx6eMnkiDS3rVhVij7+bcH+Y+EbXTrRTg
xX8l3dHmLt2sW1on7hbcdv2wMQEJDrB5CJQT7A+QgbJPIc1Mx4ucaFY99F/pQVgD
ae7IDaotJI3PIKvHQhBp6sC1wEzNLnOb1f611chcYXPzb0owiWZUff9W74jQqFhu
c/AjQG6fzb9OTew+LAthN9sDpCk4u6qMTmqtMxOZ9cBamVPf2HPuAG360v1E2s8E
dsp7/dnvev2NNlaAhNSLQjQf/nGoySDq4h7hWlrgBmhe24HL/wbtjQ8fLCKQ0MOO
ajDXZ+kCtajN2X12kDmegnv3dRMnTdmZUROvD/9qcC9oC3xTnFKZwUGRY3IIHIZn
94hS+tzAc9UVt1ZQ0zqX/dmf/UJO6298xfxbcBLc5+wPOC6I7m+ceGVf7+fdF40Y
hsWYWJhwZdPOgMhyOgutfqQTIQfVo1psaFwTg+mp9APkbh2fL0aENWl7ZnP6bXlB
w9VrVkxh+gHrmdc18UeyaXSb27bl9o7x1c7I74gVQoTQcE6AXGLMB01Sw2sqb1pv
+ZgWsQ6x+AIHa26R0WdjBUA0FuEb+gqhcUOln84TRkBQSYRd+THzpfAMszIQqhaC
hbZlwyGeZFk4h4NBQhEyf0NkNWUm46DG8/sCy/RqkZn5zcWMZuj0ZUCkw18MziDC
kPUU7Z1FsnkvG5JkazJIqs/OLDvUsokuLzbmePo4vnHUdyU+LViSJye6tXUpMH21
kKVbnBXNM4hjpVkd+2Kq8U+hA9SGTXxUTzQBx/IxZhziHP6r4YrLOpfI1UcPWvNg
edjYXKfju8ZCXX9x7hjNo4PE9AK7wvLVFMTY1KVwLWxZ4Ar80H65odphK3tGFGTL
1HOQGzAJ9WTEKhKq+qjJ6OSZ+vimlx/Cq1W6NLBLCBN8edSrCDWASyqY/DSpJdOj
1aeIwofSx2m/CwTtApUJEwUh91jD+OiR6bt+WI06rtP0EkTU/z7SxfjNqUgSttNd
OxoFmWud7UbrSJU3DV7OHOy/Ss1cbAoHeJq3SnwBQ21qp+ZpsMIyIn1Hx606+plt
3h7ywUhOEPVp1SAsCyeUtyY5wULej2LptS+VEFlqRBWvftib4IXy6DiDwogVHJ1H
VM8X5hXxtWojGm+B29Vf5axUFZidPQiawg0GnLk6bu9r8hMo2opl4jzuiOW39KdX
4sS3QGVIg0z+POGeQcK72IS1ZiT1KMdh/8EyW0dk0qcu/CpzMJ9UzVQ5NGKZheEU
xm9+7OCSZJCHSUWKF01s28j+9u8f1IA6QFJturZ2jWGITjUi/Q07QU9r95cAXTFI
vlGAftTNyjmemB4l6MITayVLOOJ9SjlAwFgA5TObtLUde4bzRgklq/6uCcU9qtG/
eQ4ng8PAcAeQtLScU+JyAyAOCN/suzdooGvnhZ564hUe0FnBec92IFZOGb2h0+1O
PuQyZsN8XT8EXxsZK11rYAE4wjXTPcsmv5Ri4zZw7qQ5h7Poj/fAVBA8zcC5s49w
sGHwgNcxNih30CQcVo5r+61kUfmVWKA4BCNCGqjEOwW8PoEjb6ZrrhO9wWuAuwn0
0/SQIrv86/AdQDFLEoRM3p8fccj5mV4ihnxakO9x3GZy5kYNqiDQ0aoB07IZ2kb1
tCUVooToSlOCvlK02ZTEm1zANThoV6sSm213OyTzPhaqDPNuBzCYoVWIj2b/gG6C
ypiYeOQyYVUFHGJf4AbV35i6+r+d2tNxHpcyqXo66+tUy0TRF+rSuLGoFwzzIXiK
I5ipZ4dr3jxgbQHzuvEpKRygJOZYO5f9tOukx+ygWwIeE8WyXN/N5TmRAlDL7CHx
xPAAXG1KAsWhireCZAJ3b+bWqIVaCMvdQJ08u+lqF2JFsJgf6F+OxwGDyCDKOIBs
x7VcBWdBhGRxfrpFZsPNdpfGZUJda/f+X0n4rQhJc5zXTzvhvSvReD8J/BpAH++F
USHMPYORcMKTn/XffXOqNIjN5gC22fkjYnd3wOw7vezNSGBf+uy7BforlrVtI1L+
FYftyx1Tex0dsxOLCHeU77YBoiTRSqMVB3aCyvNwvnFW4lxEBLkcJkygMvLRTNht
Sx5dNESSyd7GUNjEYmKtltmRYjp1s5zxzxZTERE4Bo57YlKs0LwbVo9xqaW38meP
QM0Dd7CLkF8/7je2PJT42/3xrbs3UpZcUk/+kG78PScTP8EVwCqC9+wxU+OQjmBd
p4bS7YL3UwyMnAY0aTSgNmh9UIE/9qqQmmBcY4XxN1L3SvP8WZ48cvG+9Jy+wpen
8DciwIqV4cUIojZXX1DPSF2x2kmJYBl6zMs8ui0xzvj7xiTM83FiXkYuGwzjeUbk
N9nbe6PuxbJOZ8bADWeLmkUwHybwyXONCVWCLosEsJZ/PaIYxVVaYBXbt6upt6Kn
fvCJE96XWQQIPmwTyEZf5qg+88pIU/2kB+nErB0Xd6CvlS9ZMbn+V6ufE/8+TyH+
jpCv/5iFvLVYO0S139NbOaYJmCvEM0scMXz9mYxNnJQ7HXesCnR8iDRWzxUzh8Q3
aaOweQ1qikCybACo4UBoHuPYeHGbGpQm9+kKNB5rO3oigJdSWBLLbo+ANbgr4KsF
71I4fT5b3P9dagO7uJlR5M0Hx+RIUDrh4yCKTj6zT+cjt1arEOq+/WSSiNSmH9JS
gZfYNCgLo3MLoGNIM5/VMaBE6qNz322/NeSxYcJcKrbIBAzh7EdVnH5aImiz7qp/
JWWdUcsBdHtFVdtCzxNiR1oKzfT9BHpthaZTERE7co7nnUtwgRkWWncHaKndGjpR
ytEjhIsUugd9QoOUvzXesa7zU1mEVuoddX/lwDBNG1PuOPv8K3oO04ey/e+rkX7z
Ja3vCdi0nmRktTRLs/HwjUrH1IwFI0d/Xl1b7guF6OnhiHbRakRfnlrmeYbH1TmA
Hu8fad/hZ7wrwX02qszF25G8D5Nc4CQlRxa6ikjYcCRaxsFpL+j7hPhzsxV9vwwD
gLQLwmaavH+snJc4TQSOB5cQIDir67FV5B4DkKzWfN/dmutzt/kmjr/x1O+x4Vem
ckGT4IMrhbuXcZFVXptmtCJ3GDADjwIwzb2iVDyT3xO9EiiEkrgmNs55WRyIHFU0
z4AzlSZkMRMgBMbodH1PgFvLHVxL/ncsqCHvx7iLDHUm9aYmgGsDhPHk30gzL6XU
7RphlO5I7POAv2t//p1+sFt2Z2TYKwLK+QDEiaCs4AiraB6x6PplGJvSLz91WAaF
VYGNJ2wxRtMe7XTdqKpT8zDy05zymI4uMDU9LjrMyGq3c612V8Vp5jQU+1TlyMWI
pxfKuNmsGv/AYkioY+XaDuGSfOTqrgKpo8oU7+qfNvIGC26PtH3RV6f9IJH9MhaB
YZfzTU2MNz/s+otO7Rkb737PIJpQp9zyiXN/FSoPMWoeY/Mg50pcYaCJgkH2eDA4
dimZ78sHnadgVcb7n76Vc8LRpDlFpvld1OrhxYcbJ7U8Zvkgpko8BejBCnX89NDM
hGtnRovOYw8wFfZjW8u2Ok1HbrtXJy61jmOwbXJbSV54LNOpZnKC2j3YwgWvP/Js
xPMP7KQ05VlCUMr94T5L/patdGhtigTQmfNoTdQUqtSkaVEyWBhMT4q22/NfrCTE
dHQux07pJbXM06TtPtYBJxpYGPZWe1OfES3q1odKrexwFxsD0L9GSJRGDxXzCL5p
67KSWCKfHzNYEIasMiIZ/NUqsj1RQBhat+vkCTzf/sLR934QKR92AyFGcb9M6R85
mq+nneu5aa8iEz5pQ3oHY6KCYUaAVU+X4i78UHrdoBP3RjnWeUiAMVBchmyOA4aw
ecKLh0hRv4qD/FBmgeYu/WK7woHGI9owQzPv7rWGjdoQ+OCo4Zi4+vztPewas/PY
QVDiyzY7ArtH+4vOqOSNEkuY1S9iH9j49Ey9t0FFjVQPhOOJpALlD4T1WyX5WwUl
ToAIdR7jF/Xf2oeQ42RjKIRBNdeLDJdkBnoOQJzz0Yoqe33eeZoW1SGJYgQe5aVz
3QU8AkYVJnSQbRI8gaPj91rpCDwIMbvPMRkO4go6OvWnuCpR1/QAdFMpQZUvw8lc
oKbva3Ai7Hyah5MO8NMAUrRQ28QfWpIagcyJ9Zk7XFsmWtH9GzuRz/1MfnCJjXsl
Sz55Zins/K9ctFkHiaqXVv1nkeW+LXHI/sPe6wxVQzv+88jjVusnw0JkzMPtvpCd
qTQ/UsycDmt6N2sSXVAKqTlblwWOyTgbMGL8w8T2h9xe8B/30Kyh7MCpNRrge2vg
PZJ9P4SognEP9NtPe3Wb3nK4spxg7nYefgcOyJmQlysq2LjS8Cyrh3w4w0LtA/gr
IgIdukuL/JzziUqn2dh9Hk2ugI+/pOxo192R78AXpjrJ+ryybtk8KuCXvU4eRKcB
BNgi6HvDRipEJkbHzlc3SYN3dmStTC3rsI2sm3B+F2m8tdykLVI1sol3vW86+YQn
QqafD4I2yBMs3HdXTlUsSn5RJjJPQTH/9UrAj5NvFTtEPtd6+3SwLMsLV+nuElvN
+03hK/bC3agIxSR7i6jtk/y4bez2qjbB78Gob4mK+TrxFVWanov2pBXPh6I7j7kQ
RYIoJHwte7ckbfA3Q0aiW5dS1Z/iqLGSXt3QQg5jkob2C/8kwMtjwGEMRXahNyoo
LiOyqxthaW8x43a8MyWBpU+ZfhDVwOEiMQGo0JBRjXRZfppHyOZHhdbPHltzXuLX
P0SB0E+t18KvK7NWYPujBv5Aika036U2ViT4W5hNtp1X8XAn1WkbVhVMkPDFO29o
Z6K9JzNuKZs1DZWX7/g3cBGkcYTMQ/PIoIupT9o3ai8cuKC5QB4eVW9oDTARzTJz
Ip03U0csQOSvJDX7Q7Fb0jIYTz0hnwco4cSFMtYYekaMewJaUGr8pa5fdaeUxtU/
ebETJG9f1bEldTommVd2+S/aYvckGb37wOTIPMx6YngZao8KMj1OizTnecoxLeaU
PWAgMiN853cZaE+B1RckCS6tuNr/42WP1Ytoj33wBYPm+vU/mF2ShyIaqb3VYemQ
aqA2Bt8VCPl/nLZmM7Pmvdo/ZthrcRKeFhoxFcP/2kUp2QxDvbSXXNYuXZOvwRXB
lVirO48RzIn8+Yr2buKbnD8KaahZPsdnLHi8V/ODdfKYiShNo/Zgjl49mi2aECw4
etl/GFW0zxNK4vwds96lxuSx9KKklSVjYk6VHF26m2tQJz9Dt/24UW4WZfVRuSvD
jsyH1mY/6xM6QzXsqvgcl80QPH57agQmFXmn/8MPWqKAA0oXRw62VzaQwKmnBzla
RKGlffXv412O9/BO6IVpdIaewVMBv5MHtX25TNZQfC4JgpPVQdX8OWwDBefa3/Gn
Kb6L/r0MdGwtD70sOnRSW42ZNQ0Uhmkh082S0ioqlJzWyzYkbNRA3i3kVa0Nj77R
1WIz9+vcQp3iL+OK9l8r1UcVxVzHJYAB4Dq0SSmicSzbVnc0jmcNcW6xd030hB4d
ejwYBb6Hn9HZeK2CfZSib1JcaKMRRNgPhcpmft3bFxIRnqD3ztI8OW9/6LGKnOrB
9c87DKsH6pg7k2ljs/sq6/iBKlDL7LWmrcumyU6e81jmjl5ya+scGgWUqM6FXsEJ
75CGf8qU/t6L1iD9sVVfpqv4GAkgQgKx/B8BDP3Qb0uw2RpnPfej8534iv0knfpx
D6d/xRHP3YpeaeNCaa7BPuCKi93b6qNggsiQg9ZZ9m9/7/wulYBhXEaH0hUgfcTg
mgQOKHLQPpF5nnpv0wnlXO/GJSNbLdnqL5ENHobORGKbEG3z67kjq2Rp8ALHW2JU
w89Loc3cm3zmlVJNpWmymAm0qivcTeYtThYBKue5uf8MNQp8J9VfxIilUGORBcQ1
Yi4ehzVIJUkPStQdp0ZPT0BxHDSoxKlRCjGvEJl1IKWNV+mMe/aeRtxSjyFomXn6
wdT4hghtxAOL06R02jeoSsbFFOs46MEFjVNe375rlZb2K/O1zfzJv/GMRm6cSLYS
VLfN81OJ8W8RLqRtCOAZEHAUrnBAQeuqLdquV/Xeh18lxD+DQU2oGfM6K6P/9He6
S/0y0pn4R1sHYVdkj4CLOyB+VzjgpgPyFAdi/OtplBgPtlaCFg/TMGpxuclSWw5q
3LfR/RQNNnGxrqayGxzQ/DHJcwEzn31khB4jVPEsh/DYkQ/qKlo2thYgVhTghh4Q
hR3U9WJj9ic133YfkGiQxJBVAcWg83PAqjegBsnDDdDjkx4g6fRuFzqeiAOmYLoS
UU0FNRDaGKQNgIG74KLYJjJXqVKaXWFTy56QTOzJjc6NE8el/Q8uZpf+bFrZrAQg
N+ETsbOXGTDppWd8KaLFvkShACsOvdWD1LIXk1lvHoiLN+vKCkwfyvpcv8lwvuW6
Bk6cmc89FeajnJ0ILaL0QuxPyT6LNYxdmK8Un1xMgvkKJ9QHLrNdBuT4YTDsuYZ4
Aq73ODA6PcUyzplfO4m37AEY2jLdqclRmVnecsvd8y63IglOTI7qRZfzz+28k1K4
92Z/ei6PN77VPTnCrOrjWbuloyfD1htNxjw2rDbuNoVXPdBxyHlj/3dLtFYr9yhk
2WbMv5/xviu1ccCV+JvV/8B/g9bUko6SP1sY4bhiGgiIZDdbGOHomy9N2qBstfyT
u8Oe0UpZKc6rrOunGw6f1Yo98KTtzQTFd9J+kFpmAbBPqQCRPrscHBJTl1zNNWPv
DxQGYZmmKK+iH8lbK6k/79M0KkANbg0Ip+B1J8f3sgGlxZjFlPYc/r/mBPW0e+CY
95D7pEChrVxh2YdRAXaxDytjTCzHNSJc1QEGxtII8iwF6anPHa6Gqgkj3bT+s67V
XBVAmiqJFEzL4EuU1oPnf0QB1Ggx+DJVqdqd4iHSTYcKUqh/Bi7XZpw/BRrfMQN5
7OCrHIK3m+IxPeWRX1nTKZoRnJfq0O4ZmtTY+38EG0zeoPKJ3/TgNYu9uR9Kyp/y
27ibySzb1uS123m90X7rXyp1a24MvV8ZnTMvHMClXBau68KKUyMeywPC0cVeqImR
h6YdSN3MfccJHtmaagu8JM3tqdx6tNx24I0UZGJ0akUZccupTA6IJs76z/uZqzCk
81SGVN/Z7DUFxWP7Tnrv8ixrSEQDyP0ocloYz48klerVleEh94vViC2/gZTZPi2n
XfOsKfqu4M27IV6sodSqnLwkPUni8HZtWayQ0aZjz2EXEY724osB8DID6i5Myuoy
4VHo2Qifml427qh1sA4zAGuut6zQQPSaNPndv/1xwryHfojopLrXbKUqo0kH7EOI
NDbaFQ/Mcts7+mpBIi2r5jngH6GM+DeCaGRiCtuIhwm3k3oarLOcW1yR1x53IWvn
YKXE24Ft8dbHhZ8ySAvTFp6sLFbMFCxEBpVOyrtGwz6vSYjCHL0Whe9PM+S9y0Al
ZnVLcnmsbmIn0JJd2fbUNiLAaH2hGM3am1ZBrinPflh5H6vMzw4ugaOr7RQmlTJN
HnfpAN0XxFw/jzwQp0V5RRUsY0lFkxEgGqzT8GSKD9CRtdV+bkm/El/3ywKHqXe7
uZL+sqj2pFu6ywRzc+8Hu92mf8aXDGzwwTZ7xm7pYN/gI0CBgIXE1oee9KzgBdeo
WOA9re9fVdOwr0+DNzCOBc00r/ckKJx0DZ6bg34q4uHXNFBuRfpejfMUDJmpeL8h
VYWf+3Ae/ZAn6YBqKzTp5mNy1LrQRQ+bR8JJY0coAYFd8MOg7/lY6ZRP93NhIrGM
QotMf7SD+LbICUK9l0lMW4RIhP/1xLC6w7sx8fcm66Nvy+652BUcC9XaNTCASoPi
X5voIrYxojVOFBJsD72DRWGfOWRPnWomlvuXgiE+RGVbMj7M0/fhh4DP+AktcC3u
1lG0jj4iionWu/RdAWobw8+aApa5zimgL9boCp3SyxY0zgBScxm7XvGSqYFDff9L
Zd0sSEms0CGT9GpXy+MqQl955RKimqdLjUC4u/Nk0l1U1D10wFY6rTy1b5docsYl
s6IlXEo8w1yU/iQxC/+Ebm3e54QeHCznYHbGSgo9kyISVC9xED0IifyRJpdr4W8+
V8UgblBI4iRIFocfGDMkl1hHXS6CuUU3To7Wfj/D4q91Cv+9e+JWG0xLBvl/gNHO
l744fyBlgq+zJBX546x6Own70gvZezUZ3mKVp9GB8jtqrGjXx+Sxsrh2iE/nmUCw
udze+FBYC8roZvrgCZX5mOhcbSi5LoH04LKM3SNX5uLl9tqYXR13MOf9fQ2Dh8q4
6f06PP+mOX4sYEtts3x6w+bM5Jo/LuhUgarXHkYPfIvVQTUxZhP1EuFJ4TyMy06/
oxZPikILbe8ynMJQECgHxzKCZbS8YX0Rxi7hjzc1w9LzWVhFkCaQZvfoo0YiQzeN
AALb80C1L1i6jOP/8bFeU5kZA3L/hH/efsbzEhh2Re2CT9t2jPglgKTE59SzXd+s
g3qEmwt4Co95wwTiuHbImkdh+KfwPWlLcW9eI/fogib0HH8j9cife18SnBLFfmNL
u54xAqY5WE/pOxTYt2nTbmzeq0vT5KF4W3+tzp975n2G99jxDiLtsJIBQm+/M/cQ
cBLZEMCFTn/72EJeH3tVZ4DE6nI7QUTW/CDiUushLCspyt0tokF6iY4WqqQiBJDQ
qGWFhWUm27ZhbI7yOiN+ZdpQ4JZVbqv5/NDYsVNIFfOsxGTtioSkD0qit0BaFxw7
AjtYdpnHXmpoIqpkOiePj1ukRoJXxXxuI4Mz+YKLFyWWA27mC85meZByZi+2+DR5
KReJwgHz2KNhMbBUpOzxGn/QcrvUqDnxraij5j9N8cbKQ8GzSw2aiYKBCiXHSmb7
C9u4cROUTgZP1c/AyRpq4OlZ48j7UfHmS9avwBADAk8K3pvrXhDklQxuArsh8Dlu
NPBQt6BaFpKKopLcqKSovOKEklfDK2olLtf/WMlt2h+QP1PFlBgSETrHSjpVqx/j
+xg3nGDYe+G/VlilzxuURUT4xI4aUpTPZzPGEZPv3WKwnRmdIA3q9N6XO37VUq59
pj4WDea0Lm5hvwat4eU/x4iZ99IK30XC5nHvG4EqFxQuqHQezPZLeboaYH2gygat
CcfUMEo04MBX0K022635ckzDa+YAw2fZ+vc09GbacdqVqii8JovkbOSOVcyDqOHQ
OXaoIMMi1AvzY+89oi77afRhA0GOb4uBY5VeplZuaJzzhRDNRc0U6YQPDU+NxtFu
WvVBEIuswWVGxyYW0R83gSeeucbpFNI6HOHirJZ+Yn02zfPTSLnDg4iZaD3VvhIg
E4AvblPJBbX3WrbA9024G8fz8RNeFPqflU4Cn/lecvmdL10FWiilDa97LaKSuTEV
ZY3Rg3brimesi6UK0xc/2i6O6rScpYL6BNODjnBOyeLL7LNM58iTMV7JMWCBLu+2
qz4hdlYFuy1V3YNdC0dHc2n3T0N6vSM6w/rUXQNE5PKPoQykZg1Aa4yPA6JurJpU
jJNiivUer48/kXbcVxq14jI4Nljy/UO9bwwr1FDFgX+iVdt8CBi+jqpoAMVLUpM4
/L04MOEtF5JB6TVTx7KyT8lWyi6AetUpQwtjQJRn6v9TgRaZTssAUphkE7A0s9qd
YDtCjgEGlx9pUcaxYL0oW7yGea1w/6kSrNGL+paHQPSPtn5YO566UaRGUd8p1L3j
o4Bg0+ms8O8mR384O34uCvmKzmAqulz5ITTkmmbB5BvQWzND9wlIAT8n39EB1+sW
/vmcSZeYq7bZsfxc0AROFkjdpNV17trkMZmf2ZL4yr0eqsTAGAY0L2bUqGxxa8lp
zSJBO4ivtRTP+B+81rgvInSe3PWkxLQBvH2Xzzz74CD+SZ9emNPR24xmfUYsAuqs
1DT6Phz1tw/o8iFJ04dz3h8iPVi+3g75ORntbD4eG8Ab1HmGu+V8M8H9Sf5m/07n
pDT0wgP+U755IRIZCcPZ33HYonEL8+4wWg9FAktmn18xHL4nZfEk3ZrcuvuDIpWb
n/jO9Ry5MK/JmHOEQhvvTq4CNRStbEbt0XMZUsXLALFjmn4+DJuJ4nuRhaCZh9fe
18boL4GWW6Nw+U69lYfvkjQ+dR7cBI6ynUKt9IYhrCFLVrlw0P0d0BXlpnM1iPvH
tYuFOPU00NvJHH+JLq1UBLBAZUmWka3jxfntdEIvdJT6MqxkxlceFJjOGZ4Hxy8v
ZUn0QvSbeftx098sW5lMzHiVsbln7MdhY5oWxNVl9/UigR+dbQ1K62s46VPelf1l
r029sD/pziPbg5uM1u9MMfxN8Cev8UuOstwrCkL90R83wGbEKOivQ+0CT0JSeI8Q
1iNaTmyyCb/ltXLbdFdMK7tcBeM/+DP5gp7dFCUGu0J8RxmMCpwW4Faeo6sy8LTT
sZPLoxOCAvh1pzbGYeC6OXW22HeRdeE3V5Pu3OcrH8S60XVK9h6C/LlAFhS98nu0
mPy3fn045ImSr5ZoVLY+X9MK7S14WE3XekMjONWo7d1r5GCftwzVVirQpgsyIv7Q
VraZoUkmu68guO0GknlflHpyj0PW9M2VaZzbltpU0FauWAjF+7ELOEXQkFwzVdVa
Yg5zgXgH1dT04AyU5tKt+uIetkemIsL8vXIk/c6js5I0YZBAeqxEeC3qJZWdDGLJ
stLBnnDcpg/e7sWfqDd1lMtVGtYgfWZsDv+vo7edJfYodG4GMZ3cakquzNz1017U
M3hjB/8nlwDXIgU77wHkApDKYN7ZOMpN7lknH9/L8OzMDTabiF/RNDVqPjE+Q0fg
qJ6wQtC2DYgfSI23qrOAZyXt4D+QsHpFBIuR8z5O7YzhHznhyYAhL6ntHxqspAhO
0MlQKFcq1CMj8RzWVlK1gaoKHSY9Of76Z9D8qzY/fXOHUZpFUOxLCtkjJaKcOJAX
w536FOcVypx1Z8GW824XSGc1yqKOfmrjVW2vV0TQfIwwxGhygo1e0s7DETbyrxI7
+85nuYQ7vK61XbttwFZ+7TqtgbK4oc4lQsch65L6ztfh64FUwR6Tz9VNsmdvaj7W
FfN1PjmP+mfmvnAAM8Ao4l48jfDzfHMsJlHtbMO5GLRZr/R5AKMXWGKMvp29y2/L
Dsblk1jb8/kI6eWmaxkDyQK9Zxdp2jOarfr5tlf3TXI4eJlAesSfxIlwwuNfuTbM
XDafS7JVNUz49bEUxwcPWYYoe2iMd5nRuCqTdO5F9pnvkwOPhSdPCQAOMGsnlTML
uBLK1NQBz0wa9wQKD8UwUJM/Z6xaMhxAXbVDK7hETySZ07daVpCBCOK5rm3gKlsh
LJoAgVA94mF+LPaiwTFhB3UogE61Kg2pDvvtmqq43Hlfu3aXxgpgdKKwLlCmxATQ
gpRaliP7Y05WRMD3ZvzjdgxyCH+Yaah2I4AvbD0Q2pN939S3+YUGwqfHaLDrHvvE
6fHmq7l0gic7uC4mdT9OGMX1dKri/p1/FmUYdDwZc7qU8j1aXaX2VtbNF+1WdtyJ
nuatqScflXia+ciIuiWWUi/X8/4GFDndU5Op/mZQf1DGizpTbecrFEuH+B3HfU3T
lRFIZI1mHi0gYiK5wF0VWMs9neyAPRfEPi/S3QsJGbm0rROa8NW+9xNd3BYdfcfQ
3eLqLDxNAsCzhTSZ3U/MzSw5rEiggSKsSKRus1Sa20zZ7g26h1u8EOy7lf5MZ/w5
Iu2Shsxs+0rCl1xEBIPnfyPg4nuiNLmRQKd0+ku19GWvFkPd4L7awq5LeyirFI4z
mO+BuC1kfG0oItyk/gp61/yQYNlxIOiQpynNlpCD7IF0ZJqa/GNSkXVOoJTVuyTb
fMEJcnSd8yhIjAAfQHXP4PAcG3gvLUeK1+KwL/7nxk2J+NTTrFnYSk/a23B75JI4
YSXFL9giaQIzkD9q7Gj+I3g1tcteJRfy23E/7q74mrvl0FLm9eMCFOxpu1KjZy4t
cQuoGeqiTWxI9l/k8RkLZBQyD7LEeeOFcH78HeZGDtkN9SBrKXbDL7rQI1zaST58
cbG2lGstRNPKX7ko+Ms76vTD5tt1IXOrQKANivYPaDrSciMPowyZhdUFhfvz1eHU
BnnFeOzeJlYD1Uwz+UwTWY1kLnyD16sJj8Rh1V8fLlmDyXzrOUg2FYRgkgD0vB3V
zhlvua+UsOYEwgW6gotkYcKXQR62fSlJ5vq4161rmwDbsI2AxHy/EbpsQ5DAi9S4
JxwM7uoR3bshMnQiKPRU5qFy2Derdcdv3oyLrtISoVUHMPS/KVcpRltf0W6FWiKS
JB/wA4oNBz5bKWiNEKizW3FuulPgb0djtwZTvFZN9x7y/IP9dEjnxGF6Zx8cGSgJ
SnyjFl3B+5ydwRJNW8tAPHoi0NHAeVMoTgg28GoWz6omST74jxzl1suS90SrKKgX
oVZ927zo4CoEnFGpk82i/lp03Y7sHjaYjEsNnYjK70luppuR0nT6ZnwPUXFvunZg
OVpIPkdCb5c3T78D0ceEo0CS2Uzx69BrVA6gASiMmo8W7LRpuTXtquPtbSaTwHNw
8gnMsOCFhTKXias5WHBXRWkMMtO7hUPD6uzwo2kgGLLjgw68qwo2utuCuKKNvpiq
NL/bXi8ag/dMncMWv7eZL2r8OzTY1lQ2hBDnxWoYqZYupJwcWbQ4PPF8wfQK+RRJ
cZPveIpShHuMhSVSp3dAgE98CbwSFMMWA0VsXs/2pVQvVojQXRpA0U+69e4NMPe1
lHCtOUXQTtH/eSJz9dBE3Qcpf0ku9ZupLyddw310rN/Ijr3zYmBb8ArmthfHvtab
l4xgXRyBCpX0Q4HAZXpkdRPvP0XW/Md09Zq9TYlG9/he9j+8ukHBYlzZyLkI68io
KolUVZXY0JlhVcinANv6+pK2ah/YgETWpIwp9tIFTuB7XRVoI5NnJCxJIT1jxebz
T3o76uhS339j0A1JNEDfuklYotGyq223btv5U+f6Cl+vfu0YkTi+aBg+H7V5x6yW
1vpHHnWEx6Dm9zeq5iMXuK1oPtkcGuMwrc4uOmERO98r3iLRaACKe05KCtnI8+kI
Y2EHxi/FMlJ2PX7svk7wYbbJ8PQ+hYiZZEXQH8BBnVDzHuTdKcMhAwtHMKzS6jjP
oCtqsbFvfQ8PLIYffgyoKlj2Moc1EaHlW58+m/Gu7/73Bknf4FHCfkit7XzcIHYH
/vuhCkHDL96fNE6AGLIC0t7im8/8ISv4g6vx409WswRz+dygvfzkSEt40QT7N2rx
toh1TrbwVoyCbUgvvLfouV4xk0MG1YEePm36oAriicVl/fRdwnV7KutBcEh0x2zW
Gp9pjqF3glBpC/RpK7Vtwzzw1+rb0HJDuw/OamThnHlSNplIp9iU4WiKHxOxiqru
41Mlcv8QJ7pTadVYx0ubTW6Bc2Im0boi1NIzg4nvtA64sNyOqAWVUc45DykXyTmb
32h7D4Q/KJFp6dRvuTgiLXpqZDBJ5385jrZ/rHLrZhpHKHmy9Se2Tym/zQ6vYLB8
hou1hPQRIGapRjT1rtZgLOP7D/JjurR9fgBdr9HAbNFLQhQt1AxigtynaTECSfGu
ID+MFehQ9VGu//n+7pv6GlownWzymX6qa0BdnbyiMclaRLZsCI3wTR65IeBLm+Lw
dryH3rHSHyfqTEqT4LXSz0qThkYJSwOWnbM2SsEMrvFYeFXdp0y8/wjkHNdNmps3
rbUj85QPSw1ggW50H0DY39/xqxFDtXQ94vLqn+xs/B71ftoKWBa0QES/xohoGIjn
lNajjTOdNJtYKR2XFNWP6dmxb9o5x1hi1jcuXUwkfFLMLa+RUGsiMIUvbaZePgR5
qSSHn8AqtLA93mW22SkWmuv8OgSOMdlqeC3b5y/7IZjqlje0NOL9suaT+s/32uuW
IT1FbArQoQA5UChEfqqA1TNOCjS4fKQB/sPRKWN6rmWtGiBigCKP6nH6jMIrVMWT
AAY/5uBgQo1OyuhcOc60/qOe1AyaQ64Hrk/sBCKZyXJNWqQTA1uccHncGs2usVu1
MBQzJgF62QdzhOgiBjo87dvaw4nIHZ30bHbYYJfjV+SQFtGO3RFpYNEQK5wwZ6LC
pjTBqw+7i+O7G/Lbc3wV1Uu7HGIxIZb8pgj0yyvafsDoIse5NYoiyXK4rUAx1uSQ
Pespua9hSU2rrM0hkDLyXe7TlQpmnCI73p6mPUY+UYKniN+HOCpJk5Ywk7YfeePJ
jvhS2aXFB7N4RB3oeZ3qZATnRt3jB4mh/O2AqWt3T57ZkFwAxRBtXKpSq/MJmn/F
ITqq//11swQ3MVRJ8jBfZ/ZgPnbqtj4Emy7zUDc7epeXHicO5AAO0JobJPgdnMeW
Y7yTZbuDO/Z+YpyheOTXE8J4r6ciG9ncw3GxCht6Lv2mQln37Exh86oHscA6O/RU
HNcRH7R/Oi4wuFhNS0KIYr/ONKf92YI7/IpbES3wlAHhjLK7zPc6lG7YL6Tq/4qB
ZntFApj2kdkljCaAfUXdrrc/JkNgc8Y9j/PlbgCqez1q5PgB6j+CvWgaIYASNJxx
2dLJw1lbtEnSAsDKwBvl1QRrPm6lSkSWl0O7AhQWGJifb+c1k6vDZLfw9hE24i0u
aian7CPMORiBXQ9jHCSZfjuAU1+YxC559PO329hQjgQLRkKcKx03kdOalXLhs9fg
MoR3CCoHizh+v85x0PuvKp1bGwqly59hqRWBQ927sEFuPXYoNXznYC7IK3TmegZV
TIn1Lc+t9aeenUlGpBYdugrdGdNAnD22Gxzp1ZDN4daImteKzXIpHU5+t4phSkEr
Kj7qLuKx2g+OhWTeAF6t77+vHreoCQsopHOXlDsQc/jfoLL8mKdu6FdTsvS4hZ7u
GVSePTLZrr1+zyJ6s7RLeOochZ089+UOOJb1HKV8QbPmA4tOkXsKeg1wxGoIRvie
hNqVUwqV14RUiCUgSZ7LK9KhK4mOkjhhq32rMzYlugRucEcjY09qPXPF96WhbZm9
q29PWOIajSzrb25AzzYSXhaovFQ1OCOwlvBj9skamvVVHI8IPAVel4s6G4DwPuGs
Pa8xIPJyc7E2dMfraaLwACWO1JgdcklrH9qkTA48Xb6jr/AT4Pi0oy6FsMRBxvxl
aCrzu6PDXzkiZqOytCO3CDHxb4iWVACiCaPzY9GjM4i5aOPR2pgD8T+xPdNlLqY2
eQeeQ6r8bywehLd9fGWvmjzRbH58afSYncPDcJouyzMR3F2+O9Nm10fslwAZd4h7
35NKLHXgdamk6X5TXWGwuQWdY88DOY0bmzeGRvs1hehbiEQMIewGdwYPKNmjIFQw
sDLodjq429ErA5qfo/LVPjj1S0BYvz33DKTznvkN7I0fXNKbqzPIstlAXxmYAI5X
0BzzMPyU+Yrl304OuohDmm+eP3k9EJkqoyX4UZMeiDMSqKkPG/KHmn4el4n2U0vl
kkJqKK78qxde81KObltAjuZlNFWl3bUFv9qxiCJE2daPPZokkEgxEAJnkuVSLlBX
sBtfJK8bjSoKaGOGuUNc54uRH7ePItpXns53lYRyjVs9JwCc2rEljRG5wtmt7MSz
Zq0LVe5HhONA6TeoFHLHDp69VrH1PXIYJZOayMbqEBxN897bFqzGXMIUNaQLV+c9
qiPA1wYzxSqOOClVs7ONJpg1C4GlPtM+J/tO02CNgk3UlRCuJNAlSXZbfQfro1ZR
G6Ec3SabXInP/hP/JysBqtK2IMnArCPedWsEZEGY0/WcspRjRsiUJXhYlgglijFh
aGYF/VK8dPmYxbqou7/E3LI0+N3GvJnG0kyx3WjAFyoawQEfZ9+gSZAVvAFNzwwp
/t0KdXflx4/23hacvLtpAZatFAfLwgXo/6Joiby9cjC69yVNYtqPyzXd8Z5gFfAs
1uo09N7BBebrw0i3LYBHX2rD6haryYD12djba7nLx4UsBUGYGFjajRC9A/LwMpTr
5hkzLBwXISAsBDvozmDxluwjSIy33uhh1wCi2IHpe4OcXjEZ0k7cD9KAxwh/xlV/
h7r372Mw6XZlzP8kg69arm4holXhS0weGJbDgO/Qirfu8hKmj4u/Uo45arbUiinC
TRbuLgiRWkf7jSwqKZo7KNxpj+ONDzQoQj0sbztC8BWQj2wubTgbnVj7vBt3AHEl
UtnCZalnIxFbDYGs+bERiG/v+2V8eN/1XnZYkoo+vO/XfpuZUEsTepsgdnWgLfmQ
R3zu3IS/7Imau8EVuK0qM/VDSnwwJ64wNnv0E3iCIZZeV6BRcgxmDFhjIiAnMycW
8vHSh069NtgfMvTXpMJK+gD1WH16qQcx4VpWL23rex4B+vHgYctgt82OpcuP3v+o
wAkzR73aav7N7PJMFJH+MOJY2cwfa/ODBF6BbmlCD41YIE5RufliLERZVdlvOIwe
1uxhrTNOjuXpgd1GXm878V1fSGBDYlQ2f5kq1d5783oBOjhJq46QIU/lcLgD2dzv
UNdfZ1WGVEdCe5YnKDuOblE3cSyJOZ/lscQDZaJNzURPuchVVQ65UcqmAH8KT0yM
IJFMYQ4YtEXNh0Ir3iciSDHVomY2uQMs8ldeA+7I49m63aE17FyvuwoQAx2QcINV
hzJbm0o3S1E1/4R4gHxzM59nbIbJQTOLFMaef5SA3eywZvlK7IS5XvLBSKkMGXoC
SMthS3CyHQiu4Xz+8+uv3VS3thoR77IBE0Mgy7pxCGOXi21v/AY3eToXr0tou391
8ULxC2w5MwKRd5zXFKUhvO669eU3W/q/K/pKvAZR7OH49tUYmp15CYdLx4oBQL6C
E8LKQrLfY47BJH25S9C6Yt1bs8HuvsKDbKazMkAXhX0rD1Ny6abhJvceZsAxUbit
Tbbw4cyMI60GB0eOFeXmF2YNqcjeZfDiLL5n+xwEA764Ja2uSBNk70XMzlDKlMBn
RX1M2Cv7jlrsW1BxWQ2EFRS9Ycr+swPhDosnHM4c1PMjOjwNGMXZS89uZiteLri6
QRuBcxzcobbFC2AtBp6IanhwhC8M1RZLI28ed/U5j2gIZpyU/UZBUFX1qzb70cpm
wUSxeS2DfmG+sZDpYEvGe1x2zZS6zh1GL0rFOeRDOtEVOAMZ/7YSfWR5xuVjKudB
ie7ApFanA2fMRvnkF1QVfdgZhEC3YOCzxAxMaQt1iJ8RlJoJjueWYQgJQg+nCgG4
4Cln/hZJZkP8UNEVh8B4r1C5aQUWRbp90a5VhKQ2AoEj9g3UjG8glK2mVBM5WCIK
UtMISKFTCtL8yiQhlTJXyLiFHGS+CwVTTFe+nh244nK2mo77Jkk3XAu3eHQ08s9d
Qc+ScqlSD1JtuYy4JviEYRwr/TIQzOfrc4RcYkjuNT0C2rd3bctEPB1fj1Oaxbqi
I7F6rgC2IK1b0QVjU+kDFR9DZN07LJOK/OBus86anaVbElSc0A6EyUoNzcQBoLQe
BuY8i3wKIJj8AbNnyxN0ZfJnR6253Ie9PAVYgIS8rvG8oUmjNtPIX0dI2wF5KDyv
8D9x1X9Ee+qO200KnR+IZXbmOAuUm3W0w86BmNKIYS5WpfzaQvqG2kBa7fygHQhd
emJ4miQGWN3OkurIkluBom6UrtGy5JTYst7PY0u4eXku5qjCUJXMIupRO1vG3/4o
nJ6rdU5AW7thATH2e0AJCofNVTfnH9gquE5tnwjkdXVZNqEH9n+i5OoPMWyKOWV1
nEyaBjTvXvLIVHvyAsBb4lgf3bytzpTiCimqhXJ0EBoNPogkxqfN9trzruMKD1Cg
YsDJMSd5iwiOmBjNzOnGRpabqZFFwmGiGAJPtS/oQA6fGDWwC02zFtPu+wTeXyeR
X0u1lkL5uReaxJPCiagabe0VkO90aspY284qLWRVde0s3ScR0+reteXft3vmBmR7
QU7UYn8BICFskF2+odfpiRGOVMjqSo2TEpwLI71T50RTNFwhXi8ATzCXc/u26rwm
8HEmEHC9+BpJnO0Ehr/2mSfCJ9RgpRMPwC/SMOG7z03kN85y92YQREYnOAj6gzRR
NnY8kg2Btj10kdhDLzG3wGxOrW+tGcX3ybzCpiPrL6odMVH+ap0WureBLH1bhSkw
6AVpXK1FwE7U62NXEfAhEBERoMNeZzJhOfofp4/Pmw/Z6Qidb6jve9db2hZRL9h9
LV+JKUYEhNKVGfiEy0DizztDCjJ2N+IbFBU2IYB5mCSJuWuoaCiSgqW8FAdn0oYP
/htt3/M4wAabOAeEcGRl6mC6wugjNUW8+N0+5Q0kmsGwosylGwKHnNYtgFZSI04d
SVP8n6QYe1XLdRCqxbePUhGQ1cQdzYTdmKZnYlUS14fcjLtQmoPRed+8V3wxZy05
XLXARpNAIg6ygdsxY83Oj+mIuS5sDPbnX6MwoIOTjFWQ3EUq6dlIbRBm9JDCtkwg
sbrmgCrGQ8fGTm4EnobUFhmXLm7k4D4bvkjA2hNKtqpjZ427b6MtR+c260IUJTWS
+z/58VBFQRGt0TrrBeEoqsNZZq6Nw/4pksPE6M+a5fPSf1MsqgBRC/Y9+e8zSs3M
anKdl7uYvsPyQeUjudpVwtdGPzFivzQ6gmuWtNMIohQ3UAvZ101weGoPtQvWe77K
DYW65+idbjy9EtZ7Mw1yIMnH3xQZF1yo/8KeIGIp4EUgb0byCcwIo2SLatcWNHih
qfupcwq8EnYFvOGqD46JTUG4IQi1deeXa8/FXitNrDJbOd2LhTVKDpacLkPTiGwZ
K/UIAst2UgpLRvxv2y9jUtjIVqjPJB+FNUCEP2AfLf83Enz2hJb6OqEPCsJmzjp0
cJsTixZo/BrJTsXu7icT1rk8RofGmi7kz2Yf+s1UoDJLa37Nvi5NQ4hYY7czuw9+
npkeEgCaziy+l2NJ2k5NbqX+4CWdqWOlYiDoFz2j/9vwsGrbEBg8cLDOmum8MhgZ
06PF7WhZwYvXjSoeLJIFsEoFC9WkXUU6m6kaM/gRw192VDefCrT69wS2SHF7mCEb
kQgfwkWAH2RdK6x/hyJBrqC+DuDCNh1Bw9F+cdom5giat4biLJbgk0fCMCMCLqD6
fwdNkf7pwMEDJtSbH3mrkf2oA8mhvuS1aZOpEl7siFgQQNxtKdlw/GIccP0KNg4W
/JzFTauF/AJ45M53Rzp9f3m9laZwUCIfpANzssGTdxk1EDMlllzDn2Bi5wYN/quW
LxdHcjFj+83P/DrJLv+nnJqVoHs6VdxaeVXk5DQlayw4wco1xptHpKz8KFqiSPuf
nX+xyNGP3gBMVoqP3UPRgll1Jntshfsgo9CtJ8hK+T+XjxZMZZJaqPO7RDj0N+qY
1tEGwJ6SFyT2gHFqEC1g3n5PZeLQjUYeE8DMM+aNuLTIUkBQUgHXhlxPo2DJBCna
lVHlpaaspkkQlYRtyQOydPMC26uRsyYD/blDzrnGiJKD5WQbHPa3qbGlCDJa147d
Azpv8G6IsGu19DCqeQyV0NiOxqx9GjXBHKEtuykzHTOkPWM7+r4Mbn0MMrWm+hLI
48TH0TN0VAjDL/ypOlbmRZ0Kk7QF/pLg/jdo131eocyhfxfv0H6BQENKX7JTiQq+
rt93/4GVkLnGWjQ5Nsq8fxt4V6mAeyI6zaOh8VWRwsQq0LS07yQWxzs0Fas7szTL
CoOSa76MqBIrt5dG80e6A5Rx4dJ/rwJyGkwBymdSQK9Bp/Gl5az0WzTmiBzvB5Wa
Kahsvu9dPWdACwxqTBiLMFkoTRauoOjM7J2GhnRYmZbpXqyCUGmu4SPHiCk4NQl/
2ypJXC4ycPNpw0m2WQxRtm5GJy1Rq1OeChffMlwUL2qcGOk/hFU9ExfPQ23xG0Y4
UnfsSPOOL4jjmbcpbO18nq+0hsZDy9n5UtUDse+afI1LzpCNVFOPJH77KrAUhsHZ
0ogWIW7DWo/1krz8J2lSC56NHoltcH5tiFvwQlbtYWhKUthfwFJfUz7Gxa9yw0Vm
QMOuAfi0tO0K11f0mDPwxmPNyGHOsaFwpwDNVKxyVMhURUvA1VV1JXe5CHGhEaXF
X7v5L5bbr0bBSVsBatlbncFzq0gvlv7aEErRI63YkN5M6NF1FKYhKtCJVtF038iL
PmXARytDDpvq+t92jAzl7qEsk3U0uNDMePlp7FgeHGqN07zAi3D5WBzWWFT4lC4+
vpXBGsrQkg1SxG3cKX7wYWY+rbrvafjSF6mT98+GQicNOPwjTiyHzijtiGCjerCC
8j3RmKm3vasxvZLMby8l/1Pemoc+D60P3YZxu5W7nKLNiLTw2Jl4G1N6BSqDWqnD
dTGQoReCXo27s5eiAqlt8eNdjUaJe7nbG1C0Ia6zw6TnVkgV0IoI+RzGGwpI38W0
R3pVy5RIlpLHzD3W8RxL2+jxSmB29B995A7RJV2xG7fGiaetkHDJwKYNXVZrpDHT
3dFpBnEbZn0l0RnGEwyoReQBPq8DF8uvmqqsAXinekEORV5bfhwj8v6plD8ex+Sj
D4KDZHtXczX+EapeCqzy8lPzQu1PgKyh1ErfPQQT7OMRJ6GQYQiYZBHzRnYVrUGM
oDBokoZYwDH+t+KZAssR+hKBh1JddQKpfRFgXPZXRKLyyr5suOKW/h7TW43LwXRo
njTvdDSA1oDPMn3KUb5Bgdqjufnw9fnHVfeYKETVSHYNteFNJ/YdU1B6O0mEOy9E
+6u+VK5Na7IQwHW6dLpTQiUe4ZIyozgzCQxcTg5efkhB5vH+xNzKK0EGDoU29yS1
TlDG5KZ6xz0CnHLSTJrOsCRTlZyvSaKdF9Nrzrp1wJpMxxiyzhKJPI0vAlFbPKZq
F81wgZ6AcI2gZlUpypfIEj/xJJhMAgNTcbtBxLXPvLkV5P5CkoLcCQnilemeJOGC
CFyMTKTUgFER5Z4xOPyFdjZoYUQdB0JaQY7cdZfp8vDyJF3kev2KrmmJT+3eanux
7Aa5+VJ+BfY27TRdFYrafMsycUVkuGHZ79mo5CXoHuZgOkFLBRF3vSEJD++B1K5E
xMugO0Pic7HaDAnRkSMfm1+7TsbYleWaLapoFrblFd9Fnm+//cHEL4Ve7NbpNhhB
5j7Eb2FgP7ot01NLfIzWVkYntu4hvmQO8Xn2bJ+tSVijde94tfxO1o34sdoOaKVz
hYiYvONaSevwncEjZV9eBFeyYdNw9lGQATQ66+Wmbl9jBiTByHEjF2iamIKqb5VG
+YN95R0VWtXxbs/NKcE4NwM+nSMMopVaAw5eITuvrgdSAcD9/OqQWwOPo9y2sp6P
ZONHzj45PBZ8ek7aCAQgiAxvyK5pg0eqw2y4hVND80c4/Xpvi7coMXEmD7TBiSxt
uoHG7VSLXruJzYCmUymNUDmB/LcNnYxp8RHfK9VHyeRav+O5yXugIAc3CWqpCwdN
d0H9l+/nZxKMP5HBwPUjAsK+KemTwvkSFI21HRTzPCnEIRYylrGofow5cIE0UiFh
jICk5HYeUjLfpKY7wL8M6C5JFQRTnOSIDpw9TzEfXK91LGdVdvCFKSpEu2/1XcRW
SgGzsCkATG48j6t0kf9jpb++Jjlce8CY6y5qYc9pGvuIv/AKi586NDCBgLqDCyNn
4EP3QWEk52SITxv/fB0hKcqNLBbdN5KH2eUR3oK6EIRaYUGpnFRB9rNU5fGiBbD4
0z8GYvFVSFYOL7DwHb294I6uHeYopE8lKUosAfhj7cr9BwSQ8LC4K1hC0SwHCaCl
LZsJxCpn+TM3DLGT2hoSnSrlW2ylYcliaFCKxgvTc9PBX6KPk3dWeV8CiPvHWCFk
TaqbKDWL3bOBh0xvjAupxfI3HtuhMO7VBDuuiPGVU1HzlQpY/9knm1vyO/sTReV/
QZ1aEbIVxjJ3yq5gX8ZDj0Gh+OJ1UFD535TmXcv+/qGKMccGJcKoLYmk4bveebTI
JSve9bS++pHpuPOA3imUujamFNM9XpBoO9SlQGO6vacsPFcHOfiE99Nr3jD5sYYv
JGI77+xgt4CB56SYHh1bdGHNksL4IWmiLifvZDFSq2esAG8M0JvVXg7akJSJTaa6
ZBDFbDvme0fcjL0gKi+Iaes9iRBQhndSilqhF5NVyLXxc0slyHj9NkesJELqeeK+
zlhgBf8I5tcc0UoResUKlaCyH0pMmze2tHIdDZ9a1X8K82E8ZHbYMDcRXEIqwYAV
4v5b5bK32S5ZdqiUWBVlGNWEaoExquW0NQzGYfjol3qVh9ia6oT2GrviiyzPLDEm
QoQP2rdprM5rq2fJBTEE+EsFVejmXd6vW1AdToBuZOtDg+h/Qbc5O1HU9iwKkMmv
/F9NtzvT12d+M7sE6QLv5WV6SqERxxMGxj8qlFtRvKni58IxL1DDvDUYbbUuzM7J
7rEP2sUlQhF02YJgPtKUSUIBGoE3jSVK9Qa+CN/gF4VQWtdzDRnTfm09a2fldex0
dCZXNV8517v0uZEZd8GKTw+ZZZZvofpWF99W+AjGeBpfX4A/No92POuFyamaJ4OE
5f6yG5cIIDFpPEWTO0kxKWT8y5BZ9r7i2MXglCNUhxzhsAQfdxTKIcrbR/p29L7Y
Y6hpbjqzM8pRl5PGZhibQYdKXE/5Y/HF9DF3ZGUF0GRvmmTzV1JmXqGXvCgkHVsN
ZjLhz9ltoarvj69dHHlLJg0zhvF11or5HxW5CPNtNCFK4/vXNgaE3wFm2oFPHpS/
82OSnF9yxbZuwWtF1lfgWrnhNYIeYmOcs0Lt9c2alNSfHyF5PKujIGjG6LRN4Vj9
Wz+Va0Yb3yVpMQLqSajWi3oZslSfPqthx2I97+Tbd6WCCrYaVwS8s2wqSVIa+NmF
UXDugQu/KUvePm0NDxTqcWlMuzZH/EkhL2Mv6v0a583V/6ax0uTFtqKK8G5U0C/6
61c/veK+SQ47nPsAnGvilQ5CQZGqlXK2qTEkAsAwMr/pAynztnoMnJR7ux7kiDaK
wazeHv1Ncf8jIXYJymSaMVQF4TyFYfir1+w9DtDMuKRvpGpnDj6Se1SuWgYLjQwF
8mchN5M1Ucu7iNZMSNNBKpFbmAmDOl13D/MRtx7GIMIcNNpkm/8ZeyVhCrdjSK1S
KdSRWO4mzkxKOogdiuIfryX+547yPBDNpeh28+f20FcMB9/nNcFJIgRRHOXdoiJe
JSvCVtY23cGvJ11XXfgdJpFTlbTSh3JYgVWcBCLZCe1GrdDLTuTuxGOyNQ05AJ7t
8qIZf2k5P0301Lt0t/3FBmn2vgWxopM9Pgzb6dmRYNhzxAsut5E5hBlHQwjFPOmm
9FNax+yszGOPuipkPjmPZIvf9miZM/dg19n8RkRRWGnu3P1TNBzsAdGzgjrXcJoX
aosxVnI0gLEyzh1Mfx++XZopnZt4jhiRG7uLd+g0aUPZJk95zOUG9J+HyOgsYawf
BODeIAJ2/NixaER1MGeJwNsCELfrn1YtdTBMwkRRG4jqhAXMn8izvGbQYcSwoWK+
9ZWB3Ho0eCzOV4FcmP7Wz/9/19//jD8tnUlylD0z7WYp/MX2oRThTsuYNv2jmI5Z
iyH6ZBfnbiSPr+a3Zw/ofovoDdt+agD6Hgjp0+VxEdiSgNjBVhV1XpnCg/ZlNVzF
2bdD1jVJRkeMnxNDc3AF6wmXTcebqfTKplRNMTBnwVn0FJ0+4Y6x/g7CYUqg8n7z
KGUtNgl0pT0pazAtBKiwdsso5SDRifQCjryL8g9EH5Y/en0l8xIEtfTJgHxdsn0w
J4920yHl9zGpE4cS6S0KyZo7flG8LIpBuTFxS3lR6MfC978PVRFoivYWFS1u0Uyn
dmshLP83B7xRzDDD+9FZ7/QVKGRYNtlOPTLj8QlcRmKZclIbG8DaU+mplVlvw5f0
HsV8NNCLLrRy0U/xFKXZi/39GhCrbj0t9AwB6tpecp50/cQ/LWJOa1gAkVrtOs/O
EYgYjdsJd3cI48TOmqGay+ayc4ZwkyciI1agbnbQDPv2sE0uvD9QfltiCwWz2hfT
nNwvgjWSEcw2EG9dN9rWZ5mHCCAk9PjmBdxgv1vaACr6ZyijrtMyZ6/YEVoF5nyl
it3zAW7fS018Pi7YV1I7sYTR+seXsfJWX8OU3THWxPMw6Sm/1H5plcnuHgazlsiS
SHDr8ipt4RZBY+/wpk/2fqDqoEzK6I+nfWuZ/qmBtwOt7KMqzayf77qpl7X9HbAf
4ibfnk1cJ6uscbiognNh2IUjrOPyLU5wqzE7faW6V5P8pyVnNANK7oeCu/m1XlMh
m+LYTG4OIFYvCX5ek4xE5IarAfEfUFRXklowz7xNV5tsr1UkJfO0hebcOhvHY2Fk
WB5WcBuCigPGJHhvXpDpKe0C87XaL1L/FduJHELHNc/T4j048ixreTfdGE4OVgCb
sAbyFeI7sDVo7IwCq6JbMACPXitn48NLOzwYp5Nsh0PRMQlrNST3GTfwxZM0dVzj
yQez5hNOQE8xxS7rysN51b5vlrhkNnGmkVYLsLERc2ckNIYFeVvLAZ0fV6oh50RM
DCUK+wdI+fOtbZtIzqnKqBlHPY0EpDb6qLRTC6QFtm5CcaKCOqP+u6LUlNNi02xh
adwBMG0L2DYeph2ZJva/b51XI4s7dhLZfjK1MFTBFzCaG1vek8PByhbKw2NObx2N
ayv8M4+/DfLnyRqsK9RydkQaC8eUzBl9J+M7seT9PlnikVDadjt/PKnpZHSikp8n
Wb2F3/0JDy/ensKpTb+rcqFM9GV6qTeCJqmyrbEg1SROVsqk+x1lqIjgUmLZn9i0
/PkCnRL7jR3tWFwPB4IcbWJdnjbfo6EPz0lV4evXYki0Tg3ZW01Cuj0eQlJ2aAaU
oMoWk8JbGbDysov8f4PlbqsobVXs4Buhqi96WR+Fvvo18CEi6I7XlZkvlknHXut/
AEeD18pYhhDUHFO+tcfMEjxmcZ6X66ioOJmcJZI/4WhMcnJ5t/d5dISmGpChPkWt
Pkd6NTeZOyMUir9wyN38gN2JiLOHXQFRgnm2AeyRl4/hjFNfBHf14ctEzgQE9i5x
QO2ERRX8Fs6Gi33qPcRid7uEykj7B1yvdvmh7r4o+f1z3JSZnq0bPmp169/2Qthr
v6CHwsfq8KG9qA6Bq18wHrmefir3HPEprO0iN4FHUIm2UW5oWbpMXgKzzfBg1DE7
f1zqLI6Wlvl6JLQwbLNGvng3XJGXagjG/z2Ak8hoDMUBTnNtS9cJsm80a0V+brmV
/DKieQPFfRyWIpTBNYpN0WyBS9W4nkSKSHbzcJj01kmHjrTrjaWr7cIO7GZTiM1L
2GVsqw39hRNIVAklmT7UH4xVxrMRoYwgy0WL1MrgLhwSp6UsD0h9Izo2p8qKBoL9
XF9TFHmkEaleBA1QpdRY9CXmlt6WTnZYGoW9SUKIpZ6e2u0diIlU/OXab84yVRGU
s2uDP4VkhZx0eqJlM6xmHFueGRNcn4uWCANYHlr1s4kVGSMPth0JA7/tBHCJph0f
TVweoPjK6lA5iNLu4N0iYS12qeUzqW/vDOQ4Gt6rXqO0pMmWTM4fXGRarvJlF6Wn
ViOm1Ez1OdWJu74uOWuV84rNd5u9Unl2vQ188LhiVBfpsZAVLZND8UKA+GC3uvTO
XCyFePRHc4bNt+2EodGapnFdbnkKZPojiR7Iq7W4XNlpM07DA6YJ86IXihix1WYA
5eBVxTXlL36HtBVk+9XrAIJfBEf351zWBg13LdWu3WuAacU5xIhWrDLscNjTrfCr
0QjoRX5MRsM0Qk9K3cqq9fHoCTzi3nvsUImNpCQpqkiuCbRQtDTFBzCywJ2bF9Wx
TytCyFbqBnisple83dsbXcS00aGQST406lWJQU1E9WZC/9AhOQS5n1WNcM056VM6
11H26UhBaZsBLYiGb3emjDe1ocLZe3o0x6W0J6mz7LFWTDXQA8dd/KrDxLz+3gye
EI+hXw1InY1C4PAdilBAL4y46Al13jM2KT2GUe2r7NvgOAsKKRZm8Gp47bt9c8F3
OHugfRf62QDt2DNba/RRbT0s+hCMHDMyGdPRyMVkSOUXFwOLXHym47FkCxBZ/Xzh
dN3ET6fqjwuZeK8bZNod1jR+a4y+AKFxVhyvks/D4/Euf/pdbxHl/6Mhhq/OSd2s
H4PbAeT3oWsLQumpvaa0oo5YSVQ5MxpILtuIdfODRDRFURyfQ8IfX6PlLLbG/DJ4
r1hQvXEXslrpDzCpjO+Y9N0ZO+gSvGbub+pIGbfS5+OssdKXAditM5MO/e2hmNCO
wk2VsDmq5IRxrRsiZ1py6R+fZ3whpZu3DQrhpNfLjCybHj+XEILKelOlLKVPZhac
pVooabA1eW7Z/JjDTnKZESBt3Lp+dFmIcfeBYlDQIK5nu9hq2P7irQ1SYYqt4ebz
HmEpZXXhQrGQzDQzDdMggECWeFA2xmWn6QG2t0po8qcOqPfJssnKYsrAu8b8+blx
Xr9mmKbAdOMtHxyUQd0KF4AzS9/UvqPtJhZ1zHgPJW92iknmDmp1YRFMUJA4mlPj
Xf4sa6clnQFCZ6HNMjgfygWyc/dQxhJylV32Jj4gQ24X/TkvogbzZOX6wtF5C/Q0
bTlHb+KWwwDFDE822LtXB9gpBrFY0YV0iLN9lAtqlXS4CRJNmEJXDCrqD04UH8IL
jtZYJ6DoEtj7ityKrQNIiZsgcrjdIZVicRC2EX00s/rjrr7f9dtQ/kZOvttLlS9o
yaiyfWok4otT4LU6ZQkLRJPbQJNcCn1cnwwkc8kpO6TbJmRAH5BHHAtj6NANL6lR
X96d+KRozIBgkPArhrKbiIWZg7f7eBpNPEeaiN0VquBmnVZk0aClkHipcYoqEbkN
GvYmCY8GrIyVQarafipTwNVPJlkHGN06SL1lR5uH/R/eCPsf0ASrWtvv4w3FWgoe
dWClG5AIwCtIuRh+0nmIuWCJNEUppxwQQrq01IaIfDMR7sjSX3emDxfw304oCNKy
eIrYqUtxrN3FKFg5s1wcrGGd4HurPlb1fjNV+y1ljx/7Kas9RlHnxBub54m6eQVP
4gPZbBM2YOiBd7yEsvyQFpBFwpUtI15KIQF5iQza2cmc/bFWTZh6tSKfNZpjS8xx
k6+YLyaCv/BMXgFlxdqfh7D0mDkW+qDeqA6n2Ic8IlxJLRoF5sP2hx5UDQ/iY1sc
ij+LVAXi6AnVOls5ErfcuZL2sWx+gVSSTtgVzZ3W48JYG9zF4crwxe74Y4tbnciS
AGtl4kF3zFxe3lyfSjbGAwk1pEX/5xRZkzEtiu6v5ZIl9vag4MZUw1ltBb3z0AAN
M5mHXthSgmQ0kp1+u5q7+A/+A1X3O4EPy5ebJEzUna7PiuFdakVlqWQzmGlFdGrg
ORDZFmi2s1DHYcngTY+MkfZIS+6aRatBhD9dBA7mxVxWiVdIXeL9ihBQiyS+D6uh
cRrcNIQUm9ES8Hu9NXuTkXccalh8YXXfArzv7ebKzfITenRHT0wopHaFhWqWEQRg
yEtYxNSUbBExyf5apcQ/NJM+EHNuOUr2mJGyR0ltVnSSXGqK87EJooEopH6Cu4c6
vGKbMFyewv61QoNnliZNXlIBGs/haNgwM6m26Hb/j8qT5lEtexNjAvOC8hbz1JBR
Z1IlptT2HsolPtNUJz3S+88/pszSGzZ0EmfUbSOAUqeOinO8OpXga+l3WkSPbZ43
+biMTFAilrtHZ+v+xtpWfW3TH9rxLKlQ/Ay32czoLmLkUUaLGxLCTT2W+4QaJzGF
dgTc4GZXSRs63k7OUwjf7XExQSnXbp7Nwi47CKgeoPev87L68aW/hvzw40mX9Qhq
BNGcXy5Akttd7hUrD/ufGMUH2H7eJISkZP16/e+Zx82XNGQZaJ/tY4ej6a4+E4k4
uErkliR8gDqFbS8YMjalDcZE+xyRpGCW7MhA9vdfGnnheNzml/vhjZg/R5oSfp1a
Kydi4aF7dsx47Xv0lNKcUss7Vb6O5iE9di8Hx5IVwDiTZ67YUrqpG/bTBemlHb5G
zyLWSXJMUOvOJBteuLhtkWYp9+hBylbFVIaw2hYSzm3MKA/A3GLpcJVOzuJixpg3
YXLHnFEE8jkiEPBF5e2udJB+9dCzq2/pTS/aElnr8dlhoizvL93UzPurPY/1NVT9
mmwx/nquNx8Bjf1tXayfnsvZFSFeeNeOsDfx5BIXLiGGN6c54YKxdYHf2JeiBOAQ
2diDB5uz91h2jS1lYq0GWTgw5EW5jI51ASNClFzvzq6VdlSa5fEvfybNm0YKnP0c
J9/Oj174T3U9QBht260ZLuvHGX4UFbwEo2UYRcvQiWxFW8a48MLU7JVkzv0Zjvul
o8x8QFdTRgz/OU/Hrg1okx0Vy2TbhrQrPT4FeD22gd816WZf/CBogmcqoZ3JfQ9y
YTlzmXB2SXZ4yFBrrXonmor/IDgKHUU64/53rcx6m8S0PfFpe5WWMVSW/Em51MF0
AJ6d6ljUYV2bGWXLtTav7x1L94ShxZMDXFoTx6Do3+3u3sIjMwllpeEslq+g4udA
Rgd6qvZaY7ycIokk8tCTs3VRiAtVFTF0IIrd/Ed4gVNDJWEHCPfyyfF5xwVX+pSY
bCDTgIEAEsQQIuhV3eco8Xux0eln+RYfVGfMXEMh3qfDs2DS9cDgmXRj3Rd9Sb9t
mPfnKS9tZiNZR9uhrZpavfQxcFGRYuU9sTlsB2Q8jfGI6kL1bQyUrR/tbIhDZLyE
sOaQovsCuH4D83IyCKGvCUQp0Vxh6oNi6hcJEMazW4sP4v/e+kD7LUxmtIe8LEc5
e+BURZgOtFT5C8Ij2r285HE7IrGNTcQUB2EJvGg7C5Ivt6fBST1akt8oJuK/XTSn
94wPi+oLrTGaQ0AsqucCVqClI4a6HoiJUM663QXZfh1I//kK94bSL3SsSPiqKRSQ
z4gfi/d6icOJXfWu2YMRAErsTyZx1CG7lvM1eFuIT/ilZbFDRhDW2HM7Lue8hBVH
8bY0uzYq4VVbOwTz/7UTWTGGF7OMFCytO7anaKa1sUpSsdTMzU4G41fuNDHP+IYx
AvqC0VbCYeLvUTJ3jwFjWricXcLQGsgZIsAuL8dSN5E6J/EHIfisKe/RG4zX8SA6
tmH6a1EuVxU6yR/EqMsJWG1Hec2xN++6Roqy3ectZmPRsnCMJCqRFzV4X3xcPF8I
FBuqtXQ0hZayiKPNsuJSYbl9v6gAE+dTb9kiObDuC+fMVJvxf1u1Vi1ICAvEyqX1
Q6vUsmWsY+l3qLZXQtKvPy77GdeLclD8DaECe0emicxHL5G2z5/1VyJDKpAMB489
NspS5DFKsW8kX9SJKYPPKbkfWGscDDBXInotlB0FA5fo1pbVTDbFfYVDbeeuN8DE
1rHHKD5IMKP2og+WO4fvAfa0y2zmhw9zts+/VthiOHtaKvkrOm91VA6l61aYAkta
fqmxdqRAkgN8ORmULd3ZdyMh80xxT/wByhnckNiedf5fWo9rT2fNwh3wMy/S0G/C
UGiFzGMpcx3YrvT/dBZZgn2JnKorZ8HMeBJHW24QFtsQs3sgLdrKZQyxxXPunv6t
49jegVGWBN37XOEVOxYO6kT4DgDjL9YuJmakr5RsxISuuxT5yazViAaXmimmRNFo
8+fJ+jPq05fTwYfS6QA0A128urCJoVb35Al7YQ677sfnC3/KCPlJodkP0Nd1DhgB
RkRb4QTZBb4adGC/7Dxcg2C79KsdpPDpfhKenV3uqabutVtPUD1Fgi7k0bnoAQP0
PVthh3J5oG9RFxKMcVyNJyJRpuAMphsDuompWaZDOmiy6h7FPQ25pE+Ck/rs6HfN
I6Z+A4N4nLtxSG5BTxRQAsRilrdgU2H32SzgPlYg1wqNsW51dvAw3a5QPJ6PKIA2
i+s/eb0pjDxqyqX9guMsHBgbvyKPsXfcIvm/Gj8FyHfLB8S8lJ4PKss2G6/zNbWF
o87OD+JrwhVG7h8gWfoymM1ldaWviehfgB1JVe1aseuf0JsNaxFLSMEvsbk97HlS
PH9I8FFOUktekfd7rZH0WSz6thuMhl/lyF/m02bwBKkoEuZjjVmOXra9wnxIGBgV
ghyq25ULibdXmtJe5ArN/F4rAjYKWSLLnvhS0r39Xc+uYonY6jF1QIXm4n8BZxey
hfb4apAbTFmwxYCpytmsGxFCFzSgUv7GpZgbJPII5GdN0oliF1cqVoJoCOOz8WaQ
OvRRzApV40LrT7Ye7IG29x6co1LogkqO5Gxg+XqS9kI=
`protect END_PROTECTED
