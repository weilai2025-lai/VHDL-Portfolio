`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28lVuhx575tW3ji1PqY+mRB7+/Zw4MIJs2rIoLA6oK/weBxluLb7Fm8n++fCZsR/
HomEdiKGmZx7N++3OgYz2cabF9UwuK0nvxZYssGrMW1KJxsV5u0wbzXtrRk6vSuY
eb3mLfCcV5s30iwKNuXDtl/zDDoo35N+AulkYz8q6iTCN9sM4EkGfocNgtr0dhG7
iXSiac1/59MTKgr+i/TvK4Z+RuNlsTfCaYQVwvUbZ1BZgYDVmbLhH5SXjL0fRsE7
f8girWc668fe+7HcVrbyJc4dAoYGX1mu8brw1OhG4FcvlTX+u97CK172CtkbJGjz
Ol08bfjfKwqtoYX1vdHIDZPsv66wGfOfqxcQNEPGGUrdiF/7vA3lgkY+BnXreOoj
IBGentDbNkrKrNlagZpzxdH92JfdiofDleW8W/ClGDlBVoSBVU4lD1uz+Th2oNMK
KnMrMHxi7IrCIgc8RMHYAYPSB+GeT+Ah3OE1BqeLqTM0nogwMilMwUB75b7iA7gz
SJJHaSqj0eV6/4OeXLfKeNZTEE0WPdTem9fZyOcjAMZsU0OkS8YbLk6P10TGQXn9
BUR+e+OqRc2L9PeBcPkGom9/9/Yu9r0845z9ncxFf6zQ8NguIjOxJwIJM1yoeXbc
DwVFCIf2uuSumSfdbJAVy0P6QoF8pJano5cyUzLbNdx8y+oSyzP7xwqtUGQwGzLI
SsSf4yQRLrwAsFPMTlJ0TFnzU6aS8gORU0o7/EikGMIMaKw0UbLwUNcX+qMmiUra
1OfZP5g8Xi3YRN4vfP5qUw==
`protect END_PROTECTED
