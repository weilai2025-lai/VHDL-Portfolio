`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qA1WewfPxxL5Dp4hq/4h2HVZo2W+3yMrR3UOvO3IpIWin98jO7kuc6EEhQhupx52
9rSXrvhiRxoWzSvQ0MZu0Wk3yXJ7Zm9Gt30Qfe6Z2APFmPZmHcXKqrugW57goGZB
vYWsmrlzPpB+fKgX/O4loQ0fJUTRrwIpTxJ4s+jud44ffwxB0S42f8UY2C0vp+u6
Sd06TYaNPd+7T7PinQHI4V0FE3Kezoz0RzBEqXatDPWfGIFejyXrOaecjTRIT3ur
hKQRWxcFJHndk+A5WA/b3guREDBgBGwUIJtT3gzkXNx3FQIyNpbc0f0RsTFv7eVP
7Qqm+o+DQLP8LvjGo9YOnK9qiLiEbqfLZ2P4ustYi8WJgjLPskqtqLyfpv7BnWes
ZLeU+IKx8clej4XwsA4E6onTzyqSCO0mC89txr0oO3BZAkJngzz22iFhLizys9zV
/3Ha1gf8sNT4KzWMs+UupjWa7+7pupHRXdOOmVmoanV9lxqvkjMJF7Eeoh3KrHLt
Fak5+DEaVFKLUkhsXzkR8Tpzyj4rlVlFVdnEnIh437ownYlxWBQcN3TtADU2lQFN
27/rHvr1Eu92FJGbIzsnoBKdo0SnJYQGeKyvC/Z33sY8xhbsSmYFQhKCbueJo8JX
cViflJvw6unKJUANAx7fVbJskbv+vDcqkNunJZCNHWzdn9wOnUpUj5/NSY+GuVfe
qMvbNOdvBPxGhpvtd8e/akkR0UjsE6ZzHACu5HNEGsF3L7gz3pd4soQ59eRrzqJA
eZBvvhabauOTyGoJtbEpKb7zH9G1KNUCDjXjezsvCXXRu1hBvY5BwiEXyGr9E9Wy
QEAxB198atLA2v4O+qD7kAN/FAC9mlocInAiJviW/J4+55FqizU96YuyI2Vc7fcM
8OLUf3lyDh4rS4fckTrhgY4AOj6ZdVs+7+e1Ft3pVDIfrpK32EhITJIHBO3fFKJP
yFrq9EeBwPOsXFPYTn3pJG6AVO2uPX7grn206kohK3mEvV0DWgRTJCpl0nKTcGqZ
aCopE8MrGw6vK0nB+Nfkr0ztWmLJS/oSxtw+uBrxl0L7npma+ZO/jeIxzbCpH9tR
Ic/2ngZ0Lii+TH7od29YL4NM/WCSKUR1jBdiXc8P6Xz2LGwALnEph9R3YGk2NgB5
UR+c5ureEnnDeFLdtuoniPfAaxeJ3xYUge3Dbus6TgZIQl9FToTEYmMEmk3p8p+B
og5tEIPN3gLKGOeJRpgX1dIvpgZ2Zyoh5eB7YSmqnLnneF4/Q+1h5wbk/4ixKFTH
fJ7uVTM64YLKRySkadTjlE5Ddmwz3yibOpN40HSW86roypucl2XVV3FXC7h0QkuL
ODibyW32gOEWrb+jJTHexIcJp7fSdKiJNJyE6ArxRNuNzzdsOItJCMzs9c8KySFy
NhdYkJ1j1jBVkX2/DFjvP6uNF/MFuHOJiwEhgtkM7omwYs9UikY469s3VTv6Yx5f
11ugfzLYrWfKjvxtE9mhE4jfmhF/7ZecXE5GggEE4mOaab6dlDCzqF2cRlUfNeW5
p0cRXuaH14dhdI3+4vvlV3rmBmWYRD70XbgHz9Ui/g6mFdv48O93OvFJjMH0kB2J
n1Ruu7rMVF31/SxYEB4ovXE75BoGWxlWsMG6GG7BNs5y596Kq4cSt/Jq6eXUcPHx
SpB26PrGch3X4srFjLq306dY42gHwQIf5EkMFmSWMgZJq7yg+5oG3wx6655mz6BK
h7nqk+gSxo7ynHOj12s3m7IT/Q+3lJvGv/aWaiuEdlgeRm4Cn8pqpNLUyMT273x0
QkfZGPuZN8vZwDV2I8pfRGqaErVPv//cD2dGbAS/FJpoE/JbpnYDb/f4xcZgkFN2
2f6IdlV2KuvcxhR0rLbZNGzt6nY8fp7laRsDhAwwd0hDb0GBvJSjGEoPuHBb4o9D
34TuEBdqBBQU7U1OStBR7sedG3Zn5hvEV2SncgIp/gDl0z1uje55agoAFC+v6R9F
GH+J7PfiyxNBE6SV+2RATHi4NUQ1VEXO43aBbrI1xpZw4xP48IUTEsvqn+RVtkfD
ayq4er08ouFZzfFndPh7fvTlaG9Af8nb1x/uacB2ye23BSnTgslwS1c25xsudN50
jm1yc6nSp+3pzs21pZkcLidwvv6kgaBl+JN1g09dypMS2670Arl0oxYDXdTHC/dq
20V2aU1QPVe/3UPwXO5oW6nysdVpi/X3XBGpJ8A2I8YzfSCBhj7fnQByv//unjdD
srHgFLx0Mc9TFxSUK3wDWZz70Hg+YUKWnyZX7smtJ00LuUIH769v4kEkplMGBfhi
iyT6ogQWM5tj5SStQ0xZ+ZRs+rXimvoERy8VlsVunacVYYU0qI5kghoyt4S57dkR
ZOM8lxOQc1EXLPZKLqZSBrt24iWJ7CyKfi+xDOZA974bjcVl844/f7kNHOs8hk7a
QkFZ8JRCbEo0+bv1NReEsr+d/JGNAalTdwSlpyVzYZpuEzKrkcZ4p522xV0v3sJU
gvzm0qhzkZKuNPBS1XH+6jGW7ykZVu4cEeEtTPABKhQ=
`protect END_PROTECTED
