`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
55H6LvAKP1ysVKPJ7jx2h7uS0UTlP5EJ0l5ghpT1q4G98d0dAXTsqyJ/TUxbw4FP
ZDQyyDx3JIhHu/pPGZItWscez9J4W6CUyqPbukiwdLCVodz6NBjxf0vdeHU8EEBF
CHkWD7b5p8E7yTJU5Q6ow51mfWi8rQVYzj8onsl5kPC3qFdP2fDHbQ2Zv44Kj+Pc
moxbodVXJVIH2vDhUU9cr2d5zG0dMoPyQpER29+3JqXk6fnwfSyr0FqmOVjm5Ut4
caeSaucK3bUfgHepbHbFQtVYqfafrV5Y/rzITf8AhSOruBR1z6fQ76ITMVBjlC1k
ON7oMlSTXJadxRV3sDUq4m3xkxR88hyL8KxC3/RI+XrbVD22tMdjIo8gjAaMJo2q
AK8uj6OSpSkgmQorFlfWo6N54V+jhcu+jNfB6ElHnFh3WAAvhUpyM4023gZpzMzz
fitVyVm+3j4XksoXzJnAOJVZaaecAr6ib4PvhD5+45MzjNZdMxgU3fuGzfCfTIPS
tCM/gBm8DZ57Oi+qsYlIzTtgKriJcf7Zvw50EOpSdGvgSv77cHqlMMNOj5kV4rMc
HU6zgPKfPR3tCu/nHnXJ45QVpkHH6TkiVYhpCOiRW/fTeR1iBRZsbS/E8h/uZxNO
DHsxDNOU/csABu5C67sVwNL7OT/Q/WmuO641LZV/HTIrNRsX4Hv1dh5YqTm3eumk
Jpy3Ad8SkeqfWo+wINMbisieM+4qNj7QVKZsb8214AlLD5h+FtymnQ0w8t6XD/BN
AttVIfvYNPI1dalPdT6f2lZnQuzjQaBakYbGrjugrpz2We//ZQ/4P3rST2C7jQ4/
qyOINTHpzFJsrcYyZeAiuoxBUQJkyV3TASCebPedCzm8emBH9/a35wya1pXSaqrT
+vYo8pSP1ZIcp8UWEANLLGTzErwBsiVfelX6YBD1W0TYGm7jDpDLtAO8poYDHiUx
qYuR8VW7N9uFCWjsVZITUZihsnPiuu5CyoAT9WsmNRFf8uI9GQLJwizpYb8ertTC
D3nfanCs+a6mHkNY26nZbyKkkC20wpjQFxDiYj9aj2ZsxvXk7Z+qN26WiQxuUE+s
j6uU7ldRCKaI+GkYM9XxKUYVm/fvOj3ujEu/dtXGftkUbgUdFjSZXMRQHKBvYIwI
xN/JKZzvbMGF4EA/J/johFv5ZgvmB4qr7LPUqlloCBT1B1dJnCHMn8dbjPP6BTIv
JmMZq58bX4jBgUVjnWyE8A==
`protect END_PROTECTED
