`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kPtYiwXrSziFRYN7OQnoA2ozqKfnevPLOU1agfvnSZzr98apRFqeO9Yi67S1Fol
nQ904fPHYYrHHP/WIT3WJLWlDPrdBIsEy02uWrCzz6qWMNOfJrpSqdEBCxoLGoR2
qVNpzDoIfebEJmQr7B15Jj/g7Dk1/ad/aEPmWy2PFdfR428AUqv2YuspVaaDLYFC
a0LTH83tPzt9yU2pnvD6yaPpvNPTKkrnHqOJca7EcnefAHs3O+Bs86W3cZL+Ex1i
X5zGxhTCXRTKRpMcwwByvRQAiukBkCSXnaU+z8i1RAQSbTrNJpl/SCw7qoOtgrLY
yZyo7Yyo4ipBTkSw+xch7eP17/apRWj8kPkIASDfGJlom5avPBYMW2YqUDjhDqAM
+zyMOMTrQHhZ2sHY4m9XzHaiEK39S6rdPYhzT72ngz7WK2zIaC/pMAUvNJB7il6H
ZT6DO9SzTgNL1mQSlPuiFux4UNwtQPQ0jlpTSihS2jb2koV8fZtza2GPjou7haE5
M/6i6ac5SuyAee6HwCgRRnJWga3AwXwJcBmJvyDA4JsD4TjTSjg8wOlUnYk3KMnI
YECdl1xMkgCJzzb6rRzp42fEO2kdf2GwNd+2/GRaomDo48pQlsxY0ki3OZNnq9z8
xFNrH7NkLZGHoLio4o1BEVey7N6N1EQFMbAIfWdM53bFPWewPzk0/52C6ScYzrqv
0wiDm+zNV9hQ5Ui677okZY8XeHGWvrfqfp8BpGEwdIYak7aLKtYQgI1wYoq/cv+2
miMejC/FaK2D3TRFnVFCQ1CnUG08eV0oHhxYbwN9ayJ6x73BM2jjQdSiR7XG1VR2
J38bRDzUSJDVl99145cU6AQl4OaVmMt/F9IZV5kY+NP+sC228mXanIn4sXZbjmE+
tvzH98HQyKyQ/sHQ/M6jCKhY45+Y8FvHdSWZ88g9irOB+33CDYFBIITUs/CjWm1V
sPtPN1YBNmlu5+5TFzawKVqNQq/eNxQqVDXf5uu9L8jbCWfGcPvExu0ZuQQlfJ5V
MHh94tpVlwyjEQ703Fgyevs6gIOsqTEb0YY9UHouujAaik29qpNg2RfoWeNHnYS6
8CDSnaz7oK0etlqsJPa7q3RrXOawnNWqofHQ38bXOzOk2zIF4GFfwKmYz9CKQrqZ
LQCaeD6wkdbC+InPI2pa9n53SJ2PsLlKBM+OHB6TcYoHRI1YMiBbH1I/o9qVwL23
UfSZPKXDwa9AaqE0DVRGftYfFtqDjbNW9l89Tv2m2zg=
`protect END_PROTECTED
