`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CMD3XzWeMvisKINNnobHXijIwQcavYYABsMtpcmXTUyOoWjDXX10dV3fL6YPOCG
wfXL/tqms8+6fnvHF2f0oio63lajEgYT8mHtOYa72c0nKCJq2e7H/TbmH+701Yts
Iucw4zOLx4nEg4PTvRaLR4BBTbOxkU4UmQTa9ryKDWSN346GVhWPRjtoI97MBWuI
iMwMTJkMdCGf2+pzMx8g0shaKIe3PJ41YPanerCCKjSndQYbWgc3/JF40DAlckQ2
NszNjAUIDghUwFJcwNO/T6K/kagx0cHFfA61soozSi7CrpIVdWyV7zcyNm8zaJHp
oBtXdoaeyWbqXK/TnptrPN0m9+BmtzbkuDeEFA1IOyYUQFQubdd9iF6+P5CZDifv
LHCkNNyKbAP0DCXiaFZQpgotBv7OgOMpfT82aT7d0vFKYdhaAxEXJ7ioCP7a7ixV
lkMnuKjKo2JIiJ7nkWN+qIvcQlIz2zp+tkELYgKSM7EKWPqP7UJMUQVoHAmNlA5P
3F67/2tn4ss5OymC44VBM6sG2xVyQNtlymTOin2nyRfCd9QQS22z+fbWz9pFePaZ
vbBEcMHgWYPPU3HY29OU0eF+1kNniKshXLYsBU+3qlk9xeD2/CW2W7K6E4S5vo32
zhTseeSjrwKbYGnfAeGqZoqAlc1NnHdblw+zPCIsyJO5uZoj4djFXLjD7rRHXUiJ
OtPbhwgJnADCwMrqI7AFOnd0p0cGPN1DpT/AKUnkieul/saYWvEFWllEHwkPctbN
nCuYL1P/CLtrnAfDAuAE1wuZ/Bj7t+dzeUc8Tfu9b4Ym6FJKCR9+ybsmCYxfZ9fx
Cf8zqWWX9zXCFOITrdJ28qxjJ/HX7Un9gEG4Jikss9Ux19EyyzjoZNEOTGfdoD04
FGcHxYclg36XvSH8HVcz7tC1c1AgmfyEUMtw+02n1Dw0ufInlsQAWXkG2g7pBu/z
sXSZ9/wK5CRQ1qYZiLJNk9lK1uJ4zRpDBflmLL25iTrMa6HQKiY9AwE3oQ1YGiI8
U+zXD6LnN0Isdo1FC/7H0ifvm7EwTqqZgZo6r7O+gNV2rnrrTRHlQIoFT/HdsP3e
8H+MuZsoQEGjuRdEENlFnH2+botW0uZrDx1Dg75CwT7CwILO/HFswqAtjl1ogrtL
4bQ6s8UgJCOugLismTVeGWBSLuc9F1Rf4tjF+yLonYdK9vMc5dS8H67GhIFeKE+0
6eJAlX7R3J1wndcmD3nOfQeSKCTC4DZciQgymrbdHdA57E2eaC+CQrsBYtlIU0cE
g7MXraXa8KgADz/xkU6DyBOvZr+v8d7pfNXVEd9rhK7JSG8XPDLVM2vXOdpuXP9e
et6OiIcSp5fN31HB7/48NNWdvmBHk1IzIC9hOJCYdzADv1OGaYP+dbrJa+5UYyaH
OnKIlzsAY0M2cLBAy2A3hBzvMi7cxorY0KqJ72kKPEQNthMMKlfWHsEEn3eUT24e
KK6yJ4Rp9ctaDJAI42Me76rf9Rr3bY9R/JCmCpzN/Tqd/Z8TRorYFS/3XHjtX5ja
1+Jn9B/8Bru2u5UeTYrGgLhfQ9i3oSMSAyiczktJNln6TAgVZM2gAhKhVQ2rZxDX
LseBp1DYJFDeINT85ikAEw2pswjrJcLwvNkxqLTD08ZlNPsn8IoMlX0AoYUOo047
U1DhQxOEd+WxrFz1EM1mP/kwxFl3GFTH9aGQ/O4fGq99PziZHla60BJD9ZpotRtz
fHmRDeDWq//h+Pef8P2Lafs172iXFTsDEBXc73DxIoXSFeecpF6suy3HxlRuhIiX
nLNwJ+o6WQvD302BOTZJmNFGlp4sBOl/QI6T4lSpkAhJc3RTix+g1ri7566GuJqL
BvAxzuxOcKx3KhOKbP9kuCiL8Q3byKD49LvoUVJ0+6sqTuKB+7bpE2Rf0f4SficC
0htHStXoJkZeLaiBfS8xFoaGOt2nqRT0U8BrkWzn0PrPnF/Fgg8LO/kVPf6RFx9U
bjmlxEURP732ZjNVQA91LT1GL3IYrV4J+BAP2sSWtDT+b0biBczZzG4In4tAOCax
EoG41lgRMjBdNofV3uJFscsQwJboYZjzTPfWbUvcvAak8XpSyKiLW0fIh+fFGG9G
vLXMDqHZs7rbu5kj+gb3OWRhlPTqjzI1mOFnaiQ6gkxq9G77LYU2MOaVjoBkiSRj
n8yQK23Kt5X+wdVZjq0N1zCIpaZh245xcdwJRVJ80QMaFB2GC6RYeK2CEue+pYV5
ou9VpXgVAaSIqBV2gmZ8IlAl8c8b2A3NqZsKNPEb4UcnPronhCwzJY4nfeZyMqLP
vEkii8xPANu+AlWUuBqgaW4jiPGw1knaTX3QMba20hW8GUJrvZtavGIayWC0VIf+
F5PIPzzMEy7xQm+TKXJqEDIgwdYYLWTr77OVktdAXxAuHe2h57JOlVjpWtyt8+gj
Uq1DuCdDyCQev6mXRKstmuVIxsU2OImqoApHWhmSvNyU0TxWI0xy2Q5yf8Sra4Zt
UltDQxEclGM530o1QNs7oZfwre1Np3JTaxFIpd1Y9T/2EjxHgZKjL8c/Tbt7YNcH
mY8SbsP4oI1I6kC3zBqGQFy+kdPuDEdyt5BhNg0Om4pDXOCz3KZ7H2rm9rJts+Yg
KxD2nFYKX63dpXSLS7ZXlGoVZ236JWKe2z2eaul3r2AE1FbNEb6MKaJqYztac1tf
dYBHjhfAUKs4ZPcBJ/5r21O+lgLIU8wmzVw33IPdB+6LFAWRkNOT08qaUqbTR6/X
Q5dgflSOEvhgkLqfWxWEswEnqq/Hi3JECStdZ/CqfFRhI29u5xKhtmTRJriJLxSX
O28WnD2L8RaBmyqcqlxVNnhU70kJzy8u/ZQ2zA7Tmy11dREydvHtkugg/Nmwv1Ln
riReXM6OLmg/OXIGb1JSUNpobU+jGRQn5raIy6wsjEpV8U+0u+SyFvlPRGQGsUAH
oiZfVkCefnWi9slgc17DlyhOW/gWJtFKt0aBwJxC+/JH4h1jtZVaWLLE78P7bx4y
cNDTPZdh7/gei7HjsKfb42o9tXx8qDtIQLwBTqL8qtokr3clySY0DZY34DrUErG3
7kx0U4ItMfWCAUO5w9cx+X7S2rndThpcMUI9TwqEjyPi6VsiExktG1xbOSoZ4dXa
xe4uQ8kT/hUNJM2TBEgsuo8ow7AFeo4NqxFl2vGsdoOuWwy7acqzxz6E0Pf+0Wpi
Nk0jHm60Nih5hVNWEuNDv0IsHpKOTh6BvIVRTHA8fNXwggnay6CX1uT6fRiMyVSd
3Y4VW92C338YUKjrgLdUO1MoxhYiHELBCKpYqnyw0trQH+1rw8hC3aFB8JGMbVrA
yXEfS/zSAaKG6F7GdOObpmcRM1kZNzu8/4hf/i/QhWwBFNKLGE2el4ZoKXjaE/8c
UszjOm+PENeaYrz+RO4tbXkU7E0apJEu0IeH40uMPW9PJ0VBMwuc2GDXOoVHYTSI
Q9vMtvq8utH79q8pEIoCt3WbgOv/EGbr/GRZ3rkxL7znYhJvpkcqWiK/K+ffS2UR
goi9wOq8tmnO4k5FnpOUmBPi7I+i+Ksb+WU3KwIUOQ9mbpDwcTkX00BK9CIjGedu
ACvTGzRAlDtqt5SxIY+OoHQ3tEGal14ZdwUL+xagrXmUnM7sKCiOysOpkdvI5Onf
o/uMYUMy/l3WF48aKiV1enJWcyk4eUQAQOAPseguAv8kPrJIW0PBSeCGAEkrmSuK
ljaNsWtyJfsQttoT1b2X7ul9DXIQ1ek9td3NMCETy4k22qNUZUN3L/ln+kG5/RSS
URknVCcl4q5y6nfdyLtL8EZaeO1jSRoeAbw+bqdN0Va+Ee1xrdSA4uOCJXstw+2F
PNRuEWa3uEjUBC8LbSzj2wb8neT9yjjjxuCc2mm//uo0t8PRVIvsJQST4KRyF9h6
zSlnywlmhi5GeEMBC8ToS6MNAIW5lYudYMezcz7dzkQdbULG8yt1Y9KIEbjf3WVP
34qKjhBAG52Vl0jtGjkGa6q2/naLyW2BWkWnDQxia7I4IMR/8goGdjsGCH7q6MPE
dzKjl3hgGP5macWHmXN2kUkmqX4k0NOC2ElqO4CmOafZmF/xFNgGq936Vc+VI9S7
y9DTcVLL+TZpoB2kVMCJZSYL6MtMZK+7PSeUes92td+ymo3gDZSL0Y7eifmYjUPX
PiK55AW1iO0WMAXExEa1ortVg3U2US99P/PcUe/f0jT39JRHmEsBSGzvgzZLf7Ld
HyCEva3LIMO0CzJMEFaDJMIkec/jgrct55iEpbMe97OIUCeyhaQaSub+6QfHW5ZQ
IQp7T/jhnIy0U7TdcKQvJAYbDzak54ukruifgHGx8Kw8ETDepm3RMFUcTIsR8UYK
K4FUobTZWqTct4w77E2N1wHtOICHk0dt2VWOMMrr6UVmlwZiGGzSjnUwG9p3Z0Xb
N4d4dPjYQ1iZ/kmbfIVolzffl/WQrn+n0UOIVzUZZg/niThdgLJ6+agKY1a258/i
YSttVZCKqtFDpbOlgTfhOR+Xs0UXwmYFz8MCdzVxpDGI0QZu8urknYsyL3ucRAAU
MaCrEKauC/KBRsPAUxpPrLo0rLt9q0AQFNbXoZwHMusA2pnnpn436FEme862W0Qx
enKwAkt5gj46QHXDr5VBueH7M1AwuZCTYppWIzCe+Mkf0WqNgRrsXSQSCuSOl8Ul
Ro0Udnh/thg4F82hTHzoV/F1IDVcE6nhpfdVtKeU5+OxUPpHLoo9lGZDQBnoTdL5
F2zCquA/XYgrLM+V5cvnC/6RL+2udaj7a0d0AnXaYZmj0Mx4oBsPPdSy38dgjWws
ZRjAC9BkLxRFmOX0zNlbK+cU/++EYClSwwQEDLU/6vk3YIKAWacW8dsh72rfhZRN
F8xnyv1h4a86CaUBeUpOADeKsL4wZfHbUfvLV/pLekwkrfQJTUx/4p0dTjzencnI
amQfTO9iV7W3HCBDJ1IAaCLjPbBq/02oZnB51X4ldF2XnOVIaTIkCCPna8keHFus
v+ZBIrAhcsOmSiRINtjrQPhZ7GNRTxIXDdIiqJf6PBvneCfut3i9jil0b+RWkSy6
jrKhKq7tJZdlttj/a3poFIPaFGjDmSS3EqHRukuY7Zq5MoVKHhOoQt5nOJtwg4j6
Cms744F6NYMvORV7RJQC3s2bjtTXENSk2P3ddT8KDBGdDFC7ga1UT91qps6u8Dvs
5nw7QOtsjJ2wP/mGTUh03dmL1djdQzVVipgUgEH9rq8IZBdBcKRw8H/YGjjaxoeH
yZH2TYZUp7vPjbE3/VF1bv6tvnFgGy+ac1P1amsUDLQASDVSQRalsh4Zc8rOi8BV
pOEju1z7g5DbeIjJJXe8zyLkKKnJWI+HyRuMocNMJUyaYgNXLHRDybb4UrYA+lAb
5aEg2HMOKXisonbaycXJcCeyjVLYmIHOWKfmfmm+Z/XHTn/dIVCt6Wt7U69asKG7
aHnEZqzDaeEVjzA7o8rOS9guEKD+qFT+bULB3RAPwpmXySy9kwC1z0DqboaTABTc
5osXa5teNR8R+Pfkisl+Xmgsy29KjOJdwrn+MJTdm2toDcf5NSifi9UfSTTy+l7k
vl6tPJivuvt1D2tnmzd/Fh+pqsAY0LGzcA8NPAwtz0o670r5YJyCVG9miSN7G/3+
5uA7AnAMCUdQ3zfSuWpr3asi52t5BSRToIbNWZdgIMM+naOigTgkxSM02pFvDNHJ
9/uscgvaEbn2PDr3YLW3mvDXlp/7iLuXloJbFD1ftghsoEOemLwBbHMZZww02ixr
d6CS51xDzcRnX8PCRlYDSNbdsbyYE3bPNObP7JBGbvC05H3TkPoQES7uVeg3rF85
Vt20oZWft8aaTi68Rr0slA4L+qwfX32V006uPASm0XwnJnTjVr+3KucLId+YD3LE
+GkDPbVTB0JbmGqKmKdshGhwlOPhINdmxpHwiumBMZPmMAQIe0H46Mt8RB37KKxI
M5l2dBrrurttIwjOhRc3mOoj+hL5N3V7H5AL3fK1xB77RaNk0XNBmEcxAI2mLceO
3G3yPcq5FASe3QcoesWfUW3H6+vpU3Z3h61GrezkselbPKLkJTxJ00i3P0cuUW+I
/k6IWruZpIoYiWOpOzYKaXW+Hut3NfSFUREUXZ+gwIyV1dZtM7LoRbxy+fAJ2kPM
uyvKLQtQx/0VyYJPgIEKaHQAqID+05K5ae3OJ2ddHivsfddG38qIwJ4mAy1+voDk
udBlKjZI7pFbQAXYwK7076SmKBxoI5TWCarsquYLKcMVpt658WNnVjx1exgcLYIv
MKW5Oegca2lcf4sVTar7M+z5d1srkzJY7hmlhIgCoK2zQNInZPJlhagU5/ZmFgjk
3TkjB90RyAEFtKAwCNqFfIJxNYST1wV5form4W54SY7P/5DS3ty+rXZ1fv4L4rar
wTQh+/gvFMBHp5y4k0e0IkdGBmx5UNKF7h7GcqB9O75Hrh8+Zh7P1UzL6LVizm2W
lvxMYTLqo9GAcu7Qlux1PXBlDJ76dQG1TSZaRzO61tw2zG8dNf7uIiYwE/ZnZs1/
7Ycwr9/n8HzxiRQzibSwOld4YtiG+nPcG5v6yCWRS9n6z2403eHKRZmvZmrz933C
fuTufKQf1JquwI9yz/RgiIeBEHIhv1G0hLuqHf8nfnTv77IOc042CBMSNb/lGCcs
p4zeCvODt75jREPy829pIvy7K5Dst/9jQame1yqv6i9k7mkAeZLB6msi06A5/ZYP
QldgY9L+6tuPSBMSJCdMZ22o2yPuogprMn5EnDQS1rNM+fkxpdj6yv3gNe6RtRjM
GD6x5sKr5asFEhOSK/0uXIdGL4l8s5OhNRw0q3yAY6fovULf4OWCiH4ju/tPpXm5
lxNIiqrr/OYRpp7NM3jSTR9dWfhhEXr2vDv69chXY5cqL21l/rIaHOqiuLaYe1KB
64vZNCiL7eywM7Yg1Bgr4hw9zAPHYTI2bwO+4dGSQllvWiJLKEQWs58qMj58xe1C
a0tfqlgyqDbz/A7dv+8inrspmBsR6SbuBDGSbzC4XWGS0U85eLHSUaRIimGmJrPx
g4qs6ag6i9icAi7sPSRzBWXc/2UfOmkp1ckX/dWu6Y8BvSEtAr0wrHP60aWRpXaX
L5wJkjsG7DVvImDht/6Z6lrMrXSbICp379BVAyyXt77EQp1UodRJYlyPPripFEQO
uFo761RkeDp7rUVJhwXrxQ4iCQajWSlIVAwfdO4Fl4V/LnLqS3EdSEh9E5SGdDdy
xxE5VIF/cNinZuZrQilK496MIDUjAn+4DZ/IDG8iSPkWwu/9J4bW7bC4anvqQ3a1
0yEHSaBTZcIVz5XSV0EwtcuiwQBjvcTxT96H3C4YibPURw40a6AxGjZa+csxMVl1
iIzs98YWnYTIoQOK0mBArULdMjnj2CWsvX+Euw/xQ9c7BHrwa6yx8q9wxefNHl1o
D+1v1CieFcqh5lgMekG43MYjPbz8fE6ImaZgfylVdrojE7ocO19ISrPV34XLSUxx
taB/KcWa0Z9WDlJ+DggIhrH4HKCJoCXiiBP3GlvYB5BIeJMwqbOzi6Zweph0JFnw
Xklx0IjKwF/gq9VOSEIeo3JkHXj2zO5J4pvSx8z4oaqgBG/DdD3d16+a17GsGkS9
uKTAMiQYUrOv0ucGQjciq3NM6TgW1a6urOUDi3952VwqMVO4CtVo3ofl2hUGINtm
+fPRFX9eCtzl5RiMIIKkMh7s5yUgLzWU3upTUnFbTztsPrETfcvCS3HoiUShfQ21
BSELQjY2kjyzw1kvkkFCBSYS1pbga+xTM5x/yTknaf+PGjjeO5fkGvMBBELqtI+F
4en4bIdtz5aGFpZfGpU+P5GVNjF8FBL5gJ8GqOyTceMLm37zOXAtYFN7ArZM/9CA
m3YTR/lpZVT3xJp87BncdeLLufafeiy2UzERD8p4BZ2rWqPx7NOssXQQ/1PJmcyU
2dHUvxMUO4q1I34oln7r10PS+4gIP/iGU+P7difHZonCyWXmt5XSYEYSmxz7smQJ
ajASXXJSyCm8aPAl9CDdhej0tQ7NbwWFzCC0tt5khlEGrkZE2NROwiGz/OjqqeD2
/QaLg2MZEntPY1AO2fPzZd6+SvTrmzUGtaIwTyXnd+qb8PV27fqED2MOyOScn4Wm
jay5o2R5OZEZo5NujBANvMzZ5IqBYQBdf/c9bsG0QCKzo7EcB9psFjEdbaCb2KWB
8VoB6OJeh69PgugRsC913v2HS5oIoDmbjLYzdCFIZaRiHwivdMUspfj/8ICUb+3F
8aTKNJdv70dTy0/b+AKT4CSyegp5C6APcXMDkHatBhhzZu4m6nMNxPgUul4UzOWh
Sfkt4vFWx6LvtoaNf92kW71qVkUwpOpRJRGBEQfsyblLXMZsTj54n9aLM9K3kEHp
P+Rp5/0B+e1oXsf/wCHXiv8F+dOtJShiXIvxIJH+QvOIsx7qLRIw9aHMP5QU13V8
qPBdnxG5YVvMPPAtiknQUW9Xdww5k8nA1VbzuLM8vwOsWGezA3YNrFtwJw5h26dl
DPR2o5jD/Qv3z7kdAq6p/yxufE1W70SCMasT07D6IsHCKhYn8NpKAhY2SYSJAU/Y
uE3cZAFzTqsP7txmZDSuS2up8hWqubSXg5mzqQxUG5Gb87hybROi/C5Nq1kxxBpl
uK8J1yiaDourpzVWOoomgaSkbPgXvw0rGCO/l3DgtlIIYAhY7pd2KeNQod8mNjrm
JbElh5ybXyIBd2a3ZS5EqqEJvrKcrYLGa8appV+S/PiwIKsKclHmC7o+FM6f1nGl
ZR1QoetWDYuqYHgPLr7BF8sek+i7uIyOz+8lLxtJlReE5KY40PpjhrDKWXtO6OZn
LfNRqns3F85utXg+qWH3imylEvmADZt0FcuaaSOW+6DtnfXz7+LbPIE8xWSDPXuA
vnZaUONLdep/cGvbQ9ycbMgsWa1EKUY6qieEb+darxHhLwWiXuXHPqmXOBG3iZBE
0LsREkvShULDueKrIm8s/xWl4sImFAm4k9pJdHtN24nevvXpFEbPBaANxc1EyeTD
X0GcsNc3CgW7p367kmHMarIiFTD+O4Wr2YAPklWUSalHMbefuQw978sZcAGP3X7D
Xp1NUUp8r/BY7Lfo2oeevYPidCSs0d9hL+gQJzlKImJ7EMFHUL2ECTxlbeUrdP9l
iKJZo3K9eXQeHPXVMWGnLB0miZ0dJ3+iaLebM1DR0x2459ViuK3FTeSSdIHANjuI
tigguvFiwfJfpcPQ+o6omoCKu36DCU+pNVvSJZa/vSeIAKXoLiAhQIgj3ra9iuAb
kRlWOSryJ9tadNrzMyt3FFmVcBrVUmgw6ANgk9CQFrUJStjCu/g++Cdvc2A+CsGh
+DhfTAru9XV5BUNRQuCIiXfTvCAAuElSLkvJTP83p6/rEMmRlJyS66op5JUfw5W+
H4yrGsYg5090gF8kvqSSWUITJ+DE+iVaVLXlj6E3H7y+bAd7IMaxVHqitltYJ/9/
ULjNiuucvl4tRUD6K/3M/fxWr/vqvlcZDmVJl9V9zxPoAEfw5M7uI49gZ3ThGivo
+pDyMmjVUFlzocyWS0B8n2tTIJ+qsLzUMyz6GR9i+v328s53vcjnwzRvh3iQIe8R
qB3euP/VQ1nYHg6kfnKPKXlESc+BsrZndMQ9Wg0AB0jRyp0//8HVA25wwPDN5F7l
bbPJXGQO9JOPp9bO1S549hRxd7+/taJobcKTzmCH+n9eKoFk23jv1jdBrbLlruQw
q2RwtJQP2HMZcS5IXBxloGW2eMkEPW023c9mTjaFu5Q2v4G11fwDvfaaBDWvVz+k
VZr9b+cWyejI+pi7xq+7Mfgzb4mGI40vAoKIarZ4RVMb7aInZs73mDY1/JzlLRwv
zZPYJmMK+MDhBM7Np2cOQjIcr6g2jRVpI9/Hune/0uIB1ygiP2VBiSHCIkFKLSBs
QyqIv4WA4zKEIuU6eDwVVgemURq57yeCy4C20wXNLisoVr5P4KTYQS3MmB00rpGC
bD2cJZs+Rv9Icef2VKrceF1UAHuvG11jFR/Pe+VGlcLpF+QFgv746LTTLfC7ETxa
KWOuJqmyyHS6spPnZITSptsN6eVJTyUF4ozfQkulp1fOx/bIdo60vDhTcI3P1EMD
GlBmdI184wQkxwZHnmzu9wtuF74KK+k5sIAzaqnSx1l5+xDzOWCkV/vYicsdX04b
Vi5ctBzblhBs2xxioIz9ZyljKi/qZZv5iGQNy3sb6KvVjug0ZOzdZ+sPrqjILkWr
eEEZa+mQduYJGvBh0LyeO3mT18OvDDuMljR+OKlfBGNh3bfbyDu+2dQpFlw03pn7
/+zhXQj0xwWZrSv5a0A9UisgxkzNSLIvoElOMruPPraRiahUXvYxFzwXmuci128m
s9s1K7FSLCWzRNlsRrsypVGoBGE8D2sPs4wklcsTRyzNpO/5ZHkEHMdrdktPyHir
HIUc0awgqpVD4P9tW+NIuJaBKO2kegWDg58UWMu2Bl/X1qu921Ekf2ae+t1bnwks
mRlFhzenSpYg+EYr3yMxkFfxWSwjbSpe5/Bhlzug7ynDbkqMxDzQdubPbnSbd12l
N2R0ntO2i3cqp5zFsye4VaY1ZPY1tswsuLqY9Rvzq4AwsDmyxfmEModLtrYqgLnC
2ObBTQtiPAHJZ9l3HayKmpNGie3XgCfo/4u2QzitSYYfZ1bL1HO3Rvxeuq7+dEI0
hAktt+Rh/5qxu1T8uJcBmvIxhXon46hYC5RrpHlmU950qVMQEEjlT7BARNUHwxa2
xwLYmITvX4IchZUYiSG2dXP5KTZIg0Xp2z3wuHBVZepw6C5HEIkZzCw3dULX1zOA
3/k97wjXcvYZ0R7PBYBHTdDy9MNgaTOWqHyLTQ/Myg1nY+TkGE7GXWPunuK2X8s6
9vMqDY4ucSJouwBaeP2YM/a+U8LciOIbTk5m9BjutVL1CXgMwezwZN9v1BeCY5K3
qPwPLL5alWlDxP4uQUyIimDPCNBUTxBqP7IGEl9vj3sTiKi6rHjEkLZnPTTmjORh
quyrC5HAfUZYBrHIIir9rn5SqFOEOCRcHusiX3sT3KzT5XtoOYnQzgoMf4ibZJct
NncCqDAA17rmNHYtMKiry6reza0SGylv2Jcg12eZTPtUjOAkOa9jM2oUUzFnjcVi
WDKqxI2KYcIk1+DJAFKe6RjlEYPNZEP7mnc7DC8k7x9U1ZXOvKjcYJjX1rhcbW5Z
U9bFNt7S1ZlQYcK5+ylbms7QiX9XqXGmxYVwS1YDxnD1m8zmM3p3j3e/7D+gnXvc
lOoErLhvSO3vbh8E/v+RpYMo4jWgisyBsSvKfs7H206NHrANyLcJ/myNS6iOAREk
d5igkkYAlRnF7d039Ss2/3TfEpe9Bb+llogOpQevOEoN96NFWCNAsL3l+XDb0WS8
5uzzVjZR/JhunFv+qHyOoK6gMcefybcZktF5auOBbGa+IlqM9cFhTjRKFIoW7/ye
1qVSFGVs9CvMXS8ZWlyOV4tBXboSybciPDqAaAsDYgnqMjmLhj7uPscJ3kw4nmGN
puJcxFF3ktOvCer3Lt7ZqmO84PlvOVe3VJuPZA66QEPoRfmhAdXl4VC1vs5hvyx/
vdOzgLO7g43hmS39CrZy7tr7/8Xe5IWny86VifKLuWpCENHjyrPxPph0btuQgviv
9u0shCLQKKAyn7V1s9DhOolme5f6ATI7D8SKN4LrY5UaCAOm72yCVTQOUQNibykW
//nqDLTH75OvbuP3WF2LxkOocam5PJ2mxUvXbMKtU0SuX7BvJY3DA9UygTN/8j3Z
g90lC7iVkzVeytgfDI9R14GcCzmil76ywPrYdvlZJY7d26jUlSzN87ngOFsRwc2o
6ap+AFk1aVqVDvdKI5KkbYlb8WhQCXTUJqJZ+tlj6NQqFqqEbpumVjr1v5kDC5W2
dZB5kBnW9dI3Ii2aZ+PjRuWghHy3YIJVK9VUt+wnPLMOJxcaBpIMLW3xmI6mwz0O
vv3UEnM1vQmP+n4Kh0W5xJJEcrPOHJ57nkm5Du9hYg+QQZPe7PE+qo/mCXefK+xE
lHc1PcAnqNKBNrP2pmHI9NrmEv4W76e7s4G4U6cg8owENbO7FJvK0mLY7rMrVbOZ
Hy/icLrk2sSOEtTS+cnUSERUnemM4vzi7QhgufFkqXGyHCKHfsYbUZbCtr2XLffG
OnsnF8s2oznEWq49Sm0KXhXqchjbnuL40FpqU8lEoDYMxMulKUJtioPz4ye9jfZk
Nf8JQpq5Z/Na6mnUfOGzLxQ7i+bGM7+EhcxH1IeGK3LdnxSZoABqLtOyW6yxryaE
DHz9rgxY4xDHvyhZU/aTuRtN4IoOE89mJMtQ10k/RfKl2W1ixveI3MhT/zcf92x9
YP4hIKsZYuyWcaxCDBZ7Ey4irKXG1NRF17IZnONJhgMzd02g7mMIl/YFLA8LZ2cu
BHEmxsBL8Fvtc4bevFzKUBYnY8oEgf/aMdSM5hqx1MiVh8eNK4Wp8dXNCywi0C4I
3siiR2uHE/BHrTfZ0/2MF6R3w/V8ITRaiPeD2v/xOF3EVfNC4aTZnRuMR01rzB3N
SdSWd9aVDDKcX7OQ+xoRtWoiY/7v+eAaVGM721DJmhdDi2yUn8VUiurqpd8spnQh
54zNA5GGvGC7lZxKH5A3usWxDIWXRUphAyeBRekwHGm2/BGl2YZRKfCjXvfXRGcs
dkuLFQ1avvSKZ9xwghvcmlCMX5Jo+VrR4mm8J8KfiVvB0aBcdKR8er6RS+GNnb8p
iLollS8B9k/u/VyVajs8Ic9rImGjTYIpg3d//1p9lNVqkGX1TiU/aj61nlIC8A70
otpFvkx0n57h1gzWxiRqquEMzSu+ozhy3x/EpdU7dm/OWEqwWUfNYWXO0gJDvMKH
oy3xweu5UC8bbc717NDgBtaDntHDbvXxa1goXRxakCLJZ3w/UfmDQKPIpKrmucIt
rQ/cb0QHJkc5/BCZ2ytaMe+M3/U/sAeJW6DPwCXtHHh0IptU7pm+TH61hXXXsErF
STTp71dvAtIXOUSYiU2qoUmYzHKG7HU+SBdqhKkvIGFKHKzx+NaTXR58gHLlqaLz
jjsRd8S8ZkH7q0l1TxLp9g7vpo63LQW7+48Ua6NdmA5X4Kj5rvisHED2wAz/7bzu
xkDFwWpz03JiDtBKvY00vSyjiA4tEd18Vmc0HUZwygx3MizEBj/c2OOg0W/7TAnY
8iF5kNyWLMWwhTRjarzIzaPE8sfbtWf0L2zbRry9WswcmrHlS4U1zj/dGghv7Kfg
JK2ZIGcFerX6Zqq+xwMwkrDZ3Rw358QKOk8dzGSxvLttXv+QKhkLRaI39rTbE9rt
f0QfXzF6OnOK+1nelaAuL4a3mNv7bqGKZtdffAuQ7e4CBK45IgzivFdaiapDqr/k
r/6T68Hw9C0ye/oogeKy01crCp18iP3+yO2iwLGlehW/CCICw3gGt1Tay/N5ZS7C
rT8zvbPaUdukDPd3zjMB+Ihja29bEFjkaf5qXeRcFZJtYbjScvdiDadrk8nPoQ6u
WH4cWP5g8Mzq+wCg7nxI1EcMlPBKEW6GCifVOWLhqFCoUMcOT86xZwTDOdI4DVHX
+/XiHbzqPdwtMttAGLmyd34fwZkrA3IWZEdjkiI4loZSQTCc/p4kmwx3lf3ATSGJ
BM+x1r/ZvU5HtHceP/SX09AqtMSJKrS85nsu/tLZjaAclgQJHkOFRCJFKhPepU1z
wqTKIg0KkOOQA1cznwqsvFPhdQogdIMA7+Y/5L33RASiyKWOduO57LnttZIJZrKn
huuTfJaEi1UFWUqMSvFUxzujHUHoy+d7hekfggtTocYybOF5dD/zxp16/w4e47BB
SVo6yN4UwTP5foSu1ZDs0vAWbIOGWbqqBNKEb4Pw3e9XxkgJ/5H8h+fSaSWFNhAa
TFcXi7yMXS+k9Gmit90P1dnY2NyCRDKwIW04RLycthr61gK4nHSkkpL0vQEf2zBl
p43AHzpGQ2X2VJ+saRkiTVrhezE8u0DtX3LdZqyEUgOGRVV2iJsBQquMShMGF9OQ
9fbMV4mHbopb3luBiWbA/fKStxYOylX2dgKJcSgXA0wKBJzaMb3ml7sMFhrDFmlB
FGXpTX9jC9cpaYG25u140EGajXRuB1wYcXYkOvtGQqFR+i3pkm0rukltaiirNncK
sOKBevhoQHsnNW1FT8+zCYuKMRWh/2VqFii/YNaVkOl6BzHsVZHS8MTUeqyDXBTN
mLUGMDU3JM07c9cwRceW3sSrZn6wpvcXDbGJeUGnzuJQW7f/NtwznsoX9qigb/nZ
+sRtAoE4R6vP9L/AcA/yfhxtCdCz5yw5N/ZYhLi2IcLMKl/ZRnIgRLxRFCKX2t2N
VXGUfVwuhknix1PhD6iPvRxJzEjgSJvi7iZ0LRs3k1nHHd2yjohEvMfeAejsUPSR
f8zluJt8+QCq9L5HxMvAVzejv+bVvHUawz5DggvPWaBLc1vuu4t0O3HhaADEYkG3
ke8DtK2EcTN08ZKY5Em621GRUvakcYTeQf1esBl6cb6LgfaGzxtd0Y9SqK3xm5pD
gXIQZ5eS6ZzM4nYMNSV4bWRBNDb0k+qFs/TGZRU8VjNnqthUo/BH/fzhFPgM8TMT
Sx0D5/imbYKH6ER7s7VH2W4oY+R/lLa93soizlnzbmyORCHfklcYSd8YEDpLaPsK
n5t19Vk8tz1kYQk8G0dbvLFkr5TFXQvbN77xaG8PNiFxXVU9ZJqSJczYbFeM2goo
9yU/+Q310jPdv+/tb/dlLMrvMu6WJv/2g2ip+QKzOXIhDz1JH+o3anEuOh4dCDkG
U9KP316M+pvnxWgWxh63G2FydveBh492f8oKfLwEHjrICnSzl8mb2ahRtRs1AowB
0Z2uKnkMoASjFX6IM7NiVUqyl8jayWUEAPGr1J0VubIQbQuuMsakFewbITNbtNjy
DkdUMnCgv8goq5ar1XaRJwrXjDP5qOH9rObCtIWXDLdptrwCO8lUyaOXtIDm0yk8
tTuusiZ0bzo4wDWKYQNIGjAhPifE+/DTFM72+byc4C3aPCu1SGfZWxnKxkvpdG4j
KmGvhIbA5elB4jeBHVvcnjSpl1xEbU8HNBPIQ4E9LaxuNkgfWp4ZgnNzpuoikcpC
ZWVlQ3HQZIxUPI0ZbmLnlOfub3yie6WJvAHFINnD86RiJAnElL52PeggUdmk3brd
i9s+dFc+KVjTBwG1BIMkgDH+6qNRKnbCAyQ7Qkr02dnKfMBAuZSo/kxjxMaCSUZi
IfBys3a4gHGwsNP7VZU0HVPH9ClA4cSEIXG9YNPlhaWkr8KjEVHOkdpuPNNCXQi1
XnUsvLjXlZnwTXZ6mihe9e/rIEnYQqdIliYd6tGKEEZOtnDEo98ih2vdy3gcbDHB
jzWQasYMF3ySRXcBcr8WtPyKhVRQwuTXvCbkU1YFzst1CePGnr6NWPqV8UcF70or
GBGJWC0ufc1sVKIu6/QYg+t4F1L5g+K7duXBtI63aYrg1boE+IKqlCFzuIOvscp2
1I6wxYkogwko4CkS7y4Yr4KUGHE3elzLvp97ytH16ByfoHMk/sg0ukr94GqFb3BG
xiTQ7LLIfrdh+p9s957QyssRwXG6kXv/nah8zav+ELA4smihSgETCWdjEU90leAq
MJs+iRdW5KX3Hhr/EpuBhM+4yTCJ1T30daoeS0qDq586L1lafkcGeHjus+2KE0VP
n7S4R7d/7Lvvj3QIhDxUogFiUGcpOsbOKRrs7GH9byvYAYR0UhHcQDx93zv+S2wu
sjcrsS1bp7wp+nO9etq4qSnktCrw4fQrnoe/pcP7EqJxlCzuZvUFYnU3j2bMpUhi
+6BbhylUNYa7+Ye4/6AJzq9gcjrulD9Qt2NgxE6p12XV0aNlOiRo8MlI7bH2lOJd
fT2eApVPogTStzENIvNwapHXx0MffcywItb2vN/PjoNcMCduDCsX1c5yHayyllk0
2LdvdJASVqRWCZct4sDS/A3u5qFMf8B4qC9KgQfEEloWXjbSbNaCBR5ieK/dEiGY
jsKEu2SgIjtS+AYiDPWLIwXh0NpVzTooLU22VQPJKLreTjFxhIGt+AXK1u8kStrD
Kr7VISaMaa23LaBz+Q+Jz2cjt94qLNUFvJLa21CFhDC9820vpZN1FckPZTWRM4tj
Ou0vvNsGCX59M5nCtYHo+qb3gYdFiej0Ozmv9zkvf+YU1Pq5HyRmeMw3/VHkC7sy
9Bn2XHWXC6515NMHa11jDlj/fFaRzYqtGIaIrTkhBntnwmEK/wZo1yh5T42O9d43
7dUaXiQ29xoC51W5DUYQCmlwaH1YcFpu2Z516jIJlwLUJFDhDZgiOSQmcVvhoawy
07Ibb20TFHurFF9JI3XPkShZLpQiuMyWAsfUFjS77+A5EvAbf7iwtcSMiQBdGVgG
8SGJdkUMIXFZwsoTch17PWtgBYgt3Awfd9csW6yQIO6Uf907Qh7jhcKFmeRGZfFp
y/X8IaTTL+RI2v3m6cF3AkOGZWgln2K235go7FwHE7JXQejR/sxA9P1MnjB8lHyR
GaEYmFY8gkdqVWfeifOIw3dprVstk74/wfW7AObWKZT2skU+BbYjqjMZBCatG4qR
WQ0t/FEdHOY547qTVh8Us9pMQ+uxazS1+1Rqmsz6CDKM/d1r0//+8+04KF7nK//s
p4dgZq09xfIO9AJhV82VBmvZISNqloDE2QULN7YdG06ojpaBkNfK2qkovf0sQ6Os
2wkt7MQy9G4/91eViKLVN6A2aAUY93VlyJOlaKLcYaA6DJQJfPRJkg+XrF0WPfoU
8KewhWp3f3pFQ4lJDC+3mDI0SDHZe0ma7ypkCuBF/GwoAzq5J7cbADKCZFBObign
D5XfVj4zRWZLbBc6aejJCgJ6Of4Qv7KDfulDTBw2gp+HrwuObA/+Ldzfu/vV59Jh
crUQYxPO71wX1CEjkxBXW7W0On9sITzEu4+spjEkeps1fUBTMri5iaXmsOp7bV9p
3DLcbZzeTGii1vdBrveEMtsPRTLTaDZvPhCQGFqmyY4bcG2BFZSmrOzBngJvoJJH
HFci0gV1xV8M5hNzyQziMx+K082MFAwPXvM29zjzBIjCb8fbnGNxqndoGzdlN3Ug
jQ2VhlwptgPYDZ18WyU5EdswhxL9TWEF0t/2S/VwGkf60nlN59MxeUNRz4DmoCIw
wGfObzZVTyeUg4qabQiQkWzyDiaGjA2P8etZVxRXEPSyXvavm/sbK/p66VcMTN5C
7jUNQf40FwYNiiL1PJ/y3nECVqnL9lHxK2FetHW9aMES3WIsK4ypSJFSYdgnvvqn
lITihc0NVXsQPSnIGcvdq3Z0uELaazXi5bj7AFVK9vUMpGsPLQYdX9PaahY88TIL
JheZe0Q4LJZHAfu58emAV4dKfbfvsjlOOKfpFYn5eS9/z19Gsea/YtBWRMHeivDh
rda8/xC3DfiB8Q6WcmFZnoXnb3iTCqtmUtN8UcCeinp/jQly28/HrNmC9eS4euv1
bNkfEPRRpZISag7WFSlvFVwTT2WmHKFLKiC1eqJKztQKb4lfBkaJcuSfUy1XwRIF
Z6k/AzQbLpDjIcVQOkPTt5QihaTpolZ6ByYiJhbauV0qJ0qnh1S5FyJ9DaIs3n9R
DY8/aLL99/TWpwVEp42Bp4CyzUM5lJETRZ81Sbs7WbP+GJaSG7l82RI9OKzW9ppv
+OPhJ+q4cFtzHnxauHbYefkjYXTmBDE4cPOGScf9a6e7EwnvRc+aUrswt45SUMEJ
w5BsIlSZlI7Y1yy4ED616c/uBfejCR/92A63rvalOzoX23Y+wSGVDzdtJwWAmYvV
G2Xb7z6YNQTtWbR+HbzbvfFx86PcSnGgOr3e9GHPuQF+wyLe46L4ycAWJDlPhk5C
Bns3DxYCF0FWst8xGhgqgfMDVF9BnP7OGxsFrtODjPZDzMkUk4LgHBG88rSRaype
Nt7KQeTgV4ZL9XV8ZCvqnEttAi13QKfXqfev6D9vQ5gN7h/7pVQ5GjXbVuF/AcSs
z7zYNcqhd0Y8cIOpuPpVbFFIaHPPQCpxOHEdwPlDelgiIrv5MH6NMKSKHFvs0z8M
8iPjXqgPe6zaRJQNLG+wGHeWT6wX/+3fTbmIsefrDQNbCtOQ5X/MdLL4Tw0EzTGz
ldy8Y5fO6qxk4UakvnF8CJKrgU6Y/Wv//k4XdWv+EtZ0/KgUo+lLj/89ExD16zo1
CFnuRCJLQhBhMiJEByhRxLnC//tSDvaZEdTVIoGlgwEdSkEfGgnDGhs+ZaSHbg2h
9jiOr0IVAUOIypvZrEeSkCe5ZmWffgJvYyHkfcTY+eORIy24DsWqx1xEUxQ2YFbp
6g6jk3jKjHbzU5KdUe4c8ArG4IzR5flF8FULU1+oe6Mc/r5/tC8Z/f/0cM3PFASl
PDNNIAJ6ABL34/cfL+frvvZXhNBNoX1CjcMKrk2us0ykoS1LtptCU6H+sWRO3jNZ
BC+IiRKFTsyHo1aVD/oj6ExWygJZIBaalxPTzAuJaPuycfWeWtF506C/nmayknHv
5uB17+Bt8U2nqHDJzC/aMkgkRmkdq6xshh0SdrlXHIEmZU+5YvyD2J6f0+UUDRet
3kHgL8o2JQ65FXUWo/z163D/z10QJahB3N1x4D7XAKMNZdb0vcaCw0sy8R8+p0f8
RMuupii6+I/N5v/brlCkoOO9FAGfBiJxxQCjlo6jIlujP6Q/7BAZ6tQ71EFItroH
rAZr5shUlzgVqajhmPh97xiiF85mVJzxAWeCH63w1Lv2Etcq3SLL1o5gpXmdYdDd
J+cSv1mCfXDX1HJOeAtJ65oosqkVt1/kFl9AG2JQMy9Nvi7ZKpMLI1+KZbCMCbq0
MSdJHbHCjt4DCfKXDSzZwZBiIwwO7oYZ0mxU1ttONVIBrylHkYKT0Ta3D8pCaQyu
jBztAnoa6QRdHY4iixL+TLw+pzMDv0k1J++MMamADO46yVwU68qrs4kaL+u7ftax
B28vfIY7QWdo5kl4ZK6nK1gNbASrMvLWgdJyjQzC6I/f/2gnESOB1JOqO92tW1Kp
IckNZPQyLqOcEY29/Nyzt28JdiwoDJUrPWPRnXBt2tr6NxbBAh0wJYLo2WSKY1QW
8FwgM8It/qRiOF/3BHCdE35otx114DU6btAFvYexbvFdvPDvDK2aKTs7x2d2pDLs
GTPygHj3ptBHbYPtz6Gev2VBZghMHKJsR9F6KO8eTY2aon1qHMtcMB6FQ9wUgywu
3Q05rL3QARK80dLgNu+Wn/v6kcFFjj9co+11BFAaISRS2nLK63A+4Hngqob6mhSg
gMHtHg4hMWOFtk8WuOBraV03Pp+XgnmSD/q1EML+0oMUUofH5225M/wlii7y+oDP
ECC74ua/va/7yTw0MNge9WPd+TcuvHsMOFXZmMh7Lknoyilmw8SB63kgfNo/8AMf
Q5mctuQWM3ignPHB5Ik17LGo2RixCWIqjoUl/lmh2Tn2sf8c4YgWH4xNwKFoBqyE
cpyeCI2qs4i+mZSjspVi7NVe5VUcNfF3eurZzH2CXsKNDp6n93zKXAimvmnazy7B
DhZVGqsFFg+zV0eUHB0JznJmWGdSOWqKSn6dLKLbsGFI0907RDR450b8Up0jiQlk
2hxTDJt2B4/KyxbuPiIbFMMZ/+deOTMuNKofSjgc3bj2WptVhszL880BChicLvDJ
j5AeXWkmYPOTZgpc1TGeL+bfpZj/m3ZkmWANWEl7gecEo5gO20Dmu2OugRFZhUap
K3sSx/IDqvxPUrkTVozU9h/MIxj5fNDWCVM/pa3PO2zbTGZ36n0HM8da0MxfCVy8
PJACrwTPvw0YIZZ+kvweh7bqFtII8RZhF8SSHooVrt1PpigYBGRHspfmIkN5eumF
IBkmzOfrf4MdkA/q+qQWnhVCyRjlp9lI+FgKkJtr0xIxFEzSlAjv0IGJZKxihx+R
2UsPNTLPazptEJ3Wxz5DhXyjPWooqKJOQWkrl4h7oDoR/ieGXTS4yrNAU0DgpAq3
3J9PKM4U0f+SrMspponXdFK2NyzcYJFE6U1MgS5hQl+QPeTp9IZXrsEBEFOF89Op
9BeRvqNby/M2VWWOUxEiUSdyHVo/xQ1TVhSa3e5ZVA4SJCIzL5apHpFqpH+S6z6V
hd//gd4ZjNzeK50CXULhIVipertbLKcWU/xt69M3X3+QX/qdwBzJajm0TKd5UrJo
Lg8Vx2BDuDscQCwKzsZgBE9nt6e5VQ7IKIvzGIXtAcSpjYOdoL45PhNhs8tOTaE2
xGy1J0fJvbtTZsYIYRJL2PklHyp3WcMtraWDKOHYbMdVZpaTPMCKfU4YbyjIhfu5
4in3sPkS3DKmoU4MdscqS4+JFot+W6sEu/M3EMkiuUAF/7R85tcz5pNacJwKVxrc
PcJ/NIYyYkPOGgJNzKwkyxv1naLnbmeDJSnJoCrJo/n7yhjwxys77MNiOuTYmYqW
C8vA9O5RCs4AkD3rW3F83UQmvdz9E94cXcnxKppP1dS7leya0wW1VUHaTpWffmSD
+nEBYVMGcIKjxMHE+ubRhBv7VDLkULZWCS4MD+IaSB9cYKsUebk5tKGj7QAD2yJl
LjU7UQilRvzXmgsqZlCyC9zZ25XPh0zRIG5j8HAvAmUHnL8F/q3sz25dZW8sCFFD
VlZVX5odNVQ/FNsSoQzQZhbH/grKX4Txk0of03GHgqEvzxxjaRUVXdNCEAO7qbv2
esdeXyM8RVo+aPQktIrwDe7sXWWr0/RPlgeVZU/3X8961AHKp3Uu2ml3JjhzHhZo
p+bVEKGG6GTKvE5Mio9VDlwBU9gguA86JkjqqMKMtyFBT5DVIyAtjM+SyJEZxLRH
wjhNq7PblB7NZXnM/mmK2bjfLJizRSSIAjwig2wJejQJoZAy3+xCB9JFlALd/1oB
/XIOtdA03gNBVIR+GqU/c/TmwbVNNXbdMpMaiKRXfeuXx4tuwFqwyy1sNGGmIaQe
dV2thz8eHquhwsjZp+pc4XF1efnALhndBqd1s+z4NOIqMl9pyKpg9ZXzoTpGEvRP
zlTiytFKc/eu9+2LCN9lpRXpXIcMg1n9ZecEZd9yZG2oVvR9c7HnutXuTiWyXown
2bzMYR3P2saG+8doHX7sGdQ36s6E6Ybe1Xzu+Vc0ds+hLjAaAkq8hWU7Ebei5fA8
Tr4yBZA308MQpI2KkoNWTugv0BJNkeWCcaQ9sdX6a32zSMGqyStmhTG0BdodMYSD
N4qFkX/aJIpd6KLt1aISc5vker+QFPI42dqrjU5YiC6hrlU7Ec3z2f4Me3q48zIw
HrdzlKlpuOECT2TSBcNMx0Culaj9kSDU8uiuT7+t7ry9ah9P7bZJ/gICFeCJOYhl
GfXUfn9Q0i71xR93yRJOzscp2LSAS33bQnQblRgGGZej3pd9zuH1kt9HbPL+/M0T
03Gvs2qvbrodHKaiI7u2+XeV1gepdvQTbGCMf0MFbOo9KTAdRbL4PzMSOZNcVqdO
yAmiM3+nl03FDPKqt1DwW6Js0lyPDxZHMd0OBNEVlnjrq6Zaaa55zm8D/1UIDMfe
yXoK8LlxFtt8ZbA4AHb6rhr7nADdUcACLqLVvTfgrvD6205IRn+XGUYqT8Lycee1
JOIYczuyeOiOd7ISTzS6E4w1pZvYiameJesMir9nkvujczKBhpsUtlCl+ZsUDXDe
Qo30LGj/a3g3da7FEzUNC5g2Ws1S170fWb1e6V6pVNV21Tb1Emci4b0MXlRQedOV
TKUMQl2WQ2EtBsETuGaeQNYkbiWBwYeeng2jg1Kv6fqTLPIuwWbDBsUY5IT90Bfk
8t/cXl2H2EKdoABa3wfKcQ9I0kmECpheNXaipejJr2nSMUU+8v37vFBtLVYPNozS
/CTLkZmSHQ1c2qyJU4Z3Qprd14foOOSmheuTMvYjHvW4D7IjU3R3tjGxyVriDjeK
EVT+5iKOipS+TTfGlRyaOwCY8xDOoGVbb7YCupPTsfQes8w2RI+mvyjssUTDc1Zm
4hBppUvqorNE8gBXB7ZiDlsnw2BuZYtizTj/zuzl33uxIoMGYq4ogHxbYX0XFc5K
oT/b9wYmSJkHvEQ41+syvfV9soO9GkkYqtA2KFm68LkfW/+j5TiLNSCUabDjE4Ha
fXSQVBt7DeMjvr9TsFkFBns2yfPk7ZisS+w6lyPyQYpJERLjATjEQTvjNkCo6Wh1
JQxd6v1XITzmDqJr/X6/+JO1XjA19ts/H13KvgnbRvLvI7DKyRlmXFWgg2UlOM5y
w1UK58RUeWyYux9adAky8ZC8wPJ2Wbz4j5rMBATQcrGmtiK9ef/pl1mOUkD/3sR8
EBbMyt3NFSbuyVeUThVv67Ax5guJBTEw4WoctWQ7FxeVqzDBEJBpipLUJYHiwHQD
/jzKCHqvgZ1nOnOqvGaW56df4b61/jSlDrxVb4L9JGyGOP1tfNKsPeiwnV+81NGI
eNr8zfhpM39GYHkjug8/SoUR1RXHLiogoT2hUBR6hR6kF8XIZlSpc1C/utfv7P2b
ov1zeVD6bzcYkGFEkPm9Ccy3usxlPPzlvfqOOv5FnYVjn37bAsc01Mw40g+y1egJ
NI0tpYXz7iZgWB7A5NYpu0VzzefphimknAcxnpFgIJsa3Gh0aJDwgSddCgSbIoGZ
wOKhwihsh8QCamHB52H61TUcnGddz12Cf9awOZ3FHnYnqUZ5F2m6GHuT15IQNwpw
nrf5PFTnWxaJUivt80CyN7jbVe5g+3SCkPtSgbF5H5H67RDoLMxIPo/+Nlt9DfFe
BExDGJJPD8gtOalstslU4MZKm0Szb5n8+yUOxOeT9aKNOwef/F/HZHP3884V0g9g
qawo59DxXf3SY2AdHj5ST4PhfdOHQsOiYtlHjclqqDN7c9NLM3Gl9nzW86srQkYs
nkejz9oooUiYqMvXJPsEpcQCDEXfDsva7I2cZOgrXrGp+tr0fj372Usg6HtUrgZa
BQCGauLwkAYoBDxKu7xQCb8cg/qSjURuu/LF9Zl6lz6UosakakHjilAIPV6/iEA7
VF9jz538BDJuVkURjuWyYVdxwqVqub3xtgCiW8hKk3YNHFIxQT4lvVSARmHRv42p
baNXjL0T61Sxa5XfVbmh0s0WlAGWhlnW1M2XJNYfWeL8TsWhaesXsiZa2Xi4GHU0
pfcjfnqE2xG+2EO63sR85mTl/bLHh0jFy5XmqAa1STibx19wVdj0x0LnfREbnLIF
oO/08Dmhk7aNlX9S9ghEUZduMvUjkqgqzGeQDtgxrspf8oTyzQMfrkNr5nB6osTO
YQD80UtcASvdT1KiJc9y5RNzLUnsiaY85yvmpimW2zwelLKWrFk2JEB9mI3QN9l+
J5alQx03z3/52R/yPaXCxWRIn8EN2NIHZMKirj+3mtgGXkHv3CZzHbwTUj/HXB9S
6RkcLG0KPjHheRqEMl8dHEhS11t9Y/8nOEBbbPg/9m0Lqv2svr4TYMYbmJYkxisA
bzUCKRkZxtqjqj2IvQzbLX3D06/3bvGb0uMIr/vJPOyaYz2tCwrQy5FbWoME6T5i
Cloc4426l/HLprPz0tTwfe6VvjhODm61uAtvnJzBRdA5npttmEjhfu/Pzb0fuwvF
+wuQG6mu3xLdS7sPdFcXzq83f446kU0YpBp1b/lHwKY/KhvTEI9KVRqf0HGt6/1+
Ggwaa0xce2hXgJcb7lqgvqw3SmNPrFErDVv+5/AqdimtFNOQJZBep4y8nDkn28RO
0MOpFvUtc+ghsNKnm6CrHpjcJCHnSOusAUnszp3HY5VBNzogObyCmIpqCbHLNN1q
mQ4EyR6pxe4QU273NSTeHaBO53MDt2q44uJFgbjFXyREDUQ3gp+LiGXiF9xF98NE
f5S2sWqz0exSbvgTbRaT89F+Nudp6qVS9SaTIzMAm3xgKFiXhQeIEnBnqJsdV6ju
EOjCDDCjhq5+WC2eHEvooTgmQFZMRWCbO9rtYhxkl484dvHlwm5MhgUxuYqq+7G+
CXDYMa4DpYlx3tkiSndDwhTqZ7YAG04pjMWKJn+OVEiToiu7KpYIuOPVrz251ZRd
b0IDkevrYMKsnLfStLUfVey8mWRSVHXggvX1YL+pR26HBVMbEPM2GrfhuRbopIEv
cWoUcr1+Ru3IAPb6YZcIeVIOLnIvLnrE/9ZD0/veB1DxecJcGvPExuZgXAfqoy1u
ewLTPq6VFCFZ1kx3f9Q/YGOWB8sjJMOLWooQxEPVq3AxsMmAUw1pcYtGNZ0+kZqL
pkCAF1UiXanKmHbOB/ramuu/cRbGAgwJgVzY2ill23zk+DJ04BmQsb4LEjHXhk+i
tcqe9A3YRj2y/McuZv3a7zzS/yoSU5nriy5tKLC3dKAljn7TmE5RXJW5f5A+q7Gt
ZhfbqfSVhKtNnUjWTKt+e87Ci5rcsZB42cuokPUrcJPbv6JvZN27cj9bgGx6aGep
cwTNTP8C+TtjznkonmZpdMi5XdH1fhTgOdWbCG1r6OdQ3NSodpCAZXEk0KrnVZzG
YSDSYI/x8DxxozULOvv8H8OnPgfIc8ngjN03cb9YmXz4njikivX6JN+m33nDF0ll
gZBcx6EHYmmnEyQpZr1fBwj282wfCletu0JAijvpPzik3WAtKM8wyyiSG22XCGi2
Fzf4nrNK/eoTdM4kmzGCjapABRYY4bc39vxw9PNv1hmPBBPGjYSy8GBhJK38E9C0
3Thigmfu746G9jXu5HEuroHIhy6BmEUmevTQE6chHKW9qFWn7ojLUclXeVKEynix
MsT+ZM39X9fjFx8aNkzqRYcXLvoZr4EdhPAUijP5U+rpElJ3ScYbqHoovOWD+ONQ
YaFYfNqHz8ZS6JoUPiR8t9YHKZ9dVfeOQ71xufEXtGvRYU3l04HRVndGRtycG4n1
64Zey5Bgo3k2ET+sxabSIdpcfv7zoV+cs/YuXkAb7ujZ3jC+raZyoUdmatnHld02
bVIm7ph1R7FYB65+QP0IUusoV3WYlcH0gNt0gdFYmxF9mHUU4s7Y4R+P8E/tLocI
q3Sf+2P72Aee+BleYJgTgPgwSMfpcyTjKrAOvp9lTTuDQvwON9TmhoNb/2F+0Vbf
jhkEZNr+x7mrJTX1iN+VBQtAKtcyAWraA0nFX9smLefaEeD1AVXl/3pWc2Cw6vtA
dKLOThRb7uHTLLs3GqbatcbHQruT8jQKulxChB+NL3EnZ22hUo6QQ254ng+w1sa3
Y+lr6pEk5Q+dAdFlvYORjj0MZex7AZwt8xkHIpcxal2GPFfGk5zTog5GDO2E1qiF
FMz3MTfmY6knwN3x9TzatoQFYaruRBkWgrYc4loc8+5AcOYAjoG3z0W+WZ+hzzLQ
6SoIlr0Ck0t1gd8jfY/1L2dX7V6HZ7hQ/dKJ4opFdsTs+84BncxQWw0qjbGEHtN3
UXzULNWJesbuSZh5mi22X4HAL2i7tRt5nLqsANOu9JM9dk7xvkm8d51IEBCEA7C0
bBLmUrPMCG2cLPXZSp3rYjoF5dB5erZZYxZgSc4HeUeNIjSgcwgv+3XZ+hpVEDPK
tk1qluEin4usJsUou/giOCkAcL9wZ446FBVUcFGeHO9RaJdqwjOvh/pvxnV5D5mT
ot1b8KqZY0wCfBoJs1UPp6KvvGrSj9HNKazdq8Dbbd/iRzuyMROlFB1urQknuHyj
PuuxymhOY0Ks+JiW6iPpIIriWm/+6UU1Atdog6nH0D7MggBn6wL3/fpEnflILnAx
4t6iIKGmZAapQzyVR/VyH9SB0y5/5BdEf0OQP7VQCnnx+2XaTrnoHIveKtYniXFF
JOTWe7BDXZt3fnwXb2TsW+oH/U+I2u7EQ/VvZaBV2yps1tYPB8BmctG+cG6b3lfI
jMshJhuxV8ep99MKCKN6Ia9tiZVB8Hfd0Lf7Eo8B/GCwztXA+VHg0Vt7wgFfedk+
1Lf4JecCDK2qSlwvU0p2E0u0nXAbDO0jnqQMQuS7njq+d18gX/srfa2Q23e88QZY
P9vOT9tmQZNQQ6UumBhZu9hBwJD7ROVivAlmGoBwbx48aIhRooynfk4UVGkYcfIg
s5peUk0dClfKqyLoXNn0vxeqoSwqRA+lZl2qAHniBa0iDa4+9r9nT1/fr5oACNU6
YPgHEJukbYCQr2FsktIbmlLAVsL7h+926GshE40DokYTXWP/APegtqbAONOsc4Sz
04d+ychOC2qISsktIAB9BN+9l+SfCzmVFaqlycIeF248JBfd2rzHnuluN4F7kimw
Y7R+aYQOYnbJtXr332UmRy2Q1yWNnrLjY3pbNmlV0Z7e8pu2UejDRyJS/nd6i0zl
VdJ8omepuRZ9rG4q1yQTnRizbVVsFqlrJTi23XJOjlCdg8mFdshRjsnafv++j+82
OFGo9eWebLcflc0Oco6zjvdozn0kDX2qERT2u8rblwa+OxHvBr5pRlKuOHosvobb
Ej9zAd/nSgud0CMioKVQDHFfPpGjTguDL/LBltXbU7SDAmlW0wza4GY/K4yiQR7d
j5yBjXrcSsHCklWSyhy6UEo1KiRfGIcweAJRUsZcWMwL7BRd3RYV1YEnBqm5mxoB
MwWMa9Becs3m5Ejgl4K+w6hVkk2yyJ5FLVE2ncupInm92c3BsH7behS9r70mfsru
gQbnIa0j3MY7HhuW0NkioaH0UMo2GA42NSI4L7kq85N6wJlmzVZcpkTOLuA2i7Mz
tL2lS5RenQEXSORPcU9zfoEFQxMuKBjFgrYKUKQWge8Q52ZYWDVtqjAYbVFKQQwt
MJhlQrUxa5c7WWGOGpOa5OzHF+Krrlx5Rope553myYw8SHklH/6iDp7gRd9BTYQt
Aj9dEJN1+q7gIYAmXNrxfLzs3ttz4ZPyA0+Wu1DHgmTmaSoyOeFevt7l3pYZ4/mq
S/IRm6HjlcTF2gXRpdaldkReC/yiHo0OFJhvoP5u4PpBsm1wI2OkxbQIbbUdnptu
e5CUJm4aVsgBbfvRjMsiNuB7G3VFvDfsfiuhvglhU3P73z5GXJRPWz0MvAPl+XaB
idOvKdvka7e/hwWl/gfOQYT/99NIVPwMzQKRp3aXgm+/FhwxDDqgPocT6tRqHL5T
skhUn/a4l1Naz2rekYe0RY8v/ym2buLDP2Pn7lpFXGtS1CKzfxtv0i3OPZDYou7i
9fCeHJra3GPFIAd3msLCpFy6r5vDOgpPa8zHOSFOi5aOSJ38aksupt5VLLKlHo8m
BXnMplNzis/uC5ZnkS4jEbOfGifbB58AAhFX4LG4WAZ6MLnwIMfKg/bKKVBBAh66
2dKu93g7EoEMFnvDQucyNjTW8txytUt8NGO/oPyZcUARPMkNsuSyv2ahPR2gAQxj
ii88BoY8x0rbeKh2hJL7LTdcbFNW6OZMB5Xv9EBjMnX86l6p2zkhfSthZtljfP9M
RwhiFh9jjfQHrDGduI565CejTph1wLDJBJiP0PRg7/W+V4p8ziBZ06HGTPhd30fC
ysZiWn7KZOeKB53mTANjxU/A7kiJrx5APxp6vI6GKfVUXko7znMLuuuZfraRCR9w
nUqd0Av0RiFsHkSs34jwIUz2Fo/C8UhrHC4SyNFippc70yKn+qincbOUhhZBYOLm
WWAy8hH1+qg88RpVN14TlJ793TEHzdD/DP+cCxlcQmPxBK+In6FMPjyIUl/ijP9F
kOebqft7lIVZ2L1KIJtORL74etsNVGV+uDma3kP12cr/TQIlb9WzFJFOk/isgAjf
g5LQhSv8JwM8hCeMPVynpIXWwIYT7th4qQaUdCTpsuEMb8kO0FMeT52urCLx5X67
XPNb8Y/NYMh5yL0AIWLvToW2Mz5LSfFOhWBgOjM60dAB57Pg/k5uRep+2ZMqgHBK
y1wM+Mjx4QZpz/63ujmw7dshm77fn1CTWHtWq1obGArQFMr8Bu0qqrrH6n6Ibp14
M4x1zRVwFmY/5YUJG3ENHMxRFWwbvv7bV9vDhXahlkjw5ZxvQEX7s2jgX6g7I/0M
I0HRZIz2DiNvI5T4tDtn2c3YupF200HrwKNnfzC0KGCjnnd6RY987MfLZ1eAqlJd
idJfukL978c6JBcAgQLTJB9n9BCavDoSxvnfOOwrjL7ibeUtuKudk795+PAePHgF
b2CIdzqfIPW/nxi5V/fs9HG/C9P3u560vbG7LzsEVG4hgQErLJ4z6UKAyg4XWAa0
+yefGT2VW50F3OryFMImlGY4inqm3jpayMc0jAF7L2CsPjeSPf0mRz1zgsb8btwn
QSwzp47/hr28qMbIH3iNtOTP49NtKC+rTjJJ3soToYljftU5Z6tukdYDWDOPWtIs
yXWKOVoyWT5hw0Fes0OSGkdT+Sun+9Kj7aHMod8LewBlacpplVwvnlqwTi5fnF57
unhrVCTs42mYLv9tcB+L1oxBowJgGhzYQWM39yKb42tSApJXMnhYgvQJGYZp6vB3
9uIy1sS7TpHI9Z/eLPcCzIHacnnPSN6wPdSWxlwO2tms6OEajCo8vAnXhkpfr6mI
u/fNMthPQWAXqOy7TlaARXwjEzxqj7YeG54kHKPGXRoMakKCpvrxolBg0/RlmWjl
JWJxiUCuaZ8raOQG+hw6mhB7mTVLgJ+LsK0yB7vH4sPfTi2vM4xlB/gE/8YdHi7X
Clrqc2BRM/eEIV4sS2I/pwcv4zTei18iyXGr40U7N63OsT2x6P4qAiFrqY8t5YEU
ecMshSqa+cleWJ4Q9/yRqM6TVz7yz6w9UrFgyjGDLo+mFbuILD6iLictyJD6CUaS
4sIaCBfm4QfE8q3582EeSHkVSLwIXnOjkT+7I/UikNPkSNjL8aybsmLWePJfOGa4
EgNiwiJOoRD24jZz4jCVrv326OPySO2H/BKhV/mcFZ+PjVaUsy7nA2YOffRnEe+v
HJIa8fzCboJgWY+YjEhm9nTiqRNMuQ/1hmH5iSKl3NmQdnxNVQl/4Kgd7XNAMFrN
UU+d7uxnNsHDJaUquk8IlYbKbWc250825z8R6naJpCNyZwIdtGh0RqV34pTqrH4V
POE63ekoVxi9lP0agBkb4qjk98/JLWmYjQZUFOeNk4h0s+SVe3zp0AL6npflR5dF
yAHyZSlNSWw5o/yg0/asE8BHXCVFsz2u/dmH1UiJAR8i8Bi9tKLkWaU7FHafmbj3
PSQXr/6M8CTBtjKIotbs4Fi6yLsaTU9arLo/6owXPsqS9OPvchpu25KDT22bwEex
wNQjLwosrxdsoNyGfEtqHeMJlhpZJtzLKqQud8blRvWSmQUVk8TXBtN534Y8EAm/
l7KUpz+zzlnMBWv2ETlaDUNqJ0D7n59hS8mjJyT+kZULa4d3HD3Mnvz5Yd6k2idf
CRmZzlmnWSqJG/PXBCZoqUI3T5o8wL2CGU4lLhztJZIMOUv62VQdTRXBNW4GSE66
KlDQp2S478sPb8tDxgYfr9+n1lFfq1goI8GCzg9374vPQRBLYQqbH2o91+48GIlZ
jYF+DiqvjFCdAXZw5DeQJbNtgWa5thmFucM16IaXUwju72nHjYCXUVsUj1hLdFZm
xXF5DKmnW3FLlz0UO/pZM/WitP67I8QlxgZdhb5v+L5G6v6UcRH9E0Pz3ONhnlXh
ZuqwdgkKk+j5s59C/jWHkO9zKdE/Z3L+aa+8P7+A8cw3BCypw9ITx8VuL1ffjeVJ
5R3G28pL/OarlS8+xnFTrScd6PEZa2+4FAY1cnGN8mlZ3t6+1X0Gk+Y+SojXTvwx
ciDdWpprYYqHdbIps5v7/l0JIGn82+v61y6SvEjrGoBIWFkX1lrPTMsoYIwNB3x1
akd55vNaehiNdwByHSfv+sQdiDY4vcNdh+LD34AZcz3DYbYKpvLKKCic+7GLq115
RNBaAOXoZ3oxH63grUU5GDf/DUZcOTyZzRMS21JTBF9COwmcfUDAsAXWktRtRU1/
slk7khPccquhRYgiKTypkYltSGHGzhBbrDTgTJ5BAuBY4IO3LcLSR1QEef8pnCtf
nfbdM0rOoL0Ig2aBYi2qAuCcNtZ0ph64EMOIha2pmm/2OoIqsCkLRqJYvxdIZW/N
TlisbJhsToQXosMpfoRHHlJUW6tXKW1Jz06dsuyUJpnk/l7PS827blq+DU+rkDNy
2jZuozJa2V5N5+zROT+ETzK6lG8JAiZDUVsOk6VycXHbkB/lbve/hacYi5vLA1LV
I3yXRTYnkWyv+AQ1HoauCRquddQbsHk5ACeOx07/Xo4erZ0yI82WE4aLPBZ0xozt
tQ2/MBfT7n2/9kXe02QJF4VdV3AaLtCwgnXMrQhSrhGZplVJs4sgnYy2+LXqLbB4
6clGt9sryfM9T3X/dVXpDCA1UL3xG5X2LMd4EZGbVJ6djlqQ7H4ypfusfQO+gKTX
5zRUiSR0gwmBvo2Q1fSUd+3FtFSZJ1qsRjOK3HW4vs5CJQlCpuvOgL5fGPIqEsOH
640bcUIn8s5IJEHgmtd1x0oUCXwR1aZgtUvfSXAVaEAMS9fyGqppLnVwz/3hq5pF
dy7uOdg6vS7Dwt72RmNwifGfoyg3ns5ndKO42eccDNILK/sbre3lkQ9UUJQ8yKlj
pfFQL8x0IOOpPx3UxbMI2OWM9TgFBdYSqhs/5hnGit/Ovi+x3IrT3gUMQzBDaDC+
A33PBV7GQLBVAwzfUZcMj+tmITiwctCCCR+DYezZ+6l43CbjmTmJE7oTM9hmuO/2
jgO2vARrtzQzaY3xIdn9sRC03Otfk/oqAaJYm+wXPz7QEvbs0G4NuVBuNt84ytFQ
FUdw2UC1Tl1TDkHMe+j4RWqQBUy2cajOjaJdcRgaYodmyOOwFjrl4VW4N4o8SsoV
VIVI1PhhIK2IATEDpiSzbhfVTXq4oIL1FaQQRWIbNsPLawEoAZPIMd1LpHPqP1y8
zbcE/br7wcaRj4MpD3IyRFA+V3gi5k/3YBB+OrOnd/5IqrVTf4ZDDtzqhjyGE6Jq
7u2kl+SuiWaMYLCeypEqaiN/IQqs11bpB1um9BdrOrucOWO21VnrdhQQZxrsgxpz
EmUTgCZFm3bAN2jfXnaTO1DcGLQpgI1HtuuyVDSDhuvowCrjeGQTW7FrVJzahdIG
l2hGahNb4JZ6tzb/GLnJy3CYWKWLCnKK1/6j254K/NaiYLGsJUu5V/Ryo++mBkvZ
YKnk2Nj6xGu+DvfXz/wYp7PLdU6a9jvIPS21Pi3lc9eZbJsMizs7et91GeiY0+Am
6hcgufAyiX4FeKKdR3zN23w3pf5jcUJjktREYyiqWhxuIq5pAmsqRaWWkC+nm7PV
eGI0GaM6bcQnB1kDKdhkylaOow3eLm8aXKCSfMQoVUMhOIsYWlK04ruMKEOUj5O3
Y/tUs+CrIWHrJk8q2aUedfw89R9wX8AfV9S0gAJsF6YRRHCTnya2+mCzthxBPrj4
pTgwPDY7KmYikYk//gDaOeM9zeurZ6CAprwn5xeELTYRE7HOt3ShVinUUV/ApinY
K5SxZQ6+FAgteQK8bXMWjn6xXkkkTiviPZM++6/wh0gIubepjrTsChUIcXy24e7B
X849gffA6OQKsZccQMLzL6gdc9i3hiy7NDSpK9zQkzKzG/c7Z+XKGzxt5L5sBdGY
Zkvat8zR1LNQhRSrOgF3Fq9oYRDk9RKo0RLmilgQq9c7BH1JaIGOE9y46j1Mg5gS
8f82g8T+3wDhtLIDVrZeObnaiS6Ci28wNHiw4p6rUzQWLiOBsx20BTeUF7GKXXbB
R2mPxWJ7Cjk/2vQHMjDQn/Thu4DudvRXauYgSMVjs7pn2FuX4O+KN6aeTbkdG/Lb
hUiUzbza0G0Ima9Y08iHg42lAhy/D4x+QOGgieUzcTBUm6Cj/uOfgYuvGsQfoNvO
4eWxII118HJtVAb2RVNbsjBvFjU9WfZT+PdXs3MLD4sUIcWf6sKg3DS0ontYoHtM
F3Gf7TUPMKFfGScnMf8fKeJRZUSE8pFFGzP+6oKALhssudAkkMn/oGnxajmpOj65
fVd32G17LNs2r9hfV90/CZD22CTG0FvgjOEArqezWc1RbQrGsQdPMWE84M3EU/oc
cdVzCOq1ZXXTLmTvTNLrvie5Z0/Udgw0TgT40KN/c0T02EJ0vV9ZtoaKTRVDFr1F
B9Kg70BIlfu7gCJR/aB1Mi1BvDUutkVSQRdo2R3WtXzCuJBBtGLHgP/SGhGmBIZX
DlDtUXLjYHHc0EGUVmEYIZ6CHmk5Jnl7rN0hk86vgM1BHi8qAUpNM7oli6RZeloA
hRsTMZUtDHMyrTk/wh/3QweBDDP7IsvF+XH9G3ERWzVBflWs1A7p0tODZN40oUfu
zlo/5bW38jOlgfl4hfLaD9Fsh/WI3YGFy4DJboW73lcCt8RMPVh2y3nuKjPNKUJW
3PjoLKQqfL0RR0XjcRZ/99c71a/bwGNEn09SxyZY5dwkMH8Jv9jZrpUMg3/gC0gT
18LoKBu4ovWaKApvrmv2XgEhgBBg9t6T7+HqOC/BQSCFK7Ji7A0Gz5D7Tutc0aHp
Umuhue13DfE/8v3O6sXoNfGoXSWFnJXA6lKHikJoNFDVlpizOYtlGj1+dxT7qPwT
ihqbrFtsSN+0gJe0Iul6b8w5buhHT0Vj4s4a+MzjDMYudnfK2g2t2tTslvl+2cHE
AnmYgswODQRxB/tWQE0OvxYaefkzUh3u7oUZK5SYYyUYWMAVsOg8MBmKBLUoJXX9
/6Zat/2VR5LL9kny2a/ogcZhD5wmehnm1PdHl0SdGG67Cw1e1gQUAtEIU8TfA5Ui
c5NpIpww/8OYKp8JV/VAiMj5+v24iDeAJRvj5a2VDkMO/uIoyjgYv23xZvtbuSnU
4Qxdb2QPfeVAeZhtj6I8qB6vRzKLaCSWctSpKXrEi7rghrEnnyEQk6evUVfwsK4h
yvQYAKd8CiF7oJezQWr0HMUGI7QNdGX2NJV62VPcaoOtNLvrva61QtdVVBFHLy7c
6in2Z5l4h9yDDKpcql4G5GzQ6ZjL/d8ly5tmTd7da2FjlHNSWMOcYnfIkxRNBUsD
gpV9eM1nESvSGtfUmGLksXkddmv5oN8IdVnSsIO1N96+7/g9KFJXrVD0BrblUNni
wUTZ/Co47nkT/zb54Sfa1NuVsqHJqSYiXVGtyJCfQdyel6sLsmftZ/zYmLvAAzt0
0LFVyGyoY0Ll3gxbvKmT8jmys1KCfSHWk4AytNERrhAljHm5W8OELOb+muP9l1nX
8y91cu25G3ALXRj6ut8kCgIHfdEYpTcTZNiDp1yGku4X7tTbLkHn0UqRfmQT0ydt
0U0VaF9D6AxMd/z5ivCG0n7t3jZll/T8fTt72FCQSrq0CosmexW7mMJNvBbtPhe2
k2l37EiNQTkRZQlVN9A+9SYM65J6nrPmgaaiIeJKNH6FbpqLLmIpIiqWgUEVSqhw
OjFszMhnfg4yBrcv4kwC/mO2nGVKYBvM8MrQ9H2n9q24zT0Lm8iNKiBRqLDo8DM5
yMpXgiAvfKTr36vbSTkUcLD7CIZXrC9orvHk5e7PWHhgCBzYmP4UX+mAm5hg+7fY
cnluJVj2ZoRYWXTx0Vgim84sMlEzG5cvwfuEimlnhpuGh0w1+/UFAcBwd02B8cYc
6tgqQrN67owRhNDhQSCkPxMOdTWWqDf85VITJK7cPBRqPPMNU1udDtfb0MpbA4c7
5MrjlZ2PHh61hDkENGbob29nDuV1ycAVBGcW0Xo7xboPF9IT8T0vfbc7FP64VYUz
aWvZOC/WPDeqNALYQmKov+IpgQsDYgGPac8ZMpC6S28sm5fWyKLw25nabL3mIrTm
zJfMFDtp58NOptYdBrkhr1j7oIeVVca5VZfFY1ZC0U2hqZ+5OJEL0utGokSA9r1b
so+c0FQqLoWry5Wg5FOlvq+wa9kTh64/EKmEh6x1+U8vL/r8E5i84dtBuJeoqoeu
gzMoKqLizbOkKgT+viRgfyBK39b5BDChBSWZaiNnGMqP9AZcI8YMpnJBYykTHl9c
IR3lrtfesbVr0P8kEHAfLpmVleFa9mBkFJQyNHxsAtaRjrrEDjy6btS164k+ur/8
TmVm9yDQ2z+aSnP1s8DKbDd/445BbFQE4XTcOcM+Jbf0Z1/iWzZ0pc1dtvqC89vc
QrbQuI5Wz761Gzvz5f8yQYxYYTtR7SDxbdBjNH04jvz/QM8JKUdV0iRPAS1WnZ41
Ch5mTuVrmtDClgOkgHSDpUQ3KF6khzsggw50ZImp82Yv8ZwpAtL9KBAqMmPTsIoN
fRrD9eyuxgelVLsUaFWUYFnJrZ3os/XujGI/2oHR3Fvho/gfICGthFGryHYh4zRM
3W3zh0HwHFPFSICA8wdQS4Fqpa092iElxXAT/Rah3LFYQC2zeIs2TI0dImEEBIZk
/rtvVD45QIKCSr3M9KfR02nlsJ+Mol0Ng0q3IdJjnUgGeZo+F9DdT0MxxyQSZG8s
xamcjcQvGWses0wvOfO4NmK5QA/jSnrHTwXD8Xlq6AtUE2JL8zw0NQkNSUeIU+Lg
PB1ecTZmLKQA8aMG7V5eQeHttv36xroHYGtx9rRgAm+vtYvtDHRwsmwbyEmtiJM6
UygJ0CV4h49FEf7NIY4c3Hs7esWfsa7T/jmr88km/vLnpD9Jgf4XTWNe6+EcXZrD
H9+YzMuNr0iVEbs9bbh9JF17pVCl9G2FJN+d9QXq+pCWA2LhEsgnjH6KBPgK8EsD
QryKxyFNKaoOTY7r2DDBppAJJvbPp93L2Go44IlxHSPaHeZVIC8mkA89WU925Q1k
NvidXHGQA5FC//VAN2vE7IUwLZ7aHwSTypvCJH3GMp2JUVJRmo2c8zm2lzfeKIKI
6QVih1NvwQwLP9h9Y93UJEecHja6yTA21AadjzLXA2To12iWSo8b53fznFJGj5m/
6p1IELwmW7VnJR7yEChcpOzVB6ynr2OSdEDiORR7a6Miq2X4laLljr4VvIiMLizZ
0sL401VqsuWdivUpQJeL4Z03AovCB0UTYqkjgmVKnJWuxQiiLZaKlGs8mKny3lb4
5IQxQN3llKP88ehe+eGoHhg7uBorqKNNuT0jBfcaubh4X/06VEOzZuGgwcD3BLak
qCKJyTJeR54ApQDAhbIU89HhRbPTVCA+DRabex8vUTNxm57NODApbAtEYGIJ292E
mJr2Johdpn2y6l5EEPeMvD31EsStSDI8+mt02BLdoq5HNVUExM+3OR+0wI4GMB5f
m4AkMzIVFyc1lgCfIKIMESDI9xWWfUN9qz4sOHRV4OYCmUGx/SWeMq9pTVdslHkB
JubMct3a95voqvEx8/WNffRhQWAct2fVdZNk9hl5x+1vjcMMbvTmu1Tlh2AAsRlO
4ZJUm7n/5O4IQ5FAMaIUmMvCYAmVj3461RyICMtL7ARtyZ3XVppsC2NLy76bCaXm
44eapebcE+SzYxumwJj79ca1IJT4aXZi1iRwh/Ui5VWHBkSVEi8qYB+g8OOJ79f4
KsMb8rcYtyWjU3+jHVtfC+CmGPvLPcal5QHSeBgRsV1+Uc7uzULXAPsp/UX5/YBu
dHxV3OkVO/72BFBIT+UnlDetc5VrhFkV4aBrhehnFSSO4y0NeIWAPlW6p+gKFt0q
YsjuTFn1llZLiiJE+P2hItElbFpYHfmIZ8uIiTPI2f+I6EvPy4m89sj4ayG1zEOL
4Q7simY/7SDe7dXSfHixKvVIIeTBNcPuKJk6YdQ2REB/ZHcJwVjIGzB/3hpi4Mny
WJE/zRjKQTPcly4uFlT3t9yE9oYwntfMqz5j9CwuX+0c3H2GL5fLfCLFD4J595Hv
Thmw1fDB30ww11OvOUBBvknnjfJ++GK1bxL8Y4rlMTfPvr169vrNirT0DFA07E01
a30waddV4PXjHFNI/ALvyavLhJDc5bUZ1ljjo2lLu/kpjTVC/VmKBNpCjVzsMY1Y
sq9szPheZbT0UtJ4pPyx+ICKWJ1IFYSVPU32rIDYbkZl+qM/Za8qLX7XiSielV/X
pKEz/BiIovLNYdfYJlz7+J2zbr3j+je7bLY20QqZrrsWtmTB3f2KIt6MwlIbEalH
8FnPCLz/KLk94F6BK2gphdTTHxzEFuecf+xLmQA4y4b31mV21FVe/jOyNOH8bWct
5cxnLTq8b/jQi0pLCA0UZF17QlxjUGJjtSiUBXdtIIRztKWywRbJBNmgf3XsICI3
a2xQLNh88CnEWlrxDTMGGkg6V1Tu5ok2wGJ/mPv9U3sijQZa6Tk+uyRrNtVbEbS1
vQXYG2495vItgekKRkqq4Zo8JhBgG5phqltIrGMh1vucTZhoMlAHFRd2WDaO77YV
N0wHwdZibuQybIuOl36Metd/6DlkiP8eWoGD1P7o9XwbTPtzvg3TbYGNAWcprhTt
hmG2uegA6HCxaqCSJkXREWP5Z85oStEK3iD/AY/z8cKNu1OkU9V0kikjV9L+8G1n
QIbgXGpd5t5qIImNr4MH+CRgbIWOHceOukmb/1fK7dgOCW3wXriCN2xCSckVrvY2
KkLcoz38HnuFUPt+KSsjC2F69ccT34KWIQS28wu0FCd0LTf+Aa6TLwlzG0FZ1Z0K
V+ROyzfitKnAwz5ROM1o693K7guBBYesQx0E3jXyY+tHexog5l4IZA/qmKtfa4t8
HoQzpuLKuvjddsObNrLTNuQzlHJswaJc+fg2cTMgzLiDcHs0zqDQW1Ly3uRdhVuM
k3wNzunJc2ps71ng8gtDzwFm/cWpwIOt4Uk4BFzIos/Jq0K0LcinQ/qyvEw86RUq
XaHBSKRnCKuvzRdJmgoTBpmwdcjpLOf1mAhYq2mZQA6OdPQUe8ExuwCQBf6AKv3j
NzYdI4iNdWTUmvVHg2lU5q5g7wEL3WfxK4udtQ/WS0ciFR9TJ3JJKPheUQts3s7M
dUAP0BZi6gbeOF8p05hxrOxbtObFXX5SWTwmwPShpfm1FEzzkGBLtGVNYIaxkRhS
kmVtWWToP/ua1JJ+dbL7PL0wbPSMnb09NY5cITUloL2XUfII2NWY3frXieUPTJ6B
qa5tYrFMNLSZL5MFZDWDGRxZTkEUPu5Y2Ff+r7Kvv/ULlaTssch+4MxGcVAWyVdA
07ungl9QPCi3nclIsLFcDI/q3jPAllHEHhmV1iNFZs2Zzyyh7Prw6lTXj7T6HXeA
9ZvL4I0i/VWiQb19uvJLDCIG1nSXCtWe1tBpUs+q8pIB8mL2IPc4E1OOklhG3ozw
YdFAfT1R6uinBYXjb+wvsnoK6XK7q0x1HKNdxgEmRupwSCN8uNqR+liCzsSf5sWq
STPEPENcFqmtbAICq5A3Fe2FwlnRF/Ckaw9nms4OIUG9P67bVQ+vwIIhSFlFLZxP
euEJg732hyNWr9F8RhFUSxOzBP7EObHW9Y6C/bCl6bfqZ5IdpL/tfEFwANSzz+oa
X7BoZp6jpiNB2Hsntho9c7h/dT5HoD9edujbLm8Y9yiyF7ci0NBakxKYj4+8w5iu
3l/xdJrOk4492siIwpQN/nkxvOgktxbO2hnTGr17J/LMkmuwubwuOWUDn+uyLzOW
iTap7TWQtsPz+ToeZjaGDaC5aud7Ym/JrSkvfYo3yPdjei1pL2LOgtnPg0dSE4Qb
R0i7yuwoclH3cOUFRftYlARTwbNL21uCMb22Ks1zfsNRWhbi1VSHzRozzcMMBPQc
ahrz5wRncqwnuyVP0n/oSr/hGuBR93n5Vowx2cpOD1HdkP0qgMvHiUywgMG+J7YC
FgyIZf3p+EOGH0a9watltqzxNmxilTMYck+URVN+Aq3XAs4MfJTuAf2PZmF2w4kz
sHEEbKMOs2Gfwc2GICtFBnvcZxuKqJcWrodeWTYeUmzqAgsItac/84lkPw4E7cXQ
`protect END_PROTECTED
