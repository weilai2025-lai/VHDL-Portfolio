`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRnXywyI3SgLvoStDgSLx6JviPO58vlYKpxGBEDqsbuaKjLIJ2OKQYn5Fqwdjj15
eKq+TM+ORqhODHK7kSIIrhENqYwnq1aDGp37XAe9Zcr//pGs3FHIVnpD6MEzv3kr
UeGmgZ4gfnbS531ftf9sZF2NBKH3EUvEhG8CYyVnKBE=
`protect END_PROTECTED
