`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpkLayK/oaE3yPDkiZiUnD1ph5JSTLCe27S4a2ohGY1JQfyhQGHeRh72/L6V4BPn
cjWdaWHlUJGbsmc2BLnrZQS7ZZnSviA9TY2Dtzp9HubQTFRj+3VYMj86LygNkBaf
CqJB5O+wOhVdjBibAjOZTfeaAKRTMSoAXiMlfb+nojsSq3if3dlQYZqe1J7ZnC4z
WpC32v9Nd/sq+FY6+R227cljl4sC7DOiJjkmnl1UfY7JZFwbP9hmomqYJ4QSIpJG
b8ObpGlsMxxF59b5Q+2L6d9YsR6LIQYUb6hAdzRQUL3d0cTawMgpqr496y48/LXS
FXkytnZKmYVwW4RgIOs27ii2NETbg/izW8YTRqCzxKdfvi7nTFptququDETBfIl2
iFd1lAj9NdfCE54ZezvsHu/G4RyAlDAvD39F0Ajdngx0Esz1d7gsfVojyJ4kbR58
VxErWgTmHsmlFTBfwp7a1vG6XxnlBa+zTabiU7oJnI2zYtkxMBv0Tz5kELgUFTII
oUnSf7l4Juah0Zfy7T4wX5cL6WJd0c182qkTKsB14RQTTzDd65o0FC+TW4U/qwMa
+BR5pAAsGgZq/PVsoQQfPXekxqpfFoWD11Ns9wJ8a1eEHDhGR1zetujoahIZo/Le
SzZw+NZyH4pyDvu6t3keu9CHKQzes50bhr7fzFL5xedX5nMF2oiVDCSOWtPaGIJK
5xkuQsN7G7y8AvUQNsnBJTmjgiJ+hPQHjV/3nhLpGgm99qR2AKN1jleKyc04bCQw
dtDylX+D3vdrcklaaNdMlitMLsAV2XmuOPFQQkVnieIyu+cDJFsHbzmBi3tFG3Yn
BsbBHMekX+zHWHH3u+GNAW0yqt+5YSd7DHw6m5hXMyiej5IlOK2wj+jV2yES4C5y
alWjABgdt4Jxu01oFPQW+KAwrIXD/miS+tdcnCkjAlYdi/kmlVvL31so98xCWRyQ
ZNySK5rJtS0ExfJey6x1p/kqpDidKqHpL30z4yk/pN59sui/B/JYfxnb/eoSTDBM
0CGdZGrEYNsDErpJtkxoy+eE6z+PjETrgqyzyBnQZVhnl+nx5K4kf5Kfri2ITY5a
ESTUh8fCa09/Gh0WmsvrhrRU5yUQEgUUJWV9/eTwartT2X+DDCjQ+IwSlYUefJ3n
f3SauLuPm+ggB3DGOPBW83XZYZ3Qxi3Cu+kwJfLRV0JGrIasccEdtR2DhJy5Ngcp
NCzvoFJ7V56l3GcWCKlMJXcExpMxPYWyOeCNb5W818dszNPs0V7kkkZAM0v0dmEl
8URw1vl96WTBk03cUxd0Xoh5uA2PQcqwD5cDvumX9EGyG2TgJwI/V0UUKtWSZsNP
VSg41P4SM1aU0IkgAmB4OuZUvkFtWVzM3tKrz/0U6+kQS+rlJnYBC4CsxWd8ciMy
jocltvAqbIDT2ti0tMHYEkO1c0rf3PjJYVK4IrQf8LGvy8uLhXkfC81bNeaaPq4C
OZsDGC1+dz/pm3qbowGbpd81DsUTrkfFywvzXayKrhh4lFGkfcC6XVS4iofo8pdq
W68sMtaEeWs1p36yYFJ5aDs3okGKywHDu6kEBARJIb6HlC5h9g2JRNCHZrOoeEc1
dFTg8GIfNEGCqSJLgWTjXMIOq1Xcf50qV3DM1PeUCH1vfIq3IBNN4tNU0TzaYyU1
BZeRhbK0xXgJDxoS/PukPRLn9wAczHFdBJqO0cMGBX3IZTcXyxJy5xnv234vu3iH
kUgcjPde54u7AC5mrPlNcvw4Mp5nd4YiS5CEy08uqdT3olatg39BRfdCtfzudkPv
7P1xcIAExXfnWHjrLzF3qneLSl9mnm7X4N6ZKqDI0nu7Vn154pxMWMjy4l2a3llw
NvvJJOSUxyr0FO5TjdbN9DecKliFO/6xnXB3VG1RJgb4T+EE7BlBYONMctpQsr2o
2PyUI8/foC55KEF+s+CkwTHzkofdtgW3Ot3ox6DYqIF/KfipCKKNDK+TiiVrec+m
tWgCDn2JVxBwmN/LIPqaAXT1PV3bgz+UofNTZODKDZhTYzI2UzhwV+bmVJ1QHqbl
0PXjq/Zrf6BIvnjbyl+WYdvyY4MdEJl76cZMtYYFSPxV2UlurZ0yncSb9+bLKKkI
zyM8er2DpJfdHKAnXW6oWUceT7SaN5KNRKL63QWEEtpVybdvbidNlM1gh4sEobN1
zNTZbmmMWqxmQoiCW5+srJb3cjjuY//4Gia6qpaG9QvnLHwA0O6930CzrUDsunUt
p8qgHiveE96T0no6ClrtkBlSSRb9/VzuGFRX+zVc4sQ0JVUeehNb+GTzuf6XC29U
KeSVclOZtOa/ulA0wdh+8JRU5ktPsTRYsJTeAkaszt17FOx/GOVkXIEEblaD9Jjw
lTMLCDipK6hQ8MQVlpBmuYVXSRRDqDfdX0vc9jvyGJ2GhQOrh6iOFhFlNvEhJ5RC
PyOSTgl7j30K1CcUypt7e8ZL74sIapncF263JHeV1IwDkapCz6cfqpAsgJq+KHHs
aD55kQ+mvOm6ZNYKfFOeXT4dswcyovSlKHlBNE0UupheoYO3hM3M+Ee2XbZghMYM
kTsD6HfAFRIpiy3VV4Tf+sTSPHqEM8/0NNMUBPRogxwBG0W3/SjVIF+Eaa3wnYyo
GC1jDuX2uy3SYdwZLD2l55z6YLRD4VvyoGNMkU8RP8Eh0UgvzjDK2m3MK893f9I+
xtgVhbIZbJ4O6C83Xni+QbhjjGyQI4LYfk6if6rSvo6SdwtZ2WdWtZed7JABEx1O
hFE7uGhO/mSXy/syGl2tu91w4hV7dmVdem7kpPYYP/053OpJ00vMOv4e1HGITIL3
AbYrq6dMDuvFKFnqREhIIZTvn+rwMW2Nbga4gJkTlCCTQmHwZtbnZd/zVoz4zUd1
H/BKJxlRNnAGCjD7fvLGE2/Yb+Pl7zM0Yr1w8eORM3tK27hbUl52tXt7Z+u0qFCk
q8XQqvRQ3s3K0G60n10h85+TPAxoEvADa2nWTCLSoULBP9mEubDvoFCpD4z3u0MW
5vUCOFvUlIhdqMTNEtlmVuv+ed/8RAo9oeu4bNPbsCZlOVIbhyqK1ln8QLC1zB/k
JfL3mWB+Uy+haByUa3/kfU3eIbsT5YOMjFdCsFXpR+hlGTZkg1U1gKlJ1ApMF8qJ
dLBg0kHc92wbFdBH1rzeqNxkXCZ4e7q1L/HAFcZpMF3xJq1rUYIODL6jfIrzEbsv
D8pU9HAaCeB/o6FHK01vKJk7bhYbvrxdaMvPK7frm7JA+ylS6r+GI9yFK0J1QglB
YpANJLduwp99ep1Asv7Wk5YfVL7vO8akKC0Mix2TbnLT4w7+mJcug83taRgOesfd
ECio6LzpPQJajXzbISWQ+xzvHZdoRdNEbmrD5bpcOHwipzi6wo36zaziGV+88qHg
HeMfqMyEbAjgmQ+0aZaTq2u/AhkpczXE5oI889+2WLqtJSznj3XD+CoPCbfn3go6
wAlDYPlQBJfpAU0duhB2JFdN0E471gX3EwTgkbHeI1f1zG4yMgfCt1dr7X53K2nJ
ighvnihVfaUe7kn+5iDvqu1B8UoosqxTXy1KE/QtUqUZ1PqPAigJZTTlZAjswhHT
U3bhPbfOLf5KlRBXaHmqiHD2blHBMfBBQDp0N/QdARU1buz3N1eBaubkN62zu7Rm
nUT7faHApQecR0d+DB2WUN6hTvRQPNYvUfq/NUrMiGJbCr3a1cQkd0ksdjC++MUC
Bo5jPRo+cw9g+pLjOFPkV7b+a+wGY48cSi3QeYtrXtSCvmI0/7JikCpIQDrm72I2
taJNUAt9u7XFWssaec1fQ4xGSmEB75P9dywF2lUg8j83UNmdNa4GxTgEJcKCJSpC
CFi6/GAUcqX02FN0pL2Xo0jPadjCzq+/pddiJzR31qT5/IQWQv77L2kEYvtY+C4P
fYT03DGOy6CUYohDJP9UR0xrdGiQ+FDiK9Jn4pX0+yNjQOj5AlISbAkxKh4fRk5K
MDbZrEYS+yHxuPoL6HSDgA94hquH4smj6cXewmgsTmLP431T1hZAq9M11dDs5AhW
Xn6bROw8Xkyt24gm8RozbTPwgIEjmBZ1r3PFHbYn2bC5Ao/j2XlyxhVH6yYIJISg
s/0T7t98uNv0aVlNhTbfDNis3TIAzancIEUGTgGTF79rJuiIbkBmpihZj1Ie/D+D
fVsnguAbfkyZ+rqjAq9pCOEZ8ZpBrKYyZSEvw6pEa3Mye58JN7b+0lcXhCh2Dqm5
os1XtxmrZSmetVY39+AQuR4UJpUENxWbQljDwqh0O5ejR5jRnTzAqNGCvjIVeEcS
/7PXEtAsllNMwr5iWQrrt+V/bQ1nCpFykWv8rlhg+5VVicLfcAMDhyRb+GEbJuRA
Je2DOTj6Cj7CkP0n/hvgCv8j9dqY1Kur863EqobhO16N/BXOqlebIDTWL+cFlx/B
O6a84TBIKAA8bypphtlCtSRuaUYMo8TbxBOJzRK7zyoqby3aYmU9cKRTUnSBEccQ
cbA2yfiN7gLBOcPhpDdvhZx6TSV0LRwM3gv+sYaSGNYAgO+ZuWdR+O5UmGj8Qw5W
QGxrDCCkv72wgAo/rP0yJOl6nlNfRA8M4hjSyKEnOqR3n1bpNHcBHErxg1vntWFE
vVX6LIpTmdH9A/pHxaJ0uw9l7uuoe6qOHDBODddJHduK/Fubb2DmljKhejZxtcMw
KGNbucp6A8ILQB8dTxaVTVED+DNJ+uZN3b4Z9jzHsTq0xmB7fT+Ns9Mq68CjQB7j
yTTLfwIG2JvGZFGwXIBC7XVvxLlAFIYY7fd2rNVYufFO4+a48viJ2JPzttonY6VX
SHzoUJWFGwaSw4HtQevbkqbyAMpa5RUaak4V+ek0zWcNGDl3EE34wzV6mbiYaKGL
HsgaUphnbkJLgGY/N+UdQ8zUmFzDmjP+2RZ+ephFCr5OpB1YQa6ijC5TY2N65Q7c
zmzbW6A+lirNuxRzvh2wlC++xeMxct9xozo5/JPEj3atzxUpvUb3kIDdURATQfRE
DpfT0UVMd4vYgKEPMXUDGbX5AYrnOr7M5xeQ0fIxq8tkrhvH6M58mVj62Iw5cMO9
uLMy2Qk4WmFP2/a8RnhPq7jKEGln1ro7rJbDw65XEa/OMCLFIsc59Npg07SMjGGc
rWq4TD9LK7Vag6ioC9Gv93zNk0umRACwt4Pe93N35HayrSrBidHNp77WKLU+xz4T
1SmpiMOGTpV/8gzq96D5Xltikm1gPbdZxj+l6OGbFvioAZmEPCgPeyubq+QE6NIR
Zp62oC7pGQ5OVRdZv8OD+zOS3TA3sR47yfST8FQm26hAyMehVq6XdJCx2cM4Uixh
bgoHEAb3dWNRC0410M2yHpfK3nP4UB4/fyMuhnFAhpePGHAd/o0aD8q9I4+WCmFX
0Z8WQTt9TQGHKxeWGkmc+O+45yduiZAUZLpTK04PyCELQ+XjbzrhUR3kZPUlXpDM
sxAb6L2b7Vpvde/UpGbnItPYPYWMo4X/89Mqji3SY4QLCB3bWnxBN4/FY4kGsKOg
RTCPo49QqYZ8pa9NUeL9nIrigYmjWf398JCCmkOp4yUn4wD1lOiIjfEGNo9d/5qQ
iFngOG0eF79LQMvglhXPZoAYak8z5HN5eO3SzWGC29lITlrZ8ymU/YKGyLkkPmjX
vBSVAwvPXa1a+UBgg7OF5M7KSJTa3mxoELrPFLnpL7ER8WO2L7qqDHJVcEgIn4tz
V73vLm++gMNFa1h3gwZcOmz22an5HQM/3gLkg1BdFKC7ZHwYC/QuYU9ixTiezBfZ
joLKzZVHqs8rv3TEWVybETCh3oOLO4wHWoODHujgtvnrq852va8v9ryHgYDRXYuA
OidatZqzTWPa1rj79/5KGdMIArSisoiRSLUEwfyj/+9z5eM7VeVRPmjmhBjsMiQj
Gsg86zfOkohQ+xLmwwuXrheMDhW9uavw9yI0tyVSmN//Gz5qcEKSD8ucKx3Qbfoe
ikUr1TLjpw7woXu8NhkMZ6ddz2m3pPHV/yu2g8ZnhhFU6K5ABEwJo0OzwKz/wXVL
QFBvPBCdYu4VgydaEtNSc2RG8VjWC6VtUCpFsfQS/HR6hgCEqlr9MpuryBIT61gW
hp8EYxgBaDp1k+hZU+IrNSLdC10T5oXoKKkAb6FlABnOyS3vZ8dOgSt35k3x52lx
9erqukF7WrzITd3hPHhKzg3X0SZUTe+z9sFAOcyhbFodY5RYJkjzV2nEAmQNwUgN
yn7BWZYChTI2SbgV1kMP2si1cxkTsFMAihLJozhxjiXigA1qR62MeNqDYmjsReNq
5Hl6BbsIFiHtVZbeh+YZw6KpsdAuUhyp+Z332/68cP3NkGt/3aMHIkLlwoXcFCMp
jVk8+nNln5MIohZ8tZMTXWDhb5ZMRYNIylWw1B3pxPJ8FMs7sOAOIopMmKm5c0fE
SxhRv63qGAnki0s6TvTDdWZpJHbdIArwejaZ635DCHkYkvPuJuwyd5hiQFgPdEwB
pfZcQTbuu24MMhi9RGlIXrJnSUy+dT/Xzh9e/ivGcIOdFVCcArlPtPezHe6xcMDU
D0SpuWBFpxH0XBNL5KfiOGNb4zBqormzlPHHfhg8nQ4s9nW5gaq4Apm4o4VFkbuC
IER1nK5LtOcZqQ3E3iMzg28pKmkz9XLqW2bAgZNzIo8gFizg3mYxC37rYVNYBkeV
S4aqI1MBxUzTiM+R5dAIJhizginHW8WrexcvyrmPQdfJ3U0h2AsJIan78leTyB5/
kRJm25Mrw95nldfzl59hr8U5+UJ6Rf8WLnJQcF4eG6TBkleBoZgo2NgmXR3yGnKc
OGsAYCrttTJAnpGt7HPEtucwq2XYT0jZRF6TArNdHvjN6bzWKZmWnnWmxeJxl93A
QhEZkqTagQcKq+66vx2msyPuCHERC6CHMS6tJ3gUOKBX1beTfhBcPpCAgJeQiAQt
CnJ/pUaiYk1fcqYmIxjrWdnAY1pcfRsBInKdhjIQbBSMG3EwhkTwF72RI7GENKQE
qlnmhDZBVCVzoacxw+4tcZ58knoF6d6qbg2tSWG+RFUy5J0lAm5zeCZPnQ2jc8UD
nZfal+UESXYE96isjEwoXL+GfqQFhqgx23EArAiXHYApboSJOXRkgRrK46L281bG
oxNfC4djxYZsk9e8UTTuYNU2dvdtoXnbcD1RyD9QTKkNxwPWIXSx0Jf4+p63J8qf
NwqeoczeANR4FqzjaGunf9IzZ7euL/IM5tq+9M9SiqnFfFsRIfSaXDmDqKFkauNA
SA/MFzi/nbdTzflNqrYGaCBl5ht+mu7RsqFOuaTos5DugNW3kE1gq/msRr3IbdDb
e8+SglulIJBhhQ3nNJbq/cn7nZLI9m51wYjVVO2+595f4ydGK9xcgD+pVS/vpVkK
ppRrIL++VGXd94/d1RrkevM+/nNxcB1ivB0YJrNBLRgqde2GAS45XoOP/aBu1fv1
yczFgSIo5I3VditZ+567gZBp44/mJ9FTee5oWwrXgz69EJhZcqOZ+IbKLYp6N5y9
TbcgDDE285lqMcFVNvEQpkyEmIquUnFD344d8nJu6x9aIVdIDYbwuGMNp0xMh/+X
oeww453Aoyfnrd6+VQs9YFRIJwhGf/mJ7K8Ix+6GLAXTMtY0Zfz0OLVY2pzM8VOC
mKPpRBo0VmQVeVHw5VQqjJOzmfqbJTH3EASoOcSzUc86K6vi3dUsGAhZnNIwSZH7
IeHOP2Mt6tgneiz/U12UqJJDRTYiiamiShpDarCK8cbY7HOIChwDfsqqKJnRDtdo
jUtFRFQvDsnr9HYaEpBXmkKxeCcT3y3aztBdIGTi6BnuKVG+qfF7/f9lztSZKRkw
u8FTmd8nFdmUnqpP2hgZOYD2WMWptFFsSYefd0vVOkPEbfCX2RESAoRyunpyl3Zd
mPeP17hIjJxRFSCxpXKYgbTlBUmAkeWBlad9Bis14kWxU+gHVDBgoPB0Su3O/IjM
YLzIQnxBSRDqZANonz1+Gi32i4fl6JqLnqMdpizyziyF2e8ObkQPt+mC5a+QM0sM
wZvhbHbtenaVfFErFL/a5TdliSz6zzYExLc87jmsc4xJ7R1f0OyoyA1St28Vir7U
4AVnz1fSYhHH/EJvt4chjst4zjX4oFtxPi6+Fj1Ce9ha7fx9qXOYbam3TlvgR4Yh
Ooxv4jys9gNLyXXaRfIkLDyfJfJzrZN/H/jDv7anY32SM5e3Exfdt5K0yTIcoqLF
a1qbqkLylDpTagjttBdhKhtwaot8dPa8CBYmPe1CDjVWJ8HhUdzPc7XqfNMruCpE
01IvgLCe+aDHkk6CLjwk53JYYjeyaZAyfF+lQKvteXwLcpkrBGDp9w+8AGMN0+jb
cJ6dMDO8bjYbErk5NFeTQr9Mlv6SW0CQt1c+nVSSVcalRhLqR0TM1R9BolPAM4F+
uPxT3UvBfkqEB7H+kqmMY4cWEQzCYl3GtV2QaBTFltuvWaOjxV5sT7iAy2rWBrHx
8ifp9z+cmqEeQu9IbkLtRsAHwiZ6a8R2hZZguCfFvewyftGRhFKumAmwrF3XxI5s
Mp9gjeoOrPl8o9hev+ZX/ILO6BeK4R7U2wKwxLPdPeNPpRtFoVsLwU3cYW7DJUyE
/WpY3L8Ci0y6Fn2mmDIU3y8pH9Lu1bmnjUBeG/hRmT08vgOxgxGJgFNWUf9RgheV
2eMe08JMWiNQGdyYrEQwvoxhodDqf5yA8jaY2W9YgwGQX+4vWXHlfmerASe23JLG
qa/bkXXFzxThiFGYP0ty78LQrXOfKyX0XCCDd/FUZbzKs9R8owPdzT3TI0XVIATi
C+DxB7ymPkYHIO+mOuqvIqRMqmVrtDHjYV2rn/TbAcaZoaFfzDWKykuaMC2HPDbH
+yWd+LzMIJkERlZC6GqdxLcYgZhLqpLLirLmHhQ5lsra6ZFOqCgA8M3l7ycRyOW4
OhrAhtbBWNsx1VgL7lYEJAhS6hLtAK2JD9nspM50JSEfesLlCq6zgex6Dehyn91Z
lsO+fglDwx4J+OKPKHjqoUNBT9Hbz2wKHjZO7PkH+f9gLSnHp3lV7xYAXyKX944Y
YV/15haHwA+AWQt9B/5fLfr0QkmqW3411fzr+sbjy5kU1NK0mc2n78e7ArNZEqWs
MMfZ9BbRiZnsRn3LAaKJ4tdIvmAHorUnCm5zcPScIoZm10xdNOUgcvCR2GVz/7k3
Jgz1omZML5c8zVaZCr3alGe35FTxBzamYab3KkmRuovjD+dBm3SskG9DM3CpB8NX
OoHk9t9Bhz9Pz471fm8S+hUIVfC0ofVnLqEh863r5HTQ/xY7Qm4dx4A/V10pTXqK
K7cmxra+VhTC8tOwQQtYTyikfvqSropD0X2SC11CITUjy13OXQycvbb4h4ZBG4Ev
4C6JOPdv8uKHW9aEEepU3mFj9Zeg4O3aDeJjPTpNoHCgWtm5XgjYDsRlsIbP4eZ1
gj31K50XBAESVkWBMfdO8UR9XWOaCPjf/1dxAAqklu4hT8iir0c4fqitDY6BBI1h
aB++8h0ia8MBi3LJRkIiz/+RmkaXm580qZfe+Ei+qE6TC5Dvukl4m0XG35xAVscR
dUqpkX3Q0IfnV+6fQfdmTJeTP1fnseXc/Y5Layahv7GWnbiXCj6HJXh1yOqOEpWJ
nBRvDVbEWuo6XthQ/gCtWbCAflP4ZIjGbZrSDO0BcTg2cIC7ewA74y1D5nqVnXSS
a82xMsxgHJdAYPNnrEVqrV0ClngNk2qKYDBdXT5hqDqZ1nGAltIo7J/QrLATC5ux
8Xr5ff/vDP3ESIcrtq9fgy5NMq9r1uv6SShQWg0htBwPQz9xw5XBfM2+TwCgQZMN
TT07Z1x6B5yTM3xmvbZkXV+I+h/KMJd5KgNFxQSfWmjJgW3YGOI6LB+BG9WkTLnu
KlSsHS3VsxhTvHpPBS6uDhUU/LGizbusl/1nGbmyt5FNJ+WX+Ud57DLEkpXxpdED
iPvC5gC3s2urpizcLbTwVBDnGNZj3uNjdIDiO0ndV9UppyeuQ0QKITzswvKbxThL
6ZsT2wt118NHDraZUcoAtRmiiuO85ApiEg+qJULINZdGzOGUIeKK5jhqwOKdl2Ry
2cf6l2QTmMhQbP+lOUUXGhI5MFGmgYwKgmim76CPDkTSUFcUjYA4vvD2HbLUb+wf
7oZxlHovOFwdukes6yp5jIHPOoC8WF6Kf+kZq9BD02U0iCCkeinmwvdn1XsQT3KY
QesDXO7AuWsgt+sGaBIG8qEzX6f07vM/uyNNIXm543jmPQbOExxWxbBINuTPsIbI
DADD9DBmUJGJwp3nINUmqntWJlXkyyFKZNURGpCyuJZMnsKMnpXPDBV19A+WY/w9
RpoDS/shOZkYw6QwpF5m9qA9MsQ1EtO3Dwgy2uVjAvfSTYJ7nzhfMbHymKg8Kh4d
e2veufIFpODZdNMr02RWtLpaPwP9nuw/lizXsAKFXF67Y1VyWcTwI5YLYdfuIGqw
Xs8writtPVY1PztFaq2OnBwPnJeFUxk/TTYHeyjSTSivfZsUekxMTKHmOMfk8Mbn
E+o4ual7B+rr41+4b2WG4tJJ99bk5UB1oazbeWybt4qBnxAoNNlxFaqhhLtlClre
ZalGPLsIjNXy7agTxeuZz8o6euVVbyaC2YoTddqKb2GfFhFfxVHzLc9z4eR/dY0c
Jsm1a0PnyrtP3fhVgRgrdkItpxUatv51PqpQfOafT0xdDUnJt2/QFFG4w+Qf3i8w
IutOtZspw6+Z9hnLw+L+p/eWpBIZTyqs66irkMxA47LZe3Oa5mmyMoTd/mnYIFBp
pjSzVeefxHerojxItTFKHs8ElDUFCpm19Q1Iqdvs8LdBxYRATt2jQvUA0kwjsDis
ew0ZnKpeNt1UdJIban2nlxGxaaKrh/dW9619Ub1cWQgehgJ32tcBdSrbgYfBjARj
A9BXceeWxQqqnmpG6OXTSZ4/DimZ3EIrJmwZ2T6z4v9Y69ZH7dTiORpMeYNCOBPd
MyTJ2OXSRTkUbR3v25gkLgROOVVVolTXhQ8oVfVFde8MjKglAGZTfCif5V905E41
d+YeVGyWZMrUU4xNS6zg0CgOn1lnFPJNrMotK6yaEtnF/CuyMr30B5JL+oON0XpS
afKwtjMYhKa4IMQaBI2v3NbnJuUmLfts30qUhG8dn8J3LNm5yaL9+zc5ZCtPCLHD
VBdWMVsJxKrSZ6e1qSMhLH00e2VCMRCxh/t28q8qQ/Qbi6yeUlkGCePTXk3xKREu
sGziKIp194aLVkl+Rs9pixb1cs4ti5N1L5MpjcY7e1ZCHaH1X4tqqEOrDciMKPm8
Twm3H0GoDbgF8CQatoEYDZVlWRPwYo2O2LdsRsRX8v/Boo57c9VhAiNllqyoNrCi
8tQXK6Y4DJRDRH5AkFWlYHzRbPOcoBldWBeRPeWtvIisXFYtQXxNa6EdCfu9bjho
ZpK3OxdejVstkyAII/7ZJsrU6KRGcKvz4WKjXyZcZ68glXfDV6cZMXyDqf2+Hsb1
nMKlMhrTAkD8V7K9ntDkS8M/uKy++AuQKJUPIroNu74ACIE0fZTYl85mBl1JqVFr
Km/aGkRuuXf7m5r6smP9Rn7NJnw2rcksFSSiZmiDLtci+48y9OjY8ps18d+WcrDe
cUzlpRXknhJlJE9o+aUl5ZFUPw23jYgMo9IVYFRCXLj7RJy4MXh1sATr87IrwkHK
4xUDJIchUWelvkKxluJt+jU8A2Y6iWGG6xxLjWCllyl0wEu3uKyIGEuM7dszxB/m
z/3mQBxpNhADNwP2yrqbNpas3nHbKlFL02Bh4PS2iQnfg23ygUHZWbyz1F+nvHs5
RFXqJY29zXGF6rVu6xOwLInQFxY9yft8WKaG3OYLOKyGTln04+MeDBZXvn05u9xO
EVn5GKUZp/Or2m8jLc0Pn/gWUC0lhXbZjIRKiaHUHLRAm5sqN+pitvadkOhEGxlk
UtRs3dAkagQsOtdcNV3rNqm/dA13kqEQmXkL70pfxTvzfgKQF6Ii4vFNjtAuV6ot
/1ckfBt2qMkyXdvprvZBEepxXn6oh+ae8EcQs33YCc61Y8BIShFmBom3ii5axST4
oxjVDMbOVCG0GE+T0Tzgt4lB2lRCyyGSoZD3x67pExmkL+sfYnluOGRvcYlQc1+i
z30cASq84TlKymfYQVoOsgDnYKgUU4eKV+upy1Y8R7zJ3EZ1IqfmNXIXZqQhDlWn
2B4kF+vWniks+H4rfXgXfjoSumFQndFd5Vj7folJhfyTxZfcd9ATxwe8CXHpFJ8/
OYJ96j3GKWPK6pLji7Av1uLEGMLCX3uVi9aQdfJRqLyoDMBHiuTuboG+C2ssBJOb
Diy1w1bDVovruHXMgS7jK9C+Exrqs2YZNE0g5PvAUI47zC697zjhsWTSCoIedjW6
jPVmxB/z1E+J3tbcz4kfN1jeUSd1iCabSruJAirfNI2ZbwoF9DYRbVoskMqEapwT
xJUHPufq6GAf04Yo1C07N0v7LgPj79mY0YFNPxGcGc42ySy9HPSK1McSL71fXzpO
9ftcqQ7yFJRWyxFDQiCNFsSaA/UEZSG8zNLDs2MyO8BAogNQ34lXfhyZ+Wl8gf4T
enKTqQBiy3U22GeN/ybmrkLa49JPsbN5VIPvkBJbqIobRQJsaB1ILCuoPaTfbKLg
di+rscEn0UMsGOKXGuZC9PEEN4hARYV8wfRYxlvn82h8tLu3jNXy7/k22Ba+7s0s
9B2v4gxOWhet8nFQ968zQMsNaIPiSC47Q+zyc8Pt1imqJ+7r9/AnDGpkQbKhT1ts
35SElpL1cjSEl6Dh74qieU3zhkb4HMsgOxwlwZD3ZJHwKBgET2RBbLEOa3Fdg23w
WxPJwbaGr6f9KvI8M4QZOUHN6vFh2i2cv9ol6sjdc97Exe2l+PAX8+Y9YYQJ3d8a
K2OUjMmtIGu9IATILXl6baaxDshs4go5b9ZVJ7g8ozA1noKrleMwFF6spEWEB1A7
y++stGsMPtIBVvr6KtiujQYzRc28x/q7Yr9qiE3pYObgjuStij0HD652POil6EXN
1vdF41XHLX22YZv1gmyeeZ1mV3iLl8ZywRzKoRMGz+ZZNlDL6mpCZIVBRGqkhk0g
n5xjhRMMAkv7BLRR5K0UdaWUcYjJieS7QB4rDfeU8vQKWOdFe9XsT02JPPf5kAC4
+wBmfQMUVUXeDDD0wsDVD9eLGYr9WpEm04CoUcGOWFOGU45TFYibFwGJMahZE8Yv
`protect END_PROTECTED
