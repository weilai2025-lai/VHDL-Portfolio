`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G7vVCdnieJWtQRXUVbYDFhwGsAP8t6YB6YcymLXQkqWpPFeT6CtwG8mFVqMCwHJh
LkfN0pFLOqAzuhrHEhEwjymKA/gHZ5axAi1uK/980UK5lxBatQeY+kJBriRmNsGw
Tl6m7ZJJDAeYjY8x0nj1tit6N6DdCLnm5a0P3OpIK1HEM6QqpM1YD036xbmCfHRt
VLf/nVuDR1/F0VbHqHiaQM3bFdDjXHsoMaDyDdubc7LZgukLLeZUwqQ25GWXET/r
+vG/mV7HvA0mJPIqTuktF/onQ1QpVQ4RbT1T0a8nSSUCXjkFE5m6nORMW8Wg38Zl
MQa1SsCTtwDJzjEAJgM1xRyl8CYOixGNss9r+O2ZtFgHb+nAAuINJ9u0/0fjPyCN
9KeoUyPDj7z2u3ozAob0X2N++p61Prn+JTqDmBNg0AlvpgA4unsGyly+cE9boKuJ
QaYKISWEiTFaa6azJx2o98Wd8iQ9rTxFOxfeCEQAyGYbB1Xbjo2s6D5cUK+TwBhm
iUhQOBKVg05m6JRTnc9jpdoYTrgZxGdNJod0YCqzFARi/F6SNdkIfzckttYvp52Z
jHFi0XW9jqYC0nAogTv7nPgIPda6PFR4rlDH9mlqmH0T6q0xWAsE1t5ewGzcnJE3
hzzaKWrZ39lgdFpZ2dBGOCgzn6kmTSB6Zrkt/HiNPY97tUV7pWrC9bCDrvE8j2nC
4/Sp1eEA6i5jjzj0DWPfMCzU213orNGN2qs05b3itUFj6FZh2KbAm/EfesyMHo62
gRmh1sDnsxEfsK6w919plqkBO3v12yi/CQdz+UXwzhQpxsmJ+55MwMUdZFqh/33W
aoKctau7hMy4EAEiwOktVahbjtbQ0Rl3SsqjO+0XJ7lREzJ8/XCOWzl2PdJ/zC6e
5jVdflFHmRJTjGtoGLQzyMUvLXdz5h/4D//1txHr5llKt7hMs1sIVHiS4BmRYAAn
aB7K39i+54o1GQLdZpqtOnBzyErgcYTk2y7tSYog3Hc+lWQLX0Rq3mHnO4Vlxikw
4LlEAQTTAnQfcmbiWFBBYusUoT2rfVadk9SD9MlBXOVHYucj/my/5/uoiorldrIW
nN4D+IMfUUwkYKg+mBCIMQJs6CA2RGe2CL+x67EMT1JaiC8n0/H+3WoOIsWu6R6I
sROiLlgMJ00AUIs/3Pk/YFv5WnuKV4xpQuzV6QshIXZoFxjecdqxi4pVRaA8BoSd
CzBmrsMxqPfNETmH4le88ohoD6AKvgOV9Th1IF9iYgiLZWx1NLlKh43vGvt8rj4t
71kotFUYvr1uj9VzJAPajPSzqAt1IyIuAJGKDWMjr74B6vLnnIjB6OQeySt+t8a9
G8/b318Ql5Km6BFxT7B0iufhL7cYwpXZ8g13wYRcwsJ4J5rBlWHntR/cmRQpaxbs
QV+FCSSe/pcar2bdUBYgyudJl0yV0AZUHG0N1nvJxm4loJpLOb77v/2loKq1YzHE
JcVsCVmvYyAPKJ36js+/TfhnFov5i4X25WwdFaxFZ1oSfZAClFfNv9zMC25s5ud3
7mDlT/Juu9fqzmYudaNFIQb2kKLbY2MVczDA6l6dm1V8tUL2LOACdC9666abAYPd
DQ7pw6N4QMSHLrbK0p3OmKYcHQzjxzsAj7D9k1JwknTPNDnLnt6equsep9DjzSuR
Hg64g4/0OPC7D/AR4MHWq8B8MJW6434d26AFVhvdMzMd2YQoKtv/F+JgME6e+UUJ
NXhlSCihmvMRlUdbZbpLLzI2xkD81m9r6DdgZC9wk6teeSPgffF1nbx2YyEm9NVJ
`protect END_PROTECTED
