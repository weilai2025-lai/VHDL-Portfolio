`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMS7lTr3L0fngN/gG5L6Jrjvqc15iaCqWcsXqyPaeLn4SqntiNNlZAHEgalxBpYR
/WBP1U9qaQAZcFMuP7HkG3/+v3PvCJ8PxJY0McHvDm2CwS8vz+nr7GZ88MtiBEn3
S/LtMvxfylb4VVz9ejEDdl4S+4BPcq1KMNQ8nYDazyCiXi6qixlT+xTQNyJu8Sxb
Il5DoyeN5STQmHZaZf5nA7FkH++shhq7WIVcpteO+kTPpq67O+uBV67BWLh117PN
f9sLA+KbNskZIfuO0J0S+y9ye9/2b+kKEJbOTLyTZapGLgsQdvlCBBjH924Gb2PK
2hwyBCkrWqDMA25UO7Hystczu7uEe8zD0F4vY0gEcAKianR9tjJoxttvdREioj1W
dBIqz+ppebclZRGvdxDG+yQMP/pKHtCFMiSlRWWUyIywzEicmsidEcv8swp1gHwi
25JWTtbf45SnZW7TK4v+qXwSHReosTPJOX/tSIYFQLJjSCGkVQmDsjbIRpOf/djk
69VokEFJgKz2RL3kPj5SJXF/HtukNi4oe0bO+RdLLAyoJlkpHwAOo28eGyzlA0Hg
tnon6B29ulEuaC+ZE40GKhb0IZB4vRMMJXpu9a626etfsCXnzHsTEz9PFveZJkCL
9JQKqszcfj7z6xia9Sg5fezi9xm2gzcY/tNBTo+TNiVuS/ZTdHgZNRjIA8J+UvVS
XsO39MUUHOQB+yIhLqMfurFVPB05yEUnbkTcvBeVye/ABR0AuswM6OcQSlp/wWq+
6a/MYGJeIYQkmpccaZNdKVnXLj/qA02tMiDcjPAdgdt/6Nm7i+BtTiL8ILXz3U/6
NPfJjn9kKTeOBEmKfeZrIBDmuXyXNi7Akh/pwRIUkeFzHr7YNYTSiwIZ411sh4ZB
tmNzHyPw9h/rdJRFIUaIbPT2gtfFcUfDGybUKU98GKs7TpMRb3hWLPDwvXQgSJ4f
pZRlA0TT7LUrHGVYoiOMnSBXHwTZYh/gDH5YdGtIUs9qRkH/MlOXtGOdazAFG9/x
jL3l+yxCIWbxByv1sShi1QAg7HEPVpJ1/MhXMmkYnEtVBzUqvFsBfVkY/5UaHyQw
1UP7fVLF+e8tBM/bwe0hHZO/jqiub7GSzn+zOrmhe4iv2J8yEX25lkoREwt0FrRU
5H7gd9JywyEpi1SIpyZcE0TM8ZINlopDVF9fJtfPqLEC7VAbZbh2xODMwZ5+GNqk
gEqK/YiUxo9EPZC7rWqB8lGKw1/0SXu1rg5vpSAluZy1kHUAcz201KjiRGBIwQ0C
ntq5NR+6LKDGXYMgCJ9Epe1Zt5x+Pb8aWGQO97hSaw2dlbkFMihFd6QUeZDSkJgo
Iq3hms88cZnyBLf+mCCCEcGEgOw89Sld31kUW9imYsGinpj9foN1uZ/VwNSkucVJ
sBno/BfNNf8itcIFWsGx7zy/6u3Mf+F2jkFkkTpnn0SejrR9ZQB2D9w3tIQ2nB0h
LZcw3xrdUo5r8jfyzVr5Vc6vxFcNJC5p+BOxvOlbAyAWK3hHyjyaJTbTK9KDxGb2
85Lh8mvlFJiMLje+10HMkFAKXrcFeQBdg2I6RkJTnLexsSDjuIibQRV2WiLlRjOr
/LYWV1gur08wEH9K8B6blesulIo5N/DGMijTRuKI2WeyK+jwmIT8kSH/Au0EAtOA
65+lMNNLBIZCuLAgwiN8BqQVqspk2YIhXoPs6501mDMesKvRu0ry+M/3nidvA2hO
5Kx7e3uA2H37kHN3gQqZiKGK/GdPvlrN3Gjn7OL3H9QtrIiNlqr7VmtfuyXen7IF
Bq4IzX19ELML9ug1vWcMpZATIsHMPmDojtwXOvvtPGghHnXB73YXjBUP/cn+8Ftf
UMJE7udyHbaxpfXybqBOfQDM28wG6DTuToAofK5Nb/mx0HpR2NLp8aTTQIVHaWtu
`protect END_PROTECTED
