`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YxqDuqLg1CSQRr6/wb/sI2CyEV7Rq92dR9fw1jJSOX5zVi7+ONk1UQR+yfo5RL12
lCQvM2b3h7/apvCc/fkDUfnTlNx66QUZH+h60yvKctnJzA85eGtUu0fJkyZpaDUX
CkIeVQSKxG5EUtrwNmh/feMRAf/hOGOArb2J4o9nDBY+bHUzShq+nBqmbdiBb8Kc
cpLYOmnCoF+LohOConEllhJ1Ege55FjtB/rMawnq/hxDjui4HmQ82e5XKOTROJpF
4BAjyX+RF0Sbq40qXXOTuaG3zZDXC3Ox/qUXJ4J4y5Iqs+EIb8WaDHB0+zki95tC
E5OWhTaXBMaUXWXf5wgvrZ+QKc13aKJWqX8L47xpECsGjRF4lAeXPwQhE7hwPJhN
hNOVteSbn2EFuondPCn+mg36xWnnT/Ftj6VfKsIPfPaF230+P9gpJbOmolNPckUu
f/GQBJZvq31rq8uxcQ0dg9rsTXyahCFo9VW5PyXgOGT5gV9pcTz/WL9yZMyMng3C
cjBENTkEXRMhOItXxY+d1jBlhsSIUHdgOhfqwoj1jkvBOpmGS8UDnQyXX46Ke+xQ
DEcCxRvEt/Jir+JcaV1NE1xFBpjpCKwRVTZhY+n6NE7lmXD9xj2SxHYfk9fNo+vk
4XebLj3ERe/0SZegy46/stpjRYPqJzfAEYlUyh3teJXp8YgMA+TL3nBWjAf1PPyd
fJf9sJRFAow/xyMA3XRugzf2GcP/nRdytvm0xgU9tE2dcha1M7QQM2CktaECgoA9
hb1XJEbEj8pbnZ1VuH8qS04kZYR3pHuyCw3sy4JAxowN/1gH+R6OXMPWRi2ureZb
Vn0sw3jllRHXj3JYBrNw3hfiR2faq2uCAbiQOYDMKcfvd2b61lAkPlw78iDUj1Yu
`protect END_PROTECTED
