`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7lJiLu1RnxqxsstC/uZpGCfcc8IP+eo8BQeU2QKD9SQZs+IWn/l8OgKyCZEQ/4DI
yn/wKW0nPrcWnqaELX/t1o9OHYqkik8G02Y8knZ6g9z6boKOMF4RUxwJCSricC6J
tNn4Nz+trzFYTNbST54/md7wu/Uy80pnbhg8pSqUm8LEzY5Hog5UOtwOaBqHrD7b
f7H5kfWsyisaDeMZYyvGwBHnarCxUkuYdbCWPtWvIAcxpA26novz5+Ti7+zDf4wh
tluXnlPoCGaHNZM+MZMhrJuLkS/11Bfa1JanofHOexABYazA/+asfUAik4TEZEBu
PId29hbUXReJG/VyXXPlEVxM/hjPc1hCfuJfnDxhMMPRYuu1/rhWOLiP1sTkzGAP
Q+vjBaavLi5qCmHQe2ajva0GXAqqAX9JQxeca2ZUHcES9HotFkFCt853cZhuPMrO
QU/DGvP3hvpG9AU8jjRgjojj6wQXXByp+9FIy4lKZg+eaDhZhnnqknN7CO2SrL9g
r6abCtvMf5TybmBbZM1dxguD70J+thh/DWQMa2tkp63411VYALJ7Y3oq9Rq/LOJH
Gsi6RBBwucoVJehR5lDNjfEJSRorENsUcFZySiU+nGuieFDibAIrvVLEr2ZG7XrY
AuEpIwB/bleRl3oOc3JWpM4+ck6Upn6/gYg3h84iMUiLiGZ03OV7T7aBihxnnYK4
gEgCRherDR48w2bqw5zeT9FEw7wPq3NP5TKo4Kvtr1fAB9yhXEfHc4epIObDKXUc
QjDh1ukjD1Cy3zY/KfLoLjT5F1JtoBdV/gkA8bf3lHBDc+9BCm8cl0tuh7iQofLX
pqJ0EZPMU/+ejunYammS6pXL3Gr4HWA22tCjBhMiu5ePMm7V/pWZdTmG22vIP83l
hFpYM+0MmK9nBWjmVk+92IPo8FeaBxn8pwoRUKdX8NaxC7G/mUiGhmfZGfTD32lo
DNUkHwjnsLFSDCAWTqdePFSbxig6cz3cLtSiRHTpwQi1FkPpWoj3Q1PM2hPXY+tR
XTghcQ90+dNS25Qm6fKylOhLtXpOoJBvPfu5nnOCQv7xCxGGmJ5m3rV8W2C7K150
58ntc/SI/xiQYj79vl5OS6E3+RbQi34sALFNCbGFjQv1GThx0AV2XtY/Ev5ElrUK
rMn+ZDBseFIaN6G3Ys7I2mgvb4Dqg2BmFLxDQ1b4ff8nyforezgknwn61kdV9jJJ
ceKj2gKwExMe3KsirZWZeHl9+HG6RREbKhsvO30p1fyjoOZLnUmmgubWu+n+w/xN
x1eYIW0n3MKB4XrtCFk877RsNkiWwdVunx6BLPWZC+Z3bvcRYf23g2kLvMogKfPU
IemPzTBD3ndq3u5Fc/xjGKoBdyYoiovJmVdXH454k5u2dLBo92pkNpyb86fnTdO7
QqehFDGyZlh2JXud4nJ0fMoU6Q+6XSsk2FyPAaUg3zhhfpfEsXdyVWxXip2uAnjn
lWsOkT5eV+K94WXjWhGm3wSlP3ZlMBnKOnsEgv7eqLRotE2ypUA4gJdXu6b84/FA
8HveolE5/l20bE5Td56QfOAUGcNdo6b8MSn8uA4eL7F+cBPKzjEfK4xW75nDvKGw
5NEMWTHTiEFg6NxArsdl9xaNtr0Iyd2pyvNq1326bl8lFiLIC0Or+Xxix6UuUq2R
DSChj0ivj25ctaOE0unGzhzK4xfBe1lI+1lewj2Qk90tVweRj4n+hUVRv/HjTZvl
7WD+HGS7yPYQHf3ZqRQx182cbVpNHHg/AXeLESRAUOPtL+0rwj+/Uf3cIObCMO08
nqcPWFqSoh6dQYFpPHIuyM39rvmcOBqxxsRbIiLrW81JEC4oaMcSTSo5H55AeGtF
HwUHj2vUfktgi2dfWJoP3XNnta4swglyPf2XpfOHfQvj1+Xhzn+mvp7DRZ6Brrox
lcZmmK2aEivOK/nNCjTMuXUsBFHKoxcrqbhVX11kv3VnMbO/bUfpwxOuO60XNu0P
4AV1H3t3QFe6KUmrpi1Q7PeD1N/a2Z3fWFQs+z/c10XqmejOliW3Ef+gGPE3XUm2
2TRy57pe19XmxbMFlJdf5IT7v8M6VDzfjfolFYwzXLCyUxdz3xcWU1SBDdp/aQKz
Ild7zHtZ1LbJbU23dKcbKPKyqtcfZtU7pCNhSQ1o7wWNkJ0NBYYut6WavGfRmSJe
5/S3f6teBvqaFKdHXvviO1GCaScPm+PKRDuke36QwkCTRigeRnpA6xmLGA5ogmVr
1o7Evt6QlwHyMYc9XBJA7rybfBztla2Xf0pVxhaBbBezRxD2P818jFA2WSjuE9rN
qox8AF73ZStMz+mV3u2z9JDV1RoN4UBFnDuyWsZb7YqxQh5FmKxnMeZbFWKErHu/
xF286VIbxY4qDBUwV3Hag1cDJH24+IBvO5BcAd9WPP715kZrngB8ORcfq2BPO3a/
i/e45BR2KNDQulgsnE3o0G2LfmKtHcEkrdu1Yqph6bWi+gb+tvGBE+wn1olI3fzP
FR/RNLh9Ftz1nUG2tmOqSAI0wLKgBq+ft1ZRZYSSotnM6wpXWs24WaEl+IRagYpi
8+FIlxe8r2hCvObNMP519QSC/6s8ldMBLziXGHM/rS1dJhiA6XKHtqHbUourZPQH
NwQh4ctY+0NoaBaK5BnAPPggYqvE2CdAH4WIO3C1LrQMTGTHeURaoHNDFW4dPk3h
87CVVCkT9G0BTG/wtViekzWKVgT/aYJbiBKy1u6upD4Wvm7VRUxXLoqXv+4Whruy
fPCX4p+yjCsd8xPI5RVMbc2oDtp8nID+0poytdJnaLy3GGoIzD1CQqBvUsKsk0m4
LlpG0e9EiH45BSjoFtr2rvb/KaK70wU9sCZQrtu/yR3vcAgaTlwnff1iNLzGsasI
6RSnguEjkuhqerPdNNO02AmEfZqMkBXdJQLOKhz/DAW7QcjzwIjdPMXX8jdALEal
39FMxtg7UiHyorSAUxWzKI9e8j17mv9mO7/hElWU33C5Q+hhMRBM1GHZPf7+n9lt
SeQrXC6ZuRt79SU4uLZiVsC2dsnzMSmYT7Hb+XNO2wWcFtA6VeB+u8+/8qmEx7Ah
Iy7SygNSdExMPjcBFqK3qlenZWbHNB7y4kvfVxBWOTv0uHXNm508w/Iq6RAA2dQX
BLYhzJTkr+d2oRH7E5gLCAs5pCGtuJHAMbHU0Pq4KgTOFYfd2VOZ+BxhIPGRmIqB
S//ZdKnKOMO0s8G1HIZAeQX5SVHaWXP0i+AYeb29Tx6JvCyQCFms+c/tvkycEwqz
750m29sB+ndQ8Of4dU9S+K50O8IdvUChPecbDzOzA/y3yO/gsob+SZRz8qu1tIOP
/JVmuKOTz7SjN0hYhRFxUMLLsSRi52br4w9MoD6TionYedYpAMzGCy97pW/LS6xt
TYd72BSAjUWyumAljtyTCFNPJtF8u71OgF7Gv1v7O3ZCl92hiig/kXJr6Ts2eJqO
u+/pn9tsqJ7Iyj+hAooJ1yf48S+3gUE73QYzwgb+xynMS5OukSJ7CwN/E70D5aZV
IJMhD1uRB4s0JO/ClfvVMiTxaTUo7S+hzTbtYVvomVbNGuXNvnh6eNWNRFRW62Oy
48qoLdKYAPJJ9DLCoHV4QlZD1sxApJn5ju6yCNxUJ0Mp9t4nvFVm5iMEf4W7pxCf
+sSfMyelAjC3jKDJ8rjXKayhRisPhJfRK/QTcRA8Pxwelyce0OLtwq98o/NPIM3U
ifxAdejqYugmMX4ca8Y/KXV6q27L7bSPcQdUvrbUfFkuYFWdIy0WLicz/NNpOtFD
w5ZqU5d0eHmT3cKylB3Ql5/EdzcJDd4jrKAiGk+3P1SlbhxWVop4zHQhOiE3/XeV
3XRPGaBFyYpLHXLiw5egEAclevmJZp6GOcZ9ckeaIyEE3mVQ0cAip9D79mFvqnBT
jkqy2BlWLLDj2dOQP3+dgbbF9cvrocesGOHHmupThyLrqXnpU3WHJ5VGKzBtmUex
AA2PjTbW9IvrltC4rYmf9R7/r5pNoXCrKCH/FHkICTNqrUZxBrzKOgOVuEnfLmq5
vtumY2kgpdT20euBTBN8hIUJXdtgqxYT/F/ABwUkbCJs3jJ00IqcikL90MiVVhiB
HcGYUEqeX4n9ELcGzwOWqBBGJOqVrBdy+2CEsvaeDPH3ENdNip+9shsWFooeZ2rL
41gXTwRtvqI8g/VfOFXumNGIk+vdxiatq4LlefgCFM3fY8ShXY62irwUXNxwA8yg
y42bX4bkKGzhTXWdhrIhejAggUDdPINDJ8bK3MWl+Vh6zFTaSiQ5doqPiBsOgXdb
8su+CK2NwIlxhBDovfL6VYKBH1bt0VtCkJM3mO6lAZgrTfaF+q+Jhyi6EJJQftPD
0q8m82eUgx29mQTlGqWQeFXRgAAhYXN2Vklyt/pVqYqmiP3qQTMewmwy9395mjpu
JsiUp5Sr1LXuhiL0yQ9jJxi+FrTGk2HRGzip2cxCYy69H7v9x+1j2XfXEmyuWQDt
AZmSm4gFdnJvZsbGMZYO6lD0DvkgKwpeCrTceXVvFkH5byWoUrd9AWp2uJ2V2Uii
XkmDCFPmXMuT+rb02hVUFkLvVyxI/IYkqZd+a4BNxEU5Mv3MHRiOkiZuKhYBcVKs
S6xpHN0WeGfsepuWtH5xeGYkIRuyiz9SPGDlgIg3cyAdGy2cKa5kKl4IV5xbBwk+
qPeB+buh+wCrQbwFmMy2sHIr8mmDSUL8piM1gQJGnV0a7uuZPL4EVIsq3OKCeJ6a
P/JRW3I4388TLEofcp84d+WUUvEm6nUwkPpbXHfZmGXVAuTX38YLR5VKpBALG0tP
nLkjmRAEmZtC4rtFhVU/tEREGJhTyARKddGgxDCXYS1Nl3FUneqvZwuPckX01D1p
L5ZKpuhoG+wJRjjb7fk30waMnIS+KsaUjxV/x94Hovx3+/ooI0cgyy4kvElpc6lE
W0LJk1JtiLOMmd+R5grtBu3UzTQjS3WfJf9jZeBtqtfTWsw45jLbKaxyj8myIyoW
wRm8wb4mU3aYZflHiZXtd8WRrMXItv4GpZKgKLmrsHCU3JbOcDN3fmpU1RswHwIt
ZqStB2bHSzh8VhuDHojEQTQpJTCEt7onMNrdGfMxmdO2WMAwNkMekkPmNYfjxqN7
0uOodzPbefNMJMsdz4c5Ubcig9vyX3VXsVCpdrHJG0Re8MGSxwcZkHoPDVm3mp4G
Ka0nTC+/XLnHFw8ZSXc8SqC6wRFUNhXcpJVJqdQv2YlXNaH2LCzMnS6oJMVAOR5G
e702mexXVRs3tnBbp65vnQioYJADKyL+hA8RSoegoFRchd5Yh4p9pQt6N1fsgZNj
d3pgdE0wX8SwfuPgqak4xfA5WZj6L/lIQNmy2t4LhhB0dwbtF9+vXnbCokH+msIx
X9avwcmfnKHeaMPgsuV9dEfWbuWNR9mugTSFYz121mNIH/z4iyDhkCf2NsLQVjGm
7tI2IcI7AYNyo6VQDn8BcSMlT7uYiBTa7GHL38yQQPU2U/2A+25Q1Ud1VC5rKSQ9
+TbFDxb3jIj5aUgOGB4unhLLavxzBsq40ejVh2LxgE1/Yt49RfMwFzWq+v0OPiTO
LzqtalhTHG3rruA2CpeEpO+k3vIwFJylCMb6opfcSNZwSDonYsiO7/ADgjJm58uw
rdFc3CsEvZTLf+Olzxrq9FPJCajGWpwPuCreFsdjt2Azwee39eYdp39ng3od8yst
CEv67oS3Owy0Kyjc4nuytqTPP7KeUVX3ZpPrnRb/VxoSG8sPCENBiOyfCaiUNNQ2
FAoavJFUC5GuVdsnV5p+gCHdOUWKEftkuAWqQJ/cQx3Zk17NFvsAfJYQLA0V5wCt
PCRJXkyIIbPjR/MShriLGsbjBxUhSsVSuF3fm0Pz/nsbu4J6Z2Xhe72MKbp4vV0Y
h0bm15ZGDIqa0joTuxTokqRTfA/JAsL2YxmZHC3SID5D03btrOmDNADMkPwVya0T
j37HL4zMwKIzjrmJEi/EZKMKA5zQJM41WrbbE1gZz/7CF6mAIstvEe2p+NUiJL81
GOJlsx8aQ1GDL0Dd6LsXWx/7CxwELrXIb0nuYVQ7LVzDELp3Tmiy1ntFykzSCudb
aAv65p/C5Xb6UjOQtjVeD7JBN+n06ooZfWPrRI5PYNf+5Kwir6Z85jM3NRhXrqiQ
i6nqGjgI0rqpeUrxGFZhwd7rqr+9Kf1QspOMIDAdhe6sr3+dehTntQFVANOxG0xO
U8+943yeuycevKKGgHxJvs9RWR0tr9Kn1e33bTaTE1ZwDWT+34BWEFNNwdGL1YG6
Fouq/acs8pM+XEer+24mmLtDCTJjt8wtTCOT3mDcDay0fAeVZu5tXpS+DPgjyk3n
CzANV4YyVc2SLCEvyZT5ynhwQroWceFqm6wKEdBETPbjgXYXjeMSKksymW7W7p2e
rXunXBSScKTWB+MKaYSzUHf1YY96khpsny/V1qOCTKu836Zf0YP0FQZXc5LJ3YSx
mxMj9aMPPMfDiReJ+LTx95cEYRpHpKHUGrW+a6y566BmFXuZLlEwDYbLDstsCeVW
X8loLyJfbhHLz2W0wFdS8TGGqDnBkZKzr30N2GlROmVMAPj8DPeWPgUDBxZBjIqm
u/4L+XXeRuDLBNG/0p3TppwvaJAiMibMm+6aZiL4in+UkLQeEaDSodhk+CkIVdWc
wpOtj41reRf1HMsLXIp9Sc6pyY6NnDyCYHaLCDkcWFMDWB+eSaH5AmP/QV6DMuZa
f/eE/JJP9NiBGz/i7RbNBKi2kfQ1glhDxE8mO0iDMI4Z++8p2Esr2Q6cYWA+cSeT
kR0dOlRVps3QmUprggTNC0jSWAViBtZD0BmOqkqzRME2ChS56CLARbG/aWV7GzCa
IrrdAWwJS8P7Rd3jSNvnobzVDiUvTTBnVoFVgrR3zWtx21r0sWgz2el3OKJcCjCj
7R5nuswrZMFbasI01Ng+SiwV4QIAMcExLov+TjCDXrJDgQ/wjUC6/pDQav7Y0wdS
BODAheIGZagkemGUb8nU4+GwzHeZdCdgLeR4FPa5R5JEWknMzC2IdCewro4o2y2k
LyzSHxY9QJQoN8uaBTR3sbDFgPQyT/Kt2UEkd6pYu+0XbdgCoTdNyUpWAkLnU85c
2dKvc3T0P4mr1kE0WH/+Jab+g8sXsy2AURTkh0AA0piCfj237ltqVx1GqEv8hYLL
B2R1A7Ei9vpHHfqMqbcFTQqc4hCxQvWJ4ZagPN3bz49e7CHu5/OOJdN5pMDBqIDj
IJimuXXOpab7deIFxsb9ypzDs1XeBMBZGE9MCB9RzYTaWGtN/NbP07YEGczmZgnI
QJJhTTbvCQheuPhpy8xh5VfOf48RvMzGTXq4NBQcCOJY2YeaImZ6kHeWwT9JDN85
N3i2mJFDdQc7BdV77kzWYB2pM8DusQoA341zvmUSpZsDWge4P4aJWdZUqftDmzLX
lxE00kV8PwrxQojAkJcwrEH/mJrHLKhuxbuE67Le8xPsRY+KySxjthdje/JDFAqX
H0hz5MEH2x0pYgM+Q/UjX5ELW2fFCU4aFBrxv+d+9Wtlp9vhaqTqBaO+uosogtRR
Wu0EnDfrSnoOqhZI+zoIFPnuqQdFWN2K16/CYJ82JICNsx1Bq9cZwsV2wuE4If2j
fZAUdmxE7khTh8TKbVMiHNexn6D20DKc+qGnF0d+pMwHadu37bzVkYEKxi1ENyJO
y2XbodGdJtD0TfoDxnh0wPqEMK9QgMw2YFPver+nHifF7BAGScqzjaK3ZWmH0Tlc
S2zejhWPRJsolKZNTxuZ5X3cg7jCXF4wJwZOS95Iaqae8QqsrlLNIdkcXyZ79Cjo
mgmdVknZXfcd82zruwzKp1B2/qc1iSaxFP3WPeGJj6EBLj2zFTOejNaub9vc6VcL
R1ys3pmyD1HqxQBph5phGpxMNFVt/hXmi8N5GX1O2dO+kDzJ5pbf11QQFKTHbLyF
L/i0/mW7OqWvDoGcOzZLCbgRay7y0vQmfU83CzVbj929fHhCIqEImW61B1RuFORn
1OoOxBiBEt85IgzT1Q6POM3zhIKcg8W18Qpn4etr6LYH50OpsjUhW+1sVB76DilA
H/bQHSdf5Kd/E2kKBU+gBq65FGyTJ/kaO68Bi9MMtwyxvb+s+Xb2Gyrnw508QkJT
TGQUCpZYzcJoPh4glDFPEgJd6Mi1DSESNPuWMhHAkiqA+9/S8vq27FVLxxjRa2XP
PmFJ30mNRvm5iCjab7c/PX97yyk8bhhvtAgbg1N2xiMjVI3KRaTx/lacajT9/uW2
aGhPkAXfDFYg85sLYsFR6gH0LJBmXYT3McQpt8L0358fddDk7Ac7KDpClSMOpGlL
ckDfvQThtJJdui0LDamsNJJphs5OkZp+I5AvHr9UzE4lHczDBSPy++Bt7raPEK+7
FW9aLW/RFjkBjQwcqOCLFxEEgcSjQ8d4QfUPZH0PG0h2DQaGbdLsmFLd7VCwlQr1
eQUHsRNGGQtxLvnA6+7RBezVFyRfLBKe+3JqeCuCB1hIz1sj8dYuOMTxR3Fld8WU
rL7dailNS+v7SDFSBkz0CvqiuYA+LD3uWZ68hUB6PGsBXtmMpUZaCt+nxT6lhfSG
/4rB1A5yrVlHHVGoM5yO53bSaFYzJc136MO0Jv/O2b3Up/p1xsFgybwlYOVhNebT
wQwMb1jpbMgLElVYetMHC6wYjN6uQj3mZ3l+WvPNI+7sLLMsYXMnlkAJPmJ4KVRJ
xiGTaRhz58vZ4CzdiCjmTWnrMH6AcdPhDOit9hJy1160Cz8frL5PyODTaPHZ6Xi2
e88iFJp3grFT5e4Lyf3RX9psxWB5y/ARcWFDhB00n0mI7YqMRSjJZ0aApbqpYALg
wIQnhsnrUbwTOSOXcCDCzkRpqruyHw3G/dY1Q+GEjTAUnUxbDPomGpLNQ6894VI0
ch74LdRU/oW4eBr+G2LPAdivVt+QA9OZ/TvEnWoF/MHlRHSZDCIEthfcucbF5Vex
Hp4k/4foai3QURwyD8NU8cBgDaHDVVXq/liB9oU63jPib2cEqggRh4PzNnVOCBqz
SPgT26peHd//dMTkAyj9rrqX8wRAq4+jTOPkFsA6DYDuiR365t5yQ8e+5h2/jnnt
ij1MAbVlzyK+yptkSX05XdZhPdqlXEf3Ct/u6RFZ60Cx5NCsKIMpLKg/9yLaZhtu
DJLXUcNTYK1sqzeghttr6UyTilVNhe009adUv4Fks2irDMRTnGKgS65CbQtOM04f
Bmzbcw4HIgWkQufO1ZX1GhJ16QUA+yWSSpbh/4psfFlQuvURXpXy5InC65xd8vxt
P+w5D9Bi/Hty+3cmCGNNEB0RxpPGgbOAXAzoPjpzkHkhL+lfhBS0ORU2uhzgXrmg
heyZBGKThuHc4C9ay9t6Qh9ztR4Gp679gUOjToBBnmTOCn6xUFnnOUs7Fn+0fa3M
HlRMlZnKmQqyYUce8a2GGmzrKNkzTXsUDHbyQbb/NYxnpLt1pj5OVY+8JpGH+Pdb
+KQq5HALExPUIhaonaCNQKpE1I7Yx3GyYSlVobc3ElbMTz2JDGiD2xTXsdyr5++r
yrVwuakaL1gcvIQuHR9PcuE95yFxt5+VLFxjZG8Qo/lVy3KLkScC1MmqiTYeoDVx
0MolgdXxaugpVVY7iZhIckQuVnbCmLIFVMd2raoQW4L4Z6VJceNklfT0VtiJWekK
rDTqGZ65fyMdY/WA5Cw44k/wSK6WwyWzc7odLoc8mEW63y6c+5udSXFrBM3o9yu7
a6NoAPsyy1KubKoXYf2jBlaos4vxNzapj5KSYNgiTrWykdIBYU+UqEoyTJ5YT7rC
7bhvZweV4s2Dq+PKN1Pr41/oB0kINi1cW83O6fu8dr3XfYAwYq7q4/+HHNWEWVAl
a51pdzfLAYsZTuGTf0xKaMAEKplU/KKw5gNDWcwWhiHtAW0i43Zv7fg4xNpt/Mp9
jdEk1GGL4OlPu2O/7A0OOU66ey8br6NVx+4e5E2GyNPD0nNE2Gbk/DlsJDNM/XC7
N7hYLdkbceIWWkGGV0Vx337EddMdx2mFyqYRHNMqzGaT0P82FWl5Zfy3WlLfz2Fi
NQChSHMWDZk8EpdSnbw7vD4ee9CFV9YWcnNLGpgCtfSzlr4CdA9vRR7m00XGF1lK
h+TBWJdYBrVJGrH9Y8TTs4f/Y612IbAhQWUOMs0uRLybCQhjDEFA7vXqKZ91K0MU
6CamN+Ec2i1eS3TxtjhbW3hy6TpIOfDDNZb1oVRbRtwFia62VtM/yfvu3nVa2eCX
RVKjMOAWx5tHYzQhF6qinpRP4gQ/g/ekXB/nV6augltPESv0afCOwhz49zf3Mq9I
HxQ1vsdbtx+ta7Mc3Z3DyZQ9+eorvzh2bN4qG78b8w/iJP4/4uadcyAS/CEWhRGf
CRn2u0rm0LZFlN+tZ7KotY00EFDN5rV37xXZRfLR2JLc1cgKmRHqGzaosfr2Zzye
u3f8lPC88OxnIe0GJdrd5NmZkPa6JUQD9hFm4S4gdUan3bvo3EY6TMJ0VJ8Dq0gA
kL0A1Gv5v34I7J+B7eYSU0eaxJRjw2ZDFDo4umMrubL2n7BebvNpR4e/8rJ5XtlV
AxxvF+en1ZqPTZUeTJY5/wyJWSop99BO2kSG+4dnO5APoV431ehe3AgjoAXKXNUk
hoPAGAasfnb+DgjGYxsKE8mbvxriHGMLPMobwvtL7+drTmy0eOLaEoHbNbVvRss3
Ysy+gzzatp78S99l4gYYRA==
`protect END_PROTECTED
