`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7Jz4WFEEGlCJOWCCwQygLR9qX2oQ96Ykp1WJTI8n+s9BSNL1Sm/lRl5k1T806hf
PoJFQkl31/h9+AY2xrq9+8v+/Mg8t+bZMTeCVFbq+5JWXEpZGgZckoNEdUtJ9tlB
L2OSCvU8Ordpy47pGflTd4Ytya0L6/nkHOx2kG7ozAYAkPtYBdky9jWrchsexz5U
bl25mlRIh3wlVwWQUOL1N3fEuiULGKte8bD7uVt+qvygUsZdhNotFl6LcTScTbbn
tCjou/TSJamhnPedQYH5S6wi5heujm8CPdL9JngFF8PxB+FSD17jIrY/m4/DI1k+
dnzfPKrYn9fPgxtPZZeBwQWyNHSfupuGjR+s8tkDlZ3OEYn6IZF41uet9pVEIwPi
8vsL8UZQ2MiYc0gbWWfXr5bQLsloHSaQztAiH1wfPWko/usJRTCGWNltTKKOqSAD
eX490a1UrwBy7yjpA1JtK/EWcc/ErXo5fXP45+Hc4gRWKomAXDVDqpLQ9bhrbLAK
QP4zLSK1lYDvL7rUj/CGw0p6GQztwqe636ZXvrLR3AkytyRvd7g8LYyQPGRNiK5d
J7/LIJreTB4RnUHnojJvCEw6eBocAXXc8231rH0QrMyhAzHaT1hhBZh1sJeF9YZB
TFcaD9L8NL5USiL0uONZSE30tPL8s3SCcRoy3cQJAvMwS622tL2IVG+6ZJvWjyAC
USqkQnZ8kzcHUptY/WWqGwIj7DcqI9NnAWjWofLvNrzEfirC+eB7Fdw5eqBU23eA
9nbpF/eMoirK+CUr0DB7tmUxxCCRH24GiJK5gAqOP6HGQhgkoyDDPuAIlzWosrWt
483FEokt3+3aBnMT/33fctwKmEyyBdjjgcAjq9kfIhS+jjeQtw1BYFmfV7BVqpa5
tGxa434lerAqZ9E5KHzSeke/VHwOlKh+jLu0w15+75p/mynL+o+owD9kTX/Er50k
Uv8VPBixQlNQmwuoWDWGbJnqyMJGH49U95knLAJIis8Y1zF12SG+jUF2WoXNTo7f
kdXFvm1D+RkjgZFE3ju0glZY2SiD/dy513318maQZXuEtppzMe5p9RguBBQp/GBY
ZvnV/0JTfbXNk+uXKGDyEKHgm2EL5sYREYqgjvyCPs+kJWN4Ubby20Pu/aSJqbCV
pMtv302/cUh0hnJ/KjaGmis1FVMNUfecUpTn469N3QTgzEfhEaufDieNApXreKdq
M6z7IWsiPbn9bWsxm/3fYBm+ckrXxt0rql+gvmAGmL7/ajTcrSS7z1IJQammVqTz
ssd0H3vNuB6WDNt9CkZfq7Qy8Fb8e+yE/0NitCsAE7aYYbxMziiH3pLDWVQ3f3Oi
kMXuNbl+EIehQGteboL0jit5NcVCS6xjgNvT7oZyQIMFlajk2v+vPniVZs04NM9x
GGE+yuq4kZWcCFXlmoN8NypubQrvfD6nxVMsp3kzbUcf7uiJJGvfz0g0baPqyJxL
xet4lnFsUNJrOOkiNJhx7BsDt5ZG3kM/SruFMusOcnYNMWziHK0NDjRM70H8Mvcs
k9rlEXkY6Upb3XprR3wYKNCWs0SWjO1rkg4UKhTJ4sW5gYE/72qks8FOXPuMh8uZ
HywEeTnUWi9quuvBAX+hw6enRFhlFKTzMKigh7Zfih2mceOjZwLyH2arOCBq9sjb
OvRMy3Yy97XSFabAdrDzIq7g9lNLnDbtCMU0r2dujtjm7Bo/u5Z0m3LhcEwk7AQ9
hultcolFr09oyNmlrpkJ8dbNU8SrQgHFZ9QizIOLghQ40RHCEoKEuFFeyyxfvefJ
b325qUDFioXeS2aGVaQ5OV8Xp6yyIalpovRrXSisBSi4uLgrg2OJPU9EMF0sSq5N
nr1SomRaxetEfqvoUqyxHkoEY6iHdNPnokmXBDiIYM+/ddcbx0+Nq+JiOpIrGr3D
x4zC1d3fnKr7wpceASuXwLbNdiS//yddFlkTw4bPHQJN+aulYWDosNjloZnN4Z34
jRQh+JB5LGBYLv1FLLCvqPVgjAPAjsxufFpz4JpPbE0PkG2vDkv0Qp48xjGbaFcT
Rt3PMTMQ9iVS76m7LFfVkVcRMOt9EG086GYgxp0imbmcdeRHfegNsUMYtTeKcoVB
rNkDhaeUeonCAZfrVjC0Qh18LWYj8GwXc0UfHeOEM/o=
`protect END_PROTECTED
