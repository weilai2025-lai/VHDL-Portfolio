`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OiyruDyFOi6eVz8APXoG+YlfXPv9ovdMQmuy/b2k83xXfMmFZShGWqoEMqyL0+Rv
Y1Q4RjKQZXIBCPYLnNjPLZCXBSF6y+qB+nXBYad9sc+tcPQUU9WFWljkoRmHWeHS
PGgXs6vlbMvJ0mt7ZuVp+SfTSBrBJUEb1v3u6vxZyPYHpDG/kdDcBrA+z8KjFl+L
NhesyLtVej4AaLWVJppwtRAdPiMK/gKkTA4bwclntNbu8CSfWQkjPnm2brcS5kJ2
mW9Cqcr9IDxYWwxNWF9mf6jko53ZXnY85tc7biT4EOv5UT6diioG7PLfdeUy5Hfa
7vdrD0eYfJYRUiwBkqz8qAg/PY+us8OWbM3E7n9W1GoB0MQUIDEWQ1QqBKr+JMdr
WieBvEVPsUaBkmKDq2TVvd6AcvQTioXFS5sNR1GoPo4s+G3RD4HNYGE3CJz5LV18
1+WIe+BFytmkpaJI3QfLiwkEpKFpgpo9p/fEuzNnbJpk3hqE/3jk3MeB+EK4qgSJ
2m091CcKcmplo1LWBeqmN8hR5R5+ah8HYzUQSMIh/PYYUfkVVw61kqzl9jTTyNM1
eBREAbqdqnqMfNUs5DGrK+W/LFnpabOVAM9UrdDw0+b9bdr+8WP9Y9n8VWysiLD3
s7+w8DOtHKd3Qr9VzNj6oqbMUIlJwgvsev3FOlACZ4ng3zlhJTFj8vIkOrtCliRp
2USkL6BR3adFby0du2zjl3iGXK/PmsGlCtaJbIHsNrH0vdgKvQFailu+V9gsQOyE
C/LuWrAPDuXvc107B0foC2zbtP/ltCBEV77TFL0lrlCoYOdhX+4hlDYLhFe4rP8Z
MiyC0mTPZ0nkod/FRAOJfsOICl8mbDa0j/pCyCAbStCZzn85wKr9e7sUAqoSY0Jc
REWjNzHPCn4VQpqjcAMYqQjxvdKeTOmQeI0gYWOZ5hsvyIfwfSBgo26J5xw6p2Vo
hg4scAeGIHS8fSRAdZ4V3Khgz+6uLPj5WlK1N/YQ5OY1lfdYRXmdJzi0MkTorchK
RTkqIyn4byP1Y7P/Kvf5uWxW3xngyHai680zbF4+bkZp4PnI5oYYEmTtQjUFcA+Z
g/p2qSWdS4heWGsJ05IewKXBMs2F8ZH961M1051AjG0KNwsLF/Sw03U7rE0Fn/8d
FNnPF/3UxxrVpwS6Y9VB5pev85+LTNheRl0GXOstJDdMY+0s9LiY+ZFhWhmXvafy
HBbxoAvRoCLwnuLzdG1rXHrWgRdctizR4vkl7hR1fit+p1XS4iAeCHZ05Gbru0Pz
tr/QMp/l12bJG5oY9cUZYOBMbQ4PvLj1fTnM6X2komfB/SSLp2rlbzZhwFSYTwGR
LIc3X/BY0lQrWcrThWykvoskIPh7LjRpIf6cYY1AMgyMaQRHns8TBs2jAfzgtgbJ
SLbOjgfOQOOWJgAv5G2ttKF8PO9oAJS7aXBW48C9hF8at3dVYbrClVtowMfUzcN7
QT0rP9vgFqh9pcBUni4XvwdhsT3ESgaklt3/eQgw/tvrF3REw8cF1O76rhrWMnjI
8DztZyx1RCd8DMHw3bRTBqE07z4K/RqTo+EQ/y7KRGDq/YfFO5KZijv/n7StD5IN
tUNGVwM/a/VzJxe2YD6rOgCKJQKDdgY9G9CXyUQdF1Xh7y1WFOK6TMQvCpTSPmk+
H42JXOvEcML68tn9ARZtCjFn0MXXeej8QyWWPg4vNag+Q/vRTsK+fq2tzDKgnewH
JLwuDfRNkontoa1ePQ5riTgQFhW6IMcfyX0v+sFBrf7uq2gXNwN4gDSNmi1JOyhn
`protect END_PROTECTED
