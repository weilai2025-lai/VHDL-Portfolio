`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61j2R4/iS3InfCe4FM/IvHdaxwLr3Hpr56ADMP3d4QOYdRGlofxe4GYhVSxAJNsf
Nn5zIC0axOcMRjCyqIMQIbyB8avAqAKNSucA1+jJ3bk7b3snaHQOYVRCZ4hJMTrf
jOtOSqnQ9/O3YLFJynRe9dxrOud5/k/ZxTdTkI80PzEwvOqbT9AWPzbCxP0axMOU
kKCTaYNNSNNh8qDctxqT+pnNNw6q5LBL68aegzGq2TTKVICnoQFMgwutdENzlXM6
T6a+1M+VyMtI+RW5IpaaTlB9mnHZgjMjygY5KrOHStx/gnslGUtetHseYPA+Ho82
gULgnBfmQ+YjrKPLI7i7iNGK19xtgZAJuhm93A6G+6B0pDUSjFgcpSXBH3X5anWY
upqNGMZHqYDs+02KILSHrKSktRmS6L2WR5xt7QjfktCv2r2uS02uompnRCXV+VLJ
Qvz0aJ/jLJUxMgIJVObazjp1FyaiJXVnqqJVNrkYLUdLe4tVFO68kGH0694XYIls
G+LkjTAHzSp32zZD5shqp0gx9HtVo5PnzW/y9OjNA2VD8SvHia1C4BWjrOLk3WXa
9a4XzRbNu2zCBLpV+DTeLgCQ3jl9vTMrV96mpjFE6FCk3LYmmSQU69P4LLNRN+bY
kxugbH9nm3v4Loz6A7Rjg4j1NOJ81pm1ioJLqySFy7n6j7qbrzJSGa/K8Gb1MegU
+UFkx7w+TrS+v5rKzErEYkwCFRVOIRkbvwdpdDMKsQkvosnkG75tZ1zUagD1+ZBU
xtyzxCutq/vu4Vk5+eRJGG1vpogqrws0WXPA3vtnyFNATTqv/C3O+mpyLehv2Y6t
b18eksyzeHc75kD5fmis5OUrF4fHHLcVF6Wkp1ZwsZfPE96QXLBg08aX6Q1wHA8c
EDOKEz3eX1Ljo0RT1mJr8gHJBhbO/rxFlF4VemkHx3/fi4KugfOFm1+yXgrdrjud
m/aYf2/yAHiYEMxWSiKf2jC+GNs2LMRLgpvllKOsrLI+nqUSZ9yDCYKA8hwUt9Db
xL5MKEDdzOwgyAwgihJRIe5eBUtO/tU+MDRdiF79YjXCbHzsZxWPp8yjMOh+4b4c
xpOoRy0xWlJJgZuBCjXTW08pU0NlSXyG3dEA3wYuCsCIrrz6aUBrWrJb5WCbYOhL
RzoRF/DjiGdtC+eW/Fcl2Eg44GpfFbcVUO0EnfSkJydNFz2UqM4ne0eyegssU/Hp
wM83DS+A1A+r2WSCZorcQ8LxGfWfwJDo9OdC5WvS2XdGv9HkQLj/xmZoQa1SjX3y
tgW7LYoSpWdXDO5ujvvB3b3pw/NAp7x96CqmuKgMykqh62NvATcJFsZE7XO4Uz2T
rUGjQWMW//dV2Wf8tPsakU0H7BG+FhJai4dxklSjttcVedYWg+8mAZMrbb16t/6g
24JsFKHm3JbE9vCo9Kg3xeUV4S2Pzu57s0BHmzDmecUftLAyT1mx6PV1LjmWjILP
Fw2EIW6GdL9d6CPJFw+a7void4HiYWb7JqOBDvFlVCUHDQ8J79yRUqSxZgepHcqW
hSZnXmy7OJwo8mo3TbeQNg+VuZodi9CIa1o/b9NorlOCg+G2mJKDg6xP8FImuQMX
oI4thKtSHUZg8/BPmmsnQS2W/XK5iD2hijoXX8Zyir5YTyJby+IvRrfD+/AF30Yb
b/NX6Yk0SgRmF2SW88Wy2azZ76umQqEk66zEwZrfJVACSBO1YQu3x+6lwrUK+vL9
4jISEJLrMQr2g758aKOfJEpAiayD2jaEVNkt7qMv6neo33pFABAVJAY7Vk901chU
jKe3c+fNgVKejN2P3izwk5W1LACYuNrJVgkCiBDodCxxC6UixnXmiYKWYeqdnurg
DtwGvDNKW0UVQJ4I9fwRRqSNbRcNk6cdeil2fVg/XfR8dgGgo8FtfTZOPsjTAXon
GOHJzbknnDWDB6mD3P2sEpwFmr00v+fvF/g2atohYHQM95tRkDC7JItnL3VzejOY
eZeDTwP4r526PdvNw4hoplF3AEqRt5S1A9ne/vuFVsG2UiklK1JDjJAiJwSjzZYp
TfdBk3BTTW3T39cjD2D7xm4SRAqfJ5fIgsMM/ZLvAy3aoeU9m8o4OOmZ8dOpLli8
V0FW6xXIvOZDwlYqdzZ+Abpy6TNnxw4QZw5B6zpoUkmpzfNmcrCoRqIHoPvBZKMa
8Ui+T+23r1//BtGwrWAHJoIsFv6Bx9lpmEfumoSE8Zm5NoCtRbfYZ9kD9Q+KJc3Q
E8xznH5eSeurTMc2zagv/+h48xwOYo8iAk71lLo1H4XbwYYluhKJFOwQsXFrpFuo
kUkD3MXBHJVt4ivYvsV1SfXyYEmi5IijYUAuIn3f7m5e1pheBloqKHefO3sTaJtx
2jVXTDhkd0EvQvLpHxV8rxzo0gxIKXC5d8Gcdyc2EgILdhU7raSX50MuM5m4CilC
Sn36O3rX6OX5DcGMa8/fx/6cVPg6X8A8IKpzBFTP1qPK7Mdsvb4/CFks8ZI3o7//
nB3Dda5CiNJfxjAoaZjaAbV1T9T4n9RQwGvLP+e4Qsc/SMpJcVhs/xMGhXTG965U
DB3U8BxV9fQJp8KGMv/NhgtrbZKmlOwPYmO7q5yi71hBUVRHBtc8hnXSDG3Wv7VK
VuUdGG9keJWthSPWtP6lNGQ6NZPCBk992mzG5C+pq0DrtknnWJ//Cw2OOCTI1yAI
`protect END_PROTECTED
