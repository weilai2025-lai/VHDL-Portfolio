`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TyrdpUIqdqjggXCVTvr3gbsRgOVcSZG4ZAE0Pp6iyomsUWhhcVwgzoKYQCsWP3ao
oZBUky2wPSxaYyR5L0HgG/IAQv0sa1BgRUu6Vi5HRDG9IFkJMmgBtXupcEnHa9On
gxlTHkrC+vzwSLTW6setl+u8GcUprFbOsjZVS2AxElqeZnZh3kvTm09Biu6a9hV9
vWhQ7lmF0ZHSIsrYc2M9MKfKhTqzQmpzh1arsBgi+NO5C9o9J4sOl/gMs84Gvjsp
m+u8gZBIy/I/1Gelsv30W6T6/Ob3eY3emXARj2PDvFeXSW9CxZojwmFKPLrkus7Y
8aBkdHOExTQTmRKfsgqmQYz8EbbAHsTIRPEmEdUk3LBW2uvOxXQVR2iY/Np34b5d
NJTU/yMx6CFh6b1mCJnKsuuWG+/h+MuovZi0vITx6FMoVyoRDhPo2mnCL+BIhxoZ
TVxg4JCqupjFwpujUGZwQPqMyj7ab7HLlof3xsTzvNgMf0Ir3zMFMTC1hgmi0TEV
keFZadEmvjCmVqlWqk3Q3A2yTF4+RDJAPV+fGJZq0YPCOo8gWMD9SvpXSOfwsCrU
4pnwzZjZWP61T4X9oYW4dYCT55CPghe39t65UXv3nSNSKiwGArjTgGGXhVHGiEca
nM3YOzzZay2vC4xrU/fII3RQLu5DKJhptMoeg7HsQFi1j3FtNniKfUcgHeWG3Z0U
qbYWaAjdbWvjkfayAh0lHcbXegF4BA5nAS5LR4PoWkc/FHQMa/2upTO+IgeSL12c
uY7gx1FxjwXBxOAg14dOHMbZm8X188EpzsIUtm8b65Q094DJvxKwgvIGv3yFivwr
aWf2qMbg6MnBLpwaePi6QxUkORMOwUvEPnXpH8KEfrC2zQ8ADM/VyZTOOTHEuhLI
CK4jqmNWHE5SG2es+qN6ZkGi6q1suJ4RGU9FK/hHGEF5Q104757aWQtFhjFq/HfF
/ojpJ//G/EVIQfsRhqCG/c6FF7NLHRYuVnSIMg+gHCz2wfdDo4WmQtHIRzMP0p9c
nC3s2Ds1mxv8foIDntQZgj2q7MpytY958w9Adcm9L57ft17sSQJOYN5D9Wn+UOWt
R5JszW5GoDgAuEZimxdkhVtRWMH2VsVoLaIIbKTdtR2Bpjlw6jtPWOcxy/vFOMg0
2Zxd5jNOol7TPNfPVXW8dsIyOk35FEs1atFH4B/GzxUg53Z74PYqxg1BbtuXH2dh
tvNrhUMFcryB1P2lSA3j1dZfBtqhJ4N9f/u9Rk/AUvX03+Yr2Bg3QNceace9Xk/M
ZdM9jKaO9SXBylDIaPHYFbGHC0Kfe87hSbYt2G8//3cu4opFiC2l6fH8v+G1brAc
Iyj/1mAqFdzPTDxPaqCwv2QX4yT0qo5wpCwmzRvMewIcz6fF+AsjJ+b2Hg7KP9rv
T2fnnwTnIGHp61ZRSFxMrFliMNLiWYL3jjmmxbWfYbQbR1NnFUt6CI2m3yGgK+HY
G5ep//ZMiKgLpP+lSkV3NGL2ebOE9YBOlpMe9hC/bTqFbR8m7y8b+eTcKMBLWbJO
s2E20Kg3CjK4cTymavZDy/8FvGYVHgjhaQM78KHXzhX515HBb/bPlv9tJ8RGZZGc
C+lzVobIGYzKzGLJ3uYLB9Bwv+olnsxHXg2vt6eWlvaqvBZqQj61UkjiBTMKeCxK
zYrVbaMUz2MDye1FutKKkfAQ+vX6d72MzkW751b6NEIBEw1byPmzD3nOHh/gY5xn
7xrzfd0lyWFR+YwIT+8fNNp5egJWA/vpxTDFRMZS1ng9seC05u3iuWaQuZFecrxU
RIy38Qcm86M+3gk5Wc4xXNaz1Ma8V0RndR53krpdNfccsuRcqqQKckzdoiOmDPz4
97qHjKsRB4SB/PilETBj+6dtVkKPBYOT3+KG94SSyuHN4D3qdTrKrc24/71cHKhe
+qJ3ROGunRTr5mOhU/xYG6146MPTKzZmoxdrvP/WSVm+pylyJiLjIAHXo7bmZbYC
T8D0UraP/TomrIpOBQUrunBOD+PPMAX2UmlQYYTdWgj3BSezQYbETliQsLK45MjO
C1g3xesWWv55piIJcEEMrM12A29z+xHb/u2omqunff0pvn7+9U6pNlTj3W5Sv0EA
E1B1qJQSI4NkFIKilZ4Bj3x3DXxKpKjPwxac2D41t1t/kRIqeD2mRx5H2dX1dbfw
/1L5bT+d8q8B1IdC+bXHwFRUTWErW5N47qLThODo+2/NFtfmpSaUkrLJ72ue47cj
lBfDN4LCQ8+tcPi2Q5w0RJAI6Q31/Gcq8W7gwk7KOYQdXqZccxGud7rbo9kM/V75
bWtFGVNn5cDMjZsPGbBtkpVBTc1RNsi2efyd64P5qFHVW422PYoyQsrAeE8Ps7pD
IV9G+o3XmGb/R6sX5THYb1lngUgKLlmj5dDkTbM2Ceylw4tgXdFy/kdjjvwfXrQZ
3NfAI/PB5SCu9NCUZ8y28LBGXcvMgoDFw+rnfyLNSN1EuAcNGrkTshiGMs18F9K7
NJMLYwHsirmjoUEA01wnNRZWL5gNdu0uE2GOaHbTLpYm8pJZeNxURL2Oqweqjg1S
zgYZCJqbtY+Tnbnf+9j1VX22Nfa9xK6CBYA9ePKlJiISqCMSMSBCokA3UhFrEolF
VmxHTNs230C7G5dhqXe3gRPr1LyE6sduW5oW2infc8Gcih59t6FHMKqATFazpHBL
Q9IOaiBr87bRYL/GC/KD3N5+5Wsp10AW6fZs3oA25obadPiry4a3Z2MDG76Al+NK
A1eClX8Ww/H5Cg5H040iYaFWwgaHW3xjZpvqPk1Lp/h+mEdfhW/b7n9mUb2OoJeR
iWbpYdnX7N1Bb4u2BvRV3onMMR0PD4Q4wxcXwY1+x8HL1JndAWiBWBc221iRLsOk
8AENvMbJcF8YtqHeUFG6+8UiuWs46rI3CpQ3oeVX6UpCf8/pERdUAHx7xsEwTUiN
s8VYSX4BecEWJRtKtyZTogaHrorU5iNaH6/1J8muqK2jG4JoEgTTTwAK4n2hJ8rt
OJx+w7VRgRqyqnE4++Hwq5ySnfYPPTyk1YhhQmmAri5TuzLoG2BiKa9zZR4RjkSa
KA5X1owmzI7QafU4EWxk9dDbMAJpQBtBQP2KS+YKTOYbGRcX9NQL4h4Kgn0IpIFn
kcopszULH3PFthFxrcjzVX0f3xALg0vyXNipOqoTvJEERIGtS2XC2n7xt/ZhUwFD
2qgKISGhQdxlN8/ePwh7Aof3Cm+0umlEVgMLGSyVdPdACwzyHbDcAfXvsV2l17CC
ENnn6YQPJY5l5+O3rO8aq4iILITwex6de3kSmT0470XYPGo1Abgggr9VuBA0T4wS
jj98SYm2uOoG7gfY014zS+d+ovBlH6+1NAnNA0iuYOLURTijkgUFvlE+NB4L7hNa
Bb6/O8GFmXwEudWOtXRBVruyEZuFhKjItkUoQNm4H/U71Z2XqCaWWGSSfFDNmajK
8yeR1OjgzttiHOuyXaXObcpQ9vYCYJ9v0pv2L6WuWqFOnfdHx+GQzD+4/diSSv3N
FOjkhqpTuBiakR8roK0ubFPm+9FR7L30LC4v3Fd+0bEpHrqa1sF1j7Oa1nPUbs7M
IZNLX/DrErHtpxvjTqicoUHXsNRpDeZnyP9LtrhBEP66YZhKAIcdzwbUtzrTE+KQ
DEMTm4vAh+F3+bDyGcvnnLOGtAWsO0Xm6etIlXKucH5rNj09ytuQOw+UlMTDbN4E
VPBrIuthBiMqpB8WBqABIt5W+tZ7LZYxzLVzlfGS0X157TA3pEPGdrdH2yJGHNFk
qcIrT+hXQYLbMCnBQnqnn0mxw8WWx3ZVYQsmUHW8cxhVhTHWmnTeD/pXUkLHG5kq
11YpguDDnToifjacUEUa2hwOrkRDDmLMyHin+JqorWBZgextUmzHN8T6JA/Av376
VI1VojdI9AwjjUvVkS+ivG5rOZc/zVgzB8I3c3KwJuhvLLHOHmyk4vlBr6p+k1Su
iFXQ0wdMI5eV8HUJRLY3DCo78MymqaealSiGA6dHKl08BW025txXhzG4JsVrsr8s
Ts5vnJeMbin1jwMkXToDEKDSpGov+QnnYI/w5agETcpm2ioxWPV/omyssXJKuvBg
ExrASyi89g8nmsPqgkfdfdTa6AdYnsVsvaWxAC5H4n+jcf4LdO3DrVRLgwKnBvDf
3Y4/rCDjvsoQU5Mn8v9xouZrHJtcDeBJmc57RJrNE6LpK+atgzyHbCYHlRO7L/vr
`protect END_PROTECTED
