`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yW4VIRiIahWJnzXn06kqWhVdG5W38qTA7/6HhGJ8TS8B0uerdnA4O1G1OJNEfwCW
4mfJkEKfUnwSfqTs2H0tu+Mp8VfGrOevAOqidHIrnG5YLX/G44yb9U9tlu3XO+Qn
vP6MoLeVc7xarSqK2l4Re6gHsshYA+SAcF8m+YGxurZ2M45h/A/IVfXQAXSL/kug
Hyln+us3p3fpyU/uK0G3PV1fiuUiheQyVE0uWeUxhLlc4vqiXmhmUi8iypN6xlkE
k6fUirmGh08j952c8D1z2AvgzJAudO5YU5APa2WiuOrmoQn2V/qtEoFUq0tl8er2
Q593s13EnwgBP81ANuUsNMw83F31P16emxmGl4VKl4BQoHgDBmMVQZJ7VhkJCXzC
2VcbIrjT+CE7jFeoUpOCajNROBy3OKenuWiGxJhj4CducjgBA5sRoWUbre8R/K/3
i2sYktKlexPSyAuw6PlWipG8Af0q620fx2unSiAT6Ii2rtmHn8zFSRdZNxL5JkRs
isTHeNIbWcMmG16L7hAaphcyVaJC77PS2fQRiUbIUBGduMJ0oA34dkzS5VtB+iOW
C5mKcZZo4KrTZgaCrPGNwVomz/jciQTBttEx28vFRPd2MWu6PH+4SokF39V06Xcc
BPfVo5iCfajE6dm/GEC8ZqW/lBSJs6TJfOMFb+VYfvJDljWOC+2T+QrEnKyW7rzy
fI6uNl2HIIk36+VSJVDsQjPDpZEj6UKBeUv2SC7czQxPeDL5EKZ0ImgkRbW0Wbvk
1Z/xHI8j/yldC9Nqpq6xIVJl3ThoMajFWqn6NcYBHOvUg5LYdVN2nDAEUro2x35q
XCP79z0WMUI9NnY9/bvQqsuLmN2c81wKqSzdkBUUgdE=
`protect END_PROTECTED
