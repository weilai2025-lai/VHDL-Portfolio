`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vktALp4AverGG3/rZaG7KwAnIUsCSJ43ltrEJN37XqN31edP1j3H96oo9gcWrveF
e+v3oq6RcKel+M574dEniX64ysPk1hqVUCwrCm+zNsZoEmh7obLrQdhCngHGLGWq
ZrO9A9QtrREltd3SDJKRZrr9j65exvfKduQUgVZE+lBiX6kwGJXjKpAYKe6gJrHT
aTMMJKAeStG57sPY2dSgYfmyFHi35QG8X2rFDLOia+YHvSjgy0UA7OFrXip/DaGJ
jA1COWRay2w3Q2cppfWIRwPLZBXhe5gScGqu9Wmr+pAYzLBzquTtFBHinManYz7h
zC3Ipxb/9zXDetIOL1wn4OQuO5xr8Xy3nFjCYUpvzRs3PGIuAtuon8FaA7jADl+f
lZ7G/Yw16fcwRSHhWtj8Xn4UeXNLtbYuV3gukmNuq//KMi5tpp+i7nyzr+EGeMjU
Dk4o/KPFyJ5KZE1EXfyc3XpQ9AD9DUtdYg0VxZn838nlehE6aOpnTMmJuxPVzpjo
sfok5FP5qxNjtROl+50N9Lj2ZVIqkkR2Pvu30jgzg0u2nblAaWiCr7eAr+1xO/AD
lnIYa0AFTWFI/GHPISZ+o1UVLVUU8FTQZFiN1QfA40DS89Rx2sxlkrKA4bYTR2UL
wdirPQ9g6mNSsqioVQAkaCf6EnBBMBwYOAH2kCv9DzYWGT7TFvo2uq8ZbAU0Y1LD
L/vx/Ca/UnJ1Zki3xxwWfqvg02M7cGjaX5g3wnZHuag=
`protect END_PROTECTED
