`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuZUotw5LziT4Zo1iUiFzwelB1v3hLgxR8V89e6q7HTNUozuiD3let3iObMQarKJ
aDHA0+ow9oOChXv39Yis30akDixoGLFRuaUVWrC8wPlds7YfUOwVCIF21LkQew5Y
cQZh9cBEsTO9zdiqqXkp5zdBd1PRR3nMx3kNHez9Gjs8is5Yk/l+46IpJ2iHKiQw
Lek+Bp0N6iGs0z9bAOlAMot618A51JVJAc1Onuw5YhwMX9HAO9HjsV01KWuhd/QI
OXt6Fd0mBkAOsH72KfbD8V/2gIpK+sgzj2Qk6e51mJcByGpQ27SXQbzYXTNC6SLE
cfXVPKAbniCrveo37FdkX99vgrNDmBSx9fl8F5TIMDA8aBVkd20EvxymakVmAYhF
9QIlPUQwp/g68ycZbje456NxmcyA5oEE3NBBG+G5w3W6SWMLCYAwPF0dWtsQfjE0
pc6akNGKG9hgBvbmrs9F/m1cv06etj7CFd3NrYtgSsq6tvyGpYCt6qBGN02qHwMu
sVxryO/GBNQvVVhhwpheeQr5W7xqdZlkFqfGCCFB5Ef4MfZYDyxdklA5upnkasNU
LvPSJBoLrC/URySa/OgBOlOPDefi+BNBZYDHe4xlLHbzcqpnTz3NVAUgncxJ8sHl
r0j16n46Rw4zRu2pO965Ne2wIimNb20OiXpnVQkEPFg5XBvby/tyo9rJKAS0/bgU
`protect END_PROTECTED
