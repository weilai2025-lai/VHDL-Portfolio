`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0nvHML/Is0bPCtsSfAULwTCDcFPCPian9pt1GPi+BzNhZdTQfU8aAsreK/rp9mcl
/RLCYYAD9j3Z9o/lF1qaiJRiS0hHE8tOw38IDUtbm99x58IoZ+/yCoOeXTX3itna
Kb9EG4RzDiWS6N1AAobbmhLAgFzy0+e8AY47xHxWgI8YyPxgl4R9BzNEAVYW1IJO
0c0UkIHdBfmO8DdptY6p76KImZ2GE4lOD7wiysgBaXUouYktCbYFW0F46xUzcJQ1
zQ1tH9Ye8aESJfHwg/yhbPoLrvf+GX7npSNVIl82NIdUwPjJY424ZHVecr/iCZme
wN/n50K2sX9FX1fVgsQrc8YUQQqVQLD4o/mxHrDxnFGeoWGpHrrfu4S/pFzqAEle
rdQshlcEk5KIcoDiEypdTX/OCIO4FHA+cpZ1VNweDAv16WTU8yRVqKl6C4yUK5QE
DbbPq0mMyK3VeHNxG3eAQe+qv8xJGUz2YHb4SRFIJ8/lWAjDiGmclAurUTOf/Lki
Y5/fGN7AYLpm7c8TRp8kxvCl5NJAgRsHSaVz1dVbgpguiF3LvFTfocICIC2Wohew
WrXHtNPX5AiMoCDcLdCrXxlYMmKPEm3oHGAITMVyuANBpGWpltsFrm1v6POeep8V
Z136P3IRELtmO0/X+IFoELgeoaJQUKyG+NNoC/IJDjS9Ktmpz7Ez7ASsqG4uCsYO
O5OQyHyYm2rNkCoOE+j3iuTp9EtiTXt6DGF8S/x+mbVMumFGlFp50bYOLzDt666h
pFCDA7mw5FQQjqZg+IV9LXryJdLPLt4K/er+SMEXc0erZQj+uJCTVhDiBRbcHlrW
f7BK4QTDqd1GN7WTK3vcePXEiG1z2m4q0F8OUo8qSceqdcg7WqG7zkyfhDzebE2C
r/7yKO68f+uD53tZnx2mqqC4gFvVzC9Ema/EO9ADYbOo3M4SbI59D/DfEkM3/WC7
9dEX2/Vt9+d+ii4rGrwgQtlux93wbtNjXbHDykOofcb8psGko74UchUKGV6huCak
dE8Te25enxQBSBttNpQRAxOqgxNdeOUrM0cU62CC9k0P/EeJ4y5C0ijtqEglQO+w
ERzOMgz/I8EifYOrNW6ChvkcMm3WpcryC26LHofI3ym5hXaf/cMOihxMRtLPWdu5
yD61B355yGqFZnr97tEQgL1SZaoQP5nOD4Efx+O9HruQn2fIpt4rLFAiq0TSEpwa
qKyzN/DbshPbNsLI2esOXCQpAFpAkFHuaw4Ckf9+lrQP8iiITMz3PIBWfq8Go8MX
aj8wRLnkhbFoipB97Rcxx9Y6UWDnTyrdfirhYMmghzcKeZ+z1dk4cZInV2z8hXtp
3A/eD3+HjeJPDt+DGVt6DkOG0DVn4b/iw1NbzCTpwkcu5dmzq0Wt60Afydrog3wr
bNGm67ER4xsuVwUcAabaGmMJkVOO8ZGn27ddGAA3NYJY69B8mE+vMH8IQptoWPSw
ffHSoWWP7+dP3c7/m95fp+QwieKA/9cQc7A98aKH/edy9gG2w7z9r57G8seNfYac
CRKhkpFBQil+AmRLL8SulNkEfIm8Y8AiDYyJie7qtYM9CLWrgWbryZoDLu8CLT4x
M07wLHxhQuAohZg/amBHLXqWo0vYoHmbfP4+J57H5xoq+0nb1mg2Tpkgy5Pakghm
In149/2/fyQoaorL7lsNAZaX+HSK/CLEM0Dt8O0nobmBDSWHJiNYeEXkmqqwjIdz
LPu3mYdhbzwAgYyZAE+GrlJjz6OwyPi0uRkFlVNze29P65Z56n+GuUKg6gkrgtiB
qGFHiyiGDK48fXq3qVcsYQFWgJA2lRr8BIs6bBtlbRfLJbv9Ne4fT4at7WldQZRd
jABRGium68EmnJ6Y8k2kNo3CeOpmYYVDIyzyiLHCvVNPUR3yD0CwjX8T+uk0up21
U3DYk1LgIG/7vHFPu/AzEZRS+GhOMbqneVAFA7XNAMNwTUZYukB2c4dBsQeROKU5
Vp902fumYvL9R+BNntfMeP9JhVTY29Hb6L2DhRGt4E3uk7aBQxPZdb0dkXkY7bdn
zjwCQu+5oxG7WUCCTWuXDJk5RgAsvtvUieAJ5X0OaaDWQrCKS8luLxTgDIYFnhc9
9BNS9M8S7Wpexljcwz9qY87OwaijEVaR9gjAzVvvOPSeYY5VyvS4ZZbb3wDwnUHL
kFFRKuC73bj6T+3uaJJh89asuyhuuTG9BhX/7PNx/HJJsrzEWlbrxbOqYznSTmWr
toPjweHp5Ix5uCB3JgMHnhjut+jhnDD6npLPxafd7sIpr/ha/ExSQZMoAPqvquib
quwuXHyYWf5rx/4VNddg89GA5PAMal0CcrRmf19B0OuCU5+SUj+yiTml81zTPXpl
XzpxkJtW135cK7v75yi0KVkVsT7dteqWmZB0BoXpA4LlfC/z042jxbZzWVgWp29t
`protect END_PROTECTED
