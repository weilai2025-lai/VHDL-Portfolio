`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4abpJlbs8/ofLdyp8xy38JFC+/xaXJw4G5Mr+Ofzx8GfJW9bVAoxDg8XJZRIJyYd
tCEfTz/QkWXpecCptDtzXhVlwy9ifa6J6gzMubh6BCyXEJHuerxM+T8IN5SiewLF
6VX12rEPjVhv5R/4GvdamUFuKHMUYRj7FVN4L19YHoZyqZJcOfaASUJfKqotHsa/
rcNGmh9ig/2RFFkCqbUTxk5bx0q/wBA1k8EZzDsFQ9h1fmEDc9ieX6vUjraPS0kh
ET/n7JhMiUupDzBGJlFhf8TfKO7NBaJzqVQ9745fLoO1ye25KQ+Pc1JaLiRVTM4K
Tx5QnWwO9ANnwIYr4rJPwcD8GJrwHfuJIYT+G//jVvoG5HwQpYjiF67bbTDhjDAa
PK5CXgFes6l5wE4m3Z2qx2SzFJF8k2zE2pvgGWzZ9VDcLqr8f28iu82/9zwWa3zo
950e6Cxiru1L8dPcUSNjEOcm14WGiKgaGKUZGQ8KNyHHN3MvQtl1Z0EaccZK0IPA
pvD3Lb5IMBzrJzC2ixLwRwS7LF31CwQ1mHMZdLgHoxTiNfOJLEhaOsLOYPuak6Qb
NQ6g4FSjOrX9bSIUSaAgsaJWiREnuecDA/B4q1xaoIC0JriCQD4p+l0vN8V34nF5
IEUCiDJ224WbNs5fZ5nO1OMzRSg2o3JxAfRlywDY92DmAD2GiTKJ7AbLswf9O2dI
09Pcx6PmrepUmCQJQrVtxQo9svfmmk1YJoMA5logkkKek2VTFK6zmfImoSac5CB1
g2A/ojxVJW1EBHayqhFL4lGnLRQNmQgq/xzkOXSeJvxOpazkpoWLex4fUjPWRXcP
fmSNfyEp6CSLz+uJI6IYOq8lBbqnvL4HBQYS67NcnaTfLLd/Juy0xgtysvxnomha
XxMD/6EB+n3MH320k1vyzt6IH848LYVtxVqD+TiWlLCCVkXf2pDwNWTfXwZDA9cA
//7FJu0F4TgpDgLH7d+Ca05/5R1iiItOjXda0CoXK99bV101Q49Kagl7aGDSJGHQ
KeW1HdTgkE8Ty9A00ZAaTja+l6rg132QAv5l3ieVynHyV16or2+iCTBF41S9CQ0z
F0h8TYMES104hC4noZxsUhVMFC0D9LSVxvYFqrsvPv6n3RjCUNyYmSN5MwlgjemX
LVBLgWqnAeYuHKXNUrWj55nU4xWO2Fw1wUosDf9VY5vxdjwYvXvQS9uIT+uNShNc
bmsGN23BKJ1P1wEvFcGSLShrH9We6AhLGoy69Fi3Wsf+K2qL7cLYITQuCVg4xzmw
vWZ0Q1aNViGHL4dlU+2oawOF0GAjZIgnMOdnDPuvGcKr49vLhLax9xb46nAWMU6B
1Wd5Oifik8K9UOK3NUJFCxayYy8UDkMHUEgyX00NG8zsarl8ErAWBW2GqVWjA98J
ebTV4cR9YW92+Erx9Psx8EwCSAtFEFYtC1e1PPX0Ty/qEVijAguLwArgX6/4aZ4I
pB4Arj+wlSAShlO/2NRPZmrFtBWFT3fmRuKz5wVWBiftPcdHaM5O4/PFpJv21w17
Z6q+Ml4u/tXAtLY0pasy4g6L7VPI2By45RYxBj4vK9hMbT6zbjp2YNV8CdANL/tN
p/GjxJ/B3yCgPMaDxBtDhbo2aeN4M+A4x+hSxyFgxAMKftPuDLSShSkA+3Ugi/zq
mCa3EDeSzSsCuluRNq4zk3Dq8CQHOd4zHjbwf+JluQU6aQgLsyUxSVBp8yz6cOhV
+0Mhkrr3CfS1m7JzcXPqjEptSFGDK5ETHcKIN9fkI4sFhZIj2b8FgdPY21OWeKb2
6YZn6TgYpRUg5meQ5OA/lGR0qKMhyraNnmFII/E0QZIf3AbU+d6XN12dHKzT/n2U
YGh728WDgpIPD1EnLesagyNr4o5Ka2JHYj403qsLjpbu+wbN63ADG3325UBIavzj
X50Yj0o6W6/UjpwhGH7fzreT7x0SUJhfnGxIM6C3K1OS+l/6Eq5eqmAmXDR9Bjlr
yL7w5x72SMUTyWQ9ioFP8/W1LFhljx7J8LahmBOqrhyB/766pEdqfu+OX70zT6k6
WlLwbXYl9UvU7M4uFZQX3XD4rs+bhIeDlDUe1B+wSYmVnJfiptiY6z5sN3jBx+Nk
TeD9SXMYuRRK/elf9300RV06r4ykoS5t+IvG8FecOclRsUSeV7/vQAUGRc6xvBUR
sjI5MNhylSkezvBwDtsBgnkdyJBNT9wFGsNluqeo8fcNdhTOTadwGNh3KEbBV28G
wOeQfsBTfg9d8i7wpOWzP5mzU4xwj8WO5MDyFPqzMD+3lZ9GIWfjIJ3+PfuLKlBJ
YRDlVzfI5sHej4Qdo0Lp2co0iUI9UQgtg879Pr2MAZf6HZH1H8/b7SXx1digtki+
/lHLt6toqZY4fFDJb3ypGP2j8ev7GardL/jIh+btiD8M3br0hDShgGwgPB1dmgvF
RaOCLf3wz5h2tQPHV/BPVqsDM1nm2FhhRNDgbb5ZO5Hy52FE8zeRjFSefzcooRiX
KAd5aVyk7JaiMY/7RqIxIKH/+chKQ0LXt+pL+YVVwV5sofII0RnOh8K+XzZneAkO
VHitx4szEeE5FdMh27VjIWkT0SdHPy7rE9xeTRwr1EtdABbvXrpQ5UcppbiWbQ+6
ERnpVdvt+xS9OussUtrSARzYZwfLDivYmFangWD8F+DZHgegoIm+lkD+MLEtmfYV
r3CqlP9txZlIif3fYCxvdSxyOXQ3lnnARWoDW4guWPzBvOYe22mtukZpXEjiUKvE
pIgnDIH8+eIlxfoLrG2/RV+zhGIgMkW3OqH19DdM0Io4xhMdyyQ5keEoQ58mYqkP
aJH4SGrNdxqbc8cPjKkhn5lr8x+XATPadp2pa6VSRiemsWY780uazAZCMq3oKOSK
StayB5GbIQD6cMd2TjduX1DgIYAo/Bz3DeETa795U0s0wbHGauNUl0vWbHySk78d
bAEIN33GU3dRQE8d61Y829/RTvUIceJDS2rEXfoO0/w7qXf+8MImI+NqVOzLz7kq
IgLf+iDQ/LBQY2wSK/14QKtslYxYf3sbnxUpAPGuI1K9q6CIy0uNezcM/NZmYVxi
vW/230S0Wc0R3ItTlvirYlabUmm6SFdH4tcUjo5U8bCkYZDzc2dubM7SJ54hEsmS
yzzpk/UwKiCZVpx73v8l3kKmC684Z79+dQJsjnKVndtWUgWTJG6l/Ai6EqyNBYbv
pb2UC2C3qwjZyyIdPMK8PdruWnpn2I+yJRyVeZdGU7KRXlwtyw0b9vQ3Ltv6fKbV
kasOS/F9Opzbn+rAaZzdacaqGCcZGuX7qQOCvzrUw/jMRwyj4KhXKnTiqZztNx+A
TLp6+5Klm0PvQ0u3uKlWtrp+NdL5XtIRMz2JdcNCiPkw+kz56dOhIntGioYshaHB
UsFAM04oTLOjLUHvH8QQvMa+cnXw7GFS7jeCciDAebkWhH5qcyhO7Xnj5IlWJLxg
ELHmQ9EHkKMoeDvoOkozZkWPCSTmpiLm0zDgc7f4MAbYuU2plXLv4O4TKgmbjqGn
`protect END_PROTECTED
