`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uToEmSQxwi6aguAbdyVTsdNkdFti6Pwi55+Qq7Mgb/SgQ0SBm9g+ZCW4F17CToK0
bhzZPoXxFx2bTsi+1Irbczi2mVyGepwortTrv/8DcI6xIeIKOpCVO+dE1lEmUoCH
UlQ9H7XkLzSMldBnG22ITLUDk4BVdLvYGx1tSOXb7YxOTS8BQUcNGFXxistBK9Fx
fCYCHM65edUGcA1PjB/pnCYLesiMl2PLia4Ml7VWyw5FjjNKEmiVgYALBkqIHr0j
1FU88cogGTYAXtR4cfaBYv1vECpzlc2n9MXnmJBKDYeL6KlSVhp0u02mCy1MLjAG
8+ApJ/fQjpcHA99FNsfFNx5TACAbo14XJ+xX5j5RTSTU9dJvzLkvezezHMe2Spnt
`protect END_PROTECTED
