`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Et2VTRb1zsGo54f+VctdnVtM3uRcGT3ytHlbKRIS2hum+vpcLNad4A1aj+sTpilL
GNBDck/Ae+4F93LpX7GYePgsuEJ0Zcg7hamZlazjE3zbcbLoJ+OaOTpq0adZ4sdH
n8kaQJ64nFIxyLw6AoXd7cwtsQ7RQS1SkIAFc1dGdc+QC9/1JquoynmFqsYRUMsJ
Q4EbfocEb3wkqI0dJOkHmZzC6Kxs/0C19iJzUHKPYuo7NPqBUAmQQfg+1LtXVafU
3FwumgUakJje1lCuVnkk4btuyV2zA67xnn5pTIzK2WWpcSe4g4+xICW62CbbCVEw
82DvxqXDA0grPsvv1ylnEans7A/Q89f0dD04uz51+i9r3GREPAKcn2WwifM/Douw
gV5E34VSAZgFlmppPhVWwDVQ4V2s1NE/rJb+4nJvejQ6RbUlpJ9oVVjHdNSkdEXy
n9sGupPSrFlSbGolrMW+2jllAUcLR7cXXJTwbY2Ex1kc2+sdyXFl21dNkJVrKFtk
5/TQhAfvLTfOB5G0l0K3nWODaPpRwVuvFZtcOn/Gb9elagcMPIo98bAxU37a+8kZ
GFsEI4J02zA9swePn/62ediTB9hP7XMFittlI+lBsFJajE5M6h0fuxgOagke0tCw
CLiFkQ3rqlR9HviRRJ6f8esmZQ3o7+NXZ5GD/c0GJHDRter5Ehj1us0EU/vPTE2+
MVx57Vt4S5D9UEPg0xnsTrBn3jYXQHn82U+TkJfsE7qnZ/LfEHKHYlBXOLuh0pnu
V5ZSHd7CovY6Em4i4tTe1/BHM1mLatcnikUga7m2OukhidPgGH1L8W5AVHHgP5cm
CulXg3bhc1Fwnuabh4ZM/WXfE1O98+1x54B9FEHoxAlWtaefLcVb373GgNVx3XAS
OySLqT5du2pKcRm1owoAFAyVWsNX2y1DfazTApvlh1UEVOcJkI0Su4dHTQuwK10u
KhFeaeKEHqVGeJU7jBbmh3RsyP9Y52i9wpFe6TWEDPONAfJWors8mVPCNvg2OunU
ovjmftQE6X7WP6B9MnCpiOBtoxsrV6hYK+fTLSBOKdKtvHTD9B3jM4PtFiq/ofZE
BaqCuG1D6u8od7Qsy1mNqhWTFqSez0gGRsWC0B28VO6NiqNUqooTMc4S4QLCKVlQ
ied2Zkcjw6/PKIWZsNMvPwULBFgp/B5K4Akw2KJGQH0wLxv1lBlkoY2VOEXZHZ2d
rzx26Yag5TIgCIAiLiWOgyHAYcCicjwsIQ4/cTxjwLgdFPL8g19B8QjP4olgNLc2
5ZOVocaisULGfbDnBD1UGceZhNFqwDn0Lvu35AgCiUpXqlFZlwC6rXss7Fi+Pp4A
nfPbxjFFFe8mTRmr2ZY4Vre3+abj72ee0VI8VspMm/BMdRLChh/GGP1dSTFASyLt
bzY8X4biuMV2RPMCZ9JpReh7KZ8LeN9znEKzyxeImDinSHTw/wYSSOC0iLZp6tt7
wk7akcywzZhjKjJcEhHAEx5I85zR0Vn8P3qM8N+XYwnyHmrqg28n+DPbYIkwvNL4
HHiNRq2W/1vHvS7Jm1osMTCURPymdn5J9s9FGM2Sb8BCz88mZFdK+izFrO3cXXUB
Q7WwIUMUn2B2DVAjDzW09JVreNUGiVOAMh5qQHbpVuw6rtrHYaZ8PR1o05qon8TX
y7xoLGueSOX8cxYwShji2xKbCCkhTbNXgKArsWEuaZkum58lFw38lTCk7fG0eE0X
PLwCzbESpVBOxf7Z7xa1JhlJOH0v0qQDHaAublpTbWZLpFvUrEdV5Rba+ueygudD
0hvv3y+ThFbQ6iTTzUmGpvxsvYpY/bW7aEDwlnBMitEJIxJfNCkw2wJMLms556gQ
11wt3p9whcVvEoB2E1BsKsDeDyjs9BAXEI+2fHLyQpSgQcjlE0CqChJntimjbG3n
O8YQTCJpyzVOIcq9xp2imb4Z0Or+h0DPNaO7VHdYYKSHMm0s0HTgaQMgOAGqR2xS
yG7h/VH0RNzW7WH0yo5Eza/VH3qYj/9klHuu4OPfbLt8uwJYa/KA/u+duYpvzhyN
/ocTee5TL08xzcgGjb+rOONtuP/XorvsGRLxHMB3q74lHRswL5Qeex4Pq9PwTURD
eP1luXbqYDJhJMo8QW3r86oMUERxYgUpX9z2bqWVA0a2RBsRxsdeAfVueDSfZw98
wjUTcCjnFpaQTGsQuEuk2o3jPyxsx/h59D9foTgFcC/G8rlAg6aWgmAOzBLDHKgv
SKz2tjCFBvfb7W9bMbvJV6ajf9uy4zUd5s/ooKF1wAf743ddC2NBVKQdqpxjXvuH
cazJyhTuhzUXUya6j+2xRm+qmwv464eLyTgl81hRBZ5DCr2KG1XzwFzBodUy0ycV
wfMouK0YpP5Ofu32SxJD//SrNYpmmJA7q4X2Im6qoTmHZngpWBChBNZ/2gbNPnXn
r4sJUDQrgkvYCqe4zxjRwCU9i5Kvx2ovKbqscUAJk25hTKrZqVBjm5y/QoPNwrQ6
yVv2QGIgbe112oYTe+zEKvEAM/ABzoIcbf28ylIbx9143BKJxWvcXclcBIRXLthn
1GGziQzx1AvGe52UsZam/tDyNYWuCbNNjtJa9fj/h0wDzmrArqfYLMjfpw1qDpRz
tN3DgPKpLnEqU25r0FzlOKkytHywwFZ1qYMTPToZ1uqUpS2D0trkO87KXnqYfrtW
O/ISEio/oAH6dwL0aSf0GM1Kv3qYCYLjlkqd2GyLpKKw99Ck5kZ2zqOvtkO1rVKF
XJTbecoU86L8fF6V7kT/TC9KTn7iixFhDNddz18rqZR8ufVYXR8eXe2KigjCmYJ0
Q+Xk9sTpaJgHwrgHHloD5ktc4UxuX6hoRY9HfmhfGDL1s+VE8s+PxAWtpDdDxSh0
Oh0UMIPaDPoovENPVEpGMd7Pp/1zW2S6JKBtiNLbIF4nSXYJtQ9i3E8wWwpDELQt
RZBNSdeH/UUnwoOxTsXlsfdiQdglUp35Vxa4qEV2G01KcLDtT7l4LYw8HBWFLn39
qz+E0LoOH3pFlqiSStQ81ThQab+DEuqfC8Bx20cB25t8GPJUf59ZNUIoFxrXy+2W
Bso0nMsdJ2Sy4D7SjxkgN9H86Y5rR/qdA/8yofF4M2TNqNMI1WaOPV9UJa13sejo
eOxbwpeghQlu5VcgrH6r0OPZTWxZX8rnx7nqAkXmx/vFduGleRSEEp8lRqj3NHDQ
HT33pXAMplfnHxlyK1xcWR+o42Yn/72EIhl8eGY2M8ofZOzjw/avTdmvdm1eQyuU
cFUS5VDGN4kCDMhRHi1JhlADWnuEUhzmYgR7viWPr5K3lqbBhVS/KMadtOVU93vy
zN6xOiAen+eABfQUd7OUVtvLD6IrJqNlUTBGeoz2Pt6Hqsv68w1XyDODyrRbTTHI
S+su9xChQ/SjjOYK2UDbUtd4xNBvICNF/HcbYNKQMnhmvdT7snXiHmtkCQIIYTWb
L02y1vzLprLMgWIvv/PSg+5m+avakRVAVDmLMfjomBG2edCf39cMCEs8jV54kYk3
lPNkyD0E7bdWHay1Wlt1VuBYsNPk57eSnhJVst3nVKAjZ/NWH2yBzKkXoibxBEO8
zrIFeBjIiDuYAS/dP2TikyMtdvddRRS4BY0WRbvNupeHA/yXxKP2aPqNtq/N4ton
XI5kt7A8jyrJ6Nog+y1OB7tReV5ZQwfoSKr+ksfxmP5+7MRBWN+/Lxe9YXnEE+wL
X328TprltqVyQRei98J0S7nU0TFcfXkHT3ip7sUR0RxXYxPdrlzmZfebidyzjleH
fd/Sh/x8sb/whAG4tgGF3YpGfT69IuaMJ65rtc8+Ka979s1a//2ctPnG4PyuKIPF
CMSK8pO58XAJ5tZWaeSFCH+rDGgICZcFIxKvs0LMsUItn0Se9fIgo4qNOZHwmaig
OOrv8j4/hEox71XQAGneLEB5m0/ZHAMVtjS8OUWUpLRYAA/57wZWlH87YlGP2Ars
ZvDoWLLEc1SVbaHZmzrXNdrvodGG2ZRE6zxrpFCK65iDHxA4JQcKbRwpZSF+FCJK
5zz4rPJYno5uZ7Ob4owJRGA6mBmABlM0GE0CyKzStSq/o4cNU4uNjNtoUnN1W87G
EhN5xlDOqq6Iih0z24p024SARy6ToQV8GvirDxQIaGRoXaztTfM30AGL23u8BNwa
yX5iE/TN0ZATashqSJj0uwqpmHzgpSW2LCx3y8n3fHuvufwFpJaSQxG7tBnxLuLS
3s1/rBpbvyjp0anwUwDxB3HSSu/KVqmNIrOGuvk9s5a4JDVjxfU/c/xE9H8xjQQV
RTK2rrPT5DQ1PQCS8DzQlJPa9VOg/BKZLKW+EJSkQ7iOpduIBPkB6S/8LoJcv/h8
diJF+z0paWu7q1ASgbt0hvhAa23pHhV971gHJy5Ek7DBMIIFD4zDsHo30Vp4lxND
Tj6YHIdDefy8nc5MYdpFsTocrnLnuLiBxdTtbNHlpLAV2cA2X5lsF/yNHHhojS3w
DZkHEKh1YyDQyVlVT0gATF8xjCap4KHQHBo/EhyR111jS9nUOTmsz6Q5THj+qUs7
c+0Vky80PcZg8viNqruQqrIBvrITXqxjuFUuoa2NcT8sGetUq3PGDTE53+ZdtPG4
AtS2wI13NmvZ7+8a1JHdnUaNX3ze4m0buRjBD/d9HJBqccL7csRwrCLdiBmg105u
nzClqaHuJ0NC5wYUmX9RPDcdL24l0im7/xam/2TzhHY+cUAcOzn5nOOT8SznfE5T
L4bTyRhJ4DVIgtHZwNi77ZscRej+XArgIqK+XTfj3uNt+00vH3MMGAhIMb36wZw+
lT+jgZcLycX2XZOS1ObHMvD6nQp+S8FEarboCd77Z2nkZAb4XODXyoHND2S5hELC
Aykvck918z315BoXlhKhOxHooPW9JoqQoi988XQ8PAapkmFO3fUK0Ti7Iv7dSaL1
wD7vJIEKlAvIOxBuTBj7VQ8taCb6Rzi8b8lJRN4hvu3DuQP0tyF28dBwIJVrnxdn
u/l9yP6h8GyRTVXVE59oXlwnpb1ljiXgXYjRE3mQhVT6n0psj9wxDCa49U3Fjqm6
l1B6IUYtR678WLwQPJqAIR17OnpzoBW4ViBIWt7pXI4g+ZonPsSfaeLs2OwPlA77
dra5y9kqY6U3iWSZKpajqQf8nPIXBErgUe5iKBEwie58eyoOXkLHtw+kwGGyIiX3
beAjhBnkudcKiTjbtCBpzAdJXBIzJPgbPXi1FgNEpPxVy8s8GXa8yfYmXrUAdLrx
edNMRZ05wk2IBIm46SbZ0A==
`protect END_PROTECTED
