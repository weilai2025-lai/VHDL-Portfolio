`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4SPcvHP9/VkEUl8cMirry/21Y1K8BlLGjFn0UMg5fSdwV/+RlcMhDbJW+49zfDIv
gH8KBvoLwQa/6QN+56zzLf0yIfpBZ4CvCTBEJoE5kKJnjqW3LJJPfpYV0Fb5+4om
GcqngfO8f7CF6uvuUI7iA1lp/ywqeKVqFkZQjULr8HndTTsh+fhoh6MtmB94/MSR
LQSCVHqEozOF9ZPYGBRfjO7ItYp+gJBaLN/B2ct9e1fgt1MDuXWIqTFCkEVM5wO0
JLVkIEG5gTCGnxOFXxX4bQ/RDH3py3liqGFCQDaCRecRukGQR/xYYnY35FIkjEqk
FvqKbZcZV5h4cyAMzTxyj/Odf9aLd7XPFns9RYMgNgkmFcBHU8u31ZOU2R0Fp7F/
Cvo2JCsFlnXBEHQd1YlEGmzJYTjSWeUWYjnw7ULKVma9wUiDdFhekYUmNrXS9n1C
eKEanT8JKQY1ceo1AGPR+QXp6vIo8cU+POJtqyZm3bNQH3h53nLUlOikwMtPOn3T
WPWG4shGDj4QcxwAJRJGpmI/TIh110g/ITYLfjoK4tX57Z3XXYE70/BzBPZKjJMV
krbTTfJPjyNO16E+g7YmvNWnUB/kiDqobgJf7pRaiXxvA/jlZ1D/5NRtysr/9SdT
jB+8qTWojEAi4MyRjUib1waVtyZFObIyGnP4DkFmU326qRz89yUf4YCrVjbzAzQ1
RH1a0ARu04Go6jX8yDfjeVgNhskg29JkCDJl/r73nAiVtGF2JmxNjNOD9KZ15Wqd
5ARXPvxbRuujBaoKqkXewNWlGc/ZOj24Ymq/ByqiIfHH1rxhckLXs6oKCDxhoOsL
8yEhxFwsvyzqAD/nqw8IE81nO2Lht4Z8NoThfqJPfiG3uuFHGRmiT1KslTqPY1AM
tXJ/tbyjI2h37xZQNZftIMCxR7zUil7r4OOgnpDR9LWI46nMjsLsD3XmEy1gsm7k
`protect END_PROTECTED
