`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k2/pFTQuHGNZOUU3XCGOttHRDqkmIru8WmmpqrgnULB3HHZa47F+oZ12uf67xso0
FPzNZdTHV1KHUobGHBVaeehIJFTadR3a88R2fBrTlV/kOrXocRx8WohlNSwomRxc
zFJ3r8Z+Uaav8WmZV3qVQa1V7gZ0rGk/sM4w7FiMZ51LZEsDp1o3KHAG030y6anl
U9eTni8Jh2lS/aOBIiZghN9Y5K3AgiBNA/r7IoKJEwVgumiHSr2pIJFkIuBLcdSj
etzOyImcd9/8ouGfzBXdIfLa7Th0+y3sMbDZYt4b2tqP4ijPOJaE3PY7AKL3vSMI
5foLnRE+blA1RdcnzlqwPWebSHtUczhaylbd9jolf0M+fBCwF1ERX3UCCZIfIyXs
JEDDOHvsPZYDqJqZd7ATmOi7AmLlBSq0dRrsr2Gs4wjFo7wPqgTJL+oeCbHjVKhl
g7wkqLfq+tYvduWfO4wxJD/3HqWDQgKDB42uRAWXBtx42shvUEj70UkW76xT7FbR
6zp0WSp9jUHVbM61qf15hwEBlfpfQP4dLcWg6yHZ2jWxp6A/pzF0A9pHPVHooq69
MuOOthTs2I4ONVbT9b96Kg==
`protect END_PROTECTED
