`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0LmD2vWQMRPgD6S5WwCkl6x8BmZ3YR8pOJi0Vjx261nnrluLHouPsSKB1SSmmvL
njJh7hdR8idJ7TgOkyC59YIH4QPMfjOeNuSqcHfktkQIR2yX9jmPV0bz6dMsr3YK
9JkjEGp24m37RIQx5lz7t6Wm6LThe3OVe9G1t+kbUdh30DPr/z4FsyVicRD7+Zl/
IFp/5OmOlLFMVNsJayOWi8oiAoLQUZJxhZHZhIykYZYPELUdu/3gIae6khLW9REp
7USlLwyAwrYW+VwrXMF8+DeovM2/Y/C35rw2mi4s9mLWK1gA6V0Sd5WhBo2K67mm
tw97Mz3eOV1wELN7zeEtL9e73WIRcQEqQCESfZhP1tR1yNqk91rNVrHLpXVT21ng
R583vcTxs5mmpOCrOaZs/yBbSTM8AlWwjR9hTOID45JRVJ+790i2GCqu11c0sej+
tB4fFSCwxzfwzf2cjgmJEefcbkIcO5RrVyvKLkkTV3chiZ7XI6XUXmh/Y4RxUvTi
J/yL1yeaB6uCaVDh6+sBWcJkv2W4isp1nEXb1MCJuyYoN7chQZZB13sOZOqSp9Dd
VuuBfHecqovFAuKkOeeus6wbuBTMOJi4BWRMLNGaKS3T+ikvy198n1NHOapw7sWc
rQ04rnPXiunaLazdmDtAopQtvRQM+eY30Q5AjzfvlNbAgxzYhQXkw3CpqhQ3oQqe
d82NVd8Br7tc5hnCArZXSjWGlI2WZruO+dMe/4PwafgATMAwqISnvbetbVaJcUfc
P+69t2sINu+8BZ6NaG7qpxcykkQIr1OTFiQWeog66OAsgTDixBtiBt6ibBQVcnK8
1kb1EI/CgiSP0YtowM1kam5I+VrkyGXCVQ9RmZcSJgTUriCSHg4gzjnr78qFQUPs
OwH29UgDtvnW67e8rI+uvvz4RmUSky3CDMeRkzDubOejCJ8DNWjwZnS0dx7Yafs5
ZKT1PkMzRwGGmB2uB+QlFpqqCziKQSV8CI0wuwSMoA2XVbP/H3xHhGlKsjZ0mmSO
jFo4r2IR90s+mELW8VdpgIDpkMMSy/LNkQ7JiGgFDxL85GAu4w19PDAjokPcNdjy
T2B6HO262ztUCnk4X3xxLpvgUFNuN7SQU8ThfNGz8il+ffVdfU3SjxCDd1TmbkjO
aG1iJ7QMRHldjuo7owEpsCjhBSYP0NLDtPsHZhA0v47LOoJhmvYWKaiPIiVbIWrs
Avq6boH2BlGO+zAFXFd08W9SbRIiA2E18KDqaFotNnaxrlYCzUu/KwsKpiaa5ONM
GsHoc9vIGx/uVlIDiYKn72/RzgmFEooX9+N9Cy7daUPi+qfNkTzwnta7HZHvOcQf
aUJ6Grn6evfKVbrHQuPHsnHJZmwN8B+78oyL7BRX5tzTkn6DQI+eOKlbF+unoO1+
zmCknkwEGIvW4neDXbfu6XHD5UiwLkQZCb2eu7vps2RGtR44nj3nvBa1Kta5L0zH
k6N6VnqDC0ZtWzbHVcxVDNjcYc1sEC/okRvhS5CbfxnDC+w9+sf0eLSGHolZFgag
9lbnQ3ZwJnHU0yY0n1rHSzaZAtgcwA3uSxiIGrx1ke5RlhDZD2WY53Ev8p3/zXFT
ENVdZ81mGfuGAAtoUORU1qwqZsd816p7FUDdh/uzkrRxO1IP1Rvu8FrpMXlJsSIX
f/7FJjnUcRM4L9PlYbvH0xkR4F2gqR0ygy9e+v6JVN5GBON5EJZzTPLpqU9znU6V
XkHYPftDpetwkOL07kJNfCmPu5hgwpij2bMEGX+daYELznHRCo6+KbkwRw4MRM2Q
2WBDN/ree0tX786mdveU5rOqBbdQdPRDOUju+1GUZK/mF0Q8ZLStKPDaYJknoMxe
2fyaTt0GcQbp80x23zl+7zSw1zEGkSHdFDJgEriSy4qRXnJCI8JxhPWJ2p/tZ8oH
JmB0cniTc3Xbm8lM7XBK9MiEOr44mSep98xu6M8ZgUYuBADn+YRv2lHMgLQCu/w4
T8FnrtoNs9KiuZQsfi9zeFXu/k3E7MmV0Ob2ju7+Q+mtgWogw0BewPc7JpDMSSY1
kvjfOwoS3GG5IS3E63AYtNXCjVbAK2jNH8FLxqQbKtWXjDzzzWA+TIfEjpnyRmTd
K/duyQrcWcW3163JDae3M8uRFMifKejYRqSvXH3Vot94/RKILEXWp2qu4el+rzf4
Sxhgsblh6mEmBzBvDOH0ZYRTIbzmY2Ct+GV1vbkqWO0t4BGhuQytlfEyGU+uz1qI
xytgvznjPdkcb0blGwu84VzVnNMF1okjxLjS4fd80AQF5yy+MFGJy59FCsr/yOsK
8QVC9MUxnsVpOWMAzWFOcy22o3McY8hEvJUalZkdaw3f8onYsCWX+2yawYoxrNkB
Zy9s2fh7+AVsMZgtMp8rFaTe6BpLIALrlpoXhqPdeAs67NgghGRgcofamq4Spio6
+MR2DeOl/XMpRTE9byePanwtJZr2mF2VPYsY43oaysC7r72tZ/9K6AbYA/Y8NpCc
mkeumsm8G8YUDWzIEZOFE1ltLYPwRrv2cI355z+sECAc9t5/u40peXnD29W4bMiQ
2iFBBVkYslGWkPyqtTlIsu7jSRSMkEUgMemoz6KoM7BSi0HpAuXywmL0E+Buh8nz
UACTs2lxxKqhY9ZcbKbKYAS+UwyKvC8S6HO8aspnMy3CRnGKAWSVn2ewoshhHt09
riTU/1dMUcOTDgy/4v3jxlh4zvUgHAikDR3225VyRVS/12ImtkVXU2L9lqkhq3Nh
lY306JAu4YjmWM+DczzLerVp3vUlyzXQ9J3MCZvh2Tx3YOqEpgF/DYEXHkkkUDXJ
VfVkMEERQgFiBoB7QNm9SCCQtTs5BygByQTjTWSFZNEj0LC2uNuI8hEUtnFGSmUF
WLVvbOnUx19YK3J0eSSb2dmf6UQbpSmlNU5RocnDkTfe528MRsYNrVrrtrO8aY9Q
g5ogpyuOK/RhEyxCsYg2KTslukIOfueb/gamqokePHVyx+VTIwzuwGG5QNM/WDY+
yx7M1qPE8vAUyXRBq5wgBaIR7ixrN9c3P3bVT+brmAL9wNfeO5a+hRTwuGullytu
YrWV36Tt8cIcv5NC84oGTYDK5JhcL/341v4lHwJOdP4AFPYnuqwiOc83Oq8cFlhV
6nYus+eLryL4Bz0+14vs/W39iKgwEEoX41jJU8/OgaOMVoal3OC7o9jKRhm4YMSw
iYw5DP0gIIZKEYu1UziAKENLcc1Wof271zQIzvx4E/1qP7AOJl32h+4LXJ5pH/wr
NSwk6WkSJUcvPZyc0ky+xeHFR21wnyobF5rZravZkf//bIIfc6csXGm3DIWzZePT
TCKnOarqzOTWpx0h/zHiFshNjfariq5bwTbxDYBqMTXvw6GzjXt/4wvsqnKxmy+n
aFiZg1JKEkerAV8LabG2XLgN3kT4B2yotx4a0Gxz93P8u9mgZ+e8iqXToKBxHcMw
Nw4ePPuyerjkqkqPWYd+YIzZusUdFfhRX9QcbMgITA3gR0ItP3pd3N70c4DVFkRO
`protect END_PROTECTED
