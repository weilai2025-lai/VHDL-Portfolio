`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOCYEMB7qfteUFeoNV2jdPj76ghYO8TLOalSGVQFNNYeRTr0w94LfyfvohwrS5Gs
J0hWdxMt7N4OXoybuD6I4atqzYMncagTPjp7Bg4O+jbGHdmlp65xPLscGPCbom17
v9Q+LOqrql1V+LUAev7mjosex9kWbmeAbLg6ZkoL1YP44JvQhLecppiwRG18ZVd4
j9xCne9gkMCB1C3gSkZ8w/PHd7G5x2mtJkITBIh6PuAdKxG0oUNON6bmnyOWxOh8
Q8eATwhEJKDY8cDsiR6F/O/yx+FJGqmf5wmXYl6z0cWAtWMDT2X9kRuYr1q+0Zkc
HEQeYI4yuQrWb6RLjmceZG1TQIUrMdSw4b6tTMNHGMX1pKifWF6o7kVA5WpEF8yb
RUc3NrcBrY9b4ncXK64cTnobdIttyiet0R9XMzpBQBZ9ozX0IV+zptB8NMGbSfN7
n6X8VvIhwJH9lYEWzCq3dYRdwWWaC6/sZ0+cfsQl1lmtxHgcbhT17hVPsBn4uU/5
jBCxoxxBPKImfToQCCSSy528FSD52t2g/JxHuE4UXEF3uRnbU7i/d6IgIOXUc12R
eFb1ZBjXrkwuHnWj+Hqh2WhlaT1QSHxesndotoJWtv/YRkLjXs11uUwdvp0qbP/5
DTLOpG9XGxVd75lNIqYNTEWAIY+pxNzCJx99PNWLKxCT32vhZxtjiZKlI3+I4FxD
imlrHUNldcd/KUULOiNJcR8eByBm0nXmDdHiLZQ4MAkMds3EFsv4JviiJp92KGci
5GLd99Or8pArHEJIohIegwbkpEzmEqGZO3BbHt0KEt/NwoB9V/Qihb+JpUA4gvr+
PHJ0TqMP7OQiV9opVrnJxPoqcPK5qxdBtknnJQcajKUx3wFOK8t4xsoOvYWAxgTD
P9xBSjWzuzC1jUKqdvlBZihaGDaErKLgtlvZOiKWM3A30RM6wgLqmN/qrn70TAsr
1mIUCTL3kIRQStNMKFsAo2I+vmYVgNrh2jtEu7ynKw5dPVKBZApaPklPZ/uxaCNG
vHUleSaqlZ7hR0aADrh9a0ptBWCqzWfSflUxvnrIrODz8Cno/OhpQ6cRvevGVCrb
vNPtC23vvD6Ftow2ZCDiWlI8AZlVcZxxoHSoK//FUebjIIsAGc1HELI33YecsXzp
q3JnIw1gSZ5gr4J4q0tT96bktWMuBhnW2DotLHGga6IFlYJHP6g/NOxnAGLwMyzy
1VZkfkbQzIXUBrIoXE7iofz6oHsLC//9nsKT7aP7QSm9PaubMRmkyWnX/uv3toKU
t3ypFJTWso99Oe0r9kEWHvHiL3UyhfBAX+Gf+0Bo2mJJHTn3PXKjAWy8fSamaiMy
6p2emNaRnu30znEHtLNTdFDBuFAyNT7Eo9WviNXlWgS7RIgt7LjdxYZTbFmgsL/M
8BXCsKWsCxkmABPEolmBSm45rGmnaSavmDon0m8TYwfCuf/MYfeoNO0hyp3lyM6C
1E2KhHlOrRYALBUpn7JXqEMIq81w7N4P088KYMImQoW6sS6wgn0nnV20ZVype8mD
xsKc+Sgn5vNBnbcbvhREPPibKjYikRc4VyetH+OeZ0wJpRw6yxgRdVnykOqIzdFe
VBOMpf7rbPYqWZW9/gmIs6rEHTIP2jugpZjlZEbsx9c=
`protect END_PROTECTED
