`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0WFPBevCqkiRoww4AxGb4eJsp/agj0GvsaMyi+w8GtgqUNzeCcTH4LoJ536yPLM
SrIz5YWkvCxd63kKL90wGvhiDMl5pP5sXQAwchnAsj3oSzKrJA4zxjDlEvB5cT5Z
JX+sJqKr225S8MC82R0lKcxbHNuUGbZ379R9kl8Svpope5wxPSnCzqvpEFlgu2bB
NP7WM+0mccMpHD3wHc1hLph2cYXtCowDAmZdPpfIJWRKoXy6rUc8IUc46bZC6FJP
kDQ724Douaxv1UaEdc5iHIwh9xALwhPpoEMX+xy89D5igGsfD0zdsjAzhCpvCXJM
XLpcKSGgrlql8GEzqmYQw9YS4RcvvoWzAjMV+WgFBs/NGaUvn0xi1SAIs163YqQM
azuwnyytjRTKNxH5KulBe1amRcSZaNjxBQxammLQOLTjOzuw/fZgRe/Bp6c2NS38
331s52NB8AHvSDhwjgOBZ7Rx/+G4tzC/kfXzbXm/vxplmXFLfy9HPPF/JWd07Qi2
ON53lRz9Sc8egIF3l6+KtgxwzwE/zi1W8oBiQLQzIvB5MLlWhJXZOqjxhHWCItYT
fvpCsWj2twW2eMeKenkEZcLkrC61Pjg3QFO4YpLcpKIw6IIXgKCmKu2TqVWfHRSz
UjsTSw+Om1M/ZpJIjM6/GLgcjOvEQTNFr0dSj7CJpGweODpoyNaO3FKlcrNY9Et3
g4+yZCxlHwC9byV5dGlwM47teTHMRp1CdrUEa7a7ezAnstgkr5UzdsRi+jgxiPqh
bDZ5AkbtC+ebIsYtpKinLAh54OX5iwlsJsKRBLa22MAAxq1s6G+Kzk307Tk2gDyX
85X7y1E81Lb3opa+W8pKLCoFsRR2mxLSZS+DkiCQKrxU8L1T/x7j7VuuUM2PHvWK
hkz0jrun5YGIW9y4xzvN7NLcAqJ91EO/WD/LMWKmzVFoUt2/8gRqQGkAJWFcZzsK
b831PZQrzNbd9Zb8HAHZA5C35Bho8vEnUMcWVK3Cy3urkFpAh4lL7L8fGr385Noe
ne9+WmvVNWsjw5qvjc1fCcdPALLKiDGvZ0CcdcwrSiE=
`protect END_PROTECTED
