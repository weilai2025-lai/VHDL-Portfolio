`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8j5KJQPgsbCH1jOzvA8jbY1y+OjkI2g5QAkvEljf7cnQ+Mu6d95WD7ZoadZd9tiu
n4a4RsiwgwnPCPzBZ+8jkpGOzTPHObdBePFnB3wlQsgOIk2ApcZUHWkq1yG/dOqG
GQr8sKU9tiAkPCA7tO+HJ0TbppDalShXztmvTP//2vvqN7k9+rtpDo89e8gdV5cu
RGNF4b6mzmg4duSle2DvRi0g7JAZyFH6NeDm942SWMKQztdo7nAxEeDGOuFJogPj
mefSbJni9ZRExpnUcCFXJ8waQ4wxbt/xf1GP4pHeB7lQ9pIqTA6d+VIUMB0slOHL
Hrcfgdm7Oc5cyeu3e0uRqVjfBrIR45lhCUzxkZ7ZLjiDL22yf3qUj4fuyYGLx4j0
9vCOw4Yio0uwcb9/pG3Saip/xI4+7cngVf8svKhwMwG0fVe9RJC7rA9dgACNf4Vu
mRloObQA4T6Ya1Q5oKTZKOwsph9BEBGlitjBeGvVXtSYJ88rrj8EOMwK+reBp+tw
HUM6Qhpn9e/HA6cGh6JnP9l/U5E3YMn3os3uGjFmi/DO6jhoPfV6hBIlMPhiHIR4
0ovTwwoQ6XIKDDxzkxk6pywRnPp4m4Q3xM70kr/Xp3yes6wAGbeuB1TXzS6MFpFR
VYcX9MOUq8PoVvG0A8tDjS3dg47RNRXQjFHB/2A6eo4RmQq/VTfR3be7AInB+6iF
bJRWQHSzFwL+wVh/UGTIWWhYR1Sz3JSJxscJLTpikPbwVMbUeLxw0Cx57hL9tCin
/MtIzzR34HU1TIVErAwsxGykON+JKlOF5iYlxJhGJIcboNWXOD2rxJMi78mtaJeH
uGYur+xi2lATpPA3ooz+88lGTmDPlZ4ALnwCI3J2NRGPpETlah/303jKQCN9iKcR
WlXkb7N/sZJwgMBcRrtObWPVQacfennDKtnX5Isu7jJO4ivQH6sMpx4WRlvyw3Rv
d5zu8/F70V/24/63ID8/x7bKplsryHAdy2ZzpZh5I4LBULQjIAywWhV/4Jrmv1lP
gHZ8ekWRilLDh3263VtXx+S0PI8nqgQ3Jei4r9k/x3ZLmySqAUbi5zRKBtP+d2ye
0YiHRTBTT3uGsWC2ZSE0lFfEqUUOukes01VoiT0ZL1BE1kbw0TWhZTVcLzIu9ObG
LXgbggKxBWOKHiJYHyWf/JbxhjtS17KfvmuN53HlpuexBH4ws22A1eV5/lIyxSOa
22VufTF3F1qt8/79Lb3C4x2E79ljs5xTGoLqynmit0nlHbqOy3tCLhTU40O1B8AI
DHqa25d1rLpFBbN4QO+eArXNgVIoPaj+YkyMbL3KHtyC4el7uPAJn463w3RIbt6L
QDmkRHnyuj9zcPGh8E0OgQCLpM9o/Px8829AXX8Dl4K+cLKIsUQAQDlVke7mmr2H
+QOu+jczuKm+R0r53X+QOUZJS117ClXSwq4frJsYcH8hfio7SZ5JE6ivqiQwndGG
klPv0b7528Q5AFaM6sXbXtXbXyK339d9+vhRsvWZTa/kRzO4pWfV7xxIwOlBG/bw
QV3QDXPr5cn5fIJuTDGIWR+3hhDmhVmgPYESjFu29FuUhPI74pocEvUPkaoXVlAi
QS5NvgLXvr5PywwrHn/wPhxq66rCITaoFKMng4jyz0tRnWfbczwL3j4Nsg/eWBdK
fUL7ORxOorTUa5Tv9JpkYTRCtsNctJaHPxYQfbbFK4GS/gsTikNT0cjnVL9G0ovO
7ofIqztW1xt+FJth+cpOQCBz+dxjGqWKjQ/6lG3AMy6NxgHja32jFS4m/WkFmOyk
guQ50XOMovoylsOeoI+nOL1n3eS4xvhbnPGgmXHQFO3kqcLmaPNQXM3lZGgxt+gt
aDHXIZZjx+wNWeGE+Jh0C6eZfPYhXjYO+dBDHOagAJbeAG6c4/9Pt2uAf5FmHAuP
LIHuMG9d4bZc5RSQPNlof3u1HUZnuxx23NEB8pk/snf2hFxxjhTFpfH9zvGem0Dk
xosvoTbtK9M6rVa7D3X9twQvRcBySEphvZKmjeDgXzUicm4d8LS54PnQQM5JMEo0
gH3yt82CsrEzZwhe7438z9zUABNWuSRkLbJWjOu7uN160QwnULr7G3NUcOpJauNm
wv3Q+gHF30w4fPlMeGuANoQzckLmkWQLviXxUaKcmLrmvX8b5Mssmuouao/+pTwM
6RUhlmNTfJZkL1I+mUwvSXHv3Vkr0a0BT/qttdvfzg/aOQ29Eubs+Z5o+ulZ3i1Y
SQwDtof0+WazKli2qNN04GX9eL9QGz9x+TeYJXEorZUpeeJMFbOoAFGmKi4L+jdO
7knWQ/xAMPjp1xVdCQdiaYcqoyFvFPnz6t+z8rNztVvfoVm4XEtkY3ySFP2lW+QT
N36ccvSqIyGPJxSIYKS83vZLPiCzwX2HZkZQe8yF+hXxlb5ZDRtQSmxwCOOP0iRM
zM4DBB38NqP+FM/nbKE6bZ1hP+Nb5bcZBgA+G1gRG4Xd7hqbsRVpfy80kdegtiP2
d1F6CDynJhTgbOVhGt/JxVSR4lVqMjFtMEj59JK03cdYCAzbvHSqQs6F+Tay1fbn
XzQtieUi1WpoaMuyjxjOqw9am9TmI4YB6FgUnONDKQCzZ+SuL4pB5qpx1UJ4m+4R
NCeIjGrvF5/1h1dkl/w2XbI3f+1HI9ZCcE3qBLRvxMs2iv3id6RLiv7gjQN7pr3A
M6uO5d3Q716ciSUhrhskM0OwZ8fXupU1PMQNyyAkZnmV/H37LmcF06eyW3NFQ/1C
K7uOR2ui9eScRPpIqhKHBY1bqVaDoT9lDL6G/Bd/6jzC+pwXrB1mDf9B/yLCsQ1n
Cnh9t5efD73zTRhQm74HN/z5C9YkYq+ubiZTgTjOTV18eZLku4tPf5xTc8w+3u9W
4olg8UfInA6aBK0KeUGHispTbN6/j4I0mRpNENRPgPr8QxL1vB7W7hj8L2UYsUpY
1dYf7EVm3RPag0frCYUMy4kOSC264aH9ssDDC3OTDMcgIHdOU+bGbjeMtFYtqrQ3
sHtzbxglKnbUP+4fhnjWDfme1UQoIsBlX64NzzNBX9h8/EchXz66fS5/xWaD0gGt
SlzOGqq6my9I3mnflRlaJ24TV0fDYA/IIoVKcQYU3UUlyDBFKjhiGR2eJRd6u25/
3m2PKAJbWXurhX2G09eYRCvIEeADUJEE3G3lvRGRXk+JjKGpTeGtqVsva5adNcpk
V2zUDD7+ZGiFPTKhhsrgArJplZPyKes35+EgYk/UhFIUg9+E55g1xwrTpDvU7Eeh
4OlPzI79R04XNekoF2VA7mwSmBq97rLeMc8KVAZZ0oO61T3WGWMgDQLl0oh3Ory0
wsWg+rndwVDzJKDYIDfPTOLQmJHwS0FU+u5IkgjS12NvgoREIp427wD7ssNcGQQH
zNSZdeGJlcpof1U0cunc+WiWfIx0O7plhB5P09LQ7DypTAFMWgyB3ztb2IcZ3cMw
aj558UGlG+h52NYn4il2tR3e8zb24pc7Gi/IftGliwPofC7IZvpyb3J71n31rHak
msYSAiUePJ+cbdVZKeWMH0/IQmyRXE2h+hmKf3oPe8bjGnUPBNyKvCaru5r4nKFZ
nwLa7LMP060YR0GKQKppAFKBjxW7LVcHT3Hi2zjgEurNr/SpCQWmwud3lUXFXZAe
fSv4e0GiVE7OWuE2u4m9Ntd9WleqoktgoFQcd6A1A6yo0z/R6EZ9x3l2RHX8TTHF
aO17pyvgZhDf26M7WoSZ/SvaK7rAHGpF+x7heNrT/yS3HadlMREXNLqUh0qDAYcr
nDV/lODCyuvLr6yDGEPvFQj4XcyUck27YbfXD5PcDi/+SopxZvmktfO90OZNqAiB
BKrcMlN2a5Wsn5GFyq6IXnsB/NFDMeJ5Kdp4qBagtWqzXFjrXGpmQf7AcfdjcFs3
1UYObe6H1W3gtwdKMqHrez2hOH8ekAb4n6XLO7Icy+Nifb8oh28V4TzSH/2+mB63
TuTju22wpzjkjPqVdJE0OWPn+mMaAAa4WwKdUW0dIWTq242CQ4JMQ7ylrS/flmDg
15oQA3IolT1qXprwN9GBuCOFiBiHax/7ITQHnU6fsTiwBE0NJybuzMJezX6tN69c
mVSIArIV9FYsJW/b95+Bl53ZZl2ZKA62pCH78Bp8kWblPN6WKwbwxa2y9eZXPv+M
pmQCO9QrUzXzz+kySqcCwkjEMTf0h2FBAdWmt5oKKReJQw+XZ8GcIPyidnVUYNrJ
dVWy9eL6OLrET+JU3tNhRCgt7Z8OWgIJBknxp42GgEUNCF8m/v/GeXHMHdmEnkG9
da2SvJri8HK53JoSgKm74fQy4rrdzZdHNjBGHO9z0UUK2JTLbdqT0vEwa/WVCCSH
L4r8DYKdHoY2dXYXjCE6ZONStAQKXrLW41IF8q88mqd4COEq/QsMmCRocB3LGKQn
F0PjyXYyOEEBIQMuiPGJUGjG5S7WaKDdh9//iODIB8Uqs8NUcBOo5/e83FKRDDkH
yjCJf0w4oKaAJ94eCqutcYvuxyR3anJyGIFtgkstk19GA5nIwConA4xq8p4h+mDg
8OqVuNeDcqFa9sG7VhrEqXc+vsHmNNAp4WP4CC4AhU2twBDhEZLS8cDLbkSLFKfE
tphXcmKzuLiq0uZE+IKUdh4SJed9PN8xHab9cu0MjyaqsiwQ0xcxuTr8QhtMZMju
u2ZHLS2dpApcuGWCXN3yZGOSr/HUyQdge8Zhizsvb+R++N7fJfr9VPZueWECJDNm
s3NOBblFn3Zcufwjcko8bxP/iHvAEiFkdybZ6Qh3eWZzPw8HKYEYLakntB+aF29p
yOTkoQj5QnJL4MuEpSMak9cUeaVP4IghQM+2ahQ3OwqGVTcgrWPQZq7KoYwIJvAk
m9WIyA4Q+Z06a8Hoo3qoUWCtAFqggKdhjGeChhgFtljr93CsScBqdsSnNVhgMBrY
WqGoFyF+LmTy6UKMzXuCNcLRfoOxoAkzu+zRoveSR1bJPRQhnmMjwBUK/nVMj1Fd
okp9KCuB+PiH/gEaRJMFYzeVQWZ/GpXGfXtUNcruQbtt5gO+VGHv/9qXaQc2fUbs
mEj14JVTYFcJfxN/DT/excFYhVEOtNjBRC+z5eepzFDRf1ur3r2K3hS7tEBsIDUR
wXPzfBy2Bah36jbYnciO4sAfhuRxmo45vCqRpCQ+pEbfawU+5pyODTOTAu7Omt/G
mn4oS2iGIM8fVxVWslLF8A9E7l38zSe5eN0yHHkByGswtDbZXcN16NHzEtLRe08M
dp2NJkcPTV7GlQdV+JOL/fVKHGANrCj3a8517Kt1lklHJ/DbWh1NSXlCYKCPb1Hp
ewpPirGeYiOTCBUzXUD/K+L4Jy6uD+G+ybWhIy43Tjavy/pQYHnVNORrh/PhChvp
nSG/VC5gQbPddoU2UzRvIz7Fx2pt5/5+dplecD4tRZJwtfWZAt8mrh3+4E1ZCgK7
8hcSzoqLbRQDe9HVKEv4fHr/IPj+Mdz7iO0UQR40vzZpwV79QDWz48YFNKVTrQDW
botzVRIPXh3YOUj4MhG6Nius04R1iKoxFbd6/UASR+bvVQfXo62rBnv7WXRZoY2s
JUB/XILTqK+/M1qw508uj3okYR6vkBlZBOGd04dIYGdueArjZ/885csXhXB/Xk2u
xos6TQtnl183qMmqX5uT0B8ZavNTCTEdvgZprBBlLiXpx/ZRZ/CgHW0EIns1Jybf
wd4HL9cGh3ysEOM5YswKDqGLinNjsEY6ecIb6hTxIuiPDh2nK3e6Sgk2AhQmJFHo
qHaCB9gZVs9GRPBfIr/2hTlKzccMks01jQucDfKO53VLcFnBfDXMN7W5J+vDIW89
ztsoNJUbKl8KdNzBU+uSdXx71EKH2S1BWjiLgLrJzzTH18Pjr4m889ro72yzik7s
ZmH4LhQ5zRMqHQzIPnGKgm9MT4Xao+P+tCW1BGuN9rnkh1nkz0riI8SIb9a6ubB0
7RAFARMcfQl7F8iYaZ5GmvpzjkfRzOdPVoteA8GtLuAHdUOH/Q9La9c3W+21tPem
E4ZwQYcDpFx/6qBHZEYgY9za7pkYUW6zDN/s/JTQZ9HhqZCnoDoVyNq289bumvxg
sG8QYV15jWnNgWyJHmN561pmoVKAu58KVVQ6XNOpPvflOiLqQMKgL2SpfqlpIuDj
/wnSTbehwllh6nKnv2NC7zNQzrAzUxOG7UKlAjStmwwLPhGHUttLK1O0Aijq7+QA
NgeIc3JauiLNDPnAlBa7o9ZxzAvXSmbnA4LFTO4M/DVBiMbXBPyufQy2KsgSp3/e
dFpfUslvb+m63XPn7Kz58LUJwpvet7nywlHEWkhFcrGnbL0Vu7w8ylDi7GuaditF
bsz0MpFIxsQjj4p3xd6S0GCPYfKoSEWQCs/SpMO5Tp6DhJ3Ct4Z1DgiWAJPItwQo
islZCdtsBKnz3M5bPdMR15zF6dfFV5EH/Sl5U3ePwUWT2fK/d/KRv2A67agzqFqJ
K+R5aP0lvEaCSybOj8zg1D9dM8iMXqDZrIt7LHC18hQfiMgB3cecugfV/AeK0r9e
gE2iEMznPQ59K9yQJGdZuHHTE2CCKBW8oRT14Gb46OMRHcPL1InNWyPHICNgoR6l
exUN76pMw2YXcUF0HAmx4/FbxrBpu/R4ST9JQzN8ltQ5xkDq0eX2jZGawmNQTskF
xtcR73DB80GV4BqJEV2tEWLtb/OR6F6aS8kBCzgeavrIDnhrageMGmo4ufK/0Cf2
VfE7tbLUhMzBLL4X7yKsEUf7qfrGVwAfv6VL0FlDFfxrQZt1r25lif8liSF7ERVi
wAV2J8Rsz/OiH78itRm1UvTzX/QaKtJpFQwLmxgKxkwm74SNXtmFoeU9tBakoCC4
c9i1WC7QUdrS3horBcbN1Nfe6Q1ST5qJiLSx7URfHeVoTlNN30pPnmr3FqqUux/A
8bIFy7oiy5R/mtvBQgQa1lhEJAn5HFhI9JUAgb8Epb6AEPlK99fXB5Sply9jYPZ7
8Vg5uBSrjKIoWNVCCmezaOAg2yhaClq0MFAdruQNhp+M7kXfrOoliSpzh9MjgNvS
rheo5toe5KSIwyiGNYIjW+wdyWmZCP/9p0898SFgPG/Ouhr0kdFaGSW/0xw/SJ0c
++FnB0HegLP6fT4Bu5AA8hXVmFUGHMGx2w5bkXVLUvhvqFhfeCUaRgEOD6/B5cFO
SpMRrKdVV+aSru5xfJqpJ5VfhCDhsMIlw/RBzG3kb0P0keJbXG5660CJaQh0M2cN
mp9YaQCPwd3EzONbtJqq5tNd8PfVV6mNfYfFg3bk6NJRqr78YzbD6QtVF09UMIAi
H3hZnj41xOQWhi9tIMkhteNeQNdyBc9et+onPbnhVg8UCHjclkWLhDhYWWOsRkys
tqZgereruYzZB1Z7R7Z4GXhnbn3/YGhghl0eBiV9SpIcWIP5iuJrlQod5sV8hROt
FKiNziihAc5/lR5/6lRrCxQlQWIRbtIEUxahGuiN5JKWXkNy4JVWxC6Tg6Aa/wWY
FREtSoAIHioueO6uhVULD5lV20JBOLKI6Iqq9FwbZZI6bDhrSdkaK5I84UWLIzOv
teTe+orTAmlJ/Xjj4ffBrHAjXCvaABvRTUeY1j39TuRmdJZ1+PaCPdwtC/dDNMZs
NUbzMPYf0VhP5I2IdsVNbsiYwYVdIporBK6za2E4ifxuCErpWhGStkBYdcApDn2V
7K4tuGdG7AHwIgvOOZ9o37vTZk3lPcguSx6891l3arjBdTkUXcjsU7mM6r8rfSrB
I9v7MRZAV2UZTLqmrP2sdLL/IJjTnSer5rze3PzdFkooxynDkl6gI6l2Mw/RCjtS
4m0LMisUsZr10nfbhFJzRGUjFRUbJvRqDNSy5Sx4xLNoATvi909UuoDqCDpIfWD0
Clbk52OP9hHAt8BIQDxTghkmE2OE11DqmdluVHt7DnOFvQwkHm6+oOMfdpChmvZx
M6a/+iq4rja5j6dto8vLaZCMoDlN/4LpZf97k2Z6i7podTlm+cwJFhtLRioTbZIA
GPdIAsQ5iF8CPLD6LgUIaTxM0jJNS2no5weprI6ev9dOi8J5L1Nkojd8ngewfiGy
UAH6CJ4m+QZRFahcBI0WEwoirAI09FT8Cf3KqWjvJ9kLsJwh7aZXNqbU11HDn2Mb
TBlOn/f7Rz0a2jq28CZSA4J+YaZ4Mw8Nwy6qd0R7BXiM6O3KDs4Z1K550dFXyj0F
JPRqi6GCBHDI2hyyzXPer1jcVduT9jtX8m6ACCpE15CCWT0ZAj6zoXW9BJYhlFvR
x9S26W+3mjQAXq5K+AdfzfxIq6FIVij6ViZovu2VrQXYk+d0fut4t/W4zS+ibudZ
iSgwJu5Gw08abtxK4D/6t2eHRfXTD5nG3d2DVfpJKdFs1Ux1GSfFsRMTsrxQ/lRY
VhcSuX0cjoDLDDQCoIMa0EamT9tnYw73XlPPaW+IHNnMk0m+d+gLEbF8JdGAe8we
J/ZkLn7D3v4NfoJcoLBB33BWQPJL1PKLQMp96H9xk2xsZQw5VJNqKloZIsXnNus5
TLqoNKfNI8g8Ce+dgw4MjiH43Zl6FjfkhCIDkmYMYg1GrBlyaqTSp46+hC5BmhQS
LbLrGOsI4x/hlEWw1js2aQ==
`protect END_PROTECTED
