`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaidUuyPNU8JrZJmrrnD9wP594qCW1F6U949dwfj0S0VkK44iqjtgDeG4t0dApMl
Op3DFX0jqT4BBLI+QYqj4haqAnWsip3D/lbKsb82C4GOj01eMIU13D2862k8Sisj
+2fYGUn+rFHh52Q53Ji73ZFZ8tS82AjV2ucRyJ8lybocmKpxr9RzNSakxVxfrItP
oFsSNZMq5jUWTPXfGKsNIoxkyOvoBysp7nO0cTTFdj7DTfz9OuvFGx6jG7OeMW6s
n513BNwEvafQJZNczdqZdmDv4PSCoryI3UHHXWUHzZy3a8q9GzeBspRosL1v1QSV
flz9xvblKwIWmrVi9DBwlv2G699aDyvbWGqze9oCUMBXMsILp1hUa7OHxz2Nn6Fl
9I407avuroazuUlqSs97Bvcf6JX2KJFJZ2EdvmsGlpDTMVgvQEPG4ef7FKh7rPnn
i70IKLI3v4856TcGu7li9NH15djOWwKuCwHdhif1TVZ4LJKppljFh34A2+qbNLOh
WGROx0A9Eq5BjHJcN/jvWWXKKaf15i3n3KxdJ08cfGVO5Fm3OitMrIdWRfDd3Wzw
jo4umP9N+OPZdMzP9KYSZSHlNV8XaEx1ojHyESZsI9Q7UPuAFRmO8dpK1xUPp0he
49T5ug3YWGg8m4oDYmIwD5RCfBxHRMX38bs4MGfPlmZSjZsHJRFOEXd0MYemxC/a
NrV9vu65u3ycK35YoMGDOVI8iwOf4i/Wgq4uNPod1bOCKQQ6jTO3E22NWUuEIuTg
7uzfwfFawgwAPSHFdwFZXbe70yIvY6Ivkwvvjw0nZMgqqDuw6Mv0qAayfQcmFASu
mozylPJXCo0IaTk47lxGCQ==
`protect END_PROTECTED
