`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mk2aNEkjLp8y9zNHyYH7qRW7+gq7pQDKi7HUIN2XZzv4H3lB0lBn+11Gi8SF+egS
sG/s0HG5oEMHtxCqoEf5OwPyFFOGC7T3UmILl5N4tCWtufmjx9l0C3lRLfs5NM/0
mld0OUaRaYpuFaQwWzkh9uhiPvGoQGG9hPMMhxvZrDv/Tf3CQgcu7TWXkAaIho+2
5O8pnl8XfUXGYYacweFVIMcWp9h+6T+zH6Nysk4QVZtsYrE2nENCS5CBFQECZTp0
ZvCWSid17ocIB9ew6I/Hymt8/D6yOIv5zERWcxFOGbJmLMO4T1fYNxKT2gh+EMKs
KapUSo14zd0dPUY9jrkU9bCoWahczIMEhwv7fix1LJAEy2A/QVMc4iqP+jBZrtLg
St5FoxqhGWcxE+R0Tvxn0bghvC56MLNmC5RYiiwdlAgoPADoR8bbhbfdF5ndKkFY
LfyBTHI5/JB9H8bf9mk5+MqPmOvYlNtdSIHlEUJSyKLc+XOie9EsHiLbKfKWix5P
X2UAkTg7BTiRe5Q4tiihE0lzdF8N5GBvYZU9zmSjqlgqsJlQiFULblxFf89bmOVM
MRH+JlxS3tAL3yYUmkWoZcnD24et9YL0ZqFUaLNdGP6GUzqtTd0xWSkUDd+yFm0y
Om3N7R6tOElX+QjFo/oezJGK975HSPgYuaB6qaWu7k+SnIQhkBHAYZaPuPqou4Bk
5rhA5Z6bxR6avYYQjgRBFuF4T2PPO61kx2wUT/axeQjioBNT5Xqsny9qfVKBsO7w
R4KU3Zc4LngY59J1J2XeJrXgC4EuyJ6jD4aq3DuQrITfTfP8bm47+QH71uDkNZbN
nuscP/uvxEbF3xl1hgA5k6jKrVZ7bmLPaV6Zp7m9XgFNq6ITBZlrFY/+YcjaQB2H
yfTiq+O5dytV8DRdJ3TPh3NubwVjOl6V6UUHTrGeFEP5LdUu2DcwrEY84ghcBNkQ
yf7I7NMTE7v3Xf4flRY5ofHCd0htZINAVJ0XF0CMG4BJX0lwMLrfpG8spfWOiww/
jsOR6t6SXR9dTcT6L58PQQ5eV83VOFR64i0bf4KkGhP3b6tqdHSjQ4Dm7DPt6bQk
qVdsGcwwASofoeWp9J2OLzzfTDIsprLzJc6TPmMvOfcZqTtZZkT2BKtmAt7zMDxM
Cuzin8fKFoWNpbwoHtMH/sDSje7Dp3av7HsUe44ZCjohBkzPZBDSoRgLhgIjuXDs
`protect END_PROTECTED
