`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjmpoboyFrXy5xJ4740/F/XDWkzCPeaREQEhFCb0v+vge8NuLehudhkJKAq3XddP
Hn82gkA4a4MvLvGMU2/yTdkZ4vLCsMkcHnmfB5k4PLUzxSsApHg3d/bC/nQfeJmx
JDPcBrg9d6xtG1vnlCy/SmvIBgmgtPsk6EZIsm+wJF8+0Y+aDH9s+pvWgsmP1grC
ZmMmLuI7O8B5uwbYWS+XgOYNJPnfSwpDtwbxQV9YXi9+H98X8+0+j5XYb4h+H/gC
cFh3LWts3V+H2BaD+dyxbZEWVWta9MT1tfcIgTz4ebZOYht18apoGjArxO4iFLk6
y00zABshqXJRXJOLpi9If9Lt33MnCErtDrffZ5YREnetjF2b/aMs4mF1xVZRL3d2
aK9KP2EysAo7bRH0fTDvKibNdgZILvHWZJSizO30cwwtuWOfOtqHzdvzESrosQKz
FuBEHO7wvL16h2H1qf7rrDKX+wkNQIxI+2dssOQQsOL4NoLffnFKIFc4+SN4rI9z
KdTwQxr2MkemYRsAbqCdlqXwOw2ZD4KzG0yDLGQVscxYWMrm/1bycUHtPrmog1FH
pT/IrE1kZgzK2YoNWSYpnvCqyX3eGmuR9JyF6j9PBxRMYn696JRwH6rXIUy4cKpI
heqh2PqT233D682cTR1Zy0zt0x6Nop7pQsRIlzg+KssGn4hXNQIf2mPS/cjsZ09U
oSqIfluiFpkv8rfSPvlixVPXIo4BudmXicRZsiJa212YBriWFNZ06ZIyMOgDDeG8
XIvd9mXEH4gG0HdiWkJGEw==
`protect END_PROTECTED
