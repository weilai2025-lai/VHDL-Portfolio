`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTeMgzdjLb7B2znLKC3HGk74PqFLbKDO+kjGB3VoVIsVrm6oSC2VGMHn0BW47EO3
WX99Asam3OaMXF9ofEd7dksUMMdKEIpkzy4WJdsJ8855H9L6zMhhHqqO8INKyxij
Frmy2f9lmSZS95xrXDWbYK8wqOoPiWZLcKk59HUSaR+Iae8SFuyEPE4BxDM+XuJp
z/j9UZAJyGZhKSbAimgOrQI3i7q5egjyo2xp48wwmorpVF/Noi0JrJe8UwN6bc1C
aqY6xw3tmaXHFLSeMxmEgplRagWKcAFeG7KG/0e72Volmgm7iYHeACxyyP9Bl73V
qYZnVgutVTt+x+AZmVSPJWsKZUt3fkhSxJRdTdwXWKiiEos6+o2mhfYsDAjEpQhn
HNpzBCeptn90YUryxfRiKRo11gNoUv4g8/52R5oviQ7IqnSEAgGFx6hGIP8afkDz
VS8hWuzJcA1YhAheVHSTR+Xu8pwmb8RSUsv4VN80D3JWKuwBJe/aKuug1eo2bhTM
laGpDu08PQNlmL+wGbHg/i++i/LbwULLROLsIZALIJe7kgMjhLGRP7CMiXUuIIsH
2HHsMXap1U+fbfEWY+mU3vM3sFL/1meKwILy+6AHfTuQdLKGTmV0pBSZBAbeBuVf
AELj1rjlEnAi9xtW3dDZNYAfddtKbruPXHE5rAxa58qzh4L5LOoGGXmW0D0HV7VW
NTg3nLLmp6E/YTeG70rMFc+Dy4YZ49MNQTB+uKSRh0qEeU8XsJ43CYfRDD3H7a6e
Z737Wg9Sy4i+TeLiiM1Q+K85Yx8U1jFN0xAgsgwT364NYNpZAV2J5yeZkZDOkaxD
4Cmpw0XT2z+yMRI/n6brcgig28XQb75LonuZuHP2eWsQjAY83s+FcSGUX7nCBciH
hJVSuy4/5nk8xIaHXJF2WN3dbjnP0DgqrtqGhFS/xng7Ztp1EJZQWtnoeCjpUnDi
4PMgFYItCDYpq7oJ1NGHzw/WVHHkepNfetWMX0blTdSRPT4XK0+tgxQf+eDnUMuj
1WgQdHEfmbhGgghPnnIM8LK6CT39lnJwgZ6S0luCrKCQRX/I3R519oNMqDdfVmJW
97et/dm55QeDfVD0YWriIAxONWc49mchZ6goZPS4EeOQp4xnApsDnPA0z4f29WGO
fBsBqIJUCVB2XBu/UXfCAndNz34qEIvt8w520fepwdltOSaPi/T0wcq83GavkSzA
sWGJufTkeVw4Jql/jiKfwfPp7xMQSgYrd0gcULfs+HTphLi+/r6Xqa7nPc1z4u/t
0OJEIC7BCv02QfcVR96KOKbwaW38sQ7HBXNqnR4PYGMJmBbqgD+9uUxOZ9mRKLdl
8bnAFEC/jJk7leY58+AIjum726n9EpwGoQ/DWNCjcw/4hu0BWJd8vqt4tgUinz1h
siSbizZLxh/kRggB4kvWOc68YUee2sePB6ypvF6R0YZM7FOWG049DF9KhfGOVayR
TT7iLavmc4xanFIcC8UNug==
`protect END_PROTECTED
