`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/RtioTI45tcmQuSSG3JTIU6G+GOTQLi3wN8x7XrtczHQswIHoJjwMhTZ/6Br4Ge
WqjcgmyCzrOwqV0zbRxDYB3WrSlj/1EtQ5CAuoDyQknWkQhEcTBj4iT0I0DqPxgq
v3P5Mc/idW4d9ClBjPuO1lSA6/UOivRE0gs8okP9y+96yEOAsCDJm2+2BV1A/J15
BdwtLjgwNriTaPXiE4ldvpb5ek4Y+eFbuwcehVLHRYne2X61dhPnhaKpW8ziM/e8
K/XR8fnOvJznIjhW78+fxj9QQ8hDi1D7NkmPkCSPK2cceXBJASWzNvKC0di74+sE
StFyD7wQRlqZeNAC+oGa1c19FTo8rp6YD/6IN81TZ/g2vSExUKo/APtEcgjtTQF8
aqZe9MGexs6kmvoQuSRRQJm2WJ8afNlQ4nf7ucc4qlvjwON++peTVMSx69RC4qQR
AFAiKeZ2Y2aw2CosY8kgfEfewzQDTiqsw6gD/bukesLsIMrH6O925RdlJcayVa4R
NgFu8nF4Hnxx6fxjoMoLZqespBlZ/8b9CfPwP+4e4uTXJ43dAB48d+SUY7exIb8S
kjPforFQU2MZorJpBRIGxOHJjbQPvvm1qutIylJ1rVyKgcE16ZnP7FCBee+dVrY8
08MeUfbPM1uWArqkyBlE1CaqZ6uocx+QDb7Qh9lxkXoEZNDdvcITElNhPOHjhbTJ
eZN4auQ2MuJL2Pwnn+YZJEQpL4ZTFfZEAMgLnrOC8SE4wTXsqttozfFatbrrAq5B
vET0+CWAsNqBp4c0xIh4jNUNfnGn6ae8U5tCEZUI3oa78LARsKiXv7rWS82fP+It
B4oZ9LXMWHjdn2HokwfjTZKTAtX2mLjNAVlmqvLUuZaVgK1GsA/WrZjMZvlFJj9T
`protect END_PROTECTED
