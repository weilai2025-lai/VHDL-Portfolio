`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
plqLChhgGYTXPstu9fa3kH9Kvfbrim3dsvIpfndBd3wzOfTp8zRgd8LqCbaYfVno
zyD3bu3vS2+czriSDCJi+kThSLeo08+EYORDFsPoXGvvxSfRTuy21d2T97chaGLc
2KeHvRpGaZksQxQ2t5X2rKcbgWt/hbsyyphF5Jby8dvG/ZwehNHTtfcwKCe3dVYR
gJVIO0Ur2ucVbKCucBRBbrIMHSa+4hC0rRncE1v0mMnvulBI5ztzU00kV533PGlA
xyayqgpwV32C5flQOpQ2oZHvtSwGH21mu8PvSLpTtgrzQGZ/b2MIVtOMAuT2Q8Tr
PyfshMON1J+cat7jhRFult2gSlHlXB0I65wL8rJl8Htv0obrOE+wXoX56bnYDlt4
0kVGnLkEtEoNM2LXfREa5s/bQDKg439tYsIG8oiOkRNYc09n73cq2WslGJw+zhvx
uV70n49z8vr5U4HFPnBHm8tSwWrQuR/HKyQLfU+p8kNKDTVCqySSbaRfJl3+4UuB
+douVqfzlUPSIBqNNf6lmVkbqdhgxs+cT93S0276CXfU7zXWataoS4dd7aFfI8lZ
swfDLudq2GkM9i6/Ty0YMaNH4I3JblDnYCPcnfWaKrev22VEaX2jwdZZuakVdlvP
eYpn2fby+EgjT+mpaxSaj6Y/dkfmrrQ4mz79vsXZBIN9DSHJtCqIEB3/rHrsbKcB
Uop3ThhkWyhc8j01WQEg+bwYnEkVqBt7Y9HV+zmjJMA93C9ghweV/UCv3idaFjOx
cTz6MSjIlzmjI0xRat5sQwcNSlafHuDnw7sjPXCuGxXCA2Yq8AiWfprb3BQchJAC
oSL61/slfO5qKHLd3hb1tCU/opTY95XPmRDSWCrBbJyPmg3GGq8PilC0PcQG1kiC
lBZJQQT74DFjB9zRCD4WZQ9jjd8/gtvQXaxkqRDvWuSZ9tEvv4JFiwaFwoqplwog
gJxJi9maJL6lagLWoaka78C/GzYlo/vGRMiFl4hSCvvJjQCJrPNTZEQZEVx74fHZ
15/DPlr3sx7sw3gbecPic3pDKtG+9J95SpkDpdmZ4eEUC+knStj1m1VPKKR0m4L8
t0tEoxQ7JU9nsYu//lNUb03Ik9jb+ZcwrymlhBTaRyLKdxuflxIc6WmY+jETwf1O
ibQEK8MhOJmUKK81NuQqh06Ezv7ctPp5i2OI0xD9bbWVACjnd76j3D3Ju/t5+U8I
wNxLA+eHTkoTgIK7AWX48D2qEwTqHC6+zW6VHfxfnuo0kcNWKKCaPubKVGMVFYOW
d2PpaeWaaOmp02nWKsms1wJos8T0FaiDwBjsDDMiSrVhfa9EE1p+BukH0o69/xK+
/eHnXeT0pKXM+ikARnxhSd/kByUTwwBVxatrtWjGTa3f9hDuXDFUCo74dxKPbHPp
ecMnK5iPNBzmo+mExiIKn79OFAa2UrbyFboWoEhXRO16l2USrkHnujUDeMex5zqh
sEkqEcjc8f0d/LOe6krL8g3goQU3ijpUq1g40SmUPjwntzu7wZEOQc/keKeNmyuo
z6INf+OXXvZngZpzOr7qyMjTgZzkjMk7ycUS7xcKb9F/9c5qH9tIPKMXL22hiQV6
kBbqGt77A2ICy8zYqdmg6QptxVT/OAB00dI1qr/48q9Ypo+Yv755NfpRCPbzmobp
dvwMyPu7JSIbUOg1ojtlVc342HUx+1CSxb8QhwG703xNfXt5gD41SLTAUoCN0ti4
uhvy9Zjds3qGipKcLHn9X1fzDwaytFXdNqmTQQJYHSVc2lDgmBEYt9f0YCtft4LE
8oHg8cyfL58FzAQhz0dZpYhpCMpbXd+KrKXhyPB5Pc9MBjnQ8ArkvzCwDkgBftpX
iBBuP6305EXJsRfAeSZUc8SJ7Lew+/JsXjTc5KvMggXoZsmPYhWivNZKlNbNq3Id
Ku6SDciatYosOA+tYcWX1EebmkMxI/B/Um9ILrkR6IjXnV1yF2RAApWfB2z4BUXm
J6sNkFVqAJQLxPtR23TbBYLo4HhmOYBGosKnXY6NhUKfLev2U5pU7EfrpabYgWsm
8RbqgEJEqpUoI6rdBor7gTp8ioYguVBK8koF5x68XDgX5VF69fFJRAzv9/X8/Our
wi3mfFCOYIpdVXrVGTbJs1LYTB3X4RkV/n5Jw1K/4QF3ND35JrVGZLW3eHEmEF28
StQnPV1OGty1LsdtPwE/uG695s57Rr/xUOo5dPyAe+qeyLm07UjJ5yJj+i8Q342K
2HlcLae20vmXt3IRVBAm6mcDfc5X529VMU3WComU+EoSomzVCbo27AyvuPWwyXUB
q/hIzPRLleWVtnktxTzTrEStbUV0CTUj40Tpnd3ZZbf8nsIriZqJ+vj9JrK/NvgI
DS36nifZiO38tFPTyeEm9xHPoUabybtsj8muQ/6rOIHPueQRC2VkVL2X4MSX6ZLM
SSgtkipKsizgY+SZrJEoQFv3DO4amY9RZw7OgbT//IcLvYJCpEJSgBnxhVPxx1Cr
SzQPj450Risse5FLMUclBTGMl8YkpkynkhFxHSAwPMk3YKnIk+eg0twX3YW3dQkQ
OBCy11KR8m8HXob8JAUtknYjyQfJ8CEf2qiYaK7xqZ9X2NhEnnSHzCDXQfTWwLgS
+XxwJ0c2b+ItOyq1zsgxM4INo7DVPsH5G76nlQB+07NT+rXQgjjm3Bb8cu5A6xzt
zBurHl1jzeEgv1X4ECv6ir9H12yB/e6XJWXwxMKeBpjhe1ce1RFdoMCD7DX8XpGe
0HBplUjrzl8rQw2KZT86rbW0LWtJsksQaSUIudcK/j4qATRvd30CMj3svjkcAYgc
9FH91+2NpeYG0Mqs9nhm1Ue53sQVGQvTCiISuC2YJyZ+v86hSgi46Z07iljJwTZl
8R4DC3TiKRQ6VAKHm6BKw0Rk1xNxWgz6eA6kV8NxFNO39s7NZ8lq479ppfzTDK2R
xGqDVaOTu4zVbJPUt7oCCjP7MyI3pzCgOL4IZ6uZqk1mMpDYSZY4uy1HXYOVfMct
lEZhroeGC6MHUbNmJYtvFj3pIb8CX3GpKhwLq4Sjum2F6qsHhy0hRMtu3jrzTfaX
avBCPATCyp2fXJNz0tj3uZamRbUkOaQIE5nZer3ay4xQja6kr/01toRReg29qGT0
nkHJfOilWHx7IM0+jBSofkDwxLxuGkRUkWJTIUmuUJx3F9WOoNzL7TooMTQKaNcE
dQcV5FpjGbxIsuEhEx1z2gKPrsFUyUX2BpvXaYtwwAwyN7d+QhxhC266ulmx4s3F
fk8JMzmXtO0tsjwATDRbWyxiWnbvV6zWAS87aFc9khpVbtkfu1hizcIrEAh9IuSw
KEf6p84hoQsAXV22k6XqjbjxVwcRxQbQ7cZr5o3dHqc38b1ZYEaK7KECe1/5RoQL
UHp/OZhL55rgxr5WpHWY6lTdeGHshCCbNOZid99dlY9XFQ/HL2X5CV6TK7Lk4SWB
8XVeX9/cwGcDQrPrPpLuGXM4vVPVCo+LcvCdgwSa4K2+ctaXHyr/EQuDW0cBXy01
nFkA+kqagYpTPgkNrW6mk6CsO6nhw7zBs5g3EbF0C4xN/4mcPl7/G9HZOGCWD92n
FFO0juYFT/wXXtnn9o9PMzNGbhO0b2Z0FkqOBA9ryshwcgTbHj1Occ6C4MWGC8k8
qqK87q22RN7y8nUGsK019g76PEWvXXEd7buMU6zxPsnJTGbG1phR9/ED68ny5ZHg
wQH54XUW2k7JZRIXBn1nMJO9cMMORZ6zXgsZuErqv9mDGOOCrpbduVUK5QoeuTgz
OXuwVhkpc+XanCHFIWLAYuHMVn+TC+UH7I4wulASbT6HCsx6VCNSnLJ9l0yaLq2h
U0Ii54a3FvyUZfFufmUj8Loy7Z/6OBVOFvqm7eOBZiSqI+oNC6aXBK2YHm9yJast
OsZpFz19eYf2xIP2XvwON5U2cU5J6kkYn9ut84KGrJ56zR3eEaSKanxMOYkd5mlZ
Bw+0jYjLAGjyvpS+YIGwt+Xz+YEvhNV8qM6LeV+vtz2Go6TVI8C+NZynLkRtZRYy
hM6b8ZWMEhn7T+qqaDtSnzAakd6ZFUW3aHpQ9Xeq+9NfTG5efAXLqa8pPFIdmvw1
h6FHiM3qnaMf0QJPgQsxRrjords1Dbkq8CPJNLPpIDscj8Ld5IRPSwNaKISgtrMW
cUNVr0McmEOko/Zntvbg4LxvdlvBQiiPA+GjS9tppAP1qm+Y/CKVEmMbxBzxbC1O
rLQeT3nk3GKXK4Hp/FoMLDZ7U305oCOW9ZEBC8jtjOe54XhS7ziQu0l+WnPSbL0G
x0K6Du/v5CS5+BwcLvu0XXHYTeoq3wie0cupkPPewVZg6Ubm403wvsXFDX7uKjih
MOtmLhYociWggyMAE8733KZ5fovRWix0eeM5ocUEIyG7qvkk9WBELPHfLXPZ8bzb
rCYQMgUW5t35oniEJqrLUnpb3n61uLbi6FttzDMXmVLZTBS/KnBsvX2iC4FamLzN
uIvYfQkem5UNIR+xk7aZLi35OjPSNmmmWoFEu0dahpUuiV4lipAR5aJkHUJxMPEK
g0utTVsa1OONjp8uq7Zx2h080k6MHVXjQVhX8fVeJ+2adnkCtVf9ko29nQE3n7vD
7XYYGNxx0qJd0izWcqvOUkvgZ+/D7hexunUzkaker7Vv50JWtYySvh4nWgQgoyiD
RGlVvhlwC1zINfFTCUTIbzi+lGZxOAVT/9nlLq3YyxWdQYVPC5ylexH06H9edhgY
rH24moLDDcQuw+q4qQrV1OhzjfcSHcnpKssrOaftv/lT+uDSez6/6tYLBxuGwfg/
AZ/4c0gNClUZN360i0FelqndXM2Zz0iTJOvAX0HceEA+R6QUEG4t+B6RXApmhftM
GDiEceR8DIVzddpParnAzRCIV1FIgR/u+K5SereNDmH/H+xrYWhOpBaWsaHzEHHv
51kqFc7WA+sVeEcl6o+s26JPXQtXuSUuNJmD6qgyoYWFluFuLgqcCA7Gk8iKX9uN
FdJOFntMt8q1v/DP53qsBs+TTHI3TxWbZhuajup5TdEP0UFg7TyCNgXYrhxd51aY
nVVtoM5ZMZ9wJfcfRvrfOL00SmDanEWDNhoc2sMmYStxxgcMWFE6/V0HkvcCLfFg
JnR1os8YlsgQktNtJtFt1BancLvDJCTBwqVgQ+X9LF0/fDu5ViWfFJASZclSxxe9
/w/uV/OJx86AGsQ8wcDLMTVQAak78fa2xXcAFkpvEEYptEbCjqWQp7d/GLhyd7LG
SN0AfQLk8YkSY9tBvSPy9JIzSCYqjOEuJYgMWvsG7UX9aCnZ647kXD39QEmMuLXc
t9Pgj7UKGLLC46AmrnfGV50UAlzChoBfkOAYuVtuz05nvFxChDY1Mn6QvL4Qx3QY
sTXxy3bQ9JLgTWKzU1n63PpYLuu0iK9DiGfWb897VTx/FeP/VT0yEoAe0B0uHCWY
B4eFrV15mZmaHbGP68FphA==
`protect END_PROTECTED
