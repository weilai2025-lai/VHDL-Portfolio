`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CuGRrRihqZ5rQfEyMb5uBnf8Qq1U242HA73nYFz54ScxPjE/ZrbNvdG6TPhLvRg+
rioXc8BKXmiulhqPPnIeY3bZirsagKGKiKvmEGrI7vMXd9+ee4T7O8qVe+puwYS1
+4V0q4IJ0eNb9TxZrWPQWXimiGCXskVeLBnLMIwtoDkQqHB/Os4RkXK2qOom5Hw2
rwlSYU3RNfFkkL0KjxTsLrbPvlKhxsHplDEehF1TYXjo/uPtI2CqagFFjYedPlPm
vdSdrJr7XYUAK8/ICyrAjnb7JJtXrADxVUk861lm6aN5dDLP8WApUrkXMFiGCPaq
kaPL2+fayaxvGr/qCzLYh5qB6pdtVGBKoK9bY46pfI7VPY88k4x+98v2KLUTHG5Y
MSx1++Mc/kqIxLQMGDRNkWWSyoVyOhWg5kk0tavycRqiiJ7adbFlmbFLIP8xHLc6
hs4X0XmIR/wr7iFsZDekeqcP/1sA0T1KvFzyf6UAAkv7Y94niCsxOtGBr+9X3+jD
m7nqxngFFa3ta6gay0a56/TbfOV62nNNihdd9Eb9F7wgEJG37gL78xzD5njScrY8
otBbBg4w/D1DGfMQ3i0R+A==
`protect END_PROTECTED
