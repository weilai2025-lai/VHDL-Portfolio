`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wnnFwxTRxVb0sWaF8ubecvVYtsTfbMsD9+6QFZjcwj8gjRxOqvlX7OYFGqUDTO22
MGWwXzDFFN2s/QRSHwTAK9x5t2PT2GxJ4xK1VEjUZ9WCYltWD7RdkZBzZKMaV9Bo
vxYsY2csUDcmBFI8ns+/liy7n3YI+aU5/QTZhvs/6K6OzIWkIvM9J4EODXoRb7kd
mjAodKPYmDtpUHZBGK5kBL5ayTYZeHrWqsu2ggq+Z0AzLKIRWipiOKX+7ltCHJB1
FoAVow/q/rUqBUTSQ1eti9oNJGKAzBf5qGRcrncn1VjqC/ovzcB5dw8fsaedGpkM
3Sc4OHwyX3Nd6hadTcLvmLEZ0IaAnooqDAh3INU/EWr8YiNQBtvhpcFXlzaaXROu
6iWXONIVQgjvb4aYGvLIX8yzymHJlNk7uPIU/0JcNo8XjmBX4nwYzWjc8wJgVDUN
zgAYNsM3pultK87P8VS1Ni44kh3p1uXUjFzQTdjUG36Ew5cQPkgTrwHmFHemtvzw
LLTRzJ0JsngTeOpOLs/WkuTR3cXZIC7q5X8Tn0WHitObKswxxXQmhNnvoAP5AsFB
d2Ta3Oh/EALzU0+eQHW+jDmbsaQuCNb4QTIsrj5Egui6AeQbqdmRxkTojH+/BmKs
PDPPq3sA1h/JHHXqVphwqdQ5w8LcBFuZzTWcfDelhwYP64sevatFcNHFeB/ohW1i
NtrriN6KouHIU42Rk5wzbbvU40N76Zd+/1bsouGcJX3InJf//JEluftHDzEJDZxq
0inr4EhxdaWwfDg7MJRzhlfyufi0hU8qwDsdu0MdtJbbVu/RkHoyCfidoCLggzAx
GmHFiJXpn9ZdfssBVxtYwMbg8PbT4ncDLg1dCVmY9LNrCKVKNQjBQwdfDTLzN8IB
HQvDAwwHxcYob3Ihk3DFTvk9dxaZrZ/mX+WQ7ukl8uvsNcz3WpwtVVZ2P1Tguv8A
LPmuWBeQRbfbLnovz5HC4dAYZjs8tA+YDtCTlfDSnvy5XubiDDQsM3H06OK1+/kx
Mn+0R4HafMZJYx4A4fNOtcxvxfiAFmf3Sp4PIxJmljvhz/ppebEsON/nn53x1IPz
IvvHnha+1BpyIm3kVv7HT7fI+SmJzzON+bNc/Kp4k6fGsuEYx8ytXdnT99Te75UP
X1FlQE5WJcME3O3Edyk7tiN0he4RA2EjTqHpxS+26mDesL/0xWrbpdYnT6KMWs8z
S4jBeFdVRN65dPBs5S1XNDO15CTNldBPE3XFaWvhrRIBSyhvLiJKSrS/GfmFJRRC
yiAcFiesQ1uyzy7P9yoyF3bN43FljOP6HnjXeNag9hOJPy1xgO/jCVoRxBSlCJbn
CzOIRJLaQMhHJiQzUijWVosMt/I6yTyJtbhjotr+SUrY0ezYFVOcSdCZFUPpYm+b
o1wnRCXAdJ1Hex6+fXoi57H3mqbbGycpN+6MTEksMIcnFRkoXCdxkAgHdZY8I3Ee
gqXq9/6z+9MPcif10DNIfL7AJr8NK7Zkl1JT+CFYOJd4TU52VVBkXMG7QWs1pGoC
VNk7Mgm+46zQdurW9U4YmPrYW2K27zyo3IfX0yKS0xgge3N8BXsOaMGKSkfma42c
axxD1UXveOEFND5mOuLwnx2JApFkR+K/OAINl5Dh5iFm1lxVcHHqcKtK0P4LJcQl
BQIYHCoKM+644es09Dl3FpScD04LImRVJuRdVuWwSCDZ0jRB4FAF4+ksTPOfYx4h
oIrvwXluU9Bwibvq/IG+tEpAT7WdELkPfHoc6v63Xnffvu+zWE1gjHA5jWiDOXsT
Ys02iGeDQgoBBhxJabozJ0KfYq8ndeYUNhnsPqwKaljGWoFFJ/pArYv75/vEBLwr
SJEyAXYQGIOOAc78Qg2C9cOmj8JvW10dCRedQ6yWSfti+kN6S71H4NiVvrEtYNtX
lDWv4QImSgjSuJzHM0PzSHctCyvuBmPauFcDPEAAColYWtMwfK1dTs6+oHgg31M+
p38roik7Ohdrc12f04kyPh9pOGSiRvyCtLEYNnn75Y00bdxZ73P3rUJw5h9sSnDr
DiCq71sKIfyjwBN7HQZA4h3lIEm9ASaVgSN72mLvSVsChsktPnrFM8XRLdAHK1Ga
MaIBBWAOyZsCwViTnBZTuDOwwYQAxbDgRz+7+lV0BXVln2fUUfbXlDEdm88OPL3j
eZ/M48BvxwP8l2uIwzjWEUedWebCscoMc0GAe1/z7UYluc8QW6LyJ2KrQth8A+1l
oYw4U68U69PIGbFigduS6KodKZQEpsf0Dcx2iv3Nf75GQbCWffltu3pwKeSFaw3C
tl/YGXZcT71eoMuIDlP2UsEHQqwXk1t+1K+VKwZAC8Ge39RTvHesnhVwv8BYEmSK
XiPZHnWnUadmKXbsdyxnvJZBRjm2SXHW4O+w98ywu6vniaPRwRgNHl0+iUMtnZ4g
ZerSEu5x/g+ryzt3CYMlK5qh0e6u6Cle+l4SIn2HvPAC69qQthGkEPQ/Sgd+Qv0F
bGt5uyVZkCbbbFIT0C+XbT0CN+zTAg1/Bz1W2dOYgBerPuaITimpnUcMI/tttxIB
H8bo2jlsNUvmvRJBXpofGvSFQPuU4Ux0dWrRr4JkaFKBTPUH/2j4nhkAiyd/aJhu
kiOcVyGBjC/Tcgz/88B1YtBvcFxa+7DHwlnkHkNyozA=
`protect END_PROTECTED
