`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QbRwvWXiX4xxAhtOu1VZ/+rSLdhkdftzhBzGjGgoVQsCj2OBrHjQvYG9NcQgSffV
fw4aVg26JdsV2SEwBsLiwzMBtO4dKT1/uq1qxfRaTv/DIXMEyoVSkvMzHLdCs6Fr
dy+E6cNI3oypJvL9FoOHfcRRR1PgCWrl5vmDiX2093tGW8m+rkSto52Rvx8a/DLi
L4bAnPsNP3QWCrNIrOxiyvu4lN5YzEnRu0dMCTOXSOt/hUrJ3w0jtENzsYYzyXct
Q68drDEzaWLdgT4xSnCTrHsSVQD9TkSYOm3bSpUANZEFOxZWRulaD0ZsxlLNVB9S
GZbcLUeFqgCphyZMW/NNs0/QPep9I7+XeAqPN8PuBdeDzbjZxEqLQ1bPRzPIgc/9
1FX3veqhtqqmaFoup0U6MjAc+ZGUaGLmrwSjVOZ5l08iU/K3gOZ4WUdmJbHDGAkH
bg6xicWKmzAR02IQ0bSEMJIjQdhhK3WigimaNjB7R1aEAWIcBqGowngGZ8MCWPYS
OguXTrUSqvz70CU44VlB3tW1H0lvi2yvRxWiQD5e25qNDwHUXp9AP9pZTZ7Qw73t
/jJJIYDvyF33W+T8YLhCed07RvqR96gKE+NjNqYTUi8xMYWsF6oi4f2WwJoava6K
eautqIxIN0KRPTryAHc7FJDxoyvD556YqJjbJXXnFEEYI9lkg/Z0ogssL6A6ROpw
tsZ1HzhbZsU9I6HLfZx2jwvYBZ5Ras6wpcwWZU/tzNijYG2uAzufOegsfeMMVAe5
yaZe0O24G1Rq/3qIbhhOQA/kuwJZYVzYpjlMJRWvURrJ+rvPbvf9UOIPny7GRHfp
Wvqmn2gu9mTA6/IT6RXmbFOS2XRM69i1NQHFvmsF2XECBjeVFwqOhGDWq0CvDZYI
nfePxc17yLATZbwjeCA/kVIZ+Vxr5ATvoNehtITRNPUEXl0E/0yHv/HdOYGgua94
xXTrJh26o8PPHCpMr8tFtDGcxcmr0dsissT4Lz0Fl2TMAQIoRzN0TMk7QiOwgABN
VEecaJVLbyR0Ap7w1Gb9paAHIvHbfNDJUg8K75l3ARiS9YbxMyAZEYjaAxTLDciq
sWAk/EL4KXGbEPQsdIChT5dCJlQ11GD+Nx5XDUYz7dHW7q7wXctgSpUT+YzyCtTe
C6FRDu9CJDdV7E878RRTnAcJxQsS70/HB4nIceKGCdAs75LRYsfxHC42kUGYsZxS
FyY4iCn2PH1bjTAranIt1VHBlwFRCWb757gqGTSvkqCjT/xc/KehhSggSKEc4lmf
J+Jn4MDWdp1jX7fQsBKmuWqDZbElXIhIDOfWadyJJtGhxcBkS26QKXj3cvKgqx/j
5VpHxaK5cuSu8l/jN1oN7yccv7tcWu79rttoL7bWfmgYIkFwDMWBuektLrCL83hg
Ek4BYHj3tUMaK9gmqVRbP+Cd9uYMJqxr2qc0XzLiRecbdIdGHnE1lfUbtrwdaCUP
elMhGtxm+U/i6fYQESP+ZiA84wBPmgEAsdLXxTOKkGHt4YQnbxgKXz5JQEZ4UMzc
01CLU+sB1npPaaAkM7xCiT1SsxO4j19xvTjQA1oh//QjoNa7wgkf7fUcV/fTe1yq
tpUJdSAgsBaF3/QAIzewjgjNVmhhOulIjOa2v4t0kJMWdLdxf7gwK2hRatZH9G7Z
6kfbjt/wlPIrFpFj9VqQPE+PgQlaWQ0eDU7qAVZzt16VoGXovISJalElHxW9oTF9
8jsXeCsc7FsuA+kASeywlPkaLriKVIIFXugQdDXhb9Whd/eorYQMBDQhaQucGRtt
DCSqh+QcJMjqR4x7CxHnDL98711cSyRYFRF3ekDepb3rP0if9fXLqXGT3S/Mnepm
9UjSvql1kGreVihk/RhtC4+/MVyZ5Ku1wa298ycMjeIgczZc2sns6gwrIRb1zq4I
AZufeCbHFZyqNSxy5FK14O13Mw2i9Nq5CycvbGviy/MWeBJDcGL0MjRByWeFO9/x
Ao18AMQ4zSM/fjZByMv2Upe8vYUE3/VMcrze1Vzz5S4V8oF+T/Kf2y8s4d4EkEKN
JcOohrflAX80f/Qa2QuogIx95Ep1jjTp3gBwjpbN1YAVeYcN3+A6QCiD9PUOUHl2
agzR6ZRD/+pD7wXENqrVFMeMaxkm3dljguj1HaozjykOUWN3ZZYjZL/8DVmaArI8
Jm7OCIvmNKDnJ9WEelRTDCH018sVwNyCOpmudJoKzSORAg4dgZVg/N1G7fDK2ys0
wxiWYNrrGTqRgsp24hPtYpsnBIsxV6MTx+ZT5Epq+E+ZgpUqKJT271abnlpzU1Rj
9kLzGjIaMxGKRBzNcKtb0GTSPDlxnWQdZ19YSAc7XeF50VeClvQ10DPkmI/LvVww
9PqHRRS+ti/gJc6+CHgzk4VYvcJA76DmOJ8cGG/SqVsggxTq5UPfd09ytOQhK89A
rb4tgYNc5L2HHFhWY/IXhjG5jCllqRJ79f+lZx1lnHWrVl/FS3I6YuAGPPt9LGW2
ozTzqoCoa73rNxUGDdO4mosiK5EUAl2WDS9dHpUWEiudIjKGYHhaoOYgkiHt/DE8
oRrqAOSQMtxa63/yhdQFbgl4/MfXURX8URn6ISea3qzs9eVHD5yGhFYKLN9o6Y96
gRsTmiw+E+TlSpyGGGra/XbfEqKjZqEHgX+V4C5O04Xcm/j4to7jes64F8tdel7D
mDLFGkMO5aEr5B/RN1SSChsTrUqmlJv/ltOy3+Bb132017akmPJ82rUutffKtm7d
dGFf8v1V0PSfw8ipnCSaTJdCuG9roL2OULc6NVjDiAmzJ4uPQ9R0niV/kRMZt926
zr1GtRXXgMARHK3BTf3goYfCY1zUM7Xx2iT7xbSEIVYzakfnhfVgD5Suk8Q4AVPm
aDJsW4x6QAESlbh4K6xwSMZrBWyzZVoRuGa0ellB1Z7DRSWpihaPMsgiLCMPHazp
AgP/D3hrb+qC9QJIf7b8hg==
`protect END_PROTECTED
