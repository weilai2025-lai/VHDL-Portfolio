`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldVC4DPI1NttsmbI4zoUUM4qaT+8B8EgWJkl+zW1+WISvCithJtJtYqUO+k2AjNy
R+8rhpu0KSm5ddDPPzfN1ZLwNOn9FFhX3svhKvdOjNMmDoo6kjU5cK0g2U1MMCyw
bPM2lrSFkpxCAHJgp9VzU65IRCN68w9corQuxYnoOc7gd1g120mRf1wYDQjKTK8f
xkh89nWx1SHIV1EwZ+fk/UWKBMw4CqLnkgdnI2yGhhY/fLnjdbJjeXfKpIblPZXY
bqOR1aV4ZV7CiMGCm+nvwUAmBkudgHn0kKuTevJnXXvOfln04EOVer8HK36xNl9w
o5DD3iBS2KTcr/dt5J9zBAtPje5zVpyLGTxlloGJNdLgyuqerewskt3Is2hHZGMq
I2NMdT/1w2XS1SdNjYFB7OnPIA3wLBN6pFQGwacB85Wzaj1Zo69O7JL/F9K4OZF8
6DcPun1YdL1QTHNJLEMmqt9Pe4mr9HG5jpibvwyeefFaOUIpXo5rA1Aqaxoo4WMg
kCk8V02lOP6JJy7oFc2wXAZ5a13cm7vKyBwstmhv0sMaA3pfXtp6su1cBkcK1rNA
4NDBc+mZMQ1kQUOR5bRKVL9ag5kLUKauWsiycXtg3UFxYgUUzNjio8dPgWO8Td/3
dSZ6ejy4XCwiiLcdHZ8/XGIPUHerVP7OJpwRZKmp0pOMNSsmNrGeNi+h1sol9BXi
nNg4Xff5AsL5qXzJA2rMqGZUKi5RC//jJkFXNOui1kA3hhxA1Y4Os/XQKvFEzrl4
NiOLly83RD/2l4cosPdVch1jZDpy6YvcSDRXMoQYEGwXL++hGm72yeu2azMmIFue
/kCJjnUKplcTM7AsnjZL2eR+XSeIIYNuoeYmIiuuXSL0OiLmlAFbOxVYuWE5rtfn
hnFwW+joUp2gtFiAN+QNWD8jN0oPS9cg7K6euIVeyBw1DHVW3uWk7ZqS8N0/INOM
8ZnHWaizRr3WPdikU8a2JyGNeief6Yrntg2lCwEJEyPOB2aKwcZo4s+feXrLkvv3
yCa0hX9KkmQ2jxAFjva3TvsosGOkXilXsn7naAyw9aUOSBfiaJilVo6z1pTif9ok
FGOPKX3S+Hof5PikrWDSIrXs5IA3OND6ZbjJ1fToJREes/5Ph81xNORKqw0Z0XoM
n5OB/ZStrrSIW6NpKg2LFA==
`protect END_PROTECTED
