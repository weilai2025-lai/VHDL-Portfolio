`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHxqxIYkoVYQawT6vllmm0B9Ain8/DzcMrcD0R2ySEtU53ymc1bItoty7jj1/tGW
A6X+kRDtnvBQUJniJ4sRc3ymDBX5LRGHUYcsOCkvZiprBpHlUJMzBFdZtPxqLZpD
rWGfuScqi78tYnuoADscR+7Gtnjn0shvhnLy0E8KeNhv0ozyJygEZXxaVVU1+Y97
K4U27cpK4Xn+fLQiMIDD/NrRy7yL2rY59OGsK5UlJ8aORY7D/e7glHd1WeQW38ei
5EVVdnMV0xpxqEXMZrwFclJyHXOX6Kt/9OaJpGrMYPX5VqGDV51o5c/U834gfxl8
uSjc4c2UmYsA8LtqjWYn3jOzYqYElhW3K1ZV4Jw54Zy1T22DDVdlicmKj+AqaqYf
ECW8yyecyT46RzLOYlKzYStA0lrCPtQA6+GaV79z2TeIts/57y3S0QsbnDnze/CM
emMkM2vBeyHA6XlGhWbWLQAaQ3X5BiuQw+vNc5ViN1k+w+OGI4taEz3EGBQai0vo
7PK94LfTCLIEaoXAs8LmTCYlYaLqGRh4ao/ZVd4pOY5vVc8Ax0IRQse9EVM3Q49D
DcAl2eB3Z1EEfC3epvEGwJbenMHiWu5Wnf+Jc1LaUaJnsXCEkrXal1QoAZo3JQ5+
Liu5xlSWRUL/MHFQGA3tRc4FX3RxXUs35dOhAOYENfWWTObTVNIjZ+urNK9E4BAQ
MRRVdLh3g7grax/0dIjrFmKs+v2aODx9LjEfimJJe91jfb9kxWBg4pYlI+W3Qj39
JYj6oy04K9Iz1BaaBnSKnhJ+BvGfYRvLMmlBzH6m16LB+Kf7UJqpvzt2bZ1r7eJd
Cb1oF0b76fIZbzgXzrdiOHfg56Ou+xIlZkBfjh7SX0i6V7XuKwksO+rWu8qkQcLv
j7a6/GAxIZ5YuYzYneSMHP6evyCE8qF5F+SJLJlYBRNvLWfM3HBJaWnbw61Dgkeq
B5s03NG62qjc4BhdLvC7hpV+/4ThJcpzFdMGKPznlJWxIakXg+OMaznJ3z3+UY7j
oowyaSUK6dya12P4dCM57ZvSiDSh0ITeTTL1jS3apkEHQ0A0inTy+usdvSkF/WaO
M/lB6VCQ5+8hnFuXt4gGjwHZslh87mNGbzQ1QcM8sEWwrNStJP9fCx+goMQJoHyu
GytyR761NojcUalHJFW9/C8x0c/MlRtmmyjboKNarSWdWkIs/KhBM2IsiL5qGFrI
4iZNS/6NnwieaIGgkAqEYMPpv4hW4cjr+fSlC9b8igO/69o3LX734RyGWv+GVyRv
fLoU7PxwWBuUUGcoO9SJCYm0Q1Ptu5+ShxHuDpvHQ6xOF1esRebKY88IG2fJbPTU
AkPUZup7BRgIsVPAul7sqP10MjjSKBM2MxAbyWP1V48okmJyqprduPfcuRF4A1Xk
gzeeqwqhaMaSQHvU3IXszGlaA+lfqkp5ZVcWYBIbCjJPwbts3vX14kw54cHfyoCo
DCgdBlmanT3tpxd6k+PXp13+BrghxGB4oTXBc+7TekrAqNp7h/EBqYS0B5LkEnFF
GOxflOIrQkY0VQ7Nfx5w11xYyNGTPHwey+TyaA3rJnZatTzmdyn/bbSanq2uPTrb
wWps6HIo7PUKKGlkPqzZVJS72NlwoUPxSe1fiNVuyQwgpKuHs5H6mGVGSaNXjlH3
0yfqkmU6dH+ANcnJVEE06oYbjdPgUp04XNnzME2kEClSrpqFQ3xID1TrurO5m2dj
dBWKgfadNyUVhNYCqmAWnZBEb7VjsedDz0o4vUi4TINKtDlJWNa8nczKwxLWe4a1
eYq+KAeZamkHmXpmWuxXE+IAVQxoVPEhoubXNlKDvWCachX5qOQLHjZCxmsZiDyM
IwCh6nL6Irxb/cZVLSRHmuPFGEfJm7P+pS8SaHzDckKodFzfyyBUVA3lorwjMrkj
gmtpfSQbtJZh7UhKhUA4C1FX5UXYkg5GRUPc3/gjyjc154sSvel2O4yisyqnA99z
OeVlmrcdns0KLbld300SMaO/LNMuQ0rg0lvQ4YEwr318xxkajn74RUX6E153Ge15
H0CsIZb7/Kbm97vtygyxEgJdt0K69GevFe7n+TLm2WPoshhWDF8xl2Huqz4MpKKG
Me7XKexvPImC7tS05hRuWgJ+nR1JMa8Ta6/nQ5wWtUS/OMKrcHyMbMWYR3C9rXB6
LIiwqi/fqxZLu3wNVB6oHPpqBayGHKmTDq9PNl7wFFy4xdmAea/GuTsfBcKioeL5
JcGy1BG2BFx5XqmcouRWtqrvm7giZvCoyRFxC22KiREICI+HNnFxIiVigvGfGFXq
tw1nHMbHWxOpZSVyL/C+SQ3YFxX/NVb5n2HtnjdhuB9o8srFM3SFIRXV8UYndZsV
BzDehP1rCbxxjBzT1EinF47lzmRYlZZbr7u8C9KChYLKo5YK7zBh4Xvhb2cLnq0h
3ntrzobtHO9xggoprhdN6rd+b5BroDMhJj3st5wL1ktuaqqOS4Me92/tnm9ON6yz
WbxxBRkEHYBCxRfnBK9Tns01wxh8hv/HGOpmClosO5e2AVzN+YkY1OPKJ2ZuE+72
lgTBK65tOYqGrYbRKB2D6yqZ44XLd+pThJffqhCJIqrosMseFmOX4h0FqaKkT9/6
gurJKSRPtI0TUjoF2Odw7+hg07fyqPwo4Bh5R0W6jW7b9tsgLBDfk0sb7T7aXcCj
WznJlUljUpRbM6MvFFXx/f+yM8i2ol6jAy4UVjX6IDxCCR4wvBpnDNMT0E29BsJe
DX8HpHUxV8duWTMuJ+GyWq/Yxg5UWtxCf56e/frRbCEoBxq/sYR6jgzrEuw5iRxl
VxRl6TP7w3cBzd/aJfXoTxXYSq3wJAvgvZGytu71lh2PONJmJEi/AYKzC8vOQ5xo
xVgphaLxOcVNl68D6MAjhQEKO7opnHm0nr401sPx6PySTsOz+lT8qfFezIkem4Fi
cQ8kA6qbCKt3mtFtePrIHEvKbrXUxGQ2M8ce6eO/zKNyL6ZlFc3EWzzSWpPSIVQm
eqtDiu+UjYGpKmKfS3bHtuIdh8UEvcIznCmQS2dKA2zprVcM7dMDtpLnqhMqxFR9
UTd9CEEq8vLNm8aKtZeUnzfG2EnhjX36Mj3pKc2krcQ0NViybmbKcDs6+vm0NZuf
bvnu18gSWIAIXYtrLNpBwtKV0abcJV9DgDwHM+iPRShJzDzk3gJLtK+bqP4bHroN
F6NophM0sXpDe088MyzV8e1+UKi5fuvx95x+9fpLGl1/Iw4oe8/QEOaUTg74QP5X
3BjqsBsNpGMj5h8x7zf/yv/0nMc44/mRuAgU5/tOK33lv8D7+cUeXFK6rOtYNrIs
mjK/V4FcMln+UOhw/RvhI3QXTgTnDPNvy3yKbDReBMUblxciJoXoHGdeFN0qgCFG
gXVH7F3O5rDLdiw7JjWLgJaKJSu+AN8pQVzK3SzlTYRhWskUIrD4Pm5mSzOIHnBe
jHuRs4yokjIYmzbxu58NfZSzB90mm5T4WZ+Su1rwj1MjuivNoenesVBQ2hxyn6+s
tkquPlMGDGX36QiOk/3gkf9OoIZ1FwpI2z2U8WaLr/Lgrzr9nv+/sf3HI5mAdHm5
2363s5Ps2+9TyHKYhKfI9RDc9eK74vk8oHzW2+MZ6SJgrNJSMxaXXpZsDsaE4XNz
AvcA622TxtRGUqrJlcgFdhTElZ4Symk3pEvYWgBREhpflyaFA6iMADIY4eTJ4LuW
wpXOzZCS6taCIrlk04Py2h0AXs/OMRCgN3ihH56t+rqqD1W6p7db/yzJPKLIbprt
PmZILmgxkmxjfDOvnSwhTEWWKewbsmiNmGdZQ56XEx9ghW+XpJ4pOjqtlmvTAwu6
l5hFtieLOVUiHbKIXkarKrnT/OwbWtMMDn2qoukph8LKQ/Eubk32S5y/Id5WNbXz
DFAOrGn4yChAa6y7olzRI8d46hEUhCNb+QjeZiSGe7IjnlLgg6BZqR/lcYvEhVYC
j6u40ruNBEt5c0Y0H11P6doKcncgVo2egPjYjD1ICrvMNMmLPp8jqmtOi5pUvFIy
avuJ5LyWzyss12fjjh1IMgHfqOD6xGV3jca329cPlivk/Vh99QBC4rFG7gHW0X1p
1Btop/lO3YLiPfa0EP+p3aVVwkIozDhcmNufe9ksKlGJg53Xmqn+169brKzMgk6J
p3TNxOWhueVwQS6hvYnkPfiVqOZXZrDKMBBdvIZtF2V8g26HweCwL0ai8Awi9wfY
0IvqBQf27WGi954jt7MgZ0JQwNKGirUQv+zqKo9Xw6IdwSZyhF9tn1ldh8sR9NOs
WGF7VkrfTw/aTUhukdzt5rGw/zol/7S4PtGiCKKdm4m1JaU9dl6jsyVTeeRlE+1E
fvwNTm0WlgQmvydNrmzZwAZmNTxnV5luQhHES00INS8/4Ozz3aiLm1A2RUsAt7jA
2INizndhQXctry1giTvhEkh5r2uuRDlUerxxhwgXekaLcB+NQd0l1NTnAeaXkmW6
EsLbpwPuRu4h+Nl32Q+P/GBAeiMgg6fZfidUlHuyp4k3ockY1UOvRWwCTqV7WIvW
jeb/R7TTcb2sFDuqccJbp9uHBSgSskY2UcvghPRx+tRDNzg7zWCNVx4VDbXiXJcR
L3OblPmL2QFSHdefqUuxWeptnukXgkwXr8O+U6Nve5hsO5dMAhQI8E0RWxGwRpW6
8FhZi/wVLInVLl8rvU4TWW4BW96enNxMbntFPjRXwFU8idq+hJOvqW96uhROwvBb
j9+f2ALOX7J0VFz1YGcBGlfz+U9GwoFs+P+lx9rASPw9OVjOdTK8T3gzNTH9e+fT
Z/+KT9iYQ+3Nhbsdw7koNifmQxxq9NkgEHsJfyD7vjzUnO/6jH4gNxFC3UhMLdct
+bOpfenZ5foZ0Hj+CXMCLTuzgnOZSXJLnVvwsaSsG4tZftHwS7V3629ACgQFbIay
ib/1ML6x164klVrqo5WQAJINB8fXvGUyLlwng07KpYINT15OmZp0L1LGTKGRg8Fz
v38ejl73AQVKw2+Bz5nJzad6mYJZdUuubwboMHl+Dnwvkr+8/JOb13AVXrHcvwDP
tBeWw7hetv/RQEMGBeXku59FGxgOLEqjnHsyy8nrMFF9fQ5ouqAglkoSScQ4oQJC
mglD3dj9/Xo+BgVA5+zC4GqIvpeswPzupKKrU/JErmfjPrDXO97zPHtAoa4uJqZU
ZzIsw9Nx6/1iiSl2a9DeDHTw3TimQ8/z29soUbsDDzRH0hIlDruI8ud2AHcpCJBX
/KQ0sxIAHOmFPRivkAc0EWoRd4hbMCI3BKaEVpLQKFsz0e/D9g/s32se8OZZSP6P
1PHoQB5NqbtLxR26BBu6nVT4uJDngSvLOkmfKxJh2k9Vvd1w/wMdJd4U7LStgc5J
icE8G3sitO+COPl7x95aV3PrOC2mmo/YqOvnzD+MQ3ES0wKO5pvwyAc3dHE4jKGe
DoPaneu3Ju0iOSpHd0Oalvf60uRaz4crBzNrDBhrwR7Q3bKI01rjsZPI7IxYjcSB
6DdhoYLlhDTWbt11aPFDE+BwLTTFlhG0PM7nSaoa1Knigm2ZEzRouxzDx89ffj2G
J4+HYSQyDa60hLdW6rb/GNZtuqzm/BCHvK8D+q61Q/J47f3eIoEBHbTZfZWwIXf/
V7Lv1Z5mJ9rKBd4RzmCI5j3jAfT74lujS2G2NRifPywucjoCizvXLIDCocQ72NGA
sPFBjcdekNEIoq7JGw2Liz3cylc3UvTbMoKHyZMLA0X09QF5N7FK0W/jAu8+DOTM
fz/glWebn/UgzLkoNSBJkzpfOepDrQDslnMyMi7eDSjb2BulhMqeifDsul5XCQ+W
gEhq0+LfrQ2rQFTWzpGCQ6fDe5HHTKDwgx69OHHMazH37Mh6mr/sRTVEf99m8880
szGJUjSllxph0aIVDjPbLM2CWO23bs9XfTC5gtyiYq51VNJeenCGd4u3BoETgkYL
23WiiO6HDoi/E1M1hV87yM/mmKxM4UT01e75QBby1EINA+Ja8Q4r+TeCNK0ieTjU
wHOoQDW9PP8b/p205acoSSqXB00CtyJ4DBBj+Oh8ORwu5PqYS/UoP3AH994Y/UR2
5jbD0fN/O5DgwSYbprrVxW67FDeFwRcXv8B97AHBwgamGFCuytoJDI4Y39pGDHws
PO24ugc6ci7mo5CR6LjkVveCsAbmkyyEcX3jmDpoea4nAMNAFfCAxNSROvAfsqPt
ig7+G5ZdRP8E1yYxg+l7J9yq+uagQKsBX6StsVSqpFrTx6HLGN4oUWNHoDlO4PLo
sgj3L18tUpovRG4Ata8YUBaR9ZMrVlzqZh8EaoPxeSMAez4SnerJMWOrWoq+ed8p
PwJoPlvA2u2ij7dloeo0HDTRRxoTZFo0hrVwNY1+M8aop+gT7XD0Dt1wRtCDmB0s
omX0NmEmXuMuLTeCLc2SnktRixqksOFR5NHMiitwcmn8TTMepxnO6QvHzDcDSw9C
bA5aHxpIMvkKcPmxOOkHcKsY9zjo1V3y0chBsu26Q/YRfh9ly93SrbE+BwoxR/7Y
ebi4f1hjBSDezGbd9fV/8uvHXTH20bf6Pwgq7OlLWuYCYquXwFVP+zjGY1WkoJDd
c3mCrYGYQ2V33Lv71nfsHayRPpAE7Pt7BhFlvbkrB/2YnEXPbE+2ocdVcw8CPLao
AkOursBL0/NESEvxlZZNPvxXwHvoU7cvB+HIu9TbP9UkMtwzAbElmht8Io0r2cXH
rhiFVOxh2IJl2cAf5LqcHWIcnmtDI87XBroje8d76kbhze9mCLDxPqBBA6+CVVbC
stpqjZVdiQo+bJOKmAsQ77lgskMgBic9OfCOTu+RcbWESukUm62GG4jDrwfIS9VC
WnWYZsyl6Ol8P/Ti5GvDi4v75jB6MfOUuYeUKe5sEiS9VjCtNtPrf+++ijoXz6RC
NyG95pPrkmvhGVXHewo8lsgLY0bVQ0LAC5hfeYUqJl4pA7vhz3BbMRW/BzKdi8Mh
BzX/bPIs30LuhStrPxJ2vsVewM6FTY1jEkEh5Z5c0oYsYGLRavZgT4m/DfuI8Mux
b9A+E9SkeLGKPVDzzayYreRCg7VXHN7x90zedK8ciZALB4ezgZKoZZVzLd272he8
lq1dLM1bVjbdaKrTJMvcyjcdzO86mpAOtFxtDFTeaFauEg7oJOYvW20qooKeZXEZ
duOWkiFny6zNhgnD5hUeuWz3Aqf66fhpIzjXJX3BkrMUu/i/rVbGUJwNONXMJQQw
tF/0/f7cBVMSBHFZqWdEqP2cdR7ZWmkZIhKlK/GsfQ3WkuWkNKn1RdM6GMhpvaKb
C+5fJuZs+dT3z4yu/dH1T/x0gsGFUTk6w2qEd0labTwqOD+aktTDp3IZILysr402
OWs40RgdCHRYOcqGRjDeYASWoLRzfpdYXC2LM/YEouwEawBu1DydhNsAtofdVB5t
jde4F+CXIFySnzgDEDa+ILIColkHWfj3aC6aFNqNw48a+bgp9nK6L0Wn1KlofEIL
jLJ3lP70kkSwZCKt373sG/Z4pxziuCVL73WRM684OkKLh0KXrejZaCdXFod9qi2e
SfhOjpktvX0eretfqGnD5lHRnHNIrj9f9kN/v+omqLDVAEXbWp1Au2fIOycvtOBb
zmeql6jItyoxUjYOrTxahy1s+xy4TUwTSP+3yz0OA601paYpug19hdeVTF4bOnZE
qc1PWXVva8y9BF9vLn1B6VHFMwCUL3xhpR0j9GkM+N3QOimRwZ2QJi8Ss34QnCgA
GQYu6vq+tKVAs67B5qPQSAOUUNy5SosVqv3Ui+1B5j3HM4yxD5+jsnWbGwUivagV
vRe0GkRTE4rm8ByjiBAk8d1UqntgDsjzuYZGMjsFLdIovBz1t1czJBj14Uwe5rxC
mPdcLx6uG0TUV9U9j8knxHasQWP/L4qNtl1vTt2cCBH2lzNxI9yMG7FeJ5gZMj11
RxdSRs0Xf7W8+rQFrnqZJHtG2CGabcyiRl6CpT+RPHmrhg99ANwciJDiPeAMPJlk
p/P1ei/1kKmmTXtNVHlxUOr2BJ6J0mhl6eZus+tVTHPTuFh8Yf9y9G4ztipYDeix
3nq2lVC/Q4ayg9rtNNZt7JbNiukygqGj8G/MsTFj5v2hYspAuPvNqZEH/zqlCUdw
IbOIfpXv1RYfvlCzpNMSm87J38KZmujbIMI7IgF00kVp87a5mIk4lXB7ZI/e7lkO
FIOSpjB4N3M/2dCNRCJQTECnIYgdRKFZIQCrsn6W/tmHasiqSvf5Z7z4MkmS8v4n
EZ8nBdhK3ohzGo2t80fb+Sr9fKpSFR9aezDvJDCsP1Wyqkh/8MQcTDscH2DGcIEX
I//Ep9MA5vjtoPfEwtrskq8l2uHe0XMEt0B3VjzKBAmOq5lNbVVG2xQqLca1oBDd
bWDMkmxTBQAQVJ07ACWhs+EGeBTbETD3WlgCqB21vXD7BJ0c1e60tSyFXQQt3cVh
ZWx2EgIuhcG33Ebe3yDYz7bulxh+kkzASXXVgrV9NnwmqqRM3YwtMcaZISuzPNXI
Fddqi1e3HpjtPnZo8iy3/m+3Q9tl3TN9+vznwes7fliKW+klmGuRL2Fr+FmuA8mp
WApWNAUZCinNwo92JjtkfT2Jk/oAJa9Hqe7OdGKKJT6qKSq9CeeDa8skrER5BHBq
5WBWbY1gCbVu51VoeOyiyQ3v3vbwyDM4nP86LxMuQOjNRhBcs0IGGs6igCrovA89
S4DcGwIQgRwpmsJrugxVMMoMu9qiGu2/pBxzUZeQCtIRFa8uu/fOPfeK7qw2w1z7
BkpLpB76VA7AYxAld4cllQrdnSuq5d6Sy/IO/s06ZTYf7WRRxQTEgLvy8LbstH/c
9v7xaMedc7Cd+vRhX0kf08FPDuZjZX8RBUWcAzbJV/AcND+2XCuv4t2w6ImPXGlc
WWgTULm3hb6NEjd1R14WFdbA4GePQMF9H3eqCQyz+e5M91EncxAH1YKyx1SXAzN8
+Aktbux3w6b4nbEnJiMqApI4j0RpyGF6WBgyi0Mq8CUTJiH/QjzlZgnu75m5pz2M
7kih/KWrmGuDVDFmtxt8EEbOlMV65ZYoN0DAttlS+AfFbFbJG7W9SnRNHoMS6yyJ
K9ah5TqIv8haWZsM1g0RS2o3ZTX7VNHZoc1cIR3u9LXTWG9JKN6U40Ok9CgwT9Xt
Gs35B3xeul7XGBnarF/+pwFiAxUQXaJUdkmE+7nlzSFVt74dnz2gfNLhx7O6xuOv
GaNJq8mrznVSH/pgrtzMFQ58Qw1pfNMeeAt2lCySxiiY2vjVZ1LsL+gz/vO2fRdO
mJLkt0UB2PhZjm8zKxPH41t9nqpQBjgKBQHuNutB01Dj5Ns0Uy55p0S+BNcGSLSC
oysbwLsEKkyZeViEUhhU0wBXHBOjhVQwoQ2pFjnTBrhfPFR5ZNJT8PToSYtUxj9j
P2eIeLes3udhYBpZY0tYJNCcgGpNKBiTfk3PmrpEuNpLHIZEeWB8aq+auzOaspXp
jbJqH7ExEp21JVaQVvYUzyFkrRkq044xl3ennGeQ4k0fqRV6yrzLrsTIoUeATdG6
1FH+wUlzZrfsuRug7LQvGJnFRl5JZzSRhD+X1/nt0r2WBglF1oqKLVFrVGFBqidi
l3rF964bMbLH3gTXiKZeMovgrBbjb1ucbbCAWpJsvdP/Fr1BJfJDHXt68Zzy4UbS
b5iyjNWMX0L7mNOR9OKHFKku1c82zukmHEMXXaKFT9j9Nc3Mwd+8sbK62QzTslee
7fbPt5SMFDQ5aCm7FA8F+8wHW3re3ySwPmncnifVlsMf5tDWR6AhnjyYwXWruDQv
nUy2itjRkxc0JNndVRO9Cm2Uh/C3laxN71ADDrwV2eEzRxoButDtpDAJaY/6G69J
NeVNLjfow7/739KBrQzQEfM6cZXGbUsSWvCV2IiZaQZ2/ip6pj7gfLb/HralXY3m
HTkB91p2MgDXVNo2UiNgCetC+R6achErA0EtgNUMgYgEYAdoMB9Z8AArzV9pidPv
Wq+YndylV226F4/Y/3vVakZx6jMlO5ybZo7RFsYu0yzdV4hF/kG57wzejkVj2c2+
LM9FQN9kC3ctRISPZeWvaybSEnhlvdUZZJIqxvjgEwXsZwkQEoslDG3HmnDwD+vW
OA8m92n074Ro2+wzKvhaG+9tbRTqLN6D11569XiVd9/RjvWO+ZLBtx2jevz8Zev6
sjkWtl+jo99S7XEWw8BqDRvlKRFCZit/TnB/jfHw47L5BrbNUm2a0TKE+T6x5xhl
faieX1FvVGkXo9Ueu1pMA86rBufjTURHTs1HkKb7mGV5Wj6KxS1v3GF7TxvIsdrL
J+b8g65G6id2rMM+eEc/FdwNht+0lOIZS4jeJPuqJvrU1Q0RQ4DF3cDDt2HhB88a
09AXRi8K5e81P5Wwcn4atX+NmiFej2FaMOIM9lDGKigM8tsuA8m7r8POjU/lTBsH
SmEeo8fZryv3gmPXrk6cTdW5D3/e3V9V0Awb8b5esqD6gwFr70XHF1yYfNe/L4ab
/SpHlPfpwE2dMihQch+ETgGaFsm75kwoDM1lyOyQtneXZiPikeHTKo+ybDtShhc7
Yvw2XZuY4IEjJ3ApuosTTs08CxvQgz69UxRPCWEPe3nbjimVIvmmfNZAdBnATb0i
bxkz1tERgn/dR3UXj0vaylJ/TfhOtc0Kg3o1Fc/lnW2nu1Dp8/WKyDaaTnpOMZp3
OTxVM4MC8Rxxw7UizUbgo8/m5EFY6Co9HRabZJ6LuTzRleQD2++5UWn0qqhGDH+M
xeaJ6sTEOrQXrGMgCs6JygzYaTJOqJ0mSo9zrxZ3Q/+URUa9sOTGkfQiG3W3RzBv
eRLah5QDxmXqz8D5ytq0UN2vEb5W0bEH6aaZ5D3dgMPUc+kB+l+cnWhlMSJcxExi
K5xVHCuGXpBADZD75vL62/PUEbvT46j6Ua4C5ACxES1i7BV/AaHluMvw0+E52Wls
oRp2ypz01oJYxNxLQDxPIrwk/2uVsi2NKcfhjlIGmYwXc7GKurGxng2H4ijMtB+r
uxttOEgyTruj4mCmu6Wwsn0Ir8n4fFghu4YJNbuM1B9YWOFIZHUe0gV71dcajgGp
HobaFqUqCIn55KzSewm0Wj2eH6iUkycG3beOkt6V+RvNC1Pkc+1R/hhPby8/XTHB
rqbImMsYktJU6XuWicBA6i8qFo7Zbla2xUo7+uZ2+oK20Ex3Rnkdrinvc06RKd1H
zN9UbGUk09CXE5urjg7nPypOR+ZWXj09rIG3x2BY0XpakIwzDBFJBMACKip0TPe2
VUVsOJU2HzcGOaFIsrwNI+Soj58dbEc+1mcRJEjYpD5bBEPP//lTaVye41ciPjEK
2/kr3ayA/9dM5o31BCrJctetM5mJf+fvsjh7IEn2NGqpD7gKBUQ2DYDaIPoaNGnm
m4ctakz/dZS9DeeF9qdb5njhcfPGMIscbpQruyh++ZaigTi2xclk38oo2RcI6Yvc
9WAR56AcGsk9t26ipS5ewI4iwb94n5T//OiiTsq2REWhJF3KfoJPVX2r952jbpNo
egCgVMeyuSoojJhKYiO1uYa5ESMDQFlGN/53ZiPIJk+j6wZMQ9CS/uTduBfTkK4q
pxHmouqXyABmqkChULZP6rc8okEZnf/+jse1yb+cU20oneLr6fCFNgpA4oT9DZEx
Paf+t5HKVTZZunlgNv14Oa5RhWIJA5QjYGx4iJRHGc3bej47cSymoNjhKkKkw71U
oV3nE6isTRrbKzwp/8bnG3nhRW2deIxNkcrSaezI/3WDFnEQJ26vlHVxjev4WlMj
Wqrz8iNmpmUEBvIfYLc0O4CnOPTuMMQrW1KMV1LG9nqmvrHVqVC+g9s6FL8yl70S
vtyzghSFIpc76XlJbm+QthGuxUm+hHWeLrSMtS7lXry0RqlEJvax2mQl+m6dpTDN
3fEJUs02P7ZXvZ7JCR2rZwWe5PmXHNBDgax+oJr+Fb8yzGi3Rv8+pvd9vL/1B2BS
qcijrC4X/6p6g6/M+UGFQu+8aQbPts99MSkff5OLEaakAcnA0zDn9A8ItjzGSfqo
IBCM782zH7r0HjTd3zWDaogD5E0eomnDuj6VnRxW/XNtUU/FSqRN7qXEvAwBYmJy
QaEM/2IVtcT+BQ5QW9GAAKhdFam6LPhrEBekEBhwNAO6Z70dIbKdV00JPKl5YIP0
YXes5nv1EC5vMWoLzT6JW8/16ixQr6dlR6SYX5fw5pwLo38OZ8mZ0AA51RXZPOVg
plXaH5D12TGlunZLUGMf8efy71/U0PYKrk5sYMFWC84n2SOH9DeAuo/+r+IPAOTK
t8GwMq/T2ot6N/Rad8keorBkC39+W9VWaKGtS9Y/cr24CMl7DV607UnBGYxr3vq2
iFMQq61mnvX6PHn3Znm3Uhl2yHWSuH2krNaTm/umOGqTYj0ahrCJBBcvQ8GjCuUq
SpfNB+j9dLgt9gRiKtWPMbnPa4Gw2UTUg3pDnEDdYjhCgMpGEkufWL9Ra/xGAeBw
VupKQw1iOk3Tpt+ZzuaGWe4mmhwRY+cI2VeNgnw5w75nPsIiYMrB+TZ3q3Vk/QcL
464MWrTsFy9aQ7e9PzcnJxg7jczk8BqgbUwokIOm2hitcullQe+h1s4ObaVIFVA/
NoWzaryi5zWNQgU0c3HEb0OrOuVb3l0fAnNVpCE4ZKvs/HOL/n3vtLhc8Qnd8y6P
4aXUsOtY8z/8t+wBlW+17wVQ0+YRuUs2ZFbWPICawDnV16js+52/9qDWUNfr3NyU
XANhGaLAXPa4e2tBJcPWtLJf73qowED4rpQIQvCNVFra21TRhdEwbQbjU0cSZ1iX
fJ5NxDmBHHG36pQvtJqA1ADzBE+cxDpqZrAPiDJWumK+7AidCIeh39Af6jsJyP7R
9k8KxTyeLK1ik8Jvf8Ffkfi1VGZBU3izpk0TK0LHYULelmnMiGoiLIGZqQoUIjUk
10TOS9ducrNnpTfOvsZZKr5WO3QakKfYK4NcY4tIG4wkPmZotGn2JKA1lqqVMyoi
aIRbdLRcXYhuA6trM502bdP1Z22VXso0qiOHS0G9Kj5Adgwy9LiLzpT7BYcH2/ne
loM5DD0e9GcZsrTwGpCLMzSdTJAV0mp8q/Kxgn2wuhVDgXLuQ6GWUB8LZp/YXU9K
mXaKLfrJua/wC7NZxhosgLjBhyBTDi58qBtxjYL3f3Sx3Bh67li+oK0Mwvje2I+X
bhoBIMns8BuHpmmIeLJvX+TWvkM7YGIs6jFsV7NuWvdtB8mxVvxQYRBqT5CWfa08
nN0GaC0WiCRzV5aeg2E7+ytu5kSK1lwVnTjSPN9i7f3SRLRC5sBg5evp8jv7K7qj
i6OT9K3LfFl406thCpw0TIDYhQaglraoma9hiKsd7XuTZ95+QSurc4jTnV8I6sSE
8BX5V/4g/W/xBpeIj/d2X0xZlyyDfay4zc4BX/OaksPYbYLGBmQxjn5uDc2bZelO
vqK+A8y+iR0SUgfuVX38tiyOropQLe09MmOFm/TM1SlVqPNWb7Yy9MGlB7Ci9BY2
E9Oiw5ZprXZDu1jVtlOxFbTy42aQ0gXa7v+BVCUL5Ug9BPMfsrxq1Jt2yg742OYq
nIYUIfKU2bGAtl2zn3dWDBgra2CtSoUzhYjF96wbs2fLNU3KfCMhJY9Q14HqpRid
8vUVxaim0kKktT4lKQwWw511Xy9xmKkkX4Add1GlzeSJNv2PA8gdlRh/n3okryHv
QtlFmO466YBlvG2LyOLfTdOyKRvLXwzxUYO4hN05TTxtif06sWOKNyHDaMvcLGre
/K57s4r45Arn6SlNeRr8p8XdovnMT/lHDkIdUPftDImwAkSmExTwTDZ0oOu/RF8V
v64ZjYQfEqzNQDH+BZ+02WYg56figVeyyXD1onIJ4ogxJZLrTsztTzXKfVQS5VDn
2gR46Z0gT+iePuQhgmnLds/FuC0sqKsd1y/UrSd0nLSAUiNEZJUVdhyv9SKQunRP
XPULZgrPLqc9nQVexn25LsdYs5F041c2A4lGZNBUGdzo/JDSxi7V1jYcauA9W47F
qTCklIGc/3IIxuVSyql9SmA2+0mLkvZwqSlwhA2RW/jF+ihzf3T1qgRhl492BdQi
x74EglHShRZ/mT6r3gHXZsvILJi3cNiZL3a30uYm5qMZw4xyBtvV9wasGTUIdkWV
aUg4G0y6RBnaxfaV7QqDLUUSu9qfHn4RKnUWBn78s06Yao8r1VfZhrGqdjF6QAld
rtBuYbuwsUnC9kWAsXtSxJrr1qVZWQtsA7d7iP5ehqgsgYNhvnuQsdPsKuWJ+i/F
Ioo99SJsIvlz9hBU+Ueqpw7jDEI+JwVi+yHEs+KJHexa8Cz4EH3sBDdbg0z6UVhH
7VsykUjCSEWy+ig5WOzBGKlYM031rK79V1Do/MEPRGjjhwEWXAWwbi8ShF/0Aj3/
kS5X9YZUBuPrsSiY5k3z0OXmH1Cu9dNKzCwcA89UUFXYsQYS8x3JslPH0Oc2n3xW
XgXS4ncat4GjDTSm2qVgeFtUSyFb5xnHA/HJeQCoYNveGoHRSQRcgB4RqCioJcM5
XFTHSdTXpI1PdSvJSlFsi1/iAcyE5Ef86UVoPKeUs2nDOCfxiicKXYgmJwbGYbnR
xpAGnZoyFIrnUppHOofq3lKUe4SZn/6w0B4h9tRRxoEVRCmjRxFtAQEG05zdeC0C
yn2BiqlQt1hMPq5OltHqtOdoyD+27ib4yP5w0Wa0LSw5vfS5l3Z01txVBt4FcrSW
ZxjFfTj0KTZwbL74JfMygi5m5iB1oQWlR9bpOCdXvVuGDStcE1ZcpvTgsTU27bBi
lCDYsd8UO/5nlbPpXplVnKJ2weYdqx01ezxeV+q2VJWEc3N12EwADW3RNsUp3oNi
6HMHe/GyAV/Ukf3sjGN5jSI4u4ytQzb+IaRpzz8hOdsMlbnqsIJKh/KTcLZYJn/u
t3mvt70CP3cwKlAfQeud8K3Ik8XA1+nId3yb9O4nZPmd7omDxImhZWcS63YDXUAB
You1mSvK6Mdg0JP7zYcazAhQQne5uzxFYdjlNwo4QKa0gwjiDi7d20Q7miWriZ7F
75LFT1f5Esl5FpcwfijMmq5Kic53H1Uw6EmCI7OQgEzakxEGO/7IgtAUEAYT9l52
Elp57Q6w0la/M59Fz6FOJOlLAHMN8RfR42e1tZkKTuADnVEPZl5p9lYJYo2mOr+a
ikRfExWT1mp4zl2dSJw2fkdxavaV8VRO6UY+1CzYMbXqrdmMDIyiRAyMYWEKFuNO
vNbOHe1h1HTyx11vkzofviMclCUNkodyEzrvGvaFpfM6ZsfboocBR8jkGRfYqY1Z
LnHwWQ0paeKOfcyi6c0Ze0a3aUkDCZ6O+Iad3oUSzTQv1Q195bH0R1mhtb6M64Tj
t5UcexPiwy4auH9fEBxxwfYh2edweUXq4fKKJlH/S2JmTLcTj9W0JZkeTc5n4AG4
24rMlCX2+ruQGrDU5o3GTsbcL+bUzCXoPUdFGkU85+NYwFDGRWVUk2/Z/GaUu5zk
Pl9C438GTNyydjc1ZIGvhxBUsl9zlr/J/12k3P9i1D2b5BH+D68oQuUTR6Lb8mLo
MVC/SDQNdHUUJdWfeHCs74p6Y9AGJYHQLSffHUrGy0StI4M9RTd/Itx26fiXc65T
PnyosVDM+fuWi5fkHPzmk7mK5SKx1BAAegujzPUZbD/YsZsTEgzBSlc/zTg20Wx7
U/DoEEE0ZoY4N44IwxeZ5ExkQdHWJ/tzi6LTtwwRcW6fg2/HinY2dcKnzbGcciVT
yPGbBm07TijM1W991bj3m1w2j84JWJ+w2mEU4SRsuN+esfUtHaqnh0cLSBzTu63k
Diaw+uvgQgtX5q30QjeWt5OoQCwWp5KHuM8uzdwdPCosgwdfF6IJVAWFAgBS5HDe
eG5+A/kkmHbnVqPthKxaxEt9+PFZnw5V/7E57R3dKzEYYKTjxxyWMO8LLDCQ2jbV
OP8MJKZj8ycNZh/Mb4WwVV109VjgNyRnafr/+rZJ6V4LMTnbrlA3BVDrlZXeAFPY
+pnhftbyYHJRU1k4Zshu6mHvK6YkqrsRDa1QH9fOjtXLB1/96FnVexigHBFAs5Ka
2rc5V8zu5d9K51qEABQnR2//hgOL33J+ChrAFQiAXM05a6fB5LJH0llJxIB1mJ9p
Q7Bw3WhEeBxCkDvBdtnms8geEd0tBYPZzvMoYbpznl5hrQ8YapRAzZ5/CmJHd0aq
p/OCJuST9X2Ij1XGAiQIEnBY0TEtpTMXYXmjkQeAGbIu17XrWocLrrm8P2tCCxe2
fMCcXa53BMHrYa0vEOz1GAAaoB5yq9BQVhJTQCWdh8leWb2kFKb6UFD+RjxdtB4m
ACfvpfuITkdWExlIfXLA4T3fkydnWCfrRRouamNA4doahuqwuqq/xyg0jD76qR6H
Old+fDn1ydxqWZP6z5wswY2du8GdoCNYWX5cM/QbpNw8DzDUQrqt2APUE0Er2KY2
6iyXAPWlrcP0fNZuNM6Ln9JVqJRJXz4knJ/0M7ZyrsUOQH5RuBA952mm4UVHV1XC
1pqdLB25RN9h8uq691bPvBmT0ZjUtKeGeYTzwGeH7zSjqquBsQYFw897Ly2zWgC1
loHXbFYHxzoUkHYbZ3Fy3i97TLUY16oSD1wcbYNm1rYRdv5f2B87hd9Pydi6BmcF
K8AR9ebMyT2/AEW02KyIth8JKizeS3+hxCetgTx0Z3/RmZmfE7zFuhSjQe/jaD/v
EPm0WO0bzWw/+V0bvQCXnQ9r8JCpgd8NuPpvzxTJmzOru2FaoxtvYWb3gsO1FPJK
ma++OQCjR8/2jRkQ1KEDXXHnvPEewM9u+vRx9Y/SPOHs+wmxsySobShFNfOt/Rmk
BRQ8OmOgYfnRZ2tKamlXjJMv40JjF9W/B/1BzX80qBdf07Hrz/nk++b2CIH1Apyr
L8UUTp1aoCdLqzSh2qGtijOW4/ymAH7R9//dRZ6sNyHdU5yIwbZuf9NnbG1a8JVC
fRou2N/0KKvUXcsqApxolvzhxv+Q0uj5pPTaI2veD3785qyKleKw+tTo4cO8uA5Q
ONXDhGk2kFnMUMiT8pYQM4IMxlW4FMqLYUOtS9VZWWojgF/3qSUquiGBOHPNm07y
d5cFQeEpso8HsFQJQ+xsbTJkSQzkyKIZpq9jcx18pKYOUDIm+mtEHh4M7JodIbkN
UaU7UDLYtlM6c7I9unY2GzuQhSyHy2I0TB2FqIG7s+UIPoGTVHgUq+DFQ2LCcZCn
OCUPLFPSd47GxOtf1LWwxLz2SUNiusZ0Gxq6+fE9EJz1ZdT6+VFPREGxc/KnTD71
1QfiikEnfR7z+CIxKr/fwjf9gmOOUYTSzyYnzKa/MztY57GiPlPhLrdP19xY+YTf
Hw00BY+VY7WKu2ctApCmV5IGvrzVpLzoJpqv5iH5GNDeODgBUoVKtfkZy6s8Swwf
4jQjOXYh0ln9WmPNIXCls1Hc6BMP+hKs3uAfc+3o6EBHvfL8CS2ZC6yWXR+biOEQ
StVXnsx1lTWIC5LDsfelFxgzkDlgg1LYUpWAVfoLcX+x2cnu3hQLJUjt8c/nSNOY
fHXFVjJ7tDG8/OHPFk5LcZNOwBsnPFb7siDxKEoA+Tvbe2ScirQG0a8KgZyLDYCJ
3SUnoDCYja+0KugtQLbYNv6WxeG5q56aBokhNVJcJAl33XlC9bE5keo3SilFqs+N
sHFHst5GYFZtojWlKPEjH/79VHVGqU4/l01ICJ85j2CLWXBw7I4BU2LeL+TyOG+A
7GozfYjKDEt/Xsal4qBbgOK3M6mwQAv81rVW7JddhVLeuYFsCydSdCilbpiCVMHu
MJ7MKTh3iU7YP724FEDHlW2ph4oZEep6ImR4HH43JdScfkScTl/qt719jgrYISle
pGRQqsgIBnwATEE7GFgXOpsOnA1hW/1NgSN7I9Igkmq/2PY7FpBZqQ4l3lYEji8C
a6G2M5iIoAvVvAOon+J3fZGJfJjNOA5WjbMbZ5R1XweGQwzpthQGRa29xg3i08tM
E9GuviUenwN3ix4vrV8Ml/01gpqCkQrdrgHsKtKZjcYG0S0AdLwtVYFpytvyZtoD
a7+HcpsAlhDWIy3bT8/ZScX43OEBwPLYf83entaFhHaNffMkjsuQaRuo3nyqdFIm
TGx2ZSydK9KtLKrHHDo+Yu/xDUscVkOW1ezY4pNnL4ZwQ+XuvXOo2nzHSTYJJd2/
uIAiFn9GFkVrJspMyWctyNUTcSN+s9+/JS63Fxn8CdZ2O6wBc54TJKGD1Xe4vReB
V8aqjmPF2Ilw+Iqfg648oF2axpdE0gMckdZwhex4toPQb/wVYGc28lpldSUn772k
3mPh9o3vzG0WhZ4MJXbTCIAxbex/bswKXsBBXj8KmPAWdiIfOmFg4wax2Nc4D2Jc
fq1zF+vmqHzTT7TV5goIZIsIOXBr2QPZEc+OOpgboYp3jwfgomAMcu34wzz2jQrL
Yn5+rverYtUuhirSZXe7TfGqPpDYoXJ77+f2K45iwauiFsvsZcrBq+DTYjfSjxVL
Uz8IHf522fR3qqLKOnVDk1Vl7LvyVMaSNh4bC6W2Lp1ERI9b3If9D3sOJGFB+oWp
botzj3LLbdr1XTFOpVmObEKAyvrKw4pJyXykD6St1Wa5yaac497KSji8bsC4NMtN
Bm5sLTpBfe0yPRQirmigT6xC4UbDVK/DlE6EXsRbmC3v2FanuPgXupn/4vVK65Th
DQ6EGzXr0dy3nujuFIE1fGFy7et0dIYiuie79E5CUurdM60s78bCUDeZdYsHSCRC
LfT058wqjEkoE7Npy7VnaSgEH/ZsSYYrnbxSuuibYgOI2iNcjZIB3wcdi+8FqZXk
KWEedY9qsZe3ljV3TOEoWIvdz5511nP5QuUiDhfRTX0/mtzX108DmX7AZNBrae9U
BYf5RlYx9v/wwZ1sXQeHhhsnZZnw5g5EoX/IDod6DvDA9EniZrXg8aGDny5jUIoQ
Dbtl3LRymaCVzes5jnIb7n9nE3wL01WpAk1/8itdi59kxcdM76F8GJ6NwSpDwezc
wGJ9rmal33Lfs7NYcIMvjOdPmNu53VgL/v5RbJF6tyWk6qdqh4wA1/MJS0WbFdwg
CwLxa3byyv61dLaFbwxWrDl6EuDC/gzIByanIajVtW/azUDIBlY1shyuluSOT6Vs
MV76xWq5JRPhX1AN+HYYhLqHtHDGYNo/rVZVOdHUkkZv0ia+kkUvw+j9cszTIS4d
KV45vcXiGCAoausDy2BoCj6Aw8O5nhAq2r5n+RqZZ6kl+8dSYOZLU3BzCZvnaFIT
ZDH/WMxVAZxxjoR/8cL/1+vn2NvcIA1XdsIWH8NpeyXen3XHcnGshuiv9Tcw1tOV
Ct1bQaRclCGdAlLMTICJ4c+p2av0iG87ZY6EZmHxp+bp+6h/EQvxO0BeJUu4C82z
vrhOwQVqDT4HhvdUE88T1aYWbVa5VJwTjgmdj0LqwVSbrv9uGY9m50/67i2J74K6
ZEByS7wFOQ0wpXbjoBzTRC0IIiBMTHMLOaNFbOnsGHqJfrrw5xmZRkAr5NldeSA3
ViIuHxB5B6cOwOJTnUPhmIY5bwSYujqbNknTJkqUXFmwEit8mGkjqC63Q85MVysf
Cveva2otESEPTXxbpzYrZiyD/ecQ0OYUrC7RNev94EF4UUj/hv2rQS+djyRzM3F+
bdmZRlRpEMudyKsBcQsA/RCbB/5YsyKTe6+2coxT9ip9HdUBuUi0Q2oDEF4LEO6r
zzBrn8GbapQSKgpiiZ4FSqax453rMgNQk+YqQv6gYfmMPORxxFo2Le3jC+5Bs9P4
YEm3mYoutEsFtCkmPkqohuW6wuGkCbUPDWBi0PCYYVlTfxYodwuE3+4ppynZJ9/q
b6LfBsDHqGCcmUkqLCdLxFMz4zq2VjYMeTlqeF7rj2I+oRTiL+0s0x+S/kvMOVGw
l09oFSak74U8y2UyQBA09r1dblbiWmjicS88+ks94xUAaz0gzhx2ZWJeYZ2OF1BC
MJp7RPH+WyPFqUVjy9fclPSiLDeQ0omOt4i5udIYHm7VImjPOrxvG5AGoEdJJPWj
65f19EhiyU1fmD+YUDkiGqngkNxvydldvMiSLJ4HOVgjOl2EiILYQO4/ihzRaD+4
8jNsZR69G9dI8nyKVNGoYGQd9BmTlIZVR6ByzHIdv5/zGGRaW9J67VeZG5n1iMCD
I1fU15dX9aT7+nF+r3R7fJFYfMx18StZVzy7qK0T01itSGMWuf3uhvEEop/5DdG0
a/wldkpuIWtaEMEGgI8tHkz2TXFMUimWyAL1RXUkl2ds+kmH4K5DLlgoekLsOIL0
VNcrlWEgzBD0MdCrBNn5aiI1pSOpCD/JNqncNPIIiouqU/i2zjdNqHl/4i9jKUjS
HcvQP2h2eZPG6eNAfKEedYW0U43tIy+OlczlYjGZ8OhZdyeNBr0Q4y8MOc6RF/WF
/5HGuGBcwEEBDk6KltRqlvvF8FBWXoAod0Lz0+87IossOuzQuTCNkWBKv61nA6iG
NgHjLNj5ULKKKavr/ofwwR0pXjHHydgtMgXW0y7BOqupKBIIp27XW3Q/VcEPTt9C
vIarH9H3TuvTnUmAU0DDQQd4JbitN78h/q389YnxwaEDA0s+tAeI1JQFhDqlXF/6
mddFeRfe9BINGMBgncXESLDtny/nvdCmlwXhOfQUkD9CaIIYTAJRyUF3I/qjSgWP
1ZGxhNF1dwgdgIxjA6blszwIGsb1JETL5gs40NpW6UfEDceKJ3HHqSJ26FBsfP/n
jj8mVU0nQYBJHld/MzhRD/yZDfNzvarYUe6L8IpR0qK9q9Lmbn25sEuBdBdS0VG1
sbojBEmioJuUG5eNTFq7+ER/kO2mwrv12VyYsln6KckXm4vpNNm2MGrxKdOVhG07
XXHb0kTLlVuVngYV2sN7oYGxxOv72tsf56456HIU03QS5cnPLVoMmb9lRY10OzJS
W4EGgQBBAJYkIt2pBX2IJruFJuhgLThSAlUC42MnzPud5xKu4CWbM4Azt5oXAKnx
HTYcwQRndIcYjTWd9iVuQWyFbrQ0qfY1zxNqxe/naHC3pVQg1ilkcEMGIrN3upDH
36JxHVlwdZbY/dDHbRmx2bdersuhOPsnv3YJcruBdx1YBYNzDnHul/b2x0q9ECGs
+XDY+gwtYbXVnmmwLA+J42NBAkCUnYsAlf3ZFy44G/QAU8X/b47PcchUyAl9hO8I
YR+knrNhrYoS7nxZjcgYpVYBIsT1wA8B5XVQtpRMWvomFvw9D8b+oL8w3zaOBjZP
ej2j3RDpjSkPmRbuJMhQaXD/+5ieDg4hfGJrvJJDddTRejGbmrOCEJMp/mK/WmVZ
dKeA+EV6d95EiwHc2pmA36jGGRsZlUBSFXyV0Lm42QpX/1aHwLI2JnGwVBzk4rWt
Uwf2iqmtOhiKgHEiTN6azCj8hAsBYgtiRwS4Z+AWGV/rC4gKasLNU3p6NkoocDzX
xxxbQSFXKuWAZixdfyq4PR9g0Mwfr0R0eUzdLcTOF0TAbgibBDk/CsT3Lhcr8N5p
D2h9Hqf81nS0X96C7jNx8CrAzyyJGmupsUHkCrVqT0UkeLN9fGujlBLWQgxqbgqC
+RxZnpfdzvcvYEEgbSbEybXATCQDH3ae6vK8KBPCDvxhbI9PVZ8zyFhkHbgRujQG
OG5TBFpWFrEgGAXl+EEYQFBTiGiys/4eE+7raDww022AI5VoCt4v45giCEkJmczb
G1Xy9NxxGveY5o07e/r2QIqOYpmf0Y2lCLESgP5asTZ6zO/Jsd8IhYX/j/yb/6Zz
rD6MSoqct3Q4cIbj0B2YER6JFq0Ewr/EmHk0y8tmgQ9ToqYAAYfp+TAm5PXhxVn2
1YO2RR9bFG9uDcqAz4B2y11+RwGwt2oC4b2naCCut2JMOLvocad7dyCqP0mXBcrF
jinJzy3tjfSdKxvLcr3oDsqPUiy1JxtEas5qyfEqPCGqPl/Bs6EVBeORRa8V/Xs4
P+ItjnO8Rd3ZzvGU7HgV900DyKJqbwNwsaR9OU/gweoqi5B+75gNDjVtR+T3aQQ3
NkMatZbrtqoOn0HzSvWH1bPauadqK8FUSAKnfzkvgyxYn7CYLBScLxAnibL2qGaU
CPhF3F4LgiKdL5IVqxBCgrdPguNtzMqgp/t9GwTeact+OZbrwsqXZ1yRTYP275bi
YJsbsPvR6Hay7cy9XEyAa40/MKYRsnyl4LxmGj2+usZLmIIujdRYMi9bwls4cYBx
v8jmI01qZRJqY/CVJoJkdrSSkPWhQzcJqKYpZo3WJrqAoUf/vYwlPhA9HDjzMynQ
uoruEVfqnjuRzwlT62nbVw==
`protect END_PROTECTED
