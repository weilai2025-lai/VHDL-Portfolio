`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mU5NXOW9sDLZlgG/bmaEQhzAf0ugBND11/pMkrVQKRIpfs8188kTowgkBREkOd1N
16itdBVYimGmHn0jyU8cA+uDudany3GoSWd1sIjqW349iyn3FSbC/GOV2ReNRU87
Spq9+nLxhAPEUXukvVRdGxE8wDgQsDAQW6jT9s/hrz9Q2aNFS27OmcNJyJPCFuZ9
Q6I18ZTtNAXM5WzGN5elIuDOQTotxvNL8+tlRQFyZREH5PvgB4I/T4d5C1XJ3t91
huYMRUQCnKZO+MFeXCOzpbPLpb2WTAJIj46YXokCtQKI+TaDUVkIJILCD1MY8FFU
9CgHMm8S7l0jmfhSW6bJcgxKUmO9ANJsXu0+t940KEpyrgsD5xOAiSh2DCYF58Gx
K45RJShccYqRuuRrH6LVuN4+wbtyRzEoIBFe5721EMT2yCDRg2i34yUXPMOPACNq
D46qlIODDjZX95ynZtTc3bqyhEuwWU6433aP3aaEvYyevlOdeBpTObgUXR9q/wO0
9rKcl+Pa60JFI7iJVc8Rq7ho78SansLNlGhNWlRIWhPRecyUJoadQRjfgw3vyUcD
PIDQdGBsGdj1P3KyTg3EcEcJjf3Xpk043e3HV0CCM9mZfVqtPLDnnhJd0ALsXW42
f6mKDNGV2dWE+I2yeBihRzZiaI//OG9ZGzy/xgUM2MG6WFqO5uC/7ZisSEoUIGgq
59O9O1razsH/bZBnx1e4FuSCD3NN7lYyEyH1WygVH7aRD3jQdkxSbKxFOO5R6u3n
4LJFzIw0tzEu929MAJGT0IQz5K3FKYtOaT+TcukVkd9gBq8Cxs0Zyve/VtYSxnOD
I0JEmTh5wmoELcmo5MwsRbGWfDQemDP+IvvYclftQt6M2wvC7UPkViTUSxM/I0Wb
E5V5piATCvJuQrErwH6tH2Fl1X9F+sgMXU2yKKJO2LDUx2O0lPopkSLv+mXGfWub
0irf1PuKMH7AF0Cf5ZcmoAvZ6aLouKI5HdmbGlIjQvlektNxRFvH17JiheUbLGGh
gpyZaKNn7V390vDMwjMx1IMT5hRYkSq96+t7s1T2Sy07o1993wW1U4YqTTwJBIFS
Yxsgc6eiEF1uDwA6POcs+ijJNts8sGtl6VNaPROyYGLh/FlUCk1Fnr2xXpKgYHRL
rX7gDJ8ZlYhBpu2jQv91CEgQQXpujbaRfJfCAVm5XA1avNwOiR/Y/P1w9zAO1ZsW
ebFtSnCBfZmCT0OlqsrlK6l25h5KRY+ltrc/tnlRNbpRwJMHvUz9lQstwFAnVraP
1GYWDsS9suoGWLj1j0xJ6CHujdBl4wiCNz50vl4WcxMUzsGYzhqMnn+wZFRlGVhl
fL5BUKIPJmRz7LC4QZ9bTOMnGAudIkizkuyOFM5guqPobjOFdVmTfRJTwHpdZ69h
SlTIuOfLmZ3B8WTTFi9cH0fzXRcTgxUkYSlvjIYrfupUVPU2YVb6mO1WMjNaSuB4
OR+dM11g7cObiIAQMqAFs0A7O7PSsxZzpFMlHQBUY0e/lxNjQow+gYtOpJp8M6A4
NA5/cUQOBpJTQJS7m0oxuuXCJWtpM71A9jOce3+nCldsq5hy2PYu4saXJyhB2B8Q
t8MlINBYz1s+pJrat4N9kt6FLMeOUu1IxiGXiu1p9SRoIf9X85Gnc8L99htzGg3N
iXYIyLVmqzCWuk5kO6JyQjY9ljeDRjnXLn5Pg69ATqCQhqhA+z9bcfbviwBMBQbP
PooiJ5Hw8h3KOmavxDPN9NIVEv5Q6fEk4NjwW373HcbqHQ1j0R4YTCrQ4b6TGolu
V0XLnrHKJ5EvzV4ycKqlN9ry6rM4Wgew3/LmVdKRUjAn9zKtHjkjxTFAlazAWGPs
QBr5550juD3skysvPMQW3n9k7iD69zB6eR3GP00F9MJC9Th37L6trpgAzkqe7MEa
HCuZOVBa6yBit1NrXqjZ37o9oe3FjQSoTSwt17zYYGLZjVJH2KOPMuuZKpn5k5Ft
oS4ilD12RoSGpSktdUoywYWoajhSTzGmbZnLL7ITscetjYf/bbxf1+pMxn++hItr
D99REJwd8BrpA1IZP+nXcUtRRFqQcxMOyfwdvWad6qO5Ud3o7UDeCmPSi/HN7UBn
+hEQhecLR8yNdBMKukWItPxenvyHbhYtOGcRW+VSHuH4XLpUAuPbGW+hEHIrvwFj
PmT7+n8WjTTvxuTN5QitJvp2+1hJRQZQfDGu5wlFiyvTzxcjTQW/PJ4kcnlOc25T
A8n85vT2s1apDMrTHGMk3Z6u4WFPKgCdjAxxe6ZzIIOLkjj4osIkgbagTTozWhcw
kPhmQYb+aAbA0UlwrwNlcmy5SfU4DSH+Y7Jom/w7ON3IV68OlNf+5oFlAQ5/fxXf
7tDLXlvmebs0yexDa3NTImBWTN0MpwPMeL4PpYwevgbCRpLnWPBAKGZI0nRgKDq6
xAE3vs25dQAqErkng/lojXzRSFpNmGjDa3usr4hJ2md6qS4zlR06Rmf616tScHvk
s4bdPkNtyhwXCyT9Ea3F2nGZ9EJGt5jcHBUSZtWEluiUr7+E/tEvHH+vwDdG+90h
bLKr/KvgnZIPi2n+Vq2q5KzqCaqVmOJijr2AGpTFgdJpCSKm2DExuKbKcNpk4tbG
2zSBgTF7XPwVbwoosX9+ct2EkQ+MtiuC3uQC+rYuL/hNSK141wypg4FQDavgstez
1SoBoYqotKULpMrDRo2mgt8nnDqzjWDm6g+FwTFG/jwr53ziLCA/B1JKCI6OKwjE
lZ3qOrQDkUULRld1EnsQWBUrnUSgo/pjSKFI53nioYvdrWyHqbLstzqjIW3ncOVZ
jWybv82TSDrpMsUB5TJ64vYTkBBkkjg02ZrkrYeVOgQYECw03wU2GodpOoAxt2Ka
IcTkisJoxo/djjGGGeahbitxmSDe8lNzkkmBg5/ufs8pZK8aqtOFV4DxunLiQ0VY
/jPE6U24KhB9jakWvLiVtQe1ADbXHB2YTj6YuIZUtjZ4pXh7HKy+/hqUHzsMkjTt
mqPg4ryDy4uwniRlSyvAkXDmiMfO41oSzBUn79rlLBZP4M+m15GYseBYH560Njop
LnNx3UeW4ea2yG8z6Cx09iOUP0gJbYSfqR3vIRRgI98ISGNXm6atnv5MZvl+Uxby
SaQNKRwbrQZy7BqUQBBjfxpsoKw717bOmo8GJNFYX9JHux2gxZxXFgoB+VMf2/5s
bfrEMRQblNRfbS2zL5kid2yY1RsZbRsu2O2s4D/fuktV0MtgTHJPQdg7m2KcIP68
UhqSO4WfUIWbagiLmOQMArJVLfQpYlzxwQQl1zE6WeHEj/QzoC8i0iPML9T02UUI
sriZ99ur8x5rc5MP9dX+VfmX4555RD5/3+dIDSlz3lNSyfnIvkkGo95swvIucVKG
S1BYu/nzFeir4QAwlOujamXIrXGmTO8C68DQw19WFpyKIp/ZrINZlrK3c3RINk4p
f6m5xW1RQMycWUQP2YYLGjF6YfaY7afQ33gYfFYH7xvR+egYj+ntEW71aMiW/8Hi
u2MXj1BHCYVH5dW8ZVMXvbMRrbCnXuISF9poJMG25vHJJuObXJ5oHUY/5clmd2sh
aRzMFPiNFdtCsQhTYWQGKoFljSDzGkhg32A56Oh875wv+e2QTZJXfKutfQuKvcEI
PJX3A+VGLBoSB+HOwKoBiiCd4eLBwbiV7eQTi0LI/CwX05mKLTdd1cR65VM5ejsE
iLLGjPTdEjMbwFElLKVs91jpPZe6rhy8f7MIbAN3S3etchphJbZMcQcMlZIVrPpO
QyE7ojZvoOd+I0yhksBnjzHAyYufTnYklCeA6ScHUb9jFotJk5dtih7NBCe4suy5
PxAI+TQtOn3nJrPEeqrZcg3PfI1RCAqSpHlaHiWqwfL4FJwRh6McyyyV4ztduI68
3RF90tAQxTNc2eaFdzhdq5ZoD9kRbybXMlSgILCZYUT8Hehkd1LUaziVolIUBdNa
Rk/hT8j6hdPC+foDbWwmHAmtekINalg6W2rBh2diNNtJEMGIJOZa9aVzSJT5D9rb
79aI1//Yc7arS48MrQDEPQY+mCmX/BHd2HGRCakXjNAXF4ybJX4tWFdWxDXWznGe
PCga5HZB40ZwTYtucCwwaYPsW0rzPtKLyfi9oTX9h/B9iL+JSmGIeba8JrnjSU/8
S6G2D88MM9uor4HiHbpRlxmGA9GQM5iI+KgZwK6DOqSIwmANW9zSDZiHPKBPKO3S
Bxv04u8sa1Q1YyA0eSXFQLAtnDrGp1opK2hEYW7hmqrSDCARMPFLbrZp4uhPQ1lq
a7s5DUTe8sGN7Jg1qMSB4aTNAFVZ9lVPxhW6hC+dQxM/MZdoOCZyrSde1z0Cl60i
YAY2WjBTxQzWgWuWW2FngFn3vcOQohl8E14q8V93V9jjkSoeTwwL8wqMJJay6Jkb
0EMFW2VRrNkyBOrNkaKs6Aav6+YpbqsAoxyE5PVTyDdrZhlQGZ5PZyeW3iGpSESf
2c15zZYe4fmstOZrNtiEqUM8we4HzNrwIPqVB3dUtu17KN0sXEK0Dkdl3I2tMmLR
86ggYfzmRgMKr3g/BVRb8WtcQ+6BQl08IQ6t5oexyhFixR/+giMx8Kj3PUNsHSBL
/cIj0woowcHuUPlB4BXjkmlVmpDGtTh1YepgVYyt4mRmpDcujguJK0jgdQckm8Uq
WynbEFILAUzb2f6fdqKMWiDEpHdhxrafTpyHsEOx30taeE4Phk97NebHc9awjsjF
CnyUUao/Jw13qs9Y04xf7ofJrB6q2C1nNYEVWZ+t45snTt6zZEyPBnULHFr31y0N
u6cjG/4Z4HW6X1nJsjsmKo341a1Pz6zkfTWb6qkEKKWSfiNP3XG5oxXA3ZYpgBIB
UIXq0rxz8rpUsvEZanFU3BXcRFpKo8HSIBrXTdNM1txBrFVRRCMPxTGV071ODER7
aLScCFkQEjosAR/45l0At8Ilv/dRaSO6mfhXmtVwcycZ7ONauWec+zESepAG8zID
PEIiWQ1Wa3fqfF1A1Fa1lx9/3x1RNK8Lvfmk3GnMiDlF1by54bPmy8d9nEz1TbkN
nVWyVQQIbNUEDN+4LyNxyI++AbOo6MzSvSaw4YRz22LBMg9z7h2kIYpvy2zUjqyd
dBj60Ry63CkztVmoV2HMdT1V7UpVab7kLkhWadBWJ6bRhx+uEUxmHopdVmG5bKaD
u2PxEWGwiQAaWZX/WzlbeX8ipLsw9mkF8L3yq9egFUrFo+2GcSoW6ydZmE9fW5+3
z2xNDWbi3Dj8F64U4yzTqSlqVi0exWrAiQ6aMQb13/B2Pupr6FvdGhQdPcNRypZY
j1w/thf/HTOa2DgT8YG8dw13EbjANjQUHFt5hVcz0Kizx4s2Tqfo4yQ6HyR4/vCv
rCJznkewaSd1GEhXnnJjNuwK7JH5E0m+Eyu/FuUIeSBEBYAYhIqpn+PnN1G21gq8
j/JVrXNilBH2Or/vFqQZOmQni0vur6zHjjoZu+VfEhYM4oTd2H6XIjYHrLI5pAmM
YbHU+64ys5EqDxPJO+N9xFBFYoKFkA30w1Bu05UVZ975p8bLrxMR3b6cyQkCWe19
FLGre0DRGeU6nG5OMjXslyiX1/CT7hFTg+yBb/SFQu8dXnNXYVttc41aZ1jHdQpD
r0IQ4pSK94BibOTRjOmPiN4PQcFLjf/cRaAnH39uJQJ2tISnxQO7/asdizlihDIB
1Pg/INxuxcieqbsF+kXGjDMN2ccEGSHbfzWzYEEredxaPVSS1rI1/MaRHFzgw7/E
7281v+ANsJcZiBtvAF26uLcy8mBmy44pVIyU0EOmtRjmGJaUbWzdWUUhyq5Zn/lS
wsIULDSSQvh9Od5GR3LnfSHvjjMlZkxnWPjok0V8AC8VMLgvFEjRDu7WU2HkwPE3
0BS3dBi9u5/OprbVTMP5Mj/s+9ivj/0UkBl4D1rohbt9o83hsK+J2df6l2GQSnXt
+VRlHekJGbESNSc7E/1bFd5h+amtpg/wKxggdtK47ENQ/sWpMZBl2iOJ3h0fCYNY
51BmP755+lgpsAjrLqanijrWCsbVY6P3UnCa9Zs+1HAWTWF8S40tHAn0KCyJwJcC
KQvA7tdl2h+lelJv2/Fp7VFp6/0LbXeDhZBURv19to73gkBxvMOGohIm8ZHwFez0
PW9VPAQGqGTQ6J3YObgFKpwM1rJlqpQYss7QR5LFsSS9Yp7j/BSFT7BzxCpqTmOq
E6MWljjBHhg0ncGE4GACi68Clama/n2BXiMLwmiM/QRGIiHOUKOaC1TYlqlNkgWK
T1Q1UXvQp0QLpiL49G+WN4kKHWv8qMzpUjj6xdMKkNG1GWKaWQXkZ3lRrjAQL1gy
gtpsAEHo8lJKTeweTP1vaObBuImJNb5af7wOoWTcydKnqMUVG2rZWAeUcQx6XH+l
nm+hiH7d0C/PREc71x/X6TqZ5GvT/iVSUvBlKGPDfMACXvTr6IpUNgF6Vx78DXRU
oOKxZlY1kgGSampLL56dhnGP5Ycr5mKiEnH76vAqug68j2HXkG9rPEN/3DtGDbxQ
3PvZrCSagGU5k968F1nROKD4n6LHeeX5zj4N0XWNBRMe83Lvk2erWSregF5fuAfA
Zm6Pi7dWeoFgGVGK/o4KPDSAbCWl5F04/CM9/lPzImefgy2rmhPLeoog2OVhwlGm
4TeAE7JbTyB0XDIC5R2zKoxV1isKPXGYfWMnIQM+i07pdnRwsdd46utZD3Bk33JF
26+cPDGVN1ZdqkE/DXYKrB3lulX0R8qQiCuEJqDO0PVBIesMuBfJG/dqWdUKBbnk
9znT7wkPUUF7zPafXrfp34WU1FLlYM6o88TR0bZMQtoeoy/0rSFAU6acfBVv/TC8
TEHq6Z8guThV/V7l3WzexIG2IdOqoqWodbwkca+Re1gVb9XTKskre3N5AEVXQgos
gAW22LLzAgsBX5xB6gJC5q/0cKhp9CRUE5D7liwYr6tT0J/WH6I4TzTEev6frO1J
IVThaTdTaMZyiLgxCcumgDkmN4TOpY98dfgWHCAaaHrBQNtsGfNCxvz2kLxPAMP/
hwDLON6jj3a01sddz45qGQs6+hd5Xa+ZRX9QYHu2WIX0PTjqjkA6h1FIrf0Po5BY
s4XzlzbBg722+Ie73sySYo9g/wHCARup7k4mHpUg3AYIDFasPRTkOJeS0QrBso5w
PllD1n4M6ECTvcnpkwCjO/9yNhFNA5yw8nIhFZ2SPxKLfniPHcJb8kOWjU0m/wGC
Ra/9ATihZ8TChrajn4K0elAn4j+WC2Sg0j+/9Bi3yLWPw4dLq77jNP89+Gn6p4md
JcCtIvj2gsshBfPVnFJdOOENNT+ZJ7xrRpXW9r+4UAoQrOKiM7U4jx+WIC1HYVxF
3cYyP+1yt26KHkN9aHmLgOtB+Ul9roMoni+Eukzg++Dx/ZpY3ZI4IGs42cEG1QwY
20ScFK9hox1JIg+TuKYrdp9rnFENDJPjsbVRWsXbaFuEswnRuY+9gDZzPA5X6bsZ
ICSrUyGTF3UDVhZ1TwS0COsYZ9R/yt6aNcHuXrwh0k1FNch+5Y2LTKUWV0KRGEbe
7kATeITJ/lP6WV9PzUomaCOlqnbFitB9+EL1g2+Qv0LbD9ppquDYGkTN01/G6voG
d6S3Adk79u6M9FqiCWrEwar6MwY8yibE9km0Py5V6NsixVMOGRojtDo/h6WXAosb
KAkJCLmP7QSGR/aMBezOvbEsOWaqPYR6JdHTzur0bxwKXlxO54Qv/jYhoiYO9Uno
lAgjMbxu2+Fn391N727n57iG20qA7aYeiVPzwEiNzpnHmSUNyB9LVgJGBwanK1ed
4dX/f3H4KNuNSA59ZxtuCeUlHzeN9C6RVd64/SlbNDKU3NssvZxYRwQmHTjepw1A
OZV6dvJf4b82oZx2/zVaPn3n23D4mY1u/TvYRNb+tKac2PIBYnnim7kFcUyBY5bk
b0A29zbNiqlVhGy0zTf2SK7qG9wM8deJAucAlVkRoBSKnntHqfeOaMLPzdI5z9ou
Z2XveiGqPrfMGmc5JEetum5UCoGZQb3lNgjCPmgG/u17cd5OMPHJN7ERpf7NRgsI
QTyTfe2TaXnwwNBiSH7ugTT8DOsMSqd+sDiPmhf+hlaGO4Ok1q0ZB3uMPKxfabVk
aonydI35+cBjsDiaZNX3AnUgIAwvEQhausDnqnt5sXSoyRK9crtBtOr23p7ZVYV6
3w2qgShGixUH9QAXEvXG6OI4SazRgWNG37wpaj/95B/X/VSYrwWOwHi8kDFTDFWu
oWh3gdPrYD2Z2FTJUcq1v4MNjkZPdrw5cCR+d2r259myKtLu6cbEq5i0qHyRmXm/
VG4ns2VrcLxqHCi36c5yVsvmnjCHTFO0KLw1aBFbh7w5+m/9oFSCPsUelVf4s3sY
gteQahV5zTt8zxZbA0276v7jK7a5Q4ZIKvTsrMvh2rdW0L7jF+ikPrl6KUk0HM0Q
BJ3yHnxVamREFdnp+F4mpSkWEGORdNXxy21BLBiMvekph9+SSESIfsGap1dUm6fH
UuHUHJrOBrUVyU9GagU6wUyqoKWhdMJOmbTz5meqwSfa3DEKfNukt0se4IEP5M8W
aJ3YRDakn/xn8AU/YD/EOeJOOJXMlcib0ASWurFyoeaq9xbtAgDrxABiry1peU8A
FAnLSW0EJg3ZFkIW0GJt3c5Fxf1NZiHTvPTk3rbPjQbUr5gHCEgBBT5hiqfGkBK2
V82KEC4yFsD2vCL/4CY8MhLsKDksulDxNqLxrDK1lIpaQQ6Uh7okUKle7DE3f+Xv
mg/czpOqXXtap6Iowfh86widaJuoEMwQxImF9oAJPQKMTZ1w4/zvddTQyKRQFa5z
JScMKrylGodMucBsfPU1NQhrIuib7LIoKkGquW39xUNOoZ1cXhVhoz7sx+l8BgtM
cycteIkipVN3p9kBECdtG9K8Pp6Nu6V76kQIIcbvI6rv+dyM0ibalgVFppOFiczv
Z0o23ZkSq5MFYtON9JipUR3wEkixET3X8NZSrGkKHSr40E5RYhtsgE92O5h+mvm9
YrKt39XF3zMnMNa4EaYqFdSxdi1IluxtJ7Ey3NNSPUawnri5ColDlrUfwUZJLEqa
VfYup3Be2GSV099XTC5cLHBdcjJRLqT95KondloG5h/YZJGxGezxSaEHexcrrGgd
Q4JarVh4WYUt3cYmrOY8IWw81ETJ3YFkxysihUUYYN304/ZgZiM+5FX8a6sBmQOF
7Oa6eOOYl4vK/R5SpwqniHnqUSQGrM6mUQ0erPZBochReFtA6gUoOPBVyKYqrycH
BDjCN5zgJBOufGlaj/ROyVRhPaEXumh51xi00WDNLeQrcr2Ydj/pnAbYtiGWguJf
HIPBgCMPnswZuEL3CwSGr9Uo/oE9yEmeyxVUTC2YK/S+9qjdaHxyOSjWj6ZkXqEB
tIDOT3nJnmhg31wqwrEvj37uuuhiuuvxHG5U1YHCyixuO3ctMCOr/V/sz4sdz27/
ZpvNoP0opjRh8OXnGY8jyztL9NlLRIHKQGRCOxq99A3YNWx+LyWGH0aJbUkMqocB
H2Ql1EBrI7KQw2kxWevNAo94MnG0dMIfq7tjXhCkaZrsRtzx3PYpSU2eJuC0nWsU
r/t1hSEIubXgtMkHpDWiYQHC4Y3Oxz9PjWKvehLtPtCa5hSODRnouGQRJIuiAWEH
bNywJYwJ2eTBacNvH9apGs5i8y7tbGc1MqQXdB87jABNw1zxjNF0WRFYkB8HvCSJ
ZZOjHlh4MAJGL3UXs+EbsHNA5WEV2X3N6IWg9iq+OJNo/od/RVsQE6fvPAK53Tot
SpT1zNBabzOEkakWePuAvyfz2uV16hfxV/Y7KyO9wgb/xtNZx3Bpha4YDmM+fib4
TRUlVv56Ulhpfpk8FUiUVAxThW2tYgCOXHuutULeU7LcR49LNlQHuOitV2yrqCJE
ND2AMl0Fbn9LFBtwOfusRaoLzc+4lrE/9p9Rmew3940CqTBgJZwD55m5EqOL2Ohl
id1thPsfoTZvD+NUMYXjsMrT/jfHhm53rIxekGaOfnQP77audZlF4BdwQ4AEvR7i
PzvtOtf2KLDgp1SqWOBkU933mITACIR7mVSUfI3Pl+dq2hnCIiUPCsN+Zpl1EwtA
BELtyePIMKKrdxwI/9jueNPKD/oockBGrjSHOkbBcT5CYbHliplS/kiPxN1MXeGE
F9FfTb4cOuYNO8t9pM5HWCBSMjjmriU9iQUx+rTISb1sXyo71Pv3v2zrtpbqc8wM
V/6VSHBVDZHJeoG/nnkwKQR/xd54sQzebKpKGK5/eoVQecvK5xTau7aYzOV5cqrz
/4GjjrjE5VjoQxEXM81VLDgYAOL7BpYFBbHxh4JW/Uv1hWNOR1b6QK26rOkCP/SE
+lJXVouuTIPtsoxmgLlyQLf6RlpIf3KbAVucBg4jiaVA6sCmy4pRqNo+P3NGoQ9S
IxiCjqLkTEMX+W0db/0NYGRR9by7eOfVJn7tkiCcc+PVUeZJG8Thx7CxeT8lyVWk
7DLnd8KqlQ0NqLDNGX4twXJoA/IRZcbWeb+bS1Wv9TgtfnSSrOhLle4Q3pIqYN6z
eBQnQjLGC+7bFmRf9Q91g5VLSwhEnkUGf2QkmQ4mUTroxkP/XVcYfOmvOcgy2Isu
BjCbPobSFZAw6rVvnD5WyW5J1gb7+TQlYhR+t0uqsvGTqnAxWK6W+Ihujif/upd/
6+/Pc1zYfL2UytdtyX9Zei9cmo/m/VmIHqAn0SdsipFYQjiFQoIaWAnF7HHMCpcL
o5vs83RLnZKH5fx2HE1IFvHSRqLk92AJNSChWm5f3XQdoZVbILjO3rbjbOIVODRG
oEcSBJ2sEldOZsA4OaE/vTklfP8bdxr6GMrEBjtrIcLOqeWD5BMYxQZlEx/46Rci
XQWXfoJkJ6rTvPDQh9c10X1XMqFdtv+yaN8l8duzGRWL7DMRtuz0sgmOsSSPl5Xd
gCPxegqZ6cLCItlGSihU3wMwexNHPMivZQBKk/ibtyaAMxNgZtlgzZrOeodk/NoC
LFnFItRiBipkYnhoFwRu097kqC7Y0ioApcg/eiGtJc2oQ0IavI0qGqA4AHwJe/5T
4CIic+2kcQZcTzggiYnlntsGH1U4DUQWYeD/PK1PfTWtzkkyrb4bODIXMpoje++Y
7hsvSOvwC3f7jPRcQdR8fvG/xPYgCiepfaO7UCibvr0sT+yAk91ND32O5d+I/29X
L1UxHZRMhbKm5AV5IYADuEa5joowFMq/XJLFykAiaE7RF2gxHR8Y0Jcsg9hvPrPo
EkZNd+3aU+VErsNk/NohqnrLvOl+tpVA5WBPuJy3AORnKIGFnf5sim/Jw9BCXlLH
s9+EIrMMyUhrMSHRKlItihPxr1d6jjdjplf5GTGN6A/wmZ2Yk4cWbn9rftsA3mdI
NklzeutTdkAKpH0aDyqnQkPFXw+jcs/9ReJINRj+wiPsnSOdIMwiqSt4CDi2+5Pf
g0f+hJFtH3PIdMhd+1JOj7GhX0vjnxlpnM6ff8cSN5eW26B3xhYzgea9dUvKVfIz
iTHGaRsbu5fKcgN8F6fVxrSbk1MDvn++SDsfl1clQgJj8LquTI7iaPJcoO10VLLd
ytTitJixKr2+qJYWORCaZrV1s1Z7j9uzanAQo+sSlcW68MCSOBN2rD4S/ONPxYz3
GMO0yn5zHqoEvMPgGMwCOgpOXfqzE/ntJRLg2JJNnJ72wvRJz/+6JdZj2dgmPjCJ
XkK7PJxknJeWRK5iOLMvoGlWIQ08megTRZi/z5HyckvgpXeUp37BwQ/CrnCZWpLN
IqIZ6X5UVitYOYJKkKG37D8Zc4FyK22xpqVDdMP8M9GfpVf3rJUEd+8yjxMCxTBR
umGfyPrC7yhVV4+anSg9mF5QipewsuwcK/++26fFfER47HtEoEVS4gGTf954PmSS
QE9HX8PRVyAnSHKeMLaRlSc0CkzqEVJWke+8Yr7ap0My5SOGU+C9BTughyfpHb9m
/J9iC2/dnTtCkX2eXzTwcir3twMdSb1mVl12g90N7GnqXW8WNhV/pu0RtVrNXNhF
+RGf9wIlm3LMo8JtC5E9rM/Q058bOKcW1GVObzOU9BhdPOroBoA45ZZWG+Ct16vQ
F9SngnHxsP8/EmJWkq0xcrQwgL4WsauNG18PvCfLdSh/AaEhzuZTRPqOuVSEaBiy
DJa5peXCsUfr9gda4TBOzzxR09VB8pp9AaExZ+6s3JuuGfveOqN/b7cZPVxtgvuP
YhBjAysgtEaMv1mADZagpuVw3HhyfrASCP9Qz9aOtUOfi67erSxFzSoIkpCTXkTJ
4mZ9mN05FQCbpGba04YRges6Pmi2WT67B8GzABv4i8kwnLxI4e01hV8LJfn3RSL1
XvUvFblAQt+emyPuSx4Mtd/0m2NImafDe+k0tXzeItYu9RpqRANqPvNva26vYjuQ
6w/hmtT7OXpJVpTJOLwXWaeFsRTeYXELL8Qm+mJZNbbAkrW9YWvjtkHndTol4jSs
cRc3MZnilDXLIhnf5LYOePnY9gVp7I3GGMYNw89bbyrVUXtnompkCxYOEZpOBViy
ls1APHE5caTHuKZeRRe6eIIKd0cT3ks4IA4hj04nn2yJ02r456GSU5XTPNhOCpTZ
aV4Q1j84V47yXOKQWcNuswe1VXZ288eR4z886XAfBMiVurz9v8p5S8XITTxAvu6v
NI0NGPJCGvalVup5xmw/tt7LdcMqsm1tpEB3iqYPXeutZaO+al4ow+1wD0f4jls9
T7vuyI8YB8sZvAp4/NXEJvT2qO3yRHGKbtEzwctfSrhXwCDXxEjgxu/itkbya6+a
5nOaGB1z0O6Wrb1XJuV71gE+gCYoNjOoPl0h9IdBRscLpUTIN7FhrcGhkxERY04J
THUdoe0VCAvWYqLlK4yHww6FWIKBpyGXCtJd28fZUwgnkALL16B4IKMP4wsNEZKa
PdC9D7bBwp6oC8Trswb4B65oA7mgPnLdLpoqQCwAM2Rr+pTgqD3kJtJQZUnkOwON
8aaXbbQwa8K2qXzCbODRhjYafNje8lzjV3MDWjBlzhMUfjfVM+2qPqaKtDcvN0qo
3kwxY/5OK/62Ug55difedHTdq3Ziic/sp4gRzUHmysDK1GW0p2IsH5/URHBTLyIQ
PYhuww95I+bU9yJ1ER6aytzP6R3K/1735ncomcNLK64sif8PZ05+JxZPEIb2HSjS
HNGK5evY3+RQ7U8zu/LrkdfzZHzQebvPpOmdp/Z48c4PGsFjZaC0wLMQt797dXJ3
h35WOH6zO6Of7BFAZAu75tleY1n25v9Z1SpmrKip3uPkTmOfPCXll490MMXJEbZE
puq8OE7p97wVJ34DIUdo2py/8u/dS7Mhars1RgWzGNlPiR1W4mX8JaaU5486V86L
AqHq2BOVhU4YihH0ki4NWhvs/7pYNbvewHB6AenbtnydHCrPSr5MhVzjlKvLOgc5
WCLk4L+dC3x1/LWkhmupEc8I66vzA6+kga9nKpVXar/4RVP4N6ptJ40d3IpyoFyj
odfLjUmBR6w0WKTzoLqReeJIckGXiMNJkehNiwYgXYSv3Bg3wbLlyD288F2znegW
NhlzFHfNXiNGWRJoALMWALc4NGHh0SADbneWKNdqYOnUx2nvoro1ZizMGEd0ZLLy
gYjhr04+EhmBCOvCxAulzSbqXAwNrD7+jkzuLpIaKESFpoo5RFCZJmy0OI8g1ANn
J1ayCSSuNg9HbmJ+N86wLcHfxDMLK5wd7RoKe6gj/S5YARP0toWbLw9uUMfeq/8s
6lELFEuDAP2rOjP1AWCzFGKuulE71rMAHksoYu92iZqhRh12BSz3yxmLEjKQYfXQ
mGFyiHyhQ+qqMeT/+ZsKAYsdtWJ+w2q7QMe03L1iY+KoA24/xTBo3xD18j8SqkgZ
uHt3Km3hskEXidn12KPH9D+UOb4zBdDDL1ADmB1nrDhhaDgTsjZO8hL7Mmt+9ykl
DrI+su/waYfzj302EWnQChV9Rt2qmotoV7o1eZc+gjpF7QPPA4/Vj3F6u4PplZlG
3IBX/YqWxat3hvOrDwX9lkwfIbAwziYf1YCm9k/l6zi088Yn3oSXf3eajdivSlKF
HtHcJ3lFPo0lHmA/bYCZstbnx2hUpYmPScVpe70Z7CdAHvwIHXTrAB3XrFFsiEY7
5lSla6vtdoh71ffRqsG3BAnCWtbyHtxwooedc8Gd85mpbNujSm2Q6L+skTDeHxtf
swXGJ313oWdX8M1c02E33UdFPMyC+RqfG2lZEKlH98f5YHg0tiVkD0AHGGJ+sRBI
5UKq+g1zunRI6kdnKGkDQ6gSP4/uw2ObZy1MFK61Cf86faYeshufiMYzFf2s/hPg
UzSdk746nu5iV3Gdb8BC2DAH9l8FiVk6gl+sVEf3Eay6+LbMy2kgtejFQ9L2rwmj
ctT0sgzcvAAxSafjIUf2M1iWEfJMIl2KGIqYd5dxgNBJzASc8wg4DNplaXDAZXZI
pZCdwXrBH9QMIgI9Zf6NGlNpabcPF0CFrVsBHg6pKW57SBqnoZF0XKYhBzkQ4U45
hoLc2SMxJ665OgW8Zddo2aqey8yjdPhQxMSPsYuOMwq3sKmiZHdiy6zmb++t5mGm
W0anWOVFZjrYaaJJCMnAsS9MwsydosWnuokXoqIixiOQGaFsOh9AOuEEVg4jS5xw
AQPWysFQiHeFpIZLpytBGK1uHPg6Ks2iW70ZvQUlyYt57dAmMgAjDz/9t+lI+FII
mOXsvEAj520TXTZDieiIMw/5qwVeSeTQI3U2Eg2K+0+/1T/77zclrcMFfvBg4cRP
yvY8Rc4cNUsm/LiDwY0Xp9Ceh7Uw1ddFdAb2roBZQVpTgCooSVyKgJaLAixIiRka
aL8u3gX//FbtPxBWNu4Yya8TFHj9zV11fMDxrNPVkZ+fKGxwSoJC29lZz1djAR0I
QKms1JijNPK6yGIup0sFtfKWwh5+ZAe4alIaIfftZNgVpySoPXXMoRqL5AmOL8l+
g0/Hw23ps0PC7osrLAcws86Ti4h8a9+NGeQXEpPv6sGcm2DtcXrBjQJdHl1ZCPLG
WWhrrlq9kAOiZ95thfDGYTXy860Gf5mOE7y6zsemNLCm4xBt8OhMCZIecTLxjqxU
Iq5RBbCvcE7o6VkQyeW1fekC6EC+5jR/aEJJi+1vGStEoaNQ27tQC6FgBuvdZpib
NX/BUVwHQMP9CXbkeqKCoABPzLXagmwC2UX0UaMgg39MTmCAoTKIAMzNSz3Ugr7w
wReSZr5kvy8wZnx56GJuNefkDyo6ZMZwb4NPg4ryBeG2KqTXBoSWYRjbjFBkcwcA
tfkF1BHlr9mbKRfzjJKet1FCbXqE4JuI+cdnB0Sc5Wz3JhejRp25ZOoUPGi7U+th
zPwYNsdhEQlbajdBOzWC9+/bQUIZyD+25jx+2DG7fcmj3CxzSQ7uv+ZR/rmTJMJb
da7EtFLpvXjhCq/Xy/dHpD934e7mRSrz0Cec8srII7IfMBZVOG87q4rpawUeH7kC
tvRFXaMf2nVycpn4KmrHqh6j7zNVHedtTKSoYE7KfEZcoNxIdIrDg5N3LrKlaZao
5GSxdo9Qif987IiwS0qGgd359zaBQqy8qIpk5kquYKYnKly33qcLwUh+mDYfepc+
K1YBCIqWYgjlkEPM9mKDddhOJR1M447z1XYSHaGWlMypGtIkJbFRfYNzwdWuIwuS
qscvyTcadEtMG5ysP0cNd4ApSvmXvvz5YHXCGVS3pZZE3sS0gM8IwslEwxuyC/+m
k7tLk6P0kx5fYCjOuuXSdZ/i0GfZOWqvpNfHGbpI4NW3gRCEe+iHCJjhkaq0qwyE
jhmNaZbwHoJa4+fFboXR8AGneZfSbk9p37Qped0TGP84dbMHQau4tghU1Y1Von5H
G2cDMBo5CKEEo1BAlCeCnFHnE7c5UTnggFWx3xMRqTKVQtJ1F14HXaDX2Slmmf2r
janUF9dqGk78LtyOLBeHrchhHjPTzBDZFTAYGwnaBUfaz7zvb8k3LHw6S4lQfJkJ
zeHQCXkJZ9QQKnu6mKl+VEod0ZrZTv91XKH7uOICSHjVBtFNOjkI9jfvzJvAdTy/
g5YunvXBjKyyjX6G7pjD+64p14BKo21En+AeeTcjYvt+LhHUyCm/G0dGr9E4dQ5+
dQZWNwp9JkDpUdKmsQU6Gri0JVJcX6+Z/hoTlI6Lwpse+bF9ss5o8KGCrI9Hc6oK
4HbkkOBBbg5oWdk27cZONmm6jqxfFPjmkMTvfwyVMtEQENOF6x4Ys8DdukViMTvC
xTDQkMyox2G2op0XwC+it9Wtnr+OjzE7Vj7RP3JopWuynahgLIE0Kvqhsusw7EIz
8QKqQMBWljZRCK2F+S1UthaeHp3Hqiaq5Xu/0NNPECPafDWgJ+xeMmyAvpLnxBk4
hoZjM3N9pKSpq3KINJyeVxVLzODFuGuzNOOoYYWWLHEXADZbDbSB7PaBEE8ozeS1
4XUIYkQKwa6HCtBnfHlYlprtu0o6Nu2ZPCCap9Ug4i4flTZlvOPopz9Uc7rVwQhr
vCkOQxe3xmQcZabrS3C4PdSvW6FynYUsLaCcHybV+6BvCyqpV0AgzE+V9QZVrdhq
dBTtqAwzxK3SSfISY9227Gvlzv869X3flb9sU7js1QEG/ELwxNdmlcKRXVlU3whd
TEmz1zkE+ZJwZqxTVJCtHRhiktxJotC02OEA3lIjmh5xNjTex1pckUYFaBOskQ0w
s4bKqiTgXUZfwFGqy1csL+xat2T8C2C4n22Zw8VquRDn2dwsEkwxY0bqTnv09vxg
KhZnvuQqMDhXkTNk5SzNnnHxgL4/6FhvwMosyt9Y624+vmQENjXV8zj1qvZK9cia
/JbaksrN615Q8CDN1WLO5uhijK/ARuaQdpSsHhgqtG5qpf3Lyd91CCDn/EixCJmJ
y6hPJEHjMfuj0l04/bYpQNwCQzsw0Zkcqm3xRIuzwxPG2z4mHOdELfBXvzaLpzdr
PiR+Vy5HZVHXoIOApkEZmQYG5hT7OW09sat3dECyZIDHv9t1aVtb8hDeVidcGfCD
sZ/egHzOG9KLeDEIvtnwdbROOGyxYXm0NzFoM60wfOcoIicQozsjkh4fUhLynyl6
lRdYJYFon6eaCh5Y+TPLbfGz7LW+sfqU1dNadklb+Sl75Bt4VoDcO6pvhk64AZ9A
FL5mBbA+majQ3qTA3HwmPqOJEVLz2YEob9jxd+wJ3ku4CvHQyg7kX4jIgsGJLA5g
X8h8Cpym5aF1TS75APSX8a/y7QUL2alC84DITvLHHDs34wZTIMJw+jlSLItWfktT
OBRxqjp3eU5s4XXpn9Y6x+shMy67tPVUG9QIByNDHat4SbKqGMfKPftdU8CqLlNT
PJR0rWhtGi46lvpQp1kR5jCSfOlC3sB9ddtvBQ9hP4Axt4Xc07r/cK2yQF1/elv+
yGo0janbQZTUW9pNFGOSnBPjIXciQ05Argpcns9wDVKu5P6zj27TXNYjnRyBnc60
t9shixqlb176XvSzAsU8cSdj70HFDFTfa3D23rneJVigk03Pwtn3U0tvDkWXu7Qc
FRBYDIAKD5hK/0FhKQaNWtPL25Qm1Yyfi26LQQe2t/NetbWSNjHtPWSBmbHCK9X7
KHKOJOJOjjs7kXC7oXH016D1E/6mkcc6c5Qxr8JsiRmeL6U5ZflR/or9uvm7HhwJ
PR0EXk396igbgT3EN0nAqUPvbQI2iigtsWFwCGt9OYqmkVvVCwbhOxwK5L/ROL9S
kohNZZ4NYiVij7YImXGp/F8BurcaEwUpKXyVypEEkRU0nTSaoodVuozG07zGOWhk
/lpfxM7dILPJjpFA1WReSbYCjZotFHhV7qOTPWuEY67AUow/ViIeD3eEK3La32Cw
IRdxdaS8Mdg+d9GAvqBkoprXHO7bXnOpRZI/9A1tTO5NrK3CDMf13NKupfp1UBuR
lQmftVzu4Mtmu2IdxslsIdrwZ0z5vthTdHvU7RN64ZJY4nJ7Pwj0Jr/k8+gaYphv
LwcUAZ/q/OIJzoxeT+Wn105ktbpQxqIteAQoFSVSVP300ajLQk+qEismsEEi0dMg
p5dMCWIjASuQXY3FWLayM4Y61nOqFwqSU4iFyi/mpCRF5w3HN34uB5R1Jx1kK1aW
f1Kor5BtQ43df3RzGv7+LhJsLtGUYLWWSogIje8LmgbIteIWC4dhusI2o1kyLLTn
AU9/+Ny+TeGC2IXS21LNRxLeHQMNMgWGRzn9S2oDKekS6AHvnRm8EFTdZWqa6Xn5
8Jn0XsoMaf5OezkX49WJnd6NoWau2N3dtAt7rVEBuyZxNKcWeSGZvsUc347s2uu2
9fYGWKE/gtsBbCikfCCd0sa7HWktev789+ZuTaQM3QbDWOY0Cx0RkPkge4nxDfXO
FLRhGg1MwqLyMznyeqhNMTiGqbl0A1CThng5pzlPHq/+HwQwEeZIRT7AkR7kU932
FQ+Au/AKJYSR5NtVRnQ1669WuVqVKQiqOfKb2Laac6pNOeVQqImcEbcpK9Jm6kNc
ZzE1Krs9GAy2d/su0+gnp3kOiwzZx62wRLn8XEkqCB8DbMZKJprBSJtm2b/CAfWV
RAvOxNxor68BD98QZcOUR49disxaJBkScnvgGWhAqMFZW/H4ZbWaKZ501S47zUtv
OCz+KEAdsZBIoVMKaw/oza2H7Q4QXc2LoDZxshZ6Tf/Xl+d0THbET41x9v6yY0j/
Od/GXePIMqSEx2C+BKhnk2o8NjbRiR+Jq443E+KL8NLop+x0PsH/bIuQ136aLyXy
VqB7KX6n/wNg+B1PzwRaXtwtOsNXtnmvVGHngSzV9hBWd29TGLuL2qlhrLtcL/+F
/3UW3XvnZtbMRNpD8FY7qTakAbC3Pn22eAIzoXCEMWn3HuktN+ERfShpp5UEyb5K
1tddRVhInyIqmhIzMrS0M4MnpweLS1zx+ppwFMrrCKiJs+2QodeFJ5mj8kuBGalv
uB5J5Avx5sTVrfoId3eR+ELhbtfOW/5QSYMFk3dofQxv1VOp8vj0Y1KPZlaoX8T2
UfamFiuQ+mfVBZQgXpnM8ktIM7t334gmkAyyuJBo1g3MYFsS3qj4nCFCtu+C+tB6
Dpye9YS652ZO6CCoOqVPbFwn1vUt0wyEPmRMYw6XqbuizD6uQmDRMdaQ9FTSnKJ6
MkjEVYsG9guTOyy9WZ8XVev6wE3J6383Ba85wdW0ihCH9F9fz2jYJxtGFVH61twS
x/sxmIk8cYQcU3rK4h5KvJag1tSv36tVrvjvX0JE3EoK3QpdLkR8VxBkdBMEFZ9W
iCZSQTTwRm6wzC+8ft7xkVNHWNbdEsr8JD5fSS7SUfIw9htouUFiN/5kQogHJYJL
kqEO56aGh1Vv6kN+judbqXQBsJL2YptLg6+yCtjY/98dfY42eKY5LyNVwl3BPUs6
voCliU5sCP3ZMPT2JeNBAzMJuryKHUWucJc2FLH0sFOYVM4aoIgDNoCLPMqn4ja1
9Dds4EEY4Hp6GOWakCOYT6N9O6Bp28EniKi2RE3rk8GjZHE6e4t9bptnNR+bP1Eu
xMkI2l8GzqwLoIktev37J2cQqCvH69GkZiaBAtB6pexreZdGyI0l1zTzcxau7ROJ
vu7bvo9x8vhsJ0mRCSNB1KJcL3AT7xB8w7+3FRIagjXJTX+n5XDvWKRvuapzPeO3
Ju71dwdRC9uTo0+TBM3ebOXi/J67iezUhvcUY9UJIvjHwzxHq0JdxWfes37LaDgs
3u1IVHWlARcwMu0C+9kMbKOd3oIB1ImT7okHvag7vnbkAehWsy/uNsxFGfDBbqPJ
ykPIE/996nHvUeoiSSmovqDcTgZSY3z+4UZyJr1UqyAut0aFSCFyHPtZ4rIXhPBn
CSaGH9IRQaMCORpxa5+2TPjG5FEPtzu0vmt9h/XC6Gqq/Efkj8Afk6g08GD+EjW+
tb4AmZlmbz5cB4AV2NiDbjr9RAlTcUPBn9QQSqVUeQOjQCvHPqAOEy7oCa0t/O6d
PNEUpvl5xCeDO28nT53nKrOCm5x6RLhSZXzb4DukkIfMO7Bq+NNKjE2Cp6J9e9IX
zwVZU3EHgTprnrCut2lYzeOhaX8ThPj4KwANE5+M0N5yMHgWmFyyPDFTqEC9wYfd
qhpfpc1jxKJRCsF5ssjyQRd+uRGoodztg2ZILou3qXvloYpO5UDkd1lJ+CDvx3KS
oOi3Qu0NiUKUX7rg5fPe1UtArv9VMnPBxNGPDHkxjLYIIYHNROkhMZjBywnVUinY
i0xihuxl5mnEFcxPZEvghBQUbdNXM3R19iz7DpN83NLheeeLW5DRYfzGkg7NsWFT
EuPuGUH5WzHCRs8aKuXIpiAGrGU7H2iJsqlend61ERMIQmsPKOcTPSCUZCmuPy21
2aDLjYJsLfllkx8VldJm1ThSFS/lxfp7RjyDAK03BpBurMXUtthtPxmigC40sDjw
nXqR1pyO9nICT1e0EKCTVU44juLb39aFz/efZDsktG4vRIACi6dzKWJmT1vkqTsn
XxbIXyptgGBdUAsZDT2NrB294+XA3mKGfw21HTXMfmZUxl5ePz1fj2le80rKheUb
lpRFGHK/3wnV8AtqOgeB/aWSb7CfnCgU26U1PZ9wdToYGsiiXnmpIKTV2zaHoyAU
mC5l4Y4Mrbty1eYCdh1GOXPM/wYX8QdQ2HQkhN9t6KQRDHFXFtubx8fXnjHYj+JO
JZZKwzgaX7Wp06cQqXwmzUjgx4GvK1f8BfnOMLkYiZSW6ZYiONVR3nrcj1szKX7u
Ov2WMb8odhR+legM2kg2/s31Kyz9ME5LMgKf92+SodAVmsWfiI5J7TYwj370wAwo
u9i4An5d+QPr8b6/gVcydaNTAnmUs4K4ZKv+XiJAbtqRZ8WSYFMsrR9R7/l4IDwb
/ig25Tv7wyGepuga5obpVV3uxBocVN1DGQ16kPYibBApVGx5BUcxV4JtEvFLQNse
WcmK6PzAEX1QOrGFj6GfOrpn6MNFYHBZFGt4HzIOmqqW6x2KsRvCJckiD/k6fncq
cjE0KNifJOmvnyqhhhGVapGRhMKxqSqGEzgENcMSN28HT6ynGcFm5eODb5QdPn+S
zjW9e/PcU6e4Ffy9SIGp5J3C21ULB93thOhZRZQJiDeFbkWM2aYkanNxDAu+9pNN
SoELJAVAiFb10c+rG63GlayhEsNygeA2SSta192ZY0JEd/3Hix9sEolWYt+f3T2z
jJXdM2UxJEToj4SqtpTPCAfDMJNyjq/I7Lp/mPDFuSVsmycI2UXgTikR9BlZmbIR
dCUCfYLyLmSlmKgBMEUyX4AkHcVTOiWlk5HcOnzcrt//qdE+yhpon3oRKIFM4B64
sDpmKp5cp5pTJH/tIgyHBCrpNrQ5UwfZ4wUDqPJc4WwbZZPULl5diGNCnRe8IAdL
mLONml7pKLUm4lq1xl1owtKKhDT378QnWulMno7DmWzISPFQNlM6K11vn7PS0DN7
EiEzgvPSQl/g7M2zxJ3j69iImhNr8D3roAi6GwjgPekkbU4zsYlLrMG6do90w7Jr
h5G3QxnOh3HEr8NY+9FQZ/xvdyK12j8CEi9TUkpW1L1gItPFmQPnonqZJzdt4+iD
019Oe9lQ8cGIj5i7HXhEw4qvFwbSHiG9KpmIg9UK/3Zg34i3BSPcxGDgiFwZ/tp9
ad5uSQqbhbD3zmAfZEcpaRnut/j+wQ7+iAbQIex+psF1aCXSadhNlD3X3NKATQyF
R9GHlKGs9R7wS10lRzFsG/EMNt3CKvcbANYgcPppbniJmhkzRFHgdcEgiiMhmdAL
Tu3C9Yhjh4izPRLf3InO34OCPLoDAT8kUmkdDfq+92NbeFzVcAcxyxOSReriXPYy
AItX9IRWqX6/IktBtVyDT/AdFHsjUd/MiF/YUKJlV0Ftk1KKA39joYn0jydp7PHy
hZFDyaWBBscyjbFjJ9iHlf0cnSpA4UmIUhF2fK9gBaMoLV6yx4n5eZY46wnXamqN
pMRfwv1RUjpledZvy+G9k4A+2jRPnUKpqe0GT7hUuodvlby71x5gPgIvtF4tiYUI
FZprA3bqsRqC4RWBT4W9Ip0bYLZCz2MqY7oo8tsgaxlsxrbFlsm3vwr2a+Yivchd
m8R7cbftWIaeJlJ9GZKmTYJJiH0LtldCYnyDEs5RnPAnvXQNXXIBvNhrbZyexL/5
cQeBn6c/d7xzcY4IOr631IPj0tnGe1Rus2MuAqcR8+1TMZ5gdtfFfXVp3qNl1AKP
1+YCIYCkh4feW2iW7hSSmauIFacttdjsFarOtlB2D5mjc/Lo21JSu7TyGhyAR/6V
jWkwl6+5ekZuGwXUZUAZi5Ui6PizNF2M92d35ZnYiLbbCNNNeZdQrrIpywI0OWJR
k9UasiKEC/oyeNrBfdALNyBzobe1kD+oa1blXO3v+BntLB0LOLYyGKb1EqMSiLuT
S7wMXPlUoVAauiTxvkbcJGpGn1QFldi5lCRIZE8rM7Le53BFWXiWzdpLrFzQRsBb
ubeSi9LMdn53La3R3W29fzDaK6SSkyWEsASfNSffXq/N964vdb9xbvtVi3Bb1ceQ
x53nJNNrF2IC/YTkNIffN3HQbAvWHvk/L8paVw+RRbH9DuNN+LlGN5T+gniZxRzK
AzQ1rwS51SS4HzjuQI2yNJrmGyRGGA8N5VOcJc7X2KKZKY5DYOJW9k7E1jDM5Mzo
ZsO+gQPYkmyi/+GvQbBrtbFu8+Rn/emyL6Adn0kueXlDJZEcYc3x1AFN6LAMBi5g
LT9FxxMUzd+x2rZO6u4j0qMW/DGtyfVTELnLeNfx5tAN4H/IScNYr2BqE89oawpZ
C6RU+vw8b1u9tQ+1lNVSNtEvJm2zQSOHojLcbZzpQq7/5oH+erosGpP1YOLoeWhh
xX4ExxMdbyHnuBmQWo5FHtBYH3igfA0EjID/KuNAfrVbvHdi0DFxOeIXryJEg2JT
OZu1wYv4zOiHbpY3vfrvkXKdfmfCUQ0q6cSZCGOiRgm7m1E0nZnB3GQV+fAd/3gb
68XhJr8vKnYSK+MP84Ia3OopYMREtHsVKuWRr2ZZSoH3qhS6lF7nCefHjIEYP5Y5
EloydvFanNiisMzd/MWNsP7gwekTv0gTnvw06seuXJLkORG1prqLNCc/yIsbrZO6
/QiUudw24g5EO+mE1ciOHBgSc3wCrHfdJ9w/5SiXYrP/wKO+p4ZQqstDdZNYpYaF
xQWtTHAtuEVuvTrZmnx5EOZwZ6UbUrvM9xn1JtDeMOEbCuNJk+t0oaC8864W1OP+
P7rDUgWD6TXqDoMokC7gjxt/f42GeE6KuBqAevcvFSRScAFasOWhT2FmLfEkjAqo
WGJFQY+M7tigtV1kYtr3o33wF6nbfDsA+AEW+qbt1LSgaFZ5KxYkxBwjw9CNywa8
nD/mCMyu0AJEmtBW/b/kkitmebrvAH0dbCPA8IDtLiG6T8KtRupJ1zFP2VxVScDU
MdN9ZRjl47oMtKAQlULC5qypjAaA+zHjHjAKTCtZQtluDSyhpmoihFbCHIx2cC9b
SDkV+UKhucQG45dw5UP8UkYt/OBX55NENi/rQZI4ggtaLO2S/XB3oNF4af3YPqTD
KHeOdxNIz1yn/mrMIdEiVT6f5R8UKVZaEt2wIpD1bLnwv3Z15mlVASnsZLHiD3Cp
8xN3d3wucmpcCXLPMk2A07Jll6minNemRRzn40TCfdEayr0YkKZwbVO312LBgpnw
9auk8akJfbxHW1nraPkgUvxfJBkKm4hN1ELe6p88k03SFKRXPCnSIQmptfQjQbPD
FQLVeFtTYjATUfZrdKS9BFAG+a8rzXHhb4uWkFk2ZizAbZ7mgZlkDUSYMT+0ZKFH
nRriw29Zs25CscsxMpnIyzZlOx9I6R9lpd/EZleEOene7ufrq3NOW1hBD1/Uls/B
5QEbYT6QdyjXqBlda0Rwc673021Mst+P/6hDhm/NaGdatnwyNhHMgfzc+h7mMzCg
rkLGXQQ8vhFWHf368JhtcWhh2m3jKCuE+VK0XMn5GRGxKvo88vTjoCxXG026Yq2E
6YA4HBxPFYty6k76bCiGYN25XOv/mpawJRbnobNa+KmTIwfnPigMI3wcxYYW3GXg
f2mMdi3cn5So482u0pSdyzTuic/Fo7SPkQ+6/n3cImKKmDD09dTFzeOFleFQ3vDD
YC7dKo3xmEDWnoRueFLoJto7ZAzCaityJU6+gTvfmdwcTwCi9eN/esX0ZD8Eqt8e
AdI0iPrgq0NVOexTj29NXf6GNqZQjGYi7LY3Fzc76GVhX4MfOMxGKerLvEsOX7ys
/ONjGOoeEaxr0VHUN/XGRz131REylebzyQn8oljJM2Jh6yoESelnJ1XWmNY9cMPJ
1nBhdD3YBFlY1mUL//yfvEGd3UUDupUPIg00HxCSdAzeYpcXST7mm7oHz+F9uT89
kOfl0uWhpRHfMfRSEROHLHHTB9ERMTbQGpqopo5NoeiqEw8WtBH5gfQ/Lkdb/Q9S
pn8xSMOqr/LrMYyvSfNNKs1JwHUQmtX5sfXBThz1EuSZAlTIJQJyFuToinjaSbOH
pIk9ttoiwSK6BIL8ZcoesV3agSNS7uz7osIYwCHsH6M4UH6LfqC657wHigPutU1y
XUOP6wgY9sDCHnLqxOk4OV55JoJJE1jEF2WcHC9GSIX+ObHunDRPqJahN8+vtb6L
6eYk9DmEErNl9oMTfW65OUp+vKUKGpxCZ6yIrRwPRFkccK7qfYnbSHeOp+nPwv9A
33u6gC3FHSz80ARIG2Fph/5eY/lALhi34OLLV1YFwHgznAkRIwyV/kh5/NkzRqTI
0LL0t/SSjg0k5UdIrgXMolY1HaaAXOh96XHDk8f2PdZAtqciNtMkE3xRgiVHmWUf
cC9GoapuJ2IzVh0LP2oNZtaeZDuVv3GGe6XGAsS1Qkze7Q9Z/YRdKbtagyCIj+8P
JeBovT7C+q9xPoJcKprfmjvLXjAacHBE0GS1Y2EXYem/sHR/RKliAHOGflN4puZp
vr2Jt89kpWK5AN4YQaW7Whm8ciphahMWH46C4paz3RU6FF+lCQ2PvhT4aRprLK/k
4vG/EwkFe5cnFOWKXIWXn01NwnkEo6Oae7oYF/w/fAaxFFsrH9E1ObQxZiytRUfc
CGG5TIYUMiLmwRZcgZ9W1o/GBC6dmsd11ordDk1094hwwASeuJNMQ4sp0nWz5/F6
G9pm9VrBFkjIHtIx6IRcW+uM4vjDpS5M1y8mVd9hIUFKVvZKzjhuBo8qvc204bvE
JzEsMBTkgY9T63omtLpZVzrYpP04Tc0R86tgSg8lAIMamGpPWxN62o11xlYvNSaY
vA7+nkEIfZdrjK74GfAhCktyyFVtMAVWTbQwAnssUSOXqvPojaCxHZMwjexDdA8n
gBLDcmWd+BhtPhyb6eIsiYer0l+UxXqf3hMIHeF3RV9S+/LN2EfKUMtcy4JZzppQ
rq6AiVPimkrdBGmLPNE1KIp3pQxQU7MndRW8XbOFM8W1t/Zq0Sq94l+D7nhi+JnR
WOSlM1nOoXv5bjGrOrxQ60ykH30dwGAnTEFouYJwP4aBteswt0ZFHK4xyOQoLICt
KusRTiih4rfqzf2UwqhI2A3SZcO+NQ4uCkn83LXUVT+R2gQBpCf2KwtRuLsu/7qI
pLeejka7YrAzpu3SAkyUiRMn1LsuIIhNQNhmaHV3FFmAOAFlCKqp+jRBRTu4rTpb
X2zlguf2Hs2syIQlL5B/LZu2xDklYRa0QmGQq05KHl/cKPoNg1YZxMMfn+KvG4ze
S2DmktwMupec1QL8sRkN0RXPu/jb2Bb0MVRPv74FdzhBQTiuNnK7X6dmI7fU33SF
wWX45sYWUvvH88NYO3USPmX7GeR/oh9+yym1UMGeLmZh3KI72t5O6kC69LlDuyn0
o6NOJLoo4Yu1V220iUTkqFcow4OcMi1dKqOAyHRpEM2IZ8mOjtD4gQr9vARJos87
VXnqrclajXoE8o9BuvhQzLC5Jk4fu8i8dZoL81dhWQtdDnBEgNXM86hsCSweu90G
ykZUMGnHMBOaBlx3kSNAhDtOPn6OvhW0i2Sf+PHkg9EopCxYg21fBpbj9L8n74Eo
tvNiPktm0bKuJoAXWGvnLRYZb5ub2rKTcZ3756Wh3DSSc0aZybUqsCkOo6Nf6jaA
dTgPTHr9FptkZ1r53YSCxNBZS6GqARhXP7L8UWBRp1ewsY8vMmEJ6bk++Ih5+ecH
40oi1VbB/T6ijE9hQDWGLelKrgNaYU2eCoJ6OJs//Mi5Gn5JS0V22Onu5Bn31aXk
EOQSFGXa9lPM6XBlG3Ma31d4PEbyvp/yvIQnNvXNmavJnUXzwmSqcLmHLEMK5C2l
/5FdL4keRAVAKenVHE61X/z/aPQGOzjvKyKt7AL/AIk0flP9XygILFcxlhWkIOQY
41BJ0avlRyp4BJ9d1Q9ecGOzUgtSyu8mij8KQEzBExoVeKczhZnRHs+DqoA4QQw9
dF4lbxaI9kEQqc/UNXPx7xhab1xq4x3iKstIcWUjOa+/3FidbyCifyQLMurO/flS
GxnE6Vwp4OTVJO/8Vn6juS3MqVCnFrBDmgQgdLUSqvKJILxUQZN6wRnQd2S4V8Z0
amtwZ/KGxAaTfrkYJIt6KtroZA3hoBVVr1LulZKLVx88izxYGZsID6B9iwtN5eY8
aJbgZMIfBa23az3xSCNR4u4egfOPnUfFP89ggE3s9K94Yq430AQ9JF2nwbcdZP9c
FUYVWRo7onwj68yCh/hBTSgm80dwguJdlItIuU0eg207X2lYR5hD920tQY+hYDlF
936zd8UznRJCY3+jxV2iEDQtP9ycEbqHFg04uF++zVtlBnXfU1FkDT7wJ7A8W7As
4g1qC7xDr1Q6jGTBvqCF/jNaxMpZbQXnEEeNYqXB0e4N7ToQTcXgQcko63A6f/jd
0CZKFtFv4s/hTtfXYnXlHMJ/JDWoK7+qny3q4x/5rKzws3cg+I0N8Feh3LZF+wgn
SMhfhFkvBdF9p0QXvvrmDJ/1kSpPLh1T62ZtzZZYhn8JqFc8WthfT07m4ofr27XK
D/3zRN1VP/F0m9F1tRsfbzvb8TPaZHsbAyHV9YkCpaNCYMDgUOT//yb0jhd9uqFR
6m9sFDvx4mSA0IswNbHEweZHgfqBvoeO4Dvt6LMHhSE8hbDL1w/5kbHDObbrMswv
CnZkknTU3Q8smmkwyqvRs3lVoTu/k3sU6JgeH4eJhFRF7iVH79VZeeC8Pm8PsySR
kFODq9hz5jkegT9P2UKnfqaZYB2Vuy9GryBjzmxqToaRmWwoX0AyODDeclRBN9O4
YMzmWKQWiQvyMX/Lqa+0Mzb+Ebsyb5e6PRxR3kdVB1Z0sjleD7+4GqiflnLIX6Cq
VhiFHduIHGJzrzLQmALR2jWUEbLuSHHnl0QfWuzzqDNOcZ90qjuEVwSTqglmU/fj
2a+maacvp8iisrcSQvJGKK+inp1F3tnCJcHLRaLBfaXMtFjhkcaZOpwYuFLvN1SP
OBu10SXlLQzLErKc9fLCrAzzWwT8KGsiwDkfSUU7DTZ+jnwEYcOU6d2/sr0UzARv
J9rFu7ITXjX+FzpZd1uS6+FywaIafx7TnsyJdQ4tJa8x8P2o4g/ItX+R2mKZpmvO
BSiS/bsFi7GXwGKKY01XfDEI1EW8lyTL/BvoMuxeST5tJyuhlw8iwetZhn4SYNvd
PC+etcy5lBJfU512MUJZwfnvT/ujhB00P7Uprm9z5eRfj1DDcJnrPLj0YwqcYCzK
yX+SR4z06YnRKjq2dX4htOb60pklMllkfjmYPJkJCIKnrvZ8edWN4n3MQQgqQydL
gEg7RijsovINsjcSFtXnmi7Teo/LqKktds/gI7FwbPkrsA+58XJHsq753/3xy/Q1
AFdQnwA0AVWk+a/31+fnkDUDAhP7rDTpu+TaGCUlmfO7B88E2iwt7xlBezyX6M1U
LYnanE3vC/E9UylfGU+5Lb34HZAcUFhfSbszM1TUMsNfG98LjKhCzlE7dFbDVZRI
B1/Vi8jt1A/8Ce8YRpjzosYOT070Pwnd/fpix6wYCidvrewCy0Au3w4BhcoJjp/c
QvZrr7nOfrKatduikch8Tz+Aej7w/qD9mCva28eUtauzXDYlSOTdOLFAfOovhKu4
T5XC64vw3wdlGv5GwmpccQkr+2wluPMi3sevtnppP1dGa+JWiEKeS1djRVeUMW1H
t4mD0kwkxVKTPfJhZAnBbLknyo75bj6xgaLzDacI0ihS3S+8s9comP/tSGPNLHZu
igyRpU4XDcTlw0k2K7+RW+ABCwWnrwpFqg6PkYL8CIXd+IZcnNzboiWyS4L46qM+
94JzoKZV6WF8+4IR9CD8STUXUS95+UJgSvseu/nXtlgkqhtejT9gYC4lob/AsXMk
23Rc9dM56yEddndy7yFGHoTE+8tmS0kZGXDakGzGEbqChhpfCCoxvwC/yxXNnHgH
duckF8hc4gLhHPlmhhvo/03qkN0Y5ZN/JK928B0lBYqeEMsQjWtE/FMSoPd/F6Ej
os98fLF47b6uLndY9qDxheuPYYs4mT1eL4sZ68GZZIUdfNdfauWr8+Of7cKknbLJ
n5QlM9dQgTPTVLeqclf+Sf47s65Q4/LyD7ycH8FAmNTUMhWNuSV/4yyNM5s8TX5R
ncDkoLj6Fl7i2eZHYx8/CY+vTSWwhuVQVPJ2ARwAqgK9nFfu1E6W37H3wClYkCF6
ptoINj8Xb+BKpVzWyG8ZzG41Z7JG1hRx/dBAbzuDDjsZ8SSg8b+yCv3PktcHc6i4
8lOh9yXUrfqpcVv0PJM3IbWND+Fo+LZJFiAtJjwUV68PCowwaedhga4cV4nye3BC
HsO/ca/68ZGXxzrzeRXAlTLxKhBDv68rGToy34HV+2jDoakISIXW22Z9NKA/HY2L
chTFXg3nwgvCZgYieiXw+ciLUT/9GP2mb0hd0ufwl8Js6/k6an3sy1DYNR4t2Qnk
OoxiTPjD+U7igck/G5ESnZDdvUTqEGtciCoZNnN6Oki4jr7TKJ+KI4L09QBCMoUA
SyotSU6YJ4Ws5Jva9082u3n0CfXU8ict0OyiuiIHD/Bysb8AGob9bdWHbRbbmgOr
PY7fhOWrzunNU6bIp/JunvfCcfzE10bUxMVP0jKPK6R7nM2d08Zc6IuggC9TSQpf
4ovNhXtgGrZn7+MMSLee5DZ0jbz4RebTUjQzsVhKeWriKntEJ2ivjr9u5QaSzGIJ
fINXDc1YK0jE14hBCjDX3OMnViUoTFcajEjpI0Lt0bCGeMUcQTWMfTG74oXGyZbb
FnXsXs7o4oh4uBbzxAPrdXRQ7eGq+GpLMstKvvHylQrVTJIe5+EWz4xqqglvpaOc
gPDq7nw9t7KOyJ3QDyU8AoZdexs1c7nG6cS8HDDS37m4vBKKmIqF9x7GSTIyhKoS
HXqFx0rhuTxpYZTNHEImpDwCFz0DanyoiYwSb7GKYGbdy9ZSi8mtmlrGoXqQYqLM
7beDuECTPRkOM3PoXk25YqCJ057z9fxXeG4iv325gDEJiirXTr2FOxn/EOSWDmBl
insh7ws4U295a3hiwU+L/aqZki3lpS4b0a3EtZ3jqjlPPwADYQQUl1lHlXowUcqi
tz53d5Ca188VU3fe3XWmlYNxy/QEyFequ+z0VI0nA8DSHq4pgAPeJml22LqHfoe5
dfjNsnHwKPjHfY8uMr1FNjZ943YMD3L1aPqVlzWzNpVp//1y43E8+79BLWRLhvvc
4Nko+2UFZWxnUNM2iREcA0sPsW1nJrHo/AR0PDqzDL2NRp7MMapIA6HjugZxwpJq
iDlBbEAVUuGp/zWNFxMwnrQ9/BJ3jZWXyxm9jyvyfjATQ7Ht1WBB50PcModHXFRc
vE/iHNV+Cm5e2mhsi19fGOsNxMOClaBJ07iqw+v1HKlcl0X5pX6LY5el1uZNml4+
Fk5C3jy+LuuLXZQ98leAiCunKw27NCRdFI2tkbzw7RBHmrz+TP7rvnCUoka96WVn
cXfbMv99fzwXUfGuShnyiplmQl8naQEwnUxHp2ZuURT8eGXlF0owi9tIKJndT4Or
gxJw20raz5pAQzzZ9WQGjmNPxu7CCiBKgtfZgmEcE3F+6r0ICGZryejZfLJ/mjV8
p5F6cUotH22ZGEIa17ykFaL26MbFL6zbDOyQx1RsQF7VTivUXWZSHzPm/6mSZO43
jP2UTIrwXpADwYTdeVUJzbDbb+esZPiuLAtUg7UJNSYOd6y3U4holYp0clfUFTgQ
kCzCVNrziP6oMJpfgErxLki1fWtNXxLDUiP7zsFCC2HiJO1QCUIchz/57vOf3iBZ
VEHXs+vuZ6V5d5zB2OzvSEGJRke9JnBslUouuypoHFD9T/6cuE1VgiHJ8uDwa6Ml
FfGoLjrfF0kg8SCGB3dRrF1Nk5yJiy1aGvZox+BLyHNQ1JLGMxKFsSCI8pmNbtDp
5gz1LJReE577qkWXn7VSrTPEzT5HEY3i8D1yADHor+hOZV3DJ7vVZg6qZWQfAWNZ
/qZZUDjbnVhb6nQ+dlYUhBlV4mRO7tmA/2mpNczV4EvOEkkPbcr+5OLP9h2CFsaK
oKQ3XG3Lf8CXrp/piIOGUwRONJvQPJTPF+nT+HWZMJEqWOsdQKBn75btncipci0p
2Pl/JdB19fAOgaNcgI/aVQ5vkFh5X0bnmn9X2IVEjvKQQjESWQwrEl1EuFbDzJRi
Zuh+OHBbDeX8AYRBVKqKjqoKBxMizc4U+SZV1AUYuuFKodMIuWWT698hUuyiAVt4
fTBRldLYw689BzNj+KhcwFNcSP8Il8c3BdQ59WGDP2SDsF+Y9PsEms7RKS8Nekqc
UU6UZiaRraeAQnWR9e8zidF6HktUDx7/fh+HhpMWUBkJzvMhIjQma/PbaJwCzteS
GjfMmfCnwoOUNDZB/UNC4g2/iMs5GFIuZBHlEGOa0tVtopYDBFEwc12k7qfCGBGb
dQ/6JS3CCHhkP/No/ln5O6pTWXFBE7J51NQZZOS8sB9xjlkAsZBdai7ZC/DssU19
r2oBmW9hn/Mcx83gRAH7Bv1G0wiwV7VpQb6tKTiwTkImp4GQOx0Q2zTd58/+HruD
loOryZHBNJivHcdTIJh00HwrvF7Vt5QV+3mtvDc1vmz+nf9KiMyptFvoqpvVMf2l
eHz0iuwwIXFa2XR2Ju3jO9OkwdveEmSUWflXGAvMsHiCqfughj3OgDNWte05Cy0E
vuCkfsajnamxAYhKVEuw0DcDryU21nshSK7lIK+9VuiMM+E9xTv89cm4QvBSKZhL
L7aHl3lvZ2Av5Ilgsz0TNnmInNqwUw4CuEAVQAibBIjsWHDNEPqV+5EGGkEcnlAq
+Dz/IxwPkyb4W9W40flvgKu0RZDiaxY7934HKZvVJikiLTvv9aNxrJdNTMkP6wfn
nNf5sSiEo2+PCpvpDBjvuhrK/w7Oion4m0uBJH6Dtc4ySMsga56f+nVWqhO0Apbi
4L9d/XOsZ4idTOjp4Cqs6WMCYI9MCiG36DFXLl5lVwDBwe6zR3rTjVS1ezjjSxZu
g6NE/j16UZxXqfnQcvGoI6mFu8Sm58VARut6H+t4W6REWvmoGmEe7fStX+HHsbfo
nFYvbXWZUjSrIYX13USimYSiJoRnH4H52ekbqkvWYva+DtvaRYn6EGUSADeadXun
EKY+AkxTXN8Oj5jVaSev4bArHKLxgiBLjVC94cxYSCLXMb1EfMaoklM6adYhiNwv
5NVCUdWf3/n71b0q0wOuTinDYyXcppHPvgYbtkLnfM0gfOjm5LaDVolFHWIOE7bt
oiRipHJeOo1aG1MqGYQRoPZjWRlCDGiPMa9tL6GSgTzI2q3VDZHRe5h3O6XxRUaJ
FVUDBuA6qIgd8M0TLCazXtkFIQT4552/fELJrQwkFsiXaMDyHsx5sy/MJQhWsFya
zETXLO/jevxZra+qKyeyUrbSCVaOorDkjkp6DOAfDciYo+JlMOGNA0em+Ho8p9uf
JadDuktAKqd4ejcMyzpTjvRBnz8MUlNhjlpalMug7NRuGvBzgY07MrHZ2Pa7L/ux
Ydl2tKl00wbxKbC+V70a18GTY9/tHHLJvr4lHcdVmcybHtYeyZXJLhymaZO1YT7u
vU+Ux36YUQIIevqv1o04Xned64xr3NeyOTZKR64quHSsl/ro1JvUaEOnSvya6E+K
0kbUY47MNXOVNomj+EHW58/FqzPjXZg4HJLkN6m31K/IgyR2OttRMUfZZjFWoQaK
k+WohKSrzvR+B/0FeXaBDTf4akmR6KFtLamCo14+my0Nre+urThGrkSO5L3r/fKR
nGijiOKxpNC72vBBvSsvEkX/aiUWUADmIJ4zZRI796OGQMWzlajkwPoEW3s4dVRl
+XclqlLORl9SmfDEbcvHCTzXqhFfZRKur9GtumLDMsPjkOsOIAv+/P7BD52Vvnzm
j31LHk1y/ocnQSznbwTwrbiEQODZJh48H0EezSVshYmeXHPHAFBf5/YG+cqGHdvB
ewy/dVlCLZkKwJrOwUcpDG47mbARilZenubk1/C4CviQkQPN3v/U5G982GYf0wl/
3o+UVknANwb1EJxajG0yori8DtHDFv6XmDuqQ49z2zbE3roNuPeGw/M+6vCIVri7
SHeusbu/tASmcuUHaVWBxGSsuU8mWkx6Yc2ncFNBnCJ7QNM3YYIlWt2bE9sz6h0Y
31A/6fG9nZ1fL4lRkoCF+oRJ5gMWQHIYh3pKpsLFVl4GOcliUWzM9qCh+0mrmPia
1TyNr/XFrVQiEOMC/4q5M1/jxDyTT2u4F0JnY650Gmta/Ti/nwRWFbWPeudZIoA5
/EaVh93o1k19vPxZP5ak7+ic4xPpLYfThyh3kY5xKARQDk7Y3aWiFpREmoaJ6JaC
RIwffnQZIM4E/1cB0yaM+sl76xwrq2Tc2DDDBnTCeabJEZGee4e7bNpxDe9o+SX8
M6Us9mAfNu/RGeDThCC3rlhohXcsx1teBt6Z3iO2/ylFDq3QP8ZmyCMG2YkXqjCv
ylnculMzzq9ZPU8EUXhVMEUjrJDc/tb8jAyLrioprz0wKrcg98iCEoA0YsAMvFmc
0AWf8y/+TdeC3/T62GmM1LsNEcfQ3Off+JHfjoN3VgtIJZAszR+Jl+IOcS75bVKP
6IHH3ctsanxv3NYQYTDcupKawOlt73NcHXoU6Ua+oHRDHkozfNkV7BoG/ORPLgk+
TRv5pPS4yIMqL6TaRAKree2D013ENPOA/4L+EYh8NUaeGikbkZTJ8m823pORNgEO
NJWmluznxgDsSivncDD2Cw2y8zw6oYf/lbrewQ98mdLUoaFkU9AuOPzbUPar123I
s6OJ24dLtwhAe4ttM9YS2Ut50RdlxDI28J3qnOKDXYilWVroVLd5L2dmglCe+mxD
D0ayGdFcbM66DnhC2r8uX1WsfNE3XSsH6ttklL/STYjmOsTq9pWtVD/hc2csewj8
93N8usxKDadqU1KrS8AA3OOkeJ9giDwZyJDFi2B8f1B8Bm8R5Y5+aVv31W+DxYrT
tALgLZz5KDZ25tReQxMtTAqwQ55UeSKhJWOznO+tFqTXYOg/Y3EktNe5KHjfw679
Lpmr4b+pZZf3NPukSU0eMksgkdL1lut/2KQ/ZYvWlWY2FS52tnP8kzowuCmp1of1
KgbfPeMWZyjS7CypXQCGWghHwGiBdV0nStcNtV0PElt0ZlTswAvLhiWBn8TbFZZV
HoNURPcXXTDbFjaX1b/40wwmjh9mgzwCfYz4l7UDoz/o/9QONKbhBRFGbMeBfFeI
uLZqhtnQpEfxUtO0XIpI4iFstLTm356XRfI348tgCfVMAph94j+plbFzxlUAAEus
QEiPrUhMmbTkuPG5jRMU7fw0yz7Yw8NNif7k1KtZL3hSewu2G3Mx1JuCN61oRX4H
t6nb5UmS9b1aIOZ8RJAmbnTentAiO6472mKFQtSAp6gF3Yysvsx+9uXnz9DpCLWA
blqYzGf2WyZf+fJ0zw2Gu4tcV4+Y+LyU90dSGFE1wqd7FWFJ1NeGmvwylAifwJfi
qkoU7DCuM0lkwDeazoCNaoAh/D3dYDuvOeAPeZ7hUnqKfA3Vu2aUPhBU6ZOP8tHD
yr06rEpIgcpD4M7HSnrqU0UMatRkZfB9UH0VmXMpcUByu7G3UQ8C6ZFPyb1WqAsV
KnlKh+36A7O9CAvHXE88joJdBAnKmtYqGcvXKFC/mEmMKeye+Xwx/9FOKpmzvsRn
pTPQPG/2ksAcH2BCUH3ANX0vTtto+vZNjO5uDLhzg5rq2CKrtvBj7EzNMD0U824d
CGgyHL2QgbqWZPpCmq5FM8IUh6FvPNmFp6H2ByKuGE/WLmDNlI/6Am3DsQ9nTyj3
bSyICYQVBzdMEEKog2i6YSYQt8PYUmjn2m2wFk1L7iDk1BpulqDWA2Ot0P+MdqAW
iSqQqp0vAlB6I+jKZP9Vq8B6OGb9p0weqK8mbCdQuvaBemgD0Wruv3nk7/giJZgF
9jNICJpuokQ7aLUttJkFJI6Yr4XKKv/ADrfpmy3DX3NhHQoDxwZ2H0eApUFwdIs4
BXalcpANM8z589C+Wuu68a19elPRSP4SF+hToZwQtBatBktTh/iUf9k0KU2+KrsD
NLTwBRqN3ZxJSSfdUvRgSoNEHPGQZxurFqPCwvHUtPN2+PWycBiOGwQWwF1jO6LZ
hFONmMd/UxEQPbqtdDA2FZQ3d1ZqpK9D7RVfTlQFWBrrSObPsHdWd3KZkh0lK8Xa
oK4lMYDoo0gnX9WtGHSkLMnvHxHtfkXyBcjmiYhpHWmUcMUeeeQ59qC6c/ZIAOM2
j6xm0NHZ9LmXLp+HjyRLIrayoDzQF7OmW5WPY7u+aU3mdfdkuwVkB7QzUm0rjAYI
wkooOr5XGQTVmD8u/CCSq4dzguGn4SsMA3YBaw7s3lFCvqksvujQwDCXIjVuG/a/
aYDtY2BXxBXJbq+gww+gM9BZIlGOzou5NUvhnP0qwLSZlOvC5HH9c41lRD7dKaGA
nBfiiIzD87nFU3kFEJ9FOMKa1cn6cwFSKL9/W9qEDr9A8Dr779XNTTgf1HRn8TQ2
wFpS1Skojoyb+YH2ciwW418XYfSe/mnvub+f0eOGcys7tOtI+9M6/HS5BBP9CGF6
S6H7bZEzOCKjLo/CQ/DN5iLWTgSPaHf5aFsz9f3SuZ+qi8JnMskYUo5mnJ+SwAvA
/Nj3FwP3Btj9vAD9MY/TsOMTnPYhQnT+uciA/3hkJZMA957GyWIMCOHiCbQI75ga
CWIp7VrO3OlqCyKF1TVJMnDIJjspBuq2jPHIr7Xb1Ir/WIciCXJPHw8yq8iOybSV
AsEGdGd0K712S0bT7dJhDzx+nxAoQxznBPg8KUS11US8Z54up1VhZG6dXEczx+wB
ERqYOrWLfhFefxSSr3+hjSKnq42aA+U2BBUXFkvsN4dYvKkMtTE1/WrYXr7Mdy0L
MiDaU7d+U+L+D/GoScyIQUm+czCm5g5b/M8vh/qVfEWJ8V//SFjhwkttwoOBVoHR
gUh8tCJY+1mpodH6PuAZFJqlWhzEKyM09ro7On0axOHiQxPc8xRE2li81uIEQxz/
RmYP4ii9vV4mlCRcTQPUEqLmWI0edy4t4XXbf1Cy7Yfz+2kqG3aY1sSKs1OBekQQ
bwdX8zo12M0v05VGBW4FsQJaibox9RyuR8Ya5H0qjL76z5d6PQ20oFfCeEr6WlfA
yc3JO/SPok3qCRjZmnSfklIXLO/AHZNNU9udwdEYwcLF8CLftd5y+Tbam2ytn2H7
7HRcCDMB73VweQ0YkCeY/XItePKm9VYsy+sxfFL5afbdBVLDu8bzXCDQjPwrx8Bx
YCbPDUPVZfjK5iUViATPQGkGZdRSwr9PBPPhLU8t1Jkxkz/vakAsRtOYK7JtkvFn
q2dtTMeme0fCxHn/kqYJaBr3U5ry27bJhSMIP96S9qNB0tLNiW9mfh7muP6ZxK3o
PfOjEn/gAAeS/tBQgaN3d9eGdy769MQ+g/wyITFWiGxwjJOaFAQMZ9S3OIxlOXk2
6puKknVnrdCo5fbO8lN2mbhgDNfXVcNpCHfPprMNfnDAchF4cDoDa9fetVdQQCuQ
L6s2BSVuBddEcmlJSF2t0upGKVkKlRf6Q/QbWORZD1w0ww5bO6G5dl1KgHeyXqMb
m6cC1I//zaxI59jg2Hl5wyGhMehVh8UHaBL7ZTjtTJBJZrl+hMvJzRVBGbQj0N2u
1vq/pwtOs6jbB5Tx7apDGwWPIABW/3HU0sQvmsmFbOUB+klBFrmNIrrDZjnHz3xI
0QqxkKnbyT/IxnACVLBCVO35PleDDvWxjmDV+ZfmOq5pJqhKrIbIauvpzHOFd0Ts
TNgOFgZsIMBZm5WT1RiE8ivXH8oEsy/Ax/0DLKNPF16cpkVOKd0rypCtXm/F1YVb
4r2yzlHg20SjOdLGpulR6huC/eGONDOeuMhk2MP0Jh4F/HC4QQyi7NYjvWmS8+04
fjOqkV1ucS9LW+ov0WySbH6Kkzdq2/Czi3nWUIGxhIFyZUm6o97V1lUoRnWM3e5T
A5jOu8/psBjLpeZ/czvMYz1u74cNMzUDkEoAtHaeQtZjCmooE7jKEXABHMrUGl3c
Hc8xIQixCW6eetnchMAaBqjF891T7uCHuCoVzmnQB4Phgy+FPXPb424g/cz1SHWg
pr06Pp6DPkYoaw3CWpGtlKlOwMTXaXAf8UwXvNyMpHa/bxp7sUVbbF7ejvbZCjvA
D0xJiMG4JvDF3jF7DwIPfnrLenNzDfdCXcwEg+jcap5cU6nJcXoYKtl70+B+pYtd
ybOf4F5lCsYJVRpqYLqkORniJpbPBwq9LZgf0JCmOBo2aXoUnM3FDYtkmyjdQREH
554xd1LkSSocOo3rYjU80TGFj5sTnoy7LuVmasErzmzlI0GCMzsYCTRgkyRo0KvJ
SBcfWj0TFqlLiGFcxtmBRUeA0firpUKD29hl+OrZuGWKrLUh7TtmlAYJCXnTTQCf
R1ChOJHjpcYdlFt0mYZUithx7uGB6fpGcwk+s4ZRHxOD4S8+GmREy7z8N0qzqD6I
7Uot0Sav8AKTVqqoHxOe69n4zcyGV9R88j4/kTfor1k7I9uNOICPOOAnML8V796M
6vPJuddcpYN35MWzB8FO0Modm4jYvGPUnTGBsY9HYA7yyFyI+kte3FhySEuoQ7x3
4w19mYZfb86K2FaO/+oGb+mSmM+RheWan9qwwmq/bAie1bmesmGci5I4eZHubhPm
aGW4psC5vpqCxxdu3HXVtdoQlXN2PLYZ86LRN0+QCSl+PnXUGnI9kxBMfQ6Tno+Y
ivn/u06SXVW0KKa7sR3kVD2pb3KIk4tFKS4Ang16ArcYsnPMz/DTZbtPfvYGc1kT
C6T/3OHKXcGrv1OWTAouzkxcnyQI9Xq6Eqj+6jJglEf2jVGKPwsVrWa6iieoK6x2
I2AxC37Cu28+FmMbpOIjiNeemTxH7u7/l7Hv4iWJmXuiYZJ4MmUX53Ayt9BGSA12
SgF5yBHInixphJ5jMTdXku7ctZaeU3zsZeCiTIq/dAy6sIOWpWPhX4+uKLX2gO2C
ARI7nEyUwmzBs2u3NIP+KRoK7GuC/+gGip6V9vfubZ+qdMVWbl5jyMvzE2yzNBHl
S5MMUhec+rNdnJ7J5lY7cONo05nHnriweqGEqZdp8hodYFlDLEkzzaQp0Td5Hnyr
l5k3SOyBr0IYYvg7YfCdjodyFmmbKUgFxeVMB8aClPQA9FgUxb9fE07BVk/z9fF6
/Hfgz6UtvKaPLjrpMdGJnEY5FxIbOiukojQQaLX1OImiFohTBGP20ey+1hC3Mnp9
HGCvFEi0vmRy8MNVJGthXgffdSUht2MpxY7UIB+tm4topSiTtKxLAHXkTkoAKVrA
IwKcFaZwT66U1HQCHd4TX7VeoEXzS1LIz+fLRvzgGSJdQ8+X5mDYxUb02WM3GzEm
C0lOM7gImNgVsdqE2CUb4jxNXPZcxmVNPO0Ooz4RBzZPw61laqSNqhvwx7phXszt
vtUWePqfX04zeq/VRr7sFh/9x1DI3NSk3Gb+2ta/avdIu056roIrmgHT3vM3QWi1
o4Yw7hd+JC3xyTrOsoHitQmtUUIXFyrQxA/JsLgnyoVUpT0O3yxzQTMQQOMvwDXs
HEUhtt1HgEBdIGPZPYz+d8qJogC3iIdwODBNVmGhU+D/ZC5rxWt+MkoT0+YIfZWi
zLdXEI/QmI+xYxecFiqx8Z4Cbt+v5teLdy16dFlnrRY2VzO6JiEaIHm2skCjowr+
FAAEjOw8R9NQpyNMbK1eU4bArBjUEaqI8wruF41jMWcnmb751HqQs3IXXN0n/umX
9bajU/zk/pQnEcGEmyRac0IrMVjUTVgZGP3oFWkjPlHmqDnWLMauXlaogyPdLbeM
EPTJPJJddqp5Eus07Xp4qKRle5hbBa/HUTNIFIJAEqhznUB4w/LKrr44BA2adh9G
hhgzuP93JMAk+uLtl1sqwHh5XcfXzlPjoPWN7eOLMDEVntsoHO0F8JnotFRvWc3w
9m9mcVw+OOaEJDnPqDsHEXiVOZq6xCmsnJi13kQNQopfEcF5oIaLNloAYTVxWg24
SlazykVThmruVe0e5yOHNYwt8rZIUp2Bep+5U+tXUPfKWWwYO43WtUpe86EKPURg
dNUgti6maOSjsBi5jtV+L8SnJfPi/LuRVIpKnAClWBB6WxgLCb8GUPK/lD5gvjR1
iSTGA5YnJaNeG9aSTbPsA1vDffc9uxSuHrh0it7zkCjNkdcnAFrUHCvxVayXt4ma
IZOBUjf8hilRC/2T6RO1ukr78AiBh3OrZOT7QSlQSl16x+AFm7OpNmbxWn9UYJn+
gJKV8OMxUHIafjYGAozQASXAs1SOPWH/wkBBjDHdhCPWbnPRbHxhb+mokD8rSSbL
5BfPxANPD5T8gqhE9Dd8DSqQzh3+Z8bQt6P1a/dc9e8OzEhIQ2NbYkn6s6XICjAV
RasUVNZkzV2XVMIeS94Lv54nzOl96Vypo/KjgklXCjSNA2h8m7q9QEzcHEhTY6xI
Jm720kv+Yn9DJDLCFurMN8gVdFWbo5Ud7OIR8d4LEYy0Zqji+90JQeCy5fkkwIKI
dE1ATnE6VF1FEawAUDnXif1wpQrCgKmJ26Ylrbi+tzXLLksrZjFEp3Rg+vPf64Db
v/AiBmx8GldMZNf0Kzvip4yVQ88stySNxN5RpdVPdPc6BJnILUM/dz20z9T/oLDp
O4MDpk6D2gv7h8vTrpMdWQWnV9q7/2Eft/a0R6qFBRhzWWSZKd1VO1diB3HNuAI3
Y3Mdr6NDbdw4zV53Vq/TFCjk1nhAR+1pTZmSU3wqXUxGZdA3BogWlUhzpNkIDxGv
eQJ+8gzv6CQqvcXpe8iBI1/+kNpcU7u9Q9abAl/y8duLpWsr5gfbrGqRyloZjD+3
91JCx/FeJtVhWAHIvTUnWupJpw2bgQJYv3b2wTUW4skVTxwYOTVfe4Xnn/8tNPTs
WmwLtz9HsZxJSVvsoWgYSRPwPakSszOKnS6qn1LxC5NBV/gQeIMSSDH8eOuYgdFx
HXR+ijrMeJ3GUnXm5LJnBuCbHMuTFKfjeEdiXkIIOAlS75uJ51VKWaEPtvIh2cg5
4dduMLCkmEeEQrGMQe7Pg4PLu+3LjNmHCUdqOfx9lHC8QNlKrE0i5sJyR2gZvPuo
is2MMZ6CVAWGZCwMhV65ujtbPJ4AAkXOOm/uhAgIVGSovPwaA/A4B3GB5hO5ohEk
OlrDWdF+Vtfhc7f48hiqZKVuytKUk0XRbeW6LNPqVOshMiRxTUqW2Ut14WrzwWlS
bKKKZPrrHiHfsKkGPivBuvtEvsCIZUyjA0RnGzxH7nk1LDCcdbFw00X0wq31lf7o
ly4bTrxiYnuECKzyFHrkpNwov40chzlFtqX/m6cHc9SFwMmLIK/PuAeo6T2Kf7hB
dMamlftZnahEi6D+OE017odjYCtjexlbImySiAN7zDBVvREGZ2UMY156GbxYp0qA
qPiFX5G0l3iEWJm1GRU3nIQ/ED5MbEO7fURaWDqIqOF7jKH+8PROIHdEtriEtFeX
mSStOBnbAiqdtfK6o5XsfSxZaajQ+6+r4PGjcNdazeaF0BIo2rxCSGL0NfT/+FvM
GXIgfttT2FQE8nlpi/udKvCKM8rYVHsQ6g4CwrqAoHE3qo7/WU6oFRanpMQoc5q2
Eix+VR9Xe42RKknbqah3qLUBbII99yHwFGgO4/jZ/vblOSSycdD/1gY1KfmVagEE
fLHhGXg49xWu7rI6Wz6hZY4qG664xwYeGLQ5PBOW14/aU50BAAg2rmSMoQ97HaNF
f+zTDHcD5KRzVtR99z3AHxz5eiZOTGNxUX5KzslT//ejEK24EB9BKb20/hR78JAe
v34DqnOhTodpk64NVGDnzm/ZmTbuTcSWGcOERAEHDFfwPE4DdxYcP40XElKVWBz/
ioecSR4ra9mQPm+0gwS9kYOKxiosP4RG/f8cDbFXFrEP3hVhIaD2NsUEE7Xo12VO
4/Qsl80QziWd5otR0LaluHvbWlkrm9b707NoY2yJ5Fa1dk7wfmEme2Z7XmzU2PWH
RDBCE+rXoPXMnQ6+lvgA4g5OdenGqrqLQqmTpWILaZy6fVy+BSmvO2tInQNh0Yr5
VjkG68XI8xzoAqcA4GbBqSv6Yv/pSapnVpXkhNccm8lInI7JIeYr/7BujWwHGoMS
+ToGftOuNFLpjvQBxDv25wh1GXdfx4B2L72hmEaat+WdCuUFihdy/kdl9RQBMN+v
qG/F/T3GDOYKXHELSK/COkFZSaQsohNWiGCrs9iKmTPb8wCbsgZMPX8pKBrU3NDR
5zJFMWMcHv8yIFdUNQjzuuTRIpHy1ZjGwCCqKmxMmgKkbnwsCZsxuYtSTgESRT2N
a60v3ppGwFHChhvZSlZpxZXRvP6g/utbfbbW1LF/My6NK/3ALPkuxpl0GSQClsiJ
H3ivQC/q/f3Px6q+9SCdTCA7US6wI2sjMUqAQ8BUrvztpx286BJtaOK2uwWCdLzz
qpvKTQgCOCNqugTXXlGU6T0E8+APyuuI6Dfqqr+/6Rc90IwOwxqQNT0pTnRRVxQ4
S0Iv7YYK2RYIkEQgecMUlg5tvMcA8atrVAOwtA1vrME+MKm26WLxy3X0ETTcR39C
bWSF99dY0CrDonnCUWVRpV6RVY0w2DgTKwstl8qWPnTByNwVyjDePYSldMcNVjVs
CX152gu2pDYSnS0UTr3q6scqURIgz4BTuSYk+iNsoMu16as+m6/XSGBizCTyoFDm
dVFfClSbT8UiXeNMA/gPbbO/q22LcULUw7hvWlzsjoTBXJx+buAMsSn/Ja4U9BL4
o3hiep9sBvesdnnippxBQ5WNFLN94q+CgncqGf6hUxm2PFm7AcdhPmjOcJZWFp+T
tGoImN5371NadcTUetVJ+OpOB+lkkIjFFGYvY1wkN6Gt6hX2O/LkYiPDN44FG5zz
qMBScaS98zqYfz6GtkL4/lus1t4n5bCJylYyB3bkhN1f18m0fa8yr1wRPr4zVKWV
J3w2BIqc3cZx2DOlXagXp2KCPq6vD2eflCa1IKZMYr7MD2UAdrlttrDpng4dBuP3
aHOZQ3oLVF7X9aVuq1B8FIbMLzRvLs6mg6kMvqsncqSgE8gMf0hUlUkztHdQixS9
TaknWwPpHCaYpSEmbXVwJY+3B4eZBiidosTLrNwgoOdjRM1yNWGda1XnNEq9xW/9
m2uli3Dd7s2rWdgnCRxW7N76zyfyBUsnZ7P3KCaeSOY9hD0F4hHDDi5eHT1shU6p
PipqcfhVEkHxAMZyYrdPqnnOJX/dsMN/UcosT6avXtzZy7vwlz0+ltdxyJH92k8/
FPngOJPECndhRYNNM1AhQaptFa13diNZGWuVEOuG18CRIEEfe02xetPSLmyaZ2Mq
fv1nXOIhicEuxl01jS1cT0u0ffC3KUDyWX1tRpdhmRunV5Bg7EV4kKsBdt1x7Ba4
lRzWi/2CfAjcQ9cEKyiLCNzbHLWMe++YVOKAK+/x8etMzAhdr2OlpdabwJBsIGXp
xG3P6guEN1oKyQ6gOw+v0HCQAYqaFx6MzsBwqE8X9W/lUN6EOfF0gNAsiiQ59zAz
Cr2pHk6P7uG6Lv+lxvzTXaPHZdhO+BHhVvqdrbv99h8yq+XZxNSDES3vd4Z1qtPF
7Ee4vdSttedNO/alJpNB0AgREEDNxCCPzy2810Hfu4c8YhcMSwvvos7naH4I8JMp
bRfHJuy9LEYA+ulIv1UMfk7nf0HFt9s4hDrCYTeYlFJaMRJ2J/oSsKCeqsT0RaQP
cf+LkyFleMFAg5LYtU2KcbkmRLH2dH5SHXIrhoGqsu0zaGinEQPKKmhZXl4hv95F
ChHA3Dtae5L9DAoz1z7iAEoFMh1C/TT7ETF3NG4W08MlBvSQcB0ge7wcY9xtg0qs
d448k5SQfuJclIGvm29DmAtcSY9ctluJX5wErgXNfz6AfjyB9jv2WsWN5cObJ2sK
08duiOYhIy+UL3buPcpHJh7GhqMavakm42U5Rvn9YP2mf9QnNYkolLTmrX6EdJVd
Rg/hxynvzyT1A8qMkCeO4jlKRM9y8JLIqFz9KtKks8hmkraLVTK4afCJQlClmyv0
pNxxo3g2ctC3onlCkVAjaFxl8jcAigRFKi7A1KoO7fxg1OHJYNG3gmShkSJ8qipC
k5LWlXmrSOmjgmlKMfU3X1nhLMjIcjHJ5AhBqOT21z8VGYG8053MsDZrt8rRkNXs
osFj7Nl5P1c50XEgJdDhn+d6lw9Ia/shypoJcb3vS0nEVJpI+t5qXx3EblSc64bK
sfI8CWm7Zl7F3TCdzsNQlmHeVieFp1zF7FFj9vNIN+jSMgfEZ1EjrxJSMi0aRPS3
yvaNexz7fmRvNrybxq7/xd5JvDduMIJFJdyrLW7piDaZtEex/p/TrOWvaaJO89KJ
k0Ha3EEQGdqo8ugoNiiWfJ9qFB52R6+JVB9++ar5YYvsq89shbE6gllgGZojQzwy
hG4Oze44vFlJLdSww+iv4WWaE3hmgm9gK0rE7HXoP4E13NbySWFJjLVmmG/EDHAt
VrXotKH8yieCN6qL0jhYOl+vE3wiySsC8S6n14MfrGi4pwZqmjwXvvWABDAQLAma
swxPvzwKKqfVJkj9GGVuZV7hMGsDEcBeUuhB7u2r8BRXDQJ4jRARq/0ddmiaSVAk
hBS2AX+IaAOjp3hURrdh8GXsPTXRPraSLuTdMuBVygRwnxUq/LhAk/FzVkZ7A/oj
7M2q3//ejziNRNlRBxLwLdvNKsOvVaXLpEjuWeG/1eO1Qf1AZg0+7YUfdGCPUt5M
0dTN62d5LkLVwM7A0eSD1A1JUmiXTHHpNSb9x05yD87/ek8zSoJrYGUC7tk3J+S6
BnQYiEIhg+aVPiuCm0GnvAjKM9Z1Qq91WfTL78YL4chLQ9OB0EmkfxTGvoTPI2j9
kZEYCNCjM4KhXjfWJVAchAZ/Hw9g0jiXnl8JQjNiRDSnB3CZJQZJyitZ0mcxUQUT
LtijB+I2aXJ3cA+GnyyQ7tP+MpmTjOj9vnkZySFpxvV5s7wUg8J+w2SJOW/NuKYW
yznQuruIpZmXgQZS2jFi69j+KZfuBB2j1RdTM3FBuPZQSDm/rTaZ4Ba2Cmv53mQ+
SpsdC5zv6ikns/TWYLMZUy9LaFF28f5g5/Xae3zcFJRa5DWxzEtg9A9WV7xw5uzS
xpFLWohsN5YD5Mxvk5J+T0k5I9VrKafzFSSvVVxK3MoA9vK2q9i1f+s8Ek3lM+qm
wFFmLnrazOP28vHl4A4RN8n5W8Eb1OmSdDgmCItw0b9Wvv+YTdeaiIfiVNnRD8P5
ogfemkUD2UWQVuTpf5A1cgAhpfmhTRi+eWJqd7jrzUNlgcRO81BxKiHOs+BYrQ35
knCvhZg6Iyw0Hd0zNVSW2TfwD/CUgfyWB+tGx239BJKw78pVedO1GeQ+8nJg92ez
jXtb9va6qyNZ8akb8NOtPnWZ2uVBGB/oXy1M40kO2/8wZxXYDup17hYuckZlZsx2
wvaGKhG1OU2CxWjxjJD9QM/ptImhG5BR6wk080Z+4wjGP29zLXeLknGNsO2uWPQf
D96O8+9J/kuPKjGLHFnCRtmKgFSiT7HU3G8fgco8TrExHsyOPIS80IKh70LWBSfa
VXxVxcRA/c0YqGJlyP+VdXSa/QZ91IcgaIlBjMewb4Tfed7mmfMa+5suw/zS+rfB
bdMmq1lbrKdsI+LQlIsiG3SM6wv3hE1QNZ4Y4ZRPPGcA0TUAriwouW4QPuahfGT0
KigaIoOMCRb6NqERZj8CQ2id07LWq9XY4YbjdylYyqImmUzKbnp14Lsj8Mg7bnBR
haRvVesXEaLZPb1toJN4KBNVdVyCgGcH5i6uphnix616sRWRSLVFzuNiMMDLi0/A
E9iGVbdqL5IUk23pO6YLzK9beuHDuIXQKQz97ZqAyYV0RukNfVu66eFtHITlJPB2
2DxfhYWxkVnFqJ3ietYA2YQ9FUDi4IHIEl6ZKWdK54e9tqxYG6wc3I9/4+XUEZHU
NUc14AugGl2ufZXIZJ5kCtlHBDEe64iUuUdpvd8lOTvFVdrHRmFZOtoCpeaMqiGn
co126Xt1zZCBbW4UvccscofxXaljqdqVYzXStNxXGlo/TiaavDUVIJyXUBivzDQL
KKg3dm2G9h3eb/FRtCpHg28WC8smLU8t//yZETUkm2RlxiJe9PXUSKkHeks4eyf8
aavannyyQDui937wXmJRkCTBOcUVitzb2dOYtEj58LlCOn4JxCQw/irVbQusXT5p
myZh3ueD3B0uH4gj4H7H+kJ9HnQ/l3TUqZr2QhNt04a83drIjSgIRZw3sEOMk31e
BsidhToMmTKnmfJt1yPZZLYnqbhhGy6IaywOgVfvRvWbZ7KefrzCYJG023j7sHcM
h7mJ4cmtq+GJERroba8uG9EFoiCOxHJaVB81d3QiE62qs6YA8WZUkgiIDNBu9ITD
oZlttiSo9XpjFDd7/uwpV+Mb56yI3nwfqntfFg71e0SKWnA0k3IGm+IC7kemwUWu
XAYdaFD12RkzeLRpQH9wKmoHklgZAuntZTmyp9zNUHA5TX+Atu7ZPBJOejJ5DHmC
TGq237GSxJs5k4w8HQP9KoNUPCFBul3zHmzFrEuTCDWUiQtZliWoHmkJG8WyLK2c
0ThhJWHTKYURrVx933XiQiPFk+dsefb/twQLNpRkkY/aXSq4sQ4O8M9ojuFVNye2
o68Cd5XtI86uUqTN52d7qcnrlbQgTkS3Dihd1/3ZNQE47dkPm8JERbHorbR+w0ij
WjBFWWOFVZNWBOpuLTROOGccS4GnhqG8jEB/+PEvT43TsGgYxrH93ccKHev4obfb
qeXBU5axVWY8lStsmha1KiaKleVepNJwK/U/Z6OLzvp7D5sYn+f6HHNWgPpm+Sqt
BXHTcaO9VwHDVvAt9uv09aINYR05WW8dXm47UqO53d3AjLI3fEKUohma44Mnl5ml
zcqGCIW+k4tXjbIw9k0KcM0d5HA68/jH/Niq8QayDzxYmG10KXk+Zur/3IBZtqTu
1YlSBVbJ5adtlFGNMOSfInQ3vLZMEVv8v34FGb/k10TnqArRu17wo8Np3cwvo2Am
aUkk7YDeuL9CnDoDRdWXUIt018uldXtQJazDT3RuJM/t7cIInJNaB7sJOP1XLAE0
3v02FjSkulUm2OHAltmwGUP92jyIw1qv55EMKxzs0iO7j22ItU190aTvD8r7PtX3
5bVMpnKoxCSsanLq8BC6UnaEZvA5P+KVDn86ZX3YFujpd66VqyJR9aQOC5zx9ykz
0MFfD5DkGL7WzOSQhEPTlK7wicbbqBVzGqA2iYqv/+nxWBnZFmQya1h4JWiykh8m
qzyQPfdv/FmVQ0LcjS6+ONBVeK2SrPBCTdP14poJug4szaXR0ZNMkO6o/1cCln0l
5TZHHijLB18Mg24FN8G1N7hUTUgUWB/i+o5SSjwKLoLZrKfbarBZ+vahCCAzrzgZ
8I6WsbjQHfcu5322/yg9s1aFxLIh4Pu2sEt8CAy5Bn2baK1VRtahDdUCUvbN9zN+
Pa4bdVrvBF6wzU9Qv/KdGQo/OzzyvRqBYJtTlvYKi3V9H+K3QEN86ns1lQYRbuZU
BsG7TO6mgB4PRgUA5SG3kbHWywLaLI1q4a5/c26uarRi+/K7W5TwD8kMOl0b6cZF
6Gw79+/BNSlQYL4eE8ciYnS/CP8svvlIf0Iderl+7VUZbtYWR28o1Ea7Kps6pV5q
vxsnZ4eQSQ/54/XM6seAbVQRJYPFfLnD48/cDeEzYxAM/rfVG9oYlSLaLcSon+PM
gZ3GN0yPVbN4BEFp5ao9g6zkC3py/aWQMthcwD1/ZhQLHKkp+SSJkE2pmGf/3wS0
HRrPj7XiA2vb0Qsd9wp+6wp+6cVR2Q5W79L3/2A7oIiAQaPgrnI9cimSzGpCCPVM
tnfBjiGUxxkpeIyQdeG3HnnGCRtFCrB2HtyquTiBMw5b1q3kCPzB9tCuRoQcwnkj
SZRiyrqvUBJBpeq5q/zl6ccz+QeaF2l0MJ+8DFwOAgtqhyetYNc0JEc99FPydNf4
KTRn+Q9jPDXpAcoD4xdHqFNUvq5kKmnKmLjNdPtZZgs0QfoWNynOCq2TH+lyzyEJ
v+8ZRklfJA6Fas1Hw9usv8EP1ALs8jL1uv0DD2+emgSTAw2OzuF6z/yj8KuZoXAD
od2a7LUvZPmg8p24awngfEblqWmrKFNK80mMhTFhfSGhfG4/uw5FOf4kdPMRa3t4
aEGT2eW2FaapEAVmd6/otKZiJ/Z4uhpQZC7IIjWYXbqOQyztoF8Kkdm7Z8uSl2ek
siciboAbY13afUJ8tLAbDiRJXhvv5kzzcKchAZPU+IJtTCghyJwn40lTzcYN4PPm
f19f6cR9HUSk43HV+0pF61leEsP9x2v6sx5HcqdegnLr0t6ctPMvkODuTEwMHR8B
PRPYDpxTQW2VPFtt8XzLZeA5xZdTATXbPenCxujTUXnsYR006dxxDJG6un8c86lq
IsXmapQhukmTwQZ8MnkLMkC+EaTKZ9muhZpechf5j2SxrB0tp4RfFxvnBVkDsAE8
dUqHDyNz/8V7cKMGdHIKgZoh8zcuO1fi6kE8waMO5/2LyYv6a1H1KgjEKJRF1miS
7He/B2913L2QSjXRekD2SI4rdhYimszxRKL76zAjpTzUuycqlj80MXToC+bef7O0
dZfDIoxL2iJjIHtdgTPGIZDanVIORekLmTY+smXfX/4JIAxLGEcqbwnzSVToQgG7
vdnVc71GMK+m1QsTxshtWeCmUUrrO+zpTp8Rfy+AsQBnhDfWDu4UrMK32Xpko+Mf
QVUYjNJr5lPBCLBd+8Z/BoTzmmAP8J6q9JPLqKg5d2WQ/4TSPTKGo9ZXYgWKCrcn
2QJsyeotfbAcqvFFh+d/r2ds1ZK7+NNY0GQ7oq/F97fzSiQEh4Z1eNI14mkV7MK6
7HG/N4p5fSkACQlGkwsVPETJGw+BlPSO3V4aTMLi4+7//vHK5LiZHiNn8FLHBJHr
mo38+mHQAe9zf6Yqua0nvdZ9FuxuWU4sUy91siyF3sjuMiY8Qhh+/FSXzKruZ8oz
MSh1PGLnL5efw/C4gNOKKPqfBPFhVaPTbPbGGGVJqySP6TKe+RpA6mBbA1lnfc6G
U55WLv0/ZvSfdkJmTwXwEUWZPDPXqLiAK4tONbCSJW84g2OL7aS56N93AViPgtmq
HcYY0C/59MIBX3KF4Mle+wJUwDs4dHFD1NPXKbL9RUeCY720ZYc1usWnevbB/1zn
wnhuaoH0Xg2zxteMQ1A6X/mtd1MGEcWLrdJfn/e5oirhqgdP+UroU2d50LYs7tjr
cMfPDG/d6/5EXhr8x7oUTKZc6ACCSwlWFM0MBpfDJvvCN97VVRRc2UxMLEM+cG5P
LDOKtf3R4g7npxmBFW+OVPbnaL+9y6PPBK95uZNs7nKXgU66WQ0zIiMeCwwutNix
ThkWbYKuflMzB7dT/uOGHs2A517CT4W1nhxQ7rVRUvKLnTlhpisIHpPeu2sk9S9x
tn7S8rYWvXNkc1YaF5zdYXA6pMtKPjyQnm8ngnhnFqvpkNV+RwLHs9+BpV+XfMOO
2J9cY1pzjHR4WAInDD+tocRA9ZUGAuRXjSGyQDDpZQ71hM9O/mYINgsaJCWIDBhb
EvFZJZagtRCBaTkKgDBra6hZu8dtbAdZDSJvJslM4F1JDkLh1lUZjAJ+jE0lSEop
R9wnWwOKLTWLQGmVQESZ5n7+UcnEQr4//MqfiJV2cNylCYVMeFTnJ1TEymBXslfX
xz1OiQwnez05jtoDp7hiD6ShSLsPpZXS94kFNT1bsF1iJyoe3Nnx5bKr0l4gOGw1
zLB3T1qoJ30Z32KU9rtCRIIH4Eh+vAffYGWVX1xPbuFVd90OMXOHyVLKsejorsOM
DdefMInAb3qSe8WeqwWMx4uGQ1crtr4iBDoaH1iPeUAzmz7YxWV8e+/fG7AwrKFx
SFZMR2IFXopC+LY4bC4jiLjbZ+xuG6K66ZHlzK3IJp1UZZAI8lvP2JH3w2YYfBa+
t5nJCB7nc+NyedFsy5ioYAYjOXSP/H39wLPtO4uxfWcETk6c6H1vBknbaUB73rRQ
VIElLL7C1oOUDCzRJjZJiRxn4ttWuRlbjxlC6TOmrHM5x2zqdE0GxkFAz4SqLu9m
/nvCPJddf2OGmwqTPXQX2HM2Za6ZFtbbypD21Jom53ury5Mtn3wnuZ1L5Ij3tCeZ
nrjF6Dh8n8u8ufq8SgWtf3rMnlARoi5SOjVWdNNwFuxz6dXfH102/9KPgDTo4R9D
sSTN74SGd58AIYxZHQresnUdGDj/aANUa9tOyMFQwoCWALVKmRqwjxDWb1tybk7U
wpToqfb/f9B2ZFnNxk2ZRT405V5xbvCi+5bk/OtfUETWO/bHY5yvHfmsWY6zi+eS
V0F9NAS8FteN7NObxhmB4DgtfQfMzs1blvIZRENiD9DG+yLQpIN5CYqqtT++z17k
xDa1dTNiua7XqrAuT9OHLkWogE7DUiEsWYZ7W1luyW1gGOw+5OWmrXoYZeu9rPh8
XNz5VUWl3if4mXVXaj8XkBBdVjDqm6J5YF5Q0c8RioJZ/cwXP1LcBO0ZS5VbTAbv
oDuGZiV2REnRGFHwpLJBrA6bscpV5jx1iXH2f+EikXkbFFEtk/ciX+fP65hEWKmt
iKll8xm6dt3LzMU1myToEwHIUrYLAy22/IS7iWCdp/l2qvVkd1zMgx/2PEo+G0fS
jqKdhBKu/DnqTfPcOjSfVARyiTKUMRl+77nou/ovTJqxw63VgBdL5C3XzIyVPsPj
7irXZbcfEs0zkRn9A5Aqx1t4h5mIX57FGp9Jru35tSbfhEy0xhdluujXg46r5iQB
K0BFF/zbH5qRKZzYeGjMkDgK/ABdqc+wpNoFIWtd+CMrwGufEWK0Y3TY1qmSGsZ+
2bX4afZk8AI4cIBMyn8+3yRYNWfNs85XUXPBCfmog7eh8346LQ0iu8pbsQ3VLbph
5MsbsylpgW4EiXrP3XCxVQU9jp3bhXWYf4Pcu0pfNnB1nLiBX7HF7pkaJQtpPSJ+
VW97b7CwXlrOFltqfgkB5Z2ewZOcfjrpvogYLAKXX/qYZdUbe3n6pAgZJinAFNG0
1xIdoYflScOvvmJu8un4inNt/SV/UR9AN6fbxL9E5ZzOETjrqyOBVmXcydLr8PD2
24g0ias7kL3HI9ocRo2shwZUgzrW9GLSyrYChFaT2aby9DLIhQ4cru3menIKrcyp
w5rdCjTzPE1EaA8P/NBS+V96eSdyWndpHIorx8N4j60u6kuLapQnWpUeTENDjkVX
o4p6jhl2DcCgrKR4DN2yIulLabnJL/7ECnb1HENSy9zx890edu5fseV/TZAz+nTJ
BsFEICvMLbITrGS6fwK2w4t3KI4zfnYrp7+zB9oMHw0ww9+Mv0X5b+JKv6z3ahTv
oRl/pE50KsBt053I01MUEfTt2mVEUBbYqWeYOHVwWQjKE+R2nh+iM5dV/NVkxuXI
aYxp6jer5LF1SdBPL7eq4wUghiw6STvsuJuUsNrJijuQlB/nVYeeQ5p/0pyj7mHO
nz/ARPcRdAg8Fct/OQlNIsOdZlqUYibMzF+wiAjohrajWc7n9DH8aRf+mYPpGYVu
+sUa4er++s+le0MzHItT8nF7a2OzoKB8Dmwit6RyuYlzESvJrunStakYYZst0xUK
GvJEkLfV6dnMT3kZ4yHBwI835AzNzCqiikxNEcwole/JmArwl2qgz86wPDtWfhfI
o3RJuwX/xMqOjQKQkoBrWKdllQyhK/pxYfwRs/M82hiA6q1lihVoL5DstEt568CR
MiUqNdelEvsUVDOKKHTv8KegrZbOvdjrMOOcbPNiFEFTBuj4ywg+dOso1B//A+PB
/ByytdPRflRjgy2Y9t6zMpY+pOKB0A58lJsmT4ckCVXN54muwYT6l12k1Q5Ym2K6
qzLmjyIJ6En56WDEOLXl6boUs7Zz93af1xd5bVQ46e3ONTY+ob8x/pkdQtN2V/Sw
BNf5+/xLIWlOP4RuTmnV5IVi6nOrnZCG2ilR2jZPbSirVap+c/DEQ5lMfhkD7fg6
aJaSiFnk4gxAxl0z3DKBnBxcTY4UcqAI8KwiqTT9tstk57NL3/PBeJfjN9QrTs5K
kqEUw+cV2fBQ0hM3k/m+swCvaAwMH/PGUlWXjL43QZrZJNlJlq1QXpG6LK3UoWrE
7HPoXK72+e1gjD156oDG4ohOj3WcCJ1SwwNDG1bMhboD8YlNu/F+fk/Lt2m13jvT
HZojRG8OBh/QVP4ScG3/9k7xqT9pTJTAugfD0VGKuE3Fqned0slrs55+OO0V1mVW
cOScGsJhdTG5LFfSI99Irx608qdINci0queiDVXGdGHRL0tzSE42ZQm6rbSYHBK8
Z14YOVtUPRIIvzC4YIeS7v9Z4hz4wHvo8cWSybGWIqnEjo7DNljathgZYiPrvpcA
BPyA+OT59s0d7ajkdWVi4Zm8l8E5b1pWKmMOIwTPibbigLM+qyJ2H+EQ+5G9nwU2
8MBuAT4jtQCq8IQoAuB5X3jbU8uFSBKL00aIDevB9xRaP7VEfjhUDBTXJLpAQ1S8
dZi5J+EZ3XNBTfOfP9h7x1tyHTR6uv5EMoE7HrxS4/rq/8DcuinXQNEN9110l5RF
KUlTBqSJcO8iy2iNxEjUSXFEpLQWxbYg/aQLeKyTsBXG/aFOv3dHu4Q0qznWlIua
+Jc5oQJrNDXfpAtQGIvP79rY+SiO41JvPtOKurE9SJK88aM4hkH6Hcmk/ez8k2a5
lfXwv+k3H7QdfeMZil8jIWF+cGmTkQ0NKAVu8fX+LvgPkF+aQ7wtuNepCogNGfJY
EU7cp8ab95xzsolYh1fFz66p2I5dYzI58AwqgZ3dK3PzXjmUfS1XyVi27KufZvYd
IswYhiu0O8zM400fPZdJHA5F3J9oN7AznspMhQ84UqUpEFQyCRMRV49TXIJ26Ktx
T6RWoM3tZCUKbmMWUvMu4qewB8VPzyr9d3O0dNVyOpTCAGOOheObUxpufOHaDxfM
jQQAulyaeflsOyr6OfayEaKUMoK5NN0/KdbIwPM7kB/IM5qQu7n9zkbSC4xRBew6
Xup/eluvtP1cjTyAkkUk6MoFe2rTa5nKi1Lt1Vk9hVJpHterEMNXfHk6UYV7F1JN
z2+Xug4tVcdTdZKtHaPS4Bnax22TcnuQ47OuQlTWvU6hmcwIbdRJuxBLCiUYvP71
zmsggPUPKcJ08CCXIUeEl+3zdLFivXn+EYk1RX7gfhiVVHHFjDMrKqOtHfaXDSct
vyIufvzIAvck4I5FpFAt1ZJizfFrE0wnkgR7OpIQvKZYR5dlHJjhA7v2j0K1gBM7
6L2F4MS+zKkMIafU1QVcsre0EBk019X3Qk1KZt8Vz8AlAdqV5stK79PAdYKN++fj
MNPGsf02SnwNv7JrPM3qnlDd30/FyaHMSVXOBENKVmqyCadkb0zFmD9sDOkXWoKN
nrbqY2eTdqZmaJN1EEd+gmX8gveRy4uSGhgSov016aAmT++TW+LLtgDhI5m3akce
PsJfLN6utCYH0l/G2lcwULrqKVn8mIrVc1VdhBwLHuSe+ZjhGvLhXrGttL6Ylipq
KEvR8tjW2YhW/QX+oVKtUo7F3gd8gujMo+B9EdIPDUXVWUJWxPnIv7kPz+yRlC9J
CBSJ89VPqU5WayjRqDuLDKgCJxQvd70jLBZ0mvHHfpfLyiEOJiwpmSwFucA5+/7M
JjWcZ2xrQDwHy4OXk8+BJuDL1KkRboiPeEYSdabZOUrwGUm81gn/G02XieyDCBJb
XXF/TWrvnthEq1RFn3xz13Z9tLHL+J0CLhakqSaWch3KXLfBrZ2UbtXuFONVfM2O
VMLgR8+r/CDDoJk4pYJsA5G5+OYZ5XNd8wlquPx4P7bsfpw2P14Dy3UtzWwM4jhc
6pQ3MHIqgN4BhYs+rjdYBA/rnz4zN8K8gCKo6jMYaisRF5niFnc/YDXBMwQacdKJ
rIW7ieh9VSs2U3pBVEbU84qMA9Rl3TWFNh/mydjtao5WxmpZn4lNeWyOsMX4ZYpG
3nGSpI6268UjS8gi8drqu0von1arQDATxPR9eyFIUS+vUi/pM4bW6pxT1kYoTB31
C6uR774FnSkyR+tRRM7rmaMZyNh+e8GfX7q7NhVVrn1ujWVUD0IJSd9m0r9axANl
PAo7Irro6W1sO/DCZl/tHcYBn7RaiTONOByLuIMYZnIw0i/78++4gSXUYSx8j9Xs
7JcWkcNTY/7eAqSKUTsKcmvwiqvLyh1G2n36e/JOheeBChoQTQyoXAkdUalUlwhI
2DbSM2Yhg6d40g9KWALki3tnqkCtUljFb4so/hGgbGQgwlDsxg1ss8O5VQ2gxoAt
Xb31U4szYhHRQfDFhTUbQNmYf/CCaLLPzaI5N4NzYGaAKIme/wJRyLLKAU6CuB74
WvkyKUUfYr34NliBF4mlfw6CuFmbtpSo+Wk/D47aCK3DTz1kPFAQPy3Rj0hDt7iC
iWL0MtRifo7oDqrfkUdKlnjJHY8rIrFAfDyi/GiaXCtA57zd41rQW019RQwr+IDX
g6GpMpOpLROPUN1WaGvFWG/DzYiuQdlR3vDftYAmAtwD81IofFmASOxUoC6cExru
rhIHm4OYs65Kod6obt+KatG3N2Jr8YNMLl6lPBdSHvfpDjJVoAwQDlwYn/pUtPXG
mORgN/EnSaTLd9OyBgxqfr+F0uTMvDK9odFcuoUPtlDoGfqXD7srU/MSTW3Dpd9Q
3ml392OTNYtbXCU3cbbftFdCY84/VjbHoe8vi+8bQbneLT0ukL5c5aY6II+D9UDH
QqhRZ+sZR9R0m7QMKSw421wmw5FuFKB0HhX55ayBf8//8lzJhkJUnhb/RHCdU7wS
/E6ldGjUFij+muA59FmHnoBOdSHv9b7+NegFb4ow1kk189NtDO/+hH35Z1+WsjsB
HDfjPxISy2qMU+SJW5dhlw9k441hP2C8UCjGKj3eGGmeF8MM1JQpCMw+d19XfmHK
qXQSdu0/d0aVCixYZp3Q+53K2Mtg5lcTFz76a7mV7s/z12CvOYDL/SUslfKjlv2J
9Hjknk7rGgnzh2tuAy+rso9frW+p2+f13k0OVReoZuoLDI3HOXqzR+il9RLpjIXk
lkAKrFVRkj3OY+g5CP022joMYv+XbvhbHDAYXq+FLivlL4lRHd33JtKDCPsThgv4
mFiJgwZjwuUDCHVQjXYK0el2lr+o9f8dNiB9ihmZ4ovQ46AUd5CItH8L/RIfgbt1
g+iXuelWCDO3/jqmiTxfpf9QsmNnmd29BQTDeI2hY/u0PCyFWEROMhRg9gVJGeTy
XreobeP9dW5KtLi0Y6U99LdWIi5CGeAkLt0n90zhGMb4y2eI7FS3sAlF0uoxbPK9
PG64LVzODptSvzNj5NlKP0FjdJeZXFD2yceDGTl4122IZOQGOr+Kl8UbgOH6ZS+U
8U5S97pi07H+8dZmGsbYOqv411gJ2rsEhBtseQ81MC3+deu6ZcdQLQ9z6jmLlmwJ
niIEzaKTp386sab54dF7unn3AhF3a5WbgknPbmOE0oGE92lfWc3zo0j3UVVqk2ws
70pIi+AW2hcssEk/uoHN8Okm0mcPlhxiy9t8RaEAo85Y2SdVk/HmUZZwLUumUjgO
VcKzc0OSsjZt1J/V5tfTixGrKtnP+jaauLdqyZOlqGr5x60MdoPUZeDmV+WlAaCf
NIZ42AhP5Tc65PcFDQNCZE+gFM5x1VnU9sfup5DsRdYppmw0rf5VTy5KDRurbogp
xFZczMK0F2150v/1TwDCjMrI10iUMjKNYRLcuJ2VeH4SpPhwN33NjcG+cOhI6eSM
PaLl1DjLRkBDMjIwzTGQqr6zAzWc8OeeBSTZmzSl9XskUPsQ1QSXf1cMd78HHqYW
YiJ+rVeEeHmPn1olA/SrwS9d+nmCXSzo2Z4uR9L5j5EOE3t2ZOnCQZrSAB1Rt51w
+KqHDNNzwh+3AEQHORWP1iFw04lnQ9Hmnz/fef3OdCBxcHRcnuA3D/pQIM6e6S2s
quHDd8Q+s7rTa1V3wpHeyx8SSGPELDN4qTHBcVYZxFrVcYsB4fJY+6SCGuWYKk88
bBblpjFOb/Z6AVCiCv4FcgUi/28LpCObxtFpVD9CS5tabH2j9xi2I1gaFTdAV54A
Dx0ZRenNS/cpuB/YYwSTta1lfF7KruUPRrSLJ26ceK2hlMacry2uWXtvrPjVMpbs
fD6jTgxjlshoQeVZzE4S4hfVzLKKF8fyxYhSnic0j5mrUClx87oCrmcE3fvQ/XXA
dpMtRn71u1gD40m+41aULqTFc2C/hFKiv1URvjFX12XZyoG24AFXSd5QbqoSVC6C
x9Qc1vhwkz7RON4ikU1gZyQc1idlG9LhRVK/XShOPiI8AyDz2aSqDdxVh3QMv1uh
NhahMsqMvqgWLQg3jSqerefHOQ9kz4ZtmYPBqkAxjS87aQ+rISwk2cKr5hUWMl98
wwXNVJ0+LyNYd2e/iV/GRDKAsMOQAUtImHTW/XOTZgpr4Pb0uJxS9xjEt0H2oV3H
rMXF1cZvFdbwev415iuK3ux6jtAOY88xIW17LwNQJQzdJw2n0jirIFKeComoo4CY
vFxxKCtAgfVa0XiYZh1QaL//1IpY11ZA1sRAlYTxISHxEyJBOdzoGsZGloU9Jx37
CAA8y/G/QeDkCOjKToVJwT5Am3BS2iPbnYrYn0oWKm6xxEwuTOrW0K5+8h1xg9rm
nOnK/DhKlampJN4AMAZfL4ltZ1iaXNg3Db5A8sIqaIdLqb6o+CbrT+H+ZN7JLMYX
THPESHAc6usXp30v2rv8KJ5NrRZWcCkNwnKuPf0rFsysUD+vMAel0kvJTifprYId
j0/tKcodLzSB0d+AY3CVHCskTrXDGITRu6Nc6+dKhfhKJBJUgzh3jay9Tp73wewm
TwN0dBREVSk0SJXxLXwzUMKkqxvaWODe02RSFM4/7HzIYLL0PeEs/kvEZTx5Mi3Q
bglYTDM49nSTryCBANxBlKL3W/yg9f0PU5wgyywk3HKSl7cvfC9mzxkqnmhdt3mx
8OROr5cVCaWwvhVKVUtpB7XwsO+Db7wBzJ4+/b8FDEaHzX+YlZtlbvaqF0L9zxIY
aFtcz8ZdsObWcN1kmieH9tdYkI7pY3OSTVTCqPJQdatDNhgBuFwW2gMOqF3v4z+e
IiB5M2zvO5wX2c94UtwbZQo6xN+1RQliTP6Jqow1Tsln9jMBg/39SHkIy98SZepo
WOkCi+EybEcf/GnFnUEZbRGFxOtDtF7/blE6UJTv8SGfoVqFrTinIYv7rJ2He70w
tYZIb8K5xJuwJ3OdzqcCEgSP+AtNI51qMHr/PMzVPGFqTjcratT/XPtj5EKFijX0
PyEO1SiFdAM2cNJkN9wyjpWLnmZdINLZ4++SBUcwQJXXzQtl9YRsysUsz/BARcST
IekiCkfOvKstVDcZhAbjWQVJsFiTdCTJiMVKTMSypxP69ccdy6fFmvpVlf/nDMd1
vwROS+zGloRR9T+YVfE8plXsnhf3PZkEDI/lewJuFnoMuFK+aaaMPyP/Ro4VKwyX
MqoL0qZhCyhRy4CjIDbCAHyEHFxz2OKxKMy52SXAqevFn8BRG10caq4TARIZm7By
S9JJ0eyY1Ts0rOtYA0gavjKZO4wpvNDr6b3rPAf5G0ZXAcnuf8Ert9pVpng6/tX1
JyYq5nh4xR58HkOnZ1J/p73zgMyowrE1nClB0hdWR28KbQXtkerl7wSWIuTcPmis
N5NTjcGTp3p2rGGScPxcchREe7ttjsgeH603MShEjkVXlRt8GqGEES+qh8HrJtXp
0IXkfUQIx8+ni9MsXzRc9fuHXez751aS9TdwpW/cOxwn52tEPBHxjO/P+b9QrrX7
ecq3FXoBMERMlok6sPyczxBTHb2DC+fdMkuxx/YrpI33YH0NKpvLRWO6E3brmBgf
arzSixuLPlhOPuLYkHjgvf1SrDI7Bojh7q73SBZjKiByLIM4VO8TpWyGSJAt15Kf
zwvLsav6SJUvhGd3L3JNt5SyZsJMb7SY7Js9jWeir6PlRjfP9ELEOZwcEVlcrzVm
7y17IaDGvGxRkmGdWAHaINW1CsAiQzm3YyOSLY6CdIDo6zgD+DOoKlr/suDlcKmj
v4apbp/9cRLyRIYPANyxmY6E8/duTN4f7CWhePaY/7Vtk6Lx/2jGb/+zKExPzkbZ
T/vbZUDgj0pI5s5qIBkTYnlMXjcLzWRVeFgggN7cN4u04DlrMJlL2aUbHqgeV3sj
xmZy5LIVRAyi59pPh8DKF9eMJu5xBK8SmY9GhSPQc9NdhBoXp1S+ZkqZltMbOeB0
aG13MRqCZPpnS3CI1QzoVY1dsNc0kbduTNboZGnAPNCkiyfWVm8vkGpllO2KfwSm
PQMHSiMk82D2JbQc7ExhqWrKqlYcIPiiK2JjtXLNxWBHFLwfFTt4o/aKiFe3RwQ3
ruTohE8Pb7/izrU4ZC1VwYjlJPdyOTXBNDHfT0GFGOuB660Adbo07pcQ6E8mkV6l
yEJJKm7U2jnGbO+76u6K3k3jEg4NcoBYfVMe/+j8l0FxpNvCdFs48fdE2slFA+4+
wOGYVWxBmVnEeb0pmJfYNaCGuIV2W/RtQh+B28vBqrdF01rC5MFbPBk8+Oo7FE//
/O9h8gDjXtXTdP5Ny59NCJp0PRv3xikJQg+5N7ka88FaK9ukFy49J1NwVWEDesuf
suxZ5sNlMNsj8YS6CvLVydSE5hVLMAqq07JCEEbSw/RodERdGFPfqUuFDYATYFIt
X53WG+XLIWr9unGhNOTqWBbaoF5twn7rNAaEW6w0FME9heMz1WZVWt5FqBxBNvzZ
pqYvApEY8ZNcqIzbP5FstW82nXPEAB2Ogh3lQZ28HRabYc41aOzuf0VfTDyGCvkY
smFbMAH7kvg6ud4MoMcuQYHP0d/uzi+4QPf7zPKWAVrX3vLdjN9Pwl44nw7tVobd
oHlrgot41s2od8uhEMyE97k7a2wxHYgg8AveYwuGqSsCFGV4fWvhmM1jEB/Owr9J
aN5/65jaD/InT+eP4znCeGTzkTTGMlCfUP4UwvfjbQglZaJ+HEk2NRNTs4o3w2a0
4IO/JQMWd27z9ljO8TW4GQm6aBgJOy4dc6QHsFsrCOVP6RhiIg6zcPZrltHwCx9+
Hem/tc5jhPIj3QKwuSH/kK98RB4MQgG86WDsnHRpjk5JRnp2zzP+Jgjn1FC+aAG2
TqJ4Fpqle6ZliPixIKVmr/nlqXUs6aWO15vBiFoLqaHUN2VUVgBWk5nKg9wBOxyr
fmrz9nucf0jKG92Aut2ahpC2ZL+oBjjqXQ0F/bH3GmBh37f++arbnCIt+/85bpJj
mz4um7JsfSi0FArLd3rEvzTtGiOcrvS2edsYuqngEHUJlZUQBnelxDByOfoABrki
QK6srFKqCC+SXtdU7IXQSNFTrVy4cC21xYLyij+aYdrxESbYJCiMQ33Yk1/5gTcr
Qxr99c5UM6eA6lI4zoa1fvfQh98dHRpU+f3ev41ENKtUr1Fw/FJ1WmSoMirX6l2d
xsthKqtxndO4YZoJ2O2n98hesCeikk5RxoWgd9XBS3opqg45nsCnEvhlBAv2IPzJ
ir0sv7dzjuDuz565fE08iqstAi9eKTrDjg9/cAMsmA+SPqt7S53lL4NN9OggGGuI
AutrEyAN5n8npEt2yjshHFR3FsHW7jVPqy1Nf7yK8Q+qkNY1/OyUb4xygiCeI/w8
oDqwWENUsCo/RLVgOH4CV3bp1g6pCsrRtLAAabEKqBhJhG1v2p0Q0MD1oejL3fCg
aED3nsIyZwUw99QbxnWHSxYKsYk8if2/v+1SW5u3A6Wz7qOFg/DPCP1MjDJLcIaE
70u7wx2za4VXgDuVSsCf9kNqrVuF8cYg8C7sR5HS9CCIt58l1/e5flb1QJzDdnRy
IPtnkFcudmSdSaCvSEv17tRxshoZT16KZg5kWSyQUx4XQ6E9DbSBmD2I1TEtpU6d
y0PZgysKzWj3ErRtegV5EXRkhu4YA6LwAux5ouzwuksApq6Z14/LC9o1Wrp5mWIc
SJ0nSIkQazZVS0x6k7vThgfqxMKx/jE/gopM3h6fHLYH+j5Q0AKXnUzjIfvGkyN4
NME7D2vz8NZicQELnD8kBFyvK8MnMpWcTeyDKTZLM93Npju1FEUuI+bO/xbfucn3
MvFylA07NBWINklSDhvy6UxkJ04wsR+ON1qTdzW9IkbINx+mSIShU8nRNhAJudUn
FZ9UE6vRSkl7703s8z/5cxKhu76PFMd6mSufWAYz8wyAomcec5zSWc3VC4aPhJJF
KO83lhvDZARhv3Hlxy5SUHOtYwWhjVNOiTtKvWg6v72j4g6evEg9+IoWHnJYQdtM
Gbt8XrVXc72DDTSa/pEKUPZiI++XQ+EgjXg9WWbkqlG6ZJjU9eb6+1uDgDQTtJWC
BvF4n2jQg5sXlIJg8JF8niuiYOvst75KvyKNkOq0+z3cSq+ie4/PNHquJsoQq/Gl
aPnBRw9jV4O0rduYdRcxxkLTbYe0qX5L9lpYoaGP7YdtVHsADSrHWhXmdNt93zg6
Yud/9NRbkXApj3md242ALc2alstmOzdJcI52uFiM4XF5PMWb5zP04GWalPcbSW9j
HVFL2q8QBkXsJofAAltDrDatk8ww64ORx9cmZWfPIPeHVI7bZwMLYonYNefOIuQP
dx8RauxHDC5JxxdjSQl+EE8etx49d9+U9NuZ20v7U1BrV1YIl5gaHLLAm71VXPG0
oP1KysrC3TxW71kuhqOoZat+YJd1BS1cepCzcNr+q2fAMl06fUsyvK35hRMncBJB
Motid44Bf/8aj9ThCRJ5e/PHd8xGmuLrOzsYV4bdDnMdeHI5/jGgkHoG5L2uI6HY
0rIdU27wXgw0cRzPy1K7a1XbtQXyIjgOvl7eRx4K0KDD3XK2qSXQiHJkuMtpzpit
Jotoh3rZHK2Ci/0bGBGJpr+iRHycaaJYyADD0j12wh3PlbvonwwVn4KmAxBbr2D0
iCJWoi/x1zDqRe94Wf0UZx27Yhv/7ww/0q+qkPzDCgHDvj8k8VEWUQVl1Mi7f4sz
dUtFsmgqBSA5qXXzLFukT1GX8ld+7ZWwwyh2d6nza5KgORD9zGGJ9dSICATWfhjx
havtVNsuvDkca0o0FS0mtU17RqKw7DTIgrbAdI3BeKmf9PtgXxA/2FuAngDr2gDE
jpE8uNPjCdm/BoorAjW0kqIb45FAjQp/kg2aDq003Uq8JngqaUcRam86Lp3tMYwQ
NJgfQp4yTtEmYEidbWfnctuRNy3kzwvui2w//EC/nRsmd+9xmECC5+MsLnHQemUj
CbR3cF9NC4GnfeBwWVUfLkXLblxRStyp2zh1EebiVSbYh1B9mPhXo3q5EREwc/Xw
yYCwJrcAnsm6RSeqjJV2y2DahejYLRtrCPq5/orFS18vBQt2fUsfir0NxGj7xnOw
54yFzl9dX2EPMrtlL9bylcajk2CJoGAvb6Lf3R1jDfShCNG3YSKW+WrNpdb77R10
rFtw9jJLRtkk8HvcUPTZNgYlvW2nU6z28YdgslIvH98uW8zF5GNlwm+C6JXdRuWD
pwEUO8UosWWcg91MOynnIEDrsQH+0ZblXBZlmnz6r2lzk5mA6sFqIl8Kxsu4Wvnz
wgQ37Ybz9/+SFi4zU3qpBgenHlSBe/hqpkwM4f88VAZplP8rWuqq2yuUN24z5TDx
Ugih9n4MeZwYD9iz5avF83opQ/Zie3NY020JgtU19Z/BcxCmn/nYQpCad1+M4Ptv
sE+W+gI1F0mNmsFXtaaPhS4R1QEyJ5LNYuIbZQR861dvKZ8p3P17XpvZXmnlWJ0p
q7SLdD3GsYbvuc0e53Br0zwmf5O0cpQKwcniBJ/z7VlxSzXTQShJMiNJqhKYmFd3
m2+sMoLvXZT4mzPVfi9Rxx+1z3w1jBCe32XJFHUtO3gIUVjHBJzUZ9IyT2V+op+B
Y5DeuK0SsIHmdrMdAuYAPNn80wi4JiwGj9D0X+UuNtWI5qF1R/POSZ6pMftCddJy
lOK91AhkBlvLgEXMaZ+mfHkkkPc/HMhiBhqRmWuHl1ZsX750gAdvEKIHmABeD5gx
lvFKzi3rLRvBG6e/LVEhKguVJFyCgO2vvi8AfoEb3n+cbiFzXK+xPw5NYkRELu8Q
T/sl+AGu6bJz3qKkmavrNPubFhk7SMGqIxZOB7LptVHPrpt/Igw22Q3pWhHnI9YJ
/csuKjHkcr9MvqEo4l4A8NJT6R1Q3W8TkUDZWZt2rFVINhxASqXFYXbfWxdx+gnW
Byt5gkn9rS+5zCq1PCCtmCHXug2d1AYQv19b9ADGenOD4e5xezkbkFdD1t62cmyA
xyGyzKktDUJw6fhMRsYIsQbVqnoivUgS3Vph9ZF/ZWVxLF7PAKXg4tq7AFfro3so
nMmUOLUkHz9KNVnnrkV9tr5BHioTmfUpwJf6njMXrd1B98ImmIwOe10bRjtUJmJi
Y7FFS1jQrXTDltKD6moGMQds5gcbkPz3tb6l7CFlJOJuWBUIbcpaPVXMC6MZVQNf
fqtLygdZ+79YO5T4CYBOaSdQOY2r6itULm7vD4w+wxPU19pzsKcEHhVbCz7WIV24
pE+LqGWgvgcbKCocq1Mdn8ZgV+tONhqPiFLzZhMEYR9OF3fAMXTU7Ltm+p1aFkB3
uNrSazpAhNLgZUR2Gf0g+yiUNZ9RWuXZjo5/XWoayfun6g4xEZMO1AyoaLESSZEC
N1TvlcyW6uxwo8ptg4MiKWMQXfi99ar/DH3fYbjlrwps/4u1ZYWBDzcQQoSJrDHM
rUAWknJP0L7Y08qoLxm7X2njZjR9x2ucjh3rN1AwuKhBwn5SL/S0iwWIvqiUFjmD
1KbIru7NGRZxvbkyzqdAlwxNObvhNRVmhOKtSDwJGFIEvJVnPwKWHxbZhj7J4n3M
756ywm6o6TlpLYwfyu92LaRPOSuIzsg4lhhJJAF8Qb01SgR+NfrLn8OkvaJTT5YC
sHdqVWYfGqV+EjyuiaB5ukbbNpvj6S2G/KP/p1udmkatIQZx1yvndqbl5Jt50kot
tuR33ZUZ+gw/Ey14fgoO+NXqeYL0MWVo5w+k+cObsUfrisf/jwlMtEVffaEUuO+d
9U/w9rzuFM2Ic96wgwUS7C8NEeicuQUccKaHx7zW0aw1NSOddLxvgqUe0bs9M1ro
T5d2s0mhG92F/SKtBZlUNuYUnWvPQa+FCfupy2t7mIO7LaGf4TNZgoajAEeRiFK0
vaXusOBY5BmsG+2RxyGtom9YnC/gW8DjcR2CB1JsoV9Q3GGjoqdo0AQGzUQsneiM
ZC5ICyHcKtfAWFTFwSEhel9BTWD7gP1KwwQm87iCaiFneH+6+oODPK5vrqxSQrf9
8McrYCT+/NlyC1VBL1K4zxHxfuKC1w1oZieOGHjC8T2zg8Ln3OV/ZmDkw0wnoN7U
7LTymjhbMxeJ/R/FVQDBoW73LGT78vGrdEb6gn82YdBbHkaHYrNicqAUf/EEMyCK
aSrElCBtcz8SAzWktmNkUljZipGXZbwhzI2sCyDGLtWF0Wr8ybj/CT19Y7goeh1B
0mAYxujkMf5VdiUL6D48hmcK+r96BNiTYQg65bKVA9ju7mksX1eiBhI4CCSckFdb
9j+NsxSl/3b1m84ITb3R6szCAbqlz8+VmLcGhp6l7sqJL+W1mLqepraM+C3NDOaP
GDvUnsyErgYe8731WYXOIZyaiIWSAi+RNHnRLPCYgbe0CZYgGhbEiyT5GTuH0WKQ
wcX2hKiQIV3ikKSOB3KyAGo7QGyyDHI7pFCFrjqAK98cA3WKN1zWtpCBseK4lRiR
imH5RJ7P8R/grMrKdEH7XsKn8HUZ9eHOwJmeHHUEogCtv3/YJ3w3vc+PChtzsaJ1
pG2IIGyMvPOwH0cyRTRiCyP3LVRYyRiKM27jZ2gDb+9UxBtCdqCIRg5PueD63xEg
Yfxw3JvwoqmXXTfjLiyBkSFjw3ukVEC48PXVxnx5UMRqdVxaJPHi1ygx9I1zV68q
AFVJrN0U2hiPR9vrUgrh3bXTXRkRAUFjKpVAydXE6v2giL/i3iABxenC7PrcsHrY
55Aqa0tbOM9fMOvZ39odxqbC0a+rXdgvqME4DOFd5HkvFDh7BFs9vcHukGS9B9Jt
DiU7lmauMZF3bnUyAdkh8cQ7ffgGHrptKFU6044BWxtZPT60KGXbITc3KcbVkI+l
VTCRmB0kT3Tb5NkmXLqpJnYfJBx8tWy1nrSEI5X6GRsO416K08VnIyPc4lo57MjQ
4to3atyWthvFQYUCpbQit1r/unsjR/upRN0QUZDcl+/8+LbgLAoJPKuvD1MsluGh
RqN1fNHIl0M6AR8AO4zWUCEuNxoskHq1HzC8CUjyhiv8pl9d+FH++4qDrne57Wqr
SpDyPqUHzunKf5AGROTo9trRuYyCjCFMYZVKIXcM7t3mHqj4B/Nfs8nEC/h9Mj2C
2Y/y25H9pgyZLeQfsGObAUzKLzwHOBW9g4n9botVltkPaxZoe0WX8JL8nw7zJqSH
sw05hDzkpq4YZJPzYFx6AY6LxH5g9FTqlo2zS5ovXTQBelsq1sxBIgRTSm/6pVw4
tBWEeRDgIaiFVWd44xRdPEiwYkOKLTdwLWl2LRHY2qPWujpinJ7oW+dQI/wnXhsJ
oRg5Mv0IMfOGZGWxycopDTvJh7t6zFM+vGpGCsaqCc1zRZ69d3QxCOVt+ZEPWcht
DIqwau+yxT8o+/DV+My55wYThJh3Y0gv8LEJ8OsF0KlPzX0JHi0kgLg08Nx6F6ZP
fllGkj2oE0+UEeG4v97rkIwznVXQNu2ONXPWGgrO46ZO+QygyOfH4RVOB9YcNfSR
N5Iq7O+7an82xn5pPgk7SDI7lQUpmR/9eD/A+yzBzyyldSLiy12uE5EVkCHpyLcO
yEzgO0esCtOHW90Z9cYLx5DN+lE5xgVlXcmGL+Ey0drpxE/vUoqTF8jnXZeZVNQ+
yuOIzWoTi94x5EBfrfKUnRuhtA46JF+v4AOC9PWFKbt/YwtrvR2dVJ43D1t1+W1H
dXTgjyUrKrMsxE8fy703utj0qX6u7so7qHs1YI6bQVHFO8Z6H3nm8TJjizyosQ+g
yYY5dnGAnxixNVuRpVlPfno//bTSx5ITPWE8/lYtA83IS6ImcAv/67fTDqawMep9
A6JsUsjtF0gh9kQbdOHPhXxMuYKwklf+f7waamKRmBlwtWqSwfJk3SajPLLi2iVY
a9Iz6NCFWxflCZROvCOWq48b1xcugIAy8y6658+4pPvsLQ4JgpvvUGbXEXQCJkag
PquQrCQWI6TGVqfG8wTKhGztO04tbRWj4MY5TenWncEIRUMuVRCS4y0nRir4SYt3
S9yFYLOF+DOrqgHeLauflSBbTwlGq96IedO8rfw2om0HiqVEirKnxLMCsWRtOiH9
cp4DxJaVD5a4n53c2D+dssGULfcEDMjkTqm8xOtXE+NqWbVU0LthegZU17MCFB05
EgO7rSJTtI/7WO9PIGyffBTFeXdpExRXAd2KTZBl+n03rZ5d97fjSVvc03INusDT
9pyppAOaIDs4Num+r+C0Sm1x+UGNlgc8aaaTOzJvcQv1WSVkLbr63iGYIR4zqQtr
0A4JsJVIvRkMu2E+ta8Eyuk0SILUHbduR9Ahy43zUaT34iFGvJFhWqxSdWcXsh5U
w3nqBcWrLmnCD/JVoLzJT4DS9x5To39yBWk2Epgdxitc8NYUeB1OeC7UTDYUExuq
MkWOoNFYB9aZolQK/9fQpxiiMOJlqDOpX+OS3dHabmsrN19Yl/N80Y6DYbPO0Xt/
L8B9uFlZrvQEaYZyJJwUE+XCcTEm0AwQFLGiXkU2e7B41BKXRYg73RYzDsOYiKaL
6up6XA69/5Y6ig6YdPGd0EQaIaCYZSDW4ajnMWxw1pDp2iKyU2tDP1IcuCi+WnLX
7OC8CQYcgYEJhJRohtKeXs4AijafInYUeH1yMh+7VKjqCJ4pPyb6jn0PokpxJoOr
QDx+Jcjv0e+8lbZE9mmk2Ptz9K69/vmesuwoKQIEeS4AkyudfqOPEv18oxBxfn62
Prp7bn+x5cCw2qp6YIqDc+/xUlzm1HgaAiF/mqSlmVpv4au+5lPCe3pE/X9vuNnp
eZGrL2Yt2tTrMIko0znC7Trs26H8CUHcxUWcRUw0HTZKRltTL3bZoDBdhJqAJVsA
SldXmS0jJN6KySG7ITI9nseydG1+8xzNgGih4ASNjVlpeOD8nHZ/0FX0T4DQMQpj
VTVVUZLjcHt6IkGAZmdWZRKPlGMAgHxv06N4bijgOSp79Pn91FNevERSVF//yKKm
yX8He0jmfTj5dOBgsJ8gQ3iQLs/OuoXLIm2qLDa/ZjRqDREACbbQlWZ29v0SPKP4
khGp6va/pIi/jab4VBlXTJ1VuCfbeEiO3EVUyvR4gdfBRAZRc5CXOWPnlD3+Yr6B
Dpc9ISPjNkGo0nm/qViDEuY4aLzDA9xxoMQFZOMgChzeRUeXu9HEbHjYr2Chi457
P2JxDOpe65i2JsUtF76HD784Jp9hQaP2y8O5dvlYdD5u44b88we4XcusXzyoMtpJ
D9JPCa48wmOnlmAj4M10pO0MLQYzgJ5eLqMNktdtPGfsyGWriw1EZpxdZq1Wp+qX
6MyAXFxvQKNRutQJfD301NTQNpM1cETha7oN11u+UvmkYpyOcMvltUHaHAs4xkOZ
zqmpgNmagd0uU8Gn3EUJJDjPpIPtFU33NMxx7mbgQLK5Ph6v0LT1yvUyq85BcXGE
uHnuf1lT+nS9jMYJhdcN32W6KmRDOwgRqSg3ju35Sw8n64rYrOkTPGdvd4eoXlmh
2oFkRB7V8fM0XJN6OKxJ5cAgrRc/8mxBU578uOMTl2aj1MPbwdmu72qX2a3op1Bg
B6oP2ZzcRU6MFOTxT9FD16UgB9a+I5zB6+ZDP1Xp0e/2gHd/FWsgTpa0pjIbVhsm
eh/Mtz5oXHuLnnLfsz4KiDTXWhZWuf4jcItNhqikmAJMnZSVIpdk+Dy8Ahf+T1lF
o7amKPfYe/LGjq98cZsHSnZdqb/l0g9GYqt9N+DI2k7uh9UE8n41IQMDey2lZddA
JDtZdYCMVJSerErooAsLBI5qKKjrBwo2uuGk8HsI+gmevCG5/K9ZT/ZGmrI62Utm
EQEApvSwXRLYDgutRkDrSa1hjTFAnh+WCQL0fljgH/TdTZcWXN+7SXkYJAC/scVn
4BVrkwzqN9O9DT+h288wmh2MHo8NsoVL23B/Nmib54vZbnt40aI8ajC/SXRD3ink
S9oIWkKGY3PSKoaVVH3O/EAj1ng3KwFSTIAPjobAYmbh/5UWtlcZIj10Uxa+zLSi
rLrL9J5BnSRTq4RFf0KbVfIYps5zI+Ib4YIYBF9PKgIPbIot+WaRTzeLhcYN+90y
NHxRwK4H3uGen4WimjcyOK9isXdlTf+7zpAe6l+6bJubPSCZv/Z3nTanVSzgxfO6
RaKS40oRUtxv1PTZAMzpkA7Vw/1e/GoDEyIfX5vOe6gJcfo0oRys13egLvLyPuEe
xAAYclGs4nFFzVE5TdiB+5KFsE2J8/gzWQMid+xwkTpIyCghQn22BLd9bOWIiHLT
uag6aDiUViXBKkzh1zUT8rn2Z3yN9j2B9rpip9LArGBkCc4amBEYN3C69fwRLUKt
PyzZ0puq6IORr+cr1EfA6eWUKP3ipRh5UrvQYdz6d/F0ZZovX5AoJbWnFXTgjSLX
2i0JeBEBreYhLM7ivchBypjBvn4LKuATZrt0S45u4YQj7sItDMQXKdQZIOICj9Qr
ubZSL+ApVnh856QMiIiDaXWz4KTdKcyYM2jmOz3Wnqaz9xaf4mbmxZORtZ/eZGUM
tWm+hHjdRUHMvhokcsX2V4bg9sU5AB9eKOPRFzqOxX9A1cWE/60GDRMxZjYHvdgc
sF1NnUgNFqOiBhhhO7ZcHy1LNBr4vzTfKzys5cpKFuV46hmAMXszAYu1IS5FK0cX
YgM6Avtcz6TmX21oa8n//oN+qR5zGAWaG+kuSGIh91AOfSCaZmNW4HvW/5lulYMq
MPuR3RmN7fXrrwSCsCCTpm+ilt++/wo/c/LFFnFIQHDvgC8ZE/ZqVIHIlcrB9+5L
Hy8zaydRXak3ypL8WX5vrCgFkLLM2JjmLdSDbDvQOPmwJNvRO1SAkmPyTcc8R3Bj
/VBkEq2T9+ae6YZD+2OCYhVodFErZxjEsbR3xjZSyS1Dg3f37qHAVGaDneXMXTd4
k3kD9xCfD8AA2P6NJclVOki36OlCdl62qH3yD9KO8R0Dm6TAhCulvqddQPyHPX7U
Vd9/WBJx1sPKdwPSdJqReke2n5HXb5zm0hFEe50k5oIeVAtx8OJBNRELJm7Sm1KA
BBgxK3v91g7ZM8/ZScxj6mIozVjzTWIp5wVLcs2sA4VVcaIYzlmtHJQvqnQqEzyg
3ZaIIuipZanYy7X7dl8KumR6cdYegD/iDN4ITQjnAewTlFKPHxDqwOeXCfPSxWOj
FZUHTiSUMQqMt1+DnEfySXJD+o1yQMvs8Zb+BAOOz92DhP2wZD02PaGfH+VlJ2We
O+/Jg8YqpHuVkVUf5CFxrC2PJfcctep5qjelr3Yyp2HFqbfhYWsVc5nnqF1e0HxW
5jKGbw1pRdtoojDvn1H9frmh8U+6TYqepfh36VH0XgKozpNXeywdjwu1PIQVY6Up
C4L3XCm/PpvZAH3TCTez1rBA6Xbi97tCDEDS1R8qiOGDrtolkveVaBcsovBV8VCR
owSEIcW9PgtZMN4qdUK5rajMQIKVdjCQKnpu/fBWtAgTo0du05wWE+54bt9LXqjz
s6PJJR3Lef3DtHFsKYg/eDML++h2zdN6NTNBKL+ti+KOUXHfiZ54ideWxgAsg+3z
kyHe9LLaUjsELwLd7huX2Pp56QkIOQbvu9w2OIVxPJ2/CgJtKuAjyNGG86U8mADT
f9n4Ecj0ketrarLVcZU/IqVyUWXWyzL2mJq/ybsNAPPybnaN2roKx+SBLp063Otw
cLUnT0ynV2msk+RXTn2ax3pbWimt5QpD0iCKHyAhV5Suya/Zbx1cF+tqi7uvitWc
It1aNb3Go5Zue942px9thkbuYg8tMod5kP0ufSh5xrMNFogJjo1RYV6OPhouQw9e
v+QAvwcVMJmONfdrHNsHwwkRNYP0n3SsNT0oy6EYfl3l6f2RoqlzoA6pWmOeZeGR
LxqJk5TxuAOXGVs/WyVd8dcmwn7eingLMtr+pvJcPf60Uo7Q2urLsvFwp0BqDLOK
ujHPAeTsyyravxBWo7vCttcve75/Buqoz0Q+IoZbdQeaUbhm6V0TlnCW5k7qC87p
EUQRfda8YIERD3JrlopLZx+vnc0/ZEYulwD41sx/rCri+IX/8CNOGhysPV31/+aw
Pm179zw1+Tx99kE0AHAcSHfI97I5wNePYuNFddhIZlx01ZDON1t1XaS3GXaSC9kP
gGnyEu8WFbEa90TGsZ/TOXV7fDrwXBveYSmyfy0PFmie0SsaCsg4MAJivPI0ZRrm
f7m6GnQhEt0btqqS/itErO2TbMv54p7W2TMryyE3nlnEckZnKailek4RB6x5hotq
/Hn8cn9ddHRWI0I8Yg0Dxx7fq9ILGtbcPpgCF9mjzU+AwgYH5cFnPn8+NpOzufgO
8QJKeSrxXIuAE0yqSz5zrWXHY1O49BWaSSsWBpEmKg8tOM+r/JIl0LYcayaoHfBC
cGyLXUvkPCP86Gzg3wdHSVUweKZCX3If29Dy9/uH4fQ/JuZJ48gNVsGWjMakCFUq
Cmy0zhNX97FEZIHMIAQF7C4+lrVA2dXYC9oKkW9Fx7IwRI8Yns++cyTM5ZiIyByv
wLynavDN+HJrtUF4IKmD1LSTPoUZrTPp3Yw67n9xHUXNq3iFBtbB6u12yLmkWYU4
t611C6ouSDkObIvAZRqNem30fJ7YHXdVprp7JI5Ja8wk3HgG08/sb2c0nxqJDiJ6
27ezpiwhjY1UiYBcvXT12vecf6KAAmz2upo0kbzNLXPXAhUEpsN94jmDCJvrL+6l
0udoQPOfsvP62INwIBS/V7ZJ1r+BrebTjWfKephZa5EkJAYMyV7w5T6x9gwjTqc8
QKJtwVmtLhcj/VGTD9hWqI8vIbmLNtt6DL9LyxIu0fs32CN1GO2LefQExKokTlaV
CI3IxyuAbHGEgaofHXccFBUzsoABZqKM/fUfAXa+AgYpQSwJVB+9PiogaRqq3iZe
q2a6eBGXSBzVbemWQsKGqliUjaG+GeXccYmuf4MorGBc9hUJy7ZZoZtKEHqsGJYs
bLI1q8XE59dleIH/uivTBcCxkKods3DhBolCqbUCX1axNSHTXFd6AKEOVoi4L3bI
1xilzcukXYK0m4dgV6QQZTe8mGCCOqg5r7e/p4zeNhsIVTW6RxVDSoMaxGRZxNmh
o6MsJzUExIIQyS2MC2wp5xZ9tngB0oTl4P+jWNbi0RzOSQ0o3Nrf+19wzLjH3kLi
n2Upr0TLe4rmmsWOyCGVn0vqMQblQwUQBCjoa2/wjlOwc/0OUkn5SijUrv4V/CgW
nfevRmRbLUncoGpCF1WGTfxm9GzB9po8hJBKZjT0vzz22BAg9qHzZjo4u4XywuHT
vuCdEad5DU39IjzE1efbBy9CwOnVk1PfupCqx1fulqMQNxiSIGL9YTq6jaUK0Wxi
EHTLN1JyC9Y/PiEw8OnWFsZKqeIUwm7JnYhLxXbwbIbLhubRdnOnu97h0bRLyLIj
SZvh6oIL4CrBtEUggMELIB03wyBTL8N0+lMp8vGwq+Jbwv2NwI/PGTQmNhlYI6e+
wu/nkDT1NuHbEPiGVS5jCP1C/PPNNiAGXHSjrlb7NAsATNNvSi0myn11G4iK/kPN
+UdwGABS9PGKUHg7sbTZJAvWWU1Yh0SR3CAT+3NS0NUCGszUSzoD98GRPHBTIBBZ
Zr4e3yfrSNQzAtQHER2moCTps9SPCvimOPOD4kKXKqfc3gfVu25fsy/qmXZ0Yd9z
Ua4Kn48Sp8qaIVeTIEL0rCrt5kC4gABICpKnsR61ON+VrpcvtQKq3HISf73vy6aM
HzOvy8RhvpX/kCCEKremf9axyO9YL9d+/d8ndyMk/1jc1oE+rM9xJghtFJKKq5eu
tQlp2R3N9PGSi9nuucWpdicCLw/SYdMbglwK3M3AFZSQzb/BkDQgQa9wUs61bkU8
U4tzt02VLixuyip4CokWjZwzPP8wyXfCVRDhaXa45ie9U8Y09SYVOWcp90ODmVK/
leZ1jXNjBeYw6f4gku8MzWVyWugb3JbsQyCplyvxy/r/Hc59rUVUcQxo4ecvmGgP
PrikV3RISMKeGibb5I9QalN3nJafnJ1mWZ1uJlTYh0cgBCuti4/TOUr8WmamNbWP
r2QwGF8XCK1PXt7VStaXY8QGbTM1V1BQgUXsvhhsXFbSOIEbhqz/rcUdRFLJBRux
wIleHUcRizEgUCjfeFkshytQLtxD3HvbNyZ5ZMiYhds95Z0mz2BDjMEThLOXWG0Z
Zv4sYovUk8DuFUVw1o1LG86fNzq0brz8de6Pwo/S59Sa9Momqx3XhqGuLTpYXIn7
Rrsn33xjQNYY5GZWpZ1cFJyMpE+N9kiWFRYc1aKUS4OK7ILE9C9Kozlbgu7gNjA6
Bd99ZfiuKiSf18qWCFOkvxGndGHarDCXbYrRmx5/efKWQbhEzoN17l36vQaV7PvE
q/sSfkFQPBV+SDpyZPsun38TTWABPVtsl2FsutggH4tvDCKSEyZS9ulWqz9k3+0l
3kETNcT6lvRbpMgkg0lEdFyuOMuqdnGgW+KiOcEP8ZkthXihRdvRxblHUYiO9afY
mBgEQNW2DCohg3zqkfCU6E9VoSdwOs/DNFWOgnAfcNf6UOSZNilKHrd97o/PGG4j
+EsduzJ+NEXvOP/sW7cbwH4WRNjw2QCZhpfeS8egfRFmHl288gHeX89INtyLbJ/l
PtGNGN+mvhZ/UjgKsbmgH0k+mKwmyR5O3vt15tg4sCGNXl0DACqj1JMI3+GJrCf6
0B8xRkMvGDzs/uh2qjPAT0/0laavWGEvL2W0b1CalO+2+dEOOSGI75erSkC2pSTY
a5cATVWT6PfwA+l5uVFqqZ3ixujk5OOrwKU0juXz8/xah4YbeGKxZ5sZIXwuoqDx
3tBPz1IMhgAU/W4i/7xVc3LpqtXwS5mg9TGHRXUNNDYS179QrQlyroQdi6Ua77QV
l0XvcBwkcgJx4U59kC6okTWc4iFK/zBjG7WBZgM448ph6Mv1LcKPk2I/C1h5x8AP
msHkUduKgxyJ5V3LVOnerhWHBpWXKC3AmSm+Sqcgo5LcdEiTQ6Cg+YCNqc1OWJRu
9a2A4s3KrZvkuj1PK1V6c50QahDWL/fEbx5J+D9W8UlJn9x+ci5gATUEahatNCK+
BujyuVu9+zdVtckkYS7D0sxp8ymrZl6rCVch/0sg8/2a7TVj9miKxPmjWXazEqMQ
jxQBwVJKpsb2V2pHM5orKq7evpUYzNVkU0C7jmIi6zaopG+UBo4+hwTSjASlkWwS
DtEBQjn3JaqeW+ZN7L6fRRsPBl3PwtJZPiXAd5u2/pV+EXRlmSxSZ5ZporCwc8LR
x3u8BGGJRdegR0HJ+A8/THWCu2ONaS+nA5jbRLIqUqlBcmT7HcY8/G8s/aPLwaXj
qqXgoRdsbcmPvL33AgX1xNVXe1Nw66r523VQB3ap8qpD2zCDda/B/6lfrlzmighP
DagcDhyvTeQSFTJc4viYsLpRV7QTSlEYu14Jw0CQbvzS/t2ASAnFXicQ1qufBWVW
5Ogrsfl+R6gPs+7UTdioHijtrRddXRHzNBtGBwNsi7lefOpQUeIlPXxUAlwE+svz
0vLriUaexT24oJvGw6ZtYCREnhVwhbsw752PxHctLby5uYzqUWH5lq27bJxeCrZp
BO2942CfVEUb3ZLQS3fIlQVcaPxLrumRlac+NkLBFaqbRa8sVnJVmd50sxggbO2Q
/MILj+bzNbCy1Vs0dMKykrNVjAjL00gjslmKjUIQSTR5TGR0uTwCWOrRfTi8UdXX
IpX8Er2jPzTBuOtJaJItP9bKkVi2fFlfgYrUv7uSVhEPzHCebulSF7Qu2aspxobd
g8SfvCN/J+Y1ptC5m190tKqnyEDXJJAZehXphUGfz4EDugi56t6Dz10/Rocr2ypF
NgVVFdRAO6hKvG16Sv5rCpoo85oqDb+gL7DajNnE+1dY9tuYtjERdCokWsL/QQuz
CmuY9Gs777CVV/XC0BEJeyNx0Rh4IKxVmKOOnv49UetD5J8e11AE2z3gXiUHh8Gv
ZmgYxXmrvCBZViB8DxJCwnywHwf9o5KDspD+nozxTavuZfzbgmbmrYBt+xin+Jrk
UURG3uCC7ETnp49bcqI//YQ1gqoJTsT/hzt9UYudGBY0yfCORBgPGGJAq52ds62X
ZgUyW2N1hr18wfUZ07/C7XGWLMZKT7+aO2d47eFJEmVbvFZnFUcAeieewZfjV5KK
gLqhGowFYuZ2sy05CA1BFBKnvQ9zipoTrj1yATG4dCM8nUd9KrlyrBjrQxuQntD+
mcyg6ZLqowU0B5aZPYz/mZZSqEXNxOSKCYO2LRO6fNCMNPiQ7RRfvNbFRFmwKpp6
dkRpwF8S1N0jAIrgS5QHB1enH7i5vE2FDBJrrG1RUJRroMAaSyWVv081zvL/XK9I
/7GeC5wwIHtlgBQbFun2H7Ta9lqY5cjW9sJOdqfRAWB+vVJs8A68MiPqCmbcpb9h
6UJPQGQmm0/tGovcTPw9+T/YKw0kcCTfAprT9mCiKfFDv/dqr2EEWxDOWTIgwoqR
0loVdZXiqVcEWvyzW8c33vuV89F1nwenflyJGmoawYeO8Uiox5KCV42rR4W1E305
nBNEFL2U2WkQkEQlYD+4qdZFUvTDS/m93bxLZYNUMx3rTqxMGPR6eKTozvsLATbf
iWpiRvej++aXHMPF4mavR1eHPcfUFcBLMEfZjn6ijQJEAnYfoGImIe2M7KdhaHMT
o3RYFI3gSKCY6Ma95MjkYeIqUxVn0w1KnE2D+b+XY8IKsYwwyZVP4dl5cLIHGtic
taCx6YwpkZr6FBMfzZfnGNoka6Z+mOt2AZVNF2u58TqqCUIQ983Ea7ND9riHl1yx
XbmJo0F2NH+zRvpJVkKGwQBxC7di7rtuqHMD4cbOE5SCAXRZzLW1MpH4zsv9LBWF
S/4lqf21qS/UW9MpW5eQVTKEC7SQOK9xB0JrcV+/TPYaFrsmkBxx4Unr6F4h5MNv
A9mdy6Kcv/HFcJC/Zee9uAzKe8nyWWoM+5ItbeqFviVvcW0X8I5T3KYA5wBf2Rxb
Ky3jjCcB/H8NrVY9F9pEFxF0Akv6FXBFmanz0DGSzAXdr+dPe+wChxRb7ZNTLkkE
NnWa4MMs0Z6bf4ejLD6tDLO2Z60OXHOccFP48e6JPAG/D7w3uPVnRNv2I66gNDTd
oftri+ChW8Qv6yopWv/ZJ4MMMC5Se2WwdH5elJwlGOoy7DWnT+kAIUoPTsbtd7+s
x00Mp2j3w8nvIjGwvyR+pmH/AH/soFjhdh6RgmRFEAqQTLHaKyjaubTBf9mBKa4G
7y/va6tckmset1FUxZBTHG99zECFkfpX3UXFEFnF8nwZYxNiW4hrqAsUnkuT/V++
99bN465W4oRXeIU7iUkrD0FQZuR93rQESvsXwJIUR+2EM4rnro7LrO5s8uXNIE+9
9V6bHC4ezI3QzF7qGLTH2ZZ59wHuPbMuoW+D4EW1HRE72qdQM41p28b1V5l+RMB8
EwYtunetWsLy1Rh0r8cS6Tj4jO3fLxRhyj6HunREFXAXKI6sd9x06FXqPfmOhH43
iFyFLMJirUKmGmjx5znLY1xgh6dPVlVy4G35wwKiiyEknzXTfptyr/+xmtrTFSlv
50q/T6utOL+wPuBuxW0gw83yt+7UM+BPoK+w61W//0h4lyNlcZiPwhjb+3RVl5QT
MFenBfn+ueYzZvASBJ/iCOte7tLP2h+t8+b0dspkf8Q=
`protect END_PROTECTED
