`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHTaMDZy5ybBvPdsQnvmpohKO6fVI29lS6MjwATTltC4ArC/WgbIA6wq3A2OVykg
KnE50XYZ9QijN68rwkxPCBS21qeJw1wCLnl3ZT//pHIWte3gsPgkzJSqhwnRT5wq
eXk1BJuusgsx8EfkqYUvbYulAmGNXZCbqYGBs4M2ogso5g/UC6abKrsfXHSHp+ms
3zrHwP/z3mo50WiG1Lq4BO5Oq7Z0BwitjvaMtkaRnicjZ6usWG/7Kbnb/WcT4F3B
hIwfB5sXedSxp3jejPRlBHwWPgW2AR7NtJlA8HGceMbZIF6d6CXuy3NCmdWBv5AD
UWx9xzEDC40SiHbVEAacUsu31BblXGTyW3NgMLNdmuG6g/L67+hniFHk4MpDU3Rx
SvuSRbeXQn5VJUQd9wrk9l9+8BUx2yQW6O3d6Eh4sC5tTyJmokE4Ju1HtZMBvJc9
`protect END_PROTECTED
