`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7xffaLhyNuSSr0qsgOtIbICW44Xyg8K2Zcw659bJD5vvZBFhEpX032/ykrFt1Kk
C7K8y2P6N3H1BVDdhqjwuU2Df+W19I8n3mYXQ3QOwZ0D6Nhov8JmiIC56ctqDD+X
oTAkce+RcU++vJZ2BRUklCx0tGLG6JfY0DWdVoT/Sx5RxB4gAQS2ruJqkAgV5Yr6
QYoWX2oPRInfQ9KUWXghA6u7hWR1SNEVLNofb8BjyfT++2ZmGGNfYDzF8p5pE9kS
lKABQObWW4XhMhx0fAxFZV0moRLrtG/zd2gxuk/3uCVL+abEWATAzxJCbJZ9gnI6
xrIkwGZFG8GN1vH0M3rfgpyChIIW0RtFVFBCK3eYYhJJjBR2W0bMSOESpc+O99SN
N5F7ioW9pAkJJr4I34/GQmxjTBGbWEU4k5HKNAFdZ0OgMy94o/Tt1GgF25Xjr0kM
GKFLtWFQDunXIBf7uMtw8kpTx78BXANwH13mbaUEawEEzhZC7q4gVCR/5WN/lL9k
FvcvuozjzYeweJH3ITGRwSl7iyn9Z+l/LNNPgpMoSIoKynEoYkdCmReh5IuiamY3
RnXLV0SVUYkMePqWSAxldzJGL2l809eOjwmdPZIvOID5hMWP4B5LnWBndGov4oC+
uySAPBD+HdehbzZ9q6ZheqavAWAZRh1sVEhlpJOX/RaGOaUY9PQPQjCE7Swl2aoV
mIPS4c834W9uqVnDawIOUOXdFbbhrxalpKDNgSIoELrlTVxXufgGHWtYu2Gv7LEf
kpVi3kuD9r424XNTiSOKZwtkPNIppJxEV5O60Uz2mcdp9Xz/c6hQB3Mtd0gccp9y
iGFrKx9a8hICe4+VGRPhmQnb3kTWDCBJAN1AgWbk5JRMhD77PFrJVnchf3R4bPsT
kL3MTTtvrZganpZULw0nVpN61owVGRBCQnPQDYD6wlp1XZbdQWF/EUAtdGDSR8vR
cU648E+wRNRpBedUQK6vhkNsufxdICpZxQ14r2jBWmnQKbuZTlOAv4QuZMKli2yQ
KMW5JdKeUTChU4sl7LT/kGC+3837HXBFZYZ8+Ad4+xK1Jh7diNiLLwhqWe08i23u
VWPVWsxSxuQDj3NkOZGNLmZyZ3wsV6kCK7FJvJZD9qBBtyY7wEE8CCI2omRGN7Bz
eWbVxXO8jUH8ExWLS3QUv8XjFRqp7bK7W1iOEXguoUyrQY3YFfmm2uj/+BFcqS5x
LwYLFtL4++eGinmSqn90gfdNRvbhteB7xiRNe8kjO+0BWwOinO5YjH1lKxvchQdE
gX54i/3T0Y5NaHDj8pUwuYfjnX+XH5Yo7PX0AtAoMeoVw3VXAa0+687tfkLQHEP3
OEOH1OsAlHPkix51Or6BL0ARHe2WeWnfkWN7sg+qzmrFiGxQr8xt0iSRs2YDvUEe
mdn1MRo4rclSte98phhTStDFMT2EdHyLV1JkxTxntf+Z3d/XV9rFVoy2BsTrb7md
rCrg3HJorSLdhs7WkL0+2afdyRbk8FC6x07Rc2Fxc5Cpb+Awj8rbhIXWaSdfdGN1
SWQM0SFTwa9/0rbtQ4pub8ZgYrhD6fXmlWt65qrUtmRbwKgIsdJAKAAxNp7ACtcq
jBifkTW3zUu+GNH5ohOxGe6/8uQZdqLvj2HqT87ayPidEg/vxSV3+LMKHXgOxsxG
d0W6m3MYhTI8Md/fKNsN0w2MOXLlydHWQpWP1yPJSTsWBUo+PJb0TVtki6OtWgxy
iPnZRmlZyhQ5fdLL2bhMkvSqvSble6o0dR5TWxI3zxVgrZ2gXd6Xs+2YtvrUE78b
fjmAKyZ+QoNYhA6eOyhwz2fzc1P8dviJjSVKYxDM1ifBLXfMHBzGZevtmGWC86j8
F37fca22my5kH5pxbnKHw/NwGnUEvm3XkoE1QBWpC85ET252DEVJ9DbFbgL8qP/z
+New/eV3ku15hGQbOtFBMpZb4NXutzMRFaSTxOgCB9m6LXRl26MTGH7SGvHPu3nV
OnSkW3kPm0dDux0Rw3lt84QHi4GEKvIc6OUnV3Kc+OyHs9qLCHmJ8Xbal/YPu8S4
Y1U4XTqmymU/+LreoJU81v64blrc9xMdYkqRuCczGPF8Dl4yOo3hqXucwfqOUsW3
F1tJTpq0b523TRassnVQ4Ie0vETu77xnErmq6Aw1/looVybTfoqs1aS2o4iQLy8+
uBhusJCPMP83i1SbGQ/JYFJWG4SnNPNceHX2o462OKzuDVtWk+Iai+VebugsRC6E
vi3WHKkT839uY3JBCfBhcb3/GW2xx0YjePegyKm3to6YAjIUq0rXVJA3rEQ1SCsH
HKAJJVL4aBb6h01p1NoGDvb17YUuBZKOtNQlyty9VsxNENujXxmM8khyDBFth6+5
aZke/rp5OSoOlz2497m3hTfeS4wcb8gPr6X0aGLVVps8Z0yP5V5yB6YpZHmeSKaI
4cWs2RTfjr+aw3mc1mG+Bkhzy+L2ydxHOlT71/IEmDdS7h1wLin5tpWYIjN/zhM1
oXsXAQg/3HQ1LkEfUwdJVrPfsy2dFvogqz4ocZH+9J60rjCIDukMKcwU5QkdbvIa
v9cT7TUxxjDpUY+IbbJw1B7Vstfg3ZpP/qS9ExLqvmxpnqJKuqMzH1eCAQvZYgv9
AlUmEs63QTCLLf7pxTspeD0ByYdUom7TC34kln8mNHc8ODvrX1c+RknK3baNxeyU
NRUoGX8CckqmHt6I5Y3Z7vuwj+lzPwKs4L7JrXs39NUqSBzCOozCXpas1YUoO0uu
GX17DSuLexMCYdz0aQjp7f8GlFWKbHuWXV4WnBhMoDFzks2DM2ihME98E+GxGRHD
LOBKf1/YqMsdICEWjfLLi+/Yqpjwx15/mcbtMVdBJiifZ/jcOEHP1n5hZ4VXcfaX
WbZ1fFwQhlTs186XNeyGX5a8Ku05k6z765Ocdlz9H1aT9PqbeE1md0uOVr1HMkr9
K77t02OxAf2OD3BgB8XlXblW6KQ4RE/7v5P/70hLxJrHNX6sq+eZ6Dudap+W5SY9
V3J3nVr49P2wQ/OGls6w9+uoOqRR1OBORXWwiTqvm/wvx4llHpe2enppQwatQ755
tnG74F+yb5ri6QMZRKziBEH163vXyZcYt9GCvH7/pPZqQziH2l8y4qn8d0T9gJTK
q1g3/9YLyITJk1HZsEuzEsqE1/opD4kICFkIYFy2Dy98U4vWOhkvIOClLNXjn20X
RtlCoz4KzyDl2GlPQnJ56HTb8482vcbnY6X2Q2Iu86zJOJ0SBbhgHffXTs/ZTvTt
MvK8qRHcRTKVvRlr5f7SFHEYar6O22JIfQJR1jc9iuiyIbP1aXktxbKOns/0kdY6
SrSx3jxmSQK+UX22K9uIzdj4f5K7cxAARvoCNtv/SF9owF+M57KPTNUtrbIoNr2e
r3lPlFn9EZk+YwIhSsxbaoVi4Zcud060JhHj02HuU6bwvy/rmkQXOQM+gFJf+Crl
y8dDLHEJiHB3Ssv8fmH4E5fVcrq2vb0jhrt/AhbJpSJFHUheWU1K7StdkPnlKzx2
i/13xLTDZYnw7kbEkOGKJyTn8my8iiUnbmYodpx/F8r5MjKXvFqIkjS7g9lqfXHx
NhJIg7lwrgpPKOkEX8/CavhJ23n1Cxz9N4qQH1qTCLKH1MC0KSjkgKTRRyHGiR/N
j5nBlv/hhZkGO6G9yZenQoCfA+yTvFzDUhAOzvwiNQVKkWYbRbq0r7ZvHVzJTpaE
/2dLlyKPw6d77oAFCWAKGhTOOdBW86o69Nr8RAtCRd4JR6reyDwsxHfC45jAseon
RY8GJybS37sd5FicWk0cZy3s95JQ920OP95rRiki/UrfqYH2M5qACYMs9fvcgLXS
2d6g7WGk5FxcP+fTLmNeldHWoNvOINLgz4hi5luAGmj4DTZ7zwD14hthXxPbDVml
mTx5ZpO7t5IsvZCjLdcf6wA3a3cv0xmUnU5pp0wSihOqjhor28z1dZZ94wvl8qlE
BEFIF3X9mWj4LfUOW0LMkLYWNljbQRUsCSkGVkqFBKlGSIsphMuydkIpxqcSSSbV
PDn+l1c9nCI1mxFW4QWtnh0ALVZYO1I1NJF+RiIhuQJohGakxol/kTMDh6mH/o1h
rEEWFR5KEi2pHZpy2Px7wbaHbOogiB4XSgYVPpPqjuDk+YQGI30N82m+IhMtXy/l
PO0zGIxI2JaeRm156eGF6Z4i8jgJY3CfRonTOjEa9N90GVlor/9KCSRdk38mfXgW
Z3DoteiKHz6mfDDTL1Gd5ohXrvNGizSDWGBS+C6pvhPN7074uBLejGOpp+BwHbyY
6oglHIqp+tBW4blL9cjsgKkyA6uZ2tp1vmGHizD3P/JpEwKyoVec56pqqUtzexQk
w4yq2yG7qLeId30OnyOkzZeveLiloNyL/1uGZNy9mVHwHmog7kobkAKBCZLItMZE
xg41GtEEgYtRrQXZnT2803WdfCF9Ykd2Fr4f8pLUt+VJ/n4yVzmPFmkBm/Ws4XFZ
WNk1abhk1uoFXnEFRqhDiF4CnqXkUJj0Mtvg133gM5xf4M4lI1Ji7QJVIWyWg54P
9j368t+E3uicNvz2XlJLHoFb20vz3D7i/FFAbcgwzTCZyF+b4KB/zbXmac+mu/D1
XK9XJK5BiAszqAvp/pJo/e6en7bbmdUy3gWavz+LFC4o5G93NUbza/C+gpJXn1ge
3skSlOJ6DPNo9HYeS7pg9RrKk3uEaBoavlOpqTATBgl9iFLeEGMJC+qbi+9ZqwNO
GNz88N5z/dGTD/CPfVBfn09tn2kGMNEe/fgs43jamuwBD5SuTLe9LdpPA8xYzSwO
rzQww8dcgSARzvcMdKnfSI/o5e993uwP+GOhH/2WoabZIm3EK4frOQKAlDNlBdRL
SEYFnNxqR+dQw8Bs+kUM2XYknckEPigTDrsMGRs4Rs7FfFuRV412BiwhFNQYjWRH
NcC30glC+ItTzAdlW3QrgU6Y8kUJQQ7EwhF/D557TvmqqcpK8HGJVFXkv7httThm
b4cnWX6wEZcBvJu5/rEtBiGtuPfJZ1z45Hpdd8xo61SnaoAon/BwOftzfFiHGnJ/
nbd744H0vgpU3WSutybls5EkEFZe0fAh7Mn+wusG34l0QdnUlrHnXu22cVb1oJ8t
/sIa7Ur2tsNs/GNzCoG8lGrzgxY9sNTucG6dvhs6djAAMKoNDr4yzBX1tSdu0/fR
Wp6wVvN/1cGreGufee1gImJKggmw3VAqCNZ7g++BbEeJc5fOVxGunHH6mXwym8uI
EDL6CTKGnbOI7Sy1FzDI2MyK6a8FuXdBxqkwNsE84i1q6OZOlrRTaxAuTsjmZnG6
ysKi4IQNt/fOZLUCXNc/FG4Yo4H5ZzakELEVqINumvCeovuU2TX2kFs/fWDuknNu
IR7JN++Z47y5dBEsDnzs6WaH2mglv337BL8Fv/ukwnYJgxSWDnu5aqff57zOXXLE
p0N+VOPRcIVymCqepiCeFVlo468UYD01GnJV80dg0KzyxfN0iKmuYFl4GJKas+nz
zDHjkj0CmyDuO7lNXq6V2/tw/iteDr7BTDqhAkCw6ghpZTzWAxwGRAw4xEpQwMyl
IZHkEMWjOixM655g3w0yDh7VutNv+XqXatBGY49Ink6YA602uuYNhakq0SpKE2OR
LPFCf4P3F5sfPuezSkAp9H0saxF3W8MdUW5yK8Z24N6Dpb5cwKtqwBheogFnlZvZ
RmfGoTA7nmdkef+5v/Um2C0/9qoO9WRh5ynLDQyTf171CFaaKvamHfgT2M6mkYwo
YOZWUplQN/Hp8gkjU3etqPIbI4XLWbH/6BkzBcnIFoU=
`protect END_PROTECTED
